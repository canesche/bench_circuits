// Benchmark "testing" written by ABC on Thu Oct  8 22:16:30 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A76  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A76;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ , \new_[350]_ ,
    \new_[351]_ , \new_[352]_ , \new_[353]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[405]_ ,
    \new_[406]_ , \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ ,
    \new_[411]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[436]_ , \new_[437]_ , \new_[438]_ , \new_[439]_ , \new_[440]_ ,
    \new_[441]_ , \new_[442]_ , \new_[443]_ , \new_[444]_ , \new_[445]_ ,
    \new_[446]_ , \new_[447]_ , \new_[448]_ , \new_[449]_ , \new_[450]_ ,
    \new_[451]_ , \new_[452]_ , \new_[453]_ , \new_[454]_ , \new_[455]_ ,
    \new_[456]_ , \new_[457]_ , \new_[458]_ , \new_[459]_ , \new_[460]_ ,
    \new_[461]_ , \new_[462]_ , \new_[463]_ , \new_[464]_ , \new_[465]_ ,
    \new_[466]_ , \new_[467]_ , \new_[468]_ , \new_[469]_ , \new_[470]_ ,
    \new_[471]_ , \new_[472]_ , \new_[473]_ , \new_[474]_ , \new_[475]_ ,
    \new_[476]_ , \new_[477]_ , \new_[478]_ , \new_[479]_ , \new_[480]_ ,
    \new_[481]_ , \new_[482]_ , \new_[483]_ , \new_[484]_ , \new_[485]_ ,
    \new_[486]_ , \new_[487]_ , \new_[488]_ , \new_[489]_ , \new_[490]_ ,
    \new_[491]_ , \new_[492]_ , \new_[493]_ , \new_[494]_ , \new_[495]_ ,
    \new_[496]_ , \new_[497]_ , \new_[498]_ , \new_[499]_ , \new_[500]_ ,
    \new_[501]_ , \new_[502]_ , \new_[503]_ , \new_[504]_ , \new_[505]_ ,
    \new_[506]_ , \new_[507]_ , \new_[508]_ , \new_[509]_ , \new_[510]_ ,
    \new_[511]_ , \new_[512]_ , \new_[513]_ , \new_[514]_ , \new_[515]_ ,
    \new_[516]_ , \new_[517]_ , \new_[518]_ , \new_[519]_ , \new_[520]_ ,
    \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[525]_ ,
    \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ , \new_[530]_ ,
    \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ , \new_[535]_ ,
    \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ , \new_[540]_ ,
    \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ , \new_[545]_ ,
    \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ , \new_[550]_ ,
    \new_[551]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[566]_ , \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ ,
    \new_[571]_ , \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ ,
    \new_[576]_ , \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ ,
    \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[584]_ , \new_[585]_ ,
    \new_[586]_ , \new_[587]_ , \new_[588]_ , \new_[589]_ , \new_[590]_ ,
    \new_[591]_ , \new_[592]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[598]_ , \new_[599]_ , \new_[600]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ ,
    \new_[611]_ , \new_[612]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[616]_ , \new_[617]_ , \new_[618]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[626]_ , \new_[627]_ , \new_[628]_ , \new_[629]_ , \new_[630]_ ,
    \new_[631]_ , \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ ,
    \new_[636]_ , \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ ,
    \new_[641]_ , \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ ,
    \new_[646]_ , \new_[647]_ , \new_[648]_ , \new_[649]_ , \new_[650]_ ,
    \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[655]_ ,
    \new_[656]_ , \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ ,
    \new_[661]_ , \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ ,
    \new_[666]_ , \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ ,
    \new_[671]_ , \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ ,
    \new_[676]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ ,
    \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ ,
    \new_[686]_ , \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ ,
    \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ ,
    \new_[696]_ , \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ ,
    \new_[701]_ , \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ ,
    \new_[706]_ , \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ ,
    \new_[711]_ , \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ ,
    \new_[716]_ , \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ ,
    \new_[726]_ , \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ ,
    \new_[731]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[736]_ , \new_[737]_ , \new_[738]_ , \new_[739]_ , \new_[740]_ ,
    \new_[741]_ , \new_[742]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ ,
    \new_[746]_ , \new_[747]_ , \new_[748]_ , \new_[749]_ , \new_[750]_ ,
    \new_[751]_ , \new_[752]_ , \new_[753]_ , \new_[754]_ , \new_[755]_ ,
    \new_[756]_ , \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ ,
    \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ ,
    \new_[766]_ , \new_[767]_ , \new_[768]_ , \new_[769]_ , \new_[770]_ ,
    \new_[771]_ , \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ ,
    \new_[776]_ , \new_[777]_ , \new_[778]_ , \new_[779]_ , \new_[780]_ ,
    \new_[781]_ , \new_[782]_ , \new_[783]_ , \new_[784]_ , \new_[785]_ ,
    \new_[786]_ , \new_[787]_ , \new_[788]_ , \new_[789]_ , \new_[790]_ ,
    \new_[791]_ , \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ ,
    \new_[796]_ , \new_[797]_ , \new_[798]_ , \new_[799]_ , \new_[800]_ ,
    \new_[801]_ , \new_[802]_ , \new_[803]_ , \new_[804]_ , \new_[805]_ ,
    \new_[806]_ , \new_[807]_ , \new_[808]_ , \new_[809]_ , \new_[810]_ ,
    \new_[811]_ , \new_[812]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ ,
    \new_[816]_ , \new_[817]_ , \new_[818]_ , \new_[819]_ , \new_[820]_ ,
    \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[824]_ , \new_[825]_ ,
    \new_[826]_ , \new_[827]_ , \new_[828]_ , \new_[829]_ , \new_[830]_ ,
    \new_[831]_ , \new_[832]_ , \new_[833]_ , \new_[834]_ , \new_[835]_ ,
    \new_[836]_ , \new_[837]_ , \new_[838]_ , \new_[839]_ , \new_[840]_ ,
    \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[845]_ ,
    \new_[846]_ , \new_[847]_ , \new_[848]_ , \new_[849]_ , \new_[850]_ ,
    \new_[851]_ , \new_[852]_ , \new_[853]_ , \new_[854]_ , \new_[855]_ ,
    \new_[856]_ , \new_[857]_ , \new_[858]_ , \new_[859]_ , \new_[860]_ ,
    \new_[861]_ , \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[865]_ ,
    \new_[866]_ , \new_[867]_ , \new_[868]_ , \new_[869]_ , \new_[870]_ ,
    \new_[871]_ , \new_[872]_ , \new_[873]_ , \new_[874]_ , \new_[875]_ ,
    \new_[876]_ , \new_[877]_ , \new_[878]_ , \new_[879]_ , \new_[880]_ ,
    \new_[881]_ , \new_[882]_ , \new_[883]_ , \new_[884]_ , \new_[885]_ ,
    \new_[886]_ , \new_[887]_ , \new_[888]_ , \new_[889]_ , \new_[890]_ ,
    \new_[891]_ , \new_[892]_ , \new_[893]_ , \new_[894]_ , \new_[895]_ ,
    \new_[896]_ , \new_[897]_ , \new_[898]_ , \new_[899]_ , \new_[900]_ ,
    \new_[901]_ , \new_[902]_ , \new_[903]_ , \new_[904]_ , \new_[905]_ ,
    \new_[906]_ , \new_[907]_ , \new_[908]_ , \new_[909]_ , \new_[910]_ ,
    \new_[911]_ , \new_[912]_ , \new_[913]_ , \new_[914]_ , \new_[915]_ ,
    \new_[916]_ , \new_[917]_ , \new_[918]_ , \new_[919]_ , \new_[920]_ ,
    \new_[921]_ , \new_[922]_ , \new_[923]_ , \new_[924]_ , \new_[925]_ ,
    \new_[926]_ , \new_[927]_ , \new_[928]_ , \new_[929]_ , \new_[930]_ ,
    \new_[931]_ , \new_[932]_ , \new_[933]_ , \new_[934]_ , \new_[935]_ ,
    \new_[936]_ , \new_[937]_ , \new_[938]_ , \new_[939]_ , \new_[940]_ ,
    \new_[941]_ , \new_[942]_ , \new_[943]_ , \new_[944]_ , \new_[945]_ ,
    \new_[946]_ , \new_[947]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ ,
    \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[955]_ ,
    \new_[956]_ , \new_[957]_ , \new_[958]_ , \new_[959]_ , \new_[960]_ ,
    \new_[961]_ , \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ ,
    \new_[966]_ , \new_[967]_ , \new_[968]_ , \new_[969]_ , \new_[970]_ ,
    \new_[971]_ , \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[975]_ ,
    \new_[976]_ , \new_[977]_ , \new_[978]_ , \new_[979]_ , \new_[980]_ ,
    \new_[981]_ , \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ ,
    \new_[986]_ , \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ ,
    \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ ,
    \new_[996]_ , \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ ,
    \new_[1001]_ , \new_[1002]_ , \new_[1003]_ , \new_[1004]_ ,
    \new_[1005]_ , \new_[1006]_ , \new_[1007]_ , \new_[1008]_ ,
    \new_[1009]_ , \new_[1010]_ , \new_[1011]_ , \new_[1012]_ ,
    \new_[1013]_ , \new_[1014]_ , \new_[1015]_ , \new_[1016]_ ,
    \new_[1017]_ , \new_[1018]_ , \new_[1019]_ , \new_[1020]_ ,
    \new_[1021]_ , \new_[1022]_ , \new_[1023]_ , \new_[1024]_ ,
    \new_[1025]_ , \new_[1026]_ , \new_[1027]_ , \new_[1028]_ ,
    \new_[1029]_ , \new_[1030]_ , \new_[1031]_ , \new_[1032]_ ,
    \new_[1033]_ , \new_[1034]_ , \new_[1035]_ , \new_[1036]_ ,
    \new_[1037]_ , \new_[1038]_ , \new_[1039]_ , \new_[1040]_ ,
    \new_[1041]_ , \new_[1042]_ , \new_[1043]_ , \new_[1044]_ ,
    \new_[1045]_ , \new_[1046]_ , \new_[1047]_ , \new_[1048]_ ,
    \new_[1049]_ , \new_[1050]_ , \new_[1051]_ , \new_[1052]_ ,
    \new_[1053]_ , \new_[1054]_ , \new_[1055]_ , \new_[1056]_ ,
    \new_[1057]_ , \new_[1058]_ , \new_[1059]_ , \new_[1060]_ ,
    \new_[1061]_ , \new_[1062]_ , \new_[1063]_ , \new_[1064]_ ,
    \new_[1065]_ , \new_[1066]_ , \new_[1067]_ , \new_[1068]_ ,
    \new_[1069]_ , \new_[1070]_ , \new_[1071]_ , \new_[1072]_ ,
    \new_[1073]_ , \new_[1074]_ , \new_[1075]_ , \new_[1076]_ ,
    \new_[1077]_ , \new_[1078]_ , \new_[1079]_ , \new_[1080]_ ,
    \new_[1081]_ , \new_[1082]_ , \new_[1083]_ , \new_[1084]_ ,
    \new_[1085]_ , \new_[1086]_ , \new_[1087]_ , \new_[1088]_ ,
    \new_[1089]_ , \new_[1090]_ , \new_[1091]_ , \new_[1092]_ ,
    \new_[1093]_ , \new_[1094]_ , \new_[1095]_ , \new_[1096]_ ,
    \new_[1097]_ , \new_[1098]_ , \new_[1099]_ , \new_[1100]_ ,
    \new_[1101]_ , \new_[1102]_ , \new_[1103]_ , \new_[1104]_ ,
    \new_[1105]_ , \new_[1106]_ , \new_[1107]_ , \new_[1108]_ ,
    \new_[1109]_ , \new_[1110]_ , \new_[1111]_ , \new_[1112]_ ,
    \new_[1113]_ , \new_[1114]_ , \new_[1115]_ , \new_[1116]_ ,
    \new_[1117]_ , \new_[1118]_ , \new_[1119]_ , \new_[1120]_ ,
    \new_[1121]_ , \new_[1122]_ , \new_[1123]_ , \new_[1124]_ ,
    \new_[1125]_ , \new_[1126]_ , \new_[1127]_ , \new_[1128]_ ,
    \new_[1129]_ , \new_[1130]_ , \new_[1131]_ , \new_[1132]_ ,
    \new_[1133]_ , \new_[1134]_ , \new_[1135]_ , \new_[1136]_ ,
    \new_[1137]_ , \new_[1138]_ , \new_[1139]_ , \new_[1140]_ ,
    \new_[1141]_ , \new_[1142]_ , \new_[1143]_ , \new_[1144]_ ,
    \new_[1145]_ , \new_[1146]_ , \new_[1147]_ , \new_[1148]_ ,
    \new_[1149]_ , \new_[1150]_ , \new_[1151]_ , \new_[1152]_ ,
    \new_[1153]_ , \new_[1154]_ , \new_[1155]_ , \new_[1156]_ ,
    \new_[1157]_ , \new_[1158]_ , \new_[1159]_ , \new_[1160]_ ,
    \new_[1161]_ , \new_[1162]_ , \new_[1163]_ , \new_[1164]_ ,
    \new_[1165]_ , \new_[1166]_ , \new_[1167]_ , \new_[1168]_ ,
    \new_[1169]_ , \new_[1170]_ , \new_[1171]_ , \new_[1172]_ ,
    \new_[1173]_ , \new_[1174]_ , \new_[1175]_ , \new_[1176]_ ,
    \new_[1177]_ , \new_[1178]_ , \new_[1179]_ , \new_[1180]_ ,
    \new_[1181]_ , \new_[1182]_ , \new_[1183]_ , \new_[1184]_ ,
    \new_[1185]_ , \new_[1186]_ , \new_[1187]_ , \new_[1188]_ ,
    \new_[1189]_ , \new_[1190]_ , \new_[1191]_ , \new_[1192]_ ,
    \new_[1193]_ , \new_[1194]_ , \new_[1195]_ , \new_[1196]_ ,
    \new_[1197]_ , \new_[1198]_ , \new_[1199]_ , \new_[1200]_ ,
    \new_[1201]_ , \new_[1202]_ , \new_[1203]_ , \new_[1204]_ ,
    \new_[1205]_ , \new_[1206]_ , \new_[1207]_ , \new_[1208]_ ,
    \new_[1209]_ , \new_[1210]_ , \new_[1211]_ , \new_[1212]_ ,
    \new_[1213]_ , \new_[1214]_ , \new_[1215]_ , \new_[1216]_ ,
    \new_[1217]_ , \new_[1218]_ , \new_[1219]_ , \new_[1220]_ ,
    \new_[1221]_ , \new_[1222]_ , \new_[1223]_ , \new_[1224]_ ,
    \new_[1225]_ , \new_[1226]_ , \new_[1227]_ , \new_[1228]_ ,
    \new_[1229]_ , \new_[1230]_ , \new_[1231]_ , \new_[1232]_ ,
    \new_[1233]_ , \new_[1234]_ , \new_[1235]_ , \new_[1236]_ ,
    \new_[1237]_ , \new_[1238]_ , \new_[1239]_ , \new_[1240]_ ,
    \new_[1241]_ , \new_[1242]_ , \new_[1243]_ , \new_[1244]_ ,
    \new_[1245]_ , \new_[1246]_ , \new_[1247]_ , \new_[1248]_ ,
    \new_[1249]_ , \new_[1250]_ , \new_[1251]_ , \new_[1252]_ ,
    \new_[1253]_ , \new_[1254]_ , \new_[1255]_ , \new_[1256]_ ,
    \new_[1257]_ , \new_[1258]_ , \new_[1259]_ , \new_[1260]_ ,
    \new_[1261]_ , \new_[1262]_ , \new_[1263]_ , \new_[1264]_ ,
    \new_[1265]_ , \new_[1266]_ , \new_[1267]_ , \new_[1268]_ ,
    \new_[1269]_ , \new_[1270]_ , \new_[1271]_ , \new_[1272]_ ,
    \new_[1273]_ , \new_[1274]_ , \new_[1275]_ , \new_[1276]_ ,
    \new_[1277]_ , \new_[1278]_ , \new_[1279]_ , \new_[1280]_ ,
    \new_[1281]_ , \new_[1282]_ , \new_[1283]_ , \new_[1284]_ ,
    \new_[1285]_ , \new_[1286]_ , \new_[1287]_ , \new_[1288]_ ,
    \new_[1289]_ , \new_[1290]_ , \new_[1291]_ , \new_[1292]_ ,
    \new_[1293]_ , \new_[1294]_ , \new_[1295]_ , \new_[1296]_ ,
    \new_[1297]_ , \new_[1298]_ , \new_[1299]_ , \new_[1300]_ ,
    \new_[1301]_ , \new_[1302]_ , \new_[1303]_ , \new_[1304]_ ,
    \new_[1305]_ , \new_[1306]_ , \new_[1307]_ , \new_[1308]_ ,
    \new_[1309]_ , \new_[1310]_ , \new_[1311]_ , \new_[1312]_ ,
    \new_[1313]_ , \new_[1314]_ , \new_[1315]_ , \new_[1316]_ ,
    \new_[1317]_ , \new_[1318]_ , \new_[1319]_ , \new_[1320]_ ,
    \new_[1321]_ , \new_[1322]_ , \new_[1323]_ , \new_[1324]_ ,
    \new_[1325]_ , \new_[1326]_ , \new_[1327]_ , \new_[1328]_ ,
    \new_[1329]_ , \new_[1330]_ , \new_[1331]_ , \new_[1332]_ ,
    \new_[1333]_ , \new_[1334]_ , \new_[1335]_ , \new_[1336]_ ,
    \new_[1337]_ , \new_[1338]_ , \new_[1339]_ , \new_[1340]_ ,
    \new_[1341]_ , \new_[1342]_ , \new_[1343]_ , \new_[1344]_ ,
    \new_[1345]_ , \new_[1346]_ , \new_[1347]_ , \new_[1348]_ ,
    \new_[1349]_ , \new_[1350]_ , \new_[1351]_ , \new_[1352]_ ,
    \new_[1353]_ , \new_[1354]_ , \new_[1355]_ , \new_[1356]_ ,
    \new_[1357]_ , \new_[1358]_ , \new_[1359]_ , \new_[1360]_ ,
    \new_[1361]_ , \new_[1362]_ , \new_[1363]_ , \new_[1364]_ ,
    \new_[1365]_ , \new_[1366]_ , \new_[1367]_ , \new_[1368]_ ,
    \new_[1369]_ , \new_[1370]_ , \new_[1371]_ , \new_[1372]_ ,
    \new_[1373]_ , \new_[1374]_ , \new_[1375]_ , \new_[1376]_ ,
    \new_[1377]_ , \new_[1378]_ , \new_[1379]_ , \new_[1380]_ ,
    \new_[1381]_ , \new_[1382]_ , \new_[1383]_ , \new_[1384]_ ,
    \new_[1385]_ , \new_[1386]_ , \new_[1387]_ , \new_[1388]_ ,
    \new_[1389]_ , \new_[1390]_ , \new_[1391]_ , \new_[1392]_ ,
    \new_[1393]_ , \new_[1394]_ , \new_[1395]_ , \new_[1396]_ ,
    \new_[1397]_ , \new_[1398]_ , \new_[1399]_ , \new_[1400]_ ,
    \new_[1401]_ , \new_[1402]_ , \new_[1403]_ , \new_[1404]_ ,
    \new_[1405]_ , \new_[1406]_ , \new_[1407]_ , \new_[1408]_ ,
    \new_[1409]_ , \new_[1410]_ , \new_[1411]_ , \new_[1412]_ ,
    \new_[1413]_ , \new_[1414]_ , \new_[1415]_ , \new_[1416]_ ,
    \new_[1417]_ , \new_[1418]_ , \new_[1419]_ , \new_[1420]_ ,
    \new_[1421]_ , \new_[1422]_ , \new_[1423]_ , \new_[1424]_ ,
    \new_[1425]_ , \new_[1426]_ , \new_[1427]_ , \new_[1428]_ ,
    \new_[1429]_ , \new_[1430]_ , \new_[1431]_ , \new_[1432]_ ,
    \new_[1433]_ , \new_[1434]_ , \new_[1435]_ , \new_[1436]_ ,
    \new_[1437]_ , \new_[1438]_ , \new_[1439]_ , \new_[1440]_ ,
    \new_[1441]_ , \new_[1442]_ , \new_[1443]_ , \new_[1444]_ ,
    \new_[1445]_ , \new_[1446]_ , \new_[1447]_ , \new_[1448]_ ,
    \new_[1449]_ , \new_[1450]_ , \new_[1451]_ , \new_[1452]_ ,
    \new_[1453]_ , \new_[1454]_ , \new_[1455]_ , \new_[1456]_ ,
    \new_[1457]_ , \new_[1458]_ , \new_[1459]_ , \new_[1460]_ ,
    \new_[1461]_ , \new_[1462]_ , \new_[1463]_ , \new_[1464]_ ,
    \new_[1465]_ , \new_[1466]_ , \new_[1467]_ , \new_[1468]_ ,
    \new_[1469]_ , \new_[1470]_ , \new_[1471]_ , \new_[1472]_ ,
    \new_[1473]_ , \new_[1474]_ , \new_[1475]_ , \new_[1476]_ ,
    \new_[1477]_ , \new_[1478]_ , \new_[1479]_ , \new_[1480]_ ,
    \new_[1481]_ , \new_[1482]_ , \new_[1483]_ , \new_[1484]_ ,
    \new_[1485]_ , \new_[1486]_ , \new_[1487]_ , \new_[1488]_ ,
    \new_[1489]_ , \new_[1490]_ , \new_[1491]_ , \new_[1492]_ ,
    \new_[1493]_ , \new_[1494]_ , \new_[1495]_ , \new_[1496]_ ,
    \new_[1497]_ , \new_[1498]_ , \new_[1499]_ , \new_[1500]_ ,
    \new_[1501]_ , \new_[1502]_ , \new_[1503]_ , \new_[1504]_ ,
    \new_[1505]_ , \new_[1506]_ , \new_[1507]_ , \new_[1508]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1512]_ ,
    \new_[1513]_ , \new_[1514]_ , \new_[1515]_ , \new_[1516]_ ,
    \new_[1517]_ , \new_[1518]_ , \new_[1519]_ , \new_[1520]_ ,
    \new_[1521]_ , \new_[1522]_ , \new_[1523]_ , \new_[1524]_ ,
    \new_[1525]_ , \new_[1526]_ , \new_[1527]_ , \new_[1528]_ ,
    \new_[1529]_ , \new_[1530]_ , \new_[1531]_ , \new_[1532]_ ,
    \new_[1533]_ , \new_[1534]_ , \new_[1535]_ , \new_[1536]_ ,
    \new_[1537]_ , \new_[1538]_ , \new_[1539]_ , \new_[1540]_ ,
    \new_[1541]_ , \new_[1542]_ , \new_[1543]_ , \new_[1544]_ ,
    \new_[1545]_ , \new_[1546]_ , \new_[1547]_ , \new_[1548]_ ,
    \new_[1549]_ , \new_[1550]_ , \new_[1551]_ , \new_[1552]_ ,
    \new_[1553]_ , \new_[1554]_ , \new_[1555]_ , \new_[1556]_ ,
    \new_[1557]_ , \new_[1558]_ , \new_[1559]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1562]_ , \new_[1563]_ , \new_[1564]_ ,
    \new_[1565]_ , \new_[1566]_ , \new_[1567]_ , \new_[1568]_ ,
    \new_[1569]_ , \new_[1570]_ , \new_[1571]_ , \new_[1572]_ ,
    \new_[1573]_ , \new_[1574]_ , \new_[1575]_ , \new_[1576]_ ,
    \new_[1577]_ , \new_[1578]_ , \new_[1579]_ , \new_[1580]_ ,
    \new_[1581]_ , \new_[1582]_ , \new_[1583]_ , \new_[1584]_ ,
    \new_[1585]_ , \new_[1586]_ , \new_[1587]_ , \new_[1588]_ ,
    \new_[1589]_ , \new_[1590]_ , \new_[1591]_ , \new_[1592]_ ,
    \new_[1593]_ , \new_[1594]_ , \new_[1595]_ , \new_[1596]_ ,
    \new_[1597]_ , \new_[1598]_ , \new_[1599]_ , \new_[1600]_ ,
    \new_[1601]_ , \new_[1602]_ , \new_[1603]_ , \new_[1604]_ ,
    \new_[1605]_ , \new_[1606]_ , \new_[1607]_ , \new_[1608]_ ,
    \new_[1609]_ , \new_[1610]_ , \new_[1611]_ , \new_[1612]_ ,
    \new_[1613]_ , \new_[1614]_ , \new_[1615]_ , \new_[1616]_ ,
    \new_[1617]_ , \new_[1618]_ , \new_[1619]_ , \new_[1620]_ ,
    \new_[1621]_ , \new_[1622]_ , \new_[1623]_ , \new_[1624]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1627]_ , \new_[1628]_ ,
    \new_[1629]_ , \new_[1630]_ , \new_[1631]_ , \new_[1632]_ ,
    \new_[1633]_ , \new_[1634]_ , \new_[1635]_ , \new_[1636]_ ,
    \new_[1637]_ , \new_[1638]_ , \new_[1639]_ , \new_[1640]_ ,
    \new_[1641]_ , \new_[1642]_ , \new_[1643]_ , \new_[1644]_ ,
    \new_[1645]_ , \new_[1646]_ , \new_[1647]_ , \new_[1648]_ ,
    \new_[1649]_ , \new_[1650]_ , \new_[1651]_ , \new_[1652]_ ,
    \new_[1653]_ , \new_[1654]_ , \new_[1655]_ , \new_[1656]_ ,
    \new_[1657]_ , \new_[1658]_ , \new_[1659]_ , \new_[1660]_ ,
    \new_[1661]_ , \new_[1662]_ , \new_[1663]_ , \new_[1664]_ ,
    \new_[1665]_ , \new_[1666]_ , \new_[1667]_ , \new_[1668]_ ,
    \new_[1669]_ , \new_[1670]_ , \new_[1671]_ , \new_[1672]_ ,
    \new_[1673]_ , \new_[1674]_ , \new_[1675]_ , \new_[1676]_ ,
    \new_[1677]_ , \new_[1678]_ , \new_[1679]_ , \new_[1680]_ ,
    \new_[1681]_ , \new_[1682]_ , \new_[1683]_ , \new_[1684]_ ,
    \new_[1685]_ , \new_[1686]_ , \new_[1687]_ , \new_[1688]_ ,
    \new_[1689]_ , \new_[1690]_ , \new_[1691]_ , \new_[1692]_ ,
    \new_[1693]_ , \new_[1694]_ , \new_[1695]_ , \new_[1696]_ ,
    \new_[1697]_ , \new_[1698]_ , \new_[1699]_ , \new_[1700]_ ,
    \new_[1701]_ , \new_[1702]_ , \new_[1703]_ , \new_[1704]_ ,
    \new_[1705]_ , \new_[1706]_ , \new_[1707]_ , \new_[1708]_ ,
    \new_[1709]_ , \new_[1710]_ , \new_[1711]_ , \new_[1712]_ ,
    \new_[1713]_ , \new_[1714]_ , \new_[1715]_ , \new_[1716]_ ,
    \new_[1717]_ , \new_[1718]_ , \new_[1719]_ , \new_[1720]_ ,
    \new_[1721]_ , \new_[1722]_ , \new_[1723]_ , \new_[1724]_ ,
    \new_[1725]_ , \new_[1726]_ , \new_[1727]_ , \new_[1728]_ ,
    \new_[1729]_ , \new_[1730]_ , \new_[1731]_ , \new_[1732]_ ,
    \new_[1733]_ , \new_[1734]_ , \new_[1735]_ , \new_[1736]_ ,
    \new_[1737]_ , \new_[1738]_ , \new_[1739]_ , \new_[1740]_ ,
    \new_[1741]_ , \new_[1742]_ , \new_[1743]_ , \new_[1744]_ ,
    \new_[1745]_ , \new_[1746]_ , \new_[1747]_ , \new_[1748]_ ,
    \new_[1749]_ , \new_[1750]_ , \new_[1751]_ , \new_[1752]_ ,
    \new_[1753]_ , \new_[1754]_ , \new_[1755]_ , \new_[1756]_ ,
    \new_[1757]_ , \new_[1758]_ , \new_[1759]_ , \new_[1760]_ ,
    \new_[1761]_ , \new_[1762]_ , \new_[1763]_ , \new_[1764]_ ,
    \new_[1765]_ , \new_[1766]_ , \new_[1767]_ , \new_[1768]_ ,
    \new_[1769]_ , \new_[1770]_ , \new_[1771]_ , \new_[1772]_ ,
    \new_[1773]_ , \new_[1774]_ , \new_[1775]_ , \new_[1776]_ ,
    \new_[1777]_ , \new_[1778]_ , \new_[1779]_ , \new_[1780]_ ,
    \new_[1781]_ , \new_[1782]_ , \new_[1783]_ , \new_[1784]_ ,
    \new_[1785]_ , \new_[1786]_ , \new_[1787]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1791]_ , \new_[1792]_ ,
    \new_[1793]_ , \new_[1794]_ , \new_[1795]_ , \new_[1796]_ ,
    \new_[1797]_ , \new_[1798]_ , \new_[1799]_ , \new_[1800]_ ,
    \new_[1801]_ , \new_[1802]_ , \new_[1803]_ , \new_[1804]_ ,
    \new_[1805]_ , \new_[1806]_ , \new_[1807]_ , \new_[1808]_ ,
    \new_[1809]_ , \new_[1810]_ , \new_[1811]_ , \new_[1812]_ ,
    \new_[1813]_ , \new_[1814]_ , \new_[1815]_ , \new_[1816]_ ,
    \new_[1817]_ , \new_[1818]_ , \new_[1819]_ , \new_[1820]_ ,
    \new_[1821]_ , \new_[1822]_ , \new_[1823]_ , \new_[1824]_ ,
    \new_[1825]_ , \new_[1826]_ , \new_[1827]_ , \new_[1828]_ ,
    \new_[1829]_ , \new_[1830]_ , \new_[1831]_ , \new_[1832]_ ,
    \new_[1833]_ , \new_[1834]_ , \new_[1835]_ , \new_[1836]_ ,
    \new_[1837]_ , \new_[1838]_ , \new_[1839]_ , \new_[1840]_ ,
    \new_[1841]_ , \new_[1842]_ , \new_[1843]_ , \new_[1844]_ ,
    \new_[1845]_ , \new_[1846]_ , \new_[1847]_ , \new_[1848]_ ,
    \new_[1849]_ , \new_[1850]_ , \new_[1851]_ , \new_[1852]_ ,
    \new_[1853]_ , \new_[1854]_ , \new_[1855]_ , \new_[1856]_ ,
    \new_[1857]_ , \new_[1858]_ , \new_[1859]_ , \new_[1860]_ ,
    \new_[1861]_ , \new_[1862]_ , \new_[1863]_ , \new_[1864]_ ,
    \new_[1865]_ , \new_[1866]_ , \new_[1867]_ , \new_[1868]_ ,
    \new_[1869]_ , \new_[1870]_ , \new_[1871]_ , \new_[1872]_ ,
    \new_[1873]_ , \new_[1874]_ , \new_[1875]_ , \new_[1876]_ ,
    \new_[1877]_ , \new_[1878]_ , \new_[1879]_ , \new_[1880]_ ,
    \new_[1881]_ , \new_[1882]_ , \new_[1883]_ , \new_[1884]_ ,
    \new_[1885]_ , \new_[1886]_ , \new_[1887]_ , \new_[1888]_ ,
    \new_[1889]_ , \new_[1890]_ , \new_[1891]_ , \new_[1892]_ ,
    \new_[1893]_ , \new_[1894]_ , \new_[1895]_ , \new_[1896]_ ,
    \new_[1897]_ , \new_[1898]_ , \new_[1899]_ , \new_[1900]_ ,
    \new_[1901]_ , \new_[1902]_ , \new_[1903]_ , \new_[1904]_ ,
    \new_[1905]_ , \new_[1906]_ , \new_[1907]_ , \new_[1908]_ ,
    \new_[1909]_ , \new_[1910]_ , \new_[1911]_ , \new_[1912]_ ,
    \new_[1913]_ , \new_[1914]_ , \new_[1915]_ , \new_[1916]_ ,
    \new_[1917]_ , \new_[1918]_ , \new_[1919]_ , \new_[1920]_ ,
    \new_[1921]_ , \new_[1922]_ , \new_[1923]_ , \new_[1924]_ ,
    \new_[1925]_ , \new_[1926]_ , \new_[1927]_ , \new_[1928]_ ,
    \new_[1929]_ , \new_[1930]_ , \new_[1931]_ , \new_[1932]_ ,
    \new_[1933]_ , \new_[1934]_ , \new_[1935]_ , \new_[1936]_ ,
    \new_[1937]_ , \new_[1938]_ , \new_[1939]_ , \new_[1940]_ ,
    \new_[1941]_ , \new_[1942]_ , \new_[1943]_ , \new_[1944]_ ,
    \new_[1945]_ , \new_[1946]_ , \new_[1947]_ , \new_[1948]_ ,
    \new_[1949]_ , \new_[1950]_ , \new_[1951]_ , \new_[1952]_ ,
    \new_[1953]_ , \new_[1954]_ , \new_[1955]_ , \new_[1956]_ ,
    \new_[1957]_ , \new_[1958]_ , \new_[1959]_ , \new_[1960]_ ,
    \new_[1961]_ , \new_[1962]_ , \new_[1963]_ , \new_[1964]_ ,
    \new_[1965]_ , \new_[1966]_ , \new_[1967]_ , \new_[1968]_ ,
    \new_[1969]_ , \new_[1970]_ , \new_[1971]_ , \new_[1972]_ ,
    \new_[1973]_ , \new_[1974]_ , \new_[1975]_ , \new_[1976]_ ,
    \new_[1977]_ , \new_[1978]_ , \new_[1979]_ , \new_[1980]_ ,
    \new_[1981]_ , \new_[1982]_ , \new_[1983]_ , \new_[1984]_ ,
    \new_[1985]_ , \new_[1986]_ , \new_[1987]_ , \new_[1988]_ ,
    \new_[1989]_ , \new_[1990]_ , \new_[1991]_ , \new_[1992]_ ,
    \new_[1993]_ , \new_[1994]_ , \new_[1995]_ , \new_[1996]_ ,
    \new_[1997]_ , \new_[1998]_ , \new_[1999]_ , \new_[2000]_ ,
    \new_[2001]_ , \new_[2002]_ , \new_[2003]_ , \new_[2004]_ ,
    \new_[2005]_ , \new_[2006]_ , \new_[2007]_ , \new_[2008]_ ,
    \new_[2009]_ , \new_[2010]_ , \new_[2011]_ , \new_[2012]_ ,
    \new_[2013]_ , \new_[2014]_ , \new_[2015]_ , \new_[2016]_ ,
    \new_[2017]_ , \new_[2018]_ , \new_[2019]_ , \new_[2020]_ ,
    \new_[2021]_ , \new_[2022]_ , \new_[2023]_ , \new_[2024]_ ,
    \new_[2025]_ , \new_[2026]_ , \new_[2027]_ , \new_[2028]_ ,
    \new_[2029]_ , \new_[2030]_ , \new_[2031]_ , \new_[2032]_ ,
    \new_[2033]_ , \new_[2034]_ , \new_[2035]_ , \new_[2036]_ ,
    \new_[2037]_ , \new_[2038]_ , \new_[2039]_ , \new_[2040]_ ,
    \new_[2041]_ , \new_[2042]_ , \new_[2043]_ , \new_[2044]_ ,
    \new_[2045]_ , \new_[2046]_ , \new_[2047]_ , \new_[2048]_ ,
    \new_[2049]_ , \new_[2050]_ , \new_[2051]_ , \new_[2052]_ ,
    \new_[2053]_ , \new_[2054]_ , \new_[2055]_ , \new_[2056]_ ,
    \new_[2057]_ , \new_[2058]_ , \new_[2059]_ , \new_[2060]_ ,
    \new_[2061]_ , \new_[2062]_ , \new_[2063]_ , \new_[2064]_ ,
    \new_[2065]_ , \new_[2066]_ , \new_[2067]_ , \new_[2068]_ ,
    \new_[2069]_ , \new_[2070]_ , \new_[2071]_ , \new_[2072]_ ,
    \new_[2073]_ , \new_[2074]_ , \new_[2075]_ , \new_[2076]_ ,
    \new_[2077]_ , \new_[2078]_ , \new_[2079]_ , \new_[2080]_ ,
    \new_[2081]_ , \new_[2082]_ , \new_[2083]_ , \new_[2084]_ ,
    \new_[2085]_ , \new_[2086]_ , \new_[2087]_ , \new_[2088]_ ,
    \new_[2089]_ , \new_[2090]_ , \new_[2091]_ , \new_[2092]_ ,
    \new_[2093]_ , \new_[2094]_ , \new_[2095]_ , \new_[2096]_ ,
    \new_[2097]_ , \new_[2098]_ , \new_[2099]_ , \new_[2100]_ ,
    \new_[2101]_ , \new_[2102]_ , \new_[2103]_ , \new_[2104]_ ,
    \new_[2105]_ , \new_[2106]_ , \new_[2107]_ , \new_[2108]_ ,
    \new_[2109]_ , \new_[2110]_ , \new_[2111]_ , \new_[2112]_ ,
    \new_[2113]_ , \new_[2114]_ , \new_[2115]_ , \new_[2116]_ ,
    \new_[2117]_ , \new_[2118]_ , \new_[2119]_ , \new_[2120]_ ,
    \new_[2121]_ , \new_[2122]_ , \new_[2123]_ , \new_[2124]_ ,
    \new_[2125]_ , \new_[2126]_ , \new_[2127]_ , \new_[2128]_ ,
    \new_[2129]_ , \new_[2130]_ , \new_[2131]_ , \new_[2132]_ ,
    \new_[2133]_ , \new_[2134]_ , \new_[2135]_ , \new_[2136]_ ,
    \new_[2137]_ , \new_[2138]_ , \new_[2139]_ , \new_[2140]_ ,
    \new_[2141]_ , \new_[2142]_ , \new_[2143]_ , \new_[2144]_ ,
    \new_[2145]_ , \new_[2146]_ , \new_[2147]_ , \new_[2148]_ ,
    \new_[2149]_ , \new_[2150]_ , \new_[2151]_ , \new_[2152]_ ,
    \new_[2153]_ , \new_[2154]_ , \new_[2155]_ , \new_[2156]_ ,
    \new_[2157]_ , \new_[2158]_ , \new_[2159]_ , \new_[2160]_ ,
    \new_[2161]_ , \new_[2162]_ , \new_[2163]_ , \new_[2164]_ ,
    \new_[2165]_ , \new_[2166]_ , \new_[2167]_ , \new_[2168]_ ,
    \new_[2169]_ , \new_[2170]_ , \new_[2171]_ , \new_[2172]_ ,
    \new_[2173]_ , \new_[2174]_ , \new_[2175]_ , \new_[2176]_ ,
    \new_[2177]_ , \new_[2178]_ , \new_[2179]_ , \new_[2180]_ ,
    \new_[2181]_ , \new_[2182]_ , \new_[2183]_ , \new_[2184]_ ,
    \new_[2185]_ , \new_[2186]_ , \new_[2187]_ , \new_[2188]_ ,
    \new_[2189]_ , \new_[2190]_ , \new_[2191]_ , \new_[2192]_ ,
    \new_[2193]_ , \new_[2194]_ , \new_[2195]_ , \new_[2196]_ ,
    \new_[2197]_ , \new_[2198]_ , \new_[2199]_ , \new_[2200]_ ,
    \new_[2201]_ , \new_[2202]_ , \new_[2203]_ , \new_[2204]_ ,
    \new_[2205]_ , \new_[2206]_ , \new_[2207]_ , \new_[2208]_ ,
    \new_[2209]_ , \new_[2210]_ , \new_[2211]_ , \new_[2212]_ ,
    \new_[2213]_ , \new_[2214]_ , \new_[2215]_ , \new_[2216]_ ,
    \new_[2217]_ , \new_[2218]_ , \new_[2219]_ , \new_[2220]_ ,
    \new_[2221]_ , \new_[2222]_ , \new_[2223]_ , \new_[2224]_ ,
    \new_[2225]_ , \new_[2226]_ , \new_[2227]_ , \new_[2228]_ ,
    \new_[2229]_ , \new_[2230]_ , \new_[2231]_ , \new_[2232]_ ,
    \new_[2233]_ , \new_[2234]_ , \new_[2235]_ , \new_[2236]_ ,
    \new_[2237]_ , \new_[2238]_ , \new_[2239]_ , \new_[2240]_ ,
    \new_[2241]_ , \new_[2242]_ , \new_[2243]_ , \new_[2244]_ ,
    \new_[2245]_ , \new_[2246]_ , \new_[2247]_ , \new_[2248]_ ,
    \new_[2249]_ , \new_[2250]_ , \new_[2251]_ , \new_[2252]_ ,
    \new_[2253]_ , \new_[2254]_ , \new_[2255]_ , \new_[2256]_ ,
    \new_[2257]_ , \new_[2258]_ , \new_[2259]_ , \new_[2260]_ ,
    \new_[2261]_ , \new_[2262]_ , \new_[2263]_ , \new_[2264]_ ,
    \new_[2265]_ , \new_[2266]_ , \new_[2267]_ , \new_[2268]_ ,
    \new_[2269]_ , \new_[2270]_ , \new_[2271]_ , \new_[2272]_ ,
    \new_[2273]_ , \new_[2274]_ , \new_[2275]_ , \new_[2276]_ ,
    \new_[2277]_ , \new_[2278]_ , \new_[2279]_ , \new_[2280]_ ,
    \new_[2281]_ , \new_[2282]_ , \new_[2283]_ , \new_[2284]_ ,
    \new_[2285]_ , \new_[2286]_ , \new_[2287]_ , \new_[2288]_ ,
    \new_[2289]_ , \new_[2290]_ , \new_[2291]_ , \new_[2292]_ ,
    \new_[2293]_ , \new_[2294]_ , \new_[2295]_ , \new_[2296]_ ,
    \new_[2297]_ , \new_[2298]_ , \new_[2299]_ , \new_[2300]_ ,
    \new_[2301]_ , \new_[2302]_ , \new_[2303]_ , \new_[2304]_ ,
    \new_[2305]_ , \new_[2306]_ , \new_[2307]_ , \new_[2308]_ ,
    \new_[2309]_ , \new_[2310]_ , \new_[2313]_ , \new_[2316]_ ,
    \new_[2317]_ , \new_[2320]_ , \new_[2324]_ , \new_[2325]_ ,
    \new_[2326]_ , \new_[2327]_ , \new_[2330]_ , \new_[2333]_ ,
    \new_[2334]_ , \new_[2337]_ , \new_[2341]_ , \new_[2342]_ ,
    \new_[2343]_ , \new_[2344]_ , \new_[2345]_ , \new_[2348]_ ,
    \new_[2351]_ , \new_[2352]_ , \new_[2355]_ , \new_[2359]_ ,
    \new_[2360]_ , \new_[2361]_ , \new_[2362]_ , \new_[2365]_ ,
    \new_[2368]_ , \new_[2369]_ , \new_[2372]_ , \new_[2376]_ ,
    \new_[2377]_ , \new_[2378]_ , \new_[2379]_ , \new_[2380]_ ,
    \new_[2381]_ , \new_[2384]_ , \new_[2387]_ , \new_[2388]_ ,
    \new_[2391]_ , \new_[2395]_ , \new_[2396]_ , \new_[2397]_ ,
    \new_[2398]_ , \new_[2401]_ , \new_[2404]_ , \new_[2405]_ ,
    \new_[2408]_ , \new_[2412]_ , \new_[2413]_ , \new_[2414]_ ,
    \new_[2415]_ , \new_[2416]_ , \new_[2419]_ , \new_[2422]_ ,
    \new_[2423]_ , \new_[2426]_ , \new_[2430]_ , \new_[2431]_ ,
    \new_[2432]_ , \new_[2433]_ , \new_[2436]_ , \new_[2439]_ ,
    \new_[2440]_ , \new_[2443]_ , \new_[2447]_ , \new_[2448]_ ,
    \new_[2449]_ , \new_[2450]_ , \new_[2451]_ , \new_[2452]_ ,
    \new_[2453]_ , \new_[2456]_ , \new_[2459]_ , \new_[2460]_ ,
    \new_[2463]_ , \new_[2467]_ , \new_[2468]_ , \new_[2469]_ ,
    \new_[2470]_ , \new_[2473]_ , \new_[2476]_ , \new_[2477]_ ,
    \new_[2480]_ , \new_[2484]_ , \new_[2485]_ , \new_[2486]_ ,
    \new_[2487]_ , \new_[2488]_ , \new_[2491]_ , \new_[2494]_ ,
    \new_[2495]_ , \new_[2498]_ , \new_[2502]_ , \new_[2503]_ ,
    \new_[2504]_ , \new_[2505]_ , \new_[2508]_ , \new_[2511]_ ,
    \new_[2512]_ , \new_[2515]_ , \new_[2519]_ , \new_[2520]_ ,
    \new_[2521]_ , \new_[2522]_ , \new_[2523]_ , \new_[2524]_ ,
    \new_[2527]_ , \new_[2530]_ , \new_[2531]_ , \new_[2534]_ ,
    \new_[2538]_ , \new_[2539]_ , \new_[2540]_ , \new_[2541]_ ,
    \new_[2544]_ , \new_[2547]_ , \new_[2548]_ , \new_[2551]_ ,
    \new_[2555]_ , \new_[2556]_ , \new_[2557]_ , \new_[2558]_ ,
    \new_[2559]_ , \new_[2562]_ , \new_[2565]_ , \new_[2566]_ ,
    \new_[2569]_ , \new_[2573]_ , \new_[2574]_ , \new_[2575]_ ,
    \new_[2576]_ , \new_[2579]_ , \new_[2582]_ , \new_[2583]_ ,
    \new_[2586]_ , \new_[2590]_ , \new_[2591]_ , \new_[2592]_ ,
    \new_[2593]_ , \new_[2594]_ , \new_[2595]_ , \new_[2596]_ ,
    \new_[2597]_ , \new_[2600]_ , \new_[2603]_ , \new_[2604]_ ,
    \new_[2607]_ , \new_[2611]_ , \new_[2612]_ , \new_[2613]_ ,
    \new_[2614]_ , \new_[2617]_ , \new_[2620]_ , \new_[2621]_ ,
    \new_[2624]_ , \new_[2628]_ , \new_[2629]_ , \new_[2630]_ ,
    \new_[2631]_ , \new_[2632]_ , \new_[2635]_ , \new_[2638]_ ,
    \new_[2639]_ , \new_[2642]_ , \new_[2646]_ , \new_[2647]_ ,
    \new_[2648]_ , \new_[2649]_ , \new_[2652]_ , \new_[2655]_ ,
    \new_[2656]_ , \new_[2659]_ , \new_[2663]_ , \new_[2664]_ ,
    \new_[2665]_ , \new_[2666]_ , \new_[2667]_ , \new_[2668]_ ,
    \new_[2671]_ , \new_[2674]_ , \new_[2675]_ , \new_[2678]_ ,
    \new_[2682]_ , \new_[2683]_ , \new_[2684]_ , \new_[2685]_ ,
    \new_[2688]_ , \new_[2691]_ , \new_[2692]_ , \new_[2695]_ ,
    \new_[2699]_ , \new_[2700]_ , \new_[2701]_ , \new_[2702]_ ,
    \new_[2703]_ , \new_[2706]_ , \new_[2709]_ , \new_[2710]_ ,
    \new_[2713]_ , \new_[2717]_ , \new_[2718]_ , \new_[2719]_ ,
    \new_[2720]_ , \new_[2723]_ , \new_[2726]_ , \new_[2727]_ ,
    \new_[2730]_ , \new_[2734]_ , \new_[2735]_ , \new_[2736]_ ,
    \new_[2737]_ , \new_[2738]_ , \new_[2739]_ , \new_[2740]_ ,
    \new_[2743]_ , \new_[2746]_ , \new_[2747]_ , \new_[2750]_ ,
    \new_[2754]_ , \new_[2755]_ , \new_[2756]_ , \new_[2757]_ ,
    \new_[2760]_ , \new_[2763]_ , \new_[2764]_ , \new_[2767]_ ,
    \new_[2771]_ , \new_[2772]_ , \new_[2773]_ , \new_[2774]_ ,
    \new_[2775]_ , \new_[2778]_ , \new_[2781]_ , \new_[2782]_ ,
    \new_[2785]_ , \new_[2789]_ , \new_[2790]_ , \new_[2791]_ ,
    \new_[2792]_ , \new_[2795]_ , \new_[2798]_ , \new_[2799]_ ,
    \new_[2802]_ , \new_[2806]_ , \new_[2807]_ , \new_[2808]_ ,
    \new_[2809]_ , \new_[2810]_ , \new_[2811]_ , \new_[2814]_ ,
    \new_[2817]_ , \new_[2818]_ , \new_[2821]_ , \new_[2825]_ ,
    \new_[2826]_ , \new_[2827]_ , \new_[2828]_ , \new_[2831]_ ,
    \new_[2834]_ , \new_[2835]_ , \new_[2838]_ , \new_[2842]_ ,
    \new_[2843]_ , \new_[2844]_ , \new_[2845]_ , \new_[2846]_ ,
    \new_[2849]_ , \new_[2852]_ , \new_[2853]_ , \new_[2856]_ ,
    \new_[2860]_ , \new_[2861]_ , \new_[2862]_ , \new_[2863]_ ,
    \new_[2866]_ , \new_[2869]_ , \new_[2870]_ , \new_[2873]_ ,
    \new_[2877]_ , \new_[2878]_ , \new_[2879]_ , \new_[2880]_ ,
    \new_[2881]_ , \new_[2882]_ , \new_[2883]_ , \new_[2884]_ ,
    \new_[2885]_ , \new_[2888]_ , \new_[2891]_ , \new_[2892]_ ,
    \new_[2895]_ , \new_[2899]_ , \new_[2900]_ , \new_[2901]_ ,
    \new_[2902]_ , \new_[2905]_ , \new_[2908]_ , \new_[2909]_ ,
    \new_[2912]_ , \new_[2916]_ , \new_[2917]_ , \new_[2918]_ ,
    \new_[2919]_ , \new_[2920]_ , \new_[2923]_ , \new_[2926]_ ,
    \new_[2927]_ , \new_[2930]_ , \new_[2934]_ , \new_[2935]_ ,
    \new_[2936]_ , \new_[2937]_ , \new_[2940]_ , \new_[2943]_ ,
    \new_[2944]_ , \new_[2947]_ , \new_[2951]_ , \new_[2952]_ ,
    \new_[2953]_ , \new_[2954]_ , \new_[2955]_ , \new_[2956]_ ,
    \new_[2959]_ , \new_[2962]_ , \new_[2963]_ , \new_[2966]_ ,
    \new_[2970]_ , \new_[2971]_ , \new_[2972]_ , \new_[2973]_ ,
    \new_[2976]_ , \new_[2979]_ , \new_[2980]_ , \new_[2983]_ ,
    \new_[2987]_ , \new_[2988]_ , \new_[2989]_ , \new_[2990]_ ,
    \new_[2991]_ , \new_[2994]_ , \new_[2997]_ , \new_[2998]_ ,
    \new_[3001]_ , \new_[3005]_ , \new_[3006]_ , \new_[3007]_ ,
    \new_[3008]_ , \new_[3011]_ , \new_[3014]_ , \new_[3015]_ ,
    \new_[3018]_ , \new_[3022]_ , \new_[3023]_ , \new_[3024]_ ,
    \new_[3025]_ , \new_[3026]_ , \new_[3027]_ , \new_[3028]_ ,
    \new_[3031]_ , \new_[3034]_ , \new_[3035]_ , \new_[3038]_ ,
    \new_[3042]_ , \new_[3043]_ , \new_[3044]_ , \new_[3045]_ ,
    \new_[3048]_ , \new_[3051]_ , \new_[3052]_ , \new_[3055]_ ,
    \new_[3059]_ , \new_[3060]_ , \new_[3061]_ , \new_[3062]_ ,
    \new_[3063]_ , \new_[3066]_ , \new_[3069]_ , \new_[3070]_ ,
    \new_[3073]_ , \new_[3077]_ , \new_[3078]_ , \new_[3079]_ ,
    \new_[3080]_ , \new_[3083]_ , \new_[3086]_ , \new_[3087]_ ,
    \new_[3090]_ , \new_[3094]_ , \new_[3095]_ , \new_[3096]_ ,
    \new_[3097]_ , \new_[3098]_ , \new_[3099]_ , \new_[3102]_ ,
    \new_[3105]_ , \new_[3106]_ , \new_[3109]_ , \new_[3113]_ ,
    \new_[3114]_ , \new_[3115]_ , \new_[3116]_ , \new_[3119]_ ,
    \new_[3122]_ , \new_[3123]_ , \new_[3126]_ , \new_[3130]_ ,
    \new_[3131]_ , \new_[3132]_ , \new_[3133]_ , \new_[3134]_ ,
    \new_[3137]_ , \new_[3140]_ , \new_[3141]_ , \new_[3144]_ ,
    \new_[3148]_ , \new_[3149]_ , \new_[3150]_ , \new_[3151]_ ,
    \new_[3154]_ , \new_[3157]_ , \new_[3158]_ , \new_[3161]_ ,
    \new_[3165]_ , \new_[3166]_ , \new_[3167]_ , \new_[3168]_ ,
    \new_[3169]_ , \new_[3170]_ , \new_[3171]_ , \new_[3172]_ ,
    \new_[3175]_ , \new_[3178]_ , \new_[3179]_ , \new_[3182]_ ,
    \new_[3186]_ , \new_[3187]_ , \new_[3188]_ , \new_[3189]_ ,
    \new_[3192]_ , \new_[3195]_ , \new_[3196]_ , \new_[3199]_ ,
    \new_[3203]_ , \new_[3204]_ , \new_[3205]_ , \new_[3206]_ ,
    \new_[3207]_ , \new_[3210]_ , \new_[3213]_ , \new_[3214]_ ,
    \new_[3217]_ , \new_[3221]_ , \new_[3222]_ , \new_[3223]_ ,
    \new_[3224]_ , \new_[3227]_ , \new_[3230]_ , \new_[3231]_ ,
    \new_[3234]_ , \new_[3238]_ , \new_[3239]_ , \new_[3240]_ ,
    \new_[3241]_ , \new_[3242]_ , \new_[3243]_ , \new_[3246]_ ,
    \new_[3249]_ , \new_[3250]_ , \new_[3253]_ , \new_[3257]_ ,
    \new_[3258]_ , \new_[3259]_ , \new_[3260]_ , \new_[3263]_ ,
    \new_[3266]_ , \new_[3267]_ , \new_[3270]_ , \new_[3274]_ ,
    \new_[3275]_ , \new_[3276]_ , \new_[3277]_ , \new_[3278]_ ,
    \new_[3281]_ , \new_[3284]_ , \new_[3285]_ , \new_[3288]_ ,
    \new_[3292]_ , \new_[3293]_ , \new_[3294]_ , \new_[3295]_ ,
    \new_[3298]_ , \new_[3301]_ , \new_[3302]_ , \new_[3305]_ ,
    \new_[3309]_ , \new_[3310]_ , \new_[3311]_ , \new_[3312]_ ,
    \new_[3313]_ , \new_[3314]_ , \new_[3315]_ , \new_[3318]_ ,
    \new_[3321]_ , \new_[3322]_ , \new_[3325]_ , \new_[3329]_ ,
    \new_[3330]_ , \new_[3331]_ , \new_[3332]_ , \new_[3335]_ ,
    \new_[3338]_ , \new_[3339]_ , \new_[3342]_ , \new_[3346]_ ,
    \new_[3347]_ , \new_[3348]_ , \new_[3349]_ , \new_[3350]_ ,
    \new_[3353]_ , \new_[3356]_ , \new_[3357]_ , \new_[3360]_ ,
    \new_[3364]_ , \new_[3365]_ , \new_[3366]_ , \new_[3367]_ ,
    \new_[3370]_ , \new_[3373]_ , \new_[3374]_ , \new_[3377]_ ,
    \new_[3381]_ , \new_[3382]_ , \new_[3383]_ , \new_[3384]_ ,
    \new_[3385]_ , \new_[3386]_ , \new_[3389]_ , \new_[3392]_ ,
    \new_[3393]_ , \new_[3396]_ , \new_[3400]_ , \new_[3401]_ ,
    \new_[3402]_ , \new_[3403]_ , \new_[3406]_ , \new_[3409]_ ,
    \new_[3410]_ , \new_[3413]_ , \new_[3417]_ , \new_[3418]_ ,
    \new_[3419]_ , \new_[3420]_ , \new_[3421]_ , \new_[3424]_ ,
    \new_[3427]_ , \new_[3428]_ , \new_[3431]_ , \new_[3435]_ ,
    \new_[3436]_ , \new_[3437]_ , \new_[3438]_ , \new_[3441]_ ,
    \new_[3445]_ , \new_[3446]_ , \new_[3447]_ , \new_[3450]_ ,
    \new_[3454]_ , \new_[3455]_ , \new_[3456]_ , \new_[3457]_ ,
    \new_[3458]_ , \new_[3459]_ , \new_[3460]_ , \new_[3461]_ ,
    \new_[3462]_ , \new_[3463]_ , \new_[3466]_ , \new_[3469]_ ,
    \new_[3470]_ , \new_[3473]_ , \new_[3477]_ , \new_[3478]_ ,
    \new_[3479]_ , \new_[3480]_ , \new_[3483]_ , \new_[3486]_ ,
    \new_[3487]_ , \new_[3490]_ , \new_[3494]_ , \new_[3495]_ ,
    \new_[3496]_ , \new_[3497]_ , \new_[3498]_ , \new_[3501]_ ,
    \new_[3504]_ , \new_[3505]_ , \new_[3508]_ , \new_[3512]_ ,
    \new_[3513]_ , \new_[3514]_ , \new_[3515]_ , \new_[3518]_ ,
    \new_[3521]_ , \new_[3522]_ , \new_[3525]_ , \new_[3529]_ ,
    \new_[3530]_ , \new_[3531]_ , \new_[3532]_ , \new_[3533]_ ,
    \new_[3534]_ , \new_[3537]_ , \new_[3540]_ , \new_[3541]_ ,
    \new_[3544]_ , \new_[3548]_ , \new_[3549]_ , \new_[3550]_ ,
    \new_[3551]_ , \new_[3554]_ , \new_[3557]_ , \new_[3558]_ ,
    \new_[3561]_ , \new_[3565]_ , \new_[3566]_ , \new_[3567]_ ,
    \new_[3568]_ , \new_[3569]_ , \new_[3572]_ , \new_[3575]_ ,
    \new_[3576]_ , \new_[3579]_ , \new_[3583]_ , \new_[3584]_ ,
    \new_[3585]_ , \new_[3586]_ , \new_[3589]_ , \new_[3592]_ ,
    \new_[3593]_ , \new_[3596]_ , \new_[3600]_ , \new_[3601]_ ,
    \new_[3602]_ , \new_[3603]_ , \new_[3604]_ , \new_[3605]_ ,
    \new_[3606]_ , \new_[3609]_ , \new_[3612]_ , \new_[3613]_ ,
    \new_[3616]_ , \new_[3620]_ , \new_[3621]_ , \new_[3622]_ ,
    \new_[3623]_ , \new_[3626]_ , \new_[3629]_ , \new_[3630]_ ,
    \new_[3633]_ , \new_[3637]_ , \new_[3638]_ , \new_[3639]_ ,
    \new_[3640]_ , \new_[3641]_ , \new_[3644]_ , \new_[3647]_ ,
    \new_[3648]_ , \new_[3651]_ , \new_[3655]_ , \new_[3656]_ ,
    \new_[3657]_ , \new_[3658]_ , \new_[3661]_ , \new_[3664]_ ,
    \new_[3665]_ , \new_[3668]_ , \new_[3672]_ , \new_[3673]_ ,
    \new_[3674]_ , \new_[3675]_ , \new_[3676]_ , \new_[3677]_ ,
    \new_[3680]_ , \new_[3683]_ , \new_[3684]_ , \new_[3687]_ ,
    \new_[3691]_ , \new_[3692]_ , \new_[3693]_ , \new_[3694]_ ,
    \new_[3697]_ , \new_[3700]_ , \new_[3701]_ , \new_[3704]_ ,
    \new_[3708]_ , \new_[3709]_ , \new_[3710]_ , \new_[3711]_ ,
    \new_[3712]_ , \new_[3715]_ , \new_[3718]_ , \new_[3719]_ ,
    \new_[3722]_ , \new_[3726]_ , \new_[3727]_ , \new_[3728]_ ,
    \new_[3729]_ , \new_[3732]_ , \new_[3735]_ , \new_[3736]_ ,
    \new_[3739]_ , \new_[3743]_ , \new_[3744]_ , \new_[3745]_ ,
    \new_[3746]_ , \new_[3747]_ , \new_[3748]_ , \new_[3749]_ ,
    \new_[3750]_ , \new_[3753]_ , \new_[3756]_ , \new_[3757]_ ,
    \new_[3760]_ , \new_[3764]_ , \new_[3765]_ , \new_[3766]_ ,
    \new_[3767]_ , \new_[3770]_ , \new_[3773]_ , \new_[3774]_ ,
    \new_[3777]_ , \new_[3781]_ , \new_[3782]_ , \new_[3783]_ ,
    \new_[3784]_ , \new_[3785]_ , \new_[3788]_ , \new_[3791]_ ,
    \new_[3792]_ , \new_[3795]_ , \new_[3799]_ , \new_[3800]_ ,
    \new_[3801]_ , \new_[3802]_ , \new_[3805]_ , \new_[3808]_ ,
    \new_[3809]_ , \new_[3812]_ , \new_[3816]_ , \new_[3817]_ ,
    \new_[3818]_ , \new_[3819]_ , \new_[3820]_ , \new_[3821]_ ,
    \new_[3824]_ , \new_[3827]_ , \new_[3828]_ , \new_[3831]_ ,
    \new_[3835]_ , \new_[3836]_ , \new_[3837]_ , \new_[3838]_ ,
    \new_[3841]_ , \new_[3844]_ , \new_[3845]_ , \new_[3848]_ ,
    \new_[3852]_ , \new_[3853]_ , \new_[3854]_ , \new_[3855]_ ,
    \new_[3856]_ , \new_[3859]_ , \new_[3862]_ , \new_[3863]_ ,
    \new_[3866]_ , \new_[3870]_ , \new_[3871]_ , \new_[3872]_ ,
    \new_[3873]_ , \new_[3876]_ , \new_[3879]_ , \new_[3880]_ ,
    \new_[3883]_ , \new_[3887]_ , \new_[3888]_ , \new_[3889]_ ,
    \new_[3890]_ , \new_[3891]_ , \new_[3892]_ , \new_[3893]_ ,
    \new_[3896]_ , \new_[3899]_ , \new_[3900]_ , \new_[3903]_ ,
    \new_[3907]_ , \new_[3908]_ , \new_[3909]_ , \new_[3910]_ ,
    \new_[3913]_ , \new_[3916]_ , \new_[3917]_ , \new_[3920]_ ,
    \new_[3924]_ , \new_[3925]_ , \new_[3926]_ , \new_[3927]_ ,
    \new_[3928]_ , \new_[3931]_ , \new_[3934]_ , \new_[3935]_ ,
    \new_[3938]_ , \new_[3942]_ , \new_[3943]_ , \new_[3944]_ ,
    \new_[3945]_ , \new_[3948]_ , \new_[3951]_ , \new_[3952]_ ,
    \new_[3955]_ , \new_[3959]_ , \new_[3960]_ , \new_[3961]_ ,
    \new_[3962]_ , \new_[3963]_ , \new_[3964]_ , \new_[3967]_ ,
    \new_[3970]_ , \new_[3971]_ , \new_[3974]_ , \new_[3978]_ ,
    \new_[3979]_ , \new_[3980]_ , \new_[3981]_ , \new_[3984]_ ,
    \new_[3987]_ , \new_[3988]_ , \new_[3991]_ , \new_[3995]_ ,
    \new_[3996]_ , \new_[3997]_ , \new_[3998]_ , \new_[3999]_ ,
    \new_[4002]_ , \new_[4005]_ , \new_[4006]_ , \new_[4009]_ ,
    \new_[4013]_ , \new_[4014]_ , \new_[4015]_ , \new_[4016]_ ,
    \new_[4019]_ , \new_[4023]_ , \new_[4024]_ , \new_[4025]_ ,
    \new_[4028]_ , \new_[4032]_ , \new_[4033]_ , \new_[4034]_ ,
    \new_[4035]_ , \new_[4036]_ , \new_[4037]_ , \new_[4038]_ ,
    \new_[4039]_ , \new_[4040]_ , \new_[4043]_ , \new_[4046]_ ,
    \new_[4047]_ , \new_[4050]_ , \new_[4054]_ , \new_[4055]_ ,
    \new_[4056]_ , \new_[4057]_ , \new_[4060]_ , \new_[4063]_ ,
    \new_[4064]_ , \new_[4067]_ , \new_[4071]_ , \new_[4072]_ ,
    \new_[4073]_ , \new_[4074]_ , \new_[4075]_ , \new_[4078]_ ,
    \new_[4081]_ , \new_[4082]_ , \new_[4085]_ , \new_[4089]_ ,
    \new_[4090]_ , \new_[4091]_ , \new_[4092]_ , \new_[4095]_ ,
    \new_[4098]_ , \new_[4099]_ , \new_[4102]_ , \new_[4106]_ ,
    \new_[4107]_ , \new_[4108]_ , \new_[4109]_ , \new_[4110]_ ,
    \new_[4111]_ , \new_[4114]_ , \new_[4117]_ , \new_[4118]_ ,
    \new_[4121]_ , \new_[4125]_ , \new_[4126]_ , \new_[4127]_ ,
    \new_[4128]_ , \new_[4131]_ , \new_[4134]_ , \new_[4135]_ ,
    \new_[4138]_ , \new_[4142]_ , \new_[4143]_ , \new_[4144]_ ,
    \new_[4145]_ , \new_[4146]_ , \new_[4149]_ , \new_[4152]_ ,
    \new_[4153]_ , \new_[4156]_ , \new_[4160]_ , \new_[4161]_ ,
    \new_[4162]_ , \new_[4163]_ , \new_[4166]_ , \new_[4169]_ ,
    \new_[4170]_ , \new_[4173]_ , \new_[4177]_ , \new_[4178]_ ,
    \new_[4179]_ , \new_[4180]_ , \new_[4181]_ , \new_[4182]_ ,
    \new_[4183]_ , \new_[4186]_ , \new_[4189]_ , \new_[4190]_ ,
    \new_[4193]_ , \new_[4197]_ , \new_[4198]_ , \new_[4199]_ ,
    \new_[4200]_ , \new_[4203]_ , \new_[4206]_ , \new_[4207]_ ,
    \new_[4210]_ , \new_[4214]_ , \new_[4215]_ , \new_[4216]_ ,
    \new_[4217]_ , \new_[4218]_ , \new_[4221]_ , \new_[4224]_ ,
    \new_[4225]_ , \new_[4228]_ , \new_[4232]_ , \new_[4233]_ ,
    \new_[4234]_ , \new_[4235]_ , \new_[4238]_ , \new_[4241]_ ,
    \new_[4242]_ , \new_[4245]_ , \new_[4249]_ , \new_[4250]_ ,
    \new_[4251]_ , \new_[4252]_ , \new_[4253]_ , \new_[4254]_ ,
    \new_[4257]_ , \new_[4260]_ , \new_[4261]_ , \new_[4264]_ ,
    \new_[4268]_ , \new_[4269]_ , \new_[4270]_ , \new_[4271]_ ,
    \new_[4274]_ , \new_[4277]_ , \new_[4278]_ , \new_[4281]_ ,
    \new_[4285]_ , \new_[4286]_ , \new_[4287]_ , \new_[4288]_ ,
    \new_[4289]_ , \new_[4292]_ , \new_[4295]_ , \new_[4296]_ ,
    \new_[4299]_ , \new_[4303]_ , \new_[4304]_ , \new_[4305]_ ,
    \new_[4306]_ , \new_[4309]_ , \new_[4312]_ , \new_[4313]_ ,
    \new_[4316]_ , \new_[4320]_ , \new_[4321]_ , \new_[4322]_ ,
    \new_[4323]_ , \new_[4324]_ , \new_[4325]_ , \new_[4326]_ ,
    \new_[4327]_ , \new_[4330]_ , \new_[4333]_ , \new_[4334]_ ,
    \new_[4337]_ , \new_[4341]_ , \new_[4342]_ , \new_[4343]_ ,
    \new_[4344]_ , \new_[4347]_ , \new_[4350]_ , \new_[4351]_ ,
    \new_[4354]_ , \new_[4358]_ , \new_[4359]_ , \new_[4360]_ ,
    \new_[4361]_ , \new_[4362]_ , \new_[4365]_ , \new_[4368]_ ,
    \new_[4369]_ , \new_[4372]_ , \new_[4376]_ , \new_[4377]_ ,
    \new_[4378]_ , \new_[4379]_ , \new_[4382]_ , \new_[4385]_ ,
    \new_[4386]_ , \new_[4389]_ , \new_[4393]_ , \new_[4394]_ ,
    \new_[4395]_ , \new_[4396]_ , \new_[4397]_ , \new_[4398]_ ,
    \new_[4401]_ , \new_[4404]_ , \new_[4405]_ , \new_[4408]_ ,
    \new_[4412]_ , \new_[4413]_ , \new_[4414]_ , \new_[4415]_ ,
    \new_[4418]_ , \new_[4421]_ , \new_[4422]_ , \new_[4425]_ ,
    \new_[4429]_ , \new_[4430]_ , \new_[4431]_ , \new_[4432]_ ,
    \new_[4433]_ , \new_[4436]_ , \new_[4439]_ , \new_[4440]_ ,
    \new_[4443]_ , \new_[4447]_ , \new_[4448]_ , \new_[4449]_ ,
    \new_[4450]_ , \new_[4453]_ , \new_[4456]_ , \new_[4457]_ ,
    \new_[4460]_ , \new_[4464]_ , \new_[4465]_ , \new_[4466]_ ,
    \new_[4467]_ , \new_[4468]_ , \new_[4469]_ , \new_[4470]_ ,
    \new_[4473]_ , \new_[4476]_ , \new_[4477]_ , \new_[4480]_ ,
    \new_[4484]_ , \new_[4485]_ , \new_[4486]_ , \new_[4487]_ ,
    \new_[4490]_ , \new_[4493]_ , \new_[4494]_ , \new_[4497]_ ,
    \new_[4501]_ , \new_[4502]_ , \new_[4503]_ , \new_[4504]_ ,
    \new_[4505]_ , \new_[4508]_ , \new_[4511]_ , \new_[4512]_ ,
    \new_[4515]_ , \new_[4519]_ , \new_[4520]_ , \new_[4521]_ ,
    \new_[4522]_ , \new_[4525]_ , \new_[4528]_ , \new_[4529]_ ,
    \new_[4532]_ , \new_[4536]_ , \new_[4537]_ , \new_[4538]_ ,
    \new_[4539]_ , \new_[4540]_ , \new_[4541]_ , \new_[4544]_ ,
    \new_[4547]_ , \new_[4548]_ , \new_[4551]_ , \new_[4555]_ ,
    \new_[4556]_ , \new_[4557]_ , \new_[4558]_ , \new_[4561]_ ,
    \new_[4564]_ , \new_[4565]_ , \new_[4568]_ , \new_[4572]_ ,
    \new_[4573]_ , \new_[4574]_ , \new_[4575]_ , \new_[4576]_ ,
    \new_[4579]_ , \new_[4582]_ , \new_[4583]_ , \new_[4586]_ ,
    \new_[4590]_ , \new_[4591]_ , \new_[4592]_ , \new_[4593]_ ,
    \new_[4596]_ , \new_[4600]_ , \new_[4601]_ , \new_[4602]_ ,
    \new_[4605]_ , \new_[4609]_ , \new_[4610]_ , \new_[4611]_ ,
    \new_[4612]_ , \new_[4613]_ , \new_[4614]_ , \new_[4615]_ ,
    \new_[4616]_ , \new_[4617]_ , \new_[4618]_ , \new_[4619]_ ,
    \new_[4622]_ , \new_[4625]_ , \new_[4626]_ , \new_[4629]_ ,
    \new_[4633]_ , \new_[4634]_ , \new_[4635]_ , \new_[4636]_ ,
    \new_[4639]_ , \new_[4642]_ , \new_[4643]_ , \new_[4646]_ ,
    \new_[4650]_ , \new_[4651]_ , \new_[4652]_ , \new_[4653]_ ,
    \new_[4654]_ , \new_[4657]_ , \new_[4660]_ , \new_[4661]_ ,
    \new_[4664]_ , \new_[4668]_ , \new_[4669]_ , \new_[4670]_ ,
    \new_[4671]_ , \new_[4674]_ , \new_[4677]_ , \new_[4678]_ ,
    \new_[4681]_ , \new_[4685]_ , \new_[4686]_ , \new_[4687]_ ,
    \new_[4688]_ , \new_[4689]_ , \new_[4690]_ , \new_[4693]_ ,
    \new_[4696]_ , \new_[4697]_ , \new_[4700]_ , \new_[4704]_ ,
    \new_[4705]_ , \new_[4706]_ , \new_[4707]_ , \new_[4710]_ ,
    \new_[4713]_ , \new_[4714]_ , \new_[4717]_ , \new_[4721]_ ,
    \new_[4722]_ , \new_[4723]_ , \new_[4724]_ , \new_[4725]_ ,
    \new_[4728]_ , \new_[4731]_ , \new_[4732]_ , \new_[4735]_ ,
    \new_[4739]_ , \new_[4740]_ , \new_[4741]_ , \new_[4742]_ ,
    \new_[4745]_ , \new_[4748]_ , \new_[4749]_ , \new_[4752]_ ,
    \new_[4756]_ , \new_[4757]_ , \new_[4758]_ , \new_[4759]_ ,
    \new_[4760]_ , \new_[4761]_ , \new_[4762]_ , \new_[4765]_ ,
    \new_[4768]_ , \new_[4769]_ , \new_[4772]_ , \new_[4776]_ ,
    \new_[4777]_ , \new_[4778]_ , \new_[4779]_ , \new_[4782]_ ,
    \new_[4785]_ , \new_[4786]_ , \new_[4789]_ , \new_[4793]_ ,
    \new_[4794]_ , \new_[4795]_ , \new_[4796]_ , \new_[4797]_ ,
    \new_[4800]_ , \new_[4803]_ , \new_[4804]_ , \new_[4807]_ ,
    \new_[4811]_ , \new_[4812]_ , \new_[4813]_ , \new_[4814]_ ,
    \new_[4817]_ , \new_[4820]_ , \new_[4821]_ , \new_[4824]_ ,
    \new_[4828]_ , \new_[4829]_ , \new_[4830]_ , \new_[4831]_ ,
    \new_[4832]_ , \new_[4833]_ , \new_[4836]_ , \new_[4839]_ ,
    \new_[4840]_ , \new_[4843]_ , \new_[4847]_ , \new_[4848]_ ,
    \new_[4849]_ , \new_[4850]_ , \new_[4853]_ , \new_[4856]_ ,
    \new_[4857]_ , \new_[4860]_ , \new_[4864]_ , \new_[4865]_ ,
    \new_[4866]_ , \new_[4867]_ , \new_[4868]_ , \new_[4871]_ ,
    \new_[4874]_ , \new_[4875]_ , \new_[4878]_ , \new_[4882]_ ,
    \new_[4883]_ , \new_[4884]_ , \new_[4885]_ , \new_[4888]_ ,
    \new_[4891]_ , \new_[4892]_ , \new_[4895]_ , \new_[4899]_ ,
    \new_[4900]_ , \new_[4901]_ , \new_[4902]_ , \new_[4903]_ ,
    \new_[4904]_ , \new_[4905]_ , \new_[4906]_ , \new_[4909]_ ,
    \new_[4912]_ , \new_[4913]_ , \new_[4916]_ , \new_[4920]_ ,
    \new_[4921]_ , \new_[4922]_ , \new_[4923]_ , \new_[4926]_ ,
    \new_[4929]_ , \new_[4930]_ , \new_[4933]_ , \new_[4937]_ ,
    \new_[4938]_ , \new_[4939]_ , \new_[4940]_ , \new_[4941]_ ,
    \new_[4944]_ , \new_[4947]_ , \new_[4948]_ , \new_[4951]_ ,
    \new_[4955]_ , \new_[4956]_ , \new_[4957]_ , \new_[4958]_ ,
    \new_[4961]_ , \new_[4964]_ , \new_[4965]_ , \new_[4968]_ ,
    \new_[4972]_ , \new_[4973]_ , \new_[4974]_ , \new_[4975]_ ,
    \new_[4976]_ , \new_[4977]_ , \new_[4980]_ , \new_[4983]_ ,
    \new_[4984]_ , \new_[4987]_ , \new_[4991]_ , \new_[4992]_ ,
    \new_[4993]_ , \new_[4994]_ , \new_[4997]_ , \new_[5000]_ ,
    \new_[5001]_ , \new_[5004]_ , \new_[5008]_ , \new_[5009]_ ,
    \new_[5010]_ , \new_[5011]_ , \new_[5012]_ , \new_[5015]_ ,
    \new_[5018]_ , \new_[5019]_ , \new_[5022]_ , \new_[5026]_ ,
    \new_[5027]_ , \new_[5028]_ , \new_[5029]_ , \new_[5032]_ ,
    \new_[5035]_ , \new_[5036]_ , \new_[5039]_ , \new_[5043]_ ,
    \new_[5044]_ , \new_[5045]_ , \new_[5046]_ , \new_[5047]_ ,
    \new_[5048]_ , \new_[5049]_ , \new_[5052]_ , \new_[5055]_ ,
    \new_[5056]_ , \new_[5059]_ , \new_[5063]_ , \new_[5064]_ ,
    \new_[5065]_ , \new_[5066]_ , \new_[5069]_ , \new_[5072]_ ,
    \new_[5073]_ , \new_[5076]_ , \new_[5080]_ , \new_[5081]_ ,
    \new_[5082]_ , \new_[5083]_ , \new_[5084]_ , \new_[5087]_ ,
    \new_[5090]_ , \new_[5091]_ , \new_[5094]_ , \new_[5098]_ ,
    \new_[5099]_ , \new_[5100]_ , \new_[5101]_ , \new_[5104]_ ,
    \new_[5107]_ , \new_[5108]_ , \new_[5111]_ , \new_[5115]_ ,
    \new_[5116]_ , \new_[5117]_ , \new_[5118]_ , \new_[5119]_ ,
    \new_[5120]_ , \new_[5123]_ , \new_[5126]_ , \new_[5127]_ ,
    \new_[5130]_ , \new_[5134]_ , \new_[5135]_ , \new_[5136]_ ,
    \new_[5137]_ , \new_[5140]_ , \new_[5143]_ , \new_[5144]_ ,
    \new_[5147]_ , \new_[5151]_ , \new_[5152]_ , \new_[5153]_ ,
    \new_[5154]_ , \new_[5155]_ , \new_[5158]_ , \new_[5161]_ ,
    \new_[5162]_ , \new_[5165]_ , \new_[5169]_ , \new_[5170]_ ,
    \new_[5171]_ , \new_[5172]_ , \new_[5175]_ , \new_[5178]_ ,
    \new_[5179]_ , \new_[5182]_ , \new_[5186]_ , \new_[5187]_ ,
    \new_[5188]_ , \new_[5189]_ , \new_[5190]_ , \new_[5191]_ ,
    \new_[5192]_ , \new_[5193]_ , \new_[5194]_ , \new_[5197]_ ,
    \new_[5200]_ , \new_[5201]_ , \new_[5204]_ , \new_[5208]_ ,
    \new_[5209]_ , \new_[5210]_ , \new_[5211]_ , \new_[5214]_ ,
    \new_[5217]_ , \new_[5218]_ , \new_[5221]_ , \new_[5225]_ ,
    \new_[5226]_ , \new_[5227]_ , \new_[5228]_ , \new_[5229]_ ,
    \new_[5232]_ , \new_[5235]_ , \new_[5236]_ , \new_[5239]_ ,
    \new_[5243]_ , \new_[5244]_ , \new_[5245]_ , \new_[5246]_ ,
    \new_[5249]_ , \new_[5252]_ , \new_[5253]_ , \new_[5256]_ ,
    \new_[5260]_ , \new_[5261]_ , \new_[5262]_ , \new_[5263]_ ,
    \new_[5264]_ , \new_[5265]_ , \new_[5268]_ , \new_[5271]_ ,
    \new_[5272]_ , \new_[5275]_ , \new_[5279]_ , \new_[5280]_ ,
    \new_[5281]_ , \new_[5282]_ , \new_[5285]_ , \new_[5288]_ ,
    \new_[5289]_ , \new_[5292]_ , \new_[5296]_ , \new_[5297]_ ,
    \new_[5298]_ , \new_[5299]_ , \new_[5300]_ , \new_[5303]_ ,
    \new_[5306]_ , \new_[5307]_ , \new_[5310]_ , \new_[5314]_ ,
    \new_[5315]_ , \new_[5316]_ , \new_[5317]_ , \new_[5320]_ ,
    \new_[5323]_ , \new_[5324]_ , \new_[5327]_ , \new_[5331]_ ,
    \new_[5332]_ , \new_[5333]_ , \new_[5334]_ , \new_[5335]_ ,
    \new_[5336]_ , \new_[5337]_ , \new_[5340]_ , \new_[5343]_ ,
    \new_[5344]_ , \new_[5347]_ , \new_[5351]_ , \new_[5352]_ ,
    \new_[5353]_ , \new_[5354]_ , \new_[5357]_ , \new_[5360]_ ,
    \new_[5361]_ , \new_[5364]_ , \new_[5368]_ , \new_[5369]_ ,
    \new_[5370]_ , \new_[5371]_ , \new_[5372]_ , \new_[5375]_ ,
    \new_[5378]_ , \new_[5379]_ , \new_[5382]_ , \new_[5386]_ ,
    \new_[5387]_ , \new_[5388]_ , \new_[5389]_ , \new_[5392]_ ,
    \new_[5395]_ , \new_[5396]_ , \new_[5399]_ , \new_[5403]_ ,
    \new_[5404]_ , \new_[5405]_ , \new_[5406]_ , \new_[5407]_ ,
    \new_[5408]_ , \new_[5411]_ , \new_[5414]_ , \new_[5415]_ ,
    \new_[5418]_ , \new_[5422]_ , \new_[5423]_ , \new_[5424]_ ,
    \new_[5425]_ , \new_[5428]_ , \new_[5431]_ , \new_[5432]_ ,
    \new_[5435]_ , \new_[5439]_ , \new_[5440]_ , \new_[5441]_ ,
    \new_[5442]_ , \new_[5443]_ , \new_[5446]_ , \new_[5449]_ ,
    \new_[5450]_ , \new_[5453]_ , \new_[5457]_ , \new_[5458]_ ,
    \new_[5459]_ , \new_[5460]_ , \new_[5463]_ , \new_[5466]_ ,
    \new_[5467]_ , \new_[5470]_ , \new_[5474]_ , \new_[5475]_ ,
    \new_[5476]_ , \new_[5477]_ , \new_[5478]_ , \new_[5479]_ ,
    \new_[5480]_ , \new_[5481]_ , \new_[5484]_ , \new_[5487]_ ,
    \new_[5488]_ , \new_[5491]_ , \new_[5495]_ , \new_[5496]_ ,
    \new_[5497]_ , \new_[5498]_ , \new_[5501]_ , \new_[5504]_ ,
    \new_[5505]_ , \new_[5508]_ , \new_[5512]_ , \new_[5513]_ ,
    \new_[5514]_ , \new_[5515]_ , \new_[5516]_ , \new_[5519]_ ,
    \new_[5522]_ , \new_[5523]_ , \new_[5526]_ , \new_[5530]_ ,
    \new_[5531]_ , \new_[5532]_ , \new_[5533]_ , \new_[5536]_ ,
    \new_[5539]_ , \new_[5540]_ , \new_[5543]_ , \new_[5547]_ ,
    \new_[5548]_ , \new_[5549]_ , \new_[5550]_ , \new_[5551]_ ,
    \new_[5552]_ , \new_[5555]_ , \new_[5558]_ , \new_[5559]_ ,
    \new_[5562]_ , \new_[5566]_ , \new_[5567]_ , \new_[5568]_ ,
    \new_[5569]_ , \new_[5572]_ , \new_[5575]_ , \new_[5576]_ ,
    \new_[5579]_ , \new_[5583]_ , \new_[5584]_ , \new_[5585]_ ,
    \new_[5586]_ , \new_[5587]_ , \new_[5590]_ , \new_[5593]_ ,
    \new_[5594]_ , \new_[5597]_ , \new_[5601]_ , \new_[5602]_ ,
    \new_[5603]_ , \new_[5604]_ , \new_[5607]_ , \new_[5610]_ ,
    \new_[5611]_ , \new_[5614]_ , \new_[5618]_ , \new_[5619]_ ,
    \new_[5620]_ , \new_[5621]_ , \new_[5622]_ , \new_[5623]_ ,
    \new_[5624]_ , \new_[5627]_ , \new_[5630]_ , \new_[5631]_ ,
    \new_[5634]_ , \new_[5638]_ , \new_[5639]_ , \new_[5640]_ ,
    \new_[5641]_ , \new_[5644]_ , \new_[5647]_ , \new_[5648]_ ,
    \new_[5651]_ , \new_[5655]_ , \new_[5656]_ , \new_[5657]_ ,
    \new_[5658]_ , \new_[5659]_ , \new_[5662]_ , \new_[5665]_ ,
    \new_[5666]_ , \new_[5669]_ , \new_[5673]_ , \new_[5674]_ ,
    \new_[5675]_ , \new_[5676]_ , \new_[5679]_ , \new_[5682]_ ,
    \new_[5683]_ , \new_[5686]_ , \new_[5690]_ , \new_[5691]_ ,
    \new_[5692]_ , \new_[5693]_ , \new_[5694]_ , \new_[5695]_ ,
    \new_[5698]_ , \new_[5701]_ , \new_[5702]_ , \new_[5705]_ ,
    \new_[5709]_ , \new_[5710]_ , \new_[5711]_ , \new_[5712]_ ,
    \new_[5715]_ , \new_[5718]_ , \new_[5719]_ , \new_[5722]_ ,
    \new_[5726]_ , \new_[5727]_ , \new_[5728]_ , \new_[5729]_ ,
    \new_[5730]_ , \new_[5733]_ , \new_[5736]_ , \new_[5737]_ ,
    \new_[5740]_ , \new_[5744]_ , \new_[5745]_ , \new_[5746]_ ,
    \new_[5747]_ , \new_[5750]_ , \new_[5754]_ , \new_[5755]_ ,
    \new_[5756]_ , \new_[5759]_ , \new_[5763]_ , \new_[5764]_ ,
    \new_[5765]_ , \new_[5766]_ , \new_[5767]_ , \new_[5768]_ ,
    \new_[5769]_ , \new_[5770]_ , \new_[5771]_ , \new_[5772]_ ,
    \new_[5775]_ , \new_[5778]_ , \new_[5779]_ , \new_[5782]_ ,
    \new_[5786]_ , \new_[5787]_ , \new_[5788]_ , \new_[5789]_ ,
    \new_[5792]_ , \new_[5795]_ , \new_[5796]_ , \new_[5799]_ ,
    \new_[5803]_ , \new_[5804]_ , \new_[5805]_ , \new_[5806]_ ,
    \new_[5807]_ , \new_[5810]_ , \new_[5813]_ , \new_[5814]_ ,
    \new_[5817]_ , \new_[5821]_ , \new_[5822]_ , \new_[5823]_ ,
    \new_[5824]_ , \new_[5827]_ , \new_[5830]_ , \new_[5831]_ ,
    \new_[5834]_ , \new_[5838]_ , \new_[5839]_ , \new_[5840]_ ,
    \new_[5841]_ , \new_[5842]_ , \new_[5843]_ , \new_[5846]_ ,
    \new_[5849]_ , \new_[5850]_ , \new_[5853]_ , \new_[5857]_ ,
    \new_[5858]_ , \new_[5859]_ , \new_[5860]_ , \new_[5863]_ ,
    \new_[5866]_ , \new_[5867]_ , \new_[5870]_ , \new_[5874]_ ,
    \new_[5875]_ , \new_[5876]_ , \new_[5877]_ , \new_[5878]_ ,
    \new_[5881]_ , \new_[5884]_ , \new_[5885]_ , \new_[5888]_ ,
    \new_[5892]_ , \new_[5893]_ , \new_[5894]_ , \new_[5895]_ ,
    \new_[5898]_ , \new_[5901]_ , \new_[5902]_ , \new_[5905]_ ,
    \new_[5909]_ , \new_[5910]_ , \new_[5911]_ , \new_[5912]_ ,
    \new_[5913]_ , \new_[5914]_ , \new_[5915]_ , \new_[5918]_ ,
    \new_[5921]_ , \new_[5922]_ , \new_[5925]_ , \new_[5929]_ ,
    \new_[5930]_ , \new_[5931]_ , \new_[5932]_ , \new_[5935]_ ,
    \new_[5938]_ , \new_[5939]_ , \new_[5942]_ , \new_[5946]_ ,
    \new_[5947]_ , \new_[5948]_ , \new_[5949]_ , \new_[5950]_ ,
    \new_[5953]_ , \new_[5956]_ , \new_[5957]_ , \new_[5960]_ ,
    \new_[5964]_ , \new_[5965]_ , \new_[5966]_ , \new_[5967]_ ,
    \new_[5970]_ , \new_[5973]_ , \new_[5974]_ , \new_[5977]_ ,
    \new_[5981]_ , \new_[5982]_ , \new_[5983]_ , \new_[5984]_ ,
    \new_[5985]_ , \new_[5986]_ , \new_[5989]_ , \new_[5992]_ ,
    \new_[5993]_ , \new_[5996]_ , \new_[6000]_ , \new_[6001]_ ,
    \new_[6002]_ , \new_[6003]_ , \new_[6006]_ , \new_[6009]_ ,
    \new_[6010]_ , \new_[6013]_ , \new_[6017]_ , \new_[6018]_ ,
    \new_[6019]_ , \new_[6020]_ , \new_[6021]_ , \new_[6024]_ ,
    \new_[6027]_ , \new_[6028]_ , \new_[6031]_ , \new_[6035]_ ,
    \new_[6036]_ , \new_[6037]_ , \new_[6038]_ , \new_[6041]_ ,
    \new_[6044]_ , \new_[6045]_ , \new_[6048]_ , \new_[6052]_ ,
    \new_[6053]_ , \new_[6054]_ , \new_[6055]_ , \new_[6056]_ ,
    \new_[6057]_ , \new_[6058]_ , \new_[6059]_ , \new_[6062]_ ,
    \new_[6065]_ , \new_[6066]_ , \new_[6069]_ , \new_[6073]_ ,
    \new_[6074]_ , \new_[6075]_ , \new_[6076]_ , \new_[6079]_ ,
    \new_[6082]_ , \new_[6083]_ , \new_[6086]_ , \new_[6090]_ ,
    \new_[6091]_ , \new_[6092]_ , \new_[6093]_ , \new_[6094]_ ,
    \new_[6097]_ , \new_[6100]_ , \new_[6101]_ , \new_[6104]_ ,
    \new_[6108]_ , \new_[6109]_ , \new_[6110]_ , \new_[6111]_ ,
    \new_[6114]_ , \new_[6117]_ , \new_[6118]_ , \new_[6121]_ ,
    \new_[6125]_ , \new_[6126]_ , \new_[6127]_ , \new_[6128]_ ,
    \new_[6129]_ , \new_[6130]_ , \new_[6133]_ , \new_[6136]_ ,
    \new_[6137]_ , \new_[6140]_ , \new_[6144]_ , \new_[6145]_ ,
    \new_[6146]_ , \new_[6147]_ , \new_[6150]_ , \new_[6153]_ ,
    \new_[6154]_ , \new_[6157]_ , \new_[6161]_ , \new_[6162]_ ,
    \new_[6163]_ , \new_[6164]_ , \new_[6165]_ , \new_[6168]_ ,
    \new_[6171]_ , \new_[6172]_ , \new_[6175]_ , \new_[6179]_ ,
    \new_[6180]_ , \new_[6181]_ , \new_[6182]_ , \new_[6185]_ ,
    \new_[6188]_ , \new_[6189]_ , \new_[6192]_ , \new_[6196]_ ,
    \new_[6197]_ , \new_[6198]_ , \new_[6199]_ , \new_[6200]_ ,
    \new_[6201]_ , \new_[6202]_ , \new_[6205]_ , \new_[6208]_ ,
    \new_[6209]_ , \new_[6212]_ , \new_[6216]_ , \new_[6217]_ ,
    \new_[6218]_ , \new_[6219]_ , \new_[6222]_ , \new_[6225]_ ,
    \new_[6226]_ , \new_[6229]_ , \new_[6233]_ , \new_[6234]_ ,
    \new_[6235]_ , \new_[6236]_ , \new_[6237]_ , \new_[6240]_ ,
    \new_[6243]_ , \new_[6244]_ , \new_[6247]_ , \new_[6251]_ ,
    \new_[6252]_ , \new_[6253]_ , \new_[6254]_ , \new_[6257]_ ,
    \new_[6260]_ , \new_[6261]_ , \new_[6264]_ , \new_[6268]_ ,
    \new_[6269]_ , \new_[6270]_ , \new_[6271]_ , \new_[6272]_ ,
    \new_[6273]_ , \new_[6276]_ , \new_[6279]_ , \new_[6280]_ ,
    \new_[6283]_ , \new_[6287]_ , \new_[6288]_ , \new_[6289]_ ,
    \new_[6290]_ , \new_[6293]_ , \new_[6296]_ , \new_[6297]_ ,
    \new_[6300]_ , \new_[6304]_ , \new_[6305]_ , \new_[6306]_ ,
    \new_[6307]_ , \new_[6308]_ , \new_[6311]_ , \new_[6314]_ ,
    \new_[6315]_ , \new_[6318]_ , \new_[6322]_ , \new_[6323]_ ,
    \new_[6324]_ , \new_[6325]_ , \new_[6328]_ , \new_[6332]_ ,
    \new_[6333]_ , \new_[6334]_ , \new_[6337]_ , \new_[6341]_ ,
    \new_[6342]_ , \new_[6343]_ , \new_[6344]_ , \new_[6345]_ ,
    \new_[6346]_ , \new_[6347]_ , \new_[6348]_ , \new_[6349]_ ,
    \new_[6352]_ , \new_[6355]_ , \new_[6356]_ , \new_[6359]_ ,
    \new_[6363]_ , \new_[6364]_ , \new_[6365]_ , \new_[6366]_ ,
    \new_[6369]_ , \new_[6372]_ , \new_[6373]_ , \new_[6376]_ ,
    \new_[6380]_ , \new_[6381]_ , \new_[6382]_ , \new_[6383]_ ,
    \new_[6384]_ , \new_[6387]_ , \new_[6390]_ , \new_[6391]_ ,
    \new_[6394]_ , \new_[6398]_ , \new_[6399]_ , \new_[6400]_ ,
    \new_[6401]_ , \new_[6404]_ , \new_[6407]_ , \new_[6408]_ ,
    \new_[6411]_ , \new_[6415]_ , \new_[6416]_ , \new_[6417]_ ,
    \new_[6418]_ , \new_[6419]_ , \new_[6420]_ , \new_[6423]_ ,
    \new_[6426]_ , \new_[6427]_ , \new_[6430]_ , \new_[6434]_ ,
    \new_[6435]_ , \new_[6436]_ , \new_[6437]_ , \new_[6440]_ ,
    \new_[6443]_ , \new_[6444]_ , \new_[6447]_ , \new_[6451]_ ,
    \new_[6452]_ , \new_[6453]_ , \new_[6454]_ , \new_[6455]_ ,
    \new_[6458]_ , \new_[6461]_ , \new_[6462]_ , \new_[6465]_ ,
    \new_[6469]_ , \new_[6470]_ , \new_[6471]_ , \new_[6472]_ ,
    \new_[6475]_ , \new_[6478]_ , \new_[6479]_ , \new_[6482]_ ,
    \new_[6486]_ , \new_[6487]_ , \new_[6488]_ , \new_[6489]_ ,
    \new_[6490]_ , \new_[6491]_ , \new_[6492]_ , \new_[6495]_ ,
    \new_[6498]_ , \new_[6499]_ , \new_[6502]_ , \new_[6506]_ ,
    \new_[6507]_ , \new_[6508]_ , \new_[6509]_ , \new_[6512]_ ,
    \new_[6515]_ , \new_[6516]_ , \new_[6519]_ , \new_[6523]_ ,
    \new_[6524]_ , \new_[6525]_ , \new_[6526]_ , \new_[6527]_ ,
    \new_[6530]_ , \new_[6533]_ , \new_[6534]_ , \new_[6537]_ ,
    \new_[6541]_ , \new_[6542]_ , \new_[6543]_ , \new_[6544]_ ,
    \new_[6547]_ , \new_[6550]_ , \new_[6551]_ , \new_[6554]_ ,
    \new_[6558]_ , \new_[6559]_ , \new_[6560]_ , \new_[6561]_ ,
    \new_[6562]_ , \new_[6563]_ , \new_[6566]_ , \new_[6569]_ ,
    \new_[6570]_ , \new_[6573]_ , \new_[6577]_ , \new_[6578]_ ,
    \new_[6579]_ , \new_[6580]_ , \new_[6583]_ , \new_[6586]_ ,
    \new_[6587]_ , \new_[6590]_ , \new_[6594]_ , \new_[6595]_ ,
    \new_[6596]_ , \new_[6597]_ , \new_[6598]_ , \new_[6601]_ ,
    \new_[6604]_ , \new_[6605]_ , \new_[6608]_ , \new_[6612]_ ,
    \new_[6613]_ , \new_[6614]_ , \new_[6615]_ , \new_[6618]_ ,
    \new_[6621]_ , \new_[6622]_ , \new_[6625]_ , \new_[6629]_ ,
    \new_[6630]_ , \new_[6631]_ , \new_[6632]_ , \new_[6633]_ ,
    \new_[6634]_ , \new_[6635]_ , \new_[6636]_ , \new_[6639]_ ,
    \new_[6642]_ , \new_[6643]_ , \new_[6646]_ , \new_[6650]_ ,
    \new_[6651]_ , \new_[6652]_ , \new_[6653]_ , \new_[6656]_ ,
    \new_[6659]_ , \new_[6660]_ , \new_[6663]_ , \new_[6667]_ ,
    \new_[6668]_ , \new_[6669]_ , \new_[6670]_ , \new_[6671]_ ,
    \new_[6674]_ , \new_[6677]_ , \new_[6678]_ , \new_[6681]_ ,
    \new_[6685]_ , \new_[6686]_ , \new_[6687]_ , \new_[6688]_ ,
    \new_[6691]_ , \new_[6694]_ , \new_[6695]_ , \new_[6698]_ ,
    \new_[6702]_ , \new_[6703]_ , \new_[6704]_ , \new_[6705]_ ,
    \new_[6706]_ , \new_[6707]_ , \new_[6710]_ , \new_[6713]_ ,
    \new_[6714]_ , \new_[6717]_ , \new_[6721]_ , \new_[6722]_ ,
    \new_[6723]_ , \new_[6724]_ , \new_[6727]_ , \new_[6730]_ ,
    \new_[6731]_ , \new_[6734]_ , \new_[6738]_ , \new_[6739]_ ,
    \new_[6740]_ , \new_[6741]_ , \new_[6742]_ , \new_[6745]_ ,
    \new_[6748]_ , \new_[6749]_ , \new_[6752]_ , \new_[6756]_ ,
    \new_[6757]_ , \new_[6758]_ , \new_[6759]_ , \new_[6762]_ ,
    \new_[6765]_ , \new_[6766]_ , \new_[6769]_ , \new_[6773]_ ,
    \new_[6774]_ , \new_[6775]_ , \new_[6776]_ , \new_[6777]_ ,
    \new_[6778]_ , \new_[6779]_ , \new_[6782]_ , \new_[6785]_ ,
    \new_[6786]_ , \new_[6789]_ , \new_[6793]_ , \new_[6794]_ ,
    \new_[6795]_ , \new_[6796]_ , \new_[6799]_ , \new_[6802]_ ,
    \new_[6803]_ , \new_[6806]_ , \new_[6810]_ , \new_[6811]_ ,
    \new_[6812]_ , \new_[6813]_ , \new_[6814]_ , \new_[6817]_ ,
    \new_[6820]_ , \new_[6821]_ , \new_[6824]_ , \new_[6828]_ ,
    \new_[6829]_ , \new_[6830]_ , \new_[6831]_ , \new_[6834]_ ,
    \new_[6837]_ , \new_[6838]_ , \new_[6841]_ , \new_[6845]_ ,
    \new_[6846]_ , \new_[6847]_ , \new_[6848]_ , \new_[6849]_ ,
    \new_[6850]_ , \new_[6853]_ , \new_[6856]_ , \new_[6857]_ ,
    \new_[6860]_ , \new_[6864]_ , \new_[6865]_ , \new_[6866]_ ,
    \new_[6867]_ , \new_[6870]_ , \new_[6873]_ , \new_[6874]_ ,
    \new_[6877]_ , \new_[6881]_ , \new_[6882]_ , \new_[6883]_ ,
    \new_[6884]_ , \new_[6885]_ , \new_[6888]_ , \new_[6891]_ ,
    \new_[6892]_ , \new_[6895]_ , \new_[6899]_ , \new_[6900]_ ,
    \new_[6901]_ , \new_[6902]_ , \new_[6905]_ , \new_[6909]_ ,
    \new_[6910]_ , \new_[6911]_ , \new_[6914]_ , \new_[6918]_ ,
    \new_[6919]_ , \new_[6920]_ , \new_[6921]_ , \new_[6922]_ ,
    \new_[6923]_ , \new_[6924]_ , \new_[6925]_ , \new_[6926]_ ,
    \new_[6927]_ , \new_[6928]_ , \new_[6932]_ , \new_[6933]_ ,
    \new_[6937]_ , \new_[6938]_ , \new_[6942]_ , \new_[6943]_ ,
    \new_[6947]_ , \new_[6948]_ , \new_[6952]_ , \new_[6953]_ ,
    \new_[6957]_ , \new_[6958]_ , \new_[6962]_ , \new_[6963]_ ,
    \new_[6967]_ , \new_[6968]_ , \new_[6972]_ , \new_[6973]_ ,
    \new_[6977]_ , \new_[6978]_ , \new_[6982]_ , \new_[6983]_ ,
    \new_[6987]_ , \new_[6988]_ , \new_[6992]_ , \new_[6993]_ ,
    \new_[6997]_ , \new_[6998]_ , \new_[7002]_ , \new_[7003]_ ,
    \new_[7007]_ , \new_[7008]_ , \new_[7012]_ , \new_[7013]_ ,
    \new_[7016]_ , \new_[7019]_ , \new_[7020]_ , \new_[7024]_ ,
    \new_[7025]_ , \new_[7028]_ , \new_[7031]_ , \new_[7032]_ ,
    \new_[7036]_ , \new_[7037]_ , \new_[7040]_ , \new_[7043]_ ,
    \new_[7044]_ , \new_[7048]_ , \new_[7049]_ , \new_[7052]_ ,
    \new_[7055]_ , \new_[7056]_ , \new_[7060]_ , \new_[7061]_ ,
    \new_[7064]_ , \new_[7067]_ , \new_[7068]_ , \new_[7072]_ ,
    \new_[7073]_ , \new_[7076]_ , \new_[7079]_ , \new_[7080]_ ,
    \new_[7084]_ , \new_[7085]_ , \new_[7088]_ , \new_[7091]_ ,
    \new_[7092]_ , \new_[7096]_ , \new_[7097]_ , \new_[7100]_ ,
    \new_[7103]_ , \new_[7104]_ , \new_[7108]_ , \new_[7109]_ ,
    \new_[7112]_ , \new_[7115]_ , \new_[7116]_ , \new_[7120]_ ,
    \new_[7121]_ , \new_[7124]_ , \new_[7127]_ , \new_[7128]_ ,
    \new_[7132]_ , \new_[7133]_ , \new_[7136]_ , \new_[7139]_ ,
    \new_[7140]_ , \new_[7144]_ , \new_[7145]_ , \new_[7148]_ ,
    \new_[7151]_ , \new_[7152]_ , \new_[7156]_ , \new_[7157]_ ,
    \new_[7160]_ , \new_[7163]_ , \new_[7164]_ , \new_[7168]_ ,
    \new_[7169]_ , \new_[7172]_ , \new_[7175]_ , \new_[7176]_ ,
    \new_[7180]_ , \new_[7181]_ , \new_[7184]_ , \new_[7187]_ ,
    \new_[7188]_ , \new_[7192]_ , \new_[7193]_ , \new_[7196]_ ,
    \new_[7199]_ , \new_[7200]_ , \new_[7204]_ , \new_[7205]_ ,
    \new_[7208]_ , \new_[7211]_ , \new_[7212]_ , \new_[7216]_ ,
    \new_[7217]_ , \new_[7220]_ , \new_[7223]_ , \new_[7224]_ ,
    \new_[7228]_ , \new_[7229]_ , \new_[7232]_ , \new_[7235]_ ,
    \new_[7236]_ , \new_[7240]_ , \new_[7241]_ , \new_[7244]_ ,
    \new_[7247]_ , \new_[7248]_ , \new_[7252]_ , \new_[7253]_ ,
    \new_[7256]_ , \new_[7259]_ , \new_[7260]_ , \new_[7264]_ ,
    \new_[7265]_ , \new_[7268]_ , \new_[7271]_ , \new_[7272]_ ,
    \new_[7276]_ , \new_[7277]_ , \new_[7280]_ , \new_[7283]_ ,
    \new_[7284]_ , \new_[7288]_ , \new_[7289]_ , \new_[7292]_ ,
    \new_[7295]_ , \new_[7296]_ , \new_[7300]_ , \new_[7301]_ ,
    \new_[7304]_ , \new_[7307]_ , \new_[7308]_ , \new_[7312]_ ,
    \new_[7313]_ , \new_[7316]_ , \new_[7319]_ , \new_[7320]_ ,
    \new_[7324]_ , \new_[7325]_ , \new_[7328]_ , \new_[7331]_ ,
    \new_[7332]_ , \new_[7336]_ , \new_[7337]_ , \new_[7340]_ ,
    \new_[7343]_ , \new_[7344]_ , \new_[7348]_ , \new_[7349]_ ,
    \new_[7352]_ , \new_[7355]_ , \new_[7356]_ , \new_[7360]_ ,
    \new_[7361]_ , \new_[7364]_ , \new_[7367]_ , \new_[7368]_ ,
    \new_[7372]_ , \new_[7373]_ , \new_[7376]_ , \new_[7379]_ ,
    \new_[7380]_ , \new_[7384]_ , \new_[7385]_ , \new_[7388]_ ,
    \new_[7391]_ , \new_[7392]_ , \new_[7396]_ , \new_[7397]_ ,
    \new_[7400]_ , \new_[7403]_ , \new_[7404]_ , \new_[7408]_ ,
    \new_[7409]_ , \new_[7412]_ , \new_[7415]_ , \new_[7416]_ ,
    \new_[7420]_ , \new_[7421]_ , \new_[7424]_ , \new_[7427]_ ,
    \new_[7428]_ , \new_[7432]_ , \new_[7433]_ , \new_[7436]_ ,
    \new_[7439]_ , \new_[7440]_ , \new_[7444]_ , \new_[7445]_ ,
    \new_[7448]_ , \new_[7451]_ , \new_[7452]_ , \new_[7456]_ ,
    \new_[7457]_ , \new_[7460]_ , \new_[7463]_ , \new_[7464]_ ,
    \new_[7468]_ , \new_[7469]_ , \new_[7472]_ , \new_[7475]_ ,
    \new_[7476]_ , \new_[7480]_ , \new_[7481]_ , \new_[7484]_ ,
    \new_[7487]_ , \new_[7488]_ , \new_[7492]_ , \new_[7493]_ ,
    \new_[7496]_ , \new_[7499]_ , \new_[7500]_ , \new_[7504]_ ,
    \new_[7505]_ , \new_[7508]_ , \new_[7511]_ , \new_[7512]_ ,
    \new_[7516]_ , \new_[7517]_ , \new_[7520]_ , \new_[7523]_ ,
    \new_[7524]_ , \new_[7528]_ , \new_[7529]_ , \new_[7532]_ ,
    \new_[7535]_ , \new_[7536]_ , \new_[7540]_ , \new_[7541]_ ,
    \new_[7544]_ , \new_[7547]_ , \new_[7548]_ , \new_[7552]_ ,
    \new_[7553]_ , \new_[7556]_ , \new_[7559]_ , \new_[7560]_ ,
    \new_[7564]_ , \new_[7565]_ , \new_[7568]_ , \new_[7571]_ ,
    \new_[7572]_ , \new_[7576]_ , \new_[7577]_ , \new_[7580]_ ,
    \new_[7583]_ , \new_[7584]_ , \new_[7588]_ , \new_[7589]_ ,
    \new_[7592]_ , \new_[7595]_ , \new_[7596]_ , \new_[7600]_ ,
    \new_[7601]_ , \new_[7604]_ , \new_[7607]_ , \new_[7608]_ ,
    \new_[7612]_ , \new_[7613]_ , \new_[7616]_ , \new_[7619]_ ,
    \new_[7620]_ , \new_[7624]_ , \new_[7625]_ , \new_[7628]_ ,
    \new_[7631]_ , \new_[7632]_ , \new_[7635]_ , \new_[7638]_ ,
    \new_[7639]_ , \new_[7642]_ , \new_[7645]_ , \new_[7646]_ ,
    \new_[7649]_ , \new_[7652]_ , \new_[7653]_ , \new_[7656]_ ,
    \new_[7659]_ , \new_[7660]_ , \new_[7663]_ , \new_[7666]_ ,
    \new_[7667]_ , \new_[7670]_ , \new_[7673]_ , \new_[7674]_ ,
    \new_[7677]_ , \new_[7680]_ , \new_[7681]_ , \new_[7684]_ ,
    \new_[7687]_ , \new_[7688]_ , \new_[7691]_ , \new_[7694]_ ,
    \new_[7695]_ , \new_[7698]_ , \new_[7701]_ , \new_[7702]_ ,
    \new_[7705]_ , \new_[7708]_ , \new_[7709]_ , \new_[7712]_ ,
    \new_[7715]_ , \new_[7716]_ , \new_[7719]_ , \new_[7722]_ ,
    \new_[7723]_ , \new_[7726]_ , \new_[7729]_ , \new_[7730]_ ,
    \new_[7733]_ , \new_[7736]_ , \new_[7737]_ , \new_[7740]_ ,
    \new_[7743]_ , \new_[7744]_ , \new_[7747]_ , \new_[7750]_ ,
    \new_[7751]_ , \new_[7754]_ , \new_[7757]_ , \new_[7758]_ ,
    \new_[7761]_ , \new_[7764]_ , \new_[7765]_ , \new_[7768]_ ,
    \new_[7771]_ , \new_[7772]_ , \new_[7775]_ , \new_[7778]_ ,
    \new_[7779]_ , \new_[7782]_ , \new_[7785]_ , \new_[7786]_ ,
    \new_[7789]_ , \new_[7792]_ , \new_[7793]_ , \new_[7796]_ ,
    \new_[7799]_ , \new_[7800]_ , \new_[7803]_ , \new_[7806]_ ,
    \new_[7807]_ , \new_[7810]_ , \new_[7813]_ , \new_[7814]_ ,
    \new_[7817]_ , \new_[7820]_ , \new_[7821]_ , \new_[7824]_ ,
    \new_[7827]_ , \new_[7828]_ , \new_[7831]_ , \new_[7834]_ ,
    \new_[7835]_ , \new_[7838]_ , \new_[7841]_ , \new_[7842]_ ,
    \new_[7845]_ , \new_[7848]_ , \new_[7849]_ , \new_[7852]_ ,
    \new_[7855]_ , \new_[7856]_ , \new_[7859]_ , \new_[7862]_ ,
    \new_[7863]_ , \new_[7866]_ , \new_[7869]_ , \new_[7870]_ ,
    \new_[7873]_ , \new_[7876]_ , \new_[7877]_ , \new_[7880]_ ,
    \new_[7883]_ , \new_[7884]_ , \new_[7887]_ , \new_[7890]_ ,
    \new_[7891]_ , \new_[7894]_ , \new_[7897]_ , \new_[7898]_ ,
    \new_[7901]_ , \new_[7904]_ , \new_[7905]_ , \new_[7908]_ ,
    \new_[7911]_ , \new_[7912]_ , \new_[7915]_ , \new_[7918]_ ,
    \new_[7919]_ , \new_[7922]_ , \new_[7925]_ , \new_[7926]_ ,
    \new_[7929]_ , \new_[7932]_ , \new_[7933]_ , \new_[7936]_ ,
    \new_[7939]_ , \new_[7940]_ , \new_[7943]_ , \new_[7946]_ ,
    \new_[7947]_ , \new_[7950]_ , \new_[7953]_ , \new_[7954]_ ,
    \new_[7957]_ , \new_[7960]_ , \new_[7961]_ , \new_[7964]_ ,
    \new_[7967]_ , \new_[7968]_ , \new_[7971]_ , \new_[7974]_ ,
    \new_[7975]_ , \new_[7978]_ , \new_[7981]_ , \new_[7982]_ ,
    \new_[7985]_ , \new_[7988]_ , \new_[7989]_ , \new_[7992]_ ,
    \new_[7995]_ , \new_[7996]_ , \new_[7999]_ , \new_[8002]_ ,
    \new_[8003]_ , \new_[8006]_ , \new_[8009]_ , \new_[8010]_ ,
    \new_[8013]_ , \new_[8016]_ , \new_[8017]_ , \new_[8020]_ ,
    \new_[8023]_ , \new_[8024]_ , \new_[8027]_ , \new_[8030]_ ,
    \new_[8031]_ , \new_[8034]_ , \new_[8037]_ , \new_[8038]_ ,
    \new_[8041]_ , \new_[8044]_ , \new_[8045]_ , \new_[8048]_ ,
    \new_[8051]_ , \new_[8052]_ , \new_[8055]_ , \new_[8058]_ ,
    \new_[8059]_ , \new_[8062]_ , \new_[8065]_ , \new_[8066]_ ,
    \new_[8069]_ , \new_[8072]_ , \new_[8073]_ , \new_[8076]_ ,
    \new_[8079]_ , \new_[8080]_ , \new_[8083]_ , \new_[8086]_ ,
    \new_[8087]_ , \new_[8090]_ , \new_[8093]_ , \new_[8094]_ ,
    \new_[8097]_ , \new_[8100]_ , \new_[8101]_ , \new_[8104]_ ,
    \new_[8107]_ , \new_[8108]_ , \new_[8111]_ , \new_[8114]_ ,
    \new_[8115]_ , \new_[8118]_ , \new_[8121]_ , \new_[8122]_ ,
    \new_[8125]_ , \new_[8128]_ , \new_[8129]_ , \new_[8132]_ ,
    \new_[8135]_ , \new_[8136]_ , \new_[8139]_ , \new_[8142]_ ,
    \new_[8143]_ , \new_[8146]_ , \new_[8149]_ , \new_[8150]_ ,
    \new_[8153]_ , \new_[8156]_ , \new_[8157]_ , \new_[8160]_ ,
    \new_[8163]_ , \new_[8164]_ , \new_[8167]_ , \new_[8170]_ ,
    \new_[8171]_ , \new_[8174]_ , \new_[8177]_ , \new_[8178]_ ,
    \new_[8181]_ , \new_[8184]_ , \new_[8185]_ , \new_[8188]_ ,
    \new_[8191]_ , \new_[8192]_ , \new_[8195]_ , \new_[8198]_ ,
    \new_[8199]_ , \new_[8202]_ , \new_[8205]_ , \new_[8206]_ ,
    \new_[8209]_ , \new_[8212]_ , \new_[8213]_ , \new_[8216]_ ,
    \new_[8219]_ , \new_[8220]_ , \new_[8223]_ , \new_[8226]_ ,
    \new_[8227]_ , \new_[8230]_ , \new_[8233]_ , \new_[8234]_ ,
    \new_[8237]_ , \new_[8240]_ , \new_[8241]_ , \new_[8244]_ ,
    \new_[8247]_ , \new_[8248]_ , \new_[8251]_ , \new_[8254]_ ,
    \new_[8255]_ , \new_[8258]_ , \new_[8261]_ , \new_[8262]_ ,
    \new_[8265]_ , \new_[8268]_ , \new_[8269]_ , \new_[8272]_ ,
    \new_[8275]_ , \new_[8276]_ , \new_[8279]_ , \new_[8282]_ ,
    \new_[8283]_ , \new_[8286]_ , \new_[8289]_ , \new_[8290]_ ,
    \new_[8293]_ , \new_[8296]_ , \new_[8297]_ , \new_[8300]_ ,
    \new_[8303]_ , \new_[8304]_ , \new_[8307]_ , \new_[8310]_ ,
    \new_[8311]_ , \new_[8314]_ , \new_[8317]_ , \new_[8318]_ ,
    \new_[8321]_ , \new_[8324]_ , \new_[8325]_ , \new_[8328]_ ,
    \new_[8331]_ , \new_[8332]_ , \new_[8335]_ , \new_[8338]_ ,
    \new_[8339]_ , \new_[8342]_ , \new_[8345]_ , \new_[8346]_ ,
    \new_[8349]_ , \new_[8352]_ , \new_[8353]_ , \new_[8356]_ ,
    \new_[8359]_ , \new_[8360]_ , \new_[8363]_ , \new_[8366]_ ,
    \new_[8367]_ , \new_[8370]_ , \new_[8373]_ , \new_[8374]_ ,
    \new_[8377]_ , \new_[8380]_ , \new_[8381]_ , \new_[8384]_ ,
    \new_[8387]_ , \new_[8388]_ , \new_[8391]_ , \new_[8394]_ ,
    \new_[8395]_ , \new_[8398]_ , \new_[8401]_ , \new_[8402]_ ,
    \new_[8405]_ , \new_[8408]_ , \new_[8409]_ , \new_[8412]_ ,
    \new_[8415]_ , \new_[8416]_ , \new_[8419]_ , \new_[8422]_ ,
    \new_[8423]_ , \new_[8426]_ , \new_[8429]_ , \new_[8430]_ ,
    \new_[8433]_ , \new_[8436]_ , \new_[8437]_ , \new_[8440]_ ,
    \new_[8443]_ , \new_[8444]_ , \new_[8447]_ , \new_[8450]_ ,
    \new_[8451]_ , \new_[8454]_ , \new_[8457]_ , \new_[8458]_ ,
    \new_[8461]_ , \new_[8464]_ , \new_[8465]_ , \new_[8468]_ ,
    \new_[8471]_ , \new_[8472]_ , \new_[8475]_ , \new_[8478]_ ,
    \new_[8479]_ , \new_[8482]_ , \new_[8485]_ , \new_[8486]_ ,
    \new_[8489]_ , \new_[8492]_ , \new_[8493]_ , \new_[8496]_ ,
    \new_[8499]_ , \new_[8500]_ , \new_[8503]_ , \new_[8506]_ ,
    \new_[8507]_ , \new_[8510]_ , \new_[8513]_ , \new_[8514]_ ,
    \new_[8517]_ , \new_[8520]_ , \new_[8521]_ , \new_[8524]_ ,
    \new_[8527]_ , \new_[8528]_ , \new_[8531]_ , \new_[8534]_ ,
    \new_[8535]_ , \new_[8538]_ , \new_[8541]_ , \new_[8542]_ ,
    \new_[8545]_ , \new_[8548]_ , \new_[8549]_ , \new_[8552]_ ,
    \new_[8555]_ , \new_[8556]_ , \new_[8559]_ , \new_[8562]_ ,
    \new_[8563]_ , \new_[8566]_ , \new_[8569]_ , \new_[8570]_ ,
    \new_[8573]_ , \new_[8576]_ , \new_[8577]_ , \new_[8580]_ ,
    \new_[8583]_ , \new_[8584]_ , \new_[8587]_ , \new_[8590]_ ,
    \new_[8591]_ , \new_[8594]_ , \new_[8597]_ , \new_[8598]_ ,
    \new_[8601]_ , \new_[8604]_ , \new_[8605]_ , \new_[8608]_ ,
    \new_[8611]_ , \new_[8612]_ , \new_[8615]_ , \new_[8618]_ ,
    \new_[8619]_ , \new_[8622]_ , \new_[8625]_ , \new_[8626]_ ,
    \new_[8629]_ , \new_[8632]_ , \new_[8633]_ , \new_[8636]_ ,
    \new_[8639]_ , \new_[8640]_ , \new_[8643]_ , \new_[8646]_ ,
    \new_[8647]_ , \new_[8650]_ , \new_[8653]_ , \new_[8654]_ ,
    \new_[8657]_ , \new_[8660]_ , \new_[8661]_ , \new_[8664]_ ,
    \new_[8667]_ , \new_[8668]_ , \new_[8671]_ , \new_[8674]_ ,
    \new_[8675]_ , \new_[8678]_ , \new_[8681]_ , \new_[8682]_ ,
    \new_[8685]_ , \new_[8688]_ , \new_[8689]_ , \new_[8692]_ ,
    \new_[8695]_ , \new_[8696]_ , \new_[8699]_ , \new_[8702]_ ,
    \new_[8703]_ , \new_[8706]_ , \new_[8709]_ , \new_[8710]_ ,
    \new_[8713]_ , \new_[8716]_ , \new_[8717]_ , \new_[8720]_ ,
    \new_[8723]_ , \new_[8724]_ , \new_[8727]_ , \new_[8730]_ ,
    \new_[8731]_ , \new_[8734]_ , \new_[8737]_ , \new_[8738]_ ,
    \new_[8741]_ , \new_[8744]_ , \new_[8745]_ , \new_[8748]_ ,
    \new_[8751]_ , \new_[8752]_ , \new_[8755]_ , \new_[8758]_ ,
    \new_[8759]_ , \new_[8762]_ , \new_[8765]_ , \new_[8766]_ ,
    \new_[8769]_ , \new_[8772]_ , \new_[8773]_ , \new_[8776]_ ,
    \new_[8779]_ , \new_[8780]_ , \new_[8783]_ , \new_[8786]_ ,
    \new_[8787]_ , \new_[8790]_ , \new_[8793]_ , \new_[8794]_ ,
    \new_[8797]_ , \new_[8800]_ , \new_[8801]_ , \new_[8804]_ ,
    \new_[8807]_ , \new_[8808]_ , \new_[8811]_ , \new_[8814]_ ,
    \new_[8815]_ , \new_[8818]_ , \new_[8821]_ , \new_[8822]_ ,
    \new_[8825]_ , \new_[8828]_ , \new_[8829]_ , \new_[8832]_ ,
    \new_[8835]_ , \new_[8836]_ , \new_[8839]_ , \new_[8842]_ ,
    \new_[8843]_ , \new_[8846]_ , \new_[8849]_ , \new_[8850]_ ,
    \new_[8853]_ , \new_[8856]_ , \new_[8857]_ , \new_[8860]_ ,
    \new_[8863]_ , \new_[8864]_ , \new_[8867]_ , \new_[8870]_ ,
    \new_[8871]_ , \new_[8874]_ , \new_[8877]_ , \new_[8878]_ ,
    \new_[8881]_ , \new_[8884]_ , \new_[8885]_ , \new_[8888]_ ,
    \new_[8891]_ , \new_[8892]_ , \new_[8895]_ , \new_[8898]_ ,
    \new_[8899]_ , \new_[8902]_ , \new_[8905]_ , \new_[8906]_ ,
    \new_[8909]_ , \new_[8912]_ , \new_[8913]_ , \new_[8916]_ ,
    \new_[8919]_ , \new_[8920]_ , \new_[8923]_ , \new_[8926]_ ,
    \new_[8927]_ , \new_[8930]_ , \new_[8933]_ , \new_[8934]_ ,
    \new_[8937]_ , \new_[8940]_ , \new_[8941]_ , \new_[8944]_ ,
    \new_[8947]_ , \new_[8948]_ , \new_[8951]_ , \new_[8954]_ ,
    \new_[8955]_ , \new_[8958]_ , \new_[8961]_ , \new_[8962]_ ,
    \new_[8965]_ , \new_[8968]_ , \new_[8969]_ , \new_[8972]_ ,
    \new_[8975]_ , \new_[8976]_ , \new_[8979]_ , \new_[8982]_ ,
    \new_[8983]_ , \new_[8986]_ , \new_[8989]_ , \new_[8990]_ ,
    \new_[8993]_ , \new_[8996]_ , \new_[8997]_ , \new_[9000]_ ,
    \new_[9003]_ , \new_[9004]_ , \new_[9007]_ , \new_[9010]_ ,
    \new_[9011]_ , \new_[9014]_ , \new_[9017]_ , \new_[9018]_ ,
    \new_[9021]_ , \new_[9024]_ , \new_[9025]_ , \new_[9028]_ ,
    \new_[9031]_ , \new_[9032]_ , \new_[9035]_ , \new_[9038]_ ,
    \new_[9039]_ , \new_[9042]_ , \new_[9045]_ , \new_[9046]_ ,
    \new_[9049]_ , \new_[9052]_ , \new_[9053]_ , \new_[9056]_ ,
    \new_[9059]_ , \new_[9060]_ , \new_[9063]_ , \new_[9066]_ ,
    \new_[9067]_ , \new_[9070]_ , \new_[9073]_ , \new_[9074]_ ,
    \new_[9077]_ , \new_[9080]_ , \new_[9081]_ , \new_[9084]_ ,
    \new_[9087]_ , \new_[9088]_ , \new_[9091]_ , \new_[9094]_ ,
    \new_[9095]_ , \new_[9098]_ , \new_[9101]_ , \new_[9102]_ ,
    \new_[9105]_ , \new_[9108]_ , \new_[9109]_ , \new_[9112]_ ,
    \new_[9115]_ , \new_[9116]_ , \new_[9119]_ , \new_[9122]_ ,
    \new_[9123]_ , \new_[9126]_ , \new_[9129]_ , \new_[9130]_ ,
    \new_[9133]_ , \new_[9136]_ , \new_[9137]_ , \new_[9140]_ ,
    \new_[9143]_ , \new_[9144]_ , \new_[9147]_ , \new_[9150]_ ,
    \new_[9151]_ , \new_[9154]_ , \new_[9157]_ , \new_[9158]_ ,
    \new_[9161]_ , \new_[9164]_ , \new_[9165]_ , \new_[9168]_ ,
    \new_[9171]_ , \new_[9172]_ , \new_[9175]_ , \new_[9178]_ ,
    \new_[9179]_ , \new_[9182]_ , \new_[9185]_ , \new_[9186]_ ,
    \new_[9189]_ , \new_[9192]_ , \new_[9193]_ , \new_[9196]_ ,
    \new_[9199]_ , \new_[9200]_ , \new_[9203]_ , \new_[9206]_ ,
    \new_[9207]_ , \new_[9210]_ , \new_[9213]_ , \new_[9214]_ ,
    \new_[9217]_ , \new_[9220]_ , \new_[9221]_ , \new_[9224]_ ,
    \new_[9227]_ , \new_[9228]_ , \new_[9231]_ , \new_[9234]_ ,
    \new_[9235]_ , \new_[9238]_ , \new_[9241]_ , \new_[9242]_ ,
    \new_[9245]_ , \new_[9248]_ , \new_[9249]_ , \new_[9252]_ ,
    \new_[9255]_ , \new_[9256]_ , \new_[9259]_ , \new_[9262]_ ,
    \new_[9263]_ , \new_[9266]_ , \new_[9269]_ , \new_[9270]_ ,
    \new_[9273]_ , \new_[9276]_ , \new_[9277]_ , \new_[9280]_ ,
    \new_[9283]_ , \new_[9284]_ , \new_[9287]_ , \new_[9290]_ ,
    \new_[9291]_ , \new_[9294]_ , \new_[9297]_ , \new_[9298]_ ,
    \new_[9301]_ , \new_[9304]_ , \new_[9305]_ , \new_[9308]_ ,
    \new_[9311]_ , \new_[9312]_ , \new_[9315]_ , \new_[9318]_ ,
    \new_[9319]_ , \new_[9322]_ , \new_[9325]_ , \new_[9326]_ ,
    \new_[9329]_ , \new_[9332]_ , \new_[9333]_ , \new_[9336]_ ,
    \new_[9339]_ , \new_[9340]_ , \new_[9343]_ , \new_[9346]_ ,
    \new_[9347]_ , \new_[9350]_ , \new_[9353]_ , \new_[9354]_ ,
    \new_[9357]_ , \new_[9360]_ , \new_[9361]_ , \new_[9364]_ ,
    \new_[9367]_ , \new_[9368]_ , \new_[9371]_ , \new_[9374]_ ,
    \new_[9375]_ , \new_[9378]_ , \new_[9381]_ , \new_[9382]_ ,
    \new_[9385]_ , \new_[9388]_ , \new_[9389]_ , \new_[9392]_ ,
    \new_[9395]_ , \new_[9396]_ , \new_[9399]_ , \new_[9402]_ ,
    \new_[9403]_ , \new_[9406]_ , \new_[9409]_ , \new_[9410]_ ,
    \new_[9413]_ , \new_[9416]_ , \new_[9417]_ , \new_[9420]_ ,
    \new_[9423]_ , \new_[9424]_ , \new_[9427]_ , \new_[9430]_ ,
    \new_[9431]_ , \new_[9434]_ , \new_[9437]_ , \new_[9438]_ ,
    \new_[9441]_ , \new_[9444]_ , \new_[9445]_ , \new_[9448]_ ,
    \new_[9451]_ , \new_[9452]_ , \new_[9455]_ , \new_[9458]_ ,
    \new_[9459]_ , \new_[9462]_ , \new_[9465]_ , \new_[9466]_ ,
    \new_[9469]_ , \new_[9472]_ , \new_[9473]_ , \new_[9476]_ ,
    \new_[9479]_ , \new_[9480]_ , \new_[9483]_ , \new_[9486]_ ,
    \new_[9487]_ , \new_[9490]_ , \new_[9493]_ , \new_[9494]_ ,
    \new_[9497]_ , \new_[9500]_ , \new_[9501]_ , \new_[9504]_ ,
    \new_[9507]_ , \new_[9508]_ , \new_[9511]_ , \new_[9514]_ ,
    \new_[9515]_ , \new_[9518]_ , \new_[9521]_ , \new_[9522]_ ,
    \new_[9525]_ , \new_[9528]_ , \new_[9529]_ , \new_[9532]_ ,
    \new_[9535]_ , \new_[9536]_ , \new_[9539]_ , \new_[9542]_ ,
    \new_[9543]_ , \new_[9546]_ , \new_[9549]_ , \new_[9550]_ ,
    \new_[9553]_ , \new_[9556]_ , \new_[9557]_ , \new_[9560]_ ,
    \new_[9563]_ , \new_[9564]_ , \new_[9567]_ , \new_[9570]_ ,
    \new_[9571]_ , \new_[9574]_ , \new_[9577]_ , \new_[9578]_ ,
    \new_[9581]_ , \new_[9584]_ , \new_[9585]_ , \new_[9588]_ ,
    \new_[9591]_ , \new_[9592]_ , \new_[9595]_ , \new_[9598]_ ,
    \new_[9599]_ , \new_[9602]_ , \new_[9605]_ , \new_[9606]_ ,
    \new_[9609]_ , \new_[9612]_ , \new_[9613]_ , \new_[9616]_ ,
    \new_[9619]_ , \new_[9620]_ , \new_[9623]_ , \new_[9626]_ ,
    \new_[9627]_ , \new_[9630]_ , \new_[9633]_ , \new_[9634]_ ,
    \new_[9637]_ , \new_[9640]_ , \new_[9641]_ , \new_[9644]_ ,
    \new_[9647]_ , \new_[9648]_ , \new_[9651]_ , \new_[9654]_ ,
    \new_[9655]_ , \new_[9658]_ , \new_[9661]_ , \new_[9662]_ ,
    \new_[9665]_ , \new_[9668]_ , \new_[9669]_ , \new_[9672]_ ,
    \new_[9675]_ , \new_[9676]_ , \new_[9679]_ , \new_[9682]_ ,
    \new_[9683]_ , \new_[9686]_ , \new_[9689]_ , \new_[9690]_ ,
    \new_[9693]_ , \new_[9696]_ , \new_[9697]_ , \new_[9700]_ ,
    \new_[9703]_ , \new_[9704]_ , \new_[9707]_ , \new_[9710]_ ,
    \new_[9711]_ , \new_[9714]_ , \new_[9717]_ , \new_[9718]_ ,
    \new_[9721]_ , \new_[9724]_ , \new_[9725]_ , \new_[9728]_ ,
    \new_[9731]_ , \new_[9732]_ , \new_[9735]_ , \new_[9738]_ ,
    \new_[9739]_ , \new_[9742]_ , \new_[9745]_ , \new_[9746]_ ,
    \new_[9749]_ , \new_[9752]_ , \new_[9753]_ , \new_[9756]_ ,
    \new_[9759]_ , \new_[9760]_ , \new_[9763]_ , \new_[9766]_ ,
    \new_[9767]_ , \new_[9770]_ , \new_[9773]_ , \new_[9774]_ ,
    \new_[9777]_ , \new_[9780]_ , \new_[9781]_ , \new_[9784]_ ,
    \new_[9787]_ , \new_[9788]_ , \new_[9791]_ , \new_[9794]_ ,
    \new_[9795]_ , \new_[9798]_ , \new_[9801]_ , \new_[9802]_ ,
    \new_[9805]_ , \new_[9808]_ , \new_[9809]_ , \new_[9812]_ ,
    \new_[9815]_ , \new_[9816]_ , \new_[9819]_ , \new_[9822]_ ,
    \new_[9823]_ , \new_[9826]_ , \new_[9829]_ , \new_[9830]_ ,
    \new_[9833]_ , \new_[9836]_ , \new_[9837]_ , \new_[9840]_ ,
    \new_[9843]_ , \new_[9844]_ , \new_[9847]_ , \new_[9850]_ ,
    \new_[9851]_ , \new_[9854]_ , \new_[9857]_ , \new_[9858]_ ,
    \new_[9861]_ , \new_[9864]_ , \new_[9865]_ , \new_[9868]_ ,
    \new_[9871]_ , \new_[9872]_ , \new_[9875]_ , \new_[9878]_ ,
    \new_[9879]_ , \new_[9882]_ , \new_[9885]_ , \new_[9886]_ ,
    \new_[9889]_ , \new_[9892]_ , \new_[9893]_ , \new_[9896]_ ,
    \new_[9899]_ , \new_[9900]_ , \new_[9903]_ , \new_[9906]_ ,
    \new_[9907]_ , \new_[9910]_ , \new_[9913]_ , \new_[9914]_ ,
    \new_[9917]_ , \new_[9920]_ , \new_[9921]_ , \new_[9924]_ ,
    \new_[9927]_ , \new_[9928]_ , \new_[9931]_ , \new_[9934]_ ,
    \new_[9935]_ , \new_[9938]_ , \new_[9941]_ , \new_[9942]_ ,
    \new_[9945]_ , \new_[9948]_ , \new_[9949]_ , \new_[9952]_ ,
    \new_[9955]_ , \new_[9956]_ , \new_[9959]_ , \new_[9962]_ ,
    \new_[9963]_ , \new_[9966]_ , \new_[9969]_ , \new_[9970]_ ,
    \new_[9973]_ , \new_[9976]_ , \new_[9977]_ , \new_[9980]_ ,
    \new_[9983]_ , \new_[9984]_ , \new_[9987]_ , \new_[9990]_ ,
    \new_[9991]_ , \new_[9994]_ , \new_[9998]_ , \new_[9999]_ ,
    \new_[10000]_ , \new_[10003]_ , \new_[10006]_ , \new_[10007]_ ,
    \new_[10010]_ , \new_[10014]_ , \new_[10015]_ , \new_[10016]_ ,
    \new_[10019]_ , \new_[10022]_ , \new_[10023]_ , \new_[10026]_ ,
    \new_[10030]_ , \new_[10031]_ , \new_[10032]_ , \new_[10035]_ ,
    \new_[10038]_ , \new_[10039]_ , \new_[10042]_ , \new_[10046]_ ,
    \new_[10047]_ , \new_[10048]_ , \new_[10051]_ , \new_[10054]_ ,
    \new_[10055]_ , \new_[10058]_ , \new_[10062]_ , \new_[10063]_ ,
    \new_[10064]_ , \new_[10067]_ , \new_[10070]_ , \new_[10071]_ ,
    \new_[10074]_ , \new_[10078]_ , \new_[10079]_ , \new_[10080]_ ,
    \new_[10083]_ , \new_[10086]_ , \new_[10087]_ , \new_[10090]_ ,
    \new_[10094]_ , \new_[10095]_ , \new_[10096]_ , \new_[10099]_ ,
    \new_[10102]_ , \new_[10103]_ , \new_[10106]_ , \new_[10110]_ ,
    \new_[10111]_ , \new_[10112]_ , \new_[10115]_ , \new_[10118]_ ,
    \new_[10119]_ , \new_[10122]_ , \new_[10126]_ , \new_[10127]_ ,
    \new_[10128]_ , \new_[10131]_ , \new_[10134]_ , \new_[10135]_ ,
    \new_[10138]_ , \new_[10142]_ , \new_[10143]_ , \new_[10144]_ ,
    \new_[10147]_ , \new_[10150]_ , \new_[10151]_ , \new_[10154]_ ,
    \new_[10158]_ , \new_[10159]_ , \new_[10160]_ , \new_[10163]_ ,
    \new_[10166]_ , \new_[10167]_ , \new_[10170]_ , \new_[10174]_ ,
    \new_[10175]_ , \new_[10176]_ , \new_[10179]_ , \new_[10182]_ ,
    \new_[10183]_ , \new_[10186]_ , \new_[10190]_ , \new_[10191]_ ,
    \new_[10192]_ , \new_[10195]_ , \new_[10198]_ , \new_[10199]_ ,
    \new_[10202]_ , \new_[10206]_ , \new_[10207]_ , \new_[10208]_ ,
    \new_[10211]_ , \new_[10214]_ , \new_[10215]_ , \new_[10218]_ ,
    \new_[10222]_ , \new_[10223]_ , \new_[10224]_ , \new_[10227]_ ,
    \new_[10230]_ , \new_[10231]_ , \new_[10234]_ , \new_[10238]_ ,
    \new_[10239]_ , \new_[10240]_ , \new_[10243]_ , \new_[10246]_ ,
    \new_[10247]_ , \new_[10250]_ , \new_[10254]_ , \new_[10255]_ ,
    \new_[10256]_ , \new_[10259]_ , \new_[10262]_ , \new_[10263]_ ,
    \new_[10266]_ , \new_[10270]_ , \new_[10271]_ , \new_[10272]_ ,
    \new_[10275]_ , \new_[10278]_ , \new_[10279]_ , \new_[10282]_ ,
    \new_[10286]_ , \new_[10287]_ , \new_[10288]_ , \new_[10291]_ ,
    \new_[10294]_ , \new_[10295]_ , \new_[10298]_ , \new_[10302]_ ,
    \new_[10303]_ , \new_[10304]_ , \new_[10307]_ , \new_[10310]_ ,
    \new_[10311]_ , \new_[10314]_ , \new_[10318]_ , \new_[10319]_ ,
    \new_[10320]_ , \new_[10323]_ , \new_[10326]_ , \new_[10327]_ ,
    \new_[10330]_ , \new_[10334]_ , \new_[10335]_ , \new_[10336]_ ,
    \new_[10339]_ , \new_[10342]_ , \new_[10343]_ , \new_[10346]_ ,
    \new_[10350]_ , \new_[10351]_ , \new_[10352]_ , \new_[10355]_ ,
    \new_[10358]_ , \new_[10359]_ , \new_[10362]_ , \new_[10366]_ ,
    \new_[10367]_ , \new_[10368]_ , \new_[10371]_ , \new_[10374]_ ,
    \new_[10375]_ , \new_[10378]_ , \new_[10382]_ , \new_[10383]_ ,
    \new_[10384]_ , \new_[10387]_ , \new_[10390]_ , \new_[10391]_ ,
    \new_[10394]_ , \new_[10398]_ , \new_[10399]_ , \new_[10400]_ ,
    \new_[10403]_ , \new_[10406]_ , \new_[10407]_ , \new_[10410]_ ,
    \new_[10414]_ , \new_[10415]_ , \new_[10416]_ , \new_[10419]_ ,
    \new_[10422]_ , \new_[10423]_ , \new_[10426]_ , \new_[10430]_ ,
    \new_[10431]_ , \new_[10432]_ , \new_[10435]_ , \new_[10438]_ ,
    \new_[10439]_ , \new_[10442]_ , \new_[10446]_ , \new_[10447]_ ,
    \new_[10448]_ , \new_[10451]_ , \new_[10454]_ , \new_[10455]_ ,
    \new_[10458]_ , \new_[10462]_ , \new_[10463]_ , \new_[10464]_ ,
    \new_[10467]_ , \new_[10470]_ , \new_[10471]_ , \new_[10474]_ ,
    \new_[10478]_ , \new_[10479]_ , \new_[10480]_ , \new_[10483]_ ,
    \new_[10486]_ , \new_[10487]_ , \new_[10490]_ , \new_[10494]_ ,
    \new_[10495]_ , \new_[10496]_ , \new_[10499]_ , \new_[10502]_ ,
    \new_[10503]_ , \new_[10506]_ , \new_[10510]_ , \new_[10511]_ ,
    \new_[10512]_ , \new_[10515]_ , \new_[10518]_ , \new_[10519]_ ,
    \new_[10522]_ , \new_[10526]_ , \new_[10527]_ , \new_[10528]_ ,
    \new_[10531]_ , \new_[10534]_ , \new_[10535]_ , \new_[10538]_ ,
    \new_[10542]_ , \new_[10543]_ , \new_[10544]_ , \new_[10547]_ ,
    \new_[10550]_ , \new_[10551]_ , \new_[10554]_ , \new_[10558]_ ,
    \new_[10559]_ , \new_[10560]_ , \new_[10563]_ , \new_[10566]_ ,
    \new_[10567]_ , \new_[10570]_ , \new_[10574]_ , \new_[10575]_ ,
    \new_[10576]_ , \new_[10579]_ , \new_[10582]_ , \new_[10583]_ ,
    \new_[10586]_ , \new_[10590]_ , \new_[10591]_ , \new_[10592]_ ,
    \new_[10595]_ , \new_[10598]_ , \new_[10599]_ , \new_[10602]_ ,
    \new_[10606]_ , \new_[10607]_ , \new_[10608]_ , \new_[10611]_ ,
    \new_[10614]_ , \new_[10615]_ , \new_[10618]_ , \new_[10622]_ ,
    \new_[10623]_ , \new_[10624]_ , \new_[10627]_ , \new_[10630]_ ,
    \new_[10631]_ , \new_[10634]_ , \new_[10638]_ , \new_[10639]_ ,
    \new_[10640]_ , \new_[10643]_ , \new_[10646]_ , \new_[10647]_ ,
    \new_[10650]_ , \new_[10654]_ , \new_[10655]_ , \new_[10656]_ ,
    \new_[10659]_ , \new_[10662]_ , \new_[10663]_ , \new_[10666]_ ,
    \new_[10670]_ , \new_[10671]_ , \new_[10672]_ , \new_[10675]_ ,
    \new_[10678]_ , \new_[10679]_ , \new_[10682]_ , \new_[10686]_ ,
    \new_[10687]_ , \new_[10688]_ , \new_[10691]_ , \new_[10694]_ ,
    \new_[10695]_ , \new_[10698]_ , \new_[10702]_ , \new_[10703]_ ,
    \new_[10704]_ , \new_[10707]_ , \new_[10710]_ , \new_[10711]_ ,
    \new_[10714]_ , \new_[10718]_ , \new_[10719]_ , \new_[10720]_ ,
    \new_[10723]_ , \new_[10726]_ , \new_[10727]_ , \new_[10730]_ ,
    \new_[10734]_ , \new_[10735]_ , \new_[10736]_ , \new_[10739]_ ,
    \new_[10742]_ , \new_[10743]_ , \new_[10746]_ , \new_[10750]_ ,
    \new_[10751]_ , \new_[10752]_ , \new_[10755]_ , \new_[10758]_ ,
    \new_[10759]_ , \new_[10762]_ , \new_[10766]_ , \new_[10767]_ ,
    \new_[10768]_ , \new_[10771]_ , \new_[10774]_ , \new_[10775]_ ,
    \new_[10778]_ , \new_[10782]_ , \new_[10783]_ , \new_[10784]_ ,
    \new_[10787]_ , \new_[10790]_ , \new_[10791]_ , \new_[10794]_ ,
    \new_[10798]_ , \new_[10799]_ , \new_[10800]_ , \new_[10803]_ ,
    \new_[10806]_ , \new_[10807]_ , \new_[10810]_ , \new_[10814]_ ,
    \new_[10815]_ , \new_[10816]_ , \new_[10819]_ , \new_[10822]_ ,
    \new_[10823]_ , \new_[10826]_ , \new_[10830]_ , \new_[10831]_ ,
    \new_[10832]_ , \new_[10835]_ , \new_[10838]_ , \new_[10839]_ ,
    \new_[10842]_ , \new_[10846]_ , \new_[10847]_ , \new_[10848]_ ,
    \new_[10851]_ , \new_[10854]_ , \new_[10855]_ , \new_[10858]_ ,
    \new_[10862]_ , \new_[10863]_ , \new_[10864]_ , \new_[10867]_ ,
    \new_[10870]_ , \new_[10871]_ , \new_[10874]_ , \new_[10878]_ ,
    \new_[10879]_ , \new_[10880]_ , \new_[10883]_ , \new_[10886]_ ,
    \new_[10887]_ , \new_[10890]_ , \new_[10894]_ , \new_[10895]_ ,
    \new_[10896]_ , \new_[10899]_ , \new_[10902]_ , \new_[10903]_ ,
    \new_[10906]_ , \new_[10910]_ , \new_[10911]_ , \new_[10912]_ ,
    \new_[10915]_ , \new_[10918]_ , \new_[10919]_ , \new_[10922]_ ,
    \new_[10926]_ , \new_[10927]_ , \new_[10928]_ , \new_[10931]_ ,
    \new_[10934]_ , \new_[10935]_ , \new_[10938]_ , \new_[10942]_ ,
    \new_[10943]_ , \new_[10944]_ , \new_[10947]_ , \new_[10950]_ ,
    \new_[10951]_ , \new_[10954]_ , \new_[10958]_ , \new_[10959]_ ,
    \new_[10960]_ , \new_[10963]_ , \new_[10966]_ , \new_[10967]_ ,
    \new_[10970]_ , \new_[10974]_ , \new_[10975]_ , \new_[10976]_ ,
    \new_[10979]_ , \new_[10982]_ , \new_[10983]_ , \new_[10986]_ ,
    \new_[10990]_ , \new_[10991]_ , \new_[10992]_ , \new_[10995]_ ,
    \new_[10998]_ , \new_[10999]_ , \new_[11002]_ , \new_[11006]_ ,
    \new_[11007]_ , \new_[11008]_ , \new_[11011]_ , \new_[11014]_ ,
    \new_[11015]_ , \new_[11018]_ , \new_[11022]_ , \new_[11023]_ ,
    \new_[11024]_ , \new_[11027]_ , \new_[11030]_ , \new_[11031]_ ,
    \new_[11034]_ , \new_[11038]_ , \new_[11039]_ , \new_[11040]_ ,
    \new_[11043]_ , \new_[11046]_ , \new_[11047]_ , \new_[11050]_ ,
    \new_[11054]_ , \new_[11055]_ , \new_[11056]_ , \new_[11059]_ ,
    \new_[11062]_ , \new_[11063]_ , \new_[11066]_ , \new_[11070]_ ,
    \new_[11071]_ , \new_[11072]_ , \new_[11075]_ , \new_[11078]_ ,
    \new_[11079]_ , \new_[11082]_ , \new_[11086]_ , \new_[11087]_ ,
    \new_[11088]_ , \new_[11091]_ , \new_[11094]_ , \new_[11095]_ ,
    \new_[11098]_ , \new_[11102]_ , \new_[11103]_ , \new_[11104]_ ,
    \new_[11107]_ , \new_[11110]_ , \new_[11111]_ , \new_[11114]_ ,
    \new_[11118]_ , \new_[11119]_ , \new_[11120]_ , \new_[11123]_ ,
    \new_[11126]_ , \new_[11127]_ , \new_[11130]_ , \new_[11134]_ ,
    \new_[11135]_ , \new_[11136]_ , \new_[11139]_ , \new_[11142]_ ,
    \new_[11143]_ , \new_[11146]_ , \new_[11150]_ , \new_[11151]_ ,
    \new_[11152]_ , \new_[11155]_ , \new_[11158]_ , \new_[11159]_ ,
    \new_[11162]_ , \new_[11166]_ , \new_[11167]_ , \new_[11168]_ ,
    \new_[11171]_ , \new_[11174]_ , \new_[11175]_ , \new_[11178]_ ,
    \new_[11182]_ , \new_[11183]_ , \new_[11184]_ , \new_[11187]_ ,
    \new_[11190]_ , \new_[11191]_ , \new_[11194]_ , \new_[11198]_ ,
    \new_[11199]_ , \new_[11200]_ , \new_[11203]_ , \new_[11206]_ ,
    \new_[11207]_ , \new_[11210]_ , \new_[11214]_ , \new_[11215]_ ,
    \new_[11216]_ , \new_[11219]_ , \new_[11222]_ , \new_[11223]_ ,
    \new_[11226]_ , \new_[11230]_ , \new_[11231]_ , \new_[11232]_ ,
    \new_[11235]_ , \new_[11238]_ , \new_[11239]_ , \new_[11242]_ ,
    \new_[11246]_ , \new_[11247]_ , \new_[11248]_ , \new_[11251]_ ,
    \new_[11254]_ , \new_[11255]_ , \new_[11258]_ , \new_[11262]_ ,
    \new_[11263]_ , \new_[11264]_ , \new_[11267]_ , \new_[11270]_ ,
    \new_[11271]_ , \new_[11274]_ , \new_[11278]_ , \new_[11279]_ ,
    \new_[11280]_ , \new_[11283]_ , \new_[11286]_ , \new_[11287]_ ,
    \new_[11290]_ , \new_[11294]_ , \new_[11295]_ , \new_[11296]_ ,
    \new_[11299]_ , \new_[11302]_ , \new_[11303]_ , \new_[11306]_ ,
    \new_[11310]_ , \new_[11311]_ , \new_[11312]_ , \new_[11315]_ ,
    \new_[11318]_ , \new_[11319]_ , \new_[11322]_ , \new_[11326]_ ,
    \new_[11327]_ , \new_[11328]_ , \new_[11331]_ , \new_[11334]_ ,
    \new_[11335]_ , \new_[11338]_ , \new_[11342]_ , \new_[11343]_ ,
    \new_[11344]_ , \new_[11347]_ , \new_[11350]_ , \new_[11351]_ ,
    \new_[11354]_ , \new_[11358]_ , \new_[11359]_ , \new_[11360]_ ,
    \new_[11363]_ , \new_[11366]_ , \new_[11367]_ , \new_[11370]_ ,
    \new_[11374]_ , \new_[11375]_ , \new_[11376]_ , \new_[11379]_ ,
    \new_[11382]_ , \new_[11383]_ , \new_[11386]_ , \new_[11390]_ ,
    \new_[11391]_ , \new_[11392]_ , \new_[11395]_ , \new_[11398]_ ,
    \new_[11399]_ , \new_[11402]_ , \new_[11406]_ , \new_[11407]_ ,
    \new_[11408]_ , \new_[11411]_ , \new_[11414]_ , \new_[11415]_ ,
    \new_[11418]_ , \new_[11422]_ , \new_[11423]_ , \new_[11424]_ ,
    \new_[11427]_ , \new_[11430]_ , \new_[11431]_ , \new_[11434]_ ,
    \new_[11438]_ , \new_[11439]_ , \new_[11440]_ , \new_[11443]_ ,
    \new_[11446]_ , \new_[11447]_ , \new_[11450]_ , \new_[11454]_ ,
    \new_[11455]_ , \new_[11456]_ , \new_[11459]_ , \new_[11462]_ ,
    \new_[11463]_ , \new_[11466]_ , \new_[11470]_ , \new_[11471]_ ,
    \new_[11472]_ , \new_[11475]_ , \new_[11478]_ , \new_[11479]_ ,
    \new_[11482]_ , \new_[11486]_ , \new_[11487]_ , \new_[11488]_ ,
    \new_[11491]_ , \new_[11494]_ , \new_[11495]_ , \new_[11498]_ ,
    \new_[11502]_ , \new_[11503]_ , \new_[11504]_ , \new_[11507]_ ,
    \new_[11510]_ , \new_[11511]_ , \new_[11514]_ , \new_[11518]_ ,
    \new_[11519]_ , \new_[11520]_ , \new_[11523]_ , \new_[11526]_ ,
    \new_[11527]_ , \new_[11530]_ , \new_[11534]_ , \new_[11535]_ ,
    \new_[11536]_ , \new_[11539]_ , \new_[11542]_ , \new_[11543]_ ,
    \new_[11546]_ , \new_[11550]_ , \new_[11551]_ , \new_[11552]_ ,
    \new_[11555]_ , \new_[11558]_ , \new_[11559]_ , \new_[11562]_ ,
    \new_[11566]_ , \new_[11567]_ , \new_[11568]_ , \new_[11571]_ ,
    \new_[11574]_ , \new_[11575]_ , \new_[11578]_ , \new_[11582]_ ,
    \new_[11583]_ , \new_[11584]_ , \new_[11587]_ , \new_[11590]_ ,
    \new_[11591]_ , \new_[11594]_ , \new_[11598]_ , \new_[11599]_ ,
    \new_[11600]_ , \new_[11603]_ , \new_[11606]_ , \new_[11607]_ ,
    \new_[11610]_ , \new_[11614]_ , \new_[11615]_ , \new_[11616]_ ,
    \new_[11619]_ , \new_[11622]_ , \new_[11623]_ , \new_[11626]_ ,
    \new_[11630]_ , \new_[11631]_ , \new_[11632]_ , \new_[11635]_ ,
    \new_[11638]_ , \new_[11639]_ , \new_[11642]_ , \new_[11646]_ ,
    \new_[11647]_ , \new_[11648]_ , \new_[11651]_ , \new_[11654]_ ,
    \new_[11655]_ , \new_[11658]_ , \new_[11662]_ , \new_[11663]_ ,
    \new_[11664]_ , \new_[11667]_ , \new_[11670]_ , \new_[11671]_ ,
    \new_[11674]_ , \new_[11678]_ , \new_[11679]_ , \new_[11680]_ ,
    \new_[11683]_ , \new_[11686]_ , \new_[11687]_ , \new_[11690]_ ,
    \new_[11694]_ , \new_[11695]_ , \new_[11696]_ , \new_[11699]_ ,
    \new_[11702]_ , \new_[11703]_ , \new_[11706]_ , \new_[11710]_ ,
    \new_[11711]_ , \new_[11712]_ , \new_[11715]_ , \new_[11718]_ ,
    \new_[11719]_ , \new_[11722]_ , \new_[11726]_ , \new_[11727]_ ,
    \new_[11728]_ , \new_[11731]_ , \new_[11734]_ , \new_[11735]_ ,
    \new_[11738]_ , \new_[11742]_ , \new_[11743]_ , \new_[11744]_ ,
    \new_[11747]_ , \new_[11750]_ , \new_[11751]_ , \new_[11754]_ ,
    \new_[11758]_ , \new_[11759]_ , \new_[11760]_ , \new_[11763]_ ,
    \new_[11766]_ , \new_[11767]_ , \new_[11770]_ , \new_[11774]_ ,
    \new_[11775]_ , \new_[11776]_ , \new_[11779]_ , \new_[11782]_ ,
    \new_[11783]_ , \new_[11786]_ , \new_[11790]_ , \new_[11791]_ ,
    \new_[11792]_ , \new_[11795]_ , \new_[11798]_ , \new_[11799]_ ,
    \new_[11802]_ , \new_[11806]_ , \new_[11807]_ , \new_[11808]_ ,
    \new_[11811]_ , \new_[11814]_ , \new_[11815]_ , \new_[11818]_ ,
    \new_[11822]_ , \new_[11823]_ , \new_[11824]_ , \new_[11827]_ ,
    \new_[11830]_ , \new_[11831]_ , \new_[11834]_ , \new_[11838]_ ,
    \new_[11839]_ , \new_[11840]_ , \new_[11843]_ , \new_[11846]_ ,
    \new_[11847]_ , \new_[11850]_ , \new_[11854]_ , \new_[11855]_ ,
    \new_[11856]_ , \new_[11859]_ , \new_[11862]_ , \new_[11863]_ ,
    \new_[11866]_ , \new_[11870]_ , \new_[11871]_ , \new_[11872]_ ,
    \new_[11875]_ , \new_[11878]_ , \new_[11879]_ , \new_[11882]_ ,
    \new_[11886]_ , \new_[11887]_ , \new_[11888]_ , \new_[11891]_ ,
    \new_[11894]_ , \new_[11895]_ , \new_[11898]_ , \new_[11902]_ ,
    \new_[11903]_ , \new_[11904]_ , \new_[11907]_ , \new_[11910]_ ,
    \new_[11911]_ , \new_[11914]_ , \new_[11918]_ , \new_[11919]_ ,
    \new_[11920]_ , \new_[11923]_ , \new_[11926]_ , \new_[11927]_ ,
    \new_[11930]_ , \new_[11934]_ , \new_[11935]_ , \new_[11936]_ ,
    \new_[11939]_ , \new_[11942]_ , \new_[11943]_ , \new_[11946]_ ,
    \new_[11950]_ , \new_[11951]_ , \new_[11952]_ , \new_[11955]_ ,
    \new_[11958]_ , \new_[11959]_ , \new_[11962]_ , \new_[11966]_ ,
    \new_[11967]_ , \new_[11968]_ , \new_[11971]_ , \new_[11974]_ ,
    \new_[11975]_ , \new_[11978]_ , \new_[11982]_ , \new_[11983]_ ,
    \new_[11984]_ , \new_[11987]_ , \new_[11990]_ , \new_[11991]_ ,
    \new_[11994]_ , \new_[11998]_ , \new_[11999]_ , \new_[12000]_ ,
    \new_[12003]_ , \new_[12006]_ , \new_[12007]_ , \new_[12010]_ ,
    \new_[12014]_ , \new_[12015]_ , \new_[12016]_ , \new_[12019]_ ,
    \new_[12022]_ , \new_[12023]_ , \new_[12026]_ , \new_[12030]_ ,
    \new_[12031]_ , \new_[12032]_ , \new_[12035]_ , \new_[12038]_ ,
    \new_[12039]_ , \new_[12042]_ , \new_[12046]_ , \new_[12047]_ ,
    \new_[12048]_ , \new_[12051]_ , \new_[12054]_ , \new_[12055]_ ,
    \new_[12058]_ , \new_[12062]_ , \new_[12063]_ , \new_[12064]_ ,
    \new_[12067]_ , \new_[12070]_ , \new_[12071]_ , \new_[12074]_ ,
    \new_[12078]_ , \new_[12079]_ , \new_[12080]_ , \new_[12083]_ ,
    \new_[12086]_ , \new_[12087]_ , \new_[12090]_ , \new_[12094]_ ,
    \new_[12095]_ , \new_[12096]_ , \new_[12099]_ , \new_[12102]_ ,
    \new_[12103]_ , \new_[12106]_ , \new_[12110]_ , \new_[12111]_ ,
    \new_[12112]_ , \new_[12115]_ , \new_[12118]_ , \new_[12119]_ ,
    \new_[12122]_ , \new_[12126]_ , \new_[12127]_ , \new_[12128]_ ,
    \new_[12131]_ , \new_[12134]_ , \new_[12135]_ , \new_[12138]_ ,
    \new_[12142]_ , \new_[12143]_ , \new_[12144]_ , \new_[12147]_ ,
    \new_[12150]_ , \new_[12151]_ , \new_[12154]_ , \new_[12158]_ ,
    \new_[12159]_ , \new_[12160]_ , \new_[12163]_ , \new_[12166]_ ,
    \new_[12167]_ , \new_[12170]_ , \new_[12174]_ , \new_[12175]_ ,
    \new_[12176]_ , \new_[12179]_ , \new_[12182]_ , \new_[12183]_ ,
    \new_[12186]_ , \new_[12190]_ , \new_[12191]_ , \new_[12192]_ ,
    \new_[12195]_ , \new_[12198]_ , \new_[12199]_ , \new_[12202]_ ,
    \new_[12206]_ , \new_[12207]_ , \new_[12208]_ , \new_[12211]_ ,
    \new_[12214]_ , \new_[12215]_ , \new_[12218]_ , \new_[12222]_ ,
    \new_[12223]_ , \new_[12224]_ , \new_[12227]_ , \new_[12230]_ ,
    \new_[12231]_ , \new_[12234]_ , \new_[12238]_ , \new_[12239]_ ,
    \new_[12240]_ , \new_[12243]_ , \new_[12246]_ , \new_[12247]_ ,
    \new_[12250]_ , \new_[12254]_ , \new_[12255]_ , \new_[12256]_ ,
    \new_[12259]_ , \new_[12262]_ , \new_[12263]_ , \new_[12266]_ ,
    \new_[12270]_ , \new_[12271]_ , \new_[12272]_ , \new_[12275]_ ,
    \new_[12278]_ , \new_[12279]_ , \new_[12282]_ , \new_[12286]_ ,
    \new_[12287]_ , \new_[12288]_ , \new_[12291]_ , \new_[12294]_ ,
    \new_[12295]_ , \new_[12298]_ , \new_[12302]_ , \new_[12303]_ ,
    \new_[12304]_ , \new_[12307]_ , \new_[12310]_ , \new_[12311]_ ,
    \new_[12314]_ , \new_[12318]_ , \new_[12319]_ , \new_[12320]_ ,
    \new_[12323]_ , \new_[12326]_ , \new_[12327]_ , \new_[12330]_ ,
    \new_[12334]_ , \new_[12335]_ , \new_[12336]_ , \new_[12339]_ ,
    \new_[12342]_ , \new_[12343]_ , \new_[12346]_ , \new_[12350]_ ,
    \new_[12351]_ , \new_[12352]_ , \new_[12355]_ , \new_[12358]_ ,
    \new_[12359]_ , \new_[12362]_ , \new_[12366]_ , \new_[12367]_ ,
    \new_[12368]_ , \new_[12371]_ , \new_[12374]_ , \new_[12375]_ ,
    \new_[12378]_ , \new_[12382]_ , \new_[12383]_ , \new_[12384]_ ,
    \new_[12387]_ , \new_[12390]_ , \new_[12391]_ , \new_[12394]_ ,
    \new_[12398]_ , \new_[12399]_ , \new_[12400]_ , \new_[12403]_ ,
    \new_[12406]_ , \new_[12407]_ , \new_[12410]_ , \new_[12414]_ ,
    \new_[12415]_ , \new_[12416]_ , \new_[12419]_ , \new_[12422]_ ,
    \new_[12423]_ , \new_[12426]_ , \new_[12430]_ , \new_[12431]_ ,
    \new_[12432]_ , \new_[12435]_ , \new_[12438]_ , \new_[12439]_ ,
    \new_[12442]_ , \new_[12446]_ , \new_[12447]_ , \new_[12448]_ ,
    \new_[12451]_ , \new_[12454]_ , \new_[12455]_ , \new_[12458]_ ,
    \new_[12462]_ , \new_[12463]_ , \new_[12464]_ , \new_[12467]_ ,
    \new_[12470]_ , \new_[12471]_ , \new_[12474]_ , \new_[12478]_ ,
    \new_[12479]_ , \new_[12480]_ , \new_[12483]_ , \new_[12486]_ ,
    \new_[12487]_ , \new_[12490]_ , \new_[12494]_ , \new_[12495]_ ,
    \new_[12496]_ , \new_[12499]_ , \new_[12502]_ , \new_[12503]_ ,
    \new_[12506]_ , \new_[12510]_ , \new_[12511]_ , \new_[12512]_ ,
    \new_[12515]_ , \new_[12518]_ , \new_[12519]_ , \new_[12522]_ ,
    \new_[12526]_ , \new_[12527]_ , \new_[12528]_ , \new_[12531]_ ,
    \new_[12534]_ , \new_[12535]_ , \new_[12538]_ , \new_[12542]_ ,
    \new_[12543]_ , \new_[12544]_ , \new_[12547]_ , \new_[12550]_ ,
    \new_[12551]_ , \new_[12554]_ , \new_[12558]_ , \new_[12559]_ ,
    \new_[12560]_ , \new_[12563]_ , \new_[12566]_ , \new_[12567]_ ,
    \new_[12570]_ , \new_[12574]_ , \new_[12575]_ , \new_[12576]_ ,
    \new_[12579]_ , \new_[12582]_ , \new_[12583]_ , \new_[12586]_ ,
    \new_[12590]_ , \new_[12591]_ , \new_[12592]_ , \new_[12595]_ ,
    \new_[12598]_ , \new_[12599]_ , \new_[12602]_ , \new_[12606]_ ,
    \new_[12607]_ , \new_[12608]_ , \new_[12611]_ , \new_[12614]_ ,
    \new_[12615]_ , \new_[12618]_ , \new_[12622]_ , \new_[12623]_ ,
    \new_[12624]_ , \new_[12627]_ , \new_[12630]_ , \new_[12631]_ ,
    \new_[12634]_ , \new_[12638]_ , \new_[12639]_ , \new_[12640]_ ,
    \new_[12643]_ , \new_[12646]_ , \new_[12647]_ , \new_[12650]_ ,
    \new_[12654]_ , \new_[12655]_ , \new_[12656]_ , \new_[12659]_ ,
    \new_[12662]_ , \new_[12663]_ , \new_[12666]_ , \new_[12670]_ ,
    \new_[12671]_ , \new_[12672]_ , \new_[12675]_ , \new_[12678]_ ,
    \new_[12679]_ , \new_[12682]_ , \new_[12686]_ , \new_[12687]_ ,
    \new_[12688]_ , \new_[12691]_ , \new_[12694]_ , \new_[12695]_ ,
    \new_[12698]_ , \new_[12702]_ , \new_[12703]_ , \new_[12704]_ ,
    \new_[12707]_ , \new_[12710]_ , \new_[12711]_ , \new_[12714]_ ,
    \new_[12718]_ , \new_[12719]_ , \new_[12720]_ , \new_[12723]_ ,
    \new_[12726]_ , \new_[12727]_ , \new_[12730]_ , \new_[12734]_ ,
    \new_[12735]_ , \new_[12736]_ , \new_[12739]_ , \new_[12742]_ ,
    \new_[12743]_ , \new_[12746]_ , \new_[12750]_ , \new_[12751]_ ,
    \new_[12752]_ , \new_[12755]_ , \new_[12758]_ , \new_[12759]_ ,
    \new_[12762]_ , \new_[12766]_ , \new_[12767]_ , \new_[12768]_ ,
    \new_[12771]_ , \new_[12774]_ , \new_[12775]_ , \new_[12778]_ ,
    \new_[12782]_ , \new_[12783]_ , \new_[12784]_ , \new_[12787]_ ,
    \new_[12790]_ , \new_[12791]_ , \new_[12794]_ , \new_[12798]_ ,
    \new_[12799]_ , \new_[12800]_ , \new_[12803]_ , \new_[12806]_ ,
    \new_[12807]_ , \new_[12810]_ , \new_[12814]_ , \new_[12815]_ ,
    \new_[12816]_ , \new_[12819]_ , \new_[12822]_ , \new_[12823]_ ,
    \new_[12826]_ , \new_[12830]_ , \new_[12831]_ , \new_[12832]_ ,
    \new_[12835]_ , \new_[12838]_ , \new_[12839]_ , \new_[12842]_ ,
    \new_[12846]_ , \new_[12847]_ , \new_[12848]_ , \new_[12851]_ ,
    \new_[12854]_ , \new_[12855]_ , \new_[12858]_ , \new_[12862]_ ,
    \new_[12863]_ , \new_[12864]_ , \new_[12867]_ , \new_[12870]_ ,
    \new_[12871]_ , \new_[12874]_ , \new_[12878]_ , \new_[12879]_ ,
    \new_[12880]_ , \new_[12883]_ , \new_[12886]_ , \new_[12887]_ ,
    \new_[12890]_ , \new_[12894]_ , \new_[12895]_ , \new_[12896]_ ,
    \new_[12899]_ , \new_[12902]_ , \new_[12903]_ , \new_[12906]_ ,
    \new_[12910]_ , \new_[12911]_ , \new_[12912]_ , \new_[12915]_ ,
    \new_[12918]_ , \new_[12919]_ , \new_[12922]_ , \new_[12926]_ ,
    \new_[12927]_ , \new_[12928]_ , \new_[12931]_ , \new_[12934]_ ,
    \new_[12935]_ , \new_[12938]_ , \new_[12942]_ , \new_[12943]_ ,
    \new_[12944]_ , \new_[12947]_ , \new_[12950]_ , \new_[12951]_ ,
    \new_[12954]_ , \new_[12958]_ , \new_[12959]_ , \new_[12960]_ ,
    \new_[12963]_ , \new_[12966]_ , \new_[12967]_ , \new_[12970]_ ,
    \new_[12974]_ , \new_[12975]_ , \new_[12976]_ , \new_[12979]_ ,
    \new_[12982]_ , \new_[12983]_ , \new_[12986]_ , \new_[12990]_ ,
    \new_[12991]_ , \new_[12992]_ , \new_[12995]_ , \new_[12998]_ ,
    \new_[12999]_ , \new_[13002]_ , \new_[13006]_ , \new_[13007]_ ,
    \new_[13008]_ , \new_[13011]_ , \new_[13014]_ , \new_[13015]_ ,
    \new_[13018]_ , \new_[13022]_ , \new_[13023]_ , \new_[13024]_ ,
    \new_[13027]_ , \new_[13030]_ , \new_[13031]_ , \new_[13034]_ ,
    \new_[13038]_ , \new_[13039]_ , \new_[13040]_ , \new_[13043]_ ,
    \new_[13046]_ , \new_[13047]_ , \new_[13050]_ , \new_[13054]_ ,
    \new_[13055]_ , \new_[13056]_ , \new_[13059]_ , \new_[13062]_ ,
    \new_[13063]_ , \new_[13066]_ , \new_[13070]_ , \new_[13071]_ ,
    \new_[13072]_ , \new_[13075]_ , \new_[13078]_ , \new_[13079]_ ,
    \new_[13082]_ , \new_[13086]_ , \new_[13087]_ , \new_[13088]_ ,
    \new_[13091]_ , \new_[13094]_ , \new_[13095]_ , \new_[13098]_ ,
    \new_[13102]_ , \new_[13103]_ , \new_[13104]_ , \new_[13107]_ ,
    \new_[13110]_ , \new_[13111]_ , \new_[13114]_ , \new_[13118]_ ,
    \new_[13119]_ , \new_[13120]_ , \new_[13123]_ , \new_[13126]_ ,
    \new_[13127]_ , \new_[13130]_ , \new_[13134]_ , \new_[13135]_ ,
    \new_[13136]_ , \new_[13139]_ , \new_[13142]_ , \new_[13143]_ ,
    \new_[13146]_ , \new_[13150]_ , \new_[13151]_ , \new_[13152]_ ,
    \new_[13155]_ , \new_[13158]_ , \new_[13159]_ , \new_[13162]_ ,
    \new_[13166]_ , \new_[13167]_ , \new_[13168]_ , \new_[13171]_ ,
    \new_[13174]_ , \new_[13175]_ , \new_[13178]_ , \new_[13182]_ ,
    \new_[13183]_ , \new_[13184]_ , \new_[13187]_ , \new_[13190]_ ,
    \new_[13191]_ , \new_[13194]_ , \new_[13198]_ , \new_[13199]_ ,
    \new_[13200]_ , \new_[13203]_ , \new_[13206]_ , \new_[13207]_ ,
    \new_[13210]_ , \new_[13214]_ , \new_[13215]_ , \new_[13216]_ ,
    \new_[13219]_ , \new_[13222]_ , \new_[13223]_ , \new_[13226]_ ,
    \new_[13230]_ , \new_[13231]_ , \new_[13232]_ , \new_[13235]_ ,
    \new_[13238]_ , \new_[13239]_ , \new_[13242]_ , \new_[13246]_ ,
    \new_[13247]_ , \new_[13248]_ , \new_[13251]_ , \new_[13254]_ ,
    \new_[13255]_ , \new_[13258]_ , \new_[13262]_ , \new_[13263]_ ,
    \new_[13264]_ , \new_[13267]_ , \new_[13270]_ , \new_[13271]_ ,
    \new_[13274]_ , \new_[13278]_ , \new_[13279]_ , \new_[13280]_ ,
    \new_[13283]_ , \new_[13286]_ , \new_[13287]_ , \new_[13290]_ ,
    \new_[13294]_ , \new_[13295]_ , \new_[13296]_ , \new_[13299]_ ,
    \new_[13302]_ , \new_[13303]_ , \new_[13306]_ , \new_[13310]_ ,
    \new_[13311]_ , \new_[13312]_ , \new_[13315]_ , \new_[13318]_ ,
    \new_[13319]_ , \new_[13322]_ , \new_[13326]_ , \new_[13327]_ ,
    \new_[13328]_ , \new_[13331]_ , \new_[13334]_ , \new_[13335]_ ,
    \new_[13338]_ , \new_[13342]_ , \new_[13343]_ , \new_[13344]_ ,
    \new_[13347]_ , \new_[13350]_ , \new_[13351]_ , \new_[13354]_ ,
    \new_[13358]_ , \new_[13359]_ , \new_[13360]_ , \new_[13363]_ ,
    \new_[13366]_ , \new_[13367]_ , \new_[13370]_ , \new_[13374]_ ,
    \new_[13375]_ , \new_[13376]_ , \new_[13379]_ , \new_[13382]_ ,
    \new_[13383]_ , \new_[13386]_ , \new_[13390]_ , \new_[13391]_ ,
    \new_[13392]_ , \new_[13395]_ , \new_[13398]_ , \new_[13399]_ ,
    \new_[13402]_ , \new_[13406]_ , \new_[13407]_ , \new_[13408]_ ,
    \new_[13411]_ , \new_[13414]_ , \new_[13415]_ , \new_[13418]_ ,
    \new_[13422]_ , \new_[13423]_ , \new_[13424]_ , \new_[13427]_ ,
    \new_[13430]_ , \new_[13431]_ , \new_[13434]_ , \new_[13438]_ ,
    \new_[13439]_ , \new_[13440]_ , \new_[13443]_ , \new_[13446]_ ,
    \new_[13447]_ , \new_[13450]_ , \new_[13454]_ , \new_[13455]_ ,
    \new_[13456]_ , \new_[13459]_ , \new_[13462]_ , \new_[13463]_ ,
    \new_[13466]_ , \new_[13470]_ , \new_[13471]_ , \new_[13472]_ ,
    \new_[13475]_ , \new_[13478]_ , \new_[13479]_ , \new_[13482]_ ,
    \new_[13486]_ , \new_[13487]_ , \new_[13488]_ , \new_[13491]_ ,
    \new_[13494]_ , \new_[13495]_ , \new_[13498]_ , \new_[13502]_ ,
    \new_[13503]_ , \new_[13504]_ , \new_[13507]_ , \new_[13510]_ ,
    \new_[13511]_ , \new_[13514]_ , \new_[13518]_ , \new_[13519]_ ,
    \new_[13520]_ , \new_[13523]_ , \new_[13526]_ , \new_[13527]_ ,
    \new_[13530]_ , \new_[13534]_ , \new_[13535]_ , \new_[13536]_ ,
    \new_[13539]_ , \new_[13542]_ , \new_[13543]_ , \new_[13546]_ ,
    \new_[13550]_ , \new_[13551]_ , \new_[13552]_ , \new_[13555]_ ,
    \new_[13558]_ , \new_[13559]_ , \new_[13562]_ , \new_[13566]_ ,
    \new_[13567]_ , \new_[13568]_ , \new_[13571]_ , \new_[13574]_ ,
    \new_[13575]_ , \new_[13578]_ , \new_[13582]_ , \new_[13583]_ ,
    \new_[13584]_ , \new_[13587]_ , \new_[13590]_ , \new_[13591]_ ,
    \new_[13594]_ , \new_[13598]_ , \new_[13599]_ , \new_[13600]_ ,
    \new_[13603]_ , \new_[13606]_ , \new_[13607]_ , \new_[13610]_ ,
    \new_[13614]_ , \new_[13615]_ , \new_[13616]_ , \new_[13619]_ ,
    \new_[13622]_ , \new_[13623]_ , \new_[13626]_ , \new_[13630]_ ,
    \new_[13631]_ , \new_[13632]_ , \new_[13635]_ , \new_[13638]_ ,
    \new_[13639]_ , \new_[13642]_ , \new_[13646]_ , \new_[13647]_ ,
    \new_[13648]_ , \new_[13651]_ , \new_[13654]_ , \new_[13655]_ ,
    \new_[13658]_ , \new_[13662]_ , \new_[13663]_ , \new_[13664]_ ,
    \new_[13667]_ , \new_[13670]_ , \new_[13671]_ , \new_[13674]_ ,
    \new_[13678]_ , \new_[13679]_ , \new_[13680]_ , \new_[13683]_ ,
    \new_[13686]_ , \new_[13687]_ , \new_[13690]_ , \new_[13694]_ ,
    \new_[13695]_ , \new_[13696]_ , \new_[13699]_ , \new_[13702]_ ,
    \new_[13703]_ , \new_[13706]_ , \new_[13710]_ , \new_[13711]_ ,
    \new_[13712]_ , \new_[13715]_ , \new_[13718]_ , \new_[13719]_ ,
    \new_[13722]_ , \new_[13726]_ , \new_[13727]_ , \new_[13728]_ ,
    \new_[13731]_ , \new_[13734]_ , \new_[13735]_ , \new_[13738]_ ,
    \new_[13742]_ , \new_[13743]_ , \new_[13744]_ , \new_[13747]_ ,
    \new_[13750]_ , \new_[13751]_ , \new_[13754]_ , \new_[13758]_ ,
    \new_[13759]_ , \new_[13760]_ , \new_[13763]_ , \new_[13766]_ ,
    \new_[13767]_ , \new_[13770]_ , \new_[13774]_ , \new_[13775]_ ,
    \new_[13776]_ , \new_[13779]_ , \new_[13782]_ , \new_[13783]_ ,
    \new_[13786]_ , \new_[13790]_ , \new_[13791]_ , \new_[13792]_ ,
    \new_[13795]_ , \new_[13798]_ , \new_[13799]_ , \new_[13802]_ ,
    \new_[13806]_ , \new_[13807]_ , \new_[13808]_ , \new_[13811]_ ,
    \new_[13814]_ , \new_[13815]_ , \new_[13818]_ , \new_[13822]_ ,
    \new_[13823]_ , \new_[13824]_ , \new_[13827]_ , \new_[13830]_ ,
    \new_[13831]_ , \new_[13834]_ , \new_[13838]_ , \new_[13839]_ ,
    \new_[13840]_ , \new_[13843]_ , \new_[13846]_ , \new_[13847]_ ,
    \new_[13850]_ , \new_[13854]_ , \new_[13855]_ , \new_[13856]_ ,
    \new_[13859]_ , \new_[13862]_ , \new_[13863]_ , \new_[13866]_ ,
    \new_[13870]_ , \new_[13871]_ , \new_[13872]_ , \new_[13875]_ ,
    \new_[13878]_ , \new_[13879]_ , \new_[13882]_ , \new_[13886]_ ,
    \new_[13887]_ , \new_[13888]_ , \new_[13891]_ , \new_[13894]_ ,
    \new_[13895]_ , \new_[13898]_ , \new_[13902]_ , \new_[13903]_ ,
    \new_[13904]_ , \new_[13907]_ , \new_[13910]_ , \new_[13911]_ ,
    \new_[13914]_ , \new_[13918]_ , \new_[13919]_ , \new_[13920]_ ,
    \new_[13923]_ , \new_[13926]_ , \new_[13927]_ , \new_[13930]_ ,
    \new_[13934]_ , \new_[13935]_ , \new_[13936]_ , \new_[13939]_ ,
    \new_[13942]_ , \new_[13943]_ , \new_[13946]_ , \new_[13950]_ ,
    \new_[13951]_ , \new_[13952]_ , \new_[13955]_ , \new_[13958]_ ,
    \new_[13959]_ , \new_[13962]_ , \new_[13966]_ , \new_[13967]_ ,
    \new_[13968]_ , \new_[13971]_ , \new_[13974]_ , \new_[13975]_ ,
    \new_[13978]_ , \new_[13982]_ , \new_[13983]_ , \new_[13984]_ ,
    \new_[13987]_ , \new_[13990]_ , \new_[13991]_ , \new_[13994]_ ,
    \new_[13998]_ , \new_[13999]_ , \new_[14000]_ , \new_[14003]_ ,
    \new_[14006]_ , \new_[14007]_ , \new_[14010]_ , \new_[14014]_ ,
    \new_[14015]_ , \new_[14016]_ , \new_[14019]_ , \new_[14022]_ ,
    \new_[14023]_ , \new_[14026]_ , \new_[14030]_ , \new_[14031]_ ,
    \new_[14032]_ , \new_[14035]_ , \new_[14038]_ , \new_[14039]_ ,
    \new_[14042]_ , \new_[14046]_ , \new_[14047]_ , \new_[14048]_ ,
    \new_[14051]_ , \new_[14054]_ , \new_[14055]_ , \new_[14058]_ ,
    \new_[14062]_ , \new_[14063]_ , \new_[14064]_ , \new_[14067]_ ,
    \new_[14070]_ , \new_[14071]_ , \new_[14074]_ , \new_[14078]_ ,
    \new_[14079]_ , \new_[14080]_ , \new_[14083]_ , \new_[14086]_ ,
    \new_[14087]_ , \new_[14090]_ , \new_[14094]_ , \new_[14095]_ ,
    \new_[14096]_ , \new_[14099]_ , \new_[14102]_ , \new_[14103]_ ,
    \new_[14106]_ , \new_[14110]_ , \new_[14111]_ , \new_[14112]_ ,
    \new_[14115]_ , \new_[14118]_ , \new_[14119]_ , \new_[14122]_ ,
    \new_[14126]_ , \new_[14127]_ , \new_[14128]_ , \new_[14131]_ ,
    \new_[14134]_ , \new_[14135]_ , \new_[14138]_ , \new_[14142]_ ,
    \new_[14143]_ , \new_[14144]_ , \new_[14147]_ , \new_[14150]_ ,
    \new_[14151]_ , \new_[14154]_ , \new_[14158]_ , \new_[14159]_ ,
    \new_[14160]_ , \new_[14163]_ , \new_[14166]_ , \new_[14167]_ ,
    \new_[14170]_ , \new_[14174]_ , \new_[14175]_ , \new_[14176]_ ,
    \new_[14179]_ , \new_[14182]_ , \new_[14183]_ , \new_[14186]_ ,
    \new_[14190]_ , \new_[14191]_ , \new_[14192]_ , \new_[14195]_ ,
    \new_[14198]_ , \new_[14199]_ , \new_[14202]_ , \new_[14206]_ ,
    \new_[14207]_ , \new_[14208]_ , \new_[14211]_ , \new_[14214]_ ,
    \new_[14215]_ , \new_[14218]_ , \new_[14222]_ , \new_[14223]_ ,
    \new_[14224]_ , \new_[14227]_ , \new_[14230]_ , \new_[14231]_ ,
    \new_[14234]_ , \new_[14238]_ , \new_[14239]_ , \new_[14240]_ ,
    \new_[14243]_ , \new_[14246]_ , \new_[14247]_ , \new_[14250]_ ,
    \new_[14254]_ , \new_[14255]_ , \new_[14256]_ , \new_[14259]_ ,
    \new_[14262]_ , \new_[14263]_ , \new_[14266]_ , \new_[14270]_ ,
    \new_[14271]_ , \new_[14272]_ , \new_[14275]_ , \new_[14278]_ ,
    \new_[14279]_ , \new_[14282]_ , \new_[14286]_ , \new_[14287]_ ,
    \new_[14288]_ , \new_[14291]_ , \new_[14294]_ , \new_[14295]_ ,
    \new_[14298]_ , \new_[14302]_ , \new_[14303]_ , \new_[14304]_ ,
    \new_[14307]_ , \new_[14310]_ , \new_[14311]_ , \new_[14314]_ ,
    \new_[14318]_ , \new_[14319]_ , \new_[14320]_ , \new_[14323]_ ,
    \new_[14326]_ , \new_[14327]_ , \new_[14330]_ , \new_[14334]_ ,
    \new_[14335]_ , \new_[14336]_ , \new_[14339]_ , \new_[14342]_ ,
    \new_[14343]_ , \new_[14346]_ , \new_[14350]_ , \new_[14351]_ ,
    \new_[14352]_ , \new_[14355]_ , \new_[14358]_ , \new_[14359]_ ,
    \new_[14362]_ , \new_[14366]_ , \new_[14367]_ , \new_[14368]_ ,
    \new_[14371]_ , \new_[14374]_ , \new_[14375]_ , \new_[14378]_ ,
    \new_[14382]_ , \new_[14383]_ , \new_[14384]_ , \new_[14387]_ ,
    \new_[14390]_ , \new_[14391]_ , \new_[14394]_ , \new_[14398]_ ,
    \new_[14399]_ , \new_[14400]_ , \new_[14403]_ , \new_[14406]_ ,
    \new_[14407]_ , \new_[14410]_ , \new_[14414]_ , \new_[14415]_ ,
    \new_[14416]_ , \new_[14419]_ , \new_[14422]_ , \new_[14423]_ ,
    \new_[14426]_ , \new_[14430]_ , \new_[14431]_ , \new_[14432]_ ,
    \new_[14435]_ , \new_[14438]_ , \new_[14439]_ , \new_[14442]_ ,
    \new_[14446]_ , \new_[14447]_ , \new_[14448]_ , \new_[14451]_ ,
    \new_[14454]_ , \new_[14455]_ , \new_[14458]_ , \new_[14462]_ ,
    \new_[14463]_ , \new_[14464]_ , \new_[14467]_ , \new_[14470]_ ,
    \new_[14471]_ , \new_[14474]_ , \new_[14478]_ , \new_[14479]_ ,
    \new_[14480]_ , \new_[14483]_ , \new_[14486]_ , \new_[14487]_ ,
    \new_[14490]_ , \new_[14494]_ , \new_[14495]_ , \new_[14496]_ ,
    \new_[14499]_ , \new_[14502]_ , \new_[14503]_ , \new_[14506]_ ,
    \new_[14510]_ , \new_[14511]_ , \new_[14512]_ , \new_[14515]_ ,
    \new_[14518]_ , \new_[14519]_ , \new_[14522]_ , \new_[14526]_ ,
    \new_[14527]_ , \new_[14528]_ , \new_[14531]_ , \new_[14534]_ ,
    \new_[14535]_ , \new_[14538]_ , \new_[14542]_ , \new_[14543]_ ,
    \new_[14544]_ , \new_[14547]_ , \new_[14550]_ , \new_[14551]_ ,
    \new_[14554]_ , \new_[14558]_ , \new_[14559]_ , \new_[14560]_ ,
    \new_[14563]_ , \new_[14566]_ , \new_[14567]_ , \new_[14570]_ ,
    \new_[14574]_ , \new_[14575]_ , \new_[14576]_ , \new_[14579]_ ,
    \new_[14582]_ , \new_[14583]_ , \new_[14586]_ , \new_[14590]_ ,
    \new_[14591]_ , \new_[14592]_ , \new_[14595]_ , \new_[14598]_ ,
    \new_[14599]_ , \new_[14602]_ , \new_[14606]_ , \new_[14607]_ ,
    \new_[14608]_ , \new_[14611]_ , \new_[14614]_ , \new_[14615]_ ,
    \new_[14618]_ , \new_[14622]_ , \new_[14623]_ , \new_[14624]_ ,
    \new_[14627]_ , \new_[14630]_ , \new_[14631]_ , \new_[14634]_ ,
    \new_[14638]_ , \new_[14639]_ , \new_[14640]_ , \new_[14643]_ ,
    \new_[14646]_ , \new_[14647]_ , \new_[14650]_ , \new_[14654]_ ,
    \new_[14655]_ , \new_[14656]_ , \new_[14659]_ , \new_[14662]_ ,
    \new_[14663]_ , \new_[14666]_ , \new_[14670]_ , \new_[14671]_ ,
    \new_[14672]_ , \new_[14675]_ , \new_[14678]_ , \new_[14679]_ ,
    \new_[14682]_ , \new_[14686]_ , \new_[14687]_ , \new_[14688]_ ,
    \new_[14691]_ , \new_[14694]_ , \new_[14695]_ , \new_[14698]_ ,
    \new_[14702]_ , \new_[14703]_ , \new_[14704]_ , \new_[14707]_ ,
    \new_[14710]_ , \new_[14711]_ , \new_[14714]_ , \new_[14718]_ ,
    \new_[14719]_ , \new_[14720]_ , \new_[14723]_ , \new_[14726]_ ,
    \new_[14727]_ , \new_[14730]_ , \new_[14734]_ , \new_[14735]_ ,
    \new_[14736]_ , \new_[14739]_ , \new_[14742]_ , \new_[14743]_ ,
    \new_[14746]_ , \new_[14750]_ , \new_[14751]_ , \new_[14752]_ ,
    \new_[14755]_ , \new_[14758]_ , \new_[14759]_ , \new_[14762]_ ,
    \new_[14766]_ , \new_[14767]_ , \new_[14768]_ , \new_[14771]_ ,
    \new_[14774]_ , \new_[14775]_ , \new_[14778]_ , \new_[14782]_ ,
    \new_[14783]_ , \new_[14784]_ , \new_[14787]_ , \new_[14790]_ ,
    \new_[14791]_ , \new_[14794]_ , \new_[14798]_ , \new_[14799]_ ,
    \new_[14800]_ , \new_[14803]_ , \new_[14806]_ , \new_[14807]_ ,
    \new_[14810]_ , \new_[14814]_ , \new_[14815]_ , \new_[14816]_ ,
    \new_[14819]_ , \new_[14822]_ , \new_[14823]_ , \new_[14826]_ ,
    \new_[14830]_ , \new_[14831]_ , \new_[14832]_ , \new_[14835]_ ,
    \new_[14838]_ , \new_[14839]_ , \new_[14842]_ , \new_[14846]_ ,
    \new_[14847]_ , \new_[14848]_ , \new_[14851]_ , \new_[14854]_ ,
    \new_[14855]_ , \new_[14858]_ , \new_[14862]_ , \new_[14863]_ ,
    \new_[14864]_ , \new_[14867]_ , \new_[14870]_ , \new_[14871]_ ,
    \new_[14874]_ , \new_[14878]_ , \new_[14879]_ , \new_[14880]_ ,
    \new_[14883]_ , \new_[14886]_ , \new_[14887]_ , \new_[14890]_ ,
    \new_[14894]_ , \new_[14895]_ , \new_[14896]_ , \new_[14899]_ ,
    \new_[14902]_ , \new_[14903]_ , \new_[14906]_ , \new_[14910]_ ,
    \new_[14911]_ , \new_[14912]_ , \new_[14915]_ , \new_[14918]_ ,
    \new_[14919]_ , \new_[14922]_ , \new_[14926]_ , \new_[14927]_ ,
    \new_[14928]_ , \new_[14931]_ , \new_[14934]_ , \new_[14935]_ ,
    \new_[14938]_ , \new_[14942]_ , \new_[14943]_ , \new_[14944]_ ,
    \new_[14947]_ , \new_[14950]_ , \new_[14951]_ , \new_[14954]_ ,
    \new_[14958]_ , \new_[14959]_ , \new_[14960]_ , \new_[14963]_ ,
    \new_[14966]_ , \new_[14967]_ , \new_[14970]_ , \new_[14974]_ ,
    \new_[14975]_ , \new_[14976]_ , \new_[14979]_ , \new_[14982]_ ,
    \new_[14983]_ , \new_[14986]_ , \new_[14990]_ , \new_[14991]_ ,
    \new_[14992]_ , \new_[14995]_ , \new_[14998]_ , \new_[14999]_ ,
    \new_[15002]_ , \new_[15006]_ , \new_[15007]_ , \new_[15008]_ ,
    \new_[15011]_ , \new_[15014]_ , \new_[15015]_ , \new_[15018]_ ,
    \new_[15022]_ , \new_[15023]_ , \new_[15024]_ , \new_[15027]_ ,
    \new_[15030]_ , \new_[15031]_ , \new_[15034]_ , \new_[15038]_ ,
    \new_[15039]_ , \new_[15040]_ , \new_[15043]_ , \new_[15046]_ ,
    \new_[15047]_ , \new_[15050]_ , \new_[15054]_ , \new_[15055]_ ,
    \new_[15056]_ , \new_[15059]_ , \new_[15062]_ , \new_[15063]_ ,
    \new_[15066]_ , \new_[15070]_ , \new_[15071]_ , \new_[15072]_ ,
    \new_[15075]_ , \new_[15078]_ , \new_[15079]_ , \new_[15082]_ ,
    \new_[15086]_ , \new_[15087]_ , \new_[15088]_ , \new_[15091]_ ,
    \new_[15094]_ , \new_[15095]_ , \new_[15098]_ , \new_[15102]_ ,
    \new_[15103]_ , \new_[15104]_ , \new_[15107]_ , \new_[15110]_ ,
    \new_[15111]_ , \new_[15114]_ , \new_[15118]_ , \new_[15119]_ ,
    \new_[15120]_ , \new_[15123]_ , \new_[15126]_ , \new_[15127]_ ,
    \new_[15130]_ , \new_[15134]_ , \new_[15135]_ , \new_[15136]_ ,
    \new_[15139]_ , \new_[15142]_ , \new_[15143]_ , \new_[15146]_ ,
    \new_[15150]_ , \new_[15151]_ , \new_[15152]_ , \new_[15155]_ ,
    \new_[15158]_ , \new_[15159]_ , \new_[15162]_ , \new_[15166]_ ,
    \new_[15167]_ , \new_[15168]_ , \new_[15171]_ , \new_[15174]_ ,
    \new_[15175]_ , \new_[15178]_ , \new_[15182]_ , \new_[15183]_ ,
    \new_[15184]_ , \new_[15187]_ , \new_[15190]_ , \new_[15191]_ ,
    \new_[15194]_ , \new_[15198]_ , \new_[15199]_ , \new_[15200]_ ,
    \new_[15203]_ , \new_[15206]_ , \new_[15207]_ , \new_[15210]_ ,
    \new_[15214]_ , \new_[15215]_ , \new_[15216]_ , \new_[15219]_ ,
    \new_[15222]_ , \new_[15223]_ , \new_[15226]_ , \new_[15230]_ ,
    \new_[15231]_ , \new_[15232]_ , \new_[15235]_ , \new_[15239]_ ,
    \new_[15240]_ , \new_[15241]_ , \new_[15244]_ , \new_[15248]_ ,
    \new_[15249]_ , \new_[15250]_ , \new_[15253]_ , \new_[15257]_ ,
    \new_[15258]_ , \new_[15259]_ , \new_[15262]_ , \new_[15266]_ ,
    \new_[15267]_ , \new_[15268]_ , \new_[15271]_ , \new_[15275]_ ,
    \new_[15276]_ , \new_[15277]_ , \new_[15280]_ , \new_[15284]_ ,
    \new_[15285]_ , \new_[15286]_ , \new_[15289]_ , \new_[15293]_ ,
    \new_[15294]_ , \new_[15295]_ , \new_[15298]_ , \new_[15302]_ ,
    \new_[15303]_ , \new_[15304]_ , \new_[15307]_ , \new_[15311]_ ,
    \new_[15312]_ , \new_[15313]_ , \new_[15316]_ , \new_[15320]_ ,
    \new_[15321]_ , \new_[15322]_ , \new_[15325]_ , \new_[15329]_ ,
    \new_[15330]_ , \new_[15331]_ , \new_[15334]_ , \new_[15338]_ ,
    \new_[15339]_ , \new_[15340]_ , \new_[15343]_ , \new_[15347]_ ,
    \new_[15348]_ , \new_[15349]_ , \new_[15352]_ , \new_[15356]_ ,
    \new_[15357]_ , \new_[15358]_ , \new_[15361]_ , \new_[15365]_ ,
    \new_[15366]_ , \new_[15367]_ , \new_[15370]_ , \new_[15374]_ ,
    \new_[15375]_ , \new_[15376]_ , \new_[15379]_ , \new_[15383]_ ,
    \new_[15384]_ , \new_[15385]_ , \new_[15388]_ , \new_[15392]_ ,
    \new_[15393]_ , \new_[15394]_ , \new_[15397]_ , \new_[15401]_ ,
    \new_[15402]_ , \new_[15403]_ , \new_[15406]_ , \new_[15410]_ ,
    \new_[15411]_ , \new_[15412]_ , \new_[15415]_ , \new_[15419]_ ,
    \new_[15420]_ , \new_[15421]_ , \new_[15424]_ , \new_[15428]_ ,
    \new_[15429]_ , \new_[15430]_ , \new_[15433]_ , \new_[15437]_ ,
    \new_[15438]_ , \new_[15439]_ , \new_[15442]_ , \new_[15446]_ ,
    \new_[15447]_ , \new_[15448]_ , \new_[15451]_ , \new_[15455]_ ,
    \new_[15456]_ , \new_[15457]_ , \new_[15460]_ , \new_[15464]_ ,
    \new_[15465]_ , \new_[15466]_ , \new_[15469]_ , \new_[15473]_ ,
    \new_[15474]_ , \new_[15475]_ , \new_[15478]_ , \new_[15482]_ ,
    \new_[15483]_ , \new_[15484]_ , \new_[15487]_ , \new_[15491]_ ,
    \new_[15492]_ , \new_[15493]_ , \new_[15496]_ , \new_[15500]_ ,
    \new_[15501]_ , \new_[15502]_ , \new_[15505]_ , \new_[15509]_ ,
    \new_[15510]_ , \new_[15511]_ , \new_[15514]_ , \new_[15518]_ ,
    \new_[15519]_ , \new_[15520]_ , \new_[15523]_ , \new_[15527]_ ,
    \new_[15528]_ , \new_[15529]_ , \new_[15532]_ , \new_[15536]_ ,
    \new_[15537]_ , \new_[15538]_ , \new_[15541]_ , \new_[15545]_ ,
    \new_[15546]_ , \new_[15547]_ , \new_[15550]_ , \new_[15554]_ ,
    \new_[15555]_ , \new_[15556]_ , \new_[15559]_ , \new_[15563]_ ,
    \new_[15564]_ , \new_[15565]_ , \new_[15568]_ , \new_[15572]_ ,
    \new_[15573]_ , \new_[15574]_ , \new_[15577]_ , \new_[15581]_ ,
    \new_[15582]_ , \new_[15583]_ , \new_[15586]_ , \new_[15590]_ ,
    \new_[15591]_ , \new_[15592]_ , \new_[15595]_ , \new_[15599]_ ,
    \new_[15600]_ , \new_[15601]_ , \new_[15604]_ , \new_[15608]_ ,
    \new_[15609]_ , \new_[15610]_ , \new_[15613]_ , \new_[15617]_ ,
    \new_[15618]_ , \new_[15619]_ , \new_[15622]_ , \new_[15626]_ ,
    \new_[15627]_ , \new_[15628]_ , \new_[15631]_ , \new_[15635]_ ,
    \new_[15636]_ , \new_[15637]_ , \new_[15640]_ , \new_[15644]_ ,
    \new_[15645]_ , \new_[15646]_ , \new_[15649]_ , \new_[15653]_ ,
    \new_[15654]_ , \new_[15655]_ , \new_[15658]_ , \new_[15662]_ ,
    \new_[15663]_ , \new_[15664]_ , \new_[15667]_ , \new_[15671]_ ,
    \new_[15672]_ , \new_[15673]_ , \new_[15676]_ , \new_[15680]_ ,
    \new_[15681]_ , \new_[15682]_ , \new_[15685]_ , \new_[15689]_ ,
    \new_[15690]_ , \new_[15691]_ , \new_[15694]_ , \new_[15698]_ ,
    \new_[15699]_ , \new_[15700]_ , \new_[15703]_ , \new_[15707]_ ,
    \new_[15708]_ , \new_[15709]_ , \new_[15712]_ , \new_[15716]_ ,
    \new_[15717]_ , \new_[15718]_ , \new_[15721]_ , \new_[15725]_ ,
    \new_[15726]_ , \new_[15727]_ , \new_[15730]_ , \new_[15734]_ ,
    \new_[15735]_ , \new_[15736]_ , \new_[15739]_ , \new_[15743]_ ,
    \new_[15744]_ , \new_[15745]_ , \new_[15748]_ , \new_[15752]_ ,
    \new_[15753]_ , \new_[15754]_ , \new_[15757]_ , \new_[15761]_ ,
    \new_[15762]_ , \new_[15763]_ , \new_[15766]_ , \new_[15770]_ ,
    \new_[15771]_ , \new_[15772]_ , \new_[15775]_ , \new_[15779]_ ,
    \new_[15780]_ , \new_[15781]_ , \new_[15784]_ , \new_[15788]_ ,
    \new_[15789]_ , \new_[15790]_ , \new_[15793]_ , \new_[15797]_ ,
    \new_[15798]_ , \new_[15799]_ , \new_[15802]_ , \new_[15806]_ ,
    \new_[15807]_ , \new_[15808]_ , \new_[15811]_ , \new_[15815]_ ,
    \new_[15816]_ , \new_[15817]_ , \new_[15820]_ , \new_[15824]_ ,
    \new_[15825]_ , \new_[15826]_ , \new_[15829]_ , \new_[15833]_ ,
    \new_[15834]_ , \new_[15835]_ , \new_[15838]_ , \new_[15842]_ ,
    \new_[15843]_ , \new_[15844]_ , \new_[15847]_ , \new_[15851]_ ,
    \new_[15852]_ , \new_[15853]_ , \new_[15856]_ , \new_[15860]_ ,
    \new_[15861]_ , \new_[15862]_ , \new_[15865]_ , \new_[15869]_ ,
    \new_[15870]_ , \new_[15871]_ , \new_[15874]_ , \new_[15878]_ ,
    \new_[15879]_ , \new_[15880]_ , \new_[15883]_ , \new_[15887]_ ,
    \new_[15888]_ , \new_[15889]_ , \new_[15892]_ , \new_[15896]_ ,
    \new_[15897]_ , \new_[15898]_ , \new_[15901]_ , \new_[15905]_ ,
    \new_[15906]_ , \new_[15907]_ , \new_[15910]_ , \new_[15914]_ ,
    \new_[15915]_ , \new_[15916]_ , \new_[15919]_ , \new_[15923]_ ,
    \new_[15924]_ , \new_[15925]_ , \new_[15928]_ , \new_[15932]_ ,
    \new_[15933]_ , \new_[15934]_ , \new_[15937]_ , \new_[15941]_ ,
    \new_[15942]_ , \new_[15943]_ , \new_[15946]_ , \new_[15950]_ ,
    \new_[15951]_ , \new_[15952]_ , \new_[15955]_ , \new_[15959]_ ,
    \new_[15960]_ , \new_[15961]_ , \new_[15964]_ , \new_[15968]_ ,
    \new_[15969]_ , \new_[15970]_ , \new_[15973]_ , \new_[15977]_ ,
    \new_[15978]_ , \new_[15979]_ , \new_[15982]_ , \new_[15986]_ ,
    \new_[15987]_ , \new_[15988]_ , \new_[15991]_ , \new_[15995]_ ,
    \new_[15996]_ , \new_[15997]_ , \new_[16000]_ , \new_[16004]_ ,
    \new_[16005]_ , \new_[16006]_ , \new_[16009]_ , \new_[16013]_ ,
    \new_[16014]_ , \new_[16015]_ , \new_[16018]_ , \new_[16022]_ ,
    \new_[16023]_ , \new_[16024]_ , \new_[16027]_ , \new_[16031]_ ,
    \new_[16032]_ , \new_[16033]_ , \new_[16036]_ , \new_[16040]_ ,
    \new_[16041]_ , \new_[16042]_ , \new_[16045]_ , \new_[16049]_ ,
    \new_[16050]_ , \new_[16051]_ , \new_[16054]_ , \new_[16058]_ ,
    \new_[16059]_ , \new_[16060]_ , \new_[16063]_ , \new_[16067]_ ,
    \new_[16068]_ , \new_[16069]_ , \new_[16072]_ , \new_[16076]_ ,
    \new_[16077]_ , \new_[16078]_ , \new_[16081]_ , \new_[16085]_ ,
    \new_[16086]_ , \new_[16087]_ , \new_[16090]_ , \new_[16094]_ ,
    \new_[16095]_ , \new_[16096]_ , \new_[16099]_ , \new_[16103]_ ,
    \new_[16104]_ , \new_[16105]_ , \new_[16108]_ , \new_[16112]_ ,
    \new_[16113]_ , \new_[16114]_ , \new_[16117]_ , \new_[16121]_ ,
    \new_[16122]_ , \new_[16123]_ , \new_[16126]_ , \new_[16130]_ ,
    \new_[16131]_ , \new_[16132]_ , \new_[16135]_ , \new_[16139]_ ,
    \new_[16140]_ , \new_[16141]_ , \new_[16144]_ , \new_[16148]_ ,
    \new_[16149]_ , \new_[16150]_ , \new_[16153]_ , \new_[16157]_ ,
    \new_[16158]_ , \new_[16159]_ , \new_[16162]_ , \new_[16166]_ ,
    \new_[16167]_ , \new_[16168]_ , \new_[16171]_ , \new_[16175]_ ,
    \new_[16176]_ , \new_[16177]_ , \new_[16180]_ , \new_[16184]_ ,
    \new_[16185]_ , \new_[16186]_ , \new_[16189]_ , \new_[16193]_ ,
    \new_[16194]_ , \new_[16195]_ , \new_[16198]_ , \new_[16202]_ ,
    \new_[16203]_ , \new_[16204]_ , \new_[16207]_ , \new_[16211]_ ,
    \new_[16212]_ , \new_[16213]_ , \new_[16216]_ , \new_[16220]_ ,
    \new_[16221]_ , \new_[16222]_ , \new_[16225]_ , \new_[16229]_ ,
    \new_[16230]_ , \new_[16231]_ , \new_[16234]_ , \new_[16238]_ ,
    \new_[16239]_ , \new_[16240]_ , \new_[16243]_ , \new_[16247]_ ,
    \new_[16248]_ , \new_[16249]_ , \new_[16252]_ , \new_[16256]_ ,
    \new_[16257]_ , \new_[16258]_ , \new_[16261]_ , \new_[16265]_ ,
    \new_[16266]_ , \new_[16267]_ , \new_[16270]_ , \new_[16274]_ ,
    \new_[16275]_ , \new_[16276]_ , \new_[16279]_ , \new_[16283]_ ,
    \new_[16284]_ , \new_[16285]_ , \new_[16288]_ , \new_[16292]_ ,
    \new_[16293]_ , \new_[16294]_ , \new_[16297]_ , \new_[16301]_ ,
    \new_[16302]_ , \new_[16303]_ , \new_[16306]_ , \new_[16310]_ ,
    \new_[16311]_ , \new_[16312]_ , \new_[16315]_ , \new_[16319]_ ,
    \new_[16320]_ , \new_[16321]_ , \new_[16324]_ , \new_[16328]_ ,
    \new_[16329]_ , \new_[16330]_ , \new_[16333]_ , \new_[16337]_ ,
    \new_[16338]_ , \new_[16339]_ , \new_[16342]_ , \new_[16346]_ ,
    \new_[16347]_ , \new_[16348]_ , \new_[16351]_ , \new_[16355]_ ,
    \new_[16356]_ , \new_[16357]_ , \new_[16360]_ , \new_[16364]_ ,
    \new_[16365]_ , \new_[16366]_ , \new_[16369]_ , \new_[16373]_ ,
    \new_[16374]_ , \new_[16375]_ , \new_[16378]_ , \new_[16382]_ ,
    \new_[16383]_ , \new_[16384]_ , \new_[16387]_ , \new_[16391]_ ,
    \new_[16392]_ , \new_[16393]_ , \new_[16396]_ , \new_[16400]_ ,
    \new_[16401]_ , \new_[16402]_ , \new_[16405]_ , \new_[16409]_ ,
    \new_[16410]_ , \new_[16411]_ , \new_[16414]_ , \new_[16418]_ ,
    \new_[16419]_ , \new_[16420]_ , \new_[16423]_ , \new_[16427]_ ,
    \new_[16428]_ , \new_[16429]_ , \new_[16432]_ , \new_[16436]_ ,
    \new_[16437]_ , \new_[16438]_ , \new_[16441]_ , \new_[16445]_ ,
    \new_[16446]_ , \new_[16447]_ , \new_[16450]_ , \new_[16454]_ ,
    \new_[16455]_ , \new_[16456]_ , \new_[16459]_ , \new_[16463]_ ,
    \new_[16464]_ , \new_[16465]_ , \new_[16468]_ , \new_[16472]_ ,
    \new_[16473]_ , \new_[16474]_ , \new_[16477]_ , \new_[16481]_ ,
    \new_[16482]_ , \new_[16483]_ , \new_[16486]_ , \new_[16490]_ ,
    \new_[16491]_ , \new_[16492]_ , \new_[16495]_ , \new_[16499]_ ,
    \new_[16500]_ , \new_[16501]_ , \new_[16504]_ , \new_[16508]_ ,
    \new_[16509]_ , \new_[16510]_ , \new_[16513]_ , \new_[16517]_ ,
    \new_[16518]_ , \new_[16519]_ , \new_[16522]_ , \new_[16526]_ ,
    \new_[16527]_ , \new_[16528]_ , \new_[16531]_ , \new_[16535]_ ,
    \new_[16536]_ , \new_[16537]_ , \new_[16540]_ , \new_[16544]_ ,
    \new_[16545]_ , \new_[16546]_ , \new_[16549]_ , \new_[16553]_ ,
    \new_[16554]_ , \new_[16555]_ , \new_[16558]_ , \new_[16562]_ ,
    \new_[16563]_ , \new_[16564]_ , \new_[16567]_ , \new_[16571]_ ,
    \new_[16572]_ , \new_[16573]_ , \new_[16576]_ , \new_[16580]_ ,
    \new_[16581]_ , \new_[16582]_ , \new_[16585]_ , \new_[16589]_ ,
    \new_[16590]_ , \new_[16591]_ , \new_[16594]_ , \new_[16598]_ ,
    \new_[16599]_ , \new_[16600]_ , \new_[16603]_ , \new_[16607]_ ,
    \new_[16608]_ , \new_[16609]_ , \new_[16612]_ , \new_[16616]_ ,
    \new_[16617]_ , \new_[16618]_ , \new_[16621]_ , \new_[16625]_ ,
    \new_[16626]_ , \new_[16627]_ , \new_[16630]_ , \new_[16634]_ ,
    \new_[16635]_ , \new_[16636]_ , \new_[16639]_ , \new_[16643]_ ,
    \new_[16644]_ , \new_[16645]_ , \new_[16648]_ , \new_[16652]_ ,
    \new_[16653]_ , \new_[16654]_ , \new_[16657]_ , \new_[16661]_ ,
    \new_[16662]_ , \new_[16663]_ , \new_[16666]_ , \new_[16670]_ ,
    \new_[16671]_ , \new_[16672]_ , \new_[16675]_ , \new_[16679]_ ,
    \new_[16680]_ , \new_[16681]_ , \new_[16684]_ , \new_[16688]_ ,
    \new_[16689]_ , \new_[16690]_ , \new_[16693]_ , \new_[16697]_ ,
    \new_[16698]_ , \new_[16699]_ , \new_[16702]_ , \new_[16706]_ ,
    \new_[16707]_ , \new_[16708]_ , \new_[16711]_ , \new_[16715]_ ,
    \new_[16716]_ , \new_[16717]_ , \new_[16720]_ , \new_[16724]_ ,
    \new_[16725]_ , \new_[16726]_ , \new_[16729]_ , \new_[16733]_ ,
    \new_[16734]_ , \new_[16735]_ , \new_[16738]_ , \new_[16742]_ ,
    \new_[16743]_ , \new_[16744]_ , \new_[16747]_ , \new_[16751]_ ,
    \new_[16752]_ , \new_[16753]_ , \new_[16756]_ , \new_[16760]_ ,
    \new_[16761]_ , \new_[16762]_ , \new_[16765]_ , \new_[16769]_ ,
    \new_[16770]_ , \new_[16771]_ , \new_[16774]_ , \new_[16778]_ ,
    \new_[16779]_ , \new_[16780]_ , \new_[16783]_ , \new_[16787]_ ,
    \new_[16788]_ , \new_[16789]_ , \new_[16792]_ , \new_[16796]_ ,
    \new_[16797]_ , \new_[16798]_ , \new_[16801]_ , \new_[16805]_ ,
    \new_[16806]_ , \new_[16807]_ , \new_[16810]_ , \new_[16814]_ ,
    \new_[16815]_ , \new_[16816]_ , \new_[16819]_ , \new_[16823]_ ,
    \new_[16824]_ , \new_[16825]_ , \new_[16828]_ , \new_[16832]_ ,
    \new_[16833]_ , \new_[16834]_ , \new_[16837]_ , \new_[16841]_ ,
    \new_[16842]_ , \new_[16843]_ , \new_[16846]_ , \new_[16850]_ ,
    \new_[16851]_ , \new_[16852]_ , \new_[16855]_ , \new_[16859]_ ,
    \new_[16860]_ , \new_[16861]_ , \new_[16864]_ , \new_[16868]_ ,
    \new_[16869]_ , \new_[16870]_ , \new_[16873]_ , \new_[16877]_ ,
    \new_[16878]_ , \new_[16879]_ , \new_[16882]_ , \new_[16886]_ ,
    \new_[16887]_ , \new_[16888]_ , \new_[16891]_ , \new_[16895]_ ,
    \new_[16896]_ , \new_[16897]_ , \new_[16900]_ , \new_[16904]_ ,
    \new_[16905]_ , \new_[16906]_ , \new_[16909]_ , \new_[16913]_ ,
    \new_[16914]_ , \new_[16915]_ , \new_[16918]_ , \new_[16922]_ ,
    \new_[16923]_ , \new_[16924]_ , \new_[16927]_ , \new_[16931]_ ,
    \new_[16932]_ , \new_[16933]_ , \new_[16936]_ , \new_[16940]_ ,
    \new_[16941]_ , \new_[16942]_ , \new_[16945]_ , \new_[16949]_ ,
    \new_[16950]_ , \new_[16951]_ , \new_[16954]_ , \new_[16958]_ ,
    \new_[16959]_ , \new_[16960]_ , \new_[16963]_ , \new_[16967]_ ,
    \new_[16968]_ , \new_[16969]_ , \new_[16972]_ , \new_[16976]_ ,
    \new_[16977]_ , \new_[16978]_ , \new_[16981]_ , \new_[16985]_ ,
    \new_[16986]_ , \new_[16987]_ , \new_[16990]_ , \new_[16994]_ ,
    \new_[16995]_ , \new_[16996]_ , \new_[16999]_ , \new_[17003]_ ,
    \new_[17004]_ , \new_[17005]_ , \new_[17008]_ , \new_[17012]_ ,
    \new_[17013]_ , \new_[17014]_ , \new_[17017]_ , \new_[17021]_ ,
    \new_[17022]_ , \new_[17023]_ , \new_[17026]_ , \new_[17030]_ ,
    \new_[17031]_ , \new_[17032]_ , \new_[17035]_ , \new_[17039]_ ,
    \new_[17040]_ , \new_[17041]_ , \new_[17044]_ , \new_[17048]_ ,
    \new_[17049]_ , \new_[17050]_ , \new_[17053]_ , \new_[17057]_ ,
    \new_[17058]_ , \new_[17059]_ , \new_[17062]_ , \new_[17066]_ ,
    \new_[17067]_ , \new_[17068]_ , \new_[17071]_ , \new_[17075]_ ,
    \new_[17076]_ , \new_[17077]_ , \new_[17080]_ , \new_[17084]_ ,
    \new_[17085]_ , \new_[17086]_ , \new_[17089]_ , \new_[17093]_ ,
    \new_[17094]_ , \new_[17095]_ , \new_[17098]_ , \new_[17102]_ ,
    \new_[17103]_ , \new_[17104]_ , \new_[17107]_ , \new_[17111]_ ,
    \new_[17112]_ , \new_[17113]_ , \new_[17116]_ , \new_[17120]_ ,
    \new_[17121]_ , \new_[17122]_ , \new_[17125]_ , \new_[17129]_ ,
    \new_[17130]_ , \new_[17131]_ , \new_[17134]_ , \new_[17138]_ ,
    \new_[17139]_ , \new_[17140]_ , \new_[17143]_ , \new_[17147]_ ,
    \new_[17148]_ , \new_[17149]_ , \new_[17152]_ , \new_[17156]_ ,
    \new_[17157]_ , \new_[17158]_ , \new_[17161]_ , \new_[17165]_ ,
    \new_[17166]_ , \new_[17167]_ , \new_[17170]_ , \new_[17174]_ ,
    \new_[17175]_ , \new_[17176]_ , \new_[17179]_ , \new_[17183]_ ,
    \new_[17184]_ , \new_[17185]_ , \new_[17188]_ , \new_[17192]_ ,
    \new_[17193]_ , \new_[17194]_ , \new_[17197]_ , \new_[17201]_ ,
    \new_[17202]_ , \new_[17203]_ , \new_[17206]_ , \new_[17210]_ ,
    \new_[17211]_ , \new_[17212]_ , \new_[17215]_ , \new_[17219]_ ,
    \new_[17220]_ , \new_[17221]_ , \new_[17224]_ , \new_[17228]_ ,
    \new_[17229]_ , \new_[17230]_ , \new_[17233]_ , \new_[17237]_ ,
    \new_[17238]_ , \new_[17239]_ , \new_[17242]_ , \new_[17246]_ ,
    \new_[17247]_ , \new_[17248]_ , \new_[17251]_ , \new_[17255]_ ,
    \new_[17256]_ , \new_[17257]_ , \new_[17260]_ , \new_[17264]_ ,
    \new_[17265]_ , \new_[17266]_ , \new_[17269]_ , \new_[17273]_ ,
    \new_[17274]_ , \new_[17275]_ , \new_[17278]_ , \new_[17282]_ ,
    \new_[17283]_ , \new_[17284]_ , \new_[17287]_ , \new_[17291]_ ,
    \new_[17292]_ , \new_[17293]_ , \new_[17296]_ , \new_[17300]_ ,
    \new_[17301]_ , \new_[17302]_ , \new_[17305]_ , \new_[17309]_ ,
    \new_[17310]_ , \new_[17311]_ , \new_[17314]_ , \new_[17318]_ ,
    \new_[17319]_ , \new_[17320]_ , \new_[17323]_ , \new_[17327]_ ,
    \new_[17328]_ , \new_[17329]_ , \new_[17332]_ , \new_[17336]_ ,
    \new_[17337]_ , \new_[17338]_ , \new_[17341]_ , \new_[17345]_ ,
    \new_[17346]_ , \new_[17347]_ , \new_[17350]_ , \new_[17354]_ ,
    \new_[17355]_ , \new_[17356]_ , \new_[17359]_ , \new_[17363]_ ,
    \new_[17364]_ , \new_[17365]_ , \new_[17368]_ , \new_[17372]_ ,
    \new_[17373]_ , \new_[17374]_ , \new_[17377]_ , \new_[17381]_ ,
    \new_[17382]_ , \new_[17383]_ , \new_[17386]_ , \new_[17390]_ ,
    \new_[17391]_ , \new_[17392]_ , \new_[17395]_ , \new_[17399]_ ,
    \new_[17400]_ , \new_[17401]_ , \new_[17404]_ , \new_[17408]_ ,
    \new_[17409]_ , \new_[17410]_ , \new_[17413]_ , \new_[17417]_ ,
    \new_[17418]_ , \new_[17419]_ , \new_[17422]_ , \new_[17426]_ ,
    \new_[17427]_ , \new_[17428]_ , \new_[17431]_ , \new_[17435]_ ,
    \new_[17436]_ , \new_[17437]_ , \new_[17440]_ , \new_[17444]_ ,
    \new_[17445]_ , \new_[17446]_ , \new_[17449]_ , \new_[17453]_ ,
    \new_[17454]_ , \new_[17455]_ , \new_[17458]_ , \new_[17462]_ ,
    \new_[17463]_ , \new_[17464]_ , \new_[17467]_ , \new_[17471]_ ,
    \new_[17472]_ , \new_[17473]_ , \new_[17476]_ , \new_[17480]_ ,
    \new_[17481]_ , \new_[17482]_ , \new_[17485]_ , \new_[17489]_ ,
    \new_[17490]_ , \new_[17491]_ , \new_[17494]_ , \new_[17498]_ ,
    \new_[17499]_ , \new_[17500]_ , \new_[17503]_ , \new_[17507]_ ,
    \new_[17508]_ , \new_[17509]_ , \new_[17512]_ , \new_[17516]_ ,
    \new_[17517]_ , \new_[17518]_ , \new_[17521]_ , \new_[17525]_ ,
    \new_[17526]_ , \new_[17527]_ , \new_[17530]_ , \new_[17534]_ ,
    \new_[17535]_ , \new_[17536]_ , \new_[17539]_ , \new_[17543]_ ,
    \new_[17544]_ , \new_[17545]_ , \new_[17548]_ , \new_[17552]_ ,
    \new_[17553]_ , \new_[17554]_ , \new_[17557]_ , \new_[17561]_ ,
    \new_[17562]_ , \new_[17563]_ , \new_[17566]_ , \new_[17570]_ ,
    \new_[17571]_ , \new_[17572]_ , \new_[17575]_ , \new_[17579]_ ,
    \new_[17580]_ , \new_[17581]_ , \new_[17584]_ , \new_[17588]_ ,
    \new_[17589]_ , \new_[17590]_ , \new_[17593]_ , \new_[17597]_ ,
    \new_[17598]_ , \new_[17599]_ , \new_[17602]_ , \new_[17606]_ ,
    \new_[17607]_ , \new_[17608]_ , \new_[17611]_ , \new_[17615]_ ,
    \new_[17616]_ , \new_[17617]_ , \new_[17620]_ , \new_[17624]_ ,
    \new_[17625]_ , \new_[17626]_ , \new_[17629]_ , \new_[17633]_ ,
    \new_[17634]_ , \new_[17635]_ , \new_[17638]_ , \new_[17642]_ ,
    \new_[17643]_ , \new_[17644]_ , \new_[17647]_ , \new_[17651]_ ,
    \new_[17652]_ , \new_[17653]_ , \new_[17656]_ , \new_[17660]_ ,
    \new_[17661]_ , \new_[17662]_ , \new_[17665]_ , \new_[17669]_ ,
    \new_[17670]_ , \new_[17671]_ , \new_[17674]_ , \new_[17678]_ ,
    \new_[17679]_ , \new_[17680]_ , \new_[17683]_ , \new_[17687]_ ,
    \new_[17688]_ , \new_[17689]_ , \new_[17692]_ , \new_[17696]_ ,
    \new_[17697]_ , \new_[17698]_ , \new_[17701]_ , \new_[17705]_ ,
    \new_[17706]_ , \new_[17707]_ , \new_[17710]_ , \new_[17714]_ ,
    \new_[17715]_ , \new_[17716]_ , \new_[17719]_ , \new_[17723]_ ,
    \new_[17724]_ , \new_[17725]_ , \new_[17728]_ , \new_[17732]_ ,
    \new_[17733]_ , \new_[17734]_ , \new_[17737]_ , \new_[17741]_ ,
    \new_[17742]_ , \new_[17743]_ , \new_[17746]_ , \new_[17750]_ ,
    \new_[17751]_ , \new_[17752]_ , \new_[17755]_ , \new_[17759]_ ,
    \new_[17760]_ , \new_[17761]_ , \new_[17764]_ , \new_[17768]_ ,
    \new_[17769]_ , \new_[17770]_ , \new_[17773]_ , \new_[17777]_ ,
    \new_[17778]_ , \new_[17779]_ , \new_[17782]_ , \new_[17786]_ ,
    \new_[17787]_ , \new_[17788]_ , \new_[17791]_ , \new_[17795]_ ,
    \new_[17796]_ , \new_[17797]_ , \new_[17800]_ , \new_[17804]_ ,
    \new_[17805]_ , \new_[17806]_ , \new_[17809]_ , \new_[17813]_ ,
    \new_[17814]_ , \new_[17815]_ , \new_[17818]_ , \new_[17822]_ ,
    \new_[17823]_ , \new_[17824]_ , \new_[17827]_ , \new_[17831]_ ,
    \new_[17832]_ , \new_[17833]_ , \new_[17836]_ , \new_[17840]_ ,
    \new_[17841]_ , \new_[17842]_ , \new_[17845]_ , \new_[17849]_ ,
    \new_[17850]_ , \new_[17851]_ , \new_[17854]_ , \new_[17858]_ ,
    \new_[17859]_ , \new_[17860]_ , \new_[17863]_ , \new_[17867]_ ,
    \new_[17868]_ , \new_[17869]_ , \new_[17872]_ , \new_[17876]_ ,
    \new_[17877]_ , \new_[17878]_ , \new_[17881]_ , \new_[17885]_ ,
    \new_[17886]_ , \new_[17887]_ , \new_[17890]_ , \new_[17894]_ ,
    \new_[17895]_ , \new_[17896]_ , \new_[17899]_ , \new_[17903]_ ,
    \new_[17904]_ , \new_[17905]_ , \new_[17908]_ , \new_[17912]_ ,
    \new_[17913]_ , \new_[17914]_ , \new_[17917]_ , \new_[17921]_ ,
    \new_[17922]_ , \new_[17923]_ , \new_[17926]_ , \new_[17930]_ ,
    \new_[17931]_ , \new_[17932]_ , \new_[17935]_ , \new_[17939]_ ,
    \new_[17940]_ , \new_[17941]_ , \new_[17944]_ , \new_[17948]_ ,
    \new_[17949]_ , \new_[17950]_ , \new_[17953]_ , \new_[17957]_ ,
    \new_[17958]_ , \new_[17959]_ , \new_[17962]_ , \new_[17966]_ ,
    \new_[17967]_ , \new_[17968]_ , \new_[17971]_ , \new_[17975]_ ,
    \new_[17976]_ , \new_[17977]_ , \new_[17980]_ , \new_[17984]_ ,
    \new_[17985]_ , \new_[17986]_ , \new_[17989]_ , \new_[17993]_ ,
    \new_[17994]_ , \new_[17995]_ , \new_[17998]_ , \new_[18002]_ ,
    \new_[18003]_ , \new_[18004]_ , \new_[18007]_ , \new_[18011]_ ,
    \new_[18012]_ , \new_[18013]_ , \new_[18016]_ , \new_[18020]_ ,
    \new_[18021]_ , \new_[18022]_ , \new_[18025]_ , \new_[18029]_ ,
    \new_[18030]_ , \new_[18031]_ , \new_[18034]_ , \new_[18038]_ ,
    \new_[18039]_ , \new_[18040]_ , \new_[18043]_ , \new_[18047]_ ,
    \new_[18048]_ , \new_[18049]_ , \new_[18052]_ , \new_[18056]_ ,
    \new_[18057]_ , \new_[18058]_ , \new_[18061]_ , \new_[18065]_ ,
    \new_[18066]_ , \new_[18067]_ , \new_[18070]_ , \new_[18074]_ ,
    \new_[18075]_ , \new_[18076]_ , \new_[18079]_ , \new_[18083]_ ,
    \new_[18084]_ , \new_[18085]_ , \new_[18088]_ , \new_[18092]_ ,
    \new_[18093]_ , \new_[18094]_ , \new_[18097]_ , \new_[18101]_ ,
    \new_[18102]_ , \new_[18103]_ , \new_[18106]_ , \new_[18110]_ ,
    \new_[18111]_ , \new_[18112]_ , \new_[18115]_ , \new_[18119]_ ,
    \new_[18120]_ , \new_[18121]_ , \new_[18124]_ , \new_[18128]_ ,
    \new_[18129]_ , \new_[18130]_ , \new_[18133]_ , \new_[18137]_ ,
    \new_[18138]_ , \new_[18139]_ , \new_[18142]_ , \new_[18146]_ ,
    \new_[18147]_ , \new_[18148]_ , \new_[18151]_ , \new_[18155]_ ,
    \new_[18156]_ , \new_[18157]_ , \new_[18160]_ , \new_[18164]_ ,
    \new_[18165]_ , \new_[18166]_ , \new_[18169]_ , \new_[18173]_ ,
    \new_[18174]_ , \new_[18175]_ , \new_[18178]_ , \new_[18182]_ ,
    \new_[18183]_ , \new_[18184]_ , \new_[18187]_ , \new_[18191]_ ,
    \new_[18192]_ , \new_[18193]_ , \new_[18196]_ , \new_[18200]_ ,
    \new_[18201]_ , \new_[18202]_ , \new_[18205]_ , \new_[18209]_ ,
    \new_[18210]_ , \new_[18211]_ , \new_[18214]_ , \new_[18218]_ ,
    \new_[18219]_ , \new_[18220]_ , \new_[18223]_ , \new_[18227]_ ,
    \new_[18228]_ , \new_[18229]_ , \new_[18232]_ , \new_[18236]_ ,
    \new_[18237]_ , \new_[18238]_ , \new_[18241]_ , \new_[18245]_ ,
    \new_[18246]_ , \new_[18247]_ , \new_[18250]_ , \new_[18254]_ ,
    \new_[18255]_ , \new_[18256]_ , \new_[18259]_ , \new_[18263]_ ,
    \new_[18264]_ , \new_[18265]_ , \new_[18268]_ , \new_[18272]_ ,
    \new_[18273]_ , \new_[18274]_ , \new_[18277]_ , \new_[18281]_ ,
    \new_[18282]_ , \new_[18283]_ , \new_[18286]_ , \new_[18290]_ ,
    \new_[18291]_ , \new_[18292]_ , \new_[18295]_ , \new_[18299]_ ,
    \new_[18300]_ , \new_[18301]_ , \new_[18304]_ , \new_[18308]_ ,
    \new_[18309]_ , \new_[18310]_ , \new_[18313]_ , \new_[18317]_ ,
    \new_[18318]_ , \new_[18319]_ , \new_[18322]_ , \new_[18326]_ ,
    \new_[18327]_ , \new_[18328]_ , \new_[18331]_ , \new_[18335]_ ,
    \new_[18336]_ , \new_[18337]_ , \new_[18340]_ , \new_[18344]_ ,
    \new_[18345]_ , \new_[18346]_ , \new_[18349]_ , \new_[18353]_ ,
    \new_[18354]_ , \new_[18355]_ , \new_[18358]_ , \new_[18362]_ ,
    \new_[18363]_ , \new_[18364]_ , \new_[18367]_ , \new_[18371]_ ,
    \new_[18372]_ , \new_[18373]_ , \new_[18376]_ , \new_[18380]_ ,
    \new_[18381]_ , \new_[18382]_ , \new_[18385]_ , \new_[18389]_ ,
    \new_[18390]_ , \new_[18391]_ , \new_[18394]_ , \new_[18398]_ ,
    \new_[18399]_ , \new_[18400]_ , \new_[18403]_ , \new_[18407]_ ,
    \new_[18408]_ , \new_[18409]_ , \new_[18412]_ , \new_[18416]_ ,
    \new_[18417]_ , \new_[18418]_ , \new_[18421]_ , \new_[18425]_ ,
    \new_[18426]_ , \new_[18427]_ , \new_[18430]_ , \new_[18434]_ ,
    \new_[18435]_ , \new_[18436]_ , \new_[18439]_ , \new_[18443]_ ,
    \new_[18444]_ , \new_[18445]_ , \new_[18448]_ , \new_[18452]_ ,
    \new_[18453]_ , \new_[18454]_ , \new_[18457]_ , \new_[18461]_ ,
    \new_[18462]_ , \new_[18463]_ , \new_[18466]_ , \new_[18470]_ ,
    \new_[18471]_ , \new_[18472]_ , \new_[18475]_ , \new_[18479]_ ,
    \new_[18480]_ , \new_[18481]_ , \new_[18484]_ , \new_[18488]_ ,
    \new_[18489]_ , \new_[18490]_ , \new_[18493]_ , \new_[18497]_ ,
    \new_[18498]_ , \new_[18499]_ , \new_[18502]_ , \new_[18506]_ ,
    \new_[18507]_ , \new_[18508]_ , \new_[18511]_ , \new_[18515]_ ,
    \new_[18516]_ , \new_[18517]_ , \new_[18520]_ , \new_[18524]_ ,
    \new_[18525]_ , \new_[18526]_ , \new_[18529]_ , \new_[18533]_ ,
    \new_[18534]_ , \new_[18535]_ , \new_[18538]_ , \new_[18542]_ ,
    \new_[18543]_ , \new_[18544]_ , \new_[18547]_ , \new_[18551]_ ,
    \new_[18552]_ , \new_[18553]_ , \new_[18556]_ , \new_[18560]_ ,
    \new_[18561]_ , \new_[18562]_ , \new_[18565]_ , \new_[18569]_ ,
    \new_[18570]_ , \new_[18571]_ , \new_[18574]_ , \new_[18578]_ ,
    \new_[18579]_ , \new_[18580]_ , \new_[18583]_ , \new_[18587]_ ,
    \new_[18588]_ , \new_[18589]_ , \new_[18592]_ , \new_[18596]_ ,
    \new_[18597]_ , \new_[18598]_ , \new_[18601]_ , \new_[18605]_ ,
    \new_[18606]_ , \new_[18607]_ , \new_[18610]_ , \new_[18614]_ ,
    \new_[18615]_ , \new_[18616]_ , \new_[18619]_ , \new_[18623]_ ,
    \new_[18624]_ , \new_[18625]_ , \new_[18628]_ , \new_[18632]_ ,
    \new_[18633]_ , \new_[18634]_ , \new_[18637]_ , \new_[18641]_ ,
    \new_[18642]_ , \new_[18643]_ , \new_[18646]_ , \new_[18650]_ ,
    \new_[18651]_ , \new_[18652]_ , \new_[18655]_ , \new_[18659]_ ,
    \new_[18660]_ , \new_[18661]_ , \new_[18664]_ , \new_[18668]_ ,
    \new_[18669]_ , \new_[18670]_ , \new_[18673]_ , \new_[18677]_ ,
    \new_[18678]_ , \new_[18679]_ , \new_[18682]_ , \new_[18686]_ ,
    \new_[18687]_ , \new_[18688]_ , \new_[18691]_ , \new_[18695]_ ,
    \new_[18696]_ , \new_[18697]_ , \new_[18700]_ , \new_[18704]_ ,
    \new_[18705]_ , \new_[18706]_ , \new_[18709]_ , \new_[18713]_ ,
    \new_[18714]_ , \new_[18715]_ , \new_[18718]_ , \new_[18722]_ ,
    \new_[18723]_ , \new_[18724]_ , \new_[18727]_ , \new_[18731]_ ,
    \new_[18732]_ , \new_[18733]_ , \new_[18736]_ , \new_[18740]_ ,
    \new_[18741]_ , \new_[18742]_ , \new_[18745]_ , \new_[18749]_ ,
    \new_[18750]_ , \new_[18751]_ , \new_[18754]_ , \new_[18758]_ ,
    \new_[18759]_ , \new_[18760]_ , \new_[18763]_ , \new_[18767]_ ,
    \new_[18768]_ , \new_[18769]_ , \new_[18772]_ , \new_[18776]_ ,
    \new_[18777]_ , \new_[18778]_ , \new_[18781]_ , \new_[18785]_ ,
    \new_[18786]_ , \new_[18787]_ , \new_[18790]_ , \new_[18794]_ ,
    \new_[18795]_ , \new_[18796]_ , \new_[18799]_ , \new_[18803]_ ,
    \new_[18804]_ , \new_[18805]_ , \new_[18808]_ , \new_[18812]_ ,
    \new_[18813]_ , \new_[18814]_ , \new_[18817]_ , \new_[18821]_ ,
    \new_[18822]_ , \new_[18823]_ , \new_[18826]_ , \new_[18830]_ ,
    \new_[18831]_ , \new_[18832]_ , \new_[18835]_ , \new_[18839]_ ,
    \new_[18840]_ , \new_[18841]_ , \new_[18844]_ , \new_[18848]_ ,
    \new_[18849]_ , \new_[18850]_ , \new_[18853]_ , \new_[18857]_ ,
    \new_[18858]_ , \new_[18859]_ , \new_[18862]_ , \new_[18866]_ ,
    \new_[18867]_ , \new_[18868]_ , \new_[18871]_ , \new_[18875]_ ,
    \new_[18876]_ , \new_[18877]_ , \new_[18880]_ , \new_[18884]_ ,
    \new_[18885]_ , \new_[18886]_ , \new_[18889]_ , \new_[18893]_ ,
    \new_[18894]_ , \new_[18895]_ , \new_[18898]_ , \new_[18902]_ ,
    \new_[18903]_ , \new_[18904]_ , \new_[18907]_ , \new_[18911]_ ,
    \new_[18912]_ , \new_[18913]_ , \new_[18916]_ , \new_[18920]_ ,
    \new_[18921]_ , \new_[18922]_ , \new_[18925]_ , \new_[18929]_ ,
    \new_[18930]_ , \new_[18931]_ , \new_[18934]_ , \new_[18938]_ ,
    \new_[18939]_ , \new_[18940]_ , \new_[18943]_ , \new_[18947]_ ,
    \new_[18948]_ , \new_[18949]_ , \new_[18952]_ , \new_[18956]_ ,
    \new_[18957]_ , \new_[18958]_ , \new_[18961]_ , \new_[18965]_ ,
    \new_[18966]_ , \new_[18967]_ , \new_[18970]_ , \new_[18974]_ ,
    \new_[18975]_ , \new_[18976]_ , \new_[18979]_ , \new_[18983]_ ,
    \new_[18984]_ , \new_[18985]_ , \new_[18988]_ , \new_[18992]_ ,
    \new_[18993]_ , \new_[18994]_ , \new_[18997]_ , \new_[19001]_ ,
    \new_[19002]_ , \new_[19003]_ , \new_[19006]_ , \new_[19010]_ ,
    \new_[19011]_ , \new_[19012]_ , \new_[19015]_ , \new_[19019]_ ,
    \new_[19020]_ , \new_[19021]_ , \new_[19024]_ , \new_[19028]_ ,
    \new_[19029]_ , \new_[19030]_ , \new_[19033]_ , \new_[19037]_ ,
    \new_[19038]_ , \new_[19039]_ , \new_[19042]_ , \new_[19046]_ ,
    \new_[19047]_ , \new_[19048]_ , \new_[19051]_ , \new_[19055]_ ,
    \new_[19056]_ , \new_[19057]_ , \new_[19060]_ , \new_[19064]_ ,
    \new_[19065]_ , \new_[19066]_ , \new_[19069]_ , \new_[19073]_ ,
    \new_[19074]_ , \new_[19075]_ , \new_[19078]_ , \new_[19082]_ ,
    \new_[19083]_ , \new_[19084]_ , \new_[19087]_ , \new_[19091]_ ,
    \new_[19092]_ , \new_[19093]_ , \new_[19096]_ , \new_[19100]_ ,
    \new_[19101]_ , \new_[19102]_ , \new_[19105]_ , \new_[19109]_ ,
    \new_[19110]_ , \new_[19111]_ , \new_[19114]_ , \new_[19118]_ ,
    \new_[19119]_ , \new_[19120]_ , \new_[19123]_ , \new_[19127]_ ,
    \new_[19128]_ , \new_[19129]_ , \new_[19132]_ , \new_[19136]_ ,
    \new_[19137]_ , \new_[19138]_ , \new_[19141]_ , \new_[19145]_ ,
    \new_[19146]_ , \new_[19147]_ , \new_[19150]_ , \new_[19154]_ ,
    \new_[19155]_ , \new_[19156]_ , \new_[19159]_ , \new_[19163]_ ,
    \new_[19164]_ , \new_[19165]_ , \new_[19168]_ , \new_[19172]_ ,
    \new_[19173]_ , \new_[19174]_ , \new_[19177]_ , \new_[19181]_ ,
    \new_[19182]_ , \new_[19183]_ , \new_[19186]_ , \new_[19190]_ ,
    \new_[19191]_ , \new_[19192]_ , \new_[19195]_ , \new_[19199]_ ,
    \new_[19200]_ , \new_[19201]_ , \new_[19204]_ , \new_[19208]_ ,
    \new_[19209]_ , \new_[19210]_ , \new_[19213]_ , \new_[19217]_ ,
    \new_[19218]_ , \new_[19219]_ , \new_[19222]_ , \new_[19226]_ ,
    \new_[19227]_ , \new_[19228]_ , \new_[19231]_ , \new_[19235]_ ,
    \new_[19236]_ , \new_[19237]_ , \new_[19240]_ , \new_[19244]_ ,
    \new_[19245]_ , \new_[19246]_ , \new_[19249]_ , \new_[19253]_ ,
    \new_[19254]_ , \new_[19255]_ , \new_[19258]_ , \new_[19262]_ ,
    \new_[19263]_ , \new_[19264]_ , \new_[19267]_ , \new_[19271]_ ,
    \new_[19272]_ , \new_[19273]_ , \new_[19276]_ , \new_[19280]_ ,
    \new_[19281]_ , \new_[19282]_ , \new_[19285]_ , \new_[19289]_ ,
    \new_[19290]_ , \new_[19291]_ , \new_[19294]_ , \new_[19298]_ ,
    \new_[19299]_ , \new_[19300]_ , \new_[19303]_ , \new_[19307]_ ,
    \new_[19308]_ , \new_[19309]_ , \new_[19312]_ , \new_[19316]_ ,
    \new_[19317]_ , \new_[19318]_ , \new_[19321]_ , \new_[19325]_ ,
    \new_[19326]_ , \new_[19327]_ , \new_[19330]_ , \new_[19334]_ ,
    \new_[19335]_ , \new_[19336]_ , \new_[19339]_ , \new_[19343]_ ,
    \new_[19344]_ , \new_[19345]_ , \new_[19348]_ , \new_[19352]_ ,
    \new_[19353]_ , \new_[19354]_ , \new_[19357]_ , \new_[19361]_ ,
    \new_[19362]_ , \new_[19363]_ , \new_[19366]_ , \new_[19370]_ ,
    \new_[19371]_ , \new_[19372]_ , \new_[19375]_ , \new_[19379]_ ,
    \new_[19380]_ , \new_[19381]_ , \new_[19384]_ , \new_[19388]_ ,
    \new_[19389]_ , \new_[19390]_ , \new_[19393]_ , \new_[19397]_ ,
    \new_[19398]_ , \new_[19399]_ , \new_[19402]_ , \new_[19406]_ ,
    \new_[19407]_ , \new_[19408]_ , \new_[19411]_ , \new_[19415]_ ,
    \new_[19416]_ , \new_[19417]_ , \new_[19420]_ , \new_[19424]_ ,
    \new_[19425]_ , \new_[19426]_ , \new_[19429]_ , \new_[19433]_ ,
    \new_[19434]_ , \new_[19435]_ , \new_[19438]_ , \new_[19442]_ ,
    \new_[19443]_ , \new_[19444]_ , \new_[19447]_ , \new_[19451]_ ,
    \new_[19452]_ , \new_[19453]_ , \new_[19456]_ , \new_[19460]_ ,
    \new_[19461]_ , \new_[19462]_ , \new_[19465]_ , \new_[19469]_ ,
    \new_[19470]_ , \new_[19471]_ , \new_[19474]_ , \new_[19478]_ ,
    \new_[19479]_ , \new_[19480]_ , \new_[19483]_ , \new_[19487]_ ,
    \new_[19488]_ , \new_[19489]_ , \new_[19492]_ , \new_[19496]_ ,
    \new_[19497]_ , \new_[19498]_ , \new_[19501]_ , \new_[19505]_ ,
    \new_[19506]_ , \new_[19507]_ , \new_[19510]_ , \new_[19514]_ ,
    \new_[19515]_ , \new_[19516]_ , \new_[19519]_ , \new_[19523]_ ,
    \new_[19524]_ , \new_[19525]_ , \new_[19528]_ , \new_[19532]_ ,
    \new_[19533]_ , \new_[19534]_ , \new_[19537]_ , \new_[19541]_ ,
    \new_[19542]_ , \new_[19543]_ , \new_[19546]_ , \new_[19550]_ ,
    \new_[19551]_ , \new_[19552]_ , \new_[19555]_ , \new_[19559]_ ,
    \new_[19560]_ , \new_[19561]_ , \new_[19564]_ , \new_[19568]_ ,
    \new_[19569]_ , \new_[19570]_ , \new_[19573]_ , \new_[19577]_ ,
    \new_[19578]_ , \new_[19579]_ , \new_[19582]_ , \new_[19586]_ ,
    \new_[19587]_ , \new_[19588]_ , \new_[19591]_ , \new_[19595]_ ,
    \new_[19596]_ , \new_[19597]_ , \new_[19600]_ , \new_[19604]_ ,
    \new_[19605]_ , \new_[19606]_ , \new_[19609]_ , \new_[19613]_ ,
    \new_[19614]_ , \new_[19615]_ , \new_[19618]_ , \new_[19622]_ ,
    \new_[19623]_ , \new_[19624]_ , \new_[19627]_ , \new_[19631]_ ,
    \new_[19632]_ , \new_[19633]_ , \new_[19636]_ , \new_[19640]_ ,
    \new_[19641]_ , \new_[19642]_ , \new_[19645]_ , \new_[19649]_ ,
    \new_[19650]_ , \new_[19651]_ , \new_[19654]_ , \new_[19658]_ ,
    \new_[19659]_ , \new_[19660]_ , \new_[19663]_ , \new_[19667]_ ,
    \new_[19668]_ , \new_[19669]_ , \new_[19672]_ , \new_[19676]_ ,
    \new_[19677]_ , \new_[19678]_ , \new_[19681]_ , \new_[19685]_ ,
    \new_[19686]_ , \new_[19687]_ , \new_[19690]_ , \new_[19694]_ ,
    \new_[19695]_ , \new_[19696]_ , \new_[19699]_ , \new_[19703]_ ,
    \new_[19704]_ , \new_[19705]_ , \new_[19708]_ , \new_[19712]_ ,
    \new_[19713]_ , \new_[19714]_ , \new_[19717]_ , \new_[19721]_ ,
    \new_[19722]_ , \new_[19723]_ , \new_[19726]_ , \new_[19730]_ ,
    \new_[19731]_ , \new_[19732]_ , \new_[19735]_ , \new_[19739]_ ,
    \new_[19740]_ , \new_[19741]_ , \new_[19744]_ , \new_[19748]_ ,
    \new_[19749]_ , \new_[19750]_ , \new_[19753]_ , \new_[19757]_ ,
    \new_[19758]_ , \new_[19759]_ , \new_[19762]_ , \new_[19766]_ ,
    \new_[19767]_ , \new_[19768]_ , \new_[19771]_ , \new_[19775]_ ,
    \new_[19776]_ , \new_[19777]_ , \new_[19780]_ , \new_[19784]_ ,
    \new_[19785]_ , \new_[19786]_ , \new_[19789]_ , \new_[19793]_ ,
    \new_[19794]_ , \new_[19795]_ , \new_[19798]_ , \new_[19802]_ ,
    \new_[19803]_ , \new_[19804]_ , \new_[19807]_ , \new_[19811]_ ,
    \new_[19812]_ , \new_[19813]_ , \new_[19816]_ , \new_[19820]_ ,
    \new_[19821]_ , \new_[19822]_ , \new_[19825]_ , \new_[19829]_ ,
    \new_[19830]_ , \new_[19831]_ , \new_[19834]_ , \new_[19838]_ ,
    \new_[19839]_ , \new_[19840]_ , \new_[19843]_ , \new_[19847]_ ,
    \new_[19848]_ , \new_[19849]_ , \new_[19852]_ , \new_[19856]_ ,
    \new_[19857]_ , \new_[19858]_ , \new_[19861]_ , \new_[19865]_ ,
    \new_[19866]_ , \new_[19867]_ , \new_[19870]_ , \new_[19874]_ ,
    \new_[19875]_ , \new_[19876]_ , \new_[19879]_ , \new_[19883]_ ,
    \new_[19884]_ , \new_[19885]_ , \new_[19888]_ , \new_[19892]_ ,
    \new_[19893]_ , \new_[19894]_ , \new_[19897]_ , \new_[19901]_ ,
    \new_[19902]_ , \new_[19903]_ , \new_[19906]_ , \new_[19910]_ ,
    \new_[19911]_ , \new_[19912]_ , \new_[19915]_ , \new_[19919]_ ,
    \new_[19920]_ , \new_[19921]_ , \new_[19924]_ , \new_[19928]_ ,
    \new_[19929]_ , \new_[19930]_ , \new_[19933]_ , \new_[19937]_ ,
    \new_[19938]_ , \new_[19939]_ , \new_[19942]_ , \new_[19946]_ ,
    \new_[19947]_ , \new_[19948]_ , \new_[19951]_ , \new_[19955]_ ,
    \new_[19956]_ , \new_[19957]_ , \new_[19960]_ , \new_[19964]_ ,
    \new_[19965]_ , \new_[19966]_ , \new_[19969]_ , \new_[19973]_ ,
    \new_[19974]_ , \new_[19975]_ , \new_[19978]_ , \new_[19982]_ ,
    \new_[19983]_ , \new_[19984]_ , \new_[19987]_ , \new_[19991]_ ,
    \new_[19992]_ , \new_[19993]_ , \new_[19996]_ , \new_[20000]_ ,
    \new_[20001]_ , \new_[20002]_ , \new_[20005]_ , \new_[20009]_ ,
    \new_[20010]_ , \new_[20011]_ , \new_[20014]_ , \new_[20018]_ ,
    \new_[20019]_ , \new_[20020]_ , \new_[20023]_ , \new_[20027]_ ,
    \new_[20028]_ , \new_[20029]_ , \new_[20032]_ , \new_[20036]_ ,
    \new_[20037]_ , \new_[20038]_ , \new_[20041]_ , \new_[20045]_ ,
    \new_[20046]_ , \new_[20047]_ , \new_[20050]_ , \new_[20054]_ ,
    \new_[20055]_ , \new_[20056]_ , \new_[20059]_ , \new_[20063]_ ,
    \new_[20064]_ , \new_[20065]_ , \new_[20068]_ , \new_[20072]_ ,
    \new_[20073]_ , \new_[20074]_ , \new_[20077]_ , \new_[20081]_ ,
    \new_[20082]_ , \new_[20083]_ , \new_[20086]_ , \new_[20090]_ ,
    \new_[20091]_ , \new_[20092]_ , \new_[20095]_ , \new_[20099]_ ,
    \new_[20100]_ , \new_[20101]_ , \new_[20104]_ , \new_[20108]_ ,
    \new_[20109]_ , \new_[20110]_ , \new_[20113]_ , \new_[20117]_ ,
    \new_[20118]_ , \new_[20119]_ , \new_[20122]_ , \new_[20126]_ ,
    \new_[20127]_ , \new_[20128]_ , \new_[20131]_ , \new_[20135]_ ,
    \new_[20136]_ , \new_[20137]_ , \new_[20140]_ , \new_[20144]_ ,
    \new_[20145]_ , \new_[20146]_ , \new_[20149]_ , \new_[20153]_ ,
    \new_[20154]_ , \new_[20155]_ , \new_[20158]_ , \new_[20162]_ ,
    \new_[20163]_ , \new_[20164]_ , \new_[20167]_ , \new_[20171]_ ,
    \new_[20172]_ , \new_[20173]_ , \new_[20176]_ , \new_[20180]_ ,
    \new_[20181]_ , \new_[20182]_ , \new_[20185]_ , \new_[20189]_ ,
    \new_[20190]_ , \new_[20191]_ , \new_[20194]_ , \new_[20198]_ ,
    \new_[20199]_ , \new_[20200]_ , \new_[20203]_ , \new_[20207]_ ,
    \new_[20208]_ , \new_[20209]_ , \new_[20212]_ , \new_[20216]_ ,
    \new_[20217]_ , \new_[20218]_ , \new_[20221]_ , \new_[20225]_ ,
    \new_[20226]_ , \new_[20227]_ , \new_[20230]_ , \new_[20234]_ ,
    \new_[20235]_ , \new_[20236]_ , \new_[20239]_ , \new_[20243]_ ,
    \new_[20244]_ , \new_[20245]_ , \new_[20248]_ , \new_[20252]_ ,
    \new_[20253]_ , \new_[20254]_ , \new_[20257]_ , \new_[20261]_ ,
    \new_[20262]_ , \new_[20263]_ , \new_[20266]_ , \new_[20270]_ ,
    \new_[20271]_ , \new_[20272]_ , \new_[20275]_ , \new_[20279]_ ,
    \new_[20280]_ , \new_[20281]_ , \new_[20284]_ , \new_[20288]_ ,
    \new_[20289]_ , \new_[20290]_ , \new_[20293]_ , \new_[20297]_ ,
    \new_[20298]_ , \new_[20299]_ , \new_[20302]_ , \new_[20306]_ ,
    \new_[20307]_ , \new_[20308]_ , \new_[20311]_ , \new_[20315]_ ,
    \new_[20316]_ , \new_[20317]_ , \new_[20320]_ , \new_[20324]_ ,
    \new_[20325]_ , \new_[20326]_ , \new_[20329]_ , \new_[20333]_ ,
    \new_[20334]_ , \new_[20335]_ , \new_[20338]_ , \new_[20342]_ ,
    \new_[20343]_ , \new_[20344]_ , \new_[20347]_ , \new_[20351]_ ,
    \new_[20352]_ , \new_[20353]_ , \new_[20356]_ , \new_[20360]_ ,
    \new_[20361]_ , \new_[20362]_ , \new_[20365]_ , \new_[20369]_ ,
    \new_[20370]_ , \new_[20371]_ , \new_[20374]_ , \new_[20378]_ ,
    \new_[20379]_ , \new_[20380]_ , \new_[20383]_ , \new_[20387]_ ,
    \new_[20388]_ , \new_[20389]_ , \new_[20392]_ , \new_[20396]_ ,
    \new_[20397]_ , \new_[20398]_ , \new_[20401]_ , \new_[20405]_ ,
    \new_[20406]_ , \new_[20407]_ , \new_[20410]_ , \new_[20414]_ ,
    \new_[20415]_ , \new_[20416]_ , \new_[20419]_ , \new_[20423]_ ,
    \new_[20424]_ , \new_[20425]_ , \new_[20428]_ , \new_[20432]_ ,
    \new_[20433]_ , \new_[20434]_ , \new_[20437]_ , \new_[20441]_ ,
    \new_[20442]_ , \new_[20443]_ , \new_[20446]_ , \new_[20450]_ ,
    \new_[20451]_ , \new_[20452]_ , \new_[20455]_ , \new_[20459]_ ,
    \new_[20460]_ , \new_[20461]_ , \new_[20464]_ , \new_[20468]_ ,
    \new_[20469]_ , \new_[20470]_ , \new_[20473]_ , \new_[20477]_ ,
    \new_[20478]_ , \new_[20479]_ , \new_[20482]_ , \new_[20486]_ ,
    \new_[20487]_ , \new_[20488]_ , \new_[20491]_ , \new_[20495]_ ,
    \new_[20496]_ , \new_[20497]_ , \new_[20500]_ , \new_[20504]_ ,
    \new_[20505]_ , \new_[20506]_ , \new_[20509]_ , \new_[20513]_ ,
    \new_[20514]_ , \new_[20515]_ , \new_[20518]_ , \new_[20522]_ ,
    \new_[20523]_ , \new_[20524]_ , \new_[20527]_ , \new_[20531]_ ,
    \new_[20532]_ , \new_[20533]_ , \new_[20536]_ , \new_[20540]_ ,
    \new_[20541]_ , \new_[20542]_ , \new_[20545]_ , \new_[20549]_ ,
    \new_[20550]_ , \new_[20551]_ , \new_[20554]_ , \new_[20558]_ ,
    \new_[20559]_ , \new_[20560]_ , \new_[20563]_ , \new_[20567]_ ,
    \new_[20568]_ , \new_[20569]_ , \new_[20572]_ , \new_[20576]_ ,
    \new_[20577]_ , \new_[20578]_ , \new_[20581]_ , \new_[20585]_ ,
    \new_[20586]_ , \new_[20587]_ , \new_[20590]_ , \new_[20594]_ ,
    \new_[20595]_ , \new_[20596]_ , \new_[20599]_ , \new_[20603]_ ,
    \new_[20604]_ , \new_[20605]_ , \new_[20608]_ , \new_[20612]_ ,
    \new_[20613]_ , \new_[20614]_ , \new_[20617]_ , \new_[20621]_ ,
    \new_[20622]_ , \new_[20623]_ , \new_[20626]_ , \new_[20630]_ ,
    \new_[20631]_ , \new_[20632]_ , \new_[20635]_ , \new_[20639]_ ,
    \new_[20640]_ , \new_[20641]_ , \new_[20644]_ , \new_[20648]_ ,
    \new_[20649]_ , \new_[20650]_ , \new_[20653]_ , \new_[20657]_ ,
    \new_[20658]_ , \new_[20659]_ , \new_[20662]_ , \new_[20666]_ ,
    \new_[20667]_ , \new_[20668]_ , \new_[20671]_ , \new_[20675]_ ,
    \new_[20676]_ , \new_[20677]_ , \new_[20680]_ , \new_[20684]_ ,
    \new_[20685]_ , \new_[20686]_ , \new_[20689]_ , \new_[20693]_ ,
    \new_[20694]_ , \new_[20695]_ , \new_[20698]_ , \new_[20702]_ ,
    \new_[20703]_ , \new_[20704]_ , \new_[20707]_ , \new_[20711]_ ,
    \new_[20712]_ , \new_[20713]_ , \new_[20716]_ , \new_[20720]_ ,
    \new_[20721]_ , \new_[20722]_ , \new_[20725]_ , \new_[20729]_ ,
    \new_[20730]_ , \new_[20731]_ , \new_[20734]_ , \new_[20738]_ ,
    \new_[20739]_ , \new_[20740]_ , \new_[20743]_ , \new_[20747]_ ,
    \new_[20748]_ , \new_[20749]_ , \new_[20752]_ , \new_[20756]_ ,
    \new_[20757]_ , \new_[20758]_ , \new_[20761]_ , \new_[20765]_ ,
    \new_[20766]_ , \new_[20767]_ , \new_[20770]_ , \new_[20774]_ ,
    \new_[20775]_ , \new_[20776]_ , \new_[20779]_ , \new_[20783]_ ,
    \new_[20784]_ , \new_[20785]_ , \new_[20788]_ , \new_[20792]_ ,
    \new_[20793]_ , \new_[20794]_ , \new_[20797]_ , \new_[20801]_ ,
    \new_[20802]_ , \new_[20803]_ , \new_[20806]_ , \new_[20810]_ ,
    \new_[20811]_ , \new_[20812]_ , \new_[20815]_ , \new_[20819]_ ,
    \new_[20820]_ , \new_[20821]_ , \new_[20824]_ , \new_[20828]_ ,
    \new_[20829]_ , \new_[20830]_ , \new_[20833]_ , \new_[20837]_ ,
    \new_[20838]_ , \new_[20839]_ , \new_[20842]_ , \new_[20846]_ ,
    \new_[20847]_ , \new_[20848]_ , \new_[20851]_ , \new_[20855]_ ,
    \new_[20856]_ , \new_[20857]_ , \new_[20860]_ , \new_[20864]_ ,
    \new_[20865]_ , \new_[20866]_ , \new_[20869]_ , \new_[20873]_ ,
    \new_[20874]_ , \new_[20875]_ , \new_[20878]_ , \new_[20882]_ ,
    \new_[20883]_ , \new_[20884]_ , \new_[20887]_ , \new_[20891]_ ,
    \new_[20892]_ , \new_[20893]_ , \new_[20896]_ , \new_[20900]_ ,
    \new_[20901]_ , \new_[20902]_ , \new_[20905]_ , \new_[20909]_ ,
    \new_[20910]_ , \new_[20911]_ , \new_[20914]_ , \new_[20918]_ ,
    \new_[20919]_ , \new_[20920]_ , \new_[20923]_ , \new_[20927]_ ,
    \new_[20928]_ , \new_[20929]_ , \new_[20932]_ , \new_[20936]_ ,
    \new_[20937]_ , \new_[20938]_ , \new_[20941]_ , \new_[20945]_ ,
    \new_[20946]_ , \new_[20947]_ , \new_[20950]_ , \new_[20954]_ ,
    \new_[20955]_ , \new_[20956]_ , \new_[20959]_ , \new_[20963]_ ,
    \new_[20964]_ , \new_[20965]_ , \new_[20968]_ , \new_[20972]_ ,
    \new_[20973]_ , \new_[20974]_ , \new_[20977]_ , \new_[20981]_ ,
    \new_[20982]_ , \new_[20983]_ , \new_[20986]_ , \new_[20990]_ ,
    \new_[20991]_ , \new_[20992]_ , \new_[20995]_ , \new_[20999]_ ,
    \new_[21000]_ , \new_[21001]_ , \new_[21004]_ , \new_[21008]_ ,
    \new_[21009]_ , \new_[21010]_ , \new_[21013]_ , \new_[21017]_ ,
    \new_[21018]_ , \new_[21019]_ , \new_[21022]_ , \new_[21026]_ ,
    \new_[21027]_ , \new_[21028]_ , \new_[21031]_ , \new_[21035]_ ,
    \new_[21036]_ , \new_[21037]_ , \new_[21040]_ , \new_[21044]_ ,
    \new_[21045]_ , \new_[21046]_ , \new_[21049]_ , \new_[21053]_ ,
    \new_[21054]_ , \new_[21055]_ , \new_[21058]_ , \new_[21062]_ ,
    \new_[21063]_ , \new_[21064]_ , \new_[21067]_ , \new_[21071]_ ,
    \new_[21072]_ , \new_[21073]_ , \new_[21076]_ , \new_[21080]_ ,
    \new_[21081]_ , \new_[21082]_ , \new_[21085]_ , \new_[21089]_ ,
    \new_[21090]_ , \new_[21091]_ , \new_[21094]_ , \new_[21098]_ ,
    \new_[21099]_ , \new_[21100]_ , \new_[21103]_ , \new_[21107]_ ,
    \new_[21108]_ , \new_[21109]_ , \new_[21112]_ , \new_[21116]_ ,
    \new_[21117]_ , \new_[21118]_ , \new_[21121]_ , \new_[21125]_ ,
    \new_[21126]_ , \new_[21127]_ , \new_[21130]_ , \new_[21134]_ ,
    \new_[21135]_ , \new_[21136]_ , \new_[21139]_ , \new_[21143]_ ,
    \new_[21144]_ , \new_[21145]_ , \new_[21148]_ , \new_[21152]_ ,
    \new_[21153]_ , \new_[21154]_ , \new_[21157]_ , \new_[21161]_ ,
    \new_[21162]_ , \new_[21163]_ , \new_[21166]_ , \new_[21170]_ ,
    \new_[21171]_ , \new_[21172]_ , \new_[21175]_ , \new_[21179]_ ,
    \new_[21180]_ , \new_[21181]_ , \new_[21184]_ , \new_[21188]_ ,
    \new_[21189]_ , \new_[21190]_ , \new_[21193]_ , \new_[21197]_ ,
    \new_[21198]_ , \new_[21199]_ , \new_[21202]_ , \new_[21206]_ ,
    \new_[21207]_ , \new_[21208]_ , \new_[21211]_ , \new_[21215]_ ,
    \new_[21216]_ , \new_[21217]_ , \new_[21220]_ , \new_[21224]_ ,
    \new_[21225]_ , \new_[21226]_ , \new_[21229]_ , \new_[21233]_ ,
    \new_[21234]_ , \new_[21235]_ , \new_[21238]_ , \new_[21242]_ ,
    \new_[21243]_ , \new_[21244]_ , \new_[21247]_ , \new_[21251]_ ,
    \new_[21252]_ , \new_[21253]_ , \new_[21256]_ , \new_[21260]_ ,
    \new_[21261]_ , \new_[21262]_ , \new_[21265]_ , \new_[21269]_ ,
    \new_[21270]_ , \new_[21271]_ , \new_[21274]_ , \new_[21278]_ ,
    \new_[21279]_ , \new_[21280]_ , \new_[21283]_ , \new_[21287]_ ,
    \new_[21288]_ , \new_[21289]_ , \new_[21292]_ , \new_[21296]_ ,
    \new_[21297]_ , \new_[21298]_ , \new_[21301]_ , \new_[21305]_ ,
    \new_[21306]_ , \new_[21307]_ , \new_[21310]_ , \new_[21314]_ ,
    \new_[21315]_ , \new_[21316]_ , \new_[21319]_ , \new_[21323]_ ,
    \new_[21324]_ , \new_[21325]_ , \new_[21328]_ , \new_[21332]_ ,
    \new_[21333]_ , \new_[21334]_ , \new_[21337]_ , \new_[21341]_ ,
    \new_[21342]_ , \new_[21343]_ , \new_[21346]_ , \new_[21350]_ ,
    \new_[21351]_ , \new_[21352]_ , \new_[21355]_ , \new_[21359]_ ,
    \new_[21360]_ , \new_[21361]_ , \new_[21364]_ , \new_[21368]_ ,
    \new_[21369]_ , \new_[21370]_ , \new_[21373]_ , \new_[21377]_ ,
    \new_[21378]_ , \new_[21379]_ , \new_[21382]_ , \new_[21386]_ ,
    \new_[21387]_ , \new_[21388]_ , \new_[21391]_ , \new_[21395]_ ,
    \new_[21396]_ , \new_[21397]_ , \new_[21400]_ , \new_[21404]_ ,
    \new_[21405]_ , \new_[21406]_ , \new_[21409]_ , \new_[21413]_ ,
    \new_[21414]_ , \new_[21415]_ , \new_[21418]_ , \new_[21422]_ ,
    \new_[21423]_ , \new_[21424]_ , \new_[21427]_ , \new_[21431]_ ,
    \new_[21432]_ , \new_[21433]_ , \new_[21436]_ , \new_[21440]_ ,
    \new_[21441]_ , \new_[21442]_ , \new_[21445]_ , \new_[21449]_ ,
    \new_[21450]_ , \new_[21451]_ , \new_[21454]_ , \new_[21458]_ ,
    \new_[21459]_ , \new_[21460]_ , \new_[21463]_ , \new_[21467]_ ,
    \new_[21468]_ , \new_[21469]_ , \new_[21472]_ , \new_[21476]_ ,
    \new_[21477]_ , \new_[21478]_ , \new_[21481]_ , \new_[21485]_ ,
    \new_[21486]_ , \new_[21487]_ , \new_[21490]_ , \new_[21494]_ ,
    \new_[21495]_ , \new_[21496]_ , \new_[21499]_ , \new_[21503]_ ,
    \new_[21504]_ , \new_[21505]_ , \new_[21508]_ , \new_[21512]_ ,
    \new_[21513]_ , \new_[21514]_ , \new_[21517]_ , \new_[21521]_ ,
    \new_[21522]_ , \new_[21523]_ , \new_[21526]_ , \new_[21530]_ ,
    \new_[21531]_ , \new_[21532]_ , \new_[21535]_ , \new_[21539]_ ,
    \new_[21540]_ , \new_[21541]_ , \new_[21544]_ , \new_[21548]_ ,
    \new_[21549]_ , \new_[21550]_ , \new_[21553]_ , \new_[21557]_ ,
    \new_[21558]_ , \new_[21559]_ , \new_[21562]_ , \new_[21566]_ ,
    \new_[21567]_ , \new_[21568]_ , \new_[21571]_ , \new_[21575]_ ,
    \new_[21576]_ , \new_[21577]_ , \new_[21580]_ , \new_[21584]_ ,
    \new_[21585]_ , \new_[21586]_ , \new_[21589]_ , \new_[21593]_ ,
    \new_[21594]_ , \new_[21595]_ , \new_[21598]_ , \new_[21602]_ ,
    \new_[21603]_ , \new_[21604]_ , \new_[21607]_ , \new_[21611]_ ,
    \new_[21612]_ , \new_[21613]_ , \new_[21616]_ , \new_[21620]_ ,
    \new_[21621]_ , \new_[21622]_ , \new_[21625]_ , \new_[21629]_ ,
    \new_[21630]_ , \new_[21631]_ , \new_[21634]_ , \new_[21638]_ ,
    \new_[21639]_ , \new_[21640]_ , \new_[21643]_ , \new_[21647]_ ,
    \new_[21648]_ , \new_[21649]_ , \new_[21652]_ , \new_[21656]_ ,
    \new_[21657]_ , \new_[21658]_ , \new_[21661]_ , \new_[21665]_ ,
    \new_[21666]_ , \new_[21667]_ , \new_[21670]_ , \new_[21674]_ ,
    \new_[21675]_ , \new_[21676]_ , \new_[21679]_ , \new_[21683]_ ,
    \new_[21684]_ , \new_[21685]_ , \new_[21688]_ , \new_[21692]_ ,
    \new_[21693]_ , \new_[21694]_ , \new_[21697]_ , \new_[21701]_ ,
    \new_[21702]_ , \new_[21703]_ , \new_[21706]_ , \new_[21710]_ ,
    \new_[21711]_ , \new_[21712]_ , \new_[21715]_ , \new_[21719]_ ,
    \new_[21720]_ , \new_[21721]_ , \new_[21724]_ , \new_[21728]_ ,
    \new_[21729]_ , \new_[21730]_ , \new_[21733]_ , \new_[21737]_ ,
    \new_[21738]_ , \new_[21739]_ , \new_[21742]_ , \new_[21746]_ ,
    \new_[21747]_ , \new_[21748]_ , \new_[21751]_ , \new_[21755]_ ,
    \new_[21756]_ , \new_[21757]_ , \new_[21760]_ , \new_[21764]_ ,
    \new_[21765]_ , \new_[21766]_ , \new_[21769]_ , \new_[21773]_ ,
    \new_[21774]_ , \new_[21775]_ , \new_[21778]_ , \new_[21782]_ ,
    \new_[21783]_ , \new_[21784]_ , \new_[21787]_ , \new_[21791]_ ,
    \new_[21792]_ , \new_[21793]_ , \new_[21796]_ , \new_[21800]_ ,
    \new_[21801]_ , \new_[21802]_ , \new_[21805]_ , \new_[21809]_ ,
    \new_[21810]_ , \new_[21811]_ , \new_[21814]_ , \new_[21818]_ ,
    \new_[21819]_ , \new_[21820]_ , \new_[21823]_ , \new_[21827]_ ,
    \new_[21828]_ , \new_[21829]_ , \new_[21832]_ , \new_[21836]_ ,
    \new_[21837]_ , \new_[21838]_ , \new_[21841]_ , \new_[21845]_ ,
    \new_[21846]_ , \new_[21847]_ , \new_[21850]_ , \new_[21854]_ ,
    \new_[21855]_ , \new_[21856]_ , \new_[21859]_ , \new_[21863]_ ,
    \new_[21864]_ , \new_[21865]_ , \new_[21868]_ , \new_[21872]_ ,
    \new_[21873]_ , \new_[21874]_ , \new_[21877]_ , \new_[21881]_ ,
    \new_[21882]_ , \new_[21883]_ , \new_[21886]_ , \new_[21890]_ ,
    \new_[21891]_ , \new_[21892]_ , \new_[21895]_ , \new_[21899]_ ,
    \new_[21900]_ , \new_[21901]_ , \new_[21904]_ , \new_[21908]_ ,
    \new_[21909]_ , \new_[21910]_ , \new_[21913]_ , \new_[21917]_ ,
    \new_[21918]_ , \new_[21919]_ , \new_[21922]_ , \new_[21926]_ ,
    \new_[21927]_ , \new_[21928]_ , \new_[21931]_ , \new_[21935]_ ,
    \new_[21936]_ , \new_[21937]_ , \new_[21940]_ , \new_[21944]_ ,
    \new_[21945]_ , \new_[21946]_ , \new_[21949]_ , \new_[21953]_ ,
    \new_[21954]_ , \new_[21955]_ , \new_[21958]_ , \new_[21962]_ ,
    \new_[21963]_ , \new_[21964]_ , \new_[21967]_ , \new_[21971]_ ,
    \new_[21972]_ , \new_[21973]_ , \new_[21976]_ , \new_[21980]_ ,
    \new_[21981]_ , \new_[21982]_ , \new_[21985]_ , \new_[21989]_ ,
    \new_[21990]_ , \new_[21991]_ , \new_[21994]_ , \new_[21998]_ ,
    \new_[21999]_ , \new_[22000]_ , \new_[22003]_ , \new_[22007]_ ,
    \new_[22008]_ , \new_[22009]_ , \new_[22012]_ , \new_[22016]_ ,
    \new_[22017]_ , \new_[22018]_ , \new_[22021]_ , \new_[22025]_ ,
    \new_[22026]_ , \new_[22027]_ , \new_[22030]_ , \new_[22034]_ ,
    \new_[22035]_ , \new_[22036]_ , \new_[22039]_ , \new_[22043]_ ,
    \new_[22044]_ , \new_[22045]_ , \new_[22048]_ , \new_[22052]_ ,
    \new_[22053]_ , \new_[22054]_ , \new_[22057]_ , \new_[22061]_ ,
    \new_[22062]_ , \new_[22063]_ , \new_[22066]_ , \new_[22070]_ ,
    \new_[22071]_ , \new_[22072]_ , \new_[22075]_ , \new_[22079]_ ,
    \new_[22080]_ , \new_[22081]_ , \new_[22084]_ , \new_[22088]_ ,
    \new_[22089]_ , \new_[22090]_ , \new_[22093]_ , \new_[22097]_ ,
    \new_[22098]_ , \new_[22099]_ , \new_[22102]_ , \new_[22106]_ ,
    \new_[22107]_ , \new_[22108]_ , \new_[22111]_ , \new_[22115]_ ,
    \new_[22116]_ , \new_[22117]_ , \new_[22120]_ , \new_[22124]_ ,
    \new_[22125]_ , \new_[22126]_ , \new_[22129]_ , \new_[22133]_ ,
    \new_[22134]_ , \new_[22135]_ , \new_[22138]_ , \new_[22142]_ ,
    \new_[22143]_ , \new_[22144]_ , \new_[22147]_ , \new_[22151]_ ,
    \new_[22152]_ , \new_[22153]_ , \new_[22156]_ , \new_[22160]_ ,
    \new_[22161]_ , \new_[22162]_ , \new_[22165]_ , \new_[22169]_ ,
    \new_[22170]_ , \new_[22171]_ , \new_[22174]_ , \new_[22178]_ ,
    \new_[22179]_ , \new_[22180]_ , \new_[22183]_ , \new_[22187]_ ,
    \new_[22188]_ , \new_[22189]_ , \new_[22192]_ , \new_[22196]_ ,
    \new_[22197]_ , \new_[22198]_ , \new_[22201]_ , \new_[22205]_ ,
    \new_[22206]_ , \new_[22207]_ , \new_[22210]_ , \new_[22214]_ ,
    \new_[22215]_ , \new_[22216]_ , \new_[22219]_ , \new_[22223]_ ,
    \new_[22224]_ , \new_[22225]_ , \new_[22228]_ , \new_[22232]_ ,
    \new_[22233]_ , \new_[22234]_ , \new_[22237]_ , \new_[22241]_ ,
    \new_[22242]_ , \new_[22243]_ , \new_[22246]_ , \new_[22250]_ ,
    \new_[22251]_ , \new_[22252]_ , \new_[22255]_ , \new_[22259]_ ,
    \new_[22260]_ , \new_[22261]_ , \new_[22264]_ , \new_[22268]_ ,
    \new_[22269]_ , \new_[22270]_ , \new_[22273]_ , \new_[22277]_ ,
    \new_[22278]_ , \new_[22279]_ , \new_[22282]_ , \new_[22286]_ ,
    \new_[22287]_ , \new_[22288]_ , \new_[22291]_ , \new_[22295]_ ,
    \new_[22296]_ , \new_[22297]_ , \new_[22300]_ , \new_[22304]_ ,
    \new_[22305]_ , \new_[22306]_ , \new_[22309]_ , \new_[22313]_ ,
    \new_[22314]_ , \new_[22315]_ , \new_[22318]_ , \new_[22322]_ ,
    \new_[22323]_ , \new_[22324]_ , \new_[22327]_ , \new_[22331]_ ,
    \new_[22332]_ , \new_[22333]_ , \new_[22336]_ , \new_[22340]_ ,
    \new_[22341]_ , \new_[22342]_ , \new_[22345]_ , \new_[22349]_ ,
    \new_[22350]_ , \new_[22351]_ , \new_[22354]_ , \new_[22358]_ ,
    \new_[22359]_ , \new_[22360]_ , \new_[22363]_ , \new_[22367]_ ,
    \new_[22368]_ , \new_[22369]_ , \new_[22372]_ , \new_[22376]_ ,
    \new_[22377]_ , \new_[22378]_ , \new_[22381]_ , \new_[22385]_ ,
    \new_[22386]_ , \new_[22387]_ , \new_[22390]_ , \new_[22394]_ ,
    \new_[22395]_ , \new_[22396]_ , \new_[22399]_ , \new_[22403]_ ,
    \new_[22404]_ , \new_[22405]_ , \new_[22408]_ , \new_[22412]_ ,
    \new_[22413]_ , \new_[22414]_ , \new_[22417]_ , \new_[22421]_ ,
    \new_[22422]_ , \new_[22423]_ , \new_[22426]_ , \new_[22430]_ ,
    \new_[22431]_ , \new_[22432]_ , \new_[22435]_ , \new_[22439]_ ,
    \new_[22440]_ , \new_[22441]_ , \new_[22444]_ , \new_[22448]_ ,
    \new_[22449]_ , \new_[22450]_ , \new_[22453]_ , \new_[22457]_ ,
    \new_[22458]_ , \new_[22459]_ , \new_[22462]_ , \new_[22466]_ ,
    \new_[22467]_ , \new_[22468]_ , \new_[22471]_ , \new_[22475]_ ,
    \new_[22476]_ , \new_[22477]_ , \new_[22480]_ , \new_[22484]_ ,
    \new_[22485]_ , \new_[22486]_ , \new_[22489]_ , \new_[22493]_ ,
    \new_[22494]_ , \new_[22495]_ , \new_[22498]_ , \new_[22502]_ ,
    \new_[22503]_ , \new_[22504]_ , \new_[22507]_ , \new_[22511]_ ,
    \new_[22512]_ , \new_[22513]_ , \new_[22516]_ , \new_[22520]_ ,
    \new_[22521]_ , \new_[22522]_ , \new_[22525]_ , \new_[22529]_ ,
    \new_[22530]_ , \new_[22531]_ , \new_[22534]_ , \new_[22538]_ ,
    \new_[22539]_ , \new_[22540]_ , \new_[22543]_ , \new_[22547]_ ,
    \new_[22548]_ , \new_[22549]_ , \new_[22552]_ , \new_[22556]_ ,
    \new_[22557]_ , \new_[22558]_ , \new_[22561]_ , \new_[22565]_ ,
    \new_[22566]_ , \new_[22567]_ , \new_[22570]_ , \new_[22574]_ ,
    \new_[22575]_ , \new_[22576]_ , \new_[22579]_ , \new_[22583]_ ,
    \new_[22584]_ , \new_[22585]_ , \new_[22588]_ , \new_[22592]_ ,
    \new_[22593]_ , \new_[22594]_ , \new_[22597]_ , \new_[22601]_ ,
    \new_[22602]_ , \new_[22603]_ , \new_[22606]_ , \new_[22610]_ ,
    \new_[22611]_ , \new_[22612]_ , \new_[22615]_ , \new_[22619]_ ,
    \new_[22620]_ , \new_[22621]_ , \new_[22624]_ , \new_[22628]_ ,
    \new_[22629]_ , \new_[22630]_ , \new_[22633]_ , \new_[22637]_ ,
    \new_[22638]_ , \new_[22639]_ , \new_[22642]_ , \new_[22646]_ ,
    \new_[22647]_ , \new_[22648]_ , \new_[22651]_ , \new_[22655]_ ,
    \new_[22656]_ , \new_[22657]_ , \new_[22660]_ , \new_[22664]_ ,
    \new_[22665]_ , \new_[22666]_ , \new_[22669]_ , \new_[22673]_ ,
    \new_[22674]_ , \new_[22675]_ , \new_[22678]_ , \new_[22682]_ ,
    \new_[22683]_ , \new_[22684]_ , \new_[22687]_ , \new_[22691]_ ,
    \new_[22692]_ , \new_[22693]_ , \new_[22696]_ , \new_[22700]_ ,
    \new_[22701]_ , \new_[22702]_ , \new_[22705]_ , \new_[22709]_ ,
    \new_[22710]_ , \new_[22711]_ , \new_[22714]_ , \new_[22718]_ ,
    \new_[22719]_ , \new_[22720]_ , \new_[22723]_ , \new_[22727]_ ,
    \new_[22728]_ , \new_[22729]_ , \new_[22733]_ , \new_[22734]_ ,
    \new_[22738]_ , \new_[22739]_ , \new_[22740]_ , \new_[22743]_ ,
    \new_[22747]_ , \new_[22748]_ , \new_[22749]_ , \new_[22753]_ ,
    \new_[22754]_ , \new_[22758]_ , \new_[22759]_ , \new_[22760]_ ,
    \new_[22763]_ , \new_[22767]_ , \new_[22768]_ , \new_[22769]_ ,
    \new_[22773]_ , \new_[22774]_ , \new_[22778]_ , \new_[22779]_ ,
    \new_[22780]_ , \new_[22783]_ , \new_[22787]_ , \new_[22788]_ ,
    \new_[22789]_ , \new_[22793]_ , \new_[22794]_ , \new_[22798]_ ,
    \new_[22799]_ , \new_[22800]_ , \new_[22803]_ , \new_[22807]_ ,
    \new_[22808]_ , \new_[22809]_ , \new_[22813]_ , \new_[22814]_ ,
    \new_[22818]_ , \new_[22819]_ , \new_[22820]_ , \new_[22823]_ ,
    \new_[22827]_ , \new_[22828]_ , \new_[22829]_ , \new_[22833]_ ,
    \new_[22834]_ , \new_[22838]_ , \new_[22839]_ , \new_[22840]_ ,
    \new_[22843]_ , \new_[22847]_ , \new_[22848]_ , \new_[22849]_ ,
    \new_[22853]_ , \new_[22854]_ , \new_[22858]_ , \new_[22859]_ ,
    \new_[22860]_ , \new_[22863]_ , \new_[22867]_ , \new_[22868]_ ,
    \new_[22869]_ , \new_[22873]_ , \new_[22874]_ , \new_[22878]_ ,
    \new_[22879]_ , \new_[22880]_ , \new_[22883]_ , \new_[22887]_ ,
    \new_[22888]_ , \new_[22889]_ , \new_[22893]_ , \new_[22894]_ ,
    \new_[22898]_ , \new_[22899]_ , \new_[22900]_ , \new_[22903]_ ,
    \new_[22907]_ , \new_[22908]_ , \new_[22909]_ , \new_[22913]_ ,
    \new_[22914]_ , \new_[22918]_ , \new_[22919]_ , \new_[22920]_ ,
    \new_[22923]_ , \new_[22927]_ , \new_[22928]_ , \new_[22929]_ ,
    \new_[22933]_ , \new_[22934]_ , \new_[22938]_ , \new_[22939]_ ,
    \new_[22940]_ , \new_[22943]_ , \new_[22947]_ , \new_[22948]_ ,
    \new_[22949]_ , \new_[22953]_ , \new_[22954]_ , \new_[22958]_ ,
    \new_[22959]_ , \new_[22960]_ , \new_[22963]_ , \new_[22967]_ ,
    \new_[22968]_ , \new_[22969]_ , \new_[22973]_ , \new_[22974]_ ,
    \new_[22978]_ , \new_[22979]_ , \new_[22980]_ , \new_[22983]_ ,
    \new_[22987]_ , \new_[22988]_ , \new_[22989]_ , \new_[22993]_ ,
    \new_[22994]_ , \new_[22998]_ , \new_[22999]_ , \new_[23000]_ ,
    \new_[23003]_ , \new_[23007]_ , \new_[23008]_ , \new_[23009]_ ,
    \new_[23013]_ , \new_[23014]_ , \new_[23018]_ , \new_[23019]_ ,
    \new_[23020]_ , \new_[23023]_ , \new_[23027]_ , \new_[23028]_ ,
    \new_[23029]_ , \new_[23033]_ , \new_[23034]_ , \new_[23038]_ ,
    \new_[23039]_ , \new_[23040]_ , \new_[23043]_ , \new_[23047]_ ,
    \new_[23048]_ , \new_[23049]_ , \new_[23053]_ , \new_[23054]_ ,
    \new_[23058]_ , \new_[23059]_ , \new_[23060]_ , \new_[23063]_ ,
    \new_[23067]_ , \new_[23068]_ , \new_[23069]_ , \new_[23073]_ ,
    \new_[23074]_ , \new_[23078]_ , \new_[23079]_ , \new_[23080]_ ,
    \new_[23083]_ , \new_[23087]_ , \new_[23088]_ , \new_[23089]_ ,
    \new_[23093]_ , \new_[23094]_ , \new_[23098]_ , \new_[23099]_ ,
    \new_[23100]_ , \new_[23103]_ , \new_[23107]_ , \new_[23108]_ ,
    \new_[23109]_ , \new_[23113]_ , \new_[23114]_ , \new_[23118]_ ,
    \new_[23119]_ , \new_[23120]_ , \new_[23123]_ , \new_[23127]_ ,
    \new_[23128]_ , \new_[23129]_ , \new_[23133]_ , \new_[23134]_ ,
    \new_[23138]_ , \new_[23139]_ , \new_[23140]_ , \new_[23143]_ ,
    \new_[23147]_ , \new_[23148]_ , \new_[23149]_ , \new_[23153]_ ,
    \new_[23154]_ , \new_[23158]_ , \new_[23159]_ , \new_[23160]_ ,
    \new_[23163]_ , \new_[23167]_ , \new_[23168]_ , \new_[23169]_ ,
    \new_[23173]_ , \new_[23174]_ , \new_[23178]_ , \new_[23179]_ ,
    \new_[23180]_ , \new_[23183]_ , \new_[23187]_ , \new_[23188]_ ,
    \new_[23189]_ , \new_[23193]_ , \new_[23194]_ , \new_[23198]_ ,
    \new_[23199]_ , \new_[23200]_ , \new_[23203]_ , \new_[23207]_ ,
    \new_[23208]_ , \new_[23209]_ , \new_[23213]_ , \new_[23214]_ ,
    \new_[23218]_ , \new_[23219]_ , \new_[23220]_ , \new_[23223]_ ,
    \new_[23227]_ , \new_[23228]_ , \new_[23229]_ , \new_[23233]_ ,
    \new_[23234]_ , \new_[23238]_ , \new_[23239]_ , \new_[23240]_ ,
    \new_[23243]_ , \new_[23247]_ , \new_[23248]_ , \new_[23249]_ ,
    \new_[23253]_ , \new_[23254]_ , \new_[23258]_ , \new_[23259]_ ,
    \new_[23260]_ , \new_[23263]_ , \new_[23267]_ , \new_[23268]_ ,
    \new_[23269]_ , \new_[23273]_ , \new_[23274]_ , \new_[23278]_ ,
    \new_[23279]_ , \new_[23280]_ , \new_[23283]_ , \new_[23287]_ ,
    \new_[23288]_ , \new_[23289]_ , \new_[23293]_ , \new_[23294]_ ,
    \new_[23298]_ , \new_[23299]_ , \new_[23300]_ , \new_[23303]_ ,
    \new_[23307]_ , \new_[23308]_ , \new_[23309]_ , \new_[23313]_ ,
    \new_[23314]_ , \new_[23318]_ , \new_[23319]_ , \new_[23320]_ ,
    \new_[23323]_ , \new_[23327]_ , \new_[23328]_ , \new_[23329]_ ,
    \new_[23333]_ , \new_[23334]_ , \new_[23338]_ , \new_[23339]_ ,
    \new_[23340]_ , \new_[23343]_ , \new_[23347]_ , \new_[23348]_ ,
    \new_[23349]_ , \new_[23353]_ , \new_[23354]_ , \new_[23358]_ ,
    \new_[23359]_ , \new_[23360]_ , \new_[23363]_ , \new_[23367]_ ,
    \new_[23368]_ , \new_[23369]_ , \new_[23373]_ , \new_[23374]_ ,
    \new_[23378]_ , \new_[23379]_ , \new_[23380]_ , \new_[23383]_ ,
    \new_[23387]_ , \new_[23388]_ , \new_[23389]_ , \new_[23393]_ ,
    \new_[23394]_ , \new_[23398]_ , \new_[23399]_ , \new_[23400]_ ,
    \new_[23403]_ , \new_[23407]_ , \new_[23408]_ , \new_[23409]_ ,
    \new_[23413]_ , \new_[23414]_ , \new_[23418]_ , \new_[23419]_ ,
    \new_[23420]_ , \new_[23423]_ , \new_[23427]_ , \new_[23428]_ ,
    \new_[23429]_ , \new_[23433]_ , \new_[23434]_ , \new_[23438]_ ,
    \new_[23439]_ , \new_[23440]_ , \new_[23443]_ , \new_[23447]_ ,
    \new_[23448]_ , \new_[23449]_ , \new_[23453]_ , \new_[23454]_ ,
    \new_[23458]_ , \new_[23459]_ , \new_[23460]_ , \new_[23463]_ ,
    \new_[23467]_ , \new_[23468]_ , \new_[23469]_ , \new_[23473]_ ,
    \new_[23474]_ , \new_[23478]_ , \new_[23479]_ , \new_[23480]_ ,
    \new_[23483]_ , \new_[23487]_ , \new_[23488]_ , \new_[23489]_ ,
    \new_[23493]_ , \new_[23494]_ , \new_[23498]_ , \new_[23499]_ ,
    \new_[23500]_ , \new_[23503]_ , \new_[23507]_ , \new_[23508]_ ,
    \new_[23509]_ , \new_[23513]_ , \new_[23514]_ , \new_[23518]_ ,
    \new_[23519]_ , \new_[23520]_ , \new_[23523]_ , \new_[23527]_ ,
    \new_[23528]_ , \new_[23529]_ , \new_[23533]_ , \new_[23534]_ ,
    \new_[23538]_ , \new_[23539]_ , \new_[23540]_ , \new_[23543]_ ,
    \new_[23547]_ , \new_[23548]_ , \new_[23549]_ , \new_[23553]_ ,
    \new_[23554]_ , \new_[23558]_ , \new_[23559]_ , \new_[23560]_ ,
    \new_[23563]_ , \new_[23567]_ , \new_[23568]_ , \new_[23569]_ ,
    \new_[23573]_ , \new_[23574]_ , \new_[23578]_ , \new_[23579]_ ,
    \new_[23580]_ , \new_[23583]_ , \new_[23587]_ , \new_[23588]_ ,
    \new_[23589]_ , \new_[23593]_ , \new_[23594]_ , \new_[23598]_ ,
    \new_[23599]_ , \new_[23600]_ , \new_[23603]_ , \new_[23607]_ ,
    \new_[23608]_ , \new_[23609]_ , \new_[23613]_ , \new_[23614]_ ,
    \new_[23618]_ , \new_[23619]_ , \new_[23620]_ , \new_[23623]_ ,
    \new_[23627]_ , \new_[23628]_ , \new_[23629]_ , \new_[23633]_ ,
    \new_[23634]_ , \new_[23638]_ , \new_[23639]_ , \new_[23640]_ ,
    \new_[23643]_ , \new_[23647]_ , \new_[23648]_ , \new_[23649]_ ,
    \new_[23653]_ , \new_[23654]_ , \new_[23658]_ , \new_[23659]_ ,
    \new_[23660]_ , \new_[23663]_ , \new_[23667]_ , \new_[23668]_ ,
    \new_[23669]_ , \new_[23673]_ , \new_[23674]_ , \new_[23678]_ ,
    \new_[23679]_ , \new_[23680]_ , \new_[23683]_ , \new_[23687]_ ,
    \new_[23688]_ , \new_[23689]_ , \new_[23693]_ , \new_[23694]_ ,
    \new_[23698]_ , \new_[23699]_ , \new_[23700]_ , \new_[23703]_ ,
    \new_[23707]_ , \new_[23708]_ , \new_[23709]_ , \new_[23713]_ ,
    \new_[23714]_ , \new_[23718]_ , \new_[23719]_ , \new_[23720]_ ,
    \new_[23723]_ , \new_[23727]_ , \new_[23728]_ , \new_[23729]_ ,
    \new_[23733]_ , \new_[23734]_ , \new_[23738]_ , \new_[23739]_ ,
    \new_[23740]_ , \new_[23743]_ , \new_[23747]_ , \new_[23748]_ ,
    \new_[23749]_ , \new_[23753]_ , \new_[23754]_ , \new_[23758]_ ,
    \new_[23759]_ , \new_[23760]_ , \new_[23763]_ , \new_[23767]_ ,
    \new_[23768]_ , \new_[23769]_ , \new_[23773]_ , \new_[23774]_ ,
    \new_[23778]_ , \new_[23779]_ , \new_[23780]_ , \new_[23783]_ ,
    \new_[23787]_ , \new_[23788]_ , \new_[23789]_ , \new_[23793]_ ,
    \new_[23794]_ , \new_[23798]_ , \new_[23799]_ , \new_[23800]_ ,
    \new_[23803]_ , \new_[23807]_ , \new_[23808]_ , \new_[23809]_ ,
    \new_[23813]_ , \new_[23814]_ , \new_[23818]_ , \new_[23819]_ ,
    \new_[23820]_ , \new_[23823]_ , \new_[23827]_ , \new_[23828]_ ,
    \new_[23829]_ , \new_[23833]_ , \new_[23834]_ , \new_[23838]_ ,
    \new_[23839]_ , \new_[23840]_ , \new_[23843]_ , \new_[23847]_ ,
    \new_[23848]_ , \new_[23849]_ , \new_[23853]_ , \new_[23854]_ ,
    \new_[23858]_ , \new_[23859]_ , \new_[23860]_ , \new_[23863]_ ,
    \new_[23867]_ , \new_[23868]_ , \new_[23869]_ , \new_[23873]_ ,
    \new_[23874]_ , \new_[23878]_ , \new_[23879]_ , \new_[23880]_ ,
    \new_[23883]_ , \new_[23887]_ , \new_[23888]_ , \new_[23889]_ ,
    \new_[23893]_ , \new_[23894]_ , \new_[23898]_ , \new_[23899]_ ,
    \new_[23900]_ , \new_[23903]_ , \new_[23907]_ , \new_[23908]_ ,
    \new_[23909]_ , \new_[23913]_ , \new_[23914]_ , \new_[23918]_ ,
    \new_[23919]_ , \new_[23920]_ , \new_[23923]_ , \new_[23927]_ ,
    \new_[23928]_ , \new_[23929]_ , \new_[23933]_ , \new_[23934]_ ,
    \new_[23938]_ , \new_[23939]_ , \new_[23940]_ , \new_[23943]_ ,
    \new_[23947]_ , \new_[23948]_ , \new_[23949]_ , \new_[23953]_ ,
    \new_[23954]_ , \new_[23958]_ , \new_[23959]_ , \new_[23960]_ ,
    \new_[23963]_ , \new_[23967]_ , \new_[23968]_ , \new_[23969]_ ,
    \new_[23973]_ , \new_[23974]_ , \new_[23978]_ , \new_[23979]_ ,
    \new_[23980]_ , \new_[23983]_ , \new_[23987]_ , \new_[23988]_ ,
    \new_[23989]_ , \new_[23993]_ , \new_[23994]_ , \new_[23998]_ ,
    \new_[23999]_ , \new_[24000]_ , \new_[24003]_ , \new_[24007]_ ,
    \new_[24008]_ , \new_[24009]_ , \new_[24013]_ , \new_[24014]_ ,
    \new_[24018]_ , \new_[24019]_ , \new_[24020]_ , \new_[24023]_ ,
    \new_[24027]_ , \new_[24028]_ , \new_[24029]_ , \new_[24033]_ ,
    \new_[24034]_ , \new_[24038]_ , \new_[24039]_ , \new_[24040]_ ,
    \new_[24043]_ , \new_[24047]_ , \new_[24048]_ , \new_[24049]_ ,
    \new_[24053]_ , \new_[24054]_ , \new_[24058]_ , \new_[24059]_ ,
    \new_[24060]_ , \new_[24063]_ , \new_[24067]_ , \new_[24068]_ ,
    \new_[24069]_ , \new_[24073]_ , \new_[24074]_ , \new_[24078]_ ,
    \new_[24079]_ , \new_[24080]_ , \new_[24083]_ , \new_[24087]_ ,
    \new_[24088]_ , \new_[24089]_ , \new_[24093]_ , \new_[24094]_ ,
    \new_[24098]_ , \new_[24099]_ , \new_[24100]_ , \new_[24103]_ ,
    \new_[24107]_ , \new_[24108]_ , \new_[24109]_ , \new_[24113]_ ,
    \new_[24114]_ , \new_[24118]_ , \new_[24119]_ , \new_[24120]_ ,
    \new_[24123]_ , \new_[24127]_ , \new_[24128]_ , \new_[24129]_ ,
    \new_[24133]_ , \new_[24134]_ , \new_[24138]_ , \new_[24139]_ ,
    \new_[24140]_ , \new_[24143]_ , \new_[24147]_ , \new_[24148]_ ,
    \new_[24149]_ , \new_[24153]_ , \new_[24154]_ , \new_[24158]_ ,
    \new_[24159]_ , \new_[24160]_ , \new_[24163]_ , \new_[24167]_ ,
    \new_[24168]_ , \new_[24169]_ , \new_[24173]_ , \new_[24174]_ ,
    \new_[24178]_ , \new_[24179]_ , \new_[24180]_ , \new_[24183]_ ,
    \new_[24187]_ , \new_[24188]_ , \new_[24189]_ , \new_[24193]_ ,
    \new_[24194]_ , \new_[24198]_ , \new_[24199]_ , \new_[24200]_ ,
    \new_[24203]_ , \new_[24207]_ , \new_[24208]_ , \new_[24209]_ ,
    \new_[24213]_ , \new_[24214]_ , \new_[24218]_ , \new_[24219]_ ,
    \new_[24220]_ , \new_[24223]_ , \new_[24227]_ , \new_[24228]_ ,
    \new_[24229]_ , \new_[24233]_ , \new_[24234]_ , \new_[24238]_ ,
    \new_[24239]_ , \new_[24240]_ , \new_[24243]_ , \new_[24247]_ ,
    \new_[24248]_ , \new_[24249]_ , \new_[24253]_ , \new_[24254]_ ,
    \new_[24258]_ , \new_[24259]_ , \new_[24260]_ , \new_[24263]_ ,
    \new_[24267]_ , \new_[24268]_ , \new_[24269]_ , \new_[24273]_ ,
    \new_[24274]_ , \new_[24278]_ , \new_[24279]_ , \new_[24280]_ ,
    \new_[24283]_ , \new_[24287]_ , \new_[24288]_ , \new_[24289]_ ,
    \new_[24293]_ , \new_[24294]_ , \new_[24298]_ , \new_[24299]_ ,
    \new_[24300]_ , \new_[24303]_ , \new_[24307]_ , \new_[24308]_ ,
    \new_[24309]_ , \new_[24313]_ , \new_[24314]_ , \new_[24318]_ ,
    \new_[24319]_ , \new_[24320]_ , \new_[24323]_ , \new_[24327]_ ,
    \new_[24328]_ , \new_[24329]_ , \new_[24333]_ , \new_[24334]_ ,
    \new_[24338]_ , \new_[24339]_ , \new_[24340]_ , \new_[24343]_ ,
    \new_[24347]_ , \new_[24348]_ , \new_[24349]_ , \new_[24353]_ ,
    \new_[24354]_ , \new_[24358]_ , \new_[24359]_ , \new_[24360]_ ,
    \new_[24363]_ , \new_[24367]_ , \new_[24368]_ , \new_[24369]_ ,
    \new_[24373]_ , \new_[24374]_ , \new_[24378]_ , \new_[24379]_ ,
    \new_[24380]_ , \new_[24383]_ , \new_[24387]_ , \new_[24388]_ ,
    \new_[24389]_ , \new_[24393]_ , \new_[24394]_ , \new_[24398]_ ,
    \new_[24399]_ , \new_[24400]_ , \new_[24403]_ , \new_[24407]_ ,
    \new_[24408]_ , \new_[24409]_ , \new_[24413]_ , \new_[24414]_ ,
    \new_[24418]_ , \new_[24419]_ , \new_[24420]_ , \new_[24423]_ ,
    \new_[24427]_ , \new_[24428]_ , \new_[24429]_ , \new_[24433]_ ,
    \new_[24434]_ , \new_[24438]_ , \new_[24439]_ , \new_[24440]_ ,
    \new_[24443]_ , \new_[24447]_ , \new_[24448]_ , \new_[24449]_ ,
    \new_[24453]_ , \new_[24454]_ , \new_[24458]_ , \new_[24459]_ ,
    \new_[24460]_ , \new_[24463]_ , \new_[24467]_ , \new_[24468]_ ,
    \new_[24469]_ , \new_[24473]_ , \new_[24474]_ , \new_[24478]_ ,
    \new_[24479]_ , \new_[24480]_ , \new_[24483]_ , \new_[24487]_ ,
    \new_[24488]_ , \new_[24489]_ , \new_[24493]_ , \new_[24494]_ ,
    \new_[24498]_ , \new_[24499]_ , \new_[24500]_ , \new_[24503]_ ,
    \new_[24507]_ , \new_[24508]_ , \new_[24509]_ , \new_[24513]_ ,
    \new_[24514]_ , \new_[24518]_ , \new_[24519]_ , \new_[24520]_ ,
    \new_[24523]_ , \new_[24527]_ , \new_[24528]_ , \new_[24529]_ ,
    \new_[24533]_ , \new_[24534]_ , \new_[24538]_ , \new_[24539]_ ,
    \new_[24540]_ , \new_[24543]_ , \new_[24547]_ , \new_[24548]_ ,
    \new_[24549]_ , \new_[24553]_ , \new_[24554]_ , \new_[24558]_ ,
    \new_[24559]_ , \new_[24560]_ , \new_[24563]_ , \new_[24567]_ ,
    \new_[24568]_ , \new_[24569]_ , \new_[24573]_ , \new_[24574]_ ,
    \new_[24578]_ , \new_[24579]_ , \new_[24580]_ , \new_[24583]_ ,
    \new_[24587]_ , \new_[24588]_ , \new_[24589]_ , \new_[24593]_ ,
    \new_[24594]_ , \new_[24598]_ , \new_[24599]_ , \new_[24600]_ ,
    \new_[24603]_ , \new_[24607]_ , \new_[24608]_ , \new_[24609]_ ,
    \new_[24613]_ , \new_[24614]_ , \new_[24618]_ , \new_[24619]_ ,
    \new_[24620]_ , \new_[24623]_ , \new_[24627]_ , \new_[24628]_ ,
    \new_[24629]_ , \new_[24633]_ , \new_[24634]_ , \new_[24638]_ ,
    \new_[24639]_ , \new_[24640]_ , \new_[24643]_ , \new_[24647]_ ,
    \new_[24648]_ , \new_[24649]_ , \new_[24653]_ , \new_[24654]_ ,
    \new_[24658]_ , \new_[24659]_ , \new_[24660]_ , \new_[24663]_ ,
    \new_[24667]_ , \new_[24668]_ , \new_[24669]_ , \new_[24673]_ ,
    \new_[24674]_ , \new_[24678]_ , \new_[24679]_ , \new_[24680]_ ,
    \new_[24683]_ , \new_[24687]_ , \new_[24688]_ , \new_[24689]_ ,
    \new_[24693]_ , \new_[24694]_ , \new_[24698]_ , \new_[24699]_ ,
    \new_[24700]_ , \new_[24703]_ , \new_[24707]_ , \new_[24708]_ ,
    \new_[24709]_ , \new_[24713]_ , \new_[24714]_ , \new_[24718]_ ,
    \new_[24719]_ , \new_[24720]_ , \new_[24723]_ , \new_[24727]_ ,
    \new_[24728]_ , \new_[24729]_ , \new_[24733]_ , \new_[24734]_ ,
    \new_[24738]_ , \new_[24739]_ , \new_[24740]_ , \new_[24743]_ ,
    \new_[24747]_ , \new_[24748]_ , \new_[24749]_ , \new_[24753]_ ,
    \new_[24754]_ , \new_[24758]_ , \new_[24759]_ , \new_[24760]_ ,
    \new_[24763]_ , \new_[24767]_ , \new_[24768]_ , \new_[24769]_ ,
    \new_[24773]_ , \new_[24774]_ , \new_[24778]_ , \new_[24779]_ ,
    \new_[24780]_ , \new_[24783]_ , \new_[24787]_ , \new_[24788]_ ,
    \new_[24789]_ , \new_[24793]_ , \new_[24794]_ , \new_[24798]_ ,
    \new_[24799]_ , \new_[24800]_ , \new_[24803]_ , \new_[24807]_ ,
    \new_[24808]_ , \new_[24809]_ , \new_[24813]_ , \new_[24814]_ ,
    \new_[24818]_ , \new_[24819]_ , \new_[24820]_ , \new_[24823]_ ,
    \new_[24827]_ , \new_[24828]_ , \new_[24829]_ , \new_[24833]_ ,
    \new_[24834]_ , \new_[24838]_ , \new_[24839]_ , \new_[24840]_ ,
    \new_[24843]_ , \new_[24847]_ , \new_[24848]_ , \new_[24849]_ ,
    \new_[24853]_ , \new_[24854]_ , \new_[24858]_ , \new_[24859]_ ,
    \new_[24860]_ , \new_[24863]_ , \new_[24867]_ , \new_[24868]_ ,
    \new_[24869]_ , \new_[24873]_ , \new_[24874]_ , \new_[24878]_ ,
    \new_[24879]_ , \new_[24880]_ , \new_[24883]_ , \new_[24887]_ ,
    \new_[24888]_ , \new_[24889]_ , \new_[24893]_ , \new_[24894]_ ,
    \new_[24898]_ , \new_[24899]_ , \new_[24900]_ , \new_[24903]_ ,
    \new_[24907]_ , \new_[24908]_ , \new_[24909]_ , \new_[24913]_ ,
    \new_[24914]_ , \new_[24918]_ , \new_[24919]_ , \new_[24920]_ ,
    \new_[24923]_ , \new_[24927]_ , \new_[24928]_ , \new_[24929]_ ,
    \new_[24933]_ , \new_[24934]_ , \new_[24938]_ , \new_[24939]_ ,
    \new_[24940]_ , \new_[24943]_ , \new_[24947]_ , \new_[24948]_ ,
    \new_[24949]_ , \new_[24953]_ , \new_[24954]_ , \new_[24958]_ ,
    \new_[24959]_ , \new_[24960]_ , \new_[24963]_ , \new_[24967]_ ,
    \new_[24968]_ , \new_[24969]_ , \new_[24973]_ , \new_[24974]_ ,
    \new_[24978]_ , \new_[24979]_ , \new_[24980]_ , \new_[24983]_ ,
    \new_[24987]_ , \new_[24988]_ , \new_[24989]_ , \new_[24993]_ ,
    \new_[24994]_ , \new_[24998]_ , \new_[24999]_ , \new_[25000]_ ,
    \new_[25003]_ , \new_[25007]_ , \new_[25008]_ , \new_[25009]_ ,
    \new_[25013]_ , \new_[25014]_ , \new_[25018]_ , \new_[25019]_ ,
    \new_[25020]_ , \new_[25023]_ , \new_[25027]_ , \new_[25028]_ ,
    \new_[25029]_ , \new_[25033]_ , \new_[25034]_ , \new_[25038]_ ,
    \new_[25039]_ , \new_[25040]_ , \new_[25043]_ , \new_[25047]_ ,
    \new_[25048]_ , \new_[25049]_ , \new_[25053]_ , \new_[25054]_ ,
    \new_[25058]_ , \new_[25059]_ , \new_[25060]_ , \new_[25063]_ ,
    \new_[25067]_ , \new_[25068]_ , \new_[25069]_ , \new_[25073]_ ,
    \new_[25074]_ , \new_[25078]_ , \new_[25079]_ , \new_[25080]_ ,
    \new_[25083]_ , \new_[25087]_ , \new_[25088]_ , \new_[25089]_ ,
    \new_[25093]_ , \new_[25094]_ , \new_[25098]_ , \new_[25099]_ ,
    \new_[25100]_ , \new_[25103]_ , \new_[25107]_ , \new_[25108]_ ,
    \new_[25109]_ , \new_[25113]_ , \new_[25114]_ , \new_[25118]_ ,
    \new_[25119]_ , \new_[25120]_ , \new_[25123]_ , \new_[25127]_ ,
    \new_[25128]_ , \new_[25129]_ , \new_[25133]_ , \new_[25134]_ ,
    \new_[25138]_ , \new_[25139]_ , \new_[25140]_ , \new_[25143]_ ,
    \new_[25147]_ , \new_[25148]_ , \new_[25149]_ , \new_[25153]_ ,
    \new_[25154]_ , \new_[25158]_ , \new_[25159]_ , \new_[25160]_ ,
    \new_[25163]_ , \new_[25167]_ , \new_[25168]_ , \new_[25169]_ ,
    \new_[25173]_ , \new_[25174]_ , \new_[25178]_ , \new_[25179]_ ,
    \new_[25180]_ , \new_[25183]_ , \new_[25187]_ , \new_[25188]_ ,
    \new_[25189]_ , \new_[25193]_ , \new_[25194]_ , \new_[25198]_ ,
    \new_[25199]_ , \new_[25200]_ , \new_[25203]_ , \new_[25207]_ ,
    \new_[25208]_ , \new_[25209]_ , \new_[25213]_ , \new_[25214]_ ,
    \new_[25218]_ , \new_[25219]_ , \new_[25220]_ , \new_[25223]_ ,
    \new_[25227]_ , \new_[25228]_ , \new_[25229]_ , \new_[25233]_ ,
    \new_[25234]_ , \new_[25238]_ , \new_[25239]_ , \new_[25240]_ ,
    \new_[25243]_ , \new_[25247]_ , \new_[25248]_ , \new_[25249]_ ,
    \new_[25253]_ , \new_[25254]_ , \new_[25258]_ , \new_[25259]_ ,
    \new_[25260]_ , \new_[25263]_ , \new_[25267]_ , \new_[25268]_ ,
    \new_[25269]_ , \new_[25273]_ , \new_[25274]_ , \new_[25278]_ ,
    \new_[25279]_ , \new_[25280]_ , \new_[25283]_ , \new_[25287]_ ,
    \new_[25288]_ , \new_[25289]_ , \new_[25293]_ , \new_[25294]_ ,
    \new_[25298]_ , \new_[25299]_ , \new_[25300]_ , \new_[25303]_ ,
    \new_[25307]_ , \new_[25308]_ , \new_[25309]_ , \new_[25313]_ ,
    \new_[25314]_ , \new_[25318]_ , \new_[25319]_ , \new_[25320]_ ,
    \new_[25323]_ , \new_[25327]_ , \new_[25328]_ , \new_[25329]_ ,
    \new_[25333]_ , \new_[25334]_ , \new_[25338]_ , \new_[25339]_ ,
    \new_[25340]_ , \new_[25343]_ , \new_[25347]_ , \new_[25348]_ ,
    \new_[25349]_ , \new_[25353]_ , \new_[25354]_ , \new_[25358]_ ,
    \new_[25359]_ , \new_[25360]_ , \new_[25363]_ , \new_[25367]_ ,
    \new_[25368]_ , \new_[25369]_ , \new_[25373]_ , \new_[25374]_ ,
    \new_[25378]_ , \new_[25379]_ , \new_[25380]_ , \new_[25383]_ ,
    \new_[25387]_ , \new_[25388]_ , \new_[25389]_ , \new_[25393]_ ,
    \new_[25394]_ , \new_[25398]_ , \new_[25399]_ , \new_[25400]_ ,
    \new_[25403]_ , \new_[25407]_ , \new_[25408]_ , \new_[25409]_ ,
    \new_[25413]_ , \new_[25414]_ , \new_[25418]_ , \new_[25419]_ ,
    \new_[25420]_ , \new_[25423]_ , \new_[25427]_ , \new_[25428]_ ,
    \new_[25429]_ , \new_[25433]_ , \new_[25434]_ , \new_[25438]_ ,
    \new_[25439]_ , \new_[25440]_ , \new_[25443]_ , \new_[25447]_ ,
    \new_[25448]_ , \new_[25449]_ , \new_[25453]_ , \new_[25454]_ ,
    \new_[25458]_ , \new_[25459]_ , \new_[25460]_ , \new_[25463]_ ,
    \new_[25467]_ , \new_[25468]_ , \new_[25469]_ , \new_[25473]_ ,
    \new_[25474]_ , \new_[25478]_ , \new_[25479]_ , \new_[25480]_ ,
    \new_[25483]_ , \new_[25487]_ , \new_[25488]_ , \new_[25489]_ ,
    \new_[25493]_ , \new_[25494]_ , \new_[25498]_ , \new_[25499]_ ,
    \new_[25500]_ , \new_[25503]_ , \new_[25507]_ , \new_[25508]_ ,
    \new_[25509]_ , \new_[25513]_ , \new_[25514]_ , \new_[25518]_ ,
    \new_[25519]_ , \new_[25520]_ , \new_[25523]_ , \new_[25527]_ ,
    \new_[25528]_ , \new_[25529]_ , \new_[25533]_ , \new_[25534]_ ,
    \new_[25538]_ , \new_[25539]_ , \new_[25540]_ , \new_[25543]_ ,
    \new_[25547]_ , \new_[25548]_ , \new_[25549]_ , \new_[25553]_ ,
    \new_[25554]_ , \new_[25558]_ , \new_[25559]_ , \new_[25560]_ ,
    \new_[25563]_ , \new_[25567]_ , \new_[25568]_ , \new_[25569]_ ,
    \new_[25573]_ , \new_[25574]_ , \new_[25578]_ , \new_[25579]_ ,
    \new_[25580]_ , \new_[25583]_ , \new_[25587]_ , \new_[25588]_ ,
    \new_[25589]_ , \new_[25593]_ , \new_[25594]_ , \new_[25598]_ ,
    \new_[25599]_ , \new_[25600]_ , \new_[25603]_ , \new_[25607]_ ,
    \new_[25608]_ , \new_[25609]_ , \new_[25613]_ , \new_[25614]_ ,
    \new_[25618]_ , \new_[25619]_ , \new_[25620]_ , \new_[25623]_ ,
    \new_[25627]_ , \new_[25628]_ , \new_[25629]_ , \new_[25633]_ ,
    \new_[25634]_ , \new_[25638]_ , \new_[25639]_ , \new_[25640]_ ,
    \new_[25643]_ , \new_[25647]_ , \new_[25648]_ , \new_[25649]_ ,
    \new_[25653]_ , \new_[25654]_ , \new_[25658]_ , \new_[25659]_ ,
    \new_[25660]_ , \new_[25663]_ , \new_[25667]_ , \new_[25668]_ ,
    \new_[25669]_ , \new_[25673]_ , \new_[25674]_ , \new_[25678]_ ,
    \new_[25679]_ , \new_[25680]_ , \new_[25683]_ , \new_[25687]_ ,
    \new_[25688]_ , \new_[25689]_ , \new_[25693]_ , \new_[25694]_ ,
    \new_[25698]_ , \new_[25699]_ , \new_[25700]_ , \new_[25703]_ ,
    \new_[25707]_ , \new_[25708]_ , \new_[25709]_ , \new_[25713]_ ,
    \new_[25714]_ , \new_[25718]_ , \new_[25719]_ , \new_[25720]_ ,
    \new_[25723]_ , \new_[25727]_ , \new_[25728]_ , \new_[25729]_ ,
    \new_[25733]_ , \new_[25734]_ , \new_[25738]_ , \new_[25739]_ ,
    \new_[25740]_ , \new_[25743]_ , \new_[25747]_ , \new_[25748]_ ,
    \new_[25749]_ , \new_[25753]_ , \new_[25754]_ , \new_[25758]_ ,
    \new_[25759]_ , \new_[25760]_ , \new_[25763]_ , \new_[25767]_ ,
    \new_[25768]_ , \new_[25769]_ , \new_[25773]_ , \new_[25774]_ ,
    \new_[25778]_ , \new_[25779]_ , \new_[25780]_ , \new_[25783]_ ,
    \new_[25787]_ , \new_[25788]_ , \new_[25789]_ , \new_[25793]_ ,
    \new_[25794]_ , \new_[25798]_ , \new_[25799]_ , \new_[25800]_ ,
    \new_[25803]_ , \new_[25807]_ , \new_[25808]_ , \new_[25809]_ ,
    \new_[25813]_ , \new_[25814]_ , \new_[25818]_ , \new_[25819]_ ,
    \new_[25820]_ , \new_[25823]_ , \new_[25827]_ , \new_[25828]_ ,
    \new_[25829]_ , \new_[25833]_ , \new_[25834]_ , \new_[25838]_ ,
    \new_[25839]_ , \new_[25840]_ , \new_[25843]_ , \new_[25847]_ ,
    \new_[25848]_ , \new_[25849]_ , \new_[25853]_ , \new_[25854]_ ,
    \new_[25858]_ , \new_[25859]_ , \new_[25860]_ , \new_[25863]_ ,
    \new_[25867]_ , \new_[25868]_ , \new_[25869]_ , \new_[25873]_ ,
    \new_[25874]_ , \new_[25878]_ , \new_[25879]_ , \new_[25880]_ ,
    \new_[25883]_ , \new_[25887]_ , \new_[25888]_ , \new_[25889]_ ,
    \new_[25893]_ , \new_[25894]_ , \new_[25898]_ , \new_[25899]_ ,
    \new_[25900]_ , \new_[25903]_ , \new_[25907]_ , \new_[25908]_ ,
    \new_[25909]_ , \new_[25913]_ , \new_[25914]_ , \new_[25918]_ ,
    \new_[25919]_ , \new_[25920]_ , \new_[25923]_ , \new_[25927]_ ,
    \new_[25928]_ , \new_[25929]_ , \new_[25933]_ , \new_[25934]_ ,
    \new_[25938]_ , \new_[25939]_ , \new_[25940]_ , \new_[25943]_ ,
    \new_[25947]_ , \new_[25948]_ , \new_[25949]_ , \new_[25953]_ ,
    \new_[25954]_ , \new_[25958]_ , \new_[25959]_ , \new_[25960]_ ,
    \new_[25963]_ , \new_[25967]_ , \new_[25968]_ , \new_[25969]_ ,
    \new_[25973]_ , \new_[25974]_ , \new_[25978]_ , \new_[25979]_ ,
    \new_[25980]_ , \new_[25983]_ , \new_[25987]_ , \new_[25988]_ ,
    \new_[25989]_ , \new_[25993]_ , \new_[25994]_ , \new_[25998]_ ,
    \new_[25999]_ , \new_[26000]_ , \new_[26003]_ , \new_[26007]_ ,
    \new_[26008]_ , \new_[26009]_ , \new_[26013]_ , \new_[26014]_ ,
    \new_[26018]_ , \new_[26019]_ , \new_[26020]_ , \new_[26023]_ ,
    \new_[26027]_ , \new_[26028]_ , \new_[26029]_ , \new_[26033]_ ,
    \new_[26034]_ , \new_[26038]_ , \new_[26039]_ , \new_[26040]_ ,
    \new_[26043]_ , \new_[26047]_ , \new_[26048]_ , \new_[26049]_ ,
    \new_[26053]_ , \new_[26054]_ , \new_[26058]_ , \new_[26059]_ ,
    \new_[26060]_ , \new_[26063]_ , \new_[26067]_ , \new_[26068]_ ,
    \new_[26069]_ , \new_[26073]_ , \new_[26074]_ , \new_[26078]_ ,
    \new_[26079]_ , \new_[26080]_ , \new_[26083]_ , \new_[26087]_ ,
    \new_[26088]_ , \new_[26089]_ , \new_[26093]_ , \new_[26094]_ ,
    \new_[26098]_ , \new_[26099]_ , \new_[26100]_ , \new_[26103]_ ,
    \new_[26107]_ , \new_[26108]_ , \new_[26109]_ , \new_[26113]_ ,
    \new_[26114]_ , \new_[26118]_ , \new_[26119]_ , \new_[26120]_ ,
    \new_[26123]_ , \new_[26127]_ , \new_[26128]_ , \new_[26129]_ ,
    \new_[26133]_ , \new_[26134]_ , \new_[26138]_ , \new_[26139]_ ,
    \new_[26140]_ , \new_[26143]_ , \new_[26147]_ , \new_[26148]_ ,
    \new_[26149]_ , \new_[26153]_ , \new_[26154]_ , \new_[26158]_ ,
    \new_[26159]_ , \new_[26160]_ , \new_[26163]_ , \new_[26167]_ ,
    \new_[26168]_ , \new_[26169]_ , \new_[26173]_ , \new_[26174]_ ,
    \new_[26178]_ , \new_[26179]_ , \new_[26180]_ , \new_[26183]_ ,
    \new_[26187]_ , \new_[26188]_ , \new_[26189]_ , \new_[26193]_ ,
    \new_[26194]_ , \new_[26198]_ , \new_[26199]_ , \new_[26200]_ ,
    \new_[26203]_ , \new_[26207]_ , \new_[26208]_ , \new_[26209]_ ,
    \new_[26213]_ , \new_[26214]_ , \new_[26218]_ , \new_[26219]_ ,
    \new_[26220]_ , \new_[26223]_ , \new_[26227]_ , \new_[26228]_ ,
    \new_[26229]_ , \new_[26233]_ , \new_[26234]_ , \new_[26238]_ ,
    \new_[26239]_ , \new_[26240]_ , \new_[26243]_ , \new_[26247]_ ,
    \new_[26248]_ , \new_[26249]_ , \new_[26253]_ , \new_[26254]_ ,
    \new_[26258]_ , \new_[26259]_ , \new_[26260]_ , \new_[26263]_ ,
    \new_[26267]_ , \new_[26268]_ , \new_[26269]_ , \new_[26273]_ ,
    \new_[26274]_ , \new_[26278]_ , \new_[26279]_ , \new_[26280]_ ,
    \new_[26283]_ , \new_[26287]_ , \new_[26288]_ , \new_[26289]_ ,
    \new_[26293]_ , \new_[26294]_ , \new_[26298]_ , \new_[26299]_ ,
    \new_[26300]_ , \new_[26303]_ , \new_[26307]_ , \new_[26308]_ ,
    \new_[26309]_ , \new_[26313]_ , \new_[26314]_ , \new_[26318]_ ,
    \new_[26319]_ , \new_[26320]_ , \new_[26323]_ , \new_[26327]_ ,
    \new_[26328]_ , \new_[26329]_ , \new_[26333]_ , \new_[26334]_ ,
    \new_[26338]_ , \new_[26339]_ , \new_[26340]_ , \new_[26343]_ ,
    \new_[26347]_ , \new_[26348]_ , \new_[26349]_ , \new_[26353]_ ,
    \new_[26354]_ , \new_[26358]_ , \new_[26359]_ , \new_[26360]_ ,
    \new_[26363]_ , \new_[26367]_ , \new_[26368]_ , \new_[26369]_ ,
    \new_[26373]_ , \new_[26374]_ , \new_[26378]_ , \new_[26379]_ ,
    \new_[26380]_ , \new_[26383]_ , \new_[26387]_ , \new_[26388]_ ,
    \new_[26389]_ , \new_[26393]_ , \new_[26394]_ , \new_[26398]_ ,
    \new_[26399]_ , \new_[26400]_ , \new_[26403]_ , \new_[26407]_ ,
    \new_[26408]_ , \new_[26409]_ , \new_[26413]_ , \new_[26414]_ ,
    \new_[26418]_ , \new_[26419]_ , \new_[26420]_ , \new_[26423]_ ,
    \new_[26427]_ , \new_[26428]_ , \new_[26429]_ , \new_[26433]_ ,
    \new_[26434]_ , \new_[26438]_ , \new_[26439]_ , \new_[26440]_ ,
    \new_[26443]_ , \new_[26447]_ , \new_[26448]_ , \new_[26449]_ ,
    \new_[26453]_ , \new_[26454]_ , \new_[26458]_ , \new_[26459]_ ,
    \new_[26460]_ , \new_[26463]_ , \new_[26467]_ , \new_[26468]_ ,
    \new_[26469]_ , \new_[26473]_ , \new_[26474]_ , \new_[26478]_ ,
    \new_[26479]_ , \new_[26480]_ , \new_[26483]_ , \new_[26487]_ ,
    \new_[26488]_ , \new_[26489]_ , \new_[26493]_ , \new_[26494]_ ,
    \new_[26498]_ , \new_[26499]_ , \new_[26500]_ , \new_[26503]_ ,
    \new_[26507]_ , \new_[26508]_ , \new_[26509]_ , \new_[26513]_ ,
    \new_[26514]_ , \new_[26518]_ , \new_[26519]_ , \new_[26520]_ ,
    \new_[26523]_ , \new_[26527]_ , \new_[26528]_ , \new_[26529]_ ,
    \new_[26533]_ , \new_[26534]_ , \new_[26538]_ , \new_[26539]_ ,
    \new_[26540]_ , \new_[26543]_ , \new_[26547]_ , \new_[26548]_ ,
    \new_[26549]_ , \new_[26553]_ , \new_[26554]_ , \new_[26558]_ ,
    \new_[26559]_ , \new_[26560]_ , \new_[26563]_ , \new_[26567]_ ,
    \new_[26568]_ , \new_[26569]_ , \new_[26573]_ , \new_[26574]_ ,
    \new_[26578]_ , \new_[26579]_ , \new_[26580]_ , \new_[26583]_ ,
    \new_[26587]_ , \new_[26588]_ , \new_[26589]_ , \new_[26593]_ ,
    \new_[26594]_ , \new_[26598]_ , \new_[26599]_ , \new_[26600]_ ,
    \new_[26603]_ , \new_[26607]_ , \new_[26608]_ , \new_[26609]_ ,
    \new_[26613]_ , \new_[26614]_ , \new_[26618]_ , \new_[26619]_ ,
    \new_[26620]_ , \new_[26623]_ , \new_[26627]_ , \new_[26628]_ ,
    \new_[26629]_ , \new_[26633]_ , \new_[26634]_ , \new_[26638]_ ,
    \new_[26639]_ , \new_[26640]_ , \new_[26643]_ , \new_[26647]_ ,
    \new_[26648]_ , \new_[26649]_ , \new_[26653]_ , \new_[26654]_ ,
    \new_[26658]_ , \new_[26659]_ , \new_[26660]_ , \new_[26663]_ ,
    \new_[26667]_ , \new_[26668]_ , \new_[26669]_ , \new_[26673]_ ,
    \new_[26674]_ , \new_[26678]_ , \new_[26679]_ , \new_[26680]_ ,
    \new_[26683]_ , \new_[26687]_ , \new_[26688]_ , \new_[26689]_ ,
    \new_[26693]_ , \new_[26694]_ , \new_[26698]_ , \new_[26699]_ ,
    \new_[26700]_ , \new_[26703]_ , \new_[26707]_ , \new_[26708]_ ,
    \new_[26709]_ , \new_[26713]_ , \new_[26714]_ , \new_[26718]_ ,
    \new_[26719]_ , \new_[26720]_ , \new_[26723]_ , \new_[26727]_ ,
    \new_[26728]_ , \new_[26729]_ , \new_[26733]_ , \new_[26734]_ ,
    \new_[26738]_ , \new_[26739]_ , \new_[26740]_ , \new_[26743]_ ,
    \new_[26747]_ , \new_[26748]_ , \new_[26749]_ , \new_[26753]_ ,
    \new_[26754]_ , \new_[26758]_ , \new_[26759]_ , \new_[26760]_ ,
    \new_[26763]_ , \new_[26767]_ , \new_[26768]_ , \new_[26769]_ ,
    \new_[26773]_ , \new_[26774]_ , \new_[26778]_ , \new_[26779]_ ,
    \new_[26780]_ , \new_[26783]_ , \new_[26787]_ , \new_[26788]_ ,
    \new_[26789]_ , \new_[26793]_ , \new_[26794]_ , \new_[26798]_ ,
    \new_[26799]_ , \new_[26800]_ , \new_[26803]_ , \new_[26807]_ ,
    \new_[26808]_ , \new_[26809]_ , \new_[26813]_ , \new_[26814]_ ,
    \new_[26818]_ , \new_[26819]_ , \new_[26820]_ , \new_[26823]_ ,
    \new_[26827]_ , \new_[26828]_ , \new_[26829]_ , \new_[26833]_ ,
    \new_[26834]_ , \new_[26838]_ , \new_[26839]_ , \new_[26840]_ ,
    \new_[26843]_ , \new_[26847]_ , \new_[26848]_ , \new_[26849]_ ,
    \new_[26853]_ , \new_[26854]_ , \new_[26858]_ , \new_[26859]_ ,
    \new_[26860]_ , \new_[26863]_ , \new_[26867]_ , \new_[26868]_ ,
    \new_[26869]_ , \new_[26873]_ , \new_[26874]_ , \new_[26878]_ ,
    \new_[26879]_ , \new_[26880]_ , \new_[26883]_ , \new_[26887]_ ,
    \new_[26888]_ , \new_[26889]_ , \new_[26893]_ , \new_[26894]_ ,
    \new_[26898]_ , \new_[26899]_ , \new_[26900]_ , \new_[26903]_ ,
    \new_[26907]_ , \new_[26908]_ , \new_[26909]_ , \new_[26913]_ ,
    \new_[26914]_ , \new_[26918]_ , \new_[26919]_ , \new_[26920]_ ,
    \new_[26923]_ , \new_[26927]_ , \new_[26928]_ , \new_[26929]_ ,
    \new_[26933]_ , \new_[26934]_ , \new_[26938]_ , \new_[26939]_ ,
    \new_[26940]_ , \new_[26943]_ , \new_[26947]_ , \new_[26948]_ ,
    \new_[26949]_ , \new_[26953]_ , \new_[26954]_ , \new_[26958]_ ,
    \new_[26959]_ , \new_[26960]_ , \new_[26963]_ , \new_[26967]_ ,
    \new_[26968]_ , \new_[26969]_ , \new_[26973]_ , \new_[26974]_ ,
    \new_[26978]_ , \new_[26979]_ , \new_[26980]_ , \new_[26983]_ ,
    \new_[26987]_ , \new_[26988]_ , \new_[26989]_ , \new_[26993]_ ,
    \new_[26994]_ , \new_[26998]_ , \new_[26999]_ , \new_[27000]_ ,
    \new_[27003]_ , \new_[27007]_ , \new_[27008]_ , \new_[27009]_ ,
    \new_[27013]_ , \new_[27014]_ , \new_[27018]_ , \new_[27019]_ ,
    \new_[27020]_ , \new_[27023]_ , \new_[27027]_ , \new_[27028]_ ,
    \new_[27029]_ , \new_[27033]_ , \new_[27034]_ , \new_[27038]_ ,
    \new_[27039]_ , \new_[27040]_ , \new_[27043]_ , \new_[27047]_ ,
    \new_[27048]_ , \new_[27049]_ , \new_[27053]_ , \new_[27054]_ ,
    \new_[27058]_ , \new_[27059]_ , \new_[27060]_ , \new_[27063]_ ,
    \new_[27067]_ , \new_[27068]_ , \new_[27069]_ , \new_[27073]_ ,
    \new_[27074]_ , \new_[27078]_ , \new_[27079]_ , \new_[27080]_ ,
    \new_[27083]_ , \new_[27087]_ , \new_[27088]_ , \new_[27089]_ ,
    \new_[27093]_ , \new_[27094]_ , \new_[27098]_ , \new_[27099]_ ,
    \new_[27100]_ , \new_[27103]_ , \new_[27107]_ , \new_[27108]_ ,
    \new_[27109]_ , \new_[27113]_ , \new_[27114]_ , \new_[27118]_ ,
    \new_[27119]_ , \new_[27120]_ , \new_[27123]_ , \new_[27127]_ ,
    \new_[27128]_ , \new_[27129]_ , \new_[27133]_ , \new_[27134]_ ,
    \new_[27138]_ , \new_[27139]_ , \new_[27140]_ , \new_[27143]_ ,
    \new_[27147]_ , \new_[27148]_ , \new_[27149]_ , \new_[27153]_ ,
    \new_[27154]_ , \new_[27158]_ , \new_[27159]_ , \new_[27160]_ ,
    \new_[27163]_ , \new_[27167]_ , \new_[27168]_ , \new_[27169]_ ,
    \new_[27173]_ , \new_[27174]_ , \new_[27178]_ , \new_[27179]_ ,
    \new_[27180]_ , \new_[27183]_ , \new_[27187]_ , \new_[27188]_ ,
    \new_[27189]_ , \new_[27193]_ , \new_[27194]_ , \new_[27198]_ ,
    \new_[27199]_ , \new_[27200]_ , \new_[27203]_ , \new_[27207]_ ,
    \new_[27208]_ , \new_[27209]_ , \new_[27213]_ , \new_[27214]_ ,
    \new_[27218]_ , \new_[27219]_ , \new_[27220]_ , \new_[27223]_ ,
    \new_[27227]_ , \new_[27228]_ , \new_[27229]_ , \new_[27233]_ ,
    \new_[27234]_ , \new_[27238]_ , \new_[27239]_ , \new_[27240]_ ,
    \new_[27243]_ , \new_[27247]_ , \new_[27248]_ , \new_[27249]_ ,
    \new_[27253]_ , \new_[27254]_ , \new_[27258]_ , \new_[27259]_ ,
    \new_[27260]_ , \new_[27263]_ , \new_[27267]_ , \new_[27268]_ ,
    \new_[27269]_ , \new_[27273]_ , \new_[27274]_ , \new_[27278]_ ,
    \new_[27279]_ , \new_[27280]_ , \new_[27283]_ , \new_[27287]_ ,
    \new_[27288]_ , \new_[27289]_ , \new_[27293]_ , \new_[27294]_ ,
    \new_[27298]_ , \new_[27299]_ , \new_[27300]_ , \new_[27303]_ ,
    \new_[27307]_ , \new_[27308]_ , \new_[27309]_ , \new_[27313]_ ,
    \new_[27314]_ , \new_[27318]_ , \new_[27319]_ , \new_[27320]_ ,
    \new_[27323]_ , \new_[27327]_ , \new_[27328]_ , \new_[27329]_ ,
    \new_[27333]_ , \new_[27334]_ , \new_[27338]_ , \new_[27339]_ ,
    \new_[27340]_ , \new_[27343]_ , \new_[27347]_ , \new_[27348]_ ,
    \new_[27349]_ , \new_[27353]_ , \new_[27354]_ , \new_[27358]_ ,
    \new_[27359]_ , \new_[27360]_ , \new_[27363]_ , \new_[27367]_ ,
    \new_[27368]_ , \new_[27369]_ , \new_[27373]_ , \new_[27374]_ ,
    \new_[27378]_ , \new_[27379]_ , \new_[27380]_ , \new_[27383]_ ,
    \new_[27387]_ , \new_[27388]_ , \new_[27389]_ , \new_[27393]_ ,
    \new_[27394]_ , \new_[27398]_ , \new_[27399]_ , \new_[27400]_ ,
    \new_[27403]_ , \new_[27407]_ , \new_[27408]_ , \new_[27409]_ ,
    \new_[27413]_ , \new_[27414]_ , \new_[27418]_ , \new_[27419]_ ,
    \new_[27420]_ , \new_[27423]_ , \new_[27427]_ , \new_[27428]_ ,
    \new_[27429]_ , \new_[27433]_ , \new_[27434]_ , \new_[27438]_ ,
    \new_[27439]_ , \new_[27440]_ , \new_[27443]_ , \new_[27447]_ ,
    \new_[27448]_ , \new_[27449]_ , \new_[27453]_ , \new_[27454]_ ,
    \new_[27458]_ , \new_[27459]_ , \new_[27460]_ , \new_[27463]_ ,
    \new_[27467]_ , \new_[27468]_ , \new_[27469]_ , \new_[27473]_ ,
    \new_[27474]_ , \new_[27478]_ , \new_[27479]_ , \new_[27480]_ ,
    \new_[27483]_ , \new_[27487]_ , \new_[27488]_ , \new_[27489]_ ,
    \new_[27493]_ , \new_[27494]_ , \new_[27498]_ , \new_[27499]_ ,
    \new_[27500]_ , \new_[27503]_ , \new_[27507]_ , \new_[27508]_ ,
    \new_[27509]_ , \new_[27513]_ , \new_[27514]_ , \new_[27518]_ ,
    \new_[27519]_ , \new_[27520]_ , \new_[27523]_ , \new_[27527]_ ,
    \new_[27528]_ , \new_[27529]_ , \new_[27533]_ , \new_[27534]_ ,
    \new_[27538]_ , \new_[27539]_ , \new_[27540]_ , \new_[27543]_ ,
    \new_[27547]_ , \new_[27548]_ , \new_[27549]_ , \new_[27553]_ ,
    \new_[27554]_ , \new_[27558]_ , \new_[27559]_ , \new_[27560]_ ,
    \new_[27563]_ , \new_[27567]_ , \new_[27568]_ , \new_[27569]_ ,
    \new_[27573]_ , \new_[27574]_ , \new_[27578]_ , \new_[27579]_ ,
    \new_[27580]_ , \new_[27583]_ , \new_[27587]_ , \new_[27588]_ ,
    \new_[27589]_ , \new_[27593]_ , \new_[27594]_ , \new_[27598]_ ,
    \new_[27599]_ , \new_[27600]_ , \new_[27603]_ , \new_[27607]_ ,
    \new_[27608]_ , \new_[27609]_ , \new_[27613]_ , \new_[27614]_ ,
    \new_[27618]_ , \new_[27619]_ , \new_[27620]_ , \new_[27623]_ ,
    \new_[27627]_ , \new_[27628]_ , \new_[27629]_ , \new_[27633]_ ,
    \new_[27634]_ , \new_[27638]_ , \new_[27639]_ , \new_[27640]_ ,
    \new_[27643]_ , \new_[27647]_ , \new_[27648]_ , \new_[27649]_ ,
    \new_[27653]_ , \new_[27654]_ , \new_[27658]_ , \new_[27659]_ ,
    \new_[27660]_ , \new_[27663]_ , \new_[27667]_ , \new_[27668]_ ,
    \new_[27669]_ , \new_[27673]_ , \new_[27674]_ , \new_[27678]_ ,
    \new_[27679]_ , \new_[27680]_ , \new_[27683]_ , \new_[27687]_ ,
    \new_[27688]_ , \new_[27689]_ , \new_[27693]_ , \new_[27694]_ ,
    \new_[27698]_ , \new_[27699]_ , \new_[27700]_ , \new_[27703]_ ,
    \new_[27707]_ , \new_[27708]_ , \new_[27709]_ , \new_[27713]_ ,
    \new_[27714]_ , \new_[27718]_ , \new_[27719]_ , \new_[27720]_ ,
    \new_[27723]_ , \new_[27727]_ , \new_[27728]_ , \new_[27729]_ ,
    \new_[27733]_ , \new_[27734]_ , \new_[27738]_ , \new_[27739]_ ,
    \new_[27740]_ , \new_[27743]_ , \new_[27747]_ , \new_[27748]_ ,
    \new_[27749]_ , \new_[27753]_ , \new_[27754]_ , \new_[27758]_ ,
    \new_[27759]_ , \new_[27760]_ , \new_[27763]_ , \new_[27767]_ ,
    \new_[27768]_ , \new_[27769]_ , \new_[27773]_ , \new_[27774]_ ,
    \new_[27778]_ , \new_[27779]_ , \new_[27780]_ , \new_[27783]_ ,
    \new_[27787]_ , \new_[27788]_ , \new_[27789]_ , \new_[27793]_ ,
    \new_[27794]_ , \new_[27798]_ , \new_[27799]_ , \new_[27800]_ ,
    \new_[27803]_ , \new_[27807]_ , \new_[27808]_ , \new_[27809]_ ,
    \new_[27813]_ , \new_[27814]_ , \new_[27818]_ , \new_[27819]_ ,
    \new_[27820]_ , \new_[27823]_ , \new_[27827]_ , \new_[27828]_ ,
    \new_[27829]_ , \new_[27833]_ , \new_[27834]_ , \new_[27838]_ ,
    \new_[27839]_ , \new_[27840]_ , \new_[27843]_ , \new_[27847]_ ,
    \new_[27848]_ , \new_[27849]_ , \new_[27853]_ , \new_[27854]_ ,
    \new_[27858]_ , \new_[27859]_ , \new_[27860]_ , \new_[27863]_ ,
    \new_[27867]_ , \new_[27868]_ , \new_[27869]_ , \new_[27873]_ ,
    \new_[27874]_ , \new_[27878]_ , \new_[27879]_ , \new_[27880]_ ,
    \new_[27883]_ , \new_[27887]_ , \new_[27888]_ , \new_[27889]_ ,
    \new_[27893]_ , \new_[27894]_ , \new_[27898]_ , \new_[27899]_ ,
    \new_[27900]_ , \new_[27903]_ , \new_[27907]_ , \new_[27908]_ ,
    \new_[27909]_ , \new_[27913]_ , \new_[27914]_ , \new_[27918]_ ,
    \new_[27919]_ , \new_[27920]_ , \new_[27923]_ , \new_[27927]_ ,
    \new_[27928]_ , \new_[27929]_ , \new_[27933]_ , \new_[27934]_ ,
    \new_[27938]_ , \new_[27939]_ , \new_[27940]_ , \new_[27943]_ ,
    \new_[27947]_ , \new_[27948]_ , \new_[27949]_ , \new_[27953]_ ,
    \new_[27954]_ , \new_[27958]_ , \new_[27959]_ , \new_[27960]_ ,
    \new_[27963]_ , \new_[27967]_ , \new_[27968]_ , \new_[27969]_ ,
    \new_[27973]_ , \new_[27974]_ , \new_[27978]_ , \new_[27979]_ ,
    \new_[27980]_ , \new_[27983]_ , \new_[27987]_ , \new_[27988]_ ,
    \new_[27989]_ , \new_[27993]_ , \new_[27994]_ , \new_[27998]_ ,
    \new_[27999]_ , \new_[28000]_ , \new_[28003]_ , \new_[28007]_ ,
    \new_[28008]_ , \new_[28009]_ , \new_[28013]_ , \new_[28014]_ ,
    \new_[28018]_ , \new_[28019]_ , \new_[28020]_ , \new_[28023]_ ,
    \new_[28027]_ , \new_[28028]_ , \new_[28029]_ , \new_[28033]_ ,
    \new_[28034]_ , \new_[28038]_ , \new_[28039]_ , \new_[28040]_ ,
    \new_[28043]_ , \new_[28047]_ , \new_[28048]_ , \new_[28049]_ ,
    \new_[28053]_ , \new_[28054]_ , \new_[28058]_ , \new_[28059]_ ,
    \new_[28060]_ , \new_[28063]_ , \new_[28067]_ , \new_[28068]_ ,
    \new_[28069]_ , \new_[28073]_ , \new_[28074]_ , \new_[28078]_ ,
    \new_[28079]_ , \new_[28080]_ , \new_[28083]_ , \new_[28087]_ ,
    \new_[28088]_ , \new_[28089]_ , \new_[28093]_ , \new_[28094]_ ,
    \new_[28098]_ , \new_[28099]_ , \new_[28100]_ , \new_[28103]_ ,
    \new_[28107]_ , \new_[28108]_ , \new_[28109]_ , \new_[28113]_ ,
    \new_[28114]_ , \new_[28118]_ , \new_[28119]_ , \new_[28120]_ ,
    \new_[28123]_ , \new_[28127]_ , \new_[28128]_ , \new_[28129]_ ,
    \new_[28133]_ , \new_[28134]_ , \new_[28138]_ , \new_[28139]_ ,
    \new_[28140]_ , \new_[28143]_ , \new_[28147]_ , \new_[28148]_ ,
    \new_[28149]_ , \new_[28153]_ , \new_[28154]_ , \new_[28158]_ ,
    \new_[28159]_ , \new_[28160]_ , \new_[28163]_ , \new_[28167]_ ,
    \new_[28168]_ , \new_[28169]_ , \new_[28173]_ , \new_[28174]_ ,
    \new_[28178]_ , \new_[28179]_ , \new_[28180]_ , \new_[28183]_ ,
    \new_[28187]_ , \new_[28188]_ , \new_[28189]_ , \new_[28193]_ ,
    \new_[28194]_ , \new_[28198]_ , \new_[28199]_ , \new_[28200]_ ,
    \new_[28203]_ , \new_[28207]_ , \new_[28208]_ , \new_[28209]_ ,
    \new_[28213]_ , \new_[28214]_ , \new_[28218]_ , \new_[28219]_ ,
    \new_[28220]_ , \new_[28223]_ , \new_[28227]_ , \new_[28228]_ ,
    \new_[28229]_ , \new_[28233]_ , \new_[28234]_ , \new_[28238]_ ,
    \new_[28239]_ , \new_[28240]_ , \new_[28243]_ , \new_[28247]_ ,
    \new_[28248]_ , \new_[28249]_ , \new_[28253]_ , \new_[28254]_ ,
    \new_[28258]_ , \new_[28259]_ , \new_[28260]_ , \new_[28263]_ ,
    \new_[28267]_ , \new_[28268]_ , \new_[28269]_ , \new_[28273]_ ,
    \new_[28274]_ , \new_[28278]_ , \new_[28279]_ , \new_[28280]_ ,
    \new_[28283]_ , \new_[28287]_ , \new_[28288]_ , \new_[28289]_ ,
    \new_[28293]_ , \new_[28294]_ , \new_[28298]_ , \new_[28299]_ ,
    \new_[28300]_ , \new_[28303]_ , \new_[28307]_ , \new_[28308]_ ,
    \new_[28309]_ , \new_[28313]_ , \new_[28314]_ , \new_[28318]_ ,
    \new_[28319]_ , \new_[28320]_ , \new_[28323]_ , \new_[28327]_ ,
    \new_[28328]_ , \new_[28329]_ , \new_[28333]_ , \new_[28334]_ ,
    \new_[28338]_ , \new_[28339]_ , \new_[28340]_ , \new_[28343]_ ,
    \new_[28347]_ , \new_[28348]_ , \new_[28349]_ , \new_[28353]_ ,
    \new_[28354]_ , \new_[28358]_ , \new_[28359]_ , \new_[28360]_ ,
    \new_[28363]_ , \new_[28367]_ , \new_[28368]_ , \new_[28369]_ ,
    \new_[28373]_ , \new_[28374]_ , \new_[28378]_ , \new_[28379]_ ,
    \new_[28380]_ , \new_[28383]_ , \new_[28387]_ , \new_[28388]_ ,
    \new_[28389]_ , \new_[28393]_ , \new_[28394]_ , \new_[28398]_ ,
    \new_[28399]_ , \new_[28400]_ , \new_[28403]_ , \new_[28407]_ ,
    \new_[28408]_ , \new_[28409]_ , \new_[28413]_ , \new_[28414]_ ,
    \new_[28418]_ , \new_[28419]_ , \new_[28420]_ , \new_[28423]_ ,
    \new_[28427]_ , \new_[28428]_ , \new_[28429]_ , \new_[28433]_ ,
    \new_[28434]_ , \new_[28438]_ , \new_[28439]_ , \new_[28440]_ ,
    \new_[28443]_ , \new_[28447]_ , \new_[28448]_ , \new_[28449]_ ,
    \new_[28453]_ , \new_[28454]_ , \new_[28458]_ , \new_[28459]_ ,
    \new_[28460]_ , \new_[28463]_ , \new_[28467]_ , \new_[28468]_ ,
    \new_[28469]_ , \new_[28473]_ , \new_[28474]_ , \new_[28478]_ ,
    \new_[28479]_ , \new_[28480]_ , \new_[28483]_ , \new_[28487]_ ,
    \new_[28488]_ , \new_[28489]_ , \new_[28493]_ , \new_[28494]_ ,
    \new_[28498]_ , \new_[28499]_ , \new_[28500]_ , \new_[28503]_ ,
    \new_[28507]_ , \new_[28508]_ , \new_[28509]_ , \new_[28513]_ ,
    \new_[28514]_ , \new_[28518]_ , \new_[28519]_ , \new_[28520]_ ,
    \new_[28523]_ , \new_[28527]_ , \new_[28528]_ , \new_[28529]_ ,
    \new_[28533]_ , \new_[28534]_ , \new_[28538]_ , \new_[28539]_ ,
    \new_[28540]_ , \new_[28543]_ , \new_[28547]_ , \new_[28548]_ ,
    \new_[28549]_ , \new_[28553]_ , \new_[28554]_ , \new_[28558]_ ,
    \new_[28559]_ , \new_[28560]_ , \new_[28563]_ , \new_[28567]_ ,
    \new_[28568]_ , \new_[28569]_ , \new_[28573]_ , \new_[28574]_ ,
    \new_[28578]_ , \new_[28579]_ , \new_[28580]_ , \new_[28583]_ ,
    \new_[28587]_ , \new_[28588]_ , \new_[28589]_ , \new_[28593]_ ,
    \new_[28594]_ , \new_[28598]_ , \new_[28599]_ , \new_[28600]_ ,
    \new_[28603]_ , \new_[28607]_ , \new_[28608]_ , \new_[28609]_ ,
    \new_[28613]_ , \new_[28614]_ , \new_[28618]_ , \new_[28619]_ ,
    \new_[28620]_ , \new_[28623]_ , \new_[28627]_ , \new_[28628]_ ,
    \new_[28629]_ , \new_[28633]_ , \new_[28634]_ , \new_[28638]_ ,
    \new_[28639]_ , \new_[28640]_ , \new_[28643]_ , \new_[28647]_ ,
    \new_[28648]_ , \new_[28649]_ , \new_[28653]_ , \new_[28654]_ ,
    \new_[28658]_ , \new_[28659]_ , \new_[28660]_ , \new_[28663]_ ,
    \new_[28667]_ , \new_[28668]_ , \new_[28669]_ , \new_[28673]_ ,
    \new_[28674]_ , \new_[28678]_ , \new_[28679]_ , \new_[28680]_ ,
    \new_[28683]_ , \new_[28687]_ , \new_[28688]_ , \new_[28689]_ ,
    \new_[28693]_ , \new_[28694]_ , \new_[28698]_ , \new_[28699]_ ,
    \new_[28700]_ , \new_[28703]_ , \new_[28707]_ , \new_[28708]_ ,
    \new_[28709]_ , \new_[28713]_ , \new_[28714]_ , \new_[28718]_ ,
    \new_[28719]_ , \new_[28720]_ , \new_[28723]_ , \new_[28727]_ ,
    \new_[28728]_ , \new_[28729]_ , \new_[28733]_ , \new_[28734]_ ,
    \new_[28738]_ , \new_[28739]_ , \new_[28740]_ , \new_[28743]_ ,
    \new_[28747]_ , \new_[28748]_ , \new_[28749]_ , \new_[28753]_ ,
    \new_[28754]_ , \new_[28758]_ , \new_[28759]_ , \new_[28760]_ ,
    \new_[28763]_ , \new_[28767]_ , \new_[28768]_ , \new_[28769]_ ,
    \new_[28773]_ , \new_[28774]_ , \new_[28778]_ , \new_[28779]_ ,
    \new_[28780]_ , \new_[28783]_ , \new_[28787]_ , \new_[28788]_ ,
    \new_[28789]_ , \new_[28793]_ , \new_[28794]_ , \new_[28798]_ ,
    \new_[28799]_ , \new_[28800]_ , \new_[28803]_ , \new_[28807]_ ,
    \new_[28808]_ , \new_[28809]_ , \new_[28813]_ , \new_[28814]_ ,
    \new_[28818]_ , \new_[28819]_ , \new_[28820]_ , \new_[28823]_ ,
    \new_[28827]_ , \new_[28828]_ , \new_[28829]_ , \new_[28833]_ ,
    \new_[28834]_ , \new_[28838]_ , \new_[28839]_ , \new_[28840]_ ,
    \new_[28843]_ , \new_[28847]_ , \new_[28848]_ , \new_[28849]_ ,
    \new_[28853]_ , \new_[28854]_ , \new_[28858]_ , \new_[28859]_ ,
    \new_[28860]_ , \new_[28863]_ , \new_[28867]_ , \new_[28868]_ ,
    \new_[28869]_ , \new_[28873]_ , \new_[28874]_ , \new_[28878]_ ,
    \new_[28879]_ , \new_[28880]_ , \new_[28883]_ , \new_[28887]_ ,
    \new_[28888]_ , \new_[28889]_ , \new_[28893]_ , \new_[28894]_ ,
    \new_[28898]_ , \new_[28899]_ , \new_[28900]_ , \new_[28903]_ ,
    \new_[28907]_ , \new_[28908]_ , \new_[28909]_ , \new_[28913]_ ,
    \new_[28914]_ , \new_[28918]_ , \new_[28919]_ , \new_[28920]_ ,
    \new_[28923]_ , \new_[28927]_ , \new_[28928]_ , \new_[28929]_ ,
    \new_[28933]_ , \new_[28934]_ , \new_[28938]_ , \new_[28939]_ ,
    \new_[28940]_ , \new_[28943]_ , \new_[28947]_ , \new_[28948]_ ,
    \new_[28949]_ , \new_[28953]_ , \new_[28954]_ , \new_[28958]_ ,
    \new_[28959]_ , \new_[28960]_ , \new_[28963]_ , \new_[28967]_ ,
    \new_[28968]_ , \new_[28969]_ , \new_[28973]_ , \new_[28974]_ ,
    \new_[28978]_ , \new_[28979]_ , \new_[28980]_ , \new_[28983]_ ,
    \new_[28987]_ , \new_[28988]_ , \new_[28989]_ , \new_[28993]_ ,
    \new_[28994]_ , \new_[28998]_ , \new_[28999]_ , \new_[29000]_ ,
    \new_[29003]_ , \new_[29007]_ , \new_[29008]_ , \new_[29009]_ ,
    \new_[29013]_ , \new_[29014]_ , \new_[29018]_ , \new_[29019]_ ,
    \new_[29020]_ , \new_[29023]_ , \new_[29027]_ , \new_[29028]_ ,
    \new_[29029]_ , \new_[29033]_ , \new_[29034]_ , \new_[29038]_ ,
    \new_[29039]_ , \new_[29040]_ , \new_[29043]_ , \new_[29047]_ ,
    \new_[29048]_ , \new_[29049]_ , \new_[29053]_ , \new_[29054]_ ,
    \new_[29058]_ , \new_[29059]_ , \new_[29060]_ , \new_[29063]_ ,
    \new_[29067]_ , \new_[29068]_ , \new_[29069]_ , \new_[29073]_ ,
    \new_[29074]_ , \new_[29078]_ , \new_[29079]_ , \new_[29080]_ ,
    \new_[29083]_ , \new_[29087]_ , \new_[29088]_ , \new_[29089]_ ,
    \new_[29093]_ , \new_[29094]_ , \new_[29098]_ , \new_[29099]_ ,
    \new_[29100]_ , \new_[29103]_ , \new_[29107]_ , \new_[29108]_ ,
    \new_[29109]_ , \new_[29113]_ , \new_[29114]_ , \new_[29118]_ ,
    \new_[29119]_ , \new_[29120]_ , \new_[29123]_ , \new_[29127]_ ,
    \new_[29128]_ , \new_[29129]_ , \new_[29133]_ , \new_[29134]_ ,
    \new_[29138]_ , \new_[29139]_ , \new_[29140]_ , \new_[29143]_ ,
    \new_[29147]_ , \new_[29148]_ , \new_[29149]_ , \new_[29153]_ ,
    \new_[29154]_ , \new_[29158]_ , \new_[29159]_ , \new_[29160]_ ,
    \new_[29163]_ , \new_[29167]_ , \new_[29168]_ , \new_[29169]_ ,
    \new_[29173]_ , \new_[29174]_ , \new_[29178]_ , \new_[29179]_ ,
    \new_[29180]_ , \new_[29183]_ , \new_[29187]_ , \new_[29188]_ ,
    \new_[29189]_ , \new_[29193]_ , \new_[29194]_ , \new_[29198]_ ,
    \new_[29199]_ , \new_[29200]_ , \new_[29203]_ , \new_[29207]_ ,
    \new_[29208]_ , \new_[29209]_ , \new_[29213]_ , \new_[29214]_ ,
    \new_[29218]_ , \new_[29219]_ , \new_[29220]_ , \new_[29223]_ ,
    \new_[29227]_ , \new_[29228]_ , \new_[29229]_ , \new_[29233]_ ,
    \new_[29234]_ , \new_[29238]_ , \new_[29239]_ , \new_[29240]_ ,
    \new_[29243]_ , \new_[29247]_ , \new_[29248]_ , \new_[29249]_ ,
    \new_[29253]_ , \new_[29254]_ , \new_[29258]_ , \new_[29259]_ ,
    \new_[29260]_ , \new_[29263]_ , \new_[29267]_ , \new_[29268]_ ,
    \new_[29269]_ , \new_[29273]_ , \new_[29274]_ , \new_[29278]_ ,
    \new_[29279]_ , \new_[29280]_ , \new_[29283]_ , \new_[29287]_ ,
    \new_[29288]_ , \new_[29289]_ , \new_[29293]_ , \new_[29294]_ ,
    \new_[29298]_ , \new_[29299]_ , \new_[29300]_ , \new_[29303]_ ,
    \new_[29307]_ , \new_[29308]_ , \new_[29309]_ , \new_[29313]_ ,
    \new_[29314]_ , \new_[29318]_ , \new_[29319]_ , \new_[29320]_ ,
    \new_[29323]_ , \new_[29327]_ , \new_[29328]_ , \new_[29329]_ ,
    \new_[29333]_ , \new_[29334]_ , \new_[29338]_ , \new_[29339]_ ,
    \new_[29340]_ , \new_[29343]_ , \new_[29347]_ , \new_[29348]_ ,
    \new_[29349]_ , \new_[29353]_ , \new_[29354]_ , \new_[29358]_ ,
    \new_[29359]_ , \new_[29360]_ , \new_[29363]_ , \new_[29367]_ ,
    \new_[29368]_ , \new_[29369]_ , \new_[29373]_ , \new_[29374]_ ,
    \new_[29378]_ , \new_[29379]_ , \new_[29380]_ , \new_[29383]_ ,
    \new_[29387]_ , \new_[29388]_ , \new_[29389]_ , \new_[29393]_ ,
    \new_[29394]_ , \new_[29398]_ , \new_[29399]_ , \new_[29400]_ ,
    \new_[29403]_ , \new_[29407]_ , \new_[29408]_ , \new_[29409]_ ,
    \new_[29413]_ , \new_[29414]_ , \new_[29418]_ , \new_[29419]_ ,
    \new_[29420]_ , \new_[29423]_ , \new_[29427]_ , \new_[29428]_ ,
    \new_[29429]_ , \new_[29433]_ , \new_[29434]_ , \new_[29438]_ ,
    \new_[29439]_ , \new_[29440]_ , \new_[29444]_ , \new_[29445]_ ,
    \new_[29449]_ , \new_[29450]_ , \new_[29451]_ , \new_[29455]_ ,
    \new_[29456]_ , \new_[29460]_ , \new_[29461]_ , \new_[29462]_ ,
    \new_[29466]_ , \new_[29467]_ , \new_[29471]_ , \new_[29472]_ ,
    \new_[29473]_ , \new_[29477]_ , \new_[29478]_ , \new_[29482]_ ,
    \new_[29483]_ , \new_[29484]_ , \new_[29488]_ , \new_[29489]_ ,
    \new_[29493]_ , \new_[29494]_ , \new_[29495]_ , \new_[29499]_ ,
    \new_[29500]_ , \new_[29504]_ , \new_[29505]_ , \new_[29506]_ ,
    \new_[29510]_ , \new_[29511]_ , \new_[29515]_ , \new_[29516]_ ,
    \new_[29517]_ , \new_[29521]_ , \new_[29522]_ , \new_[29526]_ ,
    \new_[29527]_ , \new_[29528]_ , \new_[29532]_ , \new_[29533]_ ,
    \new_[29537]_ , \new_[29538]_ , \new_[29539]_ , \new_[29543]_ ,
    \new_[29544]_ , \new_[29548]_ , \new_[29549]_ , \new_[29550]_ ,
    \new_[29554]_ , \new_[29555]_ , \new_[29559]_ , \new_[29560]_ ,
    \new_[29561]_ , \new_[29565]_ , \new_[29566]_ , \new_[29570]_ ,
    \new_[29571]_ , \new_[29572]_ , \new_[29576]_ , \new_[29577]_ ,
    \new_[29581]_ , \new_[29582]_ , \new_[29583]_ , \new_[29587]_ ,
    \new_[29588]_ , \new_[29592]_ , \new_[29593]_ , \new_[29594]_ ,
    \new_[29598]_ , \new_[29599]_ , \new_[29603]_ , \new_[29604]_ ,
    \new_[29605]_ , \new_[29609]_ , \new_[29610]_ , \new_[29614]_ ,
    \new_[29615]_ , \new_[29616]_ , \new_[29620]_ , \new_[29621]_ ,
    \new_[29625]_ , \new_[29626]_ , \new_[29627]_ , \new_[29631]_ ,
    \new_[29632]_ , \new_[29636]_ , \new_[29637]_ , \new_[29638]_ ,
    \new_[29642]_ , \new_[29643]_ , \new_[29647]_ , \new_[29648]_ ,
    \new_[29649]_ , \new_[29653]_ , \new_[29654]_ , \new_[29658]_ ,
    \new_[29659]_ , \new_[29660]_ , \new_[29664]_ , \new_[29665]_ ,
    \new_[29669]_ , \new_[29670]_ , \new_[29671]_ , \new_[29675]_ ,
    \new_[29676]_ , \new_[29680]_ , \new_[29681]_ , \new_[29682]_ ,
    \new_[29686]_ , \new_[29687]_ , \new_[29691]_ , \new_[29692]_ ,
    \new_[29693]_ , \new_[29697]_ , \new_[29698]_ , \new_[29702]_ ,
    \new_[29703]_ , \new_[29704]_ , \new_[29708]_ , \new_[29709]_ ,
    \new_[29713]_ , \new_[29714]_ , \new_[29715]_ , \new_[29719]_ ,
    \new_[29720]_ , \new_[29724]_ , \new_[29725]_ , \new_[29726]_ ,
    \new_[29730]_ , \new_[29731]_ , \new_[29735]_ , \new_[29736]_ ,
    \new_[29737]_ , \new_[29741]_ , \new_[29742]_ , \new_[29746]_ ,
    \new_[29747]_ , \new_[29748]_ , \new_[29752]_ , \new_[29753]_ ,
    \new_[29757]_ , \new_[29758]_ , \new_[29759]_ , \new_[29763]_ ,
    \new_[29764]_ , \new_[29768]_ , \new_[29769]_ , \new_[29770]_ ,
    \new_[29774]_ , \new_[29775]_ , \new_[29779]_ , \new_[29780]_ ,
    \new_[29781]_ , \new_[29785]_ , \new_[29786]_ , \new_[29790]_ ,
    \new_[29791]_ , \new_[29792]_ , \new_[29796]_ , \new_[29797]_ ,
    \new_[29801]_ , \new_[29802]_ , \new_[29803]_ , \new_[29807]_ ,
    \new_[29808]_ , \new_[29812]_ , \new_[29813]_ , \new_[29814]_ ,
    \new_[29818]_ , \new_[29819]_ , \new_[29823]_ , \new_[29824]_ ,
    \new_[29825]_ , \new_[29829]_ , \new_[29830]_ , \new_[29834]_ ,
    \new_[29835]_ , \new_[29836]_ , \new_[29840]_ , \new_[29841]_ ,
    \new_[29845]_ , \new_[29846]_ , \new_[29847]_ , \new_[29851]_ ,
    \new_[29852]_ , \new_[29856]_ , \new_[29857]_ , \new_[29858]_ ,
    \new_[29862]_ , \new_[29863]_ , \new_[29867]_ , \new_[29868]_ ,
    \new_[29869]_ , \new_[29873]_ , \new_[29874]_ , \new_[29878]_ ,
    \new_[29879]_ , \new_[29880]_ , \new_[29884]_ , \new_[29885]_ ,
    \new_[29889]_ , \new_[29890]_ , \new_[29891]_ , \new_[29895]_ ,
    \new_[29896]_ , \new_[29900]_ , \new_[29901]_ , \new_[29902]_ ,
    \new_[29906]_ , \new_[29907]_ , \new_[29911]_ , \new_[29912]_ ,
    \new_[29913]_ , \new_[29917]_ , \new_[29918]_ , \new_[29922]_ ,
    \new_[29923]_ , \new_[29924]_ , \new_[29928]_ , \new_[29929]_ ,
    \new_[29933]_ , \new_[29934]_ , \new_[29935]_ , \new_[29939]_ ,
    \new_[29940]_ , \new_[29944]_ , \new_[29945]_ , \new_[29946]_ ,
    \new_[29950]_ , \new_[29951]_ , \new_[29955]_ , \new_[29956]_ ,
    \new_[29957]_ , \new_[29961]_ , \new_[29962]_ , \new_[29966]_ ,
    \new_[29967]_ , \new_[29968]_ , \new_[29972]_ , \new_[29973]_ ,
    \new_[29977]_ , \new_[29978]_ , \new_[29979]_ , \new_[29983]_ ,
    \new_[29984]_ , \new_[29988]_ , \new_[29989]_ , \new_[29990]_ ,
    \new_[29994]_ , \new_[29995]_ , \new_[29999]_ , \new_[30000]_ ,
    \new_[30001]_ , \new_[30005]_ , \new_[30006]_ , \new_[30010]_ ,
    \new_[30011]_ , \new_[30012]_ , \new_[30016]_ , \new_[30017]_ ,
    \new_[30021]_ , \new_[30022]_ , \new_[30023]_ , \new_[30027]_ ,
    \new_[30028]_ , \new_[30032]_ , \new_[30033]_ , \new_[30034]_ ,
    \new_[30038]_ , \new_[30039]_ , \new_[30043]_ , \new_[30044]_ ,
    \new_[30045]_ , \new_[30049]_ , \new_[30050]_ , \new_[30054]_ ,
    \new_[30055]_ , \new_[30056]_ , \new_[30060]_ , \new_[30061]_ ,
    \new_[30065]_ , \new_[30066]_ , \new_[30067]_ , \new_[30071]_ ,
    \new_[30072]_ , \new_[30076]_ , \new_[30077]_ , \new_[30078]_ ,
    \new_[30082]_ , \new_[30083]_ , \new_[30087]_ , \new_[30088]_ ,
    \new_[30089]_ , \new_[30093]_ , \new_[30094]_ , \new_[30098]_ ,
    \new_[30099]_ , \new_[30100]_ , \new_[30104]_ , \new_[30105]_ ,
    \new_[30109]_ , \new_[30110]_ , \new_[30111]_ , \new_[30115]_ ,
    \new_[30116]_ , \new_[30120]_ , \new_[30121]_ , \new_[30122]_ ,
    \new_[30126]_ , \new_[30127]_ , \new_[30131]_ , \new_[30132]_ ,
    \new_[30133]_ , \new_[30137]_ , \new_[30138]_ , \new_[30142]_ ,
    \new_[30143]_ , \new_[30144]_ , \new_[30148]_ , \new_[30149]_ ,
    \new_[30153]_ , \new_[30154]_ , \new_[30155]_ , \new_[30159]_ ,
    \new_[30160]_ , \new_[30164]_ , \new_[30165]_ , \new_[30166]_ ,
    \new_[30170]_ , \new_[30171]_ , \new_[30175]_ , \new_[30176]_ ,
    \new_[30177]_ , \new_[30181]_ , \new_[30182]_ , \new_[30186]_ ,
    \new_[30187]_ , \new_[30188]_ , \new_[30192]_ , \new_[30193]_ ,
    \new_[30197]_ , \new_[30198]_ , \new_[30199]_ , \new_[30203]_ ,
    \new_[30204]_ , \new_[30208]_ , \new_[30209]_ , \new_[30210]_ ,
    \new_[30214]_ , \new_[30215]_ , \new_[30219]_ , \new_[30220]_ ,
    \new_[30221]_ , \new_[30225]_ , \new_[30226]_ , \new_[30230]_ ,
    \new_[30231]_ , \new_[30232]_ , \new_[30236]_ , \new_[30237]_ ,
    \new_[30241]_ , \new_[30242]_ , \new_[30243]_ , \new_[30247]_ ,
    \new_[30248]_ , \new_[30252]_ , \new_[30253]_ , \new_[30254]_ ,
    \new_[30258]_ , \new_[30259]_ , \new_[30263]_ , \new_[30264]_ ,
    \new_[30265]_ , \new_[30269]_ , \new_[30270]_ , \new_[30274]_ ,
    \new_[30275]_ , \new_[30276]_ , \new_[30280]_ , \new_[30281]_ ,
    \new_[30285]_ , \new_[30286]_ , \new_[30287]_ , \new_[30291]_ ,
    \new_[30292]_ , \new_[30296]_ , \new_[30297]_ , \new_[30298]_ ,
    \new_[30302]_ , \new_[30303]_ , \new_[30307]_ , \new_[30308]_ ,
    \new_[30309]_ , \new_[30313]_ , \new_[30314]_ , \new_[30318]_ ,
    \new_[30319]_ , \new_[30320]_ , \new_[30324]_ , \new_[30325]_ ,
    \new_[30329]_ , \new_[30330]_ , \new_[30331]_ , \new_[30335]_ ,
    \new_[30336]_ , \new_[30340]_ , \new_[30341]_ , \new_[30342]_ ,
    \new_[30346]_ , \new_[30347]_ , \new_[30351]_ , \new_[30352]_ ,
    \new_[30353]_ , \new_[30357]_ , \new_[30358]_ , \new_[30362]_ ,
    \new_[30363]_ , \new_[30364]_ , \new_[30368]_ , \new_[30369]_ ,
    \new_[30373]_ , \new_[30374]_ , \new_[30375]_ , \new_[30379]_ ,
    \new_[30380]_ , \new_[30384]_ , \new_[30385]_ , \new_[30386]_ ,
    \new_[30390]_ , \new_[30391]_ , \new_[30395]_ , \new_[30396]_ ,
    \new_[30397]_ , \new_[30401]_ , \new_[30402]_ , \new_[30406]_ ,
    \new_[30407]_ , \new_[30408]_ , \new_[30412]_ , \new_[30413]_ ,
    \new_[30417]_ , \new_[30418]_ , \new_[30419]_ , \new_[30423]_ ,
    \new_[30424]_ , \new_[30428]_ , \new_[30429]_ , \new_[30430]_ ,
    \new_[30434]_ , \new_[30435]_ , \new_[30439]_ , \new_[30440]_ ,
    \new_[30441]_ , \new_[30445]_ , \new_[30446]_ , \new_[30450]_ ,
    \new_[30451]_ , \new_[30452]_ , \new_[30456]_ , \new_[30457]_ ,
    \new_[30461]_ , \new_[30462]_ , \new_[30463]_ , \new_[30467]_ ,
    \new_[30468]_ , \new_[30472]_ , \new_[30473]_ , \new_[30474]_ ,
    \new_[30478]_ , \new_[30479]_ , \new_[30483]_ , \new_[30484]_ ,
    \new_[30485]_ , \new_[30489]_ , \new_[30490]_ , \new_[30494]_ ,
    \new_[30495]_ , \new_[30496]_ , \new_[30500]_ , \new_[30501]_ ,
    \new_[30505]_ , \new_[30506]_ , \new_[30507]_ , \new_[30511]_ ,
    \new_[30512]_ , \new_[30516]_ , \new_[30517]_ , \new_[30518]_ ,
    \new_[30522]_ , \new_[30523]_ , \new_[30527]_ , \new_[30528]_ ,
    \new_[30529]_ , \new_[30533]_ , \new_[30534]_ , \new_[30538]_ ,
    \new_[30539]_ , \new_[30540]_ , \new_[30544]_ , \new_[30545]_ ,
    \new_[30549]_ , \new_[30550]_ , \new_[30551]_ , \new_[30555]_ ,
    \new_[30556]_ , \new_[30560]_ , \new_[30561]_ , \new_[30562]_ ,
    \new_[30566]_ , \new_[30567]_ , \new_[30571]_ , \new_[30572]_ ,
    \new_[30573]_ , \new_[30577]_ , \new_[30578]_ , \new_[30582]_ ,
    \new_[30583]_ , \new_[30584]_ , \new_[30588]_ , \new_[30589]_ ,
    \new_[30593]_ , \new_[30594]_ , \new_[30595]_ , \new_[30599]_ ,
    \new_[30600]_ , \new_[30604]_ , \new_[30605]_ , \new_[30606]_ ,
    \new_[30610]_ , \new_[30611]_ , \new_[30615]_ , \new_[30616]_ ,
    \new_[30617]_ , \new_[30621]_ , \new_[30622]_ , \new_[30626]_ ,
    \new_[30627]_ , \new_[30628]_ , \new_[30632]_ , \new_[30633]_ ,
    \new_[30637]_ , \new_[30638]_ , \new_[30639]_ , \new_[30643]_ ,
    \new_[30644]_ , \new_[30648]_ , \new_[30649]_ , \new_[30650]_ ,
    \new_[30654]_ , \new_[30655]_ , \new_[30659]_ , \new_[30660]_ ,
    \new_[30661]_ , \new_[30665]_ , \new_[30666]_ , \new_[30670]_ ,
    \new_[30671]_ , \new_[30672]_ , \new_[30676]_ , \new_[30677]_ ,
    \new_[30681]_ , \new_[30682]_ , \new_[30683]_ , \new_[30687]_ ,
    \new_[30688]_ , \new_[30692]_ , \new_[30693]_ , \new_[30694]_ ,
    \new_[30698]_ , \new_[30699]_ , \new_[30703]_ , \new_[30704]_ ,
    \new_[30705]_ , \new_[30709]_ , \new_[30710]_ , \new_[30714]_ ,
    \new_[30715]_ , \new_[30716]_ , \new_[30720]_ , \new_[30721]_ ,
    \new_[30725]_ , \new_[30726]_ , \new_[30727]_ , \new_[30731]_ ,
    \new_[30732]_ , \new_[30736]_ , \new_[30737]_ , \new_[30738]_ ,
    \new_[30742]_ , \new_[30743]_ , \new_[30747]_ , \new_[30748]_ ,
    \new_[30749]_ , \new_[30753]_ , \new_[30754]_ , \new_[30758]_ ,
    \new_[30759]_ , \new_[30760]_ , \new_[30764]_ , \new_[30765]_ ,
    \new_[30769]_ , \new_[30770]_ , \new_[30771]_ , \new_[30775]_ ,
    \new_[30776]_ , \new_[30780]_ , \new_[30781]_ , \new_[30782]_ ,
    \new_[30786]_ , \new_[30787]_ , \new_[30791]_ , \new_[30792]_ ,
    \new_[30793]_ , \new_[30797]_ , \new_[30798]_ , \new_[30802]_ ,
    \new_[30803]_ , \new_[30804]_ , \new_[30808]_ , \new_[30809]_ ,
    \new_[30813]_ , \new_[30814]_ , \new_[30815]_ , \new_[30819]_ ,
    \new_[30820]_ , \new_[30824]_ , \new_[30825]_ , \new_[30826]_ ,
    \new_[30830]_ , \new_[30831]_ , \new_[30835]_ , \new_[30836]_ ,
    \new_[30837]_ , \new_[30841]_ , \new_[30842]_ , \new_[30846]_ ,
    \new_[30847]_ , \new_[30848]_ , \new_[30852]_ , \new_[30853]_ ,
    \new_[30857]_ , \new_[30858]_ , \new_[30859]_ , \new_[30863]_ ,
    \new_[30864]_ , \new_[30868]_ , \new_[30869]_ , \new_[30870]_ ,
    \new_[30874]_ , \new_[30875]_ , \new_[30879]_ , \new_[30880]_ ,
    \new_[30881]_ , \new_[30885]_ , \new_[30886]_ , \new_[30890]_ ,
    \new_[30891]_ , \new_[30892]_ , \new_[30896]_ , \new_[30897]_ ,
    \new_[30901]_ , \new_[30902]_ , \new_[30903]_ , \new_[30907]_ ,
    \new_[30908]_ , \new_[30912]_ , \new_[30913]_ , \new_[30914]_ ,
    \new_[30918]_ , \new_[30919]_ , \new_[30923]_ , \new_[30924]_ ,
    \new_[30925]_ , \new_[30929]_ , \new_[30930]_ , \new_[30934]_ ,
    \new_[30935]_ , \new_[30936]_ , \new_[30940]_ , \new_[30941]_ ,
    \new_[30945]_ , \new_[30946]_ , \new_[30947]_ , \new_[30951]_ ,
    \new_[30952]_ , \new_[30956]_ , \new_[30957]_ , \new_[30958]_ ,
    \new_[30962]_ , \new_[30963]_ , \new_[30967]_ , \new_[30968]_ ,
    \new_[30969]_ , \new_[30973]_ , \new_[30974]_ , \new_[30978]_ ,
    \new_[30979]_ , \new_[30980]_ , \new_[30984]_ , \new_[30985]_ ,
    \new_[30989]_ , \new_[30990]_ , \new_[30991]_ , \new_[30995]_ ,
    \new_[30996]_ , \new_[31000]_ , \new_[31001]_ , \new_[31002]_ ,
    \new_[31006]_ , \new_[31007]_ , \new_[31011]_ , \new_[31012]_ ,
    \new_[31013]_ , \new_[31017]_ , \new_[31018]_ , \new_[31022]_ ,
    \new_[31023]_ , \new_[31024]_ , \new_[31028]_ , \new_[31029]_ ,
    \new_[31033]_ , \new_[31034]_ , \new_[31035]_ , \new_[31039]_ ,
    \new_[31040]_ , \new_[31044]_ , \new_[31045]_ , \new_[31046]_ ,
    \new_[31050]_ , \new_[31051]_ , \new_[31055]_ , \new_[31056]_ ,
    \new_[31057]_ , \new_[31061]_ , \new_[31062]_ , \new_[31066]_ ,
    \new_[31067]_ , \new_[31068]_ , \new_[31072]_ , \new_[31073]_ ,
    \new_[31077]_ , \new_[31078]_ , \new_[31079]_ , \new_[31083]_ ,
    \new_[31084]_ , \new_[31088]_ , \new_[31089]_ , \new_[31090]_ ,
    \new_[31094]_ , \new_[31095]_ , \new_[31099]_ , \new_[31100]_ ,
    \new_[31101]_ , \new_[31105]_ , \new_[31106]_ , \new_[31110]_ ,
    \new_[31111]_ , \new_[31112]_ , \new_[31116]_ , \new_[31117]_ ,
    \new_[31121]_ , \new_[31122]_ , \new_[31123]_ , \new_[31127]_ ,
    \new_[31128]_ , \new_[31132]_ , \new_[31133]_ , \new_[31134]_ ,
    \new_[31138]_ , \new_[31139]_ , \new_[31143]_ , \new_[31144]_ ,
    \new_[31145]_ , \new_[31149]_ , \new_[31150]_ , \new_[31154]_ ,
    \new_[31155]_ , \new_[31156]_ , \new_[31160]_ , \new_[31161]_ ,
    \new_[31165]_ , \new_[31166]_ , \new_[31167]_ , \new_[31171]_ ,
    \new_[31172]_ , \new_[31176]_ , \new_[31177]_ , \new_[31178]_ ,
    \new_[31182]_ , \new_[31183]_ , \new_[31187]_ , \new_[31188]_ ,
    \new_[31189]_ , \new_[31193]_ , \new_[31194]_ , \new_[31198]_ ,
    \new_[31199]_ , \new_[31200]_ , \new_[31204]_ , \new_[31205]_ ,
    \new_[31209]_ , \new_[31210]_ , \new_[31211]_ , \new_[31215]_ ,
    \new_[31216]_ , \new_[31220]_ , \new_[31221]_ , \new_[31222]_ ,
    \new_[31226]_ , \new_[31227]_ , \new_[31231]_ , \new_[31232]_ ,
    \new_[31233]_ , \new_[31237]_ , \new_[31238]_ , \new_[31242]_ ,
    \new_[31243]_ , \new_[31244]_ , \new_[31248]_ , \new_[31249]_ ,
    \new_[31253]_ , \new_[31254]_ , \new_[31255]_ , \new_[31259]_ ,
    \new_[31260]_ , \new_[31264]_ , \new_[31265]_ , \new_[31266]_ ,
    \new_[31270]_ , \new_[31271]_ , \new_[31275]_ , \new_[31276]_ ,
    \new_[31277]_ , \new_[31281]_ , \new_[31282]_ , \new_[31286]_ ,
    \new_[31287]_ , \new_[31288]_ , \new_[31292]_ , \new_[31293]_ ,
    \new_[31297]_ , \new_[31298]_ , \new_[31299]_ , \new_[31303]_ ,
    \new_[31304]_ , \new_[31308]_ , \new_[31309]_ , \new_[31310]_ ,
    \new_[31314]_ , \new_[31315]_ , \new_[31319]_ , \new_[31320]_ ,
    \new_[31321]_ , \new_[31325]_ , \new_[31326]_ , \new_[31330]_ ,
    \new_[31331]_ , \new_[31332]_ , \new_[31336]_ , \new_[31337]_ ,
    \new_[31341]_ , \new_[31342]_ , \new_[31343]_ , \new_[31347]_ ,
    \new_[31348]_ , \new_[31352]_ , \new_[31353]_ , \new_[31354]_ ,
    \new_[31358]_ , \new_[31359]_ , \new_[31363]_ , \new_[31364]_ ,
    \new_[31365]_ , \new_[31369]_ , \new_[31370]_ , \new_[31374]_ ,
    \new_[31375]_ , \new_[31376]_ , \new_[31380]_ , \new_[31381]_ ,
    \new_[31385]_ , \new_[31386]_ , \new_[31387]_ , \new_[31391]_ ,
    \new_[31392]_ , \new_[31396]_ , \new_[31397]_ , \new_[31398]_ ,
    \new_[31402]_ , \new_[31403]_ , \new_[31407]_ , \new_[31408]_ ,
    \new_[31409]_ , \new_[31413]_ , \new_[31414]_ , \new_[31418]_ ,
    \new_[31419]_ , \new_[31420]_ , \new_[31424]_ , \new_[31425]_ ,
    \new_[31429]_ , \new_[31430]_ , \new_[31431]_ , \new_[31435]_ ,
    \new_[31436]_ , \new_[31440]_ , \new_[31441]_ , \new_[31442]_ ,
    \new_[31446]_ , \new_[31447]_ , \new_[31451]_ , \new_[31452]_ ,
    \new_[31453]_ , \new_[31457]_ , \new_[31458]_ , \new_[31462]_ ,
    \new_[31463]_ , \new_[31464]_ , \new_[31468]_ , \new_[31469]_ ,
    \new_[31473]_ , \new_[31474]_ , \new_[31475]_ , \new_[31479]_ ,
    \new_[31480]_ , \new_[31484]_ , \new_[31485]_ , \new_[31486]_ ,
    \new_[31490]_ , \new_[31491]_ , \new_[31495]_ , \new_[31496]_ ,
    \new_[31497]_ , \new_[31501]_ , \new_[31502]_ , \new_[31506]_ ,
    \new_[31507]_ , \new_[31508]_ , \new_[31512]_ , \new_[31513]_ ,
    \new_[31517]_ , \new_[31518]_ , \new_[31519]_ , \new_[31523]_ ,
    \new_[31524]_ , \new_[31528]_ , \new_[31529]_ , \new_[31530]_ ,
    \new_[31534]_ , \new_[31535]_ , \new_[31539]_ , \new_[31540]_ ,
    \new_[31541]_ , \new_[31545]_ , \new_[31546]_ , \new_[31550]_ ,
    \new_[31551]_ , \new_[31552]_ , \new_[31556]_ , \new_[31557]_ ,
    \new_[31561]_ , \new_[31562]_ , \new_[31563]_ , \new_[31567]_ ,
    \new_[31568]_ , \new_[31572]_ , \new_[31573]_ , \new_[31574]_ ,
    \new_[31578]_ , \new_[31579]_ , \new_[31583]_ , \new_[31584]_ ,
    \new_[31585]_ , \new_[31589]_ , \new_[31590]_ , \new_[31594]_ ,
    \new_[31595]_ , \new_[31596]_ , \new_[31600]_ , \new_[31601]_ ,
    \new_[31605]_ , \new_[31606]_ , \new_[31607]_ , \new_[31611]_ ,
    \new_[31612]_ , \new_[31616]_ , \new_[31617]_ , \new_[31618]_ ,
    \new_[31622]_ , \new_[31623]_ , \new_[31627]_ , \new_[31628]_ ,
    \new_[31629]_ , \new_[31633]_ , \new_[31634]_ , \new_[31638]_ ,
    \new_[31639]_ , \new_[31640]_ , \new_[31644]_ , \new_[31645]_ ,
    \new_[31649]_ , \new_[31650]_ , \new_[31651]_ , \new_[31655]_ ,
    \new_[31656]_ , \new_[31660]_ , \new_[31661]_ , \new_[31662]_ ,
    \new_[31666]_ , \new_[31667]_ , \new_[31671]_ , \new_[31672]_ ,
    \new_[31673]_ , \new_[31677]_ , \new_[31678]_ , \new_[31682]_ ,
    \new_[31683]_ , \new_[31684]_ , \new_[31688]_ , \new_[31689]_ ,
    \new_[31693]_ , \new_[31694]_ , \new_[31695]_ , \new_[31699]_ ,
    \new_[31700]_ , \new_[31704]_ , \new_[31705]_ , \new_[31706]_ ,
    \new_[31710]_ , \new_[31711]_ , \new_[31715]_ , \new_[31716]_ ,
    \new_[31717]_ , \new_[31721]_ , \new_[31722]_ , \new_[31726]_ ,
    \new_[31727]_ , \new_[31728]_ , \new_[31732]_ , \new_[31733]_ ,
    \new_[31737]_ , \new_[31738]_ , \new_[31739]_ , \new_[31743]_ ,
    \new_[31744]_ , \new_[31748]_ , \new_[31749]_ , \new_[31750]_ ,
    \new_[31754]_ , \new_[31755]_ , \new_[31759]_ , \new_[31760]_ ,
    \new_[31761]_ , \new_[31765]_ , \new_[31766]_ , \new_[31770]_ ,
    \new_[31771]_ , \new_[31772]_ , \new_[31776]_ , \new_[31777]_ ,
    \new_[31781]_ , \new_[31782]_ , \new_[31783]_ , \new_[31787]_ ,
    \new_[31788]_ , \new_[31792]_ , \new_[31793]_ , \new_[31794]_ ,
    \new_[31798]_ , \new_[31799]_ , \new_[31803]_ , \new_[31804]_ ,
    \new_[31805]_ , \new_[31809]_ , \new_[31810]_ , \new_[31814]_ ,
    \new_[31815]_ , \new_[31816]_ , \new_[31820]_ , \new_[31821]_ ,
    \new_[31825]_ , \new_[31826]_ , \new_[31827]_ , \new_[31831]_ ,
    \new_[31832]_ , \new_[31836]_ , \new_[31837]_ , \new_[31838]_ ,
    \new_[31842]_ , \new_[31843]_ , \new_[31847]_ , \new_[31848]_ ,
    \new_[31849]_ , \new_[31853]_ , \new_[31854]_ , \new_[31858]_ ,
    \new_[31859]_ , \new_[31860]_ , \new_[31864]_ , \new_[31865]_ ,
    \new_[31869]_ , \new_[31870]_ , \new_[31871]_ , \new_[31875]_ ,
    \new_[31876]_ , \new_[31880]_ , \new_[31881]_ , \new_[31882]_ ,
    \new_[31886]_ , \new_[31887]_ , \new_[31891]_ , \new_[31892]_ ,
    \new_[31893]_ , \new_[31897]_ , \new_[31898]_ , \new_[31902]_ ,
    \new_[31903]_ , \new_[31904]_ , \new_[31908]_ , \new_[31909]_ ,
    \new_[31913]_ , \new_[31914]_ , \new_[31915]_ , \new_[31919]_ ,
    \new_[31920]_ , \new_[31924]_ , \new_[31925]_ , \new_[31926]_ ,
    \new_[31930]_ , \new_[31931]_ , \new_[31935]_ , \new_[31936]_ ,
    \new_[31937]_ , \new_[31941]_ , \new_[31942]_ , \new_[31946]_ ,
    \new_[31947]_ , \new_[31948]_ , \new_[31952]_ , \new_[31953]_ ,
    \new_[31957]_ , \new_[31958]_ , \new_[31959]_ , \new_[31963]_ ,
    \new_[31964]_ , \new_[31968]_ , \new_[31969]_ , \new_[31970]_ ,
    \new_[31974]_ , \new_[31975]_ , \new_[31979]_ , \new_[31980]_ ,
    \new_[31981]_ , \new_[31985]_ , \new_[31986]_ , \new_[31990]_ ,
    \new_[31991]_ , \new_[31992]_ , \new_[31996]_ , \new_[31997]_ ,
    \new_[32001]_ , \new_[32002]_ , \new_[32003]_ , \new_[32007]_ ,
    \new_[32008]_ , \new_[32012]_ , \new_[32013]_ , \new_[32014]_ ,
    \new_[32018]_ , \new_[32019]_ , \new_[32023]_ , \new_[32024]_ ,
    \new_[32025]_ , \new_[32029]_ , \new_[32030]_ , \new_[32034]_ ,
    \new_[32035]_ , \new_[32036]_ , \new_[32040]_ , \new_[32041]_ ,
    \new_[32045]_ , \new_[32046]_ , \new_[32047]_ , \new_[32051]_ ,
    \new_[32052]_ , \new_[32056]_ , \new_[32057]_ , \new_[32058]_ ,
    \new_[32062]_ , \new_[32063]_ , \new_[32067]_ , \new_[32068]_ ,
    \new_[32069]_ , \new_[32073]_ , \new_[32074]_ , \new_[32078]_ ,
    \new_[32079]_ , \new_[32080]_ , \new_[32084]_ , \new_[32085]_ ,
    \new_[32089]_ , \new_[32090]_ , \new_[32091]_ , \new_[32095]_ ,
    \new_[32096]_ , \new_[32100]_ , \new_[32101]_ , \new_[32102]_ ,
    \new_[32106]_ , \new_[32107]_ , \new_[32111]_ , \new_[32112]_ ,
    \new_[32113]_ , \new_[32117]_ , \new_[32118]_ , \new_[32122]_ ,
    \new_[32123]_ , \new_[32124]_ , \new_[32128]_ , \new_[32129]_ ,
    \new_[32133]_ , \new_[32134]_ , \new_[32135]_ , \new_[32139]_ ,
    \new_[32140]_ , \new_[32144]_ , \new_[32145]_ , \new_[32146]_ ,
    \new_[32150]_ , \new_[32151]_ , \new_[32155]_ , \new_[32156]_ ,
    \new_[32157]_ , \new_[32161]_ , \new_[32162]_ , \new_[32166]_ ,
    \new_[32167]_ , \new_[32168]_ , \new_[32172]_ , \new_[32173]_ ,
    \new_[32177]_ , \new_[32178]_ , \new_[32179]_ , \new_[32183]_ ,
    \new_[32184]_ , \new_[32188]_ , \new_[32189]_ , \new_[32190]_ ,
    \new_[32194]_ , \new_[32195]_ , \new_[32199]_ , \new_[32200]_ ,
    \new_[32201]_ , \new_[32205]_ , \new_[32206]_ , \new_[32210]_ ,
    \new_[32211]_ , \new_[32212]_ , \new_[32216]_ , \new_[32217]_ ,
    \new_[32221]_ , \new_[32222]_ , \new_[32223]_ , \new_[32227]_ ,
    \new_[32228]_ , \new_[32232]_ , \new_[32233]_ , \new_[32234]_ ,
    \new_[32238]_ , \new_[32239]_ , \new_[32243]_ , \new_[32244]_ ,
    \new_[32245]_ , \new_[32249]_ , \new_[32250]_ , \new_[32254]_ ,
    \new_[32255]_ , \new_[32256]_ , \new_[32260]_ , \new_[32261]_ ,
    \new_[32265]_ , \new_[32266]_ , \new_[32267]_ , \new_[32271]_ ,
    \new_[32272]_ , \new_[32276]_ , \new_[32277]_ , \new_[32278]_ ,
    \new_[32282]_ , \new_[32283]_ , \new_[32287]_ , \new_[32288]_ ,
    \new_[32289]_ , \new_[32293]_ , \new_[32294]_ , \new_[32298]_ ,
    \new_[32299]_ , \new_[32300]_ , \new_[32304]_ , \new_[32305]_ ,
    \new_[32309]_ , \new_[32310]_ , \new_[32311]_ , \new_[32315]_ ,
    \new_[32316]_ , \new_[32320]_ , \new_[32321]_ , \new_[32322]_ ,
    \new_[32326]_ , \new_[32327]_ , \new_[32331]_ , \new_[32332]_ ,
    \new_[32333]_ , \new_[32337]_ , \new_[32338]_ , \new_[32342]_ ,
    \new_[32343]_ , \new_[32344]_ , \new_[32348]_ , \new_[32349]_ ,
    \new_[32353]_ , \new_[32354]_ , \new_[32355]_ , \new_[32359]_ ,
    \new_[32360]_ , \new_[32364]_ , \new_[32365]_ , \new_[32366]_ ,
    \new_[32370]_ , \new_[32371]_ , \new_[32375]_ , \new_[32376]_ ,
    \new_[32377]_ , \new_[32381]_ , \new_[32382]_ , \new_[32386]_ ,
    \new_[32387]_ , \new_[32388]_ , \new_[32392]_ , \new_[32393]_ ,
    \new_[32397]_ , \new_[32398]_ , \new_[32399]_ , \new_[32403]_ ,
    \new_[32404]_ , \new_[32408]_ , \new_[32409]_ , \new_[32410]_ ,
    \new_[32414]_ , \new_[32415]_ , \new_[32419]_ , \new_[32420]_ ,
    \new_[32421]_ , \new_[32425]_ , \new_[32426]_ , \new_[32430]_ ,
    \new_[32431]_ , \new_[32432]_ , \new_[32436]_ , \new_[32437]_ ,
    \new_[32441]_ , \new_[32442]_ , \new_[32443]_ , \new_[32447]_ ,
    \new_[32448]_ , \new_[32452]_ , \new_[32453]_ , \new_[32454]_ ,
    \new_[32458]_ , \new_[32459]_ , \new_[32463]_ , \new_[32464]_ ,
    \new_[32465]_ , \new_[32469]_ , \new_[32470]_ , \new_[32474]_ ,
    \new_[32475]_ , \new_[32476]_ , \new_[32480]_ , \new_[32481]_ ,
    \new_[32485]_ , \new_[32486]_ , \new_[32487]_ , \new_[32491]_ ,
    \new_[32492]_ , \new_[32496]_ , \new_[32497]_ , \new_[32498]_ ,
    \new_[32502]_ , \new_[32503]_ , \new_[32507]_ , \new_[32508]_ ,
    \new_[32509]_ , \new_[32513]_ , \new_[32514]_ , \new_[32518]_ ,
    \new_[32519]_ , \new_[32520]_ , \new_[32524]_ , \new_[32525]_ ,
    \new_[32529]_ , \new_[32530]_ , \new_[32531]_ , \new_[32535]_ ,
    \new_[32536]_ , \new_[32540]_ , \new_[32541]_ , \new_[32542]_ ,
    \new_[32546]_ , \new_[32547]_ , \new_[32551]_ , \new_[32552]_ ,
    \new_[32553]_ , \new_[32557]_ , \new_[32558]_ , \new_[32562]_ ,
    \new_[32563]_ , \new_[32564]_ , \new_[32568]_ , \new_[32569]_ ,
    \new_[32573]_ , \new_[32574]_ , \new_[32575]_ , \new_[32579]_ ,
    \new_[32580]_ , \new_[32584]_ , \new_[32585]_ , \new_[32586]_ ,
    \new_[32590]_ , \new_[32591]_ , \new_[32595]_ , \new_[32596]_ ,
    \new_[32597]_ , \new_[32601]_ , \new_[32602]_ , \new_[32606]_ ,
    \new_[32607]_ , \new_[32608]_ , \new_[32612]_ , \new_[32613]_ ,
    \new_[32617]_ , \new_[32618]_ , \new_[32619]_ , \new_[32623]_ ,
    \new_[32624]_ , \new_[32628]_ , \new_[32629]_ , \new_[32630]_ ,
    \new_[32634]_ , \new_[32635]_ , \new_[32639]_ , \new_[32640]_ ,
    \new_[32641]_ , \new_[32645]_ , \new_[32646]_ , \new_[32650]_ ,
    \new_[32651]_ , \new_[32652]_ , \new_[32656]_ , \new_[32657]_ ,
    \new_[32661]_ , \new_[32662]_ , \new_[32663]_ , \new_[32667]_ ,
    \new_[32668]_ , \new_[32672]_ , \new_[32673]_ , \new_[32674]_ ,
    \new_[32678]_ , \new_[32679]_ , \new_[32683]_ , \new_[32684]_ ,
    \new_[32685]_ , \new_[32689]_ , \new_[32690]_ , \new_[32694]_ ,
    \new_[32695]_ , \new_[32696]_ , \new_[32700]_ , \new_[32701]_ ,
    \new_[32705]_ , \new_[32706]_ , \new_[32707]_ , \new_[32711]_ ,
    \new_[32712]_ , \new_[32716]_ , \new_[32717]_ , \new_[32718]_ ,
    \new_[32722]_ , \new_[32723]_ , \new_[32727]_ , \new_[32728]_ ,
    \new_[32729]_ , \new_[32733]_ , \new_[32734]_ , \new_[32738]_ ,
    \new_[32739]_ , \new_[32740]_ , \new_[32744]_ , \new_[32745]_ ,
    \new_[32749]_ , \new_[32750]_ , \new_[32751]_ , \new_[32755]_ ,
    \new_[32756]_ , \new_[32760]_ , \new_[32761]_ , \new_[32762]_ ,
    \new_[32766]_ , \new_[32767]_ , \new_[32771]_ , \new_[32772]_ ,
    \new_[32773]_ , \new_[32777]_ , \new_[32778]_ , \new_[32782]_ ,
    \new_[32783]_ , \new_[32784]_ , \new_[32788]_ , \new_[32789]_ ,
    \new_[32793]_ , \new_[32794]_ , \new_[32795]_ , \new_[32799]_ ,
    \new_[32800]_ , \new_[32804]_ , \new_[32805]_ , \new_[32806]_ ,
    \new_[32810]_ , \new_[32811]_ , \new_[32815]_ , \new_[32816]_ ,
    \new_[32817]_ , \new_[32821]_ , \new_[32822]_ , \new_[32826]_ ,
    \new_[32827]_ , \new_[32828]_ , \new_[32832]_ , \new_[32833]_ ,
    \new_[32837]_ , \new_[32838]_ , \new_[32839]_ , \new_[32843]_ ,
    \new_[32844]_ , \new_[32848]_ , \new_[32849]_ , \new_[32850]_ ,
    \new_[32854]_ , \new_[32855]_ , \new_[32859]_ , \new_[32860]_ ,
    \new_[32861]_ , \new_[32865]_ , \new_[32866]_ , \new_[32870]_ ,
    \new_[32871]_ , \new_[32872]_ , \new_[32876]_ , \new_[32877]_ ,
    \new_[32881]_ , \new_[32882]_ , \new_[32883]_ , \new_[32887]_ ,
    \new_[32888]_ , \new_[32892]_ , \new_[32893]_ , \new_[32894]_ ,
    \new_[32898]_ , \new_[32899]_ , \new_[32903]_ , \new_[32904]_ ,
    \new_[32905]_ , \new_[32909]_ , \new_[32910]_ , \new_[32914]_ ,
    \new_[32915]_ , \new_[32916]_ , \new_[32920]_ , \new_[32921]_ ,
    \new_[32925]_ , \new_[32926]_ , \new_[32927]_ , \new_[32931]_ ,
    \new_[32932]_ , \new_[32936]_ , \new_[32937]_ , \new_[32938]_ ,
    \new_[32942]_ , \new_[32943]_ , \new_[32947]_ , \new_[32948]_ ,
    \new_[32949]_ , \new_[32953]_ , \new_[32954]_ , \new_[32958]_ ,
    \new_[32959]_ , \new_[32960]_ , \new_[32964]_ , \new_[32965]_ ,
    \new_[32969]_ , \new_[32970]_ , \new_[32971]_ , \new_[32975]_ ,
    \new_[32976]_ , \new_[32979]_ , \new_[32982]_ , \new_[32983]_ ,
    \new_[32984]_ , \new_[32988]_ , \new_[32989]_ , \new_[32993]_ ,
    \new_[32994]_ , \new_[32995]_ , \new_[32999]_ , \new_[33000]_ ,
    \new_[33003]_ , \new_[33006]_ , \new_[33007]_ , \new_[33008]_ ,
    \new_[33012]_ , \new_[33013]_ , \new_[33017]_ , \new_[33018]_ ,
    \new_[33019]_ , \new_[33023]_ , \new_[33024]_ , \new_[33027]_ ,
    \new_[33030]_ , \new_[33031]_ , \new_[33032]_ , \new_[33036]_ ,
    \new_[33037]_ , \new_[33041]_ , \new_[33042]_ , \new_[33043]_ ,
    \new_[33047]_ , \new_[33048]_ , \new_[33051]_ , \new_[33054]_ ,
    \new_[33055]_ , \new_[33056]_ , \new_[33060]_ , \new_[33061]_ ,
    \new_[33065]_ , \new_[33066]_ , \new_[33067]_ , \new_[33071]_ ,
    \new_[33072]_ , \new_[33075]_ , \new_[33078]_ , \new_[33079]_ ,
    \new_[33080]_ , \new_[33084]_ , \new_[33085]_ , \new_[33089]_ ,
    \new_[33090]_ , \new_[33091]_ , \new_[33095]_ , \new_[33096]_ ,
    \new_[33099]_ , \new_[33102]_ , \new_[33103]_ , \new_[33104]_ ,
    \new_[33108]_ , \new_[33109]_ , \new_[33113]_ , \new_[33114]_ ,
    \new_[33115]_ , \new_[33119]_ , \new_[33120]_ , \new_[33123]_ ,
    \new_[33126]_ , \new_[33127]_ , \new_[33128]_ , \new_[33132]_ ,
    \new_[33133]_ , \new_[33137]_ , \new_[33138]_ , \new_[33139]_ ,
    \new_[33143]_ , \new_[33144]_ , \new_[33147]_ , \new_[33150]_ ,
    \new_[33151]_ , \new_[33152]_ , \new_[33156]_ , \new_[33157]_ ,
    \new_[33161]_ , \new_[33162]_ , \new_[33163]_ , \new_[33167]_ ,
    \new_[33168]_ , \new_[33171]_ , \new_[33174]_ , \new_[33175]_ ,
    \new_[33176]_ , \new_[33180]_ , \new_[33181]_ , \new_[33185]_ ,
    \new_[33186]_ , \new_[33187]_ , \new_[33191]_ , \new_[33192]_ ,
    \new_[33195]_ , \new_[33198]_ , \new_[33199]_ , \new_[33200]_ ,
    \new_[33204]_ , \new_[33205]_ , \new_[33209]_ , \new_[33210]_ ,
    \new_[33211]_ , \new_[33215]_ , \new_[33216]_ , \new_[33219]_ ,
    \new_[33222]_ , \new_[33223]_ , \new_[33224]_ , \new_[33228]_ ,
    \new_[33229]_ , \new_[33233]_ , \new_[33234]_ , \new_[33235]_ ,
    \new_[33239]_ , \new_[33240]_ , \new_[33243]_ , \new_[33246]_ ,
    \new_[33247]_ , \new_[33248]_ , \new_[33252]_ , \new_[33253]_ ,
    \new_[33257]_ , \new_[33258]_ , \new_[33259]_ , \new_[33263]_ ,
    \new_[33264]_ , \new_[33267]_ , \new_[33270]_ , \new_[33271]_ ,
    \new_[33272]_ , \new_[33276]_ , \new_[33277]_ , \new_[33281]_ ,
    \new_[33282]_ , \new_[33283]_ , \new_[33287]_ , \new_[33288]_ ,
    \new_[33291]_ , \new_[33294]_ , \new_[33295]_ , \new_[33296]_ ,
    \new_[33300]_ , \new_[33301]_ , \new_[33305]_ , \new_[33306]_ ,
    \new_[33307]_ , \new_[33311]_ , \new_[33312]_ , \new_[33315]_ ,
    \new_[33318]_ , \new_[33319]_ , \new_[33320]_ , \new_[33324]_ ,
    \new_[33325]_ , \new_[33329]_ , \new_[33330]_ , \new_[33331]_ ,
    \new_[33335]_ , \new_[33336]_ , \new_[33339]_ , \new_[33342]_ ,
    \new_[33343]_ , \new_[33344]_ , \new_[33348]_ , \new_[33349]_ ,
    \new_[33353]_ , \new_[33354]_ , \new_[33355]_ , \new_[33359]_ ,
    \new_[33360]_ , \new_[33363]_ , \new_[33366]_ , \new_[33367]_ ,
    \new_[33368]_ , \new_[33372]_ , \new_[33373]_ , \new_[33377]_ ,
    \new_[33378]_ , \new_[33379]_ , \new_[33383]_ , \new_[33384]_ ,
    \new_[33387]_ , \new_[33390]_ , \new_[33391]_ , \new_[33392]_ ,
    \new_[33396]_ , \new_[33397]_ , \new_[33401]_ , \new_[33402]_ ,
    \new_[33403]_ , \new_[33407]_ , \new_[33408]_ , \new_[33411]_ ,
    \new_[33414]_ , \new_[33415]_ , \new_[33416]_ , \new_[33420]_ ,
    \new_[33421]_ , \new_[33425]_ , \new_[33426]_ , \new_[33427]_ ,
    \new_[33431]_ , \new_[33432]_ , \new_[33435]_ , \new_[33438]_ ,
    \new_[33439]_ , \new_[33440]_ , \new_[33444]_ , \new_[33445]_ ,
    \new_[33449]_ , \new_[33450]_ , \new_[33451]_ , \new_[33455]_ ,
    \new_[33456]_ , \new_[33459]_ , \new_[33462]_ , \new_[33463]_ ,
    \new_[33464]_ , \new_[33468]_ , \new_[33469]_ , \new_[33473]_ ,
    \new_[33474]_ , \new_[33475]_ , \new_[33479]_ , \new_[33480]_ ,
    \new_[33483]_ , \new_[33486]_ , \new_[33487]_ , \new_[33488]_ ,
    \new_[33492]_ , \new_[33493]_ , \new_[33497]_ , \new_[33498]_ ,
    \new_[33499]_ , \new_[33503]_ , \new_[33504]_ , \new_[33507]_ ,
    \new_[33510]_ , \new_[33511]_ , \new_[33512]_ , \new_[33516]_ ,
    \new_[33517]_ , \new_[33521]_ , \new_[33522]_ , \new_[33523]_ ,
    \new_[33527]_ , \new_[33528]_ , \new_[33531]_ , \new_[33534]_ ,
    \new_[33535]_ , \new_[33536]_ , \new_[33540]_ , \new_[33541]_ ,
    \new_[33545]_ , \new_[33546]_ , \new_[33547]_ , \new_[33551]_ ,
    \new_[33552]_ , \new_[33555]_ , \new_[33558]_ , \new_[33559]_ ,
    \new_[33560]_ , \new_[33564]_ , \new_[33565]_ , \new_[33569]_ ,
    \new_[33570]_ , \new_[33571]_ , \new_[33575]_ , \new_[33576]_ ,
    \new_[33579]_ , \new_[33582]_ , \new_[33583]_ , \new_[33584]_ ,
    \new_[33588]_ , \new_[33589]_ , \new_[33593]_ , \new_[33594]_ ,
    \new_[33595]_ , \new_[33599]_ , \new_[33600]_ , \new_[33603]_ ,
    \new_[33606]_ , \new_[33607]_ , \new_[33608]_ , \new_[33612]_ ,
    \new_[33613]_ , \new_[33617]_ , \new_[33618]_ , \new_[33619]_ ,
    \new_[33623]_ , \new_[33624]_ , \new_[33627]_ , \new_[33630]_ ,
    \new_[33631]_ , \new_[33632]_ , \new_[33636]_ , \new_[33637]_ ,
    \new_[33641]_ , \new_[33642]_ , \new_[33643]_ , \new_[33647]_ ,
    \new_[33648]_ , \new_[33651]_ , \new_[33654]_ , \new_[33655]_ ,
    \new_[33656]_ , \new_[33660]_ , \new_[33661]_ , \new_[33665]_ ,
    \new_[33666]_ , \new_[33667]_ , \new_[33671]_ , \new_[33672]_ ,
    \new_[33675]_ , \new_[33678]_ , \new_[33679]_ , \new_[33680]_ ,
    \new_[33684]_ , \new_[33685]_ , \new_[33689]_ , \new_[33690]_ ,
    \new_[33691]_ , \new_[33695]_ , \new_[33696]_ , \new_[33699]_ ,
    \new_[33702]_ , \new_[33703]_ , \new_[33704]_ , \new_[33708]_ ,
    \new_[33709]_ , \new_[33713]_ , \new_[33714]_ , \new_[33715]_ ,
    \new_[33719]_ , \new_[33720]_ , \new_[33723]_ , \new_[33726]_ ,
    \new_[33727]_ , \new_[33728]_ , \new_[33732]_ , \new_[33733]_ ,
    \new_[33737]_ , \new_[33738]_ , \new_[33739]_ , \new_[33743]_ ,
    \new_[33744]_ , \new_[33747]_ , \new_[33750]_ , \new_[33751]_ ,
    \new_[33752]_ , \new_[33756]_ , \new_[33757]_ , \new_[33761]_ ,
    \new_[33762]_ , \new_[33763]_ , \new_[33767]_ , \new_[33768]_ ,
    \new_[33771]_ , \new_[33774]_ , \new_[33775]_ , \new_[33776]_ ,
    \new_[33780]_ , \new_[33781]_ , \new_[33785]_ , \new_[33786]_ ,
    \new_[33787]_ , \new_[33791]_ , \new_[33792]_ , \new_[33795]_ ,
    \new_[33798]_ , \new_[33799]_ , \new_[33800]_ , \new_[33804]_ ,
    \new_[33805]_ , \new_[33809]_ , \new_[33810]_ , \new_[33811]_ ,
    \new_[33815]_ , \new_[33816]_ , \new_[33819]_ , \new_[33822]_ ,
    \new_[33823]_ , \new_[33824]_ , \new_[33828]_ , \new_[33829]_ ,
    \new_[33833]_ , \new_[33834]_ , \new_[33835]_ , \new_[33839]_ ,
    \new_[33840]_ , \new_[33843]_ , \new_[33846]_ , \new_[33847]_ ,
    \new_[33848]_ , \new_[33852]_ , \new_[33853]_ , \new_[33857]_ ,
    \new_[33858]_ , \new_[33859]_ , \new_[33863]_ , \new_[33864]_ ,
    \new_[33867]_ , \new_[33870]_ , \new_[33871]_ , \new_[33872]_ ,
    \new_[33876]_ , \new_[33877]_ , \new_[33881]_ , \new_[33882]_ ,
    \new_[33883]_ , \new_[33887]_ , \new_[33888]_ , \new_[33891]_ ,
    \new_[33894]_ , \new_[33895]_ , \new_[33896]_ , \new_[33900]_ ,
    \new_[33901]_ , \new_[33905]_ , \new_[33906]_ , \new_[33907]_ ,
    \new_[33911]_ , \new_[33912]_ , \new_[33915]_ , \new_[33918]_ ,
    \new_[33919]_ , \new_[33920]_ , \new_[33924]_ , \new_[33925]_ ,
    \new_[33929]_ , \new_[33930]_ , \new_[33931]_ , \new_[33935]_ ,
    \new_[33936]_ , \new_[33939]_ , \new_[33942]_ , \new_[33943]_ ,
    \new_[33944]_ , \new_[33948]_ , \new_[33949]_ , \new_[33953]_ ,
    \new_[33954]_ , \new_[33955]_ , \new_[33959]_ , \new_[33960]_ ,
    \new_[33963]_ , \new_[33966]_ , \new_[33967]_ , \new_[33968]_ ,
    \new_[33972]_ , \new_[33973]_ , \new_[33977]_ , \new_[33978]_ ,
    \new_[33979]_ , \new_[33983]_ , \new_[33984]_ , \new_[33987]_ ,
    \new_[33990]_ , \new_[33991]_ , \new_[33992]_ , \new_[33996]_ ,
    \new_[33997]_ , \new_[34001]_ , \new_[34002]_ , \new_[34003]_ ,
    \new_[34007]_ , \new_[34008]_ , \new_[34011]_ , \new_[34014]_ ,
    \new_[34015]_ , \new_[34016]_ , \new_[34020]_ , \new_[34021]_ ,
    \new_[34025]_ , \new_[34026]_ , \new_[34027]_ , \new_[34031]_ ,
    \new_[34032]_ , \new_[34035]_ , \new_[34038]_ , \new_[34039]_ ,
    \new_[34040]_ , \new_[34044]_ , \new_[34045]_ , \new_[34049]_ ,
    \new_[34050]_ , \new_[34051]_ , \new_[34055]_ , \new_[34056]_ ,
    \new_[34059]_ , \new_[34062]_ , \new_[34063]_ , \new_[34064]_ ,
    \new_[34068]_ , \new_[34069]_ , \new_[34073]_ , \new_[34074]_ ,
    \new_[34075]_ , \new_[34079]_ , \new_[34080]_ , \new_[34083]_ ,
    \new_[34086]_ , \new_[34087]_ , \new_[34088]_ , \new_[34092]_ ,
    \new_[34093]_ , \new_[34097]_ , \new_[34098]_ , \new_[34099]_ ,
    \new_[34103]_ , \new_[34104]_ , \new_[34107]_ , \new_[34110]_ ,
    \new_[34111]_ , \new_[34112]_ , \new_[34116]_ , \new_[34117]_ ,
    \new_[34121]_ , \new_[34122]_ , \new_[34123]_ , \new_[34127]_ ,
    \new_[34128]_ , \new_[34131]_ , \new_[34134]_ , \new_[34135]_ ,
    \new_[34136]_ , \new_[34140]_ , \new_[34141]_ , \new_[34145]_ ,
    \new_[34146]_ , \new_[34147]_ , \new_[34151]_ , \new_[34152]_ ,
    \new_[34155]_ , \new_[34158]_ , \new_[34159]_ , \new_[34160]_ ,
    \new_[34164]_ , \new_[34165]_ , \new_[34169]_ , \new_[34170]_ ,
    \new_[34171]_ , \new_[34175]_ , \new_[34176]_ , \new_[34179]_ ,
    \new_[34182]_ , \new_[34183]_ , \new_[34184]_ , \new_[34188]_ ,
    \new_[34189]_ , \new_[34193]_ , \new_[34194]_ , \new_[34195]_ ,
    \new_[34199]_ , \new_[34200]_ , \new_[34203]_ , \new_[34206]_ ,
    \new_[34207]_ , \new_[34208]_ , \new_[34212]_ , \new_[34213]_ ,
    \new_[34217]_ , \new_[34218]_ , \new_[34219]_ , \new_[34223]_ ,
    \new_[34224]_ , \new_[34227]_ , \new_[34230]_ , \new_[34231]_ ,
    \new_[34232]_ , \new_[34236]_ , \new_[34237]_ , \new_[34241]_ ,
    \new_[34242]_ , \new_[34243]_ , \new_[34247]_ , \new_[34248]_ ,
    \new_[34251]_ , \new_[34254]_ , \new_[34255]_ , \new_[34256]_ ,
    \new_[34260]_ , \new_[34261]_ , \new_[34265]_ , \new_[34266]_ ,
    \new_[34267]_ , \new_[34271]_ , \new_[34272]_ , \new_[34275]_ ,
    \new_[34278]_ , \new_[34279]_ , \new_[34280]_ , \new_[34284]_ ,
    \new_[34285]_ , \new_[34289]_ , \new_[34290]_ , \new_[34291]_ ,
    \new_[34295]_ , \new_[34296]_ , \new_[34299]_ , \new_[34302]_ ,
    \new_[34303]_ , \new_[34304]_ , \new_[34308]_ , \new_[34309]_ ,
    \new_[34313]_ , \new_[34314]_ , \new_[34315]_ , \new_[34319]_ ,
    \new_[34320]_ , \new_[34323]_ , \new_[34326]_ , \new_[34327]_ ,
    \new_[34328]_ , \new_[34332]_ , \new_[34333]_ , \new_[34337]_ ,
    \new_[34338]_ , \new_[34339]_ , \new_[34343]_ , \new_[34344]_ ,
    \new_[34347]_ , \new_[34350]_ , \new_[34351]_ , \new_[34352]_ ,
    \new_[34356]_ , \new_[34357]_ , \new_[34361]_ , \new_[34362]_ ,
    \new_[34363]_ , \new_[34367]_ , \new_[34368]_ , \new_[34371]_ ,
    \new_[34374]_ , \new_[34375]_ , \new_[34376]_ , \new_[34380]_ ,
    \new_[34381]_ , \new_[34385]_ , \new_[34386]_ , \new_[34387]_ ,
    \new_[34391]_ , \new_[34392]_ , \new_[34395]_ , \new_[34398]_ ,
    \new_[34399]_ , \new_[34400]_ , \new_[34404]_ , \new_[34405]_ ,
    \new_[34409]_ , \new_[34410]_ , \new_[34411]_ , \new_[34415]_ ,
    \new_[34416]_ , \new_[34419]_ , \new_[34422]_ , \new_[34423]_ ,
    \new_[34424]_ , \new_[34428]_ , \new_[34429]_ , \new_[34433]_ ,
    \new_[34434]_ , \new_[34435]_ , \new_[34439]_ , \new_[34440]_ ,
    \new_[34443]_ , \new_[34446]_ , \new_[34447]_ , \new_[34448]_ ,
    \new_[34452]_ , \new_[34453]_ , \new_[34457]_ , \new_[34458]_ ,
    \new_[34459]_ , \new_[34463]_ , \new_[34464]_ , \new_[34467]_ ,
    \new_[34470]_ , \new_[34471]_ , \new_[34472]_ , \new_[34476]_ ,
    \new_[34477]_ , \new_[34481]_ , \new_[34482]_ , \new_[34483]_ ,
    \new_[34487]_ , \new_[34488]_ , \new_[34491]_ , \new_[34494]_ ,
    \new_[34495]_ , \new_[34496]_ , \new_[34500]_ , \new_[34501]_ ,
    \new_[34504]_ , \new_[34507]_ , \new_[34508]_ , \new_[34509]_ ,
    \new_[34513]_ , \new_[34514]_ , \new_[34517]_ , \new_[34520]_ ,
    \new_[34521]_ , \new_[34522]_ , \new_[34526]_ , \new_[34527]_ ,
    \new_[34530]_ , \new_[34533]_ , \new_[34534]_ , \new_[34535]_ ,
    \new_[34539]_ , \new_[34540]_ , \new_[34543]_ , \new_[34546]_ ,
    \new_[34547]_ , \new_[34548]_ , \new_[34552]_ , \new_[34553]_ ,
    \new_[34556]_ , \new_[34559]_ , \new_[34560]_ , \new_[34561]_ ,
    \new_[34565]_ , \new_[34566]_ , \new_[34569]_ , \new_[34572]_ ,
    \new_[34573]_ , \new_[34574]_ , \new_[34578]_ , \new_[34579]_ ,
    \new_[34582]_ , \new_[34585]_ , \new_[34586]_ , \new_[34587]_ ,
    \new_[34591]_ , \new_[34592]_ , \new_[34595]_ , \new_[34598]_ ,
    \new_[34599]_ , \new_[34600]_ , \new_[34604]_ , \new_[34605]_ ,
    \new_[34608]_ , \new_[34611]_ , \new_[34612]_ , \new_[34613]_ ,
    \new_[34617]_ , \new_[34618]_ , \new_[34621]_ , \new_[34624]_ ,
    \new_[34625]_ , \new_[34626]_ , \new_[34630]_ , \new_[34631]_ ,
    \new_[34634]_ , \new_[34637]_ , \new_[34638]_ , \new_[34639]_ ,
    \new_[34643]_ , \new_[34644]_ , \new_[34647]_ , \new_[34650]_ ,
    \new_[34651]_ , \new_[34652]_ , \new_[34656]_ , \new_[34657]_ ,
    \new_[34660]_ , \new_[34663]_ , \new_[34664]_ , \new_[34665]_ ,
    \new_[34669]_ , \new_[34670]_ , \new_[34673]_ , \new_[34676]_ ,
    \new_[34677]_ , \new_[34678]_ , \new_[34682]_ , \new_[34683]_ ,
    \new_[34686]_ , \new_[34689]_ , \new_[34690]_ , \new_[34691]_ ,
    \new_[34695]_ , \new_[34696]_ , \new_[34699]_ , \new_[34702]_ ,
    \new_[34703]_ , \new_[34704]_ , \new_[34708]_ , \new_[34709]_ ,
    \new_[34712]_ , \new_[34715]_ , \new_[34716]_ , \new_[34717]_ ,
    \new_[34721]_ , \new_[34722]_ , \new_[34725]_ , \new_[34728]_ ,
    \new_[34729]_ , \new_[34730]_ , \new_[34734]_ , \new_[34735]_ ,
    \new_[34738]_ , \new_[34741]_ , \new_[34742]_ , \new_[34743]_ ,
    \new_[34747]_ , \new_[34748]_ , \new_[34751]_ , \new_[34754]_ ,
    \new_[34755]_ , \new_[34756]_ , \new_[34760]_ , \new_[34761]_ ,
    \new_[34764]_ , \new_[34767]_ , \new_[34768]_ , \new_[34769]_ ,
    \new_[34773]_ , \new_[34774]_ , \new_[34777]_ , \new_[34780]_ ,
    \new_[34781]_ , \new_[34782]_ , \new_[34786]_ , \new_[34787]_ ,
    \new_[34790]_ , \new_[34793]_ , \new_[34794]_ , \new_[34795]_ ,
    \new_[34799]_ , \new_[34800]_ , \new_[34803]_ , \new_[34806]_ ,
    \new_[34807]_ , \new_[34808]_ , \new_[34812]_ , \new_[34813]_ ,
    \new_[34816]_ , \new_[34819]_ , \new_[34820]_ , \new_[34821]_ ,
    \new_[34825]_ , \new_[34826]_ , \new_[34829]_ , \new_[34832]_ ,
    \new_[34833]_ , \new_[34834]_ , \new_[34838]_ , \new_[34839]_ ,
    \new_[34842]_ , \new_[34845]_ , \new_[34846]_ , \new_[34847]_ ,
    \new_[34851]_ , \new_[34852]_ , \new_[34855]_ , \new_[34858]_ ,
    \new_[34859]_ , \new_[34860]_ , \new_[34864]_ , \new_[34865]_ ,
    \new_[34868]_ , \new_[34871]_ , \new_[34872]_ , \new_[34873]_ ,
    \new_[34877]_ , \new_[34878]_ , \new_[34881]_ , \new_[34884]_ ,
    \new_[34885]_ , \new_[34886]_ , \new_[34890]_ , \new_[34891]_ ,
    \new_[34894]_ , \new_[34897]_ , \new_[34898]_ , \new_[34899]_ ,
    \new_[34903]_ , \new_[34904]_ , \new_[34907]_ , \new_[34910]_ ,
    \new_[34911]_ , \new_[34912]_ , \new_[34916]_ , \new_[34917]_ ,
    \new_[34920]_ , \new_[34923]_ , \new_[34924]_ , \new_[34925]_ ,
    \new_[34929]_ , \new_[34930]_ , \new_[34933]_ , \new_[34936]_ ,
    \new_[34937]_ , \new_[34938]_ , \new_[34942]_ , \new_[34943]_ ,
    \new_[34946]_ , \new_[34949]_ , \new_[34950]_ , \new_[34951]_ ,
    \new_[34955]_ , \new_[34956]_ , \new_[34959]_ , \new_[34962]_ ,
    \new_[34963]_ , \new_[34964]_ , \new_[34968]_ , \new_[34969]_ ,
    \new_[34972]_ , \new_[34975]_ , \new_[34976]_ , \new_[34977]_ ,
    \new_[34981]_ , \new_[34982]_ , \new_[34985]_ , \new_[34988]_ ,
    \new_[34989]_ , \new_[34990]_ , \new_[34994]_ , \new_[34995]_ ,
    \new_[34998]_ , \new_[35001]_ , \new_[35002]_ , \new_[35003]_ ,
    \new_[35007]_ , \new_[35008]_ , \new_[35011]_ , \new_[35014]_ ,
    \new_[35015]_ , \new_[35016]_ , \new_[35020]_ , \new_[35021]_ ,
    \new_[35024]_ , \new_[35027]_ , \new_[35028]_ , \new_[35029]_ ,
    \new_[35033]_ , \new_[35034]_ , \new_[35037]_ , \new_[35040]_ ,
    \new_[35041]_ , \new_[35042]_ , \new_[35046]_ , \new_[35047]_ ,
    \new_[35050]_ , \new_[35053]_ , \new_[35054]_ , \new_[35055]_ ,
    \new_[35059]_ , \new_[35060]_ , \new_[35063]_ , \new_[35066]_ ,
    \new_[35067]_ , \new_[35068]_ , \new_[35072]_ , \new_[35073]_ ,
    \new_[35076]_ , \new_[35079]_ , \new_[35080]_ , \new_[35081]_ ,
    \new_[35085]_ , \new_[35086]_ , \new_[35089]_ , \new_[35092]_ ,
    \new_[35093]_ , \new_[35094]_ , \new_[35098]_ , \new_[35099]_ ,
    \new_[35102]_ , \new_[35105]_ , \new_[35106]_ , \new_[35107]_ ,
    \new_[35111]_ , \new_[35112]_ , \new_[35115]_ , \new_[35118]_ ,
    \new_[35119]_ , \new_[35120]_ , \new_[35124]_ , \new_[35125]_ ,
    \new_[35128]_ , \new_[35131]_ , \new_[35132]_ , \new_[35133]_ ,
    \new_[35137]_ , \new_[35138]_ , \new_[35141]_ , \new_[35144]_ ,
    \new_[35145]_ , \new_[35146]_ , \new_[35150]_ , \new_[35151]_ ,
    \new_[35154]_ , \new_[35157]_ , \new_[35158]_ , \new_[35159]_ ,
    \new_[35163]_ , \new_[35164]_ , \new_[35167]_ , \new_[35170]_ ,
    \new_[35171]_ , \new_[35172]_ , \new_[35176]_ , \new_[35177]_ ,
    \new_[35180]_ , \new_[35183]_ , \new_[35184]_ , \new_[35185]_ ,
    \new_[35189]_ , \new_[35190]_ , \new_[35193]_ , \new_[35196]_ ,
    \new_[35197]_ , \new_[35198]_ , \new_[35202]_ , \new_[35203]_ ,
    \new_[35206]_ , \new_[35209]_ , \new_[35210]_ , \new_[35211]_ ,
    \new_[35215]_ , \new_[35216]_ , \new_[35219]_ , \new_[35222]_ ,
    \new_[35223]_ , \new_[35224]_ , \new_[35228]_ , \new_[35229]_ ,
    \new_[35232]_ , \new_[35235]_ , \new_[35236]_ , \new_[35237]_ ,
    \new_[35241]_ , \new_[35242]_ , \new_[35245]_ , \new_[35248]_ ,
    \new_[35249]_ , \new_[35250]_ , \new_[35254]_ , \new_[35255]_ ,
    \new_[35258]_ , \new_[35261]_ , \new_[35262]_ , \new_[35263]_ ,
    \new_[35267]_ , \new_[35268]_ , \new_[35271]_ , \new_[35274]_ ,
    \new_[35275]_ , \new_[35276]_ , \new_[35280]_ , \new_[35281]_ ,
    \new_[35284]_ , \new_[35287]_ , \new_[35288]_ , \new_[35289]_ ,
    \new_[35293]_ , \new_[35294]_ , \new_[35297]_ , \new_[35300]_ ,
    \new_[35301]_ , \new_[35302]_ , \new_[35306]_ , \new_[35307]_ ,
    \new_[35310]_ , \new_[35313]_ , \new_[35314]_ , \new_[35315]_ ,
    \new_[35319]_ , \new_[35320]_ , \new_[35323]_ , \new_[35326]_ ,
    \new_[35327]_ , \new_[35328]_ , \new_[35332]_ , \new_[35333]_ ,
    \new_[35336]_ , \new_[35339]_ , \new_[35340]_ , \new_[35341]_ ,
    \new_[35345]_ , \new_[35346]_ , \new_[35349]_ , \new_[35352]_ ,
    \new_[35353]_ , \new_[35354]_ , \new_[35358]_ , \new_[35359]_ ,
    \new_[35362]_ , \new_[35365]_ , \new_[35366]_ , \new_[35367]_ ,
    \new_[35371]_ , \new_[35372]_ , \new_[35375]_ , \new_[35378]_ ,
    \new_[35379]_ , \new_[35380]_ , \new_[35384]_ , \new_[35385]_ ,
    \new_[35388]_ , \new_[35391]_ , \new_[35392]_ , \new_[35393]_ ,
    \new_[35397]_ , \new_[35398]_ , \new_[35401]_ , \new_[35404]_ ,
    \new_[35405]_ , \new_[35406]_ , \new_[35410]_ , \new_[35411]_ ,
    \new_[35414]_ , \new_[35417]_ , \new_[35418]_ , \new_[35419]_ ,
    \new_[35423]_ , \new_[35424]_ , \new_[35427]_ , \new_[35430]_ ,
    \new_[35431]_ , \new_[35432]_ , \new_[35436]_ , \new_[35437]_ ,
    \new_[35440]_ , \new_[35443]_ , \new_[35444]_ , \new_[35445]_ ,
    \new_[35449]_ , \new_[35450]_ , \new_[35453]_ , \new_[35456]_ ,
    \new_[35457]_ , \new_[35458]_ , \new_[35462]_ , \new_[35463]_ ,
    \new_[35466]_ , \new_[35469]_ , \new_[35470]_ , \new_[35471]_ ,
    \new_[35475]_ , \new_[35476]_ , \new_[35479]_ , \new_[35482]_ ,
    \new_[35483]_ , \new_[35484]_ , \new_[35488]_ , \new_[35489]_ ,
    \new_[35492]_ , \new_[35495]_ , \new_[35496]_ , \new_[35497]_ ,
    \new_[35501]_ , \new_[35502]_ , \new_[35505]_ , \new_[35508]_ ,
    \new_[35509]_ , \new_[35510]_ , \new_[35514]_ , \new_[35515]_ ,
    \new_[35518]_ , \new_[35521]_ , \new_[35522]_ , \new_[35523]_ ,
    \new_[35527]_ , \new_[35528]_ , \new_[35531]_ , \new_[35534]_ ,
    \new_[35535]_ , \new_[35536]_ , \new_[35540]_ , \new_[35541]_ ,
    \new_[35544]_ , \new_[35547]_ , \new_[35548]_ , \new_[35549]_ ,
    \new_[35553]_ , \new_[35554]_ , \new_[35557]_ , \new_[35560]_ ,
    \new_[35561]_ , \new_[35562]_ , \new_[35566]_ , \new_[35567]_ ,
    \new_[35570]_ , \new_[35573]_ , \new_[35574]_ , \new_[35575]_ ,
    \new_[35579]_ , \new_[35580]_ , \new_[35583]_ , \new_[35586]_ ,
    \new_[35587]_ , \new_[35588]_ , \new_[35592]_ , \new_[35593]_ ,
    \new_[35596]_ , \new_[35599]_ , \new_[35600]_ , \new_[35601]_ ,
    \new_[35605]_ , \new_[35606]_ , \new_[35609]_ , \new_[35612]_ ,
    \new_[35613]_ , \new_[35614]_ , \new_[35618]_ , \new_[35619]_ ,
    \new_[35622]_ , \new_[35625]_ , \new_[35626]_ , \new_[35627]_ ,
    \new_[35631]_ , \new_[35632]_ , \new_[35635]_ , \new_[35638]_ ,
    \new_[35639]_ , \new_[35640]_ , \new_[35644]_ , \new_[35645]_ ,
    \new_[35648]_ , \new_[35651]_ , \new_[35652]_ , \new_[35653]_ ,
    \new_[35657]_ , \new_[35658]_ , \new_[35661]_ , \new_[35664]_ ,
    \new_[35665]_ , \new_[35666]_ , \new_[35670]_ , \new_[35671]_ ,
    \new_[35674]_ , \new_[35677]_ , \new_[35678]_ , \new_[35679]_ ,
    \new_[35683]_ , \new_[35684]_ , \new_[35687]_ , \new_[35690]_ ,
    \new_[35691]_ , \new_[35692]_ , \new_[35696]_ , \new_[35697]_ ,
    \new_[35700]_ , \new_[35703]_ , \new_[35704]_ , \new_[35705]_ ,
    \new_[35709]_ , \new_[35710]_ , \new_[35713]_ , \new_[35716]_ ,
    \new_[35717]_ , \new_[35718]_ , \new_[35722]_ , \new_[35723]_ ,
    \new_[35726]_ , \new_[35729]_ , \new_[35730]_ , \new_[35731]_ ,
    \new_[35735]_ , \new_[35736]_ , \new_[35739]_ , \new_[35742]_ ,
    \new_[35743]_ , \new_[35744]_ , \new_[35748]_ , \new_[35749]_ ,
    \new_[35752]_ , \new_[35755]_ , \new_[35756]_ , \new_[35757]_ ,
    \new_[35761]_ , \new_[35762]_ , \new_[35765]_ , \new_[35768]_ ,
    \new_[35769]_ , \new_[35770]_ , \new_[35774]_ , \new_[35775]_ ,
    \new_[35778]_ , \new_[35781]_ , \new_[35782]_ , \new_[35783]_ ,
    \new_[35787]_ , \new_[35788]_ , \new_[35791]_ , \new_[35794]_ ,
    \new_[35795]_ , \new_[35796]_ , \new_[35800]_ , \new_[35801]_ ,
    \new_[35804]_ , \new_[35807]_ , \new_[35808]_ , \new_[35809]_ ,
    \new_[35813]_ , \new_[35814]_ , \new_[35817]_ , \new_[35820]_ ,
    \new_[35821]_ , \new_[35822]_ , \new_[35826]_ , \new_[35827]_ ,
    \new_[35830]_ , \new_[35833]_ , \new_[35834]_ , \new_[35835]_ ,
    \new_[35839]_ , \new_[35840]_ , \new_[35843]_ , \new_[35846]_ ,
    \new_[35847]_ , \new_[35848]_ , \new_[35852]_ , \new_[35853]_ ,
    \new_[35856]_ , \new_[35859]_ , \new_[35860]_ , \new_[35861]_ ,
    \new_[35865]_ , \new_[35866]_ , \new_[35869]_ , \new_[35872]_ ,
    \new_[35873]_ , \new_[35874]_ , \new_[35878]_ , \new_[35879]_ ,
    \new_[35882]_ , \new_[35885]_ , \new_[35886]_ , \new_[35887]_ ,
    \new_[35891]_ , \new_[35892]_ , \new_[35895]_ , \new_[35898]_ ,
    \new_[35899]_ , \new_[35900]_ , \new_[35904]_ , \new_[35905]_ ,
    \new_[35908]_ , \new_[35911]_ , \new_[35912]_ , \new_[35913]_ ,
    \new_[35917]_ , \new_[35918]_ , \new_[35921]_ , \new_[35924]_ ,
    \new_[35925]_ , \new_[35926]_ , \new_[35930]_ , \new_[35931]_ ,
    \new_[35934]_ , \new_[35937]_ , \new_[35938]_ , \new_[35939]_ ,
    \new_[35943]_ , \new_[35944]_ , \new_[35947]_ , \new_[35950]_ ,
    \new_[35951]_ , \new_[35952]_ , \new_[35956]_ , \new_[35957]_ ,
    \new_[35960]_ , \new_[35963]_ , \new_[35964]_ , \new_[35965]_ ,
    \new_[35969]_ , \new_[35970]_ , \new_[35973]_ , \new_[35976]_ ,
    \new_[35977]_ , \new_[35978]_ , \new_[35982]_ , \new_[35983]_ ,
    \new_[35986]_ , \new_[35989]_ , \new_[35990]_ , \new_[35991]_ ,
    \new_[35995]_ , \new_[35996]_ , \new_[35999]_ , \new_[36002]_ ,
    \new_[36003]_ , \new_[36004]_ , \new_[36008]_ , \new_[36009]_ ,
    \new_[36012]_ , \new_[36015]_ , \new_[36016]_ , \new_[36017]_ ,
    \new_[36021]_ , \new_[36022]_ , \new_[36025]_ , \new_[36028]_ ,
    \new_[36029]_ , \new_[36030]_ , \new_[36034]_ , \new_[36035]_ ,
    \new_[36038]_ , \new_[36041]_ , \new_[36042]_ , \new_[36043]_ ,
    \new_[36047]_ , \new_[36048]_ , \new_[36051]_ , \new_[36054]_ ,
    \new_[36055]_ , \new_[36056]_ , \new_[36060]_ , \new_[36061]_ ,
    \new_[36064]_ , \new_[36067]_ , \new_[36068]_ , \new_[36069]_ ,
    \new_[36073]_ , \new_[36074]_ , \new_[36077]_ , \new_[36080]_ ,
    \new_[36081]_ , \new_[36082]_ , \new_[36086]_ , \new_[36087]_ ,
    \new_[36090]_ , \new_[36093]_ , \new_[36094]_ , \new_[36095]_ ,
    \new_[36099]_ , \new_[36100]_ , \new_[36103]_ , \new_[36106]_ ,
    \new_[36107]_ , \new_[36108]_ , \new_[36112]_ , \new_[36113]_ ,
    \new_[36116]_ , \new_[36119]_ , \new_[36120]_ , \new_[36121]_ ,
    \new_[36125]_ , \new_[36126]_ , \new_[36129]_ , \new_[36132]_ ,
    \new_[36133]_ , \new_[36134]_ , \new_[36138]_ , \new_[36139]_ ,
    \new_[36142]_ , \new_[36145]_ , \new_[36146]_ , \new_[36147]_ ,
    \new_[36151]_ , \new_[36152]_ , \new_[36155]_ , \new_[36158]_ ,
    \new_[36159]_ , \new_[36160]_ , \new_[36164]_ , \new_[36165]_ ,
    \new_[36168]_ , \new_[36171]_ , \new_[36172]_ , \new_[36173]_ ,
    \new_[36177]_ , \new_[36178]_ , \new_[36181]_ , \new_[36184]_ ,
    \new_[36185]_ , \new_[36186]_ , \new_[36190]_ , \new_[36191]_ ,
    \new_[36194]_ , \new_[36197]_ , \new_[36198]_ , \new_[36199]_ ,
    \new_[36203]_ , \new_[36204]_ , \new_[36207]_ , \new_[36210]_ ,
    \new_[36211]_ , \new_[36212]_ , \new_[36216]_ , \new_[36217]_ ,
    \new_[36220]_ , \new_[36223]_ , \new_[36224]_ , \new_[36225]_ ,
    \new_[36229]_ , \new_[36230]_ , \new_[36233]_ , \new_[36236]_ ,
    \new_[36237]_ , \new_[36238]_ , \new_[36242]_ , \new_[36243]_ ,
    \new_[36246]_ , \new_[36249]_ , \new_[36250]_ , \new_[36251]_ ,
    \new_[36255]_ , \new_[36256]_ , \new_[36259]_ , \new_[36262]_ ,
    \new_[36263]_ , \new_[36264]_ , \new_[36268]_ , \new_[36269]_ ,
    \new_[36272]_ , \new_[36275]_ , \new_[36276]_ , \new_[36277]_ ,
    \new_[36281]_ , \new_[36282]_ , \new_[36285]_ , \new_[36288]_ ,
    \new_[36289]_ , \new_[36290]_ , \new_[36294]_ , \new_[36295]_ ,
    \new_[36298]_ , \new_[36301]_ , \new_[36302]_ , \new_[36303]_ ,
    \new_[36307]_ , \new_[36308]_ , \new_[36311]_ , \new_[36314]_ ,
    \new_[36315]_ , \new_[36316]_ , \new_[36320]_ , \new_[36321]_ ,
    \new_[36324]_ , \new_[36327]_ , \new_[36328]_ , \new_[36329]_ ,
    \new_[36333]_ , \new_[36334]_ , \new_[36337]_ , \new_[36340]_ ,
    \new_[36341]_ , \new_[36342]_ , \new_[36346]_ , \new_[36347]_ ,
    \new_[36350]_ , \new_[36353]_ , \new_[36354]_ , \new_[36355]_ ,
    \new_[36359]_ , \new_[36360]_ , \new_[36363]_ , \new_[36366]_ ,
    \new_[36367]_ , \new_[36368]_ , \new_[36372]_ , \new_[36373]_ ,
    \new_[36376]_ , \new_[36379]_ , \new_[36380]_ , \new_[36381]_ ,
    \new_[36385]_ , \new_[36386]_ , \new_[36389]_ , \new_[36392]_ ,
    \new_[36393]_ , \new_[36394]_ , \new_[36398]_ , \new_[36399]_ ,
    \new_[36402]_ , \new_[36405]_ , \new_[36406]_ , \new_[36407]_ ,
    \new_[36411]_ , \new_[36412]_ , \new_[36415]_ , \new_[36418]_ ,
    \new_[36419]_ , \new_[36420]_ , \new_[36424]_ , \new_[36425]_ ,
    \new_[36428]_ , \new_[36431]_ , \new_[36432]_ , \new_[36433]_ ,
    \new_[36437]_ , \new_[36438]_ , \new_[36441]_ , \new_[36444]_ ,
    \new_[36445]_ , \new_[36446]_ , \new_[36450]_ , \new_[36451]_ ,
    \new_[36454]_ , \new_[36457]_ , \new_[36458]_ , \new_[36459]_ ,
    \new_[36463]_ , \new_[36464]_ , \new_[36467]_ , \new_[36470]_ ,
    \new_[36471]_ , \new_[36472]_ , \new_[36476]_ , \new_[36477]_ ,
    \new_[36480]_ , \new_[36483]_ , \new_[36484]_ , \new_[36485]_ ,
    \new_[36489]_ , \new_[36490]_ , \new_[36493]_ , \new_[36496]_ ,
    \new_[36497]_ , \new_[36498]_ , \new_[36502]_ , \new_[36503]_ ,
    \new_[36506]_ , \new_[36509]_ , \new_[36510]_ , \new_[36511]_ ,
    \new_[36515]_ , \new_[36516]_ , \new_[36519]_ , \new_[36522]_ ,
    \new_[36523]_ , \new_[36524]_ , \new_[36528]_ , \new_[36529]_ ,
    \new_[36532]_ , \new_[36535]_ , \new_[36536]_ , \new_[36537]_ ,
    \new_[36541]_ , \new_[36542]_ , \new_[36545]_ , \new_[36548]_ ,
    \new_[36549]_ , \new_[36550]_ , \new_[36554]_ , \new_[36555]_ ,
    \new_[36558]_ , \new_[36561]_ , \new_[36562]_ , \new_[36563]_ ,
    \new_[36567]_ , \new_[36568]_ , \new_[36571]_ , \new_[36574]_ ,
    \new_[36575]_ , \new_[36576]_ , \new_[36580]_ , \new_[36581]_ ,
    \new_[36584]_ , \new_[36587]_ , \new_[36588]_ , \new_[36589]_ ,
    \new_[36593]_ , \new_[36594]_ , \new_[36597]_ , \new_[36600]_ ,
    \new_[36601]_ , \new_[36602]_ , \new_[36606]_ , \new_[36607]_ ,
    \new_[36610]_ , \new_[36613]_ , \new_[36614]_ , \new_[36615]_ ,
    \new_[36619]_ , \new_[36620]_ , \new_[36623]_ , \new_[36626]_ ,
    \new_[36627]_ , \new_[36628]_ , \new_[36632]_ , \new_[36633]_ ,
    \new_[36636]_ , \new_[36639]_ , \new_[36640]_ , \new_[36641]_ ,
    \new_[36645]_ , \new_[36646]_ , \new_[36649]_ , \new_[36652]_ ,
    \new_[36653]_ , \new_[36654]_ , \new_[36658]_ , \new_[36659]_ ,
    \new_[36662]_ , \new_[36665]_ , \new_[36666]_ , \new_[36667]_ ,
    \new_[36671]_ , \new_[36672]_ , \new_[36675]_ , \new_[36678]_ ,
    \new_[36679]_ , \new_[36680]_ , \new_[36684]_ , \new_[36685]_ ,
    \new_[36688]_ , \new_[36691]_ , \new_[36692]_ , \new_[36693]_ ,
    \new_[36697]_ , \new_[36698]_ , \new_[36701]_ , \new_[36704]_ ,
    \new_[36705]_ , \new_[36706]_ , \new_[36710]_ , \new_[36711]_ ,
    \new_[36714]_ , \new_[36717]_ , \new_[36718]_ , \new_[36719]_ ,
    \new_[36723]_ , \new_[36724]_ , \new_[36727]_ , \new_[36730]_ ,
    \new_[36731]_ , \new_[36732]_ , \new_[36736]_ , \new_[36737]_ ,
    \new_[36740]_ , \new_[36743]_ , \new_[36744]_ , \new_[36745]_ ,
    \new_[36749]_ , \new_[36750]_ , \new_[36753]_ , \new_[36756]_ ,
    \new_[36757]_ , \new_[36758]_ , \new_[36762]_ , \new_[36763]_ ,
    \new_[36766]_ , \new_[36769]_ , \new_[36770]_ , \new_[36771]_ ,
    \new_[36775]_ , \new_[36776]_ , \new_[36779]_ , \new_[36782]_ ,
    \new_[36783]_ , \new_[36784]_ , \new_[36788]_ , \new_[36789]_ ,
    \new_[36792]_ , \new_[36795]_ , \new_[36796]_ , \new_[36797]_ ,
    \new_[36801]_ , \new_[36802]_ , \new_[36805]_ , \new_[36808]_ ,
    \new_[36809]_ , \new_[36810]_ , \new_[36814]_ , \new_[36815]_ ,
    \new_[36818]_ , \new_[36821]_ , \new_[36822]_ , \new_[36823]_ ,
    \new_[36827]_ , \new_[36828]_ , \new_[36831]_ , \new_[36834]_ ,
    \new_[36835]_ , \new_[36836]_ , \new_[36840]_ , \new_[36841]_ ,
    \new_[36844]_ , \new_[36847]_ , \new_[36848]_ , \new_[36849]_ ,
    \new_[36853]_ , \new_[36854]_ , \new_[36857]_ , \new_[36860]_ ,
    \new_[36861]_ , \new_[36862]_ , \new_[36866]_ , \new_[36867]_ ,
    \new_[36870]_ , \new_[36873]_ , \new_[36874]_ , \new_[36875]_ ,
    \new_[36879]_ , \new_[36880]_ , \new_[36883]_ , \new_[36886]_ ,
    \new_[36887]_ , \new_[36888]_ , \new_[36892]_ , \new_[36893]_ ,
    \new_[36896]_ , \new_[36899]_ , \new_[36900]_ , \new_[36901]_ ,
    \new_[36905]_ , \new_[36906]_ , \new_[36909]_ , \new_[36912]_ ,
    \new_[36913]_ , \new_[36914]_ , \new_[36918]_ , \new_[36919]_ ,
    \new_[36922]_ , \new_[36925]_ , \new_[36926]_ , \new_[36927]_ ,
    \new_[36931]_ , \new_[36932]_ , \new_[36935]_ , \new_[36938]_ ,
    \new_[36939]_ , \new_[36940]_ , \new_[36944]_ , \new_[36945]_ ,
    \new_[36948]_ , \new_[36951]_ , \new_[36952]_ , \new_[36953]_ ,
    \new_[36957]_ , \new_[36958]_ , \new_[36961]_ , \new_[36964]_ ,
    \new_[36965]_ , \new_[36966]_ , \new_[36970]_ , \new_[36971]_ ,
    \new_[36974]_ , \new_[36977]_ , \new_[36978]_ , \new_[36979]_ ,
    \new_[36983]_ , \new_[36984]_ , \new_[36987]_ , \new_[36990]_ ,
    \new_[36991]_ , \new_[36992]_ , \new_[36996]_ , \new_[36997]_ ,
    \new_[37000]_ , \new_[37003]_ , \new_[37004]_ , \new_[37005]_ ,
    \new_[37009]_ , \new_[37010]_ , \new_[37013]_ , \new_[37016]_ ,
    \new_[37017]_ , \new_[37018]_ , \new_[37022]_ , \new_[37023]_ ,
    \new_[37026]_ , \new_[37029]_ , \new_[37030]_ , \new_[37031]_ ,
    \new_[37035]_ , \new_[37036]_ , \new_[37039]_ , \new_[37042]_ ,
    \new_[37043]_ , \new_[37044]_ , \new_[37048]_ , \new_[37049]_ ,
    \new_[37052]_ , \new_[37055]_ , \new_[37056]_ , \new_[37057]_ ,
    \new_[37061]_ , \new_[37062]_ , \new_[37065]_ , \new_[37068]_ ,
    \new_[37069]_ , \new_[37070]_ , \new_[37074]_ , \new_[37075]_ ,
    \new_[37078]_ , \new_[37081]_ , \new_[37082]_ , \new_[37083]_ ,
    \new_[37087]_ , \new_[37088]_ , \new_[37091]_ , \new_[37094]_ ,
    \new_[37095]_ , \new_[37096]_ , \new_[37100]_ , \new_[37101]_ ,
    \new_[37104]_ , \new_[37107]_ , \new_[37108]_ , \new_[37109]_ ,
    \new_[37113]_ , \new_[37114]_ , \new_[37117]_ , \new_[37120]_ ,
    \new_[37121]_ , \new_[37122]_ , \new_[37126]_ , \new_[37127]_ ,
    \new_[37130]_ , \new_[37133]_ , \new_[37134]_ , \new_[37135]_ ,
    \new_[37139]_ , \new_[37140]_ , \new_[37143]_ , \new_[37146]_ ,
    \new_[37147]_ , \new_[37148]_ , \new_[37152]_ , \new_[37153]_ ,
    \new_[37156]_ , \new_[37159]_ , \new_[37160]_ , \new_[37161]_ ,
    \new_[37165]_ , \new_[37166]_ , \new_[37169]_ , \new_[37172]_ ,
    \new_[37173]_ , \new_[37174]_ , \new_[37178]_ , \new_[37179]_ ,
    \new_[37182]_ , \new_[37185]_ , \new_[37186]_ , \new_[37187]_ ,
    \new_[37191]_ , \new_[37192]_ , \new_[37195]_ , \new_[37198]_ ,
    \new_[37199]_ , \new_[37200]_ , \new_[37204]_ , \new_[37205]_ ,
    \new_[37208]_ , \new_[37211]_ , \new_[37212]_ , \new_[37213]_ ,
    \new_[37217]_ , \new_[37218]_ , \new_[37221]_ , \new_[37224]_ ,
    \new_[37225]_ , \new_[37226]_ , \new_[37230]_ , \new_[37231]_ ,
    \new_[37234]_ , \new_[37237]_ , \new_[37238]_ , \new_[37239]_ ,
    \new_[37243]_ , \new_[37244]_ , \new_[37247]_ , \new_[37250]_ ,
    \new_[37251]_ , \new_[37252]_ , \new_[37256]_ , \new_[37257]_ ,
    \new_[37260]_ , \new_[37263]_ , \new_[37264]_ , \new_[37265]_ ,
    \new_[37269]_ , \new_[37270]_ , \new_[37273]_ , \new_[37276]_ ,
    \new_[37277]_ , \new_[37278]_ , \new_[37282]_ , \new_[37283]_ ,
    \new_[37286]_ , \new_[37289]_ , \new_[37290]_ , \new_[37291]_ ,
    \new_[37295]_ , \new_[37296]_ , \new_[37299]_ , \new_[37302]_ ,
    \new_[37303]_ , \new_[37304]_ , \new_[37308]_ , \new_[37309]_ ,
    \new_[37312]_ , \new_[37315]_ , \new_[37316]_ , \new_[37317]_ ,
    \new_[37321]_ , \new_[37322]_ , \new_[37325]_ , \new_[37328]_ ,
    \new_[37329]_ , \new_[37330]_ , \new_[37334]_ , \new_[37335]_ ,
    \new_[37338]_ , \new_[37341]_ , \new_[37342]_ , \new_[37343]_ ,
    \new_[37347]_ , \new_[37348]_ , \new_[37351]_ , \new_[37354]_ ,
    \new_[37355]_ , \new_[37356]_ , \new_[37360]_ , \new_[37361]_ ,
    \new_[37364]_ , \new_[37367]_ , \new_[37368]_ , \new_[37369]_ ,
    \new_[37373]_ , \new_[37374]_ , \new_[37377]_ , \new_[37380]_ ,
    \new_[37381]_ , \new_[37382]_ , \new_[37386]_ , \new_[37387]_ ,
    \new_[37390]_ , \new_[37393]_ , \new_[37394]_ , \new_[37395]_ ,
    \new_[37399]_ , \new_[37400]_ , \new_[37403]_ , \new_[37406]_ ,
    \new_[37407]_ , \new_[37408]_ , \new_[37412]_ , \new_[37413]_ ,
    \new_[37416]_ , \new_[37419]_ , \new_[37420]_ , \new_[37421]_ ,
    \new_[37425]_ , \new_[37426]_ , \new_[37429]_ , \new_[37432]_ ,
    \new_[37433]_ , \new_[37434]_ , \new_[37438]_ , \new_[37439]_ ,
    \new_[37442]_ , \new_[37445]_ , \new_[37446]_ , \new_[37447]_ ,
    \new_[37451]_ , \new_[37452]_ , \new_[37455]_ , \new_[37458]_ ,
    \new_[37459]_ , \new_[37460]_ , \new_[37464]_ , \new_[37465]_ ,
    \new_[37468]_ , \new_[37471]_ , \new_[37472]_ , \new_[37473]_ ,
    \new_[37477]_ , \new_[37478]_ , \new_[37481]_ , \new_[37484]_ ,
    \new_[37485]_ , \new_[37486]_ , \new_[37490]_ , \new_[37491]_ ,
    \new_[37494]_ , \new_[37497]_ , \new_[37498]_ , \new_[37499]_ ,
    \new_[37503]_ , \new_[37504]_ , \new_[37507]_ , \new_[37510]_ ,
    \new_[37511]_ , \new_[37512]_ , \new_[37516]_ , \new_[37517]_ ,
    \new_[37520]_ , \new_[37523]_ , \new_[37524]_ , \new_[37525]_ ,
    \new_[37529]_ , \new_[37530]_ , \new_[37533]_ , \new_[37536]_ ,
    \new_[37537]_ , \new_[37538]_ , \new_[37542]_ , \new_[37543]_ ,
    \new_[37546]_ , \new_[37549]_ , \new_[37550]_ , \new_[37551]_ ,
    \new_[37555]_ , \new_[37556]_ , \new_[37559]_ , \new_[37562]_ ,
    \new_[37563]_ , \new_[37564]_ , \new_[37568]_ , \new_[37569]_ ,
    \new_[37572]_ , \new_[37575]_ , \new_[37576]_ , \new_[37577]_ ,
    \new_[37581]_ , \new_[37582]_ , \new_[37585]_ , \new_[37588]_ ,
    \new_[37589]_ , \new_[37590]_ , \new_[37594]_ , \new_[37595]_ ,
    \new_[37598]_ , \new_[37601]_ , \new_[37602]_ , \new_[37603]_ ,
    \new_[37607]_ , \new_[37608]_ , \new_[37611]_ , \new_[37614]_ ,
    \new_[37615]_ , \new_[37616]_ , \new_[37620]_ , \new_[37621]_ ,
    \new_[37624]_ , \new_[37627]_ , \new_[37628]_ , \new_[37629]_ ,
    \new_[37633]_ , \new_[37634]_ , \new_[37637]_ , \new_[37640]_ ,
    \new_[37641]_ , \new_[37642]_ , \new_[37646]_ , \new_[37647]_ ,
    \new_[37650]_ , \new_[37653]_ , \new_[37654]_ , \new_[37655]_ ,
    \new_[37659]_ , \new_[37660]_ , \new_[37663]_ , \new_[37666]_ ,
    \new_[37667]_ , \new_[37668]_ , \new_[37672]_ , \new_[37673]_ ,
    \new_[37676]_ , \new_[37679]_ , \new_[37680]_ , \new_[37681]_ ,
    \new_[37685]_ , \new_[37686]_ , \new_[37689]_ , \new_[37692]_ ,
    \new_[37693]_ , \new_[37694]_ , \new_[37698]_ , \new_[37699]_ ,
    \new_[37702]_ , \new_[37705]_ , \new_[37706]_ , \new_[37707]_ ,
    \new_[37711]_ , \new_[37712]_ , \new_[37715]_ , \new_[37718]_ ,
    \new_[37719]_ , \new_[37720]_ , \new_[37724]_ , \new_[37725]_ ,
    \new_[37728]_ , \new_[37731]_ , \new_[37732]_ , \new_[37733]_ ,
    \new_[37737]_ , \new_[37738]_ , \new_[37741]_ , \new_[37744]_ ,
    \new_[37745]_ , \new_[37746]_ , \new_[37750]_ , \new_[37751]_ ,
    \new_[37754]_ , \new_[37757]_ , \new_[37758]_ , \new_[37759]_ ,
    \new_[37763]_ , \new_[37764]_ , \new_[37767]_ , \new_[37770]_ ,
    \new_[37771]_ , \new_[37772]_ , \new_[37776]_ , \new_[37777]_ ,
    \new_[37780]_ , \new_[37783]_ , \new_[37784]_ , \new_[37785]_ ,
    \new_[37789]_ , \new_[37790]_ , \new_[37793]_ , \new_[37796]_ ,
    \new_[37797]_ , \new_[37798]_ , \new_[37802]_ , \new_[37803]_ ,
    \new_[37806]_ , \new_[37809]_ , \new_[37810]_ , \new_[37811]_ ,
    \new_[37815]_ , \new_[37816]_ , \new_[37819]_ , \new_[37822]_ ,
    \new_[37823]_ , \new_[37824]_ , \new_[37828]_ , \new_[37829]_ ,
    \new_[37832]_ , \new_[37835]_ , \new_[37836]_ , \new_[37837]_ ,
    \new_[37840]_ , \new_[37843]_ , \new_[37844]_ , \new_[37847]_ ,
    \new_[37850]_ , \new_[37851]_ , \new_[37852]_ , \new_[37856]_ ,
    \new_[37857]_ , \new_[37860]_ , \new_[37863]_ , \new_[37864]_ ,
    \new_[37865]_ , \new_[37868]_ , \new_[37871]_ , \new_[37872]_ ,
    \new_[37875]_ , \new_[37878]_ , \new_[37879]_ , \new_[37880]_ ,
    \new_[37884]_ , \new_[37885]_ , \new_[37888]_ , \new_[37891]_ ,
    \new_[37892]_ , \new_[37893]_ , \new_[37896]_ , \new_[37899]_ ,
    \new_[37900]_ , \new_[37903]_ , \new_[37906]_ , \new_[37907]_ ,
    \new_[37908]_ , \new_[37912]_ , \new_[37913]_ , \new_[37916]_ ,
    \new_[37919]_ , \new_[37920]_ , \new_[37921]_ , \new_[37924]_ ,
    \new_[37927]_ , \new_[37928]_ , \new_[37931]_ , \new_[37934]_ ,
    \new_[37935]_ , \new_[37936]_ , \new_[37940]_ , \new_[37941]_ ,
    \new_[37944]_ , \new_[37947]_ , \new_[37948]_ , \new_[37949]_ ,
    \new_[37952]_ , \new_[37955]_ , \new_[37956]_ , \new_[37959]_ ,
    \new_[37962]_ , \new_[37963]_ , \new_[37964]_ , \new_[37968]_ ,
    \new_[37969]_ , \new_[37972]_ , \new_[37975]_ , \new_[37976]_ ,
    \new_[37977]_ , \new_[37980]_ , \new_[37983]_ , \new_[37984]_ ,
    \new_[37987]_ , \new_[37990]_ , \new_[37991]_ , \new_[37992]_ ,
    \new_[37996]_ , \new_[37997]_ , \new_[38000]_ , \new_[38003]_ ,
    \new_[38004]_ , \new_[38005]_ , \new_[38008]_ , \new_[38011]_ ,
    \new_[38012]_ , \new_[38015]_ , \new_[38018]_ , \new_[38019]_ ,
    \new_[38020]_ , \new_[38024]_ , \new_[38025]_ , \new_[38028]_ ,
    \new_[38031]_ , \new_[38032]_ , \new_[38033]_ , \new_[38036]_ ,
    \new_[38039]_ , \new_[38040]_ , \new_[38043]_ , \new_[38046]_ ,
    \new_[38047]_ , \new_[38048]_ , \new_[38052]_ , \new_[38053]_ ,
    \new_[38056]_ , \new_[38059]_ , \new_[38060]_ , \new_[38061]_ ,
    \new_[38064]_ , \new_[38067]_ , \new_[38068]_ , \new_[38071]_ ,
    \new_[38074]_ , \new_[38075]_ , \new_[38076]_ , \new_[38080]_ ,
    \new_[38081]_ , \new_[38084]_ , \new_[38087]_ , \new_[38088]_ ,
    \new_[38089]_ , \new_[38092]_ , \new_[38095]_ , \new_[38096]_ ,
    \new_[38099]_ , \new_[38102]_ , \new_[38103]_ , \new_[38104]_ ,
    \new_[38108]_ , \new_[38109]_ , \new_[38112]_ , \new_[38115]_ ,
    \new_[38116]_ , \new_[38117]_ , \new_[38120]_ , \new_[38123]_ ,
    \new_[38124]_ , \new_[38127]_ , \new_[38130]_ , \new_[38131]_ ,
    \new_[38132]_ , \new_[38136]_ , \new_[38137]_ , \new_[38140]_ ,
    \new_[38143]_ , \new_[38144]_ , \new_[38145]_ , \new_[38148]_ ,
    \new_[38151]_ , \new_[38152]_ , \new_[38155]_ , \new_[38158]_ ,
    \new_[38159]_ , \new_[38160]_ , \new_[38164]_ , \new_[38165]_ ,
    \new_[38168]_ , \new_[38171]_ , \new_[38172]_ , \new_[38173]_ ,
    \new_[38176]_ , \new_[38179]_ , \new_[38180]_ , \new_[38183]_ ,
    \new_[38186]_ , \new_[38187]_ , \new_[38188]_ , \new_[38192]_ ,
    \new_[38193]_ , \new_[38196]_ , \new_[38199]_ , \new_[38200]_ ,
    \new_[38201]_ , \new_[38204]_ , \new_[38207]_ , \new_[38208]_ ,
    \new_[38211]_ , \new_[38214]_ , \new_[38215]_ , \new_[38216]_ ,
    \new_[38220]_ , \new_[38221]_ , \new_[38224]_ , \new_[38227]_ ,
    \new_[38228]_ , \new_[38229]_ , \new_[38232]_ , \new_[38235]_ ,
    \new_[38236]_ , \new_[38239]_ , \new_[38242]_ , \new_[38243]_ ,
    \new_[38244]_ , \new_[38248]_ , \new_[38249]_ , \new_[38252]_ ,
    \new_[38255]_ , \new_[38256]_ , \new_[38257]_ , \new_[38260]_ ,
    \new_[38263]_ , \new_[38264]_ , \new_[38267]_ , \new_[38270]_ ,
    \new_[38271]_ , \new_[38272]_ , \new_[38276]_ , \new_[38277]_ ,
    \new_[38280]_ , \new_[38283]_ , \new_[38284]_ , \new_[38285]_ ,
    \new_[38288]_ , \new_[38291]_ , \new_[38292]_ , \new_[38295]_ ,
    \new_[38298]_ , \new_[38299]_ , \new_[38300]_ , \new_[38304]_ ,
    \new_[38305]_ , \new_[38308]_ , \new_[38311]_ , \new_[38312]_ ,
    \new_[38313]_ , \new_[38316]_ , \new_[38319]_ , \new_[38320]_ ,
    \new_[38323]_ , \new_[38326]_ , \new_[38327]_ , \new_[38328]_ ,
    \new_[38332]_ , \new_[38333]_ , \new_[38336]_ , \new_[38339]_ ,
    \new_[38340]_ , \new_[38341]_ , \new_[38344]_ , \new_[38347]_ ,
    \new_[38348]_ , \new_[38351]_ , \new_[38354]_ , \new_[38355]_ ,
    \new_[38356]_ , \new_[38360]_ , \new_[38361]_ , \new_[38364]_ ,
    \new_[38367]_ , \new_[38368]_ , \new_[38369]_ , \new_[38372]_ ,
    \new_[38375]_ , \new_[38376]_ , \new_[38379]_ , \new_[38382]_ ,
    \new_[38383]_ , \new_[38384]_ , \new_[38388]_ , \new_[38389]_ ,
    \new_[38392]_ , \new_[38395]_ , \new_[38396]_ , \new_[38397]_ ,
    \new_[38400]_ , \new_[38403]_ , \new_[38404]_ , \new_[38407]_ ,
    \new_[38410]_ , \new_[38411]_ , \new_[38412]_ , \new_[38416]_ ,
    \new_[38417]_ , \new_[38420]_ , \new_[38423]_ , \new_[38424]_ ,
    \new_[38425]_ , \new_[38428]_ , \new_[38431]_ , \new_[38432]_ ,
    \new_[38435]_ , \new_[38438]_ , \new_[38439]_ , \new_[38440]_ ,
    \new_[38444]_ , \new_[38445]_ , \new_[38448]_ , \new_[38451]_ ,
    \new_[38452]_ , \new_[38453]_ , \new_[38456]_ , \new_[38459]_ ,
    \new_[38460]_ , \new_[38463]_ , \new_[38466]_ , \new_[38467]_ ,
    \new_[38468]_ , \new_[38472]_ , \new_[38473]_ , \new_[38476]_ ,
    \new_[38479]_ , \new_[38480]_ , \new_[38481]_ , \new_[38484]_ ,
    \new_[38487]_ , \new_[38488]_ , \new_[38491]_ , \new_[38494]_ ,
    \new_[38495]_ , \new_[38496]_ , \new_[38500]_ , \new_[38501]_ ,
    \new_[38504]_ , \new_[38507]_ , \new_[38508]_ , \new_[38509]_ ,
    \new_[38512]_ , \new_[38515]_ , \new_[38516]_ , \new_[38519]_ ,
    \new_[38522]_ , \new_[38523]_ , \new_[38524]_ , \new_[38528]_ ,
    \new_[38529]_ , \new_[38532]_ , \new_[38535]_ , \new_[38536]_ ,
    \new_[38537]_ , \new_[38540]_ , \new_[38543]_ , \new_[38544]_ ,
    \new_[38547]_ , \new_[38550]_ , \new_[38551]_ , \new_[38552]_ ,
    \new_[38556]_ , \new_[38557]_ , \new_[38560]_ , \new_[38563]_ ,
    \new_[38564]_ , \new_[38565]_ , \new_[38568]_ , \new_[38571]_ ,
    \new_[38572]_ , \new_[38575]_ , \new_[38578]_ , \new_[38579]_ ,
    \new_[38580]_ , \new_[38584]_ , \new_[38585]_ , \new_[38588]_ ,
    \new_[38591]_ , \new_[38592]_ , \new_[38593]_ , \new_[38596]_ ,
    \new_[38599]_ , \new_[38600]_ , \new_[38603]_ , \new_[38606]_ ,
    \new_[38607]_ , \new_[38608]_ , \new_[38612]_ , \new_[38613]_ ,
    \new_[38616]_ , \new_[38619]_ , \new_[38620]_ , \new_[38621]_ ,
    \new_[38624]_ , \new_[38627]_ , \new_[38628]_ , \new_[38631]_ ,
    \new_[38634]_ , \new_[38635]_ , \new_[38636]_ , \new_[38640]_ ,
    \new_[38641]_ , \new_[38644]_ , \new_[38647]_ , \new_[38648]_ ,
    \new_[38649]_ , \new_[38652]_ , \new_[38655]_ , \new_[38656]_ ,
    \new_[38659]_ , \new_[38662]_ , \new_[38663]_ , \new_[38664]_ ,
    \new_[38668]_ , \new_[38669]_ , \new_[38672]_ , \new_[38675]_ ,
    \new_[38676]_ , \new_[38677]_ , \new_[38680]_ , \new_[38683]_ ,
    \new_[38684]_ , \new_[38687]_ , \new_[38690]_ , \new_[38691]_ ,
    \new_[38692]_ , \new_[38696]_ , \new_[38697]_ , \new_[38700]_ ,
    \new_[38703]_ , \new_[38704]_ , \new_[38705]_ , \new_[38708]_ ,
    \new_[38711]_ , \new_[38712]_ , \new_[38715]_ , \new_[38718]_ ,
    \new_[38719]_ , \new_[38720]_ , \new_[38724]_ , \new_[38725]_ ,
    \new_[38728]_ , \new_[38731]_ , \new_[38732]_ , \new_[38733]_ ,
    \new_[38736]_ , \new_[38739]_ , \new_[38740]_ , \new_[38743]_ ,
    \new_[38746]_ , \new_[38747]_ , \new_[38748]_ , \new_[38752]_ ,
    \new_[38753]_ , \new_[38756]_ , \new_[38759]_ , \new_[38760]_ ,
    \new_[38761]_ , \new_[38764]_ , \new_[38767]_ , \new_[38768]_ ,
    \new_[38771]_ , \new_[38774]_ , \new_[38775]_ , \new_[38776]_ ,
    \new_[38780]_ , \new_[38781]_ , \new_[38784]_ , \new_[38787]_ ,
    \new_[38788]_ , \new_[38789]_ , \new_[38792]_ , \new_[38795]_ ,
    \new_[38796]_ , \new_[38799]_ , \new_[38802]_ , \new_[38803]_ ,
    \new_[38804]_ , \new_[38808]_ , \new_[38809]_ , \new_[38812]_ ,
    \new_[38815]_ , \new_[38816]_ , \new_[38817]_ , \new_[38820]_ ,
    \new_[38823]_ , \new_[38824]_ , \new_[38827]_ , \new_[38830]_ ,
    \new_[38831]_ , \new_[38832]_ , \new_[38836]_ , \new_[38837]_ ,
    \new_[38840]_ , \new_[38843]_ , \new_[38844]_ , \new_[38845]_ ,
    \new_[38848]_ , \new_[38851]_ , \new_[38852]_ , \new_[38855]_ ,
    \new_[38858]_ , \new_[38859]_ , \new_[38860]_ , \new_[38864]_ ,
    \new_[38865]_ , \new_[38868]_ , \new_[38871]_ , \new_[38872]_ ,
    \new_[38873]_ , \new_[38876]_ , \new_[38879]_ , \new_[38880]_ ,
    \new_[38883]_ , \new_[38886]_ , \new_[38887]_ , \new_[38888]_ ,
    \new_[38892]_ , \new_[38893]_ , \new_[38896]_ , \new_[38899]_ ,
    \new_[38900]_ , \new_[38901]_ , \new_[38904]_ , \new_[38907]_ ,
    \new_[38908]_ , \new_[38911]_ , \new_[38914]_ , \new_[38915]_ ,
    \new_[38916]_ , \new_[38920]_ , \new_[38921]_ , \new_[38924]_ ,
    \new_[38927]_ , \new_[38928]_ , \new_[38929]_ , \new_[38932]_ ,
    \new_[38935]_ , \new_[38936]_ , \new_[38939]_ , \new_[38942]_ ,
    \new_[38943]_ , \new_[38944]_ , \new_[38948]_ , \new_[38949]_ ,
    \new_[38952]_ , \new_[38955]_ , \new_[38956]_ , \new_[38957]_ ,
    \new_[38960]_ , \new_[38963]_ , \new_[38964]_ , \new_[38967]_ ,
    \new_[38970]_ , \new_[38971]_ , \new_[38972]_ , \new_[38976]_ ,
    \new_[38977]_ , \new_[38980]_ , \new_[38983]_ , \new_[38984]_ ,
    \new_[38985]_ , \new_[38988]_ , \new_[38991]_ , \new_[38992]_ ,
    \new_[38995]_ , \new_[38998]_ , \new_[38999]_ , \new_[39000]_ ,
    \new_[39004]_ , \new_[39005]_ , \new_[39008]_ , \new_[39011]_ ,
    \new_[39012]_ , \new_[39013]_ , \new_[39016]_ , \new_[39019]_ ,
    \new_[39020]_ , \new_[39023]_ , \new_[39026]_ , \new_[39027]_ ,
    \new_[39028]_ , \new_[39032]_ , \new_[39033]_ , \new_[39036]_ ,
    \new_[39039]_ , \new_[39040]_ , \new_[39041]_ , \new_[39044]_ ,
    \new_[39047]_ , \new_[39048]_ , \new_[39051]_ , \new_[39054]_ ,
    \new_[39055]_ , \new_[39056]_ , \new_[39060]_ , \new_[39061]_ ,
    \new_[39064]_ , \new_[39067]_ , \new_[39068]_ , \new_[39069]_ ,
    \new_[39072]_ , \new_[39075]_ , \new_[39076]_ , \new_[39079]_ ,
    \new_[39082]_ , \new_[39083]_ , \new_[39084]_ , \new_[39088]_ ,
    \new_[39089]_ , \new_[39092]_ , \new_[39095]_ , \new_[39096]_ ,
    \new_[39097]_ , \new_[39100]_ , \new_[39103]_ , \new_[39104]_ ,
    \new_[39107]_ , \new_[39110]_ , \new_[39111]_ , \new_[39112]_ ,
    \new_[39116]_ , \new_[39117]_ , \new_[39120]_ , \new_[39123]_ ,
    \new_[39124]_ , \new_[39125]_ , \new_[39128]_ , \new_[39131]_ ,
    \new_[39132]_ , \new_[39135]_ , \new_[39138]_ , \new_[39139]_ ,
    \new_[39140]_ , \new_[39144]_ , \new_[39145]_ , \new_[39148]_ ,
    \new_[39151]_ , \new_[39152]_ , \new_[39153]_ , \new_[39156]_ ,
    \new_[39159]_ , \new_[39160]_ , \new_[39163]_ , \new_[39166]_ ,
    \new_[39167]_ , \new_[39168]_ , \new_[39172]_ , \new_[39173]_ ,
    \new_[39176]_ , \new_[39179]_ , \new_[39180]_ , \new_[39181]_ ,
    \new_[39184]_ , \new_[39187]_ , \new_[39188]_ , \new_[39191]_ ,
    \new_[39194]_ , \new_[39195]_ , \new_[39196]_ , \new_[39200]_ ,
    \new_[39201]_ , \new_[39204]_ , \new_[39207]_ , \new_[39208]_ ,
    \new_[39209]_ , \new_[39212]_ , \new_[39215]_ , \new_[39216]_ ,
    \new_[39219]_ , \new_[39222]_ , \new_[39223]_ , \new_[39224]_ ,
    \new_[39228]_ , \new_[39229]_ , \new_[39232]_ , \new_[39235]_ ,
    \new_[39236]_ , \new_[39237]_ , \new_[39240]_ , \new_[39243]_ ,
    \new_[39244]_ , \new_[39247]_ , \new_[39250]_ , \new_[39251]_ ,
    \new_[39252]_ , \new_[39256]_ , \new_[39257]_ , \new_[39260]_ ,
    \new_[39263]_ , \new_[39264]_ , \new_[39265]_ , \new_[39268]_ ,
    \new_[39271]_ , \new_[39272]_ , \new_[39275]_ , \new_[39278]_ ,
    \new_[39279]_ , \new_[39280]_ , \new_[39284]_ , \new_[39285]_ ,
    \new_[39288]_ , \new_[39291]_ , \new_[39292]_ , \new_[39293]_ ,
    \new_[39296]_ , \new_[39299]_ , \new_[39300]_ , \new_[39303]_ ,
    \new_[39306]_ , \new_[39307]_ , \new_[39308]_ , \new_[39312]_ ,
    \new_[39313]_ , \new_[39316]_ , \new_[39319]_ , \new_[39320]_ ,
    \new_[39321]_ , \new_[39324]_ , \new_[39327]_ , \new_[39328]_ ,
    \new_[39331]_ , \new_[39334]_ , \new_[39335]_ , \new_[39336]_ ,
    \new_[39340]_ , \new_[39341]_ , \new_[39344]_ , \new_[39347]_ ,
    \new_[39348]_ , \new_[39349]_ , \new_[39352]_ , \new_[39355]_ ,
    \new_[39356]_ , \new_[39359]_ , \new_[39362]_ , \new_[39363]_ ,
    \new_[39364]_ , \new_[39368]_ , \new_[39369]_ , \new_[39372]_ ,
    \new_[39375]_ , \new_[39376]_ , \new_[39377]_ , \new_[39380]_ ,
    \new_[39383]_ , \new_[39384]_ , \new_[39387]_ , \new_[39390]_ ,
    \new_[39391]_ , \new_[39392]_ , \new_[39396]_ , \new_[39397]_ ,
    \new_[39400]_ , \new_[39403]_ , \new_[39404]_ , \new_[39405]_ ,
    \new_[39408]_ , \new_[39411]_ , \new_[39412]_ , \new_[39415]_ ,
    \new_[39418]_ , \new_[39419]_ , \new_[39420]_ , \new_[39424]_ ,
    \new_[39425]_ , \new_[39428]_ , \new_[39431]_ , \new_[39432]_ ,
    \new_[39433]_ , \new_[39436]_ , \new_[39439]_ , \new_[39440]_ ,
    \new_[39443]_ , \new_[39446]_ , \new_[39447]_ , \new_[39448]_ ,
    \new_[39452]_ , \new_[39453]_ , \new_[39456]_ , \new_[39459]_ ,
    \new_[39460]_ , \new_[39461]_ , \new_[39464]_ , \new_[39467]_ ,
    \new_[39468]_ , \new_[39471]_ , \new_[39474]_ , \new_[39475]_ ,
    \new_[39476]_ , \new_[39480]_ , \new_[39481]_ , \new_[39484]_ ,
    \new_[39487]_ , \new_[39488]_ , \new_[39489]_ , \new_[39492]_ ,
    \new_[39495]_ , \new_[39496]_ , \new_[39499]_ , \new_[39502]_ ,
    \new_[39503]_ , \new_[39504]_ , \new_[39508]_ , \new_[39509]_ ,
    \new_[39512]_ , \new_[39515]_ , \new_[39516]_ , \new_[39517]_ ,
    \new_[39520]_ , \new_[39523]_ , \new_[39524]_ , \new_[39527]_ ,
    \new_[39530]_ , \new_[39531]_ , \new_[39532]_ , \new_[39536]_ ,
    \new_[39537]_ , \new_[39540]_ , \new_[39543]_ , \new_[39544]_ ,
    \new_[39545]_ , \new_[39548]_ , \new_[39551]_ , \new_[39552]_ ,
    \new_[39555]_ , \new_[39558]_ , \new_[39559]_ , \new_[39560]_ ,
    \new_[39564]_ , \new_[39565]_ , \new_[39568]_ , \new_[39571]_ ,
    \new_[39572]_ , \new_[39573]_ , \new_[39576]_ , \new_[39579]_ ,
    \new_[39580]_ , \new_[39583]_ , \new_[39586]_ , \new_[39587]_ ,
    \new_[39588]_ , \new_[39592]_ , \new_[39593]_ , \new_[39596]_ ,
    \new_[39599]_ , \new_[39600]_ , \new_[39601]_ , \new_[39604]_ ,
    \new_[39607]_ , \new_[39608]_ , \new_[39611]_ , \new_[39614]_ ,
    \new_[39615]_ , \new_[39616]_ , \new_[39620]_ , \new_[39621]_ ,
    \new_[39624]_ , \new_[39627]_ , \new_[39628]_ , \new_[39629]_ ,
    \new_[39632]_ , \new_[39635]_ , \new_[39636]_ , \new_[39639]_ ,
    \new_[39642]_ , \new_[39643]_ , \new_[39644]_ , \new_[39648]_ ,
    \new_[39649]_ , \new_[39652]_ , \new_[39655]_ , \new_[39656]_ ,
    \new_[39657]_ , \new_[39660]_ , \new_[39663]_ , \new_[39664]_ ,
    \new_[39667]_ , \new_[39670]_ , \new_[39671]_ , \new_[39672]_ ,
    \new_[39676]_ , \new_[39677]_ , \new_[39680]_ , \new_[39683]_ ,
    \new_[39684]_ , \new_[39685]_ , \new_[39688]_ , \new_[39691]_ ,
    \new_[39692]_ , \new_[39695]_ , \new_[39698]_ , \new_[39699]_ ,
    \new_[39700]_ , \new_[39704]_ , \new_[39705]_ , \new_[39708]_ ,
    \new_[39711]_ , \new_[39712]_ , \new_[39713]_ , \new_[39716]_ ,
    \new_[39719]_ , \new_[39720]_ , \new_[39723]_ , \new_[39726]_ ,
    \new_[39727]_ , \new_[39728]_ , \new_[39732]_ , \new_[39733]_ ,
    \new_[39736]_ , \new_[39739]_ , \new_[39740]_ , \new_[39741]_ ,
    \new_[39744]_ , \new_[39747]_ , \new_[39748]_ , \new_[39751]_ ,
    \new_[39754]_ , \new_[39755]_ , \new_[39756]_ , \new_[39760]_ ,
    \new_[39761]_ , \new_[39764]_ , \new_[39767]_ , \new_[39768]_ ,
    \new_[39769]_ , \new_[39772]_ , \new_[39775]_ , \new_[39776]_ ,
    \new_[39779]_ , \new_[39782]_ , \new_[39783]_ , \new_[39784]_ ,
    \new_[39788]_ , \new_[39789]_ , \new_[39792]_ , \new_[39795]_ ,
    \new_[39796]_ , \new_[39797]_ , \new_[39800]_ , \new_[39803]_ ,
    \new_[39804]_ , \new_[39807]_ , \new_[39810]_ , \new_[39811]_ ,
    \new_[39812]_ , \new_[39816]_ , \new_[39817]_ , \new_[39820]_ ,
    \new_[39823]_ , \new_[39824]_ , \new_[39825]_ , \new_[39828]_ ,
    \new_[39831]_ , \new_[39832]_ , \new_[39835]_ , \new_[39838]_ ,
    \new_[39839]_ , \new_[39840]_ , \new_[39844]_ , \new_[39845]_ ,
    \new_[39848]_ , \new_[39851]_ , \new_[39852]_ , \new_[39853]_ ,
    \new_[39856]_ , \new_[39859]_ , \new_[39860]_ , \new_[39863]_ ,
    \new_[39866]_ , \new_[39867]_ , \new_[39868]_ , \new_[39872]_ ,
    \new_[39873]_ , \new_[39876]_ , \new_[39879]_ , \new_[39880]_ ,
    \new_[39881]_ , \new_[39884]_ , \new_[39887]_ , \new_[39888]_ ,
    \new_[39891]_ , \new_[39894]_ , \new_[39895]_ , \new_[39896]_ ,
    \new_[39900]_ , \new_[39901]_ , \new_[39904]_ , \new_[39907]_ ,
    \new_[39908]_ , \new_[39909]_ , \new_[39912]_ , \new_[39915]_ ,
    \new_[39916]_ , \new_[39919]_ , \new_[39922]_ , \new_[39923]_ ,
    \new_[39924]_ , \new_[39928]_ , \new_[39929]_ , \new_[39932]_ ,
    \new_[39935]_ , \new_[39936]_ , \new_[39937]_ , \new_[39940]_ ,
    \new_[39943]_ , \new_[39944]_ , \new_[39947]_ , \new_[39950]_ ,
    \new_[39951]_ , \new_[39952]_ , \new_[39956]_ , \new_[39957]_ ,
    \new_[39960]_ , \new_[39963]_ , \new_[39964]_ , \new_[39965]_ ,
    \new_[39968]_ , \new_[39971]_ , \new_[39972]_ , \new_[39975]_ ,
    \new_[39978]_ , \new_[39979]_ , \new_[39980]_ , \new_[39984]_ ,
    \new_[39985]_ , \new_[39988]_ , \new_[39991]_ , \new_[39992]_ ,
    \new_[39993]_ , \new_[39996]_ , \new_[39999]_ , \new_[40000]_ ,
    \new_[40003]_ , \new_[40006]_ , \new_[40007]_ , \new_[40008]_ ,
    \new_[40012]_ , \new_[40013]_ , \new_[40016]_ , \new_[40019]_ ,
    \new_[40020]_ , \new_[40021]_ , \new_[40024]_ , \new_[40027]_ ,
    \new_[40028]_ , \new_[40031]_ , \new_[40034]_ , \new_[40035]_ ,
    \new_[40036]_ , \new_[40040]_ , \new_[40041]_ , \new_[40044]_ ,
    \new_[40047]_ , \new_[40048]_ , \new_[40049]_ , \new_[40052]_ ,
    \new_[40055]_ , \new_[40056]_ , \new_[40059]_ , \new_[40062]_ ,
    \new_[40063]_ , \new_[40064]_ , \new_[40068]_ , \new_[40069]_ ,
    \new_[40072]_ , \new_[40075]_ , \new_[40076]_ , \new_[40077]_ ,
    \new_[40080]_ , \new_[40083]_ , \new_[40084]_ , \new_[40087]_ ,
    \new_[40090]_ , \new_[40091]_ , \new_[40092]_ , \new_[40096]_ ,
    \new_[40097]_ , \new_[40100]_ , \new_[40103]_ , \new_[40104]_ ,
    \new_[40105]_ , \new_[40108]_ , \new_[40111]_ , \new_[40112]_ ,
    \new_[40115]_ , \new_[40118]_ , \new_[40119]_ , \new_[40120]_ ,
    \new_[40124]_ , \new_[40125]_ , \new_[40128]_ , \new_[40131]_ ,
    \new_[40132]_ , \new_[40133]_ , \new_[40136]_ , \new_[40139]_ ,
    \new_[40140]_ , \new_[40143]_ , \new_[40146]_ , \new_[40147]_ ,
    \new_[40148]_ , \new_[40152]_ , \new_[40153]_ , \new_[40156]_ ,
    \new_[40159]_ , \new_[40160]_ , \new_[40161]_ , \new_[40164]_ ,
    \new_[40167]_ , \new_[40168]_ , \new_[40171]_ , \new_[40174]_ ,
    \new_[40175]_ , \new_[40176]_ , \new_[40180]_ , \new_[40181]_ ,
    \new_[40184]_ , \new_[40187]_ , \new_[40188]_ , \new_[40189]_ ,
    \new_[40192]_ , \new_[40195]_ , \new_[40196]_ , \new_[40199]_ ,
    \new_[40202]_ , \new_[40203]_ , \new_[40204]_ , \new_[40208]_ ,
    \new_[40209]_ , \new_[40212]_ , \new_[40215]_ , \new_[40216]_ ,
    \new_[40217]_ , \new_[40220]_ , \new_[40223]_ , \new_[40224]_ ,
    \new_[40227]_ , \new_[40230]_ , \new_[40231]_ , \new_[40232]_ ,
    \new_[40236]_ , \new_[40237]_ , \new_[40240]_ , \new_[40243]_ ,
    \new_[40244]_ , \new_[40245]_ , \new_[40248]_ , \new_[40251]_ ,
    \new_[40252]_ , \new_[40255]_ , \new_[40258]_ , \new_[40259]_ ,
    \new_[40260]_ , \new_[40264]_ , \new_[40265]_ , \new_[40268]_ ,
    \new_[40271]_ , \new_[40272]_ , \new_[40273]_ , \new_[40276]_ ,
    \new_[40279]_ , \new_[40280]_ , \new_[40283]_ , \new_[40286]_ ,
    \new_[40287]_ , \new_[40288]_ , \new_[40292]_ , \new_[40293]_ ,
    \new_[40296]_ , \new_[40299]_ , \new_[40300]_ , \new_[40301]_ ,
    \new_[40304]_ , \new_[40307]_ , \new_[40308]_ , \new_[40311]_ ,
    \new_[40314]_ , \new_[40315]_ , \new_[40316]_ , \new_[40320]_ ,
    \new_[40321]_ , \new_[40324]_ , \new_[40327]_ , \new_[40328]_ ,
    \new_[40329]_ , \new_[40332]_ , \new_[40335]_ , \new_[40336]_ ,
    \new_[40339]_ , \new_[40342]_ , \new_[40343]_ , \new_[40344]_ ,
    \new_[40348]_ , \new_[40349]_ , \new_[40352]_ , \new_[40355]_ ,
    \new_[40356]_ , \new_[40357]_ , \new_[40360]_ , \new_[40363]_ ,
    \new_[40364]_ , \new_[40367]_ , \new_[40370]_ , \new_[40371]_ ,
    \new_[40372]_ , \new_[40376]_ , \new_[40377]_ , \new_[40380]_ ,
    \new_[40383]_ , \new_[40384]_ , \new_[40385]_ , \new_[40388]_ ,
    \new_[40391]_ , \new_[40392]_ , \new_[40395]_ , \new_[40398]_ ,
    \new_[40399]_ , \new_[40400]_ , \new_[40404]_ , \new_[40405]_ ,
    \new_[40408]_ , \new_[40411]_ , \new_[40412]_ , \new_[40413]_ ,
    \new_[40416]_ , \new_[40419]_ , \new_[40420]_ , \new_[40423]_ ,
    \new_[40426]_ , \new_[40427]_ , \new_[40428]_ , \new_[40432]_ ,
    \new_[40433]_ , \new_[40436]_ , \new_[40439]_ , \new_[40440]_ ,
    \new_[40441]_ , \new_[40444]_ , \new_[40447]_ , \new_[40448]_ ,
    \new_[40451]_ , \new_[40454]_ , \new_[40455]_ , \new_[40456]_ ,
    \new_[40460]_ , \new_[40461]_ , \new_[40464]_ , \new_[40467]_ ,
    \new_[40468]_ , \new_[40469]_ , \new_[40472]_ , \new_[40475]_ ,
    \new_[40476]_ , \new_[40479]_ , \new_[40482]_ , \new_[40483]_ ,
    \new_[40484]_ , \new_[40488]_ , \new_[40489]_ , \new_[40492]_ ,
    \new_[40495]_ , \new_[40496]_ , \new_[40497]_ , \new_[40500]_ ,
    \new_[40503]_ , \new_[40504]_ , \new_[40507]_ , \new_[40510]_ ,
    \new_[40511]_ , \new_[40512]_ , \new_[40516]_ , \new_[40517]_ ,
    \new_[40520]_ , \new_[40523]_ , \new_[40524]_ , \new_[40525]_ ,
    \new_[40528]_ , \new_[40531]_ , \new_[40532]_ , \new_[40535]_ ,
    \new_[40538]_ , \new_[40539]_ , \new_[40540]_ , \new_[40544]_ ,
    \new_[40545]_ , \new_[40548]_ , \new_[40551]_ , \new_[40552]_ ,
    \new_[40553]_ , \new_[40556]_ , \new_[40559]_ , \new_[40560]_ ,
    \new_[40563]_ , \new_[40566]_ , \new_[40567]_ , \new_[40568]_ ,
    \new_[40572]_ , \new_[40573]_ , \new_[40576]_ , \new_[40579]_ ,
    \new_[40580]_ , \new_[40581]_ , \new_[40584]_ , \new_[40587]_ ,
    \new_[40588]_ , \new_[40591]_ , \new_[40594]_ , \new_[40595]_ ,
    \new_[40596]_ , \new_[40600]_ , \new_[40601]_ , \new_[40604]_ ,
    \new_[40607]_ , \new_[40608]_ , \new_[40609]_ , \new_[40612]_ ,
    \new_[40615]_ , \new_[40616]_ , \new_[40619]_ , \new_[40622]_ ,
    \new_[40623]_ , \new_[40624]_ , \new_[40628]_ , \new_[40629]_ ,
    \new_[40632]_ , \new_[40635]_ , \new_[40636]_ , \new_[40637]_ ,
    \new_[40640]_ , \new_[40643]_ , \new_[40644]_ , \new_[40647]_ ,
    \new_[40650]_ , \new_[40651]_ , \new_[40652]_ , \new_[40656]_ ,
    \new_[40657]_ , \new_[40660]_ , \new_[40663]_ , \new_[40664]_ ,
    \new_[40665]_ , \new_[40668]_ , \new_[40671]_ , \new_[40672]_ ,
    \new_[40675]_ , \new_[40678]_ , \new_[40679]_ , \new_[40680]_ ,
    \new_[40684]_ , \new_[40685]_ , \new_[40688]_ , \new_[40691]_ ,
    \new_[40692]_ , \new_[40693]_ , \new_[40696]_ , \new_[40699]_ ,
    \new_[40700]_ , \new_[40703]_ , \new_[40706]_ , \new_[40707]_ ,
    \new_[40708]_ , \new_[40712]_ , \new_[40713]_ , \new_[40716]_ ,
    \new_[40719]_ , \new_[40720]_ , \new_[40721]_ , \new_[40724]_ ,
    \new_[40727]_ , \new_[40728]_ , \new_[40731]_ , \new_[40734]_ ,
    \new_[40735]_ , \new_[40736]_ , \new_[40740]_ , \new_[40741]_ ,
    \new_[40744]_ , \new_[40747]_ , \new_[40748]_ , \new_[40749]_ ,
    \new_[40752]_ , \new_[40755]_ , \new_[40756]_ , \new_[40759]_ ,
    \new_[40762]_ , \new_[40763]_ , \new_[40764]_ , \new_[40768]_ ,
    \new_[40769]_ , \new_[40772]_ , \new_[40775]_ , \new_[40776]_ ,
    \new_[40777]_ , \new_[40780]_ , \new_[40783]_ , \new_[40784]_ ,
    \new_[40787]_ , \new_[40790]_ , \new_[40791]_ , \new_[40792]_ ,
    \new_[40796]_ , \new_[40797]_ , \new_[40800]_ , \new_[40803]_ ,
    \new_[40804]_ , \new_[40805]_ , \new_[40808]_ , \new_[40811]_ ,
    \new_[40812]_ , \new_[40815]_ , \new_[40818]_ , \new_[40819]_ ,
    \new_[40820]_ , \new_[40824]_ , \new_[40825]_ , \new_[40828]_ ,
    \new_[40831]_ , \new_[40832]_ , \new_[40833]_ , \new_[40836]_ ,
    \new_[40839]_ , \new_[40840]_ , \new_[40843]_ , \new_[40846]_ ,
    \new_[40847]_ , \new_[40848]_ , \new_[40852]_ , \new_[40853]_ ,
    \new_[40856]_ , \new_[40859]_ , \new_[40860]_ , \new_[40861]_ ,
    \new_[40864]_ , \new_[40867]_ , \new_[40868]_ , \new_[40871]_ ,
    \new_[40874]_ , \new_[40875]_ , \new_[40876]_ , \new_[40880]_ ,
    \new_[40881]_ , \new_[40884]_ , \new_[40887]_ , \new_[40888]_ ,
    \new_[40889]_ , \new_[40892]_ , \new_[40895]_ , \new_[40896]_ ,
    \new_[40899]_ , \new_[40902]_ , \new_[40903]_ , \new_[40904]_ ,
    \new_[40908]_ , \new_[40909]_ , \new_[40912]_ , \new_[40915]_ ,
    \new_[40916]_ , \new_[40917]_ , \new_[40920]_ , \new_[40923]_ ,
    \new_[40924]_ , \new_[40927]_ , \new_[40930]_ , \new_[40931]_ ,
    \new_[40932]_ , \new_[40936]_ , \new_[40937]_ , \new_[40940]_ ,
    \new_[40943]_ , \new_[40944]_ , \new_[40945]_ , \new_[40948]_ ,
    \new_[40951]_ , \new_[40952]_ , \new_[40955]_ , \new_[40958]_ ,
    \new_[40959]_ , \new_[40960]_ , \new_[40964]_ , \new_[40965]_ ,
    \new_[40968]_ , \new_[40971]_ , \new_[40972]_ , \new_[40973]_ ,
    \new_[40976]_ , \new_[40979]_ , \new_[40980]_ , \new_[40983]_ ,
    \new_[40986]_ , \new_[40987]_ , \new_[40988]_ , \new_[40992]_ ,
    \new_[40993]_ , \new_[40996]_ , \new_[40999]_ , \new_[41000]_ ,
    \new_[41001]_ , \new_[41004]_ , \new_[41007]_ , \new_[41008]_ ,
    \new_[41011]_ , \new_[41014]_ , \new_[41015]_ , \new_[41016]_ ,
    \new_[41020]_ , \new_[41021]_ , \new_[41024]_ , \new_[41027]_ ,
    \new_[41028]_ , \new_[41029]_ , \new_[41032]_ , \new_[41035]_ ,
    \new_[41036]_ , \new_[41039]_ , \new_[41042]_ , \new_[41043]_ ,
    \new_[41044]_ , \new_[41048]_ , \new_[41049]_ , \new_[41052]_ ,
    \new_[41055]_ , \new_[41056]_ , \new_[41057]_ , \new_[41060]_ ,
    \new_[41063]_ , \new_[41064]_ , \new_[41067]_ , \new_[41070]_ ,
    \new_[41071]_ , \new_[41072]_ , \new_[41076]_ , \new_[41077]_ ,
    \new_[41080]_ , \new_[41083]_ , \new_[41084]_ , \new_[41085]_ ,
    \new_[41088]_ , \new_[41091]_ , \new_[41092]_ , \new_[41095]_ ,
    \new_[41098]_ , \new_[41099]_ , \new_[41100]_ , \new_[41104]_ ,
    \new_[41105]_ , \new_[41108]_ , \new_[41111]_ , \new_[41112]_ ,
    \new_[41113]_ , \new_[41116]_ , \new_[41119]_ , \new_[41120]_ ,
    \new_[41123]_ , \new_[41126]_ , \new_[41127]_ , \new_[41128]_ ,
    \new_[41132]_ , \new_[41133]_ , \new_[41136]_ , \new_[41139]_ ,
    \new_[41140]_ , \new_[41141]_ , \new_[41144]_ , \new_[41147]_ ,
    \new_[41148]_ , \new_[41151]_ , \new_[41154]_ , \new_[41155]_ ,
    \new_[41156]_ , \new_[41160]_ , \new_[41161]_ , \new_[41164]_ ,
    \new_[41167]_ , \new_[41168]_ , \new_[41169]_ , \new_[41172]_ ,
    \new_[41175]_ , \new_[41176]_ , \new_[41179]_ , \new_[41182]_ ,
    \new_[41183]_ , \new_[41184]_ , \new_[41188]_ , \new_[41189]_ ,
    \new_[41192]_ , \new_[41195]_ , \new_[41196]_ , \new_[41197]_ ,
    \new_[41200]_ , \new_[41203]_ , \new_[41204]_ , \new_[41207]_ ,
    \new_[41210]_ , \new_[41211]_ , \new_[41212]_ , \new_[41216]_ ,
    \new_[41217]_ , \new_[41220]_ , \new_[41223]_ , \new_[41224]_ ,
    \new_[41225]_ , \new_[41228]_ , \new_[41231]_ , \new_[41232]_ ,
    \new_[41235]_ , \new_[41238]_ , \new_[41239]_ , \new_[41240]_ ,
    \new_[41244]_ , \new_[41245]_ , \new_[41248]_ , \new_[41251]_ ,
    \new_[41252]_ , \new_[41253]_ , \new_[41256]_ , \new_[41259]_ ,
    \new_[41260]_ , \new_[41263]_ , \new_[41266]_ , \new_[41267]_ ,
    \new_[41268]_ , \new_[41272]_ , \new_[41273]_ , \new_[41276]_ ,
    \new_[41279]_ , \new_[41280]_ , \new_[41281]_ , \new_[41284]_ ,
    \new_[41287]_ , \new_[41288]_ , \new_[41291]_ , \new_[41294]_ ,
    \new_[41295]_ , \new_[41296]_ , \new_[41300]_ , \new_[41301]_ ,
    \new_[41304]_ , \new_[41307]_ , \new_[41308]_ , \new_[41309]_ ,
    \new_[41312]_ , \new_[41315]_ , \new_[41316]_ , \new_[41319]_ ,
    \new_[41322]_ , \new_[41323]_ , \new_[41324]_ , \new_[41328]_ ,
    \new_[41329]_ , \new_[41332]_ , \new_[41335]_ , \new_[41336]_ ,
    \new_[41337]_ , \new_[41340]_ , \new_[41343]_ , \new_[41344]_ ,
    \new_[41347]_ , \new_[41350]_ , \new_[41351]_ , \new_[41352]_ ,
    \new_[41356]_ , \new_[41357]_ , \new_[41360]_ , \new_[41363]_ ,
    \new_[41364]_ , \new_[41365]_ , \new_[41368]_ , \new_[41371]_ ,
    \new_[41372]_ , \new_[41375]_ , \new_[41378]_ , \new_[41379]_ ,
    \new_[41380]_ , \new_[41384]_ , \new_[41385]_ , \new_[41388]_ ,
    \new_[41391]_ , \new_[41392]_ , \new_[41393]_ , \new_[41396]_ ,
    \new_[41399]_ , \new_[41400]_ , \new_[41403]_ , \new_[41406]_ ,
    \new_[41407]_ , \new_[41408]_ , \new_[41412]_ , \new_[41413]_ ,
    \new_[41416]_ , \new_[41419]_ , \new_[41420]_ , \new_[41421]_ ,
    \new_[41424]_ , \new_[41427]_ , \new_[41428]_ , \new_[41431]_ ,
    \new_[41434]_ , \new_[41435]_ , \new_[41436]_ , \new_[41440]_ ,
    \new_[41441]_ , \new_[41444]_ , \new_[41447]_ , \new_[41448]_ ,
    \new_[41449]_ , \new_[41452]_ , \new_[41455]_ , \new_[41456]_ ,
    \new_[41459]_ , \new_[41462]_ , \new_[41463]_ , \new_[41464]_ ,
    \new_[41468]_ , \new_[41469]_ , \new_[41472]_ , \new_[41475]_ ,
    \new_[41476]_ , \new_[41477]_ , \new_[41480]_ , \new_[41483]_ ,
    \new_[41484]_ , \new_[41487]_ , \new_[41490]_ , \new_[41491]_ ,
    \new_[41492]_ , \new_[41496]_ , \new_[41497]_ , \new_[41500]_ ,
    \new_[41503]_ , \new_[41504]_ , \new_[41505]_ , \new_[41508]_ ,
    \new_[41511]_ , \new_[41512]_ , \new_[41515]_ , \new_[41518]_ ,
    \new_[41519]_ , \new_[41520]_ , \new_[41524]_ , \new_[41525]_ ,
    \new_[41528]_ , \new_[41531]_ , \new_[41532]_ , \new_[41533]_ ,
    \new_[41536]_ , \new_[41539]_ , \new_[41540]_ , \new_[41543]_ ,
    \new_[41546]_ , \new_[41547]_ , \new_[41548]_ , \new_[41552]_ ,
    \new_[41553]_ , \new_[41556]_ , \new_[41559]_ , \new_[41560]_ ,
    \new_[41561]_ , \new_[41564]_ , \new_[41567]_ , \new_[41568]_ ,
    \new_[41571]_ , \new_[41574]_ , \new_[41575]_ , \new_[41576]_ ,
    \new_[41580]_ , \new_[41581]_ , \new_[41584]_ , \new_[41587]_ ,
    \new_[41588]_ , \new_[41589]_ , \new_[41592]_ , \new_[41595]_ ,
    \new_[41596]_ , \new_[41599]_ , \new_[41602]_ , \new_[41603]_ ,
    \new_[41604]_ , \new_[41608]_ , \new_[41609]_ , \new_[41612]_ ,
    \new_[41615]_ , \new_[41616]_ , \new_[41617]_ , \new_[41620]_ ,
    \new_[41623]_ , \new_[41624]_ , \new_[41627]_ , \new_[41630]_ ,
    \new_[41631]_ , \new_[41632]_ , \new_[41636]_ , \new_[41637]_ ,
    \new_[41640]_ , \new_[41643]_ , \new_[41644]_ , \new_[41645]_ ,
    \new_[41648]_ , \new_[41651]_ , \new_[41652]_ , \new_[41655]_ ,
    \new_[41658]_ , \new_[41659]_ , \new_[41660]_ , \new_[41664]_ ,
    \new_[41665]_ , \new_[41668]_ , \new_[41671]_ , \new_[41672]_ ,
    \new_[41673]_ , \new_[41676]_ , \new_[41679]_ , \new_[41680]_ ,
    \new_[41683]_ , \new_[41686]_ , \new_[41687]_ , \new_[41688]_ ,
    \new_[41692]_ , \new_[41693]_ , \new_[41696]_ , \new_[41699]_ ,
    \new_[41700]_ , \new_[41701]_ , \new_[41704]_ , \new_[41707]_ ,
    \new_[41708]_ , \new_[41711]_ , \new_[41714]_ , \new_[41715]_ ,
    \new_[41716]_ , \new_[41720]_ , \new_[41721]_ , \new_[41724]_ ,
    \new_[41727]_ , \new_[41728]_ , \new_[41729]_ , \new_[41732]_ ,
    \new_[41735]_ , \new_[41736]_ , \new_[41739]_ , \new_[41742]_ ,
    \new_[41743]_ , \new_[41744]_ , \new_[41748]_ , \new_[41749]_ ,
    \new_[41752]_ , \new_[41755]_ , \new_[41756]_ , \new_[41757]_ ,
    \new_[41760]_ , \new_[41763]_ , \new_[41764]_ , \new_[41767]_ ,
    \new_[41770]_ , \new_[41771]_ , \new_[41772]_ , \new_[41776]_ ,
    \new_[41777]_ , \new_[41780]_ , \new_[41783]_ , \new_[41784]_ ,
    \new_[41785]_ , \new_[41788]_ , \new_[41791]_ , \new_[41792]_ ,
    \new_[41795]_ , \new_[41798]_ , \new_[41799]_ , \new_[41800]_ ,
    \new_[41804]_ , \new_[41805]_ , \new_[41808]_ , \new_[41811]_ ,
    \new_[41812]_ , \new_[41813]_ , \new_[41816]_ , \new_[41819]_ ,
    \new_[41820]_ , \new_[41823]_ , \new_[41826]_ , \new_[41827]_ ,
    \new_[41828]_ , \new_[41832]_ , \new_[41833]_ , \new_[41836]_ ,
    \new_[41839]_ , \new_[41840]_ , \new_[41841]_ , \new_[41844]_ ,
    \new_[41847]_ , \new_[41848]_ , \new_[41851]_ , \new_[41854]_ ,
    \new_[41855]_ , \new_[41856]_ , \new_[41860]_ , \new_[41861]_ ,
    \new_[41864]_ , \new_[41867]_ , \new_[41868]_ , \new_[41869]_ ,
    \new_[41872]_ , \new_[41875]_ , \new_[41876]_ , \new_[41879]_ ,
    \new_[41882]_ , \new_[41883]_ , \new_[41884]_ , \new_[41888]_ ,
    \new_[41889]_ , \new_[41892]_ , \new_[41895]_ , \new_[41896]_ ,
    \new_[41897]_ , \new_[41900]_ , \new_[41903]_ , \new_[41904]_ ,
    \new_[41907]_ , \new_[41910]_ , \new_[41911]_ , \new_[41912]_ ,
    \new_[41916]_ , \new_[41917]_ , \new_[41920]_ , \new_[41923]_ ,
    \new_[41924]_ , \new_[41925]_ , \new_[41928]_ , \new_[41931]_ ,
    \new_[41932]_ , \new_[41935]_ , \new_[41938]_ , \new_[41939]_ ,
    \new_[41940]_ , \new_[41944]_ , \new_[41945]_ , \new_[41948]_ ,
    \new_[41951]_ , \new_[41952]_ , \new_[41953]_ , \new_[41956]_ ,
    \new_[41959]_ , \new_[41960]_ , \new_[41963]_ , \new_[41966]_ ,
    \new_[41967]_ , \new_[41968]_ , \new_[41972]_ , \new_[41973]_ ,
    \new_[41976]_ , \new_[41979]_ , \new_[41980]_ , \new_[41981]_ ,
    \new_[41984]_ , \new_[41987]_ , \new_[41988]_ , \new_[41991]_ ,
    \new_[41994]_ , \new_[41995]_ , \new_[41996]_ , \new_[42000]_ ,
    \new_[42001]_ , \new_[42004]_ , \new_[42007]_ , \new_[42008]_ ,
    \new_[42009]_ , \new_[42012]_ , \new_[42015]_ , \new_[42016]_ ,
    \new_[42019]_ , \new_[42022]_ , \new_[42023]_ , \new_[42024]_ ,
    \new_[42028]_ , \new_[42029]_ , \new_[42032]_ , \new_[42035]_ ,
    \new_[42036]_ , \new_[42037]_ , \new_[42040]_ , \new_[42043]_ ,
    \new_[42044]_ , \new_[42047]_ , \new_[42050]_ , \new_[42051]_ ,
    \new_[42052]_ , \new_[42056]_ , \new_[42057]_ , \new_[42060]_ ,
    \new_[42063]_ , \new_[42064]_ , \new_[42065]_ , \new_[42068]_ ,
    \new_[42071]_ , \new_[42072]_ , \new_[42075]_ , \new_[42078]_ ,
    \new_[42079]_ , \new_[42080]_ , \new_[42084]_ , \new_[42085]_ ,
    \new_[42088]_ , \new_[42091]_ , \new_[42092]_ , \new_[42093]_ ,
    \new_[42096]_ , \new_[42099]_ , \new_[42100]_ , \new_[42103]_ ,
    \new_[42106]_ , \new_[42107]_ , \new_[42108]_ , \new_[42112]_ ,
    \new_[42113]_ , \new_[42116]_ , \new_[42119]_ , \new_[42120]_ ,
    \new_[42121]_ , \new_[42124]_ , \new_[42127]_ , \new_[42128]_ ,
    \new_[42131]_ , \new_[42134]_ , \new_[42135]_ , \new_[42136]_ ,
    \new_[42140]_ , \new_[42141]_ , \new_[42144]_ , \new_[42147]_ ,
    \new_[42148]_ , \new_[42149]_ , \new_[42152]_ , \new_[42155]_ ,
    \new_[42156]_ , \new_[42159]_ , \new_[42162]_ , \new_[42163]_ ,
    \new_[42164]_ , \new_[42168]_ , \new_[42169]_ , \new_[42172]_ ,
    \new_[42175]_ , \new_[42176]_ , \new_[42177]_ , \new_[42180]_ ,
    \new_[42183]_ , \new_[42184]_ , \new_[42187]_ , \new_[42190]_ ,
    \new_[42191]_ , \new_[42192]_ , \new_[42196]_ , \new_[42197]_ ,
    \new_[42200]_ , \new_[42203]_ , \new_[42204]_ , \new_[42205]_ ,
    \new_[42208]_ , \new_[42211]_ , \new_[42212]_ , \new_[42215]_ ,
    \new_[42218]_ , \new_[42219]_ , \new_[42220]_ , \new_[42224]_ ,
    \new_[42225]_ , \new_[42228]_ , \new_[42231]_ , \new_[42232]_ ,
    \new_[42233]_ , \new_[42236]_ , \new_[42239]_ , \new_[42240]_ ,
    \new_[42243]_ , \new_[42246]_ , \new_[42247]_ , \new_[42248]_ ,
    \new_[42252]_ , \new_[42253]_ , \new_[42256]_ , \new_[42259]_ ,
    \new_[42260]_ , \new_[42261]_ , \new_[42264]_ , \new_[42267]_ ,
    \new_[42268]_ , \new_[42271]_ , \new_[42274]_ , \new_[42275]_ ,
    \new_[42276]_ , \new_[42280]_ , \new_[42281]_ , \new_[42284]_ ,
    \new_[42287]_ , \new_[42288]_ , \new_[42289]_ , \new_[42292]_ ,
    \new_[42295]_ , \new_[42296]_ , \new_[42299]_ , \new_[42302]_ ,
    \new_[42303]_ , \new_[42304]_ , \new_[42308]_ , \new_[42309]_ ,
    \new_[42312]_ , \new_[42315]_ , \new_[42316]_ , \new_[42317]_ ,
    \new_[42320]_ , \new_[42323]_ , \new_[42324]_ , \new_[42327]_ ,
    \new_[42330]_ , \new_[42331]_ , \new_[42332]_ , \new_[42336]_ ,
    \new_[42337]_ , \new_[42340]_ , \new_[42343]_ , \new_[42344]_ ,
    \new_[42345]_ , \new_[42348]_ , \new_[42351]_ , \new_[42352]_ ,
    \new_[42355]_ , \new_[42358]_ , \new_[42359]_ , \new_[42360]_ ,
    \new_[42364]_ , \new_[42365]_ , \new_[42368]_ , \new_[42371]_ ,
    \new_[42372]_ , \new_[42373]_ , \new_[42376]_ , \new_[42379]_ ,
    \new_[42380]_ , \new_[42383]_ , \new_[42386]_ , \new_[42387]_ ,
    \new_[42388]_ , \new_[42392]_ , \new_[42393]_ , \new_[42396]_ ,
    \new_[42399]_ , \new_[42400]_ , \new_[42401]_ , \new_[42404]_ ,
    \new_[42407]_ , \new_[42408]_ , \new_[42411]_ , \new_[42414]_ ,
    \new_[42415]_ , \new_[42416]_ , \new_[42420]_ , \new_[42421]_ ,
    \new_[42424]_ , \new_[42427]_ , \new_[42428]_ , \new_[42429]_ ,
    \new_[42432]_ , \new_[42435]_ , \new_[42436]_ , \new_[42439]_ ,
    \new_[42442]_ , \new_[42443]_ , \new_[42444]_ , \new_[42448]_ ,
    \new_[42449]_ , \new_[42452]_ , \new_[42455]_ , \new_[42456]_ ,
    \new_[42457]_ , \new_[42460]_ , \new_[42463]_ , \new_[42464]_ ,
    \new_[42467]_ , \new_[42470]_ , \new_[42471]_ , \new_[42472]_ ,
    \new_[42476]_ , \new_[42477]_ , \new_[42480]_ , \new_[42483]_ ,
    \new_[42484]_ , \new_[42485]_ , \new_[42488]_ , \new_[42491]_ ,
    \new_[42492]_ , \new_[42495]_ , \new_[42498]_ , \new_[42499]_ ,
    \new_[42500]_ , \new_[42504]_ , \new_[42505]_ , \new_[42508]_ ,
    \new_[42511]_ , \new_[42512]_ , \new_[42513]_ , \new_[42516]_ ,
    \new_[42519]_ , \new_[42520]_ , \new_[42523]_ , \new_[42526]_ ,
    \new_[42527]_ , \new_[42528]_ , \new_[42532]_ , \new_[42533]_ ,
    \new_[42536]_ , \new_[42539]_ , \new_[42540]_ , \new_[42541]_ ,
    \new_[42544]_ , \new_[42547]_ , \new_[42548]_ , \new_[42551]_ ,
    \new_[42554]_ , \new_[42555]_ , \new_[42556]_ , \new_[42560]_ ,
    \new_[42561]_ , \new_[42564]_ , \new_[42567]_ , \new_[42568]_ ,
    \new_[42569]_ , \new_[42572]_ , \new_[42575]_ , \new_[42576]_ ,
    \new_[42579]_ , \new_[42582]_ , \new_[42583]_ , \new_[42584]_ ,
    \new_[42588]_ , \new_[42589]_ , \new_[42592]_ , \new_[42595]_ ,
    \new_[42596]_ , \new_[42597]_ , \new_[42600]_ , \new_[42603]_ ,
    \new_[42604]_ , \new_[42607]_ , \new_[42610]_ , \new_[42611]_ ,
    \new_[42612]_ , \new_[42616]_ , \new_[42617]_ , \new_[42620]_ ,
    \new_[42623]_ , \new_[42624]_ , \new_[42625]_ , \new_[42628]_ ,
    \new_[42631]_ , \new_[42632]_ , \new_[42635]_ , \new_[42638]_ ,
    \new_[42639]_ , \new_[42640]_ , \new_[42644]_ , \new_[42645]_ ,
    \new_[42648]_ , \new_[42651]_ , \new_[42652]_ , \new_[42653]_ ,
    \new_[42656]_ , \new_[42659]_ , \new_[42660]_ , \new_[42663]_ ,
    \new_[42666]_ , \new_[42667]_ , \new_[42668]_ , \new_[42672]_ ,
    \new_[42673]_ , \new_[42676]_ , \new_[42679]_ , \new_[42680]_ ,
    \new_[42681]_ , \new_[42684]_ , \new_[42687]_ , \new_[42688]_ ,
    \new_[42691]_ , \new_[42694]_ , \new_[42695]_ , \new_[42696]_ ,
    \new_[42700]_ , \new_[42701]_ , \new_[42704]_ , \new_[42707]_ ,
    \new_[42708]_ , \new_[42709]_ , \new_[42712]_ , \new_[42715]_ ,
    \new_[42716]_ , \new_[42719]_ , \new_[42722]_ , \new_[42723]_ ,
    \new_[42724]_ , \new_[42728]_ , \new_[42729]_ , \new_[42732]_ ,
    \new_[42735]_ , \new_[42736]_ , \new_[42737]_ , \new_[42740]_ ,
    \new_[42743]_ , \new_[42744]_ , \new_[42747]_ , \new_[42750]_ ,
    \new_[42751]_ , \new_[42752]_ , \new_[42756]_ , \new_[42757]_ ,
    \new_[42760]_ , \new_[42763]_ , \new_[42764]_ , \new_[42765]_ ,
    \new_[42768]_ , \new_[42771]_ , \new_[42772]_ , \new_[42775]_ ,
    \new_[42778]_ , \new_[42779]_ , \new_[42780]_ , \new_[42784]_ ,
    \new_[42785]_ , \new_[42788]_ , \new_[42791]_ , \new_[42792]_ ,
    \new_[42793]_ , \new_[42796]_ , \new_[42799]_ , \new_[42800]_ ,
    \new_[42803]_ , \new_[42806]_ , \new_[42807]_ , \new_[42808]_ ,
    \new_[42812]_ , \new_[42813]_ , \new_[42816]_ , \new_[42819]_ ,
    \new_[42820]_ , \new_[42821]_ , \new_[42824]_ , \new_[42827]_ ,
    \new_[42828]_ , \new_[42831]_ , \new_[42834]_ , \new_[42835]_ ,
    \new_[42836]_ , \new_[42840]_ , \new_[42841]_ , \new_[42844]_ ,
    \new_[42847]_ , \new_[42848]_ , \new_[42849]_ , \new_[42852]_ ,
    \new_[42855]_ , \new_[42856]_ , \new_[42859]_ , \new_[42862]_ ,
    \new_[42863]_ , \new_[42864]_ , \new_[42868]_ , \new_[42869]_ ,
    \new_[42872]_ , \new_[42875]_ , \new_[42876]_ , \new_[42877]_ ,
    \new_[42880]_ , \new_[42883]_ , \new_[42884]_ , \new_[42887]_ ,
    \new_[42890]_ , \new_[42891]_ , \new_[42892]_ , \new_[42896]_ ,
    \new_[42897]_ , \new_[42900]_ , \new_[42903]_ , \new_[42904]_ ,
    \new_[42905]_ , \new_[42908]_ , \new_[42911]_ , \new_[42912]_ ,
    \new_[42915]_ , \new_[42918]_ , \new_[42919]_ , \new_[42920]_ ,
    \new_[42924]_ , \new_[42925]_ , \new_[42928]_ , \new_[42931]_ ,
    \new_[42932]_ , \new_[42933]_ , \new_[42936]_ , \new_[42939]_ ,
    \new_[42940]_ , \new_[42943]_ , \new_[42946]_ , \new_[42947]_ ,
    \new_[42948]_ , \new_[42952]_ , \new_[42953]_ , \new_[42956]_ ,
    \new_[42959]_ , \new_[42960]_ , \new_[42961]_ , \new_[42964]_ ,
    \new_[42967]_ , \new_[42968]_ , \new_[42971]_ , \new_[42974]_ ,
    \new_[42975]_ , \new_[42976]_ , \new_[42980]_ , \new_[42981]_ ,
    \new_[42984]_ , \new_[42987]_ , \new_[42988]_ , \new_[42989]_ ,
    \new_[42992]_ , \new_[42995]_ , \new_[42996]_ , \new_[42999]_ ,
    \new_[43002]_ , \new_[43003]_ , \new_[43004]_ , \new_[43008]_ ,
    \new_[43009]_ , \new_[43012]_ , \new_[43015]_ , \new_[43016]_ ,
    \new_[43017]_ , \new_[43020]_ , \new_[43023]_ , \new_[43024]_ ,
    \new_[43027]_ , \new_[43030]_ , \new_[43031]_ , \new_[43032]_ ,
    \new_[43036]_ , \new_[43037]_ , \new_[43040]_ , \new_[43043]_ ,
    \new_[43044]_ , \new_[43045]_ , \new_[43048]_ , \new_[43051]_ ,
    \new_[43052]_ , \new_[43055]_ , \new_[43058]_ , \new_[43059]_ ,
    \new_[43060]_ , \new_[43064]_ , \new_[43065]_ , \new_[43068]_ ,
    \new_[43071]_ , \new_[43072]_ , \new_[43073]_ , \new_[43076]_ ,
    \new_[43079]_ , \new_[43080]_ , \new_[43083]_ , \new_[43086]_ ,
    \new_[43087]_ , \new_[43088]_ , \new_[43092]_ , \new_[43093]_ ,
    \new_[43096]_ , \new_[43099]_ , \new_[43100]_ , \new_[43101]_ ,
    \new_[43104]_ , \new_[43107]_ , \new_[43108]_ , \new_[43111]_ ,
    \new_[43114]_ , \new_[43115]_ , \new_[43116]_ , \new_[43120]_ ,
    \new_[43121]_ , \new_[43124]_ , \new_[43127]_ , \new_[43128]_ ,
    \new_[43129]_ , \new_[43132]_ , \new_[43135]_ , \new_[43136]_ ,
    \new_[43139]_ , \new_[43142]_ , \new_[43143]_ , \new_[43144]_ ,
    \new_[43148]_ , \new_[43149]_ , \new_[43152]_ , \new_[43155]_ ,
    \new_[43156]_ , \new_[43157]_ , \new_[43160]_ , \new_[43163]_ ,
    \new_[43164]_ , \new_[43167]_ , \new_[43170]_ , \new_[43171]_ ,
    \new_[43172]_ , \new_[43176]_ , \new_[43177]_ , \new_[43180]_ ,
    \new_[43183]_ , \new_[43184]_ , \new_[43185]_ , \new_[43188]_ ,
    \new_[43191]_ , \new_[43192]_ , \new_[43195]_ , \new_[43198]_ ,
    \new_[43199]_ , \new_[43200]_ , \new_[43204]_ , \new_[43205]_ ,
    \new_[43208]_ , \new_[43211]_ , \new_[43212]_ , \new_[43213]_ ,
    \new_[43216]_ , \new_[43219]_ , \new_[43220]_ , \new_[43223]_ ,
    \new_[43226]_ , \new_[43227]_ , \new_[43228]_ , \new_[43232]_ ,
    \new_[43233]_ , \new_[43236]_ , \new_[43239]_ , \new_[43240]_ ,
    \new_[43241]_ , \new_[43244]_ , \new_[43247]_ , \new_[43248]_ ,
    \new_[43251]_ , \new_[43254]_ , \new_[43255]_ , \new_[43256]_ ,
    \new_[43260]_ , \new_[43261]_ , \new_[43264]_ , \new_[43267]_ ,
    \new_[43268]_ , \new_[43269]_ , \new_[43272]_ , \new_[43275]_ ,
    \new_[43276]_ , \new_[43279]_ , \new_[43282]_ , \new_[43283]_ ,
    \new_[43284]_ , \new_[43288]_ , \new_[43289]_ , \new_[43292]_ ,
    \new_[43295]_ , \new_[43296]_ , \new_[43297]_ , \new_[43300]_ ,
    \new_[43303]_ , \new_[43304]_ , \new_[43307]_ , \new_[43310]_ ,
    \new_[43311]_ , \new_[43312]_ , \new_[43316]_ , \new_[43317]_ ,
    \new_[43320]_ , \new_[43323]_ , \new_[43324]_ , \new_[43325]_ ,
    \new_[43328]_ , \new_[43331]_ , \new_[43332]_ , \new_[43335]_ ,
    \new_[43338]_ , \new_[43339]_ , \new_[43340]_ , \new_[43344]_ ,
    \new_[43345]_ , \new_[43348]_ , \new_[43351]_ , \new_[43352]_ ,
    \new_[43353]_ , \new_[43356]_ , \new_[43359]_ , \new_[43360]_ ,
    \new_[43363]_ , \new_[43366]_ , \new_[43367]_ , \new_[43368]_ ,
    \new_[43372]_ , \new_[43373]_ , \new_[43376]_ , \new_[43379]_ ,
    \new_[43380]_ , \new_[43381]_ , \new_[43384]_ , \new_[43387]_ ,
    \new_[43388]_ , \new_[43391]_ , \new_[43394]_ , \new_[43395]_ ,
    \new_[43396]_ , \new_[43400]_ , \new_[43401]_ , \new_[43404]_ ,
    \new_[43407]_ , \new_[43408]_ , \new_[43409]_ , \new_[43412]_ ,
    \new_[43415]_ , \new_[43416]_ , \new_[43419]_ , \new_[43422]_ ,
    \new_[43423]_ , \new_[43424]_ , \new_[43428]_ , \new_[43429]_ ,
    \new_[43432]_ , \new_[43435]_ , \new_[43436]_ , \new_[43437]_ ,
    \new_[43440]_ , \new_[43443]_ , \new_[43444]_ , \new_[43447]_ ,
    \new_[43450]_ , \new_[43451]_ , \new_[43452]_ , \new_[43456]_ ,
    \new_[43457]_ , \new_[43460]_ , \new_[43463]_ , \new_[43464]_ ,
    \new_[43465]_ , \new_[43468]_ , \new_[43471]_ , \new_[43472]_ ,
    \new_[43475]_ , \new_[43478]_ , \new_[43479]_ , \new_[43480]_ ,
    \new_[43484]_ , \new_[43485]_ , \new_[43488]_ , \new_[43491]_ ,
    \new_[43492]_ , \new_[43493]_ , \new_[43496]_ , \new_[43499]_ ,
    \new_[43500]_ , \new_[43503]_ , \new_[43506]_ , \new_[43507]_ ,
    \new_[43508]_ , \new_[43512]_ , \new_[43513]_ , \new_[43516]_ ,
    \new_[43519]_ , \new_[43520]_ , \new_[43521]_ , \new_[43524]_ ,
    \new_[43527]_ , \new_[43528]_ , \new_[43531]_ , \new_[43534]_ ,
    \new_[43535]_ , \new_[43536]_ , \new_[43540]_ , \new_[43541]_ ,
    \new_[43544]_ , \new_[43547]_ , \new_[43548]_ , \new_[43549]_ ,
    \new_[43552]_ , \new_[43555]_ , \new_[43556]_ , \new_[43559]_ ,
    \new_[43562]_ , \new_[43563]_ , \new_[43564]_ , \new_[43568]_ ,
    \new_[43569]_ , \new_[43572]_ , \new_[43575]_ , \new_[43576]_ ,
    \new_[43577]_ , \new_[43580]_ , \new_[43583]_ , \new_[43584]_ ,
    \new_[43587]_ , \new_[43590]_ , \new_[43591]_ , \new_[43592]_ ,
    \new_[43596]_ , \new_[43597]_ , \new_[43600]_ , \new_[43603]_ ,
    \new_[43604]_ , \new_[43605]_ , \new_[43608]_ , \new_[43611]_ ,
    \new_[43612]_ , \new_[43615]_ , \new_[43618]_ , \new_[43619]_ ,
    \new_[43620]_ , \new_[43624]_ , \new_[43625]_ , \new_[43628]_ ,
    \new_[43631]_ , \new_[43632]_ , \new_[43633]_ , \new_[43636]_ ,
    \new_[43639]_ , \new_[43640]_ , \new_[43643]_ , \new_[43646]_ ,
    \new_[43647]_ , \new_[43648]_ , \new_[43652]_ , \new_[43653]_ ,
    \new_[43656]_ , \new_[43659]_ , \new_[43660]_ , \new_[43661]_ ,
    \new_[43664]_ , \new_[43667]_ , \new_[43668]_ , \new_[43671]_ ,
    \new_[43674]_ , \new_[43675]_ , \new_[43676]_ , \new_[43680]_ ,
    \new_[43681]_ , \new_[43684]_ , \new_[43687]_ , \new_[43688]_ ,
    \new_[43689]_ , \new_[43692]_ , \new_[43695]_ , \new_[43696]_ ,
    \new_[43699]_ , \new_[43702]_ , \new_[43703]_ , \new_[43704]_ ,
    \new_[43708]_ , \new_[43709]_ , \new_[43712]_ , \new_[43715]_ ,
    \new_[43716]_ , \new_[43717]_ , \new_[43720]_ , \new_[43723]_ ,
    \new_[43724]_ , \new_[43727]_ , \new_[43730]_ , \new_[43731]_ ,
    \new_[43732]_ , \new_[43736]_ , \new_[43737]_ , \new_[43740]_ ,
    \new_[43743]_ , \new_[43744]_ , \new_[43745]_ , \new_[43748]_ ,
    \new_[43751]_ , \new_[43752]_ , \new_[43755]_ , \new_[43758]_ ,
    \new_[43759]_ , \new_[43760]_ , \new_[43764]_ , \new_[43765]_ ,
    \new_[43768]_ , \new_[43771]_ , \new_[43772]_ , \new_[43773]_ ,
    \new_[43776]_ , \new_[43779]_ , \new_[43780]_ , \new_[43783]_ ,
    \new_[43786]_ , \new_[43787]_ , \new_[43788]_ , \new_[43792]_ ,
    \new_[43793]_ , \new_[43796]_ , \new_[43799]_ , \new_[43800]_ ,
    \new_[43801]_ , \new_[43804]_ , \new_[43807]_ , \new_[43808]_ ,
    \new_[43811]_ , \new_[43814]_ , \new_[43815]_ , \new_[43816]_ ,
    \new_[43820]_ , \new_[43821]_ , \new_[43824]_ , \new_[43827]_ ,
    \new_[43828]_ , \new_[43829]_ , \new_[43832]_ , \new_[43835]_ ,
    \new_[43836]_ , \new_[43839]_ , \new_[43842]_ , \new_[43843]_ ,
    \new_[43844]_ , \new_[43848]_ , \new_[43849]_ , \new_[43852]_ ,
    \new_[43855]_ , \new_[43856]_ , \new_[43857]_ , \new_[43860]_ ,
    \new_[43863]_ , \new_[43864]_ , \new_[43867]_ , \new_[43870]_ ,
    \new_[43871]_ , \new_[43872]_ , \new_[43876]_ , \new_[43877]_ ,
    \new_[43880]_ , \new_[43883]_ , \new_[43884]_ , \new_[43885]_ ,
    \new_[43888]_ , \new_[43891]_ , \new_[43892]_ , \new_[43895]_ ,
    \new_[43898]_ , \new_[43899]_ , \new_[43900]_ , \new_[43904]_ ,
    \new_[43905]_ , \new_[43908]_ , \new_[43911]_ , \new_[43912]_ ,
    \new_[43913]_ , \new_[43916]_ , \new_[43919]_ , \new_[43920]_ ,
    \new_[43923]_ , \new_[43926]_ , \new_[43927]_ , \new_[43928]_ ,
    \new_[43932]_ , \new_[43933]_ , \new_[43936]_ , \new_[43939]_ ,
    \new_[43940]_ , \new_[43941]_ , \new_[43944]_ , \new_[43947]_ ,
    \new_[43948]_ , \new_[43951]_ , \new_[43954]_ , \new_[43955]_ ,
    \new_[43956]_ , \new_[43960]_ , \new_[43961]_ , \new_[43964]_ ,
    \new_[43967]_ , \new_[43968]_ , \new_[43969]_ , \new_[43972]_ ,
    \new_[43975]_ , \new_[43976]_ , \new_[43979]_ , \new_[43982]_ ,
    \new_[43983]_ , \new_[43984]_ , \new_[43988]_ , \new_[43989]_ ,
    \new_[43992]_ , \new_[43995]_ , \new_[43996]_ , \new_[43997]_ ,
    \new_[44000]_ , \new_[44003]_ , \new_[44004]_ , \new_[44007]_ ,
    \new_[44010]_ , \new_[44011]_ , \new_[44012]_ , \new_[44016]_ ,
    \new_[44017]_ , \new_[44020]_ , \new_[44023]_ , \new_[44024]_ ,
    \new_[44025]_ , \new_[44028]_ , \new_[44031]_ , \new_[44032]_ ,
    \new_[44035]_ , \new_[44038]_ , \new_[44039]_ , \new_[44040]_ ,
    \new_[44044]_ , \new_[44045]_ , \new_[44048]_ , \new_[44051]_ ,
    \new_[44052]_ , \new_[44053]_ , \new_[44056]_ , \new_[44059]_ ,
    \new_[44060]_ , \new_[44063]_ , \new_[44066]_ , \new_[44067]_ ,
    \new_[44068]_ , \new_[44072]_ , \new_[44073]_ , \new_[44076]_ ,
    \new_[44079]_ , \new_[44080]_ , \new_[44081]_ , \new_[44084]_ ,
    \new_[44087]_ , \new_[44088]_ , \new_[44091]_ , \new_[44094]_ ,
    \new_[44095]_ , \new_[44096]_ , \new_[44100]_ , \new_[44101]_ ,
    \new_[44104]_ , \new_[44107]_ , \new_[44108]_ , \new_[44109]_ ,
    \new_[44112]_ , \new_[44115]_ , \new_[44116]_ , \new_[44119]_ ,
    \new_[44122]_ , \new_[44123]_ , \new_[44124]_ , \new_[44128]_ ,
    \new_[44129]_ , \new_[44132]_ , \new_[44135]_ , \new_[44136]_ ,
    \new_[44137]_ , \new_[44140]_ , \new_[44143]_ , \new_[44144]_ ,
    \new_[44147]_ , \new_[44150]_ , \new_[44151]_ , \new_[44152]_ ,
    \new_[44156]_ , \new_[44157]_ , \new_[44160]_ , \new_[44163]_ ,
    \new_[44164]_ , \new_[44165]_ , \new_[44168]_ , \new_[44171]_ ,
    \new_[44172]_ , \new_[44175]_ , \new_[44178]_ , \new_[44179]_ ,
    \new_[44180]_ , \new_[44184]_ , \new_[44185]_ , \new_[44188]_ ,
    \new_[44191]_ , \new_[44192]_ , \new_[44193]_ , \new_[44196]_ ,
    \new_[44199]_ , \new_[44200]_ , \new_[44203]_ , \new_[44206]_ ,
    \new_[44207]_ , \new_[44208]_ , \new_[44212]_ , \new_[44213]_ ,
    \new_[44216]_ , \new_[44219]_ , \new_[44220]_ , \new_[44221]_ ,
    \new_[44224]_ , \new_[44227]_ , \new_[44228]_ , \new_[44231]_ ,
    \new_[44234]_ , \new_[44235]_ , \new_[44236]_ , \new_[44240]_ ,
    \new_[44241]_ , \new_[44244]_ , \new_[44247]_ , \new_[44248]_ ,
    \new_[44249]_ , \new_[44252]_ , \new_[44255]_ , \new_[44256]_ ,
    \new_[44259]_ , \new_[44262]_ , \new_[44263]_ , \new_[44264]_ ,
    \new_[44268]_ , \new_[44269]_ , \new_[44272]_ , \new_[44275]_ ,
    \new_[44276]_ , \new_[44277]_ , \new_[44280]_ , \new_[44283]_ ,
    \new_[44284]_ , \new_[44287]_ , \new_[44290]_ , \new_[44291]_ ,
    \new_[44292]_ , \new_[44296]_ , \new_[44297]_ , \new_[44300]_ ,
    \new_[44303]_ , \new_[44304]_ , \new_[44305]_ , \new_[44308]_ ,
    \new_[44311]_ , \new_[44312]_ , \new_[44315]_ , \new_[44318]_ ,
    \new_[44319]_ , \new_[44320]_ , \new_[44324]_ , \new_[44325]_ ,
    \new_[44328]_ , \new_[44331]_ , \new_[44332]_ , \new_[44333]_ ,
    \new_[44336]_ , \new_[44339]_ , \new_[44340]_ , \new_[44343]_ ,
    \new_[44346]_ , \new_[44347]_ , \new_[44348]_ , \new_[44352]_ ,
    \new_[44353]_ , \new_[44356]_ , \new_[44359]_ , \new_[44360]_ ,
    \new_[44361]_ , \new_[44364]_ , \new_[44367]_ , \new_[44368]_ ,
    \new_[44371]_ , \new_[44374]_ , \new_[44375]_ , \new_[44376]_ ,
    \new_[44380]_ , \new_[44381]_ , \new_[44384]_ , \new_[44387]_ ,
    \new_[44388]_ , \new_[44389]_ , \new_[44392]_ , \new_[44395]_ ,
    \new_[44396]_ , \new_[44399]_ , \new_[44402]_ , \new_[44403]_ ,
    \new_[44404]_ , \new_[44408]_ , \new_[44409]_ , \new_[44412]_ ,
    \new_[44415]_ , \new_[44416]_ , \new_[44417]_ , \new_[44420]_ ,
    \new_[44423]_ , \new_[44424]_ , \new_[44427]_ , \new_[44430]_ ,
    \new_[44431]_ , \new_[44432]_ , \new_[44436]_ , \new_[44437]_ ,
    \new_[44440]_ , \new_[44443]_ , \new_[44444]_ , \new_[44445]_ ,
    \new_[44448]_ , \new_[44451]_ , \new_[44452]_ , \new_[44455]_ ,
    \new_[44458]_ , \new_[44459]_ , \new_[44460]_ , \new_[44464]_ ,
    \new_[44465]_ , \new_[44468]_ , \new_[44471]_ , \new_[44472]_ ,
    \new_[44473]_ , \new_[44476]_ , \new_[44479]_ , \new_[44480]_ ,
    \new_[44483]_ , \new_[44486]_ , \new_[44487]_ , \new_[44488]_ ,
    \new_[44492]_ , \new_[44493]_ , \new_[44496]_ , \new_[44499]_ ,
    \new_[44500]_ , \new_[44501]_ , \new_[44504]_ , \new_[44507]_ ,
    \new_[44508]_ , \new_[44511]_ , \new_[44514]_ , \new_[44515]_ ,
    \new_[44516]_ , \new_[44520]_ , \new_[44521]_ , \new_[44524]_ ,
    \new_[44527]_ , \new_[44528]_ , \new_[44529]_ , \new_[44532]_ ,
    \new_[44535]_ , \new_[44536]_ , \new_[44539]_ , \new_[44542]_ ,
    \new_[44543]_ , \new_[44544]_ , \new_[44547]_ , \new_[44550]_ ,
    \new_[44551]_ , \new_[44554]_ , \new_[44557]_ , \new_[44558]_ ,
    \new_[44559]_ , \new_[44562]_ , \new_[44565]_ , \new_[44566]_ ,
    \new_[44569]_ , \new_[44572]_ , \new_[44573]_ , \new_[44574]_ ,
    \new_[44577]_ , \new_[44580]_ , \new_[44581]_ , \new_[44584]_ ,
    \new_[44587]_ , \new_[44588]_ , \new_[44589]_ , \new_[44592]_ ,
    \new_[44595]_ , \new_[44596]_ , \new_[44599]_ , \new_[44602]_ ,
    \new_[44603]_ , \new_[44604]_ , \new_[44607]_ , \new_[44610]_ ,
    \new_[44611]_ , \new_[44614]_ , \new_[44617]_ , \new_[44618]_ ,
    \new_[44619]_ , \new_[44622]_ , \new_[44625]_ , \new_[44626]_ ,
    \new_[44629]_ , \new_[44632]_ , \new_[44633]_ , \new_[44634]_ ,
    \new_[44637]_ , \new_[44640]_ , \new_[44641]_ , \new_[44644]_ ,
    \new_[44647]_ , \new_[44648]_ , \new_[44649]_ , \new_[44652]_ ,
    \new_[44655]_ , \new_[44656]_ , \new_[44659]_ , \new_[44662]_ ,
    \new_[44663]_ , \new_[44664]_ , \new_[44667]_ , \new_[44670]_ ,
    \new_[44671]_ , \new_[44674]_ , \new_[44677]_ , \new_[44678]_ ,
    \new_[44679]_ , \new_[44682]_ , \new_[44685]_ , \new_[44686]_ ,
    \new_[44689]_ , \new_[44692]_ , \new_[44693]_ , \new_[44694]_ ,
    \new_[44697]_ , \new_[44700]_ , \new_[44701]_ , \new_[44704]_ ,
    \new_[44707]_ , \new_[44708]_ , \new_[44709]_ , \new_[44712]_ ,
    \new_[44715]_ , \new_[44716]_ , \new_[44719]_ , \new_[44722]_ ,
    \new_[44723]_ , \new_[44724]_ , \new_[44727]_ , \new_[44730]_ ,
    \new_[44731]_ , \new_[44734]_ , \new_[44737]_ , \new_[44738]_ ,
    \new_[44739]_ , \new_[44742]_ , \new_[44745]_ , \new_[44746]_ ,
    \new_[44749]_ , \new_[44752]_ , \new_[44753]_ , \new_[44754]_ ,
    \new_[44757]_ , \new_[44760]_ , \new_[44761]_ , \new_[44764]_ ,
    \new_[44767]_ , \new_[44768]_ , \new_[44769]_ , \new_[44772]_ ,
    \new_[44775]_ , \new_[44776]_ , \new_[44779]_ , \new_[44782]_ ,
    \new_[44783]_ , \new_[44784]_ , \new_[44787]_ , \new_[44790]_ ,
    \new_[44791]_ , \new_[44794]_ , \new_[44797]_ , \new_[44798]_ ,
    \new_[44799]_ , \new_[44802]_ , \new_[44805]_ , \new_[44806]_ ,
    \new_[44809]_ , \new_[44812]_ , \new_[44813]_ , \new_[44814]_ ,
    \new_[44817]_ , \new_[44820]_ , \new_[44821]_ , \new_[44824]_ ,
    \new_[44827]_ , \new_[44828]_ , \new_[44829]_ , \new_[44832]_ ,
    \new_[44835]_ , \new_[44836]_ , \new_[44839]_ , \new_[44842]_ ,
    \new_[44843]_ , \new_[44844]_ , \new_[44847]_ , \new_[44850]_ ,
    \new_[44851]_ , \new_[44854]_ , \new_[44857]_ , \new_[44858]_ ,
    \new_[44859]_ , \new_[44862]_ , \new_[44865]_ , \new_[44866]_ ,
    \new_[44869]_ , \new_[44872]_ , \new_[44873]_ , \new_[44874]_ ,
    \new_[44877]_ , \new_[44880]_ , \new_[44881]_ , \new_[44884]_ ,
    \new_[44887]_ , \new_[44888]_ , \new_[44889]_ , \new_[44892]_ ,
    \new_[44895]_ , \new_[44896]_ , \new_[44899]_ , \new_[44902]_ ,
    \new_[44903]_ , \new_[44904]_ , \new_[44907]_ , \new_[44910]_ ,
    \new_[44911]_ , \new_[44914]_ , \new_[44917]_ , \new_[44918]_ ,
    \new_[44919]_ , \new_[44922]_ , \new_[44925]_ , \new_[44926]_ ,
    \new_[44929]_ , \new_[44932]_ , \new_[44933]_ , \new_[44934]_ ,
    \new_[44937]_ , \new_[44940]_ , \new_[44941]_ , \new_[44944]_ ,
    \new_[44947]_ , \new_[44948]_ , \new_[44949]_ , \new_[44952]_ ,
    \new_[44955]_ , \new_[44956]_ , \new_[44959]_ , \new_[44962]_ ,
    \new_[44963]_ , \new_[44964]_ , \new_[44967]_ , \new_[44970]_ ,
    \new_[44971]_ , \new_[44974]_ , \new_[44977]_ , \new_[44978]_ ,
    \new_[44979]_ , \new_[44982]_ , \new_[44985]_ , \new_[44986]_ ,
    \new_[44989]_ , \new_[44992]_ , \new_[44993]_ , \new_[44994]_ ,
    \new_[44997]_ , \new_[45000]_ , \new_[45001]_ , \new_[45004]_ ,
    \new_[45007]_ , \new_[45008]_ , \new_[45009]_ , \new_[45012]_ ,
    \new_[45015]_ , \new_[45016]_ , \new_[45019]_ , \new_[45022]_ ,
    \new_[45023]_ , \new_[45024]_ , \new_[45027]_ , \new_[45030]_ ,
    \new_[45031]_ , \new_[45034]_ , \new_[45037]_ , \new_[45038]_ ,
    \new_[45039]_ , \new_[45042]_ , \new_[45045]_ , \new_[45046]_ ,
    \new_[45049]_ , \new_[45052]_ , \new_[45053]_ , \new_[45054]_ ,
    \new_[45057]_ , \new_[45060]_ , \new_[45061]_ , \new_[45064]_ ,
    \new_[45067]_ , \new_[45068]_ , \new_[45069]_ , \new_[45072]_ ,
    \new_[45075]_ , \new_[45076]_ , \new_[45079]_ , \new_[45082]_ ,
    \new_[45083]_ , \new_[45084]_ , \new_[45087]_ , \new_[45090]_ ,
    \new_[45091]_ , \new_[45094]_ , \new_[45097]_ , \new_[45098]_ ,
    \new_[45099]_ , \new_[45102]_ , \new_[45105]_ , \new_[45106]_ ,
    \new_[45109]_ , \new_[45112]_ , \new_[45113]_ , \new_[45114]_ ,
    \new_[45117]_ , \new_[45120]_ , \new_[45121]_ , \new_[45124]_ ,
    \new_[45127]_ , \new_[45128]_ , \new_[45129]_ , \new_[45132]_ ,
    \new_[45135]_ , \new_[45136]_ , \new_[45139]_ , \new_[45142]_ ,
    \new_[45143]_ , \new_[45144]_ , \new_[45147]_ , \new_[45150]_ ,
    \new_[45151]_ , \new_[45154]_ , \new_[45157]_ , \new_[45158]_ ,
    \new_[45159]_ , \new_[45162]_ , \new_[45165]_ , \new_[45166]_ ,
    \new_[45169]_ , \new_[45172]_ , \new_[45173]_ , \new_[45174]_ ,
    \new_[45177]_ , \new_[45180]_ , \new_[45181]_ , \new_[45184]_ ,
    \new_[45187]_ , \new_[45188]_ , \new_[45189]_ , \new_[45192]_ ,
    \new_[45195]_ , \new_[45196]_ , \new_[45199]_ , \new_[45202]_ ,
    \new_[45203]_ , \new_[45204]_ , \new_[45207]_ , \new_[45210]_ ,
    \new_[45211]_ , \new_[45214]_ , \new_[45217]_ , \new_[45218]_ ,
    \new_[45219]_ , \new_[45222]_ , \new_[45225]_ , \new_[45226]_ ,
    \new_[45229]_ , \new_[45232]_ , \new_[45233]_ , \new_[45234]_ ,
    \new_[45237]_ , \new_[45240]_ , \new_[45241]_ , \new_[45244]_ ,
    \new_[45247]_ , \new_[45248]_ , \new_[45249]_ , \new_[45252]_ ,
    \new_[45255]_ , \new_[45256]_ , \new_[45259]_ , \new_[45262]_ ,
    \new_[45263]_ , \new_[45264]_ , \new_[45267]_ , \new_[45270]_ ,
    \new_[45271]_ , \new_[45274]_ , \new_[45277]_ , \new_[45278]_ ,
    \new_[45279]_ , \new_[45282]_ , \new_[45285]_ , \new_[45286]_ ,
    \new_[45289]_ , \new_[45292]_ , \new_[45293]_ , \new_[45294]_ ,
    \new_[45297]_ , \new_[45300]_ , \new_[45301]_ , \new_[45304]_ ,
    \new_[45307]_ , \new_[45308]_ , \new_[45309]_ , \new_[45312]_ ,
    \new_[45315]_ , \new_[45316]_ , \new_[45319]_ , \new_[45322]_ ,
    \new_[45323]_ , \new_[45324]_ , \new_[45327]_ , \new_[45330]_ ,
    \new_[45331]_ , \new_[45334]_ , \new_[45337]_ , \new_[45338]_ ,
    \new_[45339]_ , \new_[45342]_ , \new_[45345]_ , \new_[45346]_ ,
    \new_[45349]_ , \new_[45352]_ , \new_[45353]_ , \new_[45354]_ ,
    \new_[45357]_ , \new_[45360]_ , \new_[45361]_ , \new_[45364]_ ,
    \new_[45367]_ , \new_[45368]_ , \new_[45369]_ , \new_[45372]_ ,
    \new_[45375]_ , \new_[45376]_ , \new_[45379]_ , \new_[45382]_ ,
    \new_[45383]_ , \new_[45384]_ , \new_[45387]_ , \new_[45390]_ ,
    \new_[45391]_ , \new_[45394]_ , \new_[45397]_ , \new_[45398]_ ,
    \new_[45399]_ , \new_[45402]_ , \new_[45405]_ , \new_[45406]_ ,
    \new_[45409]_ , \new_[45412]_ , \new_[45413]_ , \new_[45414]_ ,
    \new_[45417]_ , \new_[45420]_ , \new_[45421]_ , \new_[45424]_ ,
    \new_[45427]_ , \new_[45428]_ , \new_[45429]_ , \new_[45432]_ ,
    \new_[45435]_ , \new_[45436]_ , \new_[45439]_ , \new_[45442]_ ,
    \new_[45443]_ , \new_[45444]_ , \new_[45447]_ , \new_[45450]_ ,
    \new_[45451]_ , \new_[45454]_ , \new_[45457]_ , \new_[45458]_ ,
    \new_[45459]_ , \new_[45462]_ , \new_[45465]_ , \new_[45466]_ ,
    \new_[45469]_ , \new_[45472]_ , \new_[45473]_ , \new_[45474]_ ,
    \new_[45477]_ , \new_[45480]_ , \new_[45481]_ , \new_[45484]_ ,
    \new_[45487]_ , \new_[45488]_ , \new_[45489]_ , \new_[45492]_ ,
    \new_[45495]_ , \new_[45496]_ , \new_[45499]_ , \new_[45502]_ ,
    \new_[45503]_ , \new_[45504]_ , \new_[45507]_ , \new_[45510]_ ,
    \new_[45511]_ , \new_[45514]_ , \new_[45517]_ , \new_[45518]_ ,
    \new_[45519]_ , \new_[45522]_ , \new_[45525]_ , \new_[45526]_ ,
    \new_[45529]_ , \new_[45532]_ , \new_[45533]_ , \new_[45534]_ ,
    \new_[45537]_ , \new_[45540]_ , \new_[45541]_ , \new_[45544]_ ,
    \new_[45547]_ , \new_[45548]_ , \new_[45549]_ , \new_[45552]_ ,
    \new_[45555]_ , \new_[45556]_ , \new_[45559]_ , \new_[45562]_ ,
    \new_[45563]_ , \new_[45564]_ , \new_[45567]_ , \new_[45570]_ ,
    \new_[45571]_ , \new_[45574]_ , \new_[45577]_ , \new_[45578]_ ,
    \new_[45579]_ , \new_[45582]_ , \new_[45585]_ , \new_[45586]_ ,
    \new_[45589]_ , \new_[45592]_ , \new_[45593]_ , \new_[45594]_ ,
    \new_[45597]_ , \new_[45600]_ , \new_[45601]_ , \new_[45604]_ ,
    \new_[45607]_ , \new_[45608]_ , \new_[45609]_ , \new_[45612]_ ,
    \new_[45615]_ , \new_[45616]_ , \new_[45619]_ , \new_[45622]_ ,
    \new_[45623]_ , \new_[45624]_ , \new_[45627]_ , \new_[45630]_ ,
    \new_[45631]_ , \new_[45634]_ , \new_[45637]_ , \new_[45638]_ ,
    \new_[45639]_ , \new_[45642]_ , \new_[45645]_ , \new_[45646]_ ,
    \new_[45649]_ , \new_[45652]_ , \new_[45653]_ , \new_[45654]_ ,
    \new_[45657]_ , \new_[45660]_ , \new_[45661]_ , \new_[45664]_ ,
    \new_[45667]_ , \new_[45668]_ , \new_[45669]_ , \new_[45672]_ ,
    \new_[45675]_ , \new_[45676]_ , \new_[45679]_ , \new_[45682]_ ,
    \new_[45683]_ , \new_[45684]_ , \new_[45687]_ , \new_[45690]_ ,
    \new_[45691]_ , \new_[45694]_ , \new_[45697]_ , \new_[45698]_ ,
    \new_[45699]_ , \new_[45702]_ , \new_[45705]_ , \new_[45706]_ ,
    \new_[45709]_ , \new_[45712]_ , \new_[45713]_ , \new_[45714]_ ,
    \new_[45717]_ , \new_[45720]_ , \new_[45721]_ , \new_[45724]_ ,
    \new_[45727]_ , \new_[45728]_ , \new_[45729]_ , \new_[45732]_ ,
    \new_[45735]_ , \new_[45736]_ , \new_[45739]_ , \new_[45742]_ ,
    \new_[45743]_ , \new_[45744]_ , \new_[45747]_ , \new_[45750]_ ,
    \new_[45751]_ , \new_[45754]_ , \new_[45757]_ , \new_[45758]_ ,
    \new_[45759]_ , \new_[45762]_ , \new_[45765]_ , \new_[45766]_ ,
    \new_[45769]_ , \new_[45772]_ , \new_[45773]_ , \new_[45774]_ ,
    \new_[45777]_ , \new_[45780]_ , \new_[45781]_ , \new_[45784]_ ,
    \new_[45787]_ , \new_[45788]_ , \new_[45789]_ , \new_[45792]_ ,
    \new_[45795]_ , \new_[45796]_ , \new_[45799]_ , \new_[45802]_ ,
    \new_[45803]_ , \new_[45804]_ , \new_[45807]_ , \new_[45810]_ ,
    \new_[45811]_ , \new_[45814]_ , \new_[45817]_ , \new_[45818]_ ,
    \new_[45819]_ , \new_[45822]_ , \new_[45825]_ , \new_[45826]_ ,
    \new_[45829]_ , \new_[45832]_ , \new_[45833]_ , \new_[45834]_ ,
    \new_[45837]_ , \new_[45840]_ , \new_[45841]_ , \new_[45844]_ ,
    \new_[45847]_ , \new_[45848]_ , \new_[45849]_ , \new_[45852]_ ,
    \new_[45855]_ , \new_[45856]_ , \new_[45859]_ , \new_[45862]_ ,
    \new_[45863]_ , \new_[45864]_ , \new_[45867]_ , \new_[45870]_ ,
    \new_[45871]_ , \new_[45874]_ , \new_[45877]_ , \new_[45878]_ ,
    \new_[45879]_ , \new_[45882]_ , \new_[45885]_ , \new_[45886]_ ,
    \new_[45889]_ , \new_[45892]_ , \new_[45893]_ , \new_[45894]_ ,
    \new_[45897]_ , \new_[45900]_ , \new_[45901]_ , \new_[45904]_ ,
    \new_[45907]_ , \new_[45908]_ , \new_[45909]_ , \new_[45912]_ ,
    \new_[45915]_ , \new_[45916]_ , \new_[45919]_ , \new_[45922]_ ,
    \new_[45923]_ , \new_[45924]_ , \new_[45927]_ , \new_[45930]_ ,
    \new_[45931]_ , \new_[45934]_ , \new_[45937]_ , \new_[45938]_ ,
    \new_[45939]_ , \new_[45942]_ , \new_[45945]_ , \new_[45946]_ ,
    \new_[45949]_ , \new_[45952]_ , \new_[45953]_ , \new_[45954]_ ,
    \new_[45957]_ , \new_[45960]_ , \new_[45961]_ , \new_[45964]_ ,
    \new_[45967]_ , \new_[45968]_ , \new_[45969]_ , \new_[45972]_ ,
    \new_[45975]_ , \new_[45976]_ , \new_[45979]_ , \new_[45982]_ ,
    \new_[45983]_ , \new_[45984]_ , \new_[45987]_ , \new_[45990]_ ,
    \new_[45991]_ , \new_[45994]_ , \new_[45997]_ , \new_[45998]_ ,
    \new_[45999]_ , \new_[46002]_ , \new_[46005]_ , \new_[46006]_ ,
    \new_[46009]_ , \new_[46012]_ , \new_[46013]_ , \new_[46014]_ ,
    \new_[46017]_ , \new_[46020]_ , \new_[46021]_ , \new_[46024]_ ,
    \new_[46027]_ , \new_[46028]_ , \new_[46029]_ , \new_[46032]_ ,
    \new_[46035]_ , \new_[46036]_ , \new_[46039]_ , \new_[46042]_ ,
    \new_[46043]_ , \new_[46044]_ , \new_[46047]_ , \new_[46050]_ ,
    \new_[46051]_ , \new_[46054]_ , \new_[46057]_ , \new_[46058]_ ,
    \new_[46059]_ , \new_[46062]_ , \new_[46065]_ , \new_[46066]_ ,
    \new_[46069]_ , \new_[46072]_ , \new_[46073]_ , \new_[46074]_ ,
    \new_[46077]_ , \new_[46080]_ , \new_[46081]_ , \new_[46084]_ ,
    \new_[46087]_ , \new_[46088]_ , \new_[46089]_ , \new_[46092]_ ,
    \new_[46095]_ , \new_[46096]_ , \new_[46099]_ , \new_[46102]_ ,
    \new_[46103]_ , \new_[46104]_ , \new_[46107]_ , \new_[46110]_ ,
    \new_[46111]_ , \new_[46114]_ , \new_[46117]_ , \new_[46118]_ ,
    \new_[46119]_ , \new_[46122]_ , \new_[46125]_ , \new_[46126]_ ,
    \new_[46129]_ , \new_[46132]_ , \new_[46133]_ , \new_[46134]_ ,
    \new_[46137]_ , \new_[46140]_ , \new_[46141]_ , \new_[46144]_ ,
    \new_[46147]_ , \new_[46148]_ , \new_[46149]_ , \new_[46152]_ ,
    \new_[46155]_ , \new_[46156]_ , \new_[46159]_ , \new_[46162]_ ,
    \new_[46163]_ , \new_[46164]_ , \new_[46167]_ , \new_[46170]_ ,
    \new_[46171]_ , \new_[46174]_ , \new_[46177]_ , \new_[46178]_ ,
    \new_[46179]_ , \new_[46182]_ , \new_[46185]_ , \new_[46186]_ ,
    \new_[46189]_ , \new_[46192]_ , \new_[46193]_ , \new_[46194]_ ,
    \new_[46197]_ , \new_[46200]_ , \new_[46201]_ , \new_[46204]_ ,
    \new_[46207]_ , \new_[46208]_ , \new_[46209]_ , \new_[46212]_ ,
    \new_[46215]_ , \new_[46216]_ , \new_[46219]_ , \new_[46222]_ ,
    \new_[46223]_ , \new_[46224]_ , \new_[46227]_ , \new_[46230]_ ,
    \new_[46231]_ , \new_[46234]_ , \new_[46237]_ , \new_[46238]_ ,
    \new_[46239]_ , \new_[46242]_ , \new_[46245]_ , \new_[46246]_ ,
    \new_[46249]_ , \new_[46252]_ , \new_[46253]_ , \new_[46254]_ ,
    \new_[46257]_ , \new_[46260]_ , \new_[46261]_ , \new_[46264]_ ,
    \new_[46267]_ , \new_[46268]_ , \new_[46269]_ , \new_[46272]_ ,
    \new_[46275]_ , \new_[46276]_ , \new_[46279]_ , \new_[46282]_ ,
    \new_[46283]_ , \new_[46284]_ , \new_[46287]_ , \new_[46290]_ ,
    \new_[46291]_ , \new_[46294]_ , \new_[46297]_ , \new_[46298]_ ,
    \new_[46299]_ , \new_[46302]_ , \new_[46305]_ , \new_[46306]_ ,
    \new_[46309]_ , \new_[46312]_ , \new_[46313]_ , \new_[46314]_ ,
    \new_[46317]_ , \new_[46320]_ , \new_[46321]_ , \new_[46324]_ ,
    \new_[46327]_ , \new_[46328]_ , \new_[46329]_ , \new_[46332]_ ,
    \new_[46335]_ , \new_[46336]_ , \new_[46339]_ , \new_[46342]_ ,
    \new_[46343]_ , \new_[46344]_ , \new_[46347]_ , \new_[46350]_ ,
    \new_[46351]_ , \new_[46354]_ , \new_[46357]_ , \new_[46358]_ ,
    \new_[46359]_ , \new_[46362]_ , \new_[46365]_ , \new_[46366]_ ,
    \new_[46369]_ , \new_[46372]_ , \new_[46373]_ , \new_[46374]_ ,
    \new_[46377]_ , \new_[46380]_ , \new_[46381]_ , \new_[46384]_ ,
    \new_[46387]_ , \new_[46388]_ , \new_[46389]_ , \new_[46392]_ ,
    \new_[46395]_ , \new_[46396]_ , \new_[46399]_ , \new_[46402]_ ,
    \new_[46403]_ , \new_[46404]_ , \new_[46407]_ , \new_[46410]_ ,
    \new_[46411]_ , \new_[46414]_ , \new_[46417]_ , \new_[46418]_ ,
    \new_[46419]_ , \new_[46422]_ , \new_[46425]_ , \new_[46426]_ ,
    \new_[46429]_ , \new_[46432]_ , \new_[46433]_ , \new_[46434]_ ,
    \new_[46437]_ , \new_[46440]_ , \new_[46441]_ , \new_[46444]_ ,
    \new_[46447]_ , \new_[46448]_ , \new_[46449]_ , \new_[46452]_ ,
    \new_[46455]_ , \new_[46456]_ , \new_[46459]_ , \new_[46462]_ ,
    \new_[46463]_ , \new_[46464]_ , \new_[46467]_ , \new_[46470]_ ,
    \new_[46471]_ , \new_[46474]_ , \new_[46477]_ , \new_[46478]_ ,
    \new_[46479]_ , \new_[46482]_ , \new_[46485]_ , \new_[46486]_ ,
    \new_[46489]_ , \new_[46492]_ , \new_[46493]_ , \new_[46494]_ ,
    \new_[46497]_ , \new_[46500]_ , \new_[46501]_ , \new_[46504]_ ,
    \new_[46507]_ , \new_[46508]_ , \new_[46509]_ , \new_[46512]_ ,
    \new_[46515]_ , \new_[46516]_ , \new_[46519]_ , \new_[46522]_ ,
    \new_[46523]_ , \new_[46524]_ , \new_[46527]_ , \new_[46530]_ ,
    \new_[46531]_ , \new_[46534]_ , \new_[46537]_ , \new_[46538]_ ,
    \new_[46539]_ , \new_[46542]_ , \new_[46545]_ , \new_[46546]_ ,
    \new_[46549]_ , \new_[46552]_ , \new_[46553]_ , \new_[46554]_ ,
    \new_[46557]_ , \new_[46560]_ , \new_[46561]_ , \new_[46564]_ ,
    \new_[46567]_ , \new_[46568]_ , \new_[46569]_ , \new_[46572]_ ,
    \new_[46575]_ , \new_[46576]_ , \new_[46579]_ , \new_[46582]_ ,
    \new_[46583]_ , \new_[46584]_ , \new_[46587]_ , \new_[46590]_ ,
    \new_[46591]_ , \new_[46594]_ , \new_[46597]_ , \new_[46598]_ ,
    \new_[46599]_ , \new_[46602]_ , \new_[46605]_ , \new_[46606]_ ,
    \new_[46609]_ , \new_[46612]_ , \new_[46613]_ , \new_[46614]_ ,
    \new_[46617]_ , \new_[46620]_ , \new_[46621]_ , \new_[46624]_ ,
    \new_[46627]_ , \new_[46628]_ , \new_[46629]_ , \new_[46632]_ ,
    \new_[46635]_ , \new_[46636]_ , \new_[46639]_ , \new_[46642]_ ,
    \new_[46643]_ , \new_[46644]_ , \new_[46647]_ , \new_[46650]_ ,
    \new_[46651]_ , \new_[46654]_ , \new_[46657]_ , \new_[46658]_ ,
    \new_[46659]_ , \new_[46662]_ , \new_[46665]_ , \new_[46666]_ ,
    \new_[46669]_ , \new_[46672]_ , \new_[46673]_ , \new_[46674]_ ,
    \new_[46677]_ , \new_[46680]_ , \new_[46681]_ , \new_[46684]_ ,
    \new_[46687]_ , \new_[46688]_ , \new_[46689]_ , \new_[46692]_ ,
    \new_[46695]_ , \new_[46696]_ , \new_[46699]_ , \new_[46702]_ ,
    \new_[46703]_ , \new_[46704]_ , \new_[46707]_ , \new_[46710]_ ,
    \new_[46711]_ , \new_[46714]_ , \new_[46717]_ , \new_[46718]_ ,
    \new_[46719]_ , \new_[46722]_ , \new_[46725]_ , \new_[46726]_ ,
    \new_[46729]_ , \new_[46732]_ , \new_[46733]_ , \new_[46734]_ ,
    \new_[46737]_ , \new_[46740]_ , \new_[46741]_ , \new_[46744]_ ,
    \new_[46747]_ , \new_[46748]_ , \new_[46749]_ , \new_[46752]_ ,
    \new_[46755]_ , \new_[46756]_ , \new_[46759]_ , \new_[46762]_ ,
    \new_[46763]_ , \new_[46764]_ , \new_[46767]_ , \new_[46770]_ ,
    \new_[46771]_ , \new_[46774]_ , \new_[46777]_ , \new_[46778]_ ,
    \new_[46779]_ , \new_[46782]_ , \new_[46785]_ , \new_[46786]_ ,
    \new_[46789]_ , \new_[46792]_ , \new_[46793]_ , \new_[46794]_ ,
    \new_[46797]_ , \new_[46800]_ , \new_[46801]_ , \new_[46804]_ ,
    \new_[46807]_ , \new_[46808]_ , \new_[46809]_ , \new_[46812]_ ,
    \new_[46815]_ , \new_[46816]_ , \new_[46819]_ , \new_[46822]_ ,
    \new_[46823]_ , \new_[46824]_ , \new_[46827]_ , \new_[46830]_ ,
    \new_[46831]_ , \new_[46834]_ , \new_[46837]_ , \new_[46838]_ ,
    \new_[46839]_ , \new_[46842]_ , \new_[46845]_ , \new_[46846]_ ,
    \new_[46849]_ , \new_[46852]_ , \new_[46853]_ , \new_[46854]_ ,
    \new_[46857]_ , \new_[46860]_ , \new_[46861]_ , \new_[46864]_ ,
    \new_[46867]_ , \new_[46868]_ , \new_[46869]_ , \new_[46872]_ ,
    \new_[46875]_ , \new_[46876]_ , \new_[46879]_ , \new_[46882]_ ,
    \new_[46883]_ , \new_[46884]_ , \new_[46887]_ , \new_[46890]_ ,
    \new_[46891]_ , \new_[46894]_ , \new_[46897]_ , \new_[46898]_ ,
    \new_[46899]_ , \new_[46902]_ , \new_[46905]_ , \new_[46906]_ ,
    \new_[46909]_ , \new_[46912]_ , \new_[46913]_ , \new_[46914]_ ,
    \new_[46917]_ , \new_[46920]_ , \new_[46921]_ , \new_[46924]_ ,
    \new_[46927]_ , \new_[46928]_ , \new_[46929]_ , \new_[46932]_ ,
    \new_[46935]_ , \new_[46936]_ , \new_[46939]_ , \new_[46942]_ ,
    \new_[46943]_ , \new_[46944]_ , \new_[46947]_ , \new_[46950]_ ,
    \new_[46951]_ , \new_[46954]_ , \new_[46957]_ , \new_[46958]_ ,
    \new_[46959]_ , \new_[46962]_ , \new_[46965]_ , \new_[46966]_ ,
    \new_[46969]_ , \new_[46972]_ , \new_[46973]_ , \new_[46974]_ ,
    \new_[46977]_ , \new_[46980]_ , \new_[46981]_ , \new_[46984]_ ,
    \new_[46987]_ , \new_[46988]_ , \new_[46989]_ , \new_[46992]_ ,
    \new_[46995]_ , \new_[46996]_ , \new_[46999]_ , \new_[47002]_ ,
    \new_[47003]_ , \new_[47004]_ , \new_[47007]_ , \new_[47010]_ ,
    \new_[47011]_ , \new_[47014]_ , \new_[47017]_ , \new_[47018]_ ,
    \new_[47019]_ , \new_[47022]_ , \new_[47025]_ , \new_[47026]_ ,
    \new_[47029]_ , \new_[47032]_ , \new_[47033]_ , \new_[47034]_ ,
    \new_[47037]_ , \new_[47040]_ , \new_[47041]_ , \new_[47044]_ ,
    \new_[47047]_ , \new_[47048]_ , \new_[47049]_ , \new_[47052]_ ,
    \new_[47055]_ , \new_[47056]_ , \new_[47059]_ , \new_[47062]_ ,
    \new_[47063]_ , \new_[47064]_ , \new_[47067]_ , \new_[47070]_ ,
    \new_[47071]_ , \new_[47074]_ , \new_[47077]_ , \new_[47078]_ ,
    \new_[47079]_ , \new_[47082]_ , \new_[47085]_ , \new_[47086]_ ,
    \new_[47089]_ , \new_[47092]_ , \new_[47093]_ , \new_[47094]_ ,
    \new_[47097]_ , \new_[47100]_ , \new_[47101]_ , \new_[47104]_ ,
    \new_[47107]_ , \new_[47108]_ , \new_[47109]_ , \new_[47112]_ ,
    \new_[47115]_ , \new_[47116]_ , \new_[47119]_ , \new_[47122]_ ,
    \new_[47123]_ , \new_[47124]_ , \new_[47127]_ , \new_[47130]_ ,
    \new_[47131]_ , \new_[47134]_ , \new_[47137]_ , \new_[47138]_ ,
    \new_[47139]_ , \new_[47142]_ , \new_[47145]_ , \new_[47146]_ ,
    \new_[47149]_ , \new_[47152]_ , \new_[47153]_ , \new_[47154]_ ,
    \new_[47157]_ , \new_[47160]_ , \new_[47161]_ , \new_[47164]_ ,
    \new_[47167]_ , \new_[47168]_ , \new_[47169]_ , \new_[47172]_ ,
    \new_[47175]_ , \new_[47176]_ , \new_[47179]_ , \new_[47182]_ ,
    \new_[47183]_ , \new_[47184]_ , \new_[47187]_ , \new_[47190]_ ,
    \new_[47191]_ , \new_[47194]_ , \new_[47197]_ , \new_[47198]_ ,
    \new_[47199]_ , \new_[47202]_ , \new_[47205]_ , \new_[47206]_ ,
    \new_[47209]_ , \new_[47212]_ , \new_[47213]_ , \new_[47214]_ ,
    \new_[47217]_ , \new_[47220]_ , \new_[47221]_ , \new_[47224]_ ,
    \new_[47227]_ , \new_[47228]_ , \new_[47229]_ , \new_[47232]_ ,
    \new_[47235]_ , \new_[47236]_ , \new_[47239]_ , \new_[47242]_ ,
    \new_[47243]_ , \new_[47244]_ , \new_[47247]_ , \new_[47250]_ ,
    \new_[47251]_ , \new_[47254]_ , \new_[47257]_ , \new_[47258]_ ,
    \new_[47259]_ , \new_[47262]_ , \new_[47265]_ , \new_[47266]_ ,
    \new_[47269]_ , \new_[47272]_ , \new_[47273]_ , \new_[47274]_ ,
    \new_[47277]_ , \new_[47280]_ , \new_[47281]_ , \new_[47284]_ ,
    \new_[47287]_ , \new_[47288]_ , \new_[47289]_ , \new_[47292]_ ,
    \new_[47295]_ , \new_[47296]_ , \new_[47299]_ , \new_[47302]_ ,
    \new_[47303]_ , \new_[47304]_ , \new_[47307]_ , \new_[47310]_ ,
    \new_[47311]_ , \new_[47314]_ , \new_[47317]_ , \new_[47318]_ ,
    \new_[47319]_ , \new_[47322]_ , \new_[47325]_ , \new_[47326]_ ,
    \new_[47329]_ , \new_[47332]_ , \new_[47333]_ , \new_[47334]_ ,
    \new_[47337]_ , \new_[47340]_ , \new_[47341]_ , \new_[47344]_ ,
    \new_[47347]_ , \new_[47348]_ , \new_[47349]_ , \new_[47352]_ ,
    \new_[47355]_ , \new_[47356]_ , \new_[47359]_ , \new_[47362]_ ,
    \new_[47363]_ , \new_[47364]_ , \new_[47367]_ , \new_[47370]_ ,
    \new_[47371]_ , \new_[47374]_ , \new_[47377]_ , \new_[47378]_ ,
    \new_[47379]_ , \new_[47382]_ , \new_[47385]_ , \new_[47386]_ ,
    \new_[47389]_ , \new_[47392]_ , \new_[47393]_ , \new_[47394]_ ,
    \new_[47397]_ , \new_[47400]_ , \new_[47401]_ , \new_[47404]_ ,
    \new_[47407]_ , \new_[47408]_ , \new_[47409]_ , \new_[47412]_ ,
    \new_[47415]_ , \new_[47416]_ , \new_[47419]_ , \new_[47422]_ ,
    \new_[47423]_ , \new_[47424]_ , \new_[47427]_ , \new_[47430]_ ,
    \new_[47431]_ , \new_[47434]_ , \new_[47437]_ , \new_[47438]_ ,
    \new_[47439]_ , \new_[47442]_ , \new_[47445]_ , \new_[47446]_ ,
    \new_[47449]_ , \new_[47452]_ , \new_[47453]_ , \new_[47454]_ ,
    \new_[47457]_ , \new_[47460]_ , \new_[47461]_ , \new_[47464]_ ,
    \new_[47467]_ , \new_[47468]_ , \new_[47469]_ , \new_[47472]_ ,
    \new_[47475]_ , \new_[47476]_ , \new_[47479]_ , \new_[47482]_ ,
    \new_[47483]_ , \new_[47484]_ , \new_[47487]_ , \new_[47490]_ ,
    \new_[47491]_ , \new_[47494]_ , \new_[47497]_ , \new_[47498]_ ,
    \new_[47499]_ , \new_[47502]_ , \new_[47505]_ , \new_[47506]_ ,
    \new_[47509]_ , \new_[47512]_ , \new_[47513]_ , \new_[47514]_ ,
    \new_[47517]_ , \new_[47520]_ , \new_[47521]_ , \new_[47524]_ ,
    \new_[47527]_ , \new_[47528]_ , \new_[47529]_ , \new_[47532]_ ,
    \new_[47535]_ , \new_[47536]_ , \new_[47539]_ , \new_[47542]_ ,
    \new_[47543]_ , \new_[47544]_ , \new_[47547]_ , \new_[47550]_ ,
    \new_[47551]_ , \new_[47554]_ , \new_[47557]_ , \new_[47558]_ ,
    \new_[47559]_ , \new_[47562]_ , \new_[47565]_ , \new_[47566]_ ,
    \new_[47569]_ , \new_[47572]_ , \new_[47573]_ , \new_[47574]_ ,
    \new_[47577]_ , \new_[47580]_ , \new_[47581]_ , \new_[47584]_ ,
    \new_[47587]_ , \new_[47588]_ , \new_[47589]_ , \new_[47592]_ ,
    \new_[47595]_ , \new_[47596]_ , \new_[47599]_ , \new_[47602]_ ,
    \new_[47603]_ , \new_[47604]_ , \new_[47607]_ , \new_[47610]_ ,
    \new_[47611]_ , \new_[47614]_ , \new_[47617]_ , \new_[47618]_ ,
    \new_[47619]_ , \new_[47622]_ , \new_[47625]_ , \new_[47626]_ ,
    \new_[47629]_ , \new_[47632]_ , \new_[47633]_ , \new_[47634]_ ,
    \new_[47637]_ , \new_[47640]_ , \new_[47641]_ , \new_[47644]_ ,
    \new_[47647]_ , \new_[47648]_ , \new_[47649]_ , \new_[47652]_ ,
    \new_[47655]_ , \new_[47656]_ , \new_[47659]_ , \new_[47662]_ ,
    \new_[47663]_ , \new_[47664]_ , \new_[47667]_ , \new_[47670]_ ,
    \new_[47671]_ , \new_[47674]_ , \new_[47677]_ , \new_[47678]_ ,
    \new_[47679]_ , \new_[47682]_ , \new_[47685]_ , \new_[47686]_ ,
    \new_[47689]_ , \new_[47692]_ , \new_[47693]_ , \new_[47694]_ ,
    \new_[47697]_ , \new_[47700]_ , \new_[47701]_ , \new_[47704]_ ,
    \new_[47707]_ , \new_[47708]_ , \new_[47709]_ , \new_[47712]_ ,
    \new_[47715]_ , \new_[47716]_ , \new_[47719]_ , \new_[47722]_ ,
    \new_[47723]_ , \new_[47724]_ , \new_[47727]_ , \new_[47730]_ ,
    \new_[47731]_ , \new_[47734]_ , \new_[47737]_ , \new_[47738]_ ,
    \new_[47739]_ , \new_[47742]_ , \new_[47745]_ , \new_[47746]_ ,
    \new_[47749]_ , \new_[47752]_ , \new_[47753]_ , \new_[47754]_ ,
    \new_[47757]_ , \new_[47760]_ , \new_[47761]_ , \new_[47764]_ ,
    \new_[47767]_ , \new_[47768]_ , \new_[47769]_ , \new_[47772]_ ,
    \new_[47775]_ , \new_[47776]_ , \new_[47779]_ , \new_[47782]_ ,
    \new_[47783]_ , \new_[47784]_ , \new_[47787]_ , \new_[47790]_ ,
    \new_[47791]_ , \new_[47794]_ , \new_[47797]_ , \new_[47798]_ ,
    \new_[47799]_ , \new_[47802]_ , \new_[47805]_ , \new_[47806]_ ,
    \new_[47809]_ , \new_[47812]_ , \new_[47813]_ , \new_[47814]_ ,
    \new_[47817]_ , \new_[47820]_ , \new_[47821]_ , \new_[47824]_ ,
    \new_[47827]_ , \new_[47828]_ , \new_[47829]_ , \new_[47832]_ ,
    \new_[47835]_ , \new_[47836]_ , \new_[47839]_ , \new_[47842]_ ,
    \new_[47843]_ , \new_[47844]_ , \new_[47847]_ , \new_[47850]_ ,
    \new_[47851]_ , \new_[47854]_ , \new_[47857]_ , \new_[47858]_ ,
    \new_[47859]_ , \new_[47862]_ , \new_[47865]_ , \new_[47866]_ ,
    \new_[47869]_ , \new_[47872]_ , \new_[47873]_ , \new_[47874]_ ,
    \new_[47877]_ , \new_[47880]_ , \new_[47881]_ , \new_[47884]_ ,
    \new_[47887]_ , \new_[47888]_ , \new_[47889]_ , \new_[47892]_ ,
    \new_[47895]_ , \new_[47896]_ , \new_[47899]_ , \new_[47902]_ ,
    \new_[47903]_ , \new_[47904]_ , \new_[47907]_ , \new_[47910]_ ,
    \new_[47911]_ , \new_[47914]_ , \new_[47917]_ , \new_[47918]_ ,
    \new_[47919]_ , \new_[47922]_ , \new_[47925]_ , \new_[47926]_ ,
    \new_[47929]_ , \new_[47932]_ , \new_[47933]_ , \new_[47934]_ ,
    \new_[47937]_ , \new_[47940]_ , \new_[47941]_ , \new_[47944]_ ,
    \new_[47947]_ , \new_[47948]_ , \new_[47949]_ , \new_[47952]_ ,
    \new_[47955]_ , \new_[47956]_ , \new_[47959]_ , \new_[47962]_ ,
    \new_[47963]_ , \new_[47964]_ , \new_[47967]_ , \new_[47970]_ ,
    \new_[47971]_ , \new_[47974]_ , \new_[47977]_ , \new_[47978]_ ,
    \new_[47979]_ , \new_[47982]_ , \new_[47985]_ , \new_[47986]_ ,
    \new_[47989]_ , \new_[47992]_ , \new_[47993]_ , \new_[47994]_ ,
    \new_[47997]_ , \new_[48000]_ , \new_[48001]_ , \new_[48004]_ ,
    \new_[48007]_ , \new_[48008]_ , \new_[48009]_ , \new_[48012]_ ,
    \new_[48015]_ , \new_[48016]_ , \new_[48019]_ , \new_[48022]_ ,
    \new_[48023]_ , \new_[48024]_ , \new_[48027]_ , \new_[48030]_ ,
    \new_[48031]_ , \new_[48034]_ , \new_[48037]_ , \new_[48038]_ ,
    \new_[48039]_ , \new_[48042]_ , \new_[48045]_ , \new_[48046]_ ,
    \new_[48049]_ , \new_[48052]_ , \new_[48053]_ , \new_[48054]_ ,
    \new_[48057]_ , \new_[48060]_ , \new_[48061]_ , \new_[48064]_ ,
    \new_[48067]_ , \new_[48068]_ , \new_[48069]_ , \new_[48072]_ ,
    \new_[48075]_ , \new_[48076]_ , \new_[48079]_ , \new_[48082]_ ,
    \new_[48083]_ , \new_[48084]_ , \new_[48087]_ , \new_[48090]_ ,
    \new_[48091]_ , \new_[48094]_ , \new_[48097]_ , \new_[48098]_ ,
    \new_[48099]_ , \new_[48102]_ , \new_[48105]_ , \new_[48106]_ ,
    \new_[48109]_ , \new_[48112]_ , \new_[48113]_ , \new_[48114]_ ,
    \new_[48117]_ , \new_[48120]_ , \new_[48121]_ , \new_[48124]_ ,
    \new_[48127]_ , \new_[48128]_ , \new_[48129]_ , \new_[48132]_ ,
    \new_[48135]_ , \new_[48136]_ , \new_[48139]_ , \new_[48142]_ ,
    \new_[48143]_ , \new_[48144]_ , \new_[48147]_ , \new_[48150]_ ,
    \new_[48151]_ , \new_[48154]_ , \new_[48157]_ , \new_[48158]_ ,
    \new_[48159]_ , \new_[48162]_ , \new_[48165]_ , \new_[48166]_ ,
    \new_[48169]_ , \new_[48172]_ , \new_[48173]_ , \new_[48174]_ ,
    \new_[48177]_ , \new_[48180]_ , \new_[48181]_ , \new_[48184]_ ,
    \new_[48187]_ , \new_[48188]_ , \new_[48189]_ , \new_[48192]_ ,
    \new_[48195]_ , \new_[48196]_ , \new_[48199]_ , \new_[48202]_ ,
    \new_[48203]_ , \new_[48204]_ , \new_[48207]_ , \new_[48210]_ ,
    \new_[48211]_ , \new_[48214]_ , \new_[48217]_ , \new_[48218]_ ,
    \new_[48219]_ , \new_[48222]_ , \new_[48225]_ , \new_[48226]_ ,
    \new_[48229]_ , \new_[48232]_ , \new_[48233]_ , \new_[48234]_ ,
    \new_[48237]_ , \new_[48240]_ , \new_[48241]_ , \new_[48244]_ ,
    \new_[48247]_ , \new_[48248]_ , \new_[48249]_ , \new_[48252]_ ,
    \new_[48255]_ , \new_[48256]_ , \new_[48259]_ , \new_[48262]_ ,
    \new_[48263]_ , \new_[48264]_ , \new_[48267]_ , \new_[48270]_ ,
    \new_[48271]_ , \new_[48274]_ , \new_[48277]_ , \new_[48278]_ ,
    \new_[48279]_ , \new_[48282]_ , \new_[48285]_ , \new_[48286]_ ,
    \new_[48289]_ , \new_[48292]_ , \new_[48293]_ , \new_[48294]_ ,
    \new_[48297]_ , \new_[48300]_ , \new_[48301]_ , \new_[48304]_ ,
    \new_[48307]_ , \new_[48308]_ , \new_[48309]_ , \new_[48312]_ ,
    \new_[48315]_ , \new_[48316]_ , \new_[48319]_ , \new_[48322]_ ,
    \new_[48323]_ , \new_[48324]_ , \new_[48327]_ , \new_[48330]_ ,
    \new_[48331]_ , \new_[48334]_ , \new_[48337]_ , \new_[48338]_ ,
    \new_[48339]_ , \new_[48342]_ , \new_[48345]_ , \new_[48346]_ ,
    \new_[48349]_ , \new_[48352]_ , \new_[48353]_ , \new_[48354]_ ,
    \new_[48357]_ , \new_[48360]_ , \new_[48361]_ , \new_[48364]_ ,
    \new_[48367]_ , \new_[48368]_ , \new_[48369]_ , \new_[48372]_ ,
    \new_[48375]_ , \new_[48376]_ , \new_[48379]_ , \new_[48382]_ ,
    \new_[48383]_ , \new_[48384]_ , \new_[48387]_ , \new_[48390]_ ,
    \new_[48391]_ , \new_[48394]_ , \new_[48397]_ , \new_[48398]_ ,
    \new_[48399]_ , \new_[48402]_ , \new_[48405]_ , \new_[48406]_ ,
    \new_[48409]_ , \new_[48412]_ , \new_[48413]_ , \new_[48414]_ ,
    \new_[48417]_ , \new_[48420]_ , \new_[48421]_ , \new_[48424]_ ,
    \new_[48427]_ , \new_[48428]_ , \new_[48429]_ , \new_[48432]_ ,
    \new_[48435]_ , \new_[48436]_ , \new_[48439]_ , \new_[48442]_ ,
    \new_[48443]_ , \new_[48444]_ , \new_[48447]_ , \new_[48450]_ ,
    \new_[48451]_ , \new_[48454]_ , \new_[48457]_ , \new_[48458]_ ,
    \new_[48459]_ , \new_[48462]_ , \new_[48465]_ , \new_[48466]_ ,
    \new_[48469]_ , \new_[48472]_ , \new_[48473]_ , \new_[48474]_ ,
    \new_[48477]_ , \new_[48480]_ , \new_[48481]_ , \new_[48484]_ ,
    \new_[48487]_ , \new_[48488]_ , \new_[48489]_ , \new_[48492]_ ,
    \new_[48495]_ , \new_[48496]_ , \new_[48499]_ , \new_[48502]_ ,
    \new_[48503]_ , \new_[48504]_ , \new_[48507]_ , \new_[48510]_ ,
    \new_[48511]_ , \new_[48514]_ , \new_[48517]_ , \new_[48518]_ ,
    \new_[48519]_ , \new_[48522]_ , \new_[48525]_ , \new_[48526]_ ,
    \new_[48529]_ , \new_[48532]_ , \new_[48533]_ , \new_[48534]_ ,
    \new_[48537]_ , \new_[48540]_ , \new_[48541]_ , \new_[48544]_ ,
    \new_[48547]_ , \new_[48548]_ , \new_[48549]_ , \new_[48552]_ ,
    \new_[48555]_ , \new_[48556]_ , \new_[48559]_ , \new_[48562]_ ,
    \new_[48563]_ , \new_[48564]_ , \new_[48567]_ , \new_[48570]_ ,
    \new_[48571]_ , \new_[48574]_ , \new_[48577]_ , \new_[48578]_ ,
    \new_[48579]_ , \new_[48582]_ , \new_[48585]_ , \new_[48586]_ ,
    \new_[48589]_ , \new_[48592]_ , \new_[48593]_ , \new_[48594]_ ,
    \new_[48597]_ , \new_[48600]_ , \new_[48601]_ , \new_[48604]_ ,
    \new_[48607]_ , \new_[48608]_ , \new_[48609]_ , \new_[48612]_ ,
    \new_[48615]_ , \new_[48616]_ , \new_[48619]_ , \new_[48622]_ ,
    \new_[48623]_ , \new_[48624]_ , \new_[48627]_ , \new_[48630]_ ,
    \new_[48631]_ , \new_[48634]_ , \new_[48637]_ , \new_[48638]_ ,
    \new_[48639]_ , \new_[48642]_ , \new_[48645]_ , \new_[48646]_ ,
    \new_[48649]_ , \new_[48652]_ , \new_[48653]_ , \new_[48654]_ ,
    \new_[48657]_ , \new_[48660]_ , \new_[48661]_ , \new_[48664]_ ,
    \new_[48667]_ , \new_[48668]_ , \new_[48669]_ , \new_[48672]_ ,
    \new_[48675]_ , \new_[48676]_ , \new_[48679]_ , \new_[48682]_ ,
    \new_[48683]_ , \new_[48684]_ , \new_[48687]_ , \new_[48690]_ ,
    \new_[48691]_ , \new_[48694]_ , \new_[48697]_ , \new_[48698]_ ,
    \new_[48699]_ , \new_[48702]_ , \new_[48705]_ , \new_[48706]_ ,
    \new_[48709]_ , \new_[48712]_ , \new_[48713]_ , \new_[48714]_ ,
    \new_[48717]_ , \new_[48720]_ , \new_[48721]_ , \new_[48724]_ ,
    \new_[48727]_ , \new_[48728]_ , \new_[48729]_ , \new_[48732]_ ,
    \new_[48735]_ , \new_[48736]_ , \new_[48739]_ , \new_[48742]_ ,
    \new_[48743]_ , \new_[48744]_ , \new_[48747]_ , \new_[48750]_ ,
    \new_[48751]_ , \new_[48754]_ , \new_[48757]_ , \new_[48758]_ ,
    \new_[48759]_ , \new_[48762]_ , \new_[48765]_ , \new_[48766]_ ,
    \new_[48769]_ , \new_[48772]_ , \new_[48773]_ , \new_[48774]_ ,
    \new_[48777]_ , \new_[48780]_ , \new_[48781]_ , \new_[48784]_ ,
    \new_[48787]_ , \new_[48788]_ , \new_[48789]_ , \new_[48792]_ ,
    \new_[48795]_ , \new_[48796]_ , \new_[48799]_ , \new_[48802]_ ,
    \new_[48803]_ , \new_[48804]_ , \new_[48807]_ , \new_[48810]_ ,
    \new_[48811]_ , \new_[48814]_ , \new_[48817]_ , \new_[48818]_ ,
    \new_[48819]_ , \new_[48822]_ , \new_[48825]_ , \new_[48826]_ ,
    \new_[48829]_ , \new_[48832]_ , \new_[48833]_ , \new_[48834]_ ,
    \new_[48837]_ , \new_[48840]_ , \new_[48841]_ , \new_[48844]_ ,
    \new_[48847]_ , \new_[48848]_ , \new_[48849]_ , \new_[48852]_ ,
    \new_[48855]_ , \new_[48856]_ , \new_[48859]_ , \new_[48862]_ ,
    \new_[48863]_ , \new_[48864]_ , \new_[48867]_ , \new_[48870]_ ,
    \new_[48871]_ , \new_[48874]_ , \new_[48877]_ , \new_[48878]_ ,
    \new_[48879]_ , \new_[48882]_ , \new_[48885]_ , \new_[48886]_ ,
    \new_[48889]_ , \new_[48892]_ , \new_[48893]_ , \new_[48894]_ ,
    \new_[48897]_ , \new_[48900]_ , \new_[48901]_ , \new_[48904]_ ,
    \new_[48907]_ , \new_[48908]_ , \new_[48909]_ , \new_[48912]_ ,
    \new_[48915]_ , \new_[48916]_ , \new_[48919]_ , \new_[48922]_ ,
    \new_[48923]_ , \new_[48924]_ , \new_[48927]_ , \new_[48930]_ ,
    \new_[48931]_ , \new_[48934]_ , \new_[48937]_ , \new_[48938]_ ,
    \new_[48939]_ , \new_[48942]_ , \new_[48945]_ , \new_[48946]_ ,
    \new_[48949]_ , \new_[48952]_ , \new_[48953]_ , \new_[48954]_ ,
    \new_[48957]_ , \new_[48960]_ , \new_[48961]_ , \new_[48964]_ ,
    \new_[48967]_ , \new_[48968]_ , \new_[48969]_ , \new_[48972]_ ,
    \new_[48975]_ , \new_[48976]_ , \new_[48979]_ , \new_[48982]_ ,
    \new_[48983]_ , \new_[48984]_ , \new_[48987]_ , \new_[48990]_ ,
    \new_[48991]_ , \new_[48994]_ , \new_[48997]_ , \new_[48998]_ ,
    \new_[48999]_ , \new_[49002]_ , \new_[49005]_ , \new_[49006]_ ,
    \new_[49009]_ , \new_[49012]_ , \new_[49013]_ , \new_[49014]_ ,
    \new_[49017]_ , \new_[49020]_ , \new_[49021]_ , \new_[49024]_ ,
    \new_[49027]_ , \new_[49028]_ , \new_[49029]_ , \new_[49032]_ ,
    \new_[49035]_ , \new_[49036]_ , \new_[49039]_ , \new_[49042]_ ,
    \new_[49043]_ , \new_[49044]_ , \new_[49047]_ , \new_[49050]_ ,
    \new_[49051]_ , \new_[49054]_ , \new_[49057]_ , \new_[49058]_ ,
    \new_[49059]_ , \new_[49062]_ , \new_[49065]_ , \new_[49066]_ ,
    \new_[49069]_ , \new_[49072]_ , \new_[49073]_ , \new_[49074]_ ,
    \new_[49077]_ , \new_[49080]_ , \new_[49081]_ , \new_[49084]_ ,
    \new_[49087]_ , \new_[49088]_ , \new_[49089]_ , \new_[49092]_ ,
    \new_[49095]_ , \new_[49096]_ , \new_[49099]_ , \new_[49102]_ ,
    \new_[49103]_ , \new_[49104]_ , \new_[49107]_ , \new_[49110]_ ,
    \new_[49111]_ , \new_[49114]_ , \new_[49117]_ , \new_[49118]_ ,
    \new_[49119]_ , \new_[49122]_ , \new_[49125]_ , \new_[49126]_ ,
    \new_[49129]_ , \new_[49132]_ , \new_[49133]_ , \new_[49134]_ ,
    \new_[49137]_ , \new_[49140]_ , \new_[49141]_ , \new_[49144]_ ,
    \new_[49147]_ , \new_[49148]_ , \new_[49149]_ , \new_[49152]_ ,
    \new_[49155]_ , \new_[49156]_ , \new_[49159]_ , \new_[49162]_ ,
    \new_[49163]_ , \new_[49164]_ , \new_[49167]_ , \new_[49170]_ ,
    \new_[49171]_ , \new_[49174]_ , \new_[49177]_ , \new_[49178]_ ,
    \new_[49179]_ , \new_[49182]_ , \new_[49185]_ , \new_[49186]_ ,
    \new_[49189]_ , \new_[49192]_ , \new_[49193]_ , \new_[49194]_ ,
    \new_[49197]_ , \new_[49200]_ , \new_[49201]_ , \new_[49204]_ ,
    \new_[49207]_ , \new_[49208]_ , \new_[49209]_ , \new_[49212]_ ,
    \new_[49215]_ , \new_[49216]_ , \new_[49219]_ , \new_[49222]_ ,
    \new_[49223]_ , \new_[49224]_ , \new_[49227]_ , \new_[49230]_ ,
    \new_[49231]_ , \new_[49234]_ , \new_[49237]_ , \new_[49238]_ ,
    \new_[49239]_ , \new_[49242]_ , \new_[49245]_ , \new_[49246]_ ,
    \new_[49249]_ , \new_[49252]_ , \new_[49253]_ , \new_[49254]_ ,
    \new_[49257]_ , \new_[49260]_ , \new_[49261]_ , \new_[49264]_ ,
    \new_[49267]_ , \new_[49268]_ , \new_[49269]_ , \new_[49272]_ ,
    \new_[49275]_ , \new_[49276]_ , \new_[49279]_ , \new_[49282]_ ,
    \new_[49283]_ , \new_[49284]_ , \new_[49287]_ , \new_[49290]_ ,
    \new_[49291]_ , \new_[49294]_ , \new_[49297]_ , \new_[49298]_ ,
    \new_[49299]_ , \new_[49302]_ , \new_[49305]_ , \new_[49306]_ ,
    \new_[49309]_ , \new_[49312]_ , \new_[49313]_ , \new_[49314]_ ,
    \new_[49317]_ , \new_[49320]_ , \new_[49321]_ , \new_[49324]_ ,
    \new_[49327]_ , \new_[49328]_ , \new_[49329]_ , \new_[49332]_ ,
    \new_[49335]_ , \new_[49336]_ , \new_[49339]_ , \new_[49342]_ ,
    \new_[49343]_ , \new_[49344]_ , \new_[49347]_ , \new_[49350]_ ,
    \new_[49351]_ , \new_[49354]_ , \new_[49357]_ , \new_[49358]_ ,
    \new_[49359]_ , \new_[49362]_ , \new_[49365]_ , \new_[49366]_ ,
    \new_[49369]_ , \new_[49372]_ , \new_[49373]_ , \new_[49374]_ ,
    \new_[49377]_ , \new_[49380]_ , \new_[49381]_ , \new_[49384]_ ,
    \new_[49387]_ , \new_[49388]_ , \new_[49389]_ , \new_[49392]_ ,
    \new_[49395]_ , \new_[49396]_ , \new_[49399]_ , \new_[49402]_ ,
    \new_[49403]_ , \new_[49404]_ , \new_[49407]_ , \new_[49410]_ ,
    \new_[49411]_ , \new_[49414]_ , \new_[49417]_ , \new_[49418]_ ,
    \new_[49419]_ , \new_[49422]_ , \new_[49425]_ , \new_[49426]_ ,
    \new_[49429]_ , \new_[49432]_ , \new_[49433]_ , \new_[49434]_ ,
    \new_[49437]_ , \new_[49440]_ , \new_[49441]_ , \new_[49444]_ ,
    \new_[49447]_ , \new_[49448]_ , \new_[49449]_ , \new_[49452]_ ,
    \new_[49455]_ , \new_[49456]_ , \new_[49459]_ , \new_[49462]_ ,
    \new_[49463]_ , \new_[49464]_ , \new_[49467]_ , \new_[49470]_ ,
    \new_[49471]_ , \new_[49474]_ , \new_[49477]_ , \new_[49478]_ ,
    \new_[49479]_ , \new_[49482]_ , \new_[49485]_ , \new_[49486]_ ,
    \new_[49489]_ , \new_[49492]_ , \new_[49493]_ , \new_[49494]_ ,
    \new_[49497]_ , \new_[49500]_ , \new_[49501]_ , \new_[49504]_ ,
    \new_[49507]_ , \new_[49508]_ , \new_[49509]_ , \new_[49512]_ ,
    \new_[49515]_ , \new_[49516]_ , \new_[49519]_ , \new_[49522]_ ,
    \new_[49523]_ , \new_[49524]_ , \new_[49527]_ , \new_[49530]_ ,
    \new_[49531]_ , \new_[49534]_ , \new_[49537]_ , \new_[49538]_ ,
    \new_[49539]_ , \new_[49542]_ , \new_[49545]_ , \new_[49546]_ ,
    \new_[49549]_ , \new_[49552]_ , \new_[49553]_ , \new_[49554]_ ,
    \new_[49557]_ , \new_[49560]_ , \new_[49561]_ , \new_[49564]_ ,
    \new_[49567]_ , \new_[49568]_ , \new_[49569]_ , \new_[49572]_ ,
    \new_[49575]_ , \new_[49576]_ , \new_[49579]_ , \new_[49582]_ ,
    \new_[49583]_ , \new_[49584]_ , \new_[49587]_ , \new_[49590]_ ,
    \new_[49591]_ , \new_[49594]_ , \new_[49597]_ , \new_[49598]_ ,
    \new_[49599]_ , \new_[49602]_ , \new_[49605]_ , \new_[49606]_ ,
    \new_[49609]_ , \new_[49612]_ , \new_[49613]_ , \new_[49614]_ ,
    \new_[49617]_ , \new_[49620]_ , \new_[49621]_ , \new_[49624]_ ,
    \new_[49627]_ , \new_[49628]_ , \new_[49629]_ , \new_[49632]_ ,
    \new_[49635]_ , \new_[49636]_ , \new_[49639]_ , \new_[49642]_ ,
    \new_[49643]_ , \new_[49644]_ , \new_[49647]_ , \new_[49650]_ ,
    \new_[49651]_ , \new_[49654]_ , \new_[49657]_ , \new_[49658]_ ,
    \new_[49659]_ , \new_[49662]_ , \new_[49665]_ , \new_[49666]_ ,
    \new_[49669]_ , \new_[49672]_ , \new_[49673]_ , \new_[49674]_ ,
    \new_[49677]_ , \new_[49680]_ , \new_[49681]_ , \new_[49684]_ ,
    \new_[49687]_ , \new_[49688]_ , \new_[49689]_ , \new_[49692]_ ,
    \new_[49695]_ , \new_[49696]_ , \new_[49699]_ , \new_[49702]_ ,
    \new_[49703]_ , \new_[49704]_ , \new_[49707]_ , \new_[49710]_ ,
    \new_[49711]_ , \new_[49714]_ , \new_[49717]_ , \new_[49718]_ ,
    \new_[49719]_ , \new_[49722]_ , \new_[49725]_ , \new_[49726]_ ,
    \new_[49729]_ , \new_[49732]_ , \new_[49733]_ , \new_[49734]_ ,
    \new_[49737]_ , \new_[49740]_ , \new_[49741]_ , \new_[49744]_ ,
    \new_[49747]_ , \new_[49748]_ , \new_[49749]_ , \new_[49752]_ ,
    \new_[49755]_ , \new_[49756]_ , \new_[49759]_ , \new_[49762]_ ,
    \new_[49763]_ , \new_[49764]_ , \new_[49767]_ , \new_[49770]_ ,
    \new_[49771]_ , \new_[49774]_ , \new_[49777]_ , \new_[49778]_ ,
    \new_[49779]_ , \new_[49782]_ , \new_[49785]_ , \new_[49786]_ ,
    \new_[49789]_ , \new_[49792]_ , \new_[49793]_ , \new_[49794]_ ,
    \new_[49797]_ , \new_[49800]_ , \new_[49801]_ , \new_[49804]_ ,
    \new_[49807]_ , \new_[49808]_ , \new_[49809]_ , \new_[49812]_ ,
    \new_[49815]_ , \new_[49816]_ , \new_[49819]_ , \new_[49822]_ ,
    \new_[49823]_ , \new_[49824]_ , \new_[49827]_ , \new_[49830]_ ,
    \new_[49831]_ , \new_[49834]_ , \new_[49837]_ , \new_[49838]_ ,
    \new_[49839]_ , \new_[49842]_ , \new_[49845]_ , \new_[49846]_ ,
    \new_[49849]_ , \new_[49852]_ , \new_[49853]_ , \new_[49854]_ ,
    \new_[49857]_ , \new_[49860]_ , \new_[49861]_ , \new_[49864]_ ,
    \new_[49867]_ , \new_[49868]_ , \new_[49869]_ , \new_[49872]_ ,
    \new_[49875]_ , \new_[49876]_ , \new_[49879]_ , \new_[49882]_ ,
    \new_[49883]_ , \new_[49884]_ , \new_[49887]_ , \new_[49890]_ ,
    \new_[49891]_ , \new_[49894]_ , \new_[49897]_ , \new_[49898]_ ,
    \new_[49899]_ , \new_[49902]_ , \new_[49905]_ , \new_[49906]_ ,
    \new_[49909]_ , \new_[49912]_ , \new_[49913]_ , \new_[49914]_ ,
    \new_[49917]_ , \new_[49920]_ , \new_[49921]_ , \new_[49924]_ ,
    \new_[49927]_ , \new_[49928]_ , \new_[49929]_ , \new_[49932]_ ,
    \new_[49935]_ , \new_[49936]_ , \new_[49939]_ , \new_[49942]_ ,
    \new_[49943]_ , \new_[49944]_ , \new_[49947]_ , \new_[49950]_ ,
    \new_[49951]_ , \new_[49954]_ , \new_[49957]_ , \new_[49958]_ ,
    \new_[49959]_ , \new_[49962]_ , \new_[49965]_ , \new_[49966]_ ,
    \new_[49969]_ , \new_[49972]_ , \new_[49973]_ , \new_[49974]_ ,
    \new_[49977]_ , \new_[49980]_ , \new_[49981]_ , \new_[49984]_ ,
    \new_[49987]_ , \new_[49988]_ , \new_[49989]_ , \new_[49992]_ ,
    \new_[49995]_ , \new_[49996]_ , \new_[49999]_ , \new_[50002]_ ,
    \new_[50003]_ , \new_[50004]_ , \new_[50007]_ , \new_[50010]_ ,
    \new_[50011]_ , \new_[50014]_ , \new_[50017]_ , \new_[50018]_ ,
    \new_[50019]_ , \new_[50022]_ , \new_[50025]_ , \new_[50026]_ ,
    \new_[50029]_ , \new_[50032]_ , \new_[50033]_ , \new_[50034]_ ,
    \new_[50037]_ , \new_[50040]_ , \new_[50041]_ , \new_[50044]_ ,
    \new_[50047]_ , \new_[50048]_ , \new_[50049]_ , \new_[50052]_ ,
    \new_[50055]_ , \new_[50056]_ , \new_[50059]_ , \new_[50062]_ ,
    \new_[50063]_ , \new_[50064]_ , \new_[50067]_ , \new_[50070]_ ,
    \new_[50071]_ , \new_[50074]_ , \new_[50077]_ , \new_[50078]_ ,
    \new_[50079]_ , \new_[50082]_ , \new_[50085]_ , \new_[50086]_ ,
    \new_[50089]_ , \new_[50092]_ , \new_[50093]_ , \new_[50094]_ ,
    \new_[50097]_ , \new_[50100]_ , \new_[50101]_ , \new_[50104]_ ,
    \new_[50107]_ , \new_[50108]_ , \new_[50109]_ , \new_[50112]_ ,
    \new_[50115]_ , \new_[50116]_ , \new_[50119]_ , \new_[50122]_ ,
    \new_[50123]_ , \new_[50124]_ , \new_[50127]_ , \new_[50130]_ ,
    \new_[50131]_ , \new_[50134]_ , \new_[50137]_ , \new_[50138]_ ,
    \new_[50139]_ , \new_[50142]_ , \new_[50145]_ , \new_[50146]_ ,
    \new_[50149]_ , \new_[50152]_ , \new_[50153]_ , \new_[50154]_ ,
    \new_[50157]_ , \new_[50160]_ , \new_[50161]_ , \new_[50164]_ ,
    \new_[50167]_ , \new_[50168]_ , \new_[50169]_ , \new_[50172]_ ,
    \new_[50175]_ , \new_[50176]_ , \new_[50179]_ , \new_[50182]_ ,
    \new_[50183]_ , \new_[50184]_ , \new_[50187]_ , \new_[50190]_ ,
    \new_[50191]_ , \new_[50194]_ , \new_[50197]_ , \new_[50198]_ ,
    \new_[50199]_ , \new_[50202]_ , \new_[50205]_ , \new_[50206]_ ,
    \new_[50209]_ , \new_[50212]_ , \new_[50213]_ , \new_[50214]_ ,
    \new_[50217]_ , \new_[50220]_ , \new_[50221]_ , \new_[50224]_ ,
    \new_[50227]_ , \new_[50228]_ , \new_[50229]_ , \new_[50232]_ ,
    \new_[50235]_ , \new_[50236]_ , \new_[50239]_ , \new_[50242]_ ,
    \new_[50243]_ , \new_[50244]_ , \new_[50247]_ , \new_[50250]_ ,
    \new_[50251]_ , \new_[50254]_ , \new_[50257]_ , \new_[50258]_ ,
    \new_[50259]_ , \new_[50262]_ , \new_[50265]_ , \new_[50266]_ ,
    \new_[50269]_ , \new_[50272]_ , \new_[50273]_ , \new_[50274]_ ,
    \new_[50277]_ , \new_[50280]_ , \new_[50281]_ , \new_[50284]_ ,
    \new_[50287]_ , \new_[50288]_ , \new_[50289]_ , \new_[50292]_ ,
    \new_[50295]_ , \new_[50296]_ , \new_[50299]_ , \new_[50302]_ ,
    \new_[50303]_ , \new_[50304]_ , \new_[50307]_ , \new_[50310]_ ,
    \new_[50311]_ , \new_[50314]_ , \new_[50317]_ , \new_[50318]_ ,
    \new_[50319]_ , \new_[50322]_ , \new_[50325]_ , \new_[50326]_ ,
    \new_[50329]_ , \new_[50332]_ , \new_[50333]_ , \new_[50334]_ ,
    \new_[50337]_ , \new_[50340]_ , \new_[50341]_ , \new_[50344]_ ,
    \new_[50347]_ , \new_[50348]_ , \new_[50349]_ , \new_[50352]_ ,
    \new_[50355]_ , \new_[50356]_ , \new_[50359]_ , \new_[50362]_ ,
    \new_[50363]_ , \new_[50364]_ , \new_[50367]_ , \new_[50370]_ ,
    \new_[50371]_ , \new_[50374]_ , \new_[50377]_ , \new_[50378]_ ,
    \new_[50379]_ , \new_[50382]_ , \new_[50385]_ , \new_[50386]_ ,
    \new_[50389]_ , \new_[50392]_ , \new_[50393]_ , \new_[50394]_ ,
    \new_[50397]_ , \new_[50400]_ , \new_[50401]_ , \new_[50404]_ ,
    \new_[50407]_ , \new_[50408]_ , \new_[50409]_ , \new_[50412]_ ,
    \new_[50415]_ , \new_[50416]_ , \new_[50419]_ , \new_[50422]_ ,
    \new_[50423]_ , \new_[50424]_ , \new_[50427]_ , \new_[50430]_ ,
    \new_[50431]_ , \new_[50434]_ , \new_[50437]_ , \new_[50438]_ ,
    \new_[50439]_ , \new_[50442]_ , \new_[50445]_ , \new_[50446]_ ,
    \new_[50449]_ , \new_[50452]_ , \new_[50453]_ , \new_[50454]_ ,
    \new_[50457]_ , \new_[50460]_ , \new_[50461]_ , \new_[50464]_ ,
    \new_[50467]_ , \new_[50468]_ , \new_[50469]_ , \new_[50472]_ ,
    \new_[50475]_ , \new_[50476]_ , \new_[50479]_ , \new_[50482]_ ,
    \new_[50483]_ , \new_[50484]_ , \new_[50487]_ , \new_[50490]_ ,
    \new_[50491]_ , \new_[50494]_ , \new_[50497]_ , \new_[50498]_ ,
    \new_[50499]_ , \new_[50502]_ , \new_[50505]_ , \new_[50506]_ ,
    \new_[50509]_ , \new_[50512]_ , \new_[50513]_ , \new_[50514]_ ,
    \new_[50517]_ , \new_[50520]_ , \new_[50521]_ , \new_[50524]_ ,
    \new_[50527]_ , \new_[50528]_ , \new_[50529]_ , \new_[50532]_ ,
    \new_[50535]_ , \new_[50536]_ , \new_[50539]_ , \new_[50542]_ ,
    \new_[50543]_ , \new_[50544]_ , \new_[50547]_ , \new_[50550]_ ,
    \new_[50551]_ , \new_[50554]_ , \new_[50557]_ , \new_[50558]_ ,
    \new_[50559]_ , \new_[50562]_ , \new_[50565]_ , \new_[50566]_ ,
    \new_[50569]_ , \new_[50572]_ , \new_[50573]_ , \new_[50574]_ ,
    \new_[50577]_ , \new_[50580]_ , \new_[50581]_ , \new_[50584]_ ,
    \new_[50587]_ , \new_[50588]_ , \new_[50589]_ , \new_[50592]_ ,
    \new_[50595]_ , \new_[50596]_ , \new_[50599]_ , \new_[50602]_ ,
    \new_[50603]_ , \new_[50604]_ , \new_[50607]_ , \new_[50610]_ ,
    \new_[50611]_ , \new_[50614]_ , \new_[50617]_ , \new_[50618]_ ,
    \new_[50619]_ , \new_[50622]_ , \new_[50625]_ , \new_[50626]_ ,
    \new_[50629]_ , \new_[50632]_ , \new_[50633]_ , \new_[50634]_ ,
    \new_[50637]_ , \new_[50640]_ , \new_[50641]_ , \new_[50644]_ ,
    \new_[50647]_ , \new_[50648]_ , \new_[50649]_ , \new_[50652]_ ,
    \new_[50655]_ , \new_[50656]_ , \new_[50659]_ , \new_[50662]_ ,
    \new_[50663]_ , \new_[50664]_ , \new_[50667]_ , \new_[50670]_ ,
    \new_[50671]_ , \new_[50674]_ , \new_[50677]_ , \new_[50678]_ ,
    \new_[50679]_ , \new_[50682]_ , \new_[50685]_ , \new_[50686]_ ,
    \new_[50689]_ , \new_[50692]_ , \new_[50693]_ , \new_[50694]_ ,
    \new_[50697]_ , \new_[50700]_ , \new_[50701]_ , \new_[50704]_ ,
    \new_[50707]_ , \new_[50708]_ , \new_[50709]_ , \new_[50712]_ ,
    \new_[50715]_ , \new_[50716]_ , \new_[50719]_ , \new_[50722]_ ,
    \new_[50723]_ , \new_[50724]_ , \new_[50727]_ , \new_[50730]_ ,
    \new_[50731]_ , \new_[50734]_ , \new_[50737]_ , \new_[50738]_ ,
    \new_[50739]_ , \new_[50742]_ , \new_[50745]_ , \new_[50746]_ ,
    \new_[50749]_ , \new_[50752]_ , \new_[50753]_ , \new_[50754]_ ,
    \new_[50757]_ , \new_[50760]_ , \new_[50761]_ , \new_[50764]_ ,
    \new_[50767]_ , \new_[50768]_ , \new_[50769]_ , \new_[50772]_ ,
    \new_[50775]_ , \new_[50776]_ , \new_[50779]_ , \new_[50782]_ ,
    \new_[50783]_ , \new_[50784]_ , \new_[50787]_ , \new_[50790]_ ,
    \new_[50791]_ , \new_[50794]_ , \new_[50797]_ , \new_[50798]_ ,
    \new_[50799]_ , \new_[50802]_ , \new_[50805]_ , \new_[50806]_ ,
    \new_[50809]_ , \new_[50812]_ , \new_[50813]_ , \new_[50814]_ ,
    \new_[50817]_ , \new_[50820]_ , \new_[50821]_ , \new_[50824]_ ,
    \new_[50827]_ , \new_[50828]_ , \new_[50829]_ , \new_[50832]_ ,
    \new_[50835]_ , \new_[50836]_ , \new_[50839]_ , \new_[50842]_ ,
    \new_[50843]_ , \new_[50844]_ , \new_[50847]_ , \new_[50850]_ ,
    \new_[50851]_ , \new_[50854]_ , \new_[50857]_ , \new_[50858]_ ,
    \new_[50859]_ , \new_[50862]_ , \new_[50865]_ , \new_[50866]_ ,
    \new_[50869]_ , \new_[50872]_ , \new_[50873]_ , \new_[50874]_ ,
    \new_[50877]_ , \new_[50880]_ , \new_[50881]_ , \new_[50884]_ ,
    \new_[50887]_ , \new_[50888]_ , \new_[50889]_ , \new_[50892]_ ,
    \new_[50895]_ , \new_[50896]_ , \new_[50899]_ , \new_[50902]_ ,
    \new_[50903]_ , \new_[50904]_ , \new_[50907]_ , \new_[50910]_ ,
    \new_[50911]_ , \new_[50914]_ , \new_[50917]_ , \new_[50918]_ ,
    \new_[50919]_ , \new_[50922]_ , \new_[50925]_ , \new_[50926]_ ,
    \new_[50929]_ , \new_[50932]_ , \new_[50933]_ , \new_[50934]_ ,
    \new_[50937]_ , \new_[50940]_ , \new_[50941]_ , \new_[50944]_ ,
    \new_[50947]_ , \new_[50948]_ , \new_[50949]_ , \new_[50952]_ ,
    \new_[50955]_ , \new_[50956]_ , \new_[50959]_ , \new_[50962]_ ,
    \new_[50963]_ , \new_[50964]_ , \new_[50967]_ , \new_[50970]_ ,
    \new_[50971]_ , \new_[50974]_ , \new_[50977]_ , \new_[50978]_ ,
    \new_[50979]_ , \new_[50982]_ , \new_[50985]_ , \new_[50986]_ ,
    \new_[50989]_ , \new_[50992]_ , \new_[50993]_ , \new_[50994]_ ,
    \new_[50997]_ , \new_[51000]_ , \new_[51001]_ , \new_[51004]_ ,
    \new_[51007]_ , \new_[51008]_ , \new_[51009]_ , \new_[51012]_ ,
    \new_[51015]_ , \new_[51016]_ , \new_[51019]_ , \new_[51022]_ ,
    \new_[51023]_ , \new_[51024]_ , \new_[51027]_ , \new_[51030]_ ,
    \new_[51031]_ , \new_[51034]_ , \new_[51037]_ , \new_[51038]_ ,
    \new_[51039]_ , \new_[51042]_ , \new_[51045]_ , \new_[51046]_ ,
    \new_[51049]_ , \new_[51052]_ , \new_[51053]_ , \new_[51054]_ ,
    \new_[51057]_ , \new_[51060]_ , \new_[51061]_ , \new_[51064]_ ,
    \new_[51067]_ , \new_[51068]_ , \new_[51069]_ , \new_[51072]_ ,
    \new_[51075]_ , \new_[51076]_ , \new_[51079]_ , \new_[51082]_ ,
    \new_[51083]_ , \new_[51084]_ , \new_[51087]_ , \new_[51090]_ ,
    \new_[51091]_ , \new_[51094]_ , \new_[51097]_ , \new_[51098]_ ,
    \new_[51099]_ , \new_[51102]_ , \new_[51105]_ , \new_[51106]_ ,
    \new_[51109]_ , \new_[51112]_ , \new_[51113]_ , \new_[51114]_ ,
    \new_[51117]_ , \new_[51120]_ , \new_[51121]_ , \new_[51124]_ ,
    \new_[51127]_ , \new_[51128]_ , \new_[51129]_ , \new_[51132]_ ,
    \new_[51135]_ , \new_[51136]_ , \new_[51139]_ , \new_[51142]_ ,
    \new_[51143]_ , \new_[51144]_ , \new_[51147]_ , \new_[51150]_ ,
    \new_[51151]_ , \new_[51154]_ , \new_[51157]_ , \new_[51158]_ ,
    \new_[51159]_ , \new_[51162]_ , \new_[51165]_ , \new_[51166]_ ,
    \new_[51169]_ , \new_[51172]_ , \new_[51173]_ , \new_[51174]_ ,
    \new_[51177]_ , \new_[51180]_ , \new_[51181]_ , \new_[51184]_ ,
    \new_[51187]_ , \new_[51188]_ , \new_[51189]_ , \new_[51192]_ ,
    \new_[51195]_ , \new_[51196]_ , \new_[51199]_ , \new_[51202]_ ,
    \new_[51203]_ , \new_[51204]_ , \new_[51207]_ , \new_[51210]_ ,
    \new_[51211]_ , \new_[51214]_ , \new_[51217]_ , \new_[51218]_ ,
    \new_[51219]_ , \new_[51222]_ , \new_[51225]_ , \new_[51226]_ ,
    \new_[51229]_ , \new_[51232]_ , \new_[51233]_ , \new_[51234]_ ,
    \new_[51237]_ , \new_[51240]_ , \new_[51241]_ , \new_[51244]_ ,
    \new_[51247]_ , \new_[51248]_ , \new_[51249]_ , \new_[51252]_ ,
    \new_[51255]_ , \new_[51256]_ , \new_[51259]_ , \new_[51262]_ ,
    \new_[51263]_ , \new_[51264]_ , \new_[51267]_ , \new_[51270]_ ,
    \new_[51271]_ , \new_[51274]_ , \new_[51277]_ , \new_[51278]_ ,
    \new_[51279]_ , \new_[51282]_ , \new_[51285]_ , \new_[51286]_ ,
    \new_[51289]_ , \new_[51292]_ , \new_[51293]_ , \new_[51294]_ ,
    \new_[51297]_ , \new_[51300]_ , \new_[51301]_ , \new_[51304]_ ,
    \new_[51307]_ , \new_[51308]_ , \new_[51309]_ , \new_[51312]_ ,
    \new_[51315]_ , \new_[51316]_ , \new_[51319]_ , \new_[51322]_ ,
    \new_[51323]_ , \new_[51324]_ , \new_[51327]_ , \new_[51330]_ ,
    \new_[51331]_ , \new_[51334]_ , \new_[51337]_ , \new_[51338]_ ,
    \new_[51339]_ , \new_[51342]_ , \new_[51345]_ , \new_[51346]_ ,
    \new_[51349]_ , \new_[51352]_ , \new_[51353]_ , \new_[51354]_ ,
    \new_[51357]_ , \new_[51360]_ , \new_[51361]_ , \new_[51364]_ ,
    \new_[51367]_ , \new_[51368]_ , \new_[51369]_ , \new_[51372]_ ,
    \new_[51375]_ , \new_[51376]_ , \new_[51379]_ , \new_[51382]_ ,
    \new_[51383]_ , \new_[51384]_ , \new_[51387]_ , \new_[51390]_ ,
    \new_[51391]_ , \new_[51394]_ , \new_[51397]_ , \new_[51398]_ ,
    \new_[51399]_ , \new_[51402]_ , \new_[51405]_ , \new_[51406]_ ,
    \new_[51409]_ , \new_[51412]_ , \new_[51413]_ , \new_[51414]_ ,
    \new_[51417]_ , \new_[51420]_ , \new_[51421]_ , \new_[51424]_ ,
    \new_[51427]_ , \new_[51428]_ , \new_[51429]_ , \new_[51432]_ ,
    \new_[51435]_ , \new_[51436]_ , \new_[51439]_ , \new_[51442]_ ,
    \new_[51443]_ , \new_[51444]_ , \new_[51447]_ , \new_[51450]_ ,
    \new_[51451]_ , \new_[51454]_ , \new_[51457]_ , \new_[51458]_ ,
    \new_[51459]_ , \new_[51462]_ , \new_[51465]_ , \new_[51466]_ ,
    \new_[51469]_ , \new_[51472]_ , \new_[51473]_ , \new_[51474]_ ,
    \new_[51477]_ , \new_[51480]_ , \new_[51481]_ , \new_[51484]_ ,
    \new_[51487]_ , \new_[51488]_ , \new_[51489]_ , \new_[51492]_ ,
    \new_[51495]_ , \new_[51496]_ , \new_[51499]_ , \new_[51502]_ ,
    \new_[51503]_ , \new_[51504]_ , \new_[51507]_ , \new_[51510]_ ,
    \new_[51511]_ , \new_[51514]_ , \new_[51517]_ , \new_[51518]_ ,
    \new_[51519]_ , \new_[51522]_ , \new_[51525]_ , \new_[51526]_ ,
    \new_[51529]_ , \new_[51532]_ , \new_[51533]_ , \new_[51534]_ ,
    \new_[51537]_ , \new_[51540]_ , \new_[51541]_ , \new_[51544]_ ,
    \new_[51547]_ , \new_[51548]_ , \new_[51549]_ , \new_[51552]_ ,
    \new_[51555]_ , \new_[51556]_ , \new_[51559]_ , \new_[51562]_ ,
    \new_[51563]_ , \new_[51564]_ , \new_[51567]_ , \new_[51570]_ ,
    \new_[51571]_ , \new_[51574]_ , \new_[51577]_ , \new_[51578]_ ,
    \new_[51579]_ , \new_[51582]_ , \new_[51585]_ , \new_[51586]_ ,
    \new_[51589]_ , \new_[51592]_ , \new_[51593]_ , \new_[51594]_ ,
    \new_[51597]_ , \new_[51600]_ , \new_[51601]_ , \new_[51604]_ ,
    \new_[51607]_ , \new_[51608]_ , \new_[51609]_ , \new_[51612]_ ,
    \new_[51615]_ , \new_[51616]_ , \new_[51619]_ , \new_[51622]_ ,
    \new_[51623]_ , \new_[51624]_ , \new_[51627]_ , \new_[51630]_ ,
    \new_[51631]_ , \new_[51634]_ , \new_[51637]_ , \new_[51638]_ ,
    \new_[51639]_ , \new_[51642]_ , \new_[51645]_ , \new_[51646]_ ,
    \new_[51649]_ , \new_[51652]_ , \new_[51653]_ , \new_[51654]_ ,
    \new_[51657]_ , \new_[51660]_ , \new_[51661]_ , \new_[51664]_ ,
    \new_[51667]_ , \new_[51668]_ , \new_[51669]_ , \new_[51672]_ ,
    \new_[51675]_ , \new_[51676]_ , \new_[51679]_ , \new_[51682]_ ,
    \new_[51683]_ , \new_[51684]_ , \new_[51687]_ , \new_[51690]_ ,
    \new_[51691]_ , \new_[51694]_ , \new_[51697]_ , \new_[51698]_ ,
    \new_[51699]_ , \new_[51702]_ , \new_[51705]_ , \new_[51706]_ ,
    \new_[51709]_ , \new_[51712]_ , \new_[51713]_ , \new_[51714]_ ,
    \new_[51717]_ , \new_[51720]_ , \new_[51721]_ , \new_[51724]_ ,
    \new_[51727]_ , \new_[51728]_ , \new_[51729]_ , \new_[51732]_ ,
    \new_[51735]_ , \new_[51736]_ , \new_[51739]_ , \new_[51742]_ ,
    \new_[51743]_ , \new_[51744]_ , \new_[51747]_ , \new_[51750]_ ,
    \new_[51751]_ , \new_[51754]_ , \new_[51757]_ , \new_[51758]_ ,
    \new_[51759]_ , \new_[51762]_ , \new_[51765]_ , \new_[51766]_ ,
    \new_[51769]_ , \new_[51773]_ , \new_[51774]_ , \new_[51775]_ ,
    \new_[51776]_ , \new_[51779]_ , \new_[51782]_ , \new_[51783]_ ,
    \new_[51786]_ , \new_[51789]_ , \new_[51790]_ , \new_[51791]_ ,
    \new_[51794]_ , \new_[51797]_ , \new_[51798]_ , \new_[51801]_ ,
    \new_[51805]_ , \new_[51806]_ , \new_[51807]_ , \new_[51808]_ ,
    \new_[51811]_ , \new_[51814]_ , \new_[51815]_ , \new_[51818]_ ,
    \new_[51821]_ , \new_[51822]_ , \new_[51823]_ , \new_[51826]_ ,
    \new_[51829]_ , \new_[51830]_ , \new_[51833]_ , \new_[51837]_ ,
    \new_[51838]_ , \new_[51839]_ , \new_[51840]_ , \new_[51843]_ ,
    \new_[51846]_ , \new_[51847]_ , \new_[51850]_ , \new_[51853]_ ,
    \new_[51854]_ , \new_[51855]_ , \new_[51858]_ , \new_[51861]_ ,
    \new_[51862]_ , \new_[51865]_ , \new_[51869]_ , \new_[51870]_ ,
    \new_[51871]_ , \new_[51872]_ , \new_[51875]_ , \new_[51878]_ ,
    \new_[51879]_ , \new_[51882]_ , \new_[51885]_ , \new_[51886]_ ,
    \new_[51887]_ , \new_[51890]_ , \new_[51893]_ , \new_[51894]_ ,
    \new_[51897]_ , \new_[51901]_ , \new_[51902]_ , \new_[51903]_ ,
    \new_[51904]_ , \new_[51907]_ , \new_[51910]_ , \new_[51911]_ ,
    \new_[51914]_ , \new_[51917]_ , \new_[51918]_ , \new_[51919]_ ,
    \new_[51922]_ , \new_[51925]_ , \new_[51926]_ , \new_[51929]_ ,
    \new_[51933]_ , \new_[51934]_ , \new_[51935]_ , \new_[51936]_ ,
    \new_[51939]_ , \new_[51942]_ , \new_[51943]_ , \new_[51946]_ ,
    \new_[51949]_ , \new_[51950]_ , \new_[51951]_ , \new_[51954]_ ,
    \new_[51957]_ , \new_[51958]_ , \new_[51961]_ , \new_[51965]_ ,
    \new_[51966]_ , \new_[51967]_ , \new_[51968]_ , \new_[51971]_ ,
    \new_[51974]_ , \new_[51975]_ , \new_[51978]_ , \new_[51981]_ ,
    \new_[51982]_ , \new_[51983]_ , \new_[51986]_ , \new_[51989]_ ,
    \new_[51990]_ , \new_[51993]_ , \new_[51997]_ , \new_[51998]_ ,
    \new_[51999]_ , \new_[52000]_ , \new_[52003]_ , \new_[52006]_ ,
    \new_[52007]_ , \new_[52010]_ , \new_[52013]_ , \new_[52014]_ ,
    \new_[52015]_ , \new_[52018]_ , \new_[52021]_ , \new_[52022]_ ,
    \new_[52025]_ , \new_[52029]_ , \new_[52030]_ , \new_[52031]_ ,
    \new_[52032]_ , \new_[52035]_ , \new_[52038]_ , \new_[52039]_ ,
    \new_[52042]_ , \new_[52045]_ , \new_[52046]_ , \new_[52047]_ ,
    \new_[52050]_ , \new_[52053]_ , \new_[52054]_ , \new_[52057]_ ,
    \new_[52061]_ , \new_[52062]_ , \new_[52063]_ , \new_[52064]_ ,
    \new_[52067]_ , \new_[52070]_ , \new_[52071]_ , \new_[52074]_ ,
    \new_[52077]_ , \new_[52078]_ , \new_[52079]_ , \new_[52082]_ ,
    \new_[52085]_ , \new_[52086]_ , \new_[52089]_ , \new_[52093]_ ,
    \new_[52094]_ , \new_[52095]_ , \new_[52096]_ , \new_[52099]_ ,
    \new_[52102]_ , \new_[52103]_ , \new_[52106]_ , \new_[52109]_ ,
    \new_[52110]_ , \new_[52111]_ , \new_[52114]_ , \new_[52117]_ ,
    \new_[52118]_ , \new_[52121]_ , \new_[52125]_ , \new_[52126]_ ,
    \new_[52127]_ , \new_[52128]_ , \new_[52131]_ , \new_[52134]_ ,
    \new_[52135]_ , \new_[52138]_ , \new_[52141]_ , \new_[52142]_ ,
    \new_[52143]_ , \new_[52146]_ , \new_[52149]_ , \new_[52150]_ ,
    \new_[52153]_ , \new_[52157]_ , \new_[52158]_ , \new_[52159]_ ,
    \new_[52160]_ , \new_[52163]_ , \new_[52166]_ , \new_[52167]_ ,
    \new_[52170]_ , \new_[52173]_ , \new_[52174]_ , \new_[52175]_ ,
    \new_[52178]_ , \new_[52181]_ , \new_[52182]_ , \new_[52185]_ ,
    \new_[52189]_ , \new_[52190]_ , \new_[52191]_ , \new_[52192]_ ,
    \new_[52195]_ , \new_[52198]_ , \new_[52199]_ , \new_[52202]_ ,
    \new_[52205]_ , \new_[52206]_ , \new_[52207]_ , \new_[52210]_ ,
    \new_[52213]_ , \new_[52214]_ , \new_[52217]_ , \new_[52221]_ ,
    \new_[52222]_ , \new_[52223]_ , \new_[52224]_ , \new_[52227]_ ,
    \new_[52230]_ , \new_[52231]_ , \new_[52234]_ , \new_[52237]_ ,
    \new_[52238]_ , \new_[52239]_ , \new_[52242]_ , \new_[52245]_ ,
    \new_[52246]_ , \new_[52249]_ , \new_[52253]_ , \new_[52254]_ ,
    \new_[52255]_ , \new_[52256]_ , \new_[52259]_ , \new_[52262]_ ,
    \new_[52263]_ , \new_[52266]_ , \new_[52269]_ , \new_[52270]_ ,
    \new_[52271]_ , \new_[52274]_ , \new_[52277]_ , \new_[52278]_ ,
    \new_[52281]_ , \new_[52285]_ , \new_[52286]_ , \new_[52287]_ ,
    \new_[52288]_ , \new_[52291]_ , \new_[52294]_ , \new_[52295]_ ,
    \new_[52298]_ , \new_[52301]_ , \new_[52302]_ , \new_[52303]_ ,
    \new_[52306]_ , \new_[52309]_ , \new_[52310]_ , \new_[52313]_ ,
    \new_[52317]_ , \new_[52318]_ , \new_[52319]_ , \new_[52320]_ ,
    \new_[52323]_ , \new_[52326]_ , \new_[52327]_ , \new_[52330]_ ,
    \new_[52333]_ , \new_[52334]_ , \new_[52335]_ , \new_[52338]_ ,
    \new_[52341]_ , \new_[52342]_ , \new_[52345]_ , \new_[52349]_ ,
    \new_[52350]_ , \new_[52351]_ , \new_[52352]_ , \new_[52355]_ ,
    \new_[52358]_ , \new_[52359]_ , \new_[52362]_ , \new_[52365]_ ,
    \new_[52366]_ , \new_[52367]_ , \new_[52370]_ , \new_[52373]_ ,
    \new_[52374]_ , \new_[52377]_ , \new_[52381]_ , \new_[52382]_ ,
    \new_[52383]_ , \new_[52384]_ , \new_[52387]_ , \new_[52390]_ ,
    \new_[52391]_ , \new_[52394]_ , \new_[52397]_ , \new_[52398]_ ,
    \new_[52399]_ , \new_[52402]_ , \new_[52405]_ , \new_[52406]_ ,
    \new_[52409]_ , \new_[52413]_ , \new_[52414]_ , \new_[52415]_ ,
    \new_[52416]_ , \new_[52419]_ , \new_[52422]_ , \new_[52423]_ ,
    \new_[52426]_ , \new_[52429]_ , \new_[52430]_ , \new_[52431]_ ,
    \new_[52434]_ , \new_[52437]_ , \new_[52438]_ , \new_[52441]_ ,
    \new_[52445]_ , \new_[52446]_ , \new_[52447]_ , \new_[52448]_ ,
    \new_[52451]_ , \new_[52454]_ , \new_[52455]_ , \new_[52458]_ ,
    \new_[52461]_ , \new_[52462]_ , \new_[52463]_ , \new_[52466]_ ,
    \new_[52469]_ , \new_[52470]_ , \new_[52473]_ , \new_[52477]_ ,
    \new_[52478]_ , \new_[52479]_ , \new_[52480]_ , \new_[52483]_ ,
    \new_[52486]_ , \new_[52487]_ , \new_[52490]_ , \new_[52493]_ ,
    \new_[52494]_ , \new_[52495]_ , \new_[52498]_ , \new_[52501]_ ,
    \new_[52502]_ , \new_[52505]_ , \new_[52509]_ , \new_[52510]_ ,
    \new_[52511]_ , \new_[52512]_ , \new_[52515]_ , \new_[52518]_ ,
    \new_[52519]_ , \new_[52522]_ , \new_[52525]_ , \new_[52526]_ ,
    \new_[52527]_ , \new_[52530]_ , \new_[52533]_ , \new_[52534]_ ,
    \new_[52537]_ , \new_[52541]_ , \new_[52542]_ , \new_[52543]_ ,
    \new_[52544]_ , \new_[52547]_ , \new_[52550]_ , \new_[52551]_ ,
    \new_[52554]_ , \new_[52557]_ , \new_[52558]_ , \new_[52559]_ ,
    \new_[52562]_ , \new_[52565]_ , \new_[52566]_ , \new_[52569]_ ,
    \new_[52573]_ , \new_[52574]_ , \new_[52575]_ , \new_[52576]_ ,
    \new_[52579]_ , \new_[52582]_ , \new_[52583]_ , \new_[52586]_ ,
    \new_[52589]_ , \new_[52590]_ , \new_[52591]_ , \new_[52594]_ ,
    \new_[52597]_ , \new_[52598]_ , \new_[52601]_ , \new_[52605]_ ,
    \new_[52606]_ , \new_[52607]_ , \new_[52608]_ , \new_[52611]_ ,
    \new_[52614]_ , \new_[52615]_ , \new_[52618]_ , \new_[52621]_ ,
    \new_[52622]_ , \new_[52623]_ , \new_[52626]_ , \new_[52629]_ ,
    \new_[52630]_ , \new_[52633]_ , \new_[52637]_ , \new_[52638]_ ,
    \new_[52639]_ , \new_[52640]_ , \new_[52643]_ , \new_[52646]_ ,
    \new_[52647]_ , \new_[52650]_ , \new_[52653]_ , \new_[52654]_ ,
    \new_[52655]_ , \new_[52658]_ , \new_[52661]_ , \new_[52662]_ ,
    \new_[52665]_ , \new_[52669]_ , \new_[52670]_ , \new_[52671]_ ,
    \new_[52672]_ , \new_[52675]_ , \new_[52678]_ , \new_[52679]_ ,
    \new_[52682]_ , \new_[52685]_ , \new_[52686]_ , \new_[52687]_ ,
    \new_[52690]_ , \new_[52693]_ , \new_[52694]_ , \new_[52697]_ ,
    \new_[52701]_ , \new_[52702]_ , \new_[52703]_ , \new_[52704]_ ,
    \new_[52707]_ , \new_[52710]_ , \new_[52711]_ , \new_[52714]_ ,
    \new_[52717]_ , \new_[52718]_ , \new_[52719]_ , \new_[52722]_ ,
    \new_[52725]_ , \new_[52726]_ , \new_[52729]_ , \new_[52733]_ ,
    \new_[52734]_ , \new_[52735]_ , \new_[52736]_ , \new_[52739]_ ,
    \new_[52742]_ , \new_[52743]_ , \new_[52746]_ , \new_[52749]_ ,
    \new_[52750]_ , \new_[52751]_ , \new_[52754]_ , \new_[52757]_ ,
    \new_[52758]_ , \new_[52761]_ , \new_[52765]_ , \new_[52766]_ ,
    \new_[52767]_ , \new_[52768]_ , \new_[52771]_ , \new_[52774]_ ,
    \new_[52775]_ , \new_[52778]_ , \new_[52781]_ , \new_[52782]_ ,
    \new_[52783]_ , \new_[52786]_ , \new_[52789]_ , \new_[52790]_ ,
    \new_[52793]_ , \new_[52797]_ , \new_[52798]_ , \new_[52799]_ ,
    \new_[52800]_ , \new_[52803]_ , \new_[52806]_ , \new_[52807]_ ,
    \new_[52810]_ , \new_[52813]_ , \new_[52814]_ , \new_[52815]_ ,
    \new_[52818]_ , \new_[52821]_ , \new_[52822]_ , \new_[52825]_ ,
    \new_[52829]_ , \new_[52830]_ , \new_[52831]_ , \new_[52832]_ ,
    \new_[52835]_ , \new_[52838]_ , \new_[52839]_ , \new_[52842]_ ,
    \new_[52845]_ , \new_[52846]_ , \new_[52847]_ , \new_[52850]_ ,
    \new_[52853]_ , \new_[52854]_ , \new_[52857]_ , \new_[52861]_ ,
    \new_[52862]_ , \new_[52863]_ , \new_[52864]_ , \new_[52867]_ ,
    \new_[52870]_ , \new_[52871]_ , \new_[52874]_ , \new_[52877]_ ,
    \new_[52878]_ , \new_[52879]_ , \new_[52882]_ , \new_[52885]_ ,
    \new_[52886]_ , \new_[52889]_ , \new_[52893]_ , \new_[52894]_ ,
    \new_[52895]_ , \new_[52896]_ , \new_[52899]_ , \new_[52902]_ ,
    \new_[52903]_ , \new_[52906]_ , \new_[52909]_ , \new_[52910]_ ,
    \new_[52911]_ , \new_[52914]_ , \new_[52917]_ , \new_[52918]_ ,
    \new_[52921]_ , \new_[52925]_ , \new_[52926]_ , \new_[52927]_ ,
    \new_[52928]_ , \new_[52931]_ , \new_[52934]_ , \new_[52935]_ ,
    \new_[52938]_ , \new_[52941]_ , \new_[52942]_ , \new_[52943]_ ,
    \new_[52946]_ , \new_[52949]_ , \new_[52950]_ , \new_[52953]_ ,
    \new_[52957]_ , \new_[52958]_ , \new_[52959]_ , \new_[52960]_ ,
    \new_[52963]_ , \new_[52966]_ , \new_[52967]_ , \new_[52970]_ ,
    \new_[52973]_ , \new_[52974]_ , \new_[52975]_ , \new_[52978]_ ,
    \new_[52981]_ , \new_[52982]_ , \new_[52985]_ , \new_[52989]_ ,
    \new_[52990]_ , \new_[52991]_ , \new_[52992]_ , \new_[52995]_ ,
    \new_[52998]_ , \new_[52999]_ , \new_[53002]_ , \new_[53005]_ ,
    \new_[53006]_ , \new_[53007]_ , \new_[53010]_ , \new_[53013]_ ,
    \new_[53014]_ , \new_[53017]_ , \new_[53021]_ , \new_[53022]_ ,
    \new_[53023]_ , \new_[53024]_ , \new_[53027]_ , \new_[53030]_ ,
    \new_[53031]_ , \new_[53034]_ , \new_[53037]_ , \new_[53038]_ ,
    \new_[53039]_ , \new_[53042]_ , \new_[53045]_ , \new_[53046]_ ,
    \new_[53049]_ , \new_[53053]_ , \new_[53054]_ , \new_[53055]_ ,
    \new_[53056]_ , \new_[53059]_ , \new_[53062]_ , \new_[53063]_ ,
    \new_[53066]_ , \new_[53069]_ , \new_[53070]_ , \new_[53071]_ ,
    \new_[53074]_ , \new_[53077]_ , \new_[53078]_ , \new_[53081]_ ,
    \new_[53085]_ , \new_[53086]_ , \new_[53087]_ , \new_[53088]_ ,
    \new_[53091]_ , \new_[53094]_ , \new_[53095]_ , \new_[53098]_ ,
    \new_[53101]_ , \new_[53102]_ , \new_[53103]_ , \new_[53106]_ ,
    \new_[53109]_ , \new_[53110]_ , \new_[53113]_ , \new_[53117]_ ,
    \new_[53118]_ , \new_[53119]_ , \new_[53120]_ , \new_[53123]_ ,
    \new_[53126]_ , \new_[53127]_ , \new_[53130]_ , \new_[53133]_ ,
    \new_[53134]_ , \new_[53135]_ , \new_[53138]_ , \new_[53141]_ ,
    \new_[53142]_ , \new_[53145]_ , \new_[53149]_ , \new_[53150]_ ,
    \new_[53151]_ , \new_[53152]_ , \new_[53155]_ , \new_[53158]_ ,
    \new_[53159]_ , \new_[53162]_ , \new_[53165]_ , \new_[53166]_ ,
    \new_[53167]_ , \new_[53170]_ , \new_[53173]_ , \new_[53174]_ ,
    \new_[53177]_ , \new_[53181]_ , \new_[53182]_ , \new_[53183]_ ,
    \new_[53184]_ , \new_[53187]_ , \new_[53190]_ , \new_[53191]_ ,
    \new_[53194]_ , \new_[53197]_ , \new_[53198]_ , \new_[53199]_ ,
    \new_[53202]_ , \new_[53205]_ , \new_[53206]_ , \new_[53209]_ ,
    \new_[53213]_ , \new_[53214]_ , \new_[53215]_ , \new_[53216]_ ,
    \new_[53219]_ , \new_[53222]_ , \new_[53223]_ , \new_[53226]_ ,
    \new_[53229]_ , \new_[53230]_ , \new_[53231]_ , \new_[53234]_ ,
    \new_[53237]_ , \new_[53238]_ , \new_[53241]_ , \new_[53245]_ ,
    \new_[53246]_ , \new_[53247]_ , \new_[53248]_ , \new_[53251]_ ,
    \new_[53254]_ , \new_[53255]_ , \new_[53258]_ , \new_[53261]_ ,
    \new_[53262]_ , \new_[53263]_ , \new_[53266]_ , \new_[53269]_ ,
    \new_[53270]_ , \new_[53273]_ , \new_[53277]_ , \new_[53278]_ ,
    \new_[53279]_ , \new_[53280]_ , \new_[53283]_ , \new_[53286]_ ,
    \new_[53287]_ , \new_[53290]_ , \new_[53293]_ , \new_[53294]_ ,
    \new_[53295]_ , \new_[53298]_ , \new_[53301]_ , \new_[53302]_ ,
    \new_[53305]_ , \new_[53309]_ , \new_[53310]_ , \new_[53311]_ ,
    \new_[53312]_ , \new_[53315]_ , \new_[53318]_ , \new_[53319]_ ,
    \new_[53322]_ , \new_[53325]_ , \new_[53326]_ , \new_[53327]_ ,
    \new_[53330]_ , \new_[53333]_ , \new_[53334]_ , \new_[53337]_ ,
    \new_[53341]_ , \new_[53342]_ , \new_[53343]_ , \new_[53344]_ ,
    \new_[53347]_ , \new_[53350]_ , \new_[53351]_ , \new_[53354]_ ,
    \new_[53357]_ , \new_[53358]_ , \new_[53359]_ , \new_[53362]_ ,
    \new_[53365]_ , \new_[53366]_ , \new_[53369]_ , \new_[53373]_ ,
    \new_[53374]_ , \new_[53375]_ , \new_[53376]_ , \new_[53379]_ ,
    \new_[53382]_ , \new_[53383]_ , \new_[53386]_ , \new_[53389]_ ,
    \new_[53390]_ , \new_[53391]_ , \new_[53394]_ , \new_[53397]_ ,
    \new_[53398]_ , \new_[53401]_ , \new_[53405]_ , \new_[53406]_ ,
    \new_[53407]_ , \new_[53408]_ , \new_[53411]_ , \new_[53414]_ ,
    \new_[53415]_ , \new_[53418]_ , \new_[53421]_ , \new_[53422]_ ,
    \new_[53423]_ , \new_[53426]_ , \new_[53429]_ , \new_[53430]_ ,
    \new_[53433]_ , \new_[53437]_ , \new_[53438]_ , \new_[53439]_ ,
    \new_[53440]_ , \new_[53443]_ , \new_[53446]_ , \new_[53447]_ ,
    \new_[53450]_ , \new_[53453]_ , \new_[53454]_ , \new_[53455]_ ,
    \new_[53458]_ , \new_[53461]_ , \new_[53462]_ , \new_[53465]_ ,
    \new_[53469]_ , \new_[53470]_ , \new_[53471]_ , \new_[53472]_ ,
    \new_[53475]_ , \new_[53478]_ , \new_[53479]_ , \new_[53482]_ ,
    \new_[53485]_ , \new_[53486]_ , \new_[53487]_ , \new_[53490]_ ,
    \new_[53493]_ , \new_[53494]_ , \new_[53497]_ , \new_[53501]_ ,
    \new_[53502]_ , \new_[53503]_ , \new_[53504]_ , \new_[53507]_ ,
    \new_[53510]_ , \new_[53511]_ , \new_[53514]_ , \new_[53517]_ ,
    \new_[53518]_ , \new_[53519]_ , \new_[53522]_ , \new_[53525]_ ,
    \new_[53526]_ , \new_[53529]_ , \new_[53533]_ , \new_[53534]_ ,
    \new_[53535]_ , \new_[53536]_ , \new_[53539]_ , \new_[53542]_ ,
    \new_[53543]_ , \new_[53546]_ , \new_[53549]_ , \new_[53550]_ ,
    \new_[53551]_ , \new_[53554]_ , \new_[53557]_ , \new_[53558]_ ,
    \new_[53561]_ , \new_[53565]_ , \new_[53566]_ , \new_[53567]_ ,
    \new_[53568]_ , \new_[53571]_ , \new_[53574]_ , \new_[53575]_ ,
    \new_[53578]_ , \new_[53581]_ , \new_[53582]_ , \new_[53583]_ ,
    \new_[53586]_ , \new_[53589]_ , \new_[53590]_ , \new_[53593]_ ,
    \new_[53597]_ , \new_[53598]_ , \new_[53599]_ , \new_[53600]_ ,
    \new_[53603]_ , \new_[53606]_ , \new_[53607]_ , \new_[53610]_ ,
    \new_[53613]_ , \new_[53614]_ , \new_[53615]_ , \new_[53618]_ ,
    \new_[53621]_ , \new_[53622]_ , \new_[53625]_ , \new_[53629]_ ,
    \new_[53630]_ , \new_[53631]_ , \new_[53632]_ , \new_[53635]_ ,
    \new_[53638]_ , \new_[53639]_ , \new_[53642]_ , \new_[53645]_ ,
    \new_[53646]_ , \new_[53647]_ , \new_[53650]_ , \new_[53653]_ ,
    \new_[53654]_ , \new_[53657]_ , \new_[53661]_ , \new_[53662]_ ,
    \new_[53663]_ , \new_[53664]_ , \new_[53667]_ , \new_[53670]_ ,
    \new_[53671]_ , \new_[53674]_ , \new_[53677]_ , \new_[53678]_ ,
    \new_[53679]_ , \new_[53682]_ , \new_[53685]_ , \new_[53686]_ ,
    \new_[53689]_ , \new_[53693]_ , \new_[53694]_ , \new_[53695]_ ,
    \new_[53696]_ , \new_[53699]_ , \new_[53702]_ , \new_[53703]_ ,
    \new_[53706]_ , \new_[53709]_ , \new_[53710]_ , \new_[53711]_ ,
    \new_[53714]_ , \new_[53717]_ , \new_[53718]_ , \new_[53721]_ ,
    \new_[53725]_ , \new_[53726]_ , \new_[53727]_ , \new_[53728]_ ,
    \new_[53731]_ , \new_[53734]_ , \new_[53735]_ , \new_[53738]_ ,
    \new_[53741]_ , \new_[53742]_ , \new_[53743]_ , \new_[53746]_ ,
    \new_[53749]_ , \new_[53750]_ , \new_[53753]_ , \new_[53757]_ ,
    \new_[53758]_ , \new_[53759]_ , \new_[53760]_ , \new_[53763]_ ,
    \new_[53766]_ , \new_[53767]_ , \new_[53770]_ , \new_[53773]_ ,
    \new_[53774]_ , \new_[53775]_ , \new_[53778]_ , \new_[53781]_ ,
    \new_[53782]_ , \new_[53785]_ , \new_[53789]_ , \new_[53790]_ ,
    \new_[53791]_ , \new_[53792]_ , \new_[53795]_ , \new_[53798]_ ,
    \new_[53799]_ , \new_[53802]_ , \new_[53805]_ , \new_[53806]_ ,
    \new_[53807]_ , \new_[53810]_ , \new_[53813]_ , \new_[53814]_ ,
    \new_[53817]_ , \new_[53821]_ , \new_[53822]_ , \new_[53823]_ ,
    \new_[53824]_ , \new_[53827]_ , \new_[53830]_ , \new_[53831]_ ,
    \new_[53834]_ , \new_[53837]_ , \new_[53838]_ , \new_[53839]_ ,
    \new_[53842]_ , \new_[53845]_ , \new_[53846]_ , \new_[53849]_ ,
    \new_[53853]_ , \new_[53854]_ , \new_[53855]_ , \new_[53856]_ ,
    \new_[53859]_ , \new_[53862]_ , \new_[53863]_ , \new_[53866]_ ,
    \new_[53869]_ , \new_[53870]_ , \new_[53871]_ , \new_[53874]_ ,
    \new_[53877]_ , \new_[53878]_ , \new_[53881]_ , \new_[53885]_ ,
    \new_[53886]_ , \new_[53887]_ , \new_[53888]_ , \new_[53891]_ ,
    \new_[53894]_ , \new_[53895]_ , \new_[53898]_ , \new_[53901]_ ,
    \new_[53902]_ , \new_[53903]_ , \new_[53906]_ , \new_[53909]_ ,
    \new_[53910]_ , \new_[53913]_ , \new_[53917]_ , \new_[53918]_ ,
    \new_[53919]_ , \new_[53920]_ , \new_[53923]_ , \new_[53926]_ ,
    \new_[53927]_ , \new_[53930]_ , \new_[53933]_ , \new_[53934]_ ,
    \new_[53935]_ , \new_[53938]_ , \new_[53941]_ , \new_[53942]_ ,
    \new_[53945]_ , \new_[53949]_ , \new_[53950]_ , \new_[53951]_ ,
    \new_[53952]_ , \new_[53955]_ , \new_[53958]_ , \new_[53959]_ ,
    \new_[53962]_ , \new_[53965]_ , \new_[53966]_ , \new_[53967]_ ,
    \new_[53970]_ , \new_[53973]_ , \new_[53974]_ , \new_[53977]_ ,
    \new_[53981]_ , \new_[53982]_ , \new_[53983]_ , \new_[53984]_ ,
    \new_[53987]_ , \new_[53990]_ , \new_[53991]_ , \new_[53994]_ ,
    \new_[53997]_ , \new_[53998]_ , \new_[53999]_ , \new_[54002]_ ,
    \new_[54005]_ , \new_[54006]_ , \new_[54009]_ , \new_[54013]_ ,
    \new_[54014]_ , \new_[54015]_ , \new_[54016]_ , \new_[54019]_ ,
    \new_[54022]_ , \new_[54023]_ , \new_[54026]_ , \new_[54029]_ ,
    \new_[54030]_ , \new_[54031]_ , \new_[54034]_ , \new_[54037]_ ,
    \new_[54038]_ , \new_[54041]_ , \new_[54045]_ , \new_[54046]_ ,
    \new_[54047]_ , \new_[54048]_ , \new_[54051]_ , \new_[54054]_ ,
    \new_[54055]_ , \new_[54058]_ , \new_[54061]_ , \new_[54062]_ ,
    \new_[54063]_ , \new_[54066]_ , \new_[54069]_ , \new_[54070]_ ,
    \new_[54073]_ , \new_[54077]_ , \new_[54078]_ , \new_[54079]_ ,
    \new_[54080]_ , \new_[54083]_ , \new_[54086]_ , \new_[54087]_ ,
    \new_[54090]_ , \new_[54093]_ , \new_[54094]_ , \new_[54095]_ ,
    \new_[54098]_ , \new_[54101]_ , \new_[54102]_ , \new_[54105]_ ,
    \new_[54109]_ , \new_[54110]_ , \new_[54111]_ , \new_[54112]_ ,
    \new_[54115]_ , \new_[54118]_ , \new_[54119]_ , \new_[54122]_ ,
    \new_[54125]_ , \new_[54126]_ , \new_[54127]_ , \new_[54130]_ ,
    \new_[54133]_ , \new_[54134]_ , \new_[54137]_ , \new_[54141]_ ,
    \new_[54142]_ , \new_[54143]_ , \new_[54144]_ , \new_[54147]_ ,
    \new_[54150]_ , \new_[54151]_ , \new_[54154]_ , \new_[54157]_ ,
    \new_[54158]_ , \new_[54159]_ , \new_[54162]_ , \new_[54165]_ ,
    \new_[54166]_ , \new_[54169]_ , \new_[54173]_ , \new_[54174]_ ,
    \new_[54175]_ , \new_[54176]_ , \new_[54179]_ , \new_[54182]_ ,
    \new_[54183]_ , \new_[54186]_ , \new_[54189]_ , \new_[54190]_ ,
    \new_[54191]_ , \new_[54194]_ , \new_[54197]_ , \new_[54198]_ ,
    \new_[54201]_ , \new_[54205]_ , \new_[54206]_ , \new_[54207]_ ,
    \new_[54208]_ , \new_[54211]_ , \new_[54214]_ , \new_[54215]_ ,
    \new_[54218]_ , \new_[54221]_ , \new_[54222]_ , \new_[54223]_ ,
    \new_[54226]_ , \new_[54229]_ , \new_[54230]_ , \new_[54233]_ ,
    \new_[54237]_ , \new_[54238]_ , \new_[54239]_ , \new_[54240]_ ,
    \new_[54243]_ , \new_[54246]_ , \new_[54247]_ , \new_[54250]_ ,
    \new_[54253]_ , \new_[54254]_ , \new_[54255]_ , \new_[54258]_ ,
    \new_[54261]_ , \new_[54262]_ , \new_[54265]_ , \new_[54269]_ ,
    \new_[54270]_ , \new_[54271]_ , \new_[54272]_ , \new_[54275]_ ,
    \new_[54278]_ , \new_[54279]_ , \new_[54282]_ , \new_[54285]_ ,
    \new_[54286]_ , \new_[54287]_ , \new_[54290]_ , \new_[54293]_ ,
    \new_[54294]_ , \new_[54297]_ , \new_[54301]_ , \new_[54302]_ ,
    \new_[54303]_ , \new_[54304]_ , \new_[54307]_ , \new_[54310]_ ,
    \new_[54311]_ , \new_[54314]_ , \new_[54317]_ , \new_[54318]_ ,
    \new_[54319]_ , \new_[54322]_ , \new_[54325]_ , \new_[54326]_ ,
    \new_[54329]_ , \new_[54333]_ , \new_[54334]_ , \new_[54335]_ ,
    \new_[54336]_ , \new_[54339]_ , \new_[54342]_ , \new_[54343]_ ,
    \new_[54346]_ , \new_[54349]_ , \new_[54350]_ , \new_[54351]_ ,
    \new_[54354]_ , \new_[54357]_ , \new_[54358]_ , \new_[54361]_ ,
    \new_[54365]_ , \new_[54366]_ , \new_[54367]_ , \new_[54368]_ ,
    \new_[54371]_ , \new_[54374]_ , \new_[54375]_ , \new_[54378]_ ,
    \new_[54381]_ , \new_[54382]_ , \new_[54383]_ , \new_[54386]_ ,
    \new_[54389]_ , \new_[54390]_ , \new_[54393]_ , \new_[54397]_ ,
    \new_[54398]_ , \new_[54399]_ , \new_[54400]_ , \new_[54403]_ ,
    \new_[54406]_ , \new_[54407]_ , \new_[54410]_ , \new_[54413]_ ,
    \new_[54414]_ , \new_[54415]_ , \new_[54418]_ , \new_[54421]_ ,
    \new_[54422]_ , \new_[54425]_ , \new_[54429]_ , \new_[54430]_ ,
    \new_[54431]_ , \new_[54432]_ , \new_[54435]_ , \new_[54438]_ ,
    \new_[54439]_ , \new_[54442]_ , \new_[54445]_ , \new_[54446]_ ,
    \new_[54447]_ , \new_[54450]_ , \new_[54453]_ , \new_[54454]_ ,
    \new_[54457]_ , \new_[54461]_ , \new_[54462]_ , \new_[54463]_ ,
    \new_[54464]_ , \new_[54467]_ , \new_[54470]_ , \new_[54471]_ ,
    \new_[54474]_ , \new_[54477]_ , \new_[54478]_ , \new_[54479]_ ,
    \new_[54482]_ , \new_[54485]_ , \new_[54486]_ , \new_[54489]_ ,
    \new_[54493]_ , \new_[54494]_ , \new_[54495]_ , \new_[54496]_ ,
    \new_[54499]_ , \new_[54502]_ , \new_[54503]_ , \new_[54506]_ ,
    \new_[54509]_ , \new_[54510]_ , \new_[54511]_ , \new_[54514]_ ,
    \new_[54517]_ , \new_[54518]_ , \new_[54521]_ , \new_[54525]_ ,
    \new_[54526]_ , \new_[54527]_ , \new_[54528]_ , \new_[54531]_ ,
    \new_[54534]_ , \new_[54535]_ , \new_[54538]_ , \new_[54541]_ ,
    \new_[54542]_ , \new_[54543]_ , \new_[54546]_ , \new_[54549]_ ,
    \new_[54550]_ , \new_[54553]_ , \new_[54557]_ , \new_[54558]_ ,
    \new_[54559]_ , \new_[54560]_ , \new_[54563]_ , \new_[54566]_ ,
    \new_[54567]_ , \new_[54570]_ , \new_[54573]_ , \new_[54574]_ ,
    \new_[54575]_ , \new_[54578]_ , \new_[54581]_ , \new_[54582]_ ,
    \new_[54585]_ , \new_[54589]_ , \new_[54590]_ , \new_[54591]_ ,
    \new_[54592]_ , \new_[54595]_ , \new_[54598]_ , \new_[54599]_ ,
    \new_[54602]_ , \new_[54605]_ , \new_[54606]_ , \new_[54607]_ ,
    \new_[54610]_ , \new_[54613]_ , \new_[54614]_ , \new_[54617]_ ,
    \new_[54621]_ , \new_[54622]_ , \new_[54623]_ , \new_[54624]_ ,
    \new_[54627]_ , \new_[54630]_ , \new_[54631]_ , \new_[54634]_ ,
    \new_[54637]_ , \new_[54638]_ , \new_[54639]_ , \new_[54642]_ ,
    \new_[54645]_ , \new_[54646]_ , \new_[54649]_ , \new_[54653]_ ,
    \new_[54654]_ , \new_[54655]_ , \new_[54656]_ , \new_[54659]_ ,
    \new_[54662]_ , \new_[54663]_ , \new_[54666]_ , \new_[54669]_ ,
    \new_[54670]_ , \new_[54671]_ , \new_[54674]_ , \new_[54677]_ ,
    \new_[54678]_ , \new_[54681]_ , \new_[54685]_ , \new_[54686]_ ,
    \new_[54687]_ , \new_[54688]_ , \new_[54691]_ , \new_[54694]_ ,
    \new_[54695]_ , \new_[54698]_ , \new_[54701]_ , \new_[54702]_ ,
    \new_[54703]_ , \new_[54706]_ , \new_[54709]_ , \new_[54710]_ ,
    \new_[54713]_ , \new_[54717]_ , \new_[54718]_ , \new_[54719]_ ,
    \new_[54720]_ , \new_[54723]_ , \new_[54726]_ , \new_[54727]_ ,
    \new_[54730]_ , \new_[54733]_ , \new_[54734]_ , \new_[54735]_ ,
    \new_[54738]_ , \new_[54741]_ , \new_[54742]_ , \new_[54745]_ ,
    \new_[54749]_ , \new_[54750]_ , \new_[54751]_ , \new_[54752]_ ,
    \new_[54755]_ , \new_[54758]_ , \new_[54759]_ , \new_[54762]_ ,
    \new_[54765]_ , \new_[54766]_ , \new_[54767]_ , \new_[54770]_ ,
    \new_[54773]_ , \new_[54774]_ , \new_[54777]_ , \new_[54781]_ ,
    \new_[54782]_ , \new_[54783]_ , \new_[54784]_ , \new_[54787]_ ,
    \new_[54790]_ , \new_[54791]_ , \new_[54794]_ , \new_[54797]_ ,
    \new_[54798]_ , \new_[54799]_ , \new_[54802]_ , \new_[54805]_ ,
    \new_[54806]_ , \new_[54809]_ , \new_[54813]_ , \new_[54814]_ ,
    \new_[54815]_ , \new_[54816]_ , \new_[54819]_ , \new_[54822]_ ,
    \new_[54823]_ , \new_[54826]_ , \new_[54829]_ , \new_[54830]_ ,
    \new_[54831]_ , \new_[54834]_ , \new_[54837]_ , \new_[54838]_ ,
    \new_[54841]_ , \new_[54845]_ , \new_[54846]_ , \new_[54847]_ ,
    \new_[54848]_ , \new_[54851]_ , \new_[54854]_ , \new_[54855]_ ,
    \new_[54858]_ , \new_[54861]_ , \new_[54862]_ , \new_[54863]_ ,
    \new_[54866]_ , \new_[54869]_ , \new_[54870]_ , \new_[54873]_ ,
    \new_[54877]_ , \new_[54878]_ , \new_[54879]_ , \new_[54880]_ ,
    \new_[54883]_ , \new_[54886]_ , \new_[54887]_ , \new_[54890]_ ,
    \new_[54893]_ , \new_[54894]_ , \new_[54895]_ , \new_[54898]_ ,
    \new_[54901]_ , \new_[54902]_ , \new_[54905]_ , \new_[54909]_ ,
    \new_[54910]_ , \new_[54911]_ , \new_[54912]_ , \new_[54915]_ ,
    \new_[54918]_ , \new_[54919]_ , \new_[54922]_ , \new_[54925]_ ,
    \new_[54926]_ , \new_[54927]_ , \new_[54930]_ , \new_[54933]_ ,
    \new_[54934]_ , \new_[54937]_ , \new_[54941]_ , \new_[54942]_ ,
    \new_[54943]_ , \new_[54944]_ , \new_[54947]_ , \new_[54950]_ ,
    \new_[54951]_ , \new_[54954]_ , \new_[54957]_ , \new_[54958]_ ,
    \new_[54959]_ , \new_[54962]_ , \new_[54965]_ , \new_[54966]_ ,
    \new_[54969]_ , \new_[54973]_ , \new_[54974]_ , \new_[54975]_ ,
    \new_[54976]_ , \new_[54979]_ , \new_[54982]_ , \new_[54983]_ ,
    \new_[54986]_ , \new_[54989]_ , \new_[54990]_ , \new_[54991]_ ,
    \new_[54994]_ , \new_[54997]_ , \new_[54998]_ , \new_[55001]_ ,
    \new_[55005]_ , \new_[55006]_ , \new_[55007]_ , \new_[55008]_ ,
    \new_[55011]_ , \new_[55014]_ , \new_[55015]_ , \new_[55018]_ ,
    \new_[55021]_ , \new_[55022]_ , \new_[55023]_ , \new_[55026]_ ,
    \new_[55029]_ , \new_[55030]_ , \new_[55033]_ , \new_[55037]_ ,
    \new_[55038]_ , \new_[55039]_ , \new_[55040]_ , \new_[55043]_ ,
    \new_[55046]_ , \new_[55047]_ , \new_[55050]_ , \new_[55053]_ ,
    \new_[55054]_ , \new_[55055]_ , \new_[55058]_ , \new_[55061]_ ,
    \new_[55062]_ , \new_[55065]_ , \new_[55069]_ , \new_[55070]_ ,
    \new_[55071]_ , \new_[55072]_ , \new_[55075]_ , \new_[55078]_ ,
    \new_[55079]_ , \new_[55082]_ , \new_[55085]_ , \new_[55086]_ ,
    \new_[55087]_ , \new_[55090]_ , \new_[55093]_ , \new_[55094]_ ,
    \new_[55097]_ , \new_[55101]_ , \new_[55102]_ , \new_[55103]_ ,
    \new_[55104]_ , \new_[55107]_ , \new_[55110]_ , \new_[55111]_ ,
    \new_[55114]_ , \new_[55117]_ , \new_[55118]_ , \new_[55119]_ ,
    \new_[55122]_ , \new_[55125]_ , \new_[55126]_ , \new_[55129]_ ,
    \new_[55133]_ , \new_[55134]_ , \new_[55135]_ , \new_[55136]_ ,
    \new_[55139]_ , \new_[55142]_ , \new_[55143]_ , \new_[55146]_ ,
    \new_[55149]_ , \new_[55150]_ , \new_[55151]_ , \new_[55154]_ ,
    \new_[55157]_ , \new_[55158]_ , \new_[55161]_ , \new_[55165]_ ,
    \new_[55166]_ , \new_[55167]_ , \new_[55168]_ , \new_[55171]_ ,
    \new_[55174]_ , \new_[55175]_ , \new_[55178]_ , \new_[55181]_ ,
    \new_[55182]_ , \new_[55183]_ , \new_[55186]_ , \new_[55189]_ ,
    \new_[55190]_ , \new_[55193]_ , \new_[55197]_ , \new_[55198]_ ,
    \new_[55199]_ , \new_[55200]_ , \new_[55203]_ , \new_[55206]_ ,
    \new_[55207]_ , \new_[55210]_ , \new_[55213]_ , \new_[55214]_ ,
    \new_[55215]_ , \new_[55218]_ , \new_[55221]_ , \new_[55222]_ ,
    \new_[55225]_ , \new_[55229]_ , \new_[55230]_ , \new_[55231]_ ,
    \new_[55232]_ , \new_[55235]_ , \new_[55238]_ , \new_[55239]_ ,
    \new_[55242]_ , \new_[55245]_ , \new_[55246]_ , \new_[55247]_ ,
    \new_[55250]_ , \new_[55253]_ , \new_[55254]_ , \new_[55257]_ ,
    \new_[55261]_ , \new_[55262]_ , \new_[55263]_ , \new_[55264]_ ,
    \new_[55267]_ , \new_[55270]_ , \new_[55271]_ , \new_[55274]_ ,
    \new_[55277]_ , \new_[55278]_ , \new_[55279]_ , \new_[55282]_ ,
    \new_[55285]_ , \new_[55286]_ , \new_[55289]_ , \new_[55293]_ ,
    \new_[55294]_ , \new_[55295]_ , \new_[55296]_ , \new_[55299]_ ,
    \new_[55302]_ , \new_[55303]_ , \new_[55306]_ , \new_[55309]_ ,
    \new_[55310]_ , \new_[55311]_ , \new_[55314]_ , \new_[55317]_ ,
    \new_[55318]_ , \new_[55321]_ , \new_[55325]_ , \new_[55326]_ ,
    \new_[55327]_ , \new_[55328]_ , \new_[55331]_ , \new_[55334]_ ,
    \new_[55335]_ , \new_[55338]_ , \new_[55341]_ , \new_[55342]_ ,
    \new_[55343]_ , \new_[55346]_ , \new_[55349]_ , \new_[55350]_ ,
    \new_[55353]_ , \new_[55357]_ , \new_[55358]_ , \new_[55359]_ ,
    \new_[55360]_ , \new_[55363]_ , \new_[55366]_ , \new_[55367]_ ,
    \new_[55370]_ , \new_[55373]_ , \new_[55374]_ , \new_[55375]_ ,
    \new_[55378]_ , \new_[55381]_ , \new_[55382]_ , \new_[55385]_ ,
    \new_[55389]_ , \new_[55390]_ , \new_[55391]_ , \new_[55392]_ ,
    \new_[55395]_ , \new_[55398]_ , \new_[55399]_ , \new_[55402]_ ,
    \new_[55405]_ , \new_[55406]_ , \new_[55407]_ , \new_[55410]_ ,
    \new_[55413]_ , \new_[55414]_ , \new_[55417]_ , \new_[55421]_ ,
    \new_[55422]_ , \new_[55423]_ , \new_[55424]_ , \new_[55427]_ ,
    \new_[55430]_ , \new_[55431]_ , \new_[55434]_ , \new_[55437]_ ,
    \new_[55438]_ , \new_[55439]_ , \new_[55442]_ , \new_[55445]_ ,
    \new_[55446]_ , \new_[55449]_ , \new_[55453]_ , \new_[55454]_ ,
    \new_[55455]_ , \new_[55456]_ , \new_[55459]_ , \new_[55462]_ ,
    \new_[55463]_ , \new_[55466]_ , \new_[55469]_ , \new_[55470]_ ,
    \new_[55471]_ , \new_[55474]_ , \new_[55477]_ , \new_[55478]_ ,
    \new_[55481]_ , \new_[55485]_ , \new_[55486]_ , \new_[55487]_ ,
    \new_[55488]_ , \new_[55491]_ , \new_[55494]_ , \new_[55495]_ ,
    \new_[55498]_ , \new_[55501]_ , \new_[55502]_ , \new_[55503]_ ,
    \new_[55506]_ , \new_[55509]_ , \new_[55510]_ , \new_[55513]_ ,
    \new_[55517]_ , \new_[55518]_ , \new_[55519]_ , \new_[55520]_ ,
    \new_[55523]_ , \new_[55526]_ , \new_[55527]_ , \new_[55530]_ ,
    \new_[55533]_ , \new_[55534]_ , \new_[55535]_ , \new_[55538]_ ,
    \new_[55541]_ , \new_[55542]_ , \new_[55545]_ , \new_[55549]_ ,
    \new_[55550]_ , \new_[55551]_ , \new_[55552]_ , \new_[55555]_ ,
    \new_[55558]_ , \new_[55559]_ , \new_[55562]_ , \new_[55565]_ ,
    \new_[55566]_ , \new_[55567]_ , \new_[55570]_ , \new_[55573]_ ,
    \new_[55574]_ , \new_[55577]_ , \new_[55581]_ , \new_[55582]_ ,
    \new_[55583]_ , \new_[55584]_ , \new_[55587]_ , \new_[55590]_ ,
    \new_[55591]_ , \new_[55594]_ , \new_[55597]_ , \new_[55598]_ ,
    \new_[55599]_ , \new_[55602]_ , \new_[55605]_ , \new_[55606]_ ,
    \new_[55609]_ , \new_[55613]_ , \new_[55614]_ , \new_[55615]_ ,
    \new_[55616]_ , \new_[55619]_ , \new_[55622]_ , \new_[55623]_ ,
    \new_[55626]_ , \new_[55629]_ , \new_[55630]_ , \new_[55631]_ ,
    \new_[55634]_ , \new_[55637]_ , \new_[55638]_ , \new_[55641]_ ,
    \new_[55645]_ , \new_[55646]_ , \new_[55647]_ , \new_[55648]_ ,
    \new_[55651]_ , \new_[55654]_ , \new_[55655]_ , \new_[55658]_ ,
    \new_[55661]_ , \new_[55662]_ , \new_[55663]_ , \new_[55666]_ ,
    \new_[55669]_ , \new_[55670]_ , \new_[55673]_ , \new_[55677]_ ,
    \new_[55678]_ , \new_[55679]_ , \new_[55680]_ , \new_[55683]_ ,
    \new_[55686]_ , \new_[55687]_ , \new_[55690]_ , \new_[55693]_ ,
    \new_[55694]_ , \new_[55695]_ , \new_[55698]_ , \new_[55701]_ ,
    \new_[55702]_ , \new_[55705]_ , \new_[55709]_ , \new_[55710]_ ,
    \new_[55711]_ , \new_[55712]_ , \new_[55715]_ , \new_[55718]_ ,
    \new_[55719]_ , \new_[55722]_ , \new_[55725]_ , \new_[55726]_ ,
    \new_[55727]_ , \new_[55730]_ , \new_[55733]_ , \new_[55734]_ ,
    \new_[55737]_ , \new_[55741]_ , \new_[55742]_ , \new_[55743]_ ,
    \new_[55744]_ , \new_[55747]_ , \new_[55750]_ , \new_[55751]_ ,
    \new_[55754]_ , \new_[55757]_ , \new_[55758]_ , \new_[55759]_ ,
    \new_[55762]_ , \new_[55765]_ , \new_[55766]_ , \new_[55769]_ ,
    \new_[55773]_ , \new_[55774]_ , \new_[55775]_ , \new_[55776]_ ,
    \new_[55779]_ , \new_[55782]_ , \new_[55783]_ , \new_[55786]_ ,
    \new_[55789]_ , \new_[55790]_ , \new_[55791]_ , \new_[55794]_ ,
    \new_[55797]_ , \new_[55798]_ , \new_[55801]_ , \new_[55805]_ ,
    \new_[55806]_ , \new_[55807]_ , \new_[55808]_ , \new_[55811]_ ,
    \new_[55814]_ , \new_[55815]_ , \new_[55818]_ , \new_[55821]_ ,
    \new_[55822]_ , \new_[55823]_ , \new_[55826]_ , \new_[55829]_ ,
    \new_[55830]_ , \new_[55833]_ , \new_[55837]_ , \new_[55838]_ ,
    \new_[55839]_ , \new_[55840]_ , \new_[55843]_ , \new_[55846]_ ,
    \new_[55847]_ , \new_[55850]_ , \new_[55853]_ , \new_[55854]_ ,
    \new_[55855]_ , \new_[55858]_ , \new_[55861]_ , \new_[55862]_ ,
    \new_[55865]_ , \new_[55869]_ , \new_[55870]_ , \new_[55871]_ ,
    \new_[55872]_ , \new_[55875]_ , \new_[55878]_ , \new_[55879]_ ,
    \new_[55882]_ , \new_[55885]_ , \new_[55886]_ , \new_[55887]_ ,
    \new_[55890]_ , \new_[55893]_ , \new_[55894]_ , \new_[55897]_ ,
    \new_[55901]_ , \new_[55902]_ , \new_[55903]_ , \new_[55904]_ ,
    \new_[55907]_ , \new_[55910]_ , \new_[55911]_ , \new_[55914]_ ,
    \new_[55918]_ , \new_[55919]_ , \new_[55920]_ , \new_[55921]_ ,
    \new_[55924]_ , \new_[55927]_ , \new_[55928]_ , \new_[55931]_ ,
    \new_[55935]_ , \new_[55936]_ , \new_[55937]_ , \new_[55938]_ ,
    \new_[55941]_ , \new_[55944]_ , \new_[55945]_ , \new_[55948]_ ,
    \new_[55952]_ , \new_[55953]_ , \new_[55954]_ , \new_[55955]_ ,
    \new_[55958]_ , \new_[55961]_ , \new_[55962]_ , \new_[55965]_ ,
    \new_[55969]_ , \new_[55970]_ , \new_[55971]_ , \new_[55972]_ ,
    \new_[55975]_ , \new_[55978]_ , \new_[55979]_ , \new_[55982]_ ,
    \new_[55986]_ , \new_[55987]_ , \new_[55988]_ , \new_[55989]_ ,
    \new_[55992]_ , \new_[55995]_ , \new_[55996]_ , \new_[55999]_ ,
    \new_[56003]_ , \new_[56004]_ , \new_[56005]_ , \new_[56006]_ ,
    \new_[56009]_ , \new_[56012]_ , \new_[56013]_ , \new_[56016]_ ,
    \new_[56020]_ , \new_[56021]_ , \new_[56022]_ , \new_[56023]_ ,
    \new_[56026]_ , \new_[56029]_ , \new_[56030]_ , \new_[56033]_ ,
    \new_[56037]_ , \new_[56038]_ , \new_[56039]_ , \new_[56040]_ ,
    \new_[56043]_ , \new_[56046]_ , \new_[56047]_ , \new_[56050]_ ,
    \new_[56054]_ , \new_[56055]_ , \new_[56056]_ , \new_[56057]_ ,
    \new_[56060]_ , \new_[56063]_ , \new_[56064]_ , \new_[56067]_ ,
    \new_[56071]_ , \new_[56072]_ , \new_[56073]_ , \new_[56074]_ ,
    \new_[56077]_ , \new_[56080]_ , \new_[56081]_ , \new_[56084]_ ,
    \new_[56088]_ , \new_[56089]_ , \new_[56090]_ , \new_[56091]_ ,
    \new_[56094]_ , \new_[56097]_ , \new_[56098]_ , \new_[56101]_ ,
    \new_[56105]_ , \new_[56106]_ , \new_[56107]_ , \new_[56108]_ ,
    \new_[56111]_ , \new_[56114]_ , \new_[56115]_ , \new_[56118]_ ,
    \new_[56122]_ , \new_[56123]_ , \new_[56124]_ , \new_[56125]_ ,
    \new_[56128]_ , \new_[56131]_ , \new_[56132]_ , \new_[56135]_ ,
    \new_[56139]_ , \new_[56140]_ , \new_[56141]_ , \new_[56142]_ ,
    \new_[56145]_ , \new_[56148]_ , \new_[56149]_ , \new_[56152]_ ,
    \new_[56156]_ , \new_[56157]_ , \new_[56158]_ , \new_[56159]_ ,
    \new_[56162]_ , \new_[56165]_ , \new_[56166]_ , \new_[56169]_ ,
    \new_[56173]_ , \new_[56174]_ , \new_[56175]_ , \new_[56176]_ ,
    \new_[56179]_ , \new_[56182]_ , \new_[56183]_ , \new_[56186]_ ,
    \new_[56190]_ , \new_[56191]_ , \new_[56192]_ , \new_[56193]_ ,
    \new_[56196]_ , \new_[56199]_ , \new_[56200]_ , \new_[56203]_ ,
    \new_[56207]_ , \new_[56208]_ , \new_[56209]_ , \new_[56210]_ ,
    \new_[56213]_ , \new_[56216]_ , \new_[56217]_ , \new_[56220]_ ,
    \new_[56224]_ , \new_[56225]_ , \new_[56226]_ , \new_[56227]_ ,
    \new_[56230]_ , \new_[56233]_ , \new_[56234]_ , \new_[56237]_ ,
    \new_[56241]_ , \new_[56242]_ , \new_[56243]_ , \new_[56244]_ ,
    \new_[56247]_ , \new_[56250]_ , \new_[56251]_ , \new_[56254]_ ,
    \new_[56258]_ , \new_[56259]_ , \new_[56260]_ , \new_[56261]_ ,
    \new_[56264]_ , \new_[56267]_ , \new_[56268]_ , \new_[56271]_ ,
    \new_[56275]_ , \new_[56276]_ , \new_[56277]_ , \new_[56278]_ ,
    \new_[56281]_ , \new_[56284]_ , \new_[56285]_ , \new_[56288]_ ,
    \new_[56292]_ , \new_[56293]_ , \new_[56294]_ , \new_[56295]_ ,
    \new_[56298]_ , \new_[56301]_ , \new_[56302]_ , \new_[56305]_ ,
    \new_[56309]_ , \new_[56310]_ , \new_[56311]_ , \new_[56312]_ ,
    \new_[56315]_ , \new_[56318]_ , \new_[56319]_ , \new_[56322]_ ,
    \new_[56326]_ , \new_[56327]_ , \new_[56328]_ , \new_[56329]_ ,
    \new_[56332]_ , \new_[56335]_ , \new_[56336]_ , \new_[56339]_ ,
    \new_[56343]_ , \new_[56344]_ , \new_[56345]_ , \new_[56346]_ ,
    \new_[56349]_ , \new_[56352]_ , \new_[56353]_ , \new_[56356]_ ,
    \new_[56360]_ , \new_[56361]_ , \new_[56362]_ , \new_[56363]_ ,
    \new_[56366]_ , \new_[56369]_ , \new_[56370]_ , \new_[56373]_ ,
    \new_[56377]_ , \new_[56378]_ , \new_[56379]_ , \new_[56380]_ ,
    \new_[56383]_ , \new_[56386]_ , \new_[56387]_ , \new_[56390]_ ,
    \new_[56394]_ , \new_[56395]_ , \new_[56396]_ , \new_[56397]_ ,
    \new_[56400]_ , \new_[56403]_ , \new_[56404]_ , \new_[56407]_ ,
    \new_[56411]_ , \new_[56412]_ , \new_[56413]_ , \new_[56414]_ ,
    \new_[56417]_ , \new_[56420]_ , \new_[56421]_ , \new_[56424]_ ,
    \new_[56428]_ , \new_[56429]_ , \new_[56430]_ , \new_[56431]_ ,
    \new_[56434]_ , \new_[56437]_ , \new_[56438]_ , \new_[56441]_ ,
    \new_[56445]_ , \new_[56446]_ , \new_[56447]_ , \new_[56448]_ ,
    \new_[56451]_ , \new_[56454]_ , \new_[56455]_ , \new_[56458]_ ,
    \new_[56462]_ , \new_[56463]_ , \new_[56464]_ , \new_[56465]_ ,
    \new_[56468]_ , \new_[56471]_ , \new_[56472]_ , \new_[56475]_ ,
    \new_[56479]_ , \new_[56480]_ , \new_[56481]_ , \new_[56482]_ ,
    \new_[56485]_ , \new_[56488]_ , \new_[56489]_ , \new_[56492]_ ,
    \new_[56496]_ , \new_[56497]_ , \new_[56498]_ , \new_[56499]_ ,
    \new_[56502]_ , \new_[56505]_ , \new_[56506]_ , \new_[56509]_ ,
    \new_[56513]_ , \new_[56514]_ , \new_[56515]_ , \new_[56516]_ ,
    \new_[56519]_ , \new_[56522]_ , \new_[56523]_ , \new_[56526]_ ,
    \new_[56530]_ , \new_[56531]_ , \new_[56532]_ , \new_[56533]_ ,
    \new_[56536]_ , \new_[56539]_ , \new_[56540]_ , \new_[56543]_ ,
    \new_[56547]_ , \new_[56548]_ , \new_[56549]_ , \new_[56550]_ ,
    \new_[56553]_ , \new_[56556]_ , \new_[56557]_ , \new_[56560]_ ,
    \new_[56564]_ , \new_[56565]_ , \new_[56566]_ , \new_[56567]_ ,
    \new_[56570]_ , \new_[56573]_ , \new_[56574]_ , \new_[56577]_ ,
    \new_[56581]_ , \new_[56582]_ , \new_[56583]_ , \new_[56584]_ ,
    \new_[56587]_ , \new_[56590]_ , \new_[56591]_ , \new_[56594]_ ,
    \new_[56598]_ , \new_[56599]_ , \new_[56600]_ , \new_[56601]_ ,
    \new_[56604]_ , \new_[56607]_ , \new_[56608]_ , \new_[56611]_ ,
    \new_[56615]_ , \new_[56616]_ , \new_[56617]_ , \new_[56618]_ ,
    \new_[56621]_ , \new_[56624]_ , \new_[56625]_ , \new_[56628]_ ,
    \new_[56632]_ , \new_[56633]_ , \new_[56634]_ , \new_[56635]_ ,
    \new_[56638]_ , \new_[56641]_ , \new_[56642]_ , \new_[56645]_ ,
    \new_[56649]_ , \new_[56650]_ , \new_[56651]_ , \new_[56652]_ ,
    \new_[56655]_ , \new_[56658]_ , \new_[56659]_ , \new_[56662]_ ,
    \new_[56666]_ , \new_[56667]_ , \new_[56668]_ , \new_[56669]_ ,
    \new_[56672]_ , \new_[56675]_ , \new_[56676]_ , \new_[56679]_ ,
    \new_[56683]_ , \new_[56684]_ , \new_[56685]_ , \new_[56686]_ ,
    \new_[56689]_ , \new_[56692]_ , \new_[56693]_ , \new_[56696]_ ,
    \new_[56700]_ , \new_[56701]_ , \new_[56702]_ , \new_[56703]_ ,
    \new_[56706]_ , \new_[56709]_ , \new_[56710]_ , \new_[56713]_ ,
    \new_[56717]_ , \new_[56718]_ , \new_[56719]_ , \new_[56720]_ ,
    \new_[56723]_ , \new_[56726]_ , \new_[56727]_ , \new_[56730]_ ,
    \new_[56734]_ , \new_[56735]_ , \new_[56736]_ , \new_[56737]_ ,
    \new_[56740]_ , \new_[56743]_ , \new_[56744]_ , \new_[56747]_ ,
    \new_[56751]_ , \new_[56752]_ , \new_[56753]_ , \new_[56754]_ ,
    \new_[56757]_ , \new_[56760]_ , \new_[56761]_ , \new_[56764]_ ,
    \new_[56768]_ , \new_[56769]_ , \new_[56770]_ , \new_[56771]_ ,
    \new_[56774]_ , \new_[56777]_ , \new_[56778]_ , \new_[56781]_ ,
    \new_[56785]_ , \new_[56786]_ , \new_[56787]_ , \new_[56788]_ ,
    \new_[56791]_ , \new_[56794]_ , \new_[56795]_ , \new_[56798]_ ,
    \new_[56802]_ , \new_[56803]_ , \new_[56804]_ , \new_[56805]_ ,
    \new_[56808]_ , \new_[56811]_ , \new_[56812]_ , \new_[56815]_ ,
    \new_[56819]_ , \new_[56820]_ , \new_[56821]_ , \new_[56822]_ ,
    \new_[56825]_ , \new_[56828]_ , \new_[56829]_ , \new_[56832]_ ,
    \new_[56836]_ , \new_[56837]_ , \new_[56838]_ , \new_[56839]_ ,
    \new_[56842]_ , \new_[56845]_ , \new_[56846]_ , \new_[56849]_ ,
    \new_[56853]_ , \new_[56854]_ , \new_[56855]_ , \new_[56856]_ ,
    \new_[56859]_ , \new_[56862]_ , \new_[56863]_ , \new_[56866]_ ,
    \new_[56870]_ , \new_[56871]_ , \new_[56872]_ , \new_[56873]_ ,
    \new_[56876]_ , \new_[56879]_ , \new_[56880]_ , \new_[56883]_ ,
    \new_[56887]_ , \new_[56888]_ , \new_[56889]_ , \new_[56890]_ ,
    \new_[56893]_ , \new_[56896]_ , \new_[56897]_ , \new_[56900]_ ,
    \new_[56904]_ , \new_[56905]_ , \new_[56906]_ , \new_[56907]_ ,
    \new_[56910]_ , \new_[56913]_ , \new_[56914]_ , \new_[56917]_ ,
    \new_[56921]_ , \new_[56922]_ , \new_[56923]_ , \new_[56924]_ ,
    \new_[56927]_ , \new_[56930]_ , \new_[56931]_ , \new_[56934]_ ,
    \new_[56938]_ , \new_[56939]_ , \new_[56940]_ , \new_[56941]_ ,
    \new_[56944]_ , \new_[56947]_ , \new_[56948]_ , \new_[56951]_ ,
    \new_[56955]_ , \new_[56956]_ , \new_[56957]_ , \new_[56958]_ ,
    \new_[56961]_ , \new_[56964]_ , \new_[56965]_ , \new_[56968]_ ,
    \new_[56972]_ , \new_[56973]_ , \new_[56974]_ , \new_[56975]_ ,
    \new_[56978]_ , \new_[56981]_ , \new_[56982]_ , \new_[56985]_ ,
    \new_[56989]_ , \new_[56990]_ , \new_[56991]_ , \new_[56992]_ ,
    \new_[56995]_ , \new_[56998]_ , \new_[56999]_ , \new_[57002]_ ,
    \new_[57006]_ , \new_[57007]_ , \new_[57008]_ , \new_[57009]_ ,
    \new_[57012]_ , \new_[57015]_ , \new_[57016]_ , \new_[57019]_ ,
    \new_[57023]_ , \new_[57024]_ , \new_[57025]_ , \new_[57026]_ ,
    \new_[57029]_ , \new_[57032]_ , \new_[57033]_ , \new_[57036]_ ,
    \new_[57040]_ , \new_[57041]_ , \new_[57042]_ , \new_[57043]_ ,
    \new_[57046]_ , \new_[57049]_ , \new_[57050]_ , \new_[57053]_ ,
    \new_[57057]_ , \new_[57058]_ , \new_[57059]_ , \new_[57060]_ ,
    \new_[57063]_ , \new_[57066]_ , \new_[57067]_ , \new_[57070]_ ,
    \new_[57074]_ , \new_[57075]_ , \new_[57076]_ , \new_[57077]_ ,
    \new_[57080]_ , \new_[57083]_ , \new_[57084]_ , \new_[57087]_ ,
    \new_[57091]_ , \new_[57092]_ , \new_[57093]_ , \new_[57094]_ ,
    \new_[57097]_ , \new_[57100]_ , \new_[57101]_ , \new_[57104]_ ,
    \new_[57108]_ , \new_[57109]_ , \new_[57110]_ , \new_[57111]_ ,
    \new_[57114]_ , \new_[57117]_ , \new_[57118]_ , \new_[57121]_ ,
    \new_[57125]_ , \new_[57126]_ , \new_[57127]_ , \new_[57128]_ ,
    \new_[57131]_ , \new_[57134]_ , \new_[57135]_ , \new_[57138]_ ,
    \new_[57142]_ , \new_[57143]_ , \new_[57144]_ , \new_[57145]_ ,
    \new_[57148]_ , \new_[57152]_ , \new_[57153]_ , \new_[57154]_ ,
    \new_[57157]_ , \new_[57161]_ , \new_[57162]_ , \new_[57163]_ ,
    \new_[57164]_ , \new_[57167]_ , \new_[57170]_ , \new_[57171]_ ,
    \new_[57174]_ , \new_[57178]_ , \new_[57179]_ , \new_[57180]_ ,
    \new_[57181]_ , \new_[57184]_ , \new_[57188]_ , \new_[57189]_ ,
    \new_[57190]_ , \new_[57193]_ , \new_[57197]_ , \new_[57198]_ ,
    \new_[57199]_ , \new_[57200]_ , \new_[57203]_ , \new_[57206]_ ,
    \new_[57207]_ , \new_[57210]_ , \new_[57214]_ , \new_[57215]_ ,
    \new_[57216]_ , \new_[57217]_ , \new_[57220]_ , \new_[57224]_ ,
    \new_[57225]_ , \new_[57226]_ , \new_[57229]_ , \new_[57233]_ ,
    \new_[57234]_ , \new_[57235]_ , \new_[57236]_ , \new_[57239]_ ,
    \new_[57242]_ , \new_[57243]_ , \new_[57246]_ , \new_[57250]_ ,
    \new_[57251]_ , \new_[57252]_ , \new_[57253]_ , \new_[57256]_ ,
    \new_[57260]_ , \new_[57261]_ , \new_[57262]_ , \new_[57265]_ ,
    \new_[57269]_ , \new_[57270]_ , \new_[57271]_ , \new_[57272]_ ;
  assign A76 = \new_[6928]_  | \new_[4619]_ ;
  assign \new_[1]_  = \new_[57272]_  & \new_[57253]_ ;
  assign \new_[2]_  = \new_[57236]_  & \new_[57217]_ ;
  assign \new_[3]_  = \new_[57200]_  & \new_[57181]_ ;
  assign \new_[4]_  = \new_[57164]_  & \new_[57145]_ ;
  assign \new_[5]_  = \new_[57128]_  & \new_[57111]_ ;
  assign \new_[6]_  = \new_[57094]_  & \new_[57077]_ ;
  assign \new_[7]_  = \new_[57060]_  & \new_[57043]_ ;
  assign \new_[8]_  = \new_[57026]_  & \new_[57009]_ ;
  assign \new_[9]_  = \new_[56992]_  & \new_[56975]_ ;
  assign \new_[10]_  = \new_[56958]_  & \new_[56941]_ ;
  assign \new_[11]_  = \new_[56924]_  & \new_[56907]_ ;
  assign \new_[12]_  = \new_[56890]_  & \new_[56873]_ ;
  assign \new_[13]_  = \new_[56856]_  & \new_[56839]_ ;
  assign \new_[14]_  = \new_[56822]_  & \new_[56805]_ ;
  assign \new_[15]_  = \new_[56788]_  & \new_[56771]_ ;
  assign \new_[16]_  = \new_[56754]_  & \new_[56737]_ ;
  assign \new_[17]_  = \new_[56720]_  & \new_[56703]_ ;
  assign \new_[18]_  = \new_[56686]_  & \new_[56669]_ ;
  assign \new_[19]_  = \new_[56652]_  & \new_[56635]_ ;
  assign \new_[20]_  = \new_[56618]_  & \new_[56601]_ ;
  assign \new_[21]_  = \new_[56584]_  & \new_[56567]_ ;
  assign \new_[22]_  = \new_[56550]_  & \new_[56533]_ ;
  assign \new_[23]_  = \new_[56516]_  & \new_[56499]_ ;
  assign \new_[24]_  = \new_[56482]_  & \new_[56465]_ ;
  assign \new_[25]_  = \new_[56448]_  & \new_[56431]_ ;
  assign \new_[26]_  = \new_[56414]_  & \new_[56397]_ ;
  assign \new_[27]_  = \new_[56380]_  & \new_[56363]_ ;
  assign \new_[28]_  = \new_[56346]_  & \new_[56329]_ ;
  assign \new_[29]_  = \new_[56312]_  & \new_[56295]_ ;
  assign \new_[30]_  = \new_[56278]_  & \new_[56261]_ ;
  assign \new_[31]_  = \new_[56244]_  & \new_[56227]_ ;
  assign \new_[32]_  = \new_[56210]_  & \new_[56193]_ ;
  assign \new_[33]_  = \new_[56176]_  & \new_[56159]_ ;
  assign \new_[34]_  = \new_[56142]_  & \new_[56125]_ ;
  assign \new_[35]_  = \new_[56108]_  & \new_[56091]_ ;
  assign \new_[36]_  = \new_[56074]_  & \new_[56057]_ ;
  assign \new_[37]_  = \new_[56040]_  & \new_[56023]_ ;
  assign \new_[38]_  = \new_[56006]_  & \new_[55989]_ ;
  assign \new_[39]_  = \new_[55972]_  & \new_[55955]_ ;
  assign \new_[40]_  = \new_[55938]_  & \new_[55921]_ ;
  assign \new_[41]_  = \new_[55904]_  & \new_[55887]_ ;
  assign \new_[42]_  = \new_[55872]_  & \new_[55855]_ ;
  assign \new_[43]_  = \new_[55840]_  & \new_[55823]_ ;
  assign \new_[44]_  = \new_[55808]_  & \new_[55791]_ ;
  assign \new_[45]_  = \new_[55776]_  & \new_[55759]_ ;
  assign \new_[46]_  = \new_[55744]_  & \new_[55727]_ ;
  assign \new_[47]_  = \new_[55712]_  & \new_[55695]_ ;
  assign \new_[48]_  = \new_[55680]_  & \new_[55663]_ ;
  assign \new_[49]_  = \new_[55648]_  & \new_[55631]_ ;
  assign \new_[50]_  = \new_[55616]_  & \new_[55599]_ ;
  assign \new_[51]_  = \new_[55584]_  & \new_[55567]_ ;
  assign \new_[52]_  = \new_[55552]_  & \new_[55535]_ ;
  assign \new_[53]_  = \new_[55520]_  & \new_[55503]_ ;
  assign \new_[54]_  = \new_[55488]_  & \new_[55471]_ ;
  assign \new_[55]_  = \new_[55456]_  & \new_[55439]_ ;
  assign \new_[56]_  = \new_[55424]_  & \new_[55407]_ ;
  assign \new_[57]_  = \new_[55392]_  & \new_[55375]_ ;
  assign \new_[58]_  = \new_[55360]_  & \new_[55343]_ ;
  assign \new_[59]_  = \new_[55328]_  & \new_[55311]_ ;
  assign \new_[60]_  = \new_[55296]_  & \new_[55279]_ ;
  assign \new_[61]_  = \new_[55264]_  & \new_[55247]_ ;
  assign \new_[62]_  = \new_[55232]_  & \new_[55215]_ ;
  assign \new_[63]_  = \new_[55200]_  & \new_[55183]_ ;
  assign \new_[64]_  = \new_[55168]_  & \new_[55151]_ ;
  assign \new_[65]_  = \new_[55136]_  & \new_[55119]_ ;
  assign \new_[66]_  = \new_[55104]_  & \new_[55087]_ ;
  assign \new_[67]_  = \new_[55072]_  & \new_[55055]_ ;
  assign \new_[68]_  = \new_[55040]_  & \new_[55023]_ ;
  assign \new_[69]_  = \new_[55008]_  & \new_[54991]_ ;
  assign \new_[70]_  = \new_[54976]_  & \new_[54959]_ ;
  assign \new_[71]_  = \new_[54944]_  & \new_[54927]_ ;
  assign \new_[72]_  = \new_[54912]_  & \new_[54895]_ ;
  assign \new_[73]_  = \new_[54880]_  & \new_[54863]_ ;
  assign \new_[74]_  = \new_[54848]_  & \new_[54831]_ ;
  assign \new_[75]_  = \new_[54816]_  & \new_[54799]_ ;
  assign \new_[76]_  = \new_[54784]_  & \new_[54767]_ ;
  assign \new_[77]_  = \new_[54752]_  & \new_[54735]_ ;
  assign \new_[78]_  = \new_[54720]_  & \new_[54703]_ ;
  assign \new_[79]_  = \new_[54688]_  & \new_[54671]_ ;
  assign \new_[80]_  = \new_[54656]_  & \new_[54639]_ ;
  assign \new_[81]_  = \new_[54624]_  & \new_[54607]_ ;
  assign \new_[82]_  = \new_[54592]_  & \new_[54575]_ ;
  assign \new_[83]_  = \new_[54560]_  & \new_[54543]_ ;
  assign \new_[84]_  = \new_[54528]_  & \new_[54511]_ ;
  assign \new_[85]_  = \new_[54496]_  & \new_[54479]_ ;
  assign \new_[86]_  = \new_[54464]_  & \new_[54447]_ ;
  assign \new_[87]_  = \new_[54432]_  & \new_[54415]_ ;
  assign \new_[88]_  = \new_[54400]_  & \new_[54383]_ ;
  assign \new_[89]_  = \new_[54368]_  & \new_[54351]_ ;
  assign \new_[90]_  = \new_[54336]_  & \new_[54319]_ ;
  assign \new_[91]_  = \new_[54304]_  & \new_[54287]_ ;
  assign \new_[92]_  = \new_[54272]_  & \new_[54255]_ ;
  assign \new_[93]_  = \new_[54240]_  & \new_[54223]_ ;
  assign \new_[94]_  = \new_[54208]_  & \new_[54191]_ ;
  assign \new_[95]_  = \new_[54176]_  & \new_[54159]_ ;
  assign \new_[96]_  = \new_[54144]_  & \new_[54127]_ ;
  assign \new_[97]_  = \new_[54112]_  & \new_[54095]_ ;
  assign \new_[98]_  = \new_[54080]_  & \new_[54063]_ ;
  assign \new_[99]_  = \new_[54048]_  & \new_[54031]_ ;
  assign \new_[100]_  = \new_[54016]_  & \new_[53999]_ ;
  assign \new_[101]_  = \new_[53984]_  & \new_[53967]_ ;
  assign \new_[102]_  = \new_[53952]_  & \new_[53935]_ ;
  assign \new_[103]_  = \new_[53920]_  & \new_[53903]_ ;
  assign \new_[104]_  = \new_[53888]_  & \new_[53871]_ ;
  assign \new_[105]_  = \new_[53856]_  & \new_[53839]_ ;
  assign \new_[106]_  = \new_[53824]_  & \new_[53807]_ ;
  assign \new_[107]_  = \new_[53792]_  & \new_[53775]_ ;
  assign \new_[108]_  = \new_[53760]_  & \new_[53743]_ ;
  assign \new_[109]_  = \new_[53728]_  & \new_[53711]_ ;
  assign \new_[110]_  = \new_[53696]_  & \new_[53679]_ ;
  assign \new_[111]_  = \new_[53664]_  & \new_[53647]_ ;
  assign \new_[112]_  = \new_[53632]_  & \new_[53615]_ ;
  assign \new_[113]_  = \new_[53600]_  & \new_[53583]_ ;
  assign \new_[114]_  = \new_[53568]_  & \new_[53551]_ ;
  assign \new_[115]_  = \new_[53536]_  & \new_[53519]_ ;
  assign \new_[116]_  = \new_[53504]_  & \new_[53487]_ ;
  assign \new_[117]_  = \new_[53472]_  & \new_[53455]_ ;
  assign \new_[118]_  = \new_[53440]_  & \new_[53423]_ ;
  assign \new_[119]_  = \new_[53408]_  & \new_[53391]_ ;
  assign \new_[120]_  = \new_[53376]_  & \new_[53359]_ ;
  assign \new_[121]_  = \new_[53344]_  & \new_[53327]_ ;
  assign \new_[122]_  = \new_[53312]_  & \new_[53295]_ ;
  assign \new_[123]_  = \new_[53280]_  & \new_[53263]_ ;
  assign \new_[124]_  = \new_[53248]_  & \new_[53231]_ ;
  assign \new_[125]_  = \new_[53216]_  & \new_[53199]_ ;
  assign \new_[126]_  = \new_[53184]_  & \new_[53167]_ ;
  assign \new_[127]_  = \new_[53152]_  & \new_[53135]_ ;
  assign \new_[128]_  = \new_[53120]_  & \new_[53103]_ ;
  assign \new_[129]_  = \new_[53088]_  & \new_[53071]_ ;
  assign \new_[130]_  = \new_[53056]_  & \new_[53039]_ ;
  assign \new_[131]_  = \new_[53024]_  & \new_[53007]_ ;
  assign \new_[132]_  = \new_[52992]_  & \new_[52975]_ ;
  assign \new_[133]_  = \new_[52960]_  & \new_[52943]_ ;
  assign \new_[134]_  = \new_[52928]_  & \new_[52911]_ ;
  assign \new_[135]_  = \new_[52896]_  & \new_[52879]_ ;
  assign \new_[136]_  = \new_[52864]_  & \new_[52847]_ ;
  assign \new_[137]_  = \new_[52832]_  & \new_[52815]_ ;
  assign \new_[138]_  = \new_[52800]_  & \new_[52783]_ ;
  assign \new_[139]_  = \new_[52768]_  & \new_[52751]_ ;
  assign \new_[140]_  = \new_[52736]_  & \new_[52719]_ ;
  assign \new_[141]_  = \new_[52704]_  & \new_[52687]_ ;
  assign \new_[142]_  = \new_[52672]_  & \new_[52655]_ ;
  assign \new_[143]_  = \new_[52640]_  & \new_[52623]_ ;
  assign \new_[144]_  = \new_[52608]_  & \new_[52591]_ ;
  assign \new_[145]_  = \new_[52576]_  & \new_[52559]_ ;
  assign \new_[146]_  = \new_[52544]_  & \new_[52527]_ ;
  assign \new_[147]_  = \new_[52512]_  & \new_[52495]_ ;
  assign \new_[148]_  = \new_[52480]_  & \new_[52463]_ ;
  assign \new_[149]_  = \new_[52448]_  & \new_[52431]_ ;
  assign \new_[150]_  = \new_[52416]_  & \new_[52399]_ ;
  assign \new_[151]_  = \new_[52384]_  & \new_[52367]_ ;
  assign \new_[152]_  = \new_[52352]_  & \new_[52335]_ ;
  assign \new_[153]_  = \new_[52320]_  & \new_[52303]_ ;
  assign \new_[154]_  = \new_[52288]_  & \new_[52271]_ ;
  assign \new_[155]_  = \new_[52256]_  & \new_[52239]_ ;
  assign \new_[156]_  = \new_[52224]_  & \new_[52207]_ ;
  assign \new_[157]_  = \new_[52192]_  & \new_[52175]_ ;
  assign \new_[158]_  = \new_[52160]_  & \new_[52143]_ ;
  assign \new_[159]_  = \new_[52128]_  & \new_[52111]_ ;
  assign \new_[160]_  = \new_[52096]_  & \new_[52079]_ ;
  assign \new_[161]_  = \new_[52064]_  & \new_[52047]_ ;
  assign \new_[162]_  = \new_[52032]_  & \new_[52015]_ ;
  assign \new_[163]_  = \new_[52000]_  & \new_[51983]_ ;
  assign \new_[164]_  = \new_[51968]_  & \new_[51951]_ ;
  assign \new_[165]_  = \new_[51936]_  & \new_[51919]_ ;
  assign \new_[166]_  = \new_[51904]_  & \new_[51887]_ ;
  assign \new_[167]_  = \new_[51872]_  & \new_[51855]_ ;
  assign \new_[168]_  = \new_[51840]_  & \new_[51823]_ ;
  assign \new_[169]_  = \new_[51808]_  & \new_[51791]_ ;
  assign \new_[170]_  = \new_[51776]_  & \new_[51759]_ ;
  assign \new_[171]_  = \new_[51744]_  & \new_[51729]_ ;
  assign \new_[172]_  = \new_[51714]_  & \new_[51699]_ ;
  assign \new_[173]_  = \new_[51684]_  & \new_[51669]_ ;
  assign \new_[174]_  = \new_[51654]_  & \new_[51639]_ ;
  assign \new_[175]_  = \new_[51624]_  & \new_[51609]_ ;
  assign \new_[176]_  = \new_[51594]_  & \new_[51579]_ ;
  assign \new_[177]_  = \new_[51564]_  & \new_[51549]_ ;
  assign \new_[178]_  = \new_[51534]_  & \new_[51519]_ ;
  assign \new_[179]_  = \new_[51504]_  & \new_[51489]_ ;
  assign \new_[180]_  = \new_[51474]_  & \new_[51459]_ ;
  assign \new_[181]_  = \new_[51444]_  & \new_[51429]_ ;
  assign \new_[182]_  = \new_[51414]_  & \new_[51399]_ ;
  assign \new_[183]_  = \new_[51384]_  & \new_[51369]_ ;
  assign \new_[184]_  = \new_[51354]_  & \new_[51339]_ ;
  assign \new_[185]_  = \new_[51324]_  & \new_[51309]_ ;
  assign \new_[186]_  = \new_[51294]_  & \new_[51279]_ ;
  assign \new_[187]_  = \new_[51264]_  & \new_[51249]_ ;
  assign \new_[188]_  = \new_[51234]_  & \new_[51219]_ ;
  assign \new_[189]_  = \new_[51204]_  & \new_[51189]_ ;
  assign \new_[190]_  = \new_[51174]_  & \new_[51159]_ ;
  assign \new_[191]_  = \new_[51144]_  & \new_[51129]_ ;
  assign \new_[192]_  = \new_[51114]_  & \new_[51099]_ ;
  assign \new_[193]_  = \new_[51084]_  & \new_[51069]_ ;
  assign \new_[194]_  = \new_[51054]_  & \new_[51039]_ ;
  assign \new_[195]_  = \new_[51024]_  & \new_[51009]_ ;
  assign \new_[196]_  = \new_[50994]_  & \new_[50979]_ ;
  assign \new_[197]_  = \new_[50964]_  & \new_[50949]_ ;
  assign \new_[198]_  = \new_[50934]_  & \new_[50919]_ ;
  assign \new_[199]_  = \new_[50904]_  & \new_[50889]_ ;
  assign \new_[200]_  = \new_[50874]_  & \new_[50859]_ ;
  assign \new_[201]_  = \new_[50844]_  & \new_[50829]_ ;
  assign \new_[202]_  = \new_[50814]_  & \new_[50799]_ ;
  assign \new_[203]_  = \new_[50784]_  & \new_[50769]_ ;
  assign \new_[204]_  = \new_[50754]_  & \new_[50739]_ ;
  assign \new_[205]_  = \new_[50724]_  & \new_[50709]_ ;
  assign \new_[206]_  = \new_[50694]_  & \new_[50679]_ ;
  assign \new_[207]_  = \new_[50664]_  & \new_[50649]_ ;
  assign \new_[208]_  = \new_[50634]_  & \new_[50619]_ ;
  assign \new_[209]_  = \new_[50604]_  & \new_[50589]_ ;
  assign \new_[210]_  = \new_[50574]_  & \new_[50559]_ ;
  assign \new_[211]_  = \new_[50544]_  & \new_[50529]_ ;
  assign \new_[212]_  = \new_[50514]_  & \new_[50499]_ ;
  assign \new_[213]_  = \new_[50484]_  & \new_[50469]_ ;
  assign \new_[214]_  = \new_[50454]_  & \new_[50439]_ ;
  assign \new_[215]_  = \new_[50424]_  & \new_[50409]_ ;
  assign \new_[216]_  = \new_[50394]_  & \new_[50379]_ ;
  assign \new_[217]_  = \new_[50364]_  & \new_[50349]_ ;
  assign \new_[218]_  = \new_[50334]_  & \new_[50319]_ ;
  assign \new_[219]_  = \new_[50304]_  & \new_[50289]_ ;
  assign \new_[220]_  = \new_[50274]_  & \new_[50259]_ ;
  assign \new_[221]_  = \new_[50244]_  & \new_[50229]_ ;
  assign \new_[222]_  = \new_[50214]_  & \new_[50199]_ ;
  assign \new_[223]_  = \new_[50184]_  & \new_[50169]_ ;
  assign \new_[224]_  = \new_[50154]_  & \new_[50139]_ ;
  assign \new_[225]_  = \new_[50124]_  & \new_[50109]_ ;
  assign \new_[226]_  = \new_[50094]_  & \new_[50079]_ ;
  assign \new_[227]_  = \new_[50064]_  & \new_[50049]_ ;
  assign \new_[228]_  = \new_[50034]_  & \new_[50019]_ ;
  assign \new_[229]_  = \new_[50004]_  & \new_[49989]_ ;
  assign \new_[230]_  = \new_[49974]_  & \new_[49959]_ ;
  assign \new_[231]_  = \new_[49944]_  & \new_[49929]_ ;
  assign \new_[232]_  = \new_[49914]_  & \new_[49899]_ ;
  assign \new_[233]_  = \new_[49884]_  & \new_[49869]_ ;
  assign \new_[234]_  = \new_[49854]_  & \new_[49839]_ ;
  assign \new_[235]_  = \new_[49824]_  & \new_[49809]_ ;
  assign \new_[236]_  = \new_[49794]_  & \new_[49779]_ ;
  assign \new_[237]_  = \new_[49764]_  & \new_[49749]_ ;
  assign \new_[238]_  = \new_[49734]_  & \new_[49719]_ ;
  assign \new_[239]_  = \new_[49704]_  & \new_[49689]_ ;
  assign \new_[240]_  = \new_[49674]_  & \new_[49659]_ ;
  assign \new_[241]_  = \new_[49644]_  & \new_[49629]_ ;
  assign \new_[242]_  = \new_[49614]_  & \new_[49599]_ ;
  assign \new_[243]_  = \new_[49584]_  & \new_[49569]_ ;
  assign \new_[244]_  = \new_[49554]_  & \new_[49539]_ ;
  assign \new_[245]_  = \new_[49524]_  & \new_[49509]_ ;
  assign \new_[246]_  = \new_[49494]_  & \new_[49479]_ ;
  assign \new_[247]_  = \new_[49464]_  & \new_[49449]_ ;
  assign \new_[248]_  = \new_[49434]_  & \new_[49419]_ ;
  assign \new_[249]_  = \new_[49404]_  & \new_[49389]_ ;
  assign \new_[250]_  = \new_[49374]_  & \new_[49359]_ ;
  assign \new_[251]_  = \new_[49344]_  & \new_[49329]_ ;
  assign \new_[252]_  = \new_[49314]_  & \new_[49299]_ ;
  assign \new_[253]_  = \new_[49284]_  & \new_[49269]_ ;
  assign \new_[254]_  = \new_[49254]_  & \new_[49239]_ ;
  assign \new_[255]_  = \new_[49224]_  & \new_[49209]_ ;
  assign \new_[256]_  = \new_[49194]_  & \new_[49179]_ ;
  assign \new_[257]_  = \new_[49164]_  & \new_[49149]_ ;
  assign \new_[258]_  = \new_[49134]_  & \new_[49119]_ ;
  assign \new_[259]_  = \new_[49104]_  & \new_[49089]_ ;
  assign \new_[260]_  = \new_[49074]_  & \new_[49059]_ ;
  assign \new_[261]_  = \new_[49044]_  & \new_[49029]_ ;
  assign \new_[262]_  = \new_[49014]_  & \new_[48999]_ ;
  assign \new_[263]_  = \new_[48984]_  & \new_[48969]_ ;
  assign \new_[264]_  = \new_[48954]_  & \new_[48939]_ ;
  assign \new_[265]_  = \new_[48924]_  & \new_[48909]_ ;
  assign \new_[266]_  = \new_[48894]_  & \new_[48879]_ ;
  assign \new_[267]_  = \new_[48864]_  & \new_[48849]_ ;
  assign \new_[268]_  = \new_[48834]_  & \new_[48819]_ ;
  assign \new_[269]_  = \new_[48804]_  & \new_[48789]_ ;
  assign \new_[270]_  = \new_[48774]_  & \new_[48759]_ ;
  assign \new_[271]_  = \new_[48744]_  & \new_[48729]_ ;
  assign \new_[272]_  = \new_[48714]_  & \new_[48699]_ ;
  assign \new_[273]_  = \new_[48684]_  & \new_[48669]_ ;
  assign \new_[274]_  = \new_[48654]_  & \new_[48639]_ ;
  assign \new_[275]_  = \new_[48624]_  & \new_[48609]_ ;
  assign \new_[276]_  = \new_[48594]_  & \new_[48579]_ ;
  assign \new_[277]_  = \new_[48564]_  & \new_[48549]_ ;
  assign \new_[278]_  = \new_[48534]_  & \new_[48519]_ ;
  assign \new_[279]_  = \new_[48504]_  & \new_[48489]_ ;
  assign \new_[280]_  = \new_[48474]_  & \new_[48459]_ ;
  assign \new_[281]_  = \new_[48444]_  & \new_[48429]_ ;
  assign \new_[282]_  = \new_[48414]_  & \new_[48399]_ ;
  assign \new_[283]_  = \new_[48384]_  & \new_[48369]_ ;
  assign \new_[284]_  = \new_[48354]_  & \new_[48339]_ ;
  assign \new_[285]_  = \new_[48324]_  & \new_[48309]_ ;
  assign \new_[286]_  = \new_[48294]_  & \new_[48279]_ ;
  assign \new_[287]_  = \new_[48264]_  & \new_[48249]_ ;
  assign \new_[288]_  = \new_[48234]_  & \new_[48219]_ ;
  assign \new_[289]_  = \new_[48204]_  & \new_[48189]_ ;
  assign \new_[290]_  = \new_[48174]_  & \new_[48159]_ ;
  assign \new_[291]_  = \new_[48144]_  & \new_[48129]_ ;
  assign \new_[292]_  = \new_[48114]_  & \new_[48099]_ ;
  assign \new_[293]_  = \new_[48084]_  & \new_[48069]_ ;
  assign \new_[294]_  = \new_[48054]_  & \new_[48039]_ ;
  assign \new_[295]_  = \new_[48024]_  & \new_[48009]_ ;
  assign \new_[296]_  = \new_[47994]_  & \new_[47979]_ ;
  assign \new_[297]_  = \new_[47964]_  & \new_[47949]_ ;
  assign \new_[298]_  = \new_[47934]_  & \new_[47919]_ ;
  assign \new_[299]_  = \new_[47904]_  & \new_[47889]_ ;
  assign \new_[300]_  = \new_[47874]_  & \new_[47859]_ ;
  assign \new_[301]_  = \new_[47844]_  & \new_[47829]_ ;
  assign \new_[302]_  = \new_[47814]_  & \new_[47799]_ ;
  assign \new_[303]_  = \new_[47784]_  & \new_[47769]_ ;
  assign \new_[304]_  = \new_[47754]_  & \new_[47739]_ ;
  assign \new_[305]_  = \new_[47724]_  & \new_[47709]_ ;
  assign \new_[306]_  = \new_[47694]_  & \new_[47679]_ ;
  assign \new_[307]_  = \new_[47664]_  & \new_[47649]_ ;
  assign \new_[308]_  = \new_[47634]_  & \new_[47619]_ ;
  assign \new_[309]_  = \new_[47604]_  & \new_[47589]_ ;
  assign \new_[310]_  = \new_[47574]_  & \new_[47559]_ ;
  assign \new_[311]_  = \new_[47544]_  & \new_[47529]_ ;
  assign \new_[312]_  = \new_[47514]_  & \new_[47499]_ ;
  assign \new_[313]_  = \new_[47484]_  & \new_[47469]_ ;
  assign \new_[314]_  = \new_[47454]_  & \new_[47439]_ ;
  assign \new_[315]_  = \new_[47424]_  & \new_[47409]_ ;
  assign \new_[316]_  = \new_[47394]_  & \new_[47379]_ ;
  assign \new_[317]_  = \new_[47364]_  & \new_[47349]_ ;
  assign \new_[318]_  = \new_[47334]_  & \new_[47319]_ ;
  assign \new_[319]_  = \new_[47304]_  & \new_[47289]_ ;
  assign \new_[320]_  = \new_[47274]_  & \new_[47259]_ ;
  assign \new_[321]_  = \new_[47244]_  & \new_[47229]_ ;
  assign \new_[322]_  = \new_[47214]_  & \new_[47199]_ ;
  assign \new_[323]_  = \new_[47184]_  & \new_[47169]_ ;
  assign \new_[324]_  = \new_[47154]_  & \new_[47139]_ ;
  assign \new_[325]_  = \new_[47124]_  & \new_[47109]_ ;
  assign \new_[326]_  = \new_[47094]_  & \new_[47079]_ ;
  assign \new_[327]_  = \new_[47064]_  & \new_[47049]_ ;
  assign \new_[328]_  = \new_[47034]_  & \new_[47019]_ ;
  assign \new_[329]_  = \new_[47004]_  & \new_[46989]_ ;
  assign \new_[330]_  = \new_[46974]_  & \new_[46959]_ ;
  assign \new_[331]_  = \new_[46944]_  & \new_[46929]_ ;
  assign \new_[332]_  = \new_[46914]_  & \new_[46899]_ ;
  assign \new_[333]_  = \new_[46884]_  & \new_[46869]_ ;
  assign \new_[334]_  = \new_[46854]_  & \new_[46839]_ ;
  assign \new_[335]_  = \new_[46824]_  & \new_[46809]_ ;
  assign \new_[336]_  = \new_[46794]_  & \new_[46779]_ ;
  assign \new_[337]_  = \new_[46764]_  & \new_[46749]_ ;
  assign \new_[338]_  = \new_[46734]_  & \new_[46719]_ ;
  assign \new_[339]_  = \new_[46704]_  & \new_[46689]_ ;
  assign \new_[340]_  = \new_[46674]_  & \new_[46659]_ ;
  assign \new_[341]_  = \new_[46644]_  & \new_[46629]_ ;
  assign \new_[342]_  = \new_[46614]_  & \new_[46599]_ ;
  assign \new_[343]_  = \new_[46584]_  & \new_[46569]_ ;
  assign \new_[344]_  = \new_[46554]_  & \new_[46539]_ ;
  assign \new_[345]_  = \new_[46524]_  & \new_[46509]_ ;
  assign \new_[346]_  = \new_[46494]_  & \new_[46479]_ ;
  assign \new_[347]_  = \new_[46464]_  & \new_[46449]_ ;
  assign \new_[348]_  = \new_[46434]_  & \new_[46419]_ ;
  assign \new_[349]_  = \new_[46404]_  & \new_[46389]_ ;
  assign \new_[350]_  = \new_[46374]_  & \new_[46359]_ ;
  assign \new_[351]_  = \new_[46344]_  & \new_[46329]_ ;
  assign \new_[352]_  = \new_[46314]_  & \new_[46299]_ ;
  assign \new_[353]_  = \new_[46284]_  & \new_[46269]_ ;
  assign \new_[354]_  = \new_[46254]_  & \new_[46239]_ ;
  assign \new_[355]_  = \new_[46224]_  & \new_[46209]_ ;
  assign \new_[356]_  = \new_[46194]_  & \new_[46179]_ ;
  assign \new_[357]_  = \new_[46164]_  & \new_[46149]_ ;
  assign \new_[358]_  = \new_[46134]_  & \new_[46119]_ ;
  assign \new_[359]_  = \new_[46104]_  & \new_[46089]_ ;
  assign \new_[360]_  = \new_[46074]_  & \new_[46059]_ ;
  assign \new_[361]_  = \new_[46044]_  & \new_[46029]_ ;
  assign \new_[362]_  = \new_[46014]_  & \new_[45999]_ ;
  assign \new_[363]_  = \new_[45984]_  & \new_[45969]_ ;
  assign \new_[364]_  = \new_[45954]_  & \new_[45939]_ ;
  assign \new_[365]_  = \new_[45924]_  & \new_[45909]_ ;
  assign \new_[366]_  = \new_[45894]_  & \new_[45879]_ ;
  assign \new_[367]_  = \new_[45864]_  & \new_[45849]_ ;
  assign \new_[368]_  = \new_[45834]_  & \new_[45819]_ ;
  assign \new_[369]_  = \new_[45804]_  & \new_[45789]_ ;
  assign \new_[370]_  = \new_[45774]_  & \new_[45759]_ ;
  assign \new_[371]_  = \new_[45744]_  & \new_[45729]_ ;
  assign \new_[372]_  = \new_[45714]_  & \new_[45699]_ ;
  assign \new_[373]_  = \new_[45684]_  & \new_[45669]_ ;
  assign \new_[374]_  = \new_[45654]_  & \new_[45639]_ ;
  assign \new_[375]_  = \new_[45624]_  & \new_[45609]_ ;
  assign \new_[376]_  = \new_[45594]_  & \new_[45579]_ ;
  assign \new_[377]_  = \new_[45564]_  & \new_[45549]_ ;
  assign \new_[378]_  = \new_[45534]_  & \new_[45519]_ ;
  assign \new_[379]_  = \new_[45504]_  & \new_[45489]_ ;
  assign \new_[380]_  = \new_[45474]_  & \new_[45459]_ ;
  assign \new_[381]_  = \new_[45444]_  & \new_[45429]_ ;
  assign \new_[382]_  = \new_[45414]_  & \new_[45399]_ ;
  assign \new_[383]_  = \new_[45384]_  & \new_[45369]_ ;
  assign \new_[384]_  = \new_[45354]_  & \new_[45339]_ ;
  assign \new_[385]_  = \new_[45324]_  & \new_[45309]_ ;
  assign \new_[386]_  = \new_[45294]_  & \new_[45279]_ ;
  assign \new_[387]_  = \new_[45264]_  & \new_[45249]_ ;
  assign \new_[388]_  = \new_[45234]_  & \new_[45219]_ ;
  assign \new_[389]_  = \new_[45204]_  & \new_[45189]_ ;
  assign \new_[390]_  = \new_[45174]_  & \new_[45159]_ ;
  assign \new_[391]_  = \new_[45144]_  & \new_[45129]_ ;
  assign \new_[392]_  = \new_[45114]_  & \new_[45099]_ ;
  assign \new_[393]_  = \new_[45084]_  & \new_[45069]_ ;
  assign \new_[394]_  = \new_[45054]_  & \new_[45039]_ ;
  assign \new_[395]_  = \new_[45024]_  & \new_[45009]_ ;
  assign \new_[396]_  = \new_[44994]_  & \new_[44979]_ ;
  assign \new_[397]_  = \new_[44964]_  & \new_[44949]_ ;
  assign \new_[398]_  = \new_[44934]_  & \new_[44919]_ ;
  assign \new_[399]_  = \new_[44904]_  & \new_[44889]_ ;
  assign \new_[400]_  = \new_[44874]_  & \new_[44859]_ ;
  assign \new_[401]_  = \new_[44844]_  & \new_[44829]_ ;
  assign \new_[402]_  = \new_[44814]_  & \new_[44799]_ ;
  assign \new_[403]_  = \new_[44784]_  & \new_[44769]_ ;
  assign \new_[404]_  = \new_[44754]_  & \new_[44739]_ ;
  assign \new_[405]_  = \new_[44724]_  & \new_[44709]_ ;
  assign \new_[406]_  = \new_[44694]_  & \new_[44679]_ ;
  assign \new_[407]_  = \new_[44664]_  & \new_[44649]_ ;
  assign \new_[408]_  = \new_[44634]_  & \new_[44619]_ ;
  assign \new_[409]_  = \new_[44604]_  & \new_[44589]_ ;
  assign \new_[410]_  = \new_[44574]_  & \new_[44559]_ ;
  assign \new_[411]_  = \new_[44544]_  & \new_[44529]_ ;
  assign \new_[412]_  = \new_[44516]_  & \new_[44501]_ ;
  assign \new_[413]_  = \new_[44488]_  & \new_[44473]_ ;
  assign \new_[414]_  = \new_[44460]_  & \new_[44445]_ ;
  assign \new_[415]_  = \new_[44432]_  & \new_[44417]_ ;
  assign \new_[416]_  = \new_[44404]_  & \new_[44389]_ ;
  assign \new_[417]_  = \new_[44376]_  & \new_[44361]_ ;
  assign \new_[418]_  = \new_[44348]_  & \new_[44333]_ ;
  assign \new_[419]_  = \new_[44320]_  & \new_[44305]_ ;
  assign \new_[420]_  = \new_[44292]_  & \new_[44277]_ ;
  assign \new_[421]_  = \new_[44264]_  & \new_[44249]_ ;
  assign \new_[422]_  = \new_[44236]_  & \new_[44221]_ ;
  assign \new_[423]_  = \new_[44208]_  & \new_[44193]_ ;
  assign \new_[424]_  = \new_[44180]_  & \new_[44165]_ ;
  assign \new_[425]_  = \new_[44152]_  & \new_[44137]_ ;
  assign \new_[426]_  = \new_[44124]_  & \new_[44109]_ ;
  assign \new_[427]_  = \new_[44096]_  & \new_[44081]_ ;
  assign \new_[428]_  = \new_[44068]_  & \new_[44053]_ ;
  assign \new_[429]_  = \new_[44040]_  & \new_[44025]_ ;
  assign \new_[430]_  = \new_[44012]_  & \new_[43997]_ ;
  assign \new_[431]_  = \new_[43984]_  & \new_[43969]_ ;
  assign \new_[432]_  = \new_[43956]_  & \new_[43941]_ ;
  assign \new_[433]_  = \new_[43928]_  & \new_[43913]_ ;
  assign \new_[434]_  = \new_[43900]_  & \new_[43885]_ ;
  assign \new_[435]_  = \new_[43872]_  & \new_[43857]_ ;
  assign \new_[436]_  = \new_[43844]_  & \new_[43829]_ ;
  assign \new_[437]_  = \new_[43816]_  & \new_[43801]_ ;
  assign \new_[438]_  = \new_[43788]_  & \new_[43773]_ ;
  assign \new_[439]_  = \new_[43760]_  & \new_[43745]_ ;
  assign \new_[440]_  = \new_[43732]_  & \new_[43717]_ ;
  assign \new_[441]_  = \new_[43704]_  & \new_[43689]_ ;
  assign \new_[442]_  = \new_[43676]_  & \new_[43661]_ ;
  assign \new_[443]_  = \new_[43648]_  & \new_[43633]_ ;
  assign \new_[444]_  = \new_[43620]_  & \new_[43605]_ ;
  assign \new_[445]_  = \new_[43592]_  & \new_[43577]_ ;
  assign \new_[446]_  = \new_[43564]_  & \new_[43549]_ ;
  assign \new_[447]_  = \new_[43536]_  & \new_[43521]_ ;
  assign \new_[448]_  = \new_[43508]_  & \new_[43493]_ ;
  assign \new_[449]_  = \new_[43480]_  & \new_[43465]_ ;
  assign \new_[450]_  = \new_[43452]_  & \new_[43437]_ ;
  assign \new_[451]_  = \new_[43424]_  & \new_[43409]_ ;
  assign \new_[452]_  = \new_[43396]_  & \new_[43381]_ ;
  assign \new_[453]_  = \new_[43368]_  & \new_[43353]_ ;
  assign \new_[454]_  = \new_[43340]_  & \new_[43325]_ ;
  assign \new_[455]_  = \new_[43312]_  & \new_[43297]_ ;
  assign \new_[456]_  = \new_[43284]_  & \new_[43269]_ ;
  assign \new_[457]_  = \new_[43256]_  & \new_[43241]_ ;
  assign \new_[458]_  = \new_[43228]_  & \new_[43213]_ ;
  assign \new_[459]_  = \new_[43200]_  & \new_[43185]_ ;
  assign \new_[460]_  = \new_[43172]_  & \new_[43157]_ ;
  assign \new_[461]_  = \new_[43144]_  & \new_[43129]_ ;
  assign \new_[462]_  = \new_[43116]_  & \new_[43101]_ ;
  assign \new_[463]_  = \new_[43088]_  & \new_[43073]_ ;
  assign \new_[464]_  = \new_[43060]_  & \new_[43045]_ ;
  assign \new_[465]_  = \new_[43032]_  & \new_[43017]_ ;
  assign \new_[466]_  = \new_[43004]_  & \new_[42989]_ ;
  assign \new_[467]_  = \new_[42976]_  & \new_[42961]_ ;
  assign \new_[468]_  = \new_[42948]_  & \new_[42933]_ ;
  assign \new_[469]_  = \new_[42920]_  & \new_[42905]_ ;
  assign \new_[470]_  = \new_[42892]_  & \new_[42877]_ ;
  assign \new_[471]_  = \new_[42864]_  & \new_[42849]_ ;
  assign \new_[472]_  = \new_[42836]_  & \new_[42821]_ ;
  assign \new_[473]_  = \new_[42808]_  & \new_[42793]_ ;
  assign \new_[474]_  = \new_[42780]_  & \new_[42765]_ ;
  assign \new_[475]_  = \new_[42752]_  & \new_[42737]_ ;
  assign \new_[476]_  = \new_[42724]_  & \new_[42709]_ ;
  assign \new_[477]_  = \new_[42696]_  & \new_[42681]_ ;
  assign \new_[478]_  = \new_[42668]_  & \new_[42653]_ ;
  assign \new_[479]_  = \new_[42640]_  & \new_[42625]_ ;
  assign \new_[480]_  = \new_[42612]_  & \new_[42597]_ ;
  assign \new_[481]_  = \new_[42584]_  & \new_[42569]_ ;
  assign \new_[482]_  = \new_[42556]_  & \new_[42541]_ ;
  assign \new_[483]_  = \new_[42528]_  & \new_[42513]_ ;
  assign \new_[484]_  = \new_[42500]_  & \new_[42485]_ ;
  assign \new_[485]_  = \new_[42472]_  & \new_[42457]_ ;
  assign \new_[486]_  = \new_[42444]_  & \new_[42429]_ ;
  assign \new_[487]_  = \new_[42416]_  & \new_[42401]_ ;
  assign \new_[488]_  = \new_[42388]_  & \new_[42373]_ ;
  assign \new_[489]_  = \new_[42360]_  & \new_[42345]_ ;
  assign \new_[490]_  = \new_[42332]_  & \new_[42317]_ ;
  assign \new_[491]_  = \new_[42304]_  & \new_[42289]_ ;
  assign \new_[492]_  = \new_[42276]_  & \new_[42261]_ ;
  assign \new_[493]_  = \new_[42248]_  & \new_[42233]_ ;
  assign \new_[494]_  = \new_[42220]_  & \new_[42205]_ ;
  assign \new_[495]_  = \new_[42192]_  & \new_[42177]_ ;
  assign \new_[496]_  = \new_[42164]_  & \new_[42149]_ ;
  assign \new_[497]_  = \new_[42136]_  & \new_[42121]_ ;
  assign \new_[498]_  = \new_[42108]_  & \new_[42093]_ ;
  assign \new_[499]_  = \new_[42080]_  & \new_[42065]_ ;
  assign \new_[500]_  = \new_[42052]_  & \new_[42037]_ ;
  assign \new_[501]_  = \new_[42024]_  & \new_[42009]_ ;
  assign \new_[502]_  = \new_[41996]_  & \new_[41981]_ ;
  assign \new_[503]_  = \new_[41968]_  & \new_[41953]_ ;
  assign \new_[504]_  = \new_[41940]_  & \new_[41925]_ ;
  assign \new_[505]_  = \new_[41912]_  & \new_[41897]_ ;
  assign \new_[506]_  = \new_[41884]_  & \new_[41869]_ ;
  assign \new_[507]_  = \new_[41856]_  & \new_[41841]_ ;
  assign \new_[508]_  = \new_[41828]_  & \new_[41813]_ ;
  assign \new_[509]_  = \new_[41800]_  & \new_[41785]_ ;
  assign \new_[510]_  = \new_[41772]_  & \new_[41757]_ ;
  assign \new_[511]_  = \new_[41744]_  & \new_[41729]_ ;
  assign \new_[512]_  = \new_[41716]_  & \new_[41701]_ ;
  assign \new_[513]_  = \new_[41688]_  & \new_[41673]_ ;
  assign \new_[514]_  = \new_[41660]_  & \new_[41645]_ ;
  assign \new_[515]_  = \new_[41632]_  & \new_[41617]_ ;
  assign \new_[516]_  = \new_[41604]_  & \new_[41589]_ ;
  assign \new_[517]_  = \new_[41576]_  & \new_[41561]_ ;
  assign \new_[518]_  = \new_[41548]_  & \new_[41533]_ ;
  assign \new_[519]_  = \new_[41520]_  & \new_[41505]_ ;
  assign \new_[520]_  = \new_[41492]_  & \new_[41477]_ ;
  assign \new_[521]_  = \new_[41464]_  & \new_[41449]_ ;
  assign \new_[522]_  = \new_[41436]_  & \new_[41421]_ ;
  assign \new_[523]_  = \new_[41408]_  & \new_[41393]_ ;
  assign \new_[524]_  = \new_[41380]_  & \new_[41365]_ ;
  assign \new_[525]_  = \new_[41352]_  & \new_[41337]_ ;
  assign \new_[526]_  = \new_[41324]_  & \new_[41309]_ ;
  assign \new_[527]_  = \new_[41296]_  & \new_[41281]_ ;
  assign \new_[528]_  = \new_[41268]_  & \new_[41253]_ ;
  assign \new_[529]_  = \new_[41240]_  & \new_[41225]_ ;
  assign \new_[530]_  = \new_[41212]_  & \new_[41197]_ ;
  assign \new_[531]_  = \new_[41184]_  & \new_[41169]_ ;
  assign \new_[532]_  = \new_[41156]_  & \new_[41141]_ ;
  assign \new_[533]_  = \new_[41128]_  & \new_[41113]_ ;
  assign \new_[534]_  = \new_[41100]_  & \new_[41085]_ ;
  assign \new_[535]_  = \new_[41072]_  & \new_[41057]_ ;
  assign \new_[536]_  = \new_[41044]_  & \new_[41029]_ ;
  assign \new_[537]_  = \new_[41016]_  & \new_[41001]_ ;
  assign \new_[538]_  = \new_[40988]_  & \new_[40973]_ ;
  assign \new_[539]_  = \new_[40960]_  & \new_[40945]_ ;
  assign \new_[540]_  = \new_[40932]_  & \new_[40917]_ ;
  assign \new_[541]_  = \new_[40904]_  & \new_[40889]_ ;
  assign \new_[542]_  = \new_[40876]_  & \new_[40861]_ ;
  assign \new_[543]_  = \new_[40848]_  & \new_[40833]_ ;
  assign \new_[544]_  = \new_[40820]_  & \new_[40805]_ ;
  assign \new_[545]_  = \new_[40792]_  & \new_[40777]_ ;
  assign \new_[546]_  = \new_[40764]_  & \new_[40749]_ ;
  assign \new_[547]_  = \new_[40736]_  & \new_[40721]_ ;
  assign \new_[548]_  = \new_[40708]_  & \new_[40693]_ ;
  assign \new_[549]_  = \new_[40680]_  & \new_[40665]_ ;
  assign \new_[550]_  = \new_[40652]_  & \new_[40637]_ ;
  assign \new_[551]_  = \new_[40624]_  & \new_[40609]_ ;
  assign \new_[552]_  = \new_[40596]_  & \new_[40581]_ ;
  assign \new_[553]_  = \new_[40568]_  & \new_[40553]_ ;
  assign \new_[554]_  = \new_[40540]_  & \new_[40525]_ ;
  assign \new_[555]_  = \new_[40512]_  & \new_[40497]_ ;
  assign \new_[556]_  = \new_[40484]_  & \new_[40469]_ ;
  assign \new_[557]_  = \new_[40456]_  & \new_[40441]_ ;
  assign \new_[558]_  = \new_[40428]_  & \new_[40413]_ ;
  assign \new_[559]_  = \new_[40400]_  & \new_[40385]_ ;
  assign \new_[560]_  = \new_[40372]_  & \new_[40357]_ ;
  assign \new_[561]_  = \new_[40344]_  & \new_[40329]_ ;
  assign \new_[562]_  = \new_[40316]_  & \new_[40301]_ ;
  assign \new_[563]_  = \new_[40288]_  & \new_[40273]_ ;
  assign \new_[564]_  = \new_[40260]_  & \new_[40245]_ ;
  assign \new_[565]_  = \new_[40232]_  & \new_[40217]_ ;
  assign \new_[566]_  = \new_[40204]_  & \new_[40189]_ ;
  assign \new_[567]_  = \new_[40176]_  & \new_[40161]_ ;
  assign \new_[568]_  = \new_[40148]_  & \new_[40133]_ ;
  assign \new_[569]_  = \new_[40120]_  & \new_[40105]_ ;
  assign \new_[570]_  = \new_[40092]_  & \new_[40077]_ ;
  assign \new_[571]_  = \new_[40064]_  & \new_[40049]_ ;
  assign \new_[572]_  = \new_[40036]_  & \new_[40021]_ ;
  assign \new_[573]_  = \new_[40008]_  & \new_[39993]_ ;
  assign \new_[574]_  = \new_[39980]_  & \new_[39965]_ ;
  assign \new_[575]_  = \new_[39952]_  & \new_[39937]_ ;
  assign \new_[576]_  = \new_[39924]_  & \new_[39909]_ ;
  assign \new_[577]_  = \new_[39896]_  & \new_[39881]_ ;
  assign \new_[578]_  = \new_[39868]_  & \new_[39853]_ ;
  assign \new_[579]_  = \new_[39840]_  & \new_[39825]_ ;
  assign \new_[580]_  = \new_[39812]_  & \new_[39797]_ ;
  assign \new_[581]_  = \new_[39784]_  & \new_[39769]_ ;
  assign \new_[582]_  = \new_[39756]_  & \new_[39741]_ ;
  assign \new_[583]_  = \new_[39728]_  & \new_[39713]_ ;
  assign \new_[584]_  = \new_[39700]_  & \new_[39685]_ ;
  assign \new_[585]_  = \new_[39672]_  & \new_[39657]_ ;
  assign \new_[586]_  = \new_[39644]_  & \new_[39629]_ ;
  assign \new_[587]_  = \new_[39616]_  & \new_[39601]_ ;
  assign \new_[588]_  = \new_[39588]_  & \new_[39573]_ ;
  assign \new_[589]_  = \new_[39560]_  & \new_[39545]_ ;
  assign \new_[590]_  = \new_[39532]_  & \new_[39517]_ ;
  assign \new_[591]_  = \new_[39504]_  & \new_[39489]_ ;
  assign \new_[592]_  = \new_[39476]_  & \new_[39461]_ ;
  assign \new_[593]_  = \new_[39448]_  & \new_[39433]_ ;
  assign \new_[594]_  = \new_[39420]_  & \new_[39405]_ ;
  assign \new_[595]_  = \new_[39392]_  & \new_[39377]_ ;
  assign \new_[596]_  = \new_[39364]_  & \new_[39349]_ ;
  assign \new_[597]_  = \new_[39336]_  & \new_[39321]_ ;
  assign \new_[598]_  = \new_[39308]_  & \new_[39293]_ ;
  assign \new_[599]_  = \new_[39280]_  & \new_[39265]_ ;
  assign \new_[600]_  = \new_[39252]_  & \new_[39237]_ ;
  assign \new_[601]_  = \new_[39224]_  & \new_[39209]_ ;
  assign \new_[602]_  = \new_[39196]_  & \new_[39181]_ ;
  assign \new_[603]_  = \new_[39168]_  & \new_[39153]_ ;
  assign \new_[604]_  = \new_[39140]_  & \new_[39125]_ ;
  assign \new_[605]_  = \new_[39112]_  & \new_[39097]_ ;
  assign \new_[606]_  = \new_[39084]_  & \new_[39069]_ ;
  assign \new_[607]_  = \new_[39056]_  & \new_[39041]_ ;
  assign \new_[608]_  = \new_[39028]_  & \new_[39013]_ ;
  assign \new_[609]_  = \new_[39000]_  & \new_[38985]_ ;
  assign \new_[610]_  = \new_[38972]_  & \new_[38957]_ ;
  assign \new_[611]_  = \new_[38944]_  & \new_[38929]_ ;
  assign \new_[612]_  = \new_[38916]_  & \new_[38901]_ ;
  assign \new_[613]_  = \new_[38888]_  & \new_[38873]_ ;
  assign \new_[614]_  = \new_[38860]_  & \new_[38845]_ ;
  assign \new_[615]_  = \new_[38832]_  & \new_[38817]_ ;
  assign \new_[616]_  = \new_[38804]_  & \new_[38789]_ ;
  assign \new_[617]_  = \new_[38776]_  & \new_[38761]_ ;
  assign \new_[618]_  = \new_[38748]_  & \new_[38733]_ ;
  assign \new_[619]_  = \new_[38720]_  & \new_[38705]_ ;
  assign \new_[620]_  = \new_[38692]_  & \new_[38677]_ ;
  assign \new_[621]_  = \new_[38664]_  & \new_[38649]_ ;
  assign \new_[622]_  = \new_[38636]_  & \new_[38621]_ ;
  assign \new_[623]_  = \new_[38608]_  & \new_[38593]_ ;
  assign \new_[624]_  = \new_[38580]_  & \new_[38565]_ ;
  assign \new_[625]_  = \new_[38552]_  & \new_[38537]_ ;
  assign \new_[626]_  = \new_[38524]_  & \new_[38509]_ ;
  assign \new_[627]_  = \new_[38496]_  & \new_[38481]_ ;
  assign \new_[628]_  = \new_[38468]_  & \new_[38453]_ ;
  assign \new_[629]_  = \new_[38440]_  & \new_[38425]_ ;
  assign \new_[630]_  = \new_[38412]_  & \new_[38397]_ ;
  assign \new_[631]_  = \new_[38384]_  & \new_[38369]_ ;
  assign \new_[632]_  = \new_[38356]_  & \new_[38341]_ ;
  assign \new_[633]_  = \new_[38328]_  & \new_[38313]_ ;
  assign \new_[634]_  = \new_[38300]_  & \new_[38285]_ ;
  assign \new_[635]_  = \new_[38272]_  & \new_[38257]_ ;
  assign \new_[636]_  = \new_[38244]_  & \new_[38229]_ ;
  assign \new_[637]_  = \new_[38216]_  & \new_[38201]_ ;
  assign \new_[638]_  = \new_[38188]_  & \new_[38173]_ ;
  assign \new_[639]_  = \new_[38160]_  & \new_[38145]_ ;
  assign \new_[640]_  = \new_[38132]_  & \new_[38117]_ ;
  assign \new_[641]_  = \new_[38104]_  & \new_[38089]_ ;
  assign \new_[642]_  = \new_[38076]_  & \new_[38061]_ ;
  assign \new_[643]_  = \new_[38048]_  & \new_[38033]_ ;
  assign \new_[644]_  = \new_[38020]_  & \new_[38005]_ ;
  assign \new_[645]_  = \new_[37992]_  & \new_[37977]_ ;
  assign \new_[646]_  = \new_[37964]_  & \new_[37949]_ ;
  assign \new_[647]_  = \new_[37936]_  & \new_[37921]_ ;
  assign \new_[648]_  = \new_[37908]_  & \new_[37893]_ ;
  assign \new_[649]_  = \new_[37880]_  & \new_[37865]_ ;
  assign \new_[650]_  = \new_[37852]_  & \new_[37837]_ ;
  assign \new_[651]_  = \new_[37824]_  & \new_[37811]_ ;
  assign \new_[652]_  = \new_[37798]_  & \new_[37785]_ ;
  assign \new_[653]_  = \new_[37772]_  & \new_[37759]_ ;
  assign \new_[654]_  = \new_[37746]_  & \new_[37733]_ ;
  assign \new_[655]_  = \new_[37720]_  & \new_[37707]_ ;
  assign \new_[656]_  = \new_[37694]_  & \new_[37681]_ ;
  assign \new_[657]_  = \new_[37668]_  & \new_[37655]_ ;
  assign \new_[658]_  = \new_[37642]_  & \new_[37629]_ ;
  assign \new_[659]_  = \new_[37616]_  & \new_[37603]_ ;
  assign \new_[660]_  = \new_[37590]_  & \new_[37577]_ ;
  assign \new_[661]_  = \new_[37564]_  & \new_[37551]_ ;
  assign \new_[662]_  = \new_[37538]_  & \new_[37525]_ ;
  assign \new_[663]_  = \new_[37512]_  & \new_[37499]_ ;
  assign \new_[664]_  = \new_[37486]_  & \new_[37473]_ ;
  assign \new_[665]_  = \new_[37460]_  & \new_[37447]_ ;
  assign \new_[666]_  = \new_[37434]_  & \new_[37421]_ ;
  assign \new_[667]_  = \new_[37408]_  & \new_[37395]_ ;
  assign \new_[668]_  = \new_[37382]_  & \new_[37369]_ ;
  assign \new_[669]_  = \new_[37356]_  & \new_[37343]_ ;
  assign \new_[670]_  = \new_[37330]_  & \new_[37317]_ ;
  assign \new_[671]_  = \new_[37304]_  & \new_[37291]_ ;
  assign \new_[672]_  = \new_[37278]_  & \new_[37265]_ ;
  assign \new_[673]_  = \new_[37252]_  & \new_[37239]_ ;
  assign \new_[674]_  = \new_[37226]_  & \new_[37213]_ ;
  assign \new_[675]_  = \new_[37200]_  & \new_[37187]_ ;
  assign \new_[676]_  = \new_[37174]_  & \new_[37161]_ ;
  assign \new_[677]_  = \new_[37148]_  & \new_[37135]_ ;
  assign \new_[678]_  = \new_[37122]_  & \new_[37109]_ ;
  assign \new_[679]_  = \new_[37096]_  & \new_[37083]_ ;
  assign \new_[680]_  = \new_[37070]_  & \new_[37057]_ ;
  assign \new_[681]_  = \new_[37044]_  & \new_[37031]_ ;
  assign \new_[682]_  = \new_[37018]_  & \new_[37005]_ ;
  assign \new_[683]_  = \new_[36992]_  & \new_[36979]_ ;
  assign \new_[684]_  = \new_[36966]_  & \new_[36953]_ ;
  assign \new_[685]_  = \new_[36940]_  & \new_[36927]_ ;
  assign \new_[686]_  = \new_[36914]_  & \new_[36901]_ ;
  assign \new_[687]_  = \new_[36888]_  & \new_[36875]_ ;
  assign \new_[688]_  = \new_[36862]_  & \new_[36849]_ ;
  assign \new_[689]_  = \new_[36836]_  & \new_[36823]_ ;
  assign \new_[690]_  = \new_[36810]_  & \new_[36797]_ ;
  assign \new_[691]_  = \new_[36784]_  & \new_[36771]_ ;
  assign \new_[692]_  = \new_[36758]_  & \new_[36745]_ ;
  assign \new_[693]_  = \new_[36732]_  & \new_[36719]_ ;
  assign \new_[694]_  = \new_[36706]_  & \new_[36693]_ ;
  assign \new_[695]_  = \new_[36680]_  & \new_[36667]_ ;
  assign \new_[696]_  = \new_[36654]_  & \new_[36641]_ ;
  assign \new_[697]_  = \new_[36628]_  & \new_[36615]_ ;
  assign \new_[698]_  = \new_[36602]_  & \new_[36589]_ ;
  assign \new_[699]_  = \new_[36576]_  & \new_[36563]_ ;
  assign \new_[700]_  = \new_[36550]_  & \new_[36537]_ ;
  assign \new_[701]_  = \new_[36524]_  & \new_[36511]_ ;
  assign \new_[702]_  = \new_[36498]_  & \new_[36485]_ ;
  assign \new_[703]_  = \new_[36472]_  & \new_[36459]_ ;
  assign \new_[704]_  = \new_[36446]_  & \new_[36433]_ ;
  assign \new_[705]_  = \new_[36420]_  & \new_[36407]_ ;
  assign \new_[706]_  = \new_[36394]_  & \new_[36381]_ ;
  assign \new_[707]_  = \new_[36368]_  & \new_[36355]_ ;
  assign \new_[708]_  = \new_[36342]_  & \new_[36329]_ ;
  assign \new_[709]_  = \new_[36316]_  & \new_[36303]_ ;
  assign \new_[710]_  = \new_[36290]_  & \new_[36277]_ ;
  assign \new_[711]_  = \new_[36264]_  & \new_[36251]_ ;
  assign \new_[712]_  = \new_[36238]_  & \new_[36225]_ ;
  assign \new_[713]_  = \new_[36212]_  & \new_[36199]_ ;
  assign \new_[714]_  = \new_[36186]_  & \new_[36173]_ ;
  assign \new_[715]_  = \new_[36160]_  & \new_[36147]_ ;
  assign \new_[716]_  = \new_[36134]_  & \new_[36121]_ ;
  assign \new_[717]_  = \new_[36108]_  & \new_[36095]_ ;
  assign \new_[718]_  = \new_[36082]_  & \new_[36069]_ ;
  assign \new_[719]_  = \new_[36056]_  & \new_[36043]_ ;
  assign \new_[720]_  = \new_[36030]_  & \new_[36017]_ ;
  assign \new_[721]_  = \new_[36004]_  & \new_[35991]_ ;
  assign \new_[722]_  = \new_[35978]_  & \new_[35965]_ ;
  assign \new_[723]_  = \new_[35952]_  & \new_[35939]_ ;
  assign \new_[724]_  = \new_[35926]_  & \new_[35913]_ ;
  assign \new_[725]_  = \new_[35900]_  & \new_[35887]_ ;
  assign \new_[726]_  = \new_[35874]_  & \new_[35861]_ ;
  assign \new_[727]_  = \new_[35848]_  & \new_[35835]_ ;
  assign \new_[728]_  = \new_[35822]_  & \new_[35809]_ ;
  assign \new_[729]_  = \new_[35796]_  & \new_[35783]_ ;
  assign \new_[730]_  = \new_[35770]_  & \new_[35757]_ ;
  assign \new_[731]_  = \new_[35744]_  & \new_[35731]_ ;
  assign \new_[732]_  = \new_[35718]_  & \new_[35705]_ ;
  assign \new_[733]_  = \new_[35692]_  & \new_[35679]_ ;
  assign \new_[734]_  = \new_[35666]_  & \new_[35653]_ ;
  assign \new_[735]_  = \new_[35640]_  & \new_[35627]_ ;
  assign \new_[736]_  = \new_[35614]_  & \new_[35601]_ ;
  assign \new_[737]_  = \new_[35588]_  & \new_[35575]_ ;
  assign \new_[738]_  = \new_[35562]_  & \new_[35549]_ ;
  assign \new_[739]_  = \new_[35536]_  & \new_[35523]_ ;
  assign \new_[740]_  = \new_[35510]_  & \new_[35497]_ ;
  assign \new_[741]_  = \new_[35484]_  & \new_[35471]_ ;
  assign \new_[742]_  = \new_[35458]_  & \new_[35445]_ ;
  assign \new_[743]_  = \new_[35432]_  & \new_[35419]_ ;
  assign \new_[744]_  = \new_[35406]_  & \new_[35393]_ ;
  assign \new_[745]_  = \new_[35380]_  & \new_[35367]_ ;
  assign \new_[746]_  = \new_[35354]_  & \new_[35341]_ ;
  assign \new_[747]_  = \new_[35328]_  & \new_[35315]_ ;
  assign \new_[748]_  = \new_[35302]_  & \new_[35289]_ ;
  assign \new_[749]_  = \new_[35276]_  & \new_[35263]_ ;
  assign \new_[750]_  = \new_[35250]_  & \new_[35237]_ ;
  assign \new_[751]_  = \new_[35224]_  & \new_[35211]_ ;
  assign \new_[752]_  = \new_[35198]_  & \new_[35185]_ ;
  assign \new_[753]_  = \new_[35172]_  & \new_[35159]_ ;
  assign \new_[754]_  = \new_[35146]_  & \new_[35133]_ ;
  assign \new_[755]_  = \new_[35120]_  & \new_[35107]_ ;
  assign \new_[756]_  = \new_[35094]_  & \new_[35081]_ ;
  assign \new_[757]_  = \new_[35068]_  & \new_[35055]_ ;
  assign \new_[758]_  = \new_[35042]_  & \new_[35029]_ ;
  assign \new_[759]_  = \new_[35016]_  & \new_[35003]_ ;
  assign \new_[760]_  = \new_[34990]_  & \new_[34977]_ ;
  assign \new_[761]_  = \new_[34964]_  & \new_[34951]_ ;
  assign \new_[762]_  = \new_[34938]_  & \new_[34925]_ ;
  assign \new_[763]_  = \new_[34912]_  & \new_[34899]_ ;
  assign \new_[764]_  = \new_[34886]_  & \new_[34873]_ ;
  assign \new_[765]_  = \new_[34860]_  & \new_[34847]_ ;
  assign \new_[766]_  = \new_[34834]_  & \new_[34821]_ ;
  assign \new_[767]_  = \new_[34808]_  & \new_[34795]_ ;
  assign \new_[768]_  = \new_[34782]_  & \new_[34769]_ ;
  assign \new_[769]_  = \new_[34756]_  & \new_[34743]_ ;
  assign \new_[770]_  = \new_[34730]_  & \new_[34717]_ ;
  assign \new_[771]_  = \new_[34704]_  & \new_[34691]_ ;
  assign \new_[772]_  = \new_[34678]_  & \new_[34665]_ ;
  assign \new_[773]_  = \new_[34652]_  & \new_[34639]_ ;
  assign \new_[774]_  = \new_[34626]_  & \new_[34613]_ ;
  assign \new_[775]_  = \new_[34600]_  & \new_[34587]_ ;
  assign \new_[776]_  = \new_[34574]_  & \new_[34561]_ ;
  assign \new_[777]_  = \new_[34548]_  & \new_[34535]_ ;
  assign \new_[778]_  = \new_[34522]_  & \new_[34509]_ ;
  assign \new_[779]_  = \new_[34496]_  & \new_[34483]_ ;
  assign \new_[780]_  = \new_[34472]_  & \new_[34459]_ ;
  assign \new_[781]_  = \new_[34448]_  & \new_[34435]_ ;
  assign \new_[782]_  = \new_[34424]_  & \new_[34411]_ ;
  assign \new_[783]_  = \new_[34400]_  & \new_[34387]_ ;
  assign \new_[784]_  = \new_[34376]_  & \new_[34363]_ ;
  assign \new_[785]_  = \new_[34352]_  & \new_[34339]_ ;
  assign \new_[786]_  = \new_[34328]_  & \new_[34315]_ ;
  assign \new_[787]_  = \new_[34304]_  & \new_[34291]_ ;
  assign \new_[788]_  = \new_[34280]_  & \new_[34267]_ ;
  assign \new_[789]_  = \new_[34256]_  & \new_[34243]_ ;
  assign \new_[790]_  = \new_[34232]_  & \new_[34219]_ ;
  assign \new_[791]_  = \new_[34208]_  & \new_[34195]_ ;
  assign \new_[792]_  = \new_[34184]_  & \new_[34171]_ ;
  assign \new_[793]_  = \new_[34160]_  & \new_[34147]_ ;
  assign \new_[794]_  = \new_[34136]_  & \new_[34123]_ ;
  assign \new_[795]_  = \new_[34112]_  & \new_[34099]_ ;
  assign \new_[796]_  = \new_[34088]_  & \new_[34075]_ ;
  assign \new_[797]_  = \new_[34064]_  & \new_[34051]_ ;
  assign \new_[798]_  = \new_[34040]_  & \new_[34027]_ ;
  assign \new_[799]_  = \new_[34016]_  & \new_[34003]_ ;
  assign \new_[800]_  = \new_[33992]_  & \new_[33979]_ ;
  assign \new_[801]_  = \new_[33968]_  & \new_[33955]_ ;
  assign \new_[802]_  = \new_[33944]_  & \new_[33931]_ ;
  assign \new_[803]_  = \new_[33920]_  & \new_[33907]_ ;
  assign \new_[804]_  = \new_[33896]_  & \new_[33883]_ ;
  assign \new_[805]_  = \new_[33872]_  & \new_[33859]_ ;
  assign \new_[806]_  = \new_[33848]_  & \new_[33835]_ ;
  assign \new_[807]_  = \new_[33824]_  & \new_[33811]_ ;
  assign \new_[808]_  = \new_[33800]_  & \new_[33787]_ ;
  assign \new_[809]_  = \new_[33776]_  & \new_[33763]_ ;
  assign \new_[810]_  = \new_[33752]_  & \new_[33739]_ ;
  assign \new_[811]_  = \new_[33728]_  & \new_[33715]_ ;
  assign \new_[812]_  = \new_[33704]_  & \new_[33691]_ ;
  assign \new_[813]_  = \new_[33680]_  & \new_[33667]_ ;
  assign \new_[814]_  = \new_[33656]_  & \new_[33643]_ ;
  assign \new_[815]_  = \new_[33632]_  & \new_[33619]_ ;
  assign \new_[816]_  = \new_[33608]_  & \new_[33595]_ ;
  assign \new_[817]_  = \new_[33584]_  & \new_[33571]_ ;
  assign \new_[818]_  = \new_[33560]_  & \new_[33547]_ ;
  assign \new_[819]_  = \new_[33536]_  & \new_[33523]_ ;
  assign \new_[820]_  = \new_[33512]_  & \new_[33499]_ ;
  assign \new_[821]_  = \new_[33488]_  & \new_[33475]_ ;
  assign \new_[822]_  = \new_[33464]_  & \new_[33451]_ ;
  assign \new_[823]_  = \new_[33440]_  & \new_[33427]_ ;
  assign \new_[824]_  = \new_[33416]_  & \new_[33403]_ ;
  assign \new_[825]_  = \new_[33392]_  & \new_[33379]_ ;
  assign \new_[826]_  = \new_[33368]_  & \new_[33355]_ ;
  assign \new_[827]_  = \new_[33344]_  & \new_[33331]_ ;
  assign \new_[828]_  = \new_[33320]_  & \new_[33307]_ ;
  assign \new_[829]_  = \new_[33296]_  & \new_[33283]_ ;
  assign \new_[830]_  = \new_[33272]_  & \new_[33259]_ ;
  assign \new_[831]_  = \new_[33248]_  & \new_[33235]_ ;
  assign \new_[832]_  = \new_[33224]_  & \new_[33211]_ ;
  assign \new_[833]_  = \new_[33200]_  & \new_[33187]_ ;
  assign \new_[834]_  = \new_[33176]_  & \new_[33163]_ ;
  assign \new_[835]_  = \new_[33152]_  & \new_[33139]_ ;
  assign \new_[836]_  = \new_[33128]_  & \new_[33115]_ ;
  assign \new_[837]_  = \new_[33104]_  & \new_[33091]_ ;
  assign \new_[838]_  = \new_[33080]_  & \new_[33067]_ ;
  assign \new_[839]_  = \new_[33056]_  & \new_[33043]_ ;
  assign \new_[840]_  = \new_[33032]_  & \new_[33019]_ ;
  assign \new_[841]_  = \new_[33008]_  & \new_[32995]_ ;
  assign \new_[842]_  = \new_[32984]_  & \new_[32971]_ ;
  assign \new_[843]_  = \new_[32960]_  & \new_[32949]_ ;
  assign \new_[844]_  = \new_[32938]_  & \new_[32927]_ ;
  assign \new_[845]_  = \new_[32916]_  & \new_[32905]_ ;
  assign \new_[846]_  = \new_[32894]_  & \new_[32883]_ ;
  assign \new_[847]_  = \new_[32872]_  & \new_[32861]_ ;
  assign \new_[848]_  = \new_[32850]_  & \new_[32839]_ ;
  assign \new_[849]_  = \new_[32828]_  & \new_[32817]_ ;
  assign \new_[850]_  = \new_[32806]_  & \new_[32795]_ ;
  assign \new_[851]_  = \new_[32784]_  & \new_[32773]_ ;
  assign \new_[852]_  = \new_[32762]_  & \new_[32751]_ ;
  assign \new_[853]_  = \new_[32740]_  & \new_[32729]_ ;
  assign \new_[854]_  = \new_[32718]_  & \new_[32707]_ ;
  assign \new_[855]_  = \new_[32696]_  & \new_[32685]_ ;
  assign \new_[856]_  = \new_[32674]_  & \new_[32663]_ ;
  assign \new_[857]_  = \new_[32652]_  & \new_[32641]_ ;
  assign \new_[858]_  = \new_[32630]_  & \new_[32619]_ ;
  assign \new_[859]_  = \new_[32608]_  & \new_[32597]_ ;
  assign \new_[860]_  = \new_[32586]_  & \new_[32575]_ ;
  assign \new_[861]_  = \new_[32564]_  & \new_[32553]_ ;
  assign \new_[862]_  = \new_[32542]_  & \new_[32531]_ ;
  assign \new_[863]_  = \new_[32520]_  & \new_[32509]_ ;
  assign \new_[864]_  = \new_[32498]_  & \new_[32487]_ ;
  assign \new_[865]_  = \new_[32476]_  & \new_[32465]_ ;
  assign \new_[866]_  = \new_[32454]_  & \new_[32443]_ ;
  assign \new_[867]_  = \new_[32432]_  & \new_[32421]_ ;
  assign \new_[868]_  = \new_[32410]_  & \new_[32399]_ ;
  assign \new_[869]_  = \new_[32388]_  & \new_[32377]_ ;
  assign \new_[870]_  = \new_[32366]_  & \new_[32355]_ ;
  assign \new_[871]_  = \new_[32344]_  & \new_[32333]_ ;
  assign \new_[872]_  = \new_[32322]_  & \new_[32311]_ ;
  assign \new_[873]_  = \new_[32300]_  & \new_[32289]_ ;
  assign \new_[874]_  = \new_[32278]_  & \new_[32267]_ ;
  assign \new_[875]_  = \new_[32256]_  & \new_[32245]_ ;
  assign \new_[876]_  = \new_[32234]_  & \new_[32223]_ ;
  assign \new_[877]_  = \new_[32212]_  & \new_[32201]_ ;
  assign \new_[878]_  = \new_[32190]_  & \new_[32179]_ ;
  assign \new_[879]_  = \new_[32168]_  & \new_[32157]_ ;
  assign \new_[880]_  = \new_[32146]_  & \new_[32135]_ ;
  assign \new_[881]_  = \new_[32124]_  & \new_[32113]_ ;
  assign \new_[882]_  = \new_[32102]_  & \new_[32091]_ ;
  assign \new_[883]_  = \new_[32080]_  & \new_[32069]_ ;
  assign \new_[884]_  = \new_[32058]_  & \new_[32047]_ ;
  assign \new_[885]_  = \new_[32036]_  & \new_[32025]_ ;
  assign \new_[886]_  = \new_[32014]_  & \new_[32003]_ ;
  assign \new_[887]_  = \new_[31992]_  & \new_[31981]_ ;
  assign \new_[888]_  = \new_[31970]_  & \new_[31959]_ ;
  assign \new_[889]_  = \new_[31948]_  & \new_[31937]_ ;
  assign \new_[890]_  = \new_[31926]_  & \new_[31915]_ ;
  assign \new_[891]_  = \new_[31904]_  & \new_[31893]_ ;
  assign \new_[892]_  = \new_[31882]_  & \new_[31871]_ ;
  assign \new_[893]_  = \new_[31860]_  & \new_[31849]_ ;
  assign \new_[894]_  = \new_[31838]_  & \new_[31827]_ ;
  assign \new_[895]_  = \new_[31816]_  & \new_[31805]_ ;
  assign \new_[896]_  = \new_[31794]_  & \new_[31783]_ ;
  assign \new_[897]_  = \new_[31772]_  & \new_[31761]_ ;
  assign \new_[898]_  = \new_[31750]_  & \new_[31739]_ ;
  assign \new_[899]_  = \new_[31728]_  & \new_[31717]_ ;
  assign \new_[900]_  = \new_[31706]_  & \new_[31695]_ ;
  assign \new_[901]_  = \new_[31684]_  & \new_[31673]_ ;
  assign \new_[902]_  = \new_[31662]_  & \new_[31651]_ ;
  assign \new_[903]_  = \new_[31640]_  & \new_[31629]_ ;
  assign \new_[904]_  = \new_[31618]_  & \new_[31607]_ ;
  assign \new_[905]_  = \new_[31596]_  & \new_[31585]_ ;
  assign \new_[906]_  = \new_[31574]_  & \new_[31563]_ ;
  assign \new_[907]_  = \new_[31552]_  & \new_[31541]_ ;
  assign \new_[908]_  = \new_[31530]_  & \new_[31519]_ ;
  assign \new_[909]_  = \new_[31508]_  & \new_[31497]_ ;
  assign \new_[910]_  = \new_[31486]_  & \new_[31475]_ ;
  assign \new_[911]_  = \new_[31464]_  & \new_[31453]_ ;
  assign \new_[912]_  = \new_[31442]_  & \new_[31431]_ ;
  assign \new_[913]_  = \new_[31420]_  & \new_[31409]_ ;
  assign \new_[914]_  = \new_[31398]_  & \new_[31387]_ ;
  assign \new_[915]_  = \new_[31376]_  & \new_[31365]_ ;
  assign \new_[916]_  = \new_[31354]_  & \new_[31343]_ ;
  assign \new_[917]_  = \new_[31332]_  & \new_[31321]_ ;
  assign \new_[918]_  = \new_[31310]_  & \new_[31299]_ ;
  assign \new_[919]_  = \new_[31288]_  & \new_[31277]_ ;
  assign \new_[920]_  = \new_[31266]_  & \new_[31255]_ ;
  assign \new_[921]_  = \new_[31244]_  & \new_[31233]_ ;
  assign \new_[922]_  = \new_[31222]_  & \new_[31211]_ ;
  assign \new_[923]_  = \new_[31200]_  & \new_[31189]_ ;
  assign \new_[924]_  = \new_[31178]_  & \new_[31167]_ ;
  assign \new_[925]_  = \new_[31156]_  & \new_[31145]_ ;
  assign \new_[926]_  = \new_[31134]_  & \new_[31123]_ ;
  assign \new_[927]_  = \new_[31112]_  & \new_[31101]_ ;
  assign \new_[928]_  = \new_[31090]_  & \new_[31079]_ ;
  assign \new_[929]_  = \new_[31068]_  & \new_[31057]_ ;
  assign \new_[930]_  = \new_[31046]_  & \new_[31035]_ ;
  assign \new_[931]_  = \new_[31024]_  & \new_[31013]_ ;
  assign \new_[932]_  = \new_[31002]_  & \new_[30991]_ ;
  assign \new_[933]_  = \new_[30980]_  & \new_[30969]_ ;
  assign \new_[934]_  = \new_[30958]_  & \new_[30947]_ ;
  assign \new_[935]_  = \new_[30936]_  & \new_[30925]_ ;
  assign \new_[936]_  = \new_[30914]_  & \new_[30903]_ ;
  assign \new_[937]_  = \new_[30892]_  & \new_[30881]_ ;
  assign \new_[938]_  = \new_[30870]_  & \new_[30859]_ ;
  assign \new_[939]_  = \new_[30848]_  & \new_[30837]_ ;
  assign \new_[940]_  = \new_[30826]_  & \new_[30815]_ ;
  assign \new_[941]_  = \new_[30804]_  & \new_[30793]_ ;
  assign \new_[942]_  = \new_[30782]_  & \new_[30771]_ ;
  assign \new_[943]_  = \new_[30760]_  & \new_[30749]_ ;
  assign \new_[944]_  = \new_[30738]_  & \new_[30727]_ ;
  assign \new_[945]_  = \new_[30716]_  & \new_[30705]_ ;
  assign \new_[946]_  = \new_[30694]_  & \new_[30683]_ ;
  assign \new_[947]_  = \new_[30672]_  & \new_[30661]_ ;
  assign \new_[948]_  = \new_[30650]_  & \new_[30639]_ ;
  assign \new_[949]_  = \new_[30628]_  & \new_[30617]_ ;
  assign \new_[950]_  = \new_[30606]_  & \new_[30595]_ ;
  assign \new_[951]_  = \new_[30584]_  & \new_[30573]_ ;
  assign \new_[952]_  = \new_[30562]_  & \new_[30551]_ ;
  assign \new_[953]_  = \new_[30540]_  & \new_[30529]_ ;
  assign \new_[954]_  = \new_[30518]_  & \new_[30507]_ ;
  assign \new_[955]_  = \new_[30496]_  & \new_[30485]_ ;
  assign \new_[956]_  = \new_[30474]_  & \new_[30463]_ ;
  assign \new_[957]_  = \new_[30452]_  & \new_[30441]_ ;
  assign \new_[958]_  = \new_[30430]_  & \new_[30419]_ ;
  assign \new_[959]_  = \new_[30408]_  & \new_[30397]_ ;
  assign \new_[960]_  = \new_[30386]_  & \new_[30375]_ ;
  assign \new_[961]_  = \new_[30364]_  & \new_[30353]_ ;
  assign \new_[962]_  = \new_[30342]_  & \new_[30331]_ ;
  assign \new_[963]_  = \new_[30320]_  & \new_[30309]_ ;
  assign \new_[964]_  = \new_[30298]_  & \new_[30287]_ ;
  assign \new_[965]_  = \new_[30276]_  & \new_[30265]_ ;
  assign \new_[966]_  = \new_[30254]_  & \new_[30243]_ ;
  assign \new_[967]_  = \new_[30232]_  & \new_[30221]_ ;
  assign \new_[968]_  = \new_[30210]_  & \new_[30199]_ ;
  assign \new_[969]_  = \new_[30188]_  & \new_[30177]_ ;
  assign \new_[970]_  = \new_[30166]_  & \new_[30155]_ ;
  assign \new_[971]_  = \new_[30144]_  & \new_[30133]_ ;
  assign \new_[972]_  = \new_[30122]_  & \new_[30111]_ ;
  assign \new_[973]_  = \new_[30100]_  & \new_[30089]_ ;
  assign \new_[974]_  = \new_[30078]_  & \new_[30067]_ ;
  assign \new_[975]_  = \new_[30056]_  & \new_[30045]_ ;
  assign \new_[976]_  = \new_[30034]_  & \new_[30023]_ ;
  assign \new_[977]_  = \new_[30012]_  & \new_[30001]_ ;
  assign \new_[978]_  = \new_[29990]_  & \new_[29979]_ ;
  assign \new_[979]_  = \new_[29968]_  & \new_[29957]_ ;
  assign \new_[980]_  = \new_[29946]_  & \new_[29935]_ ;
  assign \new_[981]_  = \new_[29924]_  & \new_[29913]_ ;
  assign \new_[982]_  = \new_[29902]_  & \new_[29891]_ ;
  assign \new_[983]_  = \new_[29880]_  & \new_[29869]_ ;
  assign \new_[984]_  = \new_[29858]_  & \new_[29847]_ ;
  assign \new_[985]_  = \new_[29836]_  & \new_[29825]_ ;
  assign \new_[986]_  = \new_[29814]_  & \new_[29803]_ ;
  assign \new_[987]_  = \new_[29792]_  & \new_[29781]_ ;
  assign \new_[988]_  = \new_[29770]_  & \new_[29759]_ ;
  assign \new_[989]_  = \new_[29748]_  & \new_[29737]_ ;
  assign \new_[990]_  = \new_[29726]_  & \new_[29715]_ ;
  assign \new_[991]_  = \new_[29704]_  & \new_[29693]_ ;
  assign \new_[992]_  = \new_[29682]_  & \new_[29671]_ ;
  assign \new_[993]_  = \new_[29660]_  & \new_[29649]_ ;
  assign \new_[994]_  = \new_[29638]_  & \new_[29627]_ ;
  assign \new_[995]_  = \new_[29616]_  & \new_[29605]_ ;
  assign \new_[996]_  = \new_[29594]_  & \new_[29583]_ ;
  assign \new_[997]_  = \new_[29572]_  & \new_[29561]_ ;
  assign \new_[998]_  = \new_[29550]_  & \new_[29539]_ ;
  assign \new_[999]_  = \new_[29528]_  & \new_[29517]_ ;
  assign \new_[1000]_  = \new_[29506]_  & \new_[29495]_ ;
  assign \new_[1001]_  = \new_[29484]_  & \new_[29473]_ ;
  assign \new_[1002]_  = \new_[29462]_  & \new_[29451]_ ;
  assign \new_[1003]_  = \new_[29440]_  & \new_[29429]_ ;
  assign \new_[1004]_  = \new_[29420]_  & \new_[29409]_ ;
  assign \new_[1005]_  = \new_[29400]_  & \new_[29389]_ ;
  assign \new_[1006]_  = \new_[29380]_  & \new_[29369]_ ;
  assign \new_[1007]_  = \new_[29360]_  & \new_[29349]_ ;
  assign \new_[1008]_  = \new_[29340]_  & \new_[29329]_ ;
  assign \new_[1009]_  = \new_[29320]_  & \new_[29309]_ ;
  assign \new_[1010]_  = \new_[29300]_  & \new_[29289]_ ;
  assign \new_[1011]_  = \new_[29280]_  & \new_[29269]_ ;
  assign \new_[1012]_  = \new_[29260]_  & \new_[29249]_ ;
  assign \new_[1013]_  = \new_[29240]_  & \new_[29229]_ ;
  assign \new_[1014]_  = \new_[29220]_  & \new_[29209]_ ;
  assign \new_[1015]_  = \new_[29200]_  & \new_[29189]_ ;
  assign \new_[1016]_  = \new_[29180]_  & \new_[29169]_ ;
  assign \new_[1017]_  = \new_[29160]_  & \new_[29149]_ ;
  assign \new_[1018]_  = \new_[29140]_  & \new_[29129]_ ;
  assign \new_[1019]_  = \new_[29120]_  & \new_[29109]_ ;
  assign \new_[1020]_  = \new_[29100]_  & \new_[29089]_ ;
  assign \new_[1021]_  = \new_[29080]_  & \new_[29069]_ ;
  assign \new_[1022]_  = \new_[29060]_  & \new_[29049]_ ;
  assign \new_[1023]_  = \new_[29040]_  & \new_[29029]_ ;
  assign \new_[1024]_  = \new_[29020]_  & \new_[29009]_ ;
  assign \new_[1025]_  = \new_[29000]_  & \new_[28989]_ ;
  assign \new_[1026]_  = \new_[28980]_  & \new_[28969]_ ;
  assign \new_[1027]_  = \new_[28960]_  & \new_[28949]_ ;
  assign \new_[1028]_  = \new_[28940]_  & \new_[28929]_ ;
  assign \new_[1029]_  = \new_[28920]_  & \new_[28909]_ ;
  assign \new_[1030]_  = \new_[28900]_  & \new_[28889]_ ;
  assign \new_[1031]_  = \new_[28880]_  & \new_[28869]_ ;
  assign \new_[1032]_  = \new_[28860]_  & \new_[28849]_ ;
  assign \new_[1033]_  = \new_[28840]_  & \new_[28829]_ ;
  assign \new_[1034]_  = \new_[28820]_  & \new_[28809]_ ;
  assign \new_[1035]_  = \new_[28800]_  & \new_[28789]_ ;
  assign \new_[1036]_  = \new_[28780]_  & \new_[28769]_ ;
  assign \new_[1037]_  = \new_[28760]_  & \new_[28749]_ ;
  assign \new_[1038]_  = \new_[28740]_  & \new_[28729]_ ;
  assign \new_[1039]_  = \new_[28720]_  & \new_[28709]_ ;
  assign \new_[1040]_  = \new_[28700]_  & \new_[28689]_ ;
  assign \new_[1041]_  = \new_[28680]_  & \new_[28669]_ ;
  assign \new_[1042]_  = \new_[28660]_  & \new_[28649]_ ;
  assign \new_[1043]_  = \new_[28640]_  & \new_[28629]_ ;
  assign \new_[1044]_  = \new_[28620]_  & \new_[28609]_ ;
  assign \new_[1045]_  = \new_[28600]_  & \new_[28589]_ ;
  assign \new_[1046]_  = \new_[28580]_  & \new_[28569]_ ;
  assign \new_[1047]_  = \new_[28560]_  & \new_[28549]_ ;
  assign \new_[1048]_  = \new_[28540]_  & \new_[28529]_ ;
  assign \new_[1049]_  = \new_[28520]_  & \new_[28509]_ ;
  assign \new_[1050]_  = \new_[28500]_  & \new_[28489]_ ;
  assign \new_[1051]_  = \new_[28480]_  & \new_[28469]_ ;
  assign \new_[1052]_  = \new_[28460]_  & \new_[28449]_ ;
  assign \new_[1053]_  = \new_[28440]_  & \new_[28429]_ ;
  assign \new_[1054]_  = \new_[28420]_  & \new_[28409]_ ;
  assign \new_[1055]_  = \new_[28400]_  & \new_[28389]_ ;
  assign \new_[1056]_  = \new_[28380]_  & \new_[28369]_ ;
  assign \new_[1057]_  = \new_[28360]_  & \new_[28349]_ ;
  assign \new_[1058]_  = \new_[28340]_  & \new_[28329]_ ;
  assign \new_[1059]_  = \new_[28320]_  & \new_[28309]_ ;
  assign \new_[1060]_  = \new_[28300]_  & \new_[28289]_ ;
  assign \new_[1061]_  = \new_[28280]_  & \new_[28269]_ ;
  assign \new_[1062]_  = \new_[28260]_  & \new_[28249]_ ;
  assign \new_[1063]_  = \new_[28240]_  & \new_[28229]_ ;
  assign \new_[1064]_  = \new_[28220]_  & \new_[28209]_ ;
  assign \new_[1065]_  = \new_[28200]_  & \new_[28189]_ ;
  assign \new_[1066]_  = \new_[28180]_  & \new_[28169]_ ;
  assign \new_[1067]_  = \new_[28160]_  & \new_[28149]_ ;
  assign \new_[1068]_  = \new_[28140]_  & \new_[28129]_ ;
  assign \new_[1069]_  = \new_[28120]_  & \new_[28109]_ ;
  assign \new_[1070]_  = \new_[28100]_  & \new_[28089]_ ;
  assign \new_[1071]_  = \new_[28080]_  & \new_[28069]_ ;
  assign \new_[1072]_  = \new_[28060]_  & \new_[28049]_ ;
  assign \new_[1073]_  = \new_[28040]_  & \new_[28029]_ ;
  assign \new_[1074]_  = \new_[28020]_  & \new_[28009]_ ;
  assign \new_[1075]_  = \new_[28000]_  & \new_[27989]_ ;
  assign \new_[1076]_  = \new_[27980]_  & \new_[27969]_ ;
  assign \new_[1077]_  = \new_[27960]_  & \new_[27949]_ ;
  assign \new_[1078]_  = \new_[27940]_  & \new_[27929]_ ;
  assign \new_[1079]_  = \new_[27920]_  & \new_[27909]_ ;
  assign \new_[1080]_  = \new_[27900]_  & \new_[27889]_ ;
  assign \new_[1081]_  = \new_[27880]_  & \new_[27869]_ ;
  assign \new_[1082]_  = \new_[27860]_  & \new_[27849]_ ;
  assign \new_[1083]_  = \new_[27840]_  & \new_[27829]_ ;
  assign \new_[1084]_  = \new_[27820]_  & \new_[27809]_ ;
  assign \new_[1085]_  = \new_[27800]_  & \new_[27789]_ ;
  assign \new_[1086]_  = \new_[27780]_  & \new_[27769]_ ;
  assign \new_[1087]_  = \new_[27760]_  & \new_[27749]_ ;
  assign \new_[1088]_  = \new_[27740]_  & \new_[27729]_ ;
  assign \new_[1089]_  = \new_[27720]_  & \new_[27709]_ ;
  assign \new_[1090]_  = \new_[27700]_  & \new_[27689]_ ;
  assign \new_[1091]_  = \new_[27680]_  & \new_[27669]_ ;
  assign \new_[1092]_  = \new_[27660]_  & \new_[27649]_ ;
  assign \new_[1093]_  = \new_[27640]_  & \new_[27629]_ ;
  assign \new_[1094]_  = \new_[27620]_  & \new_[27609]_ ;
  assign \new_[1095]_  = \new_[27600]_  & \new_[27589]_ ;
  assign \new_[1096]_  = \new_[27580]_  & \new_[27569]_ ;
  assign \new_[1097]_  = \new_[27560]_  & \new_[27549]_ ;
  assign \new_[1098]_  = \new_[27540]_  & \new_[27529]_ ;
  assign \new_[1099]_  = \new_[27520]_  & \new_[27509]_ ;
  assign \new_[1100]_  = \new_[27500]_  & \new_[27489]_ ;
  assign \new_[1101]_  = \new_[27480]_  & \new_[27469]_ ;
  assign \new_[1102]_  = \new_[27460]_  & \new_[27449]_ ;
  assign \new_[1103]_  = \new_[27440]_  & \new_[27429]_ ;
  assign \new_[1104]_  = \new_[27420]_  & \new_[27409]_ ;
  assign \new_[1105]_  = \new_[27400]_  & \new_[27389]_ ;
  assign \new_[1106]_  = \new_[27380]_  & \new_[27369]_ ;
  assign \new_[1107]_  = \new_[27360]_  & \new_[27349]_ ;
  assign \new_[1108]_  = \new_[27340]_  & \new_[27329]_ ;
  assign \new_[1109]_  = \new_[27320]_  & \new_[27309]_ ;
  assign \new_[1110]_  = \new_[27300]_  & \new_[27289]_ ;
  assign \new_[1111]_  = \new_[27280]_  & \new_[27269]_ ;
  assign \new_[1112]_  = \new_[27260]_  & \new_[27249]_ ;
  assign \new_[1113]_  = \new_[27240]_  & \new_[27229]_ ;
  assign \new_[1114]_  = \new_[27220]_  & \new_[27209]_ ;
  assign \new_[1115]_  = \new_[27200]_  & \new_[27189]_ ;
  assign \new_[1116]_  = \new_[27180]_  & \new_[27169]_ ;
  assign \new_[1117]_  = \new_[27160]_  & \new_[27149]_ ;
  assign \new_[1118]_  = \new_[27140]_  & \new_[27129]_ ;
  assign \new_[1119]_  = \new_[27120]_  & \new_[27109]_ ;
  assign \new_[1120]_  = \new_[27100]_  & \new_[27089]_ ;
  assign \new_[1121]_  = \new_[27080]_  & \new_[27069]_ ;
  assign \new_[1122]_  = \new_[27060]_  & \new_[27049]_ ;
  assign \new_[1123]_  = \new_[27040]_  & \new_[27029]_ ;
  assign \new_[1124]_  = \new_[27020]_  & \new_[27009]_ ;
  assign \new_[1125]_  = \new_[27000]_  & \new_[26989]_ ;
  assign \new_[1126]_  = \new_[26980]_  & \new_[26969]_ ;
  assign \new_[1127]_  = \new_[26960]_  & \new_[26949]_ ;
  assign \new_[1128]_  = \new_[26940]_  & \new_[26929]_ ;
  assign \new_[1129]_  = \new_[26920]_  & \new_[26909]_ ;
  assign \new_[1130]_  = \new_[26900]_  & \new_[26889]_ ;
  assign \new_[1131]_  = \new_[26880]_  & \new_[26869]_ ;
  assign \new_[1132]_  = \new_[26860]_  & \new_[26849]_ ;
  assign \new_[1133]_  = \new_[26840]_  & \new_[26829]_ ;
  assign \new_[1134]_  = \new_[26820]_  & \new_[26809]_ ;
  assign \new_[1135]_  = \new_[26800]_  & \new_[26789]_ ;
  assign \new_[1136]_  = \new_[26780]_  & \new_[26769]_ ;
  assign \new_[1137]_  = \new_[26760]_  & \new_[26749]_ ;
  assign \new_[1138]_  = \new_[26740]_  & \new_[26729]_ ;
  assign \new_[1139]_  = \new_[26720]_  & \new_[26709]_ ;
  assign \new_[1140]_  = \new_[26700]_  & \new_[26689]_ ;
  assign \new_[1141]_  = \new_[26680]_  & \new_[26669]_ ;
  assign \new_[1142]_  = \new_[26660]_  & \new_[26649]_ ;
  assign \new_[1143]_  = \new_[26640]_  & \new_[26629]_ ;
  assign \new_[1144]_  = \new_[26620]_  & \new_[26609]_ ;
  assign \new_[1145]_  = \new_[26600]_  & \new_[26589]_ ;
  assign \new_[1146]_  = \new_[26580]_  & \new_[26569]_ ;
  assign \new_[1147]_  = \new_[26560]_  & \new_[26549]_ ;
  assign \new_[1148]_  = \new_[26540]_  & \new_[26529]_ ;
  assign \new_[1149]_  = \new_[26520]_  & \new_[26509]_ ;
  assign \new_[1150]_  = \new_[26500]_  & \new_[26489]_ ;
  assign \new_[1151]_  = \new_[26480]_  & \new_[26469]_ ;
  assign \new_[1152]_  = \new_[26460]_  & \new_[26449]_ ;
  assign \new_[1153]_  = \new_[26440]_  & \new_[26429]_ ;
  assign \new_[1154]_  = \new_[26420]_  & \new_[26409]_ ;
  assign \new_[1155]_  = \new_[26400]_  & \new_[26389]_ ;
  assign \new_[1156]_  = \new_[26380]_  & \new_[26369]_ ;
  assign \new_[1157]_  = \new_[26360]_  & \new_[26349]_ ;
  assign \new_[1158]_  = \new_[26340]_  & \new_[26329]_ ;
  assign \new_[1159]_  = \new_[26320]_  & \new_[26309]_ ;
  assign \new_[1160]_  = \new_[26300]_  & \new_[26289]_ ;
  assign \new_[1161]_  = \new_[26280]_  & \new_[26269]_ ;
  assign \new_[1162]_  = \new_[26260]_  & \new_[26249]_ ;
  assign \new_[1163]_  = \new_[26240]_  & \new_[26229]_ ;
  assign \new_[1164]_  = \new_[26220]_  & \new_[26209]_ ;
  assign \new_[1165]_  = \new_[26200]_  & \new_[26189]_ ;
  assign \new_[1166]_  = \new_[26180]_  & \new_[26169]_ ;
  assign \new_[1167]_  = \new_[26160]_  & \new_[26149]_ ;
  assign \new_[1168]_  = \new_[26140]_  & \new_[26129]_ ;
  assign \new_[1169]_  = \new_[26120]_  & \new_[26109]_ ;
  assign \new_[1170]_  = \new_[26100]_  & \new_[26089]_ ;
  assign \new_[1171]_  = \new_[26080]_  & \new_[26069]_ ;
  assign \new_[1172]_  = \new_[26060]_  & \new_[26049]_ ;
  assign \new_[1173]_  = \new_[26040]_  & \new_[26029]_ ;
  assign \new_[1174]_  = \new_[26020]_  & \new_[26009]_ ;
  assign \new_[1175]_  = \new_[26000]_  & \new_[25989]_ ;
  assign \new_[1176]_  = \new_[25980]_  & \new_[25969]_ ;
  assign \new_[1177]_  = \new_[25960]_  & \new_[25949]_ ;
  assign \new_[1178]_  = \new_[25940]_  & \new_[25929]_ ;
  assign \new_[1179]_  = \new_[25920]_  & \new_[25909]_ ;
  assign \new_[1180]_  = \new_[25900]_  & \new_[25889]_ ;
  assign \new_[1181]_  = \new_[25880]_  & \new_[25869]_ ;
  assign \new_[1182]_  = \new_[25860]_  & \new_[25849]_ ;
  assign \new_[1183]_  = \new_[25840]_  & \new_[25829]_ ;
  assign \new_[1184]_  = \new_[25820]_  & \new_[25809]_ ;
  assign \new_[1185]_  = \new_[25800]_  & \new_[25789]_ ;
  assign \new_[1186]_  = \new_[25780]_  & \new_[25769]_ ;
  assign \new_[1187]_  = \new_[25760]_  & \new_[25749]_ ;
  assign \new_[1188]_  = \new_[25740]_  & \new_[25729]_ ;
  assign \new_[1189]_  = \new_[25720]_  & \new_[25709]_ ;
  assign \new_[1190]_  = \new_[25700]_  & \new_[25689]_ ;
  assign \new_[1191]_  = \new_[25680]_  & \new_[25669]_ ;
  assign \new_[1192]_  = \new_[25660]_  & \new_[25649]_ ;
  assign \new_[1193]_  = \new_[25640]_  & \new_[25629]_ ;
  assign \new_[1194]_  = \new_[25620]_  & \new_[25609]_ ;
  assign \new_[1195]_  = \new_[25600]_  & \new_[25589]_ ;
  assign \new_[1196]_  = \new_[25580]_  & \new_[25569]_ ;
  assign \new_[1197]_  = \new_[25560]_  & \new_[25549]_ ;
  assign \new_[1198]_  = \new_[25540]_  & \new_[25529]_ ;
  assign \new_[1199]_  = \new_[25520]_  & \new_[25509]_ ;
  assign \new_[1200]_  = \new_[25500]_  & \new_[25489]_ ;
  assign \new_[1201]_  = \new_[25480]_  & \new_[25469]_ ;
  assign \new_[1202]_  = \new_[25460]_  & \new_[25449]_ ;
  assign \new_[1203]_  = \new_[25440]_  & \new_[25429]_ ;
  assign \new_[1204]_  = \new_[25420]_  & \new_[25409]_ ;
  assign \new_[1205]_  = \new_[25400]_  & \new_[25389]_ ;
  assign \new_[1206]_  = \new_[25380]_  & \new_[25369]_ ;
  assign \new_[1207]_  = \new_[25360]_  & \new_[25349]_ ;
  assign \new_[1208]_  = \new_[25340]_  & \new_[25329]_ ;
  assign \new_[1209]_  = \new_[25320]_  & \new_[25309]_ ;
  assign \new_[1210]_  = \new_[25300]_  & \new_[25289]_ ;
  assign \new_[1211]_  = \new_[25280]_  & \new_[25269]_ ;
  assign \new_[1212]_  = \new_[25260]_  & \new_[25249]_ ;
  assign \new_[1213]_  = \new_[25240]_  & \new_[25229]_ ;
  assign \new_[1214]_  = \new_[25220]_  & \new_[25209]_ ;
  assign \new_[1215]_  = \new_[25200]_  & \new_[25189]_ ;
  assign \new_[1216]_  = \new_[25180]_  & \new_[25169]_ ;
  assign \new_[1217]_  = \new_[25160]_  & \new_[25149]_ ;
  assign \new_[1218]_  = \new_[25140]_  & \new_[25129]_ ;
  assign \new_[1219]_  = \new_[25120]_  & \new_[25109]_ ;
  assign \new_[1220]_  = \new_[25100]_  & \new_[25089]_ ;
  assign \new_[1221]_  = \new_[25080]_  & \new_[25069]_ ;
  assign \new_[1222]_  = \new_[25060]_  & \new_[25049]_ ;
  assign \new_[1223]_  = \new_[25040]_  & \new_[25029]_ ;
  assign \new_[1224]_  = \new_[25020]_  & \new_[25009]_ ;
  assign \new_[1225]_  = \new_[25000]_  & \new_[24989]_ ;
  assign \new_[1226]_  = \new_[24980]_  & \new_[24969]_ ;
  assign \new_[1227]_  = \new_[24960]_  & \new_[24949]_ ;
  assign \new_[1228]_  = \new_[24940]_  & \new_[24929]_ ;
  assign \new_[1229]_  = \new_[24920]_  & \new_[24909]_ ;
  assign \new_[1230]_  = \new_[24900]_  & \new_[24889]_ ;
  assign \new_[1231]_  = \new_[24880]_  & \new_[24869]_ ;
  assign \new_[1232]_  = \new_[24860]_  & \new_[24849]_ ;
  assign \new_[1233]_  = \new_[24840]_  & \new_[24829]_ ;
  assign \new_[1234]_  = \new_[24820]_  & \new_[24809]_ ;
  assign \new_[1235]_  = \new_[24800]_  & \new_[24789]_ ;
  assign \new_[1236]_  = \new_[24780]_  & \new_[24769]_ ;
  assign \new_[1237]_  = \new_[24760]_  & \new_[24749]_ ;
  assign \new_[1238]_  = \new_[24740]_  & \new_[24729]_ ;
  assign \new_[1239]_  = \new_[24720]_  & \new_[24709]_ ;
  assign \new_[1240]_  = \new_[24700]_  & \new_[24689]_ ;
  assign \new_[1241]_  = \new_[24680]_  & \new_[24669]_ ;
  assign \new_[1242]_  = \new_[24660]_  & \new_[24649]_ ;
  assign \new_[1243]_  = \new_[24640]_  & \new_[24629]_ ;
  assign \new_[1244]_  = \new_[24620]_  & \new_[24609]_ ;
  assign \new_[1245]_  = \new_[24600]_  & \new_[24589]_ ;
  assign \new_[1246]_  = \new_[24580]_  & \new_[24569]_ ;
  assign \new_[1247]_  = \new_[24560]_  & \new_[24549]_ ;
  assign \new_[1248]_  = \new_[24540]_  & \new_[24529]_ ;
  assign \new_[1249]_  = \new_[24520]_  & \new_[24509]_ ;
  assign \new_[1250]_  = \new_[24500]_  & \new_[24489]_ ;
  assign \new_[1251]_  = \new_[24480]_  & \new_[24469]_ ;
  assign \new_[1252]_  = \new_[24460]_  & \new_[24449]_ ;
  assign \new_[1253]_  = \new_[24440]_  & \new_[24429]_ ;
  assign \new_[1254]_  = \new_[24420]_  & \new_[24409]_ ;
  assign \new_[1255]_  = \new_[24400]_  & \new_[24389]_ ;
  assign \new_[1256]_  = \new_[24380]_  & \new_[24369]_ ;
  assign \new_[1257]_  = \new_[24360]_  & \new_[24349]_ ;
  assign \new_[1258]_  = \new_[24340]_  & \new_[24329]_ ;
  assign \new_[1259]_  = \new_[24320]_  & \new_[24309]_ ;
  assign \new_[1260]_  = \new_[24300]_  & \new_[24289]_ ;
  assign \new_[1261]_  = \new_[24280]_  & \new_[24269]_ ;
  assign \new_[1262]_  = \new_[24260]_  & \new_[24249]_ ;
  assign \new_[1263]_  = \new_[24240]_  & \new_[24229]_ ;
  assign \new_[1264]_  = \new_[24220]_  & \new_[24209]_ ;
  assign \new_[1265]_  = \new_[24200]_  & \new_[24189]_ ;
  assign \new_[1266]_  = \new_[24180]_  & \new_[24169]_ ;
  assign \new_[1267]_  = \new_[24160]_  & \new_[24149]_ ;
  assign \new_[1268]_  = \new_[24140]_  & \new_[24129]_ ;
  assign \new_[1269]_  = \new_[24120]_  & \new_[24109]_ ;
  assign \new_[1270]_  = \new_[24100]_  & \new_[24089]_ ;
  assign \new_[1271]_  = \new_[24080]_  & \new_[24069]_ ;
  assign \new_[1272]_  = \new_[24060]_  & \new_[24049]_ ;
  assign \new_[1273]_  = \new_[24040]_  & \new_[24029]_ ;
  assign \new_[1274]_  = \new_[24020]_  & \new_[24009]_ ;
  assign \new_[1275]_  = \new_[24000]_  & \new_[23989]_ ;
  assign \new_[1276]_  = \new_[23980]_  & \new_[23969]_ ;
  assign \new_[1277]_  = \new_[23960]_  & \new_[23949]_ ;
  assign \new_[1278]_  = \new_[23940]_  & \new_[23929]_ ;
  assign \new_[1279]_  = \new_[23920]_  & \new_[23909]_ ;
  assign \new_[1280]_  = \new_[23900]_  & \new_[23889]_ ;
  assign \new_[1281]_  = \new_[23880]_  & \new_[23869]_ ;
  assign \new_[1282]_  = \new_[23860]_  & \new_[23849]_ ;
  assign \new_[1283]_  = \new_[23840]_  & \new_[23829]_ ;
  assign \new_[1284]_  = \new_[23820]_  & \new_[23809]_ ;
  assign \new_[1285]_  = \new_[23800]_  & \new_[23789]_ ;
  assign \new_[1286]_  = \new_[23780]_  & \new_[23769]_ ;
  assign \new_[1287]_  = \new_[23760]_  & \new_[23749]_ ;
  assign \new_[1288]_  = \new_[23740]_  & \new_[23729]_ ;
  assign \new_[1289]_  = \new_[23720]_  & \new_[23709]_ ;
  assign \new_[1290]_  = \new_[23700]_  & \new_[23689]_ ;
  assign \new_[1291]_  = \new_[23680]_  & \new_[23669]_ ;
  assign \new_[1292]_  = \new_[23660]_  & \new_[23649]_ ;
  assign \new_[1293]_  = \new_[23640]_  & \new_[23629]_ ;
  assign \new_[1294]_  = \new_[23620]_  & \new_[23609]_ ;
  assign \new_[1295]_  = \new_[23600]_  & \new_[23589]_ ;
  assign \new_[1296]_  = \new_[23580]_  & \new_[23569]_ ;
  assign \new_[1297]_  = \new_[23560]_  & \new_[23549]_ ;
  assign \new_[1298]_  = \new_[23540]_  & \new_[23529]_ ;
  assign \new_[1299]_  = \new_[23520]_  & \new_[23509]_ ;
  assign \new_[1300]_  = \new_[23500]_  & \new_[23489]_ ;
  assign \new_[1301]_  = \new_[23480]_  & \new_[23469]_ ;
  assign \new_[1302]_  = \new_[23460]_  & \new_[23449]_ ;
  assign \new_[1303]_  = \new_[23440]_  & \new_[23429]_ ;
  assign \new_[1304]_  = \new_[23420]_  & \new_[23409]_ ;
  assign \new_[1305]_  = \new_[23400]_  & \new_[23389]_ ;
  assign \new_[1306]_  = \new_[23380]_  & \new_[23369]_ ;
  assign \new_[1307]_  = \new_[23360]_  & \new_[23349]_ ;
  assign \new_[1308]_  = \new_[23340]_  & \new_[23329]_ ;
  assign \new_[1309]_  = \new_[23320]_  & \new_[23309]_ ;
  assign \new_[1310]_  = \new_[23300]_  & \new_[23289]_ ;
  assign \new_[1311]_  = \new_[23280]_  & \new_[23269]_ ;
  assign \new_[1312]_  = \new_[23260]_  & \new_[23249]_ ;
  assign \new_[1313]_  = \new_[23240]_  & \new_[23229]_ ;
  assign \new_[1314]_  = \new_[23220]_  & \new_[23209]_ ;
  assign \new_[1315]_  = \new_[23200]_  & \new_[23189]_ ;
  assign \new_[1316]_  = \new_[23180]_  & \new_[23169]_ ;
  assign \new_[1317]_  = \new_[23160]_  & \new_[23149]_ ;
  assign \new_[1318]_  = \new_[23140]_  & \new_[23129]_ ;
  assign \new_[1319]_  = \new_[23120]_  & \new_[23109]_ ;
  assign \new_[1320]_  = \new_[23100]_  & \new_[23089]_ ;
  assign \new_[1321]_  = \new_[23080]_  & \new_[23069]_ ;
  assign \new_[1322]_  = \new_[23060]_  & \new_[23049]_ ;
  assign \new_[1323]_  = \new_[23040]_  & \new_[23029]_ ;
  assign \new_[1324]_  = \new_[23020]_  & \new_[23009]_ ;
  assign \new_[1325]_  = \new_[23000]_  & \new_[22989]_ ;
  assign \new_[1326]_  = \new_[22980]_  & \new_[22969]_ ;
  assign \new_[1327]_  = \new_[22960]_  & \new_[22949]_ ;
  assign \new_[1328]_  = \new_[22940]_  & \new_[22929]_ ;
  assign \new_[1329]_  = \new_[22920]_  & \new_[22909]_ ;
  assign \new_[1330]_  = \new_[22900]_  & \new_[22889]_ ;
  assign \new_[1331]_  = \new_[22880]_  & \new_[22869]_ ;
  assign \new_[1332]_  = \new_[22860]_  & \new_[22849]_ ;
  assign \new_[1333]_  = \new_[22840]_  & \new_[22829]_ ;
  assign \new_[1334]_  = \new_[22820]_  & \new_[22809]_ ;
  assign \new_[1335]_  = \new_[22800]_  & \new_[22789]_ ;
  assign \new_[1336]_  = \new_[22780]_  & \new_[22769]_ ;
  assign \new_[1337]_  = \new_[22760]_  & \new_[22749]_ ;
  assign \new_[1338]_  = \new_[22740]_  & \new_[22729]_ ;
  assign \new_[1339]_  = \new_[22720]_  & \new_[22711]_ ;
  assign \new_[1340]_  = \new_[22702]_  & \new_[22693]_ ;
  assign \new_[1341]_  = \new_[22684]_  & \new_[22675]_ ;
  assign \new_[1342]_  = \new_[22666]_  & \new_[22657]_ ;
  assign \new_[1343]_  = \new_[22648]_  & \new_[22639]_ ;
  assign \new_[1344]_  = \new_[22630]_  & \new_[22621]_ ;
  assign \new_[1345]_  = \new_[22612]_  & \new_[22603]_ ;
  assign \new_[1346]_  = \new_[22594]_  & \new_[22585]_ ;
  assign \new_[1347]_  = \new_[22576]_  & \new_[22567]_ ;
  assign \new_[1348]_  = \new_[22558]_  & \new_[22549]_ ;
  assign \new_[1349]_  = \new_[22540]_  & \new_[22531]_ ;
  assign \new_[1350]_  = \new_[22522]_  & \new_[22513]_ ;
  assign \new_[1351]_  = \new_[22504]_  & \new_[22495]_ ;
  assign \new_[1352]_  = \new_[22486]_  & \new_[22477]_ ;
  assign \new_[1353]_  = \new_[22468]_  & \new_[22459]_ ;
  assign \new_[1354]_  = \new_[22450]_  & \new_[22441]_ ;
  assign \new_[1355]_  = \new_[22432]_  & \new_[22423]_ ;
  assign \new_[1356]_  = \new_[22414]_  & \new_[22405]_ ;
  assign \new_[1357]_  = \new_[22396]_  & \new_[22387]_ ;
  assign \new_[1358]_  = \new_[22378]_  & \new_[22369]_ ;
  assign \new_[1359]_  = \new_[22360]_  & \new_[22351]_ ;
  assign \new_[1360]_  = \new_[22342]_  & \new_[22333]_ ;
  assign \new_[1361]_  = \new_[22324]_  & \new_[22315]_ ;
  assign \new_[1362]_  = \new_[22306]_  & \new_[22297]_ ;
  assign \new_[1363]_  = \new_[22288]_  & \new_[22279]_ ;
  assign \new_[1364]_  = \new_[22270]_  & \new_[22261]_ ;
  assign \new_[1365]_  = \new_[22252]_  & \new_[22243]_ ;
  assign \new_[1366]_  = \new_[22234]_  & \new_[22225]_ ;
  assign \new_[1367]_  = \new_[22216]_  & \new_[22207]_ ;
  assign \new_[1368]_  = \new_[22198]_  & \new_[22189]_ ;
  assign \new_[1369]_  = \new_[22180]_  & \new_[22171]_ ;
  assign \new_[1370]_  = \new_[22162]_  & \new_[22153]_ ;
  assign \new_[1371]_  = \new_[22144]_  & \new_[22135]_ ;
  assign \new_[1372]_  = \new_[22126]_  & \new_[22117]_ ;
  assign \new_[1373]_  = \new_[22108]_  & \new_[22099]_ ;
  assign \new_[1374]_  = \new_[22090]_  & \new_[22081]_ ;
  assign \new_[1375]_  = \new_[22072]_  & \new_[22063]_ ;
  assign \new_[1376]_  = \new_[22054]_  & \new_[22045]_ ;
  assign \new_[1377]_  = \new_[22036]_  & \new_[22027]_ ;
  assign \new_[1378]_  = \new_[22018]_  & \new_[22009]_ ;
  assign \new_[1379]_  = \new_[22000]_  & \new_[21991]_ ;
  assign \new_[1380]_  = \new_[21982]_  & \new_[21973]_ ;
  assign \new_[1381]_  = \new_[21964]_  & \new_[21955]_ ;
  assign \new_[1382]_  = \new_[21946]_  & \new_[21937]_ ;
  assign \new_[1383]_  = \new_[21928]_  & \new_[21919]_ ;
  assign \new_[1384]_  = \new_[21910]_  & \new_[21901]_ ;
  assign \new_[1385]_  = \new_[21892]_  & \new_[21883]_ ;
  assign \new_[1386]_  = \new_[21874]_  & \new_[21865]_ ;
  assign \new_[1387]_  = \new_[21856]_  & \new_[21847]_ ;
  assign \new_[1388]_  = \new_[21838]_  & \new_[21829]_ ;
  assign \new_[1389]_  = \new_[21820]_  & \new_[21811]_ ;
  assign \new_[1390]_  = \new_[21802]_  & \new_[21793]_ ;
  assign \new_[1391]_  = \new_[21784]_  & \new_[21775]_ ;
  assign \new_[1392]_  = \new_[21766]_  & \new_[21757]_ ;
  assign \new_[1393]_  = \new_[21748]_  & \new_[21739]_ ;
  assign \new_[1394]_  = \new_[21730]_  & \new_[21721]_ ;
  assign \new_[1395]_  = \new_[21712]_  & \new_[21703]_ ;
  assign \new_[1396]_  = \new_[21694]_  & \new_[21685]_ ;
  assign \new_[1397]_  = \new_[21676]_  & \new_[21667]_ ;
  assign \new_[1398]_  = \new_[21658]_  & \new_[21649]_ ;
  assign \new_[1399]_  = \new_[21640]_  & \new_[21631]_ ;
  assign \new_[1400]_  = \new_[21622]_  & \new_[21613]_ ;
  assign \new_[1401]_  = \new_[21604]_  & \new_[21595]_ ;
  assign \new_[1402]_  = \new_[21586]_  & \new_[21577]_ ;
  assign \new_[1403]_  = \new_[21568]_  & \new_[21559]_ ;
  assign \new_[1404]_  = \new_[21550]_  & \new_[21541]_ ;
  assign \new_[1405]_  = \new_[21532]_  & \new_[21523]_ ;
  assign \new_[1406]_  = \new_[21514]_  & \new_[21505]_ ;
  assign \new_[1407]_  = \new_[21496]_  & \new_[21487]_ ;
  assign \new_[1408]_  = \new_[21478]_  & \new_[21469]_ ;
  assign \new_[1409]_  = \new_[21460]_  & \new_[21451]_ ;
  assign \new_[1410]_  = \new_[21442]_  & \new_[21433]_ ;
  assign \new_[1411]_  = \new_[21424]_  & \new_[21415]_ ;
  assign \new_[1412]_  = \new_[21406]_  & \new_[21397]_ ;
  assign \new_[1413]_  = \new_[21388]_  & \new_[21379]_ ;
  assign \new_[1414]_  = \new_[21370]_  & \new_[21361]_ ;
  assign \new_[1415]_  = \new_[21352]_  & \new_[21343]_ ;
  assign \new_[1416]_  = \new_[21334]_  & \new_[21325]_ ;
  assign \new_[1417]_  = \new_[21316]_  & \new_[21307]_ ;
  assign \new_[1418]_  = \new_[21298]_  & \new_[21289]_ ;
  assign \new_[1419]_  = \new_[21280]_  & \new_[21271]_ ;
  assign \new_[1420]_  = \new_[21262]_  & \new_[21253]_ ;
  assign \new_[1421]_  = \new_[21244]_  & \new_[21235]_ ;
  assign \new_[1422]_  = \new_[21226]_  & \new_[21217]_ ;
  assign \new_[1423]_  = \new_[21208]_  & \new_[21199]_ ;
  assign \new_[1424]_  = \new_[21190]_  & \new_[21181]_ ;
  assign \new_[1425]_  = \new_[21172]_  & \new_[21163]_ ;
  assign \new_[1426]_  = \new_[21154]_  & \new_[21145]_ ;
  assign \new_[1427]_  = \new_[21136]_  & \new_[21127]_ ;
  assign \new_[1428]_  = \new_[21118]_  & \new_[21109]_ ;
  assign \new_[1429]_  = \new_[21100]_  & \new_[21091]_ ;
  assign \new_[1430]_  = \new_[21082]_  & \new_[21073]_ ;
  assign \new_[1431]_  = \new_[21064]_  & \new_[21055]_ ;
  assign \new_[1432]_  = \new_[21046]_  & \new_[21037]_ ;
  assign \new_[1433]_  = \new_[21028]_  & \new_[21019]_ ;
  assign \new_[1434]_  = \new_[21010]_  & \new_[21001]_ ;
  assign \new_[1435]_  = \new_[20992]_  & \new_[20983]_ ;
  assign \new_[1436]_  = \new_[20974]_  & \new_[20965]_ ;
  assign \new_[1437]_  = \new_[20956]_  & \new_[20947]_ ;
  assign \new_[1438]_  = \new_[20938]_  & \new_[20929]_ ;
  assign \new_[1439]_  = \new_[20920]_  & \new_[20911]_ ;
  assign \new_[1440]_  = \new_[20902]_  & \new_[20893]_ ;
  assign \new_[1441]_  = \new_[20884]_  & \new_[20875]_ ;
  assign \new_[1442]_  = \new_[20866]_  & \new_[20857]_ ;
  assign \new_[1443]_  = \new_[20848]_  & \new_[20839]_ ;
  assign \new_[1444]_  = \new_[20830]_  & \new_[20821]_ ;
  assign \new_[1445]_  = \new_[20812]_  & \new_[20803]_ ;
  assign \new_[1446]_  = \new_[20794]_  & \new_[20785]_ ;
  assign \new_[1447]_  = \new_[20776]_  & \new_[20767]_ ;
  assign \new_[1448]_  = \new_[20758]_  & \new_[20749]_ ;
  assign \new_[1449]_  = \new_[20740]_  & \new_[20731]_ ;
  assign \new_[1450]_  = \new_[20722]_  & \new_[20713]_ ;
  assign \new_[1451]_  = \new_[20704]_  & \new_[20695]_ ;
  assign \new_[1452]_  = \new_[20686]_  & \new_[20677]_ ;
  assign \new_[1453]_  = \new_[20668]_  & \new_[20659]_ ;
  assign \new_[1454]_  = \new_[20650]_  & \new_[20641]_ ;
  assign \new_[1455]_  = \new_[20632]_  & \new_[20623]_ ;
  assign \new_[1456]_  = \new_[20614]_  & \new_[20605]_ ;
  assign \new_[1457]_  = \new_[20596]_  & \new_[20587]_ ;
  assign \new_[1458]_  = \new_[20578]_  & \new_[20569]_ ;
  assign \new_[1459]_  = \new_[20560]_  & \new_[20551]_ ;
  assign \new_[1460]_  = \new_[20542]_  & \new_[20533]_ ;
  assign \new_[1461]_  = \new_[20524]_  & \new_[20515]_ ;
  assign \new_[1462]_  = \new_[20506]_  & \new_[20497]_ ;
  assign \new_[1463]_  = \new_[20488]_  & \new_[20479]_ ;
  assign \new_[1464]_  = \new_[20470]_  & \new_[20461]_ ;
  assign \new_[1465]_  = \new_[20452]_  & \new_[20443]_ ;
  assign \new_[1466]_  = \new_[20434]_  & \new_[20425]_ ;
  assign \new_[1467]_  = \new_[20416]_  & \new_[20407]_ ;
  assign \new_[1468]_  = \new_[20398]_  & \new_[20389]_ ;
  assign \new_[1469]_  = \new_[20380]_  & \new_[20371]_ ;
  assign \new_[1470]_  = \new_[20362]_  & \new_[20353]_ ;
  assign \new_[1471]_  = \new_[20344]_  & \new_[20335]_ ;
  assign \new_[1472]_  = \new_[20326]_  & \new_[20317]_ ;
  assign \new_[1473]_  = \new_[20308]_  & \new_[20299]_ ;
  assign \new_[1474]_  = \new_[20290]_  & \new_[20281]_ ;
  assign \new_[1475]_  = \new_[20272]_  & \new_[20263]_ ;
  assign \new_[1476]_  = \new_[20254]_  & \new_[20245]_ ;
  assign \new_[1477]_  = \new_[20236]_  & \new_[20227]_ ;
  assign \new_[1478]_  = \new_[20218]_  & \new_[20209]_ ;
  assign \new_[1479]_  = \new_[20200]_  & \new_[20191]_ ;
  assign \new_[1480]_  = \new_[20182]_  & \new_[20173]_ ;
  assign \new_[1481]_  = \new_[20164]_  & \new_[20155]_ ;
  assign \new_[1482]_  = \new_[20146]_  & \new_[20137]_ ;
  assign \new_[1483]_  = \new_[20128]_  & \new_[20119]_ ;
  assign \new_[1484]_  = \new_[20110]_  & \new_[20101]_ ;
  assign \new_[1485]_  = \new_[20092]_  & \new_[20083]_ ;
  assign \new_[1486]_  = \new_[20074]_  & \new_[20065]_ ;
  assign \new_[1487]_  = \new_[20056]_  & \new_[20047]_ ;
  assign \new_[1488]_  = \new_[20038]_  & \new_[20029]_ ;
  assign \new_[1489]_  = \new_[20020]_  & \new_[20011]_ ;
  assign \new_[1490]_  = \new_[20002]_  & \new_[19993]_ ;
  assign \new_[1491]_  = \new_[19984]_  & \new_[19975]_ ;
  assign \new_[1492]_  = \new_[19966]_  & \new_[19957]_ ;
  assign \new_[1493]_  = \new_[19948]_  & \new_[19939]_ ;
  assign \new_[1494]_  = \new_[19930]_  & \new_[19921]_ ;
  assign \new_[1495]_  = \new_[19912]_  & \new_[19903]_ ;
  assign \new_[1496]_  = \new_[19894]_  & \new_[19885]_ ;
  assign \new_[1497]_  = \new_[19876]_  & \new_[19867]_ ;
  assign \new_[1498]_  = \new_[19858]_  & \new_[19849]_ ;
  assign \new_[1499]_  = \new_[19840]_  & \new_[19831]_ ;
  assign \new_[1500]_  = \new_[19822]_  & \new_[19813]_ ;
  assign \new_[1501]_  = \new_[19804]_  & \new_[19795]_ ;
  assign \new_[1502]_  = \new_[19786]_  & \new_[19777]_ ;
  assign \new_[1503]_  = \new_[19768]_  & \new_[19759]_ ;
  assign \new_[1504]_  = \new_[19750]_  & \new_[19741]_ ;
  assign \new_[1505]_  = \new_[19732]_  & \new_[19723]_ ;
  assign \new_[1506]_  = \new_[19714]_  & \new_[19705]_ ;
  assign \new_[1507]_  = \new_[19696]_  & \new_[19687]_ ;
  assign \new_[1508]_  = \new_[19678]_  & \new_[19669]_ ;
  assign \new_[1509]_  = \new_[19660]_  & \new_[19651]_ ;
  assign \new_[1510]_  = \new_[19642]_  & \new_[19633]_ ;
  assign \new_[1511]_  = \new_[19624]_  & \new_[19615]_ ;
  assign \new_[1512]_  = \new_[19606]_  & \new_[19597]_ ;
  assign \new_[1513]_  = \new_[19588]_  & \new_[19579]_ ;
  assign \new_[1514]_  = \new_[19570]_  & \new_[19561]_ ;
  assign \new_[1515]_  = \new_[19552]_  & \new_[19543]_ ;
  assign \new_[1516]_  = \new_[19534]_  & \new_[19525]_ ;
  assign \new_[1517]_  = \new_[19516]_  & \new_[19507]_ ;
  assign \new_[1518]_  = \new_[19498]_  & \new_[19489]_ ;
  assign \new_[1519]_  = \new_[19480]_  & \new_[19471]_ ;
  assign \new_[1520]_  = \new_[19462]_  & \new_[19453]_ ;
  assign \new_[1521]_  = \new_[19444]_  & \new_[19435]_ ;
  assign \new_[1522]_  = \new_[19426]_  & \new_[19417]_ ;
  assign \new_[1523]_  = \new_[19408]_  & \new_[19399]_ ;
  assign \new_[1524]_  = \new_[19390]_  & \new_[19381]_ ;
  assign \new_[1525]_  = \new_[19372]_  & \new_[19363]_ ;
  assign \new_[1526]_  = \new_[19354]_  & \new_[19345]_ ;
  assign \new_[1527]_  = \new_[19336]_  & \new_[19327]_ ;
  assign \new_[1528]_  = \new_[19318]_  & \new_[19309]_ ;
  assign \new_[1529]_  = \new_[19300]_  & \new_[19291]_ ;
  assign \new_[1530]_  = \new_[19282]_  & \new_[19273]_ ;
  assign \new_[1531]_  = \new_[19264]_  & \new_[19255]_ ;
  assign \new_[1532]_  = \new_[19246]_  & \new_[19237]_ ;
  assign \new_[1533]_  = \new_[19228]_  & \new_[19219]_ ;
  assign \new_[1534]_  = \new_[19210]_  & \new_[19201]_ ;
  assign \new_[1535]_  = \new_[19192]_  & \new_[19183]_ ;
  assign \new_[1536]_  = \new_[19174]_  & \new_[19165]_ ;
  assign \new_[1537]_  = \new_[19156]_  & \new_[19147]_ ;
  assign \new_[1538]_  = \new_[19138]_  & \new_[19129]_ ;
  assign \new_[1539]_  = \new_[19120]_  & \new_[19111]_ ;
  assign \new_[1540]_  = \new_[19102]_  & \new_[19093]_ ;
  assign \new_[1541]_  = \new_[19084]_  & \new_[19075]_ ;
  assign \new_[1542]_  = \new_[19066]_  & \new_[19057]_ ;
  assign \new_[1543]_  = \new_[19048]_  & \new_[19039]_ ;
  assign \new_[1544]_  = \new_[19030]_  & \new_[19021]_ ;
  assign \new_[1545]_  = \new_[19012]_  & \new_[19003]_ ;
  assign \new_[1546]_  = \new_[18994]_  & \new_[18985]_ ;
  assign \new_[1547]_  = \new_[18976]_  & \new_[18967]_ ;
  assign \new_[1548]_  = \new_[18958]_  & \new_[18949]_ ;
  assign \new_[1549]_  = \new_[18940]_  & \new_[18931]_ ;
  assign \new_[1550]_  = \new_[18922]_  & \new_[18913]_ ;
  assign \new_[1551]_  = \new_[18904]_  & \new_[18895]_ ;
  assign \new_[1552]_  = \new_[18886]_  & \new_[18877]_ ;
  assign \new_[1553]_  = \new_[18868]_  & \new_[18859]_ ;
  assign \new_[1554]_  = \new_[18850]_  & \new_[18841]_ ;
  assign \new_[1555]_  = \new_[18832]_  & \new_[18823]_ ;
  assign \new_[1556]_  = \new_[18814]_  & \new_[18805]_ ;
  assign \new_[1557]_  = \new_[18796]_  & \new_[18787]_ ;
  assign \new_[1558]_  = \new_[18778]_  & \new_[18769]_ ;
  assign \new_[1559]_  = \new_[18760]_  & \new_[18751]_ ;
  assign \new_[1560]_  = \new_[18742]_  & \new_[18733]_ ;
  assign \new_[1561]_  = \new_[18724]_  & \new_[18715]_ ;
  assign \new_[1562]_  = \new_[18706]_  & \new_[18697]_ ;
  assign \new_[1563]_  = \new_[18688]_  & \new_[18679]_ ;
  assign \new_[1564]_  = \new_[18670]_  & \new_[18661]_ ;
  assign \new_[1565]_  = \new_[18652]_  & \new_[18643]_ ;
  assign \new_[1566]_  = \new_[18634]_  & \new_[18625]_ ;
  assign \new_[1567]_  = \new_[18616]_  & \new_[18607]_ ;
  assign \new_[1568]_  = \new_[18598]_  & \new_[18589]_ ;
  assign \new_[1569]_  = \new_[18580]_  & \new_[18571]_ ;
  assign \new_[1570]_  = \new_[18562]_  & \new_[18553]_ ;
  assign \new_[1571]_  = \new_[18544]_  & \new_[18535]_ ;
  assign \new_[1572]_  = \new_[18526]_  & \new_[18517]_ ;
  assign \new_[1573]_  = \new_[18508]_  & \new_[18499]_ ;
  assign \new_[1574]_  = \new_[18490]_  & \new_[18481]_ ;
  assign \new_[1575]_  = \new_[18472]_  & \new_[18463]_ ;
  assign \new_[1576]_  = \new_[18454]_  & \new_[18445]_ ;
  assign \new_[1577]_  = \new_[18436]_  & \new_[18427]_ ;
  assign \new_[1578]_  = \new_[18418]_  & \new_[18409]_ ;
  assign \new_[1579]_  = \new_[18400]_  & \new_[18391]_ ;
  assign \new_[1580]_  = \new_[18382]_  & \new_[18373]_ ;
  assign \new_[1581]_  = \new_[18364]_  & \new_[18355]_ ;
  assign \new_[1582]_  = \new_[18346]_  & \new_[18337]_ ;
  assign \new_[1583]_  = \new_[18328]_  & \new_[18319]_ ;
  assign \new_[1584]_  = \new_[18310]_  & \new_[18301]_ ;
  assign \new_[1585]_  = \new_[18292]_  & \new_[18283]_ ;
  assign \new_[1586]_  = \new_[18274]_  & \new_[18265]_ ;
  assign \new_[1587]_  = \new_[18256]_  & \new_[18247]_ ;
  assign \new_[1588]_  = \new_[18238]_  & \new_[18229]_ ;
  assign \new_[1589]_  = \new_[18220]_  & \new_[18211]_ ;
  assign \new_[1590]_  = \new_[18202]_  & \new_[18193]_ ;
  assign \new_[1591]_  = \new_[18184]_  & \new_[18175]_ ;
  assign \new_[1592]_  = \new_[18166]_  & \new_[18157]_ ;
  assign \new_[1593]_  = \new_[18148]_  & \new_[18139]_ ;
  assign \new_[1594]_  = \new_[18130]_  & \new_[18121]_ ;
  assign \new_[1595]_  = \new_[18112]_  & \new_[18103]_ ;
  assign \new_[1596]_  = \new_[18094]_  & \new_[18085]_ ;
  assign \new_[1597]_  = \new_[18076]_  & \new_[18067]_ ;
  assign \new_[1598]_  = \new_[18058]_  & \new_[18049]_ ;
  assign \new_[1599]_  = \new_[18040]_  & \new_[18031]_ ;
  assign \new_[1600]_  = \new_[18022]_  & \new_[18013]_ ;
  assign \new_[1601]_  = \new_[18004]_  & \new_[17995]_ ;
  assign \new_[1602]_  = \new_[17986]_  & \new_[17977]_ ;
  assign \new_[1603]_  = \new_[17968]_  & \new_[17959]_ ;
  assign \new_[1604]_  = \new_[17950]_  & \new_[17941]_ ;
  assign \new_[1605]_  = \new_[17932]_  & \new_[17923]_ ;
  assign \new_[1606]_  = \new_[17914]_  & \new_[17905]_ ;
  assign \new_[1607]_  = \new_[17896]_  & \new_[17887]_ ;
  assign \new_[1608]_  = \new_[17878]_  & \new_[17869]_ ;
  assign \new_[1609]_  = \new_[17860]_  & \new_[17851]_ ;
  assign \new_[1610]_  = \new_[17842]_  & \new_[17833]_ ;
  assign \new_[1611]_  = \new_[17824]_  & \new_[17815]_ ;
  assign \new_[1612]_  = \new_[17806]_  & \new_[17797]_ ;
  assign \new_[1613]_  = \new_[17788]_  & \new_[17779]_ ;
  assign \new_[1614]_  = \new_[17770]_  & \new_[17761]_ ;
  assign \new_[1615]_  = \new_[17752]_  & \new_[17743]_ ;
  assign \new_[1616]_  = \new_[17734]_  & \new_[17725]_ ;
  assign \new_[1617]_  = \new_[17716]_  & \new_[17707]_ ;
  assign \new_[1618]_  = \new_[17698]_  & \new_[17689]_ ;
  assign \new_[1619]_  = \new_[17680]_  & \new_[17671]_ ;
  assign \new_[1620]_  = \new_[17662]_  & \new_[17653]_ ;
  assign \new_[1621]_  = \new_[17644]_  & \new_[17635]_ ;
  assign \new_[1622]_  = \new_[17626]_  & \new_[17617]_ ;
  assign \new_[1623]_  = \new_[17608]_  & \new_[17599]_ ;
  assign \new_[1624]_  = \new_[17590]_  & \new_[17581]_ ;
  assign \new_[1625]_  = \new_[17572]_  & \new_[17563]_ ;
  assign \new_[1626]_  = \new_[17554]_  & \new_[17545]_ ;
  assign \new_[1627]_  = \new_[17536]_  & \new_[17527]_ ;
  assign \new_[1628]_  = \new_[17518]_  & \new_[17509]_ ;
  assign \new_[1629]_  = \new_[17500]_  & \new_[17491]_ ;
  assign \new_[1630]_  = \new_[17482]_  & \new_[17473]_ ;
  assign \new_[1631]_  = \new_[17464]_  & \new_[17455]_ ;
  assign \new_[1632]_  = \new_[17446]_  & \new_[17437]_ ;
  assign \new_[1633]_  = \new_[17428]_  & \new_[17419]_ ;
  assign \new_[1634]_  = \new_[17410]_  & \new_[17401]_ ;
  assign \new_[1635]_  = \new_[17392]_  & \new_[17383]_ ;
  assign \new_[1636]_  = \new_[17374]_  & \new_[17365]_ ;
  assign \new_[1637]_  = \new_[17356]_  & \new_[17347]_ ;
  assign \new_[1638]_  = \new_[17338]_  & \new_[17329]_ ;
  assign \new_[1639]_  = \new_[17320]_  & \new_[17311]_ ;
  assign \new_[1640]_  = \new_[17302]_  & \new_[17293]_ ;
  assign \new_[1641]_  = \new_[17284]_  & \new_[17275]_ ;
  assign \new_[1642]_  = \new_[17266]_  & \new_[17257]_ ;
  assign \new_[1643]_  = \new_[17248]_  & \new_[17239]_ ;
  assign \new_[1644]_  = \new_[17230]_  & \new_[17221]_ ;
  assign \new_[1645]_  = \new_[17212]_  & \new_[17203]_ ;
  assign \new_[1646]_  = \new_[17194]_  & \new_[17185]_ ;
  assign \new_[1647]_  = \new_[17176]_  & \new_[17167]_ ;
  assign \new_[1648]_  = \new_[17158]_  & \new_[17149]_ ;
  assign \new_[1649]_  = \new_[17140]_  & \new_[17131]_ ;
  assign \new_[1650]_  = \new_[17122]_  & \new_[17113]_ ;
  assign \new_[1651]_  = \new_[17104]_  & \new_[17095]_ ;
  assign \new_[1652]_  = \new_[17086]_  & \new_[17077]_ ;
  assign \new_[1653]_  = \new_[17068]_  & \new_[17059]_ ;
  assign \new_[1654]_  = \new_[17050]_  & \new_[17041]_ ;
  assign \new_[1655]_  = \new_[17032]_  & \new_[17023]_ ;
  assign \new_[1656]_  = \new_[17014]_  & \new_[17005]_ ;
  assign \new_[1657]_  = \new_[16996]_  & \new_[16987]_ ;
  assign \new_[1658]_  = \new_[16978]_  & \new_[16969]_ ;
  assign \new_[1659]_  = \new_[16960]_  & \new_[16951]_ ;
  assign \new_[1660]_  = \new_[16942]_  & \new_[16933]_ ;
  assign \new_[1661]_  = \new_[16924]_  & \new_[16915]_ ;
  assign \new_[1662]_  = \new_[16906]_  & \new_[16897]_ ;
  assign \new_[1663]_  = \new_[16888]_  & \new_[16879]_ ;
  assign \new_[1664]_  = \new_[16870]_  & \new_[16861]_ ;
  assign \new_[1665]_  = \new_[16852]_  & \new_[16843]_ ;
  assign \new_[1666]_  = \new_[16834]_  & \new_[16825]_ ;
  assign \new_[1667]_  = \new_[16816]_  & \new_[16807]_ ;
  assign \new_[1668]_  = \new_[16798]_  & \new_[16789]_ ;
  assign \new_[1669]_  = \new_[16780]_  & \new_[16771]_ ;
  assign \new_[1670]_  = \new_[16762]_  & \new_[16753]_ ;
  assign \new_[1671]_  = \new_[16744]_  & \new_[16735]_ ;
  assign \new_[1672]_  = \new_[16726]_  & \new_[16717]_ ;
  assign \new_[1673]_  = \new_[16708]_  & \new_[16699]_ ;
  assign \new_[1674]_  = \new_[16690]_  & \new_[16681]_ ;
  assign \new_[1675]_  = \new_[16672]_  & \new_[16663]_ ;
  assign \new_[1676]_  = \new_[16654]_  & \new_[16645]_ ;
  assign \new_[1677]_  = \new_[16636]_  & \new_[16627]_ ;
  assign \new_[1678]_  = \new_[16618]_  & \new_[16609]_ ;
  assign \new_[1679]_  = \new_[16600]_  & \new_[16591]_ ;
  assign \new_[1680]_  = \new_[16582]_  & \new_[16573]_ ;
  assign \new_[1681]_  = \new_[16564]_  & \new_[16555]_ ;
  assign \new_[1682]_  = \new_[16546]_  & \new_[16537]_ ;
  assign \new_[1683]_  = \new_[16528]_  & \new_[16519]_ ;
  assign \new_[1684]_  = \new_[16510]_  & \new_[16501]_ ;
  assign \new_[1685]_  = \new_[16492]_  & \new_[16483]_ ;
  assign \new_[1686]_  = \new_[16474]_  & \new_[16465]_ ;
  assign \new_[1687]_  = \new_[16456]_  & \new_[16447]_ ;
  assign \new_[1688]_  = \new_[16438]_  & \new_[16429]_ ;
  assign \new_[1689]_  = \new_[16420]_  & \new_[16411]_ ;
  assign \new_[1690]_  = \new_[16402]_  & \new_[16393]_ ;
  assign \new_[1691]_  = \new_[16384]_  & \new_[16375]_ ;
  assign \new_[1692]_  = \new_[16366]_  & \new_[16357]_ ;
  assign \new_[1693]_  = \new_[16348]_  & \new_[16339]_ ;
  assign \new_[1694]_  = \new_[16330]_  & \new_[16321]_ ;
  assign \new_[1695]_  = \new_[16312]_  & \new_[16303]_ ;
  assign \new_[1696]_  = \new_[16294]_  & \new_[16285]_ ;
  assign \new_[1697]_  = \new_[16276]_  & \new_[16267]_ ;
  assign \new_[1698]_  = \new_[16258]_  & \new_[16249]_ ;
  assign \new_[1699]_  = \new_[16240]_  & \new_[16231]_ ;
  assign \new_[1700]_  = \new_[16222]_  & \new_[16213]_ ;
  assign \new_[1701]_  = \new_[16204]_  & \new_[16195]_ ;
  assign \new_[1702]_  = \new_[16186]_  & \new_[16177]_ ;
  assign \new_[1703]_  = \new_[16168]_  & \new_[16159]_ ;
  assign \new_[1704]_  = \new_[16150]_  & \new_[16141]_ ;
  assign \new_[1705]_  = \new_[16132]_  & \new_[16123]_ ;
  assign \new_[1706]_  = \new_[16114]_  & \new_[16105]_ ;
  assign \new_[1707]_  = \new_[16096]_  & \new_[16087]_ ;
  assign \new_[1708]_  = \new_[16078]_  & \new_[16069]_ ;
  assign \new_[1709]_  = \new_[16060]_  & \new_[16051]_ ;
  assign \new_[1710]_  = \new_[16042]_  & \new_[16033]_ ;
  assign \new_[1711]_  = \new_[16024]_  & \new_[16015]_ ;
  assign \new_[1712]_  = \new_[16006]_  & \new_[15997]_ ;
  assign \new_[1713]_  = \new_[15988]_  & \new_[15979]_ ;
  assign \new_[1714]_  = \new_[15970]_  & \new_[15961]_ ;
  assign \new_[1715]_  = \new_[15952]_  & \new_[15943]_ ;
  assign \new_[1716]_  = \new_[15934]_  & \new_[15925]_ ;
  assign \new_[1717]_  = \new_[15916]_  & \new_[15907]_ ;
  assign \new_[1718]_  = \new_[15898]_  & \new_[15889]_ ;
  assign \new_[1719]_  = \new_[15880]_  & \new_[15871]_ ;
  assign \new_[1720]_  = \new_[15862]_  & \new_[15853]_ ;
  assign \new_[1721]_  = \new_[15844]_  & \new_[15835]_ ;
  assign \new_[1722]_  = \new_[15826]_  & \new_[15817]_ ;
  assign \new_[1723]_  = \new_[15808]_  & \new_[15799]_ ;
  assign \new_[1724]_  = \new_[15790]_  & \new_[15781]_ ;
  assign \new_[1725]_  = \new_[15772]_  & \new_[15763]_ ;
  assign \new_[1726]_  = \new_[15754]_  & \new_[15745]_ ;
  assign \new_[1727]_  = \new_[15736]_  & \new_[15727]_ ;
  assign \new_[1728]_  = \new_[15718]_  & \new_[15709]_ ;
  assign \new_[1729]_  = \new_[15700]_  & \new_[15691]_ ;
  assign \new_[1730]_  = \new_[15682]_  & \new_[15673]_ ;
  assign \new_[1731]_  = \new_[15664]_  & \new_[15655]_ ;
  assign \new_[1732]_  = \new_[15646]_  & \new_[15637]_ ;
  assign \new_[1733]_  = \new_[15628]_  & \new_[15619]_ ;
  assign \new_[1734]_  = \new_[15610]_  & \new_[15601]_ ;
  assign \new_[1735]_  = \new_[15592]_  & \new_[15583]_ ;
  assign \new_[1736]_  = \new_[15574]_  & \new_[15565]_ ;
  assign \new_[1737]_  = \new_[15556]_  & \new_[15547]_ ;
  assign \new_[1738]_  = \new_[15538]_  & \new_[15529]_ ;
  assign \new_[1739]_  = \new_[15520]_  & \new_[15511]_ ;
  assign \new_[1740]_  = \new_[15502]_  & \new_[15493]_ ;
  assign \new_[1741]_  = \new_[15484]_  & \new_[15475]_ ;
  assign \new_[1742]_  = \new_[15466]_  & \new_[15457]_ ;
  assign \new_[1743]_  = \new_[15448]_  & \new_[15439]_ ;
  assign \new_[1744]_  = \new_[15430]_  & \new_[15421]_ ;
  assign \new_[1745]_  = \new_[15412]_  & \new_[15403]_ ;
  assign \new_[1746]_  = \new_[15394]_  & \new_[15385]_ ;
  assign \new_[1747]_  = \new_[15376]_  & \new_[15367]_ ;
  assign \new_[1748]_  = \new_[15358]_  & \new_[15349]_ ;
  assign \new_[1749]_  = \new_[15340]_  & \new_[15331]_ ;
  assign \new_[1750]_  = \new_[15322]_  & \new_[15313]_ ;
  assign \new_[1751]_  = \new_[15304]_  & \new_[15295]_ ;
  assign \new_[1752]_  = \new_[15286]_  & \new_[15277]_ ;
  assign \new_[1753]_  = \new_[15268]_  & \new_[15259]_ ;
  assign \new_[1754]_  = \new_[15250]_  & \new_[15241]_ ;
  assign \new_[1755]_  = \new_[15232]_  & \new_[15223]_ ;
  assign \new_[1756]_  = \new_[15216]_  & \new_[15207]_ ;
  assign \new_[1757]_  = \new_[15200]_  & \new_[15191]_ ;
  assign \new_[1758]_  = \new_[15184]_  & \new_[15175]_ ;
  assign \new_[1759]_  = \new_[15168]_  & \new_[15159]_ ;
  assign \new_[1760]_  = \new_[15152]_  & \new_[15143]_ ;
  assign \new_[1761]_  = \new_[15136]_  & \new_[15127]_ ;
  assign \new_[1762]_  = \new_[15120]_  & \new_[15111]_ ;
  assign \new_[1763]_  = \new_[15104]_  & \new_[15095]_ ;
  assign \new_[1764]_  = \new_[15088]_  & \new_[15079]_ ;
  assign \new_[1765]_  = \new_[15072]_  & \new_[15063]_ ;
  assign \new_[1766]_  = \new_[15056]_  & \new_[15047]_ ;
  assign \new_[1767]_  = \new_[15040]_  & \new_[15031]_ ;
  assign \new_[1768]_  = \new_[15024]_  & \new_[15015]_ ;
  assign \new_[1769]_  = \new_[15008]_  & \new_[14999]_ ;
  assign \new_[1770]_  = \new_[14992]_  & \new_[14983]_ ;
  assign \new_[1771]_  = \new_[14976]_  & \new_[14967]_ ;
  assign \new_[1772]_  = \new_[14960]_  & \new_[14951]_ ;
  assign \new_[1773]_  = \new_[14944]_  & \new_[14935]_ ;
  assign \new_[1774]_  = \new_[14928]_  & \new_[14919]_ ;
  assign \new_[1775]_  = \new_[14912]_  & \new_[14903]_ ;
  assign \new_[1776]_  = \new_[14896]_  & \new_[14887]_ ;
  assign \new_[1777]_  = \new_[14880]_  & \new_[14871]_ ;
  assign \new_[1778]_  = \new_[14864]_  & \new_[14855]_ ;
  assign \new_[1779]_  = \new_[14848]_  & \new_[14839]_ ;
  assign \new_[1780]_  = \new_[14832]_  & \new_[14823]_ ;
  assign \new_[1781]_  = \new_[14816]_  & \new_[14807]_ ;
  assign \new_[1782]_  = \new_[14800]_  & \new_[14791]_ ;
  assign \new_[1783]_  = \new_[14784]_  & \new_[14775]_ ;
  assign \new_[1784]_  = \new_[14768]_  & \new_[14759]_ ;
  assign \new_[1785]_  = \new_[14752]_  & \new_[14743]_ ;
  assign \new_[1786]_  = \new_[14736]_  & \new_[14727]_ ;
  assign \new_[1787]_  = \new_[14720]_  & \new_[14711]_ ;
  assign \new_[1788]_  = \new_[14704]_  & \new_[14695]_ ;
  assign \new_[1789]_  = \new_[14688]_  & \new_[14679]_ ;
  assign \new_[1790]_  = \new_[14672]_  & \new_[14663]_ ;
  assign \new_[1791]_  = \new_[14656]_  & \new_[14647]_ ;
  assign \new_[1792]_  = \new_[14640]_  & \new_[14631]_ ;
  assign \new_[1793]_  = \new_[14624]_  & \new_[14615]_ ;
  assign \new_[1794]_  = \new_[14608]_  & \new_[14599]_ ;
  assign \new_[1795]_  = \new_[14592]_  & \new_[14583]_ ;
  assign \new_[1796]_  = \new_[14576]_  & \new_[14567]_ ;
  assign \new_[1797]_  = \new_[14560]_  & \new_[14551]_ ;
  assign \new_[1798]_  = \new_[14544]_  & \new_[14535]_ ;
  assign \new_[1799]_  = \new_[14528]_  & \new_[14519]_ ;
  assign \new_[1800]_  = \new_[14512]_  & \new_[14503]_ ;
  assign \new_[1801]_  = \new_[14496]_  & \new_[14487]_ ;
  assign \new_[1802]_  = \new_[14480]_  & \new_[14471]_ ;
  assign \new_[1803]_  = \new_[14464]_  & \new_[14455]_ ;
  assign \new_[1804]_  = \new_[14448]_  & \new_[14439]_ ;
  assign \new_[1805]_  = \new_[14432]_  & \new_[14423]_ ;
  assign \new_[1806]_  = \new_[14416]_  & \new_[14407]_ ;
  assign \new_[1807]_  = \new_[14400]_  & \new_[14391]_ ;
  assign \new_[1808]_  = \new_[14384]_  & \new_[14375]_ ;
  assign \new_[1809]_  = \new_[14368]_  & \new_[14359]_ ;
  assign \new_[1810]_  = \new_[14352]_  & \new_[14343]_ ;
  assign \new_[1811]_  = \new_[14336]_  & \new_[14327]_ ;
  assign \new_[1812]_  = \new_[14320]_  & \new_[14311]_ ;
  assign \new_[1813]_  = \new_[14304]_  & \new_[14295]_ ;
  assign \new_[1814]_  = \new_[14288]_  & \new_[14279]_ ;
  assign \new_[1815]_  = \new_[14272]_  & \new_[14263]_ ;
  assign \new_[1816]_  = \new_[14256]_  & \new_[14247]_ ;
  assign \new_[1817]_  = \new_[14240]_  & \new_[14231]_ ;
  assign \new_[1818]_  = \new_[14224]_  & \new_[14215]_ ;
  assign \new_[1819]_  = \new_[14208]_  & \new_[14199]_ ;
  assign \new_[1820]_  = \new_[14192]_  & \new_[14183]_ ;
  assign \new_[1821]_  = \new_[14176]_  & \new_[14167]_ ;
  assign \new_[1822]_  = \new_[14160]_  & \new_[14151]_ ;
  assign \new_[1823]_  = \new_[14144]_  & \new_[14135]_ ;
  assign \new_[1824]_  = \new_[14128]_  & \new_[14119]_ ;
  assign \new_[1825]_  = \new_[14112]_  & \new_[14103]_ ;
  assign \new_[1826]_  = \new_[14096]_  & \new_[14087]_ ;
  assign \new_[1827]_  = \new_[14080]_  & \new_[14071]_ ;
  assign \new_[1828]_  = \new_[14064]_  & \new_[14055]_ ;
  assign \new_[1829]_  = \new_[14048]_  & \new_[14039]_ ;
  assign \new_[1830]_  = \new_[14032]_  & \new_[14023]_ ;
  assign \new_[1831]_  = \new_[14016]_  & \new_[14007]_ ;
  assign \new_[1832]_  = \new_[14000]_  & \new_[13991]_ ;
  assign \new_[1833]_  = \new_[13984]_  & \new_[13975]_ ;
  assign \new_[1834]_  = \new_[13968]_  & \new_[13959]_ ;
  assign \new_[1835]_  = \new_[13952]_  & \new_[13943]_ ;
  assign \new_[1836]_  = \new_[13936]_  & \new_[13927]_ ;
  assign \new_[1837]_  = \new_[13920]_  & \new_[13911]_ ;
  assign \new_[1838]_  = \new_[13904]_  & \new_[13895]_ ;
  assign \new_[1839]_  = \new_[13888]_  & \new_[13879]_ ;
  assign \new_[1840]_  = \new_[13872]_  & \new_[13863]_ ;
  assign \new_[1841]_  = \new_[13856]_  & \new_[13847]_ ;
  assign \new_[1842]_  = \new_[13840]_  & \new_[13831]_ ;
  assign \new_[1843]_  = \new_[13824]_  & \new_[13815]_ ;
  assign \new_[1844]_  = \new_[13808]_  & \new_[13799]_ ;
  assign \new_[1845]_  = \new_[13792]_  & \new_[13783]_ ;
  assign \new_[1846]_  = \new_[13776]_  & \new_[13767]_ ;
  assign \new_[1847]_  = \new_[13760]_  & \new_[13751]_ ;
  assign \new_[1848]_  = \new_[13744]_  & \new_[13735]_ ;
  assign \new_[1849]_  = \new_[13728]_  & \new_[13719]_ ;
  assign \new_[1850]_  = \new_[13712]_  & \new_[13703]_ ;
  assign \new_[1851]_  = \new_[13696]_  & \new_[13687]_ ;
  assign \new_[1852]_  = \new_[13680]_  & \new_[13671]_ ;
  assign \new_[1853]_  = \new_[13664]_  & \new_[13655]_ ;
  assign \new_[1854]_  = \new_[13648]_  & \new_[13639]_ ;
  assign \new_[1855]_  = \new_[13632]_  & \new_[13623]_ ;
  assign \new_[1856]_  = \new_[13616]_  & \new_[13607]_ ;
  assign \new_[1857]_  = \new_[13600]_  & \new_[13591]_ ;
  assign \new_[1858]_  = \new_[13584]_  & \new_[13575]_ ;
  assign \new_[1859]_  = \new_[13568]_  & \new_[13559]_ ;
  assign \new_[1860]_  = \new_[13552]_  & \new_[13543]_ ;
  assign \new_[1861]_  = \new_[13536]_  & \new_[13527]_ ;
  assign \new_[1862]_  = \new_[13520]_  & \new_[13511]_ ;
  assign \new_[1863]_  = \new_[13504]_  & \new_[13495]_ ;
  assign \new_[1864]_  = \new_[13488]_  & \new_[13479]_ ;
  assign \new_[1865]_  = \new_[13472]_  & \new_[13463]_ ;
  assign \new_[1866]_  = \new_[13456]_  & \new_[13447]_ ;
  assign \new_[1867]_  = \new_[13440]_  & \new_[13431]_ ;
  assign \new_[1868]_  = \new_[13424]_  & \new_[13415]_ ;
  assign \new_[1869]_  = \new_[13408]_  & \new_[13399]_ ;
  assign \new_[1870]_  = \new_[13392]_  & \new_[13383]_ ;
  assign \new_[1871]_  = \new_[13376]_  & \new_[13367]_ ;
  assign \new_[1872]_  = \new_[13360]_  & \new_[13351]_ ;
  assign \new_[1873]_  = \new_[13344]_  & \new_[13335]_ ;
  assign \new_[1874]_  = \new_[13328]_  & \new_[13319]_ ;
  assign \new_[1875]_  = \new_[13312]_  & \new_[13303]_ ;
  assign \new_[1876]_  = \new_[13296]_  & \new_[13287]_ ;
  assign \new_[1877]_  = \new_[13280]_  & \new_[13271]_ ;
  assign \new_[1878]_  = \new_[13264]_  & \new_[13255]_ ;
  assign \new_[1879]_  = \new_[13248]_  & \new_[13239]_ ;
  assign \new_[1880]_  = \new_[13232]_  & \new_[13223]_ ;
  assign \new_[1881]_  = \new_[13216]_  & \new_[13207]_ ;
  assign \new_[1882]_  = \new_[13200]_  & \new_[13191]_ ;
  assign \new_[1883]_  = \new_[13184]_  & \new_[13175]_ ;
  assign \new_[1884]_  = \new_[13168]_  & \new_[13159]_ ;
  assign \new_[1885]_  = \new_[13152]_  & \new_[13143]_ ;
  assign \new_[1886]_  = \new_[13136]_  & \new_[13127]_ ;
  assign \new_[1887]_  = \new_[13120]_  & \new_[13111]_ ;
  assign \new_[1888]_  = \new_[13104]_  & \new_[13095]_ ;
  assign \new_[1889]_  = \new_[13088]_  & \new_[13079]_ ;
  assign \new_[1890]_  = \new_[13072]_  & \new_[13063]_ ;
  assign \new_[1891]_  = \new_[13056]_  & \new_[13047]_ ;
  assign \new_[1892]_  = \new_[13040]_  & \new_[13031]_ ;
  assign \new_[1893]_  = \new_[13024]_  & \new_[13015]_ ;
  assign \new_[1894]_  = \new_[13008]_  & \new_[12999]_ ;
  assign \new_[1895]_  = \new_[12992]_  & \new_[12983]_ ;
  assign \new_[1896]_  = \new_[12976]_  & \new_[12967]_ ;
  assign \new_[1897]_  = \new_[12960]_  & \new_[12951]_ ;
  assign \new_[1898]_  = \new_[12944]_  & \new_[12935]_ ;
  assign \new_[1899]_  = \new_[12928]_  & \new_[12919]_ ;
  assign \new_[1900]_  = \new_[12912]_  & \new_[12903]_ ;
  assign \new_[1901]_  = \new_[12896]_  & \new_[12887]_ ;
  assign \new_[1902]_  = \new_[12880]_  & \new_[12871]_ ;
  assign \new_[1903]_  = \new_[12864]_  & \new_[12855]_ ;
  assign \new_[1904]_  = \new_[12848]_  & \new_[12839]_ ;
  assign \new_[1905]_  = \new_[12832]_  & \new_[12823]_ ;
  assign \new_[1906]_  = \new_[12816]_  & \new_[12807]_ ;
  assign \new_[1907]_  = \new_[12800]_  & \new_[12791]_ ;
  assign \new_[1908]_  = \new_[12784]_  & \new_[12775]_ ;
  assign \new_[1909]_  = \new_[12768]_  & \new_[12759]_ ;
  assign \new_[1910]_  = \new_[12752]_  & \new_[12743]_ ;
  assign \new_[1911]_  = \new_[12736]_  & \new_[12727]_ ;
  assign \new_[1912]_  = \new_[12720]_  & \new_[12711]_ ;
  assign \new_[1913]_  = \new_[12704]_  & \new_[12695]_ ;
  assign \new_[1914]_  = \new_[12688]_  & \new_[12679]_ ;
  assign \new_[1915]_  = \new_[12672]_  & \new_[12663]_ ;
  assign \new_[1916]_  = \new_[12656]_  & \new_[12647]_ ;
  assign \new_[1917]_  = \new_[12640]_  & \new_[12631]_ ;
  assign \new_[1918]_  = \new_[12624]_  & \new_[12615]_ ;
  assign \new_[1919]_  = \new_[12608]_  & \new_[12599]_ ;
  assign \new_[1920]_  = \new_[12592]_  & \new_[12583]_ ;
  assign \new_[1921]_  = \new_[12576]_  & \new_[12567]_ ;
  assign \new_[1922]_  = \new_[12560]_  & \new_[12551]_ ;
  assign \new_[1923]_  = \new_[12544]_  & \new_[12535]_ ;
  assign \new_[1924]_  = \new_[12528]_  & \new_[12519]_ ;
  assign \new_[1925]_  = \new_[12512]_  & \new_[12503]_ ;
  assign \new_[1926]_  = \new_[12496]_  & \new_[12487]_ ;
  assign \new_[1927]_  = \new_[12480]_  & \new_[12471]_ ;
  assign \new_[1928]_  = \new_[12464]_  & \new_[12455]_ ;
  assign \new_[1929]_  = \new_[12448]_  & \new_[12439]_ ;
  assign \new_[1930]_  = \new_[12432]_  & \new_[12423]_ ;
  assign \new_[1931]_  = \new_[12416]_  & \new_[12407]_ ;
  assign \new_[1932]_  = \new_[12400]_  & \new_[12391]_ ;
  assign \new_[1933]_  = \new_[12384]_  & \new_[12375]_ ;
  assign \new_[1934]_  = \new_[12368]_  & \new_[12359]_ ;
  assign \new_[1935]_  = \new_[12352]_  & \new_[12343]_ ;
  assign \new_[1936]_  = \new_[12336]_  & \new_[12327]_ ;
  assign \new_[1937]_  = \new_[12320]_  & \new_[12311]_ ;
  assign \new_[1938]_  = \new_[12304]_  & \new_[12295]_ ;
  assign \new_[1939]_  = \new_[12288]_  & \new_[12279]_ ;
  assign \new_[1940]_  = \new_[12272]_  & \new_[12263]_ ;
  assign \new_[1941]_  = \new_[12256]_  & \new_[12247]_ ;
  assign \new_[1942]_  = \new_[12240]_  & \new_[12231]_ ;
  assign \new_[1943]_  = \new_[12224]_  & \new_[12215]_ ;
  assign \new_[1944]_  = \new_[12208]_  & \new_[12199]_ ;
  assign \new_[1945]_  = \new_[12192]_  & \new_[12183]_ ;
  assign \new_[1946]_  = \new_[12176]_  & \new_[12167]_ ;
  assign \new_[1947]_  = \new_[12160]_  & \new_[12151]_ ;
  assign \new_[1948]_  = \new_[12144]_  & \new_[12135]_ ;
  assign \new_[1949]_  = \new_[12128]_  & \new_[12119]_ ;
  assign \new_[1950]_  = \new_[12112]_  & \new_[12103]_ ;
  assign \new_[1951]_  = \new_[12096]_  & \new_[12087]_ ;
  assign \new_[1952]_  = \new_[12080]_  & \new_[12071]_ ;
  assign \new_[1953]_  = \new_[12064]_  & \new_[12055]_ ;
  assign \new_[1954]_  = \new_[12048]_  & \new_[12039]_ ;
  assign \new_[1955]_  = \new_[12032]_  & \new_[12023]_ ;
  assign \new_[1956]_  = \new_[12016]_  & \new_[12007]_ ;
  assign \new_[1957]_  = \new_[12000]_  & \new_[11991]_ ;
  assign \new_[1958]_  = \new_[11984]_  & \new_[11975]_ ;
  assign \new_[1959]_  = \new_[11968]_  & \new_[11959]_ ;
  assign \new_[1960]_  = \new_[11952]_  & \new_[11943]_ ;
  assign \new_[1961]_  = \new_[11936]_  & \new_[11927]_ ;
  assign \new_[1962]_  = \new_[11920]_  & \new_[11911]_ ;
  assign \new_[1963]_  = \new_[11904]_  & \new_[11895]_ ;
  assign \new_[1964]_  = \new_[11888]_  & \new_[11879]_ ;
  assign \new_[1965]_  = \new_[11872]_  & \new_[11863]_ ;
  assign \new_[1966]_  = \new_[11856]_  & \new_[11847]_ ;
  assign \new_[1967]_  = \new_[11840]_  & \new_[11831]_ ;
  assign \new_[1968]_  = \new_[11824]_  & \new_[11815]_ ;
  assign \new_[1969]_  = \new_[11808]_  & \new_[11799]_ ;
  assign \new_[1970]_  = \new_[11792]_  & \new_[11783]_ ;
  assign \new_[1971]_  = \new_[11776]_  & \new_[11767]_ ;
  assign \new_[1972]_  = \new_[11760]_  & \new_[11751]_ ;
  assign \new_[1973]_  = \new_[11744]_  & \new_[11735]_ ;
  assign \new_[1974]_  = \new_[11728]_  & \new_[11719]_ ;
  assign \new_[1975]_  = \new_[11712]_  & \new_[11703]_ ;
  assign \new_[1976]_  = \new_[11696]_  & \new_[11687]_ ;
  assign \new_[1977]_  = \new_[11680]_  & \new_[11671]_ ;
  assign \new_[1978]_  = \new_[11664]_  & \new_[11655]_ ;
  assign \new_[1979]_  = \new_[11648]_  & \new_[11639]_ ;
  assign \new_[1980]_  = \new_[11632]_  & \new_[11623]_ ;
  assign \new_[1981]_  = \new_[11616]_  & \new_[11607]_ ;
  assign \new_[1982]_  = \new_[11600]_  & \new_[11591]_ ;
  assign \new_[1983]_  = \new_[11584]_  & \new_[11575]_ ;
  assign \new_[1984]_  = \new_[11568]_  & \new_[11559]_ ;
  assign \new_[1985]_  = \new_[11552]_  & \new_[11543]_ ;
  assign \new_[1986]_  = \new_[11536]_  & \new_[11527]_ ;
  assign \new_[1987]_  = \new_[11520]_  & \new_[11511]_ ;
  assign \new_[1988]_  = \new_[11504]_  & \new_[11495]_ ;
  assign \new_[1989]_  = \new_[11488]_  & \new_[11479]_ ;
  assign \new_[1990]_  = \new_[11472]_  & \new_[11463]_ ;
  assign \new_[1991]_  = \new_[11456]_  & \new_[11447]_ ;
  assign \new_[1992]_  = \new_[11440]_  & \new_[11431]_ ;
  assign \new_[1993]_  = \new_[11424]_  & \new_[11415]_ ;
  assign \new_[1994]_  = \new_[11408]_  & \new_[11399]_ ;
  assign \new_[1995]_  = \new_[11392]_  & \new_[11383]_ ;
  assign \new_[1996]_  = \new_[11376]_  & \new_[11367]_ ;
  assign \new_[1997]_  = \new_[11360]_  & \new_[11351]_ ;
  assign \new_[1998]_  = \new_[11344]_  & \new_[11335]_ ;
  assign \new_[1999]_  = \new_[11328]_  & \new_[11319]_ ;
  assign \new_[2000]_  = \new_[11312]_  & \new_[11303]_ ;
  assign \new_[2001]_  = \new_[11296]_  & \new_[11287]_ ;
  assign \new_[2002]_  = \new_[11280]_  & \new_[11271]_ ;
  assign \new_[2003]_  = \new_[11264]_  & \new_[11255]_ ;
  assign \new_[2004]_  = \new_[11248]_  & \new_[11239]_ ;
  assign \new_[2005]_  = \new_[11232]_  & \new_[11223]_ ;
  assign \new_[2006]_  = \new_[11216]_  & \new_[11207]_ ;
  assign \new_[2007]_  = \new_[11200]_  & \new_[11191]_ ;
  assign \new_[2008]_  = \new_[11184]_  & \new_[11175]_ ;
  assign \new_[2009]_  = \new_[11168]_  & \new_[11159]_ ;
  assign \new_[2010]_  = \new_[11152]_  & \new_[11143]_ ;
  assign \new_[2011]_  = \new_[11136]_  & \new_[11127]_ ;
  assign \new_[2012]_  = \new_[11120]_  & \new_[11111]_ ;
  assign \new_[2013]_  = \new_[11104]_  & \new_[11095]_ ;
  assign \new_[2014]_  = \new_[11088]_  & \new_[11079]_ ;
  assign \new_[2015]_  = \new_[11072]_  & \new_[11063]_ ;
  assign \new_[2016]_  = \new_[11056]_  & \new_[11047]_ ;
  assign \new_[2017]_  = \new_[11040]_  & \new_[11031]_ ;
  assign \new_[2018]_  = \new_[11024]_  & \new_[11015]_ ;
  assign \new_[2019]_  = \new_[11008]_  & \new_[10999]_ ;
  assign \new_[2020]_  = \new_[10992]_  & \new_[10983]_ ;
  assign \new_[2021]_  = \new_[10976]_  & \new_[10967]_ ;
  assign \new_[2022]_  = \new_[10960]_  & \new_[10951]_ ;
  assign \new_[2023]_  = \new_[10944]_  & \new_[10935]_ ;
  assign \new_[2024]_  = \new_[10928]_  & \new_[10919]_ ;
  assign \new_[2025]_  = \new_[10912]_  & \new_[10903]_ ;
  assign \new_[2026]_  = \new_[10896]_  & \new_[10887]_ ;
  assign \new_[2027]_  = \new_[10880]_  & \new_[10871]_ ;
  assign \new_[2028]_  = \new_[10864]_  & \new_[10855]_ ;
  assign \new_[2029]_  = \new_[10848]_  & \new_[10839]_ ;
  assign \new_[2030]_  = \new_[10832]_  & \new_[10823]_ ;
  assign \new_[2031]_  = \new_[10816]_  & \new_[10807]_ ;
  assign \new_[2032]_  = \new_[10800]_  & \new_[10791]_ ;
  assign \new_[2033]_  = \new_[10784]_  & \new_[10775]_ ;
  assign \new_[2034]_  = \new_[10768]_  & \new_[10759]_ ;
  assign \new_[2035]_  = \new_[10752]_  & \new_[10743]_ ;
  assign \new_[2036]_  = \new_[10736]_  & \new_[10727]_ ;
  assign \new_[2037]_  = \new_[10720]_  & \new_[10711]_ ;
  assign \new_[2038]_  = \new_[10704]_  & \new_[10695]_ ;
  assign \new_[2039]_  = \new_[10688]_  & \new_[10679]_ ;
  assign \new_[2040]_  = \new_[10672]_  & \new_[10663]_ ;
  assign \new_[2041]_  = \new_[10656]_  & \new_[10647]_ ;
  assign \new_[2042]_  = \new_[10640]_  & \new_[10631]_ ;
  assign \new_[2043]_  = \new_[10624]_  & \new_[10615]_ ;
  assign \new_[2044]_  = \new_[10608]_  & \new_[10599]_ ;
  assign \new_[2045]_  = \new_[10592]_  & \new_[10583]_ ;
  assign \new_[2046]_  = \new_[10576]_  & \new_[10567]_ ;
  assign \new_[2047]_  = \new_[10560]_  & \new_[10551]_ ;
  assign \new_[2048]_  = \new_[10544]_  & \new_[10535]_ ;
  assign \new_[2049]_  = \new_[10528]_  & \new_[10519]_ ;
  assign \new_[2050]_  = \new_[10512]_  & \new_[10503]_ ;
  assign \new_[2051]_  = \new_[10496]_  & \new_[10487]_ ;
  assign \new_[2052]_  = \new_[10480]_  & \new_[10471]_ ;
  assign \new_[2053]_  = \new_[10464]_  & \new_[10455]_ ;
  assign \new_[2054]_  = \new_[10448]_  & \new_[10439]_ ;
  assign \new_[2055]_  = \new_[10432]_  & \new_[10423]_ ;
  assign \new_[2056]_  = \new_[10416]_  & \new_[10407]_ ;
  assign \new_[2057]_  = \new_[10400]_  & \new_[10391]_ ;
  assign \new_[2058]_  = \new_[10384]_  & \new_[10375]_ ;
  assign \new_[2059]_  = \new_[10368]_  & \new_[10359]_ ;
  assign \new_[2060]_  = \new_[10352]_  & \new_[10343]_ ;
  assign \new_[2061]_  = \new_[10336]_  & \new_[10327]_ ;
  assign \new_[2062]_  = \new_[10320]_  & \new_[10311]_ ;
  assign \new_[2063]_  = \new_[10304]_  & \new_[10295]_ ;
  assign \new_[2064]_  = \new_[10288]_  & \new_[10279]_ ;
  assign \new_[2065]_  = \new_[10272]_  & \new_[10263]_ ;
  assign \new_[2066]_  = \new_[10256]_  & \new_[10247]_ ;
  assign \new_[2067]_  = \new_[10240]_  & \new_[10231]_ ;
  assign \new_[2068]_  = \new_[10224]_  & \new_[10215]_ ;
  assign \new_[2069]_  = \new_[10208]_  & \new_[10199]_ ;
  assign \new_[2070]_  = \new_[10192]_  & \new_[10183]_ ;
  assign \new_[2071]_  = \new_[10176]_  & \new_[10167]_ ;
  assign \new_[2072]_  = \new_[10160]_  & \new_[10151]_ ;
  assign \new_[2073]_  = \new_[10144]_  & \new_[10135]_ ;
  assign \new_[2074]_  = \new_[10128]_  & \new_[10119]_ ;
  assign \new_[2075]_  = \new_[10112]_  & \new_[10103]_ ;
  assign \new_[2076]_  = \new_[10096]_  & \new_[10087]_ ;
  assign \new_[2077]_  = \new_[10080]_  & \new_[10071]_ ;
  assign \new_[2078]_  = \new_[10064]_  & \new_[10055]_ ;
  assign \new_[2079]_  = \new_[10048]_  & \new_[10039]_ ;
  assign \new_[2080]_  = \new_[10032]_  & \new_[10023]_ ;
  assign \new_[2081]_  = \new_[10016]_  & \new_[10007]_ ;
  assign \new_[2082]_  = \new_[10000]_  & \new_[9991]_ ;
  assign \new_[2083]_  = \new_[9984]_  & \new_[9977]_ ;
  assign \new_[2084]_  = \new_[9970]_  & \new_[9963]_ ;
  assign \new_[2085]_  = \new_[9956]_  & \new_[9949]_ ;
  assign \new_[2086]_  = \new_[9942]_  & \new_[9935]_ ;
  assign \new_[2087]_  = \new_[9928]_  & \new_[9921]_ ;
  assign \new_[2088]_  = \new_[9914]_  & \new_[9907]_ ;
  assign \new_[2089]_  = \new_[9900]_  & \new_[9893]_ ;
  assign \new_[2090]_  = \new_[9886]_  & \new_[9879]_ ;
  assign \new_[2091]_  = \new_[9872]_  & \new_[9865]_ ;
  assign \new_[2092]_  = \new_[9858]_  & \new_[9851]_ ;
  assign \new_[2093]_  = \new_[9844]_  & \new_[9837]_ ;
  assign \new_[2094]_  = \new_[9830]_  & \new_[9823]_ ;
  assign \new_[2095]_  = \new_[9816]_  & \new_[9809]_ ;
  assign \new_[2096]_  = \new_[9802]_  & \new_[9795]_ ;
  assign \new_[2097]_  = \new_[9788]_  & \new_[9781]_ ;
  assign \new_[2098]_  = \new_[9774]_  & \new_[9767]_ ;
  assign \new_[2099]_  = \new_[9760]_  & \new_[9753]_ ;
  assign \new_[2100]_  = \new_[9746]_  & \new_[9739]_ ;
  assign \new_[2101]_  = \new_[9732]_  & \new_[9725]_ ;
  assign \new_[2102]_  = \new_[9718]_  & \new_[9711]_ ;
  assign \new_[2103]_  = \new_[9704]_  & \new_[9697]_ ;
  assign \new_[2104]_  = \new_[9690]_  & \new_[9683]_ ;
  assign \new_[2105]_  = \new_[9676]_  & \new_[9669]_ ;
  assign \new_[2106]_  = \new_[9662]_  & \new_[9655]_ ;
  assign \new_[2107]_  = \new_[9648]_  & \new_[9641]_ ;
  assign \new_[2108]_  = \new_[9634]_  & \new_[9627]_ ;
  assign \new_[2109]_  = \new_[9620]_  & \new_[9613]_ ;
  assign \new_[2110]_  = \new_[9606]_  & \new_[9599]_ ;
  assign \new_[2111]_  = \new_[9592]_  & \new_[9585]_ ;
  assign \new_[2112]_  = \new_[9578]_  & \new_[9571]_ ;
  assign \new_[2113]_  = \new_[9564]_  & \new_[9557]_ ;
  assign \new_[2114]_  = \new_[9550]_  & \new_[9543]_ ;
  assign \new_[2115]_  = \new_[9536]_  & \new_[9529]_ ;
  assign \new_[2116]_  = \new_[9522]_  & \new_[9515]_ ;
  assign \new_[2117]_  = \new_[9508]_  & \new_[9501]_ ;
  assign \new_[2118]_  = \new_[9494]_  & \new_[9487]_ ;
  assign \new_[2119]_  = \new_[9480]_  & \new_[9473]_ ;
  assign \new_[2120]_  = \new_[9466]_  & \new_[9459]_ ;
  assign \new_[2121]_  = \new_[9452]_  & \new_[9445]_ ;
  assign \new_[2122]_  = \new_[9438]_  & \new_[9431]_ ;
  assign \new_[2123]_  = \new_[9424]_  & \new_[9417]_ ;
  assign \new_[2124]_  = \new_[9410]_  & \new_[9403]_ ;
  assign \new_[2125]_  = \new_[9396]_  & \new_[9389]_ ;
  assign \new_[2126]_  = \new_[9382]_  & \new_[9375]_ ;
  assign \new_[2127]_  = \new_[9368]_  & \new_[9361]_ ;
  assign \new_[2128]_  = \new_[9354]_  & \new_[9347]_ ;
  assign \new_[2129]_  = \new_[9340]_  & \new_[9333]_ ;
  assign \new_[2130]_  = \new_[9326]_  & \new_[9319]_ ;
  assign \new_[2131]_  = \new_[9312]_  & \new_[9305]_ ;
  assign \new_[2132]_  = \new_[9298]_  & \new_[9291]_ ;
  assign \new_[2133]_  = \new_[9284]_  & \new_[9277]_ ;
  assign \new_[2134]_  = \new_[9270]_  & \new_[9263]_ ;
  assign \new_[2135]_  = \new_[9256]_  & \new_[9249]_ ;
  assign \new_[2136]_  = \new_[9242]_  & \new_[9235]_ ;
  assign \new_[2137]_  = \new_[9228]_  & \new_[9221]_ ;
  assign \new_[2138]_  = \new_[9214]_  & \new_[9207]_ ;
  assign \new_[2139]_  = \new_[9200]_  & \new_[9193]_ ;
  assign \new_[2140]_  = \new_[9186]_  & \new_[9179]_ ;
  assign \new_[2141]_  = \new_[9172]_  & \new_[9165]_ ;
  assign \new_[2142]_  = \new_[9158]_  & \new_[9151]_ ;
  assign \new_[2143]_  = \new_[9144]_  & \new_[9137]_ ;
  assign \new_[2144]_  = \new_[9130]_  & \new_[9123]_ ;
  assign \new_[2145]_  = \new_[9116]_  & \new_[9109]_ ;
  assign \new_[2146]_  = \new_[9102]_  & \new_[9095]_ ;
  assign \new_[2147]_  = \new_[9088]_  & \new_[9081]_ ;
  assign \new_[2148]_  = \new_[9074]_  & \new_[9067]_ ;
  assign \new_[2149]_  = \new_[9060]_  & \new_[9053]_ ;
  assign \new_[2150]_  = \new_[9046]_  & \new_[9039]_ ;
  assign \new_[2151]_  = \new_[9032]_  & \new_[9025]_ ;
  assign \new_[2152]_  = \new_[9018]_  & \new_[9011]_ ;
  assign \new_[2153]_  = \new_[9004]_  & \new_[8997]_ ;
  assign \new_[2154]_  = \new_[8990]_  & \new_[8983]_ ;
  assign \new_[2155]_  = \new_[8976]_  & \new_[8969]_ ;
  assign \new_[2156]_  = \new_[8962]_  & \new_[8955]_ ;
  assign \new_[2157]_  = \new_[8948]_  & \new_[8941]_ ;
  assign \new_[2158]_  = \new_[8934]_  & \new_[8927]_ ;
  assign \new_[2159]_  = \new_[8920]_  & \new_[8913]_ ;
  assign \new_[2160]_  = \new_[8906]_  & \new_[8899]_ ;
  assign \new_[2161]_  = \new_[8892]_  & \new_[8885]_ ;
  assign \new_[2162]_  = \new_[8878]_  & \new_[8871]_ ;
  assign \new_[2163]_  = \new_[8864]_  & \new_[8857]_ ;
  assign \new_[2164]_  = \new_[8850]_  & \new_[8843]_ ;
  assign \new_[2165]_  = \new_[8836]_  & \new_[8829]_ ;
  assign \new_[2166]_  = \new_[8822]_  & \new_[8815]_ ;
  assign \new_[2167]_  = \new_[8808]_  & \new_[8801]_ ;
  assign \new_[2168]_  = \new_[8794]_  & \new_[8787]_ ;
  assign \new_[2169]_  = \new_[8780]_  & \new_[8773]_ ;
  assign \new_[2170]_  = \new_[8766]_  & \new_[8759]_ ;
  assign \new_[2171]_  = \new_[8752]_  & \new_[8745]_ ;
  assign \new_[2172]_  = \new_[8738]_  & \new_[8731]_ ;
  assign \new_[2173]_  = \new_[8724]_  & \new_[8717]_ ;
  assign \new_[2174]_  = \new_[8710]_  & \new_[8703]_ ;
  assign \new_[2175]_  = \new_[8696]_  & \new_[8689]_ ;
  assign \new_[2176]_  = \new_[8682]_  & \new_[8675]_ ;
  assign \new_[2177]_  = \new_[8668]_  & \new_[8661]_ ;
  assign \new_[2178]_  = \new_[8654]_  & \new_[8647]_ ;
  assign \new_[2179]_  = \new_[8640]_  & \new_[8633]_ ;
  assign \new_[2180]_  = \new_[8626]_  & \new_[8619]_ ;
  assign \new_[2181]_  = \new_[8612]_  & \new_[8605]_ ;
  assign \new_[2182]_  = \new_[8598]_  & \new_[8591]_ ;
  assign \new_[2183]_  = \new_[8584]_  & \new_[8577]_ ;
  assign \new_[2184]_  = \new_[8570]_  & \new_[8563]_ ;
  assign \new_[2185]_  = \new_[8556]_  & \new_[8549]_ ;
  assign \new_[2186]_  = \new_[8542]_  & \new_[8535]_ ;
  assign \new_[2187]_  = \new_[8528]_  & \new_[8521]_ ;
  assign \new_[2188]_  = \new_[8514]_  & \new_[8507]_ ;
  assign \new_[2189]_  = \new_[8500]_  & \new_[8493]_ ;
  assign \new_[2190]_  = \new_[8486]_  & \new_[8479]_ ;
  assign \new_[2191]_  = \new_[8472]_  & \new_[8465]_ ;
  assign \new_[2192]_  = \new_[8458]_  & \new_[8451]_ ;
  assign \new_[2193]_  = \new_[8444]_  & \new_[8437]_ ;
  assign \new_[2194]_  = \new_[8430]_  & \new_[8423]_ ;
  assign \new_[2195]_  = \new_[8416]_  & \new_[8409]_ ;
  assign \new_[2196]_  = \new_[8402]_  & \new_[8395]_ ;
  assign \new_[2197]_  = \new_[8388]_  & \new_[8381]_ ;
  assign \new_[2198]_  = \new_[8374]_  & \new_[8367]_ ;
  assign \new_[2199]_  = \new_[8360]_  & \new_[8353]_ ;
  assign \new_[2200]_  = \new_[8346]_  & \new_[8339]_ ;
  assign \new_[2201]_  = \new_[8332]_  & \new_[8325]_ ;
  assign \new_[2202]_  = \new_[8318]_  & \new_[8311]_ ;
  assign \new_[2203]_  = \new_[8304]_  & \new_[8297]_ ;
  assign \new_[2204]_  = \new_[8290]_  & \new_[8283]_ ;
  assign \new_[2205]_  = \new_[8276]_  & \new_[8269]_ ;
  assign \new_[2206]_  = \new_[8262]_  & \new_[8255]_ ;
  assign \new_[2207]_  = \new_[8248]_  & \new_[8241]_ ;
  assign \new_[2208]_  = \new_[8234]_  & \new_[8227]_ ;
  assign \new_[2209]_  = \new_[8220]_  & \new_[8213]_ ;
  assign \new_[2210]_  = \new_[8206]_  & \new_[8199]_ ;
  assign \new_[2211]_  = \new_[8192]_  & \new_[8185]_ ;
  assign \new_[2212]_  = \new_[8178]_  & \new_[8171]_ ;
  assign \new_[2213]_  = \new_[8164]_  & \new_[8157]_ ;
  assign \new_[2214]_  = \new_[8150]_  & \new_[8143]_ ;
  assign \new_[2215]_  = \new_[8136]_  & \new_[8129]_ ;
  assign \new_[2216]_  = \new_[8122]_  & \new_[8115]_ ;
  assign \new_[2217]_  = \new_[8108]_  & \new_[8101]_ ;
  assign \new_[2218]_  = \new_[8094]_  & \new_[8087]_ ;
  assign \new_[2219]_  = \new_[8080]_  & \new_[8073]_ ;
  assign \new_[2220]_  = \new_[8066]_  & \new_[8059]_ ;
  assign \new_[2221]_  = \new_[8052]_  & \new_[8045]_ ;
  assign \new_[2222]_  = \new_[8038]_  & \new_[8031]_ ;
  assign \new_[2223]_  = \new_[8024]_  & \new_[8017]_ ;
  assign \new_[2224]_  = \new_[8010]_  & \new_[8003]_ ;
  assign \new_[2225]_  = \new_[7996]_  & \new_[7989]_ ;
  assign \new_[2226]_  = \new_[7982]_  & \new_[7975]_ ;
  assign \new_[2227]_  = \new_[7968]_  & \new_[7961]_ ;
  assign \new_[2228]_  = \new_[7954]_  & \new_[7947]_ ;
  assign \new_[2229]_  = \new_[7940]_  & \new_[7933]_ ;
  assign \new_[2230]_  = \new_[7926]_  & \new_[7919]_ ;
  assign \new_[2231]_  = \new_[7912]_  & \new_[7905]_ ;
  assign \new_[2232]_  = \new_[7898]_  & \new_[7891]_ ;
  assign \new_[2233]_  = \new_[7884]_  & \new_[7877]_ ;
  assign \new_[2234]_  = \new_[7870]_  & \new_[7863]_ ;
  assign \new_[2235]_  = \new_[7856]_  & \new_[7849]_ ;
  assign \new_[2236]_  = \new_[7842]_  & \new_[7835]_ ;
  assign \new_[2237]_  = \new_[7828]_  & \new_[7821]_ ;
  assign \new_[2238]_  = \new_[7814]_  & \new_[7807]_ ;
  assign \new_[2239]_  = \new_[7800]_  & \new_[7793]_ ;
  assign \new_[2240]_  = \new_[7786]_  & \new_[7779]_ ;
  assign \new_[2241]_  = \new_[7772]_  & \new_[7765]_ ;
  assign \new_[2242]_  = \new_[7758]_  & \new_[7751]_ ;
  assign \new_[2243]_  = \new_[7744]_  & \new_[7737]_ ;
  assign \new_[2244]_  = \new_[7730]_  & \new_[7723]_ ;
  assign \new_[2245]_  = \new_[7716]_  & \new_[7709]_ ;
  assign \new_[2246]_  = \new_[7702]_  & \new_[7695]_ ;
  assign \new_[2247]_  = \new_[7688]_  & \new_[7681]_ ;
  assign \new_[2248]_  = \new_[7674]_  & \new_[7667]_ ;
  assign \new_[2249]_  = \new_[7660]_  & \new_[7653]_ ;
  assign \new_[2250]_  = \new_[7646]_  & \new_[7639]_ ;
  assign \new_[2251]_  = \new_[7632]_  & \new_[7625]_ ;
  assign \new_[2252]_  = \new_[7620]_  & \new_[7613]_ ;
  assign \new_[2253]_  = \new_[7608]_  & \new_[7601]_ ;
  assign \new_[2254]_  = \new_[7596]_  & \new_[7589]_ ;
  assign \new_[2255]_  = \new_[7584]_  & \new_[7577]_ ;
  assign \new_[2256]_  = \new_[7572]_  & \new_[7565]_ ;
  assign \new_[2257]_  = \new_[7560]_  & \new_[7553]_ ;
  assign \new_[2258]_  = \new_[7548]_  & \new_[7541]_ ;
  assign \new_[2259]_  = \new_[7536]_  & \new_[7529]_ ;
  assign \new_[2260]_  = \new_[7524]_  & \new_[7517]_ ;
  assign \new_[2261]_  = \new_[7512]_  & \new_[7505]_ ;
  assign \new_[2262]_  = \new_[7500]_  & \new_[7493]_ ;
  assign \new_[2263]_  = \new_[7488]_  & \new_[7481]_ ;
  assign \new_[2264]_  = \new_[7476]_  & \new_[7469]_ ;
  assign \new_[2265]_  = \new_[7464]_  & \new_[7457]_ ;
  assign \new_[2266]_  = \new_[7452]_  & \new_[7445]_ ;
  assign \new_[2267]_  = \new_[7440]_  & \new_[7433]_ ;
  assign \new_[2268]_  = \new_[7428]_  & \new_[7421]_ ;
  assign \new_[2269]_  = \new_[7416]_  & \new_[7409]_ ;
  assign \new_[2270]_  = \new_[7404]_  & \new_[7397]_ ;
  assign \new_[2271]_  = \new_[7392]_  & \new_[7385]_ ;
  assign \new_[2272]_  = \new_[7380]_  & \new_[7373]_ ;
  assign \new_[2273]_  = \new_[7368]_  & \new_[7361]_ ;
  assign \new_[2274]_  = \new_[7356]_  & \new_[7349]_ ;
  assign \new_[2275]_  = \new_[7344]_  & \new_[7337]_ ;
  assign \new_[2276]_  = \new_[7332]_  & \new_[7325]_ ;
  assign \new_[2277]_  = \new_[7320]_  & \new_[7313]_ ;
  assign \new_[2278]_  = \new_[7308]_  & \new_[7301]_ ;
  assign \new_[2279]_  = \new_[7296]_  & \new_[7289]_ ;
  assign \new_[2280]_  = \new_[7284]_  & \new_[7277]_ ;
  assign \new_[2281]_  = \new_[7272]_  & \new_[7265]_ ;
  assign \new_[2282]_  = \new_[7260]_  & \new_[7253]_ ;
  assign \new_[2283]_  = \new_[7248]_  & \new_[7241]_ ;
  assign \new_[2284]_  = \new_[7236]_  & \new_[7229]_ ;
  assign \new_[2285]_  = \new_[7224]_  & \new_[7217]_ ;
  assign \new_[2286]_  = \new_[7212]_  & \new_[7205]_ ;
  assign \new_[2287]_  = \new_[7200]_  & \new_[7193]_ ;
  assign \new_[2288]_  = \new_[7188]_  & \new_[7181]_ ;
  assign \new_[2289]_  = \new_[7176]_  & \new_[7169]_ ;
  assign \new_[2290]_  = \new_[7164]_  & \new_[7157]_ ;
  assign \new_[2291]_  = \new_[7152]_  & \new_[7145]_ ;
  assign \new_[2292]_  = \new_[7140]_  & \new_[7133]_ ;
  assign \new_[2293]_  = \new_[7128]_  & \new_[7121]_ ;
  assign \new_[2294]_  = \new_[7116]_  & \new_[7109]_ ;
  assign \new_[2295]_  = \new_[7104]_  & \new_[7097]_ ;
  assign \new_[2296]_  = \new_[7092]_  & \new_[7085]_ ;
  assign \new_[2297]_  = \new_[7080]_  & \new_[7073]_ ;
  assign \new_[2298]_  = \new_[7068]_  & \new_[7061]_ ;
  assign \new_[2299]_  = \new_[7056]_  & \new_[7049]_ ;
  assign \new_[2300]_  = \new_[7044]_  & \new_[7037]_ ;
  assign \new_[2301]_  = \new_[7032]_  & \new_[7025]_ ;
  assign \new_[2302]_  = \new_[7020]_  & \new_[7013]_ ;
  assign \new_[2303]_  = \new_[7008]_  & \new_[7003]_ ;
  assign \new_[2304]_  = \new_[6998]_  & \new_[6993]_ ;
  assign \new_[2305]_  = \new_[6988]_  & \new_[6983]_ ;
  assign \new_[2306]_  = \new_[6978]_  & \new_[6973]_ ;
  assign \new_[2307]_  = \new_[6968]_  & \new_[6963]_ ;
  assign \new_[2308]_  = \new_[6958]_  & \new_[6953]_ ;
  assign \new_[2309]_  = \new_[6948]_  & \new_[6943]_ ;
  assign \new_[2310]_  = \new_[6938]_  & \new_[6933]_ ;
  assign \new_[2313]_  = \new_[2309]_  | \new_[2310]_ ;
  assign \new_[2316]_  = \new_[2307]_  | \new_[2308]_ ;
  assign \new_[2317]_  = \new_[2316]_  | \new_[2313]_ ;
  assign \new_[2320]_  = \new_[2305]_  | \new_[2306]_ ;
  assign \new_[2324]_  = \new_[2302]_  | \new_[2303]_ ;
  assign \new_[2325]_  = \new_[2304]_  | \new_[2324]_ ;
  assign \new_[2326]_  = \new_[2325]_  | \new_[2320]_ ;
  assign \new_[2327]_  = \new_[2326]_  | \new_[2317]_ ;
  assign \new_[2330]_  = \new_[2300]_  | \new_[2301]_ ;
  assign \new_[2333]_  = \new_[2298]_  | \new_[2299]_ ;
  assign \new_[2334]_  = \new_[2333]_  | \new_[2330]_ ;
  assign \new_[2337]_  = \new_[2296]_  | \new_[2297]_ ;
  assign \new_[2341]_  = \new_[2293]_  | \new_[2294]_ ;
  assign \new_[2342]_  = \new_[2295]_  | \new_[2341]_ ;
  assign \new_[2343]_  = \new_[2342]_  | \new_[2337]_ ;
  assign \new_[2344]_  = \new_[2343]_  | \new_[2334]_ ;
  assign \new_[2345]_  = \new_[2344]_  | \new_[2327]_ ;
  assign \new_[2348]_  = \new_[2291]_  | \new_[2292]_ ;
  assign \new_[2351]_  = \new_[2289]_  | \new_[2290]_ ;
  assign \new_[2352]_  = \new_[2351]_  | \new_[2348]_ ;
  assign \new_[2355]_  = \new_[2287]_  | \new_[2288]_ ;
  assign \new_[2359]_  = \new_[2284]_  | \new_[2285]_ ;
  assign \new_[2360]_  = \new_[2286]_  | \new_[2359]_ ;
  assign \new_[2361]_  = \new_[2360]_  | \new_[2355]_ ;
  assign \new_[2362]_  = \new_[2361]_  | \new_[2352]_ ;
  assign \new_[2365]_  = \new_[2282]_  | \new_[2283]_ ;
  assign \new_[2368]_  = \new_[2280]_  | \new_[2281]_ ;
  assign \new_[2369]_  = \new_[2368]_  | \new_[2365]_ ;
  assign \new_[2372]_  = \new_[2278]_  | \new_[2279]_ ;
  assign \new_[2376]_  = \new_[2275]_  | \new_[2276]_ ;
  assign \new_[2377]_  = \new_[2277]_  | \new_[2376]_ ;
  assign \new_[2378]_  = \new_[2377]_  | \new_[2372]_ ;
  assign \new_[2379]_  = \new_[2378]_  | \new_[2369]_ ;
  assign \new_[2380]_  = \new_[2379]_  | \new_[2362]_ ;
  assign \new_[2381]_  = \new_[2380]_  | \new_[2345]_ ;
  assign \new_[2384]_  = \new_[2273]_  | \new_[2274]_ ;
  assign \new_[2387]_  = \new_[2271]_  | \new_[2272]_ ;
  assign \new_[2388]_  = \new_[2387]_  | \new_[2384]_ ;
  assign \new_[2391]_  = \new_[2269]_  | \new_[2270]_ ;
  assign \new_[2395]_  = \new_[2266]_  | \new_[2267]_ ;
  assign \new_[2396]_  = \new_[2268]_  | \new_[2395]_ ;
  assign \new_[2397]_  = \new_[2396]_  | \new_[2391]_ ;
  assign \new_[2398]_  = \new_[2397]_  | \new_[2388]_ ;
  assign \new_[2401]_  = \new_[2264]_  | \new_[2265]_ ;
  assign \new_[2404]_  = \new_[2262]_  | \new_[2263]_ ;
  assign \new_[2405]_  = \new_[2404]_  | \new_[2401]_ ;
  assign \new_[2408]_  = \new_[2260]_  | \new_[2261]_ ;
  assign \new_[2412]_  = \new_[2257]_  | \new_[2258]_ ;
  assign \new_[2413]_  = \new_[2259]_  | \new_[2412]_ ;
  assign \new_[2414]_  = \new_[2413]_  | \new_[2408]_ ;
  assign \new_[2415]_  = \new_[2414]_  | \new_[2405]_ ;
  assign \new_[2416]_  = \new_[2415]_  | \new_[2398]_ ;
  assign \new_[2419]_  = \new_[2255]_  | \new_[2256]_ ;
  assign \new_[2422]_  = \new_[2253]_  | \new_[2254]_ ;
  assign \new_[2423]_  = \new_[2422]_  | \new_[2419]_ ;
  assign \new_[2426]_  = \new_[2251]_  | \new_[2252]_ ;
  assign \new_[2430]_  = \new_[2248]_  | \new_[2249]_ ;
  assign \new_[2431]_  = \new_[2250]_  | \new_[2430]_ ;
  assign \new_[2432]_  = \new_[2431]_  | \new_[2426]_ ;
  assign \new_[2433]_  = \new_[2432]_  | \new_[2423]_ ;
  assign \new_[2436]_  = \new_[2246]_  | \new_[2247]_ ;
  assign \new_[2439]_  = \new_[2244]_  | \new_[2245]_ ;
  assign \new_[2440]_  = \new_[2439]_  | \new_[2436]_ ;
  assign \new_[2443]_  = \new_[2242]_  | \new_[2243]_ ;
  assign \new_[2447]_  = \new_[2239]_  | \new_[2240]_ ;
  assign \new_[2448]_  = \new_[2241]_  | \new_[2447]_ ;
  assign \new_[2449]_  = \new_[2448]_  | \new_[2443]_ ;
  assign \new_[2450]_  = \new_[2449]_  | \new_[2440]_ ;
  assign \new_[2451]_  = \new_[2450]_  | \new_[2433]_ ;
  assign \new_[2452]_  = \new_[2451]_  | \new_[2416]_ ;
  assign \new_[2453]_  = \new_[2452]_  | \new_[2381]_ ;
  assign \new_[2456]_  = \new_[2237]_  | \new_[2238]_ ;
  assign \new_[2459]_  = \new_[2235]_  | \new_[2236]_ ;
  assign \new_[2460]_  = \new_[2459]_  | \new_[2456]_ ;
  assign \new_[2463]_  = \new_[2233]_  | \new_[2234]_ ;
  assign \new_[2467]_  = \new_[2230]_  | \new_[2231]_ ;
  assign \new_[2468]_  = \new_[2232]_  | \new_[2467]_ ;
  assign \new_[2469]_  = \new_[2468]_  | \new_[2463]_ ;
  assign \new_[2470]_  = \new_[2469]_  | \new_[2460]_ ;
  assign \new_[2473]_  = \new_[2228]_  | \new_[2229]_ ;
  assign \new_[2476]_  = \new_[2226]_  | \new_[2227]_ ;
  assign \new_[2477]_  = \new_[2476]_  | \new_[2473]_ ;
  assign \new_[2480]_  = \new_[2224]_  | \new_[2225]_ ;
  assign \new_[2484]_  = \new_[2221]_  | \new_[2222]_ ;
  assign \new_[2485]_  = \new_[2223]_  | \new_[2484]_ ;
  assign \new_[2486]_  = \new_[2485]_  | \new_[2480]_ ;
  assign \new_[2487]_  = \new_[2486]_  | \new_[2477]_ ;
  assign \new_[2488]_  = \new_[2487]_  | \new_[2470]_ ;
  assign \new_[2491]_  = \new_[2219]_  | \new_[2220]_ ;
  assign \new_[2494]_  = \new_[2217]_  | \new_[2218]_ ;
  assign \new_[2495]_  = \new_[2494]_  | \new_[2491]_ ;
  assign \new_[2498]_  = \new_[2215]_  | \new_[2216]_ ;
  assign \new_[2502]_  = \new_[2212]_  | \new_[2213]_ ;
  assign \new_[2503]_  = \new_[2214]_  | \new_[2502]_ ;
  assign \new_[2504]_  = \new_[2503]_  | \new_[2498]_ ;
  assign \new_[2505]_  = \new_[2504]_  | \new_[2495]_ ;
  assign \new_[2508]_  = \new_[2210]_  | \new_[2211]_ ;
  assign \new_[2511]_  = \new_[2208]_  | \new_[2209]_ ;
  assign \new_[2512]_  = \new_[2511]_  | \new_[2508]_ ;
  assign \new_[2515]_  = \new_[2206]_  | \new_[2207]_ ;
  assign \new_[2519]_  = \new_[2203]_  | \new_[2204]_ ;
  assign \new_[2520]_  = \new_[2205]_  | \new_[2519]_ ;
  assign \new_[2521]_  = \new_[2520]_  | \new_[2515]_ ;
  assign \new_[2522]_  = \new_[2521]_  | \new_[2512]_ ;
  assign \new_[2523]_  = \new_[2522]_  | \new_[2505]_ ;
  assign \new_[2524]_  = \new_[2523]_  | \new_[2488]_ ;
  assign \new_[2527]_  = \new_[2201]_  | \new_[2202]_ ;
  assign \new_[2530]_  = \new_[2199]_  | \new_[2200]_ ;
  assign \new_[2531]_  = \new_[2530]_  | \new_[2527]_ ;
  assign \new_[2534]_  = \new_[2197]_  | \new_[2198]_ ;
  assign \new_[2538]_  = \new_[2194]_  | \new_[2195]_ ;
  assign \new_[2539]_  = \new_[2196]_  | \new_[2538]_ ;
  assign \new_[2540]_  = \new_[2539]_  | \new_[2534]_ ;
  assign \new_[2541]_  = \new_[2540]_  | \new_[2531]_ ;
  assign \new_[2544]_  = \new_[2192]_  | \new_[2193]_ ;
  assign \new_[2547]_  = \new_[2190]_  | \new_[2191]_ ;
  assign \new_[2548]_  = \new_[2547]_  | \new_[2544]_ ;
  assign \new_[2551]_  = \new_[2188]_  | \new_[2189]_ ;
  assign \new_[2555]_  = \new_[2185]_  | \new_[2186]_ ;
  assign \new_[2556]_  = \new_[2187]_  | \new_[2555]_ ;
  assign \new_[2557]_  = \new_[2556]_  | \new_[2551]_ ;
  assign \new_[2558]_  = \new_[2557]_  | \new_[2548]_ ;
  assign \new_[2559]_  = \new_[2558]_  | \new_[2541]_ ;
  assign \new_[2562]_  = \new_[2183]_  | \new_[2184]_ ;
  assign \new_[2565]_  = \new_[2181]_  | \new_[2182]_ ;
  assign \new_[2566]_  = \new_[2565]_  | \new_[2562]_ ;
  assign \new_[2569]_  = \new_[2179]_  | \new_[2180]_ ;
  assign \new_[2573]_  = \new_[2176]_  | \new_[2177]_ ;
  assign \new_[2574]_  = \new_[2178]_  | \new_[2573]_ ;
  assign \new_[2575]_  = \new_[2574]_  | \new_[2569]_ ;
  assign \new_[2576]_  = \new_[2575]_  | \new_[2566]_ ;
  assign \new_[2579]_  = \new_[2174]_  | \new_[2175]_ ;
  assign \new_[2582]_  = \new_[2172]_  | \new_[2173]_ ;
  assign \new_[2583]_  = \new_[2582]_  | \new_[2579]_ ;
  assign \new_[2586]_  = \new_[2170]_  | \new_[2171]_ ;
  assign \new_[2590]_  = \new_[2167]_  | \new_[2168]_ ;
  assign \new_[2591]_  = \new_[2169]_  | \new_[2590]_ ;
  assign \new_[2592]_  = \new_[2591]_  | \new_[2586]_ ;
  assign \new_[2593]_  = \new_[2592]_  | \new_[2583]_ ;
  assign \new_[2594]_  = \new_[2593]_  | \new_[2576]_ ;
  assign \new_[2595]_  = \new_[2594]_  | \new_[2559]_ ;
  assign \new_[2596]_  = \new_[2595]_  | \new_[2524]_ ;
  assign \new_[2597]_  = \new_[2596]_  | \new_[2453]_ ;
  assign \new_[2600]_  = \new_[2165]_  | \new_[2166]_ ;
  assign \new_[2603]_  = \new_[2163]_  | \new_[2164]_ ;
  assign \new_[2604]_  = \new_[2603]_  | \new_[2600]_ ;
  assign \new_[2607]_  = \new_[2161]_  | \new_[2162]_ ;
  assign \new_[2611]_  = \new_[2158]_  | \new_[2159]_ ;
  assign \new_[2612]_  = \new_[2160]_  | \new_[2611]_ ;
  assign \new_[2613]_  = \new_[2612]_  | \new_[2607]_ ;
  assign \new_[2614]_  = \new_[2613]_  | \new_[2604]_ ;
  assign \new_[2617]_  = \new_[2156]_  | \new_[2157]_ ;
  assign \new_[2620]_  = \new_[2154]_  | \new_[2155]_ ;
  assign \new_[2621]_  = \new_[2620]_  | \new_[2617]_ ;
  assign \new_[2624]_  = \new_[2152]_  | \new_[2153]_ ;
  assign \new_[2628]_  = \new_[2149]_  | \new_[2150]_ ;
  assign \new_[2629]_  = \new_[2151]_  | \new_[2628]_ ;
  assign \new_[2630]_  = \new_[2629]_  | \new_[2624]_ ;
  assign \new_[2631]_  = \new_[2630]_  | \new_[2621]_ ;
  assign \new_[2632]_  = \new_[2631]_  | \new_[2614]_ ;
  assign \new_[2635]_  = \new_[2147]_  | \new_[2148]_ ;
  assign \new_[2638]_  = \new_[2145]_  | \new_[2146]_ ;
  assign \new_[2639]_  = \new_[2638]_  | \new_[2635]_ ;
  assign \new_[2642]_  = \new_[2143]_  | \new_[2144]_ ;
  assign \new_[2646]_  = \new_[2140]_  | \new_[2141]_ ;
  assign \new_[2647]_  = \new_[2142]_  | \new_[2646]_ ;
  assign \new_[2648]_  = \new_[2647]_  | \new_[2642]_ ;
  assign \new_[2649]_  = \new_[2648]_  | \new_[2639]_ ;
  assign \new_[2652]_  = \new_[2138]_  | \new_[2139]_ ;
  assign \new_[2655]_  = \new_[2136]_  | \new_[2137]_ ;
  assign \new_[2656]_  = \new_[2655]_  | \new_[2652]_ ;
  assign \new_[2659]_  = \new_[2134]_  | \new_[2135]_ ;
  assign \new_[2663]_  = \new_[2131]_  | \new_[2132]_ ;
  assign \new_[2664]_  = \new_[2133]_  | \new_[2663]_ ;
  assign \new_[2665]_  = \new_[2664]_  | \new_[2659]_ ;
  assign \new_[2666]_  = \new_[2665]_  | \new_[2656]_ ;
  assign \new_[2667]_  = \new_[2666]_  | \new_[2649]_ ;
  assign \new_[2668]_  = \new_[2667]_  | \new_[2632]_ ;
  assign \new_[2671]_  = \new_[2129]_  | \new_[2130]_ ;
  assign \new_[2674]_  = \new_[2127]_  | \new_[2128]_ ;
  assign \new_[2675]_  = \new_[2674]_  | \new_[2671]_ ;
  assign \new_[2678]_  = \new_[2125]_  | \new_[2126]_ ;
  assign \new_[2682]_  = \new_[2122]_  | \new_[2123]_ ;
  assign \new_[2683]_  = \new_[2124]_  | \new_[2682]_ ;
  assign \new_[2684]_  = \new_[2683]_  | \new_[2678]_ ;
  assign \new_[2685]_  = \new_[2684]_  | \new_[2675]_ ;
  assign \new_[2688]_  = \new_[2120]_  | \new_[2121]_ ;
  assign \new_[2691]_  = \new_[2118]_  | \new_[2119]_ ;
  assign \new_[2692]_  = \new_[2691]_  | \new_[2688]_ ;
  assign \new_[2695]_  = \new_[2116]_  | \new_[2117]_ ;
  assign \new_[2699]_  = \new_[2113]_  | \new_[2114]_ ;
  assign \new_[2700]_  = \new_[2115]_  | \new_[2699]_ ;
  assign \new_[2701]_  = \new_[2700]_  | \new_[2695]_ ;
  assign \new_[2702]_  = \new_[2701]_  | \new_[2692]_ ;
  assign \new_[2703]_  = \new_[2702]_  | \new_[2685]_ ;
  assign \new_[2706]_  = \new_[2111]_  | \new_[2112]_ ;
  assign \new_[2709]_  = \new_[2109]_  | \new_[2110]_ ;
  assign \new_[2710]_  = \new_[2709]_  | \new_[2706]_ ;
  assign \new_[2713]_  = \new_[2107]_  | \new_[2108]_ ;
  assign \new_[2717]_  = \new_[2104]_  | \new_[2105]_ ;
  assign \new_[2718]_  = \new_[2106]_  | \new_[2717]_ ;
  assign \new_[2719]_  = \new_[2718]_  | \new_[2713]_ ;
  assign \new_[2720]_  = \new_[2719]_  | \new_[2710]_ ;
  assign \new_[2723]_  = \new_[2102]_  | \new_[2103]_ ;
  assign \new_[2726]_  = \new_[2100]_  | \new_[2101]_ ;
  assign \new_[2727]_  = \new_[2726]_  | \new_[2723]_ ;
  assign \new_[2730]_  = \new_[2098]_  | \new_[2099]_ ;
  assign \new_[2734]_  = \new_[2095]_  | \new_[2096]_ ;
  assign \new_[2735]_  = \new_[2097]_  | \new_[2734]_ ;
  assign \new_[2736]_  = \new_[2735]_  | \new_[2730]_ ;
  assign \new_[2737]_  = \new_[2736]_  | \new_[2727]_ ;
  assign \new_[2738]_  = \new_[2737]_  | \new_[2720]_ ;
  assign \new_[2739]_  = \new_[2738]_  | \new_[2703]_ ;
  assign \new_[2740]_  = \new_[2739]_  | \new_[2668]_ ;
  assign \new_[2743]_  = \new_[2093]_  | \new_[2094]_ ;
  assign \new_[2746]_  = \new_[2091]_  | \new_[2092]_ ;
  assign \new_[2747]_  = \new_[2746]_  | \new_[2743]_ ;
  assign \new_[2750]_  = \new_[2089]_  | \new_[2090]_ ;
  assign \new_[2754]_  = \new_[2086]_  | \new_[2087]_ ;
  assign \new_[2755]_  = \new_[2088]_  | \new_[2754]_ ;
  assign \new_[2756]_  = \new_[2755]_  | \new_[2750]_ ;
  assign \new_[2757]_  = \new_[2756]_  | \new_[2747]_ ;
  assign \new_[2760]_  = \new_[2084]_  | \new_[2085]_ ;
  assign \new_[2763]_  = \new_[2082]_  | \new_[2083]_ ;
  assign \new_[2764]_  = \new_[2763]_  | \new_[2760]_ ;
  assign \new_[2767]_  = \new_[2080]_  | \new_[2081]_ ;
  assign \new_[2771]_  = \new_[2077]_  | \new_[2078]_ ;
  assign \new_[2772]_  = \new_[2079]_  | \new_[2771]_ ;
  assign \new_[2773]_  = \new_[2772]_  | \new_[2767]_ ;
  assign \new_[2774]_  = \new_[2773]_  | \new_[2764]_ ;
  assign \new_[2775]_  = \new_[2774]_  | \new_[2757]_ ;
  assign \new_[2778]_  = \new_[2075]_  | \new_[2076]_ ;
  assign \new_[2781]_  = \new_[2073]_  | \new_[2074]_ ;
  assign \new_[2782]_  = \new_[2781]_  | \new_[2778]_ ;
  assign \new_[2785]_  = \new_[2071]_  | \new_[2072]_ ;
  assign \new_[2789]_  = \new_[2068]_  | \new_[2069]_ ;
  assign \new_[2790]_  = \new_[2070]_  | \new_[2789]_ ;
  assign \new_[2791]_  = \new_[2790]_  | \new_[2785]_ ;
  assign \new_[2792]_  = \new_[2791]_  | \new_[2782]_ ;
  assign \new_[2795]_  = \new_[2066]_  | \new_[2067]_ ;
  assign \new_[2798]_  = \new_[2064]_  | \new_[2065]_ ;
  assign \new_[2799]_  = \new_[2798]_  | \new_[2795]_ ;
  assign \new_[2802]_  = \new_[2062]_  | \new_[2063]_ ;
  assign \new_[2806]_  = \new_[2059]_  | \new_[2060]_ ;
  assign \new_[2807]_  = \new_[2061]_  | \new_[2806]_ ;
  assign \new_[2808]_  = \new_[2807]_  | \new_[2802]_ ;
  assign \new_[2809]_  = \new_[2808]_  | \new_[2799]_ ;
  assign \new_[2810]_  = \new_[2809]_  | \new_[2792]_ ;
  assign \new_[2811]_  = \new_[2810]_  | \new_[2775]_ ;
  assign \new_[2814]_  = \new_[2057]_  | \new_[2058]_ ;
  assign \new_[2817]_  = \new_[2055]_  | \new_[2056]_ ;
  assign \new_[2818]_  = \new_[2817]_  | \new_[2814]_ ;
  assign \new_[2821]_  = \new_[2053]_  | \new_[2054]_ ;
  assign \new_[2825]_  = \new_[2050]_  | \new_[2051]_ ;
  assign \new_[2826]_  = \new_[2052]_  | \new_[2825]_ ;
  assign \new_[2827]_  = \new_[2826]_  | \new_[2821]_ ;
  assign \new_[2828]_  = \new_[2827]_  | \new_[2818]_ ;
  assign \new_[2831]_  = \new_[2048]_  | \new_[2049]_ ;
  assign \new_[2834]_  = \new_[2046]_  | \new_[2047]_ ;
  assign \new_[2835]_  = \new_[2834]_  | \new_[2831]_ ;
  assign \new_[2838]_  = \new_[2044]_  | \new_[2045]_ ;
  assign \new_[2842]_  = \new_[2041]_  | \new_[2042]_ ;
  assign \new_[2843]_  = \new_[2043]_  | \new_[2842]_ ;
  assign \new_[2844]_  = \new_[2843]_  | \new_[2838]_ ;
  assign \new_[2845]_  = \new_[2844]_  | \new_[2835]_ ;
  assign \new_[2846]_  = \new_[2845]_  | \new_[2828]_ ;
  assign \new_[2849]_  = \new_[2039]_  | \new_[2040]_ ;
  assign \new_[2852]_  = \new_[2037]_  | \new_[2038]_ ;
  assign \new_[2853]_  = \new_[2852]_  | \new_[2849]_ ;
  assign \new_[2856]_  = \new_[2035]_  | \new_[2036]_ ;
  assign \new_[2860]_  = \new_[2032]_  | \new_[2033]_ ;
  assign \new_[2861]_  = \new_[2034]_  | \new_[2860]_ ;
  assign \new_[2862]_  = \new_[2861]_  | \new_[2856]_ ;
  assign \new_[2863]_  = \new_[2862]_  | \new_[2853]_ ;
  assign \new_[2866]_  = \new_[2030]_  | \new_[2031]_ ;
  assign \new_[2869]_  = \new_[2028]_  | \new_[2029]_ ;
  assign \new_[2870]_  = \new_[2869]_  | \new_[2866]_ ;
  assign \new_[2873]_  = \new_[2026]_  | \new_[2027]_ ;
  assign \new_[2877]_  = \new_[2023]_  | \new_[2024]_ ;
  assign \new_[2878]_  = \new_[2025]_  | \new_[2877]_ ;
  assign \new_[2879]_  = \new_[2878]_  | \new_[2873]_ ;
  assign \new_[2880]_  = \new_[2879]_  | \new_[2870]_ ;
  assign \new_[2881]_  = \new_[2880]_  | \new_[2863]_ ;
  assign \new_[2882]_  = \new_[2881]_  | \new_[2846]_ ;
  assign \new_[2883]_  = \new_[2882]_  | \new_[2811]_ ;
  assign \new_[2884]_  = \new_[2883]_  | \new_[2740]_ ;
  assign \new_[2885]_  = \new_[2884]_  | \new_[2597]_ ;
  assign \new_[2888]_  = \new_[2021]_  | \new_[2022]_ ;
  assign \new_[2891]_  = \new_[2019]_  | \new_[2020]_ ;
  assign \new_[2892]_  = \new_[2891]_  | \new_[2888]_ ;
  assign \new_[2895]_  = \new_[2017]_  | \new_[2018]_ ;
  assign \new_[2899]_  = \new_[2014]_  | \new_[2015]_ ;
  assign \new_[2900]_  = \new_[2016]_  | \new_[2899]_ ;
  assign \new_[2901]_  = \new_[2900]_  | \new_[2895]_ ;
  assign \new_[2902]_  = \new_[2901]_  | \new_[2892]_ ;
  assign \new_[2905]_  = \new_[2012]_  | \new_[2013]_ ;
  assign \new_[2908]_  = \new_[2010]_  | \new_[2011]_ ;
  assign \new_[2909]_  = \new_[2908]_  | \new_[2905]_ ;
  assign \new_[2912]_  = \new_[2008]_  | \new_[2009]_ ;
  assign \new_[2916]_  = \new_[2005]_  | \new_[2006]_ ;
  assign \new_[2917]_  = \new_[2007]_  | \new_[2916]_ ;
  assign \new_[2918]_  = \new_[2917]_  | \new_[2912]_ ;
  assign \new_[2919]_  = \new_[2918]_  | \new_[2909]_ ;
  assign \new_[2920]_  = \new_[2919]_  | \new_[2902]_ ;
  assign \new_[2923]_  = \new_[2003]_  | \new_[2004]_ ;
  assign \new_[2926]_  = \new_[2001]_  | \new_[2002]_ ;
  assign \new_[2927]_  = \new_[2926]_  | \new_[2923]_ ;
  assign \new_[2930]_  = \new_[1999]_  | \new_[2000]_ ;
  assign \new_[2934]_  = \new_[1996]_  | \new_[1997]_ ;
  assign \new_[2935]_  = \new_[1998]_  | \new_[2934]_ ;
  assign \new_[2936]_  = \new_[2935]_  | \new_[2930]_ ;
  assign \new_[2937]_  = \new_[2936]_  | \new_[2927]_ ;
  assign \new_[2940]_  = \new_[1994]_  | \new_[1995]_ ;
  assign \new_[2943]_  = \new_[1992]_  | \new_[1993]_ ;
  assign \new_[2944]_  = \new_[2943]_  | \new_[2940]_ ;
  assign \new_[2947]_  = \new_[1990]_  | \new_[1991]_ ;
  assign \new_[2951]_  = \new_[1987]_  | \new_[1988]_ ;
  assign \new_[2952]_  = \new_[1989]_  | \new_[2951]_ ;
  assign \new_[2953]_  = \new_[2952]_  | \new_[2947]_ ;
  assign \new_[2954]_  = \new_[2953]_  | \new_[2944]_ ;
  assign \new_[2955]_  = \new_[2954]_  | \new_[2937]_ ;
  assign \new_[2956]_  = \new_[2955]_  | \new_[2920]_ ;
  assign \new_[2959]_  = \new_[1985]_  | \new_[1986]_ ;
  assign \new_[2962]_  = \new_[1983]_  | \new_[1984]_ ;
  assign \new_[2963]_  = \new_[2962]_  | \new_[2959]_ ;
  assign \new_[2966]_  = \new_[1981]_  | \new_[1982]_ ;
  assign \new_[2970]_  = \new_[1978]_  | \new_[1979]_ ;
  assign \new_[2971]_  = \new_[1980]_  | \new_[2970]_ ;
  assign \new_[2972]_  = \new_[2971]_  | \new_[2966]_ ;
  assign \new_[2973]_  = \new_[2972]_  | \new_[2963]_ ;
  assign \new_[2976]_  = \new_[1976]_  | \new_[1977]_ ;
  assign \new_[2979]_  = \new_[1974]_  | \new_[1975]_ ;
  assign \new_[2980]_  = \new_[2979]_  | \new_[2976]_ ;
  assign \new_[2983]_  = \new_[1972]_  | \new_[1973]_ ;
  assign \new_[2987]_  = \new_[1969]_  | \new_[1970]_ ;
  assign \new_[2988]_  = \new_[1971]_  | \new_[2987]_ ;
  assign \new_[2989]_  = \new_[2988]_  | \new_[2983]_ ;
  assign \new_[2990]_  = \new_[2989]_  | \new_[2980]_ ;
  assign \new_[2991]_  = \new_[2990]_  | \new_[2973]_ ;
  assign \new_[2994]_  = \new_[1967]_  | \new_[1968]_ ;
  assign \new_[2997]_  = \new_[1965]_  | \new_[1966]_ ;
  assign \new_[2998]_  = \new_[2997]_  | \new_[2994]_ ;
  assign \new_[3001]_  = \new_[1963]_  | \new_[1964]_ ;
  assign \new_[3005]_  = \new_[1960]_  | \new_[1961]_ ;
  assign \new_[3006]_  = \new_[1962]_  | \new_[3005]_ ;
  assign \new_[3007]_  = \new_[3006]_  | \new_[3001]_ ;
  assign \new_[3008]_  = \new_[3007]_  | \new_[2998]_ ;
  assign \new_[3011]_  = \new_[1958]_  | \new_[1959]_ ;
  assign \new_[3014]_  = \new_[1956]_  | \new_[1957]_ ;
  assign \new_[3015]_  = \new_[3014]_  | \new_[3011]_ ;
  assign \new_[3018]_  = \new_[1954]_  | \new_[1955]_ ;
  assign \new_[3022]_  = \new_[1951]_  | \new_[1952]_ ;
  assign \new_[3023]_  = \new_[1953]_  | \new_[3022]_ ;
  assign \new_[3024]_  = \new_[3023]_  | \new_[3018]_ ;
  assign \new_[3025]_  = \new_[3024]_  | \new_[3015]_ ;
  assign \new_[3026]_  = \new_[3025]_  | \new_[3008]_ ;
  assign \new_[3027]_  = \new_[3026]_  | \new_[2991]_ ;
  assign \new_[3028]_  = \new_[3027]_  | \new_[2956]_ ;
  assign \new_[3031]_  = \new_[1949]_  | \new_[1950]_ ;
  assign \new_[3034]_  = \new_[1947]_  | \new_[1948]_ ;
  assign \new_[3035]_  = \new_[3034]_  | \new_[3031]_ ;
  assign \new_[3038]_  = \new_[1945]_  | \new_[1946]_ ;
  assign \new_[3042]_  = \new_[1942]_  | \new_[1943]_ ;
  assign \new_[3043]_  = \new_[1944]_  | \new_[3042]_ ;
  assign \new_[3044]_  = \new_[3043]_  | \new_[3038]_ ;
  assign \new_[3045]_  = \new_[3044]_  | \new_[3035]_ ;
  assign \new_[3048]_  = \new_[1940]_  | \new_[1941]_ ;
  assign \new_[3051]_  = \new_[1938]_  | \new_[1939]_ ;
  assign \new_[3052]_  = \new_[3051]_  | \new_[3048]_ ;
  assign \new_[3055]_  = \new_[1936]_  | \new_[1937]_ ;
  assign \new_[3059]_  = \new_[1933]_  | \new_[1934]_ ;
  assign \new_[3060]_  = \new_[1935]_  | \new_[3059]_ ;
  assign \new_[3061]_  = \new_[3060]_  | \new_[3055]_ ;
  assign \new_[3062]_  = \new_[3061]_  | \new_[3052]_ ;
  assign \new_[3063]_  = \new_[3062]_  | \new_[3045]_ ;
  assign \new_[3066]_  = \new_[1931]_  | \new_[1932]_ ;
  assign \new_[3069]_  = \new_[1929]_  | \new_[1930]_ ;
  assign \new_[3070]_  = \new_[3069]_  | \new_[3066]_ ;
  assign \new_[3073]_  = \new_[1927]_  | \new_[1928]_ ;
  assign \new_[3077]_  = \new_[1924]_  | \new_[1925]_ ;
  assign \new_[3078]_  = \new_[1926]_  | \new_[3077]_ ;
  assign \new_[3079]_  = \new_[3078]_  | \new_[3073]_ ;
  assign \new_[3080]_  = \new_[3079]_  | \new_[3070]_ ;
  assign \new_[3083]_  = \new_[1922]_  | \new_[1923]_ ;
  assign \new_[3086]_  = \new_[1920]_  | \new_[1921]_ ;
  assign \new_[3087]_  = \new_[3086]_  | \new_[3083]_ ;
  assign \new_[3090]_  = \new_[1918]_  | \new_[1919]_ ;
  assign \new_[3094]_  = \new_[1915]_  | \new_[1916]_ ;
  assign \new_[3095]_  = \new_[1917]_  | \new_[3094]_ ;
  assign \new_[3096]_  = \new_[3095]_  | \new_[3090]_ ;
  assign \new_[3097]_  = \new_[3096]_  | \new_[3087]_ ;
  assign \new_[3098]_  = \new_[3097]_  | \new_[3080]_ ;
  assign \new_[3099]_  = \new_[3098]_  | \new_[3063]_ ;
  assign \new_[3102]_  = \new_[1913]_  | \new_[1914]_ ;
  assign \new_[3105]_  = \new_[1911]_  | \new_[1912]_ ;
  assign \new_[3106]_  = \new_[3105]_  | \new_[3102]_ ;
  assign \new_[3109]_  = \new_[1909]_  | \new_[1910]_ ;
  assign \new_[3113]_  = \new_[1906]_  | \new_[1907]_ ;
  assign \new_[3114]_  = \new_[1908]_  | \new_[3113]_ ;
  assign \new_[3115]_  = \new_[3114]_  | \new_[3109]_ ;
  assign \new_[3116]_  = \new_[3115]_  | \new_[3106]_ ;
  assign \new_[3119]_  = \new_[1904]_  | \new_[1905]_ ;
  assign \new_[3122]_  = \new_[1902]_  | \new_[1903]_ ;
  assign \new_[3123]_  = \new_[3122]_  | \new_[3119]_ ;
  assign \new_[3126]_  = \new_[1900]_  | \new_[1901]_ ;
  assign \new_[3130]_  = \new_[1897]_  | \new_[1898]_ ;
  assign \new_[3131]_  = \new_[1899]_  | \new_[3130]_ ;
  assign \new_[3132]_  = \new_[3131]_  | \new_[3126]_ ;
  assign \new_[3133]_  = \new_[3132]_  | \new_[3123]_ ;
  assign \new_[3134]_  = \new_[3133]_  | \new_[3116]_ ;
  assign \new_[3137]_  = \new_[1895]_  | \new_[1896]_ ;
  assign \new_[3140]_  = \new_[1893]_  | \new_[1894]_ ;
  assign \new_[3141]_  = \new_[3140]_  | \new_[3137]_ ;
  assign \new_[3144]_  = \new_[1891]_  | \new_[1892]_ ;
  assign \new_[3148]_  = \new_[1888]_  | \new_[1889]_ ;
  assign \new_[3149]_  = \new_[1890]_  | \new_[3148]_ ;
  assign \new_[3150]_  = \new_[3149]_  | \new_[3144]_ ;
  assign \new_[3151]_  = \new_[3150]_  | \new_[3141]_ ;
  assign \new_[3154]_  = \new_[1886]_  | \new_[1887]_ ;
  assign \new_[3157]_  = \new_[1884]_  | \new_[1885]_ ;
  assign \new_[3158]_  = \new_[3157]_  | \new_[3154]_ ;
  assign \new_[3161]_  = \new_[1882]_  | \new_[1883]_ ;
  assign \new_[3165]_  = \new_[1879]_  | \new_[1880]_ ;
  assign \new_[3166]_  = \new_[1881]_  | \new_[3165]_ ;
  assign \new_[3167]_  = \new_[3166]_  | \new_[3161]_ ;
  assign \new_[3168]_  = \new_[3167]_  | \new_[3158]_ ;
  assign \new_[3169]_  = \new_[3168]_  | \new_[3151]_ ;
  assign \new_[3170]_  = \new_[3169]_  | \new_[3134]_ ;
  assign \new_[3171]_  = \new_[3170]_  | \new_[3099]_ ;
  assign \new_[3172]_  = \new_[3171]_  | \new_[3028]_ ;
  assign \new_[3175]_  = \new_[1877]_  | \new_[1878]_ ;
  assign \new_[3178]_  = \new_[1875]_  | \new_[1876]_ ;
  assign \new_[3179]_  = \new_[3178]_  | \new_[3175]_ ;
  assign \new_[3182]_  = \new_[1873]_  | \new_[1874]_ ;
  assign \new_[3186]_  = \new_[1870]_  | \new_[1871]_ ;
  assign \new_[3187]_  = \new_[1872]_  | \new_[3186]_ ;
  assign \new_[3188]_  = \new_[3187]_  | \new_[3182]_ ;
  assign \new_[3189]_  = \new_[3188]_  | \new_[3179]_ ;
  assign \new_[3192]_  = \new_[1868]_  | \new_[1869]_ ;
  assign \new_[3195]_  = \new_[1866]_  | \new_[1867]_ ;
  assign \new_[3196]_  = \new_[3195]_  | \new_[3192]_ ;
  assign \new_[3199]_  = \new_[1864]_  | \new_[1865]_ ;
  assign \new_[3203]_  = \new_[1861]_  | \new_[1862]_ ;
  assign \new_[3204]_  = \new_[1863]_  | \new_[3203]_ ;
  assign \new_[3205]_  = \new_[3204]_  | \new_[3199]_ ;
  assign \new_[3206]_  = \new_[3205]_  | \new_[3196]_ ;
  assign \new_[3207]_  = \new_[3206]_  | \new_[3189]_ ;
  assign \new_[3210]_  = \new_[1859]_  | \new_[1860]_ ;
  assign \new_[3213]_  = \new_[1857]_  | \new_[1858]_ ;
  assign \new_[3214]_  = \new_[3213]_  | \new_[3210]_ ;
  assign \new_[3217]_  = \new_[1855]_  | \new_[1856]_ ;
  assign \new_[3221]_  = \new_[1852]_  | \new_[1853]_ ;
  assign \new_[3222]_  = \new_[1854]_  | \new_[3221]_ ;
  assign \new_[3223]_  = \new_[3222]_  | \new_[3217]_ ;
  assign \new_[3224]_  = \new_[3223]_  | \new_[3214]_ ;
  assign \new_[3227]_  = \new_[1850]_  | \new_[1851]_ ;
  assign \new_[3230]_  = \new_[1848]_  | \new_[1849]_ ;
  assign \new_[3231]_  = \new_[3230]_  | \new_[3227]_ ;
  assign \new_[3234]_  = \new_[1846]_  | \new_[1847]_ ;
  assign \new_[3238]_  = \new_[1843]_  | \new_[1844]_ ;
  assign \new_[3239]_  = \new_[1845]_  | \new_[3238]_ ;
  assign \new_[3240]_  = \new_[3239]_  | \new_[3234]_ ;
  assign \new_[3241]_  = \new_[3240]_  | \new_[3231]_ ;
  assign \new_[3242]_  = \new_[3241]_  | \new_[3224]_ ;
  assign \new_[3243]_  = \new_[3242]_  | \new_[3207]_ ;
  assign \new_[3246]_  = \new_[1841]_  | \new_[1842]_ ;
  assign \new_[3249]_  = \new_[1839]_  | \new_[1840]_ ;
  assign \new_[3250]_  = \new_[3249]_  | \new_[3246]_ ;
  assign \new_[3253]_  = \new_[1837]_  | \new_[1838]_ ;
  assign \new_[3257]_  = \new_[1834]_  | \new_[1835]_ ;
  assign \new_[3258]_  = \new_[1836]_  | \new_[3257]_ ;
  assign \new_[3259]_  = \new_[3258]_  | \new_[3253]_ ;
  assign \new_[3260]_  = \new_[3259]_  | \new_[3250]_ ;
  assign \new_[3263]_  = \new_[1832]_  | \new_[1833]_ ;
  assign \new_[3266]_  = \new_[1830]_  | \new_[1831]_ ;
  assign \new_[3267]_  = \new_[3266]_  | \new_[3263]_ ;
  assign \new_[3270]_  = \new_[1828]_  | \new_[1829]_ ;
  assign \new_[3274]_  = \new_[1825]_  | \new_[1826]_ ;
  assign \new_[3275]_  = \new_[1827]_  | \new_[3274]_ ;
  assign \new_[3276]_  = \new_[3275]_  | \new_[3270]_ ;
  assign \new_[3277]_  = \new_[3276]_  | \new_[3267]_ ;
  assign \new_[3278]_  = \new_[3277]_  | \new_[3260]_ ;
  assign \new_[3281]_  = \new_[1823]_  | \new_[1824]_ ;
  assign \new_[3284]_  = \new_[1821]_  | \new_[1822]_ ;
  assign \new_[3285]_  = \new_[3284]_  | \new_[3281]_ ;
  assign \new_[3288]_  = \new_[1819]_  | \new_[1820]_ ;
  assign \new_[3292]_  = \new_[1816]_  | \new_[1817]_ ;
  assign \new_[3293]_  = \new_[1818]_  | \new_[3292]_ ;
  assign \new_[3294]_  = \new_[3293]_  | \new_[3288]_ ;
  assign \new_[3295]_  = \new_[3294]_  | \new_[3285]_ ;
  assign \new_[3298]_  = \new_[1814]_  | \new_[1815]_ ;
  assign \new_[3301]_  = \new_[1812]_  | \new_[1813]_ ;
  assign \new_[3302]_  = \new_[3301]_  | \new_[3298]_ ;
  assign \new_[3305]_  = \new_[1810]_  | \new_[1811]_ ;
  assign \new_[3309]_  = \new_[1807]_  | \new_[1808]_ ;
  assign \new_[3310]_  = \new_[1809]_  | \new_[3309]_ ;
  assign \new_[3311]_  = \new_[3310]_  | \new_[3305]_ ;
  assign \new_[3312]_  = \new_[3311]_  | \new_[3302]_ ;
  assign \new_[3313]_  = \new_[3312]_  | \new_[3295]_ ;
  assign \new_[3314]_  = \new_[3313]_  | \new_[3278]_ ;
  assign \new_[3315]_  = \new_[3314]_  | \new_[3243]_ ;
  assign \new_[3318]_  = \new_[1805]_  | \new_[1806]_ ;
  assign \new_[3321]_  = \new_[1803]_  | \new_[1804]_ ;
  assign \new_[3322]_  = \new_[3321]_  | \new_[3318]_ ;
  assign \new_[3325]_  = \new_[1801]_  | \new_[1802]_ ;
  assign \new_[3329]_  = \new_[1798]_  | \new_[1799]_ ;
  assign \new_[3330]_  = \new_[1800]_  | \new_[3329]_ ;
  assign \new_[3331]_  = \new_[3330]_  | \new_[3325]_ ;
  assign \new_[3332]_  = \new_[3331]_  | \new_[3322]_ ;
  assign \new_[3335]_  = \new_[1796]_  | \new_[1797]_ ;
  assign \new_[3338]_  = \new_[1794]_  | \new_[1795]_ ;
  assign \new_[3339]_  = \new_[3338]_  | \new_[3335]_ ;
  assign \new_[3342]_  = \new_[1792]_  | \new_[1793]_ ;
  assign \new_[3346]_  = \new_[1789]_  | \new_[1790]_ ;
  assign \new_[3347]_  = \new_[1791]_  | \new_[3346]_ ;
  assign \new_[3348]_  = \new_[3347]_  | \new_[3342]_ ;
  assign \new_[3349]_  = \new_[3348]_  | \new_[3339]_ ;
  assign \new_[3350]_  = \new_[3349]_  | \new_[3332]_ ;
  assign \new_[3353]_  = \new_[1787]_  | \new_[1788]_ ;
  assign \new_[3356]_  = \new_[1785]_  | \new_[1786]_ ;
  assign \new_[3357]_  = \new_[3356]_  | \new_[3353]_ ;
  assign \new_[3360]_  = \new_[1783]_  | \new_[1784]_ ;
  assign \new_[3364]_  = \new_[1780]_  | \new_[1781]_ ;
  assign \new_[3365]_  = \new_[1782]_  | \new_[3364]_ ;
  assign \new_[3366]_  = \new_[3365]_  | \new_[3360]_ ;
  assign \new_[3367]_  = \new_[3366]_  | \new_[3357]_ ;
  assign \new_[3370]_  = \new_[1778]_  | \new_[1779]_ ;
  assign \new_[3373]_  = \new_[1776]_  | \new_[1777]_ ;
  assign \new_[3374]_  = \new_[3373]_  | \new_[3370]_ ;
  assign \new_[3377]_  = \new_[1774]_  | \new_[1775]_ ;
  assign \new_[3381]_  = \new_[1771]_  | \new_[1772]_ ;
  assign \new_[3382]_  = \new_[1773]_  | \new_[3381]_ ;
  assign \new_[3383]_  = \new_[3382]_  | \new_[3377]_ ;
  assign \new_[3384]_  = \new_[3383]_  | \new_[3374]_ ;
  assign \new_[3385]_  = \new_[3384]_  | \new_[3367]_ ;
  assign \new_[3386]_  = \new_[3385]_  | \new_[3350]_ ;
  assign \new_[3389]_  = \new_[1769]_  | \new_[1770]_ ;
  assign \new_[3392]_  = \new_[1767]_  | \new_[1768]_ ;
  assign \new_[3393]_  = \new_[3392]_  | \new_[3389]_ ;
  assign \new_[3396]_  = \new_[1765]_  | \new_[1766]_ ;
  assign \new_[3400]_  = \new_[1762]_  | \new_[1763]_ ;
  assign \new_[3401]_  = \new_[1764]_  | \new_[3400]_ ;
  assign \new_[3402]_  = \new_[3401]_  | \new_[3396]_ ;
  assign \new_[3403]_  = \new_[3402]_  | \new_[3393]_ ;
  assign \new_[3406]_  = \new_[1760]_  | \new_[1761]_ ;
  assign \new_[3409]_  = \new_[1758]_  | \new_[1759]_ ;
  assign \new_[3410]_  = \new_[3409]_  | \new_[3406]_ ;
  assign \new_[3413]_  = \new_[1756]_  | \new_[1757]_ ;
  assign \new_[3417]_  = \new_[1753]_  | \new_[1754]_ ;
  assign \new_[3418]_  = \new_[1755]_  | \new_[3417]_ ;
  assign \new_[3419]_  = \new_[3418]_  | \new_[3413]_ ;
  assign \new_[3420]_  = \new_[3419]_  | \new_[3410]_ ;
  assign \new_[3421]_  = \new_[3420]_  | \new_[3403]_ ;
  assign \new_[3424]_  = \new_[1751]_  | \new_[1752]_ ;
  assign \new_[3427]_  = \new_[1749]_  | \new_[1750]_ ;
  assign \new_[3428]_  = \new_[3427]_  | \new_[3424]_ ;
  assign \new_[3431]_  = \new_[1747]_  | \new_[1748]_ ;
  assign \new_[3435]_  = \new_[1744]_  | \new_[1745]_ ;
  assign \new_[3436]_  = \new_[1746]_  | \new_[3435]_ ;
  assign \new_[3437]_  = \new_[3436]_  | \new_[3431]_ ;
  assign \new_[3438]_  = \new_[3437]_  | \new_[3428]_ ;
  assign \new_[3441]_  = \new_[1742]_  | \new_[1743]_ ;
  assign \new_[3445]_  = \new_[1739]_  | \new_[1740]_ ;
  assign \new_[3446]_  = \new_[1741]_  | \new_[3445]_ ;
  assign \new_[3447]_  = \new_[3446]_  | \new_[3441]_ ;
  assign \new_[3450]_  = \new_[1737]_  | \new_[1738]_ ;
  assign \new_[3454]_  = \new_[1734]_  | \new_[1735]_ ;
  assign \new_[3455]_  = \new_[1736]_  | \new_[3454]_ ;
  assign \new_[3456]_  = \new_[3455]_  | \new_[3450]_ ;
  assign \new_[3457]_  = \new_[3456]_  | \new_[3447]_ ;
  assign \new_[3458]_  = \new_[3457]_  | \new_[3438]_ ;
  assign \new_[3459]_  = \new_[3458]_  | \new_[3421]_ ;
  assign \new_[3460]_  = \new_[3459]_  | \new_[3386]_ ;
  assign \new_[3461]_  = \new_[3460]_  | \new_[3315]_ ;
  assign \new_[3462]_  = \new_[3461]_  | \new_[3172]_ ;
  assign \new_[3463]_  = \new_[3462]_  | \new_[2885]_ ;
  assign \new_[3466]_  = \new_[1732]_  | \new_[1733]_ ;
  assign \new_[3469]_  = \new_[1730]_  | \new_[1731]_ ;
  assign \new_[3470]_  = \new_[3469]_  | \new_[3466]_ ;
  assign \new_[3473]_  = \new_[1728]_  | \new_[1729]_ ;
  assign \new_[3477]_  = \new_[1725]_  | \new_[1726]_ ;
  assign \new_[3478]_  = \new_[1727]_  | \new_[3477]_ ;
  assign \new_[3479]_  = \new_[3478]_  | \new_[3473]_ ;
  assign \new_[3480]_  = \new_[3479]_  | \new_[3470]_ ;
  assign \new_[3483]_  = \new_[1723]_  | \new_[1724]_ ;
  assign \new_[3486]_  = \new_[1721]_  | \new_[1722]_ ;
  assign \new_[3487]_  = \new_[3486]_  | \new_[3483]_ ;
  assign \new_[3490]_  = \new_[1719]_  | \new_[1720]_ ;
  assign \new_[3494]_  = \new_[1716]_  | \new_[1717]_ ;
  assign \new_[3495]_  = \new_[1718]_  | \new_[3494]_ ;
  assign \new_[3496]_  = \new_[3495]_  | \new_[3490]_ ;
  assign \new_[3497]_  = \new_[3496]_  | \new_[3487]_ ;
  assign \new_[3498]_  = \new_[3497]_  | \new_[3480]_ ;
  assign \new_[3501]_  = \new_[1714]_  | \new_[1715]_ ;
  assign \new_[3504]_  = \new_[1712]_  | \new_[1713]_ ;
  assign \new_[3505]_  = \new_[3504]_  | \new_[3501]_ ;
  assign \new_[3508]_  = \new_[1710]_  | \new_[1711]_ ;
  assign \new_[3512]_  = \new_[1707]_  | \new_[1708]_ ;
  assign \new_[3513]_  = \new_[1709]_  | \new_[3512]_ ;
  assign \new_[3514]_  = \new_[3513]_  | \new_[3508]_ ;
  assign \new_[3515]_  = \new_[3514]_  | \new_[3505]_ ;
  assign \new_[3518]_  = \new_[1705]_  | \new_[1706]_ ;
  assign \new_[3521]_  = \new_[1703]_  | \new_[1704]_ ;
  assign \new_[3522]_  = \new_[3521]_  | \new_[3518]_ ;
  assign \new_[3525]_  = \new_[1701]_  | \new_[1702]_ ;
  assign \new_[3529]_  = \new_[1698]_  | \new_[1699]_ ;
  assign \new_[3530]_  = \new_[1700]_  | \new_[3529]_ ;
  assign \new_[3531]_  = \new_[3530]_  | \new_[3525]_ ;
  assign \new_[3532]_  = \new_[3531]_  | \new_[3522]_ ;
  assign \new_[3533]_  = \new_[3532]_  | \new_[3515]_ ;
  assign \new_[3534]_  = \new_[3533]_  | \new_[3498]_ ;
  assign \new_[3537]_  = \new_[1696]_  | \new_[1697]_ ;
  assign \new_[3540]_  = \new_[1694]_  | \new_[1695]_ ;
  assign \new_[3541]_  = \new_[3540]_  | \new_[3537]_ ;
  assign \new_[3544]_  = \new_[1692]_  | \new_[1693]_ ;
  assign \new_[3548]_  = \new_[1689]_  | \new_[1690]_ ;
  assign \new_[3549]_  = \new_[1691]_  | \new_[3548]_ ;
  assign \new_[3550]_  = \new_[3549]_  | \new_[3544]_ ;
  assign \new_[3551]_  = \new_[3550]_  | \new_[3541]_ ;
  assign \new_[3554]_  = \new_[1687]_  | \new_[1688]_ ;
  assign \new_[3557]_  = \new_[1685]_  | \new_[1686]_ ;
  assign \new_[3558]_  = \new_[3557]_  | \new_[3554]_ ;
  assign \new_[3561]_  = \new_[1683]_  | \new_[1684]_ ;
  assign \new_[3565]_  = \new_[1680]_  | \new_[1681]_ ;
  assign \new_[3566]_  = \new_[1682]_  | \new_[3565]_ ;
  assign \new_[3567]_  = \new_[3566]_  | \new_[3561]_ ;
  assign \new_[3568]_  = \new_[3567]_  | \new_[3558]_ ;
  assign \new_[3569]_  = \new_[3568]_  | \new_[3551]_ ;
  assign \new_[3572]_  = \new_[1678]_  | \new_[1679]_ ;
  assign \new_[3575]_  = \new_[1676]_  | \new_[1677]_ ;
  assign \new_[3576]_  = \new_[3575]_  | \new_[3572]_ ;
  assign \new_[3579]_  = \new_[1674]_  | \new_[1675]_ ;
  assign \new_[3583]_  = \new_[1671]_  | \new_[1672]_ ;
  assign \new_[3584]_  = \new_[1673]_  | \new_[3583]_ ;
  assign \new_[3585]_  = \new_[3584]_  | \new_[3579]_ ;
  assign \new_[3586]_  = \new_[3585]_  | \new_[3576]_ ;
  assign \new_[3589]_  = \new_[1669]_  | \new_[1670]_ ;
  assign \new_[3592]_  = \new_[1667]_  | \new_[1668]_ ;
  assign \new_[3593]_  = \new_[3592]_  | \new_[3589]_ ;
  assign \new_[3596]_  = \new_[1665]_  | \new_[1666]_ ;
  assign \new_[3600]_  = \new_[1662]_  | \new_[1663]_ ;
  assign \new_[3601]_  = \new_[1664]_  | \new_[3600]_ ;
  assign \new_[3602]_  = \new_[3601]_  | \new_[3596]_ ;
  assign \new_[3603]_  = \new_[3602]_  | \new_[3593]_ ;
  assign \new_[3604]_  = \new_[3603]_  | \new_[3586]_ ;
  assign \new_[3605]_  = \new_[3604]_  | \new_[3569]_ ;
  assign \new_[3606]_  = \new_[3605]_  | \new_[3534]_ ;
  assign \new_[3609]_  = \new_[1660]_  | \new_[1661]_ ;
  assign \new_[3612]_  = \new_[1658]_  | \new_[1659]_ ;
  assign \new_[3613]_  = \new_[3612]_  | \new_[3609]_ ;
  assign \new_[3616]_  = \new_[1656]_  | \new_[1657]_ ;
  assign \new_[3620]_  = \new_[1653]_  | \new_[1654]_ ;
  assign \new_[3621]_  = \new_[1655]_  | \new_[3620]_ ;
  assign \new_[3622]_  = \new_[3621]_  | \new_[3616]_ ;
  assign \new_[3623]_  = \new_[3622]_  | \new_[3613]_ ;
  assign \new_[3626]_  = \new_[1651]_  | \new_[1652]_ ;
  assign \new_[3629]_  = \new_[1649]_  | \new_[1650]_ ;
  assign \new_[3630]_  = \new_[3629]_  | \new_[3626]_ ;
  assign \new_[3633]_  = \new_[1647]_  | \new_[1648]_ ;
  assign \new_[3637]_  = \new_[1644]_  | \new_[1645]_ ;
  assign \new_[3638]_  = \new_[1646]_  | \new_[3637]_ ;
  assign \new_[3639]_  = \new_[3638]_  | \new_[3633]_ ;
  assign \new_[3640]_  = \new_[3639]_  | \new_[3630]_ ;
  assign \new_[3641]_  = \new_[3640]_  | \new_[3623]_ ;
  assign \new_[3644]_  = \new_[1642]_  | \new_[1643]_ ;
  assign \new_[3647]_  = \new_[1640]_  | \new_[1641]_ ;
  assign \new_[3648]_  = \new_[3647]_  | \new_[3644]_ ;
  assign \new_[3651]_  = \new_[1638]_  | \new_[1639]_ ;
  assign \new_[3655]_  = \new_[1635]_  | \new_[1636]_ ;
  assign \new_[3656]_  = \new_[1637]_  | \new_[3655]_ ;
  assign \new_[3657]_  = \new_[3656]_  | \new_[3651]_ ;
  assign \new_[3658]_  = \new_[3657]_  | \new_[3648]_ ;
  assign \new_[3661]_  = \new_[1633]_  | \new_[1634]_ ;
  assign \new_[3664]_  = \new_[1631]_  | \new_[1632]_ ;
  assign \new_[3665]_  = \new_[3664]_  | \new_[3661]_ ;
  assign \new_[3668]_  = \new_[1629]_  | \new_[1630]_ ;
  assign \new_[3672]_  = \new_[1626]_  | \new_[1627]_ ;
  assign \new_[3673]_  = \new_[1628]_  | \new_[3672]_ ;
  assign \new_[3674]_  = \new_[3673]_  | \new_[3668]_ ;
  assign \new_[3675]_  = \new_[3674]_  | \new_[3665]_ ;
  assign \new_[3676]_  = \new_[3675]_  | \new_[3658]_ ;
  assign \new_[3677]_  = \new_[3676]_  | \new_[3641]_ ;
  assign \new_[3680]_  = \new_[1624]_  | \new_[1625]_ ;
  assign \new_[3683]_  = \new_[1622]_  | \new_[1623]_ ;
  assign \new_[3684]_  = \new_[3683]_  | \new_[3680]_ ;
  assign \new_[3687]_  = \new_[1620]_  | \new_[1621]_ ;
  assign \new_[3691]_  = \new_[1617]_  | \new_[1618]_ ;
  assign \new_[3692]_  = \new_[1619]_  | \new_[3691]_ ;
  assign \new_[3693]_  = \new_[3692]_  | \new_[3687]_ ;
  assign \new_[3694]_  = \new_[3693]_  | \new_[3684]_ ;
  assign \new_[3697]_  = \new_[1615]_  | \new_[1616]_ ;
  assign \new_[3700]_  = \new_[1613]_  | \new_[1614]_ ;
  assign \new_[3701]_  = \new_[3700]_  | \new_[3697]_ ;
  assign \new_[3704]_  = \new_[1611]_  | \new_[1612]_ ;
  assign \new_[3708]_  = \new_[1608]_  | \new_[1609]_ ;
  assign \new_[3709]_  = \new_[1610]_  | \new_[3708]_ ;
  assign \new_[3710]_  = \new_[3709]_  | \new_[3704]_ ;
  assign \new_[3711]_  = \new_[3710]_  | \new_[3701]_ ;
  assign \new_[3712]_  = \new_[3711]_  | \new_[3694]_ ;
  assign \new_[3715]_  = \new_[1606]_  | \new_[1607]_ ;
  assign \new_[3718]_  = \new_[1604]_  | \new_[1605]_ ;
  assign \new_[3719]_  = \new_[3718]_  | \new_[3715]_ ;
  assign \new_[3722]_  = \new_[1602]_  | \new_[1603]_ ;
  assign \new_[3726]_  = \new_[1599]_  | \new_[1600]_ ;
  assign \new_[3727]_  = \new_[1601]_  | \new_[3726]_ ;
  assign \new_[3728]_  = \new_[3727]_  | \new_[3722]_ ;
  assign \new_[3729]_  = \new_[3728]_  | \new_[3719]_ ;
  assign \new_[3732]_  = \new_[1597]_  | \new_[1598]_ ;
  assign \new_[3735]_  = \new_[1595]_  | \new_[1596]_ ;
  assign \new_[3736]_  = \new_[3735]_  | \new_[3732]_ ;
  assign \new_[3739]_  = \new_[1593]_  | \new_[1594]_ ;
  assign \new_[3743]_  = \new_[1590]_  | \new_[1591]_ ;
  assign \new_[3744]_  = \new_[1592]_  | \new_[3743]_ ;
  assign \new_[3745]_  = \new_[3744]_  | \new_[3739]_ ;
  assign \new_[3746]_  = \new_[3745]_  | \new_[3736]_ ;
  assign \new_[3747]_  = \new_[3746]_  | \new_[3729]_ ;
  assign \new_[3748]_  = \new_[3747]_  | \new_[3712]_ ;
  assign \new_[3749]_  = \new_[3748]_  | \new_[3677]_ ;
  assign \new_[3750]_  = \new_[3749]_  | \new_[3606]_ ;
  assign \new_[3753]_  = \new_[1588]_  | \new_[1589]_ ;
  assign \new_[3756]_  = \new_[1586]_  | \new_[1587]_ ;
  assign \new_[3757]_  = \new_[3756]_  | \new_[3753]_ ;
  assign \new_[3760]_  = \new_[1584]_  | \new_[1585]_ ;
  assign \new_[3764]_  = \new_[1581]_  | \new_[1582]_ ;
  assign \new_[3765]_  = \new_[1583]_  | \new_[3764]_ ;
  assign \new_[3766]_  = \new_[3765]_  | \new_[3760]_ ;
  assign \new_[3767]_  = \new_[3766]_  | \new_[3757]_ ;
  assign \new_[3770]_  = \new_[1579]_  | \new_[1580]_ ;
  assign \new_[3773]_  = \new_[1577]_  | \new_[1578]_ ;
  assign \new_[3774]_  = \new_[3773]_  | \new_[3770]_ ;
  assign \new_[3777]_  = \new_[1575]_  | \new_[1576]_ ;
  assign \new_[3781]_  = \new_[1572]_  | \new_[1573]_ ;
  assign \new_[3782]_  = \new_[1574]_  | \new_[3781]_ ;
  assign \new_[3783]_  = \new_[3782]_  | \new_[3777]_ ;
  assign \new_[3784]_  = \new_[3783]_  | \new_[3774]_ ;
  assign \new_[3785]_  = \new_[3784]_  | \new_[3767]_ ;
  assign \new_[3788]_  = \new_[1570]_  | \new_[1571]_ ;
  assign \new_[3791]_  = \new_[1568]_  | \new_[1569]_ ;
  assign \new_[3792]_  = \new_[3791]_  | \new_[3788]_ ;
  assign \new_[3795]_  = \new_[1566]_  | \new_[1567]_ ;
  assign \new_[3799]_  = \new_[1563]_  | \new_[1564]_ ;
  assign \new_[3800]_  = \new_[1565]_  | \new_[3799]_ ;
  assign \new_[3801]_  = \new_[3800]_  | \new_[3795]_ ;
  assign \new_[3802]_  = \new_[3801]_  | \new_[3792]_ ;
  assign \new_[3805]_  = \new_[1561]_  | \new_[1562]_ ;
  assign \new_[3808]_  = \new_[1559]_  | \new_[1560]_ ;
  assign \new_[3809]_  = \new_[3808]_  | \new_[3805]_ ;
  assign \new_[3812]_  = \new_[1557]_  | \new_[1558]_ ;
  assign \new_[3816]_  = \new_[1554]_  | \new_[1555]_ ;
  assign \new_[3817]_  = \new_[1556]_  | \new_[3816]_ ;
  assign \new_[3818]_  = \new_[3817]_  | \new_[3812]_ ;
  assign \new_[3819]_  = \new_[3818]_  | \new_[3809]_ ;
  assign \new_[3820]_  = \new_[3819]_  | \new_[3802]_ ;
  assign \new_[3821]_  = \new_[3820]_  | \new_[3785]_ ;
  assign \new_[3824]_  = \new_[1552]_  | \new_[1553]_ ;
  assign \new_[3827]_  = \new_[1550]_  | \new_[1551]_ ;
  assign \new_[3828]_  = \new_[3827]_  | \new_[3824]_ ;
  assign \new_[3831]_  = \new_[1548]_  | \new_[1549]_ ;
  assign \new_[3835]_  = \new_[1545]_  | \new_[1546]_ ;
  assign \new_[3836]_  = \new_[1547]_  | \new_[3835]_ ;
  assign \new_[3837]_  = \new_[3836]_  | \new_[3831]_ ;
  assign \new_[3838]_  = \new_[3837]_  | \new_[3828]_ ;
  assign \new_[3841]_  = \new_[1543]_  | \new_[1544]_ ;
  assign \new_[3844]_  = \new_[1541]_  | \new_[1542]_ ;
  assign \new_[3845]_  = \new_[3844]_  | \new_[3841]_ ;
  assign \new_[3848]_  = \new_[1539]_  | \new_[1540]_ ;
  assign \new_[3852]_  = \new_[1536]_  | \new_[1537]_ ;
  assign \new_[3853]_  = \new_[1538]_  | \new_[3852]_ ;
  assign \new_[3854]_  = \new_[3853]_  | \new_[3848]_ ;
  assign \new_[3855]_  = \new_[3854]_  | \new_[3845]_ ;
  assign \new_[3856]_  = \new_[3855]_  | \new_[3838]_ ;
  assign \new_[3859]_  = \new_[1534]_  | \new_[1535]_ ;
  assign \new_[3862]_  = \new_[1532]_  | \new_[1533]_ ;
  assign \new_[3863]_  = \new_[3862]_  | \new_[3859]_ ;
  assign \new_[3866]_  = \new_[1530]_  | \new_[1531]_ ;
  assign \new_[3870]_  = \new_[1527]_  | \new_[1528]_ ;
  assign \new_[3871]_  = \new_[1529]_  | \new_[3870]_ ;
  assign \new_[3872]_  = \new_[3871]_  | \new_[3866]_ ;
  assign \new_[3873]_  = \new_[3872]_  | \new_[3863]_ ;
  assign \new_[3876]_  = \new_[1525]_  | \new_[1526]_ ;
  assign \new_[3879]_  = \new_[1523]_  | \new_[1524]_ ;
  assign \new_[3880]_  = \new_[3879]_  | \new_[3876]_ ;
  assign \new_[3883]_  = \new_[1521]_  | \new_[1522]_ ;
  assign \new_[3887]_  = \new_[1518]_  | \new_[1519]_ ;
  assign \new_[3888]_  = \new_[1520]_  | \new_[3887]_ ;
  assign \new_[3889]_  = \new_[3888]_  | \new_[3883]_ ;
  assign \new_[3890]_  = \new_[3889]_  | \new_[3880]_ ;
  assign \new_[3891]_  = \new_[3890]_  | \new_[3873]_ ;
  assign \new_[3892]_  = \new_[3891]_  | \new_[3856]_ ;
  assign \new_[3893]_  = \new_[3892]_  | \new_[3821]_ ;
  assign \new_[3896]_  = \new_[1516]_  | \new_[1517]_ ;
  assign \new_[3899]_  = \new_[1514]_  | \new_[1515]_ ;
  assign \new_[3900]_  = \new_[3899]_  | \new_[3896]_ ;
  assign \new_[3903]_  = \new_[1512]_  | \new_[1513]_ ;
  assign \new_[3907]_  = \new_[1509]_  | \new_[1510]_ ;
  assign \new_[3908]_  = \new_[1511]_  | \new_[3907]_ ;
  assign \new_[3909]_  = \new_[3908]_  | \new_[3903]_ ;
  assign \new_[3910]_  = \new_[3909]_  | \new_[3900]_ ;
  assign \new_[3913]_  = \new_[1507]_  | \new_[1508]_ ;
  assign \new_[3916]_  = \new_[1505]_  | \new_[1506]_ ;
  assign \new_[3917]_  = \new_[3916]_  | \new_[3913]_ ;
  assign \new_[3920]_  = \new_[1503]_  | \new_[1504]_ ;
  assign \new_[3924]_  = \new_[1500]_  | \new_[1501]_ ;
  assign \new_[3925]_  = \new_[1502]_  | \new_[3924]_ ;
  assign \new_[3926]_  = \new_[3925]_  | \new_[3920]_ ;
  assign \new_[3927]_  = \new_[3926]_  | \new_[3917]_ ;
  assign \new_[3928]_  = \new_[3927]_  | \new_[3910]_ ;
  assign \new_[3931]_  = \new_[1498]_  | \new_[1499]_ ;
  assign \new_[3934]_  = \new_[1496]_  | \new_[1497]_ ;
  assign \new_[3935]_  = \new_[3934]_  | \new_[3931]_ ;
  assign \new_[3938]_  = \new_[1494]_  | \new_[1495]_ ;
  assign \new_[3942]_  = \new_[1491]_  | \new_[1492]_ ;
  assign \new_[3943]_  = \new_[1493]_  | \new_[3942]_ ;
  assign \new_[3944]_  = \new_[3943]_  | \new_[3938]_ ;
  assign \new_[3945]_  = \new_[3944]_  | \new_[3935]_ ;
  assign \new_[3948]_  = \new_[1489]_  | \new_[1490]_ ;
  assign \new_[3951]_  = \new_[1487]_  | \new_[1488]_ ;
  assign \new_[3952]_  = \new_[3951]_  | \new_[3948]_ ;
  assign \new_[3955]_  = \new_[1485]_  | \new_[1486]_ ;
  assign \new_[3959]_  = \new_[1482]_  | \new_[1483]_ ;
  assign \new_[3960]_  = \new_[1484]_  | \new_[3959]_ ;
  assign \new_[3961]_  = \new_[3960]_  | \new_[3955]_ ;
  assign \new_[3962]_  = \new_[3961]_  | \new_[3952]_ ;
  assign \new_[3963]_  = \new_[3962]_  | \new_[3945]_ ;
  assign \new_[3964]_  = \new_[3963]_  | \new_[3928]_ ;
  assign \new_[3967]_  = \new_[1480]_  | \new_[1481]_ ;
  assign \new_[3970]_  = \new_[1478]_  | \new_[1479]_ ;
  assign \new_[3971]_  = \new_[3970]_  | \new_[3967]_ ;
  assign \new_[3974]_  = \new_[1476]_  | \new_[1477]_ ;
  assign \new_[3978]_  = \new_[1473]_  | \new_[1474]_ ;
  assign \new_[3979]_  = \new_[1475]_  | \new_[3978]_ ;
  assign \new_[3980]_  = \new_[3979]_  | \new_[3974]_ ;
  assign \new_[3981]_  = \new_[3980]_  | \new_[3971]_ ;
  assign \new_[3984]_  = \new_[1471]_  | \new_[1472]_ ;
  assign \new_[3987]_  = \new_[1469]_  | \new_[1470]_ ;
  assign \new_[3988]_  = \new_[3987]_  | \new_[3984]_ ;
  assign \new_[3991]_  = \new_[1467]_  | \new_[1468]_ ;
  assign \new_[3995]_  = \new_[1464]_  | \new_[1465]_ ;
  assign \new_[3996]_  = \new_[1466]_  | \new_[3995]_ ;
  assign \new_[3997]_  = \new_[3996]_  | \new_[3991]_ ;
  assign \new_[3998]_  = \new_[3997]_  | \new_[3988]_ ;
  assign \new_[3999]_  = \new_[3998]_  | \new_[3981]_ ;
  assign \new_[4002]_  = \new_[1462]_  | \new_[1463]_ ;
  assign \new_[4005]_  = \new_[1460]_  | \new_[1461]_ ;
  assign \new_[4006]_  = \new_[4005]_  | \new_[4002]_ ;
  assign \new_[4009]_  = \new_[1458]_  | \new_[1459]_ ;
  assign \new_[4013]_  = \new_[1455]_  | \new_[1456]_ ;
  assign \new_[4014]_  = \new_[1457]_  | \new_[4013]_ ;
  assign \new_[4015]_  = \new_[4014]_  | \new_[4009]_ ;
  assign \new_[4016]_  = \new_[4015]_  | \new_[4006]_ ;
  assign \new_[4019]_  = \new_[1453]_  | \new_[1454]_ ;
  assign \new_[4023]_  = \new_[1450]_  | \new_[1451]_ ;
  assign \new_[4024]_  = \new_[1452]_  | \new_[4023]_ ;
  assign \new_[4025]_  = \new_[4024]_  | \new_[4019]_ ;
  assign \new_[4028]_  = \new_[1448]_  | \new_[1449]_ ;
  assign \new_[4032]_  = \new_[1445]_  | \new_[1446]_ ;
  assign \new_[4033]_  = \new_[1447]_  | \new_[4032]_ ;
  assign \new_[4034]_  = \new_[4033]_  | \new_[4028]_ ;
  assign \new_[4035]_  = \new_[4034]_  | \new_[4025]_ ;
  assign \new_[4036]_  = \new_[4035]_  | \new_[4016]_ ;
  assign \new_[4037]_  = \new_[4036]_  | \new_[3999]_ ;
  assign \new_[4038]_  = \new_[4037]_  | \new_[3964]_ ;
  assign \new_[4039]_  = \new_[4038]_  | \new_[3893]_ ;
  assign \new_[4040]_  = \new_[4039]_  | \new_[3750]_ ;
  assign \new_[4043]_  = \new_[1443]_  | \new_[1444]_ ;
  assign \new_[4046]_  = \new_[1441]_  | \new_[1442]_ ;
  assign \new_[4047]_  = \new_[4046]_  | \new_[4043]_ ;
  assign \new_[4050]_  = \new_[1439]_  | \new_[1440]_ ;
  assign \new_[4054]_  = \new_[1436]_  | \new_[1437]_ ;
  assign \new_[4055]_  = \new_[1438]_  | \new_[4054]_ ;
  assign \new_[4056]_  = \new_[4055]_  | \new_[4050]_ ;
  assign \new_[4057]_  = \new_[4056]_  | \new_[4047]_ ;
  assign \new_[4060]_  = \new_[1434]_  | \new_[1435]_ ;
  assign \new_[4063]_  = \new_[1432]_  | \new_[1433]_ ;
  assign \new_[4064]_  = \new_[4063]_  | \new_[4060]_ ;
  assign \new_[4067]_  = \new_[1430]_  | \new_[1431]_ ;
  assign \new_[4071]_  = \new_[1427]_  | \new_[1428]_ ;
  assign \new_[4072]_  = \new_[1429]_  | \new_[4071]_ ;
  assign \new_[4073]_  = \new_[4072]_  | \new_[4067]_ ;
  assign \new_[4074]_  = \new_[4073]_  | \new_[4064]_ ;
  assign \new_[4075]_  = \new_[4074]_  | \new_[4057]_ ;
  assign \new_[4078]_  = \new_[1425]_  | \new_[1426]_ ;
  assign \new_[4081]_  = \new_[1423]_  | \new_[1424]_ ;
  assign \new_[4082]_  = \new_[4081]_  | \new_[4078]_ ;
  assign \new_[4085]_  = \new_[1421]_  | \new_[1422]_ ;
  assign \new_[4089]_  = \new_[1418]_  | \new_[1419]_ ;
  assign \new_[4090]_  = \new_[1420]_  | \new_[4089]_ ;
  assign \new_[4091]_  = \new_[4090]_  | \new_[4085]_ ;
  assign \new_[4092]_  = \new_[4091]_  | \new_[4082]_ ;
  assign \new_[4095]_  = \new_[1416]_  | \new_[1417]_ ;
  assign \new_[4098]_  = \new_[1414]_  | \new_[1415]_ ;
  assign \new_[4099]_  = \new_[4098]_  | \new_[4095]_ ;
  assign \new_[4102]_  = \new_[1412]_  | \new_[1413]_ ;
  assign \new_[4106]_  = \new_[1409]_  | \new_[1410]_ ;
  assign \new_[4107]_  = \new_[1411]_  | \new_[4106]_ ;
  assign \new_[4108]_  = \new_[4107]_  | \new_[4102]_ ;
  assign \new_[4109]_  = \new_[4108]_  | \new_[4099]_ ;
  assign \new_[4110]_  = \new_[4109]_  | \new_[4092]_ ;
  assign \new_[4111]_  = \new_[4110]_  | \new_[4075]_ ;
  assign \new_[4114]_  = \new_[1407]_  | \new_[1408]_ ;
  assign \new_[4117]_  = \new_[1405]_  | \new_[1406]_ ;
  assign \new_[4118]_  = \new_[4117]_  | \new_[4114]_ ;
  assign \new_[4121]_  = \new_[1403]_  | \new_[1404]_ ;
  assign \new_[4125]_  = \new_[1400]_  | \new_[1401]_ ;
  assign \new_[4126]_  = \new_[1402]_  | \new_[4125]_ ;
  assign \new_[4127]_  = \new_[4126]_  | \new_[4121]_ ;
  assign \new_[4128]_  = \new_[4127]_  | \new_[4118]_ ;
  assign \new_[4131]_  = \new_[1398]_  | \new_[1399]_ ;
  assign \new_[4134]_  = \new_[1396]_  | \new_[1397]_ ;
  assign \new_[4135]_  = \new_[4134]_  | \new_[4131]_ ;
  assign \new_[4138]_  = \new_[1394]_  | \new_[1395]_ ;
  assign \new_[4142]_  = \new_[1391]_  | \new_[1392]_ ;
  assign \new_[4143]_  = \new_[1393]_  | \new_[4142]_ ;
  assign \new_[4144]_  = \new_[4143]_  | \new_[4138]_ ;
  assign \new_[4145]_  = \new_[4144]_  | \new_[4135]_ ;
  assign \new_[4146]_  = \new_[4145]_  | \new_[4128]_ ;
  assign \new_[4149]_  = \new_[1389]_  | \new_[1390]_ ;
  assign \new_[4152]_  = \new_[1387]_  | \new_[1388]_ ;
  assign \new_[4153]_  = \new_[4152]_  | \new_[4149]_ ;
  assign \new_[4156]_  = \new_[1385]_  | \new_[1386]_ ;
  assign \new_[4160]_  = \new_[1382]_  | \new_[1383]_ ;
  assign \new_[4161]_  = \new_[1384]_  | \new_[4160]_ ;
  assign \new_[4162]_  = \new_[4161]_  | \new_[4156]_ ;
  assign \new_[4163]_  = \new_[4162]_  | \new_[4153]_ ;
  assign \new_[4166]_  = \new_[1380]_  | \new_[1381]_ ;
  assign \new_[4169]_  = \new_[1378]_  | \new_[1379]_ ;
  assign \new_[4170]_  = \new_[4169]_  | \new_[4166]_ ;
  assign \new_[4173]_  = \new_[1376]_  | \new_[1377]_ ;
  assign \new_[4177]_  = \new_[1373]_  | \new_[1374]_ ;
  assign \new_[4178]_  = \new_[1375]_  | \new_[4177]_ ;
  assign \new_[4179]_  = \new_[4178]_  | \new_[4173]_ ;
  assign \new_[4180]_  = \new_[4179]_  | \new_[4170]_ ;
  assign \new_[4181]_  = \new_[4180]_  | \new_[4163]_ ;
  assign \new_[4182]_  = \new_[4181]_  | \new_[4146]_ ;
  assign \new_[4183]_  = \new_[4182]_  | \new_[4111]_ ;
  assign \new_[4186]_  = \new_[1371]_  | \new_[1372]_ ;
  assign \new_[4189]_  = \new_[1369]_  | \new_[1370]_ ;
  assign \new_[4190]_  = \new_[4189]_  | \new_[4186]_ ;
  assign \new_[4193]_  = \new_[1367]_  | \new_[1368]_ ;
  assign \new_[4197]_  = \new_[1364]_  | \new_[1365]_ ;
  assign \new_[4198]_  = \new_[1366]_  | \new_[4197]_ ;
  assign \new_[4199]_  = \new_[4198]_  | \new_[4193]_ ;
  assign \new_[4200]_  = \new_[4199]_  | \new_[4190]_ ;
  assign \new_[4203]_  = \new_[1362]_  | \new_[1363]_ ;
  assign \new_[4206]_  = \new_[1360]_  | \new_[1361]_ ;
  assign \new_[4207]_  = \new_[4206]_  | \new_[4203]_ ;
  assign \new_[4210]_  = \new_[1358]_  | \new_[1359]_ ;
  assign \new_[4214]_  = \new_[1355]_  | \new_[1356]_ ;
  assign \new_[4215]_  = \new_[1357]_  | \new_[4214]_ ;
  assign \new_[4216]_  = \new_[4215]_  | \new_[4210]_ ;
  assign \new_[4217]_  = \new_[4216]_  | \new_[4207]_ ;
  assign \new_[4218]_  = \new_[4217]_  | \new_[4200]_ ;
  assign \new_[4221]_  = \new_[1353]_  | \new_[1354]_ ;
  assign \new_[4224]_  = \new_[1351]_  | \new_[1352]_ ;
  assign \new_[4225]_  = \new_[4224]_  | \new_[4221]_ ;
  assign \new_[4228]_  = \new_[1349]_  | \new_[1350]_ ;
  assign \new_[4232]_  = \new_[1346]_  | \new_[1347]_ ;
  assign \new_[4233]_  = \new_[1348]_  | \new_[4232]_ ;
  assign \new_[4234]_  = \new_[4233]_  | \new_[4228]_ ;
  assign \new_[4235]_  = \new_[4234]_  | \new_[4225]_ ;
  assign \new_[4238]_  = \new_[1344]_  | \new_[1345]_ ;
  assign \new_[4241]_  = \new_[1342]_  | \new_[1343]_ ;
  assign \new_[4242]_  = \new_[4241]_  | \new_[4238]_ ;
  assign \new_[4245]_  = \new_[1340]_  | \new_[1341]_ ;
  assign \new_[4249]_  = \new_[1337]_  | \new_[1338]_ ;
  assign \new_[4250]_  = \new_[1339]_  | \new_[4249]_ ;
  assign \new_[4251]_  = \new_[4250]_  | \new_[4245]_ ;
  assign \new_[4252]_  = \new_[4251]_  | \new_[4242]_ ;
  assign \new_[4253]_  = \new_[4252]_  | \new_[4235]_ ;
  assign \new_[4254]_  = \new_[4253]_  | \new_[4218]_ ;
  assign \new_[4257]_  = \new_[1335]_  | \new_[1336]_ ;
  assign \new_[4260]_  = \new_[1333]_  | \new_[1334]_ ;
  assign \new_[4261]_  = \new_[4260]_  | \new_[4257]_ ;
  assign \new_[4264]_  = \new_[1331]_  | \new_[1332]_ ;
  assign \new_[4268]_  = \new_[1328]_  | \new_[1329]_ ;
  assign \new_[4269]_  = \new_[1330]_  | \new_[4268]_ ;
  assign \new_[4270]_  = \new_[4269]_  | \new_[4264]_ ;
  assign \new_[4271]_  = \new_[4270]_  | \new_[4261]_ ;
  assign \new_[4274]_  = \new_[1326]_  | \new_[1327]_ ;
  assign \new_[4277]_  = \new_[1324]_  | \new_[1325]_ ;
  assign \new_[4278]_  = \new_[4277]_  | \new_[4274]_ ;
  assign \new_[4281]_  = \new_[1322]_  | \new_[1323]_ ;
  assign \new_[4285]_  = \new_[1319]_  | \new_[1320]_ ;
  assign \new_[4286]_  = \new_[1321]_  | \new_[4285]_ ;
  assign \new_[4287]_  = \new_[4286]_  | \new_[4281]_ ;
  assign \new_[4288]_  = \new_[4287]_  | \new_[4278]_ ;
  assign \new_[4289]_  = \new_[4288]_  | \new_[4271]_ ;
  assign \new_[4292]_  = \new_[1317]_  | \new_[1318]_ ;
  assign \new_[4295]_  = \new_[1315]_  | \new_[1316]_ ;
  assign \new_[4296]_  = \new_[4295]_  | \new_[4292]_ ;
  assign \new_[4299]_  = \new_[1313]_  | \new_[1314]_ ;
  assign \new_[4303]_  = \new_[1310]_  | \new_[1311]_ ;
  assign \new_[4304]_  = \new_[1312]_  | \new_[4303]_ ;
  assign \new_[4305]_  = \new_[4304]_  | \new_[4299]_ ;
  assign \new_[4306]_  = \new_[4305]_  | \new_[4296]_ ;
  assign \new_[4309]_  = \new_[1308]_  | \new_[1309]_ ;
  assign \new_[4312]_  = \new_[1306]_  | \new_[1307]_ ;
  assign \new_[4313]_  = \new_[4312]_  | \new_[4309]_ ;
  assign \new_[4316]_  = \new_[1304]_  | \new_[1305]_ ;
  assign \new_[4320]_  = \new_[1301]_  | \new_[1302]_ ;
  assign \new_[4321]_  = \new_[1303]_  | \new_[4320]_ ;
  assign \new_[4322]_  = \new_[4321]_  | \new_[4316]_ ;
  assign \new_[4323]_  = \new_[4322]_  | \new_[4313]_ ;
  assign \new_[4324]_  = \new_[4323]_  | \new_[4306]_ ;
  assign \new_[4325]_  = \new_[4324]_  | \new_[4289]_ ;
  assign \new_[4326]_  = \new_[4325]_  | \new_[4254]_ ;
  assign \new_[4327]_  = \new_[4326]_  | \new_[4183]_ ;
  assign \new_[4330]_  = \new_[1299]_  | \new_[1300]_ ;
  assign \new_[4333]_  = \new_[1297]_  | \new_[1298]_ ;
  assign \new_[4334]_  = \new_[4333]_  | \new_[4330]_ ;
  assign \new_[4337]_  = \new_[1295]_  | \new_[1296]_ ;
  assign \new_[4341]_  = \new_[1292]_  | \new_[1293]_ ;
  assign \new_[4342]_  = \new_[1294]_  | \new_[4341]_ ;
  assign \new_[4343]_  = \new_[4342]_  | \new_[4337]_ ;
  assign \new_[4344]_  = \new_[4343]_  | \new_[4334]_ ;
  assign \new_[4347]_  = \new_[1290]_  | \new_[1291]_ ;
  assign \new_[4350]_  = \new_[1288]_  | \new_[1289]_ ;
  assign \new_[4351]_  = \new_[4350]_  | \new_[4347]_ ;
  assign \new_[4354]_  = \new_[1286]_  | \new_[1287]_ ;
  assign \new_[4358]_  = \new_[1283]_  | \new_[1284]_ ;
  assign \new_[4359]_  = \new_[1285]_  | \new_[4358]_ ;
  assign \new_[4360]_  = \new_[4359]_  | \new_[4354]_ ;
  assign \new_[4361]_  = \new_[4360]_  | \new_[4351]_ ;
  assign \new_[4362]_  = \new_[4361]_  | \new_[4344]_ ;
  assign \new_[4365]_  = \new_[1281]_  | \new_[1282]_ ;
  assign \new_[4368]_  = \new_[1279]_  | \new_[1280]_ ;
  assign \new_[4369]_  = \new_[4368]_  | \new_[4365]_ ;
  assign \new_[4372]_  = \new_[1277]_  | \new_[1278]_ ;
  assign \new_[4376]_  = \new_[1274]_  | \new_[1275]_ ;
  assign \new_[4377]_  = \new_[1276]_  | \new_[4376]_ ;
  assign \new_[4378]_  = \new_[4377]_  | \new_[4372]_ ;
  assign \new_[4379]_  = \new_[4378]_  | \new_[4369]_ ;
  assign \new_[4382]_  = \new_[1272]_  | \new_[1273]_ ;
  assign \new_[4385]_  = \new_[1270]_  | \new_[1271]_ ;
  assign \new_[4386]_  = \new_[4385]_  | \new_[4382]_ ;
  assign \new_[4389]_  = \new_[1268]_  | \new_[1269]_ ;
  assign \new_[4393]_  = \new_[1265]_  | \new_[1266]_ ;
  assign \new_[4394]_  = \new_[1267]_  | \new_[4393]_ ;
  assign \new_[4395]_  = \new_[4394]_  | \new_[4389]_ ;
  assign \new_[4396]_  = \new_[4395]_  | \new_[4386]_ ;
  assign \new_[4397]_  = \new_[4396]_  | \new_[4379]_ ;
  assign \new_[4398]_  = \new_[4397]_  | \new_[4362]_ ;
  assign \new_[4401]_  = \new_[1263]_  | \new_[1264]_ ;
  assign \new_[4404]_  = \new_[1261]_  | \new_[1262]_ ;
  assign \new_[4405]_  = \new_[4404]_  | \new_[4401]_ ;
  assign \new_[4408]_  = \new_[1259]_  | \new_[1260]_ ;
  assign \new_[4412]_  = \new_[1256]_  | \new_[1257]_ ;
  assign \new_[4413]_  = \new_[1258]_  | \new_[4412]_ ;
  assign \new_[4414]_  = \new_[4413]_  | \new_[4408]_ ;
  assign \new_[4415]_  = \new_[4414]_  | \new_[4405]_ ;
  assign \new_[4418]_  = \new_[1254]_  | \new_[1255]_ ;
  assign \new_[4421]_  = \new_[1252]_  | \new_[1253]_ ;
  assign \new_[4422]_  = \new_[4421]_  | \new_[4418]_ ;
  assign \new_[4425]_  = \new_[1250]_  | \new_[1251]_ ;
  assign \new_[4429]_  = \new_[1247]_  | \new_[1248]_ ;
  assign \new_[4430]_  = \new_[1249]_  | \new_[4429]_ ;
  assign \new_[4431]_  = \new_[4430]_  | \new_[4425]_ ;
  assign \new_[4432]_  = \new_[4431]_  | \new_[4422]_ ;
  assign \new_[4433]_  = \new_[4432]_  | \new_[4415]_ ;
  assign \new_[4436]_  = \new_[1245]_  | \new_[1246]_ ;
  assign \new_[4439]_  = \new_[1243]_  | \new_[1244]_ ;
  assign \new_[4440]_  = \new_[4439]_  | \new_[4436]_ ;
  assign \new_[4443]_  = \new_[1241]_  | \new_[1242]_ ;
  assign \new_[4447]_  = \new_[1238]_  | \new_[1239]_ ;
  assign \new_[4448]_  = \new_[1240]_  | \new_[4447]_ ;
  assign \new_[4449]_  = \new_[4448]_  | \new_[4443]_ ;
  assign \new_[4450]_  = \new_[4449]_  | \new_[4440]_ ;
  assign \new_[4453]_  = \new_[1236]_  | \new_[1237]_ ;
  assign \new_[4456]_  = \new_[1234]_  | \new_[1235]_ ;
  assign \new_[4457]_  = \new_[4456]_  | \new_[4453]_ ;
  assign \new_[4460]_  = \new_[1232]_  | \new_[1233]_ ;
  assign \new_[4464]_  = \new_[1229]_  | \new_[1230]_ ;
  assign \new_[4465]_  = \new_[1231]_  | \new_[4464]_ ;
  assign \new_[4466]_  = \new_[4465]_  | \new_[4460]_ ;
  assign \new_[4467]_  = \new_[4466]_  | \new_[4457]_ ;
  assign \new_[4468]_  = \new_[4467]_  | \new_[4450]_ ;
  assign \new_[4469]_  = \new_[4468]_  | \new_[4433]_ ;
  assign \new_[4470]_  = \new_[4469]_  | \new_[4398]_ ;
  assign \new_[4473]_  = \new_[1227]_  | \new_[1228]_ ;
  assign \new_[4476]_  = \new_[1225]_  | \new_[1226]_ ;
  assign \new_[4477]_  = \new_[4476]_  | \new_[4473]_ ;
  assign \new_[4480]_  = \new_[1223]_  | \new_[1224]_ ;
  assign \new_[4484]_  = \new_[1220]_  | \new_[1221]_ ;
  assign \new_[4485]_  = \new_[1222]_  | \new_[4484]_ ;
  assign \new_[4486]_  = \new_[4485]_  | \new_[4480]_ ;
  assign \new_[4487]_  = \new_[4486]_  | \new_[4477]_ ;
  assign \new_[4490]_  = \new_[1218]_  | \new_[1219]_ ;
  assign \new_[4493]_  = \new_[1216]_  | \new_[1217]_ ;
  assign \new_[4494]_  = \new_[4493]_  | \new_[4490]_ ;
  assign \new_[4497]_  = \new_[1214]_  | \new_[1215]_ ;
  assign \new_[4501]_  = \new_[1211]_  | \new_[1212]_ ;
  assign \new_[4502]_  = \new_[1213]_  | \new_[4501]_ ;
  assign \new_[4503]_  = \new_[4502]_  | \new_[4497]_ ;
  assign \new_[4504]_  = \new_[4503]_  | \new_[4494]_ ;
  assign \new_[4505]_  = \new_[4504]_  | \new_[4487]_ ;
  assign \new_[4508]_  = \new_[1209]_  | \new_[1210]_ ;
  assign \new_[4511]_  = \new_[1207]_  | \new_[1208]_ ;
  assign \new_[4512]_  = \new_[4511]_  | \new_[4508]_ ;
  assign \new_[4515]_  = \new_[1205]_  | \new_[1206]_ ;
  assign \new_[4519]_  = \new_[1202]_  | \new_[1203]_ ;
  assign \new_[4520]_  = \new_[1204]_  | \new_[4519]_ ;
  assign \new_[4521]_  = \new_[4520]_  | \new_[4515]_ ;
  assign \new_[4522]_  = \new_[4521]_  | \new_[4512]_ ;
  assign \new_[4525]_  = \new_[1200]_  | \new_[1201]_ ;
  assign \new_[4528]_  = \new_[1198]_  | \new_[1199]_ ;
  assign \new_[4529]_  = \new_[4528]_  | \new_[4525]_ ;
  assign \new_[4532]_  = \new_[1196]_  | \new_[1197]_ ;
  assign \new_[4536]_  = \new_[1193]_  | \new_[1194]_ ;
  assign \new_[4537]_  = \new_[1195]_  | \new_[4536]_ ;
  assign \new_[4538]_  = \new_[4537]_  | \new_[4532]_ ;
  assign \new_[4539]_  = \new_[4538]_  | \new_[4529]_ ;
  assign \new_[4540]_  = \new_[4539]_  | \new_[4522]_ ;
  assign \new_[4541]_  = \new_[4540]_  | \new_[4505]_ ;
  assign \new_[4544]_  = \new_[1191]_  | \new_[1192]_ ;
  assign \new_[4547]_  = \new_[1189]_  | \new_[1190]_ ;
  assign \new_[4548]_  = \new_[4547]_  | \new_[4544]_ ;
  assign \new_[4551]_  = \new_[1187]_  | \new_[1188]_ ;
  assign \new_[4555]_  = \new_[1184]_  | \new_[1185]_ ;
  assign \new_[4556]_  = \new_[1186]_  | \new_[4555]_ ;
  assign \new_[4557]_  = \new_[4556]_  | \new_[4551]_ ;
  assign \new_[4558]_  = \new_[4557]_  | \new_[4548]_ ;
  assign \new_[4561]_  = \new_[1182]_  | \new_[1183]_ ;
  assign \new_[4564]_  = \new_[1180]_  | \new_[1181]_ ;
  assign \new_[4565]_  = \new_[4564]_  | \new_[4561]_ ;
  assign \new_[4568]_  = \new_[1178]_  | \new_[1179]_ ;
  assign \new_[4572]_  = \new_[1175]_  | \new_[1176]_ ;
  assign \new_[4573]_  = \new_[1177]_  | \new_[4572]_ ;
  assign \new_[4574]_  = \new_[4573]_  | \new_[4568]_ ;
  assign \new_[4575]_  = \new_[4574]_  | \new_[4565]_ ;
  assign \new_[4576]_  = \new_[4575]_  | \new_[4558]_ ;
  assign \new_[4579]_  = \new_[1173]_  | \new_[1174]_ ;
  assign \new_[4582]_  = \new_[1171]_  | \new_[1172]_ ;
  assign \new_[4583]_  = \new_[4582]_  | \new_[4579]_ ;
  assign \new_[4586]_  = \new_[1169]_  | \new_[1170]_ ;
  assign \new_[4590]_  = \new_[1166]_  | \new_[1167]_ ;
  assign \new_[4591]_  = \new_[1168]_  | \new_[4590]_ ;
  assign \new_[4592]_  = \new_[4591]_  | \new_[4586]_ ;
  assign \new_[4593]_  = \new_[4592]_  | \new_[4583]_ ;
  assign \new_[4596]_  = \new_[1164]_  | \new_[1165]_ ;
  assign \new_[4600]_  = \new_[1161]_  | \new_[1162]_ ;
  assign \new_[4601]_  = \new_[1163]_  | \new_[4600]_ ;
  assign \new_[4602]_  = \new_[4601]_  | \new_[4596]_ ;
  assign \new_[4605]_  = \new_[1159]_  | \new_[1160]_ ;
  assign \new_[4609]_  = \new_[1156]_  | \new_[1157]_ ;
  assign \new_[4610]_  = \new_[1158]_  | \new_[4609]_ ;
  assign \new_[4611]_  = \new_[4610]_  | \new_[4605]_ ;
  assign \new_[4612]_  = \new_[4611]_  | \new_[4602]_ ;
  assign \new_[4613]_  = \new_[4612]_  | \new_[4593]_ ;
  assign \new_[4614]_  = \new_[4613]_  | \new_[4576]_ ;
  assign \new_[4615]_  = \new_[4614]_  | \new_[4541]_ ;
  assign \new_[4616]_  = \new_[4615]_  | \new_[4470]_ ;
  assign \new_[4617]_  = \new_[4616]_  | \new_[4327]_ ;
  assign \new_[4618]_  = \new_[4617]_  | \new_[4040]_ ;
  assign \new_[4619]_  = \new_[4618]_  | \new_[3463]_ ;
  assign \new_[4622]_  = \new_[1154]_  | \new_[1155]_ ;
  assign \new_[4625]_  = \new_[1152]_  | \new_[1153]_ ;
  assign \new_[4626]_  = \new_[4625]_  | \new_[4622]_ ;
  assign \new_[4629]_  = \new_[1150]_  | \new_[1151]_ ;
  assign \new_[4633]_  = \new_[1147]_  | \new_[1148]_ ;
  assign \new_[4634]_  = \new_[1149]_  | \new_[4633]_ ;
  assign \new_[4635]_  = \new_[4634]_  | \new_[4629]_ ;
  assign \new_[4636]_  = \new_[4635]_  | \new_[4626]_ ;
  assign \new_[4639]_  = \new_[1145]_  | \new_[1146]_ ;
  assign \new_[4642]_  = \new_[1143]_  | \new_[1144]_ ;
  assign \new_[4643]_  = \new_[4642]_  | \new_[4639]_ ;
  assign \new_[4646]_  = \new_[1141]_  | \new_[1142]_ ;
  assign \new_[4650]_  = \new_[1138]_  | \new_[1139]_ ;
  assign \new_[4651]_  = \new_[1140]_  | \new_[4650]_ ;
  assign \new_[4652]_  = \new_[4651]_  | \new_[4646]_ ;
  assign \new_[4653]_  = \new_[4652]_  | \new_[4643]_ ;
  assign \new_[4654]_  = \new_[4653]_  | \new_[4636]_ ;
  assign \new_[4657]_  = \new_[1136]_  | \new_[1137]_ ;
  assign \new_[4660]_  = \new_[1134]_  | \new_[1135]_ ;
  assign \new_[4661]_  = \new_[4660]_  | \new_[4657]_ ;
  assign \new_[4664]_  = \new_[1132]_  | \new_[1133]_ ;
  assign \new_[4668]_  = \new_[1129]_  | \new_[1130]_ ;
  assign \new_[4669]_  = \new_[1131]_  | \new_[4668]_ ;
  assign \new_[4670]_  = \new_[4669]_  | \new_[4664]_ ;
  assign \new_[4671]_  = \new_[4670]_  | \new_[4661]_ ;
  assign \new_[4674]_  = \new_[1127]_  | \new_[1128]_ ;
  assign \new_[4677]_  = \new_[1125]_  | \new_[1126]_ ;
  assign \new_[4678]_  = \new_[4677]_  | \new_[4674]_ ;
  assign \new_[4681]_  = \new_[1123]_  | \new_[1124]_ ;
  assign \new_[4685]_  = \new_[1120]_  | \new_[1121]_ ;
  assign \new_[4686]_  = \new_[1122]_  | \new_[4685]_ ;
  assign \new_[4687]_  = \new_[4686]_  | \new_[4681]_ ;
  assign \new_[4688]_  = \new_[4687]_  | \new_[4678]_ ;
  assign \new_[4689]_  = \new_[4688]_  | \new_[4671]_ ;
  assign \new_[4690]_  = \new_[4689]_  | \new_[4654]_ ;
  assign \new_[4693]_  = \new_[1118]_  | \new_[1119]_ ;
  assign \new_[4696]_  = \new_[1116]_  | \new_[1117]_ ;
  assign \new_[4697]_  = \new_[4696]_  | \new_[4693]_ ;
  assign \new_[4700]_  = \new_[1114]_  | \new_[1115]_ ;
  assign \new_[4704]_  = \new_[1111]_  | \new_[1112]_ ;
  assign \new_[4705]_  = \new_[1113]_  | \new_[4704]_ ;
  assign \new_[4706]_  = \new_[4705]_  | \new_[4700]_ ;
  assign \new_[4707]_  = \new_[4706]_  | \new_[4697]_ ;
  assign \new_[4710]_  = \new_[1109]_  | \new_[1110]_ ;
  assign \new_[4713]_  = \new_[1107]_  | \new_[1108]_ ;
  assign \new_[4714]_  = \new_[4713]_  | \new_[4710]_ ;
  assign \new_[4717]_  = \new_[1105]_  | \new_[1106]_ ;
  assign \new_[4721]_  = \new_[1102]_  | \new_[1103]_ ;
  assign \new_[4722]_  = \new_[1104]_  | \new_[4721]_ ;
  assign \new_[4723]_  = \new_[4722]_  | \new_[4717]_ ;
  assign \new_[4724]_  = \new_[4723]_  | \new_[4714]_ ;
  assign \new_[4725]_  = \new_[4724]_  | \new_[4707]_ ;
  assign \new_[4728]_  = \new_[1100]_  | \new_[1101]_ ;
  assign \new_[4731]_  = \new_[1098]_  | \new_[1099]_ ;
  assign \new_[4732]_  = \new_[4731]_  | \new_[4728]_ ;
  assign \new_[4735]_  = \new_[1096]_  | \new_[1097]_ ;
  assign \new_[4739]_  = \new_[1093]_  | \new_[1094]_ ;
  assign \new_[4740]_  = \new_[1095]_  | \new_[4739]_ ;
  assign \new_[4741]_  = \new_[4740]_  | \new_[4735]_ ;
  assign \new_[4742]_  = \new_[4741]_  | \new_[4732]_ ;
  assign \new_[4745]_  = \new_[1091]_  | \new_[1092]_ ;
  assign \new_[4748]_  = \new_[1089]_  | \new_[1090]_ ;
  assign \new_[4749]_  = \new_[4748]_  | \new_[4745]_ ;
  assign \new_[4752]_  = \new_[1087]_  | \new_[1088]_ ;
  assign \new_[4756]_  = \new_[1084]_  | \new_[1085]_ ;
  assign \new_[4757]_  = \new_[1086]_  | \new_[4756]_ ;
  assign \new_[4758]_  = \new_[4757]_  | \new_[4752]_ ;
  assign \new_[4759]_  = \new_[4758]_  | \new_[4749]_ ;
  assign \new_[4760]_  = \new_[4759]_  | \new_[4742]_ ;
  assign \new_[4761]_  = \new_[4760]_  | \new_[4725]_ ;
  assign \new_[4762]_  = \new_[4761]_  | \new_[4690]_ ;
  assign \new_[4765]_  = \new_[1082]_  | \new_[1083]_ ;
  assign \new_[4768]_  = \new_[1080]_  | \new_[1081]_ ;
  assign \new_[4769]_  = \new_[4768]_  | \new_[4765]_ ;
  assign \new_[4772]_  = \new_[1078]_  | \new_[1079]_ ;
  assign \new_[4776]_  = \new_[1075]_  | \new_[1076]_ ;
  assign \new_[4777]_  = \new_[1077]_  | \new_[4776]_ ;
  assign \new_[4778]_  = \new_[4777]_  | \new_[4772]_ ;
  assign \new_[4779]_  = \new_[4778]_  | \new_[4769]_ ;
  assign \new_[4782]_  = \new_[1073]_  | \new_[1074]_ ;
  assign \new_[4785]_  = \new_[1071]_  | \new_[1072]_ ;
  assign \new_[4786]_  = \new_[4785]_  | \new_[4782]_ ;
  assign \new_[4789]_  = \new_[1069]_  | \new_[1070]_ ;
  assign \new_[4793]_  = \new_[1066]_  | \new_[1067]_ ;
  assign \new_[4794]_  = \new_[1068]_  | \new_[4793]_ ;
  assign \new_[4795]_  = \new_[4794]_  | \new_[4789]_ ;
  assign \new_[4796]_  = \new_[4795]_  | \new_[4786]_ ;
  assign \new_[4797]_  = \new_[4796]_  | \new_[4779]_ ;
  assign \new_[4800]_  = \new_[1064]_  | \new_[1065]_ ;
  assign \new_[4803]_  = \new_[1062]_  | \new_[1063]_ ;
  assign \new_[4804]_  = \new_[4803]_  | \new_[4800]_ ;
  assign \new_[4807]_  = \new_[1060]_  | \new_[1061]_ ;
  assign \new_[4811]_  = \new_[1057]_  | \new_[1058]_ ;
  assign \new_[4812]_  = \new_[1059]_  | \new_[4811]_ ;
  assign \new_[4813]_  = \new_[4812]_  | \new_[4807]_ ;
  assign \new_[4814]_  = \new_[4813]_  | \new_[4804]_ ;
  assign \new_[4817]_  = \new_[1055]_  | \new_[1056]_ ;
  assign \new_[4820]_  = \new_[1053]_  | \new_[1054]_ ;
  assign \new_[4821]_  = \new_[4820]_  | \new_[4817]_ ;
  assign \new_[4824]_  = \new_[1051]_  | \new_[1052]_ ;
  assign \new_[4828]_  = \new_[1048]_  | \new_[1049]_ ;
  assign \new_[4829]_  = \new_[1050]_  | \new_[4828]_ ;
  assign \new_[4830]_  = \new_[4829]_  | \new_[4824]_ ;
  assign \new_[4831]_  = \new_[4830]_  | \new_[4821]_ ;
  assign \new_[4832]_  = \new_[4831]_  | \new_[4814]_ ;
  assign \new_[4833]_  = \new_[4832]_  | \new_[4797]_ ;
  assign \new_[4836]_  = \new_[1046]_  | \new_[1047]_ ;
  assign \new_[4839]_  = \new_[1044]_  | \new_[1045]_ ;
  assign \new_[4840]_  = \new_[4839]_  | \new_[4836]_ ;
  assign \new_[4843]_  = \new_[1042]_  | \new_[1043]_ ;
  assign \new_[4847]_  = \new_[1039]_  | \new_[1040]_ ;
  assign \new_[4848]_  = \new_[1041]_  | \new_[4847]_ ;
  assign \new_[4849]_  = \new_[4848]_  | \new_[4843]_ ;
  assign \new_[4850]_  = \new_[4849]_  | \new_[4840]_ ;
  assign \new_[4853]_  = \new_[1037]_  | \new_[1038]_ ;
  assign \new_[4856]_  = \new_[1035]_  | \new_[1036]_ ;
  assign \new_[4857]_  = \new_[4856]_  | \new_[4853]_ ;
  assign \new_[4860]_  = \new_[1033]_  | \new_[1034]_ ;
  assign \new_[4864]_  = \new_[1030]_  | \new_[1031]_ ;
  assign \new_[4865]_  = \new_[1032]_  | \new_[4864]_ ;
  assign \new_[4866]_  = \new_[4865]_  | \new_[4860]_ ;
  assign \new_[4867]_  = \new_[4866]_  | \new_[4857]_ ;
  assign \new_[4868]_  = \new_[4867]_  | \new_[4850]_ ;
  assign \new_[4871]_  = \new_[1028]_  | \new_[1029]_ ;
  assign \new_[4874]_  = \new_[1026]_  | \new_[1027]_ ;
  assign \new_[4875]_  = \new_[4874]_  | \new_[4871]_ ;
  assign \new_[4878]_  = \new_[1024]_  | \new_[1025]_ ;
  assign \new_[4882]_  = \new_[1021]_  | \new_[1022]_ ;
  assign \new_[4883]_  = \new_[1023]_  | \new_[4882]_ ;
  assign \new_[4884]_  = \new_[4883]_  | \new_[4878]_ ;
  assign \new_[4885]_  = \new_[4884]_  | \new_[4875]_ ;
  assign \new_[4888]_  = \new_[1019]_  | \new_[1020]_ ;
  assign \new_[4891]_  = \new_[1017]_  | \new_[1018]_ ;
  assign \new_[4892]_  = \new_[4891]_  | \new_[4888]_ ;
  assign \new_[4895]_  = \new_[1015]_  | \new_[1016]_ ;
  assign \new_[4899]_  = \new_[1012]_  | \new_[1013]_ ;
  assign \new_[4900]_  = \new_[1014]_  | \new_[4899]_ ;
  assign \new_[4901]_  = \new_[4900]_  | \new_[4895]_ ;
  assign \new_[4902]_  = \new_[4901]_  | \new_[4892]_ ;
  assign \new_[4903]_  = \new_[4902]_  | \new_[4885]_ ;
  assign \new_[4904]_  = \new_[4903]_  | \new_[4868]_ ;
  assign \new_[4905]_  = \new_[4904]_  | \new_[4833]_ ;
  assign \new_[4906]_  = \new_[4905]_  | \new_[4762]_ ;
  assign \new_[4909]_  = \new_[1010]_  | \new_[1011]_ ;
  assign \new_[4912]_  = \new_[1008]_  | \new_[1009]_ ;
  assign \new_[4913]_  = \new_[4912]_  | \new_[4909]_ ;
  assign \new_[4916]_  = \new_[1006]_  | \new_[1007]_ ;
  assign \new_[4920]_  = \new_[1003]_  | \new_[1004]_ ;
  assign \new_[4921]_  = \new_[1005]_  | \new_[4920]_ ;
  assign \new_[4922]_  = \new_[4921]_  | \new_[4916]_ ;
  assign \new_[4923]_  = \new_[4922]_  | \new_[4913]_ ;
  assign \new_[4926]_  = \new_[1001]_  | \new_[1002]_ ;
  assign \new_[4929]_  = \new_[999]_  | \new_[1000]_ ;
  assign \new_[4930]_  = \new_[4929]_  | \new_[4926]_ ;
  assign \new_[4933]_  = \new_[997]_  | \new_[998]_ ;
  assign \new_[4937]_  = \new_[994]_  | \new_[995]_ ;
  assign \new_[4938]_  = \new_[996]_  | \new_[4937]_ ;
  assign \new_[4939]_  = \new_[4938]_  | \new_[4933]_ ;
  assign \new_[4940]_  = \new_[4939]_  | \new_[4930]_ ;
  assign \new_[4941]_  = \new_[4940]_  | \new_[4923]_ ;
  assign \new_[4944]_  = \new_[992]_  | \new_[993]_ ;
  assign \new_[4947]_  = \new_[990]_  | \new_[991]_ ;
  assign \new_[4948]_  = \new_[4947]_  | \new_[4944]_ ;
  assign \new_[4951]_  = \new_[988]_  | \new_[989]_ ;
  assign \new_[4955]_  = \new_[985]_  | \new_[986]_ ;
  assign \new_[4956]_  = \new_[987]_  | \new_[4955]_ ;
  assign \new_[4957]_  = \new_[4956]_  | \new_[4951]_ ;
  assign \new_[4958]_  = \new_[4957]_  | \new_[4948]_ ;
  assign \new_[4961]_  = \new_[983]_  | \new_[984]_ ;
  assign \new_[4964]_  = \new_[981]_  | \new_[982]_ ;
  assign \new_[4965]_  = \new_[4964]_  | \new_[4961]_ ;
  assign \new_[4968]_  = \new_[979]_  | \new_[980]_ ;
  assign \new_[4972]_  = \new_[976]_  | \new_[977]_ ;
  assign \new_[4973]_  = \new_[978]_  | \new_[4972]_ ;
  assign \new_[4974]_  = \new_[4973]_  | \new_[4968]_ ;
  assign \new_[4975]_  = \new_[4974]_  | \new_[4965]_ ;
  assign \new_[4976]_  = \new_[4975]_  | \new_[4958]_ ;
  assign \new_[4977]_  = \new_[4976]_  | \new_[4941]_ ;
  assign \new_[4980]_  = \new_[974]_  | \new_[975]_ ;
  assign \new_[4983]_  = \new_[972]_  | \new_[973]_ ;
  assign \new_[4984]_  = \new_[4983]_  | \new_[4980]_ ;
  assign \new_[4987]_  = \new_[970]_  | \new_[971]_ ;
  assign \new_[4991]_  = \new_[967]_  | \new_[968]_ ;
  assign \new_[4992]_  = \new_[969]_  | \new_[4991]_ ;
  assign \new_[4993]_  = \new_[4992]_  | \new_[4987]_ ;
  assign \new_[4994]_  = \new_[4993]_  | \new_[4984]_ ;
  assign \new_[4997]_  = \new_[965]_  | \new_[966]_ ;
  assign \new_[5000]_  = \new_[963]_  | \new_[964]_ ;
  assign \new_[5001]_  = \new_[5000]_  | \new_[4997]_ ;
  assign \new_[5004]_  = \new_[961]_  | \new_[962]_ ;
  assign \new_[5008]_  = \new_[958]_  | \new_[959]_ ;
  assign \new_[5009]_  = \new_[960]_  | \new_[5008]_ ;
  assign \new_[5010]_  = \new_[5009]_  | \new_[5004]_ ;
  assign \new_[5011]_  = \new_[5010]_  | \new_[5001]_ ;
  assign \new_[5012]_  = \new_[5011]_  | \new_[4994]_ ;
  assign \new_[5015]_  = \new_[956]_  | \new_[957]_ ;
  assign \new_[5018]_  = \new_[954]_  | \new_[955]_ ;
  assign \new_[5019]_  = \new_[5018]_  | \new_[5015]_ ;
  assign \new_[5022]_  = \new_[952]_  | \new_[953]_ ;
  assign \new_[5026]_  = \new_[949]_  | \new_[950]_ ;
  assign \new_[5027]_  = \new_[951]_  | \new_[5026]_ ;
  assign \new_[5028]_  = \new_[5027]_  | \new_[5022]_ ;
  assign \new_[5029]_  = \new_[5028]_  | \new_[5019]_ ;
  assign \new_[5032]_  = \new_[947]_  | \new_[948]_ ;
  assign \new_[5035]_  = \new_[945]_  | \new_[946]_ ;
  assign \new_[5036]_  = \new_[5035]_  | \new_[5032]_ ;
  assign \new_[5039]_  = \new_[943]_  | \new_[944]_ ;
  assign \new_[5043]_  = \new_[940]_  | \new_[941]_ ;
  assign \new_[5044]_  = \new_[942]_  | \new_[5043]_ ;
  assign \new_[5045]_  = \new_[5044]_  | \new_[5039]_ ;
  assign \new_[5046]_  = \new_[5045]_  | \new_[5036]_ ;
  assign \new_[5047]_  = \new_[5046]_  | \new_[5029]_ ;
  assign \new_[5048]_  = \new_[5047]_  | \new_[5012]_ ;
  assign \new_[5049]_  = \new_[5048]_  | \new_[4977]_ ;
  assign \new_[5052]_  = \new_[938]_  | \new_[939]_ ;
  assign \new_[5055]_  = \new_[936]_  | \new_[937]_ ;
  assign \new_[5056]_  = \new_[5055]_  | \new_[5052]_ ;
  assign \new_[5059]_  = \new_[934]_  | \new_[935]_ ;
  assign \new_[5063]_  = \new_[931]_  | \new_[932]_ ;
  assign \new_[5064]_  = \new_[933]_  | \new_[5063]_ ;
  assign \new_[5065]_  = \new_[5064]_  | \new_[5059]_ ;
  assign \new_[5066]_  = \new_[5065]_  | \new_[5056]_ ;
  assign \new_[5069]_  = \new_[929]_  | \new_[930]_ ;
  assign \new_[5072]_  = \new_[927]_  | \new_[928]_ ;
  assign \new_[5073]_  = \new_[5072]_  | \new_[5069]_ ;
  assign \new_[5076]_  = \new_[925]_  | \new_[926]_ ;
  assign \new_[5080]_  = \new_[922]_  | \new_[923]_ ;
  assign \new_[5081]_  = \new_[924]_  | \new_[5080]_ ;
  assign \new_[5082]_  = \new_[5081]_  | \new_[5076]_ ;
  assign \new_[5083]_  = \new_[5082]_  | \new_[5073]_ ;
  assign \new_[5084]_  = \new_[5083]_  | \new_[5066]_ ;
  assign \new_[5087]_  = \new_[920]_  | \new_[921]_ ;
  assign \new_[5090]_  = \new_[918]_  | \new_[919]_ ;
  assign \new_[5091]_  = \new_[5090]_  | \new_[5087]_ ;
  assign \new_[5094]_  = \new_[916]_  | \new_[917]_ ;
  assign \new_[5098]_  = \new_[913]_  | \new_[914]_ ;
  assign \new_[5099]_  = \new_[915]_  | \new_[5098]_ ;
  assign \new_[5100]_  = \new_[5099]_  | \new_[5094]_ ;
  assign \new_[5101]_  = \new_[5100]_  | \new_[5091]_ ;
  assign \new_[5104]_  = \new_[911]_  | \new_[912]_ ;
  assign \new_[5107]_  = \new_[909]_  | \new_[910]_ ;
  assign \new_[5108]_  = \new_[5107]_  | \new_[5104]_ ;
  assign \new_[5111]_  = \new_[907]_  | \new_[908]_ ;
  assign \new_[5115]_  = \new_[904]_  | \new_[905]_ ;
  assign \new_[5116]_  = \new_[906]_  | \new_[5115]_ ;
  assign \new_[5117]_  = \new_[5116]_  | \new_[5111]_ ;
  assign \new_[5118]_  = \new_[5117]_  | \new_[5108]_ ;
  assign \new_[5119]_  = \new_[5118]_  | \new_[5101]_ ;
  assign \new_[5120]_  = \new_[5119]_  | \new_[5084]_ ;
  assign \new_[5123]_  = \new_[902]_  | \new_[903]_ ;
  assign \new_[5126]_  = \new_[900]_  | \new_[901]_ ;
  assign \new_[5127]_  = \new_[5126]_  | \new_[5123]_ ;
  assign \new_[5130]_  = \new_[898]_  | \new_[899]_ ;
  assign \new_[5134]_  = \new_[895]_  | \new_[896]_ ;
  assign \new_[5135]_  = \new_[897]_  | \new_[5134]_ ;
  assign \new_[5136]_  = \new_[5135]_  | \new_[5130]_ ;
  assign \new_[5137]_  = \new_[5136]_  | \new_[5127]_ ;
  assign \new_[5140]_  = \new_[893]_  | \new_[894]_ ;
  assign \new_[5143]_  = \new_[891]_  | \new_[892]_ ;
  assign \new_[5144]_  = \new_[5143]_  | \new_[5140]_ ;
  assign \new_[5147]_  = \new_[889]_  | \new_[890]_ ;
  assign \new_[5151]_  = \new_[886]_  | \new_[887]_ ;
  assign \new_[5152]_  = \new_[888]_  | \new_[5151]_ ;
  assign \new_[5153]_  = \new_[5152]_  | \new_[5147]_ ;
  assign \new_[5154]_  = \new_[5153]_  | \new_[5144]_ ;
  assign \new_[5155]_  = \new_[5154]_  | \new_[5137]_ ;
  assign \new_[5158]_  = \new_[884]_  | \new_[885]_ ;
  assign \new_[5161]_  = \new_[882]_  | \new_[883]_ ;
  assign \new_[5162]_  = \new_[5161]_  | \new_[5158]_ ;
  assign \new_[5165]_  = \new_[880]_  | \new_[881]_ ;
  assign \new_[5169]_  = \new_[877]_  | \new_[878]_ ;
  assign \new_[5170]_  = \new_[879]_  | \new_[5169]_ ;
  assign \new_[5171]_  = \new_[5170]_  | \new_[5165]_ ;
  assign \new_[5172]_  = \new_[5171]_  | \new_[5162]_ ;
  assign \new_[5175]_  = \new_[875]_  | \new_[876]_ ;
  assign \new_[5178]_  = \new_[873]_  | \new_[874]_ ;
  assign \new_[5179]_  = \new_[5178]_  | \new_[5175]_ ;
  assign \new_[5182]_  = \new_[871]_  | \new_[872]_ ;
  assign \new_[5186]_  = \new_[868]_  | \new_[869]_ ;
  assign \new_[5187]_  = \new_[870]_  | \new_[5186]_ ;
  assign \new_[5188]_  = \new_[5187]_  | \new_[5182]_ ;
  assign \new_[5189]_  = \new_[5188]_  | \new_[5179]_ ;
  assign \new_[5190]_  = \new_[5189]_  | \new_[5172]_ ;
  assign \new_[5191]_  = \new_[5190]_  | \new_[5155]_ ;
  assign \new_[5192]_  = \new_[5191]_  | \new_[5120]_ ;
  assign \new_[5193]_  = \new_[5192]_  | \new_[5049]_ ;
  assign \new_[5194]_  = \new_[5193]_  | \new_[4906]_ ;
  assign \new_[5197]_  = \new_[866]_  | \new_[867]_ ;
  assign \new_[5200]_  = \new_[864]_  | \new_[865]_ ;
  assign \new_[5201]_  = \new_[5200]_  | \new_[5197]_ ;
  assign \new_[5204]_  = \new_[862]_  | \new_[863]_ ;
  assign \new_[5208]_  = \new_[859]_  | \new_[860]_ ;
  assign \new_[5209]_  = \new_[861]_  | \new_[5208]_ ;
  assign \new_[5210]_  = \new_[5209]_  | \new_[5204]_ ;
  assign \new_[5211]_  = \new_[5210]_  | \new_[5201]_ ;
  assign \new_[5214]_  = \new_[857]_  | \new_[858]_ ;
  assign \new_[5217]_  = \new_[855]_  | \new_[856]_ ;
  assign \new_[5218]_  = \new_[5217]_  | \new_[5214]_ ;
  assign \new_[5221]_  = \new_[853]_  | \new_[854]_ ;
  assign \new_[5225]_  = \new_[850]_  | \new_[851]_ ;
  assign \new_[5226]_  = \new_[852]_  | \new_[5225]_ ;
  assign \new_[5227]_  = \new_[5226]_  | \new_[5221]_ ;
  assign \new_[5228]_  = \new_[5227]_  | \new_[5218]_ ;
  assign \new_[5229]_  = \new_[5228]_  | \new_[5211]_ ;
  assign \new_[5232]_  = \new_[848]_  | \new_[849]_ ;
  assign \new_[5235]_  = \new_[846]_  | \new_[847]_ ;
  assign \new_[5236]_  = \new_[5235]_  | \new_[5232]_ ;
  assign \new_[5239]_  = \new_[844]_  | \new_[845]_ ;
  assign \new_[5243]_  = \new_[841]_  | \new_[842]_ ;
  assign \new_[5244]_  = \new_[843]_  | \new_[5243]_ ;
  assign \new_[5245]_  = \new_[5244]_  | \new_[5239]_ ;
  assign \new_[5246]_  = \new_[5245]_  | \new_[5236]_ ;
  assign \new_[5249]_  = \new_[839]_  | \new_[840]_ ;
  assign \new_[5252]_  = \new_[837]_  | \new_[838]_ ;
  assign \new_[5253]_  = \new_[5252]_  | \new_[5249]_ ;
  assign \new_[5256]_  = \new_[835]_  | \new_[836]_ ;
  assign \new_[5260]_  = \new_[832]_  | \new_[833]_ ;
  assign \new_[5261]_  = \new_[834]_  | \new_[5260]_ ;
  assign \new_[5262]_  = \new_[5261]_  | \new_[5256]_ ;
  assign \new_[5263]_  = \new_[5262]_  | \new_[5253]_ ;
  assign \new_[5264]_  = \new_[5263]_  | \new_[5246]_ ;
  assign \new_[5265]_  = \new_[5264]_  | \new_[5229]_ ;
  assign \new_[5268]_  = \new_[830]_  | \new_[831]_ ;
  assign \new_[5271]_  = \new_[828]_  | \new_[829]_ ;
  assign \new_[5272]_  = \new_[5271]_  | \new_[5268]_ ;
  assign \new_[5275]_  = \new_[826]_  | \new_[827]_ ;
  assign \new_[5279]_  = \new_[823]_  | \new_[824]_ ;
  assign \new_[5280]_  = \new_[825]_  | \new_[5279]_ ;
  assign \new_[5281]_  = \new_[5280]_  | \new_[5275]_ ;
  assign \new_[5282]_  = \new_[5281]_  | \new_[5272]_ ;
  assign \new_[5285]_  = \new_[821]_  | \new_[822]_ ;
  assign \new_[5288]_  = \new_[819]_  | \new_[820]_ ;
  assign \new_[5289]_  = \new_[5288]_  | \new_[5285]_ ;
  assign \new_[5292]_  = \new_[817]_  | \new_[818]_ ;
  assign \new_[5296]_  = \new_[814]_  | \new_[815]_ ;
  assign \new_[5297]_  = \new_[816]_  | \new_[5296]_ ;
  assign \new_[5298]_  = \new_[5297]_  | \new_[5292]_ ;
  assign \new_[5299]_  = \new_[5298]_  | \new_[5289]_ ;
  assign \new_[5300]_  = \new_[5299]_  | \new_[5282]_ ;
  assign \new_[5303]_  = \new_[812]_  | \new_[813]_ ;
  assign \new_[5306]_  = \new_[810]_  | \new_[811]_ ;
  assign \new_[5307]_  = \new_[5306]_  | \new_[5303]_ ;
  assign \new_[5310]_  = \new_[808]_  | \new_[809]_ ;
  assign \new_[5314]_  = \new_[805]_  | \new_[806]_ ;
  assign \new_[5315]_  = \new_[807]_  | \new_[5314]_ ;
  assign \new_[5316]_  = \new_[5315]_  | \new_[5310]_ ;
  assign \new_[5317]_  = \new_[5316]_  | \new_[5307]_ ;
  assign \new_[5320]_  = \new_[803]_  | \new_[804]_ ;
  assign \new_[5323]_  = \new_[801]_  | \new_[802]_ ;
  assign \new_[5324]_  = \new_[5323]_  | \new_[5320]_ ;
  assign \new_[5327]_  = \new_[799]_  | \new_[800]_ ;
  assign \new_[5331]_  = \new_[796]_  | \new_[797]_ ;
  assign \new_[5332]_  = \new_[798]_  | \new_[5331]_ ;
  assign \new_[5333]_  = \new_[5332]_  | \new_[5327]_ ;
  assign \new_[5334]_  = \new_[5333]_  | \new_[5324]_ ;
  assign \new_[5335]_  = \new_[5334]_  | \new_[5317]_ ;
  assign \new_[5336]_  = \new_[5335]_  | \new_[5300]_ ;
  assign \new_[5337]_  = \new_[5336]_  | \new_[5265]_ ;
  assign \new_[5340]_  = \new_[794]_  | \new_[795]_ ;
  assign \new_[5343]_  = \new_[792]_  | \new_[793]_ ;
  assign \new_[5344]_  = \new_[5343]_  | \new_[5340]_ ;
  assign \new_[5347]_  = \new_[790]_  | \new_[791]_ ;
  assign \new_[5351]_  = \new_[787]_  | \new_[788]_ ;
  assign \new_[5352]_  = \new_[789]_  | \new_[5351]_ ;
  assign \new_[5353]_  = \new_[5352]_  | \new_[5347]_ ;
  assign \new_[5354]_  = \new_[5353]_  | \new_[5344]_ ;
  assign \new_[5357]_  = \new_[785]_  | \new_[786]_ ;
  assign \new_[5360]_  = \new_[783]_  | \new_[784]_ ;
  assign \new_[5361]_  = \new_[5360]_  | \new_[5357]_ ;
  assign \new_[5364]_  = \new_[781]_  | \new_[782]_ ;
  assign \new_[5368]_  = \new_[778]_  | \new_[779]_ ;
  assign \new_[5369]_  = \new_[780]_  | \new_[5368]_ ;
  assign \new_[5370]_  = \new_[5369]_  | \new_[5364]_ ;
  assign \new_[5371]_  = \new_[5370]_  | \new_[5361]_ ;
  assign \new_[5372]_  = \new_[5371]_  | \new_[5354]_ ;
  assign \new_[5375]_  = \new_[776]_  | \new_[777]_ ;
  assign \new_[5378]_  = \new_[774]_  | \new_[775]_ ;
  assign \new_[5379]_  = \new_[5378]_  | \new_[5375]_ ;
  assign \new_[5382]_  = \new_[772]_  | \new_[773]_ ;
  assign \new_[5386]_  = \new_[769]_  | \new_[770]_ ;
  assign \new_[5387]_  = \new_[771]_  | \new_[5386]_ ;
  assign \new_[5388]_  = \new_[5387]_  | \new_[5382]_ ;
  assign \new_[5389]_  = \new_[5388]_  | \new_[5379]_ ;
  assign \new_[5392]_  = \new_[767]_  | \new_[768]_ ;
  assign \new_[5395]_  = \new_[765]_  | \new_[766]_ ;
  assign \new_[5396]_  = \new_[5395]_  | \new_[5392]_ ;
  assign \new_[5399]_  = \new_[763]_  | \new_[764]_ ;
  assign \new_[5403]_  = \new_[760]_  | \new_[761]_ ;
  assign \new_[5404]_  = \new_[762]_  | \new_[5403]_ ;
  assign \new_[5405]_  = \new_[5404]_  | \new_[5399]_ ;
  assign \new_[5406]_  = \new_[5405]_  | \new_[5396]_ ;
  assign \new_[5407]_  = \new_[5406]_  | \new_[5389]_ ;
  assign \new_[5408]_  = \new_[5407]_  | \new_[5372]_ ;
  assign \new_[5411]_  = \new_[758]_  | \new_[759]_ ;
  assign \new_[5414]_  = \new_[756]_  | \new_[757]_ ;
  assign \new_[5415]_  = \new_[5414]_  | \new_[5411]_ ;
  assign \new_[5418]_  = \new_[754]_  | \new_[755]_ ;
  assign \new_[5422]_  = \new_[751]_  | \new_[752]_ ;
  assign \new_[5423]_  = \new_[753]_  | \new_[5422]_ ;
  assign \new_[5424]_  = \new_[5423]_  | \new_[5418]_ ;
  assign \new_[5425]_  = \new_[5424]_  | \new_[5415]_ ;
  assign \new_[5428]_  = \new_[749]_  | \new_[750]_ ;
  assign \new_[5431]_  = \new_[747]_  | \new_[748]_ ;
  assign \new_[5432]_  = \new_[5431]_  | \new_[5428]_ ;
  assign \new_[5435]_  = \new_[745]_  | \new_[746]_ ;
  assign \new_[5439]_  = \new_[742]_  | \new_[743]_ ;
  assign \new_[5440]_  = \new_[744]_  | \new_[5439]_ ;
  assign \new_[5441]_  = \new_[5440]_  | \new_[5435]_ ;
  assign \new_[5442]_  = \new_[5441]_  | \new_[5432]_ ;
  assign \new_[5443]_  = \new_[5442]_  | \new_[5425]_ ;
  assign \new_[5446]_  = \new_[740]_  | \new_[741]_ ;
  assign \new_[5449]_  = \new_[738]_  | \new_[739]_ ;
  assign \new_[5450]_  = \new_[5449]_  | \new_[5446]_ ;
  assign \new_[5453]_  = \new_[736]_  | \new_[737]_ ;
  assign \new_[5457]_  = \new_[733]_  | \new_[734]_ ;
  assign \new_[5458]_  = \new_[735]_  | \new_[5457]_ ;
  assign \new_[5459]_  = \new_[5458]_  | \new_[5453]_ ;
  assign \new_[5460]_  = \new_[5459]_  | \new_[5450]_ ;
  assign \new_[5463]_  = \new_[731]_  | \new_[732]_ ;
  assign \new_[5466]_  = \new_[729]_  | \new_[730]_ ;
  assign \new_[5467]_  = \new_[5466]_  | \new_[5463]_ ;
  assign \new_[5470]_  = \new_[727]_  | \new_[728]_ ;
  assign \new_[5474]_  = \new_[724]_  | \new_[725]_ ;
  assign \new_[5475]_  = \new_[726]_  | \new_[5474]_ ;
  assign \new_[5476]_  = \new_[5475]_  | \new_[5470]_ ;
  assign \new_[5477]_  = \new_[5476]_  | \new_[5467]_ ;
  assign \new_[5478]_  = \new_[5477]_  | \new_[5460]_ ;
  assign \new_[5479]_  = \new_[5478]_  | \new_[5443]_ ;
  assign \new_[5480]_  = \new_[5479]_  | \new_[5408]_ ;
  assign \new_[5481]_  = \new_[5480]_  | \new_[5337]_ ;
  assign \new_[5484]_  = \new_[722]_  | \new_[723]_ ;
  assign \new_[5487]_  = \new_[720]_  | \new_[721]_ ;
  assign \new_[5488]_  = \new_[5487]_  | \new_[5484]_ ;
  assign \new_[5491]_  = \new_[718]_  | \new_[719]_ ;
  assign \new_[5495]_  = \new_[715]_  | \new_[716]_ ;
  assign \new_[5496]_  = \new_[717]_  | \new_[5495]_ ;
  assign \new_[5497]_  = \new_[5496]_  | \new_[5491]_ ;
  assign \new_[5498]_  = \new_[5497]_  | \new_[5488]_ ;
  assign \new_[5501]_  = \new_[713]_  | \new_[714]_ ;
  assign \new_[5504]_  = \new_[711]_  | \new_[712]_ ;
  assign \new_[5505]_  = \new_[5504]_  | \new_[5501]_ ;
  assign \new_[5508]_  = \new_[709]_  | \new_[710]_ ;
  assign \new_[5512]_  = \new_[706]_  | \new_[707]_ ;
  assign \new_[5513]_  = \new_[708]_  | \new_[5512]_ ;
  assign \new_[5514]_  = \new_[5513]_  | \new_[5508]_ ;
  assign \new_[5515]_  = \new_[5514]_  | \new_[5505]_ ;
  assign \new_[5516]_  = \new_[5515]_  | \new_[5498]_ ;
  assign \new_[5519]_  = \new_[704]_  | \new_[705]_ ;
  assign \new_[5522]_  = \new_[702]_  | \new_[703]_ ;
  assign \new_[5523]_  = \new_[5522]_  | \new_[5519]_ ;
  assign \new_[5526]_  = \new_[700]_  | \new_[701]_ ;
  assign \new_[5530]_  = \new_[697]_  | \new_[698]_ ;
  assign \new_[5531]_  = \new_[699]_  | \new_[5530]_ ;
  assign \new_[5532]_  = \new_[5531]_  | \new_[5526]_ ;
  assign \new_[5533]_  = \new_[5532]_  | \new_[5523]_ ;
  assign \new_[5536]_  = \new_[695]_  | \new_[696]_ ;
  assign \new_[5539]_  = \new_[693]_  | \new_[694]_ ;
  assign \new_[5540]_  = \new_[5539]_  | \new_[5536]_ ;
  assign \new_[5543]_  = \new_[691]_  | \new_[692]_ ;
  assign \new_[5547]_  = \new_[688]_  | \new_[689]_ ;
  assign \new_[5548]_  = \new_[690]_  | \new_[5547]_ ;
  assign \new_[5549]_  = \new_[5548]_  | \new_[5543]_ ;
  assign \new_[5550]_  = \new_[5549]_  | \new_[5540]_ ;
  assign \new_[5551]_  = \new_[5550]_  | \new_[5533]_ ;
  assign \new_[5552]_  = \new_[5551]_  | \new_[5516]_ ;
  assign \new_[5555]_  = \new_[686]_  | \new_[687]_ ;
  assign \new_[5558]_  = \new_[684]_  | \new_[685]_ ;
  assign \new_[5559]_  = \new_[5558]_  | \new_[5555]_ ;
  assign \new_[5562]_  = \new_[682]_  | \new_[683]_ ;
  assign \new_[5566]_  = \new_[679]_  | \new_[680]_ ;
  assign \new_[5567]_  = \new_[681]_  | \new_[5566]_ ;
  assign \new_[5568]_  = \new_[5567]_  | \new_[5562]_ ;
  assign \new_[5569]_  = \new_[5568]_  | \new_[5559]_ ;
  assign \new_[5572]_  = \new_[677]_  | \new_[678]_ ;
  assign \new_[5575]_  = \new_[675]_  | \new_[676]_ ;
  assign \new_[5576]_  = \new_[5575]_  | \new_[5572]_ ;
  assign \new_[5579]_  = \new_[673]_  | \new_[674]_ ;
  assign \new_[5583]_  = \new_[670]_  | \new_[671]_ ;
  assign \new_[5584]_  = \new_[672]_  | \new_[5583]_ ;
  assign \new_[5585]_  = \new_[5584]_  | \new_[5579]_ ;
  assign \new_[5586]_  = \new_[5585]_  | \new_[5576]_ ;
  assign \new_[5587]_  = \new_[5586]_  | \new_[5569]_ ;
  assign \new_[5590]_  = \new_[668]_  | \new_[669]_ ;
  assign \new_[5593]_  = \new_[666]_  | \new_[667]_ ;
  assign \new_[5594]_  = \new_[5593]_  | \new_[5590]_ ;
  assign \new_[5597]_  = \new_[664]_  | \new_[665]_ ;
  assign \new_[5601]_  = \new_[661]_  | \new_[662]_ ;
  assign \new_[5602]_  = \new_[663]_  | \new_[5601]_ ;
  assign \new_[5603]_  = \new_[5602]_  | \new_[5597]_ ;
  assign \new_[5604]_  = \new_[5603]_  | \new_[5594]_ ;
  assign \new_[5607]_  = \new_[659]_  | \new_[660]_ ;
  assign \new_[5610]_  = \new_[657]_  | \new_[658]_ ;
  assign \new_[5611]_  = \new_[5610]_  | \new_[5607]_ ;
  assign \new_[5614]_  = \new_[655]_  | \new_[656]_ ;
  assign \new_[5618]_  = \new_[652]_  | \new_[653]_ ;
  assign \new_[5619]_  = \new_[654]_  | \new_[5618]_ ;
  assign \new_[5620]_  = \new_[5619]_  | \new_[5614]_ ;
  assign \new_[5621]_  = \new_[5620]_  | \new_[5611]_ ;
  assign \new_[5622]_  = \new_[5621]_  | \new_[5604]_ ;
  assign \new_[5623]_  = \new_[5622]_  | \new_[5587]_ ;
  assign \new_[5624]_  = \new_[5623]_  | \new_[5552]_ ;
  assign \new_[5627]_  = \new_[650]_  | \new_[651]_ ;
  assign \new_[5630]_  = \new_[648]_  | \new_[649]_ ;
  assign \new_[5631]_  = \new_[5630]_  | \new_[5627]_ ;
  assign \new_[5634]_  = \new_[646]_  | \new_[647]_ ;
  assign \new_[5638]_  = \new_[643]_  | \new_[644]_ ;
  assign \new_[5639]_  = \new_[645]_  | \new_[5638]_ ;
  assign \new_[5640]_  = \new_[5639]_  | \new_[5634]_ ;
  assign \new_[5641]_  = \new_[5640]_  | \new_[5631]_ ;
  assign \new_[5644]_  = \new_[641]_  | \new_[642]_ ;
  assign \new_[5647]_  = \new_[639]_  | \new_[640]_ ;
  assign \new_[5648]_  = \new_[5647]_  | \new_[5644]_ ;
  assign \new_[5651]_  = \new_[637]_  | \new_[638]_ ;
  assign \new_[5655]_  = \new_[634]_  | \new_[635]_ ;
  assign \new_[5656]_  = \new_[636]_  | \new_[5655]_ ;
  assign \new_[5657]_  = \new_[5656]_  | \new_[5651]_ ;
  assign \new_[5658]_  = \new_[5657]_  | \new_[5648]_ ;
  assign \new_[5659]_  = \new_[5658]_  | \new_[5641]_ ;
  assign \new_[5662]_  = \new_[632]_  | \new_[633]_ ;
  assign \new_[5665]_  = \new_[630]_  | \new_[631]_ ;
  assign \new_[5666]_  = \new_[5665]_  | \new_[5662]_ ;
  assign \new_[5669]_  = \new_[628]_  | \new_[629]_ ;
  assign \new_[5673]_  = \new_[625]_  | \new_[626]_ ;
  assign \new_[5674]_  = \new_[627]_  | \new_[5673]_ ;
  assign \new_[5675]_  = \new_[5674]_  | \new_[5669]_ ;
  assign \new_[5676]_  = \new_[5675]_  | \new_[5666]_ ;
  assign \new_[5679]_  = \new_[623]_  | \new_[624]_ ;
  assign \new_[5682]_  = \new_[621]_  | \new_[622]_ ;
  assign \new_[5683]_  = \new_[5682]_  | \new_[5679]_ ;
  assign \new_[5686]_  = \new_[619]_  | \new_[620]_ ;
  assign \new_[5690]_  = \new_[616]_  | \new_[617]_ ;
  assign \new_[5691]_  = \new_[618]_  | \new_[5690]_ ;
  assign \new_[5692]_  = \new_[5691]_  | \new_[5686]_ ;
  assign \new_[5693]_  = \new_[5692]_  | \new_[5683]_ ;
  assign \new_[5694]_  = \new_[5693]_  | \new_[5676]_ ;
  assign \new_[5695]_  = \new_[5694]_  | \new_[5659]_ ;
  assign \new_[5698]_  = \new_[614]_  | \new_[615]_ ;
  assign \new_[5701]_  = \new_[612]_  | \new_[613]_ ;
  assign \new_[5702]_  = \new_[5701]_  | \new_[5698]_ ;
  assign \new_[5705]_  = \new_[610]_  | \new_[611]_ ;
  assign \new_[5709]_  = \new_[607]_  | \new_[608]_ ;
  assign \new_[5710]_  = \new_[609]_  | \new_[5709]_ ;
  assign \new_[5711]_  = \new_[5710]_  | \new_[5705]_ ;
  assign \new_[5712]_  = \new_[5711]_  | \new_[5702]_ ;
  assign \new_[5715]_  = \new_[605]_  | \new_[606]_ ;
  assign \new_[5718]_  = \new_[603]_  | \new_[604]_ ;
  assign \new_[5719]_  = \new_[5718]_  | \new_[5715]_ ;
  assign \new_[5722]_  = \new_[601]_  | \new_[602]_ ;
  assign \new_[5726]_  = \new_[598]_  | \new_[599]_ ;
  assign \new_[5727]_  = \new_[600]_  | \new_[5726]_ ;
  assign \new_[5728]_  = \new_[5727]_  | \new_[5722]_ ;
  assign \new_[5729]_  = \new_[5728]_  | \new_[5719]_ ;
  assign \new_[5730]_  = \new_[5729]_  | \new_[5712]_ ;
  assign \new_[5733]_  = \new_[596]_  | \new_[597]_ ;
  assign \new_[5736]_  = \new_[594]_  | \new_[595]_ ;
  assign \new_[5737]_  = \new_[5736]_  | \new_[5733]_ ;
  assign \new_[5740]_  = \new_[592]_  | \new_[593]_ ;
  assign \new_[5744]_  = \new_[589]_  | \new_[590]_ ;
  assign \new_[5745]_  = \new_[591]_  | \new_[5744]_ ;
  assign \new_[5746]_  = \new_[5745]_  | \new_[5740]_ ;
  assign \new_[5747]_  = \new_[5746]_  | \new_[5737]_ ;
  assign \new_[5750]_  = \new_[587]_  | \new_[588]_ ;
  assign \new_[5754]_  = \new_[584]_  | \new_[585]_ ;
  assign \new_[5755]_  = \new_[586]_  | \new_[5754]_ ;
  assign \new_[5756]_  = \new_[5755]_  | \new_[5750]_ ;
  assign \new_[5759]_  = \new_[582]_  | \new_[583]_ ;
  assign \new_[5763]_  = \new_[579]_  | \new_[580]_ ;
  assign \new_[5764]_  = \new_[581]_  | \new_[5763]_ ;
  assign \new_[5765]_  = \new_[5764]_  | \new_[5759]_ ;
  assign \new_[5766]_  = \new_[5765]_  | \new_[5756]_ ;
  assign \new_[5767]_  = \new_[5766]_  | \new_[5747]_ ;
  assign \new_[5768]_  = \new_[5767]_  | \new_[5730]_ ;
  assign \new_[5769]_  = \new_[5768]_  | \new_[5695]_ ;
  assign \new_[5770]_  = \new_[5769]_  | \new_[5624]_ ;
  assign \new_[5771]_  = \new_[5770]_  | \new_[5481]_ ;
  assign \new_[5772]_  = \new_[5771]_  | \new_[5194]_ ;
  assign \new_[5775]_  = \new_[577]_  | \new_[578]_ ;
  assign \new_[5778]_  = \new_[575]_  | \new_[576]_ ;
  assign \new_[5779]_  = \new_[5778]_  | \new_[5775]_ ;
  assign \new_[5782]_  = \new_[573]_  | \new_[574]_ ;
  assign \new_[5786]_  = \new_[570]_  | \new_[571]_ ;
  assign \new_[5787]_  = \new_[572]_  | \new_[5786]_ ;
  assign \new_[5788]_  = \new_[5787]_  | \new_[5782]_ ;
  assign \new_[5789]_  = \new_[5788]_  | \new_[5779]_ ;
  assign \new_[5792]_  = \new_[568]_  | \new_[569]_ ;
  assign \new_[5795]_  = \new_[566]_  | \new_[567]_ ;
  assign \new_[5796]_  = \new_[5795]_  | \new_[5792]_ ;
  assign \new_[5799]_  = \new_[564]_  | \new_[565]_ ;
  assign \new_[5803]_  = \new_[561]_  | \new_[562]_ ;
  assign \new_[5804]_  = \new_[563]_  | \new_[5803]_ ;
  assign \new_[5805]_  = \new_[5804]_  | \new_[5799]_ ;
  assign \new_[5806]_  = \new_[5805]_  | \new_[5796]_ ;
  assign \new_[5807]_  = \new_[5806]_  | \new_[5789]_ ;
  assign \new_[5810]_  = \new_[559]_  | \new_[560]_ ;
  assign \new_[5813]_  = \new_[557]_  | \new_[558]_ ;
  assign \new_[5814]_  = \new_[5813]_  | \new_[5810]_ ;
  assign \new_[5817]_  = \new_[555]_  | \new_[556]_ ;
  assign \new_[5821]_  = \new_[552]_  | \new_[553]_ ;
  assign \new_[5822]_  = \new_[554]_  | \new_[5821]_ ;
  assign \new_[5823]_  = \new_[5822]_  | \new_[5817]_ ;
  assign \new_[5824]_  = \new_[5823]_  | \new_[5814]_ ;
  assign \new_[5827]_  = \new_[550]_  | \new_[551]_ ;
  assign \new_[5830]_  = \new_[548]_  | \new_[549]_ ;
  assign \new_[5831]_  = \new_[5830]_  | \new_[5827]_ ;
  assign \new_[5834]_  = \new_[546]_  | \new_[547]_ ;
  assign \new_[5838]_  = \new_[543]_  | \new_[544]_ ;
  assign \new_[5839]_  = \new_[545]_  | \new_[5838]_ ;
  assign \new_[5840]_  = \new_[5839]_  | \new_[5834]_ ;
  assign \new_[5841]_  = \new_[5840]_  | \new_[5831]_ ;
  assign \new_[5842]_  = \new_[5841]_  | \new_[5824]_ ;
  assign \new_[5843]_  = \new_[5842]_  | \new_[5807]_ ;
  assign \new_[5846]_  = \new_[541]_  | \new_[542]_ ;
  assign \new_[5849]_  = \new_[539]_  | \new_[540]_ ;
  assign \new_[5850]_  = \new_[5849]_  | \new_[5846]_ ;
  assign \new_[5853]_  = \new_[537]_  | \new_[538]_ ;
  assign \new_[5857]_  = \new_[534]_  | \new_[535]_ ;
  assign \new_[5858]_  = \new_[536]_  | \new_[5857]_ ;
  assign \new_[5859]_  = \new_[5858]_  | \new_[5853]_ ;
  assign \new_[5860]_  = \new_[5859]_  | \new_[5850]_ ;
  assign \new_[5863]_  = \new_[532]_  | \new_[533]_ ;
  assign \new_[5866]_  = \new_[530]_  | \new_[531]_ ;
  assign \new_[5867]_  = \new_[5866]_  | \new_[5863]_ ;
  assign \new_[5870]_  = \new_[528]_  | \new_[529]_ ;
  assign \new_[5874]_  = \new_[525]_  | \new_[526]_ ;
  assign \new_[5875]_  = \new_[527]_  | \new_[5874]_ ;
  assign \new_[5876]_  = \new_[5875]_  | \new_[5870]_ ;
  assign \new_[5877]_  = \new_[5876]_  | \new_[5867]_ ;
  assign \new_[5878]_  = \new_[5877]_  | \new_[5860]_ ;
  assign \new_[5881]_  = \new_[523]_  | \new_[524]_ ;
  assign \new_[5884]_  = \new_[521]_  | \new_[522]_ ;
  assign \new_[5885]_  = \new_[5884]_  | \new_[5881]_ ;
  assign \new_[5888]_  = \new_[519]_  | \new_[520]_ ;
  assign \new_[5892]_  = \new_[516]_  | \new_[517]_ ;
  assign \new_[5893]_  = \new_[518]_  | \new_[5892]_ ;
  assign \new_[5894]_  = \new_[5893]_  | \new_[5888]_ ;
  assign \new_[5895]_  = \new_[5894]_  | \new_[5885]_ ;
  assign \new_[5898]_  = \new_[514]_  | \new_[515]_ ;
  assign \new_[5901]_  = \new_[512]_  | \new_[513]_ ;
  assign \new_[5902]_  = \new_[5901]_  | \new_[5898]_ ;
  assign \new_[5905]_  = \new_[510]_  | \new_[511]_ ;
  assign \new_[5909]_  = \new_[507]_  | \new_[508]_ ;
  assign \new_[5910]_  = \new_[509]_  | \new_[5909]_ ;
  assign \new_[5911]_  = \new_[5910]_  | \new_[5905]_ ;
  assign \new_[5912]_  = \new_[5911]_  | \new_[5902]_ ;
  assign \new_[5913]_  = \new_[5912]_  | \new_[5895]_ ;
  assign \new_[5914]_  = \new_[5913]_  | \new_[5878]_ ;
  assign \new_[5915]_  = \new_[5914]_  | \new_[5843]_ ;
  assign \new_[5918]_  = \new_[505]_  | \new_[506]_ ;
  assign \new_[5921]_  = \new_[503]_  | \new_[504]_ ;
  assign \new_[5922]_  = \new_[5921]_  | \new_[5918]_ ;
  assign \new_[5925]_  = \new_[501]_  | \new_[502]_ ;
  assign \new_[5929]_  = \new_[498]_  | \new_[499]_ ;
  assign \new_[5930]_  = \new_[500]_  | \new_[5929]_ ;
  assign \new_[5931]_  = \new_[5930]_  | \new_[5925]_ ;
  assign \new_[5932]_  = \new_[5931]_  | \new_[5922]_ ;
  assign \new_[5935]_  = \new_[496]_  | \new_[497]_ ;
  assign \new_[5938]_  = \new_[494]_  | \new_[495]_ ;
  assign \new_[5939]_  = \new_[5938]_  | \new_[5935]_ ;
  assign \new_[5942]_  = \new_[492]_  | \new_[493]_ ;
  assign \new_[5946]_  = \new_[489]_  | \new_[490]_ ;
  assign \new_[5947]_  = \new_[491]_  | \new_[5946]_ ;
  assign \new_[5948]_  = \new_[5947]_  | \new_[5942]_ ;
  assign \new_[5949]_  = \new_[5948]_  | \new_[5939]_ ;
  assign \new_[5950]_  = \new_[5949]_  | \new_[5932]_ ;
  assign \new_[5953]_  = \new_[487]_  | \new_[488]_ ;
  assign \new_[5956]_  = \new_[485]_  | \new_[486]_ ;
  assign \new_[5957]_  = \new_[5956]_  | \new_[5953]_ ;
  assign \new_[5960]_  = \new_[483]_  | \new_[484]_ ;
  assign \new_[5964]_  = \new_[480]_  | \new_[481]_ ;
  assign \new_[5965]_  = \new_[482]_  | \new_[5964]_ ;
  assign \new_[5966]_  = \new_[5965]_  | \new_[5960]_ ;
  assign \new_[5967]_  = \new_[5966]_  | \new_[5957]_ ;
  assign \new_[5970]_  = \new_[478]_  | \new_[479]_ ;
  assign \new_[5973]_  = \new_[476]_  | \new_[477]_ ;
  assign \new_[5974]_  = \new_[5973]_  | \new_[5970]_ ;
  assign \new_[5977]_  = \new_[474]_  | \new_[475]_ ;
  assign \new_[5981]_  = \new_[471]_  | \new_[472]_ ;
  assign \new_[5982]_  = \new_[473]_  | \new_[5981]_ ;
  assign \new_[5983]_  = \new_[5982]_  | \new_[5977]_ ;
  assign \new_[5984]_  = \new_[5983]_  | \new_[5974]_ ;
  assign \new_[5985]_  = \new_[5984]_  | \new_[5967]_ ;
  assign \new_[5986]_  = \new_[5985]_  | \new_[5950]_ ;
  assign \new_[5989]_  = \new_[469]_  | \new_[470]_ ;
  assign \new_[5992]_  = \new_[467]_  | \new_[468]_ ;
  assign \new_[5993]_  = \new_[5992]_  | \new_[5989]_ ;
  assign \new_[5996]_  = \new_[465]_  | \new_[466]_ ;
  assign \new_[6000]_  = \new_[462]_  | \new_[463]_ ;
  assign \new_[6001]_  = \new_[464]_  | \new_[6000]_ ;
  assign \new_[6002]_  = \new_[6001]_  | \new_[5996]_ ;
  assign \new_[6003]_  = \new_[6002]_  | \new_[5993]_ ;
  assign \new_[6006]_  = \new_[460]_  | \new_[461]_ ;
  assign \new_[6009]_  = \new_[458]_  | \new_[459]_ ;
  assign \new_[6010]_  = \new_[6009]_  | \new_[6006]_ ;
  assign \new_[6013]_  = \new_[456]_  | \new_[457]_ ;
  assign \new_[6017]_  = \new_[453]_  | \new_[454]_ ;
  assign \new_[6018]_  = \new_[455]_  | \new_[6017]_ ;
  assign \new_[6019]_  = \new_[6018]_  | \new_[6013]_ ;
  assign \new_[6020]_  = \new_[6019]_  | \new_[6010]_ ;
  assign \new_[6021]_  = \new_[6020]_  | \new_[6003]_ ;
  assign \new_[6024]_  = \new_[451]_  | \new_[452]_ ;
  assign \new_[6027]_  = \new_[449]_  | \new_[450]_ ;
  assign \new_[6028]_  = \new_[6027]_  | \new_[6024]_ ;
  assign \new_[6031]_  = \new_[447]_  | \new_[448]_ ;
  assign \new_[6035]_  = \new_[444]_  | \new_[445]_ ;
  assign \new_[6036]_  = \new_[446]_  | \new_[6035]_ ;
  assign \new_[6037]_  = \new_[6036]_  | \new_[6031]_ ;
  assign \new_[6038]_  = \new_[6037]_  | \new_[6028]_ ;
  assign \new_[6041]_  = \new_[442]_  | \new_[443]_ ;
  assign \new_[6044]_  = \new_[440]_  | \new_[441]_ ;
  assign \new_[6045]_  = \new_[6044]_  | \new_[6041]_ ;
  assign \new_[6048]_  = \new_[438]_  | \new_[439]_ ;
  assign \new_[6052]_  = \new_[435]_  | \new_[436]_ ;
  assign \new_[6053]_  = \new_[437]_  | \new_[6052]_ ;
  assign \new_[6054]_  = \new_[6053]_  | \new_[6048]_ ;
  assign \new_[6055]_  = \new_[6054]_  | \new_[6045]_ ;
  assign \new_[6056]_  = \new_[6055]_  | \new_[6038]_ ;
  assign \new_[6057]_  = \new_[6056]_  | \new_[6021]_ ;
  assign \new_[6058]_  = \new_[6057]_  | \new_[5986]_ ;
  assign \new_[6059]_  = \new_[6058]_  | \new_[5915]_ ;
  assign \new_[6062]_  = \new_[433]_  | \new_[434]_ ;
  assign \new_[6065]_  = \new_[431]_  | \new_[432]_ ;
  assign \new_[6066]_  = \new_[6065]_  | \new_[6062]_ ;
  assign \new_[6069]_  = \new_[429]_  | \new_[430]_ ;
  assign \new_[6073]_  = \new_[426]_  | \new_[427]_ ;
  assign \new_[6074]_  = \new_[428]_  | \new_[6073]_ ;
  assign \new_[6075]_  = \new_[6074]_  | \new_[6069]_ ;
  assign \new_[6076]_  = \new_[6075]_  | \new_[6066]_ ;
  assign \new_[6079]_  = \new_[424]_  | \new_[425]_ ;
  assign \new_[6082]_  = \new_[422]_  | \new_[423]_ ;
  assign \new_[6083]_  = \new_[6082]_  | \new_[6079]_ ;
  assign \new_[6086]_  = \new_[420]_  | \new_[421]_ ;
  assign \new_[6090]_  = \new_[417]_  | \new_[418]_ ;
  assign \new_[6091]_  = \new_[419]_  | \new_[6090]_ ;
  assign \new_[6092]_  = \new_[6091]_  | \new_[6086]_ ;
  assign \new_[6093]_  = \new_[6092]_  | \new_[6083]_ ;
  assign \new_[6094]_  = \new_[6093]_  | \new_[6076]_ ;
  assign \new_[6097]_  = \new_[415]_  | \new_[416]_ ;
  assign \new_[6100]_  = \new_[413]_  | \new_[414]_ ;
  assign \new_[6101]_  = \new_[6100]_  | \new_[6097]_ ;
  assign \new_[6104]_  = \new_[411]_  | \new_[412]_ ;
  assign \new_[6108]_  = \new_[408]_  | \new_[409]_ ;
  assign \new_[6109]_  = \new_[410]_  | \new_[6108]_ ;
  assign \new_[6110]_  = \new_[6109]_  | \new_[6104]_ ;
  assign \new_[6111]_  = \new_[6110]_  | \new_[6101]_ ;
  assign \new_[6114]_  = \new_[406]_  | \new_[407]_ ;
  assign \new_[6117]_  = \new_[404]_  | \new_[405]_ ;
  assign \new_[6118]_  = \new_[6117]_  | \new_[6114]_ ;
  assign \new_[6121]_  = \new_[402]_  | \new_[403]_ ;
  assign \new_[6125]_  = \new_[399]_  | \new_[400]_ ;
  assign \new_[6126]_  = \new_[401]_  | \new_[6125]_ ;
  assign \new_[6127]_  = \new_[6126]_  | \new_[6121]_ ;
  assign \new_[6128]_  = \new_[6127]_  | \new_[6118]_ ;
  assign \new_[6129]_  = \new_[6128]_  | \new_[6111]_ ;
  assign \new_[6130]_  = \new_[6129]_  | \new_[6094]_ ;
  assign \new_[6133]_  = \new_[397]_  | \new_[398]_ ;
  assign \new_[6136]_  = \new_[395]_  | \new_[396]_ ;
  assign \new_[6137]_  = \new_[6136]_  | \new_[6133]_ ;
  assign \new_[6140]_  = \new_[393]_  | \new_[394]_ ;
  assign \new_[6144]_  = \new_[390]_  | \new_[391]_ ;
  assign \new_[6145]_  = \new_[392]_  | \new_[6144]_ ;
  assign \new_[6146]_  = \new_[6145]_  | \new_[6140]_ ;
  assign \new_[6147]_  = \new_[6146]_  | \new_[6137]_ ;
  assign \new_[6150]_  = \new_[388]_  | \new_[389]_ ;
  assign \new_[6153]_  = \new_[386]_  | \new_[387]_ ;
  assign \new_[6154]_  = \new_[6153]_  | \new_[6150]_ ;
  assign \new_[6157]_  = \new_[384]_  | \new_[385]_ ;
  assign \new_[6161]_  = \new_[381]_  | \new_[382]_ ;
  assign \new_[6162]_  = \new_[383]_  | \new_[6161]_ ;
  assign \new_[6163]_  = \new_[6162]_  | \new_[6157]_ ;
  assign \new_[6164]_  = \new_[6163]_  | \new_[6154]_ ;
  assign \new_[6165]_  = \new_[6164]_  | \new_[6147]_ ;
  assign \new_[6168]_  = \new_[379]_  | \new_[380]_ ;
  assign \new_[6171]_  = \new_[377]_  | \new_[378]_ ;
  assign \new_[6172]_  = \new_[6171]_  | \new_[6168]_ ;
  assign \new_[6175]_  = \new_[375]_  | \new_[376]_ ;
  assign \new_[6179]_  = \new_[372]_  | \new_[373]_ ;
  assign \new_[6180]_  = \new_[374]_  | \new_[6179]_ ;
  assign \new_[6181]_  = \new_[6180]_  | \new_[6175]_ ;
  assign \new_[6182]_  = \new_[6181]_  | \new_[6172]_ ;
  assign \new_[6185]_  = \new_[370]_  | \new_[371]_ ;
  assign \new_[6188]_  = \new_[368]_  | \new_[369]_ ;
  assign \new_[6189]_  = \new_[6188]_  | \new_[6185]_ ;
  assign \new_[6192]_  = \new_[366]_  | \new_[367]_ ;
  assign \new_[6196]_  = \new_[363]_  | \new_[364]_ ;
  assign \new_[6197]_  = \new_[365]_  | \new_[6196]_ ;
  assign \new_[6198]_  = \new_[6197]_  | \new_[6192]_ ;
  assign \new_[6199]_  = \new_[6198]_  | \new_[6189]_ ;
  assign \new_[6200]_  = \new_[6199]_  | \new_[6182]_ ;
  assign \new_[6201]_  = \new_[6200]_  | \new_[6165]_ ;
  assign \new_[6202]_  = \new_[6201]_  | \new_[6130]_ ;
  assign \new_[6205]_  = \new_[361]_  | \new_[362]_ ;
  assign \new_[6208]_  = \new_[359]_  | \new_[360]_ ;
  assign \new_[6209]_  = \new_[6208]_  | \new_[6205]_ ;
  assign \new_[6212]_  = \new_[357]_  | \new_[358]_ ;
  assign \new_[6216]_  = \new_[354]_  | \new_[355]_ ;
  assign \new_[6217]_  = \new_[356]_  | \new_[6216]_ ;
  assign \new_[6218]_  = \new_[6217]_  | \new_[6212]_ ;
  assign \new_[6219]_  = \new_[6218]_  | \new_[6209]_ ;
  assign \new_[6222]_  = \new_[352]_  | \new_[353]_ ;
  assign \new_[6225]_  = \new_[350]_  | \new_[351]_ ;
  assign \new_[6226]_  = \new_[6225]_  | \new_[6222]_ ;
  assign \new_[6229]_  = \new_[348]_  | \new_[349]_ ;
  assign \new_[6233]_  = \new_[345]_  | \new_[346]_ ;
  assign \new_[6234]_  = \new_[347]_  | \new_[6233]_ ;
  assign \new_[6235]_  = \new_[6234]_  | \new_[6229]_ ;
  assign \new_[6236]_  = \new_[6235]_  | \new_[6226]_ ;
  assign \new_[6237]_  = \new_[6236]_  | \new_[6219]_ ;
  assign \new_[6240]_  = \new_[343]_  | \new_[344]_ ;
  assign \new_[6243]_  = \new_[341]_  | \new_[342]_ ;
  assign \new_[6244]_  = \new_[6243]_  | \new_[6240]_ ;
  assign \new_[6247]_  = \new_[339]_  | \new_[340]_ ;
  assign \new_[6251]_  = \new_[336]_  | \new_[337]_ ;
  assign \new_[6252]_  = \new_[338]_  | \new_[6251]_ ;
  assign \new_[6253]_  = \new_[6252]_  | \new_[6247]_ ;
  assign \new_[6254]_  = \new_[6253]_  | \new_[6244]_ ;
  assign \new_[6257]_  = \new_[334]_  | \new_[335]_ ;
  assign \new_[6260]_  = \new_[332]_  | \new_[333]_ ;
  assign \new_[6261]_  = \new_[6260]_  | \new_[6257]_ ;
  assign \new_[6264]_  = \new_[330]_  | \new_[331]_ ;
  assign \new_[6268]_  = \new_[327]_  | \new_[328]_ ;
  assign \new_[6269]_  = \new_[329]_  | \new_[6268]_ ;
  assign \new_[6270]_  = \new_[6269]_  | \new_[6264]_ ;
  assign \new_[6271]_  = \new_[6270]_  | \new_[6261]_ ;
  assign \new_[6272]_  = \new_[6271]_  | \new_[6254]_ ;
  assign \new_[6273]_  = \new_[6272]_  | \new_[6237]_ ;
  assign \new_[6276]_  = \new_[325]_  | \new_[326]_ ;
  assign \new_[6279]_  = \new_[323]_  | \new_[324]_ ;
  assign \new_[6280]_  = \new_[6279]_  | \new_[6276]_ ;
  assign \new_[6283]_  = \new_[321]_  | \new_[322]_ ;
  assign \new_[6287]_  = \new_[318]_  | \new_[319]_ ;
  assign \new_[6288]_  = \new_[320]_  | \new_[6287]_ ;
  assign \new_[6289]_  = \new_[6288]_  | \new_[6283]_ ;
  assign \new_[6290]_  = \new_[6289]_  | \new_[6280]_ ;
  assign \new_[6293]_  = \new_[316]_  | \new_[317]_ ;
  assign \new_[6296]_  = \new_[314]_  | \new_[315]_ ;
  assign \new_[6297]_  = \new_[6296]_  | \new_[6293]_ ;
  assign \new_[6300]_  = \new_[312]_  | \new_[313]_ ;
  assign \new_[6304]_  = \new_[309]_  | \new_[310]_ ;
  assign \new_[6305]_  = \new_[311]_  | \new_[6304]_ ;
  assign \new_[6306]_  = \new_[6305]_  | \new_[6300]_ ;
  assign \new_[6307]_  = \new_[6306]_  | \new_[6297]_ ;
  assign \new_[6308]_  = \new_[6307]_  | \new_[6290]_ ;
  assign \new_[6311]_  = \new_[307]_  | \new_[308]_ ;
  assign \new_[6314]_  = \new_[305]_  | \new_[306]_ ;
  assign \new_[6315]_  = \new_[6314]_  | \new_[6311]_ ;
  assign \new_[6318]_  = \new_[303]_  | \new_[304]_ ;
  assign \new_[6322]_  = \new_[300]_  | \new_[301]_ ;
  assign \new_[6323]_  = \new_[302]_  | \new_[6322]_ ;
  assign \new_[6324]_  = \new_[6323]_  | \new_[6318]_ ;
  assign \new_[6325]_  = \new_[6324]_  | \new_[6315]_ ;
  assign \new_[6328]_  = \new_[298]_  | \new_[299]_ ;
  assign \new_[6332]_  = \new_[295]_  | \new_[296]_ ;
  assign \new_[6333]_  = \new_[297]_  | \new_[6332]_ ;
  assign \new_[6334]_  = \new_[6333]_  | \new_[6328]_ ;
  assign \new_[6337]_  = \new_[293]_  | \new_[294]_ ;
  assign \new_[6341]_  = \new_[290]_  | \new_[291]_ ;
  assign \new_[6342]_  = \new_[292]_  | \new_[6341]_ ;
  assign \new_[6343]_  = \new_[6342]_  | \new_[6337]_ ;
  assign \new_[6344]_  = \new_[6343]_  | \new_[6334]_ ;
  assign \new_[6345]_  = \new_[6344]_  | \new_[6325]_ ;
  assign \new_[6346]_  = \new_[6345]_  | \new_[6308]_ ;
  assign \new_[6347]_  = \new_[6346]_  | \new_[6273]_ ;
  assign \new_[6348]_  = \new_[6347]_  | \new_[6202]_ ;
  assign \new_[6349]_  = \new_[6348]_  | \new_[6059]_ ;
  assign \new_[6352]_  = \new_[288]_  | \new_[289]_ ;
  assign \new_[6355]_  = \new_[286]_  | \new_[287]_ ;
  assign \new_[6356]_  = \new_[6355]_  | \new_[6352]_ ;
  assign \new_[6359]_  = \new_[284]_  | \new_[285]_ ;
  assign \new_[6363]_  = \new_[281]_  | \new_[282]_ ;
  assign \new_[6364]_  = \new_[283]_  | \new_[6363]_ ;
  assign \new_[6365]_  = \new_[6364]_  | \new_[6359]_ ;
  assign \new_[6366]_  = \new_[6365]_  | \new_[6356]_ ;
  assign \new_[6369]_  = \new_[279]_  | \new_[280]_ ;
  assign \new_[6372]_  = \new_[277]_  | \new_[278]_ ;
  assign \new_[6373]_  = \new_[6372]_  | \new_[6369]_ ;
  assign \new_[6376]_  = \new_[275]_  | \new_[276]_ ;
  assign \new_[6380]_  = \new_[272]_  | \new_[273]_ ;
  assign \new_[6381]_  = \new_[274]_  | \new_[6380]_ ;
  assign \new_[6382]_  = \new_[6381]_  | \new_[6376]_ ;
  assign \new_[6383]_  = \new_[6382]_  | \new_[6373]_ ;
  assign \new_[6384]_  = \new_[6383]_  | \new_[6366]_ ;
  assign \new_[6387]_  = \new_[270]_  | \new_[271]_ ;
  assign \new_[6390]_  = \new_[268]_  | \new_[269]_ ;
  assign \new_[6391]_  = \new_[6390]_  | \new_[6387]_ ;
  assign \new_[6394]_  = \new_[266]_  | \new_[267]_ ;
  assign \new_[6398]_  = \new_[263]_  | \new_[264]_ ;
  assign \new_[6399]_  = \new_[265]_  | \new_[6398]_ ;
  assign \new_[6400]_  = \new_[6399]_  | \new_[6394]_ ;
  assign \new_[6401]_  = \new_[6400]_  | \new_[6391]_ ;
  assign \new_[6404]_  = \new_[261]_  | \new_[262]_ ;
  assign \new_[6407]_  = \new_[259]_  | \new_[260]_ ;
  assign \new_[6408]_  = \new_[6407]_  | \new_[6404]_ ;
  assign \new_[6411]_  = \new_[257]_  | \new_[258]_ ;
  assign \new_[6415]_  = \new_[254]_  | \new_[255]_ ;
  assign \new_[6416]_  = \new_[256]_  | \new_[6415]_ ;
  assign \new_[6417]_  = \new_[6416]_  | \new_[6411]_ ;
  assign \new_[6418]_  = \new_[6417]_  | \new_[6408]_ ;
  assign \new_[6419]_  = \new_[6418]_  | \new_[6401]_ ;
  assign \new_[6420]_  = \new_[6419]_  | \new_[6384]_ ;
  assign \new_[6423]_  = \new_[252]_  | \new_[253]_ ;
  assign \new_[6426]_  = \new_[250]_  | \new_[251]_ ;
  assign \new_[6427]_  = \new_[6426]_  | \new_[6423]_ ;
  assign \new_[6430]_  = \new_[248]_  | \new_[249]_ ;
  assign \new_[6434]_  = \new_[245]_  | \new_[246]_ ;
  assign \new_[6435]_  = \new_[247]_  | \new_[6434]_ ;
  assign \new_[6436]_  = \new_[6435]_  | \new_[6430]_ ;
  assign \new_[6437]_  = \new_[6436]_  | \new_[6427]_ ;
  assign \new_[6440]_  = \new_[243]_  | \new_[244]_ ;
  assign \new_[6443]_  = \new_[241]_  | \new_[242]_ ;
  assign \new_[6444]_  = \new_[6443]_  | \new_[6440]_ ;
  assign \new_[6447]_  = \new_[239]_  | \new_[240]_ ;
  assign \new_[6451]_  = \new_[236]_  | \new_[237]_ ;
  assign \new_[6452]_  = \new_[238]_  | \new_[6451]_ ;
  assign \new_[6453]_  = \new_[6452]_  | \new_[6447]_ ;
  assign \new_[6454]_  = \new_[6453]_  | \new_[6444]_ ;
  assign \new_[6455]_  = \new_[6454]_  | \new_[6437]_ ;
  assign \new_[6458]_  = \new_[234]_  | \new_[235]_ ;
  assign \new_[6461]_  = \new_[232]_  | \new_[233]_ ;
  assign \new_[6462]_  = \new_[6461]_  | \new_[6458]_ ;
  assign \new_[6465]_  = \new_[230]_  | \new_[231]_ ;
  assign \new_[6469]_  = \new_[227]_  | \new_[228]_ ;
  assign \new_[6470]_  = \new_[229]_  | \new_[6469]_ ;
  assign \new_[6471]_  = \new_[6470]_  | \new_[6465]_ ;
  assign \new_[6472]_  = \new_[6471]_  | \new_[6462]_ ;
  assign \new_[6475]_  = \new_[225]_  | \new_[226]_ ;
  assign \new_[6478]_  = \new_[223]_  | \new_[224]_ ;
  assign \new_[6479]_  = \new_[6478]_  | \new_[6475]_ ;
  assign \new_[6482]_  = \new_[221]_  | \new_[222]_ ;
  assign \new_[6486]_  = \new_[218]_  | \new_[219]_ ;
  assign \new_[6487]_  = \new_[220]_  | \new_[6486]_ ;
  assign \new_[6488]_  = \new_[6487]_  | \new_[6482]_ ;
  assign \new_[6489]_  = \new_[6488]_  | \new_[6479]_ ;
  assign \new_[6490]_  = \new_[6489]_  | \new_[6472]_ ;
  assign \new_[6491]_  = \new_[6490]_  | \new_[6455]_ ;
  assign \new_[6492]_  = \new_[6491]_  | \new_[6420]_ ;
  assign \new_[6495]_  = \new_[216]_  | \new_[217]_ ;
  assign \new_[6498]_  = \new_[214]_  | \new_[215]_ ;
  assign \new_[6499]_  = \new_[6498]_  | \new_[6495]_ ;
  assign \new_[6502]_  = \new_[212]_  | \new_[213]_ ;
  assign \new_[6506]_  = \new_[209]_  | \new_[210]_ ;
  assign \new_[6507]_  = \new_[211]_  | \new_[6506]_ ;
  assign \new_[6508]_  = \new_[6507]_  | \new_[6502]_ ;
  assign \new_[6509]_  = \new_[6508]_  | \new_[6499]_ ;
  assign \new_[6512]_  = \new_[207]_  | \new_[208]_ ;
  assign \new_[6515]_  = \new_[205]_  | \new_[206]_ ;
  assign \new_[6516]_  = \new_[6515]_  | \new_[6512]_ ;
  assign \new_[6519]_  = \new_[203]_  | \new_[204]_ ;
  assign \new_[6523]_  = \new_[200]_  | \new_[201]_ ;
  assign \new_[6524]_  = \new_[202]_  | \new_[6523]_ ;
  assign \new_[6525]_  = \new_[6524]_  | \new_[6519]_ ;
  assign \new_[6526]_  = \new_[6525]_  | \new_[6516]_ ;
  assign \new_[6527]_  = \new_[6526]_  | \new_[6509]_ ;
  assign \new_[6530]_  = \new_[198]_  | \new_[199]_ ;
  assign \new_[6533]_  = \new_[196]_  | \new_[197]_ ;
  assign \new_[6534]_  = \new_[6533]_  | \new_[6530]_ ;
  assign \new_[6537]_  = \new_[194]_  | \new_[195]_ ;
  assign \new_[6541]_  = \new_[191]_  | \new_[192]_ ;
  assign \new_[6542]_  = \new_[193]_  | \new_[6541]_ ;
  assign \new_[6543]_  = \new_[6542]_  | \new_[6537]_ ;
  assign \new_[6544]_  = \new_[6543]_  | \new_[6534]_ ;
  assign \new_[6547]_  = \new_[189]_  | \new_[190]_ ;
  assign \new_[6550]_  = \new_[187]_  | \new_[188]_ ;
  assign \new_[6551]_  = \new_[6550]_  | \new_[6547]_ ;
  assign \new_[6554]_  = \new_[185]_  | \new_[186]_ ;
  assign \new_[6558]_  = \new_[182]_  | \new_[183]_ ;
  assign \new_[6559]_  = \new_[184]_  | \new_[6558]_ ;
  assign \new_[6560]_  = \new_[6559]_  | \new_[6554]_ ;
  assign \new_[6561]_  = \new_[6560]_  | \new_[6551]_ ;
  assign \new_[6562]_  = \new_[6561]_  | \new_[6544]_ ;
  assign \new_[6563]_  = \new_[6562]_  | \new_[6527]_ ;
  assign \new_[6566]_  = \new_[180]_  | \new_[181]_ ;
  assign \new_[6569]_  = \new_[178]_  | \new_[179]_ ;
  assign \new_[6570]_  = \new_[6569]_  | \new_[6566]_ ;
  assign \new_[6573]_  = \new_[176]_  | \new_[177]_ ;
  assign \new_[6577]_  = \new_[173]_  | \new_[174]_ ;
  assign \new_[6578]_  = \new_[175]_  | \new_[6577]_ ;
  assign \new_[6579]_  = \new_[6578]_  | \new_[6573]_ ;
  assign \new_[6580]_  = \new_[6579]_  | \new_[6570]_ ;
  assign \new_[6583]_  = \new_[171]_  | \new_[172]_ ;
  assign \new_[6586]_  = \new_[169]_  | \new_[170]_ ;
  assign \new_[6587]_  = \new_[6586]_  | \new_[6583]_ ;
  assign \new_[6590]_  = \new_[167]_  | \new_[168]_ ;
  assign \new_[6594]_  = \new_[164]_  | \new_[165]_ ;
  assign \new_[6595]_  = \new_[166]_  | \new_[6594]_ ;
  assign \new_[6596]_  = \new_[6595]_  | \new_[6590]_ ;
  assign \new_[6597]_  = \new_[6596]_  | \new_[6587]_ ;
  assign \new_[6598]_  = \new_[6597]_  | \new_[6580]_ ;
  assign \new_[6601]_  = \new_[162]_  | \new_[163]_ ;
  assign \new_[6604]_  = \new_[160]_  | \new_[161]_ ;
  assign \new_[6605]_  = \new_[6604]_  | \new_[6601]_ ;
  assign \new_[6608]_  = \new_[158]_  | \new_[159]_ ;
  assign \new_[6612]_  = \new_[155]_  | \new_[156]_ ;
  assign \new_[6613]_  = \new_[157]_  | \new_[6612]_ ;
  assign \new_[6614]_  = \new_[6613]_  | \new_[6608]_ ;
  assign \new_[6615]_  = \new_[6614]_  | \new_[6605]_ ;
  assign \new_[6618]_  = \new_[153]_  | \new_[154]_ ;
  assign \new_[6621]_  = \new_[151]_  | \new_[152]_ ;
  assign \new_[6622]_  = \new_[6621]_  | \new_[6618]_ ;
  assign \new_[6625]_  = \new_[149]_  | \new_[150]_ ;
  assign \new_[6629]_  = \new_[146]_  | \new_[147]_ ;
  assign \new_[6630]_  = \new_[148]_  | \new_[6629]_ ;
  assign \new_[6631]_  = \new_[6630]_  | \new_[6625]_ ;
  assign \new_[6632]_  = \new_[6631]_  | \new_[6622]_ ;
  assign \new_[6633]_  = \new_[6632]_  | \new_[6615]_ ;
  assign \new_[6634]_  = \new_[6633]_  | \new_[6598]_ ;
  assign \new_[6635]_  = \new_[6634]_  | \new_[6563]_ ;
  assign \new_[6636]_  = \new_[6635]_  | \new_[6492]_ ;
  assign \new_[6639]_  = \new_[144]_  | \new_[145]_ ;
  assign \new_[6642]_  = \new_[142]_  | \new_[143]_ ;
  assign \new_[6643]_  = \new_[6642]_  | \new_[6639]_ ;
  assign \new_[6646]_  = \new_[140]_  | \new_[141]_ ;
  assign \new_[6650]_  = \new_[137]_  | \new_[138]_ ;
  assign \new_[6651]_  = \new_[139]_  | \new_[6650]_ ;
  assign \new_[6652]_  = \new_[6651]_  | \new_[6646]_ ;
  assign \new_[6653]_  = \new_[6652]_  | \new_[6643]_ ;
  assign \new_[6656]_  = \new_[135]_  | \new_[136]_ ;
  assign \new_[6659]_  = \new_[133]_  | \new_[134]_ ;
  assign \new_[6660]_  = \new_[6659]_  | \new_[6656]_ ;
  assign \new_[6663]_  = \new_[131]_  | \new_[132]_ ;
  assign \new_[6667]_  = \new_[128]_  | \new_[129]_ ;
  assign \new_[6668]_  = \new_[130]_  | \new_[6667]_ ;
  assign \new_[6669]_  = \new_[6668]_  | \new_[6663]_ ;
  assign \new_[6670]_  = \new_[6669]_  | \new_[6660]_ ;
  assign \new_[6671]_  = \new_[6670]_  | \new_[6653]_ ;
  assign \new_[6674]_  = \new_[126]_  | \new_[127]_ ;
  assign \new_[6677]_  = \new_[124]_  | \new_[125]_ ;
  assign \new_[6678]_  = \new_[6677]_  | \new_[6674]_ ;
  assign \new_[6681]_  = \new_[122]_  | \new_[123]_ ;
  assign \new_[6685]_  = \new_[119]_  | \new_[120]_ ;
  assign \new_[6686]_  = \new_[121]_  | \new_[6685]_ ;
  assign \new_[6687]_  = \new_[6686]_  | \new_[6681]_ ;
  assign \new_[6688]_  = \new_[6687]_  | \new_[6678]_ ;
  assign \new_[6691]_  = \new_[117]_  | \new_[118]_ ;
  assign \new_[6694]_  = \new_[115]_  | \new_[116]_ ;
  assign \new_[6695]_  = \new_[6694]_  | \new_[6691]_ ;
  assign \new_[6698]_  = \new_[113]_  | \new_[114]_ ;
  assign \new_[6702]_  = \new_[110]_  | \new_[111]_ ;
  assign \new_[6703]_  = \new_[112]_  | \new_[6702]_ ;
  assign \new_[6704]_  = \new_[6703]_  | \new_[6698]_ ;
  assign \new_[6705]_  = \new_[6704]_  | \new_[6695]_ ;
  assign \new_[6706]_  = \new_[6705]_  | \new_[6688]_ ;
  assign \new_[6707]_  = \new_[6706]_  | \new_[6671]_ ;
  assign \new_[6710]_  = \new_[108]_  | \new_[109]_ ;
  assign \new_[6713]_  = \new_[106]_  | \new_[107]_ ;
  assign \new_[6714]_  = \new_[6713]_  | \new_[6710]_ ;
  assign \new_[6717]_  = \new_[104]_  | \new_[105]_ ;
  assign \new_[6721]_  = \new_[101]_  | \new_[102]_ ;
  assign \new_[6722]_  = \new_[103]_  | \new_[6721]_ ;
  assign \new_[6723]_  = \new_[6722]_  | \new_[6717]_ ;
  assign \new_[6724]_  = \new_[6723]_  | \new_[6714]_ ;
  assign \new_[6727]_  = \new_[99]_  | \new_[100]_ ;
  assign \new_[6730]_  = \new_[97]_  | \new_[98]_ ;
  assign \new_[6731]_  = \new_[6730]_  | \new_[6727]_ ;
  assign \new_[6734]_  = \new_[95]_  | \new_[96]_ ;
  assign \new_[6738]_  = \new_[92]_  | \new_[93]_ ;
  assign \new_[6739]_  = \new_[94]_  | \new_[6738]_ ;
  assign \new_[6740]_  = \new_[6739]_  | \new_[6734]_ ;
  assign \new_[6741]_  = \new_[6740]_  | \new_[6731]_ ;
  assign \new_[6742]_  = \new_[6741]_  | \new_[6724]_ ;
  assign \new_[6745]_  = \new_[90]_  | \new_[91]_ ;
  assign \new_[6748]_  = \new_[88]_  | \new_[89]_ ;
  assign \new_[6749]_  = \new_[6748]_  | \new_[6745]_ ;
  assign \new_[6752]_  = \new_[86]_  | \new_[87]_ ;
  assign \new_[6756]_  = \new_[83]_  | \new_[84]_ ;
  assign \new_[6757]_  = \new_[85]_  | \new_[6756]_ ;
  assign \new_[6758]_  = \new_[6757]_  | \new_[6752]_ ;
  assign \new_[6759]_  = \new_[6758]_  | \new_[6749]_ ;
  assign \new_[6762]_  = \new_[81]_  | \new_[82]_ ;
  assign \new_[6765]_  = \new_[79]_  | \new_[80]_ ;
  assign \new_[6766]_  = \new_[6765]_  | \new_[6762]_ ;
  assign \new_[6769]_  = \new_[77]_  | \new_[78]_ ;
  assign \new_[6773]_  = \new_[74]_  | \new_[75]_ ;
  assign \new_[6774]_  = \new_[76]_  | \new_[6773]_ ;
  assign \new_[6775]_  = \new_[6774]_  | \new_[6769]_ ;
  assign \new_[6776]_  = \new_[6775]_  | \new_[6766]_ ;
  assign \new_[6777]_  = \new_[6776]_  | \new_[6759]_ ;
  assign \new_[6778]_  = \new_[6777]_  | \new_[6742]_ ;
  assign \new_[6779]_  = \new_[6778]_  | \new_[6707]_ ;
  assign \new_[6782]_  = \new_[72]_  | \new_[73]_ ;
  assign \new_[6785]_  = \new_[70]_  | \new_[71]_ ;
  assign \new_[6786]_  = \new_[6785]_  | \new_[6782]_ ;
  assign \new_[6789]_  = \new_[68]_  | \new_[69]_ ;
  assign \new_[6793]_  = \new_[65]_  | \new_[66]_ ;
  assign \new_[6794]_  = \new_[67]_  | \new_[6793]_ ;
  assign \new_[6795]_  = \new_[6794]_  | \new_[6789]_ ;
  assign \new_[6796]_  = \new_[6795]_  | \new_[6786]_ ;
  assign \new_[6799]_  = \new_[63]_  | \new_[64]_ ;
  assign \new_[6802]_  = \new_[61]_  | \new_[62]_ ;
  assign \new_[6803]_  = \new_[6802]_  | \new_[6799]_ ;
  assign \new_[6806]_  = \new_[59]_  | \new_[60]_ ;
  assign \new_[6810]_  = \new_[56]_  | \new_[57]_ ;
  assign \new_[6811]_  = \new_[58]_  | \new_[6810]_ ;
  assign \new_[6812]_  = \new_[6811]_  | \new_[6806]_ ;
  assign \new_[6813]_  = \new_[6812]_  | \new_[6803]_ ;
  assign \new_[6814]_  = \new_[6813]_  | \new_[6796]_ ;
  assign \new_[6817]_  = \new_[54]_  | \new_[55]_ ;
  assign \new_[6820]_  = \new_[52]_  | \new_[53]_ ;
  assign \new_[6821]_  = \new_[6820]_  | \new_[6817]_ ;
  assign \new_[6824]_  = \new_[50]_  | \new_[51]_ ;
  assign \new_[6828]_  = \new_[47]_  | \new_[48]_ ;
  assign \new_[6829]_  = \new_[49]_  | \new_[6828]_ ;
  assign \new_[6830]_  = \new_[6829]_  | \new_[6824]_ ;
  assign \new_[6831]_  = \new_[6830]_  | \new_[6821]_ ;
  assign \new_[6834]_  = \new_[45]_  | \new_[46]_ ;
  assign \new_[6837]_  = \new_[43]_  | \new_[44]_ ;
  assign \new_[6838]_  = \new_[6837]_  | \new_[6834]_ ;
  assign \new_[6841]_  = \new_[41]_  | \new_[42]_ ;
  assign \new_[6845]_  = \new_[38]_  | \new_[39]_ ;
  assign \new_[6846]_  = \new_[40]_  | \new_[6845]_ ;
  assign \new_[6847]_  = \new_[6846]_  | \new_[6841]_ ;
  assign \new_[6848]_  = \new_[6847]_  | \new_[6838]_ ;
  assign \new_[6849]_  = \new_[6848]_  | \new_[6831]_ ;
  assign \new_[6850]_  = \new_[6849]_  | \new_[6814]_ ;
  assign \new_[6853]_  = \new_[36]_  | \new_[37]_ ;
  assign \new_[6856]_  = \new_[34]_  | \new_[35]_ ;
  assign \new_[6857]_  = \new_[6856]_  | \new_[6853]_ ;
  assign \new_[6860]_  = \new_[32]_  | \new_[33]_ ;
  assign \new_[6864]_  = \new_[29]_  | \new_[30]_ ;
  assign \new_[6865]_  = \new_[31]_  | \new_[6864]_ ;
  assign \new_[6866]_  = \new_[6865]_  | \new_[6860]_ ;
  assign \new_[6867]_  = \new_[6866]_  | \new_[6857]_ ;
  assign \new_[6870]_  = \new_[27]_  | \new_[28]_ ;
  assign \new_[6873]_  = \new_[25]_  | \new_[26]_ ;
  assign \new_[6874]_  = \new_[6873]_  | \new_[6870]_ ;
  assign \new_[6877]_  = \new_[23]_  | \new_[24]_ ;
  assign \new_[6881]_  = \new_[20]_  | \new_[21]_ ;
  assign \new_[6882]_  = \new_[22]_  | \new_[6881]_ ;
  assign \new_[6883]_  = \new_[6882]_  | \new_[6877]_ ;
  assign \new_[6884]_  = \new_[6883]_  | \new_[6874]_ ;
  assign \new_[6885]_  = \new_[6884]_  | \new_[6867]_ ;
  assign \new_[6888]_  = \new_[18]_  | \new_[19]_ ;
  assign \new_[6891]_  = \new_[16]_  | \new_[17]_ ;
  assign \new_[6892]_  = \new_[6891]_  | \new_[6888]_ ;
  assign \new_[6895]_  = \new_[14]_  | \new_[15]_ ;
  assign \new_[6899]_  = \new_[11]_  | \new_[12]_ ;
  assign \new_[6900]_  = \new_[13]_  | \new_[6899]_ ;
  assign \new_[6901]_  = \new_[6900]_  | \new_[6895]_ ;
  assign \new_[6902]_  = \new_[6901]_  | \new_[6892]_ ;
  assign \new_[6905]_  = \new_[9]_  | \new_[10]_ ;
  assign \new_[6909]_  = \new_[6]_  | \new_[7]_ ;
  assign \new_[6910]_  = \new_[8]_  | \new_[6909]_ ;
  assign \new_[6911]_  = \new_[6910]_  | \new_[6905]_ ;
  assign \new_[6914]_  = \new_[4]_  | \new_[5]_ ;
  assign \new_[6918]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[6919]_  = \new_[3]_  | \new_[6918]_ ;
  assign \new_[6920]_  = \new_[6919]_  | \new_[6914]_ ;
  assign \new_[6921]_  = \new_[6920]_  | \new_[6911]_ ;
  assign \new_[6922]_  = \new_[6921]_  | \new_[6902]_ ;
  assign \new_[6923]_  = \new_[6922]_  | \new_[6885]_ ;
  assign \new_[6924]_  = \new_[6923]_  | \new_[6850]_ ;
  assign \new_[6925]_  = \new_[6924]_  | \new_[6779]_ ;
  assign \new_[6926]_  = \new_[6925]_  | \new_[6636]_ ;
  assign \new_[6927]_  = \new_[6926]_  | \new_[6349]_ ;
  assign \new_[6928]_  = \new_[6927]_  | \new_[5772]_ ;
  assign \new_[6932]_  = ~A202 & ~A201;
  assign \new_[6933]_  = A169 & \new_[6932]_ ;
  assign \new_[6937]_  = A301 & A235;
  assign \new_[6938]_  = ~A203 & \new_[6937]_ ;
  assign \new_[6942]_  = ~A202 & ~A201;
  assign \new_[6943]_  = A169 & \new_[6942]_ ;
  assign \new_[6947]_  = A268 & A235;
  assign \new_[6948]_  = ~A203 & \new_[6947]_ ;
  assign \new_[6952]_  = ~A200 & ~A199;
  assign \new_[6953]_  = A169 & \new_[6952]_ ;
  assign \new_[6957]_  = A301 & A235;
  assign \new_[6958]_  = ~A202 & \new_[6957]_ ;
  assign \new_[6962]_  = ~A200 & ~A199;
  assign \new_[6963]_  = A169 & \new_[6962]_ ;
  assign \new_[6967]_  = A268 & A235;
  assign \new_[6968]_  = ~A202 & \new_[6967]_ ;
  assign \new_[6972]_  = ~A166 & ~A167;
  assign \new_[6973]_  = ~A169 & \new_[6972]_ ;
  assign \new_[6977]_  = A301 & A235;
  assign \new_[6978]_  = A202 & \new_[6977]_ ;
  assign \new_[6982]_  = ~A166 & ~A167;
  assign \new_[6983]_  = ~A169 & \new_[6982]_ ;
  assign \new_[6987]_  = A268 & A235;
  assign \new_[6988]_  = A202 & \new_[6987]_ ;
  assign \new_[6992]_  = ~A168 & ~A169;
  assign \new_[6993]_  = ~A170 & \new_[6992]_ ;
  assign \new_[6997]_  = A301 & A235;
  assign \new_[6998]_  = A202 & \new_[6997]_ ;
  assign \new_[7002]_  = ~A168 & ~A169;
  assign \new_[7003]_  = ~A170 & \new_[7002]_ ;
  assign \new_[7007]_  = A268 & A235;
  assign \new_[7008]_  = A202 & \new_[7007]_ ;
  assign \new_[7012]_  = ~A201 & A166;
  assign \new_[7013]_  = A168 & \new_[7012]_ ;
  assign \new_[7016]_  = ~A203 & ~A202;
  assign \new_[7019]_  = A301 & A235;
  assign \new_[7020]_  = \new_[7019]_  & \new_[7016]_ ;
  assign \new_[7024]_  = ~A201 & A166;
  assign \new_[7025]_  = A168 & \new_[7024]_ ;
  assign \new_[7028]_  = ~A203 & ~A202;
  assign \new_[7031]_  = A268 & A235;
  assign \new_[7032]_  = \new_[7031]_  & \new_[7028]_ ;
  assign \new_[7036]_  = ~A199 & A166;
  assign \new_[7037]_  = A168 & \new_[7036]_ ;
  assign \new_[7040]_  = ~A202 & ~A200;
  assign \new_[7043]_  = A301 & A235;
  assign \new_[7044]_  = \new_[7043]_  & \new_[7040]_ ;
  assign \new_[7048]_  = ~A199 & A166;
  assign \new_[7049]_  = A168 & \new_[7048]_ ;
  assign \new_[7052]_  = ~A202 & ~A200;
  assign \new_[7055]_  = A268 & A235;
  assign \new_[7056]_  = \new_[7055]_  & \new_[7052]_ ;
  assign \new_[7060]_  = ~A201 & A167;
  assign \new_[7061]_  = A168 & \new_[7060]_ ;
  assign \new_[7064]_  = ~A203 & ~A202;
  assign \new_[7067]_  = A301 & A235;
  assign \new_[7068]_  = \new_[7067]_  & \new_[7064]_ ;
  assign \new_[7072]_  = ~A201 & A167;
  assign \new_[7073]_  = A168 & \new_[7072]_ ;
  assign \new_[7076]_  = ~A203 & ~A202;
  assign \new_[7079]_  = A268 & A235;
  assign \new_[7080]_  = \new_[7079]_  & \new_[7076]_ ;
  assign \new_[7084]_  = ~A199 & A167;
  assign \new_[7085]_  = A168 & \new_[7084]_ ;
  assign \new_[7088]_  = ~A202 & ~A200;
  assign \new_[7091]_  = A301 & A235;
  assign \new_[7092]_  = \new_[7091]_  & \new_[7088]_ ;
  assign \new_[7096]_  = ~A199 & A167;
  assign \new_[7097]_  = A168 & \new_[7096]_ ;
  assign \new_[7100]_  = ~A202 & ~A200;
  assign \new_[7103]_  = A268 & A235;
  assign \new_[7104]_  = \new_[7103]_  & \new_[7100]_ ;
  assign \new_[7108]_  = ~A202 & ~A201;
  assign \new_[7109]_  = A169 & \new_[7108]_ ;
  assign \new_[7112]_  = A235 & ~A203;
  assign \new_[7115]_  = A300 & A299;
  assign \new_[7116]_  = \new_[7115]_  & \new_[7112]_ ;
  assign \new_[7120]_  = ~A202 & ~A201;
  assign \new_[7121]_  = A169 & \new_[7120]_ ;
  assign \new_[7124]_  = A235 & ~A203;
  assign \new_[7127]_  = A300 & A298;
  assign \new_[7128]_  = \new_[7127]_  & \new_[7124]_ ;
  assign \new_[7132]_  = ~A202 & ~A201;
  assign \new_[7133]_  = A169 & \new_[7132]_ ;
  assign \new_[7136]_  = A235 & ~A203;
  assign \new_[7139]_  = A267 & A265;
  assign \new_[7140]_  = \new_[7139]_  & \new_[7136]_ ;
  assign \new_[7144]_  = ~A202 & ~A201;
  assign \new_[7145]_  = A169 & \new_[7144]_ ;
  assign \new_[7148]_  = A235 & ~A203;
  assign \new_[7151]_  = A267 & A266;
  assign \new_[7152]_  = \new_[7151]_  & \new_[7148]_ ;
  assign \new_[7156]_  = ~A202 & ~A201;
  assign \new_[7157]_  = A169 & \new_[7156]_ ;
  assign \new_[7160]_  = A232 & ~A203;
  assign \new_[7163]_  = A301 & A234;
  assign \new_[7164]_  = \new_[7163]_  & \new_[7160]_ ;
  assign \new_[7168]_  = ~A202 & ~A201;
  assign \new_[7169]_  = A169 & \new_[7168]_ ;
  assign \new_[7172]_  = A232 & ~A203;
  assign \new_[7175]_  = A268 & A234;
  assign \new_[7176]_  = \new_[7175]_  & \new_[7172]_ ;
  assign \new_[7180]_  = ~A202 & ~A201;
  assign \new_[7181]_  = A169 & \new_[7180]_ ;
  assign \new_[7184]_  = A233 & ~A203;
  assign \new_[7187]_  = A301 & A234;
  assign \new_[7188]_  = \new_[7187]_  & \new_[7184]_ ;
  assign \new_[7192]_  = ~A202 & ~A201;
  assign \new_[7193]_  = A169 & \new_[7192]_ ;
  assign \new_[7196]_  = A233 & ~A203;
  assign \new_[7199]_  = A268 & A234;
  assign \new_[7200]_  = \new_[7199]_  & \new_[7196]_ ;
  assign \new_[7204]_  = A200 & A199;
  assign \new_[7205]_  = A169 & \new_[7204]_ ;
  assign \new_[7208]_  = ~A202 & ~A201;
  assign \new_[7211]_  = A301 & A235;
  assign \new_[7212]_  = \new_[7211]_  & \new_[7208]_ ;
  assign \new_[7216]_  = A200 & A199;
  assign \new_[7217]_  = A169 & \new_[7216]_ ;
  assign \new_[7220]_  = ~A202 & ~A201;
  assign \new_[7223]_  = A268 & A235;
  assign \new_[7224]_  = \new_[7223]_  & \new_[7220]_ ;
  assign \new_[7228]_  = ~A200 & ~A199;
  assign \new_[7229]_  = A169 & \new_[7228]_ ;
  assign \new_[7232]_  = A235 & ~A202;
  assign \new_[7235]_  = A300 & A299;
  assign \new_[7236]_  = \new_[7235]_  & \new_[7232]_ ;
  assign \new_[7240]_  = ~A200 & ~A199;
  assign \new_[7241]_  = A169 & \new_[7240]_ ;
  assign \new_[7244]_  = A235 & ~A202;
  assign \new_[7247]_  = A300 & A298;
  assign \new_[7248]_  = \new_[7247]_  & \new_[7244]_ ;
  assign \new_[7252]_  = ~A200 & ~A199;
  assign \new_[7253]_  = A169 & \new_[7252]_ ;
  assign \new_[7256]_  = A235 & ~A202;
  assign \new_[7259]_  = A267 & A265;
  assign \new_[7260]_  = \new_[7259]_  & \new_[7256]_ ;
  assign \new_[7264]_  = ~A200 & ~A199;
  assign \new_[7265]_  = A169 & \new_[7264]_ ;
  assign \new_[7268]_  = A235 & ~A202;
  assign \new_[7271]_  = A267 & A266;
  assign \new_[7272]_  = \new_[7271]_  & \new_[7268]_ ;
  assign \new_[7276]_  = ~A200 & ~A199;
  assign \new_[7277]_  = A169 & \new_[7276]_ ;
  assign \new_[7280]_  = A232 & ~A202;
  assign \new_[7283]_  = A301 & A234;
  assign \new_[7284]_  = \new_[7283]_  & \new_[7280]_ ;
  assign \new_[7288]_  = ~A200 & ~A199;
  assign \new_[7289]_  = A169 & \new_[7288]_ ;
  assign \new_[7292]_  = A232 & ~A202;
  assign \new_[7295]_  = A268 & A234;
  assign \new_[7296]_  = \new_[7295]_  & \new_[7292]_ ;
  assign \new_[7300]_  = ~A200 & ~A199;
  assign \new_[7301]_  = A169 & \new_[7300]_ ;
  assign \new_[7304]_  = A233 & ~A202;
  assign \new_[7307]_  = A301 & A234;
  assign \new_[7308]_  = \new_[7307]_  & \new_[7304]_ ;
  assign \new_[7312]_  = ~A200 & ~A199;
  assign \new_[7313]_  = A169 & \new_[7312]_ ;
  assign \new_[7316]_  = A233 & ~A202;
  assign \new_[7319]_  = A268 & A234;
  assign \new_[7320]_  = \new_[7319]_  & \new_[7316]_ ;
  assign \new_[7324]_  = ~A166 & ~A167;
  assign \new_[7325]_  = ~A169 & \new_[7324]_ ;
  assign \new_[7328]_  = A235 & A202;
  assign \new_[7331]_  = A300 & A299;
  assign \new_[7332]_  = \new_[7331]_  & \new_[7328]_ ;
  assign \new_[7336]_  = ~A166 & ~A167;
  assign \new_[7337]_  = ~A169 & \new_[7336]_ ;
  assign \new_[7340]_  = A235 & A202;
  assign \new_[7343]_  = A300 & A298;
  assign \new_[7344]_  = \new_[7343]_  & \new_[7340]_ ;
  assign \new_[7348]_  = ~A166 & ~A167;
  assign \new_[7349]_  = ~A169 & \new_[7348]_ ;
  assign \new_[7352]_  = A235 & A202;
  assign \new_[7355]_  = A267 & A265;
  assign \new_[7356]_  = \new_[7355]_  & \new_[7352]_ ;
  assign \new_[7360]_  = ~A166 & ~A167;
  assign \new_[7361]_  = ~A169 & \new_[7360]_ ;
  assign \new_[7364]_  = A235 & A202;
  assign \new_[7367]_  = A267 & A266;
  assign \new_[7368]_  = \new_[7367]_  & \new_[7364]_ ;
  assign \new_[7372]_  = ~A166 & ~A167;
  assign \new_[7373]_  = ~A169 & \new_[7372]_ ;
  assign \new_[7376]_  = A232 & A202;
  assign \new_[7379]_  = A301 & A234;
  assign \new_[7380]_  = \new_[7379]_  & \new_[7376]_ ;
  assign \new_[7384]_  = ~A166 & ~A167;
  assign \new_[7385]_  = ~A169 & \new_[7384]_ ;
  assign \new_[7388]_  = A232 & A202;
  assign \new_[7391]_  = A268 & A234;
  assign \new_[7392]_  = \new_[7391]_  & \new_[7388]_ ;
  assign \new_[7396]_  = ~A166 & ~A167;
  assign \new_[7397]_  = ~A169 & \new_[7396]_ ;
  assign \new_[7400]_  = A233 & A202;
  assign \new_[7403]_  = A301 & A234;
  assign \new_[7404]_  = \new_[7403]_  & \new_[7400]_ ;
  assign \new_[7408]_  = ~A166 & ~A167;
  assign \new_[7409]_  = ~A169 & \new_[7408]_ ;
  assign \new_[7412]_  = A233 & A202;
  assign \new_[7415]_  = A268 & A234;
  assign \new_[7416]_  = \new_[7415]_  & \new_[7412]_ ;
  assign \new_[7420]_  = ~A166 & ~A167;
  assign \new_[7421]_  = ~A169 & \new_[7420]_ ;
  assign \new_[7424]_  = A201 & A199;
  assign \new_[7427]_  = A301 & A235;
  assign \new_[7428]_  = \new_[7427]_  & \new_[7424]_ ;
  assign \new_[7432]_  = ~A166 & ~A167;
  assign \new_[7433]_  = ~A169 & \new_[7432]_ ;
  assign \new_[7436]_  = A201 & A199;
  assign \new_[7439]_  = A268 & A235;
  assign \new_[7440]_  = \new_[7439]_  & \new_[7436]_ ;
  assign \new_[7444]_  = ~A166 & ~A167;
  assign \new_[7445]_  = ~A169 & \new_[7444]_ ;
  assign \new_[7448]_  = A201 & A200;
  assign \new_[7451]_  = A301 & A235;
  assign \new_[7452]_  = \new_[7451]_  & \new_[7448]_ ;
  assign \new_[7456]_  = ~A166 & ~A167;
  assign \new_[7457]_  = ~A169 & \new_[7456]_ ;
  assign \new_[7460]_  = A201 & A200;
  assign \new_[7463]_  = A268 & A235;
  assign \new_[7464]_  = \new_[7463]_  & \new_[7460]_ ;
  assign \new_[7468]_  = A167 & ~A168;
  assign \new_[7469]_  = ~A169 & \new_[7468]_ ;
  assign \new_[7472]_  = A202 & A166;
  assign \new_[7475]_  = A301 & A235;
  assign \new_[7476]_  = \new_[7475]_  & \new_[7472]_ ;
  assign \new_[7480]_  = A167 & ~A168;
  assign \new_[7481]_  = ~A169 & \new_[7480]_ ;
  assign \new_[7484]_  = A202 & A166;
  assign \new_[7487]_  = A268 & A235;
  assign \new_[7488]_  = \new_[7487]_  & \new_[7484]_ ;
  assign \new_[7492]_  = ~A168 & ~A169;
  assign \new_[7493]_  = ~A170 & \new_[7492]_ ;
  assign \new_[7496]_  = A235 & A202;
  assign \new_[7499]_  = A300 & A299;
  assign \new_[7500]_  = \new_[7499]_  & \new_[7496]_ ;
  assign \new_[7504]_  = ~A168 & ~A169;
  assign \new_[7505]_  = ~A170 & \new_[7504]_ ;
  assign \new_[7508]_  = A235 & A202;
  assign \new_[7511]_  = A300 & A298;
  assign \new_[7512]_  = \new_[7511]_  & \new_[7508]_ ;
  assign \new_[7516]_  = ~A168 & ~A169;
  assign \new_[7517]_  = ~A170 & \new_[7516]_ ;
  assign \new_[7520]_  = A235 & A202;
  assign \new_[7523]_  = A267 & A265;
  assign \new_[7524]_  = \new_[7523]_  & \new_[7520]_ ;
  assign \new_[7528]_  = ~A168 & ~A169;
  assign \new_[7529]_  = ~A170 & \new_[7528]_ ;
  assign \new_[7532]_  = A235 & A202;
  assign \new_[7535]_  = A267 & A266;
  assign \new_[7536]_  = \new_[7535]_  & \new_[7532]_ ;
  assign \new_[7540]_  = ~A168 & ~A169;
  assign \new_[7541]_  = ~A170 & \new_[7540]_ ;
  assign \new_[7544]_  = A232 & A202;
  assign \new_[7547]_  = A301 & A234;
  assign \new_[7548]_  = \new_[7547]_  & \new_[7544]_ ;
  assign \new_[7552]_  = ~A168 & ~A169;
  assign \new_[7553]_  = ~A170 & \new_[7552]_ ;
  assign \new_[7556]_  = A232 & A202;
  assign \new_[7559]_  = A268 & A234;
  assign \new_[7560]_  = \new_[7559]_  & \new_[7556]_ ;
  assign \new_[7564]_  = ~A168 & ~A169;
  assign \new_[7565]_  = ~A170 & \new_[7564]_ ;
  assign \new_[7568]_  = A233 & A202;
  assign \new_[7571]_  = A301 & A234;
  assign \new_[7572]_  = \new_[7571]_  & \new_[7568]_ ;
  assign \new_[7576]_  = ~A168 & ~A169;
  assign \new_[7577]_  = ~A170 & \new_[7576]_ ;
  assign \new_[7580]_  = A233 & A202;
  assign \new_[7583]_  = A268 & A234;
  assign \new_[7584]_  = \new_[7583]_  & \new_[7580]_ ;
  assign \new_[7588]_  = ~A168 & ~A169;
  assign \new_[7589]_  = ~A170 & \new_[7588]_ ;
  assign \new_[7592]_  = A201 & A199;
  assign \new_[7595]_  = A301 & A235;
  assign \new_[7596]_  = \new_[7595]_  & \new_[7592]_ ;
  assign \new_[7600]_  = ~A168 & ~A169;
  assign \new_[7601]_  = ~A170 & \new_[7600]_ ;
  assign \new_[7604]_  = A201 & A199;
  assign \new_[7607]_  = A268 & A235;
  assign \new_[7608]_  = \new_[7607]_  & \new_[7604]_ ;
  assign \new_[7612]_  = ~A168 & ~A169;
  assign \new_[7613]_  = ~A170 & \new_[7612]_ ;
  assign \new_[7616]_  = A201 & A200;
  assign \new_[7619]_  = A301 & A235;
  assign \new_[7620]_  = \new_[7619]_  & \new_[7616]_ ;
  assign \new_[7624]_  = ~A168 & ~A169;
  assign \new_[7625]_  = ~A170 & \new_[7624]_ ;
  assign \new_[7628]_  = A201 & A200;
  assign \new_[7631]_  = A268 & A235;
  assign \new_[7632]_  = \new_[7631]_  & \new_[7628]_ ;
  assign \new_[7635]_  = A166 & A168;
  assign \new_[7638]_  = ~A202 & ~A201;
  assign \new_[7639]_  = \new_[7638]_  & \new_[7635]_ ;
  assign \new_[7642]_  = A235 & ~A203;
  assign \new_[7645]_  = A300 & A299;
  assign \new_[7646]_  = \new_[7645]_  & \new_[7642]_ ;
  assign \new_[7649]_  = A166 & A168;
  assign \new_[7652]_  = ~A202 & ~A201;
  assign \new_[7653]_  = \new_[7652]_  & \new_[7649]_ ;
  assign \new_[7656]_  = A235 & ~A203;
  assign \new_[7659]_  = A300 & A298;
  assign \new_[7660]_  = \new_[7659]_  & \new_[7656]_ ;
  assign \new_[7663]_  = A166 & A168;
  assign \new_[7666]_  = ~A202 & ~A201;
  assign \new_[7667]_  = \new_[7666]_  & \new_[7663]_ ;
  assign \new_[7670]_  = A235 & ~A203;
  assign \new_[7673]_  = A267 & A265;
  assign \new_[7674]_  = \new_[7673]_  & \new_[7670]_ ;
  assign \new_[7677]_  = A166 & A168;
  assign \new_[7680]_  = ~A202 & ~A201;
  assign \new_[7681]_  = \new_[7680]_  & \new_[7677]_ ;
  assign \new_[7684]_  = A235 & ~A203;
  assign \new_[7687]_  = A267 & A266;
  assign \new_[7688]_  = \new_[7687]_  & \new_[7684]_ ;
  assign \new_[7691]_  = A166 & A168;
  assign \new_[7694]_  = ~A202 & ~A201;
  assign \new_[7695]_  = \new_[7694]_  & \new_[7691]_ ;
  assign \new_[7698]_  = A232 & ~A203;
  assign \new_[7701]_  = A301 & A234;
  assign \new_[7702]_  = \new_[7701]_  & \new_[7698]_ ;
  assign \new_[7705]_  = A166 & A168;
  assign \new_[7708]_  = ~A202 & ~A201;
  assign \new_[7709]_  = \new_[7708]_  & \new_[7705]_ ;
  assign \new_[7712]_  = A232 & ~A203;
  assign \new_[7715]_  = A268 & A234;
  assign \new_[7716]_  = \new_[7715]_  & \new_[7712]_ ;
  assign \new_[7719]_  = A166 & A168;
  assign \new_[7722]_  = ~A202 & ~A201;
  assign \new_[7723]_  = \new_[7722]_  & \new_[7719]_ ;
  assign \new_[7726]_  = A233 & ~A203;
  assign \new_[7729]_  = A301 & A234;
  assign \new_[7730]_  = \new_[7729]_  & \new_[7726]_ ;
  assign \new_[7733]_  = A166 & A168;
  assign \new_[7736]_  = ~A202 & ~A201;
  assign \new_[7737]_  = \new_[7736]_  & \new_[7733]_ ;
  assign \new_[7740]_  = A233 & ~A203;
  assign \new_[7743]_  = A268 & A234;
  assign \new_[7744]_  = \new_[7743]_  & \new_[7740]_ ;
  assign \new_[7747]_  = A166 & A168;
  assign \new_[7750]_  = A200 & A199;
  assign \new_[7751]_  = \new_[7750]_  & \new_[7747]_ ;
  assign \new_[7754]_  = ~A202 & ~A201;
  assign \new_[7757]_  = A301 & A235;
  assign \new_[7758]_  = \new_[7757]_  & \new_[7754]_ ;
  assign \new_[7761]_  = A166 & A168;
  assign \new_[7764]_  = A200 & A199;
  assign \new_[7765]_  = \new_[7764]_  & \new_[7761]_ ;
  assign \new_[7768]_  = ~A202 & ~A201;
  assign \new_[7771]_  = A268 & A235;
  assign \new_[7772]_  = \new_[7771]_  & \new_[7768]_ ;
  assign \new_[7775]_  = A166 & A168;
  assign \new_[7778]_  = ~A200 & ~A199;
  assign \new_[7779]_  = \new_[7778]_  & \new_[7775]_ ;
  assign \new_[7782]_  = A235 & ~A202;
  assign \new_[7785]_  = A300 & A299;
  assign \new_[7786]_  = \new_[7785]_  & \new_[7782]_ ;
  assign \new_[7789]_  = A166 & A168;
  assign \new_[7792]_  = ~A200 & ~A199;
  assign \new_[7793]_  = \new_[7792]_  & \new_[7789]_ ;
  assign \new_[7796]_  = A235 & ~A202;
  assign \new_[7799]_  = A300 & A298;
  assign \new_[7800]_  = \new_[7799]_  & \new_[7796]_ ;
  assign \new_[7803]_  = A166 & A168;
  assign \new_[7806]_  = ~A200 & ~A199;
  assign \new_[7807]_  = \new_[7806]_  & \new_[7803]_ ;
  assign \new_[7810]_  = A235 & ~A202;
  assign \new_[7813]_  = A267 & A265;
  assign \new_[7814]_  = \new_[7813]_  & \new_[7810]_ ;
  assign \new_[7817]_  = A166 & A168;
  assign \new_[7820]_  = ~A200 & ~A199;
  assign \new_[7821]_  = \new_[7820]_  & \new_[7817]_ ;
  assign \new_[7824]_  = A235 & ~A202;
  assign \new_[7827]_  = A267 & A266;
  assign \new_[7828]_  = \new_[7827]_  & \new_[7824]_ ;
  assign \new_[7831]_  = A166 & A168;
  assign \new_[7834]_  = ~A200 & ~A199;
  assign \new_[7835]_  = \new_[7834]_  & \new_[7831]_ ;
  assign \new_[7838]_  = A232 & ~A202;
  assign \new_[7841]_  = A301 & A234;
  assign \new_[7842]_  = \new_[7841]_  & \new_[7838]_ ;
  assign \new_[7845]_  = A166 & A168;
  assign \new_[7848]_  = ~A200 & ~A199;
  assign \new_[7849]_  = \new_[7848]_  & \new_[7845]_ ;
  assign \new_[7852]_  = A232 & ~A202;
  assign \new_[7855]_  = A268 & A234;
  assign \new_[7856]_  = \new_[7855]_  & \new_[7852]_ ;
  assign \new_[7859]_  = A166 & A168;
  assign \new_[7862]_  = ~A200 & ~A199;
  assign \new_[7863]_  = \new_[7862]_  & \new_[7859]_ ;
  assign \new_[7866]_  = A233 & ~A202;
  assign \new_[7869]_  = A301 & A234;
  assign \new_[7870]_  = \new_[7869]_  & \new_[7866]_ ;
  assign \new_[7873]_  = A166 & A168;
  assign \new_[7876]_  = ~A200 & ~A199;
  assign \new_[7877]_  = \new_[7876]_  & \new_[7873]_ ;
  assign \new_[7880]_  = A233 & ~A202;
  assign \new_[7883]_  = A268 & A234;
  assign \new_[7884]_  = \new_[7883]_  & \new_[7880]_ ;
  assign \new_[7887]_  = A167 & A168;
  assign \new_[7890]_  = ~A202 & ~A201;
  assign \new_[7891]_  = \new_[7890]_  & \new_[7887]_ ;
  assign \new_[7894]_  = A235 & ~A203;
  assign \new_[7897]_  = A300 & A299;
  assign \new_[7898]_  = \new_[7897]_  & \new_[7894]_ ;
  assign \new_[7901]_  = A167 & A168;
  assign \new_[7904]_  = ~A202 & ~A201;
  assign \new_[7905]_  = \new_[7904]_  & \new_[7901]_ ;
  assign \new_[7908]_  = A235 & ~A203;
  assign \new_[7911]_  = A300 & A298;
  assign \new_[7912]_  = \new_[7911]_  & \new_[7908]_ ;
  assign \new_[7915]_  = A167 & A168;
  assign \new_[7918]_  = ~A202 & ~A201;
  assign \new_[7919]_  = \new_[7918]_  & \new_[7915]_ ;
  assign \new_[7922]_  = A235 & ~A203;
  assign \new_[7925]_  = A267 & A265;
  assign \new_[7926]_  = \new_[7925]_  & \new_[7922]_ ;
  assign \new_[7929]_  = A167 & A168;
  assign \new_[7932]_  = ~A202 & ~A201;
  assign \new_[7933]_  = \new_[7932]_  & \new_[7929]_ ;
  assign \new_[7936]_  = A235 & ~A203;
  assign \new_[7939]_  = A267 & A266;
  assign \new_[7940]_  = \new_[7939]_  & \new_[7936]_ ;
  assign \new_[7943]_  = A167 & A168;
  assign \new_[7946]_  = ~A202 & ~A201;
  assign \new_[7947]_  = \new_[7946]_  & \new_[7943]_ ;
  assign \new_[7950]_  = A232 & ~A203;
  assign \new_[7953]_  = A301 & A234;
  assign \new_[7954]_  = \new_[7953]_  & \new_[7950]_ ;
  assign \new_[7957]_  = A167 & A168;
  assign \new_[7960]_  = ~A202 & ~A201;
  assign \new_[7961]_  = \new_[7960]_  & \new_[7957]_ ;
  assign \new_[7964]_  = A232 & ~A203;
  assign \new_[7967]_  = A268 & A234;
  assign \new_[7968]_  = \new_[7967]_  & \new_[7964]_ ;
  assign \new_[7971]_  = A167 & A168;
  assign \new_[7974]_  = ~A202 & ~A201;
  assign \new_[7975]_  = \new_[7974]_  & \new_[7971]_ ;
  assign \new_[7978]_  = A233 & ~A203;
  assign \new_[7981]_  = A301 & A234;
  assign \new_[7982]_  = \new_[7981]_  & \new_[7978]_ ;
  assign \new_[7985]_  = A167 & A168;
  assign \new_[7988]_  = ~A202 & ~A201;
  assign \new_[7989]_  = \new_[7988]_  & \new_[7985]_ ;
  assign \new_[7992]_  = A233 & ~A203;
  assign \new_[7995]_  = A268 & A234;
  assign \new_[7996]_  = \new_[7995]_  & \new_[7992]_ ;
  assign \new_[7999]_  = A167 & A168;
  assign \new_[8002]_  = A200 & A199;
  assign \new_[8003]_  = \new_[8002]_  & \new_[7999]_ ;
  assign \new_[8006]_  = ~A202 & ~A201;
  assign \new_[8009]_  = A301 & A235;
  assign \new_[8010]_  = \new_[8009]_  & \new_[8006]_ ;
  assign \new_[8013]_  = A167 & A168;
  assign \new_[8016]_  = A200 & A199;
  assign \new_[8017]_  = \new_[8016]_  & \new_[8013]_ ;
  assign \new_[8020]_  = ~A202 & ~A201;
  assign \new_[8023]_  = A268 & A235;
  assign \new_[8024]_  = \new_[8023]_  & \new_[8020]_ ;
  assign \new_[8027]_  = A167 & A168;
  assign \new_[8030]_  = ~A200 & ~A199;
  assign \new_[8031]_  = \new_[8030]_  & \new_[8027]_ ;
  assign \new_[8034]_  = A235 & ~A202;
  assign \new_[8037]_  = A300 & A299;
  assign \new_[8038]_  = \new_[8037]_  & \new_[8034]_ ;
  assign \new_[8041]_  = A167 & A168;
  assign \new_[8044]_  = ~A200 & ~A199;
  assign \new_[8045]_  = \new_[8044]_  & \new_[8041]_ ;
  assign \new_[8048]_  = A235 & ~A202;
  assign \new_[8051]_  = A300 & A298;
  assign \new_[8052]_  = \new_[8051]_  & \new_[8048]_ ;
  assign \new_[8055]_  = A167 & A168;
  assign \new_[8058]_  = ~A200 & ~A199;
  assign \new_[8059]_  = \new_[8058]_  & \new_[8055]_ ;
  assign \new_[8062]_  = A235 & ~A202;
  assign \new_[8065]_  = A267 & A265;
  assign \new_[8066]_  = \new_[8065]_  & \new_[8062]_ ;
  assign \new_[8069]_  = A167 & A168;
  assign \new_[8072]_  = ~A200 & ~A199;
  assign \new_[8073]_  = \new_[8072]_  & \new_[8069]_ ;
  assign \new_[8076]_  = A235 & ~A202;
  assign \new_[8079]_  = A267 & A266;
  assign \new_[8080]_  = \new_[8079]_  & \new_[8076]_ ;
  assign \new_[8083]_  = A167 & A168;
  assign \new_[8086]_  = ~A200 & ~A199;
  assign \new_[8087]_  = \new_[8086]_  & \new_[8083]_ ;
  assign \new_[8090]_  = A232 & ~A202;
  assign \new_[8093]_  = A301 & A234;
  assign \new_[8094]_  = \new_[8093]_  & \new_[8090]_ ;
  assign \new_[8097]_  = A167 & A168;
  assign \new_[8100]_  = ~A200 & ~A199;
  assign \new_[8101]_  = \new_[8100]_  & \new_[8097]_ ;
  assign \new_[8104]_  = A232 & ~A202;
  assign \new_[8107]_  = A268 & A234;
  assign \new_[8108]_  = \new_[8107]_  & \new_[8104]_ ;
  assign \new_[8111]_  = A167 & A168;
  assign \new_[8114]_  = ~A200 & ~A199;
  assign \new_[8115]_  = \new_[8114]_  & \new_[8111]_ ;
  assign \new_[8118]_  = A233 & ~A202;
  assign \new_[8121]_  = A301 & A234;
  assign \new_[8122]_  = \new_[8121]_  & \new_[8118]_ ;
  assign \new_[8125]_  = A167 & A168;
  assign \new_[8128]_  = ~A200 & ~A199;
  assign \new_[8129]_  = \new_[8128]_  & \new_[8125]_ ;
  assign \new_[8132]_  = A233 & ~A202;
  assign \new_[8135]_  = A268 & A234;
  assign \new_[8136]_  = \new_[8135]_  & \new_[8132]_ ;
  assign \new_[8139]_  = A167 & A170;
  assign \new_[8142]_  = ~A201 & ~A166;
  assign \new_[8143]_  = \new_[8142]_  & \new_[8139]_ ;
  assign \new_[8146]_  = ~A203 & ~A202;
  assign \new_[8149]_  = A301 & A235;
  assign \new_[8150]_  = \new_[8149]_  & \new_[8146]_ ;
  assign \new_[8153]_  = A167 & A170;
  assign \new_[8156]_  = ~A201 & ~A166;
  assign \new_[8157]_  = \new_[8156]_  & \new_[8153]_ ;
  assign \new_[8160]_  = ~A203 & ~A202;
  assign \new_[8163]_  = A268 & A235;
  assign \new_[8164]_  = \new_[8163]_  & \new_[8160]_ ;
  assign \new_[8167]_  = A167 & A170;
  assign \new_[8170]_  = ~A199 & ~A166;
  assign \new_[8171]_  = \new_[8170]_  & \new_[8167]_ ;
  assign \new_[8174]_  = ~A202 & ~A200;
  assign \new_[8177]_  = A301 & A235;
  assign \new_[8178]_  = \new_[8177]_  & \new_[8174]_ ;
  assign \new_[8181]_  = A167 & A170;
  assign \new_[8184]_  = ~A199 & ~A166;
  assign \new_[8185]_  = \new_[8184]_  & \new_[8181]_ ;
  assign \new_[8188]_  = ~A202 & ~A200;
  assign \new_[8191]_  = A268 & A235;
  assign \new_[8192]_  = \new_[8191]_  & \new_[8188]_ ;
  assign \new_[8195]_  = ~A167 & A170;
  assign \new_[8198]_  = ~A201 & A166;
  assign \new_[8199]_  = \new_[8198]_  & \new_[8195]_ ;
  assign \new_[8202]_  = ~A203 & ~A202;
  assign \new_[8205]_  = A301 & A235;
  assign \new_[8206]_  = \new_[8205]_  & \new_[8202]_ ;
  assign \new_[8209]_  = ~A167 & A170;
  assign \new_[8212]_  = ~A201 & A166;
  assign \new_[8213]_  = \new_[8212]_  & \new_[8209]_ ;
  assign \new_[8216]_  = ~A203 & ~A202;
  assign \new_[8219]_  = A268 & A235;
  assign \new_[8220]_  = \new_[8219]_  & \new_[8216]_ ;
  assign \new_[8223]_  = ~A167 & A170;
  assign \new_[8226]_  = ~A199 & A166;
  assign \new_[8227]_  = \new_[8226]_  & \new_[8223]_ ;
  assign \new_[8230]_  = ~A202 & ~A200;
  assign \new_[8233]_  = A301 & A235;
  assign \new_[8234]_  = \new_[8233]_  & \new_[8230]_ ;
  assign \new_[8237]_  = ~A167 & A170;
  assign \new_[8240]_  = ~A199 & A166;
  assign \new_[8241]_  = \new_[8240]_  & \new_[8237]_ ;
  assign \new_[8244]_  = ~A202 & ~A200;
  assign \new_[8247]_  = A268 & A235;
  assign \new_[8248]_  = \new_[8247]_  & \new_[8244]_ ;
  assign \new_[8251]_  = ~A201 & A169;
  assign \new_[8254]_  = ~A203 & ~A202;
  assign \new_[8255]_  = \new_[8254]_  & \new_[8251]_ ;
  assign \new_[8258]_  = A298 & A235;
  assign \new_[8261]_  = A302 & ~A299;
  assign \new_[8262]_  = \new_[8261]_  & \new_[8258]_ ;
  assign \new_[8265]_  = ~A201 & A169;
  assign \new_[8268]_  = ~A203 & ~A202;
  assign \new_[8269]_  = \new_[8268]_  & \new_[8265]_ ;
  assign \new_[8272]_  = ~A298 & A235;
  assign \new_[8275]_  = A302 & A299;
  assign \new_[8276]_  = \new_[8275]_  & \new_[8272]_ ;
  assign \new_[8279]_  = ~A201 & A169;
  assign \new_[8282]_  = ~A203 & ~A202;
  assign \new_[8283]_  = \new_[8282]_  & \new_[8279]_ ;
  assign \new_[8286]_  = ~A265 & A235;
  assign \new_[8289]_  = A269 & A266;
  assign \new_[8290]_  = \new_[8289]_  & \new_[8286]_ ;
  assign \new_[8293]_  = ~A201 & A169;
  assign \new_[8296]_  = ~A203 & ~A202;
  assign \new_[8297]_  = \new_[8296]_  & \new_[8293]_ ;
  assign \new_[8300]_  = A265 & A235;
  assign \new_[8303]_  = A269 & ~A266;
  assign \new_[8304]_  = \new_[8303]_  & \new_[8300]_ ;
  assign \new_[8307]_  = ~A201 & A169;
  assign \new_[8310]_  = ~A203 & ~A202;
  assign \new_[8311]_  = \new_[8310]_  & \new_[8307]_ ;
  assign \new_[8314]_  = A234 & A232;
  assign \new_[8317]_  = A300 & A299;
  assign \new_[8318]_  = \new_[8317]_  & \new_[8314]_ ;
  assign \new_[8321]_  = ~A201 & A169;
  assign \new_[8324]_  = ~A203 & ~A202;
  assign \new_[8325]_  = \new_[8324]_  & \new_[8321]_ ;
  assign \new_[8328]_  = A234 & A232;
  assign \new_[8331]_  = A300 & A298;
  assign \new_[8332]_  = \new_[8331]_  & \new_[8328]_ ;
  assign \new_[8335]_  = ~A201 & A169;
  assign \new_[8338]_  = ~A203 & ~A202;
  assign \new_[8339]_  = \new_[8338]_  & \new_[8335]_ ;
  assign \new_[8342]_  = A234 & A232;
  assign \new_[8345]_  = A267 & A265;
  assign \new_[8346]_  = \new_[8345]_  & \new_[8342]_ ;
  assign \new_[8349]_  = ~A201 & A169;
  assign \new_[8352]_  = ~A203 & ~A202;
  assign \new_[8353]_  = \new_[8352]_  & \new_[8349]_ ;
  assign \new_[8356]_  = A234 & A232;
  assign \new_[8359]_  = A267 & A266;
  assign \new_[8360]_  = \new_[8359]_  & \new_[8356]_ ;
  assign \new_[8363]_  = ~A201 & A169;
  assign \new_[8366]_  = ~A203 & ~A202;
  assign \new_[8367]_  = \new_[8366]_  & \new_[8363]_ ;
  assign \new_[8370]_  = A234 & A233;
  assign \new_[8373]_  = A300 & A299;
  assign \new_[8374]_  = \new_[8373]_  & \new_[8370]_ ;
  assign \new_[8377]_  = ~A201 & A169;
  assign \new_[8380]_  = ~A203 & ~A202;
  assign \new_[8381]_  = \new_[8380]_  & \new_[8377]_ ;
  assign \new_[8384]_  = A234 & A233;
  assign \new_[8387]_  = A300 & A298;
  assign \new_[8388]_  = \new_[8387]_  & \new_[8384]_ ;
  assign \new_[8391]_  = ~A201 & A169;
  assign \new_[8394]_  = ~A203 & ~A202;
  assign \new_[8395]_  = \new_[8394]_  & \new_[8391]_ ;
  assign \new_[8398]_  = A234 & A233;
  assign \new_[8401]_  = A267 & A265;
  assign \new_[8402]_  = \new_[8401]_  & \new_[8398]_ ;
  assign \new_[8405]_  = ~A201 & A169;
  assign \new_[8408]_  = ~A203 & ~A202;
  assign \new_[8409]_  = \new_[8408]_  & \new_[8405]_ ;
  assign \new_[8412]_  = A234 & A233;
  assign \new_[8415]_  = A267 & A266;
  assign \new_[8416]_  = \new_[8415]_  & \new_[8412]_ ;
  assign \new_[8419]_  = ~A201 & A169;
  assign \new_[8422]_  = ~A203 & ~A202;
  assign \new_[8423]_  = \new_[8422]_  & \new_[8419]_ ;
  assign \new_[8426]_  = A233 & ~A232;
  assign \new_[8429]_  = A301 & A236;
  assign \new_[8430]_  = \new_[8429]_  & \new_[8426]_ ;
  assign \new_[8433]_  = ~A201 & A169;
  assign \new_[8436]_  = ~A203 & ~A202;
  assign \new_[8437]_  = \new_[8436]_  & \new_[8433]_ ;
  assign \new_[8440]_  = A233 & ~A232;
  assign \new_[8443]_  = A268 & A236;
  assign \new_[8444]_  = \new_[8443]_  & \new_[8440]_ ;
  assign \new_[8447]_  = ~A201 & A169;
  assign \new_[8450]_  = ~A203 & ~A202;
  assign \new_[8451]_  = \new_[8450]_  & \new_[8447]_ ;
  assign \new_[8454]_  = ~A233 & A232;
  assign \new_[8457]_  = A301 & A236;
  assign \new_[8458]_  = \new_[8457]_  & \new_[8454]_ ;
  assign \new_[8461]_  = ~A201 & A169;
  assign \new_[8464]_  = ~A203 & ~A202;
  assign \new_[8465]_  = \new_[8464]_  & \new_[8461]_ ;
  assign \new_[8468]_  = ~A233 & A232;
  assign \new_[8471]_  = A268 & A236;
  assign \new_[8472]_  = \new_[8471]_  & \new_[8468]_ ;
  assign \new_[8475]_  = A199 & A169;
  assign \new_[8478]_  = ~A201 & A200;
  assign \new_[8479]_  = \new_[8478]_  & \new_[8475]_ ;
  assign \new_[8482]_  = A235 & ~A202;
  assign \new_[8485]_  = A300 & A299;
  assign \new_[8486]_  = \new_[8485]_  & \new_[8482]_ ;
  assign \new_[8489]_  = A199 & A169;
  assign \new_[8492]_  = ~A201 & A200;
  assign \new_[8493]_  = \new_[8492]_  & \new_[8489]_ ;
  assign \new_[8496]_  = A235 & ~A202;
  assign \new_[8499]_  = A300 & A298;
  assign \new_[8500]_  = \new_[8499]_  & \new_[8496]_ ;
  assign \new_[8503]_  = A199 & A169;
  assign \new_[8506]_  = ~A201 & A200;
  assign \new_[8507]_  = \new_[8506]_  & \new_[8503]_ ;
  assign \new_[8510]_  = A235 & ~A202;
  assign \new_[8513]_  = A267 & A265;
  assign \new_[8514]_  = \new_[8513]_  & \new_[8510]_ ;
  assign \new_[8517]_  = A199 & A169;
  assign \new_[8520]_  = ~A201 & A200;
  assign \new_[8521]_  = \new_[8520]_  & \new_[8517]_ ;
  assign \new_[8524]_  = A235 & ~A202;
  assign \new_[8527]_  = A267 & A266;
  assign \new_[8528]_  = \new_[8527]_  & \new_[8524]_ ;
  assign \new_[8531]_  = A199 & A169;
  assign \new_[8534]_  = ~A201 & A200;
  assign \new_[8535]_  = \new_[8534]_  & \new_[8531]_ ;
  assign \new_[8538]_  = A232 & ~A202;
  assign \new_[8541]_  = A301 & A234;
  assign \new_[8542]_  = \new_[8541]_  & \new_[8538]_ ;
  assign \new_[8545]_  = A199 & A169;
  assign \new_[8548]_  = ~A201 & A200;
  assign \new_[8549]_  = \new_[8548]_  & \new_[8545]_ ;
  assign \new_[8552]_  = A232 & ~A202;
  assign \new_[8555]_  = A268 & A234;
  assign \new_[8556]_  = \new_[8555]_  & \new_[8552]_ ;
  assign \new_[8559]_  = A199 & A169;
  assign \new_[8562]_  = ~A201 & A200;
  assign \new_[8563]_  = \new_[8562]_  & \new_[8559]_ ;
  assign \new_[8566]_  = A233 & ~A202;
  assign \new_[8569]_  = A301 & A234;
  assign \new_[8570]_  = \new_[8569]_  & \new_[8566]_ ;
  assign \new_[8573]_  = A199 & A169;
  assign \new_[8576]_  = ~A201 & A200;
  assign \new_[8577]_  = \new_[8576]_  & \new_[8573]_ ;
  assign \new_[8580]_  = A233 & ~A202;
  assign \new_[8583]_  = A268 & A234;
  assign \new_[8584]_  = \new_[8583]_  & \new_[8580]_ ;
  assign \new_[8587]_  = ~A199 & A169;
  assign \new_[8590]_  = ~A202 & ~A200;
  assign \new_[8591]_  = \new_[8590]_  & \new_[8587]_ ;
  assign \new_[8594]_  = A298 & A235;
  assign \new_[8597]_  = A302 & ~A299;
  assign \new_[8598]_  = \new_[8597]_  & \new_[8594]_ ;
  assign \new_[8601]_  = ~A199 & A169;
  assign \new_[8604]_  = ~A202 & ~A200;
  assign \new_[8605]_  = \new_[8604]_  & \new_[8601]_ ;
  assign \new_[8608]_  = ~A298 & A235;
  assign \new_[8611]_  = A302 & A299;
  assign \new_[8612]_  = \new_[8611]_  & \new_[8608]_ ;
  assign \new_[8615]_  = ~A199 & A169;
  assign \new_[8618]_  = ~A202 & ~A200;
  assign \new_[8619]_  = \new_[8618]_  & \new_[8615]_ ;
  assign \new_[8622]_  = ~A265 & A235;
  assign \new_[8625]_  = A269 & A266;
  assign \new_[8626]_  = \new_[8625]_  & \new_[8622]_ ;
  assign \new_[8629]_  = ~A199 & A169;
  assign \new_[8632]_  = ~A202 & ~A200;
  assign \new_[8633]_  = \new_[8632]_  & \new_[8629]_ ;
  assign \new_[8636]_  = A265 & A235;
  assign \new_[8639]_  = A269 & ~A266;
  assign \new_[8640]_  = \new_[8639]_  & \new_[8636]_ ;
  assign \new_[8643]_  = ~A199 & A169;
  assign \new_[8646]_  = ~A202 & ~A200;
  assign \new_[8647]_  = \new_[8646]_  & \new_[8643]_ ;
  assign \new_[8650]_  = A234 & A232;
  assign \new_[8653]_  = A300 & A299;
  assign \new_[8654]_  = \new_[8653]_  & \new_[8650]_ ;
  assign \new_[8657]_  = ~A199 & A169;
  assign \new_[8660]_  = ~A202 & ~A200;
  assign \new_[8661]_  = \new_[8660]_  & \new_[8657]_ ;
  assign \new_[8664]_  = A234 & A232;
  assign \new_[8667]_  = A300 & A298;
  assign \new_[8668]_  = \new_[8667]_  & \new_[8664]_ ;
  assign \new_[8671]_  = ~A199 & A169;
  assign \new_[8674]_  = ~A202 & ~A200;
  assign \new_[8675]_  = \new_[8674]_  & \new_[8671]_ ;
  assign \new_[8678]_  = A234 & A232;
  assign \new_[8681]_  = A267 & A265;
  assign \new_[8682]_  = \new_[8681]_  & \new_[8678]_ ;
  assign \new_[8685]_  = ~A199 & A169;
  assign \new_[8688]_  = ~A202 & ~A200;
  assign \new_[8689]_  = \new_[8688]_  & \new_[8685]_ ;
  assign \new_[8692]_  = A234 & A232;
  assign \new_[8695]_  = A267 & A266;
  assign \new_[8696]_  = \new_[8695]_  & \new_[8692]_ ;
  assign \new_[8699]_  = ~A199 & A169;
  assign \new_[8702]_  = ~A202 & ~A200;
  assign \new_[8703]_  = \new_[8702]_  & \new_[8699]_ ;
  assign \new_[8706]_  = A234 & A233;
  assign \new_[8709]_  = A300 & A299;
  assign \new_[8710]_  = \new_[8709]_  & \new_[8706]_ ;
  assign \new_[8713]_  = ~A199 & A169;
  assign \new_[8716]_  = ~A202 & ~A200;
  assign \new_[8717]_  = \new_[8716]_  & \new_[8713]_ ;
  assign \new_[8720]_  = A234 & A233;
  assign \new_[8723]_  = A300 & A298;
  assign \new_[8724]_  = \new_[8723]_  & \new_[8720]_ ;
  assign \new_[8727]_  = ~A199 & A169;
  assign \new_[8730]_  = ~A202 & ~A200;
  assign \new_[8731]_  = \new_[8730]_  & \new_[8727]_ ;
  assign \new_[8734]_  = A234 & A233;
  assign \new_[8737]_  = A267 & A265;
  assign \new_[8738]_  = \new_[8737]_  & \new_[8734]_ ;
  assign \new_[8741]_  = ~A199 & A169;
  assign \new_[8744]_  = ~A202 & ~A200;
  assign \new_[8745]_  = \new_[8744]_  & \new_[8741]_ ;
  assign \new_[8748]_  = A234 & A233;
  assign \new_[8751]_  = A267 & A266;
  assign \new_[8752]_  = \new_[8751]_  & \new_[8748]_ ;
  assign \new_[8755]_  = ~A199 & A169;
  assign \new_[8758]_  = ~A202 & ~A200;
  assign \new_[8759]_  = \new_[8758]_  & \new_[8755]_ ;
  assign \new_[8762]_  = A233 & ~A232;
  assign \new_[8765]_  = A301 & A236;
  assign \new_[8766]_  = \new_[8765]_  & \new_[8762]_ ;
  assign \new_[8769]_  = ~A199 & A169;
  assign \new_[8772]_  = ~A202 & ~A200;
  assign \new_[8773]_  = \new_[8772]_  & \new_[8769]_ ;
  assign \new_[8776]_  = A233 & ~A232;
  assign \new_[8779]_  = A268 & A236;
  assign \new_[8780]_  = \new_[8779]_  & \new_[8776]_ ;
  assign \new_[8783]_  = ~A199 & A169;
  assign \new_[8786]_  = ~A202 & ~A200;
  assign \new_[8787]_  = \new_[8786]_  & \new_[8783]_ ;
  assign \new_[8790]_  = ~A233 & A232;
  assign \new_[8793]_  = A301 & A236;
  assign \new_[8794]_  = \new_[8793]_  & \new_[8790]_ ;
  assign \new_[8797]_  = ~A199 & A169;
  assign \new_[8800]_  = ~A202 & ~A200;
  assign \new_[8801]_  = \new_[8800]_  & \new_[8797]_ ;
  assign \new_[8804]_  = ~A233 & A232;
  assign \new_[8807]_  = A268 & A236;
  assign \new_[8808]_  = \new_[8807]_  & \new_[8804]_ ;
  assign \new_[8811]_  = ~A167 & ~A169;
  assign \new_[8814]_  = A202 & ~A166;
  assign \new_[8815]_  = \new_[8814]_  & \new_[8811]_ ;
  assign \new_[8818]_  = A298 & A235;
  assign \new_[8821]_  = A302 & ~A299;
  assign \new_[8822]_  = \new_[8821]_  & \new_[8818]_ ;
  assign \new_[8825]_  = ~A167 & ~A169;
  assign \new_[8828]_  = A202 & ~A166;
  assign \new_[8829]_  = \new_[8828]_  & \new_[8825]_ ;
  assign \new_[8832]_  = ~A298 & A235;
  assign \new_[8835]_  = A302 & A299;
  assign \new_[8836]_  = \new_[8835]_  & \new_[8832]_ ;
  assign \new_[8839]_  = ~A167 & ~A169;
  assign \new_[8842]_  = A202 & ~A166;
  assign \new_[8843]_  = \new_[8842]_  & \new_[8839]_ ;
  assign \new_[8846]_  = ~A265 & A235;
  assign \new_[8849]_  = A269 & A266;
  assign \new_[8850]_  = \new_[8849]_  & \new_[8846]_ ;
  assign \new_[8853]_  = ~A167 & ~A169;
  assign \new_[8856]_  = A202 & ~A166;
  assign \new_[8857]_  = \new_[8856]_  & \new_[8853]_ ;
  assign \new_[8860]_  = A265 & A235;
  assign \new_[8863]_  = A269 & ~A266;
  assign \new_[8864]_  = \new_[8863]_  & \new_[8860]_ ;
  assign \new_[8867]_  = ~A167 & ~A169;
  assign \new_[8870]_  = A202 & ~A166;
  assign \new_[8871]_  = \new_[8870]_  & \new_[8867]_ ;
  assign \new_[8874]_  = A234 & A232;
  assign \new_[8877]_  = A300 & A299;
  assign \new_[8878]_  = \new_[8877]_  & \new_[8874]_ ;
  assign \new_[8881]_  = ~A167 & ~A169;
  assign \new_[8884]_  = A202 & ~A166;
  assign \new_[8885]_  = \new_[8884]_  & \new_[8881]_ ;
  assign \new_[8888]_  = A234 & A232;
  assign \new_[8891]_  = A300 & A298;
  assign \new_[8892]_  = \new_[8891]_  & \new_[8888]_ ;
  assign \new_[8895]_  = ~A167 & ~A169;
  assign \new_[8898]_  = A202 & ~A166;
  assign \new_[8899]_  = \new_[8898]_  & \new_[8895]_ ;
  assign \new_[8902]_  = A234 & A232;
  assign \new_[8905]_  = A267 & A265;
  assign \new_[8906]_  = \new_[8905]_  & \new_[8902]_ ;
  assign \new_[8909]_  = ~A167 & ~A169;
  assign \new_[8912]_  = A202 & ~A166;
  assign \new_[8913]_  = \new_[8912]_  & \new_[8909]_ ;
  assign \new_[8916]_  = A234 & A232;
  assign \new_[8919]_  = A267 & A266;
  assign \new_[8920]_  = \new_[8919]_  & \new_[8916]_ ;
  assign \new_[8923]_  = ~A167 & ~A169;
  assign \new_[8926]_  = A202 & ~A166;
  assign \new_[8927]_  = \new_[8926]_  & \new_[8923]_ ;
  assign \new_[8930]_  = A234 & A233;
  assign \new_[8933]_  = A300 & A299;
  assign \new_[8934]_  = \new_[8933]_  & \new_[8930]_ ;
  assign \new_[8937]_  = ~A167 & ~A169;
  assign \new_[8940]_  = A202 & ~A166;
  assign \new_[8941]_  = \new_[8940]_  & \new_[8937]_ ;
  assign \new_[8944]_  = A234 & A233;
  assign \new_[8947]_  = A300 & A298;
  assign \new_[8948]_  = \new_[8947]_  & \new_[8944]_ ;
  assign \new_[8951]_  = ~A167 & ~A169;
  assign \new_[8954]_  = A202 & ~A166;
  assign \new_[8955]_  = \new_[8954]_  & \new_[8951]_ ;
  assign \new_[8958]_  = A234 & A233;
  assign \new_[8961]_  = A267 & A265;
  assign \new_[8962]_  = \new_[8961]_  & \new_[8958]_ ;
  assign \new_[8965]_  = ~A167 & ~A169;
  assign \new_[8968]_  = A202 & ~A166;
  assign \new_[8969]_  = \new_[8968]_  & \new_[8965]_ ;
  assign \new_[8972]_  = A234 & A233;
  assign \new_[8975]_  = A267 & A266;
  assign \new_[8976]_  = \new_[8975]_  & \new_[8972]_ ;
  assign \new_[8979]_  = ~A167 & ~A169;
  assign \new_[8982]_  = A202 & ~A166;
  assign \new_[8983]_  = \new_[8982]_  & \new_[8979]_ ;
  assign \new_[8986]_  = A233 & ~A232;
  assign \new_[8989]_  = A301 & A236;
  assign \new_[8990]_  = \new_[8989]_  & \new_[8986]_ ;
  assign \new_[8993]_  = ~A167 & ~A169;
  assign \new_[8996]_  = A202 & ~A166;
  assign \new_[8997]_  = \new_[8996]_  & \new_[8993]_ ;
  assign \new_[9000]_  = A233 & ~A232;
  assign \new_[9003]_  = A268 & A236;
  assign \new_[9004]_  = \new_[9003]_  & \new_[9000]_ ;
  assign \new_[9007]_  = ~A167 & ~A169;
  assign \new_[9010]_  = A202 & ~A166;
  assign \new_[9011]_  = \new_[9010]_  & \new_[9007]_ ;
  assign \new_[9014]_  = ~A233 & A232;
  assign \new_[9017]_  = A301 & A236;
  assign \new_[9018]_  = \new_[9017]_  & \new_[9014]_ ;
  assign \new_[9021]_  = ~A167 & ~A169;
  assign \new_[9024]_  = A202 & ~A166;
  assign \new_[9025]_  = \new_[9024]_  & \new_[9021]_ ;
  assign \new_[9028]_  = ~A233 & A232;
  assign \new_[9031]_  = A268 & A236;
  assign \new_[9032]_  = \new_[9031]_  & \new_[9028]_ ;
  assign \new_[9035]_  = ~A167 & ~A169;
  assign \new_[9038]_  = A199 & ~A166;
  assign \new_[9039]_  = \new_[9038]_  & \new_[9035]_ ;
  assign \new_[9042]_  = A235 & A201;
  assign \new_[9045]_  = A300 & A299;
  assign \new_[9046]_  = \new_[9045]_  & \new_[9042]_ ;
  assign \new_[9049]_  = ~A167 & ~A169;
  assign \new_[9052]_  = A199 & ~A166;
  assign \new_[9053]_  = \new_[9052]_  & \new_[9049]_ ;
  assign \new_[9056]_  = A235 & A201;
  assign \new_[9059]_  = A300 & A298;
  assign \new_[9060]_  = \new_[9059]_  & \new_[9056]_ ;
  assign \new_[9063]_  = ~A167 & ~A169;
  assign \new_[9066]_  = A199 & ~A166;
  assign \new_[9067]_  = \new_[9066]_  & \new_[9063]_ ;
  assign \new_[9070]_  = A235 & A201;
  assign \new_[9073]_  = A267 & A265;
  assign \new_[9074]_  = \new_[9073]_  & \new_[9070]_ ;
  assign \new_[9077]_  = ~A167 & ~A169;
  assign \new_[9080]_  = A199 & ~A166;
  assign \new_[9081]_  = \new_[9080]_  & \new_[9077]_ ;
  assign \new_[9084]_  = A235 & A201;
  assign \new_[9087]_  = A267 & A266;
  assign \new_[9088]_  = \new_[9087]_  & \new_[9084]_ ;
  assign \new_[9091]_  = ~A167 & ~A169;
  assign \new_[9094]_  = A199 & ~A166;
  assign \new_[9095]_  = \new_[9094]_  & \new_[9091]_ ;
  assign \new_[9098]_  = A232 & A201;
  assign \new_[9101]_  = A301 & A234;
  assign \new_[9102]_  = \new_[9101]_  & \new_[9098]_ ;
  assign \new_[9105]_  = ~A167 & ~A169;
  assign \new_[9108]_  = A199 & ~A166;
  assign \new_[9109]_  = \new_[9108]_  & \new_[9105]_ ;
  assign \new_[9112]_  = A232 & A201;
  assign \new_[9115]_  = A268 & A234;
  assign \new_[9116]_  = \new_[9115]_  & \new_[9112]_ ;
  assign \new_[9119]_  = ~A167 & ~A169;
  assign \new_[9122]_  = A199 & ~A166;
  assign \new_[9123]_  = \new_[9122]_  & \new_[9119]_ ;
  assign \new_[9126]_  = A233 & A201;
  assign \new_[9129]_  = A301 & A234;
  assign \new_[9130]_  = \new_[9129]_  & \new_[9126]_ ;
  assign \new_[9133]_  = ~A167 & ~A169;
  assign \new_[9136]_  = A199 & ~A166;
  assign \new_[9137]_  = \new_[9136]_  & \new_[9133]_ ;
  assign \new_[9140]_  = A233 & A201;
  assign \new_[9143]_  = A268 & A234;
  assign \new_[9144]_  = \new_[9143]_  & \new_[9140]_ ;
  assign \new_[9147]_  = ~A167 & ~A169;
  assign \new_[9150]_  = A200 & ~A166;
  assign \new_[9151]_  = \new_[9150]_  & \new_[9147]_ ;
  assign \new_[9154]_  = A235 & A201;
  assign \new_[9157]_  = A300 & A299;
  assign \new_[9158]_  = \new_[9157]_  & \new_[9154]_ ;
  assign \new_[9161]_  = ~A167 & ~A169;
  assign \new_[9164]_  = A200 & ~A166;
  assign \new_[9165]_  = \new_[9164]_  & \new_[9161]_ ;
  assign \new_[9168]_  = A235 & A201;
  assign \new_[9171]_  = A300 & A298;
  assign \new_[9172]_  = \new_[9171]_  & \new_[9168]_ ;
  assign \new_[9175]_  = ~A167 & ~A169;
  assign \new_[9178]_  = A200 & ~A166;
  assign \new_[9179]_  = \new_[9178]_  & \new_[9175]_ ;
  assign \new_[9182]_  = A235 & A201;
  assign \new_[9185]_  = A267 & A265;
  assign \new_[9186]_  = \new_[9185]_  & \new_[9182]_ ;
  assign \new_[9189]_  = ~A167 & ~A169;
  assign \new_[9192]_  = A200 & ~A166;
  assign \new_[9193]_  = \new_[9192]_  & \new_[9189]_ ;
  assign \new_[9196]_  = A235 & A201;
  assign \new_[9199]_  = A267 & A266;
  assign \new_[9200]_  = \new_[9199]_  & \new_[9196]_ ;
  assign \new_[9203]_  = ~A167 & ~A169;
  assign \new_[9206]_  = A200 & ~A166;
  assign \new_[9207]_  = \new_[9206]_  & \new_[9203]_ ;
  assign \new_[9210]_  = A232 & A201;
  assign \new_[9213]_  = A301 & A234;
  assign \new_[9214]_  = \new_[9213]_  & \new_[9210]_ ;
  assign \new_[9217]_  = ~A167 & ~A169;
  assign \new_[9220]_  = A200 & ~A166;
  assign \new_[9221]_  = \new_[9220]_  & \new_[9217]_ ;
  assign \new_[9224]_  = A232 & A201;
  assign \new_[9227]_  = A268 & A234;
  assign \new_[9228]_  = \new_[9227]_  & \new_[9224]_ ;
  assign \new_[9231]_  = ~A167 & ~A169;
  assign \new_[9234]_  = A200 & ~A166;
  assign \new_[9235]_  = \new_[9234]_  & \new_[9231]_ ;
  assign \new_[9238]_  = A233 & A201;
  assign \new_[9241]_  = A301 & A234;
  assign \new_[9242]_  = \new_[9241]_  & \new_[9238]_ ;
  assign \new_[9245]_  = ~A167 & ~A169;
  assign \new_[9248]_  = A200 & ~A166;
  assign \new_[9249]_  = \new_[9248]_  & \new_[9245]_ ;
  assign \new_[9252]_  = A233 & A201;
  assign \new_[9255]_  = A268 & A234;
  assign \new_[9256]_  = \new_[9255]_  & \new_[9252]_ ;
  assign \new_[9259]_  = ~A167 & ~A169;
  assign \new_[9262]_  = ~A199 & ~A166;
  assign \new_[9263]_  = \new_[9262]_  & \new_[9259]_ ;
  assign \new_[9266]_  = A203 & A200;
  assign \new_[9269]_  = A301 & A235;
  assign \new_[9270]_  = \new_[9269]_  & \new_[9266]_ ;
  assign \new_[9273]_  = ~A167 & ~A169;
  assign \new_[9276]_  = ~A199 & ~A166;
  assign \new_[9277]_  = \new_[9276]_  & \new_[9273]_ ;
  assign \new_[9280]_  = A203 & A200;
  assign \new_[9283]_  = A268 & A235;
  assign \new_[9284]_  = \new_[9283]_  & \new_[9280]_ ;
  assign \new_[9287]_  = ~A167 & ~A169;
  assign \new_[9290]_  = A199 & ~A166;
  assign \new_[9291]_  = \new_[9290]_  & \new_[9287]_ ;
  assign \new_[9294]_  = A203 & ~A200;
  assign \new_[9297]_  = A301 & A235;
  assign \new_[9298]_  = \new_[9297]_  & \new_[9294]_ ;
  assign \new_[9301]_  = ~A167 & ~A169;
  assign \new_[9304]_  = A199 & ~A166;
  assign \new_[9305]_  = \new_[9304]_  & \new_[9301]_ ;
  assign \new_[9308]_  = A203 & ~A200;
  assign \new_[9311]_  = A268 & A235;
  assign \new_[9312]_  = \new_[9311]_  & \new_[9308]_ ;
  assign \new_[9315]_  = ~A168 & ~A169;
  assign \new_[9318]_  = A166 & A167;
  assign \new_[9319]_  = \new_[9318]_  & \new_[9315]_ ;
  assign \new_[9322]_  = A235 & A202;
  assign \new_[9325]_  = A300 & A299;
  assign \new_[9326]_  = \new_[9325]_  & \new_[9322]_ ;
  assign \new_[9329]_  = ~A168 & ~A169;
  assign \new_[9332]_  = A166 & A167;
  assign \new_[9333]_  = \new_[9332]_  & \new_[9329]_ ;
  assign \new_[9336]_  = A235 & A202;
  assign \new_[9339]_  = A300 & A298;
  assign \new_[9340]_  = \new_[9339]_  & \new_[9336]_ ;
  assign \new_[9343]_  = ~A168 & ~A169;
  assign \new_[9346]_  = A166 & A167;
  assign \new_[9347]_  = \new_[9346]_  & \new_[9343]_ ;
  assign \new_[9350]_  = A235 & A202;
  assign \new_[9353]_  = A267 & A265;
  assign \new_[9354]_  = \new_[9353]_  & \new_[9350]_ ;
  assign \new_[9357]_  = ~A168 & ~A169;
  assign \new_[9360]_  = A166 & A167;
  assign \new_[9361]_  = \new_[9360]_  & \new_[9357]_ ;
  assign \new_[9364]_  = A235 & A202;
  assign \new_[9367]_  = A267 & A266;
  assign \new_[9368]_  = \new_[9367]_  & \new_[9364]_ ;
  assign \new_[9371]_  = ~A168 & ~A169;
  assign \new_[9374]_  = A166 & A167;
  assign \new_[9375]_  = \new_[9374]_  & \new_[9371]_ ;
  assign \new_[9378]_  = A232 & A202;
  assign \new_[9381]_  = A301 & A234;
  assign \new_[9382]_  = \new_[9381]_  & \new_[9378]_ ;
  assign \new_[9385]_  = ~A168 & ~A169;
  assign \new_[9388]_  = A166 & A167;
  assign \new_[9389]_  = \new_[9388]_  & \new_[9385]_ ;
  assign \new_[9392]_  = A232 & A202;
  assign \new_[9395]_  = A268 & A234;
  assign \new_[9396]_  = \new_[9395]_  & \new_[9392]_ ;
  assign \new_[9399]_  = ~A168 & ~A169;
  assign \new_[9402]_  = A166 & A167;
  assign \new_[9403]_  = \new_[9402]_  & \new_[9399]_ ;
  assign \new_[9406]_  = A233 & A202;
  assign \new_[9409]_  = A301 & A234;
  assign \new_[9410]_  = \new_[9409]_  & \new_[9406]_ ;
  assign \new_[9413]_  = ~A168 & ~A169;
  assign \new_[9416]_  = A166 & A167;
  assign \new_[9417]_  = \new_[9416]_  & \new_[9413]_ ;
  assign \new_[9420]_  = A233 & A202;
  assign \new_[9423]_  = A268 & A234;
  assign \new_[9424]_  = \new_[9423]_  & \new_[9420]_ ;
  assign \new_[9427]_  = ~A168 & ~A169;
  assign \new_[9430]_  = A166 & A167;
  assign \new_[9431]_  = \new_[9430]_  & \new_[9427]_ ;
  assign \new_[9434]_  = A201 & A199;
  assign \new_[9437]_  = A301 & A235;
  assign \new_[9438]_  = \new_[9437]_  & \new_[9434]_ ;
  assign \new_[9441]_  = ~A168 & ~A169;
  assign \new_[9444]_  = A166 & A167;
  assign \new_[9445]_  = \new_[9444]_  & \new_[9441]_ ;
  assign \new_[9448]_  = A201 & A199;
  assign \new_[9451]_  = A268 & A235;
  assign \new_[9452]_  = \new_[9451]_  & \new_[9448]_ ;
  assign \new_[9455]_  = ~A168 & ~A169;
  assign \new_[9458]_  = A166 & A167;
  assign \new_[9459]_  = \new_[9458]_  & \new_[9455]_ ;
  assign \new_[9462]_  = A201 & A200;
  assign \new_[9465]_  = A301 & A235;
  assign \new_[9466]_  = \new_[9465]_  & \new_[9462]_ ;
  assign \new_[9469]_  = ~A168 & ~A169;
  assign \new_[9472]_  = A166 & A167;
  assign \new_[9473]_  = \new_[9472]_  & \new_[9469]_ ;
  assign \new_[9476]_  = A201 & A200;
  assign \new_[9479]_  = A268 & A235;
  assign \new_[9480]_  = \new_[9479]_  & \new_[9476]_ ;
  assign \new_[9483]_  = ~A169 & ~A170;
  assign \new_[9486]_  = A202 & ~A168;
  assign \new_[9487]_  = \new_[9486]_  & \new_[9483]_ ;
  assign \new_[9490]_  = A298 & A235;
  assign \new_[9493]_  = A302 & ~A299;
  assign \new_[9494]_  = \new_[9493]_  & \new_[9490]_ ;
  assign \new_[9497]_  = ~A169 & ~A170;
  assign \new_[9500]_  = A202 & ~A168;
  assign \new_[9501]_  = \new_[9500]_  & \new_[9497]_ ;
  assign \new_[9504]_  = ~A298 & A235;
  assign \new_[9507]_  = A302 & A299;
  assign \new_[9508]_  = \new_[9507]_  & \new_[9504]_ ;
  assign \new_[9511]_  = ~A169 & ~A170;
  assign \new_[9514]_  = A202 & ~A168;
  assign \new_[9515]_  = \new_[9514]_  & \new_[9511]_ ;
  assign \new_[9518]_  = ~A265 & A235;
  assign \new_[9521]_  = A269 & A266;
  assign \new_[9522]_  = \new_[9521]_  & \new_[9518]_ ;
  assign \new_[9525]_  = ~A169 & ~A170;
  assign \new_[9528]_  = A202 & ~A168;
  assign \new_[9529]_  = \new_[9528]_  & \new_[9525]_ ;
  assign \new_[9532]_  = A265 & A235;
  assign \new_[9535]_  = A269 & ~A266;
  assign \new_[9536]_  = \new_[9535]_  & \new_[9532]_ ;
  assign \new_[9539]_  = ~A169 & ~A170;
  assign \new_[9542]_  = A202 & ~A168;
  assign \new_[9543]_  = \new_[9542]_  & \new_[9539]_ ;
  assign \new_[9546]_  = A234 & A232;
  assign \new_[9549]_  = A300 & A299;
  assign \new_[9550]_  = \new_[9549]_  & \new_[9546]_ ;
  assign \new_[9553]_  = ~A169 & ~A170;
  assign \new_[9556]_  = A202 & ~A168;
  assign \new_[9557]_  = \new_[9556]_  & \new_[9553]_ ;
  assign \new_[9560]_  = A234 & A232;
  assign \new_[9563]_  = A300 & A298;
  assign \new_[9564]_  = \new_[9563]_  & \new_[9560]_ ;
  assign \new_[9567]_  = ~A169 & ~A170;
  assign \new_[9570]_  = A202 & ~A168;
  assign \new_[9571]_  = \new_[9570]_  & \new_[9567]_ ;
  assign \new_[9574]_  = A234 & A232;
  assign \new_[9577]_  = A267 & A265;
  assign \new_[9578]_  = \new_[9577]_  & \new_[9574]_ ;
  assign \new_[9581]_  = ~A169 & ~A170;
  assign \new_[9584]_  = A202 & ~A168;
  assign \new_[9585]_  = \new_[9584]_  & \new_[9581]_ ;
  assign \new_[9588]_  = A234 & A232;
  assign \new_[9591]_  = A267 & A266;
  assign \new_[9592]_  = \new_[9591]_  & \new_[9588]_ ;
  assign \new_[9595]_  = ~A169 & ~A170;
  assign \new_[9598]_  = A202 & ~A168;
  assign \new_[9599]_  = \new_[9598]_  & \new_[9595]_ ;
  assign \new_[9602]_  = A234 & A233;
  assign \new_[9605]_  = A300 & A299;
  assign \new_[9606]_  = \new_[9605]_  & \new_[9602]_ ;
  assign \new_[9609]_  = ~A169 & ~A170;
  assign \new_[9612]_  = A202 & ~A168;
  assign \new_[9613]_  = \new_[9612]_  & \new_[9609]_ ;
  assign \new_[9616]_  = A234 & A233;
  assign \new_[9619]_  = A300 & A298;
  assign \new_[9620]_  = \new_[9619]_  & \new_[9616]_ ;
  assign \new_[9623]_  = ~A169 & ~A170;
  assign \new_[9626]_  = A202 & ~A168;
  assign \new_[9627]_  = \new_[9626]_  & \new_[9623]_ ;
  assign \new_[9630]_  = A234 & A233;
  assign \new_[9633]_  = A267 & A265;
  assign \new_[9634]_  = \new_[9633]_  & \new_[9630]_ ;
  assign \new_[9637]_  = ~A169 & ~A170;
  assign \new_[9640]_  = A202 & ~A168;
  assign \new_[9641]_  = \new_[9640]_  & \new_[9637]_ ;
  assign \new_[9644]_  = A234 & A233;
  assign \new_[9647]_  = A267 & A266;
  assign \new_[9648]_  = \new_[9647]_  & \new_[9644]_ ;
  assign \new_[9651]_  = ~A169 & ~A170;
  assign \new_[9654]_  = A202 & ~A168;
  assign \new_[9655]_  = \new_[9654]_  & \new_[9651]_ ;
  assign \new_[9658]_  = A233 & ~A232;
  assign \new_[9661]_  = A301 & A236;
  assign \new_[9662]_  = \new_[9661]_  & \new_[9658]_ ;
  assign \new_[9665]_  = ~A169 & ~A170;
  assign \new_[9668]_  = A202 & ~A168;
  assign \new_[9669]_  = \new_[9668]_  & \new_[9665]_ ;
  assign \new_[9672]_  = A233 & ~A232;
  assign \new_[9675]_  = A268 & A236;
  assign \new_[9676]_  = \new_[9675]_  & \new_[9672]_ ;
  assign \new_[9679]_  = ~A169 & ~A170;
  assign \new_[9682]_  = A202 & ~A168;
  assign \new_[9683]_  = \new_[9682]_  & \new_[9679]_ ;
  assign \new_[9686]_  = ~A233 & A232;
  assign \new_[9689]_  = A301 & A236;
  assign \new_[9690]_  = \new_[9689]_  & \new_[9686]_ ;
  assign \new_[9693]_  = ~A169 & ~A170;
  assign \new_[9696]_  = A202 & ~A168;
  assign \new_[9697]_  = \new_[9696]_  & \new_[9693]_ ;
  assign \new_[9700]_  = ~A233 & A232;
  assign \new_[9703]_  = A268 & A236;
  assign \new_[9704]_  = \new_[9703]_  & \new_[9700]_ ;
  assign \new_[9707]_  = ~A169 & ~A170;
  assign \new_[9710]_  = A199 & ~A168;
  assign \new_[9711]_  = \new_[9710]_  & \new_[9707]_ ;
  assign \new_[9714]_  = A235 & A201;
  assign \new_[9717]_  = A300 & A299;
  assign \new_[9718]_  = \new_[9717]_  & \new_[9714]_ ;
  assign \new_[9721]_  = ~A169 & ~A170;
  assign \new_[9724]_  = A199 & ~A168;
  assign \new_[9725]_  = \new_[9724]_  & \new_[9721]_ ;
  assign \new_[9728]_  = A235 & A201;
  assign \new_[9731]_  = A300 & A298;
  assign \new_[9732]_  = \new_[9731]_  & \new_[9728]_ ;
  assign \new_[9735]_  = ~A169 & ~A170;
  assign \new_[9738]_  = A199 & ~A168;
  assign \new_[9739]_  = \new_[9738]_  & \new_[9735]_ ;
  assign \new_[9742]_  = A235 & A201;
  assign \new_[9745]_  = A267 & A265;
  assign \new_[9746]_  = \new_[9745]_  & \new_[9742]_ ;
  assign \new_[9749]_  = ~A169 & ~A170;
  assign \new_[9752]_  = A199 & ~A168;
  assign \new_[9753]_  = \new_[9752]_  & \new_[9749]_ ;
  assign \new_[9756]_  = A235 & A201;
  assign \new_[9759]_  = A267 & A266;
  assign \new_[9760]_  = \new_[9759]_  & \new_[9756]_ ;
  assign \new_[9763]_  = ~A169 & ~A170;
  assign \new_[9766]_  = A199 & ~A168;
  assign \new_[9767]_  = \new_[9766]_  & \new_[9763]_ ;
  assign \new_[9770]_  = A232 & A201;
  assign \new_[9773]_  = A301 & A234;
  assign \new_[9774]_  = \new_[9773]_  & \new_[9770]_ ;
  assign \new_[9777]_  = ~A169 & ~A170;
  assign \new_[9780]_  = A199 & ~A168;
  assign \new_[9781]_  = \new_[9780]_  & \new_[9777]_ ;
  assign \new_[9784]_  = A232 & A201;
  assign \new_[9787]_  = A268 & A234;
  assign \new_[9788]_  = \new_[9787]_  & \new_[9784]_ ;
  assign \new_[9791]_  = ~A169 & ~A170;
  assign \new_[9794]_  = A199 & ~A168;
  assign \new_[9795]_  = \new_[9794]_  & \new_[9791]_ ;
  assign \new_[9798]_  = A233 & A201;
  assign \new_[9801]_  = A301 & A234;
  assign \new_[9802]_  = \new_[9801]_  & \new_[9798]_ ;
  assign \new_[9805]_  = ~A169 & ~A170;
  assign \new_[9808]_  = A199 & ~A168;
  assign \new_[9809]_  = \new_[9808]_  & \new_[9805]_ ;
  assign \new_[9812]_  = A233 & A201;
  assign \new_[9815]_  = A268 & A234;
  assign \new_[9816]_  = \new_[9815]_  & \new_[9812]_ ;
  assign \new_[9819]_  = ~A169 & ~A170;
  assign \new_[9822]_  = A200 & ~A168;
  assign \new_[9823]_  = \new_[9822]_  & \new_[9819]_ ;
  assign \new_[9826]_  = A235 & A201;
  assign \new_[9829]_  = A300 & A299;
  assign \new_[9830]_  = \new_[9829]_  & \new_[9826]_ ;
  assign \new_[9833]_  = ~A169 & ~A170;
  assign \new_[9836]_  = A200 & ~A168;
  assign \new_[9837]_  = \new_[9836]_  & \new_[9833]_ ;
  assign \new_[9840]_  = A235 & A201;
  assign \new_[9843]_  = A300 & A298;
  assign \new_[9844]_  = \new_[9843]_  & \new_[9840]_ ;
  assign \new_[9847]_  = ~A169 & ~A170;
  assign \new_[9850]_  = A200 & ~A168;
  assign \new_[9851]_  = \new_[9850]_  & \new_[9847]_ ;
  assign \new_[9854]_  = A235 & A201;
  assign \new_[9857]_  = A267 & A265;
  assign \new_[9858]_  = \new_[9857]_  & \new_[9854]_ ;
  assign \new_[9861]_  = ~A169 & ~A170;
  assign \new_[9864]_  = A200 & ~A168;
  assign \new_[9865]_  = \new_[9864]_  & \new_[9861]_ ;
  assign \new_[9868]_  = A235 & A201;
  assign \new_[9871]_  = A267 & A266;
  assign \new_[9872]_  = \new_[9871]_  & \new_[9868]_ ;
  assign \new_[9875]_  = ~A169 & ~A170;
  assign \new_[9878]_  = A200 & ~A168;
  assign \new_[9879]_  = \new_[9878]_  & \new_[9875]_ ;
  assign \new_[9882]_  = A232 & A201;
  assign \new_[9885]_  = A301 & A234;
  assign \new_[9886]_  = \new_[9885]_  & \new_[9882]_ ;
  assign \new_[9889]_  = ~A169 & ~A170;
  assign \new_[9892]_  = A200 & ~A168;
  assign \new_[9893]_  = \new_[9892]_  & \new_[9889]_ ;
  assign \new_[9896]_  = A232 & A201;
  assign \new_[9899]_  = A268 & A234;
  assign \new_[9900]_  = \new_[9899]_  & \new_[9896]_ ;
  assign \new_[9903]_  = ~A169 & ~A170;
  assign \new_[9906]_  = A200 & ~A168;
  assign \new_[9907]_  = \new_[9906]_  & \new_[9903]_ ;
  assign \new_[9910]_  = A233 & A201;
  assign \new_[9913]_  = A301 & A234;
  assign \new_[9914]_  = \new_[9913]_  & \new_[9910]_ ;
  assign \new_[9917]_  = ~A169 & ~A170;
  assign \new_[9920]_  = A200 & ~A168;
  assign \new_[9921]_  = \new_[9920]_  & \new_[9917]_ ;
  assign \new_[9924]_  = A233 & A201;
  assign \new_[9927]_  = A268 & A234;
  assign \new_[9928]_  = \new_[9927]_  & \new_[9924]_ ;
  assign \new_[9931]_  = ~A169 & ~A170;
  assign \new_[9934]_  = ~A199 & ~A168;
  assign \new_[9935]_  = \new_[9934]_  & \new_[9931]_ ;
  assign \new_[9938]_  = A203 & A200;
  assign \new_[9941]_  = A301 & A235;
  assign \new_[9942]_  = \new_[9941]_  & \new_[9938]_ ;
  assign \new_[9945]_  = ~A169 & ~A170;
  assign \new_[9948]_  = ~A199 & ~A168;
  assign \new_[9949]_  = \new_[9948]_  & \new_[9945]_ ;
  assign \new_[9952]_  = A203 & A200;
  assign \new_[9955]_  = A268 & A235;
  assign \new_[9956]_  = \new_[9955]_  & \new_[9952]_ ;
  assign \new_[9959]_  = ~A169 & ~A170;
  assign \new_[9962]_  = A199 & ~A168;
  assign \new_[9963]_  = \new_[9962]_  & \new_[9959]_ ;
  assign \new_[9966]_  = A203 & ~A200;
  assign \new_[9969]_  = A301 & A235;
  assign \new_[9970]_  = \new_[9969]_  & \new_[9966]_ ;
  assign \new_[9973]_  = ~A169 & ~A170;
  assign \new_[9976]_  = A199 & ~A168;
  assign \new_[9977]_  = \new_[9976]_  & \new_[9973]_ ;
  assign \new_[9980]_  = A203 & ~A200;
  assign \new_[9983]_  = A268 & A235;
  assign \new_[9984]_  = \new_[9983]_  & \new_[9980]_ ;
  assign \new_[9987]_  = A166 & A168;
  assign \new_[9990]_  = ~A202 & ~A201;
  assign \new_[9991]_  = \new_[9990]_  & \new_[9987]_ ;
  assign \new_[9994]_  = A235 & ~A203;
  assign \new_[9998]_  = A302 & ~A299;
  assign \new_[9999]_  = A298 & \new_[9998]_ ;
  assign \new_[10000]_  = \new_[9999]_  & \new_[9994]_ ;
  assign \new_[10003]_  = A166 & A168;
  assign \new_[10006]_  = ~A202 & ~A201;
  assign \new_[10007]_  = \new_[10006]_  & \new_[10003]_ ;
  assign \new_[10010]_  = A235 & ~A203;
  assign \new_[10014]_  = A302 & A299;
  assign \new_[10015]_  = ~A298 & \new_[10014]_ ;
  assign \new_[10016]_  = \new_[10015]_  & \new_[10010]_ ;
  assign \new_[10019]_  = A166 & A168;
  assign \new_[10022]_  = ~A202 & ~A201;
  assign \new_[10023]_  = \new_[10022]_  & \new_[10019]_ ;
  assign \new_[10026]_  = A235 & ~A203;
  assign \new_[10030]_  = A269 & A266;
  assign \new_[10031]_  = ~A265 & \new_[10030]_ ;
  assign \new_[10032]_  = \new_[10031]_  & \new_[10026]_ ;
  assign \new_[10035]_  = A166 & A168;
  assign \new_[10038]_  = ~A202 & ~A201;
  assign \new_[10039]_  = \new_[10038]_  & \new_[10035]_ ;
  assign \new_[10042]_  = A235 & ~A203;
  assign \new_[10046]_  = A269 & ~A266;
  assign \new_[10047]_  = A265 & \new_[10046]_ ;
  assign \new_[10048]_  = \new_[10047]_  & \new_[10042]_ ;
  assign \new_[10051]_  = A166 & A168;
  assign \new_[10054]_  = ~A202 & ~A201;
  assign \new_[10055]_  = \new_[10054]_  & \new_[10051]_ ;
  assign \new_[10058]_  = A232 & ~A203;
  assign \new_[10062]_  = A300 & A299;
  assign \new_[10063]_  = A234 & \new_[10062]_ ;
  assign \new_[10064]_  = \new_[10063]_  & \new_[10058]_ ;
  assign \new_[10067]_  = A166 & A168;
  assign \new_[10070]_  = ~A202 & ~A201;
  assign \new_[10071]_  = \new_[10070]_  & \new_[10067]_ ;
  assign \new_[10074]_  = A232 & ~A203;
  assign \new_[10078]_  = A300 & A298;
  assign \new_[10079]_  = A234 & \new_[10078]_ ;
  assign \new_[10080]_  = \new_[10079]_  & \new_[10074]_ ;
  assign \new_[10083]_  = A166 & A168;
  assign \new_[10086]_  = ~A202 & ~A201;
  assign \new_[10087]_  = \new_[10086]_  & \new_[10083]_ ;
  assign \new_[10090]_  = A232 & ~A203;
  assign \new_[10094]_  = A267 & A265;
  assign \new_[10095]_  = A234 & \new_[10094]_ ;
  assign \new_[10096]_  = \new_[10095]_  & \new_[10090]_ ;
  assign \new_[10099]_  = A166 & A168;
  assign \new_[10102]_  = ~A202 & ~A201;
  assign \new_[10103]_  = \new_[10102]_  & \new_[10099]_ ;
  assign \new_[10106]_  = A232 & ~A203;
  assign \new_[10110]_  = A267 & A266;
  assign \new_[10111]_  = A234 & \new_[10110]_ ;
  assign \new_[10112]_  = \new_[10111]_  & \new_[10106]_ ;
  assign \new_[10115]_  = A166 & A168;
  assign \new_[10118]_  = ~A202 & ~A201;
  assign \new_[10119]_  = \new_[10118]_  & \new_[10115]_ ;
  assign \new_[10122]_  = A233 & ~A203;
  assign \new_[10126]_  = A300 & A299;
  assign \new_[10127]_  = A234 & \new_[10126]_ ;
  assign \new_[10128]_  = \new_[10127]_  & \new_[10122]_ ;
  assign \new_[10131]_  = A166 & A168;
  assign \new_[10134]_  = ~A202 & ~A201;
  assign \new_[10135]_  = \new_[10134]_  & \new_[10131]_ ;
  assign \new_[10138]_  = A233 & ~A203;
  assign \new_[10142]_  = A300 & A298;
  assign \new_[10143]_  = A234 & \new_[10142]_ ;
  assign \new_[10144]_  = \new_[10143]_  & \new_[10138]_ ;
  assign \new_[10147]_  = A166 & A168;
  assign \new_[10150]_  = ~A202 & ~A201;
  assign \new_[10151]_  = \new_[10150]_  & \new_[10147]_ ;
  assign \new_[10154]_  = A233 & ~A203;
  assign \new_[10158]_  = A267 & A265;
  assign \new_[10159]_  = A234 & \new_[10158]_ ;
  assign \new_[10160]_  = \new_[10159]_  & \new_[10154]_ ;
  assign \new_[10163]_  = A166 & A168;
  assign \new_[10166]_  = ~A202 & ~A201;
  assign \new_[10167]_  = \new_[10166]_  & \new_[10163]_ ;
  assign \new_[10170]_  = A233 & ~A203;
  assign \new_[10174]_  = A267 & A266;
  assign \new_[10175]_  = A234 & \new_[10174]_ ;
  assign \new_[10176]_  = \new_[10175]_  & \new_[10170]_ ;
  assign \new_[10179]_  = A166 & A168;
  assign \new_[10182]_  = ~A202 & ~A201;
  assign \new_[10183]_  = \new_[10182]_  & \new_[10179]_ ;
  assign \new_[10186]_  = ~A232 & ~A203;
  assign \new_[10190]_  = A301 & A236;
  assign \new_[10191]_  = A233 & \new_[10190]_ ;
  assign \new_[10192]_  = \new_[10191]_  & \new_[10186]_ ;
  assign \new_[10195]_  = A166 & A168;
  assign \new_[10198]_  = ~A202 & ~A201;
  assign \new_[10199]_  = \new_[10198]_  & \new_[10195]_ ;
  assign \new_[10202]_  = ~A232 & ~A203;
  assign \new_[10206]_  = A268 & A236;
  assign \new_[10207]_  = A233 & \new_[10206]_ ;
  assign \new_[10208]_  = \new_[10207]_  & \new_[10202]_ ;
  assign \new_[10211]_  = A166 & A168;
  assign \new_[10214]_  = ~A202 & ~A201;
  assign \new_[10215]_  = \new_[10214]_  & \new_[10211]_ ;
  assign \new_[10218]_  = A232 & ~A203;
  assign \new_[10222]_  = A301 & A236;
  assign \new_[10223]_  = ~A233 & \new_[10222]_ ;
  assign \new_[10224]_  = \new_[10223]_  & \new_[10218]_ ;
  assign \new_[10227]_  = A166 & A168;
  assign \new_[10230]_  = ~A202 & ~A201;
  assign \new_[10231]_  = \new_[10230]_  & \new_[10227]_ ;
  assign \new_[10234]_  = A232 & ~A203;
  assign \new_[10238]_  = A268 & A236;
  assign \new_[10239]_  = ~A233 & \new_[10238]_ ;
  assign \new_[10240]_  = \new_[10239]_  & \new_[10234]_ ;
  assign \new_[10243]_  = A166 & A168;
  assign \new_[10246]_  = A200 & A199;
  assign \new_[10247]_  = \new_[10246]_  & \new_[10243]_ ;
  assign \new_[10250]_  = ~A202 & ~A201;
  assign \new_[10254]_  = A300 & A299;
  assign \new_[10255]_  = A235 & \new_[10254]_ ;
  assign \new_[10256]_  = \new_[10255]_  & \new_[10250]_ ;
  assign \new_[10259]_  = A166 & A168;
  assign \new_[10262]_  = A200 & A199;
  assign \new_[10263]_  = \new_[10262]_  & \new_[10259]_ ;
  assign \new_[10266]_  = ~A202 & ~A201;
  assign \new_[10270]_  = A300 & A298;
  assign \new_[10271]_  = A235 & \new_[10270]_ ;
  assign \new_[10272]_  = \new_[10271]_  & \new_[10266]_ ;
  assign \new_[10275]_  = A166 & A168;
  assign \new_[10278]_  = A200 & A199;
  assign \new_[10279]_  = \new_[10278]_  & \new_[10275]_ ;
  assign \new_[10282]_  = ~A202 & ~A201;
  assign \new_[10286]_  = A267 & A265;
  assign \new_[10287]_  = A235 & \new_[10286]_ ;
  assign \new_[10288]_  = \new_[10287]_  & \new_[10282]_ ;
  assign \new_[10291]_  = A166 & A168;
  assign \new_[10294]_  = A200 & A199;
  assign \new_[10295]_  = \new_[10294]_  & \new_[10291]_ ;
  assign \new_[10298]_  = ~A202 & ~A201;
  assign \new_[10302]_  = A267 & A266;
  assign \new_[10303]_  = A235 & \new_[10302]_ ;
  assign \new_[10304]_  = \new_[10303]_  & \new_[10298]_ ;
  assign \new_[10307]_  = A166 & A168;
  assign \new_[10310]_  = A200 & A199;
  assign \new_[10311]_  = \new_[10310]_  & \new_[10307]_ ;
  assign \new_[10314]_  = ~A202 & ~A201;
  assign \new_[10318]_  = A301 & A234;
  assign \new_[10319]_  = A232 & \new_[10318]_ ;
  assign \new_[10320]_  = \new_[10319]_  & \new_[10314]_ ;
  assign \new_[10323]_  = A166 & A168;
  assign \new_[10326]_  = A200 & A199;
  assign \new_[10327]_  = \new_[10326]_  & \new_[10323]_ ;
  assign \new_[10330]_  = ~A202 & ~A201;
  assign \new_[10334]_  = A268 & A234;
  assign \new_[10335]_  = A232 & \new_[10334]_ ;
  assign \new_[10336]_  = \new_[10335]_  & \new_[10330]_ ;
  assign \new_[10339]_  = A166 & A168;
  assign \new_[10342]_  = A200 & A199;
  assign \new_[10343]_  = \new_[10342]_  & \new_[10339]_ ;
  assign \new_[10346]_  = ~A202 & ~A201;
  assign \new_[10350]_  = A301 & A234;
  assign \new_[10351]_  = A233 & \new_[10350]_ ;
  assign \new_[10352]_  = \new_[10351]_  & \new_[10346]_ ;
  assign \new_[10355]_  = A166 & A168;
  assign \new_[10358]_  = A200 & A199;
  assign \new_[10359]_  = \new_[10358]_  & \new_[10355]_ ;
  assign \new_[10362]_  = ~A202 & ~A201;
  assign \new_[10366]_  = A268 & A234;
  assign \new_[10367]_  = A233 & \new_[10366]_ ;
  assign \new_[10368]_  = \new_[10367]_  & \new_[10362]_ ;
  assign \new_[10371]_  = A166 & A168;
  assign \new_[10374]_  = ~A200 & ~A199;
  assign \new_[10375]_  = \new_[10374]_  & \new_[10371]_ ;
  assign \new_[10378]_  = A235 & ~A202;
  assign \new_[10382]_  = A302 & ~A299;
  assign \new_[10383]_  = A298 & \new_[10382]_ ;
  assign \new_[10384]_  = \new_[10383]_  & \new_[10378]_ ;
  assign \new_[10387]_  = A166 & A168;
  assign \new_[10390]_  = ~A200 & ~A199;
  assign \new_[10391]_  = \new_[10390]_  & \new_[10387]_ ;
  assign \new_[10394]_  = A235 & ~A202;
  assign \new_[10398]_  = A302 & A299;
  assign \new_[10399]_  = ~A298 & \new_[10398]_ ;
  assign \new_[10400]_  = \new_[10399]_  & \new_[10394]_ ;
  assign \new_[10403]_  = A166 & A168;
  assign \new_[10406]_  = ~A200 & ~A199;
  assign \new_[10407]_  = \new_[10406]_  & \new_[10403]_ ;
  assign \new_[10410]_  = A235 & ~A202;
  assign \new_[10414]_  = A269 & A266;
  assign \new_[10415]_  = ~A265 & \new_[10414]_ ;
  assign \new_[10416]_  = \new_[10415]_  & \new_[10410]_ ;
  assign \new_[10419]_  = A166 & A168;
  assign \new_[10422]_  = ~A200 & ~A199;
  assign \new_[10423]_  = \new_[10422]_  & \new_[10419]_ ;
  assign \new_[10426]_  = A235 & ~A202;
  assign \new_[10430]_  = A269 & ~A266;
  assign \new_[10431]_  = A265 & \new_[10430]_ ;
  assign \new_[10432]_  = \new_[10431]_  & \new_[10426]_ ;
  assign \new_[10435]_  = A166 & A168;
  assign \new_[10438]_  = ~A200 & ~A199;
  assign \new_[10439]_  = \new_[10438]_  & \new_[10435]_ ;
  assign \new_[10442]_  = A232 & ~A202;
  assign \new_[10446]_  = A300 & A299;
  assign \new_[10447]_  = A234 & \new_[10446]_ ;
  assign \new_[10448]_  = \new_[10447]_  & \new_[10442]_ ;
  assign \new_[10451]_  = A166 & A168;
  assign \new_[10454]_  = ~A200 & ~A199;
  assign \new_[10455]_  = \new_[10454]_  & \new_[10451]_ ;
  assign \new_[10458]_  = A232 & ~A202;
  assign \new_[10462]_  = A300 & A298;
  assign \new_[10463]_  = A234 & \new_[10462]_ ;
  assign \new_[10464]_  = \new_[10463]_  & \new_[10458]_ ;
  assign \new_[10467]_  = A166 & A168;
  assign \new_[10470]_  = ~A200 & ~A199;
  assign \new_[10471]_  = \new_[10470]_  & \new_[10467]_ ;
  assign \new_[10474]_  = A232 & ~A202;
  assign \new_[10478]_  = A267 & A265;
  assign \new_[10479]_  = A234 & \new_[10478]_ ;
  assign \new_[10480]_  = \new_[10479]_  & \new_[10474]_ ;
  assign \new_[10483]_  = A166 & A168;
  assign \new_[10486]_  = ~A200 & ~A199;
  assign \new_[10487]_  = \new_[10486]_  & \new_[10483]_ ;
  assign \new_[10490]_  = A232 & ~A202;
  assign \new_[10494]_  = A267 & A266;
  assign \new_[10495]_  = A234 & \new_[10494]_ ;
  assign \new_[10496]_  = \new_[10495]_  & \new_[10490]_ ;
  assign \new_[10499]_  = A166 & A168;
  assign \new_[10502]_  = ~A200 & ~A199;
  assign \new_[10503]_  = \new_[10502]_  & \new_[10499]_ ;
  assign \new_[10506]_  = A233 & ~A202;
  assign \new_[10510]_  = A300 & A299;
  assign \new_[10511]_  = A234 & \new_[10510]_ ;
  assign \new_[10512]_  = \new_[10511]_  & \new_[10506]_ ;
  assign \new_[10515]_  = A166 & A168;
  assign \new_[10518]_  = ~A200 & ~A199;
  assign \new_[10519]_  = \new_[10518]_  & \new_[10515]_ ;
  assign \new_[10522]_  = A233 & ~A202;
  assign \new_[10526]_  = A300 & A298;
  assign \new_[10527]_  = A234 & \new_[10526]_ ;
  assign \new_[10528]_  = \new_[10527]_  & \new_[10522]_ ;
  assign \new_[10531]_  = A166 & A168;
  assign \new_[10534]_  = ~A200 & ~A199;
  assign \new_[10535]_  = \new_[10534]_  & \new_[10531]_ ;
  assign \new_[10538]_  = A233 & ~A202;
  assign \new_[10542]_  = A267 & A265;
  assign \new_[10543]_  = A234 & \new_[10542]_ ;
  assign \new_[10544]_  = \new_[10543]_  & \new_[10538]_ ;
  assign \new_[10547]_  = A166 & A168;
  assign \new_[10550]_  = ~A200 & ~A199;
  assign \new_[10551]_  = \new_[10550]_  & \new_[10547]_ ;
  assign \new_[10554]_  = A233 & ~A202;
  assign \new_[10558]_  = A267 & A266;
  assign \new_[10559]_  = A234 & \new_[10558]_ ;
  assign \new_[10560]_  = \new_[10559]_  & \new_[10554]_ ;
  assign \new_[10563]_  = A166 & A168;
  assign \new_[10566]_  = ~A200 & ~A199;
  assign \new_[10567]_  = \new_[10566]_  & \new_[10563]_ ;
  assign \new_[10570]_  = ~A232 & ~A202;
  assign \new_[10574]_  = A301 & A236;
  assign \new_[10575]_  = A233 & \new_[10574]_ ;
  assign \new_[10576]_  = \new_[10575]_  & \new_[10570]_ ;
  assign \new_[10579]_  = A166 & A168;
  assign \new_[10582]_  = ~A200 & ~A199;
  assign \new_[10583]_  = \new_[10582]_  & \new_[10579]_ ;
  assign \new_[10586]_  = ~A232 & ~A202;
  assign \new_[10590]_  = A268 & A236;
  assign \new_[10591]_  = A233 & \new_[10590]_ ;
  assign \new_[10592]_  = \new_[10591]_  & \new_[10586]_ ;
  assign \new_[10595]_  = A166 & A168;
  assign \new_[10598]_  = ~A200 & ~A199;
  assign \new_[10599]_  = \new_[10598]_  & \new_[10595]_ ;
  assign \new_[10602]_  = A232 & ~A202;
  assign \new_[10606]_  = A301 & A236;
  assign \new_[10607]_  = ~A233 & \new_[10606]_ ;
  assign \new_[10608]_  = \new_[10607]_  & \new_[10602]_ ;
  assign \new_[10611]_  = A166 & A168;
  assign \new_[10614]_  = ~A200 & ~A199;
  assign \new_[10615]_  = \new_[10614]_  & \new_[10611]_ ;
  assign \new_[10618]_  = A232 & ~A202;
  assign \new_[10622]_  = A268 & A236;
  assign \new_[10623]_  = ~A233 & \new_[10622]_ ;
  assign \new_[10624]_  = \new_[10623]_  & \new_[10618]_ ;
  assign \new_[10627]_  = A167 & A168;
  assign \new_[10630]_  = ~A202 & ~A201;
  assign \new_[10631]_  = \new_[10630]_  & \new_[10627]_ ;
  assign \new_[10634]_  = A235 & ~A203;
  assign \new_[10638]_  = A302 & ~A299;
  assign \new_[10639]_  = A298 & \new_[10638]_ ;
  assign \new_[10640]_  = \new_[10639]_  & \new_[10634]_ ;
  assign \new_[10643]_  = A167 & A168;
  assign \new_[10646]_  = ~A202 & ~A201;
  assign \new_[10647]_  = \new_[10646]_  & \new_[10643]_ ;
  assign \new_[10650]_  = A235 & ~A203;
  assign \new_[10654]_  = A302 & A299;
  assign \new_[10655]_  = ~A298 & \new_[10654]_ ;
  assign \new_[10656]_  = \new_[10655]_  & \new_[10650]_ ;
  assign \new_[10659]_  = A167 & A168;
  assign \new_[10662]_  = ~A202 & ~A201;
  assign \new_[10663]_  = \new_[10662]_  & \new_[10659]_ ;
  assign \new_[10666]_  = A235 & ~A203;
  assign \new_[10670]_  = A269 & A266;
  assign \new_[10671]_  = ~A265 & \new_[10670]_ ;
  assign \new_[10672]_  = \new_[10671]_  & \new_[10666]_ ;
  assign \new_[10675]_  = A167 & A168;
  assign \new_[10678]_  = ~A202 & ~A201;
  assign \new_[10679]_  = \new_[10678]_  & \new_[10675]_ ;
  assign \new_[10682]_  = A235 & ~A203;
  assign \new_[10686]_  = A269 & ~A266;
  assign \new_[10687]_  = A265 & \new_[10686]_ ;
  assign \new_[10688]_  = \new_[10687]_  & \new_[10682]_ ;
  assign \new_[10691]_  = A167 & A168;
  assign \new_[10694]_  = ~A202 & ~A201;
  assign \new_[10695]_  = \new_[10694]_  & \new_[10691]_ ;
  assign \new_[10698]_  = A232 & ~A203;
  assign \new_[10702]_  = A300 & A299;
  assign \new_[10703]_  = A234 & \new_[10702]_ ;
  assign \new_[10704]_  = \new_[10703]_  & \new_[10698]_ ;
  assign \new_[10707]_  = A167 & A168;
  assign \new_[10710]_  = ~A202 & ~A201;
  assign \new_[10711]_  = \new_[10710]_  & \new_[10707]_ ;
  assign \new_[10714]_  = A232 & ~A203;
  assign \new_[10718]_  = A300 & A298;
  assign \new_[10719]_  = A234 & \new_[10718]_ ;
  assign \new_[10720]_  = \new_[10719]_  & \new_[10714]_ ;
  assign \new_[10723]_  = A167 & A168;
  assign \new_[10726]_  = ~A202 & ~A201;
  assign \new_[10727]_  = \new_[10726]_  & \new_[10723]_ ;
  assign \new_[10730]_  = A232 & ~A203;
  assign \new_[10734]_  = A267 & A265;
  assign \new_[10735]_  = A234 & \new_[10734]_ ;
  assign \new_[10736]_  = \new_[10735]_  & \new_[10730]_ ;
  assign \new_[10739]_  = A167 & A168;
  assign \new_[10742]_  = ~A202 & ~A201;
  assign \new_[10743]_  = \new_[10742]_  & \new_[10739]_ ;
  assign \new_[10746]_  = A232 & ~A203;
  assign \new_[10750]_  = A267 & A266;
  assign \new_[10751]_  = A234 & \new_[10750]_ ;
  assign \new_[10752]_  = \new_[10751]_  & \new_[10746]_ ;
  assign \new_[10755]_  = A167 & A168;
  assign \new_[10758]_  = ~A202 & ~A201;
  assign \new_[10759]_  = \new_[10758]_  & \new_[10755]_ ;
  assign \new_[10762]_  = A233 & ~A203;
  assign \new_[10766]_  = A300 & A299;
  assign \new_[10767]_  = A234 & \new_[10766]_ ;
  assign \new_[10768]_  = \new_[10767]_  & \new_[10762]_ ;
  assign \new_[10771]_  = A167 & A168;
  assign \new_[10774]_  = ~A202 & ~A201;
  assign \new_[10775]_  = \new_[10774]_  & \new_[10771]_ ;
  assign \new_[10778]_  = A233 & ~A203;
  assign \new_[10782]_  = A300 & A298;
  assign \new_[10783]_  = A234 & \new_[10782]_ ;
  assign \new_[10784]_  = \new_[10783]_  & \new_[10778]_ ;
  assign \new_[10787]_  = A167 & A168;
  assign \new_[10790]_  = ~A202 & ~A201;
  assign \new_[10791]_  = \new_[10790]_  & \new_[10787]_ ;
  assign \new_[10794]_  = A233 & ~A203;
  assign \new_[10798]_  = A267 & A265;
  assign \new_[10799]_  = A234 & \new_[10798]_ ;
  assign \new_[10800]_  = \new_[10799]_  & \new_[10794]_ ;
  assign \new_[10803]_  = A167 & A168;
  assign \new_[10806]_  = ~A202 & ~A201;
  assign \new_[10807]_  = \new_[10806]_  & \new_[10803]_ ;
  assign \new_[10810]_  = A233 & ~A203;
  assign \new_[10814]_  = A267 & A266;
  assign \new_[10815]_  = A234 & \new_[10814]_ ;
  assign \new_[10816]_  = \new_[10815]_  & \new_[10810]_ ;
  assign \new_[10819]_  = A167 & A168;
  assign \new_[10822]_  = ~A202 & ~A201;
  assign \new_[10823]_  = \new_[10822]_  & \new_[10819]_ ;
  assign \new_[10826]_  = ~A232 & ~A203;
  assign \new_[10830]_  = A301 & A236;
  assign \new_[10831]_  = A233 & \new_[10830]_ ;
  assign \new_[10832]_  = \new_[10831]_  & \new_[10826]_ ;
  assign \new_[10835]_  = A167 & A168;
  assign \new_[10838]_  = ~A202 & ~A201;
  assign \new_[10839]_  = \new_[10838]_  & \new_[10835]_ ;
  assign \new_[10842]_  = ~A232 & ~A203;
  assign \new_[10846]_  = A268 & A236;
  assign \new_[10847]_  = A233 & \new_[10846]_ ;
  assign \new_[10848]_  = \new_[10847]_  & \new_[10842]_ ;
  assign \new_[10851]_  = A167 & A168;
  assign \new_[10854]_  = ~A202 & ~A201;
  assign \new_[10855]_  = \new_[10854]_  & \new_[10851]_ ;
  assign \new_[10858]_  = A232 & ~A203;
  assign \new_[10862]_  = A301 & A236;
  assign \new_[10863]_  = ~A233 & \new_[10862]_ ;
  assign \new_[10864]_  = \new_[10863]_  & \new_[10858]_ ;
  assign \new_[10867]_  = A167 & A168;
  assign \new_[10870]_  = ~A202 & ~A201;
  assign \new_[10871]_  = \new_[10870]_  & \new_[10867]_ ;
  assign \new_[10874]_  = A232 & ~A203;
  assign \new_[10878]_  = A268 & A236;
  assign \new_[10879]_  = ~A233 & \new_[10878]_ ;
  assign \new_[10880]_  = \new_[10879]_  & \new_[10874]_ ;
  assign \new_[10883]_  = A167 & A168;
  assign \new_[10886]_  = A200 & A199;
  assign \new_[10887]_  = \new_[10886]_  & \new_[10883]_ ;
  assign \new_[10890]_  = ~A202 & ~A201;
  assign \new_[10894]_  = A300 & A299;
  assign \new_[10895]_  = A235 & \new_[10894]_ ;
  assign \new_[10896]_  = \new_[10895]_  & \new_[10890]_ ;
  assign \new_[10899]_  = A167 & A168;
  assign \new_[10902]_  = A200 & A199;
  assign \new_[10903]_  = \new_[10902]_  & \new_[10899]_ ;
  assign \new_[10906]_  = ~A202 & ~A201;
  assign \new_[10910]_  = A300 & A298;
  assign \new_[10911]_  = A235 & \new_[10910]_ ;
  assign \new_[10912]_  = \new_[10911]_  & \new_[10906]_ ;
  assign \new_[10915]_  = A167 & A168;
  assign \new_[10918]_  = A200 & A199;
  assign \new_[10919]_  = \new_[10918]_  & \new_[10915]_ ;
  assign \new_[10922]_  = ~A202 & ~A201;
  assign \new_[10926]_  = A267 & A265;
  assign \new_[10927]_  = A235 & \new_[10926]_ ;
  assign \new_[10928]_  = \new_[10927]_  & \new_[10922]_ ;
  assign \new_[10931]_  = A167 & A168;
  assign \new_[10934]_  = A200 & A199;
  assign \new_[10935]_  = \new_[10934]_  & \new_[10931]_ ;
  assign \new_[10938]_  = ~A202 & ~A201;
  assign \new_[10942]_  = A267 & A266;
  assign \new_[10943]_  = A235 & \new_[10942]_ ;
  assign \new_[10944]_  = \new_[10943]_  & \new_[10938]_ ;
  assign \new_[10947]_  = A167 & A168;
  assign \new_[10950]_  = A200 & A199;
  assign \new_[10951]_  = \new_[10950]_  & \new_[10947]_ ;
  assign \new_[10954]_  = ~A202 & ~A201;
  assign \new_[10958]_  = A301 & A234;
  assign \new_[10959]_  = A232 & \new_[10958]_ ;
  assign \new_[10960]_  = \new_[10959]_  & \new_[10954]_ ;
  assign \new_[10963]_  = A167 & A168;
  assign \new_[10966]_  = A200 & A199;
  assign \new_[10967]_  = \new_[10966]_  & \new_[10963]_ ;
  assign \new_[10970]_  = ~A202 & ~A201;
  assign \new_[10974]_  = A268 & A234;
  assign \new_[10975]_  = A232 & \new_[10974]_ ;
  assign \new_[10976]_  = \new_[10975]_  & \new_[10970]_ ;
  assign \new_[10979]_  = A167 & A168;
  assign \new_[10982]_  = A200 & A199;
  assign \new_[10983]_  = \new_[10982]_  & \new_[10979]_ ;
  assign \new_[10986]_  = ~A202 & ~A201;
  assign \new_[10990]_  = A301 & A234;
  assign \new_[10991]_  = A233 & \new_[10990]_ ;
  assign \new_[10992]_  = \new_[10991]_  & \new_[10986]_ ;
  assign \new_[10995]_  = A167 & A168;
  assign \new_[10998]_  = A200 & A199;
  assign \new_[10999]_  = \new_[10998]_  & \new_[10995]_ ;
  assign \new_[11002]_  = ~A202 & ~A201;
  assign \new_[11006]_  = A268 & A234;
  assign \new_[11007]_  = A233 & \new_[11006]_ ;
  assign \new_[11008]_  = \new_[11007]_  & \new_[11002]_ ;
  assign \new_[11011]_  = A167 & A168;
  assign \new_[11014]_  = ~A200 & ~A199;
  assign \new_[11015]_  = \new_[11014]_  & \new_[11011]_ ;
  assign \new_[11018]_  = A235 & ~A202;
  assign \new_[11022]_  = A302 & ~A299;
  assign \new_[11023]_  = A298 & \new_[11022]_ ;
  assign \new_[11024]_  = \new_[11023]_  & \new_[11018]_ ;
  assign \new_[11027]_  = A167 & A168;
  assign \new_[11030]_  = ~A200 & ~A199;
  assign \new_[11031]_  = \new_[11030]_  & \new_[11027]_ ;
  assign \new_[11034]_  = A235 & ~A202;
  assign \new_[11038]_  = A302 & A299;
  assign \new_[11039]_  = ~A298 & \new_[11038]_ ;
  assign \new_[11040]_  = \new_[11039]_  & \new_[11034]_ ;
  assign \new_[11043]_  = A167 & A168;
  assign \new_[11046]_  = ~A200 & ~A199;
  assign \new_[11047]_  = \new_[11046]_  & \new_[11043]_ ;
  assign \new_[11050]_  = A235 & ~A202;
  assign \new_[11054]_  = A269 & A266;
  assign \new_[11055]_  = ~A265 & \new_[11054]_ ;
  assign \new_[11056]_  = \new_[11055]_  & \new_[11050]_ ;
  assign \new_[11059]_  = A167 & A168;
  assign \new_[11062]_  = ~A200 & ~A199;
  assign \new_[11063]_  = \new_[11062]_  & \new_[11059]_ ;
  assign \new_[11066]_  = A235 & ~A202;
  assign \new_[11070]_  = A269 & ~A266;
  assign \new_[11071]_  = A265 & \new_[11070]_ ;
  assign \new_[11072]_  = \new_[11071]_  & \new_[11066]_ ;
  assign \new_[11075]_  = A167 & A168;
  assign \new_[11078]_  = ~A200 & ~A199;
  assign \new_[11079]_  = \new_[11078]_  & \new_[11075]_ ;
  assign \new_[11082]_  = A232 & ~A202;
  assign \new_[11086]_  = A300 & A299;
  assign \new_[11087]_  = A234 & \new_[11086]_ ;
  assign \new_[11088]_  = \new_[11087]_  & \new_[11082]_ ;
  assign \new_[11091]_  = A167 & A168;
  assign \new_[11094]_  = ~A200 & ~A199;
  assign \new_[11095]_  = \new_[11094]_  & \new_[11091]_ ;
  assign \new_[11098]_  = A232 & ~A202;
  assign \new_[11102]_  = A300 & A298;
  assign \new_[11103]_  = A234 & \new_[11102]_ ;
  assign \new_[11104]_  = \new_[11103]_  & \new_[11098]_ ;
  assign \new_[11107]_  = A167 & A168;
  assign \new_[11110]_  = ~A200 & ~A199;
  assign \new_[11111]_  = \new_[11110]_  & \new_[11107]_ ;
  assign \new_[11114]_  = A232 & ~A202;
  assign \new_[11118]_  = A267 & A265;
  assign \new_[11119]_  = A234 & \new_[11118]_ ;
  assign \new_[11120]_  = \new_[11119]_  & \new_[11114]_ ;
  assign \new_[11123]_  = A167 & A168;
  assign \new_[11126]_  = ~A200 & ~A199;
  assign \new_[11127]_  = \new_[11126]_  & \new_[11123]_ ;
  assign \new_[11130]_  = A232 & ~A202;
  assign \new_[11134]_  = A267 & A266;
  assign \new_[11135]_  = A234 & \new_[11134]_ ;
  assign \new_[11136]_  = \new_[11135]_  & \new_[11130]_ ;
  assign \new_[11139]_  = A167 & A168;
  assign \new_[11142]_  = ~A200 & ~A199;
  assign \new_[11143]_  = \new_[11142]_  & \new_[11139]_ ;
  assign \new_[11146]_  = A233 & ~A202;
  assign \new_[11150]_  = A300 & A299;
  assign \new_[11151]_  = A234 & \new_[11150]_ ;
  assign \new_[11152]_  = \new_[11151]_  & \new_[11146]_ ;
  assign \new_[11155]_  = A167 & A168;
  assign \new_[11158]_  = ~A200 & ~A199;
  assign \new_[11159]_  = \new_[11158]_  & \new_[11155]_ ;
  assign \new_[11162]_  = A233 & ~A202;
  assign \new_[11166]_  = A300 & A298;
  assign \new_[11167]_  = A234 & \new_[11166]_ ;
  assign \new_[11168]_  = \new_[11167]_  & \new_[11162]_ ;
  assign \new_[11171]_  = A167 & A168;
  assign \new_[11174]_  = ~A200 & ~A199;
  assign \new_[11175]_  = \new_[11174]_  & \new_[11171]_ ;
  assign \new_[11178]_  = A233 & ~A202;
  assign \new_[11182]_  = A267 & A265;
  assign \new_[11183]_  = A234 & \new_[11182]_ ;
  assign \new_[11184]_  = \new_[11183]_  & \new_[11178]_ ;
  assign \new_[11187]_  = A167 & A168;
  assign \new_[11190]_  = ~A200 & ~A199;
  assign \new_[11191]_  = \new_[11190]_  & \new_[11187]_ ;
  assign \new_[11194]_  = A233 & ~A202;
  assign \new_[11198]_  = A267 & A266;
  assign \new_[11199]_  = A234 & \new_[11198]_ ;
  assign \new_[11200]_  = \new_[11199]_  & \new_[11194]_ ;
  assign \new_[11203]_  = A167 & A168;
  assign \new_[11206]_  = ~A200 & ~A199;
  assign \new_[11207]_  = \new_[11206]_  & \new_[11203]_ ;
  assign \new_[11210]_  = ~A232 & ~A202;
  assign \new_[11214]_  = A301 & A236;
  assign \new_[11215]_  = A233 & \new_[11214]_ ;
  assign \new_[11216]_  = \new_[11215]_  & \new_[11210]_ ;
  assign \new_[11219]_  = A167 & A168;
  assign \new_[11222]_  = ~A200 & ~A199;
  assign \new_[11223]_  = \new_[11222]_  & \new_[11219]_ ;
  assign \new_[11226]_  = ~A232 & ~A202;
  assign \new_[11230]_  = A268 & A236;
  assign \new_[11231]_  = A233 & \new_[11230]_ ;
  assign \new_[11232]_  = \new_[11231]_  & \new_[11226]_ ;
  assign \new_[11235]_  = A167 & A168;
  assign \new_[11238]_  = ~A200 & ~A199;
  assign \new_[11239]_  = \new_[11238]_  & \new_[11235]_ ;
  assign \new_[11242]_  = A232 & ~A202;
  assign \new_[11246]_  = A301 & A236;
  assign \new_[11247]_  = ~A233 & \new_[11246]_ ;
  assign \new_[11248]_  = \new_[11247]_  & \new_[11242]_ ;
  assign \new_[11251]_  = A167 & A168;
  assign \new_[11254]_  = ~A200 & ~A199;
  assign \new_[11255]_  = \new_[11254]_  & \new_[11251]_ ;
  assign \new_[11258]_  = A232 & ~A202;
  assign \new_[11262]_  = A268 & A236;
  assign \new_[11263]_  = ~A233 & \new_[11262]_ ;
  assign \new_[11264]_  = \new_[11263]_  & \new_[11258]_ ;
  assign \new_[11267]_  = A167 & A170;
  assign \new_[11270]_  = ~A201 & ~A166;
  assign \new_[11271]_  = \new_[11270]_  & \new_[11267]_ ;
  assign \new_[11274]_  = ~A203 & ~A202;
  assign \new_[11278]_  = A300 & A299;
  assign \new_[11279]_  = A235 & \new_[11278]_ ;
  assign \new_[11280]_  = \new_[11279]_  & \new_[11274]_ ;
  assign \new_[11283]_  = A167 & A170;
  assign \new_[11286]_  = ~A201 & ~A166;
  assign \new_[11287]_  = \new_[11286]_  & \new_[11283]_ ;
  assign \new_[11290]_  = ~A203 & ~A202;
  assign \new_[11294]_  = A300 & A298;
  assign \new_[11295]_  = A235 & \new_[11294]_ ;
  assign \new_[11296]_  = \new_[11295]_  & \new_[11290]_ ;
  assign \new_[11299]_  = A167 & A170;
  assign \new_[11302]_  = ~A201 & ~A166;
  assign \new_[11303]_  = \new_[11302]_  & \new_[11299]_ ;
  assign \new_[11306]_  = ~A203 & ~A202;
  assign \new_[11310]_  = A267 & A265;
  assign \new_[11311]_  = A235 & \new_[11310]_ ;
  assign \new_[11312]_  = \new_[11311]_  & \new_[11306]_ ;
  assign \new_[11315]_  = A167 & A170;
  assign \new_[11318]_  = ~A201 & ~A166;
  assign \new_[11319]_  = \new_[11318]_  & \new_[11315]_ ;
  assign \new_[11322]_  = ~A203 & ~A202;
  assign \new_[11326]_  = A267 & A266;
  assign \new_[11327]_  = A235 & \new_[11326]_ ;
  assign \new_[11328]_  = \new_[11327]_  & \new_[11322]_ ;
  assign \new_[11331]_  = A167 & A170;
  assign \new_[11334]_  = ~A201 & ~A166;
  assign \new_[11335]_  = \new_[11334]_  & \new_[11331]_ ;
  assign \new_[11338]_  = ~A203 & ~A202;
  assign \new_[11342]_  = A301 & A234;
  assign \new_[11343]_  = A232 & \new_[11342]_ ;
  assign \new_[11344]_  = \new_[11343]_  & \new_[11338]_ ;
  assign \new_[11347]_  = A167 & A170;
  assign \new_[11350]_  = ~A201 & ~A166;
  assign \new_[11351]_  = \new_[11350]_  & \new_[11347]_ ;
  assign \new_[11354]_  = ~A203 & ~A202;
  assign \new_[11358]_  = A268 & A234;
  assign \new_[11359]_  = A232 & \new_[11358]_ ;
  assign \new_[11360]_  = \new_[11359]_  & \new_[11354]_ ;
  assign \new_[11363]_  = A167 & A170;
  assign \new_[11366]_  = ~A201 & ~A166;
  assign \new_[11367]_  = \new_[11366]_  & \new_[11363]_ ;
  assign \new_[11370]_  = ~A203 & ~A202;
  assign \new_[11374]_  = A301 & A234;
  assign \new_[11375]_  = A233 & \new_[11374]_ ;
  assign \new_[11376]_  = \new_[11375]_  & \new_[11370]_ ;
  assign \new_[11379]_  = A167 & A170;
  assign \new_[11382]_  = ~A201 & ~A166;
  assign \new_[11383]_  = \new_[11382]_  & \new_[11379]_ ;
  assign \new_[11386]_  = ~A203 & ~A202;
  assign \new_[11390]_  = A268 & A234;
  assign \new_[11391]_  = A233 & \new_[11390]_ ;
  assign \new_[11392]_  = \new_[11391]_  & \new_[11386]_ ;
  assign \new_[11395]_  = A167 & A170;
  assign \new_[11398]_  = A199 & ~A166;
  assign \new_[11399]_  = \new_[11398]_  & \new_[11395]_ ;
  assign \new_[11402]_  = ~A201 & A200;
  assign \new_[11406]_  = A301 & A235;
  assign \new_[11407]_  = ~A202 & \new_[11406]_ ;
  assign \new_[11408]_  = \new_[11407]_  & \new_[11402]_ ;
  assign \new_[11411]_  = A167 & A170;
  assign \new_[11414]_  = A199 & ~A166;
  assign \new_[11415]_  = \new_[11414]_  & \new_[11411]_ ;
  assign \new_[11418]_  = ~A201 & A200;
  assign \new_[11422]_  = A268 & A235;
  assign \new_[11423]_  = ~A202 & \new_[11422]_ ;
  assign \new_[11424]_  = \new_[11423]_  & \new_[11418]_ ;
  assign \new_[11427]_  = A167 & A170;
  assign \new_[11430]_  = ~A199 & ~A166;
  assign \new_[11431]_  = \new_[11430]_  & \new_[11427]_ ;
  assign \new_[11434]_  = ~A202 & ~A200;
  assign \new_[11438]_  = A300 & A299;
  assign \new_[11439]_  = A235 & \new_[11438]_ ;
  assign \new_[11440]_  = \new_[11439]_  & \new_[11434]_ ;
  assign \new_[11443]_  = A167 & A170;
  assign \new_[11446]_  = ~A199 & ~A166;
  assign \new_[11447]_  = \new_[11446]_  & \new_[11443]_ ;
  assign \new_[11450]_  = ~A202 & ~A200;
  assign \new_[11454]_  = A300 & A298;
  assign \new_[11455]_  = A235 & \new_[11454]_ ;
  assign \new_[11456]_  = \new_[11455]_  & \new_[11450]_ ;
  assign \new_[11459]_  = A167 & A170;
  assign \new_[11462]_  = ~A199 & ~A166;
  assign \new_[11463]_  = \new_[11462]_  & \new_[11459]_ ;
  assign \new_[11466]_  = ~A202 & ~A200;
  assign \new_[11470]_  = A267 & A265;
  assign \new_[11471]_  = A235 & \new_[11470]_ ;
  assign \new_[11472]_  = \new_[11471]_  & \new_[11466]_ ;
  assign \new_[11475]_  = A167 & A170;
  assign \new_[11478]_  = ~A199 & ~A166;
  assign \new_[11479]_  = \new_[11478]_  & \new_[11475]_ ;
  assign \new_[11482]_  = ~A202 & ~A200;
  assign \new_[11486]_  = A267 & A266;
  assign \new_[11487]_  = A235 & \new_[11486]_ ;
  assign \new_[11488]_  = \new_[11487]_  & \new_[11482]_ ;
  assign \new_[11491]_  = A167 & A170;
  assign \new_[11494]_  = ~A199 & ~A166;
  assign \new_[11495]_  = \new_[11494]_  & \new_[11491]_ ;
  assign \new_[11498]_  = ~A202 & ~A200;
  assign \new_[11502]_  = A301 & A234;
  assign \new_[11503]_  = A232 & \new_[11502]_ ;
  assign \new_[11504]_  = \new_[11503]_  & \new_[11498]_ ;
  assign \new_[11507]_  = A167 & A170;
  assign \new_[11510]_  = ~A199 & ~A166;
  assign \new_[11511]_  = \new_[11510]_  & \new_[11507]_ ;
  assign \new_[11514]_  = ~A202 & ~A200;
  assign \new_[11518]_  = A268 & A234;
  assign \new_[11519]_  = A232 & \new_[11518]_ ;
  assign \new_[11520]_  = \new_[11519]_  & \new_[11514]_ ;
  assign \new_[11523]_  = A167 & A170;
  assign \new_[11526]_  = ~A199 & ~A166;
  assign \new_[11527]_  = \new_[11526]_  & \new_[11523]_ ;
  assign \new_[11530]_  = ~A202 & ~A200;
  assign \new_[11534]_  = A301 & A234;
  assign \new_[11535]_  = A233 & \new_[11534]_ ;
  assign \new_[11536]_  = \new_[11535]_  & \new_[11530]_ ;
  assign \new_[11539]_  = A167 & A170;
  assign \new_[11542]_  = ~A199 & ~A166;
  assign \new_[11543]_  = \new_[11542]_  & \new_[11539]_ ;
  assign \new_[11546]_  = ~A202 & ~A200;
  assign \new_[11550]_  = A268 & A234;
  assign \new_[11551]_  = A233 & \new_[11550]_ ;
  assign \new_[11552]_  = \new_[11551]_  & \new_[11546]_ ;
  assign \new_[11555]_  = ~A167 & A170;
  assign \new_[11558]_  = ~A201 & A166;
  assign \new_[11559]_  = \new_[11558]_  & \new_[11555]_ ;
  assign \new_[11562]_  = ~A203 & ~A202;
  assign \new_[11566]_  = A300 & A299;
  assign \new_[11567]_  = A235 & \new_[11566]_ ;
  assign \new_[11568]_  = \new_[11567]_  & \new_[11562]_ ;
  assign \new_[11571]_  = ~A167 & A170;
  assign \new_[11574]_  = ~A201 & A166;
  assign \new_[11575]_  = \new_[11574]_  & \new_[11571]_ ;
  assign \new_[11578]_  = ~A203 & ~A202;
  assign \new_[11582]_  = A300 & A298;
  assign \new_[11583]_  = A235 & \new_[11582]_ ;
  assign \new_[11584]_  = \new_[11583]_  & \new_[11578]_ ;
  assign \new_[11587]_  = ~A167 & A170;
  assign \new_[11590]_  = ~A201 & A166;
  assign \new_[11591]_  = \new_[11590]_  & \new_[11587]_ ;
  assign \new_[11594]_  = ~A203 & ~A202;
  assign \new_[11598]_  = A267 & A265;
  assign \new_[11599]_  = A235 & \new_[11598]_ ;
  assign \new_[11600]_  = \new_[11599]_  & \new_[11594]_ ;
  assign \new_[11603]_  = ~A167 & A170;
  assign \new_[11606]_  = ~A201 & A166;
  assign \new_[11607]_  = \new_[11606]_  & \new_[11603]_ ;
  assign \new_[11610]_  = ~A203 & ~A202;
  assign \new_[11614]_  = A267 & A266;
  assign \new_[11615]_  = A235 & \new_[11614]_ ;
  assign \new_[11616]_  = \new_[11615]_  & \new_[11610]_ ;
  assign \new_[11619]_  = ~A167 & A170;
  assign \new_[11622]_  = ~A201 & A166;
  assign \new_[11623]_  = \new_[11622]_  & \new_[11619]_ ;
  assign \new_[11626]_  = ~A203 & ~A202;
  assign \new_[11630]_  = A301 & A234;
  assign \new_[11631]_  = A232 & \new_[11630]_ ;
  assign \new_[11632]_  = \new_[11631]_  & \new_[11626]_ ;
  assign \new_[11635]_  = ~A167 & A170;
  assign \new_[11638]_  = ~A201 & A166;
  assign \new_[11639]_  = \new_[11638]_  & \new_[11635]_ ;
  assign \new_[11642]_  = ~A203 & ~A202;
  assign \new_[11646]_  = A268 & A234;
  assign \new_[11647]_  = A232 & \new_[11646]_ ;
  assign \new_[11648]_  = \new_[11647]_  & \new_[11642]_ ;
  assign \new_[11651]_  = ~A167 & A170;
  assign \new_[11654]_  = ~A201 & A166;
  assign \new_[11655]_  = \new_[11654]_  & \new_[11651]_ ;
  assign \new_[11658]_  = ~A203 & ~A202;
  assign \new_[11662]_  = A301 & A234;
  assign \new_[11663]_  = A233 & \new_[11662]_ ;
  assign \new_[11664]_  = \new_[11663]_  & \new_[11658]_ ;
  assign \new_[11667]_  = ~A167 & A170;
  assign \new_[11670]_  = ~A201 & A166;
  assign \new_[11671]_  = \new_[11670]_  & \new_[11667]_ ;
  assign \new_[11674]_  = ~A203 & ~A202;
  assign \new_[11678]_  = A268 & A234;
  assign \new_[11679]_  = A233 & \new_[11678]_ ;
  assign \new_[11680]_  = \new_[11679]_  & \new_[11674]_ ;
  assign \new_[11683]_  = ~A167 & A170;
  assign \new_[11686]_  = A199 & A166;
  assign \new_[11687]_  = \new_[11686]_  & \new_[11683]_ ;
  assign \new_[11690]_  = ~A201 & A200;
  assign \new_[11694]_  = A301 & A235;
  assign \new_[11695]_  = ~A202 & \new_[11694]_ ;
  assign \new_[11696]_  = \new_[11695]_  & \new_[11690]_ ;
  assign \new_[11699]_  = ~A167 & A170;
  assign \new_[11702]_  = A199 & A166;
  assign \new_[11703]_  = \new_[11702]_  & \new_[11699]_ ;
  assign \new_[11706]_  = ~A201 & A200;
  assign \new_[11710]_  = A268 & A235;
  assign \new_[11711]_  = ~A202 & \new_[11710]_ ;
  assign \new_[11712]_  = \new_[11711]_  & \new_[11706]_ ;
  assign \new_[11715]_  = ~A167 & A170;
  assign \new_[11718]_  = ~A199 & A166;
  assign \new_[11719]_  = \new_[11718]_  & \new_[11715]_ ;
  assign \new_[11722]_  = ~A202 & ~A200;
  assign \new_[11726]_  = A300 & A299;
  assign \new_[11727]_  = A235 & \new_[11726]_ ;
  assign \new_[11728]_  = \new_[11727]_  & \new_[11722]_ ;
  assign \new_[11731]_  = ~A167 & A170;
  assign \new_[11734]_  = ~A199 & A166;
  assign \new_[11735]_  = \new_[11734]_  & \new_[11731]_ ;
  assign \new_[11738]_  = ~A202 & ~A200;
  assign \new_[11742]_  = A300 & A298;
  assign \new_[11743]_  = A235 & \new_[11742]_ ;
  assign \new_[11744]_  = \new_[11743]_  & \new_[11738]_ ;
  assign \new_[11747]_  = ~A167 & A170;
  assign \new_[11750]_  = ~A199 & A166;
  assign \new_[11751]_  = \new_[11750]_  & \new_[11747]_ ;
  assign \new_[11754]_  = ~A202 & ~A200;
  assign \new_[11758]_  = A267 & A265;
  assign \new_[11759]_  = A235 & \new_[11758]_ ;
  assign \new_[11760]_  = \new_[11759]_  & \new_[11754]_ ;
  assign \new_[11763]_  = ~A167 & A170;
  assign \new_[11766]_  = ~A199 & A166;
  assign \new_[11767]_  = \new_[11766]_  & \new_[11763]_ ;
  assign \new_[11770]_  = ~A202 & ~A200;
  assign \new_[11774]_  = A267 & A266;
  assign \new_[11775]_  = A235 & \new_[11774]_ ;
  assign \new_[11776]_  = \new_[11775]_  & \new_[11770]_ ;
  assign \new_[11779]_  = ~A167 & A170;
  assign \new_[11782]_  = ~A199 & A166;
  assign \new_[11783]_  = \new_[11782]_  & \new_[11779]_ ;
  assign \new_[11786]_  = ~A202 & ~A200;
  assign \new_[11790]_  = A301 & A234;
  assign \new_[11791]_  = A232 & \new_[11790]_ ;
  assign \new_[11792]_  = \new_[11791]_  & \new_[11786]_ ;
  assign \new_[11795]_  = ~A167 & A170;
  assign \new_[11798]_  = ~A199 & A166;
  assign \new_[11799]_  = \new_[11798]_  & \new_[11795]_ ;
  assign \new_[11802]_  = ~A202 & ~A200;
  assign \new_[11806]_  = A268 & A234;
  assign \new_[11807]_  = A232 & \new_[11806]_ ;
  assign \new_[11808]_  = \new_[11807]_  & \new_[11802]_ ;
  assign \new_[11811]_  = ~A167 & A170;
  assign \new_[11814]_  = ~A199 & A166;
  assign \new_[11815]_  = \new_[11814]_  & \new_[11811]_ ;
  assign \new_[11818]_  = ~A202 & ~A200;
  assign \new_[11822]_  = A301 & A234;
  assign \new_[11823]_  = A233 & \new_[11822]_ ;
  assign \new_[11824]_  = \new_[11823]_  & \new_[11818]_ ;
  assign \new_[11827]_  = ~A167 & A170;
  assign \new_[11830]_  = ~A199 & A166;
  assign \new_[11831]_  = \new_[11830]_  & \new_[11827]_ ;
  assign \new_[11834]_  = ~A202 & ~A200;
  assign \new_[11838]_  = A268 & A234;
  assign \new_[11839]_  = A233 & \new_[11838]_ ;
  assign \new_[11840]_  = \new_[11839]_  & \new_[11834]_ ;
  assign \new_[11843]_  = ~A201 & A169;
  assign \new_[11846]_  = ~A203 & ~A202;
  assign \new_[11847]_  = \new_[11846]_  & \new_[11843]_ ;
  assign \new_[11850]_  = A234 & A232;
  assign \new_[11854]_  = A302 & ~A299;
  assign \new_[11855]_  = A298 & \new_[11854]_ ;
  assign \new_[11856]_  = \new_[11855]_  & \new_[11850]_ ;
  assign \new_[11859]_  = ~A201 & A169;
  assign \new_[11862]_  = ~A203 & ~A202;
  assign \new_[11863]_  = \new_[11862]_  & \new_[11859]_ ;
  assign \new_[11866]_  = A234 & A232;
  assign \new_[11870]_  = A302 & A299;
  assign \new_[11871]_  = ~A298 & \new_[11870]_ ;
  assign \new_[11872]_  = \new_[11871]_  & \new_[11866]_ ;
  assign \new_[11875]_  = ~A201 & A169;
  assign \new_[11878]_  = ~A203 & ~A202;
  assign \new_[11879]_  = \new_[11878]_  & \new_[11875]_ ;
  assign \new_[11882]_  = A234 & A232;
  assign \new_[11886]_  = A269 & A266;
  assign \new_[11887]_  = ~A265 & \new_[11886]_ ;
  assign \new_[11888]_  = \new_[11887]_  & \new_[11882]_ ;
  assign \new_[11891]_  = ~A201 & A169;
  assign \new_[11894]_  = ~A203 & ~A202;
  assign \new_[11895]_  = \new_[11894]_  & \new_[11891]_ ;
  assign \new_[11898]_  = A234 & A232;
  assign \new_[11902]_  = A269 & ~A266;
  assign \new_[11903]_  = A265 & \new_[11902]_ ;
  assign \new_[11904]_  = \new_[11903]_  & \new_[11898]_ ;
  assign \new_[11907]_  = ~A201 & A169;
  assign \new_[11910]_  = ~A203 & ~A202;
  assign \new_[11911]_  = \new_[11910]_  & \new_[11907]_ ;
  assign \new_[11914]_  = A234 & A233;
  assign \new_[11918]_  = A302 & ~A299;
  assign \new_[11919]_  = A298 & \new_[11918]_ ;
  assign \new_[11920]_  = \new_[11919]_  & \new_[11914]_ ;
  assign \new_[11923]_  = ~A201 & A169;
  assign \new_[11926]_  = ~A203 & ~A202;
  assign \new_[11927]_  = \new_[11926]_  & \new_[11923]_ ;
  assign \new_[11930]_  = A234 & A233;
  assign \new_[11934]_  = A302 & A299;
  assign \new_[11935]_  = ~A298 & \new_[11934]_ ;
  assign \new_[11936]_  = \new_[11935]_  & \new_[11930]_ ;
  assign \new_[11939]_  = ~A201 & A169;
  assign \new_[11942]_  = ~A203 & ~A202;
  assign \new_[11943]_  = \new_[11942]_  & \new_[11939]_ ;
  assign \new_[11946]_  = A234 & A233;
  assign \new_[11950]_  = A269 & A266;
  assign \new_[11951]_  = ~A265 & \new_[11950]_ ;
  assign \new_[11952]_  = \new_[11951]_  & \new_[11946]_ ;
  assign \new_[11955]_  = ~A201 & A169;
  assign \new_[11958]_  = ~A203 & ~A202;
  assign \new_[11959]_  = \new_[11958]_  & \new_[11955]_ ;
  assign \new_[11962]_  = A234 & A233;
  assign \new_[11966]_  = A269 & ~A266;
  assign \new_[11967]_  = A265 & \new_[11966]_ ;
  assign \new_[11968]_  = \new_[11967]_  & \new_[11962]_ ;
  assign \new_[11971]_  = ~A201 & A169;
  assign \new_[11974]_  = ~A203 & ~A202;
  assign \new_[11975]_  = \new_[11974]_  & \new_[11971]_ ;
  assign \new_[11978]_  = A233 & ~A232;
  assign \new_[11982]_  = A300 & A299;
  assign \new_[11983]_  = A236 & \new_[11982]_ ;
  assign \new_[11984]_  = \new_[11983]_  & \new_[11978]_ ;
  assign \new_[11987]_  = ~A201 & A169;
  assign \new_[11990]_  = ~A203 & ~A202;
  assign \new_[11991]_  = \new_[11990]_  & \new_[11987]_ ;
  assign \new_[11994]_  = A233 & ~A232;
  assign \new_[11998]_  = A300 & A298;
  assign \new_[11999]_  = A236 & \new_[11998]_ ;
  assign \new_[12000]_  = \new_[11999]_  & \new_[11994]_ ;
  assign \new_[12003]_  = ~A201 & A169;
  assign \new_[12006]_  = ~A203 & ~A202;
  assign \new_[12007]_  = \new_[12006]_  & \new_[12003]_ ;
  assign \new_[12010]_  = A233 & ~A232;
  assign \new_[12014]_  = A267 & A265;
  assign \new_[12015]_  = A236 & \new_[12014]_ ;
  assign \new_[12016]_  = \new_[12015]_  & \new_[12010]_ ;
  assign \new_[12019]_  = ~A201 & A169;
  assign \new_[12022]_  = ~A203 & ~A202;
  assign \new_[12023]_  = \new_[12022]_  & \new_[12019]_ ;
  assign \new_[12026]_  = A233 & ~A232;
  assign \new_[12030]_  = A267 & A266;
  assign \new_[12031]_  = A236 & \new_[12030]_ ;
  assign \new_[12032]_  = \new_[12031]_  & \new_[12026]_ ;
  assign \new_[12035]_  = ~A201 & A169;
  assign \new_[12038]_  = ~A203 & ~A202;
  assign \new_[12039]_  = \new_[12038]_  & \new_[12035]_ ;
  assign \new_[12042]_  = ~A233 & A232;
  assign \new_[12046]_  = A300 & A299;
  assign \new_[12047]_  = A236 & \new_[12046]_ ;
  assign \new_[12048]_  = \new_[12047]_  & \new_[12042]_ ;
  assign \new_[12051]_  = ~A201 & A169;
  assign \new_[12054]_  = ~A203 & ~A202;
  assign \new_[12055]_  = \new_[12054]_  & \new_[12051]_ ;
  assign \new_[12058]_  = ~A233 & A232;
  assign \new_[12062]_  = A300 & A298;
  assign \new_[12063]_  = A236 & \new_[12062]_ ;
  assign \new_[12064]_  = \new_[12063]_  & \new_[12058]_ ;
  assign \new_[12067]_  = ~A201 & A169;
  assign \new_[12070]_  = ~A203 & ~A202;
  assign \new_[12071]_  = \new_[12070]_  & \new_[12067]_ ;
  assign \new_[12074]_  = ~A233 & A232;
  assign \new_[12078]_  = A267 & A265;
  assign \new_[12079]_  = A236 & \new_[12078]_ ;
  assign \new_[12080]_  = \new_[12079]_  & \new_[12074]_ ;
  assign \new_[12083]_  = ~A201 & A169;
  assign \new_[12086]_  = ~A203 & ~A202;
  assign \new_[12087]_  = \new_[12086]_  & \new_[12083]_ ;
  assign \new_[12090]_  = ~A233 & A232;
  assign \new_[12094]_  = A267 & A266;
  assign \new_[12095]_  = A236 & \new_[12094]_ ;
  assign \new_[12096]_  = \new_[12095]_  & \new_[12090]_ ;
  assign \new_[12099]_  = A199 & A169;
  assign \new_[12102]_  = ~A201 & A200;
  assign \new_[12103]_  = \new_[12102]_  & \new_[12099]_ ;
  assign \new_[12106]_  = A235 & ~A202;
  assign \new_[12110]_  = A302 & ~A299;
  assign \new_[12111]_  = A298 & \new_[12110]_ ;
  assign \new_[12112]_  = \new_[12111]_  & \new_[12106]_ ;
  assign \new_[12115]_  = A199 & A169;
  assign \new_[12118]_  = ~A201 & A200;
  assign \new_[12119]_  = \new_[12118]_  & \new_[12115]_ ;
  assign \new_[12122]_  = A235 & ~A202;
  assign \new_[12126]_  = A302 & A299;
  assign \new_[12127]_  = ~A298 & \new_[12126]_ ;
  assign \new_[12128]_  = \new_[12127]_  & \new_[12122]_ ;
  assign \new_[12131]_  = A199 & A169;
  assign \new_[12134]_  = ~A201 & A200;
  assign \new_[12135]_  = \new_[12134]_  & \new_[12131]_ ;
  assign \new_[12138]_  = A235 & ~A202;
  assign \new_[12142]_  = A269 & A266;
  assign \new_[12143]_  = ~A265 & \new_[12142]_ ;
  assign \new_[12144]_  = \new_[12143]_  & \new_[12138]_ ;
  assign \new_[12147]_  = A199 & A169;
  assign \new_[12150]_  = ~A201 & A200;
  assign \new_[12151]_  = \new_[12150]_  & \new_[12147]_ ;
  assign \new_[12154]_  = A235 & ~A202;
  assign \new_[12158]_  = A269 & ~A266;
  assign \new_[12159]_  = A265 & \new_[12158]_ ;
  assign \new_[12160]_  = \new_[12159]_  & \new_[12154]_ ;
  assign \new_[12163]_  = A199 & A169;
  assign \new_[12166]_  = ~A201 & A200;
  assign \new_[12167]_  = \new_[12166]_  & \new_[12163]_ ;
  assign \new_[12170]_  = A232 & ~A202;
  assign \new_[12174]_  = A300 & A299;
  assign \new_[12175]_  = A234 & \new_[12174]_ ;
  assign \new_[12176]_  = \new_[12175]_  & \new_[12170]_ ;
  assign \new_[12179]_  = A199 & A169;
  assign \new_[12182]_  = ~A201 & A200;
  assign \new_[12183]_  = \new_[12182]_  & \new_[12179]_ ;
  assign \new_[12186]_  = A232 & ~A202;
  assign \new_[12190]_  = A300 & A298;
  assign \new_[12191]_  = A234 & \new_[12190]_ ;
  assign \new_[12192]_  = \new_[12191]_  & \new_[12186]_ ;
  assign \new_[12195]_  = A199 & A169;
  assign \new_[12198]_  = ~A201 & A200;
  assign \new_[12199]_  = \new_[12198]_  & \new_[12195]_ ;
  assign \new_[12202]_  = A232 & ~A202;
  assign \new_[12206]_  = A267 & A265;
  assign \new_[12207]_  = A234 & \new_[12206]_ ;
  assign \new_[12208]_  = \new_[12207]_  & \new_[12202]_ ;
  assign \new_[12211]_  = A199 & A169;
  assign \new_[12214]_  = ~A201 & A200;
  assign \new_[12215]_  = \new_[12214]_  & \new_[12211]_ ;
  assign \new_[12218]_  = A232 & ~A202;
  assign \new_[12222]_  = A267 & A266;
  assign \new_[12223]_  = A234 & \new_[12222]_ ;
  assign \new_[12224]_  = \new_[12223]_  & \new_[12218]_ ;
  assign \new_[12227]_  = A199 & A169;
  assign \new_[12230]_  = ~A201 & A200;
  assign \new_[12231]_  = \new_[12230]_  & \new_[12227]_ ;
  assign \new_[12234]_  = A233 & ~A202;
  assign \new_[12238]_  = A300 & A299;
  assign \new_[12239]_  = A234 & \new_[12238]_ ;
  assign \new_[12240]_  = \new_[12239]_  & \new_[12234]_ ;
  assign \new_[12243]_  = A199 & A169;
  assign \new_[12246]_  = ~A201 & A200;
  assign \new_[12247]_  = \new_[12246]_  & \new_[12243]_ ;
  assign \new_[12250]_  = A233 & ~A202;
  assign \new_[12254]_  = A300 & A298;
  assign \new_[12255]_  = A234 & \new_[12254]_ ;
  assign \new_[12256]_  = \new_[12255]_  & \new_[12250]_ ;
  assign \new_[12259]_  = A199 & A169;
  assign \new_[12262]_  = ~A201 & A200;
  assign \new_[12263]_  = \new_[12262]_  & \new_[12259]_ ;
  assign \new_[12266]_  = A233 & ~A202;
  assign \new_[12270]_  = A267 & A265;
  assign \new_[12271]_  = A234 & \new_[12270]_ ;
  assign \new_[12272]_  = \new_[12271]_  & \new_[12266]_ ;
  assign \new_[12275]_  = A199 & A169;
  assign \new_[12278]_  = ~A201 & A200;
  assign \new_[12279]_  = \new_[12278]_  & \new_[12275]_ ;
  assign \new_[12282]_  = A233 & ~A202;
  assign \new_[12286]_  = A267 & A266;
  assign \new_[12287]_  = A234 & \new_[12286]_ ;
  assign \new_[12288]_  = \new_[12287]_  & \new_[12282]_ ;
  assign \new_[12291]_  = A199 & A169;
  assign \new_[12294]_  = ~A201 & A200;
  assign \new_[12295]_  = \new_[12294]_  & \new_[12291]_ ;
  assign \new_[12298]_  = ~A232 & ~A202;
  assign \new_[12302]_  = A301 & A236;
  assign \new_[12303]_  = A233 & \new_[12302]_ ;
  assign \new_[12304]_  = \new_[12303]_  & \new_[12298]_ ;
  assign \new_[12307]_  = A199 & A169;
  assign \new_[12310]_  = ~A201 & A200;
  assign \new_[12311]_  = \new_[12310]_  & \new_[12307]_ ;
  assign \new_[12314]_  = ~A232 & ~A202;
  assign \new_[12318]_  = A268 & A236;
  assign \new_[12319]_  = A233 & \new_[12318]_ ;
  assign \new_[12320]_  = \new_[12319]_  & \new_[12314]_ ;
  assign \new_[12323]_  = A199 & A169;
  assign \new_[12326]_  = ~A201 & A200;
  assign \new_[12327]_  = \new_[12326]_  & \new_[12323]_ ;
  assign \new_[12330]_  = A232 & ~A202;
  assign \new_[12334]_  = A301 & A236;
  assign \new_[12335]_  = ~A233 & \new_[12334]_ ;
  assign \new_[12336]_  = \new_[12335]_  & \new_[12330]_ ;
  assign \new_[12339]_  = A199 & A169;
  assign \new_[12342]_  = ~A201 & A200;
  assign \new_[12343]_  = \new_[12342]_  & \new_[12339]_ ;
  assign \new_[12346]_  = A232 & ~A202;
  assign \new_[12350]_  = A268 & A236;
  assign \new_[12351]_  = ~A233 & \new_[12350]_ ;
  assign \new_[12352]_  = \new_[12351]_  & \new_[12346]_ ;
  assign \new_[12355]_  = ~A199 & A169;
  assign \new_[12358]_  = ~A202 & ~A200;
  assign \new_[12359]_  = \new_[12358]_  & \new_[12355]_ ;
  assign \new_[12362]_  = A234 & A232;
  assign \new_[12366]_  = A302 & ~A299;
  assign \new_[12367]_  = A298 & \new_[12366]_ ;
  assign \new_[12368]_  = \new_[12367]_  & \new_[12362]_ ;
  assign \new_[12371]_  = ~A199 & A169;
  assign \new_[12374]_  = ~A202 & ~A200;
  assign \new_[12375]_  = \new_[12374]_  & \new_[12371]_ ;
  assign \new_[12378]_  = A234 & A232;
  assign \new_[12382]_  = A302 & A299;
  assign \new_[12383]_  = ~A298 & \new_[12382]_ ;
  assign \new_[12384]_  = \new_[12383]_  & \new_[12378]_ ;
  assign \new_[12387]_  = ~A199 & A169;
  assign \new_[12390]_  = ~A202 & ~A200;
  assign \new_[12391]_  = \new_[12390]_  & \new_[12387]_ ;
  assign \new_[12394]_  = A234 & A232;
  assign \new_[12398]_  = A269 & A266;
  assign \new_[12399]_  = ~A265 & \new_[12398]_ ;
  assign \new_[12400]_  = \new_[12399]_  & \new_[12394]_ ;
  assign \new_[12403]_  = ~A199 & A169;
  assign \new_[12406]_  = ~A202 & ~A200;
  assign \new_[12407]_  = \new_[12406]_  & \new_[12403]_ ;
  assign \new_[12410]_  = A234 & A232;
  assign \new_[12414]_  = A269 & ~A266;
  assign \new_[12415]_  = A265 & \new_[12414]_ ;
  assign \new_[12416]_  = \new_[12415]_  & \new_[12410]_ ;
  assign \new_[12419]_  = ~A199 & A169;
  assign \new_[12422]_  = ~A202 & ~A200;
  assign \new_[12423]_  = \new_[12422]_  & \new_[12419]_ ;
  assign \new_[12426]_  = A234 & A233;
  assign \new_[12430]_  = A302 & ~A299;
  assign \new_[12431]_  = A298 & \new_[12430]_ ;
  assign \new_[12432]_  = \new_[12431]_  & \new_[12426]_ ;
  assign \new_[12435]_  = ~A199 & A169;
  assign \new_[12438]_  = ~A202 & ~A200;
  assign \new_[12439]_  = \new_[12438]_  & \new_[12435]_ ;
  assign \new_[12442]_  = A234 & A233;
  assign \new_[12446]_  = A302 & A299;
  assign \new_[12447]_  = ~A298 & \new_[12446]_ ;
  assign \new_[12448]_  = \new_[12447]_  & \new_[12442]_ ;
  assign \new_[12451]_  = ~A199 & A169;
  assign \new_[12454]_  = ~A202 & ~A200;
  assign \new_[12455]_  = \new_[12454]_  & \new_[12451]_ ;
  assign \new_[12458]_  = A234 & A233;
  assign \new_[12462]_  = A269 & A266;
  assign \new_[12463]_  = ~A265 & \new_[12462]_ ;
  assign \new_[12464]_  = \new_[12463]_  & \new_[12458]_ ;
  assign \new_[12467]_  = ~A199 & A169;
  assign \new_[12470]_  = ~A202 & ~A200;
  assign \new_[12471]_  = \new_[12470]_  & \new_[12467]_ ;
  assign \new_[12474]_  = A234 & A233;
  assign \new_[12478]_  = A269 & ~A266;
  assign \new_[12479]_  = A265 & \new_[12478]_ ;
  assign \new_[12480]_  = \new_[12479]_  & \new_[12474]_ ;
  assign \new_[12483]_  = ~A199 & A169;
  assign \new_[12486]_  = ~A202 & ~A200;
  assign \new_[12487]_  = \new_[12486]_  & \new_[12483]_ ;
  assign \new_[12490]_  = A233 & ~A232;
  assign \new_[12494]_  = A300 & A299;
  assign \new_[12495]_  = A236 & \new_[12494]_ ;
  assign \new_[12496]_  = \new_[12495]_  & \new_[12490]_ ;
  assign \new_[12499]_  = ~A199 & A169;
  assign \new_[12502]_  = ~A202 & ~A200;
  assign \new_[12503]_  = \new_[12502]_  & \new_[12499]_ ;
  assign \new_[12506]_  = A233 & ~A232;
  assign \new_[12510]_  = A300 & A298;
  assign \new_[12511]_  = A236 & \new_[12510]_ ;
  assign \new_[12512]_  = \new_[12511]_  & \new_[12506]_ ;
  assign \new_[12515]_  = ~A199 & A169;
  assign \new_[12518]_  = ~A202 & ~A200;
  assign \new_[12519]_  = \new_[12518]_  & \new_[12515]_ ;
  assign \new_[12522]_  = A233 & ~A232;
  assign \new_[12526]_  = A267 & A265;
  assign \new_[12527]_  = A236 & \new_[12526]_ ;
  assign \new_[12528]_  = \new_[12527]_  & \new_[12522]_ ;
  assign \new_[12531]_  = ~A199 & A169;
  assign \new_[12534]_  = ~A202 & ~A200;
  assign \new_[12535]_  = \new_[12534]_  & \new_[12531]_ ;
  assign \new_[12538]_  = A233 & ~A232;
  assign \new_[12542]_  = A267 & A266;
  assign \new_[12543]_  = A236 & \new_[12542]_ ;
  assign \new_[12544]_  = \new_[12543]_  & \new_[12538]_ ;
  assign \new_[12547]_  = ~A199 & A169;
  assign \new_[12550]_  = ~A202 & ~A200;
  assign \new_[12551]_  = \new_[12550]_  & \new_[12547]_ ;
  assign \new_[12554]_  = ~A233 & A232;
  assign \new_[12558]_  = A300 & A299;
  assign \new_[12559]_  = A236 & \new_[12558]_ ;
  assign \new_[12560]_  = \new_[12559]_  & \new_[12554]_ ;
  assign \new_[12563]_  = ~A199 & A169;
  assign \new_[12566]_  = ~A202 & ~A200;
  assign \new_[12567]_  = \new_[12566]_  & \new_[12563]_ ;
  assign \new_[12570]_  = ~A233 & A232;
  assign \new_[12574]_  = A300 & A298;
  assign \new_[12575]_  = A236 & \new_[12574]_ ;
  assign \new_[12576]_  = \new_[12575]_  & \new_[12570]_ ;
  assign \new_[12579]_  = ~A199 & A169;
  assign \new_[12582]_  = ~A202 & ~A200;
  assign \new_[12583]_  = \new_[12582]_  & \new_[12579]_ ;
  assign \new_[12586]_  = ~A233 & A232;
  assign \new_[12590]_  = A267 & A265;
  assign \new_[12591]_  = A236 & \new_[12590]_ ;
  assign \new_[12592]_  = \new_[12591]_  & \new_[12586]_ ;
  assign \new_[12595]_  = ~A199 & A169;
  assign \new_[12598]_  = ~A202 & ~A200;
  assign \new_[12599]_  = \new_[12598]_  & \new_[12595]_ ;
  assign \new_[12602]_  = ~A233 & A232;
  assign \new_[12606]_  = A267 & A266;
  assign \new_[12607]_  = A236 & \new_[12606]_ ;
  assign \new_[12608]_  = \new_[12607]_  & \new_[12602]_ ;
  assign \new_[12611]_  = ~A167 & ~A169;
  assign \new_[12614]_  = A202 & ~A166;
  assign \new_[12615]_  = \new_[12614]_  & \new_[12611]_ ;
  assign \new_[12618]_  = A234 & A232;
  assign \new_[12622]_  = A302 & ~A299;
  assign \new_[12623]_  = A298 & \new_[12622]_ ;
  assign \new_[12624]_  = \new_[12623]_  & \new_[12618]_ ;
  assign \new_[12627]_  = ~A167 & ~A169;
  assign \new_[12630]_  = A202 & ~A166;
  assign \new_[12631]_  = \new_[12630]_  & \new_[12627]_ ;
  assign \new_[12634]_  = A234 & A232;
  assign \new_[12638]_  = A302 & A299;
  assign \new_[12639]_  = ~A298 & \new_[12638]_ ;
  assign \new_[12640]_  = \new_[12639]_  & \new_[12634]_ ;
  assign \new_[12643]_  = ~A167 & ~A169;
  assign \new_[12646]_  = A202 & ~A166;
  assign \new_[12647]_  = \new_[12646]_  & \new_[12643]_ ;
  assign \new_[12650]_  = A234 & A232;
  assign \new_[12654]_  = A269 & A266;
  assign \new_[12655]_  = ~A265 & \new_[12654]_ ;
  assign \new_[12656]_  = \new_[12655]_  & \new_[12650]_ ;
  assign \new_[12659]_  = ~A167 & ~A169;
  assign \new_[12662]_  = A202 & ~A166;
  assign \new_[12663]_  = \new_[12662]_  & \new_[12659]_ ;
  assign \new_[12666]_  = A234 & A232;
  assign \new_[12670]_  = A269 & ~A266;
  assign \new_[12671]_  = A265 & \new_[12670]_ ;
  assign \new_[12672]_  = \new_[12671]_  & \new_[12666]_ ;
  assign \new_[12675]_  = ~A167 & ~A169;
  assign \new_[12678]_  = A202 & ~A166;
  assign \new_[12679]_  = \new_[12678]_  & \new_[12675]_ ;
  assign \new_[12682]_  = A234 & A233;
  assign \new_[12686]_  = A302 & ~A299;
  assign \new_[12687]_  = A298 & \new_[12686]_ ;
  assign \new_[12688]_  = \new_[12687]_  & \new_[12682]_ ;
  assign \new_[12691]_  = ~A167 & ~A169;
  assign \new_[12694]_  = A202 & ~A166;
  assign \new_[12695]_  = \new_[12694]_  & \new_[12691]_ ;
  assign \new_[12698]_  = A234 & A233;
  assign \new_[12702]_  = A302 & A299;
  assign \new_[12703]_  = ~A298 & \new_[12702]_ ;
  assign \new_[12704]_  = \new_[12703]_  & \new_[12698]_ ;
  assign \new_[12707]_  = ~A167 & ~A169;
  assign \new_[12710]_  = A202 & ~A166;
  assign \new_[12711]_  = \new_[12710]_  & \new_[12707]_ ;
  assign \new_[12714]_  = A234 & A233;
  assign \new_[12718]_  = A269 & A266;
  assign \new_[12719]_  = ~A265 & \new_[12718]_ ;
  assign \new_[12720]_  = \new_[12719]_  & \new_[12714]_ ;
  assign \new_[12723]_  = ~A167 & ~A169;
  assign \new_[12726]_  = A202 & ~A166;
  assign \new_[12727]_  = \new_[12726]_  & \new_[12723]_ ;
  assign \new_[12730]_  = A234 & A233;
  assign \new_[12734]_  = A269 & ~A266;
  assign \new_[12735]_  = A265 & \new_[12734]_ ;
  assign \new_[12736]_  = \new_[12735]_  & \new_[12730]_ ;
  assign \new_[12739]_  = ~A167 & ~A169;
  assign \new_[12742]_  = A202 & ~A166;
  assign \new_[12743]_  = \new_[12742]_  & \new_[12739]_ ;
  assign \new_[12746]_  = A233 & ~A232;
  assign \new_[12750]_  = A300 & A299;
  assign \new_[12751]_  = A236 & \new_[12750]_ ;
  assign \new_[12752]_  = \new_[12751]_  & \new_[12746]_ ;
  assign \new_[12755]_  = ~A167 & ~A169;
  assign \new_[12758]_  = A202 & ~A166;
  assign \new_[12759]_  = \new_[12758]_  & \new_[12755]_ ;
  assign \new_[12762]_  = A233 & ~A232;
  assign \new_[12766]_  = A300 & A298;
  assign \new_[12767]_  = A236 & \new_[12766]_ ;
  assign \new_[12768]_  = \new_[12767]_  & \new_[12762]_ ;
  assign \new_[12771]_  = ~A167 & ~A169;
  assign \new_[12774]_  = A202 & ~A166;
  assign \new_[12775]_  = \new_[12774]_  & \new_[12771]_ ;
  assign \new_[12778]_  = A233 & ~A232;
  assign \new_[12782]_  = A267 & A265;
  assign \new_[12783]_  = A236 & \new_[12782]_ ;
  assign \new_[12784]_  = \new_[12783]_  & \new_[12778]_ ;
  assign \new_[12787]_  = ~A167 & ~A169;
  assign \new_[12790]_  = A202 & ~A166;
  assign \new_[12791]_  = \new_[12790]_  & \new_[12787]_ ;
  assign \new_[12794]_  = A233 & ~A232;
  assign \new_[12798]_  = A267 & A266;
  assign \new_[12799]_  = A236 & \new_[12798]_ ;
  assign \new_[12800]_  = \new_[12799]_  & \new_[12794]_ ;
  assign \new_[12803]_  = ~A167 & ~A169;
  assign \new_[12806]_  = A202 & ~A166;
  assign \new_[12807]_  = \new_[12806]_  & \new_[12803]_ ;
  assign \new_[12810]_  = ~A233 & A232;
  assign \new_[12814]_  = A300 & A299;
  assign \new_[12815]_  = A236 & \new_[12814]_ ;
  assign \new_[12816]_  = \new_[12815]_  & \new_[12810]_ ;
  assign \new_[12819]_  = ~A167 & ~A169;
  assign \new_[12822]_  = A202 & ~A166;
  assign \new_[12823]_  = \new_[12822]_  & \new_[12819]_ ;
  assign \new_[12826]_  = ~A233 & A232;
  assign \new_[12830]_  = A300 & A298;
  assign \new_[12831]_  = A236 & \new_[12830]_ ;
  assign \new_[12832]_  = \new_[12831]_  & \new_[12826]_ ;
  assign \new_[12835]_  = ~A167 & ~A169;
  assign \new_[12838]_  = A202 & ~A166;
  assign \new_[12839]_  = \new_[12838]_  & \new_[12835]_ ;
  assign \new_[12842]_  = ~A233 & A232;
  assign \new_[12846]_  = A267 & A265;
  assign \new_[12847]_  = A236 & \new_[12846]_ ;
  assign \new_[12848]_  = \new_[12847]_  & \new_[12842]_ ;
  assign \new_[12851]_  = ~A167 & ~A169;
  assign \new_[12854]_  = A202 & ~A166;
  assign \new_[12855]_  = \new_[12854]_  & \new_[12851]_ ;
  assign \new_[12858]_  = ~A233 & A232;
  assign \new_[12862]_  = A267 & A266;
  assign \new_[12863]_  = A236 & \new_[12862]_ ;
  assign \new_[12864]_  = \new_[12863]_  & \new_[12858]_ ;
  assign \new_[12867]_  = ~A167 & ~A169;
  assign \new_[12870]_  = A199 & ~A166;
  assign \new_[12871]_  = \new_[12870]_  & \new_[12867]_ ;
  assign \new_[12874]_  = A235 & A201;
  assign \new_[12878]_  = A302 & ~A299;
  assign \new_[12879]_  = A298 & \new_[12878]_ ;
  assign \new_[12880]_  = \new_[12879]_  & \new_[12874]_ ;
  assign \new_[12883]_  = ~A167 & ~A169;
  assign \new_[12886]_  = A199 & ~A166;
  assign \new_[12887]_  = \new_[12886]_  & \new_[12883]_ ;
  assign \new_[12890]_  = A235 & A201;
  assign \new_[12894]_  = A302 & A299;
  assign \new_[12895]_  = ~A298 & \new_[12894]_ ;
  assign \new_[12896]_  = \new_[12895]_  & \new_[12890]_ ;
  assign \new_[12899]_  = ~A167 & ~A169;
  assign \new_[12902]_  = A199 & ~A166;
  assign \new_[12903]_  = \new_[12902]_  & \new_[12899]_ ;
  assign \new_[12906]_  = A235 & A201;
  assign \new_[12910]_  = A269 & A266;
  assign \new_[12911]_  = ~A265 & \new_[12910]_ ;
  assign \new_[12912]_  = \new_[12911]_  & \new_[12906]_ ;
  assign \new_[12915]_  = ~A167 & ~A169;
  assign \new_[12918]_  = A199 & ~A166;
  assign \new_[12919]_  = \new_[12918]_  & \new_[12915]_ ;
  assign \new_[12922]_  = A235 & A201;
  assign \new_[12926]_  = A269 & ~A266;
  assign \new_[12927]_  = A265 & \new_[12926]_ ;
  assign \new_[12928]_  = \new_[12927]_  & \new_[12922]_ ;
  assign \new_[12931]_  = ~A167 & ~A169;
  assign \new_[12934]_  = A199 & ~A166;
  assign \new_[12935]_  = \new_[12934]_  & \new_[12931]_ ;
  assign \new_[12938]_  = A232 & A201;
  assign \new_[12942]_  = A300 & A299;
  assign \new_[12943]_  = A234 & \new_[12942]_ ;
  assign \new_[12944]_  = \new_[12943]_  & \new_[12938]_ ;
  assign \new_[12947]_  = ~A167 & ~A169;
  assign \new_[12950]_  = A199 & ~A166;
  assign \new_[12951]_  = \new_[12950]_  & \new_[12947]_ ;
  assign \new_[12954]_  = A232 & A201;
  assign \new_[12958]_  = A300 & A298;
  assign \new_[12959]_  = A234 & \new_[12958]_ ;
  assign \new_[12960]_  = \new_[12959]_  & \new_[12954]_ ;
  assign \new_[12963]_  = ~A167 & ~A169;
  assign \new_[12966]_  = A199 & ~A166;
  assign \new_[12967]_  = \new_[12966]_  & \new_[12963]_ ;
  assign \new_[12970]_  = A232 & A201;
  assign \new_[12974]_  = A267 & A265;
  assign \new_[12975]_  = A234 & \new_[12974]_ ;
  assign \new_[12976]_  = \new_[12975]_  & \new_[12970]_ ;
  assign \new_[12979]_  = ~A167 & ~A169;
  assign \new_[12982]_  = A199 & ~A166;
  assign \new_[12983]_  = \new_[12982]_  & \new_[12979]_ ;
  assign \new_[12986]_  = A232 & A201;
  assign \new_[12990]_  = A267 & A266;
  assign \new_[12991]_  = A234 & \new_[12990]_ ;
  assign \new_[12992]_  = \new_[12991]_  & \new_[12986]_ ;
  assign \new_[12995]_  = ~A167 & ~A169;
  assign \new_[12998]_  = A199 & ~A166;
  assign \new_[12999]_  = \new_[12998]_  & \new_[12995]_ ;
  assign \new_[13002]_  = A233 & A201;
  assign \new_[13006]_  = A300 & A299;
  assign \new_[13007]_  = A234 & \new_[13006]_ ;
  assign \new_[13008]_  = \new_[13007]_  & \new_[13002]_ ;
  assign \new_[13011]_  = ~A167 & ~A169;
  assign \new_[13014]_  = A199 & ~A166;
  assign \new_[13015]_  = \new_[13014]_  & \new_[13011]_ ;
  assign \new_[13018]_  = A233 & A201;
  assign \new_[13022]_  = A300 & A298;
  assign \new_[13023]_  = A234 & \new_[13022]_ ;
  assign \new_[13024]_  = \new_[13023]_  & \new_[13018]_ ;
  assign \new_[13027]_  = ~A167 & ~A169;
  assign \new_[13030]_  = A199 & ~A166;
  assign \new_[13031]_  = \new_[13030]_  & \new_[13027]_ ;
  assign \new_[13034]_  = A233 & A201;
  assign \new_[13038]_  = A267 & A265;
  assign \new_[13039]_  = A234 & \new_[13038]_ ;
  assign \new_[13040]_  = \new_[13039]_  & \new_[13034]_ ;
  assign \new_[13043]_  = ~A167 & ~A169;
  assign \new_[13046]_  = A199 & ~A166;
  assign \new_[13047]_  = \new_[13046]_  & \new_[13043]_ ;
  assign \new_[13050]_  = A233 & A201;
  assign \new_[13054]_  = A267 & A266;
  assign \new_[13055]_  = A234 & \new_[13054]_ ;
  assign \new_[13056]_  = \new_[13055]_  & \new_[13050]_ ;
  assign \new_[13059]_  = ~A167 & ~A169;
  assign \new_[13062]_  = A199 & ~A166;
  assign \new_[13063]_  = \new_[13062]_  & \new_[13059]_ ;
  assign \new_[13066]_  = ~A232 & A201;
  assign \new_[13070]_  = A301 & A236;
  assign \new_[13071]_  = A233 & \new_[13070]_ ;
  assign \new_[13072]_  = \new_[13071]_  & \new_[13066]_ ;
  assign \new_[13075]_  = ~A167 & ~A169;
  assign \new_[13078]_  = A199 & ~A166;
  assign \new_[13079]_  = \new_[13078]_  & \new_[13075]_ ;
  assign \new_[13082]_  = ~A232 & A201;
  assign \new_[13086]_  = A268 & A236;
  assign \new_[13087]_  = A233 & \new_[13086]_ ;
  assign \new_[13088]_  = \new_[13087]_  & \new_[13082]_ ;
  assign \new_[13091]_  = ~A167 & ~A169;
  assign \new_[13094]_  = A199 & ~A166;
  assign \new_[13095]_  = \new_[13094]_  & \new_[13091]_ ;
  assign \new_[13098]_  = A232 & A201;
  assign \new_[13102]_  = A301 & A236;
  assign \new_[13103]_  = ~A233 & \new_[13102]_ ;
  assign \new_[13104]_  = \new_[13103]_  & \new_[13098]_ ;
  assign \new_[13107]_  = ~A167 & ~A169;
  assign \new_[13110]_  = A199 & ~A166;
  assign \new_[13111]_  = \new_[13110]_  & \new_[13107]_ ;
  assign \new_[13114]_  = A232 & A201;
  assign \new_[13118]_  = A268 & A236;
  assign \new_[13119]_  = ~A233 & \new_[13118]_ ;
  assign \new_[13120]_  = \new_[13119]_  & \new_[13114]_ ;
  assign \new_[13123]_  = ~A167 & ~A169;
  assign \new_[13126]_  = A200 & ~A166;
  assign \new_[13127]_  = \new_[13126]_  & \new_[13123]_ ;
  assign \new_[13130]_  = A235 & A201;
  assign \new_[13134]_  = A302 & ~A299;
  assign \new_[13135]_  = A298 & \new_[13134]_ ;
  assign \new_[13136]_  = \new_[13135]_  & \new_[13130]_ ;
  assign \new_[13139]_  = ~A167 & ~A169;
  assign \new_[13142]_  = A200 & ~A166;
  assign \new_[13143]_  = \new_[13142]_  & \new_[13139]_ ;
  assign \new_[13146]_  = A235 & A201;
  assign \new_[13150]_  = A302 & A299;
  assign \new_[13151]_  = ~A298 & \new_[13150]_ ;
  assign \new_[13152]_  = \new_[13151]_  & \new_[13146]_ ;
  assign \new_[13155]_  = ~A167 & ~A169;
  assign \new_[13158]_  = A200 & ~A166;
  assign \new_[13159]_  = \new_[13158]_  & \new_[13155]_ ;
  assign \new_[13162]_  = A235 & A201;
  assign \new_[13166]_  = A269 & A266;
  assign \new_[13167]_  = ~A265 & \new_[13166]_ ;
  assign \new_[13168]_  = \new_[13167]_  & \new_[13162]_ ;
  assign \new_[13171]_  = ~A167 & ~A169;
  assign \new_[13174]_  = A200 & ~A166;
  assign \new_[13175]_  = \new_[13174]_  & \new_[13171]_ ;
  assign \new_[13178]_  = A235 & A201;
  assign \new_[13182]_  = A269 & ~A266;
  assign \new_[13183]_  = A265 & \new_[13182]_ ;
  assign \new_[13184]_  = \new_[13183]_  & \new_[13178]_ ;
  assign \new_[13187]_  = ~A167 & ~A169;
  assign \new_[13190]_  = A200 & ~A166;
  assign \new_[13191]_  = \new_[13190]_  & \new_[13187]_ ;
  assign \new_[13194]_  = A232 & A201;
  assign \new_[13198]_  = A300 & A299;
  assign \new_[13199]_  = A234 & \new_[13198]_ ;
  assign \new_[13200]_  = \new_[13199]_  & \new_[13194]_ ;
  assign \new_[13203]_  = ~A167 & ~A169;
  assign \new_[13206]_  = A200 & ~A166;
  assign \new_[13207]_  = \new_[13206]_  & \new_[13203]_ ;
  assign \new_[13210]_  = A232 & A201;
  assign \new_[13214]_  = A300 & A298;
  assign \new_[13215]_  = A234 & \new_[13214]_ ;
  assign \new_[13216]_  = \new_[13215]_  & \new_[13210]_ ;
  assign \new_[13219]_  = ~A167 & ~A169;
  assign \new_[13222]_  = A200 & ~A166;
  assign \new_[13223]_  = \new_[13222]_  & \new_[13219]_ ;
  assign \new_[13226]_  = A232 & A201;
  assign \new_[13230]_  = A267 & A265;
  assign \new_[13231]_  = A234 & \new_[13230]_ ;
  assign \new_[13232]_  = \new_[13231]_  & \new_[13226]_ ;
  assign \new_[13235]_  = ~A167 & ~A169;
  assign \new_[13238]_  = A200 & ~A166;
  assign \new_[13239]_  = \new_[13238]_  & \new_[13235]_ ;
  assign \new_[13242]_  = A232 & A201;
  assign \new_[13246]_  = A267 & A266;
  assign \new_[13247]_  = A234 & \new_[13246]_ ;
  assign \new_[13248]_  = \new_[13247]_  & \new_[13242]_ ;
  assign \new_[13251]_  = ~A167 & ~A169;
  assign \new_[13254]_  = A200 & ~A166;
  assign \new_[13255]_  = \new_[13254]_  & \new_[13251]_ ;
  assign \new_[13258]_  = A233 & A201;
  assign \new_[13262]_  = A300 & A299;
  assign \new_[13263]_  = A234 & \new_[13262]_ ;
  assign \new_[13264]_  = \new_[13263]_  & \new_[13258]_ ;
  assign \new_[13267]_  = ~A167 & ~A169;
  assign \new_[13270]_  = A200 & ~A166;
  assign \new_[13271]_  = \new_[13270]_  & \new_[13267]_ ;
  assign \new_[13274]_  = A233 & A201;
  assign \new_[13278]_  = A300 & A298;
  assign \new_[13279]_  = A234 & \new_[13278]_ ;
  assign \new_[13280]_  = \new_[13279]_  & \new_[13274]_ ;
  assign \new_[13283]_  = ~A167 & ~A169;
  assign \new_[13286]_  = A200 & ~A166;
  assign \new_[13287]_  = \new_[13286]_  & \new_[13283]_ ;
  assign \new_[13290]_  = A233 & A201;
  assign \new_[13294]_  = A267 & A265;
  assign \new_[13295]_  = A234 & \new_[13294]_ ;
  assign \new_[13296]_  = \new_[13295]_  & \new_[13290]_ ;
  assign \new_[13299]_  = ~A167 & ~A169;
  assign \new_[13302]_  = A200 & ~A166;
  assign \new_[13303]_  = \new_[13302]_  & \new_[13299]_ ;
  assign \new_[13306]_  = A233 & A201;
  assign \new_[13310]_  = A267 & A266;
  assign \new_[13311]_  = A234 & \new_[13310]_ ;
  assign \new_[13312]_  = \new_[13311]_  & \new_[13306]_ ;
  assign \new_[13315]_  = ~A167 & ~A169;
  assign \new_[13318]_  = A200 & ~A166;
  assign \new_[13319]_  = \new_[13318]_  & \new_[13315]_ ;
  assign \new_[13322]_  = ~A232 & A201;
  assign \new_[13326]_  = A301 & A236;
  assign \new_[13327]_  = A233 & \new_[13326]_ ;
  assign \new_[13328]_  = \new_[13327]_  & \new_[13322]_ ;
  assign \new_[13331]_  = ~A167 & ~A169;
  assign \new_[13334]_  = A200 & ~A166;
  assign \new_[13335]_  = \new_[13334]_  & \new_[13331]_ ;
  assign \new_[13338]_  = ~A232 & A201;
  assign \new_[13342]_  = A268 & A236;
  assign \new_[13343]_  = A233 & \new_[13342]_ ;
  assign \new_[13344]_  = \new_[13343]_  & \new_[13338]_ ;
  assign \new_[13347]_  = ~A167 & ~A169;
  assign \new_[13350]_  = A200 & ~A166;
  assign \new_[13351]_  = \new_[13350]_  & \new_[13347]_ ;
  assign \new_[13354]_  = A232 & A201;
  assign \new_[13358]_  = A301 & A236;
  assign \new_[13359]_  = ~A233 & \new_[13358]_ ;
  assign \new_[13360]_  = \new_[13359]_  & \new_[13354]_ ;
  assign \new_[13363]_  = ~A167 & ~A169;
  assign \new_[13366]_  = A200 & ~A166;
  assign \new_[13367]_  = \new_[13366]_  & \new_[13363]_ ;
  assign \new_[13370]_  = A232 & A201;
  assign \new_[13374]_  = A268 & A236;
  assign \new_[13375]_  = ~A233 & \new_[13374]_ ;
  assign \new_[13376]_  = \new_[13375]_  & \new_[13370]_ ;
  assign \new_[13379]_  = ~A167 & ~A169;
  assign \new_[13382]_  = ~A199 & ~A166;
  assign \new_[13383]_  = \new_[13382]_  & \new_[13379]_ ;
  assign \new_[13386]_  = A203 & A200;
  assign \new_[13390]_  = A300 & A299;
  assign \new_[13391]_  = A235 & \new_[13390]_ ;
  assign \new_[13392]_  = \new_[13391]_  & \new_[13386]_ ;
  assign \new_[13395]_  = ~A167 & ~A169;
  assign \new_[13398]_  = ~A199 & ~A166;
  assign \new_[13399]_  = \new_[13398]_  & \new_[13395]_ ;
  assign \new_[13402]_  = A203 & A200;
  assign \new_[13406]_  = A300 & A298;
  assign \new_[13407]_  = A235 & \new_[13406]_ ;
  assign \new_[13408]_  = \new_[13407]_  & \new_[13402]_ ;
  assign \new_[13411]_  = ~A167 & ~A169;
  assign \new_[13414]_  = ~A199 & ~A166;
  assign \new_[13415]_  = \new_[13414]_  & \new_[13411]_ ;
  assign \new_[13418]_  = A203 & A200;
  assign \new_[13422]_  = A267 & A265;
  assign \new_[13423]_  = A235 & \new_[13422]_ ;
  assign \new_[13424]_  = \new_[13423]_  & \new_[13418]_ ;
  assign \new_[13427]_  = ~A167 & ~A169;
  assign \new_[13430]_  = ~A199 & ~A166;
  assign \new_[13431]_  = \new_[13430]_  & \new_[13427]_ ;
  assign \new_[13434]_  = A203 & A200;
  assign \new_[13438]_  = A267 & A266;
  assign \new_[13439]_  = A235 & \new_[13438]_ ;
  assign \new_[13440]_  = \new_[13439]_  & \new_[13434]_ ;
  assign \new_[13443]_  = ~A167 & ~A169;
  assign \new_[13446]_  = ~A199 & ~A166;
  assign \new_[13447]_  = \new_[13446]_  & \new_[13443]_ ;
  assign \new_[13450]_  = A203 & A200;
  assign \new_[13454]_  = A301 & A234;
  assign \new_[13455]_  = A232 & \new_[13454]_ ;
  assign \new_[13456]_  = \new_[13455]_  & \new_[13450]_ ;
  assign \new_[13459]_  = ~A167 & ~A169;
  assign \new_[13462]_  = ~A199 & ~A166;
  assign \new_[13463]_  = \new_[13462]_  & \new_[13459]_ ;
  assign \new_[13466]_  = A203 & A200;
  assign \new_[13470]_  = A268 & A234;
  assign \new_[13471]_  = A232 & \new_[13470]_ ;
  assign \new_[13472]_  = \new_[13471]_  & \new_[13466]_ ;
  assign \new_[13475]_  = ~A167 & ~A169;
  assign \new_[13478]_  = ~A199 & ~A166;
  assign \new_[13479]_  = \new_[13478]_  & \new_[13475]_ ;
  assign \new_[13482]_  = A203 & A200;
  assign \new_[13486]_  = A301 & A234;
  assign \new_[13487]_  = A233 & \new_[13486]_ ;
  assign \new_[13488]_  = \new_[13487]_  & \new_[13482]_ ;
  assign \new_[13491]_  = ~A167 & ~A169;
  assign \new_[13494]_  = ~A199 & ~A166;
  assign \new_[13495]_  = \new_[13494]_  & \new_[13491]_ ;
  assign \new_[13498]_  = A203 & A200;
  assign \new_[13502]_  = A268 & A234;
  assign \new_[13503]_  = A233 & \new_[13502]_ ;
  assign \new_[13504]_  = \new_[13503]_  & \new_[13498]_ ;
  assign \new_[13507]_  = ~A167 & ~A169;
  assign \new_[13510]_  = A199 & ~A166;
  assign \new_[13511]_  = \new_[13510]_  & \new_[13507]_ ;
  assign \new_[13514]_  = A203 & ~A200;
  assign \new_[13518]_  = A300 & A299;
  assign \new_[13519]_  = A235 & \new_[13518]_ ;
  assign \new_[13520]_  = \new_[13519]_  & \new_[13514]_ ;
  assign \new_[13523]_  = ~A167 & ~A169;
  assign \new_[13526]_  = A199 & ~A166;
  assign \new_[13527]_  = \new_[13526]_  & \new_[13523]_ ;
  assign \new_[13530]_  = A203 & ~A200;
  assign \new_[13534]_  = A300 & A298;
  assign \new_[13535]_  = A235 & \new_[13534]_ ;
  assign \new_[13536]_  = \new_[13535]_  & \new_[13530]_ ;
  assign \new_[13539]_  = ~A167 & ~A169;
  assign \new_[13542]_  = A199 & ~A166;
  assign \new_[13543]_  = \new_[13542]_  & \new_[13539]_ ;
  assign \new_[13546]_  = A203 & ~A200;
  assign \new_[13550]_  = A267 & A265;
  assign \new_[13551]_  = A235 & \new_[13550]_ ;
  assign \new_[13552]_  = \new_[13551]_  & \new_[13546]_ ;
  assign \new_[13555]_  = ~A167 & ~A169;
  assign \new_[13558]_  = A199 & ~A166;
  assign \new_[13559]_  = \new_[13558]_  & \new_[13555]_ ;
  assign \new_[13562]_  = A203 & ~A200;
  assign \new_[13566]_  = A267 & A266;
  assign \new_[13567]_  = A235 & \new_[13566]_ ;
  assign \new_[13568]_  = \new_[13567]_  & \new_[13562]_ ;
  assign \new_[13571]_  = ~A167 & ~A169;
  assign \new_[13574]_  = A199 & ~A166;
  assign \new_[13575]_  = \new_[13574]_  & \new_[13571]_ ;
  assign \new_[13578]_  = A203 & ~A200;
  assign \new_[13582]_  = A301 & A234;
  assign \new_[13583]_  = A232 & \new_[13582]_ ;
  assign \new_[13584]_  = \new_[13583]_  & \new_[13578]_ ;
  assign \new_[13587]_  = ~A167 & ~A169;
  assign \new_[13590]_  = A199 & ~A166;
  assign \new_[13591]_  = \new_[13590]_  & \new_[13587]_ ;
  assign \new_[13594]_  = A203 & ~A200;
  assign \new_[13598]_  = A268 & A234;
  assign \new_[13599]_  = A232 & \new_[13598]_ ;
  assign \new_[13600]_  = \new_[13599]_  & \new_[13594]_ ;
  assign \new_[13603]_  = ~A167 & ~A169;
  assign \new_[13606]_  = A199 & ~A166;
  assign \new_[13607]_  = \new_[13606]_  & \new_[13603]_ ;
  assign \new_[13610]_  = A203 & ~A200;
  assign \new_[13614]_  = A301 & A234;
  assign \new_[13615]_  = A233 & \new_[13614]_ ;
  assign \new_[13616]_  = \new_[13615]_  & \new_[13610]_ ;
  assign \new_[13619]_  = ~A167 & ~A169;
  assign \new_[13622]_  = A199 & ~A166;
  assign \new_[13623]_  = \new_[13622]_  & \new_[13619]_ ;
  assign \new_[13626]_  = A203 & ~A200;
  assign \new_[13630]_  = A268 & A234;
  assign \new_[13631]_  = A233 & \new_[13630]_ ;
  assign \new_[13632]_  = \new_[13631]_  & \new_[13626]_ ;
  assign \new_[13635]_  = ~A168 & ~A169;
  assign \new_[13638]_  = A166 & A167;
  assign \new_[13639]_  = \new_[13638]_  & \new_[13635]_ ;
  assign \new_[13642]_  = A235 & A202;
  assign \new_[13646]_  = A302 & ~A299;
  assign \new_[13647]_  = A298 & \new_[13646]_ ;
  assign \new_[13648]_  = \new_[13647]_  & \new_[13642]_ ;
  assign \new_[13651]_  = ~A168 & ~A169;
  assign \new_[13654]_  = A166 & A167;
  assign \new_[13655]_  = \new_[13654]_  & \new_[13651]_ ;
  assign \new_[13658]_  = A235 & A202;
  assign \new_[13662]_  = A302 & A299;
  assign \new_[13663]_  = ~A298 & \new_[13662]_ ;
  assign \new_[13664]_  = \new_[13663]_  & \new_[13658]_ ;
  assign \new_[13667]_  = ~A168 & ~A169;
  assign \new_[13670]_  = A166 & A167;
  assign \new_[13671]_  = \new_[13670]_  & \new_[13667]_ ;
  assign \new_[13674]_  = A235 & A202;
  assign \new_[13678]_  = A269 & A266;
  assign \new_[13679]_  = ~A265 & \new_[13678]_ ;
  assign \new_[13680]_  = \new_[13679]_  & \new_[13674]_ ;
  assign \new_[13683]_  = ~A168 & ~A169;
  assign \new_[13686]_  = A166 & A167;
  assign \new_[13687]_  = \new_[13686]_  & \new_[13683]_ ;
  assign \new_[13690]_  = A235 & A202;
  assign \new_[13694]_  = A269 & ~A266;
  assign \new_[13695]_  = A265 & \new_[13694]_ ;
  assign \new_[13696]_  = \new_[13695]_  & \new_[13690]_ ;
  assign \new_[13699]_  = ~A168 & ~A169;
  assign \new_[13702]_  = A166 & A167;
  assign \new_[13703]_  = \new_[13702]_  & \new_[13699]_ ;
  assign \new_[13706]_  = A232 & A202;
  assign \new_[13710]_  = A300 & A299;
  assign \new_[13711]_  = A234 & \new_[13710]_ ;
  assign \new_[13712]_  = \new_[13711]_  & \new_[13706]_ ;
  assign \new_[13715]_  = ~A168 & ~A169;
  assign \new_[13718]_  = A166 & A167;
  assign \new_[13719]_  = \new_[13718]_  & \new_[13715]_ ;
  assign \new_[13722]_  = A232 & A202;
  assign \new_[13726]_  = A300 & A298;
  assign \new_[13727]_  = A234 & \new_[13726]_ ;
  assign \new_[13728]_  = \new_[13727]_  & \new_[13722]_ ;
  assign \new_[13731]_  = ~A168 & ~A169;
  assign \new_[13734]_  = A166 & A167;
  assign \new_[13735]_  = \new_[13734]_  & \new_[13731]_ ;
  assign \new_[13738]_  = A232 & A202;
  assign \new_[13742]_  = A267 & A265;
  assign \new_[13743]_  = A234 & \new_[13742]_ ;
  assign \new_[13744]_  = \new_[13743]_  & \new_[13738]_ ;
  assign \new_[13747]_  = ~A168 & ~A169;
  assign \new_[13750]_  = A166 & A167;
  assign \new_[13751]_  = \new_[13750]_  & \new_[13747]_ ;
  assign \new_[13754]_  = A232 & A202;
  assign \new_[13758]_  = A267 & A266;
  assign \new_[13759]_  = A234 & \new_[13758]_ ;
  assign \new_[13760]_  = \new_[13759]_  & \new_[13754]_ ;
  assign \new_[13763]_  = ~A168 & ~A169;
  assign \new_[13766]_  = A166 & A167;
  assign \new_[13767]_  = \new_[13766]_  & \new_[13763]_ ;
  assign \new_[13770]_  = A233 & A202;
  assign \new_[13774]_  = A300 & A299;
  assign \new_[13775]_  = A234 & \new_[13774]_ ;
  assign \new_[13776]_  = \new_[13775]_  & \new_[13770]_ ;
  assign \new_[13779]_  = ~A168 & ~A169;
  assign \new_[13782]_  = A166 & A167;
  assign \new_[13783]_  = \new_[13782]_  & \new_[13779]_ ;
  assign \new_[13786]_  = A233 & A202;
  assign \new_[13790]_  = A300 & A298;
  assign \new_[13791]_  = A234 & \new_[13790]_ ;
  assign \new_[13792]_  = \new_[13791]_  & \new_[13786]_ ;
  assign \new_[13795]_  = ~A168 & ~A169;
  assign \new_[13798]_  = A166 & A167;
  assign \new_[13799]_  = \new_[13798]_  & \new_[13795]_ ;
  assign \new_[13802]_  = A233 & A202;
  assign \new_[13806]_  = A267 & A265;
  assign \new_[13807]_  = A234 & \new_[13806]_ ;
  assign \new_[13808]_  = \new_[13807]_  & \new_[13802]_ ;
  assign \new_[13811]_  = ~A168 & ~A169;
  assign \new_[13814]_  = A166 & A167;
  assign \new_[13815]_  = \new_[13814]_  & \new_[13811]_ ;
  assign \new_[13818]_  = A233 & A202;
  assign \new_[13822]_  = A267 & A266;
  assign \new_[13823]_  = A234 & \new_[13822]_ ;
  assign \new_[13824]_  = \new_[13823]_  & \new_[13818]_ ;
  assign \new_[13827]_  = ~A168 & ~A169;
  assign \new_[13830]_  = A166 & A167;
  assign \new_[13831]_  = \new_[13830]_  & \new_[13827]_ ;
  assign \new_[13834]_  = ~A232 & A202;
  assign \new_[13838]_  = A301 & A236;
  assign \new_[13839]_  = A233 & \new_[13838]_ ;
  assign \new_[13840]_  = \new_[13839]_  & \new_[13834]_ ;
  assign \new_[13843]_  = ~A168 & ~A169;
  assign \new_[13846]_  = A166 & A167;
  assign \new_[13847]_  = \new_[13846]_  & \new_[13843]_ ;
  assign \new_[13850]_  = ~A232 & A202;
  assign \new_[13854]_  = A268 & A236;
  assign \new_[13855]_  = A233 & \new_[13854]_ ;
  assign \new_[13856]_  = \new_[13855]_  & \new_[13850]_ ;
  assign \new_[13859]_  = ~A168 & ~A169;
  assign \new_[13862]_  = A166 & A167;
  assign \new_[13863]_  = \new_[13862]_  & \new_[13859]_ ;
  assign \new_[13866]_  = A232 & A202;
  assign \new_[13870]_  = A301 & A236;
  assign \new_[13871]_  = ~A233 & \new_[13870]_ ;
  assign \new_[13872]_  = \new_[13871]_  & \new_[13866]_ ;
  assign \new_[13875]_  = ~A168 & ~A169;
  assign \new_[13878]_  = A166 & A167;
  assign \new_[13879]_  = \new_[13878]_  & \new_[13875]_ ;
  assign \new_[13882]_  = A232 & A202;
  assign \new_[13886]_  = A268 & A236;
  assign \new_[13887]_  = ~A233 & \new_[13886]_ ;
  assign \new_[13888]_  = \new_[13887]_  & \new_[13882]_ ;
  assign \new_[13891]_  = ~A168 & ~A169;
  assign \new_[13894]_  = A166 & A167;
  assign \new_[13895]_  = \new_[13894]_  & \new_[13891]_ ;
  assign \new_[13898]_  = A201 & A199;
  assign \new_[13902]_  = A300 & A299;
  assign \new_[13903]_  = A235 & \new_[13902]_ ;
  assign \new_[13904]_  = \new_[13903]_  & \new_[13898]_ ;
  assign \new_[13907]_  = ~A168 & ~A169;
  assign \new_[13910]_  = A166 & A167;
  assign \new_[13911]_  = \new_[13910]_  & \new_[13907]_ ;
  assign \new_[13914]_  = A201 & A199;
  assign \new_[13918]_  = A300 & A298;
  assign \new_[13919]_  = A235 & \new_[13918]_ ;
  assign \new_[13920]_  = \new_[13919]_  & \new_[13914]_ ;
  assign \new_[13923]_  = ~A168 & ~A169;
  assign \new_[13926]_  = A166 & A167;
  assign \new_[13927]_  = \new_[13926]_  & \new_[13923]_ ;
  assign \new_[13930]_  = A201 & A199;
  assign \new_[13934]_  = A267 & A265;
  assign \new_[13935]_  = A235 & \new_[13934]_ ;
  assign \new_[13936]_  = \new_[13935]_  & \new_[13930]_ ;
  assign \new_[13939]_  = ~A168 & ~A169;
  assign \new_[13942]_  = A166 & A167;
  assign \new_[13943]_  = \new_[13942]_  & \new_[13939]_ ;
  assign \new_[13946]_  = A201 & A199;
  assign \new_[13950]_  = A267 & A266;
  assign \new_[13951]_  = A235 & \new_[13950]_ ;
  assign \new_[13952]_  = \new_[13951]_  & \new_[13946]_ ;
  assign \new_[13955]_  = ~A168 & ~A169;
  assign \new_[13958]_  = A166 & A167;
  assign \new_[13959]_  = \new_[13958]_  & \new_[13955]_ ;
  assign \new_[13962]_  = A201 & A199;
  assign \new_[13966]_  = A301 & A234;
  assign \new_[13967]_  = A232 & \new_[13966]_ ;
  assign \new_[13968]_  = \new_[13967]_  & \new_[13962]_ ;
  assign \new_[13971]_  = ~A168 & ~A169;
  assign \new_[13974]_  = A166 & A167;
  assign \new_[13975]_  = \new_[13974]_  & \new_[13971]_ ;
  assign \new_[13978]_  = A201 & A199;
  assign \new_[13982]_  = A268 & A234;
  assign \new_[13983]_  = A232 & \new_[13982]_ ;
  assign \new_[13984]_  = \new_[13983]_  & \new_[13978]_ ;
  assign \new_[13987]_  = ~A168 & ~A169;
  assign \new_[13990]_  = A166 & A167;
  assign \new_[13991]_  = \new_[13990]_  & \new_[13987]_ ;
  assign \new_[13994]_  = A201 & A199;
  assign \new_[13998]_  = A301 & A234;
  assign \new_[13999]_  = A233 & \new_[13998]_ ;
  assign \new_[14000]_  = \new_[13999]_  & \new_[13994]_ ;
  assign \new_[14003]_  = ~A168 & ~A169;
  assign \new_[14006]_  = A166 & A167;
  assign \new_[14007]_  = \new_[14006]_  & \new_[14003]_ ;
  assign \new_[14010]_  = A201 & A199;
  assign \new_[14014]_  = A268 & A234;
  assign \new_[14015]_  = A233 & \new_[14014]_ ;
  assign \new_[14016]_  = \new_[14015]_  & \new_[14010]_ ;
  assign \new_[14019]_  = ~A168 & ~A169;
  assign \new_[14022]_  = A166 & A167;
  assign \new_[14023]_  = \new_[14022]_  & \new_[14019]_ ;
  assign \new_[14026]_  = A201 & A200;
  assign \new_[14030]_  = A300 & A299;
  assign \new_[14031]_  = A235 & \new_[14030]_ ;
  assign \new_[14032]_  = \new_[14031]_  & \new_[14026]_ ;
  assign \new_[14035]_  = ~A168 & ~A169;
  assign \new_[14038]_  = A166 & A167;
  assign \new_[14039]_  = \new_[14038]_  & \new_[14035]_ ;
  assign \new_[14042]_  = A201 & A200;
  assign \new_[14046]_  = A300 & A298;
  assign \new_[14047]_  = A235 & \new_[14046]_ ;
  assign \new_[14048]_  = \new_[14047]_  & \new_[14042]_ ;
  assign \new_[14051]_  = ~A168 & ~A169;
  assign \new_[14054]_  = A166 & A167;
  assign \new_[14055]_  = \new_[14054]_  & \new_[14051]_ ;
  assign \new_[14058]_  = A201 & A200;
  assign \new_[14062]_  = A267 & A265;
  assign \new_[14063]_  = A235 & \new_[14062]_ ;
  assign \new_[14064]_  = \new_[14063]_  & \new_[14058]_ ;
  assign \new_[14067]_  = ~A168 & ~A169;
  assign \new_[14070]_  = A166 & A167;
  assign \new_[14071]_  = \new_[14070]_  & \new_[14067]_ ;
  assign \new_[14074]_  = A201 & A200;
  assign \new_[14078]_  = A267 & A266;
  assign \new_[14079]_  = A235 & \new_[14078]_ ;
  assign \new_[14080]_  = \new_[14079]_  & \new_[14074]_ ;
  assign \new_[14083]_  = ~A168 & ~A169;
  assign \new_[14086]_  = A166 & A167;
  assign \new_[14087]_  = \new_[14086]_  & \new_[14083]_ ;
  assign \new_[14090]_  = A201 & A200;
  assign \new_[14094]_  = A301 & A234;
  assign \new_[14095]_  = A232 & \new_[14094]_ ;
  assign \new_[14096]_  = \new_[14095]_  & \new_[14090]_ ;
  assign \new_[14099]_  = ~A168 & ~A169;
  assign \new_[14102]_  = A166 & A167;
  assign \new_[14103]_  = \new_[14102]_  & \new_[14099]_ ;
  assign \new_[14106]_  = A201 & A200;
  assign \new_[14110]_  = A268 & A234;
  assign \new_[14111]_  = A232 & \new_[14110]_ ;
  assign \new_[14112]_  = \new_[14111]_  & \new_[14106]_ ;
  assign \new_[14115]_  = ~A168 & ~A169;
  assign \new_[14118]_  = A166 & A167;
  assign \new_[14119]_  = \new_[14118]_  & \new_[14115]_ ;
  assign \new_[14122]_  = A201 & A200;
  assign \new_[14126]_  = A301 & A234;
  assign \new_[14127]_  = A233 & \new_[14126]_ ;
  assign \new_[14128]_  = \new_[14127]_  & \new_[14122]_ ;
  assign \new_[14131]_  = ~A168 & ~A169;
  assign \new_[14134]_  = A166 & A167;
  assign \new_[14135]_  = \new_[14134]_  & \new_[14131]_ ;
  assign \new_[14138]_  = A201 & A200;
  assign \new_[14142]_  = A268 & A234;
  assign \new_[14143]_  = A233 & \new_[14142]_ ;
  assign \new_[14144]_  = \new_[14143]_  & \new_[14138]_ ;
  assign \new_[14147]_  = ~A168 & ~A169;
  assign \new_[14150]_  = A166 & A167;
  assign \new_[14151]_  = \new_[14150]_  & \new_[14147]_ ;
  assign \new_[14154]_  = A200 & ~A199;
  assign \new_[14158]_  = A301 & A235;
  assign \new_[14159]_  = A203 & \new_[14158]_ ;
  assign \new_[14160]_  = \new_[14159]_  & \new_[14154]_ ;
  assign \new_[14163]_  = ~A168 & ~A169;
  assign \new_[14166]_  = A166 & A167;
  assign \new_[14167]_  = \new_[14166]_  & \new_[14163]_ ;
  assign \new_[14170]_  = A200 & ~A199;
  assign \new_[14174]_  = A268 & A235;
  assign \new_[14175]_  = A203 & \new_[14174]_ ;
  assign \new_[14176]_  = \new_[14175]_  & \new_[14170]_ ;
  assign \new_[14179]_  = ~A168 & ~A169;
  assign \new_[14182]_  = A166 & A167;
  assign \new_[14183]_  = \new_[14182]_  & \new_[14179]_ ;
  assign \new_[14186]_  = ~A200 & A199;
  assign \new_[14190]_  = A301 & A235;
  assign \new_[14191]_  = A203 & \new_[14190]_ ;
  assign \new_[14192]_  = \new_[14191]_  & \new_[14186]_ ;
  assign \new_[14195]_  = ~A168 & ~A169;
  assign \new_[14198]_  = A166 & A167;
  assign \new_[14199]_  = \new_[14198]_  & \new_[14195]_ ;
  assign \new_[14202]_  = ~A200 & A199;
  assign \new_[14206]_  = A268 & A235;
  assign \new_[14207]_  = A203 & \new_[14206]_ ;
  assign \new_[14208]_  = \new_[14207]_  & \new_[14202]_ ;
  assign \new_[14211]_  = ~A169 & ~A170;
  assign \new_[14214]_  = A202 & ~A168;
  assign \new_[14215]_  = \new_[14214]_  & \new_[14211]_ ;
  assign \new_[14218]_  = A234 & A232;
  assign \new_[14222]_  = A302 & ~A299;
  assign \new_[14223]_  = A298 & \new_[14222]_ ;
  assign \new_[14224]_  = \new_[14223]_  & \new_[14218]_ ;
  assign \new_[14227]_  = ~A169 & ~A170;
  assign \new_[14230]_  = A202 & ~A168;
  assign \new_[14231]_  = \new_[14230]_  & \new_[14227]_ ;
  assign \new_[14234]_  = A234 & A232;
  assign \new_[14238]_  = A302 & A299;
  assign \new_[14239]_  = ~A298 & \new_[14238]_ ;
  assign \new_[14240]_  = \new_[14239]_  & \new_[14234]_ ;
  assign \new_[14243]_  = ~A169 & ~A170;
  assign \new_[14246]_  = A202 & ~A168;
  assign \new_[14247]_  = \new_[14246]_  & \new_[14243]_ ;
  assign \new_[14250]_  = A234 & A232;
  assign \new_[14254]_  = A269 & A266;
  assign \new_[14255]_  = ~A265 & \new_[14254]_ ;
  assign \new_[14256]_  = \new_[14255]_  & \new_[14250]_ ;
  assign \new_[14259]_  = ~A169 & ~A170;
  assign \new_[14262]_  = A202 & ~A168;
  assign \new_[14263]_  = \new_[14262]_  & \new_[14259]_ ;
  assign \new_[14266]_  = A234 & A232;
  assign \new_[14270]_  = A269 & ~A266;
  assign \new_[14271]_  = A265 & \new_[14270]_ ;
  assign \new_[14272]_  = \new_[14271]_  & \new_[14266]_ ;
  assign \new_[14275]_  = ~A169 & ~A170;
  assign \new_[14278]_  = A202 & ~A168;
  assign \new_[14279]_  = \new_[14278]_  & \new_[14275]_ ;
  assign \new_[14282]_  = A234 & A233;
  assign \new_[14286]_  = A302 & ~A299;
  assign \new_[14287]_  = A298 & \new_[14286]_ ;
  assign \new_[14288]_  = \new_[14287]_  & \new_[14282]_ ;
  assign \new_[14291]_  = ~A169 & ~A170;
  assign \new_[14294]_  = A202 & ~A168;
  assign \new_[14295]_  = \new_[14294]_  & \new_[14291]_ ;
  assign \new_[14298]_  = A234 & A233;
  assign \new_[14302]_  = A302 & A299;
  assign \new_[14303]_  = ~A298 & \new_[14302]_ ;
  assign \new_[14304]_  = \new_[14303]_  & \new_[14298]_ ;
  assign \new_[14307]_  = ~A169 & ~A170;
  assign \new_[14310]_  = A202 & ~A168;
  assign \new_[14311]_  = \new_[14310]_  & \new_[14307]_ ;
  assign \new_[14314]_  = A234 & A233;
  assign \new_[14318]_  = A269 & A266;
  assign \new_[14319]_  = ~A265 & \new_[14318]_ ;
  assign \new_[14320]_  = \new_[14319]_  & \new_[14314]_ ;
  assign \new_[14323]_  = ~A169 & ~A170;
  assign \new_[14326]_  = A202 & ~A168;
  assign \new_[14327]_  = \new_[14326]_  & \new_[14323]_ ;
  assign \new_[14330]_  = A234 & A233;
  assign \new_[14334]_  = A269 & ~A266;
  assign \new_[14335]_  = A265 & \new_[14334]_ ;
  assign \new_[14336]_  = \new_[14335]_  & \new_[14330]_ ;
  assign \new_[14339]_  = ~A169 & ~A170;
  assign \new_[14342]_  = A202 & ~A168;
  assign \new_[14343]_  = \new_[14342]_  & \new_[14339]_ ;
  assign \new_[14346]_  = A233 & ~A232;
  assign \new_[14350]_  = A300 & A299;
  assign \new_[14351]_  = A236 & \new_[14350]_ ;
  assign \new_[14352]_  = \new_[14351]_  & \new_[14346]_ ;
  assign \new_[14355]_  = ~A169 & ~A170;
  assign \new_[14358]_  = A202 & ~A168;
  assign \new_[14359]_  = \new_[14358]_  & \new_[14355]_ ;
  assign \new_[14362]_  = A233 & ~A232;
  assign \new_[14366]_  = A300 & A298;
  assign \new_[14367]_  = A236 & \new_[14366]_ ;
  assign \new_[14368]_  = \new_[14367]_  & \new_[14362]_ ;
  assign \new_[14371]_  = ~A169 & ~A170;
  assign \new_[14374]_  = A202 & ~A168;
  assign \new_[14375]_  = \new_[14374]_  & \new_[14371]_ ;
  assign \new_[14378]_  = A233 & ~A232;
  assign \new_[14382]_  = A267 & A265;
  assign \new_[14383]_  = A236 & \new_[14382]_ ;
  assign \new_[14384]_  = \new_[14383]_  & \new_[14378]_ ;
  assign \new_[14387]_  = ~A169 & ~A170;
  assign \new_[14390]_  = A202 & ~A168;
  assign \new_[14391]_  = \new_[14390]_  & \new_[14387]_ ;
  assign \new_[14394]_  = A233 & ~A232;
  assign \new_[14398]_  = A267 & A266;
  assign \new_[14399]_  = A236 & \new_[14398]_ ;
  assign \new_[14400]_  = \new_[14399]_  & \new_[14394]_ ;
  assign \new_[14403]_  = ~A169 & ~A170;
  assign \new_[14406]_  = A202 & ~A168;
  assign \new_[14407]_  = \new_[14406]_  & \new_[14403]_ ;
  assign \new_[14410]_  = ~A233 & A232;
  assign \new_[14414]_  = A300 & A299;
  assign \new_[14415]_  = A236 & \new_[14414]_ ;
  assign \new_[14416]_  = \new_[14415]_  & \new_[14410]_ ;
  assign \new_[14419]_  = ~A169 & ~A170;
  assign \new_[14422]_  = A202 & ~A168;
  assign \new_[14423]_  = \new_[14422]_  & \new_[14419]_ ;
  assign \new_[14426]_  = ~A233 & A232;
  assign \new_[14430]_  = A300 & A298;
  assign \new_[14431]_  = A236 & \new_[14430]_ ;
  assign \new_[14432]_  = \new_[14431]_  & \new_[14426]_ ;
  assign \new_[14435]_  = ~A169 & ~A170;
  assign \new_[14438]_  = A202 & ~A168;
  assign \new_[14439]_  = \new_[14438]_  & \new_[14435]_ ;
  assign \new_[14442]_  = ~A233 & A232;
  assign \new_[14446]_  = A267 & A265;
  assign \new_[14447]_  = A236 & \new_[14446]_ ;
  assign \new_[14448]_  = \new_[14447]_  & \new_[14442]_ ;
  assign \new_[14451]_  = ~A169 & ~A170;
  assign \new_[14454]_  = A202 & ~A168;
  assign \new_[14455]_  = \new_[14454]_  & \new_[14451]_ ;
  assign \new_[14458]_  = ~A233 & A232;
  assign \new_[14462]_  = A267 & A266;
  assign \new_[14463]_  = A236 & \new_[14462]_ ;
  assign \new_[14464]_  = \new_[14463]_  & \new_[14458]_ ;
  assign \new_[14467]_  = ~A169 & ~A170;
  assign \new_[14470]_  = A199 & ~A168;
  assign \new_[14471]_  = \new_[14470]_  & \new_[14467]_ ;
  assign \new_[14474]_  = A235 & A201;
  assign \new_[14478]_  = A302 & ~A299;
  assign \new_[14479]_  = A298 & \new_[14478]_ ;
  assign \new_[14480]_  = \new_[14479]_  & \new_[14474]_ ;
  assign \new_[14483]_  = ~A169 & ~A170;
  assign \new_[14486]_  = A199 & ~A168;
  assign \new_[14487]_  = \new_[14486]_  & \new_[14483]_ ;
  assign \new_[14490]_  = A235 & A201;
  assign \new_[14494]_  = A302 & A299;
  assign \new_[14495]_  = ~A298 & \new_[14494]_ ;
  assign \new_[14496]_  = \new_[14495]_  & \new_[14490]_ ;
  assign \new_[14499]_  = ~A169 & ~A170;
  assign \new_[14502]_  = A199 & ~A168;
  assign \new_[14503]_  = \new_[14502]_  & \new_[14499]_ ;
  assign \new_[14506]_  = A235 & A201;
  assign \new_[14510]_  = A269 & A266;
  assign \new_[14511]_  = ~A265 & \new_[14510]_ ;
  assign \new_[14512]_  = \new_[14511]_  & \new_[14506]_ ;
  assign \new_[14515]_  = ~A169 & ~A170;
  assign \new_[14518]_  = A199 & ~A168;
  assign \new_[14519]_  = \new_[14518]_  & \new_[14515]_ ;
  assign \new_[14522]_  = A235 & A201;
  assign \new_[14526]_  = A269 & ~A266;
  assign \new_[14527]_  = A265 & \new_[14526]_ ;
  assign \new_[14528]_  = \new_[14527]_  & \new_[14522]_ ;
  assign \new_[14531]_  = ~A169 & ~A170;
  assign \new_[14534]_  = A199 & ~A168;
  assign \new_[14535]_  = \new_[14534]_  & \new_[14531]_ ;
  assign \new_[14538]_  = A232 & A201;
  assign \new_[14542]_  = A300 & A299;
  assign \new_[14543]_  = A234 & \new_[14542]_ ;
  assign \new_[14544]_  = \new_[14543]_  & \new_[14538]_ ;
  assign \new_[14547]_  = ~A169 & ~A170;
  assign \new_[14550]_  = A199 & ~A168;
  assign \new_[14551]_  = \new_[14550]_  & \new_[14547]_ ;
  assign \new_[14554]_  = A232 & A201;
  assign \new_[14558]_  = A300 & A298;
  assign \new_[14559]_  = A234 & \new_[14558]_ ;
  assign \new_[14560]_  = \new_[14559]_  & \new_[14554]_ ;
  assign \new_[14563]_  = ~A169 & ~A170;
  assign \new_[14566]_  = A199 & ~A168;
  assign \new_[14567]_  = \new_[14566]_  & \new_[14563]_ ;
  assign \new_[14570]_  = A232 & A201;
  assign \new_[14574]_  = A267 & A265;
  assign \new_[14575]_  = A234 & \new_[14574]_ ;
  assign \new_[14576]_  = \new_[14575]_  & \new_[14570]_ ;
  assign \new_[14579]_  = ~A169 & ~A170;
  assign \new_[14582]_  = A199 & ~A168;
  assign \new_[14583]_  = \new_[14582]_  & \new_[14579]_ ;
  assign \new_[14586]_  = A232 & A201;
  assign \new_[14590]_  = A267 & A266;
  assign \new_[14591]_  = A234 & \new_[14590]_ ;
  assign \new_[14592]_  = \new_[14591]_  & \new_[14586]_ ;
  assign \new_[14595]_  = ~A169 & ~A170;
  assign \new_[14598]_  = A199 & ~A168;
  assign \new_[14599]_  = \new_[14598]_  & \new_[14595]_ ;
  assign \new_[14602]_  = A233 & A201;
  assign \new_[14606]_  = A300 & A299;
  assign \new_[14607]_  = A234 & \new_[14606]_ ;
  assign \new_[14608]_  = \new_[14607]_  & \new_[14602]_ ;
  assign \new_[14611]_  = ~A169 & ~A170;
  assign \new_[14614]_  = A199 & ~A168;
  assign \new_[14615]_  = \new_[14614]_  & \new_[14611]_ ;
  assign \new_[14618]_  = A233 & A201;
  assign \new_[14622]_  = A300 & A298;
  assign \new_[14623]_  = A234 & \new_[14622]_ ;
  assign \new_[14624]_  = \new_[14623]_  & \new_[14618]_ ;
  assign \new_[14627]_  = ~A169 & ~A170;
  assign \new_[14630]_  = A199 & ~A168;
  assign \new_[14631]_  = \new_[14630]_  & \new_[14627]_ ;
  assign \new_[14634]_  = A233 & A201;
  assign \new_[14638]_  = A267 & A265;
  assign \new_[14639]_  = A234 & \new_[14638]_ ;
  assign \new_[14640]_  = \new_[14639]_  & \new_[14634]_ ;
  assign \new_[14643]_  = ~A169 & ~A170;
  assign \new_[14646]_  = A199 & ~A168;
  assign \new_[14647]_  = \new_[14646]_  & \new_[14643]_ ;
  assign \new_[14650]_  = A233 & A201;
  assign \new_[14654]_  = A267 & A266;
  assign \new_[14655]_  = A234 & \new_[14654]_ ;
  assign \new_[14656]_  = \new_[14655]_  & \new_[14650]_ ;
  assign \new_[14659]_  = ~A169 & ~A170;
  assign \new_[14662]_  = A199 & ~A168;
  assign \new_[14663]_  = \new_[14662]_  & \new_[14659]_ ;
  assign \new_[14666]_  = ~A232 & A201;
  assign \new_[14670]_  = A301 & A236;
  assign \new_[14671]_  = A233 & \new_[14670]_ ;
  assign \new_[14672]_  = \new_[14671]_  & \new_[14666]_ ;
  assign \new_[14675]_  = ~A169 & ~A170;
  assign \new_[14678]_  = A199 & ~A168;
  assign \new_[14679]_  = \new_[14678]_  & \new_[14675]_ ;
  assign \new_[14682]_  = ~A232 & A201;
  assign \new_[14686]_  = A268 & A236;
  assign \new_[14687]_  = A233 & \new_[14686]_ ;
  assign \new_[14688]_  = \new_[14687]_  & \new_[14682]_ ;
  assign \new_[14691]_  = ~A169 & ~A170;
  assign \new_[14694]_  = A199 & ~A168;
  assign \new_[14695]_  = \new_[14694]_  & \new_[14691]_ ;
  assign \new_[14698]_  = A232 & A201;
  assign \new_[14702]_  = A301 & A236;
  assign \new_[14703]_  = ~A233 & \new_[14702]_ ;
  assign \new_[14704]_  = \new_[14703]_  & \new_[14698]_ ;
  assign \new_[14707]_  = ~A169 & ~A170;
  assign \new_[14710]_  = A199 & ~A168;
  assign \new_[14711]_  = \new_[14710]_  & \new_[14707]_ ;
  assign \new_[14714]_  = A232 & A201;
  assign \new_[14718]_  = A268 & A236;
  assign \new_[14719]_  = ~A233 & \new_[14718]_ ;
  assign \new_[14720]_  = \new_[14719]_  & \new_[14714]_ ;
  assign \new_[14723]_  = ~A169 & ~A170;
  assign \new_[14726]_  = A200 & ~A168;
  assign \new_[14727]_  = \new_[14726]_  & \new_[14723]_ ;
  assign \new_[14730]_  = A235 & A201;
  assign \new_[14734]_  = A302 & ~A299;
  assign \new_[14735]_  = A298 & \new_[14734]_ ;
  assign \new_[14736]_  = \new_[14735]_  & \new_[14730]_ ;
  assign \new_[14739]_  = ~A169 & ~A170;
  assign \new_[14742]_  = A200 & ~A168;
  assign \new_[14743]_  = \new_[14742]_  & \new_[14739]_ ;
  assign \new_[14746]_  = A235 & A201;
  assign \new_[14750]_  = A302 & A299;
  assign \new_[14751]_  = ~A298 & \new_[14750]_ ;
  assign \new_[14752]_  = \new_[14751]_  & \new_[14746]_ ;
  assign \new_[14755]_  = ~A169 & ~A170;
  assign \new_[14758]_  = A200 & ~A168;
  assign \new_[14759]_  = \new_[14758]_  & \new_[14755]_ ;
  assign \new_[14762]_  = A235 & A201;
  assign \new_[14766]_  = A269 & A266;
  assign \new_[14767]_  = ~A265 & \new_[14766]_ ;
  assign \new_[14768]_  = \new_[14767]_  & \new_[14762]_ ;
  assign \new_[14771]_  = ~A169 & ~A170;
  assign \new_[14774]_  = A200 & ~A168;
  assign \new_[14775]_  = \new_[14774]_  & \new_[14771]_ ;
  assign \new_[14778]_  = A235 & A201;
  assign \new_[14782]_  = A269 & ~A266;
  assign \new_[14783]_  = A265 & \new_[14782]_ ;
  assign \new_[14784]_  = \new_[14783]_  & \new_[14778]_ ;
  assign \new_[14787]_  = ~A169 & ~A170;
  assign \new_[14790]_  = A200 & ~A168;
  assign \new_[14791]_  = \new_[14790]_  & \new_[14787]_ ;
  assign \new_[14794]_  = A232 & A201;
  assign \new_[14798]_  = A300 & A299;
  assign \new_[14799]_  = A234 & \new_[14798]_ ;
  assign \new_[14800]_  = \new_[14799]_  & \new_[14794]_ ;
  assign \new_[14803]_  = ~A169 & ~A170;
  assign \new_[14806]_  = A200 & ~A168;
  assign \new_[14807]_  = \new_[14806]_  & \new_[14803]_ ;
  assign \new_[14810]_  = A232 & A201;
  assign \new_[14814]_  = A300 & A298;
  assign \new_[14815]_  = A234 & \new_[14814]_ ;
  assign \new_[14816]_  = \new_[14815]_  & \new_[14810]_ ;
  assign \new_[14819]_  = ~A169 & ~A170;
  assign \new_[14822]_  = A200 & ~A168;
  assign \new_[14823]_  = \new_[14822]_  & \new_[14819]_ ;
  assign \new_[14826]_  = A232 & A201;
  assign \new_[14830]_  = A267 & A265;
  assign \new_[14831]_  = A234 & \new_[14830]_ ;
  assign \new_[14832]_  = \new_[14831]_  & \new_[14826]_ ;
  assign \new_[14835]_  = ~A169 & ~A170;
  assign \new_[14838]_  = A200 & ~A168;
  assign \new_[14839]_  = \new_[14838]_  & \new_[14835]_ ;
  assign \new_[14842]_  = A232 & A201;
  assign \new_[14846]_  = A267 & A266;
  assign \new_[14847]_  = A234 & \new_[14846]_ ;
  assign \new_[14848]_  = \new_[14847]_  & \new_[14842]_ ;
  assign \new_[14851]_  = ~A169 & ~A170;
  assign \new_[14854]_  = A200 & ~A168;
  assign \new_[14855]_  = \new_[14854]_  & \new_[14851]_ ;
  assign \new_[14858]_  = A233 & A201;
  assign \new_[14862]_  = A300 & A299;
  assign \new_[14863]_  = A234 & \new_[14862]_ ;
  assign \new_[14864]_  = \new_[14863]_  & \new_[14858]_ ;
  assign \new_[14867]_  = ~A169 & ~A170;
  assign \new_[14870]_  = A200 & ~A168;
  assign \new_[14871]_  = \new_[14870]_  & \new_[14867]_ ;
  assign \new_[14874]_  = A233 & A201;
  assign \new_[14878]_  = A300 & A298;
  assign \new_[14879]_  = A234 & \new_[14878]_ ;
  assign \new_[14880]_  = \new_[14879]_  & \new_[14874]_ ;
  assign \new_[14883]_  = ~A169 & ~A170;
  assign \new_[14886]_  = A200 & ~A168;
  assign \new_[14887]_  = \new_[14886]_  & \new_[14883]_ ;
  assign \new_[14890]_  = A233 & A201;
  assign \new_[14894]_  = A267 & A265;
  assign \new_[14895]_  = A234 & \new_[14894]_ ;
  assign \new_[14896]_  = \new_[14895]_  & \new_[14890]_ ;
  assign \new_[14899]_  = ~A169 & ~A170;
  assign \new_[14902]_  = A200 & ~A168;
  assign \new_[14903]_  = \new_[14902]_  & \new_[14899]_ ;
  assign \new_[14906]_  = A233 & A201;
  assign \new_[14910]_  = A267 & A266;
  assign \new_[14911]_  = A234 & \new_[14910]_ ;
  assign \new_[14912]_  = \new_[14911]_  & \new_[14906]_ ;
  assign \new_[14915]_  = ~A169 & ~A170;
  assign \new_[14918]_  = A200 & ~A168;
  assign \new_[14919]_  = \new_[14918]_  & \new_[14915]_ ;
  assign \new_[14922]_  = ~A232 & A201;
  assign \new_[14926]_  = A301 & A236;
  assign \new_[14927]_  = A233 & \new_[14926]_ ;
  assign \new_[14928]_  = \new_[14927]_  & \new_[14922]_ ;
  assign \new_[14931]_  = ~A169 & ~A170;
  assign \new_[14934]_  = A200 & ~A168;
  assign \new_[14935]_  = \new_[14934]_  & \new_[14931]_ ;
  assign \new_[14938]_  = ~A232 & A201;
  assign \new_[14942]_  = A268 & A236;
  assign \new_[14943]_  = A233 & \new_[14942]_ ;
  assign \new_[14944]_  = \new_[14943]_  & \new_[14938]_ ;
  assign \new_[14947]_  = ~A169 & ~A170;
  assign \new_[14950]_  = A200 & ~A168;
  assign \new_[14951]_  = \new_[14950]_  & \new_[14947]_ ;
  assign \new_[14954]_  = A232 & A201;
  assign \new_[14958]_  = A301 & A236;
  assign \new_[14959]_  = ~A233 & \new_[14958]_ ;
  assign \new_[14960]_  = \new_[14959]_  & \new_[14954]_ ;
  assign \new_[14963]_  = ~A169 & ~A170;
  assign \new_[14966]_  = A200 & ~A168;
  assign \new_[14967]_  = \new_[14966]_  & \new_[14963]_ ;
  assign \new_[14970]_  = A232 & A201;
  assign \new_[14974]_  = A268 & A236;
  assign \new_[14975]_  = ~A233 & \new_[14974]_ ;
  assign \new_[14976]_  = \new_[14975]_  & \new_[14970]_ ;
  assign \new_[14979]_  = ~A169 & ~A170;
  assign \new_[14982]_  = ~A199 & ~A168;
  assign \new_[14983]_  = \new_[14982]_  & \new_[14979]_ ;
  assign \new_[14986]_  = A203 & A200;
  assign \new_[14990]_  = A300 & A299;
  assign \new_[14991]_  = A235 & \new_[14990]_ ;
  assign \new_[14992]_  = \new_[14991]_  & \new_[14986]_ ;
  assign \new_[14995]_  = ~A169 & ~A170;
  assign \new_[14998]_  = ~A199 & ~A168;
  assign \new_[14999]_  = \new_[14998]_  & \new_[14995]_ ;
  assign \new_[15002]_  = A203 & A200;
  assign \new_[15006]_  = A300 & A298;
  assign \new_[15007]_  = A235 & \new_[15006]_ ;
  assign \new_[15008]_  = \new_[15007]_  & \new_[15002]_ ;
  assign \new_[15011]_  = ~A169 & ~A170;
  assign \new_[15014]_  = ~A199 & ~A168;
  assign \new_[15015]_  = \new_[15014]_  & \new_[15011]_ ;
  assign \new_[15018]_  = A203 & A200;
  assign \new_[15022]_  = A267 & A265;
  assign \new_[15023]_  = A235 & \new_[15022]_ ;
  assign \new_[15024]_  = \new_[15023]_  & \new_[15018]_ ;
  assign \new_[15027]_  = ~A169 & ~A170;
  assign \new_[15030]_  = ~A199 & ~A168;
  assign \new_[15031]_  = \new_[15030]_  & \new_[15027]_ ;
  assign \new_[15034]_  = A203 & A200;
  assign \new_[15038]_  = A267 & A266;
  assign \new_[15039]_  = A235 & \new_[15038]_ ;
  assign \new_[15040]_  = \new_[15039]_  & \new_[15034]_ ;
  assign \new_[15043]_  = ~A169 & ~A170;
  assign \new_[15046]_  = ~A199 & ~A168;
  assign \new_[15047]_  = \new_[15046]_  & \new_[15043]_ ;
  assign \new_[15050]_  = A203 & A200;
  assign \new_[15054]_  = A301 & A234;
  assign \new_[15055]_  = A232 & \new_[15054]_ ;
  assign \new_[15056]_  = \new_[15055]_  & \new_[15050]_ ;
  assign \new_[15059]_  = ~A169 & ~A170;
  assign \new_[15062]_  = ~A199 & ~A168;
  assign \new_[15063]_  = \new_[15062]_  & \new_[15059]_ ;
  assign \new_[15066]_  = A203 & A200;
  assign \new_[15070]_  = A268 & A234;
  assign \new_[15071]_  = A232 & \new_[15070]_ ;
  assign \new_[15072]_  = \new_[15071]_  & \new_[15066]_ ;
  assign \new_[15075]_  = ~A169 & ~A170;
  assign \new_[15078]_  = ~A199 & ~A168;
  assign \new_[15079]_  = \new_[15078]_  & \new_[15075]_ ;
  assign \new_[15082]_  = A203 & A200;
  assign \new_[15086]_  = A301 & A234;
  assign \new_[15087]_  = A233 & \new_[15086]_ ;
  assign \new_[15088]_  = \new_[15087]_  & \new_[15082]_ ;
  assign \new_[15091]_  = ~A169 & ~A170;
  assign \new_[15094]_  = ~A199 & ~A168;
  assign \new_[15095]_  = \new_[15094]_  & \new_[15091]_ ;
  assign \new_[15098]_  = A203 & A200;
  assign \new_[15102]_  = A268 & A234;
  assign \new_[15103]_  = A233 & \new_[15102]_ ;
  assign \new_[15104]_  = \new_[15103]_  & \new_[15098]_ ;
  assign \new_[15107]_  = ~A169 & ~A170;
  assign \new_[15110]_  = A199 & ~A168;
  assign \new_[15111]_  = \new_[15110]_  & \new_[15107]_ ;
  assign \new_[15114]_  = A203 & ~A200;
  assign \new_[15118]_  = A300 & A299;
  assign \new_[15119]_  = A235 & \new_[15118]_ ;
  assign \new_[15120]_  = \new_[15119]_  & \new_[15114]_ ;
  assign \new_[15123]_  = ~A169 & ~A170;
  assign \new_[15126]_  = A199 & ~A168;
  assign \new_[15127]_  = \new_[15126]_  & \new_[15123]_ ;
  assign \new_[15130]_  = A203 & ~A200;
  assign \new_[15134]_  = A300 & A298;
  assign \new_[15135]_  = A235 & \new_[15134]_ ;
  assign \new_[15136]_  = \new_[15135]_  & \new_[15130]_ ;
  assign \new_[15139]_  = ~A169 & ~A170;
  assign \new_[15142]_  = A199 & ~A168;
  assign \new_[15143]_  = \new_[15142]_  & \new_[15139]_ ;
  assign \new_[15146]_  = A203 & ~A200;
  assign \new_[15150]_  = A267 & A265;
  assign \new_[15151]_  = A235 & \new_[15150]_ ;
  assign \new_[15152]_  = \new_[15151]_  & \new_[15146]_ ;
  assign \new_[15155]_  = ~A169 & ~A170;
  assign \new_[15158]_  = A199 & ~A168;
  assign \new_[15159]_  = \new_[15158]_  & \new_[15155]_ ;
  assign \new_[15162]_  = A203 & ~A200;
  assign \new_[15166]_  = A267 & A266;
  assign \new_[15167]_  = A235 & \new_[15166]_ ;
  assign \new_[15168]_  = \new_[15167]_  & \new_[15162]_ ;
  assign \new_[15171]_  = ~A169 & ~A170;
  assign \new_[15174]_  = A199 & ~A168;
  assign \new_[15175]_  = \new_[15174]_  & \new_[15171]_ ;
  assign \new_[15178]_  = A203 & ~A200;
  assign \new_[15182]_  = A301 & A234;
  assign \new_[15183]_  = A232 & \new_[15182]_ ;
  assign \new_[15184]_  = \new_[15183]_  & \new_[15178]_ ;
  assign \new_[15187]_  = ~A169 & ~A170;
  assign \new_[15190]_  = A199 & ~A168;
  assign \new_[15191]_  = \new_[15190]_  & \new_[15187]_ ;
  assign \new_[15194]_  = A203 & ~A200;
  assign \new_[15198]_  = A268 & A234;
  assign \new_[15199]_  = A232 & \new_[15198]_ ;
  assign \new_[15200]_  = \new_[15199]_  & \new_[15194]_ ;
  assign \new_[15203]_  = ~A169 & ~A170;
  assign \new_[15206]_  = A199 & ~A168;
  assign \new_[15207]_  = \new_[15206]_  & \new_[15203]_ ;
  assign \new_[15210]_  = A203 & ~A200;
  assign \new_[15214]_  = A301 & A234;
  assign \new_[15215]_  = A233 & \new_[15214]_ ;
  assign \new_[15216]_  = \new_[15215]_  & \new_[15210]_ ;
  assign \new_[15219]_  = ~A169 & ~A170;
  assign \new_[15222]_  = A199 & ~A168;
  assign \new_[15223]_  = \new_[15222]_  & \new_[15219]_ ;
  assign \new_[15226]_  = A203 & ~A200;
  assign \new_[15230]_  = A268 & A234;
  assign \new_[15231]_  = A233 & \new_[15230]_ ;
  assign \new_[15232]_  = \new_[15231]_  & \new_[15226]_ ;
  assign \new_[15235]_  = A166 & A168;
  assign \new_[15239]_  = ~A203 & ~A202;
  assign \new_[15240]_  = ~A201 & \new_[15239]_ ;
  assign \new_[15241]_  = \new_[15240]_  & \new_[15235]_ ;
  assign \new_[15244]_  = A234 & A232;
  assign \new_[15248]_  = A302 & ~A299;
  assign \new_[15249]_  = A298 & \new_[15248]_ ;
  assign \new_[15250]_  = \new_[15249]_  & \new_[15244]_ ;
  assign \new_[15253]_  = A166 & A168;
  assign \new_[15257]_  = ~A203 & ~A202;
  assign \new_[15258]_  = ~A201 & \new_[15257]_ ;
  assign \new_[15259]_  = \new_[15258]_  & \new_[15253]_ ;
  assign \new_[15262]_  = A234 & A232;
  assign \new_[15266]_  = A302 & A299;
  assign \new_[15267]_  = ~A298 & \new_[15266]_ ;
  assign \new_[15268]_  = \new_[15267]_  & \new_[15262]_ ;
  assign \new_[15271]_  = A166 & A168;
  assign \new_[15275]_  = ~A203 & ~A202;
  assign \new_[15276]_  = ~A201 & \new_[15275]_ ;
  assign \new_[15277]_  = \new_[15276]_  & \new_[15271]_ ;
  assign \new_[15280]_  = A234 & A232;
  assign \new_[15284]_  = A269 & A266;
  assign \new_[15285]_  = ~A265 & \new_[15284]_ ;
  assign \new_[15286]_  = \new_[15285]_  & \new_[15280]_ ;
  assign \new_[15289]_  = A166 & A168;
  assign \new_[15293]_  = ~A203 & ~A202;
  assign \new_[15294]_  = ~A201 & \new_[15293]_ ;
  assign \new_[15295]_  = \new_[15294]_  & \new_[15289]_ ;
  assign \new_[15298]_  = A234 & A232;
  assign \new_[15302]_  = A269 & ~A266;
  assign \new_[15303]_  = A265 & \new_[15302]_ ;
  assign \new_[15304]_  = \new_[15303]_  & \new_[15298]_ ;
  assign \new_[15307]_  = A166 & A168;
  assign \new_[15311]_  = ~A203 & ~A202;
  assign \new_[15312]_  = ~A201 & \new_[15311]_ ;
  assign \new_[15313]_  = \new_[15312]_  & \new_[15307]_ ;
  assign \new_[15316]_  = A234 & A233;
  assign \new_[15320]_  = A302 & ~A299;
  assign \new_[15321]_  = A298 & \new_[15320]_ ;
  assign \new_[15322]_  = \new_[15321]_  & \new_[15316]_ ;
  assign \new_[15325]_  = A166 & A168;
  assign \new_[15329]_  = ~A203 & ~A202;
  assign \new_[15330]_  = ~A201 & \new_[15329]_ ;
  assign \new_[15331]_  = \new_[15330]_  & \new_[15325]_ ;
  assign \new_[15334]_  = A234 & A233;
  assign \new_[15338]_  = A302 & A299;
  assign \new_[15339]_  = ~A298 & \new_[15338]_ ;
  assign \new_[15340]_  = \new_[15339]_  & \new_[15334]_ ;
  assign \new_[15343]_  = A166 & A168;
  assign \new_[15347]_  = ~A203 & ~A202;
  assign \new_[15348]_  = ~A201 & \new_[15347]_ ;
  assign \new_[15349]_  = \new_[15348]_  & \new_[15343]_ ;
  assign \new_[15352]_  = A234 & A233;
  assign \new_[15356]_  = A269 & A266;
  assign \new_[15357]_  = ~A265 & \new_[15356]_ ;
  assign \new_[15358]_  = \new_[15357]_  & \new_[15352]_ ;
  assign \new_[15361]_  = A166 & A168;
  assign \new_[15365]_  = ~A203 & ~A202;
  assign \new_[15366]_  = ~A201 & \new_[15365]_ ;
  assign \new_[15367]_  = \new_[15366]_  & \new_[15361]_ ;
  assign \new_[15370]_  = A234 & A233;
  assign \new_[15374]_  = A269 & ~A266;
  assign \new_[15375]_  = A265 & \new_[15374]_ ;
  assign \new_[15376]_  = \new_[15375]_  & \new_[15370]_ ;
  assign \new_[15379]_  = A166 & A168;
  assign \new_[15383]_  = ~A203 & ~A202;
  assign \new_[15384]_  = ~A201 & \new_[15383]_ ;
  assign \new_[15385]_  = \new_[15384]_  & \new_[15379]_ ;
  assign \new_[15388]_  = A233 & ~A232;
  assign \new_[15392]_  = A300 & A299;
  assign \new_[15393]_  = A236 & \new_[15392]_ ;
  assign \new_[15394]_  = \new_[15393]_  & \new_[15388]_ ;
  assign \new_[15397]_  = A166 & A168;
  assign \new_[15401]_  = ~A203 & ~A202;
  assign \new_[15402]_  = ~A201 & \new_[15401]_ ;
  assign \new_[15403]_  = \new_[15402]_  & \new_[15397]_ ;
  assign \new_[15406]_  = A233 & ~A232;
  assign \new_[15410]_  = A300 & A298;
  assign \new_[15411]_  = A236 & \new_[15410]_ ;
  assign \new_[15412]_  = \new_[15411]_  & \new_[15406]_ ;
  assign \new_[15415]_  = A166 & A168;
  assign \new_[15419]_  = ~A203 & ~A202;
  assign \new_[15420]_  = ~A201 & \new_[15419]_ ;
  assign \new_[15421]_  = \new_[15420]_  & \new_[15415]_ ;
  assign \new_[15424]_  = A233 & ~A232;
  assign \new_[15428]_  = A267 & A265;
  assign \new_[15429]_  = A236 & \new_[15428]_ ;
  assign \new_[15430]_  = \new_[15429]_  & \new_[15424]_ ;
  assign \new_[15433]_  = A166 & A168;
  assign \new_[15437]_  = ~A203 & ~A202;
  assign \new_[15438]_  = ~A201 & \new_[15437]_ ;
  assign \new_[15439]_  = \new_[15438]_  & \new_[15433]_ ;
  assign \new_[15442]_  = A233 & ~A232;
  assign \new_[15446]_  = A267 & A266;
  assign \new_[15447]_  = A236 & \new_[15446]_ ;
  assign \new_[15448]_  = \new_[15447]_  & \new_[15442]_ ;
  assign \new_[15451]_  = A166 & A168;
  assign \new_[15455]_  = ~A203 & ~A202;
  assign \new_[15456]_  = ~A201 & \new_[15455]_ ;
  assign \new_[15457]_  = \new_[15456]_  & \new_[15451]_ ;
  assign \new_[15460]_  = ~A233 & A232;
  assign \new_[15464]_  = A300 & A299;
  assign \new_[15465]_  = A236 & \new_[15464]_ ;
  assign \new_[15466]_  = \new_[15465]_  & \new_[15460]_ ;
  assign \new_[15469]_  = A166 & A168;
  assign \new_[15473]_  = ~A203 & ~A202;
  assign \new_[15474]_  = ~A201 & \new_[15473]_ ;
  assign \new_[15475]_  = \new_[15474]_  & \new_[15469]_ ;
  assign \new_[15478]_  = ~A233 & A232;
  assign \new_[15482]_  = A300 & A298;
  assign \new_[15483]_  = A236 & \new_[15482]_ ;
  assign \new_[15484]_  = \new_[15483]_  & \new_[15478]_ ;
  assign \new_[15487]_  = A166 & A168;
  assign \new_[15491]_  = ~A203 & ~A202;
  assign \new_[15492]_  = ~A201 & \new_[15491]_ ;
  assign \new_[15493]_  = \new_[15492]_  & \new_[15487]_ ;
  assign \new_[15496]_  = ~A233 & A232;
  assign \new_[15500]_  = A267 & A265;
  assign \new_[15501]_  = A236 & \new_[15500]_ ;
  assign \new_[15502]_  = \new_[15501]_  & \new_[15496]_ ;
  assign \new_[15505]_  = A166 & A168;
  assign \new_[15509]_  = ~A203 & ~A202;
  assign \new_[15510]_  = ~A201 & \new_[15509]_ ;
  assign \new_[15511]_  = \new_[15510]_  & \new_[15505]_ ;
  assign \new_[15514]_  = ~A233 & A232;
  assign \new_[15518]_  = A267 & A266;
  assign \new_[15519]_  = A236 & \new_[15518]_ ;
  assign \new_[15520]_  = \new_[15519]_  & \new_[15514]_ ;
  assign \new_[15523]_  = A166 & A168;
  assign \new_[15527]_  = ~A201 & A200;
  assign \new_[15528]_  = A199 & \new_[15527]_ ;
  assign \new_[15529]_  = \new_[15528]_  & \new_[15523]_ ;
  assign \new_[15532]_  = A235 & ~A202;
  assign \new_[15536]_  = A302 & ~A299;
  assign \new_[15537]_  = A298 & \new_[15536]_ ;
  assign \new_[15538]_  = \new_[15537]_  & \new_[15532]_ ;
  assign \new_[15541]_  = A166 & A168;
  assign \new_[15545]_  = ~A201 & A200;
  assign \new_[15546]_  = A199 & \new_[15545]_ ;
  assign \new_[15547]_  = \new_[15546]_  & \new_[15541]_ ;
  assign \new_[15550]_  = A235 & ~A202;
  assign \new_[15554]_  = A302 & A299;
  assign \new_[15555]_  = ~A298 & \new_[15554]_ ;
  assign \new_[15556]_  = \new_[15555]_  & \new_[15550]_ ;
  assign \new_[15559]_  = A166 & A168;
  assign \new_[15563]_  = ~A201 & A200;
  assign \new_[15564]_  = A199 & \new_[15563]_ ;
  assign \new_[15565]_  = \new_[15564]_  & \new_[15559]_ ;
  assign \new_[15568]_  = A235 & ~A202;
  assign \new_[15572]_  = A269 & A266;
  assign \new_[15573]_  = ~A265 & \new_[15572]_ ;
  assign \new_[15574]_  = \new_[15573]_  & \new_[15568]_ ;
  assign \new_[15577]_  = A166 & A168;
  assign \new_[15581]_  = ~A201 & A200;
  assign \new_[15582]_  = A199 & \new_[15581]_ ;
  assign \new_[15583]_  = \new_[15582]_  & \new_[15577]_ ;
  assign \new_[15586]_  = A235 & ~A202;
  assign \new_[15590]_  = A269 & ~A266;
  assign \new_[15591]_  = A265 & \new_[15590]_ ;
  assign \new_[15592]_  = \new_[15591]_  & \new_[15586]_ ;
  assign \new_[15595]_  = A166 & A168;
  assign \new_[15599]_  = ~A201 & A200;
  assign \new_[15600]_  = A199 & \new_[15599]_ ;
  assign \new_[15601]_  = \new_[15600]_  & \new_[15595]_ ;
  assign \new_[15604]_  = A232 & ~A202;
  assign \new_[15608]_  = A300 & A299;
  assign \new_[15609]_  = A234 & \new_[15608]_ ;
  assign \new_[15610]_  = \new_[15609]_  & \new_[15604]_ ;
  assign \new_[15613]_  = A166 & A168;
  assign \new_[15617]_  = ~A201 & A200;
  assign \new_[15618]_  = A199 & \new_[15617]_ ;
  assign \new_[15619]_  = \new_[15618]_  & \new_[15613]_ ;
  assign \new_[15622]_  = A232 & ~A202;
  assign \new_[15626]_  = A300 & A298;
  assign \new_[15627]_  = A234 & \new_[15626]_ ;
  assign \new_[15628]_  = \new_[15627]_  & \new_[15622]_ ;
  assign \new_[15631]_  = A166 & A168;
  assign \new_[15635]_  = ~A201 & A200;
  assign \new_[15636]_  = A199 & \new_[15635]_ ;
  assign \new_[15637]_  = \new_[15636]_  & \new_[15631]_ ;
  assign \new_[15640]_  = A232 & ~A202;
  assign \new_[15644]_  = A267 & A265;
  assign \new_[15645]_  = A234 & \new_[15644]_ ;
  assign \new_[15646]_  = \new_[15645]_  & \new_[15640]_ ;
  assign \new_[15649]_  = A166 & A168;
  assign \new_[15653]_  = ~A201 & A200;
  assign \new_[15654]_  = A199 & \new_[15653]_ ;
  assign \new_[15655]_  = \new_[15654]_  & \new_[15649]_ ;
  assign \new_[15658]_  = A232 & ~A202;
  assign \new_[15662]_  = A267 & A266;
  assign \new_[15663]_  = A234 & \new_[15662]_ ;
  assign \new_[15664]_  = \new_[15663]_  & \new_[15658]_ ;
  assign \new_[15667]_  = A166 & A168;
  assign \new_[15671]_  = ~A201 & A200;
  assign \new_[15672]_  = A199 & \new_[15671]_ ;
  assign \new_[15673]_  = \new_[15672]_  & \new_[15667]_ ;
  assign \new_[15676]_  = A233 & ~A202;
  assign \new_[15680]_  = A300 & A299;
  assign \new_[15681]_  = A234 & \new_[15680]_ ;
  assign \new_[15682]_  = \new_[15681]_  & \new_[15676]_ ;
  assign \new_[15685]_  = A166 & A168;
  assign \new_[15689]_  = ~A201 & A200;
  assign \new_[15690]_  = A199 & \new_[15689]_ ;
  assign \new_[15691]_  = \new_[15690]_  & \new_[15685]_ ;
  assign \new_[15694]_  = A233 & ~A202;
  assign \new_[15698]_  = A300 & A298;
  assign \new_[15699]_  = A234 & \new_[15698]_ ;
  assign \new_[15700]_  = \new_[15699]_  & \new_[15694]_ ;
  assign \new_[15703]_  = A166 & A168;
  assign \new_[15707]_  = ~A201 & A200;
  assign \new_[15708]_  = A199 & \new_[15707]_ ;
  assign \new_[15709]_  = \new_[15708]_  & \new_[15703]_ ;
  assign \new_[15712]_  = A233 & ~A202;
  assign \new_[15716]_  = A267 & A265;
  assign \new_[15717]_  = A234 & \new_[15716]_ ;
  assign \new_[15718]_  = \new_[15717]_  & \new_[15712]_ ;
  assign \new_[15721]_  = A166 & A168;
  assign \new_[15725]_  = ~A201 & A200;
  assign \new_[15726]_  = A199 & \new_[15725]_ ;
  assign \new_[15727]_  = \new_[15726]_  & \new_[15721]_ ;
  assign \new_[15730]_  = A233 & ~A202;
  assign \new_[15734]_  = A267 & A266;
  assign \new_[15735]_  = A234 & \new_[15734]_ ;
  assign \new_[15736]_  = \new_[15735]_  & \new_[15730]_ ;
  assign \new_[15739]_  = A166 & A168;
  assign \new_[15743]_  = ~A201 & A200;
  assign \new_[15744]_  = A199 & \new_[15743]_ ;
  assign \new_[15745]_  = \new_[15744]_  & \new_[15739]_ ;
  assign \new_[15748]_  = ~A232 & ~A202;
  assign \new_[15752]_  = A301 & A236;
  assign \new_[15753]_  = A233 & \new_[15752]_ ;
  assign \new_[15754]_  = \new_[15753]_  & \new_[15748]_ ;
  assign \new_[15757]_  = A166 & A168;
  assign \new_[15761]_  = ~A201 & A200;
  assign \new_[15762]_  = A199 & \new_[15761]_ ;
  assign \new_[15763]_  = \new_[15762]_  & \new_[15757]_ ;
  assign \new_[15766]_  = ~A232 & ~A202;
  assign \new_[15770]_  = A268 & A236;
  assign \new_[15771]_  = A233 & \new_[15770]_ ;
  assign \new_[15772]_  = \new_[15771]_  & \new_[15766]_ ;
  assign \new_[15775]_  = A166 & A168;
  assign \new_[15779]_  = ~A201 & A200;
  assign \new_[15780]_  = A199 & \new_[15779]_ ;
  assign \new_[15781]_  = \new_[15780]_  & \new_[15775]_ ;
  assign \new_[15784]_  = A232 & ~A202;
  assign \new_[15788]_  = A301 & A236;
  assign \new_[15789]_  = ~A233 & \new_[15788]_ ;
  assign \new_[15790]_  = \new_[15789]_  & \new_[15784]_ ;
  assign \new_[15793]_  = A166 & A168;
  assign \new_[15797]_  = ~A201 & A200;
  assign \new_[15798]_  = A199 & \new_[15797]_ ;
  assign \new_[15799]_  = \new_[15798]_  & \new_[15793]_ ;
  assign \new_[15802]_  = A232 & ~A202;
  assign \new_[15806]_  = A268 & A236;
  assign \new_[15807]_  = ~A233 & \new_[15806]_ ;
  assign \new_[15808]_  = \new_[15807]_  & \new_[15802]_ ;
  assign \new_[15811]_  = A166 & A168;
  assign \new_[15815]_  = ~A202 & ~A200;
  assign \new_[15816]_  = ~A199 & \new_[15815]_ ;
  assign \new_[15817]_  = \new_[15816]_  & \new_[15811]_ ;
  assign \new_[15820]_  = A234 & A232;
  assign \new_[15824]_  = A302 & ~A299;
  assign \new_[15825]_  = A298 & \new_[15824]_ ;
  assign \new_[15826]_  = \new_[15825]_  & \new_[15820]_ ;
  assign \new_[15829]_  = A166 & A168;
  assign \new_[15833]_  = ~A202 & ~A200;
  assign \new_[15834]_  = ~A199 & \new_[15833]_ ;
  assign \new_[15835]_  = \new_[15834]_  & \new_[15829]_ ;
  assign \new_[15838]_  = A234 & A232;
  assign \new_[15842]_  = A302 & A299;
  assign \new_[15843]_  = ~A298 & \new_[15842]_ ;
  assign \new_[15844]_  = \new_[15843]_  & \new_[15838]_ ;
  assign \new_[15847]_  = A166 & A168;
  assign \new_[15851]_  = ~A202 & ~A200;
  assign \new_[15852]_  = ~A199 & \new_[15851]_ ;
  assign \new_[15853]_  = \new_[15852]_  & \new_[15847]_ ;
  assign \new_[15856]_  = A234 & A232;
  assign \new_[15860]_  = A269 & A266;
  assign \new_[15861]_  = ~A265 & \new_[15860]_ ;
  assign \new_[15862]_  = \new_[15861]_  & \new_[15856]_ ;
  assign \new_[15865]_  = A166 & A168;
  assign \new_[15869]_  = ~A202 & ~A200;
  assign \new_[15870]_  = ~A199 & \new_[15869]_ ;
  assign \new_[15871]_  = \new_[15870]_  & \new_[15865]_ ;
  assign \new_[15874]_  = A234 & A232;
  assign \new_[15878]_  = A269 & ~A266;
  assign \new_[15879]_  = A265 & \new_[15878]_ ;
  assign \new_[15880]_  = \new_[15879]_  & \new_[15874]_ ;
  assign \new_[15883]_  = A166 & A168;
  assign \new_[15887]_  = ~A202 & ~A200;
  assign \new_[15888]_  = ~A199 & \new_[15887]_ ;
  assign \new_[15889]_  = \new_[15888]_  & \new_[15883]_ ;
  assign \new_[15892]_  = A234 & A233;
  assign \new_[15896]_  = A302 & ~A299;
  assign \new_[15897]_  = A298 & \new_[15896]_ ;
  assign \new_[15898]_  = \new_[15897]_  & \new_[15892]_ ;
  assign \new_[15901]_  = A166 & A168;
  assign \new_[15905]_  = ~A202 & ~A200;
  assign \new_[15906]_  = ~A199 & \new_[15905]_ ;
  assign \new_[15907]_  = \new_[15906]_  & \new_[15901]_ ;
  assign \new_[15910]_  = A234 & A233;
  assign \new_[15914]_  = A302 & A299;
  assign \new_[15915]_  = ~A298 & \new_[15914]_ ;
  assign \new_[15916]_  = \new_[15915]_  & \new_[15910]_ ;
  assign \new_[15919]_  = A166 & A168;
  assign \new_[15923]_  = ~A202 & ~A200;
  assign \new_[15924]_  = ~A199 & \new_[15923]_ ;
  assign \new_[15925]_  = \new_[15924]_  & \new_[15919]_ ;
  assign \new_[15928]_  = A234 & A233;
  assign \new_[15932]_  = A269 & A266;
  assign \new_[15933]_  = ~A265 & \new_[15932]_ ;
  assign \new_[15934]_  = \new_[15933]_  & \new_[15928]_ ;
  assign \new_[15937]_  = A166 & A168;
  assign \new_[15941]_  = ~A202 & ~A200;
  assign \new_[15942]_  = ~A199 & \new_[15941]_ ;
  assign \new_[15943]_  = \new_[15942]_  & \new_[15937]_ ;
  assign \new_[15946]_  = A234 & A233;
  assign \new_[15950]_  = A269 & ~A266;
  assign \new_[15951]_  = A265 & \new_[15950]_ ;
  assign \new_[15952]_  = \new_[15951]_  & \new_[15946]_ ;
  assign \new_[15955]_  = A166 & A168;
  assign \new_[15959]_  = ~A202 & ~A200;
  assign \new_[15960]_  = ~A199 & \new_[15959]_ ;
  assign \new_[15961]_  = \new_[15960]_  & \new_[15955]_ ;
  assign \new_[15964]_  = A233 & ~A232;
  assign \new_[15968]_  = A300 & A299;
  assign \new_[15969]_  = A236 & \new_[15968]_ ;
  assign \new_[15970]_  = \new_[15969]_  & \new_[15964]_ ;
  assign \new_[15973]_  = A166 & A168;
  assign \new_[15977]_  = ~A202 & ~A200;
  assign \new_[15978]_  = ~A199 & \new_[15977]_ ;
  assign \new_[15979]_  = \new_[15978]_  & \new_[15973]_ ;
  assign \new_[15982]_  = A233 & ~A232;
  assign \new_[15986]_  = A300 & A298;
  assign \new_[15987]_  = A236 & \new_[15986]_ ;
  assign \new_[15988]_  = \new_[15987]_  & \new_[15982]_ ;
  assign \new_[15991]_  = A166 & A168;
  assign \new_[15995]_  = ~A202 & ~A200;
  assign \new_[15996]_  = ~A199 & \new_[15995]_ ;
  assign \new_[15997]_  = \new_[15996]_  & \new_[15991]_ ;
  assign \new_[16000]_  = A233 & ~A232;
  assign \new_[16004]_  = A267 & A265;
  assign \new_[16005]_  = A236 & \new_[16004]_ ;
  assign \new_[16006]_  = \new_[16005]_  & \new_[16000]_ ;
  assign \new_[16009]_  = A166 & A168;
  assign \new_[16013]_  = ~A202 & ~A200;
  assign \new_[16014]_  = ~A199 & \new_[16013]_ ;
  assign \new_[16015]_  = \new_[16014]_  & \new_[16009]_ ;
  assign \new_[16018]_  = A233 & ~A232;
  assign \new_[16022]_  = A267 & A266;
  assign \new_[16023]_  = A236 & \new_[16022]_ ;
  assign \new_[16024]_  = \new_[16023]_  & \new_[16018]_ ;
  assign \new_[16027]_  = A166 & A168;
  assign \new_[16031]_  = ~A202 & ~A200;
  assign \new_[16032]_  = ~A199 & \new_[16031]_ ;
  assign \new_[16033]_  = \new_[16032]_  & \new_[16027]_ ;
  assign \new_[16036]_  = ~A233 & A232;
  assign \new_[16040]_  = A300 & A299;
  assign \new_[16041]_  = A236 & \new_[16040]_ ;
  assign \new_[16042]_  = \new_[16041]_  & \new_[16036]_ ;
  assign \new_[16045]_  = A166 & A168;
  assign \new_[16049]_  = ~A202 & ~A200;
  assign \new_[16050]_  = ~A199 & \new_[16049]_ ;
  assign \new_[16051]_  = \new_[16050]_  & \new_[16045]_ ;
  assign \new_[16054]_  = ~A233 & A232;
  assign \new_[16058]_  = A300 & A298;
  assign \new_[16059]_  = A236 & \new_[16058]_ ;
  assign \new_[16060]_  = \new_[16059]_  & \new_[16054]_ ;
  assign \new_[16063]_  = A166 & A168;
  assign \new_[16067]_  = ~A202 & ~A200;
  assign \new_[16068]_  = ~A199 & \new_[16067]_ ;
  assign \new_[16069]_  = \new_[16068]_  & \new_[16063]_ ;
  assign \new_[16072]_  = ~A233 & A232;
  assign \new_[16076]_  = A267 & A265;
  assign \new_[16077]_  = A236 & \new_[16076]_ ;
  assign \new_[16078]_  = \new_[16077]_  & \new_[16072]_ ;
  assign \new_[16081]_  = A166 & A168;
  assign \new_[16085]_  = ~A202 & ~A200;
  assign \new_[16086]_  = ~A199 & \new_[16085]_ ;
  assign \new_[16087]_  = \new_[16086]_  & \new_[16081]_ ;
  assign \new_[16090]_  = ~A233 & A232;
  assign \new_[16094]_  = A267 & A266;
  assign \new_[16095]_  = A236 & \new_[16094]_ ;
  assign \new_[16096]_  = \new_[16095]_  & \new_[16090]_ ;
  assign \new_[16099]_  = A167 & A168;
  assign \new_[16103]_  = ~A203 & ~A202;
  assign \new_[16104]_  = ~A201 & \new_[16103]_ ;
  assign \new_[16105]_  = \new_[16104]_  & \new_[16099]_ ;
  assign \new_[16108]_  = A234 & A232;
  assign \new_[16112]_  = A302 & ~A299;
  assign \new_[16113]_  = A298 & \new_[16112]_ ;
  assign \new_[16114]_  = \new_[16113]_  & \new_[16108]_ ;
  assign \new_[16117]_  = A167 & A168;
  assign \new_[16121]_  = ~A203 & ~A202;
  assign \new_[16122]_  = ~A201 & \new_[16121]_ ;
  assign \new_[16123]_  = \new_[16122]_  & \new_[16117]_ ;
  assign \new_[16126]_  = A234 & A232;
  assign \new_[16130]_  = A302 & A299;
  assign \new_[16131]_  = ~A298 & \new_[16130]_ ;
  assign \new_[16132]_  = \new_[16131]_  & \new_[16126]_ ;
  assign \new_[16135]_  = A167 & A168;
  assign \new_[16139]_  = ~A203 & ~A202;
  assign \new_[16140]_  = ~A201 & \new_[16139]_ ;
  assign \new_[16141]_  = \new_[16140]_  & \new_[16135]_ ;
  assign \new_[16144]_  = A234 & A232;
  assign \new_[16148]_  = A269 & A266;
  assign \new_[16149]_  = ~A265 & \new_[16148]_ ;
  assign \new_[16150]_  = \new_[16149]_  & \new_[16144]_ ;
  assign \new_[16153]_  = A167 & A168;
  assign \new_[16157]_  = ~A203 & ~A202;
  assign \new_[16158]_  = ~A201 & \new_[16157]_ ;
  assign \new_[16159]_  = \new_[16158]_  & \new_[16153]_ ;
  assign \new_[16162]_  = A234 & A232;
  assign \new_[16166]_  = A269 & ~A266;
  assign \new_[16167]_  = A265 & \new_[16166]_ ;
  assign \new_[16168]_  = \new_[16167]_  & \new_[16162]_ ;
  assign \new_[16171]_  = A167 & A168;
  assign \new_[16175]_  = ~A203 & ~A202;
  assign \new_[16176]_  = ~A201 & \new_[16175]_ ;
  assign \new_[16177]_  = \new_[16176]_  & \new_[16171]_ ;
  assign \new_[16180]_  = A234 & A233;
  assign \new_[16184]_  = A302 & ~A299;
  assign \new_[16185]_  = A298 & \new_[16184]_ ;
  assign \new_[16186]_  = \new_[16185]_  & \new_[16180]_ ;
  assign \new_[16189]_  = A167 & A168;
  assign \new_[16193]_  = ~A203 & ~A202;
  assign \new_[16194]_  = ~A201 & \new_[16193]_ ;
  assign \new_[16195]_  = \new_[16194]_  & \new_[16189]_ ;
  assign \new_[16198]_  = A234 & A233;
  assign \new_[16202]_  = A302 & A299;
  assign \new_[16203]_  = ~A298 & \new_[16202]_ ;
  assign \new_[16204]_  = \new_[16203]_  & \new_[16198]_ ;
  assign \new_[16207]_  = A167 & A168;
  assign \new_[16211]_  = ~A203 & ~A202;
  assign \new_[16212]_  = ~A201 & \new_[16211]_ ;
  assign \new_[16213]_  = \new_[16212]_  & \new_[16207]_ ;
  assign \new_[16216]_  = A234 & A233;
  assign \new_[16220]_  = A269 & A266;
  assign \new_[16221]_  = ~A265 & \new_[16220]_ ;
  assign \new_[16222]_  = \new_[16221]_  & \new_[16216]_ ;
  assign \new_[16225]_  = A167 & A168;
  assign \new_[16229]_  = ~A203 & ~A202;
  assign \new_[16230]_  = ~A201 & \new_[16229]_ ;
  assign \new_[16231]_  = \new_[16230]_  & \new_[16225]_ ;
  assign \new_[16234]_  = A234 & A233;
  assign \new_[16238]_  = A269 & ~A266;
  assign \new_[16239]_  = A265 & \new_[16238]_ ;
  assign \new_[16240]_  = \new_[16239]_  & \new_[16234]_ ;
  assign \new_[16243]_  = A167 & A168;
  assign \new_[16247]_  = ~A203 & ~A202;
  assign \new_[16248]_  = ~A201 & \new_[16247]_ ;
  assign \new_[16249]_  = \new_[16248]_  & \new_[16243]_ ;
  assign \new_[16252]_  = A233 & ~A232;
  assign \new_[16256]_  = A300 & A299;
  assign \new_[16257]_  = A236 & \new_[16256]_ ;
  assign \new_[16258]_  = \new_[16257]_  & \new_[16252]_ ;
  assign \new_[16261]_  = A167 & A168;
  assign \new_[16265]_  = ~A203 & ~A202;
  assign \new_[16266]_  = ~A201 & \new_[16265]_ ;
  assign \new_[16267]_  = \new_[16266]_  & \new_[16261]_ ;
  assign \new_[16270]_  = A233 & ~A232;
  assign \new_[16274]_  = A300 & A298;
  assign \new_[16275]_  = A236 & \new_[16274]_ ;
  assign \new_[16276]_  = \new_[16275]_  & \new_[16270]_ ;
  assign \new_[16279]_  = A167 & A168;
  assign \new_[16283]_  = ~A203 & ~A202;
  assign \new_[16284]_  = ~A201 & \new_[16283]_ ;
  assign \new_[16285]_  = \new_[16284]_  & \new_[16279]_ ;
  assign \new_[16288]_  = A233 & ~A232;
  assign \new_[16292]_  = A267 & A265;
  assign \new_[16293]_  = A236 & \new_[16292]_ ;
  assign \new_[16294]_  = \new_[16293]_  & \new_[16288]_ ;
  assign \new_[16297]_  = A167 & A168;
  assign \new_[16301]_  = ~A203 & ~A202;
  assign \new_[16302]_  = ~A201 & \new_[16301]_ ;
  assign \new_[16303]_  = \new_[16302]_  & \new_[16297]_ ;
  assign \new_[16306]_  = A233 & ~A232;
  assign \new_[16310]_  = A267 & A266;
  assign \new_[16311]_  = A236 & \new_[16310]_ ;
  assign \new_[16312]_  = \new_[16311]_  & \new_[16306]_ ;
  assign \new_[16315]_  = A167 & A168;
  assign \new_[16319]_  = ~A203 & ~A202;
  assign \new_[16320]_  = ~A201 & \new_[16319]_ ;
  assign \new_[16321]_  = \new_[16320]_  & \new_[16315]_ ;
  assign \new_[16324]_  = ~A233 & A232;
  assign \new_[16328]_  = A300 & A299;
  assign \new_[16329]_  = A236 & \new_[16328]_ ;
  assign \new_[16330]_  = \new_[16329]_  & \new_[16324]_ ;
  assign \new_[16333]_  = A167 & A168;
  assign \new_[16337]_  = ~A203 & ~A202;
  assign \new_[16338]_  = ~A201 & \new_[16337]_ ;
  assign \new_[16339]_  = \new_[16338]_  & \new_[16333]_ ;
  assign \new_[16342]_  = ~A233 & A232;
  assign \new_[16346]_  = A300 & A298;
  assign \new_[16347]_  = A236 & \new_[16346]_ ;
  assign \new_[16348]_  = \new_[16347]_  & \new_[16342]_ ;
  assign \new_[16351]_  = A167 & A168;
  assign \new_[16355]_  = ~A203 & ~A202;
  assign \new_[16356]_  = ~A201 & \new_[16355]_ ;
  assign \new_[16357]_  = \new_[16356]_  & \new_[16351]_ ;
  assign \new_[16360]_  = ~A233 & A232;
  assign \new_[16364]_  = A267 & A265;
  assign \new_[16365]_  = A236 & \new_[16364]_ ;
  assign \new_[16366]_  = \new_[16365]_  & \new_[16360]_ ;
  assign \new_[16369]_  = A167 & A168;
  assign \new_[16373]_  = ~A203 & ~A202;
  assign \new_[16374]_  = ~A201 & \new_[16373]_ ;
  assign \new_[16375]_  = \new_[16374]_  & \new_[16369]_ ;
  assign \new_[16378]_  = ~A233 & A232;
  assign \new_[16382]_  = A267 & A266;
  assign \new_[16383]_  = A236 & \new_[16382]_ ;
  assign \new_[16384]_  = \new_[16383]_  & \new_[16378]_ ;
  assign \new_[16387]_  = A167 & A168;
  assign \new_[16391]_  = ~A201 & A200;
  assign \new_[16392]_  = A199 & \new_[16391]_ ;
  assign \new_[16393]_  = \new_[16392]_  & \new_[16387]_ ;
  assign \new_[16396]_  = A235 & ~A202;
  assign \new_[16400]_  = A302 & ~A299;
  assign \new_[16401]_  = A298 & \new_[16400]_ ;
  assign \new_[16402]_  = \new_[16401]_  & \new_[16396]_ ;
  assign \new_[16405]_  = A167 & A168;
  assign \new_[16409]_  = ~A201 & A200;
  assign \new_[16410]_  = A199 & \new_[16409]_ ;
  assign \new_[16411]_  = \new_[16410]_  & \new_[16405]_ ;
  assign \new_[16414]_  = A235 & ~A202;
  assign \new_[16418]_  = A302 & A299;
  assign \new_[16419]_  = ~A298 & \new_[16418]_ ;
  assign \new_[16420]_  = \new_[16419]_  & \new_[16414]_ ;
  assign \new_[16423]_  = A167 & A168;
  assign \new_[16427]_  = ~A201 & A200;
  assign \new_[16428]_  = A199 & \new_[16427]_ ;
  assign \new_[16429]_  = \new_[16428]_  & \new_[16423]_ ;
  assign \new_[16432]_  = A235 & ~A202;
  assign \new_[16436]_  = A269 & A266;
  assign \new_[16437]_  = ~A265 & \new_[16436]_ ;
  assign \new_[16438]_  = \new_[16437]_  & \new_[16432]_ ;
  assign \new_[16441]_  = A167 & A168;
  assign \new_[16445]_  = ~A201 & A200;
  assign \new_[16446]_  = A199 & \new_[16445]_ ;
  assign \new_[16447]_  = \new_[16446]_  & \new_[16441]_ ;
  assign \new_[16450]_  = A235 & ~A202;
  assign \new_[16454]_  = A269 & ~A266;
  assign \new_[16455]_  = A265 & \new_[16454]_ ;
  assign \new_[16456]_  = \new_[16455]_  & \new_[16450]_ ;
  assign \new_[16459]_  = A167 & A168;
  assign \new_[16463]_  = ~A201 & A200;
  assign \new_[16464]_  = A199 & \new_[16463]_ ;
  assign \new_[16465]_  = \new_[16464]_  & \new_[16459]_ ;
  assign \new_[16468]_  = A232 & ~A202;
  assign \new_[16472]_  = A300 & A299;
  assign \new_[16473]_  = A234 & \new_[16472]_ ;
  assign \new_[16474]_  = \new_[16473]_  & \new_[16468]_ ;
  assign \new_[16477]_  = A167 & A168;
  assign \new_[16481]_  = ~A201 & A200;
  assign \new_[16482]_  = A199 & \new_[16481]_ ;
  assign \new_[16483]_  = \new_[16482]_  & \new_[16477]_ ;
  assign \new_[16486]_  = A232 & ~A202;
  assign \new_[16490]_  = A300 & A298;
  assign \new_[16491]_  = A234 & \new_[16490]_ ;
  assign \new_[16492]_  = \new_[16491]_  & \new_[16486]_ ;
  assign \new_[16495]_  = A167 & A168;
  assign \new_[16499]_  = ~A201 & A200;
  assign \new_[16500]_  = A199 & \new_[16499]_ ;
  assign \new_[16501]_  = \new_[16500]_  & \new_[16495]_ ;
  assign \new_[16504]_  = A232 & ~A202;
  assign \new_[16508]_  = A267 & A265;
  assign \new_[16509]_  = A234 & \new_[16508]_ ;
  assign \new_[16510]_  = \new_[16509]_  & \new_[16504]_ ;
  assign \new_[16513]_  = A167 & A168;
  assign \new_[16517]_  = ~A201 & A200;
  assign \new_[16518]_  = A199 & \new_[16517]_ ;
  assign \new_[16519]_  = \new_[16518]_  & \new_[16513]_ ;
  assign \new_[16522]_  = A232 & ~A202;
  assign \new_[16526]_  = A267 & A266;
  assign \new_[16527]_  = A234 & \new_[16526]_ ;
  assign \new_[16528]_  = \new_[16527]_  & \new_[16522]_ ;
  assign \new_[16531]_  = A167 & A168;
  assign \new_[16535]_  = ~A201 & A200;
  assign \new_[16536]_  = A199 & \new_[16535]_ ;
  assign \new_[16537]_  = \new_[16536]_  & \new_[16531]_ ;
  assign \new_[16540]_  = A233 & ~A202;
  assign \new_[16544]_  = A300 & A299;
  assign \new_[16545]_  = A234 & \new_[16544]_ ;
  assign \new_[16546]_  = \new_[16545]_  & \new_[16540]_ ;
  assign \new_[16549]_  = A167 & A168;
  assign \new_[16553]_  = ~A201 & A200;
  assign \new_[16554]_  = A199 & \new_[16553]_ ;
  assign \new_[16555]_  = \new_[16554]_  & \new_[16549]_ ;
  assign \new_[16558]_  = A233 & ~A202;
  assign \new_[16562]_  = A300 & A298;
  assign \new_[16563]_  = A234 & \new_[16562]_ ;
  assign \new_[16564]_  = \new_[16563]_  & \new_[16558]_ ;
  assign \new_[16567]_  = A167 & A168;
  assign \new_[16571]_  = ~A201 & A200;
  assign \new_[16572]_  = A199 & \new_[16571]_ ;
  assign \new_[16573]_  = \new_[16572]_  & \new_[16567]_ ;
  assign \new_[16576]_  = A233 & ~A202;
  assign \new_[16580]_  = A267 & A265;
  assign \new_[16581]_  = A234 & \new_[16580]_ ;
  assign \new_[16582]_  = \new_[16581]_  & \new_[16576]_ ;
  assign \new_[16585]_  = A167 & A168;
  assign \new_[16589]_  = ~A201 & A200;
  assign \new_[16590]_  = A199 & \new_[16589]_ ;
  assign \new_[16591]_  = \new_[16590]_  & \new_[16585]_ ;
  assign \new_[16594]_  = A233 & ~A202;
  assign \new_[16598]_  = A267 & A266;
  assign \new_[16599]_  = A234 & \new_[16598]_ ;
  assign \new_[16600]_  = \new_[16599]_  & \new_[16594]_ ;
  assign \new_[16603]_  = A167 & A168;
  assign \new_[16607]_  = ~A201 & A200;
  assign \new_[16608]_  = A199 & \new_[16607]_ ;
  assign \new_[16609]_  = \new_[16608]_  & \new_[16603]_ ;
  assign \new_[16612]_  = ~A232 & ~A202;
  assign \new_[16616]_  = A301 & A236;
  assign \new_[16617]_  = A233 & \new_[16616]_ ;
  assign \new_[16618]_  = \new_[16617]_  & \new_[16612]_ ;
  assign \new_[16621]_  = A167 & A168;
  assign \new_[16625]_  = ~A201 & A200;
  assign \new_[16626]_  = A199 & \new_[16625]_ ;
  assign \new_[16627]_  = \new_[16626]_  & \new_[16621]_ ;
  assign \new_[16630]_  = ~A232 & ~A202;
  assign \new_[16634]_  = A268 & A236;
  assign \new_[16635]_  = A233 & \new_[16634]_ ;
  assign \new_[16636]_  = \new_[16635]_  & \new_[16630]_ ;
  assign \new_[16639]_  = A167 & A168;
  assign \new_[16643]_  = ~A201 & A200;
  assign \new_[16644]_  = A199 & \new_[16643]_ ;
  assign \new_[16645]_  = \new_[16644]_  & \new_[16639]_ ;
  assign \new_[16648]_  = A232 & ~A202;
  assign \new_[16652]_  = A301 & A236;
  assign \new_[16653]_  = ~A233 & \new_[16652]_ ;
  assign \new_[16654]_  = \new_[16653]_  & \new_[16648]_ ;
  assign \new_[16657]_  = A167 & A168;
  assign \new_[16661]_  = ~A201 & A200;
  assign \new_[16662]_  = A199 & \new_[16661]_ ;
  assign \new_[16663]_  = \new_[16662]_  & \new_[16657]_ ;
  assign \new_[16666]_  = A232 & ~A202;
  assign \new_[16670]_  = A268 & A236;
  assign \new_[16671]_  = ~A233 & \new_[16670]_ ;
  assign \new_[16672]_  = \new_[16671]_  & \new_[16666]_ ;
  assign \new_[16675]_  = A167 & A168;
  assign \new_[16679]_  = ~A202 & ~A200;
  assign \new_[16680]_  = ~A199 & \new_[16679]_ ;
  assign \new_[16681]_  = \new_[16680]_  & \new_[16675]_ ;
  assign \new_[16684]_  = A234 & A232;
  assign \new_[16688]_  = A302 & ~A299;
  assign \new_[16689]_  = A298 & \new_[16688]_ ;
  assign \new_[16690]_  = \new_[16689]_  & \new_[16684]_ ;
  assign \new_[16693]_  = A167 & A168;
  assign \new_[16697]_  = ~A202 & ~A200;
  assign \new_[16698]_  = ~A199 & \new_[16697]_ ;
  assign \new_[16699]_  = \new_[16698]_  & \new_[16693]_ ;
  assign \new_[16702]_  = A234 & A232;
  assign \new_[16706]_  = A302 & A299;
  assign \new_[16707]_  = ~A298 & \new_[16706]_ ;
  assign \new_[16708]_  = \new_[16707]_  & \new_[16702]_ ;
  assign \new_[16711]_  = A167 & A168;
  assign \new_[16715]_  = ~A202 & ~A200;
  assign \new_[16716]_  = ~A199 & \new_[16715]_ ;
  assign \new_[16717]_  = \new_[16716]_  & \new_[16711]_ ;
  assign \new_[16720]_  = A234 & A232;
  assign \new_[16724]_  = A269 & A266;
  assign \new_[16725]_  = ~A265 & \new_[16724]_ ;
  assign \new_[16726]_  = \new_[16725]_  & \new_[16720]_ ;
  assign \new_[16729]_  = A167 & A168;
  assign \new_[16733]_  = ~A202 & ~A200;
  assign \new_[16734]_  = ~A199 & \new_[16733]_ ;
  assign \new_[16735]_  = \new_[16734]_  & \new_[16729]_ ;
  assign \new_[16738]_  = A234 & A232;
  assign \new_[16742]_  = A269 & ~A266;
  assign \new_[16743]_  = A265 & \new_[16742]_ ;
  assign \new_[16744]_  = \new_[16743]_  & \new_[16738]_ ;
  assign \new_[16747]_  = A167 & A168;
  assign \new_[16751]_  = ~A202 & ~A200;
  assign \new_[16752]_  = ~A199 & \new_[16751]_ ;
  assign \new_[16753]_  = \new_[16752]_  & \new_[16747]_ ;
  assign \new_[16756]_  = A234 & A233;
  assign \new_[16760]_  = A302 & ~A299;
  assign \new_[16761]_  = A298 & \new_[16760]_ ;
  assign \new_[16762]_  = \new_[16761]_  & \new_[16756]_ ;
  assign \new_[16765]_  = A167 & A168;
  assign \new_[16769]_  = ~A202 & ~A200;
  assign \new_[16770]_  = ~A199 & \new_[16769]_ ;
  assign \new_[16771]_  = \new_[16770]_  & \new_[16765]_ ;
  assign \new_[16774]_  = A234 & A233;
  assign \new_[16778]_  = A302 & A299;
  assign \new_[16779]_  = ~A298 & \new_[16778]_ ;
  assign \new_[16780]_  = \new_[16779]_  & \new_[16774]_ ;
  assign \new_[16783]_  = A167 & A168;
  assign \new_[16787]_  = ~A202 & ~A200;
  assign \new_[16788]_  = ~A199 & \new_[16787]_ ;
  assign \new_[16789]_  = \new_[16788]_  & \new_[16783]_ ;
  assign \new_[16792]_  = A234 & A233;
  assign \new_[16796]_  = A269 & A266;
  assign \new_[16797]_  = ~A265 & \new_[16796]_ ;
  assign \new_[16798]_  = \new_[16797]_  & \new_[16792]_ ;
  assign \new_[16801]_  = A167 & A168;
  assign \new_[16805]_  = ~A202 & ~A200;
  assign \new_[16806]_  = ~A199 & \new_[16805]_ ;
  assign \new_[16807]_  = \new_[16806]_  & \new_[16801]_ ;
  assign \new_[16810]_  = A234 & A233;
  assign \new_[16814]_  = A269 & ~A266;
  assign \new_[16815]_  = A265 & \new_[16814]_ ;
  assign \new_[16816]_  = \new_[16815]_  & \new_[16810]_ ;
  assign \new_[16819]_  = A167 & A168;
  assign \new_[16823]_  = ~A202 & ~A200;
  assign \new_[16824]_  = ~A199 & \new_[16823]_ ;
  assign \new_[16825]_  = \new_[16824]_  & \new_[16819]_ ;
  assign \new_[16828]_  = A233 & ~A232;
  assign \new_[16832]_  = A300 & A299;
  assign \new_[16833]_  = A236 & \new_[16832]_ ;
  assign \new_[16834]_  = \new_[16833]_  & \new_[16828]_ ;
  assign \new_[16837]_  = A167 & A168;
  assign \new_[16841]_  = ~A202 & ~A200;
  assign \new_[16842]_  = ~A199 & \new_[16841]_ ;
  assign \new_[16843]_  = \new_[16842]_  & \new_[16837]_ ;
  assign \new_[16846]_  = A233 & ~A232;
  assign \new_[16850]_  = A300 & A298;
  assign \new_[16851]_  = A236 & \new_[16850]_ ;
  assign \new_[16852]_  = \new_[16851]_  & \new_[16846]_ ;
  assign \new_[16855]_  = A167 & A168;
  assign \new_[16859]_  = ~A202 & ~A200;
  assign \new_[16860]_  = ~A199 & \new_[16859]_ ;
  assign \new_[16861]_  = \new_[16860]_  & \new_[16855]_ ;
  assign \new_[16864]_  = A233 & ~A232;
  assign \new_[16868]_  = A267 & A265;
  assign \new_[16869]_  = A236 & \new_[16868]_ ;
  assign \new_[16870]_  = \new_[16869]_  & \new_[16864]_ ;
  assign \new_[16873]_  = A167 & A168;
  assign \new_[16877]_  = ~A202 & ~A200;
  assign \new_[16878]_  = ~A199 & \new_[16877]_ ;
  assign \new_[16879]_  = \new_[16878]_  & \new_[16873]_ ;
  assign \new_[16882]_  = A233 & ~A232;
  assign \new_[16886]_  = A267 & A266;
  assign \new_[16887]_  = A236 & \new_[16886]_ ;
  assign \new_[16888]_  = \new_[16887]_  & \new_[16882]_ ;
  assign \new_[16891]_  = A167 & A168;
  assign \new_[16895]_  = ~A202 & ~A200;
  assign \new_[16896]_  = ~A199 & \new_[16895]_ ;
  assign \new_[16897]_  = \new_[16896]_  & \new_[16891]_ ;
  assign \new_[16900]_  = ~A233 & A232;
  assign \new_[16904]_  = A300 & A299;
  assign \new_[16905]_  = A236 & \new_[16904]_ ;
  assign \new_[16906]_  = \new_[16905]_  & \new_[16900]_ ;
  assign \new_[16909]_  = A167 & A168;
  assign \new_[16913]_  = ~A202 & ~A200;
  assign \new_[16914]_  = ~A199 & \new_[16913]_ ;
  assign \new_[16915]_  = \new_[16914]_  & \new_[16909]_ ;
  assign \new_[16918]_  = ~A233 & A232;
  assign \new_[16922]_  = A300 & A298;
  assign \new_[16923]_  = A236 & \new_[16922]_ ;
  assign \new_[16924]_  = \new_[16923]_  & \new_[16918]_ ;
  assign \new_[16927]_  = A167 & A168;
  assign \new_[16931]_  = ~A202 & ~A200;
  assign \new_[16932]_  = ~A199 & \new_[16931]_ ;
  assign \new_[16933]_  = \new_[16932]_  & \new_[16927]_ ;
  assign \new_[16936]_  = ~A233 & A232;
  assign \new_[16940]_  = A267 & A265;
  assign \new_[16941]_  = A236 & \new_[16940]_ ;
  assign \new_[16942]_  = \new_[16941]_  & \new_[16936]_ ;
  assign \new_[16945]_  = A167 & A168;
  assign \new_[16949]_  = ~A202 & ~A200;
  assign \new_[16950]_  = ~A199 & \new_[16949]_ ;
  assign \new_[16951]_  = \new_[16950]_  & \new_[16945]_ ;
  assign \new_[16954]_  = ~A233 & A232;
  assign \new_[16958]_  = A267 & A266;
  assign \new_[16959]_  = A236 & \new_[16958]_ ;
  assign \new_[16960]_  = \new_[16959]_  & \new_[16954]_ ;
  assign \new_[16963]_  = A167 & A170;
  assign \new_[16967]_  = ~A202 & ~A201;
  assign \new_[16968]_  = ~A166 & \new_[16967]_ ;
  assign \new_[16969]_  = \new_[16968]_  & \new_[16963]_ ;
  assign \new_[16972]_  = A235 & ~A203;
  assign \new_[16976]_  = A302 & ~A299;
  assign \new_[16977]_  = A298 & \new_[16976]_ ;
  assign \new_[16978]_  = \new_[16977]_  & \new_[16972]_ ;
  assign \new_[16981]_  = A167 & A170;
  assign \new_[16985]_  = ~A202 & ~A201;
  assign \new_[16986]_  = ~A166 & \new_[16985]_ ;
  assign \new_[16987]_  = \new_[16986]_  & \new_[16981]_ ;
  assign \new_[16990]_  = A235 & ~A203;
  assign \new_[16994]_  = A302 & A299;
  assign \new_[16995]_  = ~A298 & \new_[16994]_ ;
  assign \new_[16996]_  = \new_[16995]_  & \new_[16990]_ ;
  assign \new_[16999]_  = A167 & A170;
  assign \new_[17003]_  = ~A202 & ~A201;
  assign \new_[17004]_  = ~A166 & \new_[17003]_ ;
  assign \new_[17005]_  = \new_[17004]_  & \new_[16999]_ ;
  assign \new_[17008]_  = A235 & ~A203;
  assign \new_[17012]_  = A269 & A266;
  assign \new_[17013]_  = ~A265 & \new_[17012]_ ;
  assign \new_[17014]_  = \new_[17013]_  & \new_[17008]_ ;
  assign \new_[17017]_  = A167 & A170;
  assign \new_[17021]_  = ~A202 & ~A201;
  assign \new_[17022]_  = ~A166 & \new_[17021]_ ;
  assign \new_[17023]_  = \new_[17022]_  & \new_[17017]_ ;
  assign \new_[17026]_  = A235 & ~A203;
  assign \new_[17030]_  = A269 & ~A266;
  assign \new_[17031]_  = A265 & \new_[17030]_ ;
  assign \new_[17032]_  = \new_[17031]_  & \new_[17026]_ ;
  assign \new_[17035]_  = A167 & A170;
  assign \new_[17039]_  = ~A202 & ~A201;
  assign \new_[17040]_  = ~A166 & \new_[17039]_ ;
  assign \new_[17041]_  = \new_[17040]_  & \new_[17035]_ ;
  assign \new_[17044]_  = A232 & ~A203;
  assign \new_[17048]_  = A300 & A299;
  assign \new_[17049]_  = A234 & \new_[17048]_ ;
  assign \new_[17050]_  = \new_[17049]_  & \new_[17044]_ ;
  assign \new_[17053]_  = A167 & A170;
  assign \new_[17057]_  = ~A202 & ~A201;
  assign \new_[17058]_  = ~A166 & \new_[17057]_ ;
  assign \new_[17059]_  = \new_[17058]_  & \new_[17053]_ ;
  assign \new_[17062]_  = A232 & ~A203;
  assign \new_[17066]_  = A300 & A298;
  assign \new_[17067]_  = A234 & \new_[17066]_ ;
  assign \new_[17068]_  = \new_[17067]_  & \new_[17062]_ ;
  assign \new_[17071]_  = A167 & A170;
  assign \new_[17075]_  = ~A202 & ~A201;
  assign \new_[17076]_  = ~A166 & \new_[17075]_ ;
  assign \new_[17077]_  = \new_[17076]_  & \new_[17071]_ ;
  assign \new_[17080]_  = A232 & ~A203;
  assign \new_[17084]_  = A267 & A265;
  assign \new_[17085]_  = A234 & \new_[17084]_ ;
  assign \new_[17086]_  = \new_[17085]_  & \new_[17080]_ ;
  assign \new_[17089]_  = A167 & A170;
  assign \new_[17093]_  = ~A202 & ~A201;
  assign \new_[17094]_  = ~A166 & \new_[17093]_ ;
  assign \new_[17095]_  = \new_[17094]_  & \new_[17089]_ ;
  assign \new_[17098]_  = A232 & ~A203;
  assign \new_[17102]_  = A267 & A266;
  assign \new_[17103]_  = A234 & \new_[17102]_ ;
  assign \new_[17104]_  = \new_[17103]_  & \new_[17098]_ ;
  assign \new_[17107]_  = A167 & A170;
  assign \new_[17111]_  = ~A202 & ~A201;
  assign \new_[17112]_  = ~A166 & \new_[17111]_ ;
  assign \new_[17113]_  = \new_[17112]_  & \new_[17107]_ ;
  assign \new_[17116]_  = A233 & ~A203;
  assign \new_[17120]_  = A300 & A299;
  assign \new_[17121]_  = A234 & \new_[17120]_ ;
  assign \new_[17122]_  = \new_[17121]_  & \new_[17116]_ ;
  assign \new_[17125]_  = A167 & A170;
  assign \new_[17129]_  = ~A202 & ~A201;
  assign \new_[17130]_  = ~A166 & \new_[17129]_ ;
  assign \new_[17131]_  = \new_[17130]_  & \new_[17125]_ ;
  assign \new_[17134]_  = A233 & ~A203;
  assign \new_[17138]_  = A300 & A298;
  assign \new_[17139]_  = A234 & \new_[17138]_ ;
  assign \new_[17140]_  = \new_[17139]_  & \new_[17134]_ ;
  assign \new_[17143]_  = A167 & A170;
  assign \new_[17147]_  = ~A202 & ~A201;
  assign \new_[17148]_  = ~A166 & \new_[17147]_ ;
  assign \new_[17149]_  = \new_[17148]_  & \new_[17143]_ ;
  assign \new_[17152]_  = A233 & ~A203;
  assign \new_[17156]_  = A267 & A265;
  assign \new_[17157]_  = A234 & \new_[17156]_ ;
  assign \new_[17158]_  = \new_[17157]_  & \new_[17152]_ ;
  assign \new_[17161]_  = A167 & A170;
  assign \new_[17165]_  = ~A202 & ~A201;
  assign \new_[17166]_  = ~A166 & \new_[17165]_ ;
  assign \new_[17167]_  = \new_[17166]_  & \new_[17161]_ ;
  assign \new_[17170]_  = A233 & ~A203;
  assign \new_[17174]_  = A267 & A266;
  assign \new_[17175]_  = A234 & \new_[17174]_ ;
  assign \new_[17176]_  = \new_[17175]_  & \new_[17170]_ ;
  assign \new_[17179]_  = A167 & A170;
  assign \new_[17183]_  = ~A202 & ~A201;
  assign \new_[17184]_  = ~A166 & \new_[17183]_ ;
  assign \new_[17185]_  = \new_[17184]_  & \new_[17179]_ ;
  assign \new_[17188]_  = ~A232 & ~A203;
  assign \new_[17192]_  = A301 & A236;
  assign \new_[17193]_  = A233 & \new_[17192]_ ;
  assign \new_[17194]_  = \new_[17193]_  & \new_[17188]_ ;
  assign \new_[17197]_  = A167 & A170;
  assign \new_[17201]_  = ~A202 & ~A201;
  assign \new_[17202]_  = ~A166 & \new_[17201]_ ;
  assign \new_[17203]_  = \new_[17202]_  & \new_[17197]_ ;
  assign \new_[17206]_  = ~A232 & ~A203;
  assign \new_[17210]_  = A268 & A236;
  assign \new_[17211]_  = A233 & \new_[17210]_ ;
  assign \new_[17212]_  = \new_[17211]_  & \new_[17206]_ ;
  assign \new_[17215]_  = A167 & A170;
  assign \new_[17219]_  = ~A202 & ~A201;
  assign \new_[17220]_  = ~A166 & \new_[17219]_ ;
  assign \new_[17221]_  = \new_[17220]_  & \new_[17215]_ ;
  assign \new_[17224]_  = A232 & ~A203;
  assign \new_[17228]_  = A301 & A236;
  assign \new_[17229]_  = ~A233 & \new_[17228]_ ;
  assign \new_[17230]_  = \new_[17229]_  & \new_[17224]_ ;
  assign \new_[17233]_  = A167 & A170;
  assign \new_[17237]_  = ~A202 & ~A201;
  assign \new_[17238]_  = ~A166 & \new_[17237]_ ;
  assign \new_[17239]_  = \new_[17238]_  & \new_[17233]_ ;
  assign \new_[17242]_  = A232 & ~A203;
  assign \new_[17246]_  = A268 & A236;
  assign \new_[17247]_  = ~A233 & \new_[17246]_ ;
  assign \new_[17248]_  = \new_[17247]_  & \new_[17242]_ ;
  assign \new_[17251]_  = A167 & A170;
  assign \new_[17255]_  = A200 & A199;
  assign \new_[17256]_  = ~A166 & \new_[17255]_ ;
  assign \new_[17257]_  = \new_[17256]_  & \new_[17251]_ ;
  assign \new_[17260]_  = ~A202 & ~A201;
  assign \new_[17264]_  = A300 & A299;
  assign \new_[17265]_  = A235 & \new_[17264]_ ;
  assign \new_[17266]_  = \new_[17265]_  & \new_[17260]_ ;
  assign \new_[17269]_  = A167 & A170;
  assign \new_[17273]_  = A200 & A199;
  assign \new_[17274]_  = ~A166 & \new_[17273]_ ;
  assign \new_[17275]_  = \new_[17274]_  & \new_[17269]_ ;
  assign \new_[17278]_  = ~A202 & ~A201;
  assign \new_[17282]_  = A300 & A298;
  assign \new_[17283]_  = A235 & \new_[17282]_ ;
  assign \new_[17284]_  = \new_[17283]_  & \new_[17278]_ ;
  assign \new_[17287]_  = A167 & A170;
  assign \new_[17291]_  = A200 & A199;
  assign \new_[17292]_  = ~A166 & \new_[17291]_ ;
  assign \new_[17293]_  = \new_[17292]_  & \new_[17287]_ ;
  assign \new_[17296]_  = ~A202 & ~A201;
  assign \new_[17300]_  = A267 & A265;
  assign \new_[17301]_  = A235 & \new_[17300]_ ;
  assign \new_[17302]_  = \new_[17301]_  & \new_[17296]_ ;
  assign \new_[17305]_  = A167 & A170;
  assign \new_[17309]_  = A200 & A199;
  assign \new_[17310]_  = ~A166 & \new_[17309]_ ;
  assign \new_[17311]_  = \new_[17310]_  & \new_[17305]_ ;
  assign \new_[17314]_  = ~A202 & ~A201;
  assign \new_[17318]_  = A267 & A266;
  assign \new_[17319]_  = A235 & \new_[17318]_ ;
  assign \new_[17320]_  = \new_[17319]_  & \new_[17314]_ ;
  assign \new_[17323]_  = A167 & A170;
  assign \new_[17327]_  = A200 & A199;
  assign \new_[17328]_  = ~A166 & \new_[17327]_ ;
  assign \new_[17329]_  = \new_[17328]_  & \new_[17323]_ ;
  assign \new_[17332]_  = ~A202 & ~A201;
  assign \new_[17336]_  = A301 & A234;
  assign \new_[17337]_  = A232 & \new_[17336]_ ;
  assign \new_[17338]_  = \new_[17337]_  & \new_[17332]_ ;
  assign \new_[17341]_  = A167 & A170;
  assign \new_[17345]_  = A200 & A199;
  assign \new_[17346]_  = ~A166 & \new_[17345]_ ;
  assign \new_[17347]_  = \new_[17346]_  & \new_[17341]_ ;
  assign \new_[17350]_  = ~A202 & ~A201;
  assign \new_[17354]_  = A268 & A234;
  assign \new_[17355]_  = A232 & \new_[17354]_ ;
  assign \new_[17356]_  = \new_[17355]_  & \new_[17350]_ ;
  assign \new_[17359]_  = A167 & A170;
  assign \new_[17363]_  = A200 & A199;
  assign \new_[17364]_  = ~A166 & \new_[17363]_ ;
  assign \new_[17365]_  = \new_[17364]_  & \new_[17359]_ ;
  assign \new_[17368]_  = ~A202 & ~A201;
  assign \new_[17372]_  = A301 & A234;
  assign \new_[17373]_  = A233 & \new_[17372]_ ;
  assign \new_[17374]_  = \new_[17373]_  & \new_[17368]_ ;
  assign \new_[17377]_  = A167 & A170;
  assign \new_[17381]_  = A200 & A199;
  assign \new_[17382]_  = ~A166 & \new_[17381]_ ;
  assign \new_[17383]_  = \new_[17382]_  & \new_[17377]_ ;
  assign \new_[17386]_  = ~A202 & ~A201;
  assign \new_[17390]_  = A268 & A234;
  assign \new_[17391]_  = A233 & \new_[17390]_ ;
  assign \new_[17392]_  = \new_[17391]_  & \new_[17386]_ ;
  assign \new_[17395]_  = A167 & A170;
  assign \new_[17399]_  = ~A200 & ~A199;
  assign \new_[17400]_  = ~A166 & \new_[17399]_ ;
  assign \new_[17401]_  = \new_[17400]_  & \new_[17395]_ ;
  assign \new_[17404]_  = A235 & ~A202;
  assign \new_[17408]_  = A302 & ~A299;
  assign \new_[17409]_  = A298 & \new_[17408]_ ;
  assign \new_[17410]_  = \new_[17409]_  & \new_[17404]_ ;
  assign \new_[17413]_  = A167 & A170;
  assign \new_[17417]_  = ~A200 & ~A199;
  assign \new_[17418]_  = ~A166 & \new_[17417]_ ;
  assign \new_[17419]_  = \new_[17418]_  & \new_[17413]_ ;
  assign \new_[17422]_  = A235 & ~A202;
  assign \new_[17426]_  = A302 & A299;
  assign \new_[17427]_  = ~A298 & \new_[17426]_ ;
  assign \new_[17428]_  = \new_[17427]_  & \new_[17422]_ ;
  assign \new_[17431]_  = A167 & A170;
  assign \new_[17435]_  = ~A200 & ~A199;
  assign \new_[17436]_  = ~A166 & \new_[17435]_ ;
  assign \new_[17437]_  = \new_[17436]_  & \new_[17431]_ ;
  assign \new_[17440]_  = A235 & ~A202;
  assign \new_[17444]_  = A269 & A266;
  assign \new_[17445]_  = ~A265 & \new_[17444]_ ;
  assign \new_[17446]_  = \new_[17445]_  & \new_[17440]_ ;
  assign \new_[17449]_  = A167 & A170;
  assign \new_[17453]_  = ~A200 & ~A199;
  assign \new_[17454]_  = ~A166 & \new_[17453]_ ;
  assign \new_[17455]_  = \new_[17454]_  & \new_[17449]_ ;
  assign \new_[17458]_  = A235 & ~A202;
  assign \new_[17462]_  = A269 & ~A266;
  assign \new_[17463]_  = A265 & \new_[17462]_ ;
  assign \new_[17464]_  = \new_[17463]_  & \new_[17458]_ ;
  assign \new_[17467]_  = A167 & A170;
  assign \new_[17471]_  = ~A200 & ~A199;
  assign \new_[17472]_  = ~A166 & \new_[17471]_ ;
  assign \new_[17473]_  = \new_[17472]_  & \new_[17467]_ ;
  assign \new_[17476]_  = A232 & ~A202;
  assign \new_[17480]_  = A300 & A299;
  assign \new_[17481]_  = A234 & \new_[17480]_ ;
  assign \new_[17482]_  = \new_[17481]_  & \new_[17476]_ ;
  assign \new_[17485]_  = A167 & A170;
  assign \new_[17489]_  = ~A200 & ~A199;
  assign \new_[17490]_  = ~A166 & \new_[17489]_ ;
  assign \new_[17491]_  = \new_[17490]_  & \new_[17485]_ ;
  assign \new_[17494]_  = A232 & ~A202;
  assign \new_[17498]_  = A300 & A298;
  assign \new_[17499]_  = A234 & \new_[17498]_ ;
  assign \new_[17500]_  = \new_[17499]_  & \new_[17494]_ ;
  assign \new_[17503]_  = A167 & A170;
  assign \new_[17507]_  = ~A200 & ~A199;
  assign \new_[17508]_  = ~A166 & \new_[17507]_ ;
  assign \new_[17509]_  = \new_[17508]_  & \new_[17503]_ ;
  assign \new_[17512]_  = A232 & ~A202;
  assign \new_[17516]_  = A267 & A265;
  assign \new_[17517]_  = A234 & \new_[17516]_ ;
  assign \new_[17518]_  = \new_[17517]_  & \new_[17512]_ ;
  assign \new_[17521]_  = A167 & A170;
  assign \new_[17525]_  = ~A200 & ~A199;
  assign \new_[17526]_  = ~A166 & \new_[17525]_ ;
  assign \new_[17527]_  = \new_[17526]_  & \new_[17521]_ ;
  assign \new_[17530]_  = A232 & ~A202;
  assign \new_[17534]_  = A267 & A266;
  assign \new_[17535]_  = A234 & \new_[17534]_ ;
  assign \new_[17536]_  = \new_[17535]_  & \new_[17530]_ ;
  assign \new_[17539]_  = A167 & A170;
  assign \new_[17543]_  = ~A200 & ~A199;
  assign \new_[17544]_  = ~A166 & \new_[17543]_ ;
  assign \new_[17545]_  = \new_[17544]_  & \new_[17539]_ ;
  assign \new_[17548]_  = A233 & ~A202;
  assign \new_[17552]_  = A300 & A299;
  assign \new_[17553]_  = A234 & \new_[17552]_ ;
  assign \new_[17554]_  = \new_[17553]_  & \new_[17548]_ ;
  assign \new_[17557]_  = A167 & A170;
  assign \new_[17561]_  = ~A200 & ~A199;
  assign \new_[17562]_  = ~A166 & \new_[17561]_ ;
  assign \new_[17563]_  = \new_[17562]_  & \new_[17557]_ ;
  assign \new_[17566]_  = A233 & ~A202;
  assign \new_[17570]_  = A300 & A298;
  assign \new_[17571]_  = A234 & \new_[17570]_ ;
  assign \new_[17572]_  = \new_[17571]_  & \new_[17566]_ ;
  assign \new_[17575]_  = A167 & A170;
  assign \new_[17579]_  = ~A200 & ~A199;
  assign \new_[17580]_  = ~A166 & \new_[17579]_ ;
  assign \new_[17581]_  = \new_[17580]_  & \new_[17575]_ ;
  assign \new_[17584]_  = A233 & ~A202;
  assign \new_[17588]_  = A267 & A265;
  assign \new_[17589]_  = A234 & \new_[17588]_ ;
  assign \new_[17590]_  = \new_[17589]_  & \new_[17584]_ ;
  assign \new_[17593]_  = A167 & A170;
  assign \new_[17597]_  = ~A200 & ~A199;
  assign \new_[17598]_  = ~A166 & \new_[17597]_ ;
  assign \new_[17599]_  = \new_[17598]_  & \new_[17593]_ ;
  assign \new_[17602]_  = A233 & ~A202;
  assign \new_[17606]_  = A267 & A266;
  assign \new_[17607]_  = A234 & \new_[17606]_ ;
  assign \new_[17608]_  = \new_[17607]_  & \new_[17602]_ ;
  assign \new_[17611]_  = A167 & A170;
  assign \new_[17615]_  = ~A200 & ~A199;
  assign \new_[17616]_  = ~A166 & \new_[17615]_ ;
  assign \new_[17617]_  = \new_[17616]_  & \new_[17611]_ ;
  assign \new_[17620]_  = ~A232 & ~A202;
  assign \new_[17624]_  = A301 & A236;
  assign \new_[17625]_  = A233 & \new_[17624]_ ;
  assign \new_[17626]_  = \new_[17625]_  & \new_[17620]_ ;
  assign \new_[17629]_  = A167 & A170;
  assign \new_[17633]_  = ~A200 & ~A199;
  assign \new_[17634]_  = ~A166 & \new_[17633]_ ;
  assign \new_[17635]_  = \new_[17634]_  & \new_[17629]_ ;
  assign \new_[17638]_  = ~A232 & ~A202;
  assign \new_[17642]_  = A268 & A236;
  assign \new_[17643]_  = A233 & \new_[17642]_ ;
  assign \new_[17644]_  = \new_[17643]_  & \new_[17638]_ ;
  assign \new_[17647]_  = A167 & A170;
  assign \new_[17651]_  = ~A200 & ~A199;
  assign \new_[17652]_  = ~A166 & \new_[17651]_ ;
  assign \new_[17653]_  = \new_[17652]_  & \new_[17647]_ ;
  assign \new_[17656]_  = A232 & ~A202;
  assign \new_[17660]_  = A301 & A236;
  assign \new_[17661]_  = ~A233 & \new_[17660]_ ;
  assign \new_[17662]_  = \new_[17661]_  & \new_[17656]_ ;
  assign \new_[17665]_  = A167 & A170;
  assign \new_[17669]_  = ~A200 & ~A199;
  assign \new_[17670]_  = ~A166 & \new_[17669]_ ;
  assign \new_[17671]_  = \new_[17670]_  & \new_[17665]_ ;
  assign \new_[17674]_  = A232 & ~A202;
  assign \new_[17678]_  = A268 & A236;
  assign \new_[17679]_  = ~A233 & \new_[17678]_ ;
  assign \new_[17680]_  = \new_[17679]_  & \new_[17674]_ ;
  assign \new_[17683]_  = ~A167 & A170;
  assign \new_[17687]_  = ~A202 & ~A201;
  assign \new_[17688]_  = A166 & \new_[17687]_ ;
  assign \new_[17689]_  = \new_[17688]_  & \new_[17683]_ ;
  assign \new_[17692]_  = A235 & ~A203;
  assign \new_[17696]_  = A302 & ~A299;
  assign \new_[17697]_  = A298 & \new_[17696]_ ;
  assign \new_[17698]_  = \new_[17697]_  & \new_[17692]_ ;
  assign \new_[17701]_  = ~A167 & A170;
  assign \new_[17705]_  = ~A202 & ~A201;
  assign \new_[17706]_  = A166 & \new_[17705]_ ;
  assign \new_[17707]_  = \new_[17706]_  & \new_[17701]_ ;
  assign \new_[17710]_  = A235 & ~A203;
  assign \new_[17714]_  = A302 & A299;
  assign \new_[17715]_  = ~A298 & \new_[17714]_ ;
  assign \new_[17716]_  = \new_[17715]_  & \new_[17710]_ ;
  assign \new_[17719]_  = ~A167 & A170;
  assign \new_[17723]_  = ~A202 & ~A201;
  assign \new_[17724]_  = A166 & \new_[17723]_ ;
  assign \new_[17725]_  = \new_[17724]_  & \new_[17719]_ ;
  assign \new_[17728]_  = A235 & ~A203;
  assign \new_[17732]_  = A269 & A266;
  assign \new_[17733]_  = ~A265 & \new_[17732]_ ;
  assign \new_[17734]_  = \new_[17733]_  & \new_[17728]_ ;
  assign \new_[17737]_  = ~A167 & A170;
  assign \new_[17741]_  = ~A202 & ~A201;
  assign \new_[17742]_  = A166 & \new_[17741]_ ;
  assign \new_[17743]_  = \new_[17742]_  & \new_[17737]_ ;
  assign \new_[17746]_  = A235 & ~A203;
  assign \new_[17750]_  = A269 & ~A266;
  assign \new_[17751]_  = A265 & \new_[17750]_ ;
  assign \new_[17752]_  = \new_[17751]_  & \new_[17746]_ ;
  assign \new_[17755]_  = ~A167 & A170;
  assign \new_[17759]_  = ~A202 & ~A201;
  assign \new_[17760]_  = A166 & \new_[17759]_ ;
  assign \new_[17761]_  = \new_[17760]_  & \new_[17755]_ ;
  assign \new_[17764]_  = A232 & ~A203;
  assign \new_[17768]_  = A300 & A299;
  assign \new_[17769]_  = A234 & \new_[17768]_ ;
  assign \new_[17770]_  = \new_[17769]_  & \new_[17764]_ ;
  assign \new_[17773]_  = ~A167 & A170;
  assign \new_[17777]_  = ~A202 & ~A201;
  assign \new_[17778]_  = A166 & \new_[17777]_ ;
  assign \new_[17779]_  = \new_[17778]_  & \new_[17773]_ ;
  assign \new_[17782]_  = A232 & ~A203;
  assign \new_[17786]_  = A300 & A298;
  assign \new_[17787]_  = A234 & \new_[17786]_ ;
  assign \new_[17788]_  = \new_[17787]_  & \new_[17782]_ ;
  assign \new_[17791]_  = ~A167 & A170;
  assign \new_[17795]_  = ~A202 & ~A201;
  assign \new_[17796]_  = A166 & \new_[17795]_ ;
  assign \new_[17797]_  = \new_[17796]_  & \new_[17791]_ ;
  assign \new_[17800]_  = A232 & ~A203;
  assign \new_[17804]_  = A267 & A265;
  assign \new_[17805]_  = A234 & \new_[17804]_ ;
  assign \new_[17806]_  = \new_[17805]_  & \new_[17800]_ ;
  assign \new_[17809]_  = ~A167 & A170;
  assign \new_[17813]_  = ~A202 & ~A201;
  assign \new_[17814]_  = A166 & \new_[17813]_ ;
  assign \new_[17815]_  = \new_[17814]_  & \new_[17809]_ ;
  assign \new_[17818]_  = A232 & ~A203;
  assign \new_[17822]_  = A267 & A266;
  assign \new_[17823]_  = A234 & \new_[17822]_ ;
  assign \new_[17824]_  = \new_[17823]_  & \new_[17818]_ ;
  assign \new_[17827]_  = ~A167 & A170;
  assign \new_[17831]_  = ~A202 & ~A201;
  assign \new_[17832]_  = A166 & \new_[17831]_ ;
  assign \new_[17833]_  = \new_[17832]_  & \new_[17827]_ ;
  assign \new_[17836]_  = A233 & ~A203;
  assign \new_[17840]_  = A300 & A299;
  assign \new_[17841]_  = A234 & \new_[17840]_ ;
  assign \new_[17842]_  = \new_[17841]_  & \new_[17836]_ ;
  assign \new_[17845]_  = ~A167 & A170;
  assign \new_[17849]_  = ~A202 & ~A201;
  assign \new_[17850]_  = A166 & \new_[17849]_ ;
  assign \new_[17851]_  = \new_[17850]_  & \new_[17845]_ ;
  assign \new_[17854]_  = A233 & ~A203;
  assign \new_[17858]_  = A300 & A298;
  assign \new_[17859]_  = A234 & \new_[17858]_ ;
  assign \new_[17860]_  = \new_[17859]_  & \new_[17854]_ ;
  assign \new_[17863]_  = ~A167 & A170;
  assign \new_[17867]_  = ~A202 & ~A201;
  assign \new_[17868]_  = A166 & \new_[17867]_ ;
  assign \new_[17869]_  = \new_[17868]_  & \new_[17863]_ ;
  assign \new_[17872]_  = A233 & ~A203;
  assign \new_[17876]_  = A267 & A265;
  assign \new_[17877]_  = A234 & \new_[17876]_ ;
  assign \new_[17878]_  = \new_[17877]_  & \new_[17872]_ ;
  assign \new_[17881]_  = ~A167 & A170;
  assign \new_[17885]_  = ~A202 & ~A201;
  assign \new_[17886]_  = A166 & \new_[17885]_ ;
  assign \new_[17887]_  = \new_[17886]_  & \new_[17881]_ ;
  assign \new_[17890]_  = A233 & ~A203;
  assign \new_[17894]_  = A267 & A266;
  assign \new_[17895]_  = A234 & \new_[17894]_ ;
  assign \new_[17896]_  = \new_[17895]_  & \new_[17890]_ ;
  assign \new_[17899]_  = ~A167 & A170;
  assign \new_[17903]_  = ~A202 & ~A201;
  assign \new_[17904]_  = A166 & \new_[17903]_ ;
  assign \new_[17905]_  = \new_[17904]_  & \new_[17899]_ ;
  assign \new_[17908]_  = ~A232 & ~A203;
  assign \new_[17912]_  = A301 & A236;
  assign \new_[17913]_  = A233 & \new_[17912]_ ;
  assign \new_[17914]_  = \new_[17913]_  & \new_[17908]_ ;
  assign \new_[17917]_  = ~A167 & A170;
  assign \new_[17921]_  = ~A202 & ~A201;
  assign \new_[17922]_  = A166 & \new_[17921]_ ;
  assign \new_[17923]_  = \new_[17922]_  & \new_[17917]_ ;
  assign \new_[17926]_  = ~A232 & ~A203;
  assign \new_[17930]_  = A268 & A236;
  assign \new_[17931]_  = A233 & \new_[17930]_ ;
  assign \new_[17932]_  = \new_[17931]_  & \new_[17926]_ ;
  assign \new_[17935]_  = ~A167 & A170;
  assign \new_[17939]_  = ~A202 & ~A201;
  assign \new_[17940]_  = A166 & \new_[17939]_ ;
  assign \new_[17941]_  = \new_[17940]_  & \new_[17935]_ ;
  assign \new_[17944]_  = A232 & ~A203;
  assign \new_[17948]_  = A301 & A236;
  assign \new_[17949]_  = ~A233 & \new_[17948]_ ;
  assign \new_[17950]_  = \new_[17949]_  & \new_[17944]_ ;
  assign \new_[17953]_  = ~A167 & A170;
  assign \new_[17957]_  = ~A202 & ~A201;
  assign \new_[17958]_  = A166 & \new_[17957]_ ;
  assign \new_[17959]_  = \new_[17958]_  & \new_[17953]_ ;
  assign \new_[17962]_  = A232 & ~A203;
  assign \new_[17966]_  = A268 & A236;
  assign \new_[17967]_  = ~A233 & \new_[17966]_ ;
  assign \new_[17968]_  = \new_[17967]_  & \new_[17962]_ ;
  assign \new_[17971]_  = ~A167 & A170;
  assign \new_[17975]_  = A200 & A199;
  assign \new_[17976]_  = A166 & \new_[17975]_ ;
  assign \new_[17977]_  = \new_[17976]_  & \new_[17971]_ ;
  assign \new_[17980]_  = ~A202 & ~A201;
  assign \new_[17984]_  = A300 & A299;
  assign \new_[17985]_  = A235 & \new_[17984]_ ;
  assign \new_[17986]_  = \new_[17985]_  & \new_[17980]_ ;
  assign \new_[17989]_  = ~A167 & A170;
  assign \new_[17993]_  = A200 & A199;
  assign \new_[17994]_  = A166 & \new_[17993]_ ;
  assign \new_[17995]_  = \new_[17994]_  & \new_[17989]_ ;
  assign \new_[17998]_  = ~A202 & ~A201;
  assign \new_[18002]_  = A300 & A298;
  assign \new_[18003]_  = A235 & \new_[18002]_ ;
  assign \new_[18004]_  = \new_[18003]_  & \new_[17998]_ ;
  assign \new_[18007]_  = ~A167 & A170;
  assign \new_[18011]_  = A200 & A199;
  assign \new_[18012]_  = A166 & \new_[18011]_ ;
  assign \new_[18013]_  = \new_[18012]_  & \new_[18007]_ ;
  assign \new_[18016]_  = ~A202 & ~A201;
  assign \new_[18020]_  = A267 & A265;
  assign \new_[18021]_  = A235 & \new_[18020]_ ;
  assign \new_[18022]_  = \new_[18021]_  & \new_[18016]_ ;
  assign \new_[18025]_  = ~A167 & A170;
  assign \new_[18029]_  = A200 & A199;
  assign \new_[18030]_  = A166 & \new_[18029]_ ;
  assign \new_[18031]_  = \new_[18030]_  & \new_[18025]_ ;
  assign \new_[18034]_  = ~A202 & ~A201;
  assign \new_[18038]_  = A267 & A266;
  assign \new_[18039]_  = A235 & \new_[18038]_ ;
  assign \new_[18040]_  = \new_[18039]_  & \new_[18034]_ ;
  assign \new_[18043]_  = ~A167 & A170;
  assign \new_[18047]_  = A200 & A199;
  assign \new_[18048]_  = A166 & \new_[18047]_ ;
  assign \new_[18049]_  = \new_[18048]_  & \new_[18043]_ ;
  assign \new_[18052]_  = ~A202 & ~A201;
  assign \new_[18056]_  = A301 & A234;
  assign \new_[18057]_  = A232 & \new_[18056]_ ;
  assign \new_[18058]_  = \new_[18057]_  & \new_[18052]_ ;
  assign \new_[18061]_  = ~A167 & A170;
  assign \new_[18065]_  = A200 & A199;
  assign \new_[18066]_  = A166 & \new_[18065]_ ;
  assign \new_[18067]_  = \new_[18066]_  & \new_[18061]_ ;
  assign \new_[18070]_  = ~A202 & ~A201;
  assign \new_[18074]_  = A268 & A234;
  assign \new_[18075]_  = A232 & \new_[18074]_ ;
  assign \new_[18076]_  = \new_[18075]_  & \new_[18070]_ ;
  assign \new_[18079]_  = ~A167 & A170;
  assign \new_[18083]_  = A200 & A199;
  assign \new_[18084]_  = A166 & \new_[18083]_ ;
  assign \new_[18085]_  = \new_[18084]_  & \new_[18079]_ ;
  assign \new_[18088]_  = ~A202 & ~A201;
  assign \new_[18092]_  = A301 & A234;
  assign \new_[18093]_  = A233 & \new_[18092]_ ;
  assign \new_[18094]_  = \new_[18093]_  & \new_[18088]_ ;
  assign \new_[18097]_  = ~A167 & A170;
  assign \new_[18101]_  = A200 & A199;
  assign \new_[18102]_  = A166 & \new_[18101]_ ;
  assign \new_[18103]_  = \new_[18102]_  & \new_[18097]_ ;
  assign \new_[18106]_  = ~A202 & ~A201;
  assign \new_[18110]_  = A268 & A234;
  assign \new_[18111]_  = A233 & \new_[18110]_ ;
  assign \new_[18112]_  = \new_[18111]_  & \new_[18106]_ ;
  assign \new_[18115]_  = ~A167 & A170;
  assign \new_[18119]_  = ~A200 & ~A199;
  assign \new_[18120]_  = A166 & \new_[18119]_ ;
  assign \new_[18121]_  = \new_[18120]_  & \new_[18115]_ ;
  assign \new_[18124]_  = A235 & ~A202;
  assign \new_[18128]_  = A302 & ~A299;
  assign \new_[18129]_  = A298 & \new_[18128]_ ;
  assign \new_[18130]_  = \new_[18129]_  & \new_[18124]_ ;
  assign \new_[18133]_  = ~A167 & A170;
  assign \new_[18137]_  = ~A200 & ~A199;
  assign \new_[18138]_  = A166 & \new_[18137]_ ;
  assign \new_[18139]_  = \new_[18138]_  & \new_[18133]_ ;
  assign \new_[18142]_  = A235 & ~A202;
  assign \new_[18146]_  = A302 & A299;
  assign \new_[18147]_  = ~A298 & \new_[18146]_ ;
  assign \new_[18148]_  = \new_[18147]_  & \new_[18142]_ ;
  assign \new_[18151]_  = ~A167 & A170;
  assign \new_[18155]_  = ~A200 & ~A199;
  assign \new_[18156]_  = A166 & \new_[18155]_ ;
  assign \new_[18157]_  = \new_[18156]_  & \new_[18151]_ ;
  assign \new_[18160]_  = A235 & ~A202;
  assign \new_[18164]_  = A269 & A266;
  assign \new_[18165]_  = ~A265 & \new_[18164]_ ;
  assign \new_[18166]_  = \new_[18165]_  & \new_[18160]_ ;
  assign \new_[18169]_  = ~A167 & A170;
  assign \new_[18173]_  = ~A200 & ~A199;
  assign \new_[18174]_  = A166 & \new_[18173]_ ;
  assign \new_[18175]_  = \new_[18174]_  & \new_[18169]_ ;
  assign \new_[18178]_  = A235 & ~A202;
  assign \new_[18182]_  = A269 & ~A266;
  assign \new_[18183]_  = A265 & \new_[18182]_ ;
  assign \new_[18184]_  = \new_[18183]_  & \new_[18178]_ ;
  assign \new_[18187]_  = ~A167 & A170;
  assign \new_[18191]_  = ~A200 & ~A199;
  assign \new_[18192]_  = A166 & \new_[18191]_ ;
  assign \new_[18193]_  = \new_[18192]_  & \new_[18187]_ ;
  assign \new_[18196]_  = A232 & ~A202;
  assign \new_[18200]_  = A300 & A299;
  assign \new_[18201]_  = A234 & \new_[18200]_ ;
  assign \new_[18202]_  = \new_[18201]_  & \new_[18196]_ ;
  assign \new_[18205]_  = ~A167 & A170;
  assign \new_[18209]_  = ~A200 & ~A199;
  assign \new_[18210]_  = A166 & \new_[18209]_ ;
  assign \new_[18211]_  = \new_[18210]_  & \new_[18205]_ ;
  assign \new_[18214]_  = A232 & ~A202;
  assign \new_[18218]_  = A300 & A298;
  assign \new_[18219]_  = A234 & \new_[18218]_ ;
  assign \new_[18220]_  = \new_[18219]_  & \new_[18214]_ ;
  assign \new_[18223]_  = ~A167 & A170;
  assign \new_[18227]_  = ~A200 & ~A199;
  assign \new_[18228]_  = A166 & \new_[18227]_ ;
  assign \new_[18229]_  = \new_[18228]_  & \new_[18223]_ ;
  assign \new_[18232]_  = A232 & ~A202;
  assign \new_[18236]_  = A267 & A265;
  assign \new_[18237]_  = A234 & \new_[18236]_ ;
  assign \new_[18238]_  = \new_[18237]_  & \new_[18232]_ ;
  assign \new_[18241]_  = ~A167 & A170;
  assign \new_[18245]_  = ~A200 & ~A199;
  assign \new_[18246]_  = A166 & \new_[18245]_ ;
  assign \new_[18247]_  = \new_[18246]_  & \new_[18241]_ ;
  assign \new_[18250]_  = A232 & ~A202;
  assign \new_[18254]_  = A267 & A266;
  assign \new_[18255]_  = A234 & \new_[18254]_ ;
  assign \new_[18256]_  = \new_[18255]_  & \new_[18250]_ ;
  assign \new_[18259]_  = ~A167 & A170;
  assign \new_[18263]_  = ~A200 & ~A199;
  assign \new_[18264]_  = A166 & \new_[18263]_ ;
  assign \new_[18265]_  = \new_[18264]_  & \new_[18259]_ ;
  assign \new_[18268]_  = A233 & ~A202;
  assign \new_[18272]_  = A300 & A299;
  assign \new_[18273]_  = A234 & \new_[18272]_ ;
  assign \new_[18274]_  = \new_[18273]_  & \new_[18268]_ ;
  assign \new_[18277]_  = ~A167 & A170;
  assign \new_[18281]_  = ~A200 & ~A199;
  assign \new_[18282]_  = A166 & \new_[18281]_ ;
  assign \new_[18283]_  = \new_[18282]_  & \new_[18277]_ ;
  assign \new_[18286]_  = A233 & ~A202;
  assign \new_[18290]_  = A300 & A298;
  assign \new_[18291]_  = A234 & \new_[18290]_ ;
  assign \new_[18292]_  = \new_[18291]_  & \new_[18286]_ ;
  assign \new_[18295]_  = ~A167 & A170;
  assign \new_[18299]_  = ~A200 & ~A199;
  assign \new_[18300]_  = A166 & \new_[18299]_ ;
  assign \new_[18301]_  = \new_[18300]_  & \new_[18295]_ ;
  assign \new_[18304]_  = A233 & ~A202;
  assign \new_[18308]_  = A267 & A265;
  assign \new_[18309]_  = A234 & \new_[18308]_ ;
  assign \new_[18310]_  = \new_[18309]_  & \new_[18304]_ ;
  assign \new_[18313]_  = ~A167 & A170;
  assign \new_[18317]_  = ~A200 & ~A199;
  assign \new_[18318]_  = A166 & \new_[18317]_ ;
  assign \new_[18319]_  = \new_[18318]_  & \new_[18313]_ ;
  assign \new_[18322]_  = A233 & ~A202;
  assign \new_[18326]_  = A267 & A266;
  assign \new_[18327]_  = A234 & \new_[18326]_ ;
  assign \new_[18328]_  = \new_[18327]_  & \new_[18322]_ ;
  assign \new_[18331]_  = ~A167 & A170;
  assign \new_[18335]_  = ~A200 & ~A199;
  assign \new_[18336]_  = A166 & \new_[18335]_ ;
  assign \new_[18337]_  = \new_[18336]_  & \new_[18331]_ ;
  assign \new_[18340]_  = ~A232 & ~A202;
  assign \new_[18344]_  = A301 & A236;
  assign \new_[18345]_  = A233 & \new_[18344]_ ;
  assign \new_[18346]_  = \new_[18345]_  & \new_[18340]_ ;
  assign \new_[18349]_  = ~A167 & A170;
  assign \new_[18353]_  = ~A200 & ~A199;
  assign \new_[18354]_  = A166 & \new_[18353]_ ;
  assign \new_[18355]_  = \new_[18354]_  & \new_[18349]_ ;
  assign \new_[18358]_  = ~A232 & ~A202;
  assign \new_[18362]_  = A268 & A236;
  assign \new_[18363]_  = A233 & \new_[18362]_ ;
  assign \new_[18364]_  = \new_[18363]_  & \new_[18358]_ ;
  assign \new_[18367]_  = ~A167 & A170;
  assign \new_[18371]_  = ~A200 & ~A199;
  assign \new_[18372]_  = A166 & \new_[18371]_ ;
  assign \new_[18373]_  = \new_[18372]_  & \new_[18367]_ ;
  assign \new_[18376]_  = A232 & ~A202;
  assign \new_[18380]_  = A301 & A236;
  assign \new_[18381]_  = ~A233 & \new_[18380]_ ;
  assign \new_[18382]_  = \new_[18381]_  & \new_[18376]_ ;
  assign \new_[18385]_  = ~A167 & A170;
  assign \new_[18389]_  = ~A200 & ~A199;
  assign \new_[18390]_  = A166 & \new_[18389]_ ;
  assign \new_[18391]_  = \new_[18390]_  & \new_[18385]_ ;
  assign \new_[18394]_  = A232 & ~A202;
  assign \new_[18398]_  = A268 & A236;
  assign \new_[18399]_  = ~A233 & \new_[18398]_ ;
  assign \new_[18400]_  = \new_[18399]_  & \new_[18394]_ ;
  assign \new_[18403]_  = ~A201 & A169;
  assign \new_[18407]_  = ~A232 & ~A203;
  assign \new_[18408]_  = ~A202 & \new_[18407]_ ;
  assign \new_[18409]_  = \new_[18408]_  & \new_[18403]_ ;
  assign \new_[18412]_  = A236 & A233;
  assign \new_[18416]_  = A302 & ~A299;
  assign \new_[18417]_  = A298 & \new_[18416]_ ;
  assign \new_[18418]_  = \new_[18417]_  & \new_[18412]_ ;
  assign \new_[18421]_  = ~A201 & A169;
  assign \new_[18425]_  = ~A232 & ~A203;
  assign \new_[18426]_  = ~A202 & \new_[18425]_ ;
  assign \new_[18427]_  = \new_[18426]_  & \new_[18421]_ ;
  assign \new_[18430]_  = A236 & A233;
  assign \new_[18434]_  = A302 & A299;
  assign \new_[18435]_  = ~A298 & \new_[18434]_ ;
  assign \new_[18436]_  = \new_[18435]_  & \new_[18430]_ ;
  assign \new_[18439]_  = ~A201 & A169;
  assign \new_[18443]_  = ~A232 & ~A203;
  assign \new_[18444]_  = ~A202 & \new_[18443]_ ;
  assign \new_[18445]_  = \new_[18444]_  & \new_[18439]_ ;
  assign \new_[18448]_  = A236 & A233;
  assign \new_[18452]_  = A269 & A266;
  assign \new_[18453]_  = ~A265 & \new_[18452]_ ;
  assign \new_[18454]_  = \new_[18453]_  & \new_[18448]_ ;
  assign \new_[18457]_  = ~A201 & A169;
  assign \new_[18461]_  = ~A232 & ~A203;
  assign \new_[18462]_  = ~A202 & \new_[18461]_ ;
  assign \new_[18463]_  = \new_[18462]_  & \new_[18457]_ ;
  assign \new_[18466]_  = A236 & A233;
  assign \new_[18470]_  = A269 & ~A266;
  assign \new_[18471]_  = A265 & \new_[18470]_ ;
  assign \new_[18472]_  = \new_[18471]_  & \new_[18466]_ ;
  assign \new_[18475]_  = ~A201 & A169;
  assign \new_[18479]_  = A232 & ~A203;
  assign \new_[18480]_  = ~A202 & \new_[18479]_ ;
  assign \new_[18481]_  = \new_[18480]_  & \new_[18475]_ ;
  assign \new_[18484]_  = A236 & ~A233;
  assign \new_[18488]_  = A302 & ~A299;
  assign \new_[18489]_  = A298 & \new_[18488]_ ;
  assign \new_[18490]_  = \new_[18489]_  & \new_[18484]_ ;
  assign \new_[18493]_  = ~A201 & A169;
  assign \new_[18497]_  = A232 & ~A203;
  assign \new_[18498]_  = ~A202 & \new_[18497]_ ;
  assign \new_[18499]_  = \new_[18498]_  & \new_[18493]_ ;
  assign \new_[18502]_  = A236 & ~A233;
  assign \new_[18506]_  = A302 & A299;
  assign \new_[18507]_  = ~A298 & \new_[18506]_ ;
  assign \new_[18508]_  = \new_[18507]_  & \new_[18502]_ ;
  assign \new_[18511]_  = ~A201 & A169;
  assign \new_[18515]_  = A232 & ~A203;
  assign \new_[18516]_  = ~A202 & \new_[18515]_ ;
  assign \new_[18517]_  = \new_[18516]_  & \new_[18511]_ ;
  assign \new_[18520]_  = A236 & ~A233;
  assign \new_[18524]_  = A269 & A266;
  assign \new_[18525]_  = ~A265 & \new_[18524]_ ;
  assign \new_[18526]_  = \new_[18525]_  & \new_[18520]_ ;
  assign \new_[18529]_  = ~A201 & A169;
  assign \new_[18533]_  = A232 & ~A203;
  assign \new_[18534]_  = ~A202 & \new_[18533]_ ;
  assign \new_[18535]_  = \new_[18534]_  & \new_[18529]_ ;
  assign \new_[18538]_  = A236 & ~A233;
  assign \new_[18542]_  = A269 & ~A266;
  assign \new_[18543]_  = A265 & \new_[18542]_ ;
  assign \new_[18544]_  = \new_[18543]_  & \new_[18538]_ ;
  assign \new_[18547]_  = A199 & A169;
  assign \new_[18551]_  = ~A202 & ~A201;
  assign \new_[18552]_  = A200 & \new_[18551]_ ;
  assign \new_[18553]_  = \new_[18552]_  & \new_[18547]_ ;
  assign \new_[18556]_  = A234 & A232;
  assign \new_[18560]_  = A302 & ~A299;
  assign \new_[18561]_  = A298 & \new_[18560]_ ;
  assign \new_[18562]_  = \new_[18561]_  & \new_[18556]_ ;
  assign \new_[18565]_  = A199 & A169;
  assign \new_[18569]_  = ~A202 & ~A201;
  assign \new_[18570]_  = A200 & \new_[18569]_ ;
  assign \new_[18571]_  = \new_[18570]_  & \new_[18565]_ ;
  assign \new_[18574]_  = A234 & A232;
  assign \new_[18578]_  = A302 & A299;
  assign \new_[18579]_  = ~A298 & \new_[18578]_ ;
  assign \new_[18580]_  = \new_[18579]_  & \new_[18574]_ ;
  assign \new_[18583]_  = A199 & A169;
  assign \new_[18587]_  = ~A202 & ~A201;
  assign \new_[18588]_  = A200 & \new_[18587]_ ;
  assign \new_[18589]_  = \new_[18588]_  & \new_[18583]_ ;
  assign \new_[18592]_  = A234 & A232;
  assign \new_[18596]_  = A269 & A266;
  assign \new_[18597]_  = ~A265 & \new_[18596]_ ;
  assign \new_[18598]_  = \new_[18597]_  & \new_[18592]_ ;
  assign \new_[18601]_  = A199 & A169;
  assign \new_[18605]_  = ~A202 & ~A201;
  assign \new_[18606]_  = A200 & \new_[18605]_ ;
  assign \new_[18607]_  = \new_[18606]_  & \new_[18601]_ ;
  assign \new_[18610]_  = A234 & A232;
  assign \new_[18614]_  = A269 & ~A266;
  assign \new_[18615]_  = A265 & \new_[18614]_ ;
  assign \new_[18616]_  = \new_[18615]_  & \new_[18610]_ ;
  assign \new_[18619]_  = A199 & A169;
  assign \new_[18623]_  = ~A202 & ~A201;
  assign \new_[18624]_  = A200 & \new_[18623]_ ;
  assign \new_[18625]_  = \new_[18624]_  & \new_[18619]_ ;
  assign \new_[18628]_  = A234 & A233;
  assign \new_[18632]_  = A302 & ~A299;
  assign \new_[18633]_  = A298 & \new_[18632]_ ;
  assign \new_[18634]_  = \new_[18633]_  & \new_[18628]_ ;
  assign \new_[18637]_  = A199 & A169;
  assign \new_[18641]_  = ~A202 & ~A201;
  assign \new_[18642]_  = A200 & \new_[18641]_ ;
  assign \new_[18643]_  = \new_[18642]_  & \new_[18637]_ ;
  assign \new_[18646]_  = A234 & A233;
  assign \new_[18650]_  = A302 & A299;
  assign \new_[18651]_  = ~A298 & \new_[18650]_ ;
  assign \new_[18652]_  = \new_[18651]_  & \new_[18646]_ ;
  assign \new_[18655]_  = A199 & A169;
  assign \new_[18659]_  = ~A202 & ~A201;
  assign \new_[18660]_  = A200 & \new_[18659]_ ;
  assign \new_[18661]_  = \new_[18660]_  & \new_[18655]_ ;
  assign \new_[18664]_  = A234 & A233;
  assign \new_[18668]_  = A269 & A266;
  assign \new_[18669]_  = ~A265 & \new_[18668]_ ;
  assign \new_[18670]_  = \new_[18669]_  & \new_[18664]_ ;
  assign \new_[18673]_  = A199 & A169;
  assign \new_[18677]_  = ~A202 & ~A201;
  assign \new_[18678]_  = A200 & \new_[18677]_ ;
  assign \new_[18679]_  = \new_[18678]_  & \new_[18673]_ ;
  assign \new_[18682]_  = A234 & A233;
  assign \new_[18686]_  = A269 & ~A266;
  assign \new_[18687]_  = A265 & \new_[18686]_ ;
  assign \new_[18688]_  = \new_[18687]_  & \new_[18682]_ ;
  assign \new_[18691]_  = A199 & A169;
  assign \new_[18695]_  = ~A202 & ~A201;
  assign \new_[18696]_  = A200 & \new_[18695]_ ;
  assign \new_[18697]_  = \new_[18696]_  & \new_[18691]_ ;
  assign \new_[18700]_  = A233 & ~A232;
  assign \new_[18704]_  = A300 & A299;
  assign \new_[18705]_  = A236 & \new_[18704]_ ;
  assign \new_[18706]_  = \new_[18705]_  & \new_[18700]_ ;
  assign \new_[18709]_  = A199 & A169;
  assign \new_[18713]_  = ~A202 & ~A201;
  assign \new_[18714]_  = A200 & \new_[18713]_ ;
  assign \new_[18715]_  = \new_[18714]_  & \new_[18709]_ ;
  assign \new_[18718]_  = A233 & ~A232;
  assign \new_[18722]_  = A300 & A298;
  assign \new_[18723]_  = A236 & \new_[18722]_ ;
  assign \new_[18724]_  = \new_[18723]_  & \new_[18718]_ ;
  assign \new_[18727]_  = A199 & A169;
  assign \new_[18731]_  = ~A202 & ~A201;
  assign \new_[18732]_  = A200 & \new_[18731]_ ;
  assign \new_[18733]_  = \new_[18732]_  & \new_[18727]_ ;
  assign \new_[18736]_  = A233 & ~A232;
  assign \new_[18740]_  = A267 & A265;
  assign \new_[18741]_  = A236 & \new_[18740]_ ;
  assign \new_[18742]_  = \new_[18741]_  & \new_[18736]_ ;
  assign \new_[18745]_  = A199 & A169;
  assign \new_[18749]_  = ~A202 & ~A201;
  assign \new_[18750]_  = A200 & \new_[18749]_ ;
  assign \new_[18751]_  = \new_[18750]_  & \new_[18745]_ ;
  assign \new_[18754]_  = A233 & ~A232;
  assign \new_[18758]_  = A267 & A266;
  assign \new_[18759]_  = A236 & \new_[18758]_ ;
  assign \new_[18760]_  = \new_[18759]_  & \new_[18754]_ ;
  assign \new_[18763]_  = A199 & A169;
  assign \new_[18767]_  = ~A202 & ~A201;
  assign \new_[18768]_  = A200 & \new_[18767]_ ;
  assign \new_[18769]_  = \new_[18768]_  & \new_[18763]_ ;
  assign \new_[18772]_  = ~A233 & A232;
  assign \new_[18776]_  = A300 & A299;
  assign \new_[18777]_  = A236 & \new_[18776]_ ;
  assign \new_[18778]_  = \new_[18777]_  & \new_[18772]_ ;
  assign \new_[18781]_  = A199 & A169;
  assign \new_[18785]_  = ~A202 & ~A201;
  assign \new_[18786]_  = A200 & \new_[18785]_ ;
  assign \new_[18787]_  = \new_[18786]_  & \new_[18781]_ ;
  assign \new_[18790]_  = ~A233 & A232;
  assign \new_[18794]_  = A300 & A298;
  assign \new_[18795]_  = A236 & \new_[18794]_ ;
  assign \new_[18796]_  = \new_[18795]_  & \new_[18790]_ ;
  assign \new_[18799]_  = A199 & A169;
  assign \new_[18803]_  = ~A202 & ~A201;
  assign \new_[18804]_  = A200 & \new_[18803]_ ;
  assign \new_[18805]_  = \new_[18804]_  & \new_[18799]_ ;
  assign \new_[18808]_  = ~A233 & A232;
  assign \new_[18812]_  = A267 & A265;
  assign \new_[18813]_  = A236 & \new_[18812]_ ;
  assign \new_[18814]_  = \new_[18813]_  & \new_[18808]_ ;
  assign \new_[18817]_  = A199 & A169;
  assign \new_[18821]_  = ~A202 & ~A201;
  assign \new_[18822]_  = A200 & \new_[18821]_ ;
  assign \new_[18823]_  = \new_[18822]_  & \new_[18817]_ ;
  assign \new_[18826]_  = ~A233 & A232;
  assign \new_[18830]_  = A267 & A266;
  assign \new_[18831]_  = A236 & \new_[18830]_ ;
  assign \new_[18832]_  = \new_[18831]_  & \new_[18826]_ ;
  assign \new_[18835]_  = ~A199 & A169;
  assign \new_[18839]_  = ~A232 & ~A202;
  assign \new_[18840]_  = ~A200 & \new_[18839]_ ;
  assign \new_[18841]_  = \new_[18840]_  & \new_[18835]_ ;
  assign \new_[18844]_  = A236 & A233;
  assign \new_[18848]_  = A302 & ~A299;
  assign \new_[18849]_  = A298 & \new_[18848]_ ;
  assign \new_[18850]_  = \new_[18849]_  & \new_[18844]_ ;
  assign \new_[18853]_  = ~A199 & A169;
  assign \new_[18857]_  = ~A232 & ~A202;
  assign \new_[18858]_  = ~A200 & \new_[18857]_ ;
  assign \new_[18859]_  = \new_[18858]_  & \new_[18853]_ ;
  assign \new_[18862]_  = A236 & A233;
  assign \new_[18866]_  = A302 & A299;
  assign \new_[18867]_  = ~A298 & \new_[18866]_ ;
  assign \new_[18868]_  = \new_[18867]_  & \new_[18862]_ ;
  assign \new_[18871]_  = ~A199 & A169;
  assign \new_[18875]_  = ~A232 & ~A202;
  assign \new_[18876]_  = ~A200 & \new_[18875]_ ;
  assign \new_[18877]_  = \new_[18876]_  & \new_[18871]_ ;
  assign \new_[18880]_  = A236 & A233;
  assign \new_[18884]_  = A269 & A266;
  assign \new_[18885]_  = ~A265 & \new_[18884]_ ;
  assign \new_[18886]_  = \new_[18885]_  & \new_[18880]_ ;
  assign \new_[18889]_  = ~A199 & A169;
  assign \new_[18893]_  = ~A232 & ~A202;
  assign \new_[18894]_  = ~A200 & \new_[18893]_ ;
  assign \new_[18895]_  = \new_[18894]_  & \new_[18889]_ ;
  assign \new_[18898]_  = A236 & A233;
  assign \new_[18902]_  = A269 & ~A266;
  assign \new_[18903]_  = A265 & \new_[18902]_ ;
  assign \new_[18904]_  = \new_[18903]_  & \new_[18898]_ ;
  assign \new_[18907]_  = ~A199 & A169;
  assign \new_[18911]_  = A232 & ~A202;
  assign \new_[18912]_  = ~A200 & \new_[18911]_ ;
  assign \new_[18913]_  = \new_[18912]_  & \new_[18907]_ ;
  assign \new_[18916]_  = A236 & ~A233;
  assign \new_[18920]_  = A302 & ~A299;
  assign \new_[18921]_  = A298 & \new_[18920]_ ;
  assign \new_[18922]_  = \new_[18921]_  & \new_[18916]_ ;
  assign \new_[18925]_  = ~A199 & A169;
  assign \new_[18929]_  = A232 & ~A202;
  assign \new_[18930]_  = ~A200 & \new_[18929]_ ;
  assign \new_[18931]_  = \new_[18930]_  & \new_[18925]_ ;
  assign \new_[18934]_  = A236 & ~A233;
  assign \new_[18938]_  = A302 & A299;
  assign \new_[18939]_  = ~A298 & \new_[18938]_ ;
  assign \new_[18940]_  = \new_[18939]_  & \new_[18934]_ ;
  assign \new_[18943]_  = ~A199 & A169;
  assign \new_[18947]_  = A232 & ~A202;
  assign \new_[18948]_  = ~A200 & \new_[18947]_ ;
  assign \new_[18949]_  = \new_[18948]_  & \new_[18943]_ ;
  assign \new_[18952]_  = A236 & ~A233;
  assign \new_[18956]_  = A269 & A266;
  assign \new_[18957]_  = ~A265 & \new_[18956]_ ;
  assign \new_[18958]_  = \new_[18957]_  & \new_[18952]_ ;
  assign \new_[18961]_  = ~A199 & A169;
  assign \new_[18965]_  = A232 & ~A202;
  assign \new_[18966]_  = ~A200 & \new_[18965]_ ;
  assign \new_[18967]_  = \new_[18966]_  & \new_[18961]_ ;
  assign \new_[18970]_  = A236 & ~A233;
  assign \new_[18974]_  = A269 & ~A266;
  assign \new_[18975]_  = A265 & \new_[18974]_ ;
  assign \new_[18976]_  = \new_[18975]_  & \new_[18970]_ ;
  assign \new_[18979]_  = ~A167 & ~A169;
  assign \new_[18983]_  = ~A232 & A202;
  assign \new_[18984]_  = ~A166 & \new_[18983]_ ;
  assign \new_[18985]_  = \new_[18984]_  & \new_[18979]_ ;
  assign \new_[18988]_  = A236 & A233;
  assign \new_[18992]_  = A302 & ~A299;
  assign \new_[18993]_  = A298 & \new_[18992]_ ;
  assign \new_[18994]_  = \new_[18993]_  & \new_[18988]_ ;
  assign \new_[18997]_  = ~A167 & ~A169;
  assign \new_[19001]_  = ~A232 & A202;
  assign \new_[19002]_  = ~A166 & \new_[19001]_ ;
  assign \new_[19003]_  = \new_[19002]_  & \new_[18997]_ ;
  assign \new_[19006]_  = A236 & A233;
  assign \new_[19010]_  = A302 & A299;
  assign \new_[19011]_  = ~A298 & \new_[19010]_ ;
  assign \new_[19012]_  = \new_[19011]_  & \new_[19006]_ ;
  assign \new_[19015]_  = ~A167 & ~A169;
  assign \new_[19019]_  = ~A232 & A202;
  assign \new_[19020]_  = ~A166 & \new_[19019]_ ;
  assign \new_[19021]_  = \new_[19020]_  & \new_[19015]_ ;
  assign \new_[19024]_  = A236 & A233;
  assign \new_[19028]_  = A269 & A266;
  assign \new_[19029]_  = ~A265 & \new_[19028]_ ;
  assign \new_[19030]_  = \new_[19029]_  & \new_[19024]_ ;
  assign \new_[19033]_  = ~A167 & ~A169;
  assign \new_[19037]_  = ~A232 & A202;
  assign \new_[19038]_  = ~A166 & \new_[19037]_ ;
  assign \new_[19039]_  = \new_[19038]_  & \new_[19033]_ ;
  assign \new_[19042]_  = A236 & A233;
  assign \new_[19046]_  = A269 & ~A266;
  assign \new_[19047]_  = A265 & \new_[19046]_ ;
  assign \new_[19048]_  = \new_[19047]_  & \new_[19042]_ ;
  assign \new_[19051]_  = ~A167 & ~A169;
  assign \new_[19055]_  = A232 & A202;
  assign \new_[19056]_  = ~A166 & \new_[19055]_ ;
  assign \new_[19057]_  = \new_[19056]_  & \new_[19051]_ ;
  assign \new_[19060]_  = A236 & ~A233;
  assign \new_[19064]_  = A302 & ~A299;
  assign \new_[19065]_  = A298 & \new_[19064]_ ;
  assign \new_[19066]_  = \new_[19065]_  & \new_[19060]_ ;
  assign \new_[19069]_  = ~A167 & ~A169;
  assign \new_[19073]_  = A232 & A202;
  assign \new_[19074]_  = ~A166 & \new_[19073]_ ;
  assign \new_[19075]_  = \new_[19074]_  & \new_[19069]_ ;
  assign \new_[19078]_  = A236 & ~A233;
  assign \new_[19082]_  = A302 & A299;
  assign \new_[19083]_  = ~A298 & \new_[19082]_ ;
  assign \new_[19084]_  = \new_[19083]_  & \new_[19078]_ ;
  assign \new_[19087]_  = ~A167 & ~A169;
  assign \new_[19091]_  = A232 & A202;
  assign \new_[19092]_  = ~A166 & \new_[19091]_ ;
  assign \new_[19093]_  = \new_[19092]_  & \new_[19087]_ ;
  assign \new_[19096]_  = A236 & ~A233;
  assign \new_[19100]_  = A269 & A266;
  assign \new_[19101]_  = ~A265 & \new_[19100]_ ;
  assign \new_[19102]_  = \new_[19101]_  & \new_[19096]_ ;
  assign \new_[19105]_  = ~A167 & ~A169;
  assign \new_[19109]_  = A232 & A202;
  assign \new_[19110]_  = ~A166 & \new_[19109]_ ;
  assign \new_[19111]_  = \new_[19110]_  & \new_[19105]_ ;
  assign \new_[19114]_  = A236 & ~A233;
  assign \new_[19118]_  = A269 & ~A266;
  assign \new_[19119]_  = A265 & \new_[19118]_ ;
  assign \new_[19120]_  = \new_[19119]_  & \new_[19114]_ ;
  assign \new_[19123]_  = ~A167 & ~A169;
  assign \new_[19127]_  = A201 & A199;
  assign \new_[19128]_  = ~A166 & \new_[19127]_ ;
  assign \new_[19129]_  = \new_[19128]_  & \new_[19123]_ ;
  assign \new_[19132]_  = A234 & A232;
  assign \new_[19136]_  = A302 & ~A299;
  assign \new_[19137]_  = A298 & \new_[19136]_ ;
  assign \new_[19138]_  = \new_[19137]_  & \new_[19132]_ ;
  assign \new_[19141]_  = ~A167 & ~A169;
  assign \new_[19145]_  = A201 & A199;
  assign \new_[19146]_  = ~A166 & \new_[19145]_ ;
  assign \new_[19147]_  = \new_[19146]_  & \new_[19141]_ ;
  assign \new_[19150]_  = A234 & A232;
  assign \new_[19154]_  = A302 & A299;
  assign \new_[19155]_  = ~A298 & \new_[19154]_ ;
  assign \new_[19156]_  = \new_[19155]_  & \new_[19150]_ ;
  assign \new_[19159]_  = ~A167 & ~A169;
  assign \new_[19163]_  = A201 & A199;
  assign \new_[19164]_  = ~A166 & \new_[19163]_ ;
  assign \new_[19165]_  = \new_[19164]_  & \new_[19159]_ ;
  assign \new_[19168]_  = A234 & A232;
  assign \new_[19172]_  = A269 & A266;
  assign \new_[19173]_  = ~A265 & \new_[19172]_ ;
  assign \new_[19174]_  = \new_[19173]_  & \new_[19168]_ ;
  assign \new_[19177]_  = ~A167 & ~A169;
  assign \new_[19181]_  = A201 & A199;
  assign \new_[19182]_  = ~A166 & \new_[19181]_ ;
  assign \new_[19183]_  = \new_[19182]_  & \new_[19177]_ ;
  assign \new_[19186]_  = A234 & A232;
  assign \new_[19190]_  = A269 & ~A266;
  assign \new_[19191]_  = A265 & \new_[19190]_ ;
  assign \new_[19192]_  = \new_[19191]_  & \new_[19186]_ ;
  assign \new_[19195]_  = ~A167 & ~A169;
  assign \new_[19199]_  = A201 & A199;
  assign \new_[19200]_  = ~A166 & \new_[19199]_ ;
  assign \new_[19201]_  = \new_[19200]_  & \new_[19195]_ ;
  assign \new_[19204]_  = A234 & A233;
  assign \new_[19208]_  = A302 & ~A299;
  assign \new_[19209]_  = A298 & \new_[19208]_ ;
  assign \new_[19210]_  = \new_[19209]_  & \new_[19204]_ ;
  assign \new_[19213]_  = ~A167 & ~A169;
  assign \new_[19217]_  = A201 & A199;
  assign \new_[19218]_  = ~A166 & \new_[19217]_ ;
  assign \new_[19219]_  = \new_[19218]_  & \new_[19213]_ ;
  assign \new_[19222]_  = A234 & A233;
  assign \new_[19226]_  = A302 & A299;
  assign \new_[19227]_  = ~A298 & \new_[19226]_ ;
  assign \new_[19228]_  = \new_[19227]_  & \new_[19222]_ ;
  assign \new_[19231]_  = ~A167 & ~A169;
  assign \new_[19235]_  = A201 & A199;
  assign \new_[19236]_  = ~A166 & \new_[19235]_ ;
  assign \new_[19237]_  = \new_[19236]_  & \new_[19231]_ ;
  assign \new_[19240]_  = A234 & A233;
  assign \new_[19244]_  = A269 & A266;
  assign \new_[19245]_  = ~A265 & \new_[19244]_ ;
  assign \new_[19246]_  = \new_[19245]_  & \new_[19240]_ ;
  assign \new_[19249]_  = ~A167 & ~A169;
  assign \new_[19253]_  = A201 & A199;
  assign \new_[19254]_  = ~A166 & \new_[19253]_ ;
  assign \new_[19255]_  = \new_[19254]_  & \new_[19249]_ ;
  assign \new_[19258]_  = A234 & A233;
  assign \new_[19262]_  = A269 & ~A266;
  assign \new_[19263]_  = A265 & \new_[19262]_ ;
  assign \new_[19264]_  = \new_[19263]_  & \new_[19258]_ ;
  assign \new_[19267]_  = ~A167 & ~A169;
  assign \new_[19271]_  = A201 & A199;
  assign \new_[19272]_  = ~A166 & \new_[19271]_ ;
  assign \new_[19273]_  = \new_[19272]_  & \new_[19267]_ ;
  assign \new_[19276]_  = A233 & ~A232;
  assign \new_[19280]_  = A300 & A299;
  assign \new_[19281]_  = A236 & \new_[19280]_ ;
  assign \new_[19282]_  = \new_[19281]_  & \new_[19276]_ ;
  assign \new_[19285]_  = ~A167 & ~A169;
  assign \new_[19289]_  = A201 & A199;
  assign \new_[19290]_  = ~A166 & \new_[19289]_ ;
  assign \new_[19291]_  = \new_[19290]_  & \new_[19285]_ ;
  assign \new_[19294]_  = A233 & ~A232;
  assign \new_[19298]_  = A300 & A298;
  assign \new_[19299]_  = A236 & \new_[19298]_ ;
  assign \new_[19300]_  = \new_[19299]_  & \new_[19294]_ ;
  assign \new_[19303]_  = ~A167 & ~A169;
  assign \new_[19307]_  = A201 & A199;
  assign \new_[19308]_  = ~A166 & \new_[19307]_ ;
  assign \new_[19309]_  = \new_[19308]_  & \new_[19303]_ ;
  assign \new_[19312]_  = A233 & ~A232;
  assign \new_[19316]_  = A267 & A265;
  assign \new_[19317]_  = A236 & \new_[19316]_ ;
  assign \new_[19318]_  = \new_[19317]_  & \new_[19312]_ ;
  assign \new_[19321]_  = ~A167 & ~A169;
  assign \new_[19325]_  = A201 & A199;
  assign \new_[19326]_  = ~A166 & \new_[19325]_ ;
  assign \new_[19327]_  = \new_[19326]_  & \new_[19321]_ ;
  assign \new_[19330]_  = A233 & ~A232;
  assign \new_[19334]_  = A267 & A266;
  assign \new_[19335]_  = A236 & \new_[19334]_ ;
  assign \new_[19336]_  = \new_[19335]_  & \new_[19330]_ ;
  assign \new_[19339]_  = ~A167 & ~A169;
  assign \new_[19343]_  = A201 & A199;
  assign \new_[19344]_  = ~A166 & \new_[19343]_ ;
  assign \new_[19345]_  = \new_[19344]_  & \new_[19339]_ ;
  assign \new_[19348]_  = ~A233 & A232;
  assign \new_[19352]_  = A300 & A299;
  assign \new_[19353]_  = A236 & \new_[19352]_ ;
  assign \new_[19354]_  = \new_[19353]_  & \new_[19348]_ ;
  assign \new_[19357]_  = ~A167 & ~A169;
  assign \new_[19361]_  = A201 & A199;
  assign \new_[19362]_  = ~A166 & \new_[19361]_ ;
  assign \new_[19363]_  = \new_[19362]_  & \new_[19357]_ ;
  assign \new_[19366]_  = ~A233 & A232;
  assign \new_[19370]_  = A300 & A298;
  assign \new_[19371]_  = A236 & \new_[19370]_ ;
  assign \new_[19372]_  = \new_[19371]_  & \new_[19366]_ ;
  assign \new_[19375]_  = ~A167 & ~A169;
  assign \new_[19379]_  = A201 & A199;
  assign \new_[19380]_  = ~A166 & \new_[19379]_ ;
  assign \new_[19381]_  = \new_[19380]_  & \new_[19375]_ ;
  assign \new_[19384]_  = ~A233 & A232;
  assign \new_[19388]_  = A267 & A265;
  assign \new_[19389]_  = A236 & \new_[19388]_ ;
  assign \new_[19390]_  = \new_[19389]_  & \new_[19384]_ ;
  assign \new_[19393]_  = ~A167 & ~A169;
  assign \new_[19397]_  = A201 & A199;
  assign \new_[19398]_  = ~A166 & \new_[19397]_ ;
  assign \new_[19399]_  = \new_[19398]_  & \new_[19393]_ ;
  assign \new_[19402]_  = ~A233 & A232;
  assign \new_[19406]_  = A267 & A266;
  assign \new_[19407]_  = A236 & \new_[19406]_ ;
  assign \new_[19408]_  = \new_[19407]_  & \new_[19402]_ ;
  assign \new_[19411]_  = ~A167 & ~A169;
  assign \new_[19415]_  = A201 & A200;
  assign \new_[19416]_  = ~A166 & \new_[19415]_ ;
  assign \new_[19417]_  = \new_[19416]_  & \new_[19411]_ ;
  assign \new_[19420]_  = A234 & A232;
  assign \new_[19424]_  = A302 & ~A299;
  assign \new_[19425]_  = A298 & \new_[19424]_ ;
  assign \new_[19426]_  = \new_[19425]_  & \new_[19420]_ ;
  assign \new_[19429]_  = ~A167 & ~A169;
  assign \new_[19433]_  = A201 & A200;
  assign \new_[19434]_  = ~A166 & \new_[19433]_ ;
  assign \new_[19435]_  = \new_[19434]_  & \new_[19429]_ ;
  assign \new_[19438]_  = A234 & A232;
  assign \new_[19442]_  = A302 & A299;
  assign \new_[19443]_  = ~A298 & \new_[19442]_ ;
  assign \new_[19444]_  = \new_[19443]_  & \new_[19438]_ ;
  assign \new_[19447]_  = ~A167 & ~A169;
  assign \new_[19451]_  = A201 & A200;
  assign \new_[19452]_  = ~A166 & \new_[19451]_ ;
  assign \new_[19453]_  = \new_[19452]_  & \new_[19447]_ ;
  assign \new_[19456]_  = A234 & A232;
  assign \new_[19460]_  = A269 & A266;
  assign \new_[19461]_  = ~A265 & \new_[19460]_ ;
  assign \new_[19462]_  = \new_[19461]_  & \new_[19456]_ ;
  assign \new_[19465]_  = ~A167 & ~A169;
  assign \new_[19469]_  = A201 & A200;
  assign \new_[19470]_  = ~A166 & \new_[19469]_ ;
  assign \new_[19471]_  = \new_[19470]_  & \new_[19465]_ ;
  assign \new_[19474]_  = A234 & A232;
  assign \new_[19478]_  = A269 & ~A266;
  assign \new_[19479]_  = A265 & \new_[19478]_ ;
  assign \new_[19480]_  = \new_[19479]_  & \new_[19474]_ ;
  assign \new_[19483]_  = ~A167 & ~A169;
  assign \new_[19487]_  = A201 & A200;
  assign \new_[19488]_  = ~A166 & \new_[19487]_ ;
  assign \new_[19489]_  = \new_[19488]_  & \new_[19483]_ ;
  assign \new_[19492]_  = A234 & A233;
  assign \new_[19496]_  = A302 & ~A299;
  assign \new_[19497]_  = A298 & \new_[19496]_ ;
  assign \new_[19498]_  = \new_[19497]_  & \new_[19492]_ ;
  assign \new_[19501]_  = ~A167 & ~A169;
  assign \new_[19505]_  = A201 & A200;
  assign \new_[19506]_  = ~A166 & \new_[19505]_ ;
  assign \new_[19507]_  = \new_[19506]_  & \new_[19501]_ ;
  assign \new_[19510]_  = A234 & A233;
  assign \new_[19514]_  = A302 & A299;
  assign \new_[19515]_  = ~A298 & \new_[19514]_ ;
  assign \new_[19516]_  = \new_[19515]_  & \new_[19510]_ ;
  assign \new_[19519]_  = ~A167 & ~A169;
  assign \new_[19523]_  = A201 & A200;
  assign \new_[19524]_  = ~A166 & \new_[19523]_ ;
  assign \new_[19525]_  = \new_[19524]_  & \new_[19519]_ ;
  assign \new_[19528]_  = A234 & A233;
  assign \new_[19532]_  = A269 & A266;
  assign \new_[19533]_  = ~A265 & \new_[19532]_ ;
  assign \new_[19534]_  = \new_[19533]_  & \new_[19528]_ ;
  assign \new_[19537]_  = ~A167 & ~A169;
  assign \new_[19541]_  = A201 & A200;
  assign \new_[19542]_  = ~A166 & \new_[19541]_ ;
  assign \new_[19543]_  = \new_[19542]_  & \new_[19537]_ ;
  assign \new_[19546]_  = A234 & A233;
  assign \new_[19550]_  = A269 & ~A266;
  assign \new_[19551]_  = A265 & \new_[19550]_ ;
  assign \new_[19552]_  = \new_[19551]_  & \new_[19546]_ ;
  assign \new_[19555]_  = ~A167 & ~A169;
  assign \new_[19559]_  = A201 & A200;
  assign \new_[19560]_  = ~A166 & \new_[19559]_ ;
  assign \new_[19561]_  = \new_[19560]_  & \new_[19555]_ ;
  assign \new_[19564]_  = A233 & ~A232;
  assign \new_[19568]_  = A300 & A299;
  assign \new_[19569]_  = A236 & \new_[19568]_ ;
  assign \new_[19570]_  = \new_[19569]_  & \new_[19564]_ ;
  assign \new_[19573]_  = ~A167 & ~A169;
  assign \new_[19577]_  = A201 & A200;
  assign \new_[19578]_  = ~A166 & \new_[19577]_ ;
  assign \new_[19579]_  = \new_[19578]_  & \new_[19573]_ ;
  assign \new_[19582]_  = A233 & ~A232;
  assign \new_[19586]_  = A300 & A298;
  assign \new_[19587]_  = A236 & \new_[19586]_ ;
  assign \new_[19588]_  = \new_[19587]_  & \new_[19582]_ ;
  assign \new_[19591]_  = ~A167 & ~A169;
  assign \new_[19595]_  = A201 & A200;
  assign \new_[19596]_  = ~A166 & \new_[19595]_ ;
  assign \new_[19597]_  = \new_[19596]_  & \new_[19591]_ ;
  assign \new_[19600]_  = A233 & ~A232;
  assign \new_[19604]_  = A267 & A265;
  assign \new_[19605]_  = A236 & \new_[19604]_ ;
  assign \new_[19606]_  = \new_[19605]_  & \new_[19600]_ ;
  assign \new_[19609]_  = ~A167 & ~A169;
  assign \new_[19613]_  = A201 & A200;
  assign \new_[19614]_  = ~A166 & \new_[19613]_ ;
  assign \new_[19615]_  = \new_[19614]_  & \new_[19609]_ ;
  assign \new_[19618]_  = A233 & ~A232;
  assign \new_[19622]_  = A267 & A266;
  assign \new_[19623]_  = A236 & \new_[19622]_ ;
  assign \new_[19624]_  = \new_[19623]_  & \new_[19618]_ ;
  assign \new_[19627]_  = ~A167 & ~A169;
  assign \new_[19631]_  = A201 & A200;
  assign \new_[19632]_  = ~A166 & \new_[19631]_ ;
  assign \new_[19633]_  = \new_[19632]_  & \new_[19627]_ ;
  assign \new_[19636]_  = ~A233 & A232;
  assign \new_[19640]_  = A300 & A299;
  assign \new_[19641]_  = A236 & \new_[19640]_ ;
  assign \new_[19642]_  = \new_[19641]_  & \new_[19636]_ ;
  assign \new_[19645]_  = ~A167 & ~A169;
  assign \new_[19649]_  = A201 & A200;
  assign \new_[19650]_  = ~A166 & \new_[19649]_ ;
  assign \new_[19651]_  = \new_[19650]_  & \new_[19645]_ ;
  assign \new_[19654]_  = ~A233 & A232;
  assign \new_[19658]_  = A300 & A298;
  assign \new_[19659]_  = A236 & \new_[19658]_ ;
  assign \new_[19660]_  = \new_[19659]_  & \new_[19654]_ ;
  assign \new_[19663]_  = ~A167 & ~A169;
  assign \new_[19667]_  = A201 & A200;
  assign \new_[19668]_  = ~A166 & \new_[19667]_ ;
  assign \new_[19669]_  = \new_[19668]_  & \new_[19663]_ ;
  assign \new_[19672]_  = ~A233 & A232;
  assign \new_[19676]_  = A267 & A265;
  assign \new_[19677]_  = A236 & \new_[19676]_ ;
  assign \new_[19678]_  = \new_[19677]_  & \new_[19672]_ ;
  assign \new_[19681]_  = ~A167 & ~A169;
  assign \new_[19685]_  = A201 & A200;
  assign \new_[19686]_  = ~A166 & \new_[19685]_ ;
  assign \new_[19687]_  = \new_[19686]_  & \new_[19681]_ ;
  assign \new_[19690]_  = ~A233 & A232;
  assign \new_[19694]_  = A267 & A266;
  assign \new_[19695]_  = A236 & \new_[19694]_ ;
  assign \new_[19696]_  = \new_[19695]_  & \new_[19690]_ ;
  assign \new_[19699]_  = ~A167 & ~A169;
  assign \new_[19703]_  = A200 & ~A199;
  assign \new_[19704]_  = ~A166 & \new_[19703]_ ;
  assign \new_[19705]_  = \new_[19704]_  & \new_[19699]_ ;
  assign \new_[19708]_  = A235 & A203;
  assign \new_[19712]_  = A302 & ~A299;
  assign \new_[19713]_  = A298 & \new_[19712]_ ;
  assign \new_[19714]_  = \new_[19713]_  & \new_[19708]_ ;
  assign \new_[19717]_  = ~A167 & ~A169;
  assign \new_[19721]_  = A200 & ~A199;
  assign \new_[19722]_  = ~A166 & \new_[19721]_ ;
  assign \new_[19723]_  = \new_[19722]_  & \new_[19717]_ ;
  assign \new_[19726]_  = A235 & A203;
  assign \new_[19730]_  = A302 & A299;
  assign \new_[19731]_  = ~A298 & \new_[19730]_ ;
  assign \new_[19732]_  = \new_[19731]_  & \new_[19726]_ ;
  assign \new_[19735]_  = ~A167 & ~A169;
  assign \new_[19739]_  = A200 & ~A199;
  assign \new_[19740]_  = ~A166 & \new_[19739]_ ;
  assign \new_[19741]_  = \new_[19740]_  & \new_[19735]_ ;
  assign \new_[19744]_  = A235 & A203;
  assign \new_[19748]_  = A269 & A266;
  assign \new_[19749]_  = ~A265 & \new_[19748]_ ;
  assign \new_[19750]_  = \new_[19749]_  & \new_[19744]_ ;
  assign \new_[19753]_  = ~A167 & ~A169;
  assign \new_[19757]_  = A200 & ~A199;
  assign \new_[19758]_  = ~A166 & \new_[19757]_ ;
  assign \new_[19759]_  = \new_[19758]_  & \new_[19753]_ ;
  assign \new_[19762]_  = A235 & A203;
  assign \new_[19766]_  = A269 & ~A266;
  assign \new_[19767]_  = A265 & \new_[19766]_ ;
  assign \new_[19768]_  = \new_[19767]_  & \new_[19762]_ ;
  assign \new_[19771]_  = ~A167 & ~A169;
  assign \new_[19775]_  = A200 & ~A199;
  assign \new_[19776]_  = ~A166 & \new_[19775]_ ;
  assign \new_[19777]_  = \new_[19776]_  & \new_[19771]_ ;
  assign \new_[19780]_  = A232 & A203;
  assign \new_[19784]_  = A300 & A299;
  assign \new_[19785]_  = A234 & \new_[19784]_ ;
  assign \new_[19786]_  = \new_[19785]_  & \new_[19780]_ ;
  assign \new_[19789]_  = ~A167 & ~A169;
  assign \new_[19793]_  = A200 & ~A199;
  assign \new_[19794]_  = ~A166 & \new_[19793]_ ;
  assign \new_[19795]_  = \new_[19794]_  & \new_[19789]_ ;
  assign \new_[19798]_  = A232 & A203;
  assign \new_[19802]_  = A300 & A298;
  assign \new_[19803]_  = A234 & \new_[19802]_ ;
  assign \new_[19804]_  = \new_[19803]_  & \new_[19798]_ ;
  assign \new_[19807]_  = ~A167 & ~A169;
  assign \new_[19811]_  = A200 & ~A199;
  assign \new_[19812]_  = ~A166 & \new_[19811]_ ;
  assign \new_[19813]_  = \new_[19812]_  & \new_[19807]_ ;
  assign \new_[19816]_  = A232 & A203;
  assign \new_[19820]_  = A267 & A265;
  assign \new_[19821]_  = A234 & \new_[19820]_ ;
  assign \new_[19822]_  = \new_[19821]_  & \new_[19816]_ ;
  assign \new_[19825]_  = ~A167 & ~A169;
  assign \new_[19829]_  = A200 & ~A199;
  assign \new_[19830]_  = ~A166 & \new_[19829]_ ;
  assign \new_[19831]_  = \new_[19830]_  & \new_[19825]_ ;
  assign \new_[19834]_  = A232 & A203;
  assign \new_[19838]_  = A267 & A266;
  assign \new_[19839]_  = A234 & \new_[19838]_ ;
  assign \new_[19840]_  = \new_[19839]_  & \new_[19834]_ ;
  assign \new_[19843]_  = ~A167 & ~A169;
  assign \new_[19847]_  = A200 & ~A199;
  assign \new_[19848]_  = ~A166 & \new_[19847]_ ;
  assign \new_[19849]_  = \new_[19848]_  & \new_[19843]_ ;
  assign \new_[19852]_  = A233 & A203;
  assign \new_[19856]_  = A300 & A299;
  assign \new_[19857]_  = A234 & \new_[19856]_ ;
  assign \new_[19858]_  = \new_[19857]_  & \new_[19852]_ ;
  assign \new_[19861]_  = ~A167 & ~A169;
  assign \new_[19865]_  = A200 & ~A199;
  assign \new_[19866]_  = ~A166 & \new_[19865]_ ;
  assign \new_[19867]_  = \new_[19866]_  & \new_[19861]_ ;
  assign \new_[19870]_  = A233 & A203;
  assign \new_[19874]_  = A300 & A298;
  assign \new_[19875]_  = A234 & \new_[19874]_ ;
  assign \new_[19876]_  = \new_[19875]_  & \new_[19870]_ ;
  assign \new_[19879]_  = ~A167 & ~A169;
  assign \new_[19883]_  = A200 & ~A199;
  assign \new_[19884]_  = ~A166 & \new_[19883]_ ;
  assign \new_[19885]_  = \new_[19884]_  & \new_[19879]_ ;
  assign \new_[19888]_  = A233 & A203;
  assign \new_[19892]_  = A267 & A265;
  assign \new_[19893]_  = A234 & \new_[19892]_ ;
  assign \new_[19894]_  = \new_[19893]_  & \new_[19888]_ ;
  assign \new_[19897]_  = ~A167 & ~A169;
  assign \new_[19901]_  = A200 & ~A199;
  assign \new_[19902]_  = ~A166 & \new_[19901]_ ;
  assign \new_[19903]_  = \new_[19902]_  & \new_[19897]_ ;
  assign \new_[19906]_  = A233 & A203;
  assign \new_[19910]_  = A267 & A266;
  assign \new_[19911]_  = A234 & \new_[19910]_ ;
  assign \new_[19912]_  = \new_[19911]_  & \new_[19906]_ ;
  assign \new_[19915]_  = ~A167 & ~A169;
  assign \new_[19919]_  = A200 & ~A199;
  assign \new_[19920]_  = ~A166 & \new_[19919]_ ;
  assign \new_[19921]_  = \new_[19920]_  & \new_[19915]_ ;
  assign \new_[19924]_  = ~A232 & A203;
  assign \new_[19928]_  = A301 & A236;
  assign \new_[19929]_  = A233 & \new_[19928]_ ;
  assign \new_[19930]_  = \new_[19929]_  & \new_[19924]_ ;
  assign \new_[19933]_  = ~A167 & ~A169;
  assign \new_[19937]_  = A200 & ~A199;
  assign \new_[19938]_  = ~A166 & \new_[19937]_ ;
  assign \new_[19939]_  = \new_[19938]_  & \new_[19933]_ ;
  assign \new_[19942]_  = ~A232 & A203;
  assign \new_[19946]_  = A268 & A236;
  assign \new_[19947]_  = A233 & \new_[19946]_ ;
  assign \new_[19948]_  = \new_[19947]_  & \new_[19942]_ ;
  assign \new_[19951]_  = ~A167 & ~A169;
  assign \new_[19955]_  = A200 & ~A199;
  assign \new_[19956]_  = ~A166 & \new_[19955]_ ;
  assign \new_[19957]_  = \new_[19956]_  & \new_[19951]_ ;
  assign \new_[19960]_  = A232 & A203;
  assign \new_[19964]_  = A301 & A236;
  assign \new_[19965]_  = ~A233 & \new_[19964]_ ;
  assign \new_[19966]_  = \new_[19965]_  & \new_[19960]_ ;
  assign \new_[19969]_  = ~A167 & ~A169;
  assign \new_[19973]_  = A200 & ~A199;
  assign \new_[19974]_  = ~A166 & \new_[19973]_ ;
  assign \new_[19975]_  = \new_[19974]_  & \new_[19969]_ ;
  assign \new_[19978]_  = A232 & A203;
  assign \new_[19982]_  = A268 & A236;
  assign \new_[19983]_  = ~A233 & \new_[19982]_ ;
  assign \new_[19984]_  = \new_[19983]_  & \new_[19978]_ ;
  assign \new_[19987]_  = ~A167 & ~A169;
  assign \new_[19991]_  = ~A200 & A199;
  assign \new_[19992]_  = ~A166 & \new_[19991]_ ;
  assign \new_[19993]_  = \new_[19992]_  & \new_[19987]_ ;
  assign \new_[19996]_  = A235 & A203;
  assign \new_[20000]_  = A302 & ~A299;
  assign \new_[20001]_  = A298 & \new_[20000]_ ;
  assign \new_[20002]_  = \new_[20001]_  & \new_[19996]_ ;
  assign \new_[20005]_  = ~A167 & ~A169;
  assign \new_[20009]_  = ~A200 & A199;
  assign \new_[20010]_  = ~A166 & \new_[20009]_ ;
  assign \new_[20011]_  = \new_[20010]_  & \new_[20005]_ ;
  assign \new_[20014]_  = A235 & A203;
  assign \new_[20018]_  = A302 & A299;
  assign \new_[20019]_  = ~A298 & \new_[20018]_ ;
  assign \new_[20020]_  = \new_[20019]_  & \new_[20014]_ ;
  assign \new_[20023]_  = ~A167 & ~A169;
  assign \new_[20027]_  = ~A200 & A199;
  assign \new_[20028]_  = ~A166 & \new_[20027]_ ;
  assign \new_[20029]_  = \new_[20028]_  & \new_[20023]_ ;
  assign \new_[20032]_  = A235 & A203;
  assign \new_[20036]_  = A269 & A266;
  assign \new_[20037]_  = ~A265 & \new_[20036]_ ;
  assign \new_[20038]_  = \new_[20037]_  & \new_[20032]_ ;
  assign \new_[20041]_  = ~A167 & ~A169;
  assign \new_[20045]_  = ~A200 & A199;
  assign \new_[20046]_  = ~A166 & \new_[20045]_ ;
  assign \new_[20047]_  = \new_[20046]_  & \new_[20041]_ ;
  assign \new_[20050]_  = A235 & A203;
  assign \new_[20054]_  = A269 & ~A266;
  assign \new_[20055]_  = A265 & \new_[20054]_ ;
  assign \new_[20056]_  = \new_[20055]_  & \new_[20050]_ ;
  assign \new_[20059]_  = ~A167 & ~A169;
  assign \new_[20063]_  = ~A200 & A199;
  assign \new_[20064]_  = ~A166 & \new_[20063]_ ;
  assign \new_[20065]_  = \new_[20064]_  & \new_[20059]_ ;
  assign \new_[20068]_  = A232 & A203;
  assign \new_[20072]_  = A300 & A299;
  assign \new_[20073]_  = A234 & \new_[20072]_ ;
  assign \new_[20074]_  = \new_[20073]_  & \new_[20068]_ ;
  assign \new_[20077]_  = ~A167 & ~A169;
  assign \new_[20081]_  = ~A200 & A199;
  assign \new_[20082]_  = ~A166 & \new_[20081]_ ;
  assign \new_[20083]_  = \new_[20082]_  & \new_[20077]_ ;
  assign \new_[20086]_  = A232 & A203;
  assign \new_[20090]_  = A300 & A298;
  assign \new_[20091]_  = A234 & \new_[20090]_ ;
  assign \new_[20092]_  = \new_[20091]_  & \new_[20086]_ ;
  assign \new_[20095]_  = ~A167 & ~A169;
  assign \new_[20099]_  = ~A200 & A199;
  assign \new_[20100]_  = ~A166 & \new_[20099]_ ;
  assign \new_[20101]_  = \new_[20100]_  & \new_[20095]_ ;
  assign \new_[20104]_  = A232 & A203;
  assign \new_[20108]_  = A267 & A265;
  assign \new_[20109]_  = A234 & \new_[20108]_ ;
  assign \new_[20110]_  = \new_[20109]_  & \new_[20104]_ ;
  assign \new_[20113]_  = ~A167 & ~A169;
  assign \new_[20117]_  = ~A200 & A199;
  assign \new_[20118]_  = ~A166 & \new_[20117]_ ;
  assign \new_[20119]_  = \new_[20118]_  & \new_[20113]_ ;
  assign \new_[20122]_  = A232 & A203;
  assign \new_[20126]_  = A267 & A266;
  assign \new_[20127]_  = A234 & \new_[20126]_ ;
  assign \new_[20128]_  = \new_[20127]_  & \new_[20122]_ ;
  assign \new_[20131]_  = ~A167 & ~A169;
  assign \new_[20135]_  = ~A200 & A199;
  assign \new_[20136]_  = ~A166 & \new_[20135]_ ;
  assign \new_[20137]_  = \new_[20136]_  & \new_[20131]_ ;
  assign \new_[20140]_  = A233 & A203;
  assign \new_[20144]_  = A300 & A299;
  assign \new_[20145]_  = A234 & \new_[20144]_ ;
  assign \new_[20146]_  = \new_[20145]_  & \new_[20140]_ ;
  assign \new_[20149]_  = ~A167 & ~A169;
  assign \new_[20153]_  = ~A200 & A199;
  assign \new_[20154]_  = ~A166 & \new_[20153]_ ;
  assign \new_[20155]_  = \new_[20154]_  & \new_[20149]_ ;
  assign \new_[20158]_  = A233 & A203;
  assign \new_[20162]_  = A300 & A298;
  assign \new_[20163]_  = A234 & \new_[20162]_ ;
  assign \new_[20164]_  = \new_[20163]_  & \new_[20158]_ ;
  assign \new_[20167]_  = ~A167 & ~A169;
  assign \new_[20171]_  = ~A200 & A199;
  assign \new_[20172]_  = ~A166 & \new_[20171]_ ;
  assign \new_[20173]_  = \new_[20172]_  & \new_[20167]_ ;
  assign \new_[20176]_  = A233 & A203;
  assign \new_[20180]_  = A267 & A265;
  assign \new_[20181]_  = A234 & \new_[20180]_ ;
  assign \new_[20182]_  = \new_[20181]_  & \new_[20176]_ ;
  assign \new_[20185]_  = ~A167 & ~A169;
  assign \new_[20189]_  = ~A200 & A199;
  assign \new_[20190]_  = ~A166 & \new_[20189]_ ;
  assign \new_[20191]_  = \new_[20190]_  & \new_[20185]_ ;
  assign \new_[20194]_  = A233 & A203;
  assign \new_[20198]_  = A267 & A266;
  assign \new_[20199]_  = A234 & \new_[20198]_ ;
  assign \new_[20200]_  = \new_[20199]_  & \new_[20194]_ ;
  assign \new_[20203]_  = ~A167 & ~A169;
  assign \new_[20207]_  = ~A200 & A199;
  assign \new_[20208]_  = ~A166 & \new_[20207]_ ;
  assign \new_[20209]_  = \new_[20208]_  & \new_[20203]_ ;
  assign \new_[20212]_  = ~A232 & A203;
  assign \new_[20216]_  = A301 & A236;
  assign \new_[20217]_  = A233 & \new_[20216]_ ;
  assign \new_[20218]_  = \new_[20217]_  & \new_[20212]_ ;
  assign \new_[20221]_  = ~A167 & ~A169;
  assign \new_[20225]_  = ~A200 & A199;
  assign \new_[20226]_  = ~A166 & \new_[20225]_ ;
  assign \new_[20227]_  = \new_[20226]_  & \new_[20221]_ ;
  assign \new_[20230]_  = ~A232 & A203;
  assign \new_[20234]_  = A268 & A236;
  assign \new_[20235]_  = A233 & \new_[20234]_ ;
  assign \new_[20236]_  = \new_[20235]_  & \new_[20230]_ ;
  assign \new_[20239]_  = ~A167 & ~A169;
  assign \new_[20243]_  = ~A200 & A199;
  assign \new_[20244]_  = ~A166 & \new_[20243]_ ;
  assign \new_[20245]_  = \new_[20244]_  & \new_[20239]_ ;
  assign \new_[20248]_  = A232 & A203;
  assign \new_[20252]_  = A301 & A236;
  assign \new_[20253]_  = ~A233 & \new_[20252]_ ;
  assign \new_[20254]_  = \new_[20253]_  & \new_[20248]_ ;
  assign \new_[20257]_  = ~A167 & ~A169;
  assign \new_[20261]_  = ~A200 & A199;
  assign \new_[20262]_  = ~A166 & \new_[20261]_ ;
  assign \new_[20263]_  = \new_[20262]_  & \new_[20257]_ ;
  assign \new_[20266]_  = A232 & A203;
  assign \new_[20270]_  = A268 & A236;
  assign \new_[20271]_  = ~A233 & \new_[20270]_ ;
  assign \new_[20272]_  = \new_[20271]_  & \new_[20266]_ ;
  assign \new_[20275]_  = ~A168 & ~A169;
  assign \new_[20279]_  = A202 & A166;
  assign \new_[20280]_  = A167 & \new_[20279]_ ;
  assign \new_[20281]_  = \new_[20280]_  & \new_[20275]_ ;
  assign \new_[20284]_  = A234 & A232;
  assign \new_[20288]_  = A302 & ~A299;
  assign \new_[20289]_  = A298 & \new_[20288]_ ;
  assign \new_[20290]_  = \new_[20289]_  & \new_[20284]_ ;
  assign \new_[20293]_  = ~A168 & ~A169;
  assign \new_[20297]_  = A202 & A166;
  assign \new_[20298]_  = A167 & \new_[20297]_ ;
  assign \new_[20299]_  = \new_[20298]_  & \new_[20293]_ ;
  assign \new_[20302]_  = A234 & A232;
  assign \new_[20306]_  = A302 & A299;
  assign \new_[20307]_  = ~A298 & \new_[20306]_ ;
  assign \new_[20308]_  = \new_[20307]_  & \new_[20302]_ ;
  assign \new_[20311]_  = ~A168 & ~A169;
  assign \new_[20315]_  = A202 & A166;
  assign \new_[20316]_  = A167 & \new_[20315]_ ;
  assign \new_[20317]_  = \new_[20316]_  & \new_[20311]_ ;
  assign \new_[20320]_  = A234 & A232;
  assign \new_[20324]_  = A269 & A266;
  assign \new_[20325]_  = ~A265 & \new_[20324]_ ;
  assign \new_[20326]_  = \new_[20325]_  & \new_[20320]_ ;
  assign \new_[20329]_  = ~A168 & ~A169;
  assign \new_[20333]_  = A202 & A166;
  assign \new_[20334]_  = A167 & \new_[20333]_ ;
  assign \new_[20335]_  = \new_[20334]_  & \new_[20329]_ ;
  assign \new_[20338]_  = A234 & A232;
  assign \new_[20342]_  = A269 & ~A266;
  assign \new_[20343]_  = A265 & \new_[20342]_ ;
  assign \new_[20344]_  = \new_[20343]_  & \new_[20338]_ ;
  assign \new_[20347]_  = ~A168 & ~A169;
  assign \new_[20351]_  = A202 & A166;
  assign \new_[20352]_  = A167 & \new_[20351]_ ;
  assign \new_[20353]_  = \new_[20352]_  & \new_[20347]_ ;
  assign \new_[20356]_  = A234 & A233;
  assign \new_[20360]_  = A302 & ~A299;
  assign \new_[20361]_  = A298 & \new_[20360]_ ;
  assign \new_[20362]_  = \new_[20361]_  & \new_[20356]_ ;
  assign \new_[20365]_  = ~A168 & ~A169;
  assign \new_[20369]_  = A202 & A166;
  assign \new_[20370]_  = A167 & \new_[20369]_ ;
  assign \new_[20371]_  = \new_[20370]_  & \new_[20365]_ ;
  assign \new_[20374]_  = A234 & A233;
  assign \new_[20378]_  = A302 & A299;
  assign \new_[20379]_  = ~A298 & \new_[20378]_ ;
  assign \new_[20380]_  = \new_[20379]_  & \new_[20374]_ ;
  assign \new_[20383]_  = ~A168 & ~A169;
  assign \new_[20387]_  = A202 & A166;
  assign \new_[20388]_  = A167 & \new_[20387]_ ;
  assign \new_[20389]_  = \new_[20388]_  & \new_[20383]_ ;
  assign \new_[20392]_  = A234 & A233;
  assign \new_[20396]_  = A269 & A266;
  assign \new_[20397]_  = ~A265 & \new_[20396]_ ;
  assign \new_[20398]_  = \new_[20397]_  & \new_[20392]_ ;
  assign \new_[20401]_  = ~A168 & ~A169;
  assign \new_[20405]_  = A202 & A166;
  assign \new_[20406]_  = A167 & \new_[20405]_ ;
  assign \new_[20407]_  = \new_[20406]_  & \new_[20401]_ ;
  assign \new_[20410]_  = A234 & A233;
  assign \new_[20414]_  = A269 & ~A266;
  assign \new_[20415]_  = A265 & \new_[20414]_ ;
  assign \new_[20416]_  = \new_[20415]_  & \new_[20410]_ ;
  assign \new_[20419]_  = ~A168 & ~A169;
  assign \new_[20423]_  = A202 & A166;
  assign \new_[20424]_  = A167 & \new_[20423]_ ;
  assign \new_[20425]_  = \new_[20424]_  & \new_[20419]_ ;
  assign \new_[20428]_  = A233 & ~A232;
  assign \new_[20432]_  = A300 & A299;
  assign \new_[20433]_  = A236 & \new_[20432]_ ;
  assign \new_[20434]_  = \new_[20433]_  & \new_[20428]_ ;
  assign \new_[20437]_  = ~A168 & ~A169;
  assign \new_[20441]_  = A202 & A166;
  assign \new_[20442]_  = A167 & \new_[20441]_ ;
  assign \new_[20443]_  = \new_[20442]_  & \new_[20437]_ ;
  assign \new_[20446]_  = A233 & ~A232;
  assign \new_[20450]_  = A300 & A298;
  assign \new_[20451]_  = A236 & \new_[20450]_ ;
  assign \new_[20452]_  = \new_[20451]_  & \new_[20446]_ ;
  assign \new_[20455]_  = ~A168 & ~A169;
  assign \new_[20459]_  = A202 & A166;
  assign \new_[20460]_  = A167 & \new_[20459]_ ;
  assign \new_[20461]_  = \new_[20460]_  & \new_[20455]_ ;
  assign \new_[20464]_  = A233 & ~A232;
  assign \new_[20468]_  = A267 & A265;
  assign \new_[20469]_  = A236 & \new_[20468]_ ;
  assign \new_[20470]_  = \new_[20469]_  & \new_[20464]_ ;
  assign \new_[20473]_  = ~A168 & ~A169;
  assign \new_[20477]_  = A202 & A166;
  assign \new_[20478]_  = A167 & \new_[20477]_ ;
  assign \new_[20479]_  = \new_[20478]_  & \new_[20473]_ ;
  assign \new_[20482]_  = A233 & ~A232;
  assign \new_[20486]_  = A267 & A266;
  assign \new_[20487]_  = A236 & \new_[20486]_ ;
  assign \new_[20488]_  = \new_[20487]_  & \new_[20482]_ ;
  assign \new_[20491]_  = ~A168 & ~A169;
  assign \new_[20495]_  = A202 & A166;
  assign \new_[20496]_  = A167 & \new_[20495]_ ;
  assign \new_[20497]_  = \new_[20496]_  & \new_[20491]_ ;
  assign \new_[20500]_  = ~A233 & A232;
  assign \new_[20504]_  = A300 & A299;
  assign \new_[20505]_  = A236 & \new_[20504]_ ;
  assign \new_[20506]_  = \new_[20505]_  & \new_[20500]_ ;
  assign \new_[20509]_  = ~A168 & ~A169;
  assign \new_[20513]_  = A202 & A166;
  assign \new_[20514]_  = A167 & \new_[20513]_ ;
  assign \new_[20515]_  = \new_[20514]_  & \new_[20509]_ ;
  assign \new_[20518]_  = ~A233 & A232;
  assign \new_[20522]_  = A300 & A298;
  assign \new_[20523]_  = A236 & \new_[20522]_ ;
  assign \new_[20524]_  = \new_[20523]_  & \new_[20518]_ ;
  assign \new_[20527]_  = ~A168 & ~A169;
  assign \new_[20531]_  = A202 & A166;
  assign \new_[20532]_  = A167 & \new_[20531]_ ;
  assign \new_[20533]_  = \new_[20532]_  & \new_[20527]_ ;
  assign \new_[20536]_  = ~A233 & A232;
  assign \new_[20540]_  = A267 & A265;
  assign \new_[20541]_  = A236 & \new_[20540]_ ;
  assign \new_[20542]_  = \new_[20541]_  & \new_[20536]_ ;
  assign \new_[20545]_  = ~A168 & ~A169;
  assign \new_[20549]_  = A202 & A166;
  assign \new_[20550]_  = A167 & \new_[20549]_ ;
  assign \new_[20551]_  = \new_[20550]_  & \new_[20545]_ ;
  assign \new_[20554]_  = ~A233 & A232;
  assign \new_[20558]_  = A267 & A266;
  assign \new_[20559]_  = A236 & \new_[20558]_ ;
  assign \new_[20560]_  = \new_[20559]_  & \new_[20554]_ ;
  assign \new_[20563]_  = ~A168 & ~A169;
  assign \new_[20567]_  = A199 & A166;
  assign \new_[20568]_  = A167 & \new_[20567]_ ;
  assign \new_[20569]_  = \new_[20568]_  & \new_[20563]_ ;
  assign \new_[20572]_  = A235 & A201;
  assign \new_[20576]_  = A302 & ~A299;
  assign \new_[20577]_  = A298 & \new_[20576]_ ;
  assign \new_[20578]_  = \new_[20577]_  & \new_[20572]_ ;
  assign \new_[20581]_  = ~A168 & ~A169;
  assign \new_[20585]_  = A199 & A166;
  assign \new_[20586]_  = A167 & \new_[20585]_ ;
  assign \new_[20587]_  = \new_[20586]_  & \new_[20581]_ ;
  assign \new_[20590]_  = A235 & A201;
  assign \new_[20594]_  = A302 & A299;
  assign \new_[20595]_  = ~A298 & \new_[20594]_ ;
  assign \new_[20596]_  = \new_[20595]_  & \new_[20590]_ ;
  assign \new_[20599]_  = ~A168 & ~A169;
  assign \new_[20603]_  = A199 & A166;
  assign \new_[20604]_  = A167 & \new_[20603]_ ;
  assign \new_[20605]_  = \new_[20604]_  & \new_[20599]_ ;
  assign \new_[20608]_  = A235 & A201;
  assign \new_[20612]_  = A269 & A266;
  assign \new_[20613]_  = ~A265 & \new_[20612]_ ;
  assign \new_[20614]_  = \new_[20613]_  & \new_[20608]_ ;
  assign \new_[20617]_  = ~A168 & ~A169;
  assign \new_[20621]_  = A199 & A166;
  assign \new_[20622]_  = A167 & \new_[20621]_ ;
  assign \new_[20623]_  = \new_[20622]_  & \new_[20617]_ ;
  assign \new_[20626]_  = A235 & A201;
  assign \new_[20630]_  = A269 & ~A266;
  assign \new_[20631]_  = A265 & \new_[20630]_ ;
  assign \new_[20632]_  = \new_[20631]_  & \new_[20626]_ ;
  assign \new_[20635]_  = ~A168 & ~A169;
  assign \new_[20639]_  = A199 & A166;
  assign \new_[20640]_  = A167 & \new_[20639]_ ;
  assign \new_[20641]_  = \new_[20640]_  & \new_[20635]_ ;
  assign \new_[20644]_  = A232 & A201;
  assign \new_[20648]_  = A300 & A299;
  assign \new_[20649]_  = A234 & \new_[20648]_ ;
  assign \new_[20650]_  = \new_[20649]_  & \new_[20644]_ ;
  assign \new_[20653]_  = ~A168 & ~A169;
  assign \new_[20657]_  = A199 & A166;
  assign \new_[20658]_  = A167 & \new_[20657]_ ;
  assign \new_[20659]_  = \new_[20658]_  & \new_[20653]_ ;
  assign \new_[20662]_  = A232 & A201;
  assign \new_[20666]_  = A300 & A298;
  assign \new_[20667]_  = A234 & \new_[20666]_ ;
  assign \new_[20668]_  = \new_[20667]_  & \new_[20662]_ ;
  assign \new_[20671]_  = ~A168 & ~A169;
  assign \new_[20675]_  = A199 & A166;
  assign \new_[20676]_  = A167 & \new_[20675]_ ;
  assign \new_[20677]_  = \new_[20676]_  & \new_[20671]_ ;
  assign \new_[20680]_  = A232 & A201;
  assign \new_[20684]_  = A267 & A265;
  assign \new_[20685]_  = A234 & \new_[20684]_ ;
  assign \new_[20686]_  = \new_[20685]_  & \new_[20680]_ ;
  assign \new_[20689]_  = ~A168 & ~A169;
  assign \new_[20693]_  = A199 & A166;
  assign \new_[20694]_  = A167 & \new_[20693]_ ;
  assign \new_[20695]_  = \new_[20694]_  & \new_[20689]_ ;
  assign \new_[20698]_  = A232 & A201;
  assign \new_[20702]_  = A267 & A266;
  assign \new_[20703]_  = A234 & \new_[20702]_ ;
  assign \new_[20704]_  = \new_[20703]_  & \new_[20698]_ ;
  assign \new_[20707]_  = ~A168 & ~A169;
  assign \new_[20711]_  = A199 & A166;
  assign \new_[20712]_  = A167 & \new_[20711]_ ;
  assign \new_[20713]_  = \new_[20712]_  & \new_[20707]_ ;
  assign \new_[20716]_  = A233 & A201;
  assign \new_[20720]_  = A300 & A299;
  assign \new_[20721]_  = A234 & \new_[20720]_ ;
  assign \new_[20722]_  = \new_[20721]_  & \new_[20716]_ ;
  assign \new_[20725]_  = ~A168 & ~A169;
  assign \new_[20729]_  = A199 & A166;
  assign \new_[20730]_  = A167 & \new_[20729]_ ;
  assign \new_[20731]_  = \new_[20730]_  & \new_[20725]_ ;
  assign \new_[20734]_  = A233 & A201;
  assign \new_[20738]_  = A300 & A298;
  assign \new_[20739]_  = A234 & \new_[20738]_ ;
  assign \new_[20740]_  = \new_[20739]_  & \new_[20734]_ ;
  assign \new_[20743]_  = ~A168 & ~A169;
  assign \new_[20747]_  = A199 & A166;
  assign \new_[20748]_  = A167 & \new_[20747]_ ;
  assign \new_[20749]_  = \new_[20748]_  & \new_[20743]_ ;
  assign \new_[20752]_  = A233 & A201;
  assign \new_[20756]_  = A267 & A265;
  assign \new_[20757]_  = A234 & \new_[20756]_ ;
  assign \new_[20758]_  = \new_[20757]_  & \new_[20752]_ ;
  assign \new_[20761]_  = ~A168 & ~A169;
  assign \new_[20765]_  = A199 & A166;
  assign \new_[20766]_  = A167 & \new_[20765]_ ;
  assign \new_[20767]_  = \new_[20766]_  & \new_[20761]_ ;
  assign \new_[20770]_  = A233 & A201;
  assign \new_[20774]_  = A267 & A266;
  assign \new_[20775]_  = A234 & \new_[20774]_ ;
  assign \new_[20776]_  = \new_[20775]_  & \new_[20770]_ ;
  assign \new_[20779]_  = ~A168 & ~A169;
  assign \new_[20783]_  = A199 & A166;
  assign \new_[20784]_  = A167 & \new_[20783]_ ;
  assign \new_[20785]_  = \new_[20784]_  & \new_[20779]_ ;
  assign \new_[20788]_  = ~A232 & A201;
  assign \new_[20792]_  = A301 & A236;
  assign \new_[20793]_  = A233 & \new_[20792]_ ;
  assign \new_[20794]_  = \new_[20793]_  & \new_[20788]_ ;
  assign \new_[20797]_  = ~A168 & ~A169;
  assign \new_[20801]_  = A199 & A166;
  assign \new_[20802]_  = A167 & \new_[20801]_ ;
  assign \new_[20803]_  = \new_[20802]_  & \new_[20797]_ ;
  assign \new_[20806]_  = ~A232 & A201;
  assign \new_[20810]_  = A268 & A236;
  assign \new_[20811]_  = A233 & \new_[20810]_ ;
  assign \new_[20812]_  = \new_[20811]_  & \new_[20806]_ ;
  assign \new_[20815]_  = ~A168 & ~A169;
  assign \new_[20819]_  = A199 & A166;
  assign \new_[20820]_  = A167 & \new_[20819]_ ;
  assign \new_[20821]_  = \new_[20820]_  & \new_[20815]_ ;
  assign \new_[20824]_  = A232 & A201;
  assign \new_[20828]_  = A301 & A236;
  assign \new_[20829]_  = ~A233 & \new_[20828]_ ;
  assign \new_[20830]_  = \new_[20829]_  & \new_[20824]_ ;
  assign \new_[20833]_  = ~A168 & ~A169;
  assign \new_[20837]_  = A199 & A166;
  assign \new_[20838]_  = A167 & \new_[20837]_ ;
  assign \new_[20839]_  = \new_[20838]_  & \new_[20833]_ ;
  assign \new_[20842]_  = A232 & A201;
  assign \new_[20846]_  = A268 & A236;
  assign \new_[20847]_  = ~A233 & \new_[20846]_ ;
  assign \new_[20848]_  = \new_[20847]_  & \new_[20842]_ ;
  assign \new_[20851]_  = ~A168 & ~A169;
  assign \new_[20855]_  = A200 & A166;
  assign \new_[20856]_  = A167 & \new_[20855]_ ;
  assign \new_[20857]_  = \new_[20856]_  & \new_[20851]_ ;
  assign \new_[20860]_  = A235 & A201;
  assign \new_[20864]_  = A302 & ~A299;
  assign \new_[20865]_  = A298 & \new_[20864]_ ;
  assign \new_[20866]_  = \new_[20865]_  & \new_[20860]_ ;
  assign \new_[20869]_  = ~A168 & ~A169;
  assign \new_[20873]_  = A200 & A166;
  assign \new_[20874]_  = A167 & \new_[20873]_ ;
  assign \new_[20875]_  = \new_[20874]_  & \new_[20869]_ ;
  assign \new_[20878]_  = A235 & A201;
  assign \new_[20882]_  = A302 & A299;
  assign \new_[20883]_  = ~A298 & \new_[20882]_ ;
  assign \new_[20884]_  = \new_[20883]_  & \new_[20878]_ ;
  assign \new_[20887]_  = ~A168 & ~A169;
  assign \new_[20891]_  = A200 & A166;
  assign \new_[20892]_  = A167 & \new_[20891]_ ;
  assign \new_[20893]_  = \new_[20892]_  & \new_[20887]_ ;
  assign \new_[20896]_  = A235 & A201;
  assign \new_[20900]_  = A269 & A266;
  assign \new_[20901]_  = ~A265 & \new_[20900]_ ;
  assign \new_[20902]_  = \new_[20901]_  & \new_[20896]_ ;
  assign \new_[20905]_  = ~A168 & ~A169;
  assign \new_[20909]_  = A200 & A166;
  assign \new_[20910]_  = A167 & \new_[20909]_ ;
  assign \new_[20911]_  = \new_[20910]_  & \new_[20905]_ ;
  assign \new_[20914]_  = A235 & A201;
  assign \new_[20918]_  = A269 & ~A266;
  assign \new_[20919]_  = A265 & \new_[20918]_ ;
  assign \new_[20920]_  = \new_[20919]_  & \new_[20914]_ ;
  assign \new_[20923]_  = ~A168 & ~A169;
  assign \new_[20927]_  = A200 & A166;
  assign \new_[20928]_  = A167 & \new_[20927]_ ;
  assign \new_[20929]_  = \new_[20928]_  & \new_[20923]_ ;
  assign \new_[20932]_  = A232 & A201;
  assign \new_[20936]_  = A300 & A299;
  assign \new_[20937]_  = A234 & \new_[20936]_ ;
  assign \new_[20938]_  = \new_[20937]_  & \new_[20932]_ ;
  assign \new_[20941]_  = ~A168 & ~A169;
  assign \new_[20945]_  = A200 & A166;
  assign \new_[20946]_  = A167 & \new_[20945]_ ;
  assign \new_[20947]_  = \new_[20946]_  & \new_[20941]_ ;
  assign \new_[20950]_  = A232 & A201;
  assign \new_[20954]_  = A300 & A298;
  assign \new_[20955]_  = A234 & \new_[20954]_ ;
  assign \new_[20956]_  = \new_[20955]_  & \new_[20950]_ ;
  assign \new_[20959]_  = ~A168 & ~A169;
  assign \new_[20963]_  = A200 & A166;
  assign \new_[20964]_  = A167 & \new_[20963]_ ;
  assign \new_[20965]_  = \new_[20964]_  & \new_[20959]_ ;
  assign \new_[20968]_  = A232 & A201;
  assign \new_[20972]_  = A267 & A265;
  assign \new_[20973]_  = A234 & \new_[20972]_ ;
  assign \new_[20974]_  = \new_[20973]_  & \new_[20968]_ ;
  assign \new_[20977]_  = ~A168 & ~A169;
  assign \new_[20981]_  = A200 & A166;
  assign \new_[20982]_  = A167 & \new_[20981]_ ;
  assign \new_[20983]_  = \new_[20982]_  & \new_[20977]_ ;
  assign \new_[20986]_  = A232 & A201;
  assign \new_[20990]_  = A267 & A266;
  assign \new_[20991]_  = A234 & \new_[20990]_ ;
  assign \new_[20992]_  = \new_[20991]_  & \new_[20986]_ ;
  assign \new_[20995]_  = ~A168 & ~A169;
  assign \new_[20999]_  = A200 & A166;
  assign \new_[21000]_  = A167 & \new_[20999]_ ;
  assign \new_[21001]_  = \new_[21000]_  & \new_[20995]_ ;
  assign \new_[21004]_  = A233 & A201;
  assign \new_[21008]_  = A300 & A299;
  assign \new_[21009]_  = A234 & \new_[21008]_ ;
  assign \new_[21010]_  = \new_[21009]_  & \new_[21004]_ ;
  assign \new_[21013]_  = ~A168 & ~A169;
  assign \new_[21017]_  = A200 & A166;
  assign \new_[21018]_  = A167 & \new_[21017]_ ;
  assign \new_[21019]_  = \new_[21018]_  & \new_[21013]_ ;
  assign \new_[21022]_  = A233 & A201;
  assign \new_[21026]_  = A300 & A298;
  assign \new_[21027]_  = A234 & \new_[21026]_ ;
  assign \new_[21028]_  = \new_[21027]_  & \new_[21022]_ ;
  assign \new_[21031]_  = ~A168 & ~A169;
  assign \new_[21035]_  = A200 & A166;
  assign \new_[21036]_  = A167 & \new_[21035]_ ;
  assign \new_[21037]_  = \new_[21036]_  & \new_[21031]_ ;
  assign \new_[21040]_  = A233 & A201;
  assign \new_[21044]_  = A267 & A265;
  assign \new_[21045]_  = A234 & \new_[21044]_ ;
  assign \new_[21046]_  = \new_[21045]_  & \new_[21040]_ ;
  assign \new_[21049]_  = ~A168 & ~A169;
  assign \new_[21053]_  = A200 & A166;
  assign \new_[21054]_  = A167 & \new_[21053]_ ;
  assign \new_[21055]_  = \new_[21054]_  & \new_[21049]_ ;
  assign \new_[21058]_  = A233 & A201;
  assign \new_[21062]_  = A267 & A266;
  assign \new_[21063]_  = A234 & \new_[21062]_ ;
  assign \new_[21064]_  = \new_[21063]_  & \new_[21058]_ ;
  assign \new_[21067]_  = ~A168 & ~A169;
  assign \new_[21071]_  = A200 & A166;
  assign \new_[21072]_  = A167 & \new_[21071]_ ;
  assign \new_[21073]_  = \new_[21072]_  & \new_[21067]_ ;
  assign \new_[21076]_  = ~A232 & A201;
  assign \new_[21080]_  = A301 & A236;
  assign \new_[21081]_  = A233 & \new_[21080]_ ;
  assign \new_[21082]_  = \new_[21081]_  & \new_[21076]_ ;
  assign \new_[21085]_  = ~A168 & ~A169;
  assign \new_[21089]_  = A200 & A166;
  assign \new_[21090]_  = A167 & \new_[21089]_ ;
  assign \new_[21091]_  = \new_[21090]_  & \new_[21085]_ ;
  assign \new_[21094]_  = ~A232 & A201;
  assign \new_[21098]_  = A268 & A236;
  assign \new_[21099]_  = A233 & \new_[21098]_ ;
  assign \new_[21100]_  = \new_[21099]_  & \new_[21094]_ ;
  assign \new_[21103]_  = ~A168 & ~A169;
  assign \new_[21107]_  = A200 & A166;
  assign \new_[21108]_  = A167 & \new_[21107]_ ;
  assign \new_[21109]_  = \new_[21108]_  & \new_[21103]_ ;
  assign \new_[21112]_  = A232 & A201;
  assign \new_[21116]_  = A301 & A236;
  assign \new_[21117]_  = ~A233 & \new_[21116]_ ;
  assign \new_[21118]_  = \new_[21117]_  & \new_[21112]_ ;
  assign \new_[21121]_  = ~A168 & ~A169;
  assign \new_[21125]_  = A200 & A166;
  assign \new_[21126]_  = A167 & \new_[21125]_ ;
  assign \new_[21127]_  = \new_[21126]_  & \new_[21121]_ ;
  assign \new_[21130]_  = A232 & A201;
  assign \new_[21134]_  = A268 & A236;
  assign \new_[21135]_  = ~A233 & \new_[21134]_ ;
  assign \new_[21136]_  = \new_[21135]_  & \new_[21130]_ ;
  assign \new_[21139]_  = ~A168 & ~A169;
  assign \new_[21143]_  = ~A199 & A166;
  assign \new_[21144]_  = A167 & \new_[21143]_ ;
  assign \new_[21145]_  = \new_[21144]_  & \new_[21139]_ ;
  assign \new_[21148]_  = A203 & A200;
  assign \new_[21152]_  = A300 & A299;
  assign \new_[21153]_  = A235 & \new_[21152]_ ;
  assign \new_[21154]_  = \new_[21153]_  & \new_[21148]_ ;
  assign \new_[21157]_  = ~A168 & ~A169;
  assign \new_[21161]_  = ~A199 & A166;
  assign \new_[21162]_  = A167 & \new_[21161]_ ;
  assign \new_[21163]_  = \new_[21162]_  & \new_[21157]_ ;
  assign \new_[21166]_  = A203 & A200;
  assign \new_[21170]_  = A300 & A298;
  assign \new_[21171]_  = A235 & \new_[21170]_ ;
  assign \new_[21172]_  = \new_[21171]_  & \new_[21166]_ ;
  assign \new_[21175]_  = ~A168 & ~A169;
  assign \new_[21179]_  = ~A199 & A166;
  assign \new_[21180]_  = A167 & \new_[21179]_ ;
  assign \new_[21181]_  = \new_[21180]_  & \new_[21175]_ ;
  assign \new_[21184]_  = A203 & A200;
  assign \new_[21188]_  = A267 & A265;
  assign \new_[21189]_  = A235 & \new_[21188]_ ;
  assign \new_[21190]_  = \new_[21189]_  & \new_[21184]_ ;
  assign \new_[21193]_  = ~A168 & ~A169;
  assign \new_[21197]_  = ~A199 & A166;
  assign \new_[21198]_  = A167 & \new_[21197]_ ;
  assign \new_[21199]_  = \new_[21198]_  & \new_[21193]_ ;
  assign \new_[21202]_  = A203 & A200;
  assign \new_[21206]_  = A267 & A266;
  assign \new_[21207]_  = A235 & \new_[21206]_ ;
  assign \new_[21208]_  = \new_[21207]_  & \new_[21202]_ ;
  assign \new_[21211]_  = ~A168 & ~A169;
  assign \new_[21215]_  = ~A199 & A166;
  assign \new_[21216]_  = A167 & \new_[21215]_ ;
  assign \new_[21217]_  = \new_[21216]_  & \new_[21211]_ ;
  assign \new_[21220]_  = A203 & A200;
  assign \new_[21224]_  = A301 & A234;
  assign \new_[21225]_  = A232 & \new_[21224]_ ;
  assign \new_[21226]_  = \new_[21225]_  & \new_[21220]_ ;
  assign \new_[21229]_  = ~A168 & ~A169;
  assign \new_[21233]_  = ~A199 & A166;
  assign \new_[21234]_  = A167 & \new_[21233]_ ;
  assign \new_[21235]_  = \new_[21234]_  & \new_[21229]_ ;
  assign \new_[21238]_  = A203 & A200;
  assign \new_[21242]_  = A268 & A234;
  assign \new_[21243]_  = A232 & \new_[21242]_ ;
  assign \new_[21244]_  = \new_[21243]_  & \new_[21238]_ ;
  assign \new_[21247]_  = ~A168 & ~A169;
  assign \new_[21251]_  = ~A199 & A166;
  assign \new_[21252]_  = A167 & \new_[21251]_ ;
  assign \new_[21253]_  = \new_[21252]_  & \new_[21247]_ ;
  assign \new_[21256]_  = A203 & A200;
  assign \new_[21260]_  = A301 & A234;
  assign \new_[21261]_  = A233 & \new_[21260]_ ;
  assign \new_[21262]_  = \new_[21261]_  & \new_[21256]_ ;
  assign \new_[21265]_  = ~A168 & ~A169;
  assign \new_[21269]_  = ~A199 & A166;
  assign \new_[21270]_  = A167 & \new_[21269]_ ;
  assign \new_[21271]_  = \new_[21270]_  & \new_[21265]_ ;
  assign \new_[21274]_  = A203 & A200;
  assign \new_[21278]_  = A268 & A234;
  assign \new_[21279]_  = A233 & \new_[21278]_ ;
  assign \new_[21280]_  = \new_[21279]_  & \new_[21274]_ ;
  assign \new_[21283]_  = ~A168 & ~A169;
  assign \new_[21287]_  = A199 & A166;
  assign \new_[21288]_  = A167 & \new_[21287]_ ;
  assign \new_[21289]_  = \new_[21288]_  & \new_[21283]_ ;
  assign \new_[21292]_  = A203 & ~A200;
  assign \new_[21296]_  = A300 & A299;
  assign \new_[21297]_  = A235 & \new_[21296]_ ;
  assign \new_[21298]_  = \new_[21297]_  & \new_[21292]_ ;
  assign \new_[21301]_  = ~A168 & ~A169;
  assign \new_[21305]_  = A199 & A166;
  assign \new_[21306]_  = A167 & \new_[21305]_ ;
  assign \new_[21307]_  = \new_[21306]_  & \new_[21301]_ ;
  assign \new_[21310]_  = A203 & ~A200;
  assign \new_[21314]_  = A300 & A298;
  assign \new_[21315]_  = A235 & \new_[21314]_ ;
  assign \new_[21316]_  = \new_[21315]_  & \new_[21310]_ ;
  assign \new_[21319]_  = ~A168 & ~A169;
  assign \new_[21323]_  = A199 & A166;
  assign \new_[21324]_  = A167 & \new_[21323]_ ;
  assign \new_[21325]_  = \new_[21324]_  & \new_[21319]_ ;
  assign \new_[21328]_  = A203 & ~A200;
  assign \new_[21332]_  = A267 & A265;
  assign \new_[21333]_  = A235 & \new_[21332]_ ;
  assign \new_[21334]_  = \new_[21333]_  & \new_[21328]_ ;
  assign \new_[21337]_  = ~A168 & ~A169;
  assign \new_[21341]_  = A199 & A166;
  assign \new_[21342]_  = A167 & \new_[21341]_ ;
  assign \new_[21343]_  = \new_[21342]_  & \new_[21337]_ ;
  assign \new_[21346]_  = A203 & ~A200;
  assign \new_[21350]_  = A267 & A266;
  assign \new_[21351]_  = A235 & \new_[21350]_ ;
  assign \new_[21352]_  = \new_[21351]_  & \new_[21346]_ ;
  assign \new_[21355]_  = ~A168 & ~A169;
  assign \new_[21359]_  = A199 & A166;
  assign \new_[21360]_  = A167 & \new_[21359]_ ;
  assign \new_[21361]_  = \new_[21360]_  & \new_[21355]_ ;
  assign \new_[21364]_  = A203 & ~A200;
  assign \new_[21368]_  = A301 & A234;
  assign \new_[21369]_  = A232 & \new_[21368]_ ;
  assign \new_[21370]_  = \new_[21369]_  & \new_[21364]_ ;
  assign \new_[21373]_  = ~A168 & ~A169;
  assign \new_[21377]_  = A199 & A166;
  assign \new_[21378]_  = A167 & \new_[21377]_ ;
  assign \new_[21379]_  = \new_[21378]_  & \new_[21373]_ ;
  assign \new_[21382]_  = A203 & ~A200;
  assign \new_[21386]_  = A268 & A234;
  assign \new_[21387]_  = A232 & \new_[21386]_ ;
  assign \new_[21388]_  = \new_[21387]_  & \new_[21382]_ ;
  assign \new_[21391]_  = ~A168 & ~A169;
  assign \new_[21395]_  = A199 & A166;
  assign \new_[21396]_  = A167 & \new_[21395]_ ;
  assign \new_[21397]_  = \new_[21396]_  & \new_[21391]_ ;
  assign \new_[21400]_  = A203 & ~A200;
  assign \new_[21404]_  = A301 & A234;
  assign \new_[21405]_  = A233 & \new_[21404]_ ;
  assign \new_[21406]_  = \new_[21405]_  & \new_[21400]_ ;
  assign \new_[21409]_  = ~A168 & ~A169;
  assign \new_[21413]_  = A199 & A166;
  assign \new_[21414]_  = A167 & \new_[21413]_ ;
  assign \new_[21415]_  = \new_[21414]_  & \new_[21409]_ ;
  assign \new_[21418]_  = A203 & ~A200;
  assign \new_[21422]_  = A268 & A234;
  assign \new_[21423]_  = A233 & \new_[21422]_ ;
  assign \new_[21424]_  = \new_[21423]_  & \new_[21418]_ ;
  assign \new_[21427]_  = ~A169 & ~A170;
  assign \new_[21431]_  = ~A232 & A202;
  assign \new_[21432]_  = ~A168 & \new_[21431]_ ;
  assign \new_[21433]_  = \new_[21432]_  & \new_[21427]_ ;
  assign \new_[21436]_  = A236 & A233;
  assign \new_[21440]_  = A302 & ~A299;
  assign \new_[21441]_  = A298 & \new_[21440]_ ;
  assign \new_[21442]_  = \new_[21441]_  & \new_[21436]_ ;
  assign \new_[21445]_  = ~A169 & ~A170;
  assign \new_[21449]_  = ~A232 & A202;
  assign \new_[21450]_  = ~A168 & \new_[21449]_ ;
  assign \new_[21451]_  = \new_[21450]_  & \new_[21445]_ ;
  assign \new_[21454]_  = A236 & A233;
  assign \new_[21458]_  = A302 & A299;
  assign \new_[21459]_  = ~A298 & \new_[21458]_ ;
  assign \new_[21460]_  = \new_[21459]_  & \new_[21454]_ ;
  assign \new_[21463]_  = ~A169 & ~A170;
  assign \new_[21467]_  = ~A232 & A202;
  assign \new_[21468]_  = ~A168 & \new_[21467]_ ;
  assign \new_[21469]_  = \new_[21468]_  & \new_[21463]_ ;
  assign \new_[21472]_  = A236 & A233;
  assign \new_[21476]_  = A269 & A266;
  assign \new_[21477]_  = ~A265 & \new_[21476]_ ;
  assign \new_[21478]_  = \new_[21477]_  & \new_[21472]_ ;
  assign \new_[21481]_  = ~A169 & ~A170;
  assign \new_[21485]_  = ~A232 & A202;
  assign \new_[21486]_  = ~A168 & \new_[21485]_ ;
  assign \new_[21487]_  = \new_[21486]_  & \new_[21481]_ ;
  assign \new_[21490]_  = A236 & A233;
  assign \new_[21494]_  = A269 & ~A266;
  assign \new_[21495]_  = A265 & \new_[21494]_ ;
  assign \new_[21496]_  = \new_[21495]_  & \new_[21490]_ ;
  assign \new_[21499]_  = ~A169 & ~A170;
  assign \new_[21503]_  = A232 & A202;
  assign \new_[21504]_  = ~A168 & \new_[21503]_ ;
  assign \new_[21505]_  = \new_[21504]_  & \new_[21499]_ ;
  assign \new_[21508]_  = A236 & ~A233;
  assign \new_[21512]_  = A302 & ~A299;
  assign \new_[21513]_  = A298 & \new_[21512]_ ;
  assign \new_[21514]_  = \new_[21513]_  & \new_[21508]_ ;
  assign \new_[21517]_  = ~A169 & ~A170;
  assign \new_[21521]_  = A232 & A202;
  assign \new_[21522]_  = ~A168 & \new_[21521]_ ;
  assign \new_[21523]_  = \new_[21522]_  & \new_[21517]_ ;
  assign \new_[21526]_  = A236 & ~A233;
  assign \new_[21530]_  = A302 & A299;
  assign \new_[21531]_  = ~A298 & \new_[21530]_ ;
  assign \new_[21532]_  = \new_[21531]_  & \new_[21526]_ ;
  assign \new_[21535]_  = ~A169 & ~A170;
  assign \new_[21539]_  = A232 & A202;
  assign \new_[21540]_  = ~A168 & \new_[21539]_ ;
  assign \new_[21541]_  = \new_[21540]_  & \new_[21535]_ ;
  assign \new_[21544]_  = A236 & ~A233;
  assign \new_[21548]_  = A269 & A266;
  assign \new_[21549]_  = ~A265 & \new_[21548]_ ;
  assign \new_[21550]_  = \new_[21549]_  & \new_[21544]_ ;
  assign \new_[21553]_  = ~A169 & ~A170;
  assign \new_[21557]_  = A232 & A202;
  assign \new_[21558]_  = ~A168 & \new_[21557]_ ;
  assign \new_[21559]_  = \new_[21558]_  & \new_[21553]_ ;
  assign \new_[21562]_  = A236 & ~A233;
  assign \new_[21566]_  = A269 & ~A266;
  assign \new_[21567]_  = A265 & \new_[21566]_ ;
  assign \new_[21568]_  = \new_[21567]_  & \new_[21562]_ ;
  assign \new_[21571]_  = ~A169 & ~A170;
  assign \new_[21575]_  = A201 & A199;
  assign \new_[21576]_  = ~A168 & \new_[21575]_ ;
  assign \new_[21577]_  = \new_[21576]_  & \new_[21571]_ ;
  assign \new_[21580]_  = A234 & A232;
  assign \new_[21584]_  = A302 & ~A299;
  assign \new_[21585]_  = A298 & \new_[21584]_ ;
  assign \new_[21586]_  = \new_[21585]_  & \new_[21580]_ ;
  assign \new_[21589]_  = ~A169 & ~A170;
  assign \new_[21593]_  = A201 & A199;
  assign \new_[21594]_  = ~A168 & \new_[21593]_ ;
  assign \new_[21595]_  = \new_[21594]_  & \new_[21589]_ ;
  assign \new_[21598]_  = A234 & A232;
  assign \new_[21602]_  = A302 & A299;
  assign \new_[21603]_  = ~A298 & \new_[21602]_ ;
  assign \new_[21604]_  = \new_[21603]_  & \new_[21598]_ ;
  assign \new_[21607]_  = ~A169 & ~A170;
  assign \new_[21611]_  = A201 & A199;
  assign \new_[21612]_  = ~A168 & \new_[21611]_ ;
  assign \new_[21613]_  = \new_[21612]_  & \new_[21607]_ ;
  assign \new_[21616]_  = A234 & A232;
  assign \new_[21620]_  = A269 & A266;
  assign \new_[21621]_  = ~A265 & \new_[21620]_ ;
  assign \new_[21622]_  = \new_[21621]_  & \new_[21616]_ ;
  assign \new_[21625]_  = ~A169 & ~A170;
  assign \new_[21629]_  = A201 & A199;
  assign \new_[21630]_  = ~A168 & \new_[21629]_ ;
  assign \new_[21631]_  = \new_[21630]_  & \new_[21625]_ ;
  assign \new_[21634]_  = A234 & A232;
  assign \new_[21638]_  = A269 & ~A266;
  assign \new_[21639]_  = A265 & \new_[21638]_ ;
  assign \new_[21640]_  = \new_[21639]_  & \new_[21634]_ ;
  assign \new_[21643]_  = ~A169 & ~A170;
  assign \new_[21647]_  = A201 & A199;
  assign \new_[21648]_  = ~A168 & \new_[21647]_ ;
  assign \new_[21649]_  = \new_[21648]_  & \new_[21643]_ ;
  assign \new_[21652]_  = A234 & A233;
  assign \new_[21656]_  = A302 & ~A299;
  assign \new_[21657]_  = A298 & \new_[21656]_ ;
  assign \new_[21658]_  = \new_[21657]_  & \new_[21652]_ ;
  assign \new_[21661]_  = ~A169 & ~A170;
  assign \new_[21665]_  = A201 & A199;
  assign \new_[21666]_  = ~A168 & \new_[21665]_ ;
  assign \new_[21667]_  = \new_[21666]_  & \new_[21661]_ ;
  assign \new_[21670]_  = A234 & A233;
  assign \new_[21674]_  = A302 & A299;
  assign \new_[21675]_  = ~A298 & \new_[21674]_ ;
  assign \new_[21676]_  = \new_[21675]_  & \new_[21670]_ ;
  assign \new_[21679]_  = ~A169 & ~A170;
  assign \new_[21683]_  = A201 & A199;
  assign \new_[21684]_  = ~A168 & \new_[21683]_ ;
  assign \new_[21685]_  = \new_[21684]_  & \new_[21679]_ ;
  assign \new_[21688]_  = A234 & A233;
  assign \new_[21692]_  = A269 & A266;
  assign \new_[21693]_  = ~A265 & \new_[21692]_ ;
  assign \new_[21694]_  = \new_[21693]_  & \new_[21688]_ ;
  assign \new_[21697]_  = ~A169 & ~A170;
  assign \new_[21701]_  = A201 & A199;
  assign \new_[21702]_  = ~A168 & \new_[21701]_ ;
  assign \new_[21703]_  = \new_[21702]_  & \new_[21697]_ ;
  assign \new_[21706]_  = A234 & A233;
  assign \new_[21710]_  = A269 & ~A266;
  assign \new_[21711]_  = A265 & \new_[21710]_ ;
  assign \new_[21712]_  = \new_[21711]_  & \new_[21706]_ ;
  assign \new_[21715]_  = ~A169 & ~A170;
  assign \new_[21719]_  = A201 & A199;
  assign \new_[21720]_  = ~A168 & \new_[21719]_ ;
  assign \new_[21721]_  = \new_[21720]_  & \new_[21715]_ ;
  assign \new_[21724]_  = A233 & ~A232;
  assign \new_[21728]_  = A300 & A299;
  assign \new_[21729]_  = A236 & \new_[21728]_ ;
  assign \new_[21730]_  = \new_[21729]_  & \new_[21724]_ ;
  assign \new_[21733]_  = ~A169 & ~A170;
  assign \new_[21737]_  = A201 & A199;
  assign \new_[21738]_  = ~A168 & \new_[21737]_ ;
  assign \new_[21739]_  = \new_[21738]_  & \new_[21733]_ ;
  assign \new_[21742]_  = A233 & ~A232;
  assign \new_[21746]_  = A300 & A298;
  assign \new_[21747]_  = A236 & \new_[21746]_ ;
  assign \new_[21748]_  = \new_[21747]_  & \new_[21742]_ ;
  assign \new_[21751]_  = ~A169 & ~A170;
  assign \new_[21755]_  = A201 & A199;
  assign \new_[21756]_  = ~A168 & \new_[21755]_ ;
  assign \new_[21757]_  = \new_[21756]_  & \new_[21751]_ ;
  assign \new_[21760]_  = A233 & ~A232;
  assign \new_[21764]_  = A267 & A265;
  assign \new_[21765]_  = A236 & \new_[21764]_ ;
  assign \new_[21766]_  = \new_[21765]_  & \new_[21760]_ ;
  assign \new_[21769]_  = ~A169 & ~A170;
  assign \new_[21773]_  = A201 & A199;
  assign \new_[21774]_  = ~A168 & \new_[21773]_ ;
  assign \new_[21775]_  = \new_[21774]_  & \new_[21769]_ ;
  assign \new_[21778]_  = A233 & ~A232;
  assign \new_[21782]_  = A267 & A266;
  assign \new_[21783]_  = A236 & \new_[21782]_ ;
  assign \new_[21784]_  = \new_[21783]_  & \new_[21778]_ ;
  assign \new_[21787]_  = ~A169 & ~A170;
  assign \new_[21791]_  = A201 & A199;
  assign \new_[21792]_  = ~A168 & \new_[21791]_ ;
  assign \new_[21793]_  = \new_[21792]_  & \new_[21787]_ ;
  assign \new_[21796]_  = ~A233 & A232;
  assign \new_[21800]_  = A300 & A299;
  assign \new_[21801]_  = A236 & \new_[21800]_ ;
  assign \new_[21802]_  = \new_[21801]_  & \new_[21796]_ ;
  assign \new_[21805]_  = ~A169 & ~A170;
  assign \new_[21809]_  = A201 & A199;
  assign \new_[21810]_  = ~A168 & \new_[21809]_ ;
  assign \new_[21811]_  = \new_[21810]_  & \new_[21805]_ ;
  assign \new_[21814]_  = ~A233 & A232;
  assign \new_[21818]_  = A300 & A298;
  assign \new_[21819]_  = A236 & \new_[21818]_ ;
  assign \new_[21820]_  = \new_[21819]_  & \new_[21814]_ ;
  assign \new_[21823]_  = ~A169 & ~A170;
  assign \new_[21827]_  = A201 & A199;
  assign \new_[21828]_  = ~A168 & \new_[21827]_ ;
  assign \new_[21829]_  = \new_[21828]_  & \new_[21823]_ ;
  assign \new_[21832]_  = ~A233 & A232;
  assign \new_[21836]_  = A267 & A265;
  assign \new_[21837]_  = A236 & \new_[21836]_ ;
  assign \new_[21838]_  = \new_[21837]_  & \new_[21832]_ ;
  assign \new_[21841]_  = ~A169 & ~A170;
  assign \new_[21845]_  = A201 & A199;
  assign \new_[21846]_  = ~A168 & \new_[21845]_ ;
  assign \new_[21847]_  = \new_[21846]_  & \new_[21841]_ ;
  assign \new_[21850]_  = ~A233 & A232;
  assign \new_[21854]_  = A267 & A266;
  assign \new_[21855]_  = A236 & \new_[21854]_ ;
  assign \new_[21856]_  = \new_[21855]_  & \new_[21850]_ ;
  assign \new_[21859]_  = ~A169 & ~A170;
  assign \new_[21863]_  = A201 & A200;
  assign \new_[21864]_  = ~A168 & \new_[21863]_ ;
  assign \new_[21865]_  = \new_[21864]_  & \new_[21859]_ ;
  assign \new_[21868]_  = A234 & A232;
  assign \new_[21872]_  = A302 & ~A299;
  assign \new_[21873]_  = A298 & \new_[21872]_ ;
  assign \new_[21874]_  = \new_[21873]_  & \new_[21868]_ ;
  assign \new_[21877]_  = ~A169 & ~A170;
  assign \new_[21881]_  = A201 & A200;
  assign \new_[21882]_  = ~A168 & \new_[21881]_ ;
  assign \new_[21883]_  = \new_[21882]_  & \new_[21877]_ ;
  assign \new_[21886]_  = A234 & A232;
  assign \new_[21890]_  = A302 & A299;
  assign \new_[21891]_  = ~A298 & \new_[21890]_ ;
  assign \new_[21892]_  = \new_[21891]_  & \new_[21886]_ ;
  assign \new_[21895]_  = ~A169 & ~A170;
  assign \new_[21899]_  = A201 & A200;
  assign \new_[21900]_  = ~A168 & \new_[21899]_ ;
  assign \new_[21901]_  = \new_[21900]_  & \new_[21895]_ ;
  assign \new_[21904]_  = A234 & A232;
  assign \new_[21908]_  = A269 & A266;
  assign \new_[21909]_  = ~A265 & \new_[21908]_ ;
  assign \new_[21910]_  = \new_[21909]_  & \new_[21904]_ ;
  assign \new_[21913]_  = ~A169 & ~A170;
  assign \new_[21917]_  = A201 & A200;
  assign \new_[21918]_  = ~A168 & \new_[21917]_ ;
  assign \new_[21919]_  = \new_[21918]_  & \new_[21913]_ ;
  assign \new_[21922]_  = A234 & A232;
  assign \new_[21926]_  = A269 & ~A266;
  assign \new_[21927]_  = A265 & \new_[21926]_ ;
  assign \new_[21928]_  = \new_[21927]_  & \new_[21922]_ ;
  assign \new_[21931]_  = ~A169 & ~A170;
  assign \new_[21935]_  = A201 & A200;
  assign \new_[21936]_  = ~A168 & \new_[21935]_ ;
  assign \new_[21937]_  = \new_[21936]_  & \new_[21931]_ ;
  assign \new_[21940]_  = A234 & A233;
  assign \new_[21944]_  = A302 & ~A299;
  assign \new_[21945]_  = A298 & \new_[21944]_ ;
  assign \new_[21946]_  = \new_[21945]_  & \new_[21940]_ ;
  assign \new_[21949]_  = ~A169 & ~A170;
  assign \new_[21953]_  = A201 & A200;
  assign \new_[21954]_  = ~A168 & \new_[21953]_ ;
  assign \new_[21955]_  = \new_[21954]_  & \new_[21949]_ ;
  assign \new_[21958]_  = A234 & A233;
  assign \new_[21962]_  = A302 & A299;
  assign \new_[21963]_  = ~A298 & \new_[21962]_ ;
  assign \new_[21964]_  = \new_[21963]_  & \new_[21958]_ ;
  assign \new_[21967]_  = ~A169 & ~A170;
  assign \new_[21971]_  = A201 & A200;
  assign \new_[21972]_  = ~A168 & \new_[21971]_ ;
  assign \new_[21973]_  = \new_[21972]_  & \new_[21967]_ ;
  assign \new_[21976]_  = A234 & A233;
  assign \new_[21980]_  = A269 & A266;
  assign \new_[21981]_  = ~A265 & \new_[21980]_ ;
  assign \new_[21982]_  = \new_[21981]_  & \new_[21976]_ ;
  assign \new_[21985]_  = ~A169 & ~A170;
  assign \new_[21989]_  = A201 & A200;
  assign \new_[21990]_  = ~A168 & \new_[21989]_ ;
  assign \new_[21991]_  = \new_[21990]_  & \new_[21985]_ ;
  assign \new_[21994]_  = A234 & A233;
  assign \new_[21998]_  = A269 & ~A266;
  assign \new_[21999]_  = A265 & \new_[21998]_ ;
  assign \new_[22000]_  = \new_[21999]_  & \new_[21994]_ ;
  assign \new_[22003]_  = ~A169 & ~A170;
  assign \new_[22007]_  = A201 & A200;
  assign \new_[22008]_  = ~A168 & \new_[22007]_ ;
  assign \new_[22009]_  = \new_[22008]_  & \new_[22003]_ ;
  assign \new_[22012]_  = A233 & ~A232;
  assign \new_[22016]_  = A300 & A299;
  assign \new_[22017]_  = A236 & \new_[22016]_ ;
  assign \new_[22018]_  = \new_[22017]_  & \new_[22012]_ ;
  assign \new_[22021]_  = ~A169 & ~A170;
  assign \new_[22025]_  = A201 & A200;
  assign \new_[22026]_  = ~A168 & \new_[22025]_ ;
  assign \new_[22027]_  = \new_[22026]_  & \new_[22021]_ ;
  assign \new_[22030]_  = A233 & ~A232;
  assign \new_[22034]_  = A300 & A298;
  assign \new_[22035]_  = A236 & \new_[22034]_ ;
  assign \new_[22036]_  = \new_[22035]_  & \new_[22030]_ ;
  assign \new_[22039]_  = ~A169 & ~A170;
  assign \new_[22043]_  = A201 & A200;
  assign \new_[22044]_  = ~A168 & \new_[22043]_ ;
  assign \new_[22045]_  = \new_[22044]_  & \new_[22039]_ ;
  assign \new_[22048]_  = A233 & ~A232;
  assign \new_[22052]_  = A267 & A265;
  assign \new_[22053]_  = A236 & \new_[22052]_ ;
  assign \new_[22054]_  = \new_[22053]_  & \new_[22048]_ ;
  assign \new_[22057]_  = ~A169 & ~A170;
  assign \new_[22061]_  = A201 & A200;
  assign \new_[22062]_  = ~A168 & \new_[22061]_ ;
  assign \new_[22063]_  = \new_[22062]_  & \new_[22057]_ ;
  assign \new_[22066]_  = A233 & ~A232;
  assign \new_[22070]_  = A267 & A266;
  assign \new_[22071]_  = A236 & \new_[22070]_ ;
  assign \new_[22072]_  = \new_[22071]_  & \new_[22066]_ ;
  assign \new_[22075]_  = ~A169 & ~A170;
  assign \new_[22079]_  = A201 & A200;
  assign \new_[22080]_  = ~A168 & \new_[22079]_ ;
  assign \new_[22081]_  = \new_[22080]_  & \new_[22075]_ ;
  assign \new_[22084]_  = ~A233 & A232;
  assign \new_[22088]_  = A300 & A299;
  assign \new_[22089]_  = A236 & \new_[22088]_ ;
  assign \new_[22090]_  = \new_[22089]_  & \new_[22084]_ ;
  assign \new_[22093]_  = ~A169 & ~A170;
  assign \new_[22097]_  = A201 & A200;
  assign \new_[22098]_  = ~A168 & \new_[22097]_ ;
  assign \new_[22099]_  = \new_[22098]_  & \new_[22093]_ ;
  assign \new_[22102]_  = ~A233 & A232;
  assign \new_[22106]_  = A300 & A298;
  assign \new_[22107]_  = A236 & \new_[22106]_ ;
  assign \new_[22108]_  = \new_[22107]_  & \new_[22102]_ ;
  assign \new_[22111]_  = ~A169 & ~A170;
  assign \new_[22115]_  = A201 & A200;
  assign \new_[22116]_  = ~A168 & \new_[22115]_ ;
  assign \new_[22117]_  = \new_[22116]_  & \new_[22111]_ ;
  assign \new_[22120]_  = ~A233 & A232;
  assign \new_[22124]_  = A267 & A265;
  assign \new_[22125]_  = A236 & \new_[22124]_ ;
  assign \new_[22126]_  = \new_[22125]_  & \new_[22120]_ ;
  assign \new_[22129]_  = ~A169 & ~A170;
  assign \new_[22133]_  = A201 & A200;
  assign \new_[22134]_  = ~A168 & \new_[22133]_ ;
  assign \new_[22135]_  = \new_[22134]_  & \new_[22129]_ ;
  assign \new_[22138]_  = ~A233 & A232;
  assign \new_[22142]_  = A267 & A266;
  assign \new_[22143]_  = A236 & \new_[22142]_ ;
  assign \new_[22144]_  = \new_[22143]_  & \new_[22138]_ ;
  assign \new_[22147]_  = ~A169 & ~A170;
  assign \new_[22151]_  = A200 & ~A199;
  assign \new_[22152]_  = ~A168 & \new_[22151]_ ;
  assign \new_[22153]_  = \new_[22152]_  & \new_[22147]_ ;
  assign \new_[22156]_  = A235 & A203;
  assign \new_[22160]_  = A302 & ~A299;
  assign \new_[22161]_  = A298 & \new_[22160]_ ;
  assign \new_[22162]_  = \new_[22161]_  & \new_[22156]_ ;
  assign \new_[22165]_  = ~A169 & ~A170;
  assign \new_[22169]_  = A200 & ~A199;
  assign \new_[22170]_  = ~A168 & \new_[22169]_ ;
  assign \new_[22171]_  = \new_[22170]_  & \new_[22165]_ ;
  assign \new_[22174]_  = A235 & A203;
  assign \new_[22178]_  = A302 & A299;
  assign \new_[22179]_  = ~A298 & \new_[22178]_ ;
  assign \new_[22180]_  = \new_[22179]_  & \new_[22174]_ ;
  assign \new_[22183]_  = ~A169 & ~A170;
  assign \new_[22187]_  = A200 & ~A199;
  assign \new_[22188]_  = ~A168 & \new_[22187]_ ;
  assign \new_[22189]_  = \new_[22188]_  & \new_[22183]_ ;
  assign \new_[22192]_  = A235 & A203;
  assign \new_[22196]_  = A269 & A266;
  assign \new_[22197]_  = ~A265 & \new_[22196]_ ;
  assign \new_[22198]_  = \new_[22197]_  & \new_[22192]_ ;
  assign \new_[22201]_  = ~A169 & ~A170;
  assign \new_[22205]_  = A200 & ~A199;
  assign \new_[22206]_  = ~A168 & \new_[22205]_ ;
  assign \new_[22207]_  = \new_[22206]_  & \new_[22201]_ ;
  assign \new_[22210]_  = A235 & A203;
  assign \new_[22214]_  = A269 & ~A266;
  assign \new_[22215]_  = A265 & \new_[22214]_ ;
  assign \new_[22216]_  = \new_[22215]_  & \new_[22210]_ ;
  assign \new_[22219]_  = ~A169 & ~A170;
  assign \new_[22223]_  = A200 & ~A199;
  assign \new_[22224]_  = ~A168 & \new_[22223]_ ;
  assign \new_[22225]_  = \new_[22224]_  & \new_[22219]_ ;
  assign \new_[22228]_  = A232 & A203;
  assign \new_[22232]_  = A300 & A299;
  assign \new_[22233]_  = A234 & \new_[22232]_ ;
  assign \new_[22234]_  = \new_[22233]_  & \new_[22228]_ ;
  assign \new_[22237]_  = ~A169 & ~A170;
  assign \new_[22241]_  = A200 & ~A199;
  assign \new_[22242]_  = ~A168 & \new_[22241]_ ;
  assign \new_[22243]_  = \new_[22242]_  & \new_[22237]_ ;
  assign \new_[22246]_  = A232 & A203;
  assign \new_[22250]_  = A300 & A298;
  assign \new_[22251]_  = A234 & \new_[22250]_ ;
  assign \new_[22252]_  = \new_[22251]_  & \new_[22246]_ ;
  assign \new_[22255]_  = ~A169 & ~A170;
  assign \new_[22259]_  = A200 & ~A199;
  assign \new_[22260]_  = ~A168 & \new_[22259]_ ;
  assign \new_[22261]_  = \new_[22260]_  & \new_[22255]_ ;
  assign \new_[22264]_  = A232 & A203;
  assign \new_[22268]_  = A267 & A265;
  assign \new_[22269]_  = A234 & \new_[22268]_ ;
  assign \new_[22270]_  = \new_[22269]_  & \new_[22264]_ ;
  assign \new_[22273]_  = ~A169 & ~A170;
  assign \new_[22277]_  = A200 & ~A199;
  assign \new_[22278]_  = ~A168 & \new_[22277]_ ;
  assign \new_[22279]_  = \new_[22278]_  & \new_[22273]_ ;
  assign \new_[22282]_  = A232 & A203;
  assign \new_[22286]_  = A267 & A266;
  assign \new_[22287]_  = A234 & \new_[22286]_ ;
  assign \new_[22288]_  = \new_[22287]_  & \new_[22282]_ ;
  assign \new_[22291]_  = ~A169 & ~A170;
  assign \new_[22295]_  = A200 & ~A199;
  assign \new_[22296]_  = ~A168 & \new_[22295]_ ;
  assign \new_[22297]_  = \new_[22296]_  & \new_[22291]_ ;
  assign \new_[22300]_  = A233 & A203;
  assign \new_[22304]_  = A300 & A299;
  assign \new_[22305]_  = A234 & \new_[22304]_ ;
  assign \new_[22306]_  = \new_[22305]_  & \new_[22300]_ ;
  assign \new_[22309]_  = ~A169 & ~A170;
  assign \new_[22313]_  = A200 & ~A199;
  assign \new_[22314]_  = ~A168 & \new_[22313]_ ;
  assign \new_[22315]_  = \new_[22314]_  & \new_[22309]_ ;
  assign \new_[22318]_  = A233 & A203;
  assign \new_[22322]_  = A300 & A298;
  assign \new_[22323]_  = A234 & \new_[22322]_ ;
  assign \new_[22324]_  = \new_[22323]_  & \new_[22318]_ ;
  assign \new_[22327]_  = ~A169 & ~A170;
  assign \new_[22331]_  = A200 & ~A199;
  assign \new_[22332]_  = ~A168 & \new_[22331]_ ;
  assign \new_[22333]_  = \new_[22332]_  & \new_[22327]_ ;
  assign \new_[22336]_  = A233 & A203;
  assign \new_[22340]_  = A267 & A265;
  assign \new_[22341]_  = A234 & \new_[22340]_ ;
  assign \new_[22342]_  = \new_[22341]_  & \new_[22336]_ ;
  assign \new_[22345]_  = ~A169 & ~A170;
  assign \new_[22349]_  = A200 & ~A199;
  assign \new_[22350]_  = ~A168 & \new_[22349]_ ;
  assign \new_[22351]_  = \new_[22350]_  & \new_[22345]_ ;
  assign \new_[22354]_  = A233 & A203;
  assign \new_[22358]_  = A267 & A266;
  assign \new_[22359]_  = A234 & \new_[22358]_ ;
  assign \new_[22360]_  = \new_[22359]_  & \new_[22354]_ ;
  assign \new_[22363]_  = ~A169 & ~A170;
  assign \new_[22367]_  = A200 & ~A199;
  assign \new_[22368]_  = ~A168 & \new_[22367]_ ;
  assign \new_[22369]_  = \new_[22368]_  & \new_[22363]_ ;
  assign \new_[22372]_  = ~A232 & A203;
  assign \new_[22376]_  = A301 & A236;
  assign \new_[22377]_  = A233 & \new_[22376]_ ;
  assign \new_[22378]_  = \new_[22377]_  & \new_[22372]_ ;
  assign \new_[22381]_  = ~A169 & ~A170;
  assign \new_[22385]_  = A200 & ~A199;
  assign \new_[22386]_  = ~A168 & \new_[22385]_ ;
  assign \new_[22387]_  = \new_[22386]_  & \new_[22381]_ ;
  assign \new_[22390]_  = ~A232 & A203;
  assign \new_[22394]_  = A268 & A236;
  assign \new_[22395]_  = A233 & \new_[22394]_ ;
  assign \new_[22396]_  = \new_[22395]_  & \new_[22390]_ ;
  assign \new_[22399]_  = ~A169 & ~A170;
  assign \new_[22403]_  = A200 & ~A199;
  assign \new_[22404]_  = ~A168 & \new_[22403]_ ;
  assign \new_[22405]_  = \new_[22404]_  & \new_[22399]_ ;
  assign \new_[22408]_  = A232 & A203;
  assign \new_[22412]_  = A301 & A236;
  assign \new_[22413]_  = ~A233 & \new_[22412]_ ;
  assign \new_[22414]_  = \new_[22413]_  & \new_[22408]_ ;
  assign \new_[22417]_  = ~A169 & ~A170;
  assign \new_[22421]_  = A200 & ~A199;
  assign \new_[22422]_  = ~A168 & \new_[22421]_ ;
  assign \new_[22423]_  = \new_[22422]_  & \new_[22417]_ ;
  assign \new_[22426]_  = A232 & A203;
  assign \new_[22430]_  = A268 & A236;
  assign \new_[22431]_  = ~A233 & \new_[22430]_ ;
  assign \new_[22432]_  = \new_[22431]_  & \new_[22426]_ ;
  assign \new_[22435]_  = ~A169 & ~A170;
  assign \new_[22439]_  = ~A200 & A199;
  assign \new_[22440]_  = ~A168 & \new_[22439]_ ;
  assign \new_[22441]_  = \new_[22440]_  & \new_[22435]_ ;
  assign \new_[22444]_  = A235 & A203;
  assign \new_[22448]_  = A302 & ~A299;
  assign \new_[22449]_  = A298 & \new_[22448]_ ;
  assign \new_[22450]_  = \new_[22449]_  & \new_[22444]_ ;
  assign \new_[22453]_  = ~A169 & ~A170;
  assign \new_[22457]_  = ~A200 & A199;
  assign \new_[22458]_  = ~A168 & \new_[22457]_ ;
  assign \new_[22459]_  = \new_[22458]_  & \new_[22453]_ ;
  assign \new_[22462]_  = A235 & A203;
  assign \new_[22466]_  = A302 & A299;
  assign \new_[22467]_  = ~A298 & \new_[22466]_ ;
  assign \new_[22468]_  = \new_[22467]_  & \new_[22462]_ ;
  assign \new_[22471]_  = ~A169 & ~A170;
  assign \new_[22475]_  = ~A200 & A199;
  assign \new_[22476]_  = ~A168 & \new_[22475]_ ;
  assign \new_[22477]_  = \new_[22476]_  & \new_[22471]_ ;
  assign \new_[22480]_  = A235 & A203;
  assign \new_[22484]_  = A269 & A266;
  assign \new_[22485]_  = ~A265 & \new_[22484]_ ;
  assign \new_[22486]_  = \new_[22485]_  & \new_[22480]_ ;
  assign \new_[22489]_  = ~A169 & ~A170;
  assign \new_[22493]_  = ~A200 & A199;
  assign \new_[22494]_  = ~A168 & \new_[22493]_ ;
  assign \new_[22495]_  = \new_[22494]_  & \new_[22489]_ ;
  assign \new_[22498]_  = A235 & A203;
  assign \new_[22502]_  = A269 & ~A266;
  assign \new_[22503]_  = A265 & \new_[22502]_ ;
  assign \new_[22504]_  = \new_[22503]_  & \new_[22498]_ ;
  assign \new_[22507]_  = ~A169 & ~A170;
  assign \new_[22511]_  = ~A200 & A199;
  assign \new_[22512]_  = ~A168 & \new_[22511]_ ;
  assign \new_[22513]_  = \new_[22512]_  & \new_[22507]_ ;
  assign \new_[22516]_  = A232 & A203;
  assign \new_[22520]_  = A300 & A299;
  assign \new_[22521]_  = A234 & \new_[22520]_ ;
  assign \new_[22522]_  = \new_[22521]_  & \new_[22516]_ ;
  assign \new_[22525]_  = ~A169 & ~A170;
  assign \new_[22529]_  = ~A200 & A199;
  assign \new_[22530]_  = ~A168 & \new_[22529]_ ;
  assign \new_[22531]_  = \new_[22530]_  & \new_[22525]_ ;
  assign \new_[22534]_  = A232 & A203;
  assign \new_[22538]_  = A300 & A298;
  assign \new_[22539]_  = A234 & \new_[22538]_ ;
  assign \new_[22540]_  = \new_[22539]_  & \new_[22534]_ ;
  assign \new_[22543]_  = ~A169 & ~A170;
  assign \new_[22547]_  = ~A200 & A199;
  assign \new_[22548]_  = ~A168 & \new_[22547]_ ;
  assign \new_[22549]_  = \new_[22548]_  & \new_[22543]_ ;
  assign \new_[22552]_  = A232 & A203;
  assign \new_[22556]_  = A267 & A265;
  assign \new_[22557]_  = A234 & \new_[22556]_ ;
  assign \new_[22558]_  = \new_[22557]_  & \new_[22552]_ ;
  assign \new_[22561]_  = ~A169 & ~A170;
  assign \new_[22565]_  = ~A200 & A199;
  assign \new_[22566]_  = ~A168 & \new_[22565]_ ;
  assign \new_[22567]_  = \new_[22566]_  & \new_[22561]_ ;
  assign \new_[22570]_  = A232 & A203;
  assign \new_[22574]_  = A267 & A266;
  assign \new_[22575]_  = A234 & \new_[22574]_ ;
  assign \new_[22576]_  = \new_[22575]_  & \new_[22570]_ ;
  assign \new_[22579]_  = ~A169 & ~A170;
  assign \new_[22583]_  = ~A200 & A199;
  assign \new_[22584]_  = ~A168 & \new_[22583]_ ;
  assign \new_[22585]_  = \new_[22584]_  & \new_[22579]_ ;
  assign \new_[22588]_  = A233 & A203;
  assign \new_[22592]_  = A300 & A299;
  assign \new_[22593]_  = A234 & \new_[22592]_ ;
  assign \new_[22594]_  = \new_[22593]_  & \new_[22588]_ ;
  assign \new_[22597]_  = ~A169 & ~A170;
  assign \new_[22601]_  = ~A200 & A199;
  assign \new_[22602]_  = ~A168 & \new_[22601]_ ;
  assign \new_[22603]_  = \new_[22602]_  & \new_[22597]_ ;
  assign \new_[22606]_  = A233 & A203;
  assign \new_[22610]_  = A300 & A298;
  assign \new_[22611]_  = A234 & \new_[22610]_ ;
  assign \new_[22612]_  = \new_[22611]_  & \new_[22606]_ ;
  assign \new_[22615]_  = ~A169 & ~A170;
  assign \new_[22619]_  = ~A200 & A199;
  assign \new_[22620]_  = ~A168 & \new_[22619]_ ;
  assign \new_[22621]_  = \new_[22620]_  & \new_[22615]_ ;
  assign \new_[22624]_  = A233 & A203;
  assign \new_[22628]_  = A267 & A265;
  assign \new_[22629]_  = A234 & \new_[22628]_ ;
  assign \new_[22630]_  = \new_[22629]_  & \new_[22624]_ ;
  assign \new_[22633]_  = ~A169 & ~A170;
  assign \new_[22637]_  = ~A200 & A199;
  assign \new_[22638]_  = ~A168 & \new_[22637]_ ;
  assign \new_[22639]_  = \new_[22638]_  & \new_[22633]_ ;
  assign \new_[22642]_  = A233 & A203;
  assign \new_[22646]_  = A267 & A266;
  assign \new_[22647]_  = A234 & \new_[22646]_ ;
  assign \new_[22648]_  = \new_[22647]_  & \new_[22642]_ ;
  assign \new_[22651]_  = ~A169 & ~A170;
  assign \new_[22655]_  = ~A200 & A199;
  assign \new_[22656]_  = ~A168 & \new_[22655]_ ;
  assign \new_[22657]_  = \new_[22656]_  & \new_[22651]_ ;
  assign \new_[22660]_  = ~A232 & A203;
  assign \new_[22664]_  = A301 & A236;
  assign \new_[22665]_  = A233 & \new_[22664]_ ;
  assign \new_[22666]_  = \new_[22665]_  & \new_[22660]_ ;
  assign \new_[22669]_  = ~A169 & ~A170;
  assign \new_[22673]_  = ~A200 & A199;
  assign \new_[22674]_  = ~A168 & \new_[22673]_ ;
  assign \new_[22675]_  = \new_[22674]_  & \new_[22669]_ ;
  assign \new_[22678]_  = ~A232 & A203;
  assign \new_[22682]_  = A268 & A236;
  assign \new_[22683]_  = A233 & \new_[22682]_ ;
  assign \new_[22684]_  = \new_[22683]_  & \new_[22678]_ ;
  assign \new_[22687]_  = ~A169 & ~A170;
  assign \new_[22691]_  = ~A200 & A199;
  assign \new_[22692]_  = ~A168 & \new_[22691]_ ;
  assign \new_[22693]_  = \new_[22692]_  & \new_[22687]_ ;
  assign \new_[22696]_  = A232 & A203;
  assign \new_[22700]_  = A301 & A236;
  assign \new_[22701]_  = ~A233 & \new_[22700]_ ;
  assign \new_[22702]_  = \new_[22701]_  & \new_[22696]_ ;
  assign \new_[22705]_  = ~A169 & ~A170;
  assign \new_[22709]_  = ~A200 & A199;
  assign \new_[22710]_  = ~A168 & \new_[22709]_ ;
  assign \new_[22711]_  = \new_[22710]_  & \new_[22705]_ ;
  assign \new_[22714]_  = A232 & A203;
  assign \new_[22718]_  = A268 & A236;
  assign \new_[22719]_  = ~A233 & \new_[22718]_ ;
  assign \new_[22720]_  = \new_[22719]_  & \new_[22714]_ ;
  assign \new_[22723]_  = A166 & A168;
  assign \new_[22727]_  = ~A203 & ~A202;
  assign \new_[22728]_  = ~A201 & \new_[22727]_ ;
  assign \new_[22729]_  = \new_[22728]_  & \new_[22723]_ ;
  assign \new_[22733]_  = A236 & A233;
  assign \new_[22734]_  = ~A232 & \new_[22733]_ ;
  assign \new_[22738]_  = A302 & ~A299;
  assign \new_[22739]_  = A298 & \new_[22738]_ ;
  assign \new_[22740]_  = \new_[22739]_  & \new_[22734]_ ;
  assign \new_[22743]_  = A166 & A168;
  assign \new_[22747]_  = ~A203 & ~A202;
  assign \new_[22748]_  = ~A201 & \new_[22747]_ ;
  assign \new_[22749]_  = \new_[22748]_  & \new_[22743]_ ;
  assign \new_[22753]_  = A236 & A233;
  assign \new_[22754]_  = ~A232 & \new_[22753]_ ;
  assign \new_[22758]_  = A302 & A299;
  assign \new_[22759]_  = ~A298 & \new_[22758]_ ;
  assign \new_[22760]_  = \new_[22759]_  & \new_[22754]_ ;
  assign \new_[22763]_  = A166 & A168;
  assign \new_[22767]_  = ~A203 & ~A202;
  assign \new_[22768]_  = ~A201 & \new_[22767]_ ;
  assign \new_[22769]_  = \new_[22768]_  & \new_[22763]_ ;
  assign \new_[22773]_  = A236 & A233;
  assign \new_[22774]_  = ~A232 & \new_[22773]_ ;
  assign \new_[22778]_  = A269 & A266;
  assign \new_[22779]_  = ~A265 & \new_[22778]_ ;
  assign \new_[22780]_  = \new_[22779]_  & \new_[22774]_ ;
  assign \new_[22783]_  = A166 & A168;
  assign \new_[22787]_  = ~A203 & ~A202;
  assign \new_[22788]_  = ~A201 & \new_[22787]_ ;
  assign \new_[22789]_  = \new_[22788]_  & \new_[22783]_ ;
  assign \new_[22793]_  = A236 & A233;
  assign \new_[22794]_  = ~A232 & \new_[22793]_ ;
  assign \new_[22798]_  = A269 & ~A266;
  assign \new_[22799]_  = A265 & \new_[22798]_ ;
  assign \new_[22800]_  = \new_[22799]_  & \new_[22794]_ ;
  assign \new_[22803]_  = A166 & A168;
  assign \new_[22807]_  = ~A203 & ~A202;
  assign \new_[22808]_  = ~A201 & \new_[22807]_ ;
  assign \new_[22809]_  = \new_[22808]_  & \new_[22803]_ ;
  assign \new_[22813]_  = A236 & ~A233;
  assign \new_[22814]_  = A232 & \new_[22813]_ ;
  assign \new_[22818]_  = A302 & ~A299;
  assign \new_[22819]_  = A298 & \new_[22818]_ ;
  assign \new_[22820]_  = \new_[22819]_  & \new_[22814]_ ;
  assign \new_[22823]_  = A166 & A168;
  assign \new_[22827]_  = ~A203 & ~A202;
  assign \new_[22828]_  = ~A201 & \new_[22827]_ ;
  assign \new_[22829]_  = \new_[22828]_  & \new_[22823]_ ;
  assign \new_[22833]_  = A236 & ~A233;
  assign \new_[22834]_  = A232 & \new_[22833]_ ;
  assign \new_[22838]_  = A302 & A299;
  assign \new_[22839]_  = ~A298 & \new_[22838]_ ;
  assign \new_[22840]_  = \new_[22839]_  & \new_[22834]_ ;
  assign \new_[22843]_  = A166 & A168;
  assign \new_[22847]_  = ~A203 & ~A202;
  assign \new_[22848]_  = ~A201 & \new_[22847]_ ;
  assign \new_[22849]_  = \new_[22848]_  & \new_[22843]_ ;
  assign \new_[22853]_  = A236 & ~A233;
  assign \new_[22854]_  = A232 & \new_[22853]_ ;
  assign \new_[22858]_  = A269 & A266;
  assign \new_[22859]_  = ~A265 & \new_[22858]_ ;
  assign \new_[22860]_  = \new_[22859]_  & \new_[22854]_ ;
  assign \new_[22863]_  = A166 & A168;
  assign \new_[22867]_  = ~A203 & ~A202;
  assign \new_[22868]_  = ~A201 & \new_[22867]_ ;
  assign \new_[22869]_  = \new_[22868]_  & \new_[22863]_ ;
  assign \new_[22873]_  = A236 & ~A233;
  assign \new_[22874]_  = A232 & \new_[22873]_ ;
  assign \new_[22878]_  = A269 & ~A266;
  assign \new_[22879]_  = A265 & \new_[22878]_ ;
  assign \new_[22880]_  = \new_[22879]_  & \new_[22874]_ ;
  assign \new_[22883]_  = A166 & A168;
  assign \new_[22887]_  = ~A201 & A200;
  assign \new_[22888]_  = A199 & \new_[22887]_ ;
  assign \new_[22889]_  = \new_[22888]_  & \new_[22883]_ ;
  assign \new_[22893]_  = A234 & A232;
  assign \new_[22894]_  = ~A202 & \new_[22893]_ ;
  assign \new_[22898]_  = A302 & ~A299;
  assign \new_[22899]_  = A298 & \new_[22898]_ ;
  assign \new_[22900]_  = \new_[22899]_  & \new_[22894]_ ;
  assign \new_[22903]_  = A166 & A168;
  assign \new_[22907]_  = ~A201 & A200;
  assign \new_[22908]_  = A199 & \new_[22907]_ ;
  assign \new_[22909]_  = \new_[22908]_  & \new_[22903]_ ;
  assign \new_[22913]_  = A234 & A232;
  assign \new_[22914]_  = ~A202 & \new_[22913]_ ;
  assign \new_[22918]_  = A302 & A299;
  assign \new_[22919]_  = ~A298 & \new_[22918]_ ;
  assign \new_[22920]_  = \new_[22919]_  & \new_[22914]_ ;
  assign \new_[22923]_  = A166 & A168;
  assign \new_[22927]_  = ~A201 & A200;
  assign \new_[22928]_  = A199 & \new_[22927]_ ;
  assign \new_[22929]_  = \new_[22928]_  & \new_[22923]_ ;
  assign \new_[22933]_  = A234 & A232;
  assign \new_[22934]_  = ~A202 & \new_[22933]_ ;
  assign \new_[22938]_  = A269 & A266;
  assign \new_[22939]_  = ~A265 & \new_[22938]_ ;
  assign \new_[22940]_  = \new_[22939]_  & \new_[22934]_ ;
  assign \new_[22943]_  = A166 & A168;
  assign \new_[22947]_  = ~A201 & A200;
  assign \new_[22948]_  = A199 & \new_[22947]_ ;
  assign \new_[22949]_  = \new_[22948]_  & \new_[22943]_ ;
  assign \new_[22953]_  = A234 & A232;
  assign \new_[22954]_  = ~A202 & \new_[22953]_ ;
  assign \new_[22958]_  = A269 & ~A266;
  assign \new_[22959]_  = A265 & \new_[22958]_ ;
  assign \new_[22960]_  = \new_[22959]_  & \new_[22954]_ ;
  assign \new_[22963]_  = A166 & A168;
  assign \new_[22967]_  = ~A201 & A200;
  assign \new_[22968]_  = A199 & \new_[22967]_ ;
  assign \new_[22969]_  = \new_[22968]_  & \new_[22963]_ ;
  assign \new_[22973]_  = A234 & A233;
  assign \new_[22974]_  = ~A202 & \new_[22973]_ ;
  assign \new_[22978]_  = A302 & ~A299;
  assign \new_[22979]_  = A298 & \new_[22978]_ ;
  assign \new_[22980]_  = \new_[22979]_  & \new_[22974]_ ;
  assign \new_[22983]_  = A166 & A168;
  assign \new_[22987]_  = ~A201 & A200;
  assign \new_[22988]_  = A199 & \new_[22987]_ ;
  assign \new_[22989]_  = \new_[22988]_  & \new_[22983]_ ;
  assign \new_[22993]_  = A234 & A233;
  assign \new_[22994]_  = ~A202 & \new_[22993]_ ;
  assign \new_[22998]_  = A302 & A299;
  assign \new_[22999]_  = ~A298 & \new_[22998]_ ;
  assign \new_[23000]_  = \new_[22999]_  & \new_[22994]_ ;
  assign \new_[23003]_  = A166 & A168;
  assign \new_[23007]_  = ~A201 & A200;
  assign \new_[23008]_  = A199 & \new_[23007]_ ;
  assign \new_[23009]_  = \new_[23008]_  & \new_[23003]_ ;
  assign \new_[23013]_  = A234 & A233;
  assign \new_[23014]_  = ~A202 & \new_[23013]_ ;
  assign \new_[23018]_  = A269 & A266;
  assign \new_[23019]_  = ~A265 & \new_[23018]_ ;
  assign \new_[23020]_  = \new_[23019]_  & \new_[23014]_ ;
  assign \new_[23023]_  = A166 & A168;
  assign \new_[23027]_  = ~A201 & A200;
  assign \new_[23028]_  = A199 & \new_[23027]_ ;
  assign \new_[23029]_  = \new_[23028]_  & \new_[23023]_ ;
  assign \new_[23033]_  = A234 & A233;
  assign \new_[23034]_  = ~A202 & \new_[23033]_ ;
  assign \new_[23038]_  = A269 & ~A266;
  assign \new_[23039]_  = A265 & \new_[23038]_ ;
  assign \new_[23040]_  = \new_[23039]_  & \new_[23034]_ ;
  assign \new_[23043]_  = A166 & A168;
  assign \new_[23047]_  = ~A201 & A200;
  assign \new_[23048]_  = A199 & \new_[23047]_ ;
  assign \new_[23049]_  = \new_[23048]_  & \new_[23043]_ ;
  assign \new_[23053]_  = A233 & ~A232;
  assign \new_[23054]_  = ~A202 & \new_[23053]_ ;
  assign \new_[23058]_  = A300 & A299;
  assign \new_[23059]_  = A236 & \new_[23058]_ ;
  assign \new_[23060]_  = \new_[23059]_  & \new_[23054]_ ;
  assign \new_[23063]_  = A166 & A168;
  assign \new_[23067]_  = ~A201 & A200;
  assign \new_[23068]_  = A199 & \new_[23067]_ ;
  assign \new_[23069]_  = \new_[23068]_  & \new_[23063]_ ;
  assign \new_[23073]_  = A233 & ~A232;
  assign \new_[23074]_  = ~A202 & \new_[23073]_ ;
  assign \new_[23078]_  = A300 & A298;
  assign \new_[23079]_  = A236 & \new_[23078]_ ;
  assign \new_[23080]_  = \new_[23079]_  & \new_[23074]_ ;
  assign \new_[23083]_  = A166 & A168;
  assign \new_[23087]_  = ~A201 & A200;
  assign \new_[23088]_  = A199 & \new_[23087]_ ;
  assign \new_[23089]_  = \new_[23088]_  & \new_[23083]_ ;
  assign \new_[23093]_  = A233 & ~A232;
  assign \new_[23094]_  = ~A202 & \new_[23093]_ ;
  assign \new_[23098]_  = A267 & A265;
  assign \new_[23099]_  = A236 & \new_[23098]_ ;
  assign \new_[23100]_  = \new_[23099]_  & \new_[23094]_ ;
  assign \new_[23103]_  = A166 & A168;
  assign \new_[23107]_  = ~A201 & A200;
  assign \new_[23108]_  = A199 & \new_[23107]_ ;
  assign \new_[23109]_  = \new_[23108]_  & \new_[23103]_ ;
  assign \new_[23113]_  = A233 & ~A232;
  assign \new_[23114]_  = ~A202 & \new_[23113]_ ;
  assign \new_[23118]_  = A267 & A266;
  assign \new_[23119]_  = A236 & \new_[23118]_ ;
  assign \new_[23120]_  = \new_[23119]_  & \new_[23114]_ ;
  assign \new_[23123]_  = A166 & A168;
  assign \new_[23127]_  = ~A201 & A200;
  assign \new_[23128]_  = A199 & \new_[23127]_ ;
  assign \new_[23129]_  = \new_[23128]_  & \new_[23123]_ ;
  assign \new_[23133]_  = ~A233 & A232;
  assign \new_[23134]_  = ~A202 & \new_[23133]_ ;
  assign \new_[23138]_  = A300 & A299;
  assign \new_[23139]_  = A236 & \new_[23138]_ ;
  assign \new_[23140]_  = \new_[23139]_  & \new_[23134]_ ;
  assign \new_[23143]_  = A166 & A168;
  assign \new_[23147]_  = ~A201 & A200;
  assign \new_[23148]_  = A199 & \new_[23147]_ ;
  assign \new_[23149]_  = \new_[23148]_  & \new_[23143]_ ;
  assign \new_[23153]_  = ~A233 & A232;
  assign \new_[23154]_  = ~A202 & \new_[23153]_ ;
  assign \new_[23158]_  = A300 & A298;
  assign \new_[23159]_  = A236 & \new_[23158]_ ;
  assign \new_[23160]_  = \new_[23159]_  & \new_[23154]_ ;
  assign \new_[23163]_  = A166 & A168;
  assign \new_[23167]_  = ~A201 & A200;
  assign \new_[23168]_  = A199 & \new_[23167]_ ;
  assign \new_[23169]_  = \new_[23168]_  & \new_[23163]_ ;
  assign \new_[23173]_  = ~A233 & A232;
  assign \new_[23174]_  = ~A202 & \new_[23173]_ ;
  assign \new_[23178]_  = A267 & A265;
  assign \new_[23179]_  = A236 & \new_[23178]_ ;
  assign \new_[23180]_  = \new_[23179]_  & \new_[23174]_ ;
  assign \new_[23183]_  = A166 & A168;
  assign \new_[23187]_  = ~A201 & A200;
  assign \new_[23188]_  = A199 & \new_[23187]_ ;
  assign \new_[23189]_  = \new_[23188]_  & \new_[23183]_ ;
  assign \new_[23193]_  = ~A233 & A232;
  assign \new_[23194]_  = ~A202 & \new_[23193]_ ;
  assign \new_[23198]_  = A267 & A266;
  assign \new_[23199]_  = A236 & \new_[23198]_ ;
  assign \new_[23200]_  = \new_[23199]_  & \new_[23194]_ ;
  assign \new_[23203]_  = A166 & A168;
  assign \new_[23207]_  = ~A202 & ~A200;
  assign \new_[23208]_  = ~A199 & \new_[23207]_ ;
  assign \new_[23209]_  = \new_[23208]_  & \new_[23203]_ ;
  assign \new_[23213]_  = A236 & A233;
  assign \new_[23214]_  = ~A232 & \new_[23213]_ ;
  assign \new_[23218]_  = A302 & ~A299;
  assign \new_[23219]_  = A298 & \new_[23218]_ ;
  assign \new_[23220]_  = \new_[23219]_  & \new_[23214]_ ;
  assign \new_[23223]_  = A166 & A168;
  assign \new_[23227]_  = ~A202 & ~A200;
  assign \new_[23228]_  = ~A199 & \new_[23227]_ ;
  assign \new_[23229]_  = \new_[23228]_  & \new_[23223]_ ;
  assign \new_[23233]_  = A236 & A233;
  assign \new_[23234]_  = ~A232 & \new_[23233]_ ;
  assign \new_[23238]_  = A302 & A299;
  assign \new_[23239]_  = ~A298 & \new_[23238]_ ;
  assign \new_[23240]_  = \new_[23239]_  & \new_[23234]_ ;
  assign \new_[23243]_  = A166 & A168;
  assign \new_[23247]_  = ~A202 & ~A200;
  assign \new_[23248]_  = ~A199 & \new_[23247]_ ;
  assign \new_[23249]_  = \new_[23248]_  & \new_[23243]_ ;
  assign \new_[23253]_  = A236 & A233;
  assign \new_[23254]_  = ~A232 & \new_[23253]_ ;
  assign \new_[23258]_  = A269 & A266;
  assign \new_[23259]_  = ~A265 & \new_[23258]_ ;
  assign \new_[23260]_  = \new_[23259]_  & \new_[23254]_ ;
  assign \new_[23263]_  = A166 & A168;
  assign \new_[23267]_  = ~A202 & ~A200;
  assign \new_[23268]_  = ~A199 & \new_[23267]_ ;
  assign \new_[23269]_  = \new_[23268]_  & \new_[23263]_ ;
  assign \new_[23273]_  = A236 & A233;
  assign \new_[23274]_  = ~A232 & \new_[23273]_ ;
  assign \new_[23278]_  = A269 & ~A266;
  assign \new_[23279]_  = A265 & \new_[23278]_ ;
  assign \new_[23280]_  = \new_[23279]_  & \new_[23274]_ ;
  assign \new_[23283]_  = A166 & A168;
  assign \new_[23287]_  = ~A202 & ~A200;
  assign \new_[23288]_  = ~A199 & \new_[23287]_ ;
  assign \new_[23289]_  = \new_[23288]_  & \new_[23283]_ ;
  assign \new_[23293]_  = A236 & ~A233;
  assign \new_[23294]_  = A232 & \new_[23293]_ ;
  assign \new_[23298]_  = A302 & ~A299;
  assign \new_[23299]_  = A298 & \new_[23298]_ ;
  assign \new_[23300]_  = \new_[23299]_  & \new_[23294]_ ;
  assign \new_[23303]_  = A166 & A168;
  assign \new_[23307]_  = ~A202 & ~A200;
  assign \new_[23308]_  = ~A199 & \new_[23307]_ ;
  assign \new_[23309]_  = \new_[23308]_  & \new_[23303]_ ;
  assign \new_[23313]_  = A236 & ~A233;
  assign \new_[23314]_  = A232 & \new_[23313]_ ;
  assign \new_[23318]_  = A302 & A299;
  assign \new_[23319]_  = ~A298 & \new_[23318]_ ;
  assign \new_[23320]_  = \new_[23319]_  & \new_[23314]_ ;
  assign \new_[23323]_  = A166 & A168;
  assign \new_[23327]_  = ~A202 & ~A200;
  assign \new_[23328]_  = ~A199 & \new_[23327]_ ;
  assign \new_[23329]_  = \new_[23328]_  & \new_[23323]_ ;
  assign \new_[23333]_  = A236 & ~A233;
  assign \new_[23334]_  = A232 & \new_[23333]_ ;
  assign \new_[23338]_  = A269 & A266;
  assign \new_[23339]_  = ~A265 & \new_[23338]_ ;
  assign \new_[23340]_  = \new_[23339]_  & \new_[23334]_ ;
  assign \new_[23343]_  = A166 & A168;
  assign \new_[23347]_  = ~A202 & ~A200;
  assign \new_[23348]_  = ~A199 & \new_[23347]_ ;
  assign \new_[23349]_  = \new_[23348]_  & \new_[23343]_ ;
  assign \new_[23353]_  = A236 & ~A233;
  assign \new_[23354]_  = A232 & \new_[23353]_ ;
  assign \new_[23358]_  = A269 & ~A266;
  assign \new_[23359]_  = A265 & \new_[23358]_ ;
  assign \new_[23360]_  = \new_[23359]_  & \new_[23354]_ ;
  assign \new_[23363]_  = A167 & A168;
  assign \new_[23367]_  = ~A203 & ~A202;
  assign \new_[23368]_  = ~A201 & \new_[23367]_ ;
  assign \new_[23369]_  = \new_[23368]_  & \new_[23363]_ ;
  assign \new_[23373]_  = A236 & A233;
  assign \new_[23374]_  = ~A232 & \new_[23373]_ ;
  assign \new_[23378]_  = A302 & ~A299;
  assign \new_[23379]_  = A298 & \new_[23378]_ ;
  assign \new_[23380]_  = \new_[23379]_  & \new_[23374]_ ;
  assign \new_[23383]_  = A167 & A168;
  assign \new_[23387]_  = ~A203 & ~A202;
  assign \new_[23388]_  = ~A201 & \new_[23387]_ ;
  assign \new_[23389]_  = \new_[23388]_  & \new_[23383]_ ;
  assign \new_[23393]_  = A236 & A233;
  assign \new_[23394]_  = ~A232 & \new_[23393]_ ;
  assign \new_[23398]_  = A302 & A299;
  assign \new_[23399]_  = ~A298 & \new_[23398]_ ;
  assign \new_[23400]_  = \new_[23399]_  & \new_[23394]_ ;
  assign \new_[23403]_  = A167 & A168;
  assign \new_[23407]_  = ~A203 & ~A202;
  assign \new_[23408]_  = ~A201 & \new_[23407]_ ;
  assign \new_[23409]_  = \new_[23408]_  & \new_[23403]_ ;
  assign \new_[23413]_  = A236 & A233;
  assign \new_[23414]_  = ~A232 & \new_[23413]_ ;
  assign \new_[23418]_  = A269 & A266;
  assign \new_[23419]_  = ~A265 & \new_[23418]_ ;
  assign \new_[23420]_  = \new_[23419]_  & \new_[23414]_ ;
  assign \new_[23423]_  = A167 & A168;
  assign \new_[23427]_  = ~A203 & ~A202;
  assign \new_[23428]_  = ~A201 & \new_[23427]_ ;
  assign \new_[23429]_  = \new_[23428]_  & \new_[23423]_ ;
  assign \new_[23433]_  = A236 & A233;
  assign \new_[23434]_  = ~A232 & \new_[23433]_ ;
  assign \new_[23438]_  = A269 & ~A266;
  assign \new_[23439]_  = A265 & \new_[23438]_ ;
  assign \new_[23440]_  = \new_[23439]_  & \new_[23434]_ ;
  assign \new_[23443]_  = A167 & A168;
  assign \new_[23447]_  = ~A203 & ~A202;
  assign \new_[23448]_  = ~A201 & \new_[23447]_ ;
  assign \new_[23449]_  = \new_[23448]_  & \new_[23443]_ ;
  assign \new_[23453]_  = A236 & ~A233;
  assign \new_[23454]_  = A232 & \new_[23453]_ ;
  assign \new_[23458]_  = A302 & ~A299;
  assign \new_[23459]_  = A298 & \new_[23458]_ ;
  assign \new_[23460]_  = \new_[23459]_  & \new_[23454]_ ;
  assign \new_[23463]_  = A167 & A168;
  assign \new_[23467]_  = ~A203 & ~A202;
  assign \new_[23468]_  = ~A201 & \new_[23467]_ ;
  assign \new_[23469]_  = \new_[23468]_  & \new_[23463]_ ;
  assign \new_[23473]_  = A236 & ~A233;
  assign \new_[23474]_  = A232 & \new_[23473]_ ;
  assign \new_[23478]_  = A302 & A299;
  assign \new_[23479]_  = ~A298 & \new_[23478]_ ;
  assign \new_[23480]_  = \new_[23479]_  & \new_[23474]_ ;
  assign \new_[23483]_  = A167 & A168;
  assign \new_[23487]_  = ~A203 & ~A202;
  assign \new_[23488]_  = ~A201 & \new_[23487]_ ;
  assign \new_[23489]_  = \new_[23488]_  & \new_[23483]_ ;
  assign \new_[23493]_  = A236 & ~A233;
  assign \new_[23494]_  = A232 & \new_[23493]_ ;
  assign \new_[23498]_  = A269 & A266;
  assign \new_[23499]_  = ~A265 & \new_[23498]_ ;
  assign \new_[23500]_  = \new_[23499]_  & \new_[23494]_ ;
  assign \new_[23503]_  = A167 & A168;
  assign \new_[23507]_  = ~A203 & ~A202;
  assign \new_[23508]_  = ~A201 & \new_[23507]_ ;
  assign \new_[23509]_  = \new_[23508]_  & \new_[23503]_ ;
  assign \new_[23513]_  = A236 & ~A233;
  assign \new_[23514]_  = A232 & \new_[23513]_ ;
  assign \new_[23518]_  = A269 & ~A266;
  assign \new_[23519]_  = A265 & \new_[23518]_ ;
  assign \new_[23520]_  = \new_[23519]_  & \new_[23514]_ ;
  assign \new_[23523]_  = A167 & A168;
  assign \new_[23527]_  = ~A201 & A200;
  assign \new_[23528]_  = A199 & \new_[23527]_ ;
  assign \new_[23529]_  = \new_[23528]_  & \new_[23523]_ ;
  assign \new_[23533]_  = A234 & A232;
  assign \new_[23534]_  = ~A202 & \new_[23533]_ ;
  assign \new_[23538]_  = A302 & ~A299;
  assign \new_[23539]_  = A298 & \new_[23538]_ ;
  assign \new_[23540]_  = \new_[23539]_  & \new_[23534]_ ;
  assign \new_[23543]_  = A167 & A168;
  assign \new_[23547]_  = ~A201 & A200;
  assign \new_[23548]_  = A199 & \new_[23547]_ ;
  assign \new_[23549]_  = \new_[23548]_  & \new_[23543]_ ;
  assign \new_[23553]_  = A234 & A232;
  assign \new_[23554]_  = ~A202 & \new_[23553]_ ;
  assign \new_[23558]_  = A302 & A299;
  assign \new_[23559]_  = ~A298 & \new_[23558]_ ;
  assign \new_[23560]_  = \new_[23559]_  & \new_[23554]_ ;
  assign \new_[23563]_  = A167 & A168;
  assign \new_[23567]_  = ~A201 & A200;
  assign \new_[23568]_  = A199 & \new_[23567]_ ;
  assign \new_[23569]_  = \new_[23568]_  & \new_[23563]_ ;
  assign \new_[23573]_  = A234 & A232;
  assign \new_[23574]_  = ~A202 & \new_[23573]_ ;
  assign \new_[23578]_  = A269 & A266;
  assign \new_[23579]_  = ~A265 & \new_[23578]_ ;
  assign \new_[23580]_  = \new_[23579]_  & \new_[23574]_ ;
  assign \new_[23583]_  = A167 & A168;
  assign \new_[23587]_  = ~A201 & A200;
  assign \new_[23588]_  = A199 & \new_[23587]_ ;
  assign \new_[23589]_  = \new_[23588]_  & \new_[23583]_ ;
  assign \new_[23593]_  = A234 & A232;
  assign \new_[23594]_  = ~A202 & \new_[23593]_ ;
  assign \new_[23598]_  = A269 & ~A266;
  assign \new_[23599]_  = A265 & \new_[23598]_ ;
  assign \new_[23600]_  = \new_[23599]_  & \new_[23594]_ ;
  assign \new_[23603]_  = A167 & A168;
  assign \new_[23607]_  = ~A201 & A200;
  assign \new_[23608]_  = A199 & \new_[23607]_ ;
  assign \new_[23609]_  = \new_[23608]_  & \new_[23603]_ ;
  assign \new_[23613]_  = A234 & A233;
  assign \new_[23614]_  = ~A202 & \new_[23613]_ ;
  assign \new_[23618]_  = A302 & ~A299;
  assign \new_[23619]_  = A298 & \new_[23618]_ ;
  assign \new_[23620]_  = \new_[23619]_  & \new_[23614]_ ;
  assign \new_[23623]_  = A167 & A168;
  assign \new_[23627]_  = ~A201 & A200;
  assign \new_[23628]_  = A199 & \new_[23627]_ ;
  assign \new_[23629]_  = \new_[23628]_  & \new_[23623]_ ;
  assign \new_[23633]_  = A234 & A233;
  assign \new_[23634]_  = ~A202 & \new_[23633]_ ;
  assign \new_[23638]_  = A302 & A299;
  assign \new_[23639]_  = ~A298 & \new_[23638]_ ;
  assign \new_[23640]_  = \new_[23639]_  & \new_[23634]_ ;
  assign \new_[23643]_  = A167 & A168;
  assign \new_[23647]_  = ~A201 & A200;
  assign \new_[23648]_  = A199 & \new_[23647]_ ;
  assign \new_[23649]_  = \new_[23648]_  & \new_[23643]_ ;
  assign \new_[23653]_  = A234 & A233;
  assign \new_[23654]_  = ~A202 & \new_[23653]_ ;
  assign \new_[23658]_  = A269 & A266;
  assign \new_[23659]_  = ~A265 & \new_[23658]_ ;
  assign \new_[23660]_  = \new_[23659]_  & \new_[23654]_ ;
  assign \new_[23663]_  = A167 & A168;
  assign \new_[23667]_  = ~A201 & A200;
  assign \new_[23668]_  = A199 & \new_[23667]_ ;
  assign \new_[23669]_  = \new_[23668]_  & \new_[23663]_ ;
  assign \new_[23673]_  = A234 & A233;
  assign \new_[23674]_  = ~A202 & \new_[23673]_ ;
  assign \new_[23678]_  = A269 & ~A266;
  assign \new_[23679]_  = A265 & \new_[23678]_ ;
  assign \new_[23680]_  = \new_[23679]_  & \new_[23674]_ ;
  assign \new_[23683]_  = A167 & A168;
  assign \new_[23687]_  = ~A201 & A200;
  assign \new_[23688]_  = A199 & \new_[23687]_ ;
  assign \new_[23689]_  = \new_[23688]_  & \new_[23683]_ ;
  assign \new_[23693]_  = A233 & ~A232;
  assign \new_[23694]_  = ~A202 & \new_[23693]_ ;
  assign \new_[23698]_  = A300 & A299;
  assign \new_[23699]_  = A236 & \new_[23698]_ ;
  assign \new_[23700]_  = \new_[23699]_  & \new_[23694]_ ;
  assign \new_[23703]_  = A167 & A168;
  assign \new_[23707]_  = ~A201 & A200;
  assign \new_[23708]_  = A199 & \new_[23707]_ ;
  assign \new_[23709]_  = \new_[23708]_  & \new_[23703]_ ;
  assign \new_[23713]_  = A233 & ~A232;
  assign \new_[23714]_  = ~A202 & \new_[23713]_ ;
  assign \new_[23718]_  = A300 & A298;
  assign \new_[23719]_  = A236 & \new_[23718]_ ;
  assign \new_[23720]_  = \new_[23719]_  & \new_[23714]_ ;
  assign \new_[23723]_  = A167 & A168;
  assign \new_[23727]_  = ~A201 & A200;
  assign \new_[23728]_  = A199 & \new_[23727]_ ;
  assign \new_[23729]_  = \new_[23728]_  & \new_[23723]_ ;
  assign \new_[23733]_  = A233 & ~A232;
  assign \new_[23734]_  = ~A202 & \new_[23733]_ ;
  assign \new_[23738]_  = A267 & A265;
  assign \new_[23739]_  = A236 & \new_[23738]_ ;
  assign \new_[23740]_  = \new_[23739]_  & \new_[23734]_ ;
  assign \new_[23743]_  = A167 & A168;
  assign \new_[23747]_  = ~A201 & A200;
  assign \new_[23748]_  = A199 & \new_[23747]_ ;
  assign \new_[23749]_  = \new_[23748]_  & \new_[23743]_ ;
  assign \new_[23753]_  = A233 & ~A232;
  assign \new_[23754]_  = ~A202 & \new_[23753]_ ;
  assign \new_[23758]_  = A267 & A266;
  assign \new_[23759]_  = A236 & \new_[23758]_ ;
  assign \new_[23760]_  = \new_[23759]_  & \new_[23754]_ ;
  assign \new_[23763]_  = A167 & A168;
  assign \new_[23767]_  = ~A201 & A200;
  assign \new_[23768]_  = A199 & \new_[23767]_ ;
  assign \new_[23769]_  = \new_[23768]_  & \new_[23763]_ ;
  assign \new_[23773]_  = ~A233 & A232;
  assign \new_[23774]_  = ~A202 & \new_[23773]_ ;
  assign \new_[23778]_  = A300 & A299;
  assign \new_[23779]_  = A236 & \new_[23778]_ ;
  assign \new_[23780]_  = \new_[23779]_  & \new_[23774]_ ;
  assign \new_[23783]_  = A167 & A168;
  assign \new_[23787]_  = ~A201 & A200;
  assign \new_[23788]_  = A199 & \new_[23787]_ ;
  assign \new_[23789]_  = \new_[23788]_  & \new_[23783]_ ;
  assign \new_[23793]_  = ~A233 & A232;
  assign \new_[23794]_  = ~A202 & \new_[23793]_ ;
  assign \new_[23798]_  = A300 & A298;
  assign \new_[23799]_  = A236 & \new_[23798]_ ;
  assign \new_[23800]_  = \new_[23799]_  & \new_[23794]_ ;
  assign \new_[23803]_  = A167 & A168;
  assign \new_[23807]_  = ~A201 & A200;
  assign \new_[23808]_  = A199 & \new_[23807]_ ;
  assign \new_[23809]_  = \new_[23808]_  & \new_[23803]_ ;
  assign \new_[23813]_  = ~A233 & A232;
  assign \new_[23814]_  = ~A202 & \new_[23813]_ ;
  assign \new_[23818]_  = A267 & A265;
  assign \new_[23819]_  = A236 & \new_[23818]_ ;
  assign \new_[23820]_  = \new_[23819]_  & \new_[23814]_ ;
  assign \new_[23823]_  = A167 & A168;
  assign \new_[23827]_  = ~A201 & A200;
  assign \new_[23828]_  = A199 & \new_[23827]_ ;
  assign \new_[23829]_  = \new_[23828]_  & \new_[23823]_ ;
  assign \new_[23833]_  = ~A233 & A232;
  assign \new_[23834]_  = ~A202 & \new_[23833]_ ;
  assign \new_[23838]_  = A267 & A266;
  assign \new_[23839]_  = A236 & \new_[23838]_ ;
  assign \new_[23840]_  = \new_[23839]_  & \new_[23834]_ ;
  assign \new_[23843]_  = A167 & A168;
  assign \new_[23847]_  = ~A202 & ~A200;
  assign \new_[23848]_  = ~A199 & \new_[23847]_ ;
  assign \new_[23849]_  = \new_[23848]_  & \new_[23843]_ ;
  assign \new_[23853]_  = A236 & A233;
  assign \new_[23854]_  = ~A232 & \new_[23853]_ ;
  assign \new_[23858]_  = A302 & ~A299;
  assign \new_[23859]_  = A298 & \new_[23858]_ ;
  assign \new_[23860]_  = \new_[23859]_  & \new_[23854]_ ;
  assign \new_[23863]_  = A167 & A168;
  assign \new_[23867]_  = ~A202 & ~A200;
  assign \new_[23868]_  = ~A199 & \new_[23867]_ ;
  assign \new_[23869]_  = \new_[23868]_  & \new_[23863]_ ;
  assign \new_[23873]_  = A236 & A233;
  assign \new_[23874]_  = ~A232 & \new_[23873]_ ;
  assign \new_[23878]_  = A302 & A299;
  assign \new_[23879]_  = ~A298 & \new_[23878]_ ;
  assign \new_[23880]_  = \new_[23879]_  & \new_[23874]_ ;
  assign \new_[23883]_  = A167 & A168;
  assign \new_[23887]_  = ~A202 & ~A200;
  assign \new_[23888]_  = ~A199 & \new_[23887]_ ;
  assign \new_[23889]_  = \new_[23888]_  & \new_[23883]_ ;
  assign \new_[23893]_  = A236 & A233;
  assign \new_[23894]_  = ~A232 & \new_[23893]_ ;
  assign \new_[23898]_  = A269 & A266;
  assign \new_[23899]_  = ~A265 & \new_[23898]_ ;
  assign \new_[23900]_  = \new_[23899]_  & \new_[23894]_ ;
  assign \new_[23903]_  = A167 & A168;
  assign \new_[23907]_  = ~A202 & ~A200;
  assign \new_[23908]_  = ~A199 & \new_[23907]_ ;
  assign \new_[23909]_  = \new_[23908]_  & \new_[23903]_ ;
  assign \new_[23913]_  = A236 & A233;
  assign \new_[23914]_  = ~A232 & \new_[23913]_ ;
  assign \new_[23918]_  = A269 & ~A266;
  assign \new_[23919]_  = A265 & \new_[23918]_ ;
  assign \new_[23920]_  = \new_[23919]_  & \new_[23914]_ ;
  assign \new_[23923]_  = A167 & A168;
  assign \new_[23927]_  = ~A202 & ~A200;
  assign \new_[23928]_  = ~A199 & \new_[23927]_ ;
  assign \new_[23929]_  = \new_[23928]_  & \new_[23923]_ ;
  assign \new_[23933]_  = A236 & ~A233;
  assign \new_[23934]_  = A232 & \new_[23933]_ ;
  assign \new_[23938]_  = A302 & ~A299;
  assign \new_[23939]_  = A298 & \new_[23938]_ ;
  assign \new_[23940]_  = \new_[23939]_  & \new_[23934]_ ;
  assign \new_[23943]_  = A167 & A168;
  assign \new_[23947]_  = ~A202 & ~A200;
  assign \new_[23948]_  = ~A199 & \new_[23947]_ ;
  assign \new_[23949]_  = \new_[23948]_  & \new_[23943]_ ;
  assign \new_[23953]_  = A236 & ~A233;
  assign \new_[23954]_  = A232 & \new_[23953]_ ;
  assign \new_[23958]_  = A302 & A299;
  assign \new_[23959]_  = ~A298 & \new_[23958]_ ;
  assign \new_[23960]_  = \new_[23959]_  & \new_[23954]_ ;
  assign \new_[23963]_  = A167 & A168;
  assign \new_[23967]_  = ~A202 & ~A200;
  assign \new_[23968]_  = ~A199 & \new_[23967]_ ;
  assign \new_[23969]_  = \new_[23968]_  & \new_[23963]_ ;
  assign \new_[23973]_  = A236 & ~A233;
  assign \new_[23974]_  = A232 & \new_[23973]_ ;
  assign \new_[23978]_  = A269 & A266;
  assign \new_[23979]_  = ~A265 & \new_[23978]_ ;
  assign \new_[23980]_  = \new_[23979]_  & \new_[23974]_ ;
  assign \new_[23983]_  = A167 & A168;
  assign \new_[23987]_  = ~A202 & ~A200;
  assign \new_[23988]_  = ~A199 & \new_[23987]_ ;
  assign \new_[23989]_  = \new_[23988]_  & \new_[23983]_ ;
  assign \new_[23993]_  = A236 & ~A233;
  assign \new_[23994]_  = A232 & \new_[23993]_ ;
  assign \new_[23998]_  = A269 & ~A266;
  assign \new_[23999]_  = A265 & \new_[23998]_ ;
  assign \new_[24000]_  = \new_[23999]_  & \new_[23994]_ ;
  assign \new_[24003]_  = A167 & A170;
  assign \new_[24007]_  = ~A202 & ~A201;
  assign \new_[24008]_  = ~A166 & \new_[24007]_ ;
  assign \new_[24009]_  = \new_[24008]_  & \new_[24003]_ ;
  assign \new_[24013]_  = A234 & A232;
  assign \new_[24014]_  = ~A203 & \new_[24013]_ ;
  assign \new_[24018]_  = A302 & ~A299;
  assign \new_[24019]_  = A298 & \new_[24018]_ ;
  assign \new_[24020]_  = \new_[24019]_  & \new_[24014]_ ;
  assign \new_[24023]_  = A167 & A170;
  assign \new_[24027]_  = ~A202 & ~A201;
  assign \new_[24028]_  = ~A166 & \new_[24027]_ ;
  assign \new_[24029]_  = \new_[24028]_  & \new_[24023]_ ;
  assign \new_[24033]_  = A234 & A232;
  assign \new_[24034]_  = ~A203 & \new_[24033]_ ;
  assign \new_[24038]_  = A302 & A299;
  assign \new_[24039]_  = ~A298 & \new_[24038]_ ;
  assign \new_[24040]_  = \new_[24039]_  & \new_[24034]_ ;
  assign \new_[24043]_  = A167 & A170;
  assign \new_[24047]_  = ~A202 & ~A201;
  assign \new_[24048]_  = ~A166 & \new_[24047]_ ;
  assign \new_[24049]_  = \new_[24048]_  & \new_[24043]_ ;
  assign \new_[24053]_  = A234 & A232;
  assign \new_[24054]_  = ~A203 & \new_[24053]_ ;
  assign \new_[24058]_  = A269 & A266;
  assign \new_[24059]_  = ~A265 & \new_[24058]_ ;
  assign \new_[24060]_  = \new_[24059]_  & \new_[24054]_ ;
  assign \new_[24063]_  = A167 & A170;
  assign \new_[24067]_  = ~A202 & ~A201;
  assign \new_[24068]_  = ~A166 & \new_[24067]_ ;
  assign \new_[24069]_  = \new_[24068]_  & \new_[24063]_ ;
  assign \new_[24073]_  = A234 & A232;
  assign \new_[24074]_  = ~A203 & \new_[24073]_ ;
  assign \new_[24078]_  = A269 & ~A266;
  assign \new_[24079]_  = A265 & \new_[24078]_ ;
  assign \new_[24080]_  = \new_[24079]_  & \new_[24074]_ ;
  assign \new_[24083]_  = A167 & A170;
  assign \new_[24087]_  = ~A202 & ~A201;
  assign \new_[24088]_  = ~A166 & \new_[24087]_ ;
  assign \new_[24089]_  = \new_[24088]_  & \new_[24083]_ ;
  assign \new_[24093]_  = A234 & A233;
  assign \new_[24094]_  = ~A203 & \new_[24093]_ ;
  assign \new_[24098]_  = A302 & ~A299;
  assign \new_[24099]_  = A298 & \new_[24098]_ ;
  assign \new_[24100]_  = \new_[24099]_  & \new_[24094]_ ;
  assign \new_[24103]_  = A167 & A170;
  assign \new_[24107]_  = ~A202 & ~A201;
  assign \new_[24108]_  = ~A166 & \new_[24107]_ ;
  assign \new_[24109]_  = \new_[24108]_  & \new_[24103]_ ;
  assign \new_[24113]_  = A234 & A233;
  assign \new_[24114]_  = ~A203 & \new_[24113]_ ;
  assign \new_[24118]_  = A302 & A299;
  assign \new_[24119]_  = ~A298 & \new_[24118]_ ;
  assign \new_[24120]_  = \new_[24119]_  & \new_[24114]_ ;
  assign \new_[24123]_  = A167 & A170;
  assign \new_[24127]_  = ~A202 & ~A201;
  assign \new_[24128]_  = ~A166 & \new_[24127]_ ;
  assign \new_[24129]_  = \new_[24128]_  & \new_[24123]_ ;
  assign \new_[24133]_  = A234 & A233;
  assign \new_[24134]_  = ~A203 & \new_[24133]_ ;
  assign \new_[24138]_  = A269 & A266;
  assign \new_[24139]_  = ~A265 & \new_[24138]_ ;
  assign \new_[24140]_  = \new_[24139]_  & \new_[24134]_ ;
  assign \new_[24143]_  = A167 & A170;
  assign \new_[24147]_  = ~A202 & ~A201;
  assign \new_[24148]_  = ~A166 & \new_[24147]_ ;
  assign \new_[24149]_  = \new_[24148]_  & \new_[24143]_ ;
  assign \new_[24153]_  = A234 & A233;
  assign \new_[24154]_  = ~A203 & \new_[24153]_ ;
  assign \new_[24158]_  = A269 & ~A266;
  assign \new_[24159]_  = A265 & \new_[24158]_ ;
  assign \new_[24160]_  = \new_[24159]_  & \new_[24154]_ ;
  assign \new_[24163]_  = A167 & A170;
  assign \new_[24167]_  = ~A202 & ~A201;
  assign \new_[24168]_  = ~A166 & \new_[24167]_ ;
  assign \new_[24169]_  = \new_[24168]_  & \new_[24163]_ ;
  assign \new_[24173]_  = A233 & ~A232;
  assign \new_[24174]_  = ~A203 & \new_[24173]_ ;
  assign \new_[24178]_  = A300 & A299;
  assign \new_[24179]_  = A236 & \new_[24178]_ ;
  assign \new_[24180]_  = \new_[24179]_  & \new_[24174]_ ;
  assign \new_[24183]_  = A167 & A170;
  assign \new_[24187]_  = ~A202 & ~A201;
  assign \new_[24188]_  = ~A166 & \new_[24187]_ ;
  assign \new_[24189]_  = \new_[24188]_  & \new_[24183]_ ;
  assign \new_[24193]_  = A233 & ~A232;
  assign \new_[24194]_  = ~A203 & \new_[24193]_ ;
  assign \new_[24198]_  = A300 & A298;
  assign \new_[24199]_  = A236 & \new_[24198]_ ;
  assign \new_[24200]_  = \new_[24199]_  & \new_[24194]_ ;
  assign \new_[24203]_  = A167 & A170;
  assign \new_[24207]_  = ~A202 & ~A201;
  assign \new_[24208]_  = ~A166 & \new_[24207]_ ;
  assign \new_[24209]_  = \new_[24208]_  & \new_[24203]_ ;
  assign \new_[24213]_  = A233 & ~A232;
  assign \new_[24214]_  = ~A203 & \new_[24213]_ ;
  assign \new_[24218]_  = A267 & A265;
  assign \new_[24219]_  = A236 & \new_[24218]_ ;
  assign \new_[24220]_  = \new_[24219]_  & \new_[24214]_ ;
  assign \new_[24223]_  = A167 & A170;
  assign \new_[24227]_  = ~A202 & ~A201;
  assign \new_[24228]_  = ~A166 & \new_[24227]_ ;
  assign \new_[24229]_  = \new_[24228]_  & \new_[24223]_ ;
  assign \new_[24233]_  = A233 & ~A232;
  assign \new_[24234]_  = ~A203 & \new_[24233]_ ;
  assign \new_[24238]_  = A267 & A266;
  assign \new_[24239]_  = A236 & \new_[24238]_ ;
  assign \new_[24240]_  = \new_[24239]_  & \new_[24234]_ ;
  assign \new_[24243]_  = A167 & A170;
  assign \new_[24247]_  = ~A202 & ~A201;
  assign \new_[24248]_  = ~A166 & \new_[24247]_ ;
  assign \new_[24249]_  = \new_[24248]_  & \new_[24243]_ ;
  assign \new_[24253]_  = ~A233 & A232;
  assign \new_[24254]_  = ~A203 & \new_[24253]_ ;
  assign \new_[24258]_  = A300 & A299;
  assign \new_[24259]_  = A236 & \new_[24258]_ ;
  assign \new_[24260]_  = \new_[24259]_  & \new_[24254]_ ;
  assign \new_[24263]_  = A167 & A170;
  assign \new_[24267]_  = ~A202 & ~A201;
  assign \new_[24268]_  = ~A166 & \new_[24267]_ ;
  assign \new_[24269]_  = \new_[24268]_  & \new_[24263]_ ;
  assign \new_[24273]_  = ~A233 & A232;
  assign \new_[24274]_  = ~A203 & \new_[24273]_ ;
  assign \new_[24278]_  = A300 & A298;
  assign \new_[24279]_  = A236 & \new_[24278]_ ;
  assign \new_[24280]_  = \new_[24279]_  & \new_[24274]_ ;
  assign \new_[24283]_  = A167 & A170;
  assign \new_[24287]_  = ~A202 & ~A201;
  assign \new_[24288]_  = ~A166 & \new_[24287]_ ;
  assign \new_[24289]_  = \new_[24288]_  & \new_[24283]_ ;
  assign \new_[24293]_  = ~A233 & A232;
  assign \new_[24294]_  = ~A203 & \new_[24293]_ ;
  assign \new_[24298]_  = A267 & A265;
  assign \new_[24299]_  = A236 & \new_[24298]_ ;
  assign \new_[24300]_  = \new_[24299]_  & \new_[24294]_ ;
  assign \new_[24303]_  = A167 & A170;
  assign \new_[24307]_  = ~A202 & ~A201;
  assign \new_[24308]_  = ~A166 & \new_[24307]_ ;
  assign \new_[24309]_  = \new_[24308]_  & \new_[24303]_ ;
  assign \new_[24313]_  = ~A233 & A232;
  assign \new_[24314]_  = ~A203 & \new_[24313]_ ;
  assign \new_[24318]_  = A267 & A266;
  assign \new_[24319]_  = A236 & \new_[24318]_ ;
  assign \new_[24320]_  = \new_[24319]_  & \new_[24314]_ ;
  assign \new_[24323]_  = A167 & A170;
  assign \new_[24327]_  = A200 & A199;
  assign \new_[24328]_  = ~A166 & \new_[24327]_ ;
  assign \new_[24329]_  = \new_[24328]_  & \new_[24323]_ ;
  assign \new_[24333]_  = A235 & ~A202;
  assign \new_[24334]_  = ~A201 & \new_[24333]_ ;
  assign \new_[24338]_  = A302 & ~A299;
  assign \new_[24339]_  = A298 & \new_[24338]_ ;
  assign \new_[24340]_  = \new_[24339]_  & \new_[24334]_ ;
  assign \new_[24343]_  = A167 & A170;
  assign \new_[24347]_  = A200 & A199;
  assign \new_[24348]_  = ~A166 & \new_[24347]_ ;
  assign \new_[24349]_  = \new_[24348]_  & \new_[24343]_ ;
  assign \new_[24353]_  = A235 & ~A202;
  assign \new_[24354]_  = ~A201 & \new_[24353]_ ;
  assign \new_[24358]_  = A302 & A299;
  assign \new_[24359]_  = ~A298 & \new_[24358]_ ;
  assign \new_[24360]_  = \new_[24359]_  & \new_[24354]_ ;
  assign \new_[24363]_  = A167 & A170;
  assign \new_[24367]_  = A200 & A199;
  assign \new_[24368]_  = ~A166 & \new_[24367]_ ;
  assign \new_[24369]_  = \new_[24368]_  & \new_[24363]_ ;
  assign \new_[24373]_  = A235 & ~A202;
  assign \new_[24374]_  = ~A201 & \new_[24373]_ ;
  assign \new_[24378]_  = A269 & A266;
  assign \new_[24379]_  = ~A265 & \new_[24378]_ ;
  assign \new_[24380]_  = \new_[24379]_  & \new_[24374]_ ;
  assign \new_[24383]_  = A167 & A170;
  assign \new_[24387]_  = A200 & A199;
  assign \new_[24388]_  = ~A166 & \new_[24387]_ ;
  assign \new_[24389]_  = \new_[24388]_  & \new_[24383]_ ;
  assign \new_[24393]_  = A235 & ~A202;
  assign \new_[24394]_  = ~A201 & \new_[24393]_ ;
  assign \new_[24398]_  = A269 & ~A266;
  assign \new_[24399]_  = A265 & \new_[24398]_ ;
  assign \new_[24400]_  = \new_[24399]_  & \new_[24394]_ ;
  assign \new_[24403]_  = A167 & A170;
  assign \new_[24407]_  = A200 & A199;
  assign \new_[24408]_  = ~A166 & \new_[24407]_ ;
  assign \new_[24409]_  = \new_[24408]_  & \new_[24403]_ ;
  assign \new_[24413]_  = A232 & ~A202;
  assign \new_[24414]_  = ~A201 & \new_[24413]_ ;
  assign \new_[24418]_  = A300 & A299;
  assign \new_[24419]_  = A234 & \new_[24418]_ ;
  assign \new_[24420]_  = \new_[24419]_  & \new_[24414]_ ;
  assign \new_[24423]_  = A167 & A170;
  assign \new_[24427]_  = A200 & A199;
  assign \new_[24428]_  = ~A166 & \new_[24427]_ ;
  assign \new_[24429]_  = \new_[24428]_  & \new_[24423]_ ;
  assign \new_[24433]_  = A232 & ~A202;
  assign \new_[24434]_  = ~A201 & \new_[24433]_ ;
  assign \new_[24438]_  = A300 & A298;
  assign \new_[24439]_  = A234 & \new_[24438]_ ;
  assign \new_[24440]_  = \new_[24439]_  & \new_[24434]_ ;
  assign \new_[24443]_  = A167 & A170;
  assign \new_[24447]_  = A200 & A199;
  assign \new_[24448]_  = ~A166 & \new_[24447]_ ;
  assign \new_[24449]_  = \new_[24448]_  & \new_[24443]_ ;
  assign \new_[24453]_  = A232 & ~A202;
  assign \new_[24454]_  = ~A201 & \new_[24453]_ ;
  assign \new_[24458]_  = A267 & A265;
  assign \new_[24459]_  = A234 & \new_[24458]_ ;
  assign \new_[24460]_  = \new_[24459]_  & \new_[24454]_ ;
  assign \new_[24463]_  = A167 & A170;
  assign \new_[24467]_  = A200 & A199;
  assign \new_[24468]_  = ~A166 & \new_[24467]_ ;
  assign \new_[24469]_  = \new_[24468]_  & \new_[24463]_ ;
  assign \new_[24473]_  = A232 & ~A202;
  assign \new_[24474]_  = ~A201 & \new_[24473]_ ;
  assign \new_[24478]_  = A267 & A266;
  assign \new_[24479]_  = A234 & \new_[24478]_ ;
  assign \new_[24480]_  = \new_[24479]_  & \new_[24474]_ ;
  assign \new_[24483]_  = A167 & A170;
  assign \new_[24487]_  = A200 & A199;
  assign \new_[24488]_  = ~A166 & \new_[24487]_ ;
  assign \new_[24489]_  = \new_[24488]_  & \new_[24483]_ ;
  assign \new_[24493]_  = A233 & ~A202;
  assign \new_[24494]_  = ~A201 & \new_[24493]_ ;
  assign \new_[24498]_  = A300 & A299;
  assign \new_[24499]_  = A234 & \new_[24498]_ ;
  assign \new_[24500]_  = \new_[24499]_  & \new_[24494]_ ;
  assign \new_[24503]_  = A167 & A170;
  assign \new_[24507]_  = A200 & A199;
  assign \new_[24508]_  = ~A166 & \new_[24507]_ ;
  assign \new_[24509]_  = \new_[24508]_  & \new_[24503]_ ;
  assign \new_[24513]_  = A233 & ~A202;
  assign \new_[24514]_  = ~A201 & \new_[24513]_ ;
  assign \new_[24518]_  = A300 & A298;
  assign \new_[24519]_  = A234 & \new_[24518]_ ;
  assign \new_[24520]_  = \new_[24519]_  & \new_[24514]_ ;
  assign \new_[24523]_  = A167 & A170;
  assign \new_[24527]_  = A200 & A199;
  assign \new_[24528]_  = ~A166 & \new_[24527]_ ;
  assign \new_[24529]_  = \new_[24528]_  & \new_[24523]_ ;
  assign \new_[24533]_  = A233 & ~A202;
  assign \new_[24534]_  = ~A201 & \new_[24533]_ ;
  assign \new_[24538]_  = A267 & A265;
  assign \new_[24539]_  = A234 & \new_[24538]_ ;
  assign \new_[24540]_  = \new_[24539]_  & \new_[24534]_ ;
  assign \new_[24543]_  = A167 & A170;
  assign \new_[24547]_  = A200 & A199;
  assign \new_[24548]_  = ~A166 & \new_[24547]_ ;
  assign \new_[24549]_  = \new_[24548]_  & \new_[24543]_ ;
  assign \new_[24553]_  = A233 & ~A202;
  assign \new_[24554]_  = ~A201 & \new_[24553]_ ;
  assign \new_[24558]_  = A267 & A266;
  assign \new_[24559]_  = A234 & \new_[24558]_ ;
  assign \new_[24560]_  = \new_[24559]_  & \new_[24554]_ ;
  assign \new_[24563]_  = A167 & A170;
  assign \new_[24567]_  = A200 & A199;
  assign \new_[24568]_  = ~A166 & \new_[24567]_ ;
  assign \new_[24569]_  = \new_[24568]_  & \new_[24563]_ ;
  assign \new_[24573]_  = ~A232 & ~A202;
  assign \new_[24574]_  = ~A201 & \new_[24573]_ ;
  assign \new_[24578]_  = A301 & A236;
  assign \new_[24579]_  = A233 & \new_[24578]_ ;
  assign \new_[24580]_  = \new_[24579]_  & \new_[24574]_ ;
  assign \new_[24583]_  = A167 & A170;
  assign \new_[24587]_  = A200 & A199;
  assign \new_[24588]_  = ~A166 & \new_[24587]_ ;
  assign \new_[24589]_  = \new_[24588]_  & \new_[24583]_ ;
  assign \new_[24593]_  = ~A232 & ~A202;
  assign \new_[24594]_  = ~A201 & \new_[24593]_ ;
  assign \new_[24598]_  = A268 & A236;
  assign \new_[24599]_  = A233 & \new_[24598]_ ;
  assign \new_[24600]_  = \new_[24599]_  & \new_[24594]_ ;
  assign \new_[24603]_  = A167 & A170;
  assign \new_[24607]_  = A200 & A199;
  assign \new_[24608]_  = ~A166 & \new_[24607]_ ;
  assign \new_[24609]_  = \new_[24608]_  & \new_[24603]_ ;
  assign \new_[24613]_  = A232 & ~A202;
  assign \new_[24614]_  = ~A201 & \new_[24613]_ ;
  assign \new_[24618]_  = A301 & A236;
  assign \new_[24619]_  = ~A233 & \new_[24618]_ ;
  assign \new_[24620]_  = \new_[24619]_  & \new_[24614]_ ;
  assign \new_[24623]_  = A167 & A170;
  assign \new_[24627]_  = A200 & A199;
  assign \new_[24628]_  = ~A166 & \new_[24627]_ ;
  assign \new_[24629]_  = \new_[24628]_  & \new_[24623]_ ;
  assign \new_[24633]_  = A232 & ~A202;
  assign \new_[24634]_  = ~A201 & \new_[24633]_ ;
  assign \new_[24638]_  = A268 & A236;
  assign \new_[24639]_  = ~A233 & \new_[24638]_ ;
  assign \new_[24640]_  = \new_[24639]_  & \new_[24634]_ ;
  assign \new_[24643]_  = A167 & A170;
  assign \new_[24647]_  = ~A200 & ~A199;
  assign \new_[24648]_  = ~A166 & \new_[24647]_ ;
  assign \new_[24649]_  = \new_[24648]_  & \new_[24643]_ ;
  assign \new_[24653]_  = A234 & A232;
  assign \new_[24654]_  = ~A202 & \new_[24653]_ ;
  assign \new_[24658]_  = A302 & ~A299;
  assign \new_[24659]_  = A298 & \new_[24658]_ ;
  assign \new_[24660]_  = \new_[24659]_  & \new_[24654]_ ;
  assign \new_[24663]_  = A167 & A170;
  assign \new_[24667]_  = ~A200 & ~A199;
  assign \new_[24668]_  = ~A166 & \new_[24667]_ ;
  assign \new_[24669]_  = \new_[24668]_  & \new_[24663]_ ;
  assign \new_[24673]_  = A234 & A232;
  assign \new_[24674]_  = ~A202 & \new_[24673]_ ;
  assign \new_[24678]_  = A302 & A299;
  assign \new_[24679]_  = ~A298 & \new_[24678]_ ;
  assign \new_[24680]_  = \new_[24679]_  & \new_[24674]_ ;
  assign \new_[24683]_  = A167 & A170;
  assign \new_[24687]_  = ~A200 & ~A199;
  assign \new_[24688]_  = ~A166 & \new_[24687]_ ;
  assign \new_[24689]_  = \new_[24688]_  & \new_[24683]_ ;
  assign \new_[24693]_  = A234 & A232;
  assign \new_[24694]_  = ~A202 & \new_[24693]_ ;
  assign \new_[24698]_  = A269 & A266;
  assign \new_[24699]_  = ~A265 & \new_[24698]_ ;
  assign \new_[24700]_  = \new_[24699]_  & \new_[24694]_ ;
  assign \new_[24703]_  = A167 & A170;
  assign \new_[24707]_  = ~A200 & ~A199;
  assign \new_[24708]_  = ~A166 & \new_[24707]_ ;
  assign \new_[24709]_  = \new_[24708]_  & \new_[24703]_ ;
  assign \new_[24713]_  = A234 & A232;
  assign \new_[24714]_  = ~A202 & \new_[24713]_ ;
  assign \new_[24718]_  = A269 & ~A266;
  assign \new_[24719]_  = A265 & \new_[24718]_ ;
  assign \new_[24720]_  = \new_[24719]_  & \new_[24714]_ ;
  assign \new_[24723]_  = A167 & A170;
  assign \new_[24727]_  = ~A200 & ~A199;
  assign \new_[24728]_  = ~A166 & \new_[24727]_ ;
  assign \new_[24729]_  = \new_[24728]_  & \new_[24723]_ ;
  assign \new_[24733]_  = A234 & A233;
  assign \new_[24734]_  = ~A202 & \new_[24733]_ ;
  assign \new_[24738]_  = A302 & ~A299;
  assign \new_[24739]_  = A298 & \new_[24738]_ ;
  assign \new_[24740]_  = \new_[24739]_  & \new_[24734]_ ;
  assign \new_[24743]_  = A167 & A170;
  assign \new_[24747]_  = ~A200 & ~A199;
  assign \new_[24748]_  = ~A166 & \new_[24747]_ ;
  assign \new_[24749]_  = \new_[24748]_  & \new_[24743]_ ;
  assign \new_[24753]_  = A234 & A233;
  assign \new_[24754]_  = ~A202 & \new_[24753]_ ;
  assign \new_[24758]_  = A302 & A299;
  assign \new_[24759]_  = ~A298 & \new_[24758]_ ;
  assign \new_[24760]_  = \new_[24759]_  & \new_[24754]_ ;
  assign \new_[24763]_  = A167 & A170;
  assign \new_[24767]_  = ~A200 & ~A199;
  assign \new_[24768]_  = ~A166 & \new_[24767]_ ;
  assign \new_[24769]_  = \new_[24768]_  & \new_[24763]_ ;
  assign \new_[24773]_  = A234 & A233;
  assign \new_[24774]_  = ~A202 & \new_[24773]_ ;
  assign \new_[24778]_  = A269 & A266;
  assign \new_[24779]_  = ~A265 & \new_[24778]_ ;
  assign \new_[24780]_  = \new_[24779]_  & \new_[24774]_ ;
  assign \new_[24783]_  = A167 & A170;
  assign \new_[24787]_  = ~A200 & ~A199;
  assign \new_[24788]_  = ~A166 & \new_[24787]_ ;
  assign \new_[24789]_  = \new_[24788]_  & \new_[24783]_ ;
  assign \new_[24793]_  = A234 & A233;
  assign \new_[24794]_  = ~A202 & \new_[24793]_ ;
  assign \new_[24798]_  = A269 & ~A266;
  assign \new_[24799]_  = A265 & \new_[24798]_ ;
  assign \new_[24800]_  = \new_[24799]_  & \new_[24794]_ ;
  assign \new_[24803]_  = A167 & A170;
  assign \new_[24807]_  = ~A200 & ~A199;
  assign \new_[24808]_  = ~A166 & \new_[24807]_ ;
  assign \new_[24809]_  = \new_[24808]_  & \new_[24803]_ ;
  assign \new_[24813]_  = A233 & ~A232;
  assign \new_[24814]_  = ~A202 & \new_[24813]_ ;
  assign \new_[24818]_  = A300 & A299;
  assign \new_[24819]_  = A236 & \new_[24818]_ ;
  assign \new_[24820]_  = \new_[24819]_  & \new_[24814]_ ;
  assign \new_[24823]_  = A167 & A170;
  assign \new_[24827]_  = ~A200 & ~A199;
  assign \new_[24828]_  = ~A166 & \new_[24827]_ ;
  assign \new_[24829]_  = \new_[24828]_  & \new_[24823]_ ;
  assign \new_[24833]_  = A233 & ~A232;
  assign \new_[24834]_  = ~A202 & \new_[24833]_ ;
  assign \new_[24838]_  = A300 & A298;
  assign \new_[24839]_  = A236 & \new_[24838]_ ;
  assign \new_[24840]_  = \new_[24839]_  & \new_[24834]_ ;
  assign \new_[24843]_  = A167 & A170;
  assign \new_[24847]_  = ~A200 & ~A199;
  assign \new_[24848]_  = ~A166 & \new_[24847]_ ;
  assign \new_[24849]_  = \new_[24848]_  & \new_[24843]_ ;
  assign \new_[24853]_  = A233 & ~A232;
  assign \new_[24854]_  = ~A202 & \new_[24853]_ ;
  assign \new_[24858]_  = A267 & A265;
  assign \new_[24859]_  = A236 & \new_[24858]_ ;
  assign \new_[24860]_  = \new_[24859]_  & \new_[24854]_ ;
  assign \new_[24863]_  = A167 & A170;
  assign \new_[24867]_  = ~A200 & ~A199;
  assign \new_[24868]_  = ~A166 & \new_[24867]_ ;
  assign \new_[24869]_  = \new_[24868]_  & \new_[24863]_ ;
  assign \new_[24873]_  = A233 & ~A232;
  assign \new_[24874]_  = ~A202 & \new_[24873]_ ;
  assign \new_[24878]_  = A267 & A266;
  assign \new_[24879]_  = A236 & \new_[24878]_ ;
  assign \new_[24880]_  = \new_[24879]_  & \new_[24874]_ ;
  assign \new_[24883]_  = A167 & A170;
  assign \new_[24887]_  = ~A200 & ~A199;
  assign \new_[24888]_  = ~A166 & \new_[24887]_ ;
  assign \new_[24889]_  = \new_[24888]_  & \new_[24883]_ ;
  assign \new_[24893]_  = ~A233 & A232;
  assign \new_[24894]_  = ~A202 & \new_[24893]_ ;
  assign \new_[24898]_  = A300 & A299;
  assign \new_[24899]_  = A236 & \new_[24898]_ ;
  assign \new_[24900]_  = \new_[24899]_  & \new_[24894]_ ;
  assign \new_[24903]_  = A167 & A170;
  assign \new_[24907]_  = ~A200 & ~A199;
  assign \new_[24908]_  = ~A166 & \new_[24907]_ ;
  assign \new_[24909]_  = \new_[24908]_  & \new_[24903]_ ;
  assign \new_[24913]_  = ~A233 & A232;
  assign \new_[24914]_  = ~A202 & \new_[24913]_ ;
  assign \new_[24918]_  = A300 & A298;
  assign \new_[24919]_  = A236 & \new_[24918]_ ;
  assign \new_[24920]_  = \new_[24919]_  & \new_[24914]_ ;
  assign \new_[24923]_  = A167 & A170;
  assign \new_[24927]_  = ~A200 & ~A199;
  assign \new_[24928]_  = ~A166 & \new_[24927]_ ;
  assign \new_[24929]_  = \new_[24928]_  & \new_[24923]_ ;
  assign \new_[24933]_  = ~A233 & A232;
  assign \new_[24934]_  = ~A202 & \new_[24933]_ ;
  assign \new_[24938]_  = A267 & A265;
  assign \new_[24939]_  = A236 & \new_[24938]_ ;
  assign \new_[24940]_  = \new_[24939]_  & \new_[24934]_ ;
  assign \new_[24943]_  = A167 & A170;
  assign \new_[24947]_  = ~A200 & ~A199;
  assign \new_[24948]_  = ~A166 & \new_[24947]_ ;
  assign \new_[24949]_  = \new_[24948]_  & \new_[24943]_ ;
  assign \new_[24953]_  = ~A233 & A232;
  assign \new_[24954]_  = ~A202 & \new_[24953]_ ;
  assign \new_[24958]_  = A267 & A266;
  assign \new_[24959]_  = A236 & \new_[24958]_ ;
  assign \new_[24960]_  = \new_[24959]_  & \new_[24954]_ ;
  assign \new_[24963]_  = ~A167 & A170;
  assign \new_[24967]_  = ~A202 & ~A201;
  assign \new_[24968]_  = A166 & \new_[24967]_ ;
  assign \new_[24969]_  = \new_[24968]_  & \new_[24963]_ ;
  assign \new_[24973]_  = A234 & A232;
  assign \new_[24974]_  = ~A203 & \new_[24973]_ ;
  assign \new_[24978]_  = A302 & ~A299;
  assign \new_[24979]_  = A298 & \new_[24978]_ ;
  assign \new_[24980]_  = \new_[24979]_  & \new_[24974]_ ;
  assign \new_[24983]_  = ~A167 & A170;
  assign \new_[24987]_  = ~A202 & ~A201;
  assign \new_[24988]_  = A166 & \new_[24987]_ ;
  assign \new_[24989]_  = \new_[24988]_  & \new_[24983]_ ;
  assign \new_[24993]_  = A234 & A232;
  assign \new_[24994]_  = ~A203 & \new_[24993]_ ;
  assign \new_[24998]_  = A302 & A299;
  assign \new_[24999]_  = ~A298 & \new_[24998]_ ;
  assign \new_[25000]_  = \new_[24999]_  & \new_[24994]_ ;
  assign \new_[25003]_  = ~A167 & A170;
  assign \new_[25007]_  = ~A202 & ~A201;
  assign \new_[25008]_  = A166 & \new_[25007]_ ;
  assign \new_[25009]_  = \new_[25008]_  & \new_[25003]_ ;
  assign \new_[25013]_  = A234 & A232;
  assign \new_[25014]_  = ~A203 & \new_[25013]_ ;
  assign \new_[25018]_  = A269 & A266;
  assign \new_[25019]_  = ~A265 & \new_[25018]_ ;
  assign \new_[25020]_  = \new_[25019]_  & \new_[25014]_ ;
  assign \new_[25023]_  = ~A167 & A170;
  assign \new_[25027]_  = ~A202 & ~A201;
  assign \new_[25028]_  = A166 & \new_[25027]_ ;
  assign \new_[25029]_  = \new_[25028]_  & \new_[25023]_ ;
  assign \new_[25033]_  = A234 & A232;
  assign \new_[25034]_  = ~A203 & \new_[25033]_ ;
  assign \new_[25038]_  = A269 & ~A266;
  assign \new_[25039]_  = A265 & \new_[25038]_ ;
  assign \new_[25040]_  = \new_[25039]_  & \new_[25034]_ ;
  assign \new_[25043]_  = ~A167 & A170;
  assign \new_[25047]_  = ~A202 & ~A201;
  assign \new_[25048]_  = A166 & \new_[25047]_ ;
  assign \new_[25049]_  = \new_[25048]_  & \new_[25043]_ ;
  assign \new_[25053]_  = A234 & A233;
  assign \new_[25054]_  = ~A203 & \new_[25053]_ ;
  assign \new_[25058]_  = A302 & ~A299;
  assign \new_[25059]_  = A298 & \new_[25058]_ ;
  assign \new_[25060]_  = \new_[25059]_  & \new_[25054]_ ;
  assign \new_[25063]_  = ~A167 & A170;
  assign \new_[25067]_  = ~A202 & ~A201;
  assign \new_[25068]_  = A166 & \new_[25067]_ ;
  assign \new_[25069]_  = \new_[25068]_  & \new_[25063]_ ;
  assign \new_[25073]_  = A234 & A233;
  assign \new_[25074]_  = ~A203 & \new_[25073]_ ;
  assign \new_[25078]_  = A302 & A299;
  assign \new_[25079]_  = ~A298 & \new_[25078]_ ;
  assign \new_[25080]_  = \new_[25079]_  & \new_[25074]_ ;
  assign \new_[25083]_  = ~A167 & A170;
  assign \new_[25087]_  = ~A202 & ~A201;
  assign \new_[25088]_  = A166 & \new_[25087]_ ;
  assign \new_[25089]_  = \new_[25088]_  & \new_[25083]_ ;
  assign \new_[25093]_  = A234 & A233;
  assign \new_[25094]_  = ~A203 & \new_[25093]_ ;
  assign \new_[25098]_  = A269 & A266;
  assign \new_[25099]_  = ~A265 & \new_[25098]_ ;
  assign \new_[25100]_  = \new_[25099]_  & \new_[25094]_ ;
  assign \new_[25103]_  = ~A167 & A170;
  assign \new_[25107]_  = ~A202 & ~A201;
  assign \new_[25108]_  = A166 & \new_[25107]_ ;
  assign \new_[25109]_  = \new_[25108]_  & \new_[25103]_ ;
  assign \new_[25113]_  = A234 & A233;
  assign \new_[25114]_  = ~A203 & \new_[25113]_ ;
  assign \new_[25118]_  = A269 & ~A266;
  assign \new_[25119]_  = A265 & \new_[25118]_ ;
  assign \new_[25120]_  = \new_[25119]_  & \new_[25114]_ ;
  assign \new_[25123]_  = ~A167 & A170;
  assign \new_[25127]_  = ~A202 & ~A201;
  assign \new_[25128]_  = A166 & \new_[25127]_ ;
  assign \new_[25129]_  = \new_[25128]_  & \new_[25123]_ ;
  assign \new_[25133]_  = A233 & ~A232;
  assign \new_[25134]_  = ~A203 & \new_[25133]_ ;
  assign \new_[25138]_  = A300 & A299;
  assign \new_[25139]_  = A236 & \new_[25138]_ ;
  assign \new_[25140]_  = \new_[25139]_  & \new_[25134]_ ;
  assign \new_[25143]_  = ~A167 & A170;
  assign \new_[25147]_  = ~A202 & ~A201;
  assign \new_[25148]_  = A166 & \new_[25147]_ ;
  assign \new_[25149]_  = \new_[25148]_  & \new_[25143]_ ;
  assign \new_[25153]_  = A233 & ~A232;
  assign \new_[25154]_  = ~A203 & \new_[25153]_ ;
  assign \new_[25158]_  = A300 & A298;
  assign \new_[25159]_  = A236 & \new_[25158]_ ;
  assign \new_[25160]_  = \new_[25159]_  & \new_[25154]_ ;
  assign \new_[25163]_  = ~A167 & A170;
  assign \new_[25167]_  = ~A202 & ~A201;
  assign \new_[25168]_  = A166 & \new_[25167]_ ;
  assign \new_[25169]_  = \new_[25168]_  & \new_[25163]_ ;
  assign \new_[25173]_  = A233 & ~A232;
  assign \new_[25174]_  = ~A203 & \new_[25173]_ ;
  assign \new_[25178]_  = A267 & A265;
  assign \new_[25179]_  = A236 & \new_[25178]_ ;
  assign \new_[25180]_  = \new_[25179]_  & \new_[25174]_ ;
  assign \new_[25183]_  = ~A167 & A170;
  assign \new_[25187]_  = ~A202 & ~A201;
  assign \new_[25188]_  = A166 & \new_[25187]_ ;
  assign \new_[25189]_  = \new_[25188]_  & \new_[25183]_ ;
  assign \new_[25193]_  = A233 & ~A232;
  assign \new_[25194]_  = ~A203 & \new_[25193]_ ;
  assign \new_[25198]_  = A267 & A266;
  assign \new_[25199]_  = A236 & \new_[25198]_ ;
  assign \new_[25200]_  = \new_[25199]_  & \new_[25194]_ ;
  assign \new_[25203]_  = ~A167 & A170;
  assign \new_[25207]_  = ~A202 & ~A201;
  assign \new_[25208]_  = A166 & \new_[25207]_ ;
  assign \new_[25209]_  = \new_[25208]_  & \new_[25203]_ ;
  assign \new_[25213]_  = ~A233 & A232;
  assign \new_[25214]_  = ~A203 & \new_[25213]_ ;
  assign \new_[25218]_  = A300 & A299;
  assign \new_[25219]_  = A236 & \new_[25218]_ ;
  assign \new_[25220]_  = \new_[25219]_  & \new_[25214]_ ;
  assign \new_[25223]_  = ~A167 & A170;
  assign \new_[25227]_  = ~A202 & ~A201;
  assign \new_[25228]_  = A166 & \new_[25227]_ ;
  assign \new_[25229]_  = \new_[25228]_  & \new_[25223]_ ;
  assign \new_[25233]_  = ~A233 & A232;
  assign \new_[25234]_  = ~A203 & \new_[25233]_ ;
  assign \new_[25238]_  = A300 & A298;
  assign \new_[25239]_  = A236 & \new_[25238]_ ;
  assign \new_[25240]_  = \new_[25239]_  & \new_[25234]_ ;
  assign \new_[25243]_  = ~A167 & A170;
  assign \new_[25247]_  = ~A202 & ~A201;
  assign \new_[25248]_  = A166 & \new_[25247]_ ;
  assign \new_[25249]_  = \new_[25248]_  & \new_[25243]_ ;
  assign \new_[25253]_  = ~A233 & A232;
  assign \new_[25254]_  = ~A203 & \new_[25253]_ ;
  assign \new_[25258]_  = A267 & A265;
  assign \new_[25259]_  = A236 & \new_[25258]_ ;
  assign \new_[25260]_  = \new_[25259]_  & \new_[25254]_ ;
  assign \new_[25263]_  = ~A167 & A170;
  assign \new_[25267]_  = ~A202 & ~A201;
  assign \new_[25268]_  = A166 & \new_[25267]_ ;
  assign \new_[25269]_  = \new_[25268]_  & \new_[25263]_ ;
  assign \new_[25273]_  = ~A233 & A232;
  assign \new_[25274]_  = ~A203 & \new_[25273]_ ;
  assign \new_[25278]_  = A267 & A266;
  assign \new_[25279]_  = A236 & \new_[25278]_ ;
  assign \new_[25280]_  = \new_[25279]_  & \new_[25274]_ ;
  assign \new_[25283]_  = ~A167 & A170;
  assign \new_[25287]_  = A200 & A199;
  assign \new_[25288]_  = A166 & \new_[25287]_ ;
  assign \new_[25289]_  = \new_[25288]_  & \new_[25283]_ ;
  assign \new_[25293]_  = A235 & ~A202;
  assign \new_[25294]_  = ~A201 & \new_[25293]_ ;
  assign \new_[25298]_  = A302 & ~A299;
  assign \new_[25299]_  = A298 & \new_[25298]_ ;
  assign \new_[25300]_  = \new_[25299]_  & \new_[25294]_ ;
  assign \new_[25303]_  = ~A167 & A170;
  assign \new_[25307]_  = A200 & A199;
  assign \new_[25308]_  = A166 & \new_[25307]_ ;
  assign \new_[25309]_  = \new_[25308]_  & \new_[25303]_ ;
  assign \new_[25313]_  = A235 & ~A202;
  assign \new_[25314]_  = ~A201 & \new_[25313]_ ;
  assign \new_[25318]_  = A302 & A299;
  assign \new_[25319]_  = ~A298 & \new_[25318]_ ;
  assign \new_[25320]_  = \new_[25319]_  & \new_[25314]_ ;
  assign \new_[25323]_  = ~A167 & A170;
  assign \new_[25327]_  = A200 & A199;
  assign \new_[25328]_  = A166 & \new_[25327]_ ;
  assign \new_[25329]_  = \new_[25328]_  & \new_[25323]_ ;
  assign \new_[25333]_  = A235 & ~A202;
  assign \new_[25334]_  = ~A201 & \new_[25333]_ ;
  assign \new_[25338]_  = A269 & A266;
  assign \new_[25339]_  = ~A265 & \new_[25338]_ ;
  assign \new_[25340]_  = \new_[25339]_  & \new_[25334]_ ;
  assign \new_[25343]_  = ~A167 & A170;
  assign \new_[25347]_  = A200 & A199;
  assign \new_[25348]_  = A166 & \new_[25347]_ ;
  assign \new_[25349]_  = \new_[25348]_  & \new_[25343]_ ;
  assign \new_[25353]_  = A235 & ~A202;
  assign \new_[25354]_  = ~A201 & \new_[25353]_ ;
  assign \new_[25358]_  = A269 & ~A266;
  assign \new_[25359]_  = A265 & \new_[25358]_ ;
  assign \new_[25360]_  = \new_[25359]_  & \new_[25354]_ ;
  assign \new_[25363]_  = ~A167 & A170;
  assign \new_[25367]_  = A200 & A199;
  assign \new_[25368]_  = A166 & \new_[25367]_ ;
  assign \new_[25369]_  = \new_[25368]_  & \new_[25363]_ ;
  assign \new_[25373]_  = A232 & ~A202;
  assign \new_[25374]_  = ~A201 & \new_[25373]_ ;
  assign \new_[25378]_  = A300 & A299;
  assign \new_[25379]_  = A234 & \new_[25378]_ ;
  assign \new_[25380]_  = \new_[25379]_  & \new_[25374]_ ;
  assign \new_[25383]_  = ~A167 & A170;
  assign \new_[25387]_  = A200 & A199;
  assign \new_[25388]_  = A166 & \new_[25387]_ ;
  assign \new_[25389]_  = \new_[25388]_  & \new_[25383]_ ;
  assign \new_[25393]_  = A232 & ~A202;
  assign \new_[25394]_  = ~A201 & \new_[25393]_ ;
  assign \new_[25398]_  = A300 & A298;
  assign \new_[25399]_  = A234 & \new_[25398]_ ;
  assign \new_[25400]_  = \new_[25399]_  & \new_[25394]_ ;
  assign \new_[25403]_  = ~A167 & A170;
  assign \new_[25407]_  = A200 & A199;
  assign \new_[25408]_  = A166 & \new_[25407]_ ;
  assign \new_[25409]_  = \new_[25408]_  & \new_[25403]_ ;
  assign \new_[25413]_  = A232 & ~A202;
  assign \new_[25414]_  = ~A201 & \new_[25413]_ ;
  assign \new_[25418]_  = A267 & A265;
  assign \new_[25419]_  = A234 & \new_[25418]_ ;
  assign \new_[25420]_  = \new_[25419]_  & \new_[25414]_ ;
  assign \new_[25423]_  = ~A167 & A170;
  assign \new_[25427]_  = A200 & A199;
  assign \new_[25428]_  = A166 & \new_[25427]_ ;
  assign \new_[25429]_  = \new_[25428]_  & \new_[25423]_ ;
  assign \new_[25433]_  = A232 & ~A202;
  assign \new_[25434]_  = ~A201 & \new_[25433]_ ;
  assign \new_[25438]_  = A267 & A266;
  assign \new_[25439]_  = A234 & \new_[25438]_ ;
  assign \new_[25440]_  = \new_[25439]_  & \new_[25434]_ ;
  assign \new_[25443]_  = ~A167 & A170;
  assign \new_[25447]_  = A200 & A199;
  assign \new_[25448]_  = A166 & \new_[25447]_ ;
  assign \new_[25449]_  = \new_[25448]_  & \new_[25443]_ ;
  assign \new_[25453]_  = A233 & ~A202;
  assign \new_[25454]_  = ~A201 & \new_[25453]_ ;
  assign \new_[25458]_  = A300 & A299;
  assign \new_[25459]_  = A234 & \new_[25458]_ ;
  assign \new_[25460]_  = \new_[25459]_  & \new_[25454]_ ;
  assign \new_[25463]_  = ~A167 & A170;
  assign \new_[25467]_  = A200 & A199;
  assign \new_[25468]_  = A166 & \new_[25467]_ ;
  assign \new_[25469]_  = \new_[25468]_  & \new_[25463]_ ;
  assign \new_[25473]_  = A233 & ~A202;
  assign \new_[25474]_  = ~A201 & \new_[25473]_ ;
  assign \new_[25478]_  = A300 & A298;
  assign \new_[25479]_  = A234 & \new_[25478]_ ;
  assign \new_[25480]_  = \new_[25479]_  & \new_[25474]_ ;
  assign \new_[25483]_  = ~A167 & A170;
  assign \new_[25487]_  = A200 & A199;
  assign \new_[25488]_  = A166 & \new_[25487]_ ;
  assign \new_[25489]_  = \new_[25488]_  & \new_[25483]_ ;
  assign \new_[25493]_  = A233 & ~A202;
  assign \new_[25494]_  = ~A201 & \new_[25493]_ ;
  assign \new_[25498]_  = A267 & A265;
  assign \new_[25499]_  = A234 & \new_[25498]_ ;
  assign \new_[25500]_  = \new_[25499]_  & \new_[25494]_ ;
  assign \new_[25503]_  = ~A167 & A170;
  assign \new_[25507]_  = A200 & A199;
  assign \new_[25508]_  = A166 & \new_[25507]_ ;
  assign \new_[25509]_  = \new_[25508]_  & \new_[25503]_ ;
  assign \new_[25513]_  = A233 & ~A202;
  assign \new_[25514]_  = ~A201 & \new_[25513]_ ;
  assign \new_[25518]_  = A267 & A266;
  assign \new_[25519]_  = A234 & \new_[25518]_ ;
  assign \new_[25520]_  = \new_[25519]_  & \new_[25514]_ ;
  assign \new_[25523]_  = ~A167 & A170;
  assign \new_[25527]_  = A200 & A199;
  assign \new_[25528]_  = A166 & \new_[25527]_ ;
  assign \new_[25529]_  = \new_[25528]_  & \new_[25523]_ ;
  assign \new_[25533]_  = ~A232 & ~A202;
  assign \new_[25534]_  = ~A201 & \new_[25533]_ ;
  assign \new_[25538]_  = A301 & A236;
  assign \new_[25539]_  = A233 & \new_[25538]_ ;
  assign \new_[25540]_  = \new_[25539]_  & \new_[25534]_ ;
  assign \new_[25543]_  = ~A167 & A170;
  assign \new_[25547]_  = A200 & A199;
  assign \new_[25548]_  = A166 & \new_[25547]_ ;
  assign \new_[25549]_  = \new_[25548]_  & \new_[25543]_ ;
  assign \new_[25553]_  = ~A232 & ~A202;
  assign \new_[25554]_  = ~A201 & \new_[25553]_ ;
  assign \new_[25558]_  = A268 & A236;
  assign \new_[25559]_  = A233 & \new_[25558]_ ;
  assign \new_[25560]_  = \new_[25559]_  & \new_[25554]_ ;
  assign \new_[25563]_  = ~A167 & A170;
  assign \new_[25567]_  = A200 & A199;
  assign \new_[25568]_  = A166 & \new_[25567]_ ;
  assign \new_[25569]_  = \new_[25568]_  & \new_[25563]_ ;
  assign \new_[25573]_  = A232 & ~A202;
  assign \new_[25574]_  = ~A201 & \new_[25573]_ ;
  assign \new_[25578]_  = A301 & A236;
  assign \new_[25579]_  = ~A233 & \new_[25578]_ ;
  assign \new_[25580]_  = \new_[25579]_  & \new_[25574]_ ;
  assign \new_[25583]_  = ~A167 & A170;
  assign \new_[25587]_  = A200 & A199;
  assign \new_[25588]_  = A166 & \new_[25587]_ ;
  assign \new_[25589]_  = \new_[25588]_  & \new_[25583]_ ;
  assign \new_[25593]_  = A232 & ~A202;
  assign \new_[25594]_  = ~A201 & \new_[25593]_ ;
  assign \new_[25598]_  = A268 & A236;
  assign \new_[25599]_  = ~A233 & \new_[25598]_ ;
  assign \new_[25600]_  = \new_[25599]_  & \new_[25594]_ ;
  assign \new_[25603]_  = ~A167 & A170;
  assign \new_[25607]_  = ~A200 & ~A199;
  assign \new_[25608]_  = A166 & \new_[25607]_ ;
  assign \new_[25609]_  = \new_[25608]_  & \new_[25603]_ ;
  assign \new_[25613]_  = A234 & A232;
  assign \new_[25614]_  = ~A202 & \new_[25613]_ ;
  assign \new_[25618]_  = A302 & ~A299;
  assign \new_[25619]_  = A298 & \new_[25618]_ ;
  assign \new_[25620]_  = \new_[25619]_  & \new_[25614]_ ;
  assign \new_[25623]_  = ~A167 & A170;
  assign \new_[25627]_  = ~A200 & ~A199;
  assign \new_[25628]_  = A166 & \new_[25627]_ ;
  assign \new_[25629]_  = \new_[25628]_  & \new_[25623]_ ;
  assign \new_[25633]_  = A234 & A232;
  assign \new_[25634]_  = ~A202 & \new_[25633]_ ;
  assign \new_[25638]_  = A302 & A299;
  assign \new_[25639]_  = ~A298 & \new_[25638]_ ;
  assign \new_[25640]_  = \new_[25639]_  & \new_[25634]_ ;
  assign \new_[25643]_  = ~A167 & A170;
  assign \new_[25647]_  = ~A200 & ~A199;
  assign \new_[25648]_  = A166 & \new_[25647]_ ;
  assign \new_[25649]_  = \new_[25648]_  & \new_[25643]_ ;
  assign \new_[25653]_  = A234 & A232;
  assign \new_[25654]_  = ~A202 & \new_[25653]_ ;
  assign \new_[25658]_  = A269 & A266;
  assign \new_[25659]_  = ~A265 & \new_[25658]_ ;
  assign \new_[25660]_  = \new_[25659]_  & \new_[25654]_ ;
  assign \new_[25663]_  = ~A167 & A170;
  assign \new_[25667]_  = ~A200 & ~A199;
  assign \new_[25668]_  = A166 & \new_[25667]_ ;
  assign \new_[25669]_  = \new_[25668]_  & \new_[25663]_ ;
  assign \new_[25673]_  = A234 & A232;
  assign \new_[25674]_  = ~A202 & \new_[25673]_ ;
  assign \new_[25678]_  = A269 & ~A266;
  assign \new_[25679]_  = A265 & \new_[25678]_ ;
  assign \new_[25680]_  = \new_[25679]_  & \new_[25674]_ ;
  assign \new_[25683]_  = ~A167 & A170;
  assign \new_[25687]_  = ~A200 & ~A199;
  assign \new_[25688]_  = A166 & \new_[25687]_ ;
  assign \new_[25689]_  = \new_[25688]_  & \new_[25683]_ ;
  assign \new_[25693]_  = A234 & A233;
  assign \new_[25694]_  = ~A202 & \new_[25693]_ ;
  assign \new_[25698]_  = A302 & ~A299;
  assign \new_[25699]_  = A298 & \new_[25698]_ ;
  assign \new_[25700]_  = \new_[25699]_  & \new_[25694]_ ;
  assign \new_[25703]_  = ~A167 & A170;
  assign \new_[25707]_  = ~A200 & ~A199;
  assign \new_[25708]_  = A166 & \new_[25707]_ ;
  assign \new_[25709]_  = \new_[25708]_  & \new_[25703]_ ;
  assign \new_[25713]_  = A234 & A233;
  assign \new_[25714]_  = ~A202 & \new_[25713]_ ;
  assign \new_[25718]_  = A302 & A299;
  assign \new_[25719]_  = ~A298 & \new_[25718]_ ;
  assign \new_[25720]_  = \new_[25719]_  & \new_[25714]_ ;
  assign \new_[25723]_  = ~A167 & A170;
  assign \new_[25727]_  = ~A200 & ~A199;
  assign \new_[25728]_  = A166 & \new_[25727]_ ;
  assign \new_[25729]_  = \new_[25728]_  & \new_[25723]_ ;
  assign \new_[25733]_  = A234 & A233;
  assign \new_[25734]_  = ~A202 & \new_[25733]_ ;
  assign \new_[25738]_  = A269 & A266;
  assign \new_[25739]_  = ~A265 & \new_[25738]_ ;
  assign \new_[25740]_  = \new_[25739]_  & \new_[25734]_ ;
  assign \new_[25743]_  = ~A167 & A170;
  assign \new_[25747]_  = ~A200 & ~A199;
  assign \new_[25748]_  = A166 & \new_[25747]_ ;
  assign \new_[25749]_  = \new_[25748]_  & \new_[25743]_ ;
  assign \new_[25753]_  = A234 & A233;
  assign \new_[25754]_  = ~A202 & \new_[25753]_ ;
  assign \new_[25758]_  = A269 & ~A266;
  assign \new_[25759]_  = A265 & \new_[25758]_ ;
  assign \new_[25760]_  = \new_[25759]_  & \new_[25754]_ ;
  assign \new_[25763]_  = ~A167 & A170;
  assign \new_[25767]_  = ~A200 & ~A199;
  assign \new_[25768]_  = A166 & \new_[25767]_ ;
  assign \new_[25769]_  = \new_[25768]_  & \new_[25763]_ ;
  assign \new_[25773]_  = A233 & ~A232;
  assign \new_[25774]_  = ~A202 & \new_[25773]_ ;
  assign \new_[25778]_  = A300 & A299;
  assign \new_[25779]_  = A236 & \new_[25778]_ ;
  assign \new_[25780]_  = \new_[25779]_  & \new_[25774]_ ;
  assign \new_[25783]_  = ~A167 & A170;
  assign \new_[25787]_  = ~A200 & ~A199;
  assign \new_[25788]_  = A166 & \new_[25787]_ ;
  assign \new_[25789]_  = \new_[25788]_  & \new_[25783]_ ;
  assign \new_[25793]_  = A233 & ~A232;
  assign \new_[25794]_  = ~A202 & \new_[25793]_ ;
  assign \new_[25798]_  = A300 & A298;
  assign \new_[25799]_  = A236 & \new_[25798]_ ;
  assign \new_[25800]_  = \new_[25799]_  & \new_[25794]_ ;
  assign \new_[25803]_  = ~A167 & A170;
  assign \new_[25807]_  = ~A200 & ~A199;
  assign \new_[25808]_  = A166 & \new_[25807]_ ;
  assign \new_[25809]_  = \new_[25808]_  & \new_[25803]_ ;
  assign \new_[25813]_  = A233 & ~A232;
  assign \new_[25814]_  = ~A202 & \new_[25813]_ ;
  assign \new_[25818]_  = A267 & A265;
  assign \new_[25819]_  = A236 & \new_[25818]_ ;
  assign \new_[25820]_  = \new_[25819]_  & \new_[25814]_ ;
  assign \new_[25823]_  = ~A167 & A170;
  assign \new_[25827]_  = ~A200 & ~A199;
  assign \new_[25828]_  = A166 & \new_[25827]_ ;
  assign \new_[25829]_  = \new_[25828]_  & \new_[25823]_ ;
  assign \new_[25833]_  = A233 & ~A232;
  assign \new_[25834]_  = ~A202 & \new_[25833]_ ;
  assign \new_[25838]_  = A267 & A266;
  assign \new_[25839]_  = A236 & \new_[25838]_ ;
  assign \new_[25840]_  = \new_[25839]_  & \new_[25834]_ ;
  assign \new_[25843]_  = ~A167 & A170;
  assign \new_[25847]_  = ~A200 & ~A199;
  assign \new_[25848]_  = A166 & \new_[25847]_ ;
  assign \new_[25849]_  = \new_[25848]_  & \new_[25843]_ ;
  assign \new_[25853]_  = ~A233 & A232;
  assign \new_[25854]_  = ~A202 & \new_[25853]_ ;
  assign \new_[25858]_  = A300 & A299;
  assign \new_[25859]_  = A236 & \new_[25858]_ ;
  assign \new_[25860]_  = \new_[25859]_  & \new_[25854]_ ;
  assign \new_[25863]_  = ~A167 & A170;
  assign \new_[25867]_  = ~A200 & ~A199;
  assign \new_[25868]_  = A166 & \new_[25867]_ ;
  assign \new_[25869]_  = \new_[25868]_  & \new_[25863]_ ;
  assign \new_[25873]_  = ~A233 & A232;
  assign \new_[25874]_  = ~A202 & \new_[25873]_ ;
  assign \new_[25878]_  = A300 & A298;
  assign \new_[25879]_  = A236 & \new_[25878]_ ;
  assign \new_[25880]_  = \new_[25879]_  & \new_[25874]_ ;
  assign \new_[25883]_  = ~A167 & A170;
  assign \new_[25887]_  = ~A200 & ~A199;
  assign \new_[25888]_  = A166 & \new_[25887]_ ;
  assign \new_[25889]_  = \new_[25888]_  & \new_[25883]_ ;
  assign \new_[25893]_  = ~A233 & A232;
  assign \new_[25894]_  = ~A202 & \new_[25893]_ ;
  assign \new_[25898]_  = A267 & A265;
  assign \new_[25899]_  = A236 & \new_[25898]_ ;
  assign \new_[25900]_  = \new_[25899]_  & \new_[25894]_ ;
  assign \new_[25903]_  = ~A167 & A170;
  assign \new_[25907]_  = ~A200 & ~A199;
  assign \new_[25908]_  = A166 & \new_[25907]_ ;
  assign \new_[25909]_  = \new_[25908]_  & \new_[25903]_ ;
  assign \new_[25913]_  = ~A233 & A232;
  assign \new_[25914]_  = ~A202 & \new_[25913]_ ;
  assign \new_[25918]_  = A267 & A266;
  assign \new_[25919]_  = A236 & \new_[25918]_ ;
  assign \new_[25920]_  = \new_[25919]_  & \new_[25914]_ ;
  assign \new_[25923]_  = A199 & A169;
  assign \new_[25927]_  = ~A202 & ~A201;
  assign \new_[25928]_  = A200 & \new_[25927]_ ;
  assign \new_[25929]_  = \new_[25928]_  & \new_[25923]_ ;
  assign \new_[25933]_  = A236 & A233;
  assign \new_[25934]_  = ~A232 & \new_[25933]_ ;
  assign \new_[25938]_  = A302 & ~A299;
  assign \new_[25939]_  = A298 & \new_[25938]_ ;
  assign \new_[25940]_  = \new_[25939]_  & \new_[25934]_ ;
  assign \new_[25943]_  = A199 & A169;
  assign \new_[25947]_  = ~A202 & ~A201;
  assign \new_[25948]_  = A200 & \new_[25947]_ ;
  assign \new_[25949]_  = \new_[25948]_  & \new_[25943]_ ;
  assign \new_[25953]_  = A236 & A233;
  assign \new_[25954]_  = ~A232 & \new_[25953]_ ;
  assign \new_[25958]_  = A302 & A299;
  assign \new_[25959]_  = ~A298 & \new_[25958]_ ;
  assign \new_[25960]_  = \new_[25959]_  & \new_[25954]_ ;
  assign \new_[25963]_  = A199 & A169;
  assign \new_[25967]_  = ~A202 & ~A201;
  assign \new_[25968]_  = A200 & \new_[25967]_ ;
  assign \new_[25969]_  = \new_[25968]_  & \new_[25963]_ ;
  assign \new_[25973]_  = A236 & A233;
  assign \new_[25974]_  = ~A232 & \new_[25973]_ ;
  assign \new_[25978]_  = A269 & A266;
  assign \new_[25979]_  = ~A265 & \new_[25978]_ ;
  assign \new_[25980]_  = \new_[25979]_  & \new_[25974]_ ;
  assign \new_[25983]_  = A199 & A169;
  assign \new_[25987]_  = ~A202 & ~A201;
  assign \new_[25988]_  = A200 & \new_[25987]_ ;
  assign \new_[25989]_  = \new_[25988]_  & \new_[25983]_ ;
  assign \new_[25993]_  = A236 & A233;
  assign \new_[25994]_  = ~A232 & \new_[25993]_ ;
  assign \new_[25998]_  = A269 & ~A266;
  assign \new_[25999]_  = A265 & \new_[25998]_ ;
  assign \new_[26000]_  = \new_[25999]_  & \new_[25994]_ ;
  assign \new_[26003]_  = A199 & A169;
  assign \new_[26007]_  = ~A202 & ~A201;
  assign \new_[26008]_  = A200 & \new_[26007]_ ;
  assign \new_[26009]_  = \new_[26008]_  & \new_[26003]_ ;
  assign \new_[26013]_  = A236 & ~A233;
  assign \new_[26014]_  = A232 & \new_[26013]_ ;
  assign \new_[26018]_  = A302 & ~A299;
  assign \new_[26019]_  = A298 & \new_[26018]_ ;
  assign \new_[26020]_  = \new_[26019]_  & \new_[26014]_ ;
  assign \new_[26023]_  = A199 & A169;
  assign \new_[26027]_  = ~A202 & ~A201;
  assign \new_[26028]_  = A200 & \new_[26027]_ ;
  assign \new_[26029]_  = \new_[26028]_  & \new_[26023]_ ;
  assign \new_[26033]_  = A236 & ~A233;
  assign \new_[26034]_  = A232 & \new_[26033]_ ;
  assign \new_[26038]_  = A302 & A299;
  assign \new_[26039]_  = ~A298 & \new_[26038]_ ;
  assign \new_[26040]_  = \new_[26039]_  & \new_[26034]_ ;
  assign \new_[26043]_  = A199 & A169;
  assign \new_[26047]_  = ~A202 & ~A201;
  assign \new_[26048]_  = A200 & \new_[26047]_ ;
  assign \new_[26049]_  = \new_[26048]_  & \new_[26043]_ ;
  assign \new_[26053]_  = A236 & ~A233;
  assign \new_[26054]_  = A232 & \new_[26053]_ ;
  assign \new_[26058]_  = A269 & A266;
  assign \new_[26059]_  = ~A265 & \new_[26058]_ ;
  assign \new_[26060]_  = \new_[26059]_  & \new_[26054]_ ;
  assign \new_[26063]_  = A199 & A169;
  assign \new_[26067]_  = ~A202 & ~A201;
  assign \new_[26068]_  = A200 & \new_[26067]_ ;
  assign \new_[26069]_  = \new_[26068]_  & \new_[26063]_ ;
  assign \new_[26073]_  = A236 & ~A233;
  assign \new_[26074]_  = A232 & \new_[26073]_ ;
  assign \new_[26078]_  = A269 & ~A266;
  assign \new_[26079]_  = A265 & \new_[26078]_ ;
  assign \new_[26080]_  = \new_[26079]_  & \new_[26074]_ ;
  assign \new_[26083]_  = ~A167 & ~A169;
  assign \new_[26087]_  = A201 & A199;
  assign \new_[26088]_  = ~A166 & \new_[26087]_ ;
  assign \new_[26089]_  = \new_[26088]_  & \new_[26083]_ ;
  assign \new_[26093]_  = A236 & A233;
  assign \new_[26094]_  = ~A232 & \new_[26093]_ ;
  assign \new_[26098]_  = A302 & ~A299;
  assign \new_[26099]_  = A298 & \new_[26098]_ ;
  assign \new_[26100]_  = \new_[26099]_  & \new_[26094]_ ;
  assign \new_[26103]_  = ~A167 & ~A169;
  assign \new_[26107]_  = A201 & A199;
  assign \new_[26108]_  = ~A166 & \new_[26107]_ ;
  assign \new_[26109]_  = \new_[26108]_  & \new_[26103]_ ;
  assign \new_[26113]_  = A236 & A233;
  assign \new_[26114]_  = ~A232 & \new_[26113]_ ;
  assign \new_[26118]_  = A302 & A299;
  assign \new_[26119]_  = ~A298 & \new_[26118]_ ;
  assign \new_[26120]_  = \new_[26119]_  & \new_[26114]_ ;
  assign \new_[26123]_  = ~A167 & ~A169;
  assign \new_[26127]_  = A201 & A199;
  assign \new_[26128]_  = ~A166 & \new_[26127]_ ;
  assign \new_[26129]_  = \new_[26128]_  & \new_[26123]_ ;
  assign \new_[26133]_  = A236 & A233;
  assign \new_[26134]_  = ~A232 & \new_[26133]_ ;
  assign \new_[26138]_  = A269 & A266;
  assign \new_[26139]_  = ~A265 & \new_[26138]_ ;
  assign \new_[26140]_  = \new_[26139]_  & \new_[26134]_ ;
  assign \new_[26143]_  = ~A167 & ~A169;
  assign \new_[26147]_  = A201 & A199;
  assign \new_[26148]_  = ~A166 & \new_[26147]_ ;
  assign \new_[26149]_  = \new_[26148]_  & \new_[26143]_ ;
  assign \new_[26153]_  = A236 & A233;
  assign \new_[26154]_  = ~A232 & \new_[26153]_ ;
  assign \new_[26158]_  = A269 & ~A266;
  assign \new_[26159]_  = A265 & \new_[26158]_ ;
  assign \new_[26160]_  = \new_[26159]_  & \new_[26154]_ ;
  assign \new_[26163]_  = ~A167 & ~A169;
  assign \new_[26167]_  = A201 & A199;
  assign \new_[26168]_  = ~A166 & \new_[26167]_ ;
  assign \new_[26169]_  = \new_[26168]_  & \new_[26163]_ ;
  assign \new_[26173]_  = A236 & ~A233;
  assign \new_[26174]_  = A232 & \new_[26173]_ ;
  assign \new_[26178]_  = A302 & ~A299;
  assign \new_[26179]_  = A298 & \new_[26178]_ ;
  assign \new_[26180]_  = \new_[26179]_  & \new_[26174]_ ;
  assign \new_[26183]_  = ~A167 & ~A169;
  assign \new_[26187]_  = A201 & A199;
  assign \new_[26188]_  = ~A166 & \new_[26187]_ ;
  assign \new_[26189]_  = \new_[26188]_  & \new_[26183]_ ;
  assign \new_[26193]_  = A236 & ~A233;
  assign \new_[26194]_  = A232 & \new_[26193]_ ;
  assign \new_[26198]_  = A302 & A299;
  assign \new_[26199]_  = ~A298 & \new_[26198]_ ;
  assign \new_[26200]_  = \new_[26199]_  & \new_[26194]_ ;
  assign \new_[26203]_  = ~A167 & ~A169;
  assign \new_[26207]_  = A201 & A199;
  assign \new_[26208]_  = ~A166 & \new_[26207]_ ;
  assign \new_[26209]_  = \new_[26208]_  & \new_[26203]_ ;
  assign \new_[26213]_  = A236 & ~A233;
  assign \new_[26214]_  = A232 & \new_[26213]_ ;
  assign \new_[26218]_  = A269 & A266;
  assign \new_[26219]_  = ~A265 & \new_[26218]_ ;
  assign \new_[26220]_  = \new_[26219]_  & \new_[26214]_ ;
  assign \new_[26223]_  = ~A167 & ~A169;
  assign \new_[26227]_  = A201 & A199;
  assign \new_[26228]_  = ~A166 & \new_[26227]_ ;
  assign \new_[26229]_  = \new_[26228]_  & \new_[26223]_ ;
  assign \new_[26233]_  = A236 & ~A233;
  assign \new_[26234]_  = A232 & \new_[26233]_ ;
  assign \new_[26238]_  = A269 & ~A266;
  assign \new_[26239]_  = A265 & \new_[26238]_ ;
  assign \new_[26240]_  = \new_[26239]_  & \new_[26234]_ ;
  assign \new_[26243]_  = ~A167 & ~A169;
  assign \new_[26247]_  = A201 & A200;
  assign \new_[26248]_  = ~A166 & \new_[26247]_ ;
  assign \new_[26249]_  = \new_[26248]_  & \new_[26243]_ ;
  assign \new_[26253]_  = A236 & A233;
  assign \new_[26254]_  = ~A232 & \new_[26253]_ ;
  assign \new_[26258]_  = A302 & ~A299;
  assign \new_[26259]_  = A298 & \new_[26258]_ ;
  assign \new_[26260]_  = \new_[26259]_  & \new_[26254]_ ;
  assign \new_[26263]_  = ~A167 & ~A169;
  assign \new_[26267]_  = A201 & A200;
  assign \new_[26268]_  = ~A166 & \new_[26267]_ ;
  assign \new_[26269]_  = \new_[26268]_  & \new_[26263]_ ;
  assign \new_[26273]_  = A236 & A233;
  assign \new_[26274]_  = ~A232 & \new_[26273]_ ;
  assign \new_[26278]_  = A302 & A299;
  assign \new_[26279]_  = ~A298 & \new_[26278]_ ;
  assign \new_[26280]_  = \new_[26279]_  & \new_[26274]_ ;
  assign \new_[26283]_  = ~A167 & ~A169;
  assign \new_[26287]_  = A201 & A200;
  assign \new_[26288]_  = ~A166 & \new_[26287]_ ;
  assign \new_[26289]_  = \new_[26288]_  & \new_[26283]_ ;
  assign \new_[26293]_  = A236 & A233;
  assign \new_[26294]_  = ~A232 & \new_[26293]_ ;
  assign \new_[26298]_  = A269 & A266;
  assign \new_[26299]_  = ~A265 & \new_[26298]_ ;
  assign \new_[26300]_  = \new_[26299]_  & \new_[26294]_ ;
  assign \new_[26303]_  = ~A167 & ~A169;
  assign \new_[26307]_  = A201 & A200;
  assign \new_[26308]_  = ~A166 & \new_[26307]_ ;
  assign \new_[26309]_  = \new_[26308]_  & \new_[26303]_ ;
  assign \new_[26313]_  = A236 & A233;
  assign \new_[26314]_  = ~A232 & \new_[26313]_ ;
  assign \new_[26318]_  = A269 & ~A266;
  assign \new_[26319]_  = A265 & \new_[26318]_ ;
  assign \new_[26320]_  = \new_[26319]_  & \new_[26314]_ ;
  assign \new_[26323]_  = ~A167 & ~A169;
  assign \new_[26327]_  = A201 & A200;
  assign \new_[26328]_  = ~A166 & \new_[26327]_ ;
  assign \new_[26329]_  = \new_[26328]_  & \new_[26323]_ ;
  assign \new_[26333]_  = A236 & ~A233;
  assign \new_[26334]_  = A232 & \new_[26333]_ ;
  assign \new_[26338]_  = A302 & ~A299;
  assign \new_[26339]_  = A298 & \new_[26338]_ ;
  assign \new_[26340]_  = \new_[26339]_  & \new_[26334]_ ;
  assign \new_[26343]_  = ~A167 & ~A169;
  assign \new_[26347]_  = A201 & A200;
  assign \new_[26348]_  = ~A166 & \new_[26347]_ ;
  assign \new_[26349]_  = \new_[26348]_  & \new_[26343]_ ;
  assign \new_[26353]_  = A236 & ~A233;
  assign \new_[26354]_  = A232 & \new_[26353]_ ;
  assign \new_[26358]_  = A302 & A299;
  assign \new_[26359]_  = ~A298 & \new_[26358]_ ;
  assign \new_[26360]_  = \new_[26359]_  & \new_[26354]_ ;
  assign \new_[26363]_  = ~A167 & ~A169;
  assign \new_[26367]_  = A201 & A200;
  assign \new_[26368]_  = ~A166 & \new_[26367]_ ;
  assign \new_[26369]_  = \new_[26368]_  & \new_[26363]_ ;
  assign \new_[26373]_  = A236 & ~A233;
  assign \new_[26374]_  = A232 & \new_[26373]_ ;
  assign \new_[26378]_  = A269 & A266;
  assign \new_[26379]_  = ~A265 & \new_[26378]_ ;
  assign \new_[26380]_  = \new_[26379]_  & \new_[26374]_ ;
  assign \new_[26383]_  = ~A167 & ~A169;
  assign \new_[26387]_  = A201 & A200;
  assign \new_[26388]_  = ~A166 & \new_[26387]_ ;
  assign \new_[26389]_  = \new_[26388]_  & \new_[26383]_ ;
  assign \new_[26393]_  = A236 & ~A233;
  assign \new_[26394]_  = A232 & \new_[26393]_ ;
  assign \new_[26398]_  = A269 & ~A266;
  assign \new_[26399]_  = A265 & \new_[26398]_ ;
  assign \new_[26400]_  = \new_[26399]_  & \new_[26394]_ ;
  assign \new_[26403]_  = ~A167 & ~A169;
  assign \new_[26407]_  = A200 & ~A199;
  assign \new_[26408]_  = ~A166 & \new_[26407]_ ;
  assign \new_[26409]_  = \new_[26408]_  & \new_[26403]_ ;
  assign \new_[26413]_  = A234 & A232;
  assign \new_[26414]_  = A203 & \new_[26413]_ ;
  assign \new_[26418]_  = A302 & ~A299;
  assign \new_[26419]_  = A298 & \new_[26418]_ ;
  assign \new_[26420]_  = \new_[26419]_  & \new_[26414]_ ;
  assign \new_[26423]_  = ~A167 & ~A169;
  assign \new_[26427]_  = A200 & ~A199;
  assign \new_[26428]_  = ~A166 & \new_[26427]_ ;
  assign \new_[26429]_  = \new_[26428]_  & \new_[26423]_ ;
  assign \new_[26433]_  = A234 & A232;
  assign \new_[26434]_  = A203 & \new_[26433]_ ;
  assign \new_[26438]_  = A302 & A299;
  assign \new_[26439]_  = ~A298 & \new_[26438]_ ;
  assign \new_[26440]_  = \new_[26439]_  & \new_[26434]_ ;
  assign \new_[26443]_  = ~A167 & ~A169;
  assign \new_[26447]_  = A200 & ~A199;
  assign \new_[26448]_  = ~A166 & \new_[26447]_ ;
  assign \new_[26449]_  = \new_[26448]_  & \new_[26443]_ ;
  assign \new_[26453]_  = A234 & A232;
  assign \new_[26454]_  = A203 & \new_[26453]_ ;
  assign \new_[26458]_  = A269 & A266;
  assign \new_[26459]_  = ~A265 & \new_[26458]_ ;
  assign \new_[26460]_  = \new_[26459]_  & \new_[26454]_ ;
  assign \new_[26463]_  = ~A167 & ~A169;
  assign \new_[26467]_  = A200 & ~A199;
  assign \new_[26468]_  = ~A166 & \new_[26467]_ ;
  assign \new_[26469]_  = \new_[26468]_  & \new_[26463]_ ;
  assign \new_[26473]_  = A234 & A232;
  assign \new_[26474]_  = A203 & \new_[26473]_ ;
  assign \new_[26478]_  = A269 & ~A266;
  assign \new_[26479]_  = A265 & \new_[26478]_ ;
  assign \new_[26480]_  = \new_[26479]_  & \new_[26474]_ ;
  assign \new_[26483]_  = ~A167 & ~A169;
  assign \new_[26487]_  = A200 & ~A199;
  assign \new_[26488]_  = ~A166 & \new_[26487]_ ;
  assign \new_[26489]_  = \new_[26488]_  & \new_[26483]_ ;
  assign \new_[26493]_  = A234 & A233;
  assign \new_[26494]_  = A203 & \new_[26493]_ ;
  assign \new_[26498]_  = A302 & ~A299;
  assign \new_[26499]_  = A298 & \new_[26498]_ ;
  assign \new_[26500]_  = \new_[26499]_  & \new_[26494]_ ;
  assign \new_[26503]_  = ~A167 & ~A169;
  assign \new_[26507]_  = A200 & ~A199;
  assign \new_[26508]_  = ~A166 & \new_[26507]_ ;
  assign \new_[26509]_  = \new_[26508]_  & \new_[26503]_ ;
  assign \new_[26513]_  = A234 & A233;
  assign \new_[26514]_  = A203 & \new_[26513]_ ;
  assign \new_[26518]_  = A302 & A299;
  assign \new_[26519]_  = ~A298 & \new_[26518]_ ;
  assign \new_[26520]_  = \new_[26519]_  & \new_[26514]_ ;
  assign \new_[26523]_  = ~A167 & ~A169;
  assign \new_[26527]_  = A200 & ~A199;
  assign \new_[26528]_  = ~A166 & \new_[26527]_ ;
  assign \new_[26529]_  = \new_[26528]_  & \new_[26523]_ ;
  assign \new_[26533]_  = A234 & A233;
  assign \new_[26534]_  = A203 & \new_[26533]_ ;
  assign \new_[26538]_  = A269 & A266;
  assign \new_[26539]_  = ~A265 & \new_[26538]_ ;
  assign \new_[26540]_  = \new_[26539]_  & \new_[26534]_ ;
  assign \new_[26543]_  = ~A167 & ~A169;
  assign \new_[26547]_  = A200 & ~A199;
  assign \new_[26548]_  = ~A166 & \new_[26547]_ ;
  assign \new_[26549]_  = \new_[26548]_  & \new_[26543]_ ;
  assign \new_[26553]_  = A234 & A233;
  assign \new_[26554]_  = A203 & \new_[26553]_ ;
  assign \new_[26558]_  = A269 & ~A266;
  assign \new_[26559]_  = A265 & \new_[26558]_ ;
  assign \new_[26560]_  = \new_[26559]_  & \new_[26554]_ ;
  assign \new_[26563]_  = ~A167 & ~A169;
  assign \new_[26567]_  = A200 & ~A199;
  assign \new_[26568]_  = ~A166 & \new_[26567]_ ;
  assign \new_[26569]_  = \new_[26568]_  & \new_[26563]_ ;
  assign \new_[26573]_  = A233 & ~A232;
  assign \new_[26574]_  = A203 & \new_[26573]_ ;
  assign \new_[26578]_  = A300 & A299;
  assign \new_[26579]_  = A236 & \new_[26578]_ ;
  assign \new_[26580]_  = \new_[26579]_  & \new_[26574]_ ;
  assign \new_[26583]_  = ~A167 & ~A169;
  assign \new_[26587]_  = A200 & ~A199;
  assign \new_[26588]_  = ~A166 & \new_[26587]_ ;
  assign \new_[26589]_  = \new_[26588]_  & \new_[26583]_ ;
  assign \new_[26593]_  = A233 & ~A232;
  assign \new_[26594]_  = A203 & \new_[26593]_ ;
  assign \new_[26598]_  = A300 & A298;
  assign \new_[26599]_  = A236 & \new_[26598]_ ;
  assign \new_[26600]_  = \new_[26599]_  & \new_[26594]_ ;
  assign \new_[26603]_  = ~A167 & ~A169;
  assign \new_[26607]_  = A200 & ~A199;
  assign \new_[26608]_  = ~A166 & \new_[26607]_ ;
  assign \new_[26609]_  = \new_[26608]_  & \new_[26603]_ ;
  assign \new_[26613]_  = A233 & ~A232;
  assign \new_[26614]_  = A203 & \new_[26613]_ ;
  assign \new_[26618]_  = A267 & A265;
  assign \new_[26619]_  = A236 & \new_[26618]_ ;
  assign \new_[26620]_  = \new_[26619]_  & \new_[26614]_ ;
  assign \new_[26623]_  = ~A167 & ~A169;
  assign \new_[26627]_  = A200 & ~A199;
  assign \new_[26628]_  = ~A166 & \new_[26627]_ ;
  assign \new_[26629]_  = \new_[26628]_  & \new_[26623]_ ;
  assign \new_[26633]_  = A233 & ~A232;
  assign \new_[26634]_  = A203 & \new_[26633]_ ;
  assign \new_[26638]_  = A267 & A266;
  assign \new_[26639]_  = A236 & \new_[26638]_ ;
  assign \new_[26640]_  = \new_[26639]_  & \new_[26634]_ ;
  assign \new_[26643]_  = ~A167 & ~A169;
  assign \new_[26647]_  = A200 & ~A199;
  assign \new_[26648]_  = ~A166 & \new_[26647]_ ;
  assign \new_[26649]_  = \new_[26648]_  & \new_[26643]_ ;
  assign \new_[26653]_  = ~A233 & A232;
  assign \new_[26654]_  = A203 & \new_[26653]_ ;
  assign \new_[26658]_  = A300 & A299;
  assign \new_[26659]_  = A236 & \new_[26658]_ ;
  assign \new_[26660]_  = \new_[26659]_  & \new_[26654]_ ;
  assign \new_[26663]_  = ~A167 & ~A169;
  assign \new_[26667]_  = A200 & ~A199;
  assign \new_[26668]_  = ~A166 & \new_[26667]_ ;
  assign \new_[26669]_  = \new_[26668]_  & \new_[26663]_ ;
  assign \new_[26673]_  = ~A233 & A232;
  assign \new_[26674]_  = A203 & \new_[26673]_ ;
  assign \new_[26678]_  = A300 & A298;
  assign \new_[26679]_  = A236 & \new_[26678]_ ;
  assign \new_[26680]_  = \new_[26679]_  & \new_[26674]_ ;
  assign \new_[26683]_  = ~A167 & ~A169;
  assign \new_[26687]_  = A200 & ~A199;
  assign \new_[26688]_  = ~A166 & \new_[26687]_ ;
  assign \new_[26689]_  = \new_[26688]_  & \new_[26683]_ ;
  assign \new_[26693]_  = ~A233 & A232;
  assign \new_[26694]_  = A203 & \new_[26693]_ ;
  assign \new_[26698]_  = A267 & A265;
  assign \new_[26699]_  = A236 & \new_[26698]_ ;
  assign \new_[26700]_  = \new_[26699]_  & \new_[26694]_ ;
  assign \new_[26703]_  = ~A167 & ~A169;
  assign \new_[26707]_  = A200 & ~A199;
  assign \new_[26708]_  = ~A166 & \new_[26707]_ ;
  assign \new_[26709]_  = \new_[26708]_  & \new_[26703]_ ;
  assign \new_[26713]_  = ~A233 & A232;
  assign \new_[26714]_  = A203 & \new_[26713]_ ;
  assign \new_[26718]_  = A267 & A266;
  assign \new_[26719]_  = A236 & \new_[26718]_ ;
  assign \new_[26720]_  = \new_[26719]_  & \new_[26714]_ ;
  assign \new_[26723]_  = ~A167 & ~A169;
  assign \new_[26727]_  = ~A200 & A199;
  assign \new_[26728]_  = ~A166 & \new_[26727]_ ;
  assign \new_[26729]_  = \new_[26728]_  & \new_[26723]_ ;
  assign \new_[26733]_  = A234 & A232;
  assign \new_[26734]_  = A203 & \new_[26733]_ ;
  assign \new_[26738]_  = A302 & ~A299;
  assign \new_[26739]_  = A298 & \new_[26738]_ ;
  assign \new_[26740]_  = \new_[26739]_  & \new_[26734]_ ;
  assign \new_[26743]_  = ~A167 & ~A169;
  assign \new_[26747]_  = ~A200 & A199;
  assign \new_[26748]_  = ~A166 & \new_[26747]_ ;
  assign \new_[26749]_  = \new_[26748]_  & \new_[26743]_ ;
  assign \new_[26753]_  = A234 & A232;
  assign \new_[26754]_  = A203 & \new_[26753]_ ;
  assign \new_[26758]_  = A302 & A299;
  assign \new_[26759]_  = ~A298 & \new_[26758]_ ;
  assign \new_[26760]_  = \new_[26759]_  & \new_[26754]_ ;
  assign \new_[26763]_  = ~A167 & ~A169;
  assign \new_[26767]_  = ~A200 & A199;
  assign \new_[26768]_  = ~A166 & \new_[26767]_ ;
  assign \new_[26769]_  = \new_[26768]_  & \new_[26763]_ ;
  assign \new_[26773]_  = A234 & A232;
  assign \new_[26774]_  = A203 & \new_[26773]_ ;
  assign \new_[26778]_  = A269 & A266;
  assign \new_[26779]_  = ~A265 & \new_[26778]_ ;
  assign \new_[26780]_  = \new_[26779]_  & \new_[26774]_ ;
  assign \new_[26783]_  = ~A167 & ~A169;
  assign \new_[26787]_  = ~A200 & A199;
  assign \new_[26788]_  = ~A166 & \new_[26787]_ ;
  assign \new_[26789]_  = \new_[26788]_  & \new_[26783]_ ;
  assign \new_[26793]_  = A234 & A232;
  assign \new_[26794]_  = A203 & \new_[26793]_ ;
  assign \new_[26798]_  = A269 & ~A266;
  assign \new_[26799]_  = A265 & \new_[26798]_ ;
  assign \new_[26800]_  = \new_[26799]_  & \new_[26794]_ ;
  assign \new_[26803]_  = ~A167 & ~A169;
  assign \new_[26807]_  = ~A200 & A199;
  assign \new_[26808]_  = ~A166 & \new_[26807]_ ;
  assign \new_[26809]_  = \new_[26808]_  & \new_[26803]_ ;
  assign \new_[26813]_  = A234 & A233;
  assign \new_[26814]_  = A203 & \new_[26813]_ ;
  assign \new_[26818]_  = A302 & ~A299;
  assign \new_[26819]_  = A298 & \new_[26818]_ ;
  assign \new_[26820]_  = \new_[26819]_  & \new_[26814]_ ;
  assign \new_[26823]_  = ~A167 & ~A169;
  assign \new_[26827]_  = ~A200 & A199;
  assign \new_[26828]_  = ~A166 & \new_[26827]_ ;
  assign \new_[26829]_  = \new_[26828]_  & \new_[26823]_ ;
  assign \new_[26833]_  = A234 & A233;
  assign \new_[26834]_  = A203 & \new_[26833]_ ;
  assign \new_[26838]_  = A302 & A299;
  assign \new_[26839]_  = ~A298 & \new_[26838]_ ;
  assign \new_[26840]_  = \new_[26839]_  & \new_[26834]_ ;
  assign \new_[26843]_  = ~A167 & ~A169;
  assign \new_[26847]_  = ~A200 & A199;
  assign \new_[26848]_  = ~A166 & \new_[26847]_ ;
  assign \new_[26849]_  = \new_[26848]_  & \new_[26843]_ ;
  assign \new_[26853]_  = A234 & A233;
  assign \new_[26854]_  = A203 & \new_[26853]_ ;
  assign \new_[26858]_  = A269 & A266;
  assign \new_[26859]_  = ~A265 & \new_[26858]_ ;
  assign \new_[26860]_  = \new_[26859]_  & \new_[26854]_ ;
  assign \new_[26863]_  = ~A167 & ~A169;
  assign \new_[26867]_  = ~A200 & A199;
  assign \new_[26868]_  = ~A166 & \new_[26867]_ ;
  assign \new_[26869]_  = \new_[26868]_  & \new_[26863]_ ;
  assign \new_[26873]_  = A234 & A233;
  assign \new_[26874]_  = A203 & \new_[26873]_ ;
  assign \new_[26878]_  = A269 & ~A266;
  assign \new_[26879]_  = A265 & \new_[26878]_ ;
  assign \new_[26880]_  = \new_[26879]_  & \new_[26874]_ ;
  assign \new_[26883]_  = ~A167 & ~A169;
  assign \new_[26887]_  = ~A200 & A199;
  assign \new_[26888]_  = ~A166 & \new_[26887]_ ;
  assign \new_[26889]_  = \new_[26888]_  & \new_[26883]_ ;
  assign \new_[26893]_  = A233 & ~A232;
  assign \new_[26894]_  = A203 & \new_[26893]_ ;
  assign \new_[26898]_  = A300 & A299;
  assign \new_[26899]_  = A236 & \new_[26898]_ ;
  assign \new_[26900]_  = \new_[26899]_  & \new_[26894]_ ;
  assign \new_[26903]_  = ~A167 & ~A169;
  assign \new_[26907]_  = ~A200 & A199;
  assign \new_[26908]_  = ~A166 & \new_[26907]_ ;
  assign \new_[26909]_  = \new_[26908]_  & \new_[26903]_ ;
  assign \new_[26913]_  = A233 & ~A232;
  assign \new_[26914]_  = A203 & \new_[26913]_ ;
  assign \new_[26918]_  = A300 & A298;
  assign \new_[26919]_  = A236 & \new_[26918]_ ;
  assign \new_[26920]_  = \new_[26919]_  & \new_[26914]_ ;
  assign \new_[26923]_  = ~A167 & ~A169;
  assign \new_[26927]_  = ~A200 & A199;
  assign \new_[26928]_  = ~A166 & \new_[26927]_ ;
  assign \new_[26929]_  = \new_[26928]_  & \new_[26923]_ ;
  assign \new_[26933]_  = A233 & ~A232;
  assign \new_[26934]_  = A203 & \new_[26933]_ ;
  assign \new_[26938]_  = A267 & A265;
  assign \new_[26939]_  = A236 & \new_[26938]_ ;
  assign \new_[26940]_  = \new_[26939]_  & \new_[26934]_ ;
  assign \new_[26943]_  = ~A167 & ~A169;
  assign \new_[26947]_  = ~A200 & A199;
  assign \new_[26948]_  = ~A166 & \new_[26947]_ ;
  assign \new_[26949]_  = \new_[26948]_  & \new_[26943]_ ;
  assign \new_[26953]_  = A233 & ~A232;
  assign \new_[26954]_  = A203 & \new_[26953]_ ;
  assign \new_[26958]_  = A267 & A266;
  assign \new_[26959]_  = A236 & \new_[26958]_ ;
  assign \new_[26960]_  = \new_[26959]_  & \new_[26954]_ ;
  assign \new_[26963]_  = ~A167 & ~A169;
  assign \new_[26967]_  = ~A200 & A199;
  assign \new_[26968]_  = ~A166 & \new_[26967]_ ;
  assign \new_[26969]_  = \new_[26968]_  & \new_[26963]_ ;
  assign \new_[26973]_  = ~A233 & A232;
  assign \new_[26974]_  = A203 & \new_[26973]_ ;
  assign \new_[26978]_  = A300 & A299;
  assign \new_[26979]_  = A236 & \new_[26978]_ ;
  assign \new_[26980]_  = \new_[26979]_  & \new_[26974]_ ;
  assign \new_[26983]_  = ~A167 & ~A169;
  assign \new_[26987]_  = ~A200 & A199;
  assign \new_[26988]_  = ~A166 & \new_[26987]_ ;
  assign \new_[26989]_  = \new_[26988]_  & \new_[26983]_ ;
  assign \new_[26993]_  = ~A233 & A232;
  assign \new_[26994]_  = A203 & \new_[26993]_ ;
  assign \new_[26998]_  = A300 & A298;
  assign \new_[26999]_  = A236 & \new_[26998]_ ;
  assign \new_[27000]_  = \new_[26999]_  & \new_[26994]_ ;
  assign \new_[27003]_  = ~A167 & ~A169;
  assign \new_[27007]_  = ~A200 & A199;
  assign \new_[27008]_  = ~A166 & \new_[27007]_ ;
  assign \new_[27009]_  = \new_[27008]_  & \new_[27003]_ ;
  assign \new_[27013]_  = ~A233 & A232;
  assign \new_[27014]_  = A203 & \new_[27013]_ ;
  assign \new_[27018]_  = A267 & A265;
  assign \new_[27019]_  = A236 & \new_[27018]_ ;
  assign \new_[27020]_  = \new_[27019]_  & \new_[27014]_ ;
  assign \new_[27023]_  = ~A167 & ~A169;
  assign \new_[27027]_  = ~A200 & A199;
  assign \new_[27028]_  = ~A166 & \new_[27027]_ ;
  assign \new_[27029]_  = \new_[27028]_  & \new_[27023]_ ;
  assign \new_[27033]_  = ~A233 & A232;
  assign \new_[27034]_  = A203 & \new_[27033]_ ;
  assign \new_[27038]_  = A267 & A266;
  assign \new_[27039]_  = A236 & \new_[27038]_ ;
  assign \new_[27040]_  = \new_[27039]_  & \new_[27034]_ ;
  assign \new_[27043]_  = ~A168 & ~A169;
  assign \new_[27047]_  = A202 & A166;
  assign \new_[27048]_  = A167 & \new_[27047]_ ;
  assign \new_[27049]_  = \new_[27048]_  & \new_[27043]_ ;
  assign \new_[27053]_  = A236 & A233;
  assign \new_[27054]_  = ~A232 & \new_[27053]_ ;
  assign \new_[27058]_  = A302 & ~A299;
  assign \new_[27059]_  = A298 & \new_[27058]_ ;
  assign \new_[27060]_  = \new_[27059]_  & \new_[27054]_ ;
  assign \new_[27063]_  = ~A168 & ~A169;
  assign \new_[27067]_  = A202 & A166;
  assign \new_[27068]_  = A167 & \new_[27067]_ ;
  assign \new_[27069]_  = \new_[27068]_  & \new_[27063]_ ;
  assign \new_[27073]_  = A236 & A233;
  assign \new_[27074]_  = ~A232 & \new_[27073]_ ;
  assign \new_[27078]_  = A302 & A299;
  assign \new_[27079]_  = ~A298 & \new_[27078]_ ;
  assign \new_[27080]_  = \new_[27079]_  & \new_[27074]_ ;
  assign \new_[27083]_  = ~A168 & ~A169;
  assign \new_[27087]_  = A202 & A166;
  assign \new_[27088]_  = A167 & \new_[27087]_ ;
  assign \new_[27089]_  = \new_[27088]_  & \new_[27083]_ ;
  assign \new_[27093]_  = A236 & A233;
  assign \new_[27094]_  = ~A232 & \new_[27093]_ ;
  assign \new_[27098]_  = A269 & A266;
  assign \new_[27099]_  = ~A265 & \new_[27098]_ ;
  assign \new_[27100]_  = \new_[27099]_  & \new_[27094]_ ;
  assign \new_[27103]_  = ~A168 & ~A169;
  assign \new_[27107]_  = A202 & A166;
  assign \new_[27108]_  = A167 & \new_[27107]_ ;
  assign \new_[27109]_  = \new_[27108]_  & \new_[27103]_ ;
  assign \new_[27113]_  = A236 & A233;
  assign \new_[27114]_  = ~A232 & \new_[27113]_ ;
  assign \new_[27118]_  = A269 & ~A266;
  assign \new_[27119]_  = A265 & \new_[27118]_ ;
  assign \new_[27120]_  = \new_[27119]_  & \new_[27114]_ ;
  assign \new_[27123]_  = ~A168 & ~A169;
  assign \new_[27127]_  = A202 & A166;
  assign \new_[27128]_  = A167 & \new_[27127]_ ;
  assign \new_[27129]_  = \new_[27128]_  & \new_[27123]_ ;
  assign \new_[27133]_  = A236 & ~A233;
  assign \new_[27134]_  = A232 & \new_[27133]_ ;
  assign \new_[27138]_  = A302 & ~A299;
  assign \new_[27139]_  = A298 & \new_[27138]_ ;
  assign \new_[27140]_  = \new_[27139]_  & \new_[27134]_ ;
  assign \new_[27143]_  = ~A168 & ~A169;
  assign \new_[27147]_  = A202 & A166;
  assign \new_[27148]_  = A167 & \new_[27147]_ ;
  assign \new_[27149]_  = \new_[27148]_  & \new_[27143]_ ;
  assign \new_[27153]_  = A236 & ~A233;
  assign \new_[27154]_  = A232 & \new_[27153]_ ;
  assign \new_[27158]_  = A302 & A299;
  assign \new_[27159]_  = ~A298 & \new_[27158]_ ;
  assign \new_[27160]_  = \new_[27159]_  & \new_[27154]_ ;
  assign \new_[27163]_  = ~A168 & ~A169;
  assign \new_[27167]_  = A202 & A166;
  assign \new_[27168]_  = A167 & \new_[27167]_ ;
  assign \new_[27169]_  = \new_[27168]_  & \new_[27163]_ ;
  assign \new_[27173]_  = A236 & ~A233;
  assign \new_[27174]_  = A232 & \new_[27173]_ ;
  assign \new_[27178]_  = A269 & A266;
  assign \new_[27179]_  = ~A265 & \new_[27178]_ ;
  assign \new_[27180]_  = \new_[27179]_  & \new_[27174]_ ;
  assign \new_[27183]_  = ~A168 & ~A169;
  assign \new_[27187]_  = A202 & A166;
  assign \new_[27188]_  = A167 & \new_[27187]_ ;
  assign \new_[27189]_  = \new_[27188]_  & \new_[27183]_ ;
  assign \new_[27193]_  = A236 & ~A233;
  assign \new_[27194]_  = A232 & \new_[27193]_ ;
  assign \new_[27198]_  = A269 & ~A266;
  assign \new_[27199]_  = A265 & \new_[27198]_ ;
  assign \new_[27200]_  = \new_[27199]_  & \new_[27194]_ ;
  assign \new_[27203]_  = ~A168 & ~A169;
  assign \new_[27207]_  = A199 & A166;
  assign \new_[27208]_  = A167 & \new_[27207]_ ;
  assign \new_[27209]_  = \new_[27208]_  & \new_[27203]_ ;
  assign \new_[27213]_  = A234 & A232;
  assign \new_[27214]_  = A201 & \new_[27213]_ ;
  assign \new_[27218]_  = A302 & ~A299;
  assign \new_[27219]_  = A298 & \new_[27218]_ ;
  assign \new_[27220]_  = \new_[27219]_  & \new_[27214]_ ;
  assign \new_[27223]_  = ~A168 & ~A169;
  assign \new_[27227]_  = A199 & A166;
  assign \new_[27228]_  = A167 & \new_[27227]_ ;
  assign \new_[27229]_  = \new_[27228]_  & \new_[27223]_ ;
  assign \new_[27233]_  = A234 & A232;
  assign \new_[27234]_  = A201 & \new_[27233]_ ;
  assign \new_[27238]_  = A302 & A299;
  assign \new_[27239]_  = ~A298 & \new_[27238]_ ;
  assign \new_[27240]_  = \new_[27239]_  & \new_[27234]_ ;
  assign \new_[27243]_  = ~A168 & ~A169;
  assign \new_[27247]_  = A199 & A166;
  assign \new_[27248]_  = A167 & \new_[27247]_ ;
  assign \new_[27249]_  = \new_[27248]_  & \new_[27243]_ ;
  assign \new_[27253]_  = A234 & A232;
  assign \new_[27254]_  = A201 & \new_[27253]_ ;
  assign \new_[27258]_  = A269 & A266;
  assign \new_[27259]_  = ~A265 & \new_[27258]_ ;
  assign \new_[27260]_  = \new_[27259]_  & \new_[27254]_ ;
  assign \new_[27263]_  = ~A168 & ~A169;
  assign \new_[27267]_  = A199 & A166;
  assign \new_[27268]_  = A167 & \new_[27267]_ ;
  assign \new_[27269]_  = \new_[27268]_  & \new_[27263]_ ;
  assign \new_[27273]_  = A234 & A232;
  assign \new_[27274]_  = A201 & \new_[27273]_ ;
  assign \new_[27278]_  = A269 & ~A266;
  assign \new_[27279]_  = A265 & \new_[27278]_ ;
  assign \new_[27280]_  = \new_[27279]_  & \new_[27274]_ ;
  assign \new_[27283]_  = ~A168 & ~A169;
  assign \new_[27287]_  = A199 & A166;
  assign \new_[27288]_  = A167 & \new_[27287]_ ;
  assign \new_[27289]_  = \new_[27288]_  & \new_[27283]_ ;
  assign \new_[27293]_  = A234 & A233;
  assign \new_[27294]_  = A201 & \new_[27293]_ ;
  assign \new_[27298]_  = A302 & ~A299;
  assign \new_[27299]_  = A298 & \new_[27298]_ ;
  assign \new_[27300]_  = \new_[27299]_  & \new_[27294]_ ;
  assign \new_[27303]_  = ~A168 & ~A169;
  assign \new_[27307]_  = A199 & A166;
  assign \new_[27308]_  = A167 & \new_[27307]_ ;
  assign \new_[27309]_  = \new_[27308]_  & \new_[27303]_ ;
  assign \new_[27313]_  = A234 & A233;
  assign \new_[27314]_  = A201 & \new_[27313]_ ;
  assign \new_[27318]_  = A302 & A299;
  assign \new_[27319]_  = ~A298 & \new_[27318]_ ;
  assign \new_[27320]_  = \new_[27319]_  & \new_[27314]_ ;
  assign \new_[27323]_  = ~A168 & ~A169;
  assign \new_[27327]_  = A199 & A166;
  assign \new_[27328]_  = A167 & \new_[27327]_ ;
  assign \new_[27329]_  = \new_[27328]_  & \new_[27323]_ ;
  assign \new_[27333]_  = A234 & A233;
  assign \new_[27334]_  = A201 & \new_[27333]_ ;
  assign \new_[27338]_  = A269 & A266;
  assign \new_[27339]_  = ~A265 & \new_[27338]_ ;
  assign \new_[27340]_  = \new_[27339]_  & \new_[27334]_ ;
  assign \new_[27343]_  = ~A168 & ~A169;
  assign \new_[27347]_  = A199 & A166;
  assign \new_[27348]_  = A167 & \new_[27347]_ ;
  assign \new_[27349]_  = \new_[27348]_  & \new_[27343]_ ;
  assign \new_[27353]_  = A234 & A233;
  assign \new_[27354]_  = A201 & \new_[27353]_ ;
  assign \new_[27358]_  = A269 & ~A266;
  assign \new_[27359]_  = A265 & \new_[27358]_ ;
  assign \new_[27360]_  = \new_[27359]_  & \new_[27354]_ ;
  assign \new_[27363]_  = ~A168 & ~A169;
  assign \new_[27367]_  = A199 & A166;
  assign \new_[27368]_  = A167 & \new_[27367]_ ;
  assign \new_[27369]_  = \new_[27368]_  & \new_[27363]_ ;
  assign \new_[27373]_  = A233 & ~A232;
  assign \new_[27374]_  = A201 & \new_[27373]_ ;
  assign \new_[27378]_  = A300 & A299;
  assign \new_[27379]_  = A236 & \new_[27378]_ ;
  assign \new_[27380]_  = \new_[27379]_  & \new_[27374]_ ;
  assign \new_[27383]_  = ~A168 & ~A169;
  assign \new_[27387]_  = A199 & A166;
  assign \new_[27388]_  = A167 & \new_[27387]_ ;
  assign \new_[27389]_  = \new_[27388]_  & \new_[27383]_ ;
  assign \new_[27393]_  = A233 & ~A232;
  assign \new_[27394]_  = A201 & \new_[27393]_ ;
  assign \new_[27398]_  = A300 & A298;
  assign \new_[27399]_  = A236 & \new_[27398]_ ;
  assign \new_[27400]_  = \new_[27399]_  & \new_[27394]_ ;
  assign \new_[27403]_  = ~A168 & ~A169;
  assign \new_[27407]_  = A199 & A166;
  assign \new_[27408]_  = A167 & \new_[27407]_ ;
  assign \new_[27409]_  = \new_[27408]_  & \new_[27403]_ ;
  assign \new_[27413]_  = A233 & ~A232;
  assign \new_[27414]_  = A201 & \new_[27413]_ ;
  assign \new_[27418]_  = A267 & A265;
  assign \new_[27419]_  = A236 & \new_[27418]_ ;
  assign \new_[27420]_  = \new_[27419]_  & \new_[27414]_ ;
  assign \new_[27423]_  = ~A168 & ~A169;
  assign \new_[27427]_  = A199 & A166;
  assign \new_[27428]_  = A167 & \new_[27427]_ ;
  assign \new_[27429]_  = \new_[27428]_  & \new_[27423]_ ;
  assign \new_[27433]_  = A233 & ~A232;
  assign \new_[27434]_  = A201 & \new_[27433]_ ;
  assign \new_[27438]_  = A267 & A266;
  assign \new_[27439]_  = A236 & \new_[27438]_ ;
  assign \new_[27440]_  = \new_[27439]_  & \new_[27434]_ ;
  assign \new_[27443]_  = ~A168 & ~A169;
  assign \new_[27447]_  = A199 & A166;
  assign \new_[27448]_  = A167 & \new_[27447]_ ;
  assign \new_[27449]_  = \new_[27448]_  & \new_[27443]_ ;
  assign \new_[27453]_  = ~A233 & A232;
  assign \new_[27454]_  = A201 & \new_[27453]_ ;
  assign \new_[27458]_  = A300 & A299;
  assign \new_[27459]_  = A236 & \new_[27458]_ ;
  assign \new_[27460]_  = \new_[27459]_  & \new_[27454]_ ;
  assign \new_[27463]_  = ~A168 & ~A169;
  assign \new_[27467]_  = A199 & A166;
  assign \new_[27468]_  = A167 & \new_[27467]_ ;
  assign \new_[27469]_  = \new_[27468]_  & \new_[27463]_ ;
  assign \new_[27473]_  = ~A233 & A232;
  assign \new_[27474]_  = A201 & \new_[27473]_ ;
  assign \new_[27478]_  = A300 & A298;
  assign \new_[27479]_  = A236 & \new_[27478]_ ;
  assign \new_[27480]_  = \new_[27479]_  & \new_[27474]_ ;
  assign \new_[27483]_  = ~A168 & ~A169;
  assign \new_[27487]_  = A199 & A166;
  assign \new_[27488]_  = A167 & \new_[27487]_ ;
  assign \new_[27489]_  = \new_[27488]_  & \new_[27483]_ ;
  assign \new_[27493]_  = ~A233 & A232;
  assign \new_[27494]_  = A201 & \new_[27493]_ ;
  assign \new_[27498]_  = A267 & A265;
  assign \new_[27499]_  = A236 & \new_[27498]_ ;
  assign \new_[27500]_  = \new_[27499]_  & \new_[27494]_ ;
  assign \new_[27503]_  = ~A168 & ~A169;
  assign \new_[27507]_  = A199 & A166;
  assign \new_[27508]_  = A167 & \new_[27507]_ ;
  assign \new_[27509]_  = \new_[27508]_  & \new_[27503]_ ;
  assign \new_[27513]_  = ~A233 & A232;
  assign \new_[27514]_  = A201 & \new_[27513]_ ;
  assign \new_[27518]_  = A267 & A266;
  assign \new_[27519]_  = A236 & \new_[27518]_ ;
  assign \new_[27520]_  = \new_[27519]_  & \new_[27514]_ ;
  assign \new_[27523]_  = ~A168 & ~A169;
  assign \new_[27527]_  = A200 & A166;
  assign \new_[27528]_  = A167 & \new_[27527]_ ;
  assign \new_[27529]_  = \new_[27528]_  & \new_[27523]_ ;
  assign \new_[27533]_  = A234 & A232;
  assign \new_[27534]_  = A201 & \new_[27533]_ ;
  assign \new_[27538]_  = A302 & ~A299;
  assign \new_[27539]_  = A298 & \new_[27538]_ ;
  assign \new_[27540]_  = \new_[27539]_  & \new_[27534]_ ;
  assign \new_[27543]_  = ~A168 & ~A169;
  assign \new_[27547]_  = A200 & A166;
  assign \new_[27548]_  = A167 & \new_[27547]_ ;
  assign \new_[27549]_  = \new_[27548]_  & \new_[27543]_ ;
  assign \new_[27553]_  = A234 & A232;
  assign \new_[27554]_  = A201 & \new_[27553]_ ;
  assign \new_[27558]_  = A302 & A299;
  assign \new_[27559]_  = ~A298 & \new_[27558]_ ;
  assign \new_[27560]_  = \new_[27559]_  & \new_[27554]_ ;
  assign \new_[27563]_  = ~A168 & ~A169;
  assign \new_[27567]_  = A200 & A166;
  assign \new_[27568]_  = A167 & \new_[27567]_ ;
  assign \new_[27569]_  = \new_[27568]_  & \new_[27563]_ ;
  assign \new_[27573]_  = A234 & A232;
  assign \new_[27574]_  = A201 & \new_[27573]_ ;
  assign \new_[27578]_  = A269 & A266;
  assign \new_[27579]_  = ~A265 & \new_[27578]_ ;
  assign \new_[27580]_  = \new_[27579]_  & \new_[27574]_ ;
  assign \new_[27583]_  = ~A168 & ~A169;
  assign \new_[27587]_  = A200 & A166;
  assign \new_[27588]_  = A167 & \new_[27587]_ ;
  assign \new_[27589]_  = \new_[27588]_  & \new_[27583]_ ;
  assign \new_[27593]_  = A234 & A232;
  assign \new_[27594]_  = A201 & \new_[27593]_ ;
  assign \new_[27598]_  = A269 & ~A266;
  assign \new_[27599]_  = A265 & \new_[27598]_ ;
  assign \new_[27600]_  = \new_[27599]_  & \new_[27594]_ ;
  assign \new_[27603]_  = ~A168 & ~A169;
  assign \new_[27607]_  = A200 & A166;
  assign \new_[27608]_  = A167 & \new_[27607]_ ;
  assign \new_[27609]_  = \new_[27608]_  & \new_[27603]_ ;
  assign \new_[27613]_  = A234 & A233;
  assign \new_[27614]_  = A201 & \new_[27613]_ ;
  assign \new_[27618]_  = A302 & ~A299;
  assign \new_[27619]_  = A298 & \new_[27618]_ ;
  assign \new_[27620]_  = \new_[27619]_  & \new_[27614]_ ;
  assign \new_[27623]_  = ~A168 & ~A169;
  assign \new_[27627]_  = A200 & A166;
  assign \new_[27628]_  = A167 & \new_[27627]_ ;
  assign \new_[27629]_  = \new_[27628]_  & \new_[27623]_ ;
  assign \new_[27633]_  = A234 & A233;
  assign \new_[27634]_  = A201 & \new_[27633]_ ;
  assign \new_[27638]_  = A302 & A299;
  assign \new_[27639]_  = ~A298 & \new_[27638]_ ;
  assign \new_[27640]_  = \new_[27639]_  & \new_[27634]_ ;
  assign \new_[27643]_  = ~A168 & ~A169;
  assign \new_[27647]_  = A200 & A166;
  assign \new_[27648]_  = A167 & \new_[27647]_ ;
  assign \new_[27649]_  = \new_[27648]_  & \new_[27643]_ ;
  assign \new_[27653]_  = A234 & A233;
  assign \new_[27654]_  = A201 & \new_[27653]_ ;
  assign \new_[27658]_  = A269 & A266;
  assign \new_[27659]_  = ~A265 & \new_[27658]_ ;
  assign \new_[27660]_  = \new_[27659]_  & \new_[27654]_ ;
  assign \new_[27663]_  = ~A168 & ~A169;
  assign \new_[27667]_  = A200 & A166;
  assign \new_[27668]_  = A167 & \new_[27667]_ ;
  assign \new_[27669]_  = \new_[27668]_  & \new_[27663]_ ;
  assign \new_[27673]_  = A234 & A233;
  assign \new_[27674]_  = A201 & \new_[27673]_ ;
  assign \new_[27678]_  = A269 & ~A266;
  assign \new_[27679]_  = A265 & \new_[27678]_ ;
  assign \new_[27680]_  = \new_[27679]_  & \new_[27674]_ ;
  assign \new_[27683]_  = ~A168 & ~A169;
  assign \new_[27687]_  = A200 & A166;
  assign \new_[27688]_  = A167 & \new_[27687]_ ;
  assign \new_[27689]_  = \new_[27688]_  & \new_[27683]_ ;
  assign \new_[27693]_  = A233 & ~A232;
  assign \new_[27694]_  = A201 & \new_[27693]_ ;
  assign \new_[27698]_  = A300 & A299;
  assign \new_[27699]_  = A236 & \new_[27698]_ ;
  assign \new_[27700]_  = \new_[27699]_  & \new_[27694]_ ;
  assign \new_[27703]_  = ~A168 & ~A169;
  assign \new_[27707]_  = A200 & A166;
  assign \new_[27708]_  = A167 & \new_[27707]_ ;
  assign \new_[27709]_  = \new_[27708]_  & \new_[27703]_ ;
  assign \new_[27713]_  = A233 & ~A232;
  assign \new_[27714]_  = A201 & \new_[27713]_ ;
  assign \new_[27718]_  = A300 & A298;
  assign \new_[27719]_  = A236 & \new_[27718]_ ;
  assign \new_[27720]_  = \new_[27719]_  & \new_[27714]_ ;
  assign \new_[27723]_  = ~A168 & ~A169;
  assign \new_[27727]_  = A200 & A166;
  assign \new_[27728]_  = A167 & \new_[27727]_ ;
  assign \new_[27729]_  = \new_[27728]_  & \new_[27723]_ ;
  assign \new_[27733]_  = A233 & ~A232;
  assign \new_[27734]_  = A201 & \new_[27733]_ ;
  assign \new_[27738]_  = A267 & A265;
  assign \new_[27739]_  = A236 & \new_[27738]_ ;
  assign \new_[27740]_  = \new_[27739]_  & \new_[27734]_ ;
  assign \new_[27743]_  = ~A168 & ~A169;
  assign \new_[27747]_  = A200 & A166;
  assign \new_[27748]_  = A167 & \new_[27747]_ ;
  assign \new_[27749]_  = \new_[27748]_  & \new_[27743]_ ;
  assign \new_[27753]_  = A233 & ~A232;
  assign \new_[27754]_  = A201 & \new_[27753]_ ;
  assign \new_[27758]_  = A267 & A266;
  assign \new_[27759]_  = A236 & \new_[27758]_ ;
  assign \new_[27760]_  = \new_[27759]_  & \new_[27754]_ ;
  assign \new_[27763]_  = ~A168 & ~A169;
  assign \new_[27767]_  = A200 & A166;
  assign \new_[27768]_  = A167 & \new_[27767]_ ;
  assign \new_[27769]_  = \new_[27768]_  & \new_[27763]_ ;
  assign \new_[27773]_  = ~A233 & A232;
  assign \new_[27774]_  = A201 & \new_[27773]_ ;
  assign \new_[27778]_  = A300 & A299;
  assign \new_[27779]_  = A236 & \new_[27778]_ ;
  assign \new_[27780]_  = \new_[27779]_  & \new_[27774]_ ;
  assign \new_[27783]_  = ~A168 & ~A169;
  assign \new_[27787]_  = A200 & A166;
  assign \new_[27788]_  = A167 & \new_[27787]_ ;
  assign \new_[27789]_  = \new_[27788]_  & \new_[27783]_ ;
  assign \new_[27793]_  = ~A233 & A232;
  assign \new_[27794]_  = A201 & \new_[27793]_ ;
  assign \new_[27798]_  = A300 & A298;
  assign \new_[27799]_  = A236 & \new_[27798]_ ;
  assign \new_[27800]_  = \new_[27799]_  & \new_[27794]_ ;
  assign \new_[27803]_  = ~A168 & ~A169;
  assign \new_[27807]_  = A200 & A166;
  assign \new_[27808]_  = A167 & \new_[27807]_ ;
  assign \new_[27809]_  = \new_[27808]_  & \new_[27803]_ ;
  assign \new_[27813]_  = ~A233 & A232;
  assign \new_[27814]_  = A201 & \new_[27813]_ ;
  assign \new_[27818]_  = A267 & A265;
  assign \new_[27819]_  = A236 & \new_[27818]_ ;
  assign \new_[27820]_  = \new_[27819]_  & \new_[27814]_ ;
  assign \new_[27823]_  = ~A168 & ~A169;
  assign \new_[27827]_  = A200 & A166;
  assign \new_[27828]_  = A167 & \new_[27827]_ ;
  assign \new_[27829]_  = \new_[27828]_  & \new_[27823]_ ;
  assign \new_[27833]_  = ~A233 & A232;
  assign \new_[27834]_  = A201 & \new_[27833]_ ;
  assign \new_[27838]_  = A267 & A266;
  assign \new_[27839]_  = A236 & \new_[27838]_ ;
  assign \new_[27840]_  = \new_[27839]_  & \new_[27834]_ ;
  assign \new_[27843]_  = ~A168 & ~A169;
  assign \new_[27847]_  = ~A199 & A166;
  assign \new_[27848]_  = A167 & \new_[27847]_ ;
  assign \new_[27849]_  = \new_[27848]_  & \new_[27843]_ ;
  assign \new_[27853]_  = A235 & A203;
  assign \new_[27854]_  = A200 & \new_[27853]_ ;
  assign \new_[27858]_  = A302 & ~A299;
  assign \new_[27859]_  = A298 & \new_[27858]_ ;
  assign \new_[27860]_  = \new_[27859]_  & \new_[27854]_ ;
  assign \new_[27863]_  = ~A168 & ~A169;
  assign \new_[27867]_  = ~A199 & A166;
  assign \new_[27868]_  = A167 & \new_[27867]_ ;
  assign \new_[27869]_  = \new_[27868]_  & \new_[27863]_ ;
  assign \new_[27873]_  = A235 & A203;
  assign \new_[27874]_  = A200 & \new_[27873]_ ;
  assign \new_[27878]_  = A302 & A299;
  assign \new_[27879]_  = ~A298 & \new_[27878]_ ;
  assign \new_[27880]_  = \new_[27879]_  & \new_[27874]_ ;
  assign \new_[27883]_  = ~A168 & ~A169;
  assign \new_[27887]_  = ~A199 & A166;
  assign \new_[27888]_  = A167 & \new_[27887]_ ;
  assign \new_[27889]_  = \new_[27888]_  & \new_[27883]_ ;
  assign \new_[27893]_  = A235 & A203;
  assign \new_[27894]_  = A200 & \new_[27893]_ ;
  assign \new_[27898]_  = A269 & A266;
  assign \new_[27899]_  = ~A265 & \new_[27898]_ ;
  assign \new_[27900]_  = \new_[27899]_  & \new_[27894]_ ;
  assign \new_[27903]_  = ~A168 & ~A169;
  assign \new_[27907]_  = ~A199 & A166;
  assign \new_[27908]_  = A167 & \new_[27907]_ ;
  assign \new_[27909]_  = \new_[27908]_  & \new_[27903]_ ;
  assign \new_[27913]_  = A235 & A203;
  assign \new_[27914]_  = A200 & \new_[27913]_ ;
  assign \new_[27918]_  = A269 & ~A266;
  assign \new_[27919]_  = A265 & \new_[27918]_ ;
  assign \new_[27920]_  = \new_[27919]_  & \new_[27914]_ ;
  assign \new_[27923]_  = ~A168 & ~A169;
  assign \new_[27927]_  = ~A199 & A166;
  assign \new_[27928]_  = A167 & \new_[27927]_ ;
  assign \new_[27929]_  = \new_[27928]_  & \new_[27923]_ ;
  assign \new_[27933]_  = A232 & A203;
  assign \new_[27934]_  = A200 & \new_[27933]_ ;
  assign \new_[27938]_  = A300 & A299;
  assign \new_[27939]_  = A234 & \new_[27938]_ ;
  assign \new_[27940]_  = \new_[27939]_  & \new_[27934]_ ;
  assign \new_[27943]_  = ~A168 & ~A169;
  assign \new_[27947]_  = ~A199 & A166;
  assign \new_[27948]_  = A167 & \new_[27947]_ ;
  assign \new_[27949]_  = \new_[27948]_  & \new_[27943]_ ;
  assign \new_[27953]_  = A232 & A203;
  assign \new_[27954]_  = A200 & \new_[27953]_ ;
  assign \new_[27958]_  = A300 & A298;
  assign \new_[27959]_  = A234 & \new_[27958]_ ;
  assign \new_[27960]_  = \new_[27959]_  & \new_[27954]_ ;
  assign \new_[27963]_  = ~A168 & ~A169;
  assign \new_[27967]_  = ~A199 & A166;
  assign \new_[27968]_  = A167 & \new_[27967]_ ;
  assign \new_[27969]_  = \new_[27968]_  & \new_[27963]_ ;
  assign \new_[27973]_  = A232 & A203;
  assign \new_[27974]_  = A200 & \new_[27973]_ ;
  assign \new_[27978]_  = A267 & A265;
  assign \new_[27979]_  = A234 & \new_[27978]_ ;
  assign \new_[27980]_  = \new_[27979]_  & \new_[27974]_ ;
  assign \new_[27983]_  = ~A168 & ~A169;
  assign \new_[27987]_  = ~A199 & A166;
  assign \new_[27988]_  = A167 & \new_[27987]_ ;
  assign \new_[27989]_  = \new_[27988]_  & \new_[27983]_ ;
  assign \new_[27993]_  = A232 & A203;
  assign \new_[27994]_  = A200 & \new_[27993]_ ;
  assign \new_[27998]_  = A267 & A266;
  assign \new_[27999]_  = A234 & \new_[27998]_ ;
  assign \new_[28000]_  = \new_[27999]_  & \new_[27994]_ ;
  assign \new_[28003]_  = ~A168 & ~A169;
  assign \new_[28007]_  = ~A199 & A166;
  assign \new_[28008]_  = A167 & \new_[28007]_ ;
  assign \new_[28009]_  = \new_[28008]_  & \new_[28003]_ ;
  assign \new_[28013]_  = A233 & A203;
  assign \new_[28014]_  = A200 & \new_[28013]_ ;
  assign \new_[28018]_  = A300 & A299;
  assign \new_[28019]_  = A234 & \new_[28018]_ ;
  assign \new_[28020]_  = \new_[28019]_  & \new_[28014]_ ;
  assign \new_[28023]_  = ~A168 & ~A169;
  assign \new_[28027]_  = ~A199 & A166;
  assign \new_[28028]_  = A167 & \new_[28027]_ ;
  assign \new_[28029]_  = \new_[28028]_  & \new_[28023]_ ;
  assign \new_[28033]_  = A233 & A203;
  assign \new_[28034]_  = A200 & \new_[28033]_ ;
  assign \new_[28038]_  = A300 & A298;
  assign \new_[28039]_  = A234 & \new_[28038]_ ;
  assign \new_[28040]_  = \new_[28039]_  & \new_[28034]_ ;
  assign \new_[28043]_  = ~A168 & ~A169;
  assign \new_[28047]_  = ~A199 & A166;
  assign \new_[28048]_  = A167 & \new_[28047]_ ;
  assign \new_[28049]_  = \new_[28048]_  & \new_[28043]_ ;
  assign \new_[28053]_  = A233 & A203;
  assign \new_[28054]_  = A200 & \new_[28053]_ ;
  assign \new_[28058]_  = A267 & A265;
  assign \new_[28059]_  = A234 & \new_[28058]_ ;
  assign \new_[28060]_  = \new_[28059]_  & \new_[28054]_ ;
  assign \new_[28063]_  = ~A168 & ~A169;
  assign \new_[28067]_  = ~A199 & A166;
  assign \new_[28068]_  = A167 & \new_[28067]_ ;
  assign \new_[28069]_  = \new_[28068]_  & \new_[28063]_ ;
  assign \new_[28073]_  = A233 & A203;
  assign \new_[28074]_  = A200 & \new_[28073]_ ;
  assign \new_[28078]_  = A267 & A266;
  assign \new_[28079]_  = A234 & \new_[28078]_ ;
  assign \new_[28080]_  = \new_[28079]_  & \new_[28074]_ ;
  assign \new_[28083]_  = ~A168 & ~A169;
  assign \new_[28087]_  = ~A199 & A166;
  assign \new_[28088]_  = A167 & \new_[28087]_ ;
  assign \new_[28089]_  = \new_[28088]_  & \new_[28083]_ ;
  assign \new_[28093]_  = ~A232 & A203;
  assign \new_[28094]_  = A200 & \new_[28093]_ ;
  assign \new_[28098]_  = A301 & A236;
  assign \new_[28099]_  = A233 & \new_[28098]_ ;
  assign \new_[28100]_  = \new_[28099]_  & \new_[28094]_ ;
  assign \new_[28103]_  = ~A168 & ~A169;
  assign \new_[28107]_  = ~A199 & A166;
  assign \new_[28108]_  = A167 & \new_[28107]_ ;
  assign \new_[28109]_  = \new_[28108]_  & \new_[28103]_ ;
  assign \new_[28113]_  = ~A232 & A203;
  assign \new_[28114]_  = A200 & \new_[28113]_ ;
  assign \new_[28118]_  = A268 & A236;
  assign \new_[28119]_  = A233 & \new_[28118]_ ;
  assign \new_[28120]_  = \new_[28119]_  & \new_[28114]_ ;
  assign \new_[28123]_  = ~A168 & ~A169;
  assign \new_[28127]_  = ~A199 & A166;
  assign \new_[28128]_  = A167 & \new_[28127]_ ;
  assign \new_[28129]_  = \new_[28128]_  & \new_[28123]_ ;
  assign \new_[28133]_  = A232 & A203;
  assign \new_[28134]_  = A200 & \new_[28133]_ ;
  assign \new_[28138]_  = A301 & A236;
  assign \new_[28139]_  = ~A233 & \new_[28138]_ ;
  assign \new_[28140]_  = \new_[28139]_  & \new_[28134]_ ;
  assign \new_[28143]_  = ~A168 & ~A169;
  assign \new_[28147]_  = ~A199 & A166;
  assign \new_[28148]_  = A167 & \new_[28147]_ ;
  assign \new_[28149]_  = \new_[28148]_  & \new_[28143]_ ;
  assign \new_[28153]_  = A232 & A203;
  assign \new_[28154]_  = A200 & \new_[28153]_ ;
  assign \new_[28158]_  = A268 & A236;
  assign \new_[28159]_  = ~A233 & \new_[28158]_ ;
  assign \new_[28160]_  = \new_[28159]_  & \new_[28154]_ ;
  assign \new_[28163]_  = ~A168 & ~A169;
  assign \new_[28167]_  = A199 & A166;
  assign \new_[28168]_  = A167 & \new_[28167]_ ;
  assign \new_[28169]_  = \new_[28168]_  & \new_[28163]_ ;
  assign \new_[28173]_  = A235 & A203;
  assign \new_[28174]_  = ~A200 & \new_[28173]_ ;
  assign \new_[28178]_  = A302 & ~A299;
  assign \new_[28179]_  = A298 & \new_[28178]_ ;
  assign \new_[28180]_  = \new_[28179]_  & \new_[28174]_ ;
  assign \new_[28183]_  = ~A168 & ~A169;
  assign \new_[28187]_  = A199 & A166;
  assign \new_[28188]_  = A167 & \new_[28187]_ ;
  assign \new_[28189]_  = \new_[28188]_  & \new_[28183]_ ;
  assign \new_[28193]_  = A235 & A203;
  assign \new_[28194]_  = ~A200 & \new_[28193]_ ;
  assign \new_[28198]_  = A302 & A299;
  assign \new_[28199]_  = ~A298 & \new_[28198]_ ;
  assign \new_[28200]_  = \new_[28199]_  & \new_[28194]_ ;
  assign \new_[28203]_  = ~A168 & ~A169;
  assign \new_[28207]_  = A199 & A166;
  assign \new_[28208]_  = A167 & \new_[28207]_ ;
  assign \new_[28209]_  = \new_[28208]_  & \new_[28203]_ ;
  assign \new_[28213]_  = A235 & A203;
  assign \new_[28214]_  = ~A200 & \new_[28213]_ ;
  assign \new_[28218]_  = A269 & A266;
  assign \new_[28219]_  = ~A265 & \new_[28218]_ ;
  assign \new_[28220]_  = \new_[28219]_  & \new_[28214]_ ;
  assign \new_[28223]_  = ~A168 & ~A169;
  assign \new_[28227]_  = A199 & A166;
  assign \new_[28228]_  = A167 & \new_[28227]_ ;
  assign \new_[28229]_  = \new_[28228]_  & \new_[28223]_ ;
  assign \new_[28233]_  = A235 & A203;
  assign \new_[28234]_  = ~A200 & \new_[28233]_ ;
  assign \new_[28238]_  = A269 & ~A266;
  assign \new_[28239]_  = A265 & \new_[28238]_ ;
  assign \new_[28240]_  = \new_[28239]_  & \new_[28234]_ ;
  assign \new_[28243]_  = ~A168 & ~A169;
  assign \new_[28247]_  = A199 & A166;
  assign \new_[28248]_  = A167 & \new_[28247]_ ;
  assign \new_[28249]_  = \new_[28248]_  & \new_[28243]_ ;
  assign \new_[28253]_  = A232 & A203;
  assign \new_[28254]_  = ~A200 & \new_[28253]_ ;
  assign \new_[28258]_  = A300 & A299;
  assign \new_[28259]_  = A234 & \new_[28258]_ ;
  assign \new_[28260]_  = \new_[28259]_  & \new_[28254]_ ;
  assign \new_[28263]_  = ~A168 & ~A169;
  assign \new_[28267]_  = A199 & A166;
  assign \new_[28268]_  = A167 & \new_[28267]_ ;
  assign \new_[28269]_  = \new_[28268]_  & \new_[28263]_ ;
  assign \new_[28273]_  = A232 & A203;
  assign \new_[28274]_  = ~A200 & \new_[28273]_ ;
  assign \new_[28278]_  = A300 & A298;
  assign \new_[28279]_  = A234 & \new_[28278]_ ;
  assign \new_[28280]_  = \new_[28279]_  & \new_[28274]_ ;
  assign \new_[28283]_  = ~A168 & ~A169;
  assign \new_[28287]_  = A199 & A166;
  assign \new_[28288]_  = A167 & \new_[28287]_ ;
  assign \new_[28289]_  = \new_[28288]_  & \new_[28283]_ ;
  assign \new_[28293]_  = A232 & A203;
  assign \new_[28294]_  = ~A200 & \new_[28293]_ ;
  assign \new_[28298]_  = A267 & A265;
  assign \new_[28299]_  = A234 & \new_[28298]_ ;
  assign \new_[28300]_  = \new_[28299]_  & \new_[28294]_ ;
  assign \new_[28303]_  = ~A168 & ~A169;
  assign \new_[28307]_  = A199 & A166;
  assign \new_[28308]_  = A167 & \new_[28307]_ ;
  assign \new_[28309]_  = \new_[28308]_  & \new_[28303]_ ;
  assign \new_[28313]_  = A232 & A203;
  assign \new_[28314]_  = ~A200 & \new_[28313]_ ;
  assign \new_[28318]_  = A267 & A266;
  assign \new_[28319]_  = A234 & \new_[28318]_ ;
  assign \new_[28320]_  = \new_[28319]_  & \new_[28314]_ ;
  assign \new_[28323]_  = ~A168 & ~A169;
  assign \new_[28327]_  = A199 & A166;
  assign \new_[28328]_  = A167 & \new_[28327]_ ;
  assign \new_[28329]_  = \new_[28328]_  & \new_[28323]_ ;
  assign \new_[28333]_  = A233 & A203;
  assign \new_[28334]_  = ~A200 & \new_[28333]_ ;
  assign \new_[28338]_  = A300 & A299;
  assign \new_[28339]_  = A234 & \new_[28338]_ ;
  assign \new_[28340]_  = \new_[28339]_  & \new_[28334]_ ;
  assign \new_[28343]_  = ~A168 & ~A169;
  assign \new_[28347]_  = A199 & A166;
  assign \new_[28348]_  = A167 & \new_[28347]_ ;
  assign \new_[28349]_  = \new_[28348]_  & \new_[28343]_ ;
  assign \new_[28353]_  = A233 & A203;
  assign \new_[28354]_  = ~A200 & \new_[28353]_ ;
  assign \new_[28358]_  = A300 & A298;
  assign \new_[28359]_  = A234 & \new_[28358]_ ;
  assign \new_[28360]_  = \new_[28359]_  & \new_[28354]_ ;
  assign \new_[28363]_  = ~A168 & ~A169;
  assign \new_[28367]_  = A199 & A166;
  assign \new_[28368]_  = A167 & \new_[28367]_ ;
  assign \new_[28369]_  = \new_[28368]_  & \new_[28363]_ ;
  assign \new_[28373]_  = A233 & A203;
  assign \new_[28374]_  = ~A200 & \new_[28373]_ ;
  assign \new_[28378]_  = A267 & A265;
  assign \new_[28379]_  = A234 & \new_[28378]_ ;
  assign \new_[28380]_  = \new_[28379]_  & \new_[28374]_ ;
  assign \new_[28383]_  = ~A168 & ~A169;
  assign \new_[28387]_  = A199 & A166;
  assign \new_[28388]_  = A167 & \new_[28387]_ ;
  assign \new_[28389]_  = \new_[28388]_  & \new_[28383]_ ;
  assign \new_[28393]_  = A233 & A203;
  assign \new_[28394]_  = ~A200 & \new_[28393]_ ;
  assign \new_[28398]_  = A267 & A266;
  assign \new_[28399]_  = A234 & \new_[28398]_ ;
  assign \new_[28400]_  = \new_[28399]_  & \new_[28394]_ ;
  assign \new_[28403]_  = ~A168 & ~A169;
  assign \new_[28407]_  = A199 & A166;
  assign \new_[28408]_  = A167 & \new_[28407]_ ;
  assign \new_[28409]_  = \new_[28408]_  & \new_[28403]_ ;
  assign \new_[28413]_  = ~A232 & A203;
  assign \new_[28414]_  = ~A200 & \new_[28413]_ ;
  assign \new_[28418]_  = A301 & A236;
  assign \new_[28419]_  = A233 & \new_[28418]_ ;
  assign \new_[28420]_  = \new_[28419]_  & \new_[28414]_ ;
  assign \new_[28423]_  = ~A168 & ~A169;
  assign \new_[28427]_  = A199 & A166;
  assign \new_[28428]_  = A167 & \new_[28427]_ ;
  assign \new_[28429]_  = \new_[28428]_  & \new_[28423]_ ;
  assign \new_[28433]_  = ~A232 & A203;
  assign \new_[28434]_  = ~A200 & \new_[28433]_ ;
  assign \new_[28438]_  = A268 & A236;
  assign \new_[28439]_  = A233 & \new_[28438]_ ;
  assign \new_[28440]_  = \new_[28439]_  & \new_[28434]_ ;
  assign \new_[28443]_  = ~A168 & ~A169;
  assign \new_[28447]_  = A199 & A166;
  assign \new_[28448]_  = A167 & \new_[28447]_ ;
  assign \new_[28449]_  = \new_[28448]_  & \new_[28443]_ ;
  assign \new_[28453]_  = A232 & A203;
  assign \new_[28454]_  = ~A200 & \new_[28453]_ ;
  assign \new_[28458]_  = A301 & A236;
  assign \new_[28459]_  = ~A233 & \new_[28458]_ ;
  assign \new_[28460]_  = \new_[28459]_  & \new_[28454]_ ;
  assign \new_[28463]_  = ~A168 & ~A169;
  assign \new_[28467]_  = A199 & A166;
  assign \new_[28468]_  = A167 & \new_[28467]_ ;
  assign \new_[28469]_  = \new_[28468]_  & \new_[28463]_ ;
  assign \new_[28473]_  = A232 & A203;
  assign \new_[28474]_  = ~A200 & \new_[28473]_ ;
  assign \new_[28478]_  = A268 & A236;
  assign \new_[28479]_  = ~A233 & \new_[28478]_ ;
  assign \new_[28480]_  = \new_[28479]_  & \new_[28474]_ ;
  assign \new_[28483]_  = ~A169 & ~A170;
  assign \new_[28487]_  = A201 & A199;
  assign \new_[28488]_  = ~A168 & \new_[28487]_ ;
  assign \new_[28489]_  = \new_[28488]_  & \new_[28483]_ ;
  assign \new_[28493]_  = A236 & A233;
  assign \new_[28494]_  = ~A232 & \new_[28493]_ ;
  assign \new_[28498]_  = A302 & ~A299;
  assign \new_[28499]_  = A298 & \new_[28498]_ ;
  assign \new_[28500]_  = \new_[28499]_  & \new_[28494]_ ;
  assign \new_[28503]_  = ~A169 & ~A170;
  assign \new_[28507]_  = A201 & A199;
  assign \new_[28508]_  = ~A168 & \new_[28507]_ ;
  assign \new_[28509]_  = \new_[28508]_  & \new_[28503]_ ;
  assign \new_[28513]_  = A236 & A233;
  assign \new_[28514]_  = ~A232 & \new_[28513]_ ;
  assign \new_[28518]_  = A302 & A299;
  assign \new_[28519]_  = ~A298 & \new_[28518]_ ;
  assign \new_[28520]_  = \new_[28519]_  & \new_[28514]_ ;
  assign \new_[28523]_  = ~A169 & ~A170;
  assign \new_[28527]_  = A201 & A199;
  assign \new_[28528]_  = ~A168 & \new_[28527]_ ;
  assign \new_[28529]_  = \new_[28528]_  & \new_[28523]_ ;
  assign \new_[28533]_  = A236 & A233;
  assign \new_[28534]_  = ~A232 & \new_[28533]_ ;
  assign \new_[28538]_  = A269 & A266;
  assign \new_[28539]_  = ~A265 & \new_[28538]_ ;
  assign \new_[28540]_  = \new_[28539]_  & \new_[28534]_ ;
  assign \new_[28543]_  = ~A169 & ~A170;
  assign \new_[28547]_  = A201 & A199;
  assign \new_[28548]_  = ~A168 & \new_[28547]_ ;
  assign \new_[28549]_  = \new_[28548]_  & \new_[28543]_ ;
  assign \new_[28553]_  = A236 & A233;
  assign \new_[28554]_  = ~A232 & \new_[28553]_ ;
  assign \new_[28558]_  = A269 & ~A266;
  assign \new_[28559]_  = A265 & \new_[28558]_ ;
  assign \new_[28560]_  = \new_[28559]_  & \new_[28554]_ ;
  assign \new_[28563]_  = ~A169 & ~A170;
  assign \new_[28567]_  = A201 & A199;
  assign \new_[28568]_  = ~A168 & \new_[28567]_ ;
  assign \new_[28569]_  = \new_[28568]_  & \new_[28563]_ ;
  assign \new_[28573]_  = A236 & ~A233;
  assign \new_[28574]_  = A232 & \new_[28573]_ ;
  assign \new_[28578]_  = A302 & ~A299;
  assign \new_[28579]_  = A298 & \new_[28578]_ ;
  assign \new_[28580]_  = \new_[28579]_  & \new_[28574]_ ;
  assign \new_[28583]_  = ~A169 & ~A170;
  assign \new_[28587]_  = A201 & A199;
  assign \new_[28588]_  = ~A168 & \new_[28587]_ ;
  assign \new_[28589]_  = \new_[28588]_  & \new_[28583]_ ;
  assign \new_[28593]_  = A236 & ~A233;
  assign \new_[28594]_  = A232 & \new_[28593]_ ;
  assign \new_[28598]_  = A302 & A299;
  assign \new_[28599]_  = ~A298 & \new_[28598]_ ;
  assign \new_[28600]_  = \new_[28599]_  & \new_[28594]_ ;
  assign \new_[28603]_  = ~A169 & ~A170;
  assign \new_[28607]_  = A201 & A199;
  assign \new_[28608]_  = ~A168 & \new_[28607]_ ;
  assign \new_[28609]_  = \new_[28608]_  & \new_[28603]_ ;
  assign \new_[28613]_  = A236 & ~A233;
  assign \new_[28614]_  = A232 & \new_[28613]_ ;
  assign \new_[28618]_  = A269 & A266;
  assign \new_[28619]_  = ~A265 & \new_[28618]_ ;
  assign \new_[28620]_  = \new_[28619]_  & \new_[28614]_ ;
  assign \new_[28623]_  = ~A169 & ~A170;
  assign \new_[28627]_  = A201 & A199;
  assign \new_[28628]_  = ~A168 & \new_[28627]_ ;
  assign \new_[28629]_  = \new_[28628]_  & \new_[28623]_ ;
  assign \new_[28633]_  = A236 & ~A233;
  assign \new_[28634]_  = A232 & \new_[28633]_ ;
  assign \new_[28638]_  = A269 & ~A266;
  assign \new_[28639]_  = A265 & \new_[28638]_ ;
  assign \new_[28640]_  = \new_[28639]_  & \new_[28634]_ ;
  assign \new_[28643]_  = ~A169 & ~A170;
  assign \new_[28647]_  = A201 & A200;
  assign \new_[28648]_  = ~A168 & \new_[28647]_ ;
  assign \new_[28649]_  = \new_[28648]_  & \new_[28643]_ ;
  assign \new_[28653]_  = A236 & A233;
  assign \new_[28654]_  = ~A232 & \new_[28653]_ ;
  assign \new_[28658]_  = A302 & ~A299;
  assign \new_[28659]_  = A298 & \new_[28658]_ ;
  assign \new_[28660]_  = \new_[28659]_  & \new_[28654]_ ;
  assign \new_[28663]_  = ~A169 & ~A170;
  assign \new_[28667]_  = A201 & A200;
  assign \new_[28668]_  = ~A168 & \new_[28667]_ ;
  assign \new_[28669]_  = \new_[28668]_  & \new_[28663]_ ;
  assign \new_[28673]_  = A236 & A233;
  assign \new_[28674]_  = ~A232 & \new_[28673]_ ;
  assign \new_[28678]_  = A302 & A299;
  assign \new_[28679]_  = ~A298 & \new_[28678]_ ;
  assign \new_[28680]_  = \new_[28679]_  & \new_[28674]_ ;
  assign \new_[28683]_  = ~A169 & ~A170;
  assign \new_[28687]_  = A201 & A200;
  assign \new_[28688]_  = ~A168 & \new_[28687]_ ;
  assign \new_[28689]_  = \new_[28688]_  & \new_[28683]_ ;
  assign \new_[28693]_  = A236 & A233;
  assign \new_[28694]_  = ~A232 & \new_[28693]_ ;
  assign \new_[28698]_  = A269 & A266;
  assign \new_[28699]_  = ~A265 & \new_[28698]_ ;
  assign \new_[28700]_  = \new_[28699]_  & \new_[28694]_ ;
  assign \new_[28703]_  = ~A169 & ~A170;
  assign \new_[28707]_  = A201 & A200;
  assign \new_[28708]_  = ~A168 & \new_[28707]_ ;
  assign \new_[28709]_  = \new_[28708]_  & \new_[28703]_ ;
  assign \new_[28713]_  = A236 & A233;
  assign \new_[28714]_  = ~A232 & \new_[28713]_ ;
  assign \new_[28718]_  = A269 & ~A266;
  assign \new_[28719]_  = A265 & \new_[28718]_ ;
  assign \new_[28720]_  = \new_[28719]_  & \new_[28714]_ ;
  assign \new_[28723]_  = ~A169 & ~A170;
  assign \new_[28727]_  = A201 & A200;
  assign \new_[28728]_  = ~A168 & \new_[28727]_ ;
  assign \new_[28729]_  = \new_[28728]_  & \new_[28723]_ ;
  assign \new_[28733]_  = A236 & ~A233;
  assign \new_[28734]_  = A232 & \new_[28733]_ ;
  assign \new_[28738]_  = A302 & ~A299;
  assign \new_[28739]_  = A298 & \new_[28738]_ ;
  assign \new_[28740]_  = \new_[28739]_  & \new_[28734]_ ;
  assign \new_[28743]_  = ~A169 & ~A170;
  assign \new_[28747]_  = A201 & A200;
  assign \new_[28748]_  = ~A168 & \new_[28747]_ ;
  assign \new_[28749]_  = \new_[28748]_  & \new_[28743]_ ;
  assign \new_[28753]_  = A236 & ~A233;
  assign \new_[28754]_  = A232 & \new_[28753]_ ;
  assign \new_[28758]_  = A302 & A299;
  assign \new_[28759]_  = ~A298 & \new_[28758]_ ;
  assign \new_[28760]_  = \new_[28759]_  & \new_[28754]_ ;
  assign \new_[28763]_  = ~A169 & ~A170;
  assign \new_[28767]_  = A201 & A200;
  assign \new_[28768]_  = ~A168 & \new_[28767]_ ;
  assign \new_[28769]_  = \new_[28768]_  & \new_[28763]_ ;
  assign \new_[28773]_  = A236 & ~A233;
  assign \new_[28774]_  = A232 & \new_[28773]_ ;
  assign \new_[28778]_  = A269 & A266;
  assign \new_[28779]_  = ~A265 & \new_[28778]_ ;
  assign \new_[28780]_  = \new_[28779]_  & \new_[28774]_ ;
  assign \new_[28783]_  = ~A169 & ~A170;
  assign \new_[28787]_  = A201 & A200;
  assign \new_[28788]_  = ~A168 & \new_[28787]_ ;
  assign \new_[28789]_  = \new_[28788]_  & \new_[28783]_ ;
  assign \new_[28793]_  = A236 & ~A233;
  assign \new_[28794]_  = A232 & \new_[28793]_ ;
  assign \new_[28798]_  = A269 & ~A266;
  assign \new_[28799]_  = A265 & \new_[28798]_ ;
  assign \new_[28800]_  = \new_[28799]_  & \new_[28794]_ ;
  assign \new_[28803]_  = ~A169 & ~A170;
  assign \new_[28807]_  = A200 & ~A199;
  assign \new_[28808]_  = ~A168 & \new_[28807]_ ;
  assign \new_[28809]_  = \new_[28808]_  & \new_[28803]_ ;
  assign \new_[28813]_  = A234 & A232;
  assign \new_[28814]_  = A203 & \new_[28813]_ ;
  assign \new_[28818]_  = A302 & ~A299;
  assign \new_[28819]_  = A298 & \new_[28818]_ ;
  assign \new_[28820]_  = \new_[28819]_  & \new_[28814]_ ;
  assign \new_[28823]_  = ~A169 & ~A170;
  assign \new_[28827]_  = A200 & ~A199;
  assign \new_[28828]_  = ~A168 & \new_[28827]_ ;
  assign \new_[28829]_  = \new_[28828]_  & \new_[28823]_ ;
  assign \new_[28833]_  = A234 & A232;
  assign \new_[28834]_  = A203 & \new_[28833]_ ;
  assign \new_[28838]_  = A302 & A299;
  assign \new_[28839]_  = ~A298 & \new_[28838]_ ;
  assign \new_[28840]_  = \new_[28839]_  & \new_[28834]_ ;
  assign \new_[28843]_  = ~A169 & ~A170;
  assign \new_[28847]_  = A200 & ~A199;
  assign \new_[28848]_  = ~A168 & \new_[28847]_ ;
  assign \new_[28849]_  = \new_[28848]_  & \new_[28843]_ ;
  assign \new_[28853]_  = A234 & A232;
  assign \new_[28854]_  = A203 & \new_[28853]_ ;
  assign \new_[28858]_  = A269 & A266;
  assign \new_[28859]_  = ~A265 & \new_[28858]_ ;
  assign \new_[28860]_  = \new_[28859]_  & \new_[28854]_ ;
  assign \new_[28863]_  = ~A169 & ~A170;
  assign \new_[28867]_  = A200 & ~A199;
  assign \new_[28868]_  = ~A168 & \new_[28867]_ ;
  assign \new_[28869]_  = \new_[28868]_  & \new_[28863]_ ;
  assign \new_[28873]_  = A234 & A232;
  assign \new_[28874]_  = A203 & \new_[28873]_ ;
  assign \new_[28878]_  = A269 & ~A266;
  assign \new_[28879]_  = A265 & \new_[28878]_ ;
  assign \new_[28880]_  = \new_[28879]_  & \new_[28874]_ ;
  assign \new_[28883]_  = ~A169 & ~A170;
  assign \new_[28887]_  = A200 & ~A199;
  assign \new_[28888]_  = ~A168 & \new_[28887]_ ;
  assign \new_[28889]_  = \new_[28888]_  & \new_[28883]_ ;
  assign \new_[28893]_  = A234 & A233;
  assign \new_[28894]_  = A203 & \new_[28893]_ ;
  assign \new_[28898]_  = A302 & ~A299;
  assign \new_[28899]_  = A298 & \new_[28898]_ ;
  assign \new_[28900]_  = \new_[28899]_  & \new_[28894]_ ;
  assign \new_[28903]_  = ~A169 & ~A170;
  assign \new_[28907]_  = A200 & ~A199;
  assign \new_[28908]_  = ~A168 & \new_[28907]_ ;
  assign \new_[28909]_  = \new_[28908]_  & \new_[28903]_ ;
  assign \new_[28913]_  = A234 & A233;
  assign \new_[28914]_  = A203 & \new_[28913]_ ;
  assign \new_[28918]_  = A302 & A299;
  assign \new_[28919]_  = ~A298 & \new_[28918]_ ;
  assign \new_[28920]_  = \new_[28919]_  & \new_[28914]_ ;
  assign \new_[28923]_  = ~A169 & ~A170;
  assign \new_[28927]_  = A200 & ~A199;
  assign \new_[28928]_  = ~A168 & \new_[28927]_ ;
  assign \new_[28929]_  = \new_[28928]_  & \new_[28923]_ ;
  assign \new_[28933]_  = A234 & A233;
  assign \new_[28934]_  = A203 & \new_[28933]_ ;
  assign \new_[28938]_  = A269 & A266;
  assign \new_[28939]_  = ~A265 & \new_[28938]_ ;
  assign \new_[28940]_  = \new_[28939]_  & \new_[28934]_ ;
  assign \new_[28943]_  = ~A169 & ~A170;
  assign \new_[28947]_  = A200 & ~A199;
  assign \new_[28948]_  = ~A168 & \new_[28947]_ ;
  assign \new_[28949]_  = \new_[28948]_  & \new_[28943]_ ;
  assign \new_[28953]_  = A234 & A233;
  assign \new_[28954]_  = A203 & \new_[28953]_ ;
  assign \new_[28958]_  = A269 & ~A266;
  assign \new_[28959]_  = A265 & \new_[28958]_ ;
  assign \new_[28960]_  = \new_[28959]_  & \new_[28954]_ ;
  assign \new_[28963]_  = ~A169 & ~A170;
  assign \new_[28967]_  = A200 & ~A199;
  assign \new_[28968]_  = ~A168 & \new_[28967]_ ;
  assign \new_[28969]_  = \new_[28968]_  & \new_[28963]_ ;
  assign \new_[28973]_  = A233 & ~A232;
  assign \new_[28974]_  = A203 & \new_[28973]_ ;
  assign \new_[28978]_  = A300 & A299;
  assign \new_[28979]_  = A236 & \new_[28978]_ ;
  assign \new_[28980]_  = \new_[28979]_  & \new_[28974]_ ;
  assign \new_[28983]_  = ~A169 & ~A170;
  assign \new_[28987]_  = A200 & ~A199;
  assign \new_[28988]_  = ~A168 & \new_[28987]_ ;
  assign \new_[28989]_  = \new_[28988]_  & \new_[28983]_ ;
  assign \new_[28993]_  = A233 & ~A232;
  assign \new_[28994]_  = A203 & \new_[28993]_ ;
  assign \new_[28998]_  = A300 & A298;
  assign \new_[28999]_  = A236 & \new_[28998]_ ;
  assign \new_[29000]_  = \new_[28999]_  & \new_[28994]_ ;
  assign \new_[29003]_  = ~A169 & ~A170;
  assign \new_[29007]_  = A200 & ~A199;
  assign \new_[29008]_  = ~A168 & \new_[29007]_ ;
  assign \new_[29009]_  = \new_[29008]_  & \new_[29003]_ ;
  assign \new_[29013]_  = A233 & ~A232;
  assign \new_[29014]_  = A203 & \new_[29013]_ ;
  assign \new_[29018]_  = A267 & A265;
  assign \new_[29019]_  = A236 & \new_[29018]_ ;
  assign \new_[29020]_  = \new_[29019]_  & \new_[29014]_ ;
  assign \new_[29023]_  = ~A169 & ~A170;
  assign \new_[29027]_  = A200 & ~A199;
  assign \new_[29028]_  = ~A168 & \new_[29027]_ ;
  assign \new_[29029]_  = \new_[29028]_  & \new_[29023]_ ;
  assign \new_[29033]_  = A233 & ~A232;
  assign \new_[29034]_  = A203 & \new_[29033]_ ;
  assign \new_[29038]_  = A267 & A266;
  assign \new_[29039]_  = A236 & \new_[29038]_ ;
  assign \new_[29040]_  = \new_[29039]_  & \new_[29034]_ ;
  assign \new_[29043]_  = ~A169 & ~A170;
  assign \new_[29047]_  = A200 & ~A199;
  assign \new_[29048]_  = ~A168 & \new_[29047]_ ;
  assign \new_[29049]_  = \new_[29048]_  & \new_[29043]_ ;
  assign \new_[29053]_  = ~A233 & A232;
  assign \new_[29054]_  = A203 & \new_[29053]_ ;
  assign \new_[29058]_  = A300 & A299;
  assign \new_[29059]_  = A236 & \new_[29058]_ ;
  assign \new_[29060]_  = \new_[29059]_  & \new_[29054]_ ;
  assign \new_[29063]_  = ~A169 & ~A170;
  assign \new_[29067]_  = A200 & ~A199;
  assign \new_[29068]_  = ~A168 & \new_[29067]_ ;
  assign \new_[29069]_  = \new_[29068]_  & \new_[29063]_ ;
  assign \new_[29073]_  = ~A233 & A232;
  assign \new_[29074]_  = A203 & \new_[29073]_ ;
  assign \new_[29078]_  = A300 & A298;
  assign \new_[29079]_  = A236 & \new_[29078]_ ;
  assign \new_[29080]_  = \new_[29079]_  & \new_[29074]_ ;
  assign \new_[29083]_  = ~A169 & ~A170;
  assign \new_[29087]_  = A200 & ~A199;
  assign \new_[29088]_  = ~A168 & \new_[29087]_ ;
  assign \new_[29089]_  = \new_[29088]_  & \new_[29083]_ ;
  assign \new_[29093]_  = ~A233 & A232;
  assign \new_[29094]_  = A203 & \new_[29093]_ ;
  assign \new_[29098]_  = A267 & A265;
  assign \new_[29099]_  = A236 & \new_[29098]_ ;
  assign \new_[29100]_  = \new_[29099]_  & \new_[29094]_ ;
  assign \new_[29103]_  = ~A169 & ~A170;
  assign \new_[29107]_  = A200 & ~A199;
  assign \new_[29108]_  = ~A168 & \new_[29107]_ ;
  assign \new_[29109]_  = \new_[29108]_  & \new_[29103]_ ;
  assign \new_[29113]_  = ~A233 & A232;
  assign \new_[29114]_  = A203 & \new_[29113]_ ;
  assign \new_[29118]_  = A267 & A266;
  assign \new_[29119]_  = A236 & \new_[29118]_ ;
  assign \new_[29120]_  = \new_[29119]_  & \new_[29114]_ ;
  assign \new_[29123]_  = ~A169 & ~A170;
  assign \new_[29127]_  = ~A200 & A199;
  assign \new_[29128]_  = ~A168 & \new_[29127]_ ;
  assign \new_[29129]_  = \new_[29128]_  & \new_[29123]_ ;
  assign \new_[29133]_  = A234 & A232;
  assign \new_[29134]_  = A203 & \new_[29133]_ ;
  assign \new_[29138]_  = A302 & ~A299;
  assign \new_[29139]_  = A298 & \new_[29138]_ ;
  assign \new_[29140]_  = \new_[29139]_  & \new_[29134]_ ;
  assign \new_[29143]_  = ~A169 & ~A170;
  assign \new_[29147]_  = ~A200 & A199;
  assign \new_[29148]_  = ~A168 & \new_[29147]_ ;
  assign \new_[29149]_  = \new_[29148]_  & \new_[29143]_ ;
  assign \new_[29153]_  = A234 & A232;
  assign \new_[29154]_  = A203 & \new_[29153]_ ;
  assign \new_[29158]_  = A302 & A299;
  assign \new_[29159]_  = ~A298 & \new_[29158]_ ;
  assign \new_[29160]_  = \new_[29159]_  & \new_[29154]_ ;
  assign \new_[29163]_  = ~A169 & ~A170;
  assign \new_[29167]_  = ~A200 & A199;
  assign \new_[29168]_  = ~A168 & \new_[29167]_ ;
  assign \new_[29169]_  = \new_[29168]_  & \new_[29163]_ ;
  assign \new_[29173]_  = A234 & A232;
  assign \new_[29174]_  = A203 & \new_[29173]_ ;
  assign \new_[29178]_  = A269 & A266;
  assign \new_[29179]_  = ~A265 & \new_[29178]_ ;
  assign \new_[29180]_  = \new_[29179]_  & \new_[29174]_ ;
  assign \new_[29183]_  = ~A169 & ~A170;
  assign \new_[29187]_  = ~A200 & A199;
  assign \new_[29188]_  = ~A168 & \new_[29187]_ ;
  assign \new_[29189]_  = \new_[29188]_  & \new_[29183]_ ;
  assign \new_[29193]_  = A234 & A232;
  assign \new_[29194]_  = A203 & \new_[29193]_ ;
  assign \new_[29198]_  = A269 & ~A266;
  assign \new_[29199]_  = A265 & \new_[29198]_ ;
  assign \new_[29200]_  = \new_[29199]_  & \new_[29194]_ ;
  assign \new_[29203]_  = ~A169 & ~A170;
  assign \new_[29207]_  = ~A200 & A199;
  assign \new_[29208]_  = ~A168 & \new_[29207]_ ;
  assign \new_[29209]_  = \new_[29208]_  & \new_[29203]_ ;
  assign \new_[29213]_  = A234 & A233;
  assign \new_[29214]_  = A203 & \new_[29213]_ ;
  assign \new_[29218]_  = A302 & ~A299;
  assign \new_[29219]_  = A298 & \new_[29218]_ ;
  assign \new_[29220]_  = \new_[29219]_  & \new_[29214]_ ;
  assign \new_[29223]_  = ~A169 & ~A170;
  assign \new_[29227]_  = ~A200 & A199;
  assign \new_[29228]_  = ~A168 & \new_[29227]_ ;
  assign \new_[29229]_  = \new_[29228]_  & \new_[29223]_ ;
  assign \new_[29233]_  = A234 & A233;
  assign \new_[29234]_  = A203 & \new_[29233]_ ;
  assign \new_[29238]_  = A302 & A299;
  assign \new_[29239]_  = ~A298 & \new_[29238]_ ;
  assign \new_[29240]_  = \new_[29239]_  & \new_[29234]_ ;
  assign \new_[29243]_  = ~A169 & ~A170;
  assign \new_[29247]_  = ~A200 & A199;
  assign \new_[29248]_  = ~A168 & \new_[29247]_ ;
  assign \new_[29249]_  = \new_[29248]_  & \new_[29243]_ ;
  assign \new_[29253]_  = A234 & A233;
  assign \new_[29254]_  = A203 & \new_[29253]_ ;
  assign \new_[29258]_  = A269 & A266;
  assign \new_[29259]_  = ~A265 & \new_[29258]_ ;
  assign \new_[29260]_  = \new_[29259]_  & \new_[29254]_ ;
  assign \new_[29263]_  = ~A169 & ~A170;
  assign \new_[29267]_  = ~A200 & A199;
  assign \new_[29268]_  = ~A168 & \new_[29267]_ ;
  assign \new_[29269]_  = \new_[29268]_  & \new_[29263]_ ;
  assign \new_[29273]_  = A234 & A233;
  assign \new_[29274]_  = A203 & \new_[29273]_ ;
  assign \new_[29278]_  = A269 & ~A266;
  assign \new_[29279]_  = A265 & \new_[29278]_ ;
  assign \new_[29280]_  = \new_[29279]_  & \new_[29274]_ ;
  assign \new_[29283]_  = ~A169 & ~A170;
  assign \new_[29287]_  = ~A200 & A199;
  assign \new_[29288]_  = ~A168 & \new_[29287]_ ;
  assign \new_[29289]_  = \new_[29288]_  & \new_[29283]_ ;
  assign \new_[29293]_  = A233 & ~A232;
  assign \new_[29294]_  = A203 & \new_[29293]_ ;
  assign \new_[29298]_  = A300 & A299;
  assign \new_[29299]_  = A236 & \new_[29298]_ ;
  assign \new_[29300]_  = \new_[29299]_  & \new_[29294]_ ;
  assign \new_[29303]_  = ~A169 & ~A170;
  assign \new_[29307]_  = ~A200 & A199;
  assign \new_[29308]_  = ~A168 & \new_[29307]_ ;
  assign \new_[29309]_  = \new_[29308]_  & \new_[29303]_ ;
  assign \new_[29313]_  = A233 & ~A232;
  assign \new_[29314]_  = A203 & \new_[29313]_ ;
  assign \new_[29318]_  = A300 & A298;
  assign \new_[29319]_  = A236 & \new_[29318]_ ;
  assign \new_[29320]_  = \new_[29319]_  & \new_[29314]_ ;
  assign \new_[29323]_  = ~A169 & ~A170;
  assign \new_[29327]_  = ~A200 & A199;
  assign \new_[29328]_  = ~A168 & \new_[29327]_ ;
  assign \new_[29329]_  = \new_[29328]_  & \new_[29323]_ ;
  assign \new_[29333]_  = A233 & ~A232;
  assign \new_[29334]_  = A203 & \new_[29333]_ ;
  assign \new_[29338]_  = A267 & A265;
  assign \new_[29339]_  = A236 & \new_[29338]_ ;
  assign \new_[29340]_  = \new_[29339]_  & \new_[29334]_ ;
  assign \new_[29343]_  = ~A169 & ~A170;
  assign \new_[29347]_  = ~A200 & A199;
  assign \new_[29348]_  = ~A168 & \new_[29347]_ ;
  assign \new_[29349]_  = \new_[29348]_  & \new_[29343]_ ;
  assign \new_[29353]_  = A233 & ~A232;
  assign \new_[29354]_  = A203 & \new_[29353]_ ;
  assign \new_[29358]_  = A267 & A266;
  assign \new_[29359]_  = A236 & \new_[29358]_ ;
  assign \new_[29360]_  = \new_[29359]_  & \new_[29354]_ ;
  assign \new_[29363]_  = ~A169 & ~A170;
  assign \new_[29367]_  = ~A200 & A199;
  assign \new_[29368]_  = ~A168 & \new_[29367]_ ;
  assign \new_[29369]_  = \new_[29368]_  & \new_[29363]_ ;
  assign \new_[29373]_  = ~A233 & A232;
  assign \new_[29374]_  = A203 & \new_[29373]_ ;
  assign \new_[29378]_  = A300 & A299;
  assign \new_[29379]_  = A236 & \new_[29378]_ ;
  assign \new_[29380]_  = \new_[29379]_  & \new_[29374]_ ;
  assign \new_[29383]_  = ~A169 & ~A170;
  assign \new_[29387]_  = ~A200 & A199;
  assign \new_[29388]_  = ~A168 & \new_[29387]_ ;
  assign \new_[29389]_  = \new_[29388]_  & \new_[29383]_ ;
  assign \new_[29393]_  = ~A233 & A232;
  assign \new_[29394]_  = A203 & \new_[29393]_ ;
  assign \new_[29398]_  = A300 & A298;
  assign \new_[29399]_  = A236 & \new_[29398]_ ;
  assign \new_[29400]_  = \new_[29399]_  & \new_[29394]_ ;
  assign \new_[29403]_  = ~A169 & ~A170;
  assign \new_[29407]_  = ~A200 & A199;
  assign \new_[29408]_  = ~A168 & \new_[29407]_ ;
  assign \new_[29409]_  = \new_[29408]_  & \new_[29403]_ ;
  assign \new_[29413]_  = ~A233 & A232;
  assign \new_[29414]_  = A203 & \new_[29413]_ ;
  assign \new_[29418]_  = A267 & A265;
  assign \new_[29419]_  = A236 & \new_[29418]_ ;
  assign \new_[29420]_  = \new_[29419]_  & \new_[29414]_ ;
  assign \new_[29423]_  = ~A169 & ~A170;
  assign \new_[29427]_  = ~A200 & A199;
  assign \new_[29428]_  = ~A168 & \new_[29427]_ ;
  assign \new_[29429]_  = \new_[29428]_  & \new_[29423]_ ;
  assign \new_[29433]_  = ~A233 & A232;
  assign \new_[29434]_  = A203 & \new_[29433]_ ;
  assign \new_[29438]_  = A267 & A266;
  assign \new_[29439]_  = A236 & \new_[29438]_ ;
  assign \new_[29440]_  = \new_[29439]_  & \new_[29434]_ ;
  assign \new_[29444]_  = A199 & A166;
  assign \new_[29445]_  = A168 & \new_[29444]_ ;
  assign \new_[29449]_  = ~A202 & ~A201;
  assign \new_[29450]_  = A200 & \new_[29449]_ ;
  assign \new_[29451]_  = \new_[29450]_  & \new_[29445]_ ;
  assign \new_[29455]_  = A236 & A233;
  assign \new_[29456]_  = ~A232 & \new_[29455]_ ;
  assign \new_[29460]_  = A302 & ~A299;
  assign \new_[29461]_  = A298 & \new_[29460]_ ;
  assign \new_[29462]_  = \new_[29461]_  & \new_[29456]_ ;
  assign \new_[29466]_  = A199 & A166;
  assign \new_[29467]_  = A168 & \new_[29466]_ ;
  assign \new_[29471]_  = ~A202 & ~A201;
  assign \new_[29472]_  = A200 & \new_[29471]_ ;
  assign \new_[29473]_  = \new_[29472]_  & \new_[29467]_ ;
  assign \new_[29477]_  = A236 & A233;
  assign \new_[29478]_  = ~A232 & \new_[29477]_ ;
  assign \new_[29482]_  = A302 & A299;
  assign \new_[29483]_  = ~A298 & \new_[29482]_ ;
  assign \new_[29484]_  = \new_[29483]_  & \new_[29478]_ ;
  assign \new_[29488]_  = A199 & A166;
  assign \new_[29489]_  = A168 & \new_[29488]_ ;
  assign \new_[29493]_  = ~A202 & ~A201;
  assign \new_[29494]_  = A200 & \new_[29493]_ ;
  assign \new_[29495]_  = \new_[29494]_  & \new_[29489]_ ;
  assign \new_[29499]_  = A236 & A233;
  assign \new_[29500]_  = ~A232 & \new_[29499]_ ;
  assign \new_[29504]_  = A269 & A266;
  assign \new_[29505]_  = ~A265 & \new_[29504]_ ;
  assign \new_[29506]_  = \new_[29505]_  & \new_[29500]_ ;
  assign \new_[29510]_  = A199 & A166;
  assign \new_[29511]_  = A168 & \new_[29510]_ ;
  assign \new_[29515]_  = ~A202 & ~A201;
  assign \new_[29516]_  = A200 & \new_[29515]_ ;
  assign \new_[29517]_  = \new_[29516]_  & \new_[29511]_ ;
  assign \new_[29521]_  = A236 & A233;
  assign \new_[29522]_  = ~A232 & \new_[29521]_ ;
  assign \new_[29526]_  = A269 & ~A266;
  assign \new_[29527]_  = A265 & \new_[29526]_ ;
  assign \new_[29528]_  = \new_[29527]_  & \new_[29522]_ ;
  assign \new_[29532]_  = A199 & A166;
  assign \new_[29533]_  = A168 & \new_[29532]_ ;
  assign \new_[29537]_  = ~A202 & ~A201;
  assign \new_[29538]_  = A200 & \new_[29537]_ ;
  assign \new_[29539]_  = \new_[29538]_  & \new_[29533]_ ;
  assign \new_[29543]_  = A236 & ~A233;
  assign \new_[29544]_  = A232 & \new_[29543]_ ;
  assign \new_[29548]_  = A302 & ~A299;
  assign \new_[29549]_  = A298 & \new_[29548]_ ;
  assign \new_[29550]_  = \new_[29549]_  & \new_[29544]_ ;
  assign \new_[29554]_  = A199 & A166;
  assign \new_[29555]_  = A168 & \new_[29554]_ ;
  assign \new_[29559]_  = ~A202 & ~A201;
  assign \new_[29560]_  = A200 & \new_[29559]_ ;
  assign \new_[29561]_  = \new_[29560]_  & \new_[29555]_ ;
  assign \new_[29565]_  = A236 & ~A233;
  assign \new_[29566]_  = A232 & \new_[29565]_ ;
  assign \new_[29570]_  = A302 & A299;
  assign \new_[29571]_  = ~A298 & \new_[29570]_ ;
  assign \new_[29572]_  = \new_[29571]_  & \new_[29566]_ ;
  assign \new_[29576]_  = A199 & A166;
  assign \new_[29577]_  = A168 & \new_[29576]_ ;
  assign \new_[29581]_  = ~A202 & ~A201;
  assign \new_[29582]_  = A200 & \new_[29581]_ ;
  assign \new_[29583]_  = \new_[29582]_  & \new_[29577]_ ;
  assign \new_[29587]_  = A236 & ~A233;
  assign \new_[29588]_  = A232 & \new_[29587]_ ;
  assign \new_[29592]_  = A269 & A266;
  assign \new_[29593]_  = ~A265 & \new_[29592]_ ;
  assign \new_[29594]_  = \new_[29593]_  & \new_[29588]_ ;
  assign \new_[29598]_  = A199 & A166;
  assign \new_[29599]_  = A168 & \new_[29598]_ ;
  assign \new_[29603]_  = ~A202 & ~A201;
  assign \new_[29604]_  = A200 & \new_[29603]_ ;
  assign \new_[29605]_  = \new_[29604]_  & \new_[29599]_ ;
  assign \new_[29609]_  = A236 & ~A233;
  assign \new_[29610]_  = A232 & \new_[29609]_ ;
  assign \new_[29614]_  = A269 & ~A266;
  assign \new_[29615]_  = A265 & \new_[29614]_ ;
  assign \new_[29616]_  = \new_[29615]_  & \new_[29610]_ ;
  assign \new_[29620]_  = A199 & A167;
  assign \new_[29621]_  = A168 & \new_[29620]_ ;
  assign \new_[29625]_  = ~A202 & ~A201;
  assign \new_[29626]_  = A200 & \new_[29625]_ ;
  assign \new_[29627]_  = \new_[29626]_  & \new_[29621]_ ;
  assign \new_[29631]_  = A236 & A233;
  assign \new_[29632]_  = ~A232 & \new_[29631]_ ;
  assign \new_[29636]_  = A302 & ~A299;
  assign \new_[29637]_  = A298 & \new_[29636]_ ;
  assign \new_[29638]_  = \new_[29637]_  & \new_[29632]_ ;
  assign \new_[29642]_  = A199 & A167;
  assign \new_[29643]_  = A168 & \new_[29642]_ ;
  assign \new_[29647]_  = ~A202 & ~A201;
  assign \new_[29648]_  = A200 & \new_[29647]_ ;
  assign \new_[29649]_  = \new_[29648]_  & \new_[29643]_ ;
  assign \new_[29653]_  = A236 & A233;
  assign \new_[29654]_  = ~A232 & \new_[29653]_ ;
  assign \new_[29658]_  = A302 & A299;
  assign \new_[29659]_  = ~A298 & \new_[29658]_ ;
  assign \new_[29660]_  = \new_[29659]_  & \new_[29654]_ ;
  assign \new_[29664]_  = A199 & A167;
  assign \new_[29665]_  = A168 & \new_[29664]_ ;
  assign \new_[29669]_  = ~A202 & ~A201;
  assign \new_[29670]_  = A200 & \new_[29669]_ ;
  assign \new_[29671]_  = \new_[29670]_  & \new_[29665]_ ;
  assign \new_[29675]_  = A236 & A233;
  assign \new_[29676]_  = ~A232 & \new_[29675]_ ;
  assign \new_[29680]_  = A269 & A266;
  assign \new_[29681]_  = ~A265 & \new_[29680]_ ;
  assign \new_[29682]_  = \new_[29681]_  & \new_[29676]_ ;
  assign \new_[29686]_  = A199 & A167;
  assign \new_[29687]_  = A168 & \new_[29686]_ ;
  assign \new_[29691]_  = ~A202 & ~A201;
  assign \new_[29692]_  = A200 & \new_[29691]_ ;
  assign \new_[29693]_  = \new_[29692]_  & \new_[29687]_ ;
  assign \new_[29697]_  = A236 & A233;
  assign \new_[29698]_  = ~A232 & \new_[29697]_ ;
  assign \new_[29702]_  = A269 & ~A266;
  assign \new_[29703]_  = A265 & \new_[29702]_ ;
  assign \new_[29704]_  = \new_[29703]_  & \new_[29698]_ ;
  assign \new_[29708]_  = A199 & A167;
  assign \new_[29709]_  = A168 & \new_[29708]_ ;
  assign \new_[29713]_  = ~A202 & ~A201;
  assign \new_[29714]_  = A200 & \new_[29713]_ ;
  assign \new_[29715]_  = \new_[29714]_  & \new_[29709]_ ;
  assign \new_[29719]_  = A236 & ~A233;
  assign \new_[29720]_  = A232 & \new_[29719]_ ;
  assign \new_[29724]_  = A302 & ~A299;
  assign \new_[29725]_  = A298 & \new_[29724]_ ;
  assign \new_[29726]_  = \new_[29725]_  & \new_[29720]_ ;
  assign \new_[29730]_  = A199 & A167;
  assign \new_[29731]_  = A168 & \new_[29730]_ ;
  assign \new_[29735]_  = ~A202 & ~A201;
  assign \new_[29736]_  = A200 & \new_[29735]_ ;
  assign \new_[29737]_  = \new_[29736]_  & \new_[29731]_ ;
  assign \new_[29741]_  = A236 & ~A233;
  assign \new_[29742]_  = A232 & \new_[29741]_ ;
  assign \new_[29746]_  = A302 & A299;
  assign \new_[29747]_  = ~A298 & \new_[29746]_ ;
  assign \new_[29748]_  = \new_[29747]_  & \new_[29742]_ ;
  assign \new_[29752]_  = A199 & A167;
  assign \new_[29753]_  = A168 & \new_[29752]_ ;
  assign \new_[29757]_  = ~A202 & ~A201;
  assign \new_[29758]_  = A200 & \new_[29757]_ ;
  assign \new_[29759]_  = \new_[29758]_  & \new_[29753]_ ;
  assign \new_[29763]_  = A236 & ~A233;
  assign \new_[29764]_  = A232 & \new_[29763]_ ;
  assign \new_[29768]_  = A269 & A266;
  assign \new_[29769]_  = ~A265 & \new_[29768]_ ;
  assign \new_[29770]_  = \new_[29769]_  & \new_[29764]_ ;
  assign \new_[29774]_  = A199 & A167;
  assign \new_[29775]_  = A168 & \new_[29774]_ ;
  assign \new_[29779]_  = ~A202 & ~A201;
  assign \new_[29780]_  = A200 & \new_[29779]_ ;
  assign \new_[29781]_  = \new_[29780]_  & \new_[29775]_ ;
  assign \new_[29785]_  = A236 & ~A233;
  assign \new_[29786]_  = A232 & \new_[29785]_ ;
  assign \new_[29790]_  = A269 & ~A266;
  assign \new_[29791]_  = A265 & \new_[29790]_ ;
  assign \new_[29792]_  = \new_[29791]_  & \new_[29786]_ ;
  assign \new_[29796]_  = ~A166 & A167;
  assign \new_[29797]_  = A170 & \new_[29796]_ ;
  assign \new_[29801]_  = ~A203 & ~A202;
  assign \new_[29802]_  = ~A201 & \new_[29801]_ ;
  assign \new_[29803]_  = \new_[29802]_  & \new_[29797]_ ;
  assign \new_[29807]_  = A236 & A233;
  assign \new_[29808]_  = ~A232 & \new_[29807]_ ;
  assign \new_[29812]_  = A302 & ~A299;
  assign \new_[29813]_  = A298 & \new_[29812]_ ;
  assign \new_[29814]_  = \new_[29813]_  & \new_[29808]_ ;
  assign \new_[29818]_  = ~A166 & A167;
  assign \new_[29819]_  = A170 & \new_[29818]_ ;
  assign \new_[29823]_  = ~A203 & ~A202;
  assign \new_[29824]_  = ~A201 & \new_[29823]_ ;
  assign \new_[29825]_  = \new_[29824]_  & \new_[29819]_ ;
  assign \new_[29829]_  = A236 & A233;
  assign \new_[29830]_  = ~A232 & \new_[29829]_ ;
  assign \new_[29834]_  = A302 & A299;
  assign \new_[29835]_  = ~A298 & \new_[29834]_ ;
  assign \new_[29836]_  = \new_[29835]_  & \new_[29830]_ ;
  assign \new_[29840]_  = ~A166 & A167;
  assign \new_[29841]_  = A170 & \new_[29840]_ ;
  assign \new_[29845]_  = ~A203 & ~A202;
  assign \new_[29846]_  = ~A201 & \new_[29845]_ ;
  assign \new_[29847]_  = \new_[29846]_  & \new_[29841]_ ;
  assign \new_[29851]_  = A236 & A233;
  assign \new_[29852]_  = ~A232 & \new_[29851]_ ;
  assign \new_[29856]_  = A269 & A266;
  assign \new_[29857]_  = ~A265 & \new_[29856]_ ;
  assign \new_[29858]_  = \new_[29857]_  & \new_[29852]_ ;
  assign \new_[29862]_  = ~A166 & A167;
  assign \new_[29863]_  = A170 & \new_[29862]_ ;
  assign \new_[29867]_  = ~A203 & ~A202;
  assign \new_[29868]_  = ~A201 & \new_[29867]_ ;
  assign \new_[29869]_  = \new_[29868]_  & \new_[29863]_ ;
  assign \new_[29873]_  = A236 & A233;
  assign \new_[29874]_  = ~A232 & \new_[29873]_ ;
  assign \new_[29878]_  = A269 & ~A266;
  assign \new_[29879]_  = A265 & \new_[29878]_ ;
  assign \new_[29880]_  = \new_[29879]_  & \new_[29874]_ ;
  assign \new_[29884]_  = ~A166 & A167;
  assign \new_[29885]_  = A170 & \new_[29884]_ ;
  assign \new_[29889]_  = ~A203 & ~A202;
  assign \new_[29890]_  = ~A201 & \new_[29889]_ ;
  assign \new_[29891]_  = \new_[29890]_  & \new_[29885]_ ;
  assign \new_[29895]_  = A236 & ~A233;
  assign \new_[29896]_  = A232 & \new_[29895]_ ;
  assign \new_[29900]_  = A302 & ~A299;
  assign \new_[29901]_  = A298 & \new_[29900]_ ;
  assign \new_[29902]_  = \new_[29901]_  & \new_[29896]_ ;
  assign \new_[29906]_  = ~A166 & A167;
  assign \new_[29907]_  = A170 & \new_[29906]_ ;
  assign \new_[29911]_  = ~A203 & ~A202;
  assign \new_[29912]_  = ~A201 & \new_[29911]_ ;
  assign \new_[29913]_  = \new_[29912]_  & \new_[29907]_ ;
  assign \new_[29917]_  = A236 & ~A233;
  assign \new_[29918]_  = A232 & \new_[29917]_ ;
  assign \new_[29922]_  = A302 & A299;
  assign \new_[29923]_  = ~A298 & \new_[29922]_ ;
  assign \new_[29924]_  = \new_[29923]_  & \new_[29918]_ ;
  assign \new_[29928]_  = ~A166 & A167;
  assign \new_[29929]_  = A170 & \new_[29928]_ ;
  assign \new_[29933]_  = ~A203 & ~A202;
  assign \new_[29934]_  = ~A201 & \new_[29933]_ ;
  assign \new_[29935]_  = \new_[29934]_  & \new_[29929]_ ;
  assign \new_[29939]_  = A236 & ~A233;
  assign \new_[29940]_  = A232 & \new_[29939]_ ;
  assign \new_[29944]_  = A269 & A266;
  assign \new_[29945]_  = ~A265 & \new_[29944]_ ;
  assign \new_[29946]_  = \new_[29945]_  & \new_[29940]_ ;
  assign \new_[29950]_  = ~A166 & A167;
  assign \new_[29951]_  = A170 & \new_[29950]_ ;
  assign \new_[29955]_  = ~A203 & ~A202;
  assign \new_[29956]_  = ~A201 & \new_[29955]_ ;
  assign \new_[29957]_  = \new_[29956]_  & \new_[29951]_ ;
  assign \new_[29961]_  = A236 & ~A233;
  assign \new_[29962]_  = A232 & \new_[29961]_ ;
  assign \new_[29966]_  = A269 & ~A266;
  assign \new_[29967]_  = A265 & \new_[29966]_ ;
  assign \new_[29968]_  = \new_[29967]_  & \new_[29962]_ ;
  assign \new_[29972]_  = ~A166 & A167;
  assign \new_[29973]_  = A170 & \new_[29972]_ ;
  assign \new_[29977]_  = ~A201 & A200;
  assign \new_[29978]_  = A199 & \new_[29977]_ ;
  assign \new_[29979]_  = \new_[29978]_  & \new_[29973]_ ;
  assign \new_[29983]_  = A234 & A232;
  assign \new_[29984]_  = ~A202 & \new_[29983]_ ;
  assign \new_[29988]_  = A302 & ~A299;
  assign \new_[29989]_  = A298 & \new_[29988]_ ;
  assign \new_[29990]_  = \new_[29989]_  & \new_[29984]_ ;
  assign \new_[29994]_  = ~A166 & A167;
  assign \new_[29995]_  = A170 & \new_[29994]_ ;
  assign \new_[29999]_  = ~A201 & A200;
  assign \new_[30000]_  = A199 & \new_[29999]_ ;
  assign \new_[30001]_  = \new_[30000]_  & \new_[29995]_ ;
  assign \new_[30005]_  = A234 & A232;
  assign \new_[30006]_  = ~A202 & \new_[30005]_ ;
  assign \new_[30010]_  = A302 & A299;
  assign \new_[30011]_  = ~A298 & \new_[30010]_ ;
  assign \new_[30012]_  = \new_[30011]_  & \new_[30006]_ ;
  assign \new_[30016]_  = ~A166 & A167;
  assign \new_[30017]_  = A170 & \new_[30016]_ ;
  assign \new_[30021]_  = ~A201 & A200;
  assign \new_[30022]_  = A199 & \new_[30021]_ ;
  assign \new_[30023]_  = \new_[30022]_  & \new_[30017]_ ;
  assign \new_[30027]_  = A234 & A232;
  assign \new_[30028]_  = ~A202 & \new_[30027]_ ;
  assign \new_[30032]_  = A269 & A266;
  assign \new_[30033]_  = ~A265 & \new_[30032]_ ;
  assign \new_[30034]_  = \new_[30033]_  & \new_[30028]_ ;
  assign \new_[30038]_  = ~A166 & A167;
  assign \new_[30039]_  = A170 & \new_[30038]_ ;
  assign \new_[30043]_  = ~A201 & A200;
  assign \new_[30044]_  = A199 & \new_[30043]_ ;
  assign \new_[30045]_  = \new_[30044]_  & \new_[30039]_ ;
  assign \new_[30049]_  = A234 & A232;
  assign \new_[30050]_  = ~A202 & \new_[30049]_ ;
  assign \new_[30054]_  = A269 & ~A266;
  assign \new_[30055]_  = A265 & \new_[30054]_ ;
  assign \new_[30056]_  = \new_[30055]_  & \new_[30050]_ ;
  assign \new_[30060]_  = ~A166 & A167;
  assign \new_[30061]_  = A170 & \new_[30060]_ ;
  assign \new_[30065]_  = ~A201 & A200;
  assign \new_[30066]_  = A199 & \new_[30065]_ ;
  assign \new_[30067]_  = \new_[30066]_  & \new_[30061]_ ;
  assign \new_[30071]_  = A234 & A233;
  assign \new_[30072]_  = ~A202 & \new_[30071]_ ;
  assign \new_[30076]_  = A302 & ~A299;
  assign \new_[30077]_  = A298 & \new_[30076]_ ;
  assign \new_[30078]_  = \new_[30077]_  & \new_[30072]_ ;
  assign \new_[30082]_  = ~A166 & A167;
  assign \new_[30083]_  = A170 & \new_[30082]_ ;
  assign \new_[30087]_  = ~A201 & A200;
  assign \new_[30088]_  = A199 & \new_[30087]_ ;
  assign \new_[30089]_  = \new_[30088]_  & \new_[30083]_ ;
  assign \new_[30093]_  = A234 & A233;
  assign \new_[30094]_  = ~A202 & \new_[30093]_ ;
  assign \new_[30098]_  = A302 & A299;
  assign \new_[30099]_  = ~A298 & \new_[30098]_ ;
  assign \new_[30100]_  = \new_[30099]_  & \new_[30094]_ ;
  assign \new_[30104]_  = ~A166 & A167;
  assign \new_[30105]_  = A170 & \new_[30104]_ ;
  assign \new_[30109]_  = ~A201 & A200;
  assign \new_[30110]_  = A199 & \new_[30109]_ ;
  assign \new_[30111]_  = \new_[30110]_  & \new_[30105]_ ;
  assign \new_[30115]_  = A234 & A233;
  assign \new_[30116]_  = ~A202 & \new_[30115]_ ;
  assign \new_[30120]_  = A269 & A266;
  assign \new_[30121]_  = ~A265 & \new_[30120]_ ;
  assign \new_[30122]_  = \new_[30121]_  & \new_[30116]_ ;
  assign \new_[30126]_  = ~A166 & A167;
  assign \new_[30127]_  = A170 & \new_[30126]_ ;
  assign \new_[30131]_  = ~A201 & A200;
  assign \new_[30132]_  = A199 & \new_[30131]_ ;
  assign \new_[30133]_  = \new_[30132]_  & \new_[30127]_ ;
  assign \new_[30137]_  = A234 & A233;
  assign \new_[30138]_  = ~A202 & \new_[30137]_ ;
  assign \new_[30142]_  = A269 & ~A266;
  assign \new_[30143]_  = A265 & \new_[30142]_ ;
  assign \new_[30144]_  = \new_[30143]_  & \new_[30138]_ ;
  assign \new_[30148]_  = ~A166 & A167;
  assign \new_[30149]_  = A170 & \new_[30148]_ ;
  assign \new_[30153]_  = ~A201 & A200;
  assign \new_[30154]_  = A199 & \new_[30153]_ ;
  assign \new_[30155]_  = \new_[30154]_  & \new_[30149]_ ;
  assign \new_[30159]_  = A233 & ~A232;
  assign \new_[30160]_  = ~A202 & \new_[30159]_ ;
  assign \new_[30164]_  = A300 & A299;
  assign \new_[30165]_  = A236 & \new_[30164]_ ;
  assign \new_[30166]_  = \new_[30165]_  & \new_[30160]_ ;
  assign \new_[30170]_  = ~A166 & A167;
  assign \new_[30171]_  = A170 & \new_[30170]_ ;
  assign \new_[30175]_  = ~A201 & A200;
  assign \new_[30176]_  = A199 & \new_[30175]_ ;
  assign \new_[30177]_  = \new_[30176]_  & \new_[30171]_ ;
  assign \new_[30181]_  = A233 & ~A232;
  assign \new_[30182]_  = ~A202 & \new_[30181]_ ;
  assign \new_[30186]_  = A300 & A298;
  assign \new_[30187]_  = A236 & \new_[30186]_ ;
  assign \new_[30188]_  = \new_[30187]_  & \new_[30182]_ ;
  assign \new_[30192]_  = ~A166 & A167;
  assign \new_[30193]_  = A170 & \new_[30192]_ ;
  assign \new_[30197]_  = ~A201 & A200;
  assign \new_[30198]_  = A199 & \new_[30197]_ ;
  assign \new_[30199]_  = \new_[30198]_  & \new_[30193]_ ;
  assign \new_[30203]_  = A233 & ~A232;
  assign \new_[30204]_  = ~A202 & \new_[30203]_ ;
  assign \new_[30208]_  = A267 & A265;
  assign \new_[30209]_  = A236 & \new_[30208]_ ;
  assign \new_[30210]_  = \new_[30209]_  & \new_[30204]_ ;
  assign \new_[30214]_  = ~A166 & A167;
  assign \new_[30215]_  = A170 & \new_[30214]_ ;
  assign \new_[30219]_  = ~A201 & A200;
  assign \new_[30220]_  = A199 & \new_[30219]_ ;
  assign \new_[30221]_  = \new_[30220]_  & \new_[30215]_ ;
  assign \new_[30225]_  = A233 & ~A232;
  assign \new_[30226]_  = ~A202 & \new_[30225]_ ;
  assign \new_[30230]_  = A267 & A266;
  assign \new_[30231]_  = A236 & \new_[30230]_ ;
  assign \new_[30232]_  = \new_[30231]_  & \new_[30226]_ ;
  assign \new_[30236]_  = ~A166 & A167;
  assign \new_[30237]_  = A170 & \new_[30236]_ ;
  assign \new_[30241]_  = ~A201 & A200;
  assign \new_[30242]_  = A199 & \new_[30241]_ ;
  assign \new_[30243]_  = \new_[30242]_  & \new_[30237]_ ;
  assign \new_[30247]_  = ~A233 & A232;
  assign \new_[30248]_  = ~A202 & \new_[30247]_ ;
  assign \new_[30252]_  = A300 & A299;
  assign \new_[30253]_  = A236 & \new_[30252]_ ;
  assign \new_[30254]_  = \new_[30253]_  & \new_[30248]_ ;
  assign \new_[30258]_  = ~A166 & A167;
  assign \new_[30259]_  = A170 & \new_[30258]_ ;
  assign \new_[30263]_  = ~A201 & A200;
  assign \new_[30264]_  = A199 & \new_[30263]_ ;
  assign \new_[30265]_  = \new_[30264]_  & \new_[30259]_ ;
  assign \new_[30269]_  = ~A233 & A232;
  assign \new_[30270]_  = ~A202 & \new_[30269]_ ;
  assign \new_[30274]_  = A300 & A298;
  assign \new_[30275]_  = A236 & \new_[30274]_ ;
  assign \new_[30276]_  = \new_[30275]_  & \new_[30270]_ ;
  assign \new_[30280]_  = ~A166 & A167;
  assign \new_[30281]_  = A170 & \new_[30280]_ ;
  assign \new_[30285]_  = ~A201 & A200;
  assign \new_[30286]_  = A199 & \new_[30285]_ ;
  assign \new_[30287]_  = \new_[30286]_  & \new_[30281]_ ;
  assign \new_[30291]_  = ~A233 & A232;
  assign \new_[30292]_  = ~A202 & \new_[30291]_ ;
  assign \new_[30296]_  = A267 & A265;
  assign \new_[30297]_  = A236 & \new_[30296]_ ;
  assign \new_[30298]_  = \new_[30297]_  & \new_[30292]_ ;
  assign \new_[30302]_  = ~A166 & A167;
  assign \new_[30303]_  = A170 & \new_[30302]_ ;
  assign \new_[30307]_  = ~A201 & A200;
  assign \new_[30308]_  = A199 & \new_[30307]_ ;
  assign \new_[30309]_  = \new_[30308]_  & \new_[30303]_ ;
  assign \new_[30313]_  = ~A233 & A232;
  assign \new_[30314]_  = ~A202 & \new_[30313]_ ;
  assign \new_[30318]_  = A267 & A266;
  assign \new_[30319]_  = A236 & \new_[30318]_ ;
  assign \new_[30320]_  = \new_[30319]_  & \new_[30314]_ ;
  assign \new_[30324]_  = ~A166 & A167;
  assign \new_[30325]_  = A170 & \new_[30324]_ ;
  assign \new_[30329]_  = ~A202 & ~A200;
  assign \new_[30330]_  = ~A199 & \new_[30329]_ ;
  assign \new_[30331]_  = \new_[30330]_  & \new_[30325]_ ;
  assign \new_[30335]_  = A236 & A233;
  assign \new_[30336]_  = ~A232 & \new_[30335]_ ;
  assign \new_[30340]_  = A302 & ~A299;
  assign \new_[30341]_  = A298 & \new_[30340]_ ;
  assign \new_[30342]_  = \new_[30341]_  & \new_[30336]_ ;
  assign \new_[30346]_  = ~A166 & A167;
  assign \new_[30347]_  = A170 & \new_[30346]_ ;
  assign \new_[30351]_  = ~A202 & ~A200;
  assign \new_[30352]_  = ~A199 & \new_[30351]_ ;
  assign \new_[30353]_  = \new_[30352]_  & \new_[30347]_ ;
  assign \new_[30357]_  = A236 & A233;
  assign \new_[30358]_  = ~A232 & \new_[30357]_ ;
  assign \new_[30362]_  = A302 & A299;
  assign \new_[30363]_  = ~A298 & \new_[30362]_ ;
  assign \new_[30364]_  = \new_[30363]_  & \new_[30358]_ ;
  assign \new_[30368]_  = ~A166 & A167;
  assign \new_[30369]_  = A170 & \new_[30368]_ ;
  assign \new_[30373]_  = ~A202 & ~A200;
  assign \new_[30374]_  = ~A199 & \new_[30373]_ ;
  assign \new_[30375]_  = \new_[30374]_  & \new_[30369]_ ;
  assign \new_[30379]_  = A236 & A233;
  assign \new_[30380]_  = ~A232 & \new_[30379]_ ;
  assign \new_[30384]_  = A269 & A266;
  assign \new_[30385]_  = ~A265 & \new_[30384]_ ;
  assign \new_[30386]_  = \new_[30385]_  & \new_[30380]_ ;
  assign \new_[30390]_  = ~A166 & A167;
  assign \new_[30391]_  = A170 & \new_[30390]_ ;
  assign \new_[30395]_  = ~A202 & ~A200;
  assign \new_[30396]_  = ~A199 & \new_[30395]_ ;
  assign \new_[30397]_  = \new_[30396]_  & \new_[30391]_ ;
  assign \new_[30401]_  = A236 & A233;
  assign \new_[30402]_  = ~A232 & \new_[30401]_ ;
  assign \new_[30406]_  = A269 & ~A266;
  assign \new_[30407]_  = A265 & \new_[30406]_ ;
  assign \new_[30408]_  = \new_[30407]_  & \new_[30402]_ ;
  assign \new_[30412]_  = ~A166 & A167;
  assign \new_[30413]_  = A170 & \new_[30412]_ ;
  assign \new_[30417]_  = ~A202 & ~A200;
  assign \new_[30418]_  = ~A199 & \new_[30417]_ ;
  assign \new_[30419]_  = \new_[30418]_  & \new_[30413]_ ;
  assign \new_[30423]_  = A236 & ~A233;
  assign \new_[30424]_  = A232 & \new_[30423]_ ;
  assign \new_[30428]_  = A302 & ~A299;
  assign \new_[30429]_  = A298 & \new_[30428]_ ;
  assign \new_[30430]_  = \new_[30429]_  & \new_[30424]_ ;
  assign \new_[30434]_  = ~A166 & A167;
  assign \new_[30435]_  = A170 & \new_[30434]_ ;
  assign \new_[30439]_  = ~A202 & ~A200;
  assign \new_[30440]_  = ~A199 & \new_[30439]_ ;
  assign \new_[30441]_  = \new_[30440]_  & \new_[30435]_ ;
  assign \new_[30445]_  = A236 & ~A233;
  assign \new_[30446]_  = A232 & \new_[30445]_ ;
  assign \new_[30450]_  = A302 & A299;
  assign \new_[30451]_  = ~A298 & \new_[30450]_ ;
  assign \new_[30452]_  = \new_[30451]_  & \new_[30446]_ ;
  assign \new_[30456]_  = ~A166 & A167;
  assign \new_[30457]_  = A170 & \new_[30456]_ ;
  assign \new_[30461]_  = ~A202 & ~A200;
  assign \new_[30462]_  = ~A199 & \new_[30461]_ ;
  assign \new_[30463]_  = \new_[30462]_  & \new_[30457]_ ;
  assign \new_[30467]_  = A236 & ~A233;
  assign \new_[30468]_  = A232 & \new_[30467]_ ;
  assign \new_[30472]_  = A269 & A266;
  assign \new_[30473]_  = ~A265 & \new_[30472]_ ;
  assign \new_[30474]_  = \new_[30473]_  & \new_[30468]_ ;
  assign \new_[30478]_  = ~A166 & A167;
  assign \new_[30479]_  = A170 & \new_[30478]_ ;
  assign \new_[30483]_  = ~A202 & ~A200;
  assign \new_[30484]_  = ~A199 & \new_[30483]_ ;
  assign \new_[30485]_  = \new_[30484]_  & \new_[30479]_ ;
  assign \new_[30489]_  = A236 & ~A233;
  assign \new_[30490]_  = A232 & \new_[30489]_ ;
  assign \new_[30494]_  = A269 & ~A266;
  assign \new_[30495]_  = A265 & \new_[30494]_ ;
  assign \new_[30496]_  = \new_[30495]_  & \new_[30490]_ ;
  assign \new_[30500]_  = A166 & ~A167;
  assign \new_[30501]_  = A170 & \new_[30500]_ ;
  assign \new_[30505]_  = ~A203 & ~A202;
  assign \new_[30506]_  = ~A201 & \new_[30505]_ ;
  assign \new_[30507]_  = \new_[30506]_  & \new_[30501]_ ;
  assign \new_[30511]_  = A236 & A233;
  assign \new_[30512]_  = ~A232 & \new_[30511]_ ;
  assign \new_[30516]_  = A302 & ~A299;
  assign \new_[30517]_  = A298 & \new_[30516]_ ;
  assign \new_[30518]_  = \new_[30517]_  & \new_[30512]_ ;
  assign \new_[30522]_  = A166 & ~A167;
  assign \new_[30523]_  = A170 & \new_[30522]_ ;
  assign \new_[30527]_  = ~A203 & ~A202;
  assign \new_[30528]_  = ~A201 & \new_[30527]_ ;
  assign \new_[30529]_  = \new_[30528]_  & \new_[30523]_ ;
  assign \new_[30533]_  = A236 & A233;
  assign \new_[30534]_  = ~A232 & \new_[30533]_ ;
  assign \new_[30538]_  = A302 & A299;
  assign \new_[30539]_  = ~A298 & \new_[30538]_ ;
  assign \new_[30540]_  = \new_[30539]_  & \new_[30534]_ ;
  assign \new_[30544]_  = A166 & ~A167;
  assign \new_[30545]_  = A170 & \new_[30544]_ ;
  assign \new_[30549]_  = ~A203 & ~A202;
  assign \new_[30550]_  = ~A201 & \new_[30549]_ ;
  assign \new_[30551]_  = \new_[30550]_  & \new_[30545]_ ;
  assign \new_[30555]_  = A236 & A233;
  assign \new_[30556]_  = ~A232 & \new_[30555]_ ;
  assign \new_[30560]_  = A269 & A266;
  assign \new_[30561]_  = ~A265 & \new_[30560]_ ;
  assign \new_[30562]_  = \new_[30561]_  & \new_[30556]_ ;
  assign \new_[30566]_  = A166 & ~A167;
  assign \new_[30567]_  = A170 & \new_[30566]_ ;
  assign \new_[30571]_  = ~A203 & ~A202;
  assign \new_[30572]_  = ~A201 & \new_[30571]_ ;
  assign \new_[30573]_  = \new_[30572]_  & \new_[30567]_ ;
  assign \new_[30577]_  = A236 & A233;
  assign \new_[30578]_  = ~A232 & \new_[30577]_ ;
  assign \new_[30582]_  = A269 & ~A266;
  assign \new_[30583]_  = A265 & \new_[30582]_ ;
  assign \new_[30584]_  = \new_[30583]_  & \new_[30578]_ ;
  assign \new_[30588]_  = A166 & ~A167;
  assign \new_[30589]_  = A170 & \new_[30588]_ ;
  assign \new_[30593]_  = ~A203 & ~A202;
  assign \new_[30594]_  = ~A201 & \new_[30593]_ ;
  assign \new_[30595]_  = \new_[30594]_  & \new_[30589]_ ;
  assign \new_[30599]_  = A236 & ~A233;
  assign \new_[30600]_  = A232 & \new_[30599]_ ;
  assign \new_[30604]_  = A302 & ~A299;
  assign \new_[30605]_  = A298 & \new_[30604]_ ;
  assign \new_[30606]_  = \new_[30605]_  & \new_[30600]_ ;
  assign \new_[30610]_  = A166 & ~A167;
  assign \new_[30611]_  = A170 & \new_[30610]_ ;
  assign \new_[30615]_  = ~A203 & ~A202;
  assign \new_[30616]_  = ~A201 & \new_[30615]_ ;
  assign \new_[30617]_  = \new_[30616]_  & \new_[30611]_ ;
  assign \new_[30621]_  = A236 & ~A233;
  assign \new_[30622]_  = A232 & \new_[30621]_ ;
  assign \new_[30626]_  = A302 & A299;
  assign \new_[30627]_  = ~A298 & \new_[30626]_ ;
  assign \new_[30628]_  = \new_[30627]_  & \new_[30622]_ ;
  assign \new_[30632]_  = A166 & ~A167;
  assign \new_[30633]_  = A170 & \new_[30632]_ ;
  assign \new_[30637]_  = ~A203 & ~A202;
  assign \new_[30638]_  = ~A201 & \new_[30637]_ ;
  assign \new_[30639]_  = \new_[30638]_  & \new_[30633]_ ;
  assign \new_[30643]_  = A236 & ~A233;
  assign \new_[30644]_  = A232 & \new_[30643]_ ;
  assign \new_[30648]_  = A269 & A266;
  assign \new_[30649]_  = ~A265 & \new_[30648]_ ;
  assign \new_[30650]_  = \new_[30649]_  & \new_[30644]_ ;
  assign \new_[30654]_  = A166 & ~A167;
  assign \new_[30655]_  = A170 & \new_[30654]_ ;
  assign \new_[30659]_  = ~A203 & ~A202;
  assign \new_[30660]_  = ~A201 & \new_[30659]_ ;
  assign \new_[30661]_  = \new_[30660]_  & \new_[30655]_ ;
  assign \new_[30665]_  = A236 & ~A233;
  assign \new_[30666]_  = A232 & \new_[30665]_ ;
  assign \new_[30670]_  = A269 & ~A266;
  assign \new_[30671]_  = A265 & \new_[30670]_ ;
  assign \new_[30672]_  = \new_[30671]_  & \new_[30666]_ ;
  assign \new_[30676]_  = A166 & ~A167;
  assign \new_[30677]_  = A170 & \new_[30676]_ ;
  assign \new_[30681]_  = ~A201 & A200;
  assign \new_[30682]_  = A199 & \new_[30681]_ ;
  assign \new_[30683]_  = \new_[30682]_  & \new_[30677]_ ;
  assign \new_[30687]_  = A234 & A232;
  assign \new_[30688]_  = ~A202 & \new_[30687]_ ;
  assign \new_[30692]_  = A302 & ~A299;
  assign \new_[30693]_  = A298 & \new_[30692]_ ;
  assign \new_[30694]_  = \new_[30693]_  & \new_[30688]_ ;
  assign \new_[30698]_  = A166 & ~A167;
  assign \new_[30699]_  = A170 & \new_[30698]_ ;
  assign \new_[30703]_  = ~A201 & A200;
  assign \new_[30704]_  = A199 & \new_[30703]_ ;
  assign \new_[30705]_  = \new_[30704]_  & \new_[30699]_ ;
  assign \new_[30709]_  = A234 & A232;
  assign \new_[30710]_  = ~A202 & \new_[30709]_ ;
  assign \new_[30714]_  = A302 & A299;
  assign \new_[30715]_  = ~A298 & \new_[30714]_ ;
  assign \new_[30716]_  = \new_[30715]_  & \new_[30710]_ ;
  assign \new_[30720]_  = A166 & ~A167;
  assign \new_[30721]_  = A170 & \new_[30720]_ ;
  assign \new_[30725]_  = ~A201 & A200;
  assign \new_[30726]_  = A199 & \new_[30725]_ ;
  assign \new_[30727]_  = \new_[30726]_  & \new_[30721]_ ;
  assign \new_[30731]_  = A234 & A232;
  assign \new_[30732]_  = ~A202 & \new_[30731]_ ;
  assign \new_[30736]_  = A269 & A266;
  assign \new_[30737]_  = ~A265 & \new_[30736]_ ;
  assign \new_[30738]_  = \new_[30737]_  & \new_[30732]_ ;
  assign \new_[30742]_  = A166 & ~A167;
  assign \new_[30743]_  = A170 & \new_[30742]_ ;
  assign \new_[30747]_  = ~A201 & A200;
  assign \new_[30748]_  = A199 & \new_[30747]_ ;
  assign \new_[30749]_  = \new_[30748]_  & \new_[30743]_ ;
  assign \new_[30753]_  = A234 & A232;
  assign \new_[30754]_  = ~A202 & \new_[30753]_ ;
  assign \new_[30758]_  = A269 & ~A266;
  assign \new_[30759]_  = A265 & \new_[30758]_ ;
  assign \new_[30760]_  = \new_[30759]_  & \new_[30754]_ ;
  assign \new_[30764]_  = A166 & ~A167;
  assign \new_[30765]_  = A170 & \new_[30764]_ ;
  assign \new_[30769]_  = ~A201 & A200;
  assign \new_[30770]_  = A199 & \new_[30769]_ ;
  assign \new_[30771]_  = \new_[30770]_  & \new_[30765]_ ;
  assign \new_[30775]_  = A234 & A233;
  assign \new_[30776]_  = ~A202 & \new_[30775]_ ;
  assign \new_[30780]_  = A302 & ~A299;
  assign \new_[30781]_  = A298 & \new_[30780]_ ;
  assign \new_[30782]_  = \new_[30781]_  & \new_[30776]_ ;
  assign \new_[30786]_  = A166 & ~A167;
  assign \new_[30787]_  = A170 & \new_[30786]_ ;
  assign \new_[30791]_  = ~A201 & A200;
  assign \new_[30792]_  = A199 & \new_[30791]_ ;
  assign \new_[30793]_  = \new_[30792]_  & \new_[30787]_ ;
  assign \new_[30797]_  = A234 & A233;
  assign \new_[30798]_  = ~A202 & \new_[30797]_ ;
  assign \new_[30802]_  = A302 & A299;
  assign \new_[30803]_  = ~A298 & \new_[30802]_ ;
  assign \new_[30804]_  = \new_[30803]_  & \new_[30798]_ ;
  assign \new_[30808]_  = A166 & ~A167;
  assign \new_[30809]_  = A170 & \new_[30808]_ ;
  assign \new_[30813]_  = ~A201 & A200;
  assign \new_[30814]_  = A199 & \new_[30813]_ ;
  assign \new_[30815]_  = \new_[30814]_  & \new_[30809]_ ;
  assign \new_[30819]_  = A234 & A233;
  assign \new_[30820]_  = ~A202 & \new_[30819]_ ;
  assign \new_[30824]_  = A269 & A266;
  assign \new_[30825]_  = ~A265 & \new_[30824]_ ;
  assign \new_[30826]_  = \new_[30825]_  & \new_[30820]_ ;
  assign \new_[30830]_  = A166 & ~A167;
  assign \new_[30831]_  = A170 & \new_[30830]_ ;
  assign \new_[30835]_  = ~A201 & A200;
  assign \new_[30836]_  = A199 & \new_[30835]_ ;
  assign \new_[30837]_  = \new_[30836]_  & \new_[30831]_ ;
  assign \new_[30841]_  = A234 & A233;
  assign \new_[30842]_  = ~A202 & \new_[30841]_ ;
  assign \new_[30846]_  = A269 & ~A266;
  assign \new_[30847]_  = A265 & \new_[30846]_ ;
  assign \new_[30848]_  = \new_[30847]_  & \new_[30842]_ ;
  assign \new_[30852]_  = A166 & ~A167;
  assign \new_[30853]_  = A170 & \new_[30852]_ ;
  assign \new_[30857]_  = ~A201 & A200;
  assign \new_[30858]_  = A199 & \new_[30857]_ ;
  assign \new_[30859]_  = \new_[30858]_  & \new_[30853]_ ;
  assign \new_[30863]_  = A233 & ~A232;
  assign \new_[30864]_  = ~A202 & \new_[30863]_ ;
  assign \new_[30868]_  = A300 & A299;
  assign \new_[30869]_  = A236 & \new_[30868]_ ;
  assign \new_[30870]_  = \new_[30869]_  & \new_[30864]_ ;
  assign \new_[30874]_  = A166 & ~A167;
  assign \new_[30875]_  = A170 & \new_[30874]_ ;
  assign \new_[30879]_  = ~A201 & A200;
  assign \new_[30880]_  = A199 & \new_[30879]_ ;
  assign \new_[30881]_  = \new_[30880]_  & \new_[30875]_ ;
  assign \new_[30885]_  = A233 & ~A232;
  assign \new_[30886]_  = ~A202 & \new_[30885]_ ;
  assign \new_[30890]_  = A300 & A298;
  assign \new_[30891]_  = A236 & \new_[30890]_ ;
  assign \new_[30892]_  = \new_[30891]_  & \new_[30886]_ ;
  assign \new_[30896]_  = A166 & ~A167;
  assign \new_[30897]_  = A170 & \new_[30896]_ ;
  assign \new_[30901]_  = ~A201 & A200;
  assign \new_[30902]_  = A199 & \new_[30901]_ ;
  assign \new_[30903]_  = \new_[30902]_  & \new_[30897]_ ;
  assign \new_[30907]_  = A233 & ~A232;
  assign \new_[30908]_  = ~A202 & \new_[30907]_ ;
  assign \new_[30912]_  = A267 & A265;
  assign \new_[30913]_  = A236 & \new_[30912]_ ;
  assign \new_[30914]_  = \new_[30913]_  & \new_[30908]_ ;
  assign \new_[30918]_  = A166 & ~A167;
  assign \new_[30919]_  = A170 & \new_[30918]_ ;
  assign \new_[30923]_  = ~A201 & A200;
  assign \new_[30924]_  = A199 & \new_[30923]_ ;
  assign \new_[30925]_  = \new_[30924]_  & \new_[30919]_ ;
  assign \new_[30929]_  = A233 & ~A232;
  assign \new_[30930]_  = ~A202 & \new_[30929]_ ;
  assign \new_[30934]_  = A267 & A266;
  assign \new_[30935]_  = A236 & \new_[30934]_ ;
  assign \new_[30936]_  = \new_[30935]_  & \new_[30930]_ ;
  assign \new_[30940]_  = A166 & ~A167;
  assign \new_[30941]_  = A170 & \new_[30940]_ ;
  assign \new_[30945]_  = ~A201 & A200;
  assign \new_[30946]_  = A199 & \new_[30945]_ ;
  assign \new_[30947]_  = \new_[30946]_  & \new_[30941]_ ;
  assign \new_[30951]_  = ~A233 & A232;
  assign \new_[30952]_  = ~A202 & \new_[30951]_ ;
  assign \new_[30956]_  = A300 & A299;
  assign \new_[30957]_  = A236 & \new_[30956]_ ;
  assign \new_[30958]_  = \new_[30957]_  & \new_[30952]_ ;
  assign \new_[30962]_  = A166 & ~A167;
  assign \new_[30963]_  = A170 & \new_[30962]_ ;
  assign \new_[30967]_  = ~A201 & A200;
  assign \new_[30968]_  = A199 & \new_[30967]_ ;
  assign \new_[30969]_  = \new_[30968]_  & \new_[30963]_ ;
  assign \new_[30973]_  = ~A233 & A232;
  assign \new_[30974]_  = ~A202 & \new_[30973]_ ;
  assign \new_[30978]_  = A300 & A298;
  assign \new_[30979]_  = A236 & \new_[30978]_ ;
  assign \new_[30980]_  = \new_[30979]_  & \new_[30974]_ ;
  assign \new_[30984]_  = A166 & ~A167;
  assign \new_[30985]_  = A170 & \new_[30984]_ ;
  assign \new_[30989]_  = ~A201 & A200;
  assign \new_[30990]_  = A199 & \new_[30989]_ ;
  assign \new_[30991]_  = \new_[30990]_  & \new_[30985]_ ;
  assign \new_[30995]_  = ~A233 & A232;
  assign \new_[30996]_  = ~A202 & \new_[30995]_ ;
  assign \new_[31000]_  = A267 & A265;
  assign \new_[31001]_  = A236 & \new_[31000]_ ;
  assign \new_[31002]_  = \new_[31001]_  & \new_[30996]_ ;
  assign \new_[31006]_  = A166 & ~A167;
  assign \new_[31007]_  = A170 & \new_[31006]_ ;
  assign \new_[31011]_  = ~A201 & A200;
  assign \new_[31012]_  = A199 & \new_[31011]_ ;
  assign \new_[31013]_  = \new_[31012]_  & \new_[31007]_ ;
  assign \new_[31017]_  = ~A233 & A232;
  assign \new_[31018]_  = ~A202 & \new_[31017]_ ;
  assign \new_[31022]_  = A267 & A266;
  assign \new_[31023]_  = A236 & \new_[31022]_ ;
  assign \new_[31024]_  = \new_[31023]_  & \new_[31018]_ ;
  assign \new_[31028]_  = A166 & ~A167;
  assign \new_[31029]_  = A170 & \new_[31028]_ ;
  assign \new_[31033]_  = ~A202 & ~A200;
  assign \new_[31034]_  = ~A199 & \new_[31033]_ ;
  assign \new_[31035]_  = \new_[31034]_  & \new_[31029]_ ;
  assign \new_[31039]_  = A236 & A233;
  assign \new_[31040]_  = ~A232 & \new_[31039]_ ;
  assign \new_[31044]_  = A302 & ~A299;
  assign \new_[31045]_  = A298 & \new_[31044]_ ;
  assign \new_[31046]_  = \new_[31045]_  & \new_[31040]_ ;
  assign \new_[31050]_  = A166 & ~A167;
  assign \new_[31051]_  = A170 & \new_[31050]_ ;
  assign \new_[31055]_  = ~A202 & ~A200;
  assign \new_[31056]_  = ~A199 & \new_[31055]_ ;
  assign \new_[31057]_  = \new_[31056]_  & \new_[31051]_ ;
  assign \new_[31061]_  = A236 & A233;
  assign \new_[31062]_  = ~A232 & \new_[31061]_ ;
  assign \new_[31066]_  = A302 & A299;
  assign \new_[31067]_  = ~A298 & \new_[31066]_ ;
  assign \new_[31068]_  = \new_[31067]_  & \new_[31062]_ ;
  assign \new_[31072]_  = A166 & ~A167;
  assign \new_[31073]_  = A170 & \new_[31072]_ ;
  assign \new_[31077]_  = ~A202 & ~A200;
  assign \new_[31078]_  = ~A199 & \new_[31077]_ ;
  assign \new_[31079]_  = \new_[31078]_  & \new_[31073]_ ;
  assign \new_[31083]_  = A236 & A233;
  assign \new_[31084]_  = ~A232 & \new_[31083]_ ;
  assign \new_[31088]_  = A269 & A266;
  assign \new_[31089]_  = ~A265 & \new_[31088]_ ;
  assign \new_[31090]_  = \new_[31089]_  & \new_[31084]_ ;
  assign \new_[31094]_  = A166 & ~A167;
  assign \new_[31095]_  = A170 & \new_[31094]_ ;
  assign \new_[31099]_  = ~A202 & ~A200;
  assign \new_[31100]_  = ~A199 & \new_[31099]_ ;
  assign \new_[31101]_  = \new_[31100]_  & \new_[31095]_ ;
  assign \new_[31105]_  = A236 & A233;
  assign \new_[31106]_  = ~A232 & \new_[31105]_ ;
  assign \new_[31110]_  = A269 & ~A266;
  assign \new_[31111]_  = A265 & \new_[31110]_ ;
  assign \new_[31112]_  = \new_[31111]_  & \new_[31106]_ ;
  assign \new_[31116]_  = A166 & ~A167;
  assign \new_[31117]_  = A170 & \new_[31116]_ ;
  assign \new_[31121]_  = ~A202 & ~A200;
  assign \new_[31122]_  = ~A199 & \new_[31121]_ ;
  assign \new_[31123]_  = \new_[31122]_  & \new_[31117]_ ;
  assign \new_[31127]_  = A236 & ~A233;
  assign \new_[31128]_  = A232 & \new_[31127]_ ;
  assign \new_[31132]_  = A302 & ~A299;
  assign \new_[31133]_  = A298 & \new_[31132]_ ;
  assign \new_[31134]_  = \new_[31133]_  & \new_[31128]_ ;
  assign \new_[31138]_  = A166 & ~A167;
  assign \new_[31139]_  = A170 & \new_[31138]_ ;
  assign \new_[31143]_  = ~A202 & ~A200;
  assign \new_[31144]_  = ~A199 & \new_[31143]_ ;
  assign \new_[31145]_  = \new_[31144]_  & \new_[31139]_ ;
  assign \new_[31149]_  = A236 & ~A233;
  assign \new_[31150]_  = A232 & \new_[31149]_ ;
  assign \new_[31154]_  = A302 & A299;
  assign \new_[31155]_  = ~A298 & \new_[31154]_ ;
  assign \new_[31156]_  = \new_[31155]_  & \new_[31150]_ ;
  assign \new_[31160]_  = A166 & ~A167;
  assign \new_[31161]_  = A170 & \new_[31160]_ ;
  assign \new_[31165]_  = ~A202 & ~A200;
  assign \new_[31166]_  = ~A199 & \new_[31165]_ ;
  assign \new_[31167]_  = \new_[31166]_  & \new_[31161]_ ;
  assign \new_[31171]_  = A236 & ~A233;
  assign \new_[31172]_  = A232 & \new_[31171]_ ;
  assign \new_[31176]_  = A269 & A266;
  assign \new_[31177]_  = ~A265 & \new_[31176]_ ;
  assign \new_[31178]_  = \new_[31177]_  & \new_[31172]_ ;
  assign \new_[31182]_  = A166 & ~A167;
  assign \new_[31183]_  = A170 & \new_[31182]_ ;
  assign \new_[31187]_  = ~A202 & ~A200;
  assign \new_[31188]_  = ~A199 & \new_[31187]_ ;
  assign \new_[31189]_  = \new_[31188]_  & \new_[31183]_ ;
  assign \new_[31193]_  = A236 & ~A233;
  assign \new_[31194]_  = A232 & \new_[31193]_ ;
  assign \new_[31198]_  = A269 & ~A266;
  assign \new_[31199]_  = A265 & \new_[31198]_ ;
  assign \new_[31200]_  = \new_[31199]_  & \new_[31194]_ ;
  assign \new_[31204]_  = ~A166 & ~A167;
  assign \new_[31205]_  = ~A169 & \new_[31204]_ ;
  assign \new_[31209]_  = A203 & A200;
  assign \new_[31210]_  = ~A199 & \new_[31209]_ ;
  assign \new_[31211]_  = \new_[31210]_  & \new_[31205]_ ;
  assign \new_[31215]_  = A236 & A233;
  assign \new_[31216]_  = ~A232 & \new_[31215]_ ;
  assign \new_[31220]_  = A302 & ~A299;
  assign \new_[31221]_  = A298 & \new_[31220]_ ;
  assign \new_[31222]_  = \new_[31221]_  & \new_[31216]_ ;
  assign \new_[31226]_  = ~A166 & ~A167;
  assign \new_[31227]_  = ~A169 & \new_[31226]_ ;
  assign \new_[31231]_  = A203 & A200;
  assign \new_[31232]_  = ~A199 & \new_[31231]_ ;
  assign \new_[31233]_  = \new_[31232]_  & \new_[31227]_ ;
  assign \new_[31237]_  = A236 & A233;
  assign \new_[31238]_  = ~A232 & \new_[31237]_ ;
  assign \new_[31242]_  = A302 & A299;
  assign \new_[31243]_  = ~A298 & \new_[31242]_ ;
  assign \new_[31244]_  = \new_[31243]_  & \new_[31238]_ ;
  assign \new_[31248]_  = ~A166 & ~A167;
  assign \new_[31249]_  = ~A169 & \new_[31248]_ ;
  assign \new_[31253]_  = A203 & A200;
  assign \new_[31254]_  = ~A199 & \new_[31253]_ ;
  assign \new_[31255]_  = \new_[31254]_  & \new_[31249]_ ;
  assign \new_[31259]_  = A236 & A233;
  assign \new_[31260]_  = ~A232 & \new_[31259]_ ;
  assign \new_[31264]_  = A269 & A266;
  assign \new_[31265]_  = ~A265 & \new_[31264]_ ;
  assign \new_[31266]_  = \new_[31265]_  & \new_[31260]_ ;
  assign \new_[31270]_  = ~A166 & ~A167;
  assign \new_[31271]_  = ~A169 & \new_[31270]_ ;
  assign \new_[31275]_  = A203 & A200;
  assign \new_[31276]_  = ~A199 & \new_[31275]_ ;
  assign \new_[31277]_  = \new_[31276]_  & \new_[31271]_ ;
  assign \new_[31281]_  = A236 & A233;
  assign \new_[31282]_  = ~A232 & \new_[31281]_ ;
  assign \new_[31286]_  = A269 & ~A266;
  assign \new_[31287]_  = A265 & \new_[31286]_ ;
  assign \new_[31288]_  = \new_[31287]_  & \new_[31282]_ ;
  assign \new_[31292]_  = ~A166 & ~A167;
  assign \new_[31293]_  = ~A169 & \new_[31292]_ ;
  assign \new_[31297]_  = A203 & A200;
  assign \new_[31298]_  = ~A199 & \new_[31297]_ ;
  assign \new_[31299]_  = \new_[31298]_  & \new_[31293]_ ;
  assign \new_[31303]_  = A236 & ~A233;
  assign \new_[31304]_  = A232 & \new_[31303]_ ;
  assign \new_[31308]_  = A302 & ~A299;
  assign \new_[31309]_  = A298 & \new_[31308]_ ;
  assign \new_[31310]_  = \new_[31309]_  & \new_[31304]_ ;
  assign \new_[31314]_  = ~A166 & ~A167;
  assign \new_[31315]_  = ~A169 & \new_[31314]_ ;
  assign \new_[31319]_  = A203 & A200;
  assign \new_[31320]_  = ~A199 & \new_[31319]_ ;
  assign \new_[31321]_  = \new_[31320]_  & \new_[31315]_ ;
  assign \new_[31325]_  = A236 & ~A233;
  assign \new_[31326]_  = A232 & \new_[31325]_ ;
  assign \new_[31330]_  = A302 & A299;
  assign \new_[31331]_  = ~A298 & \new_[31330]_ ;
  assign \new_[31332]_  = \new_[31331]_  & \new_[31326]_ ;
  assign \new_[31336]_  = ~A166 & ~A167;
  assign \new_[31337]_  = ~A169 & \new_[31336]_ ;
  assign \new_[31341]_  = A203 & A200;
  assign \new_[31342]_  = ~A199 & \new_[31341]_ ;
  assign \new_[31343]_  = \new_[31342]_  & \new_[31337]_ ;
  assign \new_[31347]_  = A236 & ~A233;
  assign \new_[31348]_  = A232 & \new_[31347]_ ;
  assign \new_[31352]_  = A269 & A266;
  assign \new_[31353]_  = ~A265 & \new_[31352]_ ;
  assign \new_[31354]_  = \new_[31353]_  & \new_[31348]_ ;
  assign \new_[31358]_  = ~A166 & ~A167;
  assign \new_[31359]_  = ~A169 & \new_[31358]_ ;
  assign \new_[31363]_  = A203 & A200;
  assign \new_[31364]_  = ~A199 & \new_[31363]_ ;
  assign \new_[31365]_  = \new_[31364]_  & \new_[31359]_ ;
  assign \new_[31369]_  = A236 & ~A233;
  assign \new_[31370]_  = A232 & \new_[31369]_ ;
  assign \new_[31374]_  = A269 & ~A266;
  assign \new_[31375]_  = A265 & \new_[31374]_ ;
  assign \new_[31376]_  = \new_[31375]_  & \new_[31370]_ ;
  assign \new_[31380]_  = ~A166 & ~A167;
  assign \new_[31381]_  = ~A169 & \new_[31380]_ ;
  assign \new_[31385]_  = A203 & ~A200;
  assign \new_[31386]_  = A199 & \new_[31385]_ ;
  assign \new_[31387]_  = \new_[31386]_  & \new_[31381]_ ;
  assign \new_[31391]_  = A236 & A233;
  assign \new_[31392]_  = ~A232 & \new_[31391]_ ;
  assign \new_[31396]_  = A302 & ~A299;
  assign \new_[31397]_  = A298 & \new_[31396]_ ;
  assign \new_[31398]_  = \new_[31397]_  & \new_[31392]_ ;
  assign \new_[31402]_  = ~A166 & ~A167;
  assign \new_[31403]_  = ~A169 & \new_[31402]_ ;
  assign \new_[31407]_  = A203 & ~A200;
  assign \new_[31408]_  = A199 & \new_[31407]_ ;
  assign \new_[31409]_  = \new_[31408]_  & \new_[31403]_ ;
  assign \new_[31413]_  = A236 & A233;
  assign \new_[31414]_  = ~A232 & \new_[31413]_ ;
  assign \new_[31418]_  = A302 & A299;
  assign \new_[31419]_  = ~A298 & \new_[31418]_ ;
  assign \new_[31420]_  = \new_[31419]_  & \new_[31414]_ ;
  assign \new_[31424]_  = ~A166 & ~A167;
  assign \new_[31425]_  = ~A169 & \new_[31424]_ ;
  assign \new_[31429]_  = A203 & ~A200;
  assign \new_[31430]_  = A199 & \new_[31429]_ ;
  assign \new_[31431]_  = \new_[31430]_  & \new_[31425]_ ;
  assign \new_[31435]_  = A236 & A233;
  assign \new_[31436]_  = ~A232 & \new_[31435]_ ;
  assign \new_[31440]_  = A269 & A266;
  assign \new_[31441]_  = ~A265 & \new_[31440]_ ;
  assign \new_[31442]_  = \new_[31441]_  & \new_[31436]_ ;
  assign \new_[31446]_  = ~A166 & ~A167;
  assign \new_[31447]_  = ~A169 & \new_[31446]_ ;
  assign \new_[31451]_  = A203 & ~A200;
  assign \new_[31452]_  = A199 & \new_[31451]_ ;
  assign \new_[31453]_  = \new_[31452]_  & \new_[31447]_ ;
  assign \new_[31457]_  = A236 & A233;
  assign \new_[31458]_  = ~A232 & \new_[31457]_ ;
  assign \new_[31462]_  = A269 & ~A266;
  assign \new_[31463]_  = A265 & \new_[31462]_ ;
  assign \new_[31464]_  = \new_[31463]_  & \new_[31458]_ ;
  assign \new_[31468]_  = ~A166 & ~A167;
  assign \new_[31469]_  = ~A169 & \new_[31468]_ ;
  assign \new_[31473]_  = A203 & ~A200;
  assign \new_[31474]_  = A199 & \new_[31473]_ ;
  assign \new_[31475]_  = \new_[31474]_  & \new_[31469]_ ;
  assign \new_[31479]_  = A236 & ~A233;
  assign \new_[31480]_  = A232 & \new_[31479]_ ;
  assign \new_[31484]_  = A302 & ~A299;
  assign \new_[31485]_  = A298 & \new_[31484]_ ;
  assign \new_[31486]_  = \new_[31485]_  & \new_[31480]_ ;
  assign \new_[31490]_  = ~A166 & ~A167;
  assign \new_[31491]_  = ~A169 & \new_[31490]_ ;
  assign \new_[31495]_  = A203 & ~A200;
  assign \new_[31496]_  = A199 & \new_[31495]_ ;
  assign \new_[31497]_  = \new_[31496]_  & \new_[31491]_ ;
  assign \new_[31501]_  = A236 & ~A233;
  assign \new_[31502]_  = A232 & \new_[31501]_ ;
  assign \new_[31506]_  = A302 & A299;
  assign \new_[31507]_  = ~A298 & \new_[31506]_ ;
  assign \new_[31508]_  = \new_[31507]_  & \new_[31502]_ ;
  assign \new_[31512]_  = ~A166 & ~A167;
  assign \new_[31513]_  = ~A169 & \new_[31512]_ ;
  assign \new_[31517]_  = A203 & ~A200;
  assign \new_[31518]_  = A199 & \new_[31517]_ ;
  assign \new_[31519]_  = \new_[31518]_  & \new_[31513]_ ;
  assign \new_[31523]_  = A236 & ~A233;
  assign \new_[31524]_  = A232 & \new_[31523]_ ;
  assign \new_[31528]_  = A269 & A266;
  assign \new_[31529]_  = ~A265 & \new_[31528]_ ;
  assign \new_[31530]_  = \new_[31529]_  & \new_[31524]_ ;
  assign \new_[31534]_  = ~A166 & ~A167;
  assign \new_[31535]_  = ~A169 & \new_[31534]_ ;
  assign \new_[31539]_  = A203 & ~A200;
  assign \new_[31540]_  = A199 & \new_[31539]_ ;
  assign \new_[31541]_  = \new_[31540]_  & \new_[31535]_ ;
  assign \new_[31545]_  = A236 & ~A233;
  assign \new_[31546]_  = A232 & \new_[31545]_ ;
  assign \new_[31550]_  = A269 & ~A266;
  assign \new_[31551]_  = A265 & \new_[31550]_ ;
  assign \new_[31552]_  = \new_[31551]_  & \new_[31546]_ ;
  assign \new_[31556]_  = A167 & ~A168;
  assign \new_[31557]_  = ~A169 & \new_[31556]_ ;
  assign \new_[31561]_  = A201 & A199;
  assign \new_[31562]_  = A166 & \new_[31561]_ ;
  assign \new_[31563]_  = \new_[31562]_  & \new_[31557]_ ;
  assign \new_[31567]_  = A236 & A233;
  assign \new_[31568]_  = ~A232 & \new_[31567]_ ;
  assign \new_[31572]_  = A302 & ~A299;
  assign \new_[31573]_  = A298 & \new_[31572]_ ;
  assign \new_[31574]_  = \new_[31573]_  & \new_[31568]_ ;
  assign \new_[31578]_  = A167 & ~A168;
  assign \new_[31579]_  = ~A169 & \new_[31578]_ ;
  assign \new_[31583]_  = A201 & A199;
  assign \new_[31584]_  = A166 & \new_[31583]_ ;
  assign \new_[31585]_  = \new_[31584]_  & \new_[31579]_ ;
  assign \new_[31589]_  = A236 & A233;
  assign \new_[31590]_  = ~A232 & \new_[31589]_ ;
  assign \new_[31594]_  = A302 & A299;
  assign \new_[31595]_  = ~A298 & \new_[31594]_ ;
  assign \new_[31596]_  = \new_[31595]_  & \new_[31590]_ ;
  assign \new_[31600]_  = A167 & ~A168;
  assign \new_[31601]_  = ~A169 & \new_[31600]_ ;
  assign \new_[31605]_  = A201 & A199;
  assign \new_[31606]_  = A166 & \new_[31605]_ ;
  assign \new_[31607]_  = \new_[31606]_  & \new_[31601]_ ;
  assign \new_[31611]_  = A236 & A233;
  assign \new_[31612]_  = ~A232 & \new_[31611]_ ;
  assign \new_[31616]_  = A269 & A266;
  assign \new_[31617]_  = ~A265 & \new_[31616]_ ;
  assign \new_[31618]_  = \new_[31617]_  & \new_[31612]_ ;
  assign \new_[31622]_  = A167 & ~A168;
  assign \new_[31623]_  = ~A169 & \new_[31622]_ ;
  assign \new_[31627]_  = A201 & A199;
  assign \new_[31628]_  = A166 & \new_[31627]_ ;
  assign \new_[31629]_  = \new_[31628]_  & \new_[31623]_ ;
  assign \new_[31633]_  = A236 & A233;
  assign \new_[31634]_  = ~A232 & \new_[31633]_ ;
  assign \new_[31638]_  = A269 & ~A266;
  assign \new_[31639]_  = A265 & \new_[31638]_ ;
  assign \new_[31640]_  = \new_[31639]_  & \new_[31634]_ ;
  assign \new_[31644]_  = A167 & ~A168;
  assign \new_[31645]_  = ~A169 & \new_[31644]_ ;
  assign \new_[31649]_  = A201 & A199;
  assign \new_[31650]_  = A166 & \new_[31649]_ ;
  assign \new_[31651]_  = \new_[31650]_  & \new_[31645]_ ;
  assign \new_[31655]_  = A236 & ~A233;
  assign \new_[31656]_  = A232 & \new_[31655]_ ;
  assign \new_[31660]_  = A302 & ~A299;
  assign \new_[31661]_  = A298 & \new_[31660]_ ;
  assign \new_[31662]_  = \new_[31661]_  & \new_[31656]_ ;
  assign \new_[31666]_  = A167 & ~A168;
  assign \new_[31667]_  = ~A169 & \new_[31666]_ ;
  assign \new_[31671]_  = A201 & A199;
  assign \new_[31672]_  = A166 & \new_[31671]_ ;
  assign \new_[31673]_  = \new_[31672]_  & \new_[31667]_ ;
  assign \new_[31677]_  = A236 & ~A233;
  assign \new_[31678]_  = A232 & \new_[31677]_ ;
  assign \new_[31682]_  = A302 & A299;
  assign \new_[31683]_  = ~A298 & \new_[31682]_ ;
  assign \new_[31684]_  = \new_[31683]_  & \new_[31678]_ ;
  assign \new_[31688]_  = A167 & ~A168;
  assign \new_[31689]_  = ~A169 & \new_[31688]_ ;
  assign \new_[31693]_  = A201 & A199;
  assign \new_[31694]_  = A166 & \new_[31693]_ ;
  assign \new_[31695]_  = \new_[31694]_  & \new_[31689]_ ;
  assign \new_[31699]_  = A236 & ~A233;
  assign \new_[31700]_  = A232 & \new_[31699]_ ;
  assign \new_[31704]_  = A269 & A266;
  assign \new_[31705]_  = ~A265 & \new_[31704]_ ;
  assign \new_[31706]_  = \new_[31705]_  & \new_[31700]_ ;
  assign \new_[31710]_  = A167 & ~A168;
  assign \new_[31711]_  = ~A169 & \new_[31710]_ ;
  assign \new_[31715]_  = A201 & A199;
  assign \new_[31716]_  = A166 & \new_[31715]_ ;
  assign \new_[31717]_  = \new_[31716]_  & \new_[31711]_ ;
  assign \new_[31721]_  = A236 & ~A233;
  assign \new_[31722]_  = A232 & \new_[31721]_ ;
  assign \new_[31726]_  = A269 & ~A266;
  assign \new_[31727]_  = A265 & \new_[31726]_ ;
  assign \new_[31728]_  = \new_[31727]_  & \new_[31722]_ ;
  assign \new_[31732]_  = A167 & ~A168;
  assign \new_[31733]_  = ~A169 & \new_[31732]_ ;
  assign \new_[31737]_  = A201 & A200;
  assign \new_[31738]_  = A166 & \new_[31737]_ ;
  assign \new_[31739]_  = \new_[31738]_  & \new_[31733]_ ;
  assign \new_[31743]_  = A236 & A233;
  assign \new_[31744]_  = ~A232 & \new_[31743]_ ;
  assign \new_[31748]_  = A302 & ~A299;
  assign \new_[31749]_  = A298 & \new_[31748]_ ;
  assign \new_[31750]_  = \new_[31749]_  & \new_[31744]_ ;
  assign \new_[31754]_  = A167 & ~A168;
  assign \new_[31755]_  = ~A169 & \new_[31754]_ ;
  assign \new_[31759]_  = A201 & A200;
  assign \new_[31760]_  = A166 & \new_[31759]_ ;
  assign \new_[31761]_  = \new_[31760]_  & \new_[31755]_ ;
  assign \new_[31765]_  = A236 & A233;
  assign \new_[31766]_  = ~A232 & \new_[31765]_ ;
  assign \new_[31770]_  = A302 & A299;
  assign \new_[31771]_  = ~A298 & \new_[31770]_ ;
  assign \new_[31772]_  = \new_[31771]_  & \new_[31766]_ ;
  assign \new_[31776]_  = A167 & ~A168;
  assign \new_[31777]_  = ~A169 & \new_[31776]_ ;
  assign \new_[31781]_  = A201 & A200;
  assign \new_[31782]_  = A166 & \new_[31781]_ ;
  assign \new_[31783]_  = \new_[31782]_  & \new_[31777]_ ;
  assign \new_[31787]_  = A236 & A233;
  assign \new_[31788]_  = ~A232 & \new_[31787]_ ;
  assign \new_[31792]_  = A269 & A266;
  assign \new_[31793]_  = ~A265 & \new_[31792]_ ;
  assign \new_[31794]_  = \new_[31793]_  & \new_[31788]_ ;
  assign \new_[31798]_  = A167 & ~A168;
  assign \new_[31799]_  = ~A169 & \new_[31798]_ ;
  assign \new_[31803]_  = A201 & A200;
  assign \new_[31804]_  = A166 & \new_[31803]_ ;
  assign \new_[31805]_  = \new_[31804]_  & \new_[31799]_ ;
  assign \new_[31809]_  = A236 & A233;
  assign \new_[31810]_  = ~A232 & \new_[31809]_ ;
  assign \new_[31814]_  = A269 & ~A266;
  assign \new_[31815]_  = A265 & \new_[31814]_ ;
  assign \new_[31816]_  = \new_[31815]_  & \new_[31810]_ ;
  assign \new_[31820]_  = A167 & ~A168;
  assign \new_[31821]_  = ~A169 & \new_[31820]_ ;
  assign \new_[31825]_  = A201 & A200;
  assign \new_[31826]_  = A166 & \new_[31825]_ ;
  assign \new_[31827]_  = \new_[31826]_  & \new_[31821]_ ;
  assign \new_[31831]_  = A236 & ~A233;
  assign \new_[31832]_  = A232 & \new_[31831]_ ;
  assign \new_[31836]_  = A302 & ~A299;
  assign \new_[31837]_  = A298 & \new_[31836]_ ;
  assign \new_[31838]_  = \new_[31837]_  & \new_[31832]_ ;
  assign \new_[31842]_  = A167 & ~A168;
  assign \new_[31843]_  = ~A169 & \new_[31842]_ ;
  assign \new_[31847]_  = A201 & A200;
  assign \new_[31848]_  = A166 & \new_[31847]_ ;
  assign \new_[31849]_  = \new_[31848]_  & \new_[31843]_ ;
  assign \new_[31853]_  = A236 & ~A233;
  assign \new_[31854]_  = A232 & \new_[31853]_ ;
  assign \new_[31858]_  = A302 & A299;
  assign \new_[31859]_  = ~A298 & \new_[31858]_ ;
  assign \new_[31860]_  = \new_[31859]_  & \new_[31854]_ ;
  assign \new_[31864]_  = A167 & ~A168;
  assign \new_[31865]_  = ~A169 & \new_[31864]_ ;
  assign \new_[31869]_  = A201 & A200;
  assign \new_[31870]_  = A166 & \new_[31869]_ ;
  assign \new_[31871]_  = \new_[31870]_  & \new_[31865]_ ;
  assign \new_[31875]_  = A236 & ~A233;
  assign \new_[31876]_  = A232 & \new_[31875]_ ;
  assign \new_[31880]_  = A269 & A266;
  assign \new_[31881]_  = ~A265 & \new_[31880]_ ;
  assign \new_[31882]_  = \new_[31881]_  & \new_[31876]_ ;
  assign \new_[31886]_  = A167 & ~A168;
  assign \new_[31887]_  = ~A169 & \new_[31886]_ ;
  assign \new_[31891]_  = A201 & A200;
  assign \new_[31892]_  = A166 & \new_[31891]_ ;
  assign \new_[31893]_  = \new_[31892]_  & \new_[31887]_ ;
  assign \new_[31897]_  = A236 & ~A233;
  assign \new_[31898]_  = A232 & \new_[31897]_ ;
  assign \new_[31902]_  = A269 & ~A266;
  assign \new_[31903]_  = A265 & \new_[31902]_ ;
  assign \new_[31904]_  = \new_[31903]_  & \new_[31898]_ ;
  assign \new_[31908]_  = A167 & ~A168;
  assign \new_[31909]_  = ~A169 & \new_[31908]_ ;
  assign \new_[31913]_  = A200 & ~A199;
  assign \new_[31914]_  = A166 & \new_[31913]_ ;
  assign \new_[31915]_  = \new_[31914]_  & \new_[31909]_ ;
  assign \new_[31919]_  = A234 & A232;
  assign \new_[31920]_  = A203 & \new_[31919]_ ;
  assign \new_[31924]_  = A302 & ~A299;
  assign \new_[31925]_  = A298 & \new_[31924]_ ;
  assign \new_[31926]_  = \new_[31925]_  & \new_[31920]_ ;
  assign \new_[31930]_  = A167 & ~A168;
  assign \new_[31931]_  = ~A169 & \new_[31930]_ ;
  assign \new_[31935]_  = A200 & ~A199;
  assign \new_[31936]_  = A166 & \new_[31935]_ ;
  assign \new_[31937]_  = \new_[31936]_  & \new_[31931]_ ;
  assign \new_[31941]_  = A234 & A232;
  assign \new_[31942]_  = A203 & \new_[31941]_ ;
  assign \new_[31946]_  = A302 & A299;
  assign \new_[31947]_  = ~A298 & \new_[31946]_ ;
  assign \new_[31948]_  = \new_[31947]_  & \new_[31942]_ ;
  assign \new_[31952]_  = A167 & ~A168;
  assign \new_[31953]_  = ~A169 & \new_[31952]_ ;
  assign \new_[31957]_  = A200 & ~A199;
  assign \new_[31958]_  = A166 & \new_[31957]_ ;
  assign \new_[31959]_  = \new_[31958]_  & \new_[31953]_ ;
  assign \new_[31963]_  = A234 & A232;
  assign \new_[31964]_  = A203 & \new_[31963]_ ;
  assign \new_[31968]_  = A269 & A266;
  assign \new_[31969]_  = ~A265 & \new_[31968]_ ;
  assign \new_[31970]_  = \new_[31969]_  & \new_[31964]_ ;
  assign \new_[31974]_  = A167 & ~A168;
  assign \new_[31975]_  = ~A169 & \new_[31974]_ ;
  assign \new_[31979]_  = A200 & ~A199;
  assign \new_[31980]_  = A166 & \new_[31979]_ ;
  assign \new_[31981]_  = \new_[31980]_  & \new_[31975]_ ;
  assign \new_[31985]_  = A234 & A232;
  assign \new_[31986]_  = A203 & \new_[31985]_ ;
  assign \new_[31990]_  = A269 & ~A266;
  assign \new_[31991]_  = A265 & \new_[31990]_ ;
  assign \new_[31992]_  = \new_[31991]_  & \new_[31986]_ ;
  assign \new_[31996]_  = A167 & ~A168;
  assign \new_[31997]_  = ~A169 & \new_[31996]_ ;
  assign \new_[32001]_  = A200 & ~A199;
  assign \new_[32002]_  = A166 & \new_[32001]_ ;
  assign \new_[32003]_  = \new_[32002]_  & \new_[31997]_ ;
  assign \new_[32007]_  = A234 & A233;
  assign \new_[32008]_  = A203 & \new_[32007]_ ;
  assign \new_[32012]_  = A302 & ~A299;
  assign \new_[32013]_  = A298 & \new_[32012]_ ;
  assign \new_[32014]_  = \new_[32013]_  & \new_[32008]_ ;
  assign \new_[32018]_  = A167 & ~A168;
  assign \new_[32019]_  = ~A169 & \new_[32018]_ ;
  assign \new_[32023]_  = A200 & ~A199;
  assign \new_[32024]_  = A166 & \new_[32023]_ ;
  assign \new_[32025]_  = \new_[32024]_  & \new_[32019]_ ;
  assign \new_[32029]_  = A234 & A233;
  assign \new_[32030]_  = A203 & \new_[32029]_ ;
  assign \new_[32034]_  = A302 & A299;
  assign \new_[32035]_  = ~A298 & \new_[32034]_ ;
  assign \new_[32036]_  = \new_[32035]_  & \new_[32030]_ ;
  assign \new_[32040]_  = A167 & ~A168;
  assign \new_[32041]_  = ~A169 & \new_[32040]_ ;
  assign \new_[32045]_  = A200 & ~A199;
  assign \new_[32046]_  = A166 & \new_[32045]_ ;
  assign \new_[32047]_  = \new_[32046]_  & \new_[32041]_ ;
  assign \new_[32051]_  = A234 & A233;
  assign \new_[32052]_  = A203 & \new_[32051]_ ;
  assign \new_[32056]_  = A269 & A266;
  assign \new_[32057]_  = ~A265 & \new_[32056]_ ;
  assign \new_[32058]_  = \new_[32057]_  & \new_[32052]_ ;
  assign \new_[32062]_  = A167 & ~A168;
  assign \new_[32063]_  = ~A169 & \new_[32062]_ ;
  assign \new_[32067]_  = A200 & ~A199;
  assign \new_[32068]_  = A166 & \new_[32067]_ ;
  assign \new_[32069]_  = \new_[32068]_  & \new_[32063]_ ;
  assign \new_[32073]_  = A234 & A233;
  assign \new_[32074]_  = A203 & \new_[32073]_ ;
  assign \new_[32078]_  = A269 & ~A266;
  assign \new_[32079]_  = A265 & \new_[32078]_ ;
  assign \new_[32080]_  = \new_[32079]_  & \new_[32074]_ ;
  assign \new_[32084]_  = A167 & ~A168;
  assign \new_[32085]_  = ~A169 & \new_[32084]_ ;
  assign \new_[32089]_  = A200 & ~A199;
  assign \new_[32090]_  = A166 & \new_[32089]_ ;
  assign \new_[32091]_  = \new_[32090]_  & \new_[32085]_ ;
  assign \new_[32095]_  = A233 & ~A232;
  assign \new_[32096]_  = A203 & \new_[32095]_ ;
  assign \new_[32100]_  = A300 & A299;
  assign \new_[32101]_  = A236 & \new_[32100]_ ;
  assign \new_[32102]_  = \new_[32101]_  & \new_[32096]_ ;
  assign \new_[32106]_  = A167 & ~A168;
  assign \new_[32107]_  = ~A169 & \new_[32106]_ ;
  assign \new_[32111]_  = A200 & ~A199;
  assign \new_[32112]_  = A166 & \new_[32111]_ ;
  assign \new_[32113]_  = \new_[32112]_  & \new_[32107]_ ;
  assign \new_[32117]_  = A233 & ~A232;
  assign \new_[32118]_  = A203 & \new_[32117]_ ;
  assign \new_[32122]_  = A300 & A298;
  assign \new_[32123]_  = A236 & \new_[32122]_ ;
  assign \new_[32124]_  = \new_[32123]_  & \new_[32118]_ ;
  assign \new_[32128]_  = A167 & ~A168;
  assign \new_[32129]_  = ~A169 & \new_[32128]_ ;
  assign \new_[32133]_  = A200 & ~A199;
  assign \new_[32134]_  = A166 & \new_[32133]_ ;
  assign \new_[32135]_  = \new_[32134]_  & \new_[32129]_ ;
  assign \new_[32139]_  = A233 & ~A232;
  assign \new_[32140]_  = A203 & \new_[32139]_ ;
  assign \new_[32144]_  = A267 & A265;
  assign \new_[32145]_  = A236 & \new_[32144]_ ;
  assign \new_[32146]_  = \new_[32145]_  & \new_[32140]_ ;
  assign \new_[32150]_  = A167 & ~A168;
  assign \new_[32151]_  = ~A169 & \new_[32150]_ ;
  assign \new_[32155]_  = A200 & ~A199;
  assign \new_[32156]_  = A166 & \new_[32155]_ ;
  assign \new_[32157]_  = \new_[32156]_  & \new_[32151]_ ;
  assign \new_[32161]_  = A233 & ~A232;
  assign \new_[32162]_  = A203 & \new_[32161]_ ;
  assign \new_[32166]_  = A267 & A266;
  assign \new_[32167]_  = A236 & \new_[32166]_ ;
  assign \new_[32168]_  = \new_[32167]_  & \new_[32162]_ ;
  assign \new_[32172]_  = A167 & ~A168;
  assign \new_[32173]_  = ~A169 & \new_[32172]_ ;
  assign \new_[32177]_  = A200 & ~A199;
  assign \new_[32178]_  = A166 & \new_[32177]_ ;
  assign \new_[32179]_  = \new_[32178]_  & \new_[32173]_ ;
  assign \new_[32183]_  = ~A233 & A232;
  assign \new_[32184]_  = A203 & \new_[32183]_ ;
  assign \new_[32188]_  = A300 & A299;
  assign \new_[32189]_  = A236 & \new_[32188]_ ;
  assign \new_[32190]_  = \new_[32189]_  & \new_[32184]_ ;
  assign \new_[32194]_  = A167 & ~A168;
  assign \new_[32195]_  = ~A169 & \new_[32194]_ ;
  assign \new_[32199]_  = A200 & ~A199;
  assign \new_[32200]_  = A166 & \new_[32199]_ ;
  assign \new_[32201]_  = \new_[32200]_  & \new_[32195]_ ;
  assign \new_[32205]_  = ~A233 & A232;
  assign \new_[32206]_  = A203 & \new_[32205]_ ;
  assign \new_[32210]_  = A300 & A298;
  assign \new_[32211]_  = A236 & \new_[32210]_ ;
  assign \new_[32212]_  = \new_[32211]_  & \new_[32206]_ ;
  assign \new_[32216]_  = A167 & ~A168;
  assign \new_[32217]_  = ~A169 & \new_[32216]_ ;
  assign \new_[32221]_  = A200 & ~A199;
  assign \new_[32222]_  = A166 & \new_[32221]_ ;
  assign \new_[32223]_  = \new_[32222]_  & \new_[32217]_ ;
  assign \new_[32227]_  = ~A233 & A232;
  assign \new_[32228]_  = A203 & \new_[32227]_ ;
  assign \new_[32232]_  = A267 & A265;
  assign \new_[32233]_  = A236 & \new_[32232]_ ;
  assign \new_[32234]_  = \new_[32233]_  & \new_[32228]_ ;
  assign \new_[32238]_  = A167 & ~A168;
  assign \new_[32239]_  = ~A169 & \new_[32238]_ ;
  assign \new_[32243]_  = A200 & ~A199;
  assign \new_[32244]_  = A166 & \new_[32243]_ ;
  assign \new_[32245]_  = \new_[32244]_  & \new_[32239]_ ;
  assign \new_[32249]_  = ~A233 & A232;
  assign \new_[32250]_  = A203 & \new_[32249]_ ;
  assign \new_[32254]_  = A267 & A266;
  assign \new_[32255]_  = A236 & \new_[32254]_ ;
  assign \new_[32256]_  = \new_[32255]_  & \new_[32250]_ ;
  assign \new_[32260]_  = A167 & ~A168;
  assign \new_[32261]_  = ~A169 & \new_[32260]_ ;
  assign \new_[32265]_  = ~A200 & A199;
  assign \new_[32266]_  = A166 & \new_[32265]_ ;
  assign \new_[32267]_  = \new_[32266]_  & \new_[32261]_ ;
  assign \new_[32271]_  = A234 & A232;
  assign \new_[32272]_  = A203 & \new_[32271]_ ;
  assign \new_[32276]_  = A302 & ~A299;
  assign \new_[32277]_  = A298 & \new_[32276]_ ;
  assign \new_[32278]_  = \new_[32277]_  & \new_[32272]_ ;
  assign \new_[32282]_  = A167 & ~A168;
  assign \new_[32283]_  = ~A169 & \new_[32282]_ ;
  assign \new_[32287]_  = ~A200 & A199;
  assign \new_[32288]_  = A166 & \new_[32287]_ ;
  assign \new_[32289]_  = \new_[32288]_  & \new_[32283]_ ;
  assign \new_[32293]_  = A234 & A232;
  assign \new_[32294]_  = A203 & \new_[32293]_ ;
  assign \new_[32298]_  = A302 & A299;
  assign \new_[32299]_  = ~A298 & \new_[32298]_ ;
  assign \new_[32300]_  = \new_[32299]_  & \new_[32294]_ ;
  assign \new_[32304]_  = A167 & ~A168;
  assign \new_[32305]_  = ~A169 & \new_[32304]_ ;
  assign \new_[32309]_  = ~A200 & A199;
  assign \new_[32310]_  = A166 & \new_[32309]_ ;
  assign \new_[32311]_  = \new_[32310]_  & \new_[32305]_ ;
  assign \new_[32315]_  = A234 & A232;
  assign \new_[32316]_  = A203 & \new_[32315]_ ;
  assign \new_[32320]_  = A269 & A266;
  assign \new_[32321]_  = ~A265 & \new_[32320]_ ;
  assign \new_[32322]_  = \new_[32321]_  & \new_[32316]_ ;
  assign \new_[32326]_  = A167 & ~A168;
  assign \new_[32327]_  = ~A169 & \new_[32326]_ ;
  assign \new_[32331]_  = ~A200 & A199;
  assign \new_[32332]_  = A166 & \new_[32331]_ ;
  assign \new_[32333]_  = \new_[32332]_  & \new_[32327]_ ;
  assign \new_[32337]_  = A234 & A232;
  assign \new_[32338]_  = A203 & \new_[32337]_ ;
  assign \new_[32342]_  = A269 & ~A266;
  assign \new_[32343]_  = A265 & \new_[32342]_ ;
  assign \new_[32344]_  = \new_[32343]_  & \new_[32338]_ ;
  assign \new_[32348]_  = A167 & ~A168;
  assign \new_[32349]_  = ~A169 & \new_[32348]_ ;
  assign \new_[32353]_  = ~A200 & A199;
  assign \new_[32354]_  = A166 & \new_[32353]_ ;
  assign \new_[32355]_  = \new_[32354]_  & \new_[32349]_ ;
  assign \new_[32359]_  = A234 & A233;
  assign \new_[32360]_  = A203 & \new_[32359]_ ;
  assign \new_[32364]_  = A302 & ~A299;
  assign \new_[32365]_  = A298 & \new_[32364]_ ;
  assign \new_[32366]_  = \new_[32365]_  & \new_[32360]_ ;
  assign \new_[32370]_  = A167 & ~A168;
  assign \new_[32371]_  = ~A169 & \new_[32370]_ ;
  assign \new_[32375]_  = ~A200 & A199;
  assign \new_[32376]_  = A166 & \new_[32375]_ ;
  assign \new_[32377]_  = \new_[32376]_  & \new_[32371]_ ;
  assign \new_[32381]_  = A234 & A233;
  assign \new_[32382]_  = A203 & \new_[32381]_ ;
  assign \new_[32386]_  = A302 & A299;
  assign \new_[32387]_  = ~A298 & \new_[32386]_ ;
  assign \new_[32388]_  = \new_[32387]_  & \new_[32382]_ ;
  assign \new_[32392]_  = A167 & ~A168;
  assign \new_[32393]_  = ~A169 & \new_[32392]_ ;
  assign \new_[32397]_  = ~A200 & A199;
  assign \new_[32398]_  = A166 & \new_[32397]_ ;
  assign \new_[32399]_  = \new_[32398]_  & \new_[32393]_ ;
  assign \new_[32403]_  = A234 & A233;
  assign \new_[32404]_  = A203 & \new_[32403]_ ;
  assign \new_[32408]_  = A269 & A266;
  assign \new_[32409]_  = ~A265 & \new_[32408]_ ;
  assign \new_[32410]_  = \new_[32409]_  & \new_[32404]_ ;
  assign \new_[32414]_  = A167 & ~A168;
  assign \new_[32415]_  = ~A169 & \new_[32414]_ ;
  assign \new_[32419]_  = ~A200 & A199;
  assign \new_[32420]_  = A166 & \new_[32419]_ ;
  assign \new_[32421]_  = \new_[32420]_  & \new_[32415]_ ;
  assign \new_[32425]_  = A234 & A233;
  assign \new_[32426]_  = A203 & \new_[32425]_ ;
  assign \new_[32430]_  = A269 & ~A266;
  assign \new_[32431]_  = A265 & \new_[32430]_ ;
  assign \new_[32432]_  = \new_[32431]_  & \new_[32426]_ ;
  assign \new_[32436]_  = A167 & ~A168;
  assign \new_[32437]_  = ~A169 & \new_[32436]_ ;
  assign \new_[32441]_  = ~A200 & A199;
  assign \new_[32442]_  = A166 & \new_[32441]_ ;
  assign \new_[32443]_  = \new_[32442]_  & \new_[32437]_ ;
  assign \new_[32447]_  = A233 & ~A232;
  assign \new_[32448]_  = A203 & \new_[32447]_ ;
  assign \new_[32452]_  = A300 & A299;
  assign \new_[32453]_  = A236 & \new_[32452]_ ;
  assign \new_[32454]_  = \new_[32453]_  & \new_[32448]_ ;
  assign \new_[32458]_  = A167 & ~A168;
  assign \new_[32459]_  = ~A169 & \new_[32458]_ ;
  assign \new_[32463]_  = ~A200 & A199;
  assign \new_[32464]_  = A166 & \new_[32463]_ ;
  assign \new_[32465]_  = \new_[32464]_  & \new_[32459]_ ;
  assign \new_[32469]_  = A233 & ~A232;
  assign \new_[32470]_  = A203 & \new_[32469]_ ;
  assign \new_[32474]_  = A300 & A298;
  assign \new_[32475]_  = A236 & \new_[32474]_ ;
  assign \new_[32476]_  = \new_[32475]_  & \new_[32470]_ ;
  assign \new_[32480]_  = A167 & ~A168;
  assign \new_[32481]_  = ~A169 & \new_[32480]_ ;
  assign \new_[32485]_  = ~A200 & A199;
  assign \new_[32486]_  = A166 & \new_[32485]_ ;
  assign \new_[32487]_  = \new_[32486]_  & \new_[32481]_ ;
  assign \new_[32491]_  = A233 & ~A232;
  assign \new_[32492]_  = A203 & \new_[32491]_ ;
  assign \new_[32496]_  = A267 & A265;
  assign \new_[32497]_  = A236 & \new_[32496]_ ;
  assign \new_[32498]_  = \new_[32497]_  & \new_[32492]_ ;
  assign \new_[32502]_  = A167 & ~A168;
  assign \new_[32503]_  = ~A169 & \new_[32502]_ ;
  assign \new_[32507]_  = ~A200 & A199;
  assign \new_[32508]_  = A166 & \new_[32507]_ ;
  assign \new_[32509]_  = \new_[32508]_  & \new_[32503]_ ;
  assign \new_[32513]_  = A233 & ~A232;
  assign \new_[32514]_  = A203 & \new_[32513]_ ;
  assign \new_[32518]_  = A267 & A266;
  assign \new_[32519]_  = A236 & \new_[32518]_ ;
  assign \new_[32520]_  = \new_[32519]_  & \new_[32514]_ ;
  assign \new_[32524]_  = A167 & ~A168;
  assign \new_[32525]_  = ~A169 & \new_[32524]_ ;
  assign \new_[32529]_  = ~A200 & A199;
  assign \new_[32530]_  = A166 & \new_[32529]_ ;
  assign \new_[32531]_  = \new_[32530]_  & \new_[32525]_ ;
  assign \new_[32535]_  = ~A233 & A232;
  assign \new_[32536]_  = A203 & \new_[32535]_ ;
  assign \new_[32540]_  = A300 & A299;
  assign \new_[32541]_  = A236 & \new_[32540]_ ;
  assign \new_[32542]_  = \new_[32541]_  & \new_[32536]_ ;
  assign \new_[32546]_  = A167 & ~A168;
  assign \new_[32547]_  = ~A169 & \new_[32546]_ ;
  assign \new_[32551]_  = ~A200 & A199;
  assign \new_[32552]_  = A166 & \new_[32551]_ ;
  assign \new_[32553]_  = \new_[32552]_  & \new_[32547]_ ;
  assign \new_[32557]_  = ~A233 & A232;
  assign \new_[32558]_  = A203 & \new_[32557]_ ;
  assign \new_[32562]_  = A300 & A298;
  assign \new_[32563]_  = A236 & \new_[32562]_ ;
  assign \new_[32564]_  = \new_[32563]_  & \new_[32558]_ ;
  assign \new_[32568]_  = A167 & ~A168;
  assign \new_[32569]_  = ~A169 & \new_[32568]_ ;
  assign \new_[32573]_  = ~A200 & A199;
  assign \new_[32574]_  = A166 & \new_[32573]_ ;
  assign \new_[32575]_  = \new_[32574]_  & \new_[32569]_ ;
  assign \new_[32579]_  = ~A233 & A232;
  assign \new_[32580]_  = A203 & \new_[32579]_ ;
  assign \new_[32584]_  = A267 & A265;
  assign \new_[32585]_  = A236 & \new_[32584]_ ;
  assign \new_[32586]_  = \new_[32585]_  & \new_[32580]_ ;
  assign \new_[32590]_  = A167 & ~A168;
  assign \new_[32591]_  = ~A169 & \new_[32590]_ ;
  assign \new_[32595]_  = ~A200 & A199;
  assign \new_[32596]_  = A166 & \new_[32595]_ ;
  assign \new_[32597]_  = \new_[32596]_  & \new_[32591]_ ;
  assign \new_[32601]_  = ~A233 & A232;
  assign \new_[32602]_  = A203 & \new_[32601]_ ;
  assign \new_[32606]_  = A267 & A266;
  assign \new_[32607]_  = A236 & \new_[32606]_ ;
  assign \new_[32608]_  = \new_[32607]_  & \new_[32602]_ ;
  assign \new_[32612]_  = ~A168 & ~A169;
  assign \new_[32613]_  = ~A170 & \new_[32612]_ ;
  assign \new_[32617]_  = A203 & A200;
  assign \new_[32618]_  = ~A199 & \new_[32617]_ ;
  assign \new_[32619]_  = \new_[32618]_  & \new_[32613]_ ;
  assign \new_[32623]_  = A236 & A233;
  assign \new_[32624]_  = ~A232 & \new_[32623]_ ;
  assign \new_[32628]_  = A302 & ~A299;
  assign \new_[32629]_  = A298 & \new_[32628]_ ;
  assign \new_[32630]_  = \new_[32629]_  & \new_[32624]_ ;
  assign \new_[32634]_  = ~A168 & ~A169;
  assign \new_[32635]_  = ~A170 & \new_[32634]_ ;
  assign \new_[32639]_  = A203 & A200;
  assign \new_[32640]_  = ~A199 & \new_[32639]_ ;
  assign \new_[32641]_  = \new_[32640]_  & \new_[32635]_ ;
  assign \new_[32645]_  = A236 & A233;
  assign \new_[32646]_  = ~A232 & \new_[32645]_ ;
  assign \new_[32650]_  = A302 & A299;
  assign \new_[32651]_  = ~A298 & \new_[32650]_ ;
  assign \new_[32652]_  = \new_[32651]_  & \new_[32646]_ ;
  assign \new_[32656]_  = ~A168 & ~A169;
  assign \new_[32657]_  = ~A170 & \new_[32656]_ ;
  assign \new_[32661]_  = A203 & A200;
  assign \new_[32662]_  = ~A199 & \new_[32661]_ ;
  assign \new_[32663]_  = \new_[32662]_  & \new_[32657]_ ;
  assign \new_[32667]_  = A236 & A233;
  assign \new_[32668]_  = ~A232 & \new_[32667]_ ;
  assign \new_[32672]_  = A269 & A266;
  assign \new_[32673]_  = ~A265 & \new_[32672]_ ;
  assign \new_[32674]_  = \new_[32673]_  & \new_[32668]_ ;
  assign \new_[32678]_  = ~A168 & ~A169;
  assign \new_[32679]_  = ~A170 & \new_[32678]_ ;
  assign \new_[32683]_  = A203 & A200;
  assign \new_[32684]_  = ~A199 & \new_[32683]_ ;
  assign \new_[32685]_  = \new_[32684]_  & \new_[32679]_ ;
  assign \new_[32689]_  = A236 & A233;
  assign \new_[32690]_  = ~A232 & \new_[32689]_ ;
  assign \new_[32694]_  = A269 & ~A266;
  assign \new_[32695]_  = A265 & \new_[32694]_ ;
  assign \new_[32696]_  = \new_[32695]_  & \new_[32690]_ ;
  assign \new_[32700]_  = ~A168 & ~A169;
  assign \new_[32701]_  = ~A170 & \new_[32700]_ ;
  assign \new_[32705]_  = A203 & A200;
  assign \new_[32706]_  = ~A199 & \new_[32705]_ ;
  assign \new_[32707]_  = \new_[32706]_  & \new_[32701]_ ;
  assign \new_[32711]_  = A236 & ~A233;
  assign \new_[32712]_  = A232 & \new_[32711]_ ;
  assign \new_[32716]_  = A302 & ~A299;
  assign \new_[32717]_  = A298 & \new_[32716]_ ;
  assign \new_[32718]_  = \new_[32717]_  & \new_[32712]_ ;
  assign \new_[32722]_  = ~A168 & ~A169;
  assign \new_[32723]_  = ~A170 & \new_[32722]_ ;
  assign \new_[32727]_  = A203 & A200;
  assign \new_[32728]_  = ~A199 & \new_[32727]_ ;
  assign \new_[32729]_  = \new_[32728]_  & \new_[32723]_ ;
  assign \new_[32733]_  = A236 & ~A233;
  assign \new_[32734]_  = A232 & \new_[32733]_ ;
  assign \new_[32738]_  = A302 & A299;
  assign \new_[32739]_  = ~A298 & \new_[32738]_ ;
  assign \new_[32740]_  = \new_[32739]_  & \new_[32734]_ ;
  assign \new_[32744]_  = ~A168 & ~A169;
  assign \new_[32745]_  = ~A170 & \new_[32744]_ ;
  assign \new_[32749]_  = A203 & A200;
  assign \new_[32750]_  = ~A199 & \new_[32749]_ ;
  assign \new_[32751]_  = \new_[32750]_  & \new_[32745]_ ;
  assign \new_[32755]_  = A236 & ~A233;
  assign \new_[32756]_  = A232 & \new_[32755]_ ;
  assign \new_[32760]_  = A269 & A266;
  assign \new_[32761]_  = ~A265 & \new_[32760]_ ;
  assign \new_[32762]_  = \new_[32761]_  & \new_[32756]_ ;
  assign \new_[32766]_  = ~A168 & ~A169;
  assign \new_[32767]_  = ~A170 & \new_[32766]_ ;
  assign \new_[32771]_  = A203 & A200;
  assign \new_[32772]_  = ~A199 & \new_[32771]_ ;
  assign \new_[32773]_  = \new_[32772]_  & \new_[32767]_ ;
  assign \new_[32777]_  = A236 & ~A233;
  assign \new_[32778]_  = A232 & \new_[32777]_ ;
  assign \new_[32782]_  = A269 & ~A266;
  assign \new_[32783]_  = A265 & \new_[32782]_ ;
  assign \new_[32784]_  = \new_[32783]_  & \new_[32778]_ ;
  assign \new_[32788]_  = ~A168 & ~A169;
  assign \new_[32789]_  = ~A170 & \new_[32788]_ ;
  assign \new_[32793]_  = A203 & ~A200;
  assign \new_[32794]_  = A199 & \new_[32793]_ ;
  assign \new_[32795]_  = \new_[32794]_  & \new_[32789]_ ;
  assign \new_[32799]_  = A236 & A233;
  assign \new_[32800]_  = ~A232 & \new_[32799]_ ;
  assign \new_[32804]_  = A302 & ~A299;
  assign \new_[32805]_  = A298 & \new_[32804]_ ;
  assign \new_[32806]_  = \new_[32805]_  & \new_[32800]_ ;
  assign \new_[32810]_  = ~A168 & ~A169;
  assign \new_[32811]_  = ~A170 & \new_[32810]_ ;
  assign \new_[32815]_  = A203 & ~A200;
  assign \new_[32816]_  = A199 & \new_[32815]_ ;
  assign \new_[32817]_  = \new_[32816]_  & \new_[32811]_ ;
  assign \new_[32821]_  = A236 & A233;
  assign \new_[32822]_  = ~A232 & \new_[32821]_ ;
  assign \new_[32826]_  = A302 & A299;
  assign \new_[32827]_  = ~A298 & \new_[32826]_ ;
  assign \new_[32828]_  = \new_[32827]_  & \new_[32822]_ ;
  assign \new_[32832]_  = ~A168 & ~A169;
  assign \new_[32833]_  = ~A170 & \new_[32832]_ ;
  assign \new_[32837]_  = A203 & ~A200;
  assign \new_[32838]_  = A199 & \new_[32837]_ ;
  assign \new_[32839]_  = \new_[32838]_  & \new_[32833]_ ;
  assign \new_[32843]_  = A236 & A233;
  assign \new_[32844]_  = ~A232 & \new_[32843]_ ;
  assign \new_[32848]_  = A269 & A266;
  assign \new_[32849]_  = ~A265 & \new_[32848]_ ;
  assign \new_[32850]_  = \new_[32849]_  & \new_[32844]_ ;
  assign \new_[32854]_  = ~A168 & ~A169;
  assign \new_[32855]_  = ~A170 & \new_[32854]_ ;
  assign \new_[32859]_  = A203 & ~A200;
  assign \new_[32860]_  = A199 & \new_[32859]_ ;
  assign \new_[32861]_  = \new_[32860]_  & \new_[32855]_ ;
  assign \new_[32865]_  = A236 & A233;
  assign \new_[32866]_  = ~A232 & \new_[32865]_ ;
  assign \new_[32870]_  = A269 & ~A266;
  assign \new_[32871]_  = A265 & \new_[32870]_ ;
  assign \new_[32872]_  = \new_[32871]_  & \new_[32866]_ ;
  assign \new_[32876]_  = ~A168 & ~A169;
  assign \new_[32877]_  = ~A170 & \new_[32876]_ ;
  assign \new_[32881]_  = A203 & ~A200;
  assign \new_[32882]_  = A199 & \new_[32881]_ ;
  assign \new_[32883]_  = \new_[32882]_  & \new_[32877]_ ;
  assign \new_[32887]_  = A236 & ~A233;
  assign \new_[32888]_  = A232 & \new_[32887]_ ;
  assign \new_[32892]_  = A302 & ~A299;
  assign \new_[32893]_  = A298 & \new_[32892]_ ;
  assign \new_[32894]_  = \new_[32893]_  & \new_[32888]_ ;
  assign \new_[32898]_  = ~A168 & ~A169;
  assign \new_[32899]_  = ~A170 & \new_[32898]_ ;
  assign \new_[32903]_  = A203 & ~A200;
  assign \new_[32904]_  = A199 & \new_[32903]_ ;
  assign \new_[32905]_  = \new_[32904]_  & \new_[32899]_ ;
  assign \new_[32909]_  = A236 & ~A233;
  assign \new_[32910]_  = A232 & \new_[32909]_ ;
  assign \new_[32914]_  = A302 & A299;
  assign \new_[32915]_  = ~A298 & \new_[32914]_ ;
  assign \new_[32916]_  = \new_[32915]_  & \new_[32910]_ ;
  assign \new_[32920]_  = ~A168 & ~A169;
  assign \new_[32921]_  = ~A170 & \new_[32920]_ ;
  assign \new_[32925]_  = A203 & ~A200;
  assign \new_[32926]_  = A199 & \new_[32925]_ ;
  assign \new_[32927]_  = \new_[32926]_  & \new_[32921]_ ;
  assign \new_[32931]_  = A236 & ~A233;
  assign \new_[32932]_  = A232 & \new_[32931]_ ;
  assign \new_[32936]_  = A269 & A266;
  assign \new_[32937]_  = ~A265 & \new_[32936]_ ;
  assign \new_[32938]_  = \new_[32937]_  & \new_[32932]_ ;
  assign \new_[32942]_  = ~A168 & ~A169;
  assign \new_[32943]_  = ~A170 & \new_[32942]_ ;
  assign \new_[32947]_  = A203 & ~A200;
  assign \new_[32948]_  = A199 & \new_[32947]_ ;
  assign \new_[32949]_  = \new_[32948]_  & \new_[32943]_ ;
  assign \new_[32953]_  = A236 & ~A233;
  assign \new_[32954]_  = A232 & \new_[32953]_ ;
  assign \new_[32958]_  = A269 & ~A266;
  assign \new_[32959]_  = A265 & \new_[32958]_ ;
  assign \new_[32960]_  = \new_[32959]_  & \new_[32954]_ ;
  assign \new_[32964]_  = ~A166 & A167;
  assign \new_[32965]_  = A170 & \new_[32964]_ ;
  assign \new_[32969]_  = ~A201 & A200;
  assign \new_[32970]_  = A199 & \new_[32969]_ ;
  assign \new_[32971]_  = \new_[32970]_  & \new_[32965]_ ;
  assign \new_[32975]_  = A233 & ~A232;
  assign \new_[32976]_  = ~A202 & \new_[32975]_ ;
  assign \new_[32979]_  = A298 & A236;
  assign \new_[32982]_  = A302 & ~A299;
  assign \new_[32983]_  = \new_[32982]_  & \new_[32979]_ ;
  assign \new_[32984]_  = \new_[32983]_  & \new_[32976]_ ;
  assign \new_[32988]_  = ~A166 & A167;
  assign \new_[32989]_  = A170 & \new_[32988]_ ;
  assign \new_[32993]_  = ~A201 & A200;
  assign \new_[32994]_  = A199 & \new_[32993]_ ;
  assign \new_[32995]_  = \new_[32994]_  & \new_[32989]_ ;
  assign \new_[32999]_  = A233 & ~A232;
  assign \new_[33000]_  = ~A202 & \new_[32999]_ ;
  assign \new_[33003]_  = ~A298 & A236;
  assign \new_[33006]_  = A302 & A299;
  assign \new_[33007]_  = \new_[33006]_  & \new_[33003]_ ;
  assign \new_[33008]_  = \new_[33007]_  & \new_[33000]_ ;
  assign \new_[33012]_  = ~A166 & A167;
  assign \new_[33013]_  = A170 & \new_[33012]_ ;
  assign \new_[33017]_  = ~A201 & A200;
  assign \new_[33018]_  = A199 & \new_[33017]_ ;
  assign \new_[33019]_  = \new_[33018]_  & \new_[33013]_ ;
  assign \new_[33023]_  = A233 & ~A232;
  assign \new_[33024]_  = ~A202 & \new_[33023]_ ;
  assign \new_[33027]_  = ~A265 & A236;
  assign \new_[33030]_  = A269 & A266;
  assign \new_[33031]_  = \new_[33030]_  & \new_[33027]_ ;
  assign \new_[33032]_  = \new_[33031]_  & \new_[33024]_ ;
  assign \new_[33036]_  = ~A166 & A167;
  assign \new_[33037]_  = A170 & \new_[33036]_ ;
  assign \new_[33041]_  = ~A201 & A200;
  assign \new_[33042]_  = A199 & \new_[33041]_ ;
  assign \new_[33043]_  = \new_[33042]_  & \new_[33037]_ ;
  assign \new_[33047]_  = A233 & ~A232;
  assign \new_[33048]_  = ~A202 & \new_[33047]_ ;
  assign \new_[33051]_  = A265 & A236;
  assign \new_[33054]_  = A269 & ~A266;
  assign \new_[33055]_  = \new_[33054]_  & \new_[33051]_ ;
  assign \new_[33056]_  = \new_[33055]_  & \new_[33048]_ ;
  assign \new_[33060]_  = ~A166 & A167;
  assign \new_[33061]_  = A170 & \new_[33060]_ ;
  assign \new_[33065]_  = ~A201 & A200;
  assign \new_[33066]_  = A199 & \new_[33065]_ ;
  assign \new_[33067]_  = \new_[33066]_  & \new_[33061]_ ;
  assign \new_[33071]_  = ~A233 & A232;
  assign \new_[33072]_  = ~A202 & \new_[33071]_ ;
  assign \new_[33075]_  = A298 & A236;
  assign \new_[33078]_  = A302 & ~A299;
  assign \new_[33079]_  = \new_[33078]_  & \new_[33075]_ ;
  assign \new_[33080]_  = \new_[33079]_  & \new_[33072]_ ;
  assign \new_[33084]_  = ~A166 & A167;
  assign \new_[33085]_  = A170 & \new_[33084]_ ;
  assign \new_[33089]_  = ~A201 & A200;
  assign \new_[33090]_  = A199 & \new_[33089]_ ;
  assign \new_[33091]_  = \new_[33090]_  & \new_[33085]_ ;
  assign \new_[33095]_  = ~A233 & A232;
  assign \new_[33096]_  = ~A202 & \new_[33095]_ ;
  assign \new_[33099]_  = ~A298 & A236;
  assign \new_[33102]_  = A302 & A299;
  assign \new_[33103]_  = \new_[33102]_  & \new_[33099]_ ;
  assign \new_[33104]_  = \new_[33103]_  & \new_[33096]_ ;
  assign \new_[33108]_  = ~A166 & A167;
  assign \new_[33109]_  = A170 & \new_[33108]_ ;
  assign \new_[33113]_  = ~A201 & A200;
  assign \new_[33114]_  = A199 & \new_[33113]_ ;
  assign \new_[33115]_  = \new_[33114]_  & \new_[33109]_ ;
  assign \new_[33119]_  = ~A233 & A232;
  assign \new_[33120]_  = ~A202 & \new_[33119]_ ;
  assign \new_[33123]_  = ~A265 & A236;
  assign \new_[33126]_  = A269 & A266;
  assign \new_[33127]_  = \new_[33126]_  & \new_[33123]_ ;
  assign \new_[33128]_  = \new_[33127]_  & \new_[33120]_ ;
  assign \new_[33132]_  = ~A166 & A167;
  assign \new_[33133]_  = A170 & \new_[33132]_ ;
  assign \new_[33137]_  = ~A201 & A200;
  assign \new_[33138]_  = A199 & \new_[33137]_ ;
  assign \new_[33139]_  = \new_[33138]_  & \new_[33133]_ ;
  assign \new_[33143]_  = ~A233 & A232;
  assign \new_[33144]_  = ~A202 & \new_[33143]_ ;
  assign \new_[33147]_  = A265 & A236;
  assign \new_[33150]_  = A269 & ~A266;
  assign \new_[33151]_  = \new_[33150]_  & \new_[33147]_ ;
  assign \new_[33152]_  = \new_[33151]_  & \new_[33144]_ ;
  assign \new_[33156]_  = A166 & ~A167;
  assign \new_[33157]_  = A170 & \new_[33156]_ ;
  assign \new_[33161]_  = ~A201 & A200;
  assign \new_[33162]_  = A199 & \new_[33161]_ ;
  assign \new_[33163]_  = \new_[33162]_  & \new_[33157]_ ;
  assign \new_[33167]_  = A233 & ~A232;
  assign \new_[33168]_  = ~A202 & \new_[33167]_ ;
  assign \new_[33171]_  = A298 & A236;
  assign \new_[33174]_  = A302 & ~A299;
  assign \new_[33175]_  = \new_[33174]_  & \new_[33171]_ ;
  assign \new_[33176]_  = \new_[33175]_  & \new_[33168]_ ;
  assign \new_[33180]_  = A166 & ~A167;
  assign \new_[33181]_  = A170 & \new_[33180]_ ;
  assign \new_[33185]_  = ~A201 & A200;
  assign \new_[33186]_  = A199 & \new_[33185]_ ;
  assign \new_[33187]_  = \new_[33186]_  & \new_[33181]_ ;
  assign \new_[33191]_  = A233 & ~A232;
  assign \new_[33192]_  = ~A202 & \new_[33191]_ ;
  assign \new_[33195]_  = ~A298 & A236;
  assign \new_[33198]_  = A302 & A299;
  assign \new_[33199]_  = \new_[33198]_  & \new_[33195]_ ;
  assign \new_[33200]_  = \new_[33199]_  & \new_[33192]_ ;
  assign \new_[33204]_  = A166 & ~A167;
  assign \new_[33205]_  = A170 & \new_[33204]_ ;
  assign \new_[33209]_  = ~A201 & A200;
  assign \new_[33210]_  = A199 & \new_[33209]_ ;
  assign \new_[33211]_  = \new_[33210]_  & \new_[33205]_ ;
  assign \new_[33215]_  = A233 & ~A232;
  assign \new_[33216]_  = ~A202 & \new_[33215]_ ;
  assign \new_[33219]_  = ~A265 & A236;
  assign \new_[33222]_  = A269 & A266;
  assign \new_[33223]_  = \new_[33222]_  & \new_[33219]_ ;
  assign \new_[33224]_  = \new_[33223]_  & \new_[33216]_ ;
  assign \new_[33228]_  = A166 & ~A167;
  assign \new_[33229]_  = A170 & \new_[33228]_ ;
  assign \new_[33233]_  = ~A201 & A200;
  assign \new_[33234]_  = A199 & \new_[33233]_ ;
  assign \new_[33235]_  = \new_[33234]_  & \new_[33229]_ ;
  assign \new_[33239]_  = A233 & ~A232;
  assign \new_[33240]_  = ~A202 & \new_[33239]_ ;
  assign \new_[33243]_  = A265 & A236;
  assign \new_[33246]_  = A269 & ~A266;
  assign \new_[33247]_  = \new_[33246]_  & \new_[33243]_ ;
  assign \new_[33248]_  = \new_[33247]_  & \new_[33240]_ ;
  assign \new_[33252]_  = A166 & ~A167;
  assign \new_[33253]_  = A170 & \new_[33252]_ ;
  assign \new_[33257]_  = ~A201 & A200;
  assign \new_[33258]_  = A199 & \new_[33257]_ ;
  assign \new_[33259]_  = \new_[33258]_  & \new_[33253]_ ;
  assign \new_[33263]_  = ~A233 & A232;
  assign \new_[33264]_  = ~A202 & \new_[33263]_ ;
  assign \new_[33267]_  = A298 & A236;
  assign \new_[33270]_  = A302 & ~A299;
  assign \new_[33271]_  = \new_[33270]_  & \new_[33267]_ ;
  assign \new_[33272]_  = \new_[33271]_  & \new_[33264]_ ;
  assign \new_[33276]_  = A166 & ~A167;
  assign \new_[33277]_  = A170 & \new_[33276]_ ;
  assign \new_[33281]_  = ~A201 & A200;
  assign \new_[33282]_  = A199 & \new_[33281]_ ;
  assign \new_[33283]_  = \new_[33282]_  & \new_[33277]_ ;
  assign \new_[33287]_  = ~A233 & A232;
  assign \new_[33288]_  = ~A202 & \new_[33287]_ ;
  assign \new_[33291]_  = ~A298 & A236;
  assign \new_[33294]_  = A302 & A299;
  assign \new_[33295]_  = \new_[33294]_  & \new_[33291]_ ;
  assign \new_[33296]_  = \new_[33295]_  & \new_[33288]_ ;
  assign \new_[33300]_  = A166 & ~A167;
  assign \new_[33301]_  = A170 & \new_[33300]_ ;
  assign \new_[33305]_  = ~A201 & A200;
  assign \new_[33306]_  = A199 & \new_[33305]_ ;
  assign \new_[33307]_  = \new_[33306]_  & \new_[33301]_ ;
  assign \new_[33311]_  = ~A233 & A232;
  assign \new_[33312]_  = ~A202 & \new_[33311]_ ;
  assign \new_[33315]_  = ~A265 & A236;
  assign \new_[33318]_  = A269 & A266;
  assign \new_[33319]_  = \new_[33318]_  & \new_[33315]_ ;
  assign \new_[33320]_  = \new_[33319]_  & \new_[33312]_ ;
  assign \new_[33324]_  = A166 & ~A167;
  assign \new_[33325]_  = A170 & \new_[33324]_ ;
  assign \new_[33329]_  = ~A201 & A200;
  assign \new_[33330]_  = A199 & \new_[33329]_ ;
  assign \new_[33331]_  = \new_[33330]_  & \new_[33325]_ ;
  assign \new_[33335]_  = ~A233 & A232;
  assign \new_[33336]_  = ~A202 & \new_[33335]_ ;
  assign \new_[33339]_  = A265 & A236;
  assign \new_[33342]_  = A269 & ~A266;
  assign \new_[33343]_  = \new_[33342]_  & \new_[33339]_ ;
  assign \new_[33344]_  = \new_[33343]_  & \new_[33336]_ ;
  assign \new_[33348]_  = ~A202 & ~A201;
  assign \new_[33349]_  = A169 & \new_[33348]_ ;
  assign \new_[33353]_  = ~A235 & ~A234;
  assign \new_[33354]_  = ~A203 & \new_[33353]_ ;
  assign \new_[33355]_  = \new_[33354]_  & \new_[33349]_ ;
  assign \new_[33359]_  = ~A268 & ~A267;
  assign \new_[33360]_  = ~A236 & \new_[33359]_ ;
  assign \new_[33363]_  = ~A300 & ~A269;
  assign \new_[33366]_  = ~A302 & ~A301;
  assign \new_[33367]_  = \new_[33366]_  & \new_[33363]_ ;
  assign \new_[33368]_  = \new_[33367]_  & \new_[33360]_ ;
  assign \new_[33372]_  = ~A202 & ~A201;
  assign \new_[33373]_  = A169 & \new_[33372]_ ;
  assign \new_[33377]_  = ~A235 & ~A234;
  assign \new_[33378]_  = ~A203 & \new_[33377]_ ;
  assign \new_[33379]_  = \new_[33378]_  & \new_[33373]_ ;
  assign \new_[33383]_  = ~A268 & ~A267;
  assign \new_[33384]_  = ~A236 & \new_[33383]_ ;
  assign \new_[33387]_  = ~A298 & ~A269;
  assign \new_[33390]_  = ~A301 & ~A299;
  assign \new_[33391]_  = \new_[33390]_  & \new_[33387]_ ;
  assign \new_[33392]_  = \new_[33391]_  & \new_[33384]_ ;
  assign \new_[33396]_  = ~A202 & ~A201;
  assign \new_[33397]_  = A169 & \new_[33396]_ ;
  assign \new_[33401]_  = ~A235 & ~A234;
  assign \new_[33402]_  = ~A203 & \new_[33401]_ ;
  assign \new_[33403]_  = \new_[33402]_  & \new_[33397]_ ;
  assign \new_[33407]_  = ~A266 & ~A265;
  assign \new_[33408]_  = ~A236 & \new_[33407]_ ;
  assign \new_[33411]_  = ~A300 & ~A268;
  assign \new_[33414]_  = ~A302 & ~A301;
  assign \new_[33415]_  = \new_[33414]_  & \new_[33411]_ ;
  assign \new_[33416]_  = \new_[33415]_  & \new_[33408]_ ;
  assign \new_[33420]_  = ~A202 & ~A201;
  assign \new_[33421]_  = A169 & \new_[33420]_ ;
  assign \new_[33425]_  = ~A235 & ~A234;
  assign \new_[33426]_  = ~A203 & \new_[33425]_ ;
  assign \new_[33427]_  = \new_[33426]_  & \new_[33421]_ ;
  assign \new_[33431]_  = ~A266 & ~A265;
  assign \new_[33432]_  = ~A236 & \new_[33431]_ ;
  assign \new_[33435]_  = ~A298 & ~A268;
  assign \new_[33438]_  = ~A301 & ~A299;
  assign \new_[33439]_  = \new_[33438]_  & \new_[33435]_ ;
  assign \new_[33440]_  = \new_[33439]_  & \new_[33432]_ ;
  assign \new_[33444]_  = ~A202 & ~A201;
  assign \new_[33445]_  = A169 & \new_[33444]_ ;
  assign \new_[33449]_  = ~A233 & ~A232;
  assign \new_[33450]_  = ~A203 & \new_[33449]_ ;
  assign \new_[33451]_  = \new_[33450]_  & \new_[33445]_ ;
  assign \new_[33455]_  = ~A268 & ~A267;
  assign \new_[33456]_  = ~A235 & \new_[33455]_ ;
  assign \new_[33459]_  = ~A300 & ~A269;
  assign \new_[33462]_  = ~A302 & ~A301;
  assign \new_[33463]_  = \new_[33462]_  & \new_[33459]_ ;
  assign \new_[33464]_  = \new_[33463]_  & \new_[33456]_ ;
  assign \new_[33468]_  = ~A202 & ~A201;
  assign \new_[33469]_  = A169 & \new_[33468]_ ;
  assign \new_[33473]_  = ~A233 & ~A232;
  assign \new_[33474]_  = ~A203 & \new_[33473]_ ;
  assign \new_[33475]_  = \new_[33474]_  & \new_[33469]_ ;
  assign \new_[33479]_  = ~A268 & ~A267;
  assign \new_[33480]_  = ~A235 & \new_[33479]_ ;
  assign \new_[33483]_  = ~A298 & ~A269;
  assign \new_[33486]_  = ~A301 & ~A299;
  assign \new_[33487]_  = \new_[33486]_  & \new_[33483]_ ;
  assign \new_[33488]_  = \new_[33487]_  & \new_[33480]_ ;
  assign \new_[33492]_  = ~A202 & ~A201;
  assign \new_[33493]_  = A169 & \new_[33492]_ ;
  assign \new_[33497]_  = ~A233 & ~A232;
  assign \new_[33498]_  = ~A203 & \new_[33497]_ ;
  assign \new_[33499]_  = \new_[33498]_  & \new_[33493]_ ;
  assign \new_[33503]_  = ~A266 & ~A265;
  assign \new_[33504]_  = ~A235 & \new_[33503]_ ;
  assign \new_[33507]_  = ~A300 & ~A268;
  assign \new_[33510]_  = ~A302 & ~A301;
  assign \new_[33511]_  = \new_[33510]_  & \new_[33507]_ ;
  assign \new_[33512]_  = \new_[33511]_  & \new_[33504]_ ;
  assign \new_[33516]_  = ~A202 & ~A201;
  assign \new_[33517]_  = A169 & \new_[33516]_ ;
  assign \new_[33521]_  = ~A233 & ~A232;
  assign \new_[33522]_  = ~A203 & \new_[33521]_ ;
  assign \new_[33523]_  = \new_[33522]_  & \new_[33517]_ ;
  assign \new_[33527]_  = ~A266 & ~A265;
  assign \new_[33528]_  = ~A235 & \new_[33527]_ ;
  assign \new_[33531]_  = ~A298 & ~A268;
  assign \new_[33534]_  = ~A301 & ~A299;
  assign \new_[33535]_  = \new_[33534]_  & \new_[33531]_ ;
  assign \new_[33536]_  = \new_[33535]_  & \new_[33528]_ ;
  assign \new_[33540]_  = ~A200 & ~A199;
  assign \new_[33541]_  = A169 & \new_[33540]_ ;
  assign \new_[33545]_  = ~A235 & ~A234;
  assign \new_[33546]_  = ~A202 & \new_[33545]_ ;
  assign \new_[33547]_  = \new_[33546]_  & \new_[33541]_ ;
  assign \new_[33551]_  = ~A268 & ~A267;
  assign \new_[33552]_  = ~A236 & \new_[33551]_ ;
  assign \new_[33555]_  = ~A300 & ~A269;
  assign \new_[33558]_  = ~A302 & ~A301;
  assign \new_[33559]_  = \new_[33558]_  & \new_[33555]_ ;
  assign \new_[33560]_  = \new_[33559]_  & \new_[33552]_ ;
  assign \new_[33564]_  = ~A200 & ~A199;
  assign \new_[33565]_  = A169 & \new_[33564]_ ;
  assign \new_[33569]_  = ~A235 & ~A234;
  assign \new_[33570]_  = ~A202 & \new_[33569]_ ;
  assign \new_[33571]_  = \new_[33570]_  & \new_[33565]_ ;
  assign \new_[33575]_  = ~A268 & ~A267;
  assign \new_[33576]_  = ~A236 & \new_[33575]_ ;
  assign \new_[33579]_  = ~A298 & ~A269;
  assign \new_[33582]_  = ~A301 & ~A299;
  assign \new_[33583]_  = \new_[33582]_  & \new_[33579]_ ;
  assign \new_[33584]_  = \new_[33583]_  & \new_[33576]_ ;
  assign \new_[33588]_  = ~A200 & ~A199;
  assign \new_[33589]_  = A169 & \new_[33588]_ ;
  assign \new_[33593]_  = ~A235 & ~A234;
  assign \new_[33594]_  = ~A202 & \new_[33593]_ ;
  assign \new_[33595]_  = \new_[33594]_  & \new_[33589]_ ;
  assign \new_[33599]_  = ~A266 & ~A265;
  assign \new_[33600]_  = ~A236 & \new_[33599]_ ;
  assign \new_[33603]_  = ~A300 & ~A268;
  assign \new_[33606]_  = ~A302 & ~A301;
  assign \new_[33607]_  = \new_[33606]_  & \new_[33603]_ ;
  assign \new_[33608]_  = \new_[33607]_  & \new_[33600]_ ;
  assign \new_[33612]_  = ~A200 & ~A199;
  assign \new_[33613]_  = A169 & \new_[33612]_ ;
  assign \new_[33617]_  = ~A235 & ~A234;
  assign \new_[33618]_  = ~A202 & \new_[33617]_ ;
  assign \new_[33619]_  = \new_[33618]_  & \new_[33613]_ ;
  assign \new_[33623]_  = ~A266 & ~A265;
  assign \new_[33624]_  = ~A236 & \new_[33623]_ ;
  assign \new_[33627]_  = ~A298 & ~A268;
  assign \new_[33630]_  = ~A301 & ~A299;
  assign \new_[33631]_  = \new_[33630]_  & \new_[33627]_ ;
  assign \new_[33632]_  = \new_[33631]_  & \new_[33624]_ ;
  assign \new_[33636]_  = ~A200 & ~A199;
  assign \new_[33637]_  = A169 & \new_[33636]_ ;
  assign \new_[33641]_  = ~A233 & ~A232;
  assign \new_[33642]_  = ~A202 & \new_[33641]_ ;
  assign \new_[33643]_  = \new_[33642]_  & \new_[33637]_ ;
  assign \new_[33647]_  = ~A268 & ~A267;
  assign \new_[33648]_  = ~A235 & \new_[33647]_ ;
  assign \new_[33651]_  = ~A300 & ~A269;
  assign \new_[33654]_  = ~A302 & ~A301;
  assign \new_[33655]_  = \new_[33654]_  & \new_[33651]_ ;
  assign \new_[33656]_  = \new_[33655]_  & \new_[33648]_ ;
  assign \new_[33660]_  = ~A200 & ~A199;
  assign \new_[33661]_  = A169 & \new_[33660]_ ;
  assign \new_[33665]_  = ~A233 & ~A232;
  assign \new_[33666]_  = ~A202 & \new_[33665]_ ;
  assign \new_[33667]_  = \new_[33666]_  & \new_[33661]_ ;
  assign \new_[33671]_  = ~A268 & ~A267;
  assign \new_[33672]_  = ~A235 & \new_[33671]_ ;
  assign \new_[33675]_  = ~A298 & ~A269;
  assign \new_[33678]_  = ~A301 & ~A299;
  assign \new_[33679]_  = \new_[33678]_  & \new_[33675]_ ;
  assign \new_[33680]_  = \new_[33679]_  & \new_[33672]_ ;
  assign \new_[33684]_  = ~A200 & ~A199;
  assign \new_[33685]_  = A169 & \new_[33684]_ ;
  assign \new_[33689]_  = ~A233 & ~A232;
  assign \new_[33690]_  = ~A202 & \new_[33689]_ ;
  assign \new_[33691]_  = \new_[33690]_  & \new_[33685]_ ;
  assign \new_[33695]_  = ~A266 & ~A265;
  assign \new_[33696]_  = ~A235 & \new_[33695]_ ;
  assign \new_[33699]_  = ~A300 & ~A268;
  assign \new_[33702]_  = ~A302 & ~A301;
  assign \new_[33703]_  = \new_[33702]_  & \new_[33699]_ ;
  assign \new_[33704]_  = \new_[33703]_  & \new_[33696]_ ;
  assign \new_[33708]_  = ~A200 & ~A199;
  assign \new_[33709]_  = A169 & \new_[33708]_ ;
  assign \new_[33713]_  = ~A233 & ~A232;
  assign \new_[33714]_  = ~A202 & \new_[33713]_ ;
  assign \new_[33715]_  = \new_[33714]_  & \new_[33709]_ ;
  assign \new_[33719]_  = ~A266 & ~A265;
  assign \new_[33720]_  = ~A235 & \new_[33719]_ ;
  assign \new_[33723]_  = ~A298 & ~A268;
  assign \new_[33726]_  = ~A301 & ~A299;
  assign \new_[33727]_  = \new_[33726]_  & \new_[33723]_ ;
  assign \new_[33728]_  = \new_[33727]_  & \new_[33720]_ ;
  assign \new_[33732]_  = ~A166 & ~A167;
  assign \new_[33733]_  = ~A169 & \new_[33732]_ ;
  assign \new_[33737]_  = ~A235 & ~A234;
  assign \new_[33738]_  = A202 & \new_[33737]_ ;
  assign \new_[33739]_  = \new_[33738]_  & \new_[33733]_ ;
  assign \new_[33743]_  = ~A268 & ~A267;
  assign \new_[33744]_  = ~A236 & \new_[33743]_ ;
  assign \new_[33747]_  = ~A300 & ~A269;
  assign \new_[33750]_  = ~A302 & ~A301;
  assign \new_[33751]_  = \new_[33750]_  & \new_[33747]_ ;
  assign \new_[33752]_  = \new_[33751]_  & \new_[33744]_ ;
  assign \new_[33756]_  = ~A166 & ~A167;
  assign \new_[33757]_  = ~A169 & \new_[33756]_ ;
  assign \new_[33761]_  = ~A235 & ~A234;
  assign \new_[33762]_  = A202 & \new_[33761]_ ;
  assign \new_[33763]_  = \new_[33762]_  & \new_[33757]_ ;
  assign \new_[33767]_  = ~A268 & ~A267;
  assign \new_[33768]_  = ~A236 & \new_[33767]_ ;
  assign \new_[33771]_  = ~A298 & ~A269;
  assign \new_[33774]_  = ~A301 & ~A299;
  assign \new_[33775]_  = \new_[33774]_  & \new_[33771]_ ;
  assign \new_[33776]_  = \new_[33775]_  & \new_[33768]_ ;
  assign \new_[33780]_  = ~A166 & ~A167;
  assign \new_[33781]_  = ~A169 & \new_[33780]_ ;
  assign \new_[33785]_  = ~A235 & ~A234;
  assign \new_[33786]_  = A202 & \new_[33785]_ ;
  assign \new_[33787]_  = \new_[33786]_  & \new_[33781]_ ;
  assign \new_[33791]_  = ~A266 & ~A265;
  assign \new_[33792]_  = ~A236 & \new_[33791]_ ;
  assign \new_[33795]_  = ~A300 & ~A268;
  assign \new_[33798]_  = ~A302 & ~A301;
  assign \new_[33799]_  = \new_[33798]_  & \new_[33795]_ ;
  assign \new_[33800]_  = \new_[33799]_  & \new_[33792]_ ;
  assign \new_[33804]_  = ~A166 & ~A167;
  assign \new_[33805]_  = ~A169 & \new_[33804]_ ;
  assign \new_[33809]_  = ~A235 & ~A234;
  assign \new_[33810]_  = A202 & \new_[33809]_ ;
  assign \new_[33811]_  = \new_[33810]_  & \new_[33805]_ ;
  assign \new_[33815]_  = ~A266 & ~A265;
  assign \new_[33816]_  = ~A236 & \new_[33815]_ ;
  assign \new_[33819]_  = ~A298 & ~A268;
  assign \new_[33822]_  = ~A301 & ~A299;
  assign \new_[33823]_  = \new_[33822]_  & \new_[33819]_ ;
  assign \new_[33824]_  = \new_[33823]_  & \new_[33816]_ ;
  assign \new_[33828]_  = ~A166 & ~A167;
  assign \new_[33829]_  = ~A169 & \new_[33828]_ ;
  assign \new_[33833]_  = ~A233 & ~A232;
  assign \new_[33834]_  = A202 & \new_[33833]_ ;
  assign \new_[33835]_  = \new_[33834]_  & \new_[33829]_ ;
  assign \new_[33839]_  = ~A268 & ~A267;
  assign \new_[33840]_  = ~A235 & \new_[33839]_ ;
  assign \new_[33843]_  = ~A300 & ~A269;
  assign \new_[33846]_  = ~A302 & ~A301;
  assign \new_[33847]_  = \new_[33846]_  & \new_[33843]_ ;
  assign \new_[33848]_  = \new_[33847]_  & \new_[33840]_ ;
  assign \new_[33852]_  = ~A166 & ~A167;
  assign \new_[33853]_  = ~A169 & \new_[33852]_ ;
  assign \new_[33857]_  = ~A233 & ~A232;
  assign \new_[33858]_  = A202 & \new_[33857]_ ;
  assign \new_[33859]_  = \new_[33858]_  & \new_[33853]_ ;
  assign \new_[33863]_  = ~A268 & ~A267;
  assign \new_[33864]_  = ~A235 & \new_[33863]_ ;
  assign \new_[33867]_  = ~A298 & ~A269;
  assign \new_[33870]_  = ~A301 & ~A299;
  assign \new_[33871]_  = \new_[33870]_  & \new_[33867]_ ;
  assign \new_[33872]_  = \new_[33871]_  & \new_[33864]_ ;
  assign \new_[33876]_  = ~A166 & ~A167;
  assign \new_[33877]_  = ~A169 & \new_[33876]_ ;
  assign \new_[33881]_  = ~A233 & ~A232;
  assign \new_[33882]_  = A202 & \new_[33881]_ ;
  assign \new_[33883]_  = \new_[33882]_  & \new_[33877]_ ;
  assign \new_[33887]_  = ~A266 & ~A265;
  assign \new_[33888]_  = ~A235 & \new_[33887]_ ;
  assign \new_[33891]_  = ~A300 & ~A268;
  assign \new_[33894]_  = ~A302 & ~A301;
  assign \new_[33895]_  = \new_[33894]_  & \new_[33891]_ ;
  assign \new_[33896]_  = \new_[33895]_  & \new_[33888]_ ;
  assign \new_[33900]_  = ~A166 & ~A167;
  assign \new_[33901]_  = ~A169 & \new_[33900]_ ;
  assign \new_[33905]_  = ~A233 & ~A232;
  assign \new_[33906]_  = A202 & \new_[33905]_ ;
  assign \new_[33907]_  = \new_[33906]_  & \new_[33901]_ ;
  assign \new_[33911]_  = ~A266 & ~A265;
  assign \new_[33912]_  = ~A235 & \new_[33911]_ ;
  assign \new_[33915]_  = ~A298 & ~A268;
  assign \new_[33918]_  = ~A301 & ~A299;
  assign \new_[33919]_  = \new_[33918]_  & \new_[33915]_ ;
  assign \new_[33920]_  = \new_[33919]_  & \new_[33912]_ ;
  assign \new_[33924]_  = A167 & ~A168;
  assign \new_[33925]_  = ~A169 & \new_[33924]_ ;
  assign \new_[33929]_  = A200 & ~A199;
  assign \new_[33930]_  = A166 & \new_[33929]_ ;
  assign \new_[33931]_  = \new_[33930]_  & \new_[33925]_ ;
  assign \new_[33935]_  = A233 & ~A232;
  assign \new_[33936]_  = A203 & \new_[33935]_ ;
  assign \new_[33939]_  = A298 & A236;
  assign \new_[33942]_  = A302 & ~A299;
  assign \new_[33943]_  = \new_[33942]_  & \new_[33939]_ ;
  assign \new_[33944]_  = \new_[33943]_  & \new_[33936]_ ;
  assign \new_[33948]_  = A167 & ~A168;
  assign \new_[33949]_  = ~A169 & \new_[33948]_ ;
  assign \new_[33953]_  = A200 & ~A199;
  assign \new_[33954]_  = A166 & \new_[33953]_ ;
  assign \new_[33955]_  = \new_[33954]_  & \new_[33949]_ ;
  assign \new_[33959]_  = A233 & ~A232;
  assign \new_[33960]_  = A203 & \new_[33959]_ ;
  assign \new_[33963]_  = ~A298 & A236;
  assign \new_[33966]_  = A302 & A299;
  assign \new_[33967]_  = \new_[33966]_  & \new_[33963]_ ;
  assign \new_[33968]_  = \new_[33967]_  & \new_[33960]_ ;
  assign \new_[33972]_  = A167 & ~A168;
  assign \new_[33973]_  = ~A169 & \new_[33972]_ ;
  assign \new_[33977]_  = A200 & ~A199;
  assign \new_[33978]_  = A166 & \new_[33977]_ ;
  assign \new_[33979]_  = \new_[33978]_  & \new_[33973]_ ;
  assign \new_[33983]_  = A233 & ~A232;
  assign \new_[33984]_  = A203 & \new_[33983]_ ;
  assign \new_[33987]_  = ~A265 & A236;
  assign \new_[33990]_  = A269 & A266;
  assign \new_[33991]_  = \new_[33990]_  & \new_[33987]_ ;
  assign \new_[33992]_  = \new_[33991]_  & \new_[33984]_ ;
  assign \new_[33996]_  = A167 & ~A168;
  assign \new_[33997]_  = ~A169 & \new_[33996]_ ;
  assign \new_[34001]_  = A200 & ~A199;
  assign \new_[34002]_  = A166 & \new_[34001]_ ;
  assign \new_[34003]_  = \new_[34002]_  & \new_[33997]_ ;
  assign \new_[34007]_  = A233 & ~A232;
  assign \new_[34008]_  = A203 & \new_[34007]_ ;
  assign \new_[34011]_  = A265 & A236;
  assign \new_[34014]_  = A269 & ~A266;
  assign \new_[34015]_  = \new_[34014]_  & \new_[34011]_ ;
  assign \new_[34016]_  = \new_[34015]_  & \new_[34008]_ ;
  assign \new_[34020]_  = A167 & ~A168;
  assign \new_[34021]_  = ~A169 & \new_[34020]_ ;
  assign \new_[34025]_  = A200 & ~A199;
  assign \new_[34026]_  = A166 & \new_[34025]_ ;
  assign \new_[34027]_  = \new_[34026]_  & \new_[34021]_ ;
  assign \new_[34031]_  = ~A233 & A232;
  assign \new_[34032]_  = A203 & \new_[34031]_ ;
  assign \new_[34035]_  = A298 & A236;
  assign \new_[34038]_  = A302 & ~A299;
  assign \new_[34039]_  = \new_[34038]_  & \new_[34035]_ ;
  assign \new_[34040]_  = \new_[34039]_  & \new_[34032]_ ;
  assign \new_[34044]_  = A167 & ~A168;
  assign \new_[34045]_  = ~A169 & \new_[34044]_ ;
  assign \new_[34049]_  = A200 & ~A199;
  assign \new_[34050]_  = A166 & \new_[34049]_ ;
  assign \new_[34051]_  = \new_[34050]_  & \new_[34045]_ ;
  assign \new_[34055]_  = ~A233 & A232;
  assign \new_[34056]_  = A203 & \new_[34055]_ ;
  assign \new_[34059]_  = ~A298 & A236;
  assign \new_[34062]_  = A302 & A299;
  assign \new_[34063]_  = \new_[34062]_  & \new_[34059]_ ;
  assign \new_[34064]_  = \new_[34063]_  & \new_[34056]_ ;
  assign \new_[34068]_  = A167 & ~A168;
  assign \new_[34069]_  = ~A169 & \new_[34068]_ ;
  assign \new_[34073]_  = A200 & ~A199;
  assign \new_[34074]_  = A166 & \new_[34073]_ ;
  assign \new_[34075]_  = \new_[34074]_  & \new_[34069]_ ;
  assign \new_[34079]_  = ~A233 & A232;
  assign \new_[34080]_  = A203 & \new_[34079]_ ;
  assign \new_[34083]_  = ~A265 & A236;
  assign \new_[34086]_  = A269 & A266;
  assign \new_[34087]_  = \new_[34086]_  & \new_[34083]_ ;
  assign \new_[34088]_  = \new_[34087]_  & \new_[34080]_ ;
  assign \new_[34092]_  = A167 & ~A168;
  assign \new_[34093]_  = ~A169 & \new_[34092]_ ;
  assign \new_[34097]_  = A200 & ~A199;
  assign \new_[34098]_  = A166 & \new_[34097]_ ;
  assign \new_[34099]_  = \new_[34098]_  & \new_[34093]_ ;
  assign \new_[34103]_  = ~A233 & A232;
  assign \new_[34104]_  = A203 & \new_[34103]_ ;
  assign \new_[34107]_  = A265 & A236;
  assign \new_[34110]_  = A269 & ~A266;
  assign \new_[34111]_  = \new_[34110]_  & \new_[34107]_ ;
  assign \new_[34112]_  = \new_[34111]_  & \new_[34104]_ ;
  assign \new_[34116]_  = A167 & ~A168;
  assign \new_[34117]_  = ~A169 & \new_[34116]_ ;
  assign \new_[34121]_  = ~A200 & A199;
  assign \new_[34122]_  = A166 & \new_[34121]_ ;
  assign \new_[34123]_  = \new_[34122]_  & \new_[34117]_ ;
  assign \new_[34127]_  = A233 & ~A232;
  assign \new_[34128]_  = A203 & \new_[34127]_ ;
  assign \new_[34131]_  = A298 & A236;
  assign \new_[34134]_  = A302 & ~A299;
  assign \new_[34135]_  = \new_[34134]_  & \new_[34131]_ ;
  assign \new_[34136]_  = \new_[34135]_  & \new_[34128]_ ;
  assign \new_[34140]_  = A167 & ~A168;
  assign \new_[34141]_  = ~A169 & \new_[34140]_ ;
  assign \new_[34145]_  = ~A200 & A199;
  assign \new_[34146]_  = A166 & \new_[34145]_ ;
  assign \new_[34147]_  = \new_[34146]_  & \new_[34141]_ ;
  assign \new_[34151]_  = A233 & ~A232;
  assign \new_[34152]_  = A203 & \new_[34151]_ ;
  assign \new_[34155]_  = ~A298 & A236;
  assign \new_[34158]_  = A302 & A299;
  assign \new_[34159]_  = \new_[34158]_  & \new_[34155]_ ;
  assign \new_[34160]_  = \new_[34159]_  & \new_[34152]_ ;
  assign \new_[34164]_  = A167 & ~A168;
  assign \new_[34165]_  = ~A169 & \new_[34164]_ ;
  assign \new_[34169]_  = ~A200 & A199;
  assign \new_[34170]_  = A166 & \new_[34169]_ ;
  assign \new_[34171]_  = \new_[34170]_  & \new_[34165]_ ;
  assign \new_[34175]_  = A233 & ~A232;
  assign \new_[34176]_  = A203 & \new_[34175]_ ;
  assign \new_[34179]_  = ~A265 & A236;
  assign \new_[34182]_  = A269 & A266;
  assign \new_[34183]_  = \new_[34182]_  & \new_[34179]_ ;
  assign \new_[34184]_  = \new_[34183]_  & \new_[34176]_ ;
  assign \new_[34188]_  = A167 & ~A168;
  assign \new_[34189]_  = ~A169 & \new_[34188]_ ;
  assign \new_[34193]_  = ~A200 & A199;
  assign \new_[34194]_  = A166 & \new_[34193]_ ;
  assign \new_[34195]_  = \new_[34194]_  & \new_[34189]_ ;
  assign \new_[34199]_  = A233 & ~A232;
  assign \new_[34200]_  = A203 & \new_[34199]_ ;
  assign \new_[34203]_  = A265 & A236;
  assign \new_[34206]_  = A269 & ~A266;
  assign \new_[34207]_  = \new_[34206]_  & \new_[34203]_ ;
  assign \new_[34208]_  = \new_[34207]_  & \new_[34200]_ ;
  assign \new_[34212]_  = A167 & ~A168;
  assign \new_[34213]_  = ~A169 & \new_[34212]_ ;
  assign \new_[34217]_  = ~A200 & A199;
  assign \new_[34218]_  = A166 & \new_[34217]_ ;
  assign \new_[34219]_  = \new_[34218]_  & \new_[34213]_ ;
  assign \new_[34223]_  = ~A233 & A232;
  assign \new_[34224]_  = A203 & \new_[34223]_ ;
  assign \new_[34227]_  = A298 & A236;
  assign \new_[34230]_  = A302 & ~A299;
  assign \new_[34231]_  = \new_[34230]_  & \new_[34227]_ ;
  assign \new_[34232]_  = \new_[34231]_  & \new_[34224]_ ;
  assign \new_[34236]_  = A167 & ~A168;
  assign \new_[34237]_  = ~A169 & \new_[34236]_ ;
  assign \new_[34241]_  = ~A200 & A199;
  assign \new_[34242]_  = A166 & \new_[34241]_ ;
  assign \new_[34243]_  = \new_[34242]_  & \new_[34237]_ ;
  assign \new_[34247]_  = ~A233 & A232;
  assign \new_[34248]_  = A203 & \new_[34247]_ ;
  assign \new_[34251]_  = ~A298 & A236;
  assign \new_[34254]_  = A302 & A299;
  assign \new_[34255]_  = \new_[34254]_  & \new_[34251]_ ;
  assign \new_[34256]_  = \new_[34255]_  & \new_[34248]_ ;
  assign \new_[34260]_  = A167 & ~A168;
  assign \new_[34261]_  = ~A169 & \new_[34260]_ ;
  assign \new_[34265]_  = ~A200 & A199;
  assign \new_[34266]_  = A166 & \new_[34265]_ ;
  assign \new_[34267]_  = \new_[34266]_  & \new_[34261]_ ;
  assign \new_[34271]_  = ~A233 & A232;
  assign \new_[34272]_  = A203 & \new_[34271]_ ;
  assign \new_[34275]_  = ~A265 & A236;
  assign \new_[34278]_  = A269 & A266;
  assign \new_[34279]_  = \new_[34278]_  & \new_[34275]_ ;
  assign \new_[34280]_  = \new_[34279]_  & \new_[34272]_ ;
  assign \new_[34284]_  = A167 & ~A168;
  assign \new_[34285]_  = ~A169 & \new_[34284]_ ;
  assign \new_[34289]_  = ~A200 & A199;
  assign \new_[34290]_  = A166 & \new_[34289]_ ;
  assign \new_[34291]_  = \new_[34290]_  & \new_[34285]_ ;
  assign \new_[34295]_  = ~A233 & A232;
  assign \new_[34296]_  = A203 & \new_[34295]_ ;
  assign \new_[34299]_  = A265 & A236;
  assign \new_[34302]_  = A269 & ~A266;
  assign \new_[34303]_  = \new_[34302]_  & \new_[34299]_ ;
  assign \new_[34304]_  = \new_[34303]_  & \new_[34296]_ ;
  assign \new_[34308]_  = ~A168 & ~A169;
  assign \new_[34309]_  = ~A170 & \new_[34308]_ ;
  assign \new_[34313]_  = ~A235 & ~A234;
  assign \new_[34314]_  = A202 & \new_[34313]_ ;
  assign \new_[34315]_  = \new_[34314]_  & \new_[34309]_ ;
  assign \new_[34319]_  = ~A268 & ~A267;
  assign \new_[34320]_  = ~A236 & \new_[34319]_ ;
  assign \new_[34323]_  = ~A300 & ~A269;
  assign \new_[34326]_  = ~A302 & ~A301;
  assign \new_[34327]_  = \new_[34326]_  & \new_[34323]_ ;
  assign \new_[34328]_  = \new_[34327]_  & \new_[34320]_ ;
  assign \new_[34332]_  = ~A168 & ~A169;
  assign \new_[34333]_  = ~A170 & \new_[34332]_ ;
  assign \new_[34337]_  = ~A235 & ~A234;
  assign \new_[34338]_  = A202 & \new_[34337]_ ;
  assign \new_[34339]_  = \new_[34338]_  & \new_[34333]_ ;
  assign \new_[34343]_  = ~A268 & ~A267;
  assign \new_[34344]_  = ~A236 & \new_[34343]_ ;
  assign \new_[34347]_  = ~A298 & ~A269;
  assign \new_[34350]_  = ~A301 & ~A299;
  assign \new_[34351]_  = \new_[34350]_  & \new_[34347]_ ;
  assign \new_[34352]_  = \new_[34351]_  & \new_[34344]_ ;
  assign \new_[34356]_  = ~A168 & ~A169;
  assign \new_[34357]_  = ~A170 & \new_[34356]_ ;
  assign \new_[34361]_  = ~A235 & ~A234;
  assign \new_[34362]_  = A202 & \new_[34361]_ ;
  assign \new_[34363]_  = \new_[34362]_  & \new_[34357]_ ;
  assign \new_[34367]_  = ~A266 & ~A265;
  assign \new_[34368]_  = ~A236 & \new_[34367]_ ;
  assign \new_[34371]_  = ~A300 & ~A268;
  assign \new_[34374]_  = ~A302 & ~A301;
  assign \new_[34375]_  = \new_[34374]_  & \new_[34371]_ ;
  assign \new_[34376]_  = \new_[34375]_  & \new_[34368]_ ;
  assign \new_[34380]_  = ~A168 & ~A169;
  assign \new_[34381]_  = ~A170 & \new_[34380]_ ;
  assign \new_[34385]_  = ~A235 & ~A234;
  assign \new_[34386]_  = A202 & \new_[34385]_ ;
  assign \new_[34387]_  = \new_[34386]_  & \new_[34381]_ ;
  assign \new_[34391]_  = ~A266 & ~A265;
  assign \new_[34392]_  = ~A236 & \new_[34391]_ ;
  assign \new_[34395]_  = ~A298 & ~A268;
  assign \new_[34398]_  = ~A301 & ~A299;
  assign \new_[34399]_  = \new_[34398]_  & \new_[34395]_ ;
  assign \new_[34400]_  = \new_[34399]_  & \new_[34392]_ ;
  assign \new_[34404]_  = ~A168 & ~A169;
  assign \new_[34405]_  = ~A170 & \new_[34404]_ ;
  assign \new_[34409]_  = ~A233 & ~A232;
  assign \new_[34410]_  = A202 & \new_[34409]_ ;
  assign \new_[34411]_  = \new_[34410]_  & \new_[34405]_ ;
  assign \new_[34415]_  = ~A268 & ~A267;
  assign \new_[34416]_  = ~A235 & \new_[34415]_ ;
  assign \new_[34419]_  = ~A300 & ~A269;
  assign \new_[34422]_  = ~A302 & ~A301;
  assign \new_[34423]_  = \new_[34422]_  & \new_[34419]_ ;
  assign \new_[34424]_  = \new_[34423]_  & \new_[34416]_ ;
  assign \new_[34428]_  = ~A168 & ~A169;
  assign \new_[34429]_  = ~A170 & \new_[34428]_ ;
  assign \new_[34433]_  = ~A233 & ~A232;
  assign \new_[34434]_  = A202 & \new_[34433]_ ;
  assign \new_[34435]_  = \new_[34434]_  & \new_[34429]_ ;
  assign \new_[34439]_  = ~A268 & ~A267;
  assign \new_[34440]_  = ~A235 & \new_[34439]_ ;
  assign \new_[34443]_  = ~A298 & ~A269;
  assign \new_[34446]_  = ~A301 & ~A299;
  assign \new_[34447]_  = \new_[34446]_  & \new_[34443]_ ;
  assign \new_[34448]_  = \new_[34447]_  & \new_[34440]_ ;
  assign \new_[34452]_  = ~A168 & ~A169;
  assign \new_[34453]_  = ~A170 & \new_[34452]_ ;
  assign \new_[34457]_  = ~A233 & ~A232;
  assign \new_[34458]_  = A202 & \new_[34457]_ ;
  assign \new_[34459]_  = \new_[34458]_  & \new_[34453]_ ;
  assign \new_[34463]_  = ~A266 & ~A265;
  assign \new_[34464]_  = ~A235 & \new_[34463]_ ;
  assign \new_[34467]_  = ~A300 & ~A268;
  assign \new_[34470]_  = ~A302 & ~A301;
  assign \new_[34471]_  = \new_[34470]_  & \new_[34467]_ ;
  assign \new_[34472]_  = \new_[34471]_  & \new_[34464]_ ;
  assign \new_[34476]_  = ~A168 & ~A169;
  assign \new_[34477]_  = ~A170 & \new_[34476]_ ;
  assign \new_[34481]_  = ~A233 & ~A232;
  assign \new_[34482]_  = A202 & \new_[34481]_ ;
  assign \new_[34483]_  = \new_[34482]_  & \new_[34477]_ ;
  assign \new_[34487]_  = ~A266 & ~A265;
  assign \new_[34488]_  = ~A235 & \new_[34487]_ ;
  assign \new_[34491]_  = ~A298 & ~A268;
  assign \new_[34494]_  = ~A301 & ~A299;
  assign \new_[34495]_  = \new_[34494]_  & \new_[34491]_ ;
  assign \new_[34496]_  = \new_[34495]_  & \new_[34488]_ ;
  assign \new_[34500]_  = ~A201 & A166;
  assign \new_[34501]_  = A168 & \new_[34500]_ ;
  assign \new_[34504]_  = ~A203 & ~A202;
  assign \new_[34507]_  = ~A235 & ~A234;
  assign \new_[34508]_  = \new_[34507]_  & \new_[34504]_ ;
  assign \new_[34509]_  = \new_[34508]_  & \new_[34501]_ ;
  assign \new_[34513]_  = ~A268 & ~A267;
  assign \new_[34514]_  = ~A236 & \new_[34513]_ ;
  assign \new_[34517]_  = ~A300 & ~A269;
  assign \new_[34520]_  = ~A302 & ~A301;
  assign \new_[34521]_  = \new_[34520]_  & \new_[34517]_ ;
  assign \new_[34522]_  = \new_[34521]_  & \new_[34514]_ ;
  assign \new_[34526]_  = ~A201 & A166;
  assign \new_[34527]_  = A168 & \new_[34526]_ ;
  assign \new_[34530]_  = ~A203 & ~A202;
  assign \new_[34533]_  = ~A235 & ~A234;
  assign \new_[34534]_  = \new_[34533]_  & \new_[34530]_ ;
  assign \new_[34535]_  = \new_[34534]_  & \new_[34527]_ ;
  assign \new_[34539]_  = ~A268 & ~A267;
  assign \new_[34540]_  = ~A236 & \new_[34539]_ ;
  assign \new_[34543]_  = ~A298 & ~A269;
  assign \new_[34546]_  = ~A301 & ~A299;
  assign \new_[34547]_  = \new_[34546]_  & \new_[34543]_ ;
  assign \new_[34548]_  = \new_[34547]_  & \new_[34540]_ ;
  assign \new_[34552]_  = ~A201 & A166;
  assign \new_[34553]_  = A168 & \new_[34552]_ ;
  assign \new_[34556]_  = ~A203 & ~A202;
  assign \new_[34559]_  = ~A235 & ~A234;
  assign \new_[34560]_  = \new_[34559]_  & \new_[34556]_ ;
  assign \new_[34561]_  = \new_[34560]_  & \new_[34553]_ ;
  assign \new_[34565]_  = ~A266 & ~A265;
  assign \new_[34566]_  = ~A236 & \new_[34565]_ ;
  assign \new_[34569]_  = ~A300 & ~A268;
  assign \new_[34572]_  = ~A302 & ~A301;
  assign \new_[34573]_  = \new_[34572]_  & \new_[34569]_ ;
  assign \new_[34574]_  = \new_[34573]_  & \new_[34566]_ ;
  assign \new_[34578]_  = ~A201 & A166;
  assign \new_[34579]_  = A168 & \new_[34578]_ ;
  assign \new_[34582]_  = ~A203 & ~A202;
  assign \new_[34585]_  = ~A235 & ~A234;
  assign \new_[34586]_  = \new_[34585]_  & \new_[34582]_ ;
  assign \new_[34587]_  = \new_[34586]_  & \new_[34579]_ ;
  assign \new_[34591]_  = ~A266 & ~A265;
  assign \new_[34592]_  = ~A236 & \new_[34591]_ ;
  assign \new_[34595]_  = ~A298 & ~A268;
  assign \new_[34598]_  = ~A301 & ~A299;
  assign \new_[34599]_  = \new_[34598]_  & \new_[34595]_ ;
  assign \new_[34600]_  = \new_[34599]_  & \new_[34592]_ ;
  assign \new_[34604]_  = ~A201 & A166;
  assign \new_[34605]_  = A168 & \new_[34604]_ ;
  assign \new_[34608]_  = ~A203 & ~A202;
  assign \new_[34611]_  = ~A233 & ~A232;
  assign \new_[34612]_  = \new_[34611]_  & \new_[34608]_ ;
  assign \new_[34613]_  = \new_[34612]_  & \new_[34605]_ ;
  assign \new_[34617]_  = ~A268 & ~A267;
  assign \new_[34618]_  = ~A235 & \new_[34617]_ ;
  assign \new_[34621]_  = ~A300 & ~A269;
  assign \new_[34624]_  = ~A302 & ~A301;
  assign \new_[34625]_  = \new_[34624]_  & \new_[34621]_ ;
  assign \new_[34626]_  = \new_[34625]_  & \new_[34618]_ ;
  assign \new_[34630]_  = ~A201 & A166;
  assign \new_[34631]_  = A168 & \new_[34630]_ ;
  assign \new_[34634]_  = ~A203 & ~A202;
  assign \new_[34637]_  = ~A233 & ~A232;
  assign \new_[34638]_  = \new_[34637]_  & \new_[34634]_ ;
  assign \new_[34639]_  = \new_[34638]_  & \new_[34631]_ ;
  assign \new_[34643]_  = ~A268 & ~A267;
  assign \new_[34644]_  = ~A235 & \new_[34643]_ ;
  assign \new_[34647]_  = ~A298 & ~A269;
  assign \new_[34650]_  = ~A301 & ~A299;
  assign \new_[34651]_  = \new_[34650]_  & \new_[34647]_ ;
  assign \new_[34652]_  = \new_[34651]_  & \new_[34644]_ ;
  assign \new_[34656]_  = ~A201 & A166;
  assign \new_[34657]_  = A168 & \new_[34656]_ ;
  assign \new_[34660]_  = ~A203 & ~A202;
  assign \new_[34663]_  = ~A233 & ~A232;
  assign \new_[34664]_  = \new_[34663]_  & \new_[34660]_ ;
  assign \new_[34665]_  = \new_[34664]_  & \new_[34657]_ ;
  assign \new_[34669]_  = ~A266 & ~A265;
  assign \new_[34670]_  = ~A235 & \new_[34669]_ ;
  assign \new_[34673]_  = ~A300 & ~A268;
  assign \new_[34676]_  = ~A302 & ~A301;
  assign \new_[34677]_  = \new_[34676]_  & \new_[34673]_ ;
  assign \new_[34678]_  = \new_[34677]_  & \new_[34670]_ ;
  assign \new_[34682]_  = ~A201 & A166;
  assign \new_[34683]_  = A168 & \new_[34682]_ ;
  assign \new_[34686]_  = ~A203 & ~A202;
  assign \new_[34689]_  = ~A233 & ~A232;
  assign \new_[34690]_  = \new_[34689]_  & \new_[34686]_ ;
  assign \new_[34691]_  = \new_[34690]_  & \new_[34683]_ ;
  assign \new_[34695]_  = ~A266 & ~A265;
  assign \new_[34696]_  = ~A235 & \new_[34695]_ ;
  assign \new_[34699]_  = ~A298 & ~A268;
  assign \new_[34702]_  = ~A301 & ~A299;
  assign \new_[34703]_  = \new_[34702]_  & \new_[34699]_ ;
  assign \new_[34704]_  = \new_[34703]_  & \new_[34696]_ ;
  assign \new_[34708]_  = ~A199 & A166;
  assign \new_[34709]_  = A168 & \new_[34708]_ ;
  assign \new_[34712]_  = ~A202 & ~A200;
  assign \new_[34715]_  = ~A235 & ~A234;
  assign \new_[34716]_  = \new_[34715]_  & \new_[34712]_ ;
  assign \new_[34717]_  = \new_[34716]_  & \new_[34709]_ ;
  assign \new_[34721]_  = ~A268 & ~A267;
  assign \new_[34722]_  = ~A236 & \new_[34721]_ ;
  assign \new_[34725]_  = ~A300 & ~A269;
  assign \new_[34728]_  = ~A302 & ~A301;
  assign \new_[34729]_  = \new_[34728]_  & \new_[34725]_ ;
  assign \new_[34730]_  = \new_[34729]_  & \new_[34722]_ ;
  assign \new_[34734]_  = ~A199 & A166;
  assign \new_[34735]_  = A168 & \new_[34734]_ ;
  assign \new_[34738]_  = ~A202 & ~A200;
  assign \new_[34741]_  = ~A235 & ~A234;
  assign \new_[34742]_  = \new_[34741]_  & \new_[34738]_ ;
  assign \new_[34743]_  = \new_[34742]_  & \new_[34735]_ ;
  assign \new_[34747]_  = ~A268 & ~A267;
  assign \new_[34748]_  = ~A236 & \new_[34747]_ ;
  assign \new_[34751]_  = ~A298 & ~A269;
  assign \new_[34754]_  = ~A301 & ~A299;
  assign \new_[34755]_  = \new_[34754]_  & \new_[34751]_ ;
  assign \new_[34756]_  = \new_[34755]_  & \new_[34748]_ ;
  assign \new_[34760]_  = ~A199 & A166;
  assign \new_[34761]_  = A168 & \new_[34760]_ ;
  assign \new_[34764]_  = ~A202 & ~A200;
  assign \new_[34767]_  = ~A235 & ~A234;
  assign \new_[34768]_  = \new_[34767]_  & \new_[34764]_ ;
  assign \new_[34769]_  = \new_[34768]_  & \new_[34761]_ ;
  assign \new_[34773]_  = ~A266 & ~A265;
  assign \new_[34774]_  = ~A236 & \new_[34773]_ ;
  assign \new_[34777]_  = ~A300 & ~A268;
  assign \new_[34780]_  = ~A302 & ~A301;
  assign \new_[34781]_  = \new_[34780]_  & \new_[34777]_ ;
  assign \new_[34782]_  = \new_[34781]_  & \new_[34774]_ ;
  assign \new_[34786]_  = ~A199 & A166;
  assign \new_[34787]_  = A168 & \new_[34786]_ ;
  assign \new_[34790]_  = ~A202 & ~A200;
  assign \new_[34793]_  = ~A235 & ~A234;
  assign \new_[34794]_  = \new_[34793]_  & \new_[34790]_ ;
  assign \new_[34795]_  = \new_[34794]_  & \new_[34787]_ ;
  assign \new_[34799]_  = ~A266 & ~A265;
  assign \new_[34800]_  = ~A236 & \new_[34799]_ ;
  assign \new_[34803]_  = ~A298 & ~A268;
  assign \new_[34806]_  = ~A301 & ~A299;
  assign \new_[34807]_  = \new_[34806]_  & \new_[34803]_ ;
  assign \new_[34808]_  = \new_[34807]_  & \new_[34800]_ ;
  assign \new_[34812]_  = ~A199 & A166;
  assign \new_[34813]_  = A168 & \new_[34812]_ ;
  assign \new_[34816]_  = ~A202 & ~A200;
  assign \new_[34819]_  = ~A233 & ~A232;
  assign \new_[34820]_  = \new_[34819]_  & \new_[34816]_ ;
  assign \new_[34821]_  = \new_[34820]_  & \new_[34813]_ ;
  assign \new_[34825]_  = ~A268 & ~A267;
  assign \new_[34826]_  = ~A235 & \new_[34825]_ ;
  assign \new_[34829]_  = ~A300 & ~A269;
  assign \new_[34832]_  = ~A302 & ~A301;
  assign \new_[34833]_  = \new_[34832]_  & \new_[34829]_ ;
  assign \new_[34834]_  = \new_[34833]_  & \new_[34826]_ ;
  assign \new_[34838]_  = ~A199 & A166;
  assign \new_[34839]_  = A168 & \new_[34838]_ ;
  assign \new_[34842]_  = ~A202 & ~A200;
  assign \new_[34845]_  = ~A233 & ~A232;
  assign \new_[34846]_  = \new_[34845]_  & \new_[34842]_ ;
  assign \new_[34847]_  = \new_[34846]_  & \new_[34839]_ ;
  assign \new_[34851]_  = ~A268 & ~A267;
  assign \new_[34852]_  = ~A235 & \new_[34851]_ ;
  assign \new_[34855]_  = ~A298 & ~A269;
  assign \new_[34858]_  = ~A301 & ~A299;
  assign \new_[34859]_  = \new_[34858]_  & \new_[34855]_ ;
  assign \new_[34860]_  = \new_[34859]_  & \new_[34852]_ ;
  assign \new_[34864]_  = ~A199 & A166;
  assign \new_[34865]_  = A168 & \new_[34864]_ ;
  assign \new_[34868]_  = ~A202 & ~A200;
  assign \new_[34871]_  = ~A233 & ~A232;
  assign \new_[34872]_  = \new_[34871]_  & \new_[34868]_ ;
  assign \new_[34873]_  = \new_[34872]_  & \new_[34865]_ ;
  assign \new_[34877]_  = ~A266 & ~A265;
  assign \new_[34878]_  = ~A235 & \new_[34877]_ ;
  assign \new_[34881]_  = ~A300 & ~A268;
  assign \new_[34884]_  = ~A302 & ~A301;
  assign \new_[34885]_  = \new_[34884]_  & \new_[34881]_ ;
  assign \new_[34886]_  = \new_[34885]_  & \new_[34878]_ ;
  assign \new_[34890]_  = ~A199 & A166;
  assign \new_[34891]_  = A168 & \new_[34890]_ ;
  assign \new_[34894]_  = ~A202 & ~A200;
  assign \new_[34897]_  = ~A233 & ~A232;
  assign \new_[34898]_  = \new_[34897]_  & \new_[34894]_ ;
  assign \new_[34899]_  = \new_[34898]_  & \new_[34891]_ ;
  assign \new_[34903]_  = ~A266 & ~A265;
  assign \new_[34904]_  = ~A235 & \new_[34903]_ ;
  assign \new_[34907]_  = ~A298 & ~A268;
  assign \new_[34910]_  = ~A301 & ~A299;
  assign \new_[34911]_  = \new_[34910]_  & \new_[34907]_ ;
  assign \new_[34912]_  = \new_[34911]_  & \new_[34904]_ ;
  assign \new_[34916]_  = ~A201 & A167;
  assign \new_[34917]_  = A168 & \new_[34916]_ ;
  assign \new_[34920]_  = ~A203 & ~A202;
  assign \new_[34923]_  = ~A235 & ~A234;
  assign \new_[34924]_  = \new_[34923]_  & \new_[34920]_ ;
  assign \new_[34925]_  = \new_[34924]_  & \new_[34917]_ ;
  assign \new_[34929]_  = ~A268 & ~A267;
  assign \new_[34930]_  = ~A236 & \new_[34929]_ ;
  assign \new_[34933]_  = ~A300 & ~A269;
  assign \new_[34936]_  = ~A302 & ~A301;
  assign \new_[34937]_  = \new_[34936]_  & \new_[34933]_ ;
  assign \new_[34938]_  = \new_[34937]_  & \new_[34930]_ ;
  assign \new_[34942]_  = ~A201 & A167;
  assign \new_[34943]_  = A168 & \new_[34942]_ ;
  assign \new_[34946]_  = ~A203 & ~A202;
  assign \new_[34949]_  = ~A235 & ~A234;
  assign \new_[34950]_  = \new_[34949]_  & \new_[34946]_ ;
  assign \new_[34951]_  = \new_[34950]_  & \new_[34943]_ ;
  assign \new_[34955]_  = ~A268 & ~A267;
  assign \new_[34956]_  = ~A236 & \new_[34955]_ ;
  assign \new_[34959]_  = ~A298 & ~A269;
  assign \new_[34962]_  = ~A301 & ~A299;
  assign \new_[34963]_  = \new_[34962]_  & \new_[34959]_ ;
  assign \new_[34964]_  = \new_[34963]_  & \new_[34956]_ ;
  assign \new_[34968]_  = ~A201 & A167;
  assign \new_[34969]_  = A168 & \new_[34968]_ ;
  assign \new_[34972]_  = ~A203 & ~A202;
  assign \new_[34975]_  = ~A235 & ~A234;
  assign \new_[34976]_  = \new_[34975]_  & \new_[34972]_ ;
  assign \new_[34977]_  = \new_[34976]_  & \new_[34969]_ ;
  assign \new_[34981]_  = ~A266 & ~A265;
  assign \new_[34982]_  = ~A236 & \new_[34981]_ ;
  assign \new_[34985]_  = ~A300 & ~A268;
  assign \new_[34988]_  = ~A302 & ~A301;
  assign \new_[34989]_  = \new_[34988]_  & \new_[34985]_ ;
  assign \new_[34990]_  = \new_[34989]_  & \new_[34982]_ ;
  assign \new_[34994]_  = ~A201 & A167;
  assign \new_[34995]_  = A168 & \new_[34994]_ ;
  assign \new_[34998]_  = ~A203 & ~A202;
  assign \new_[35001]_  = ~A235 & ~A234;
  assign \new_[35002]_  = \new_[35001]_  & \new_[34998]_ ;
  assign \new_[35003]_  = \new_[35002]_  & \new_[34995]_ ;
  assign \new_[35007]_  = ~A266 & ~A265;
  assign \new_[35008]_  = ~A236 & \new_[35007]_ ;
  assign \new_[35011]_  = ~A298 & ~A268;
  assign \new_[35014]_  = ~A301 & ~A299;
  assign \new_[35015]_  = \new_[35014]_  & \new_[35011]_ ;
  assign \new_[35016]_  = \new_[35015]_  & \new_[35008]_ ;
  assign \new_[35020]_  = ~A201 & A167;
  assign \new_[35021]_  = A168 & \new_[35020]_ ;
  assign \new_[35024]_  = ~A203 & ~A202;
  assign \new_[35027]_  = ~A233 & ~A232;
  assign \new_[35028]_  = \new_[35027]_  & \new_[35024]_ ;
  assign \new_[35029]_  = \new_[35028]_  & \new_[35021]_ ;
  assign \new_[35033]_  = ~A268 & ~A267;
  assign \new_[35034]_  = ~A235 & \new_[35033]_ ;
  assign \new_[35037]_  = ~A300 & ~A269;
  assign \new_[35040]_  = ~A302 & ~A301;
  assign \new_[35041]_  = \new_[35040]_  & \new_[35037]_ ;
  assign \new_[35042]_  = \new_[35041]_  & \new_[35034]_ ;
  assign \new_[35046]_  = ~A201 & A167;
  assign \new_[35047]_  = A168 & \new_[35046]_ ;
  assign \new_[35050]_  = ~A203 & ~A202;
  assign \new_[35053]_  = ~A233 & ~A232;
  assign \new_[35054]_  = \new_[35053]_  & \new_[35050]_ ;
  assign \new_[35055]_  = \new_[35054]_  & \new_[35047]_ ;
  assign \new_[35059]_  = ~A268 & ~A267;
  assign \new_[35060]_  = ~A235 & \new_[35059]_ ;
  assign \new_[35063]_  = ~A298 & ~A269;
  assign \new_[35066]_  = ~A301 & ~A299;
  assign \new_[35067]_  = \new_[35066]_  & \new_[35063]_ ;
  assign \new_[35068]_  = \new_[35067]_  & \new_[35060]_ ;
  assign \new_[35072]_  = ~A201 & A167;
  assign \new_[35073]_  = A168 & \new_[35072]_ ;
  assign \new_[35076]_  = ~A203 & ~A202;
  assign \new_[35079]_  = ~A233 & ~A232;
  assign \new_[35080]_  = \new_[35079]_  & \new_[35076]_ ;
  assign \new_[35081]_  = \new_[35080]_  & \new_[35073]_ ;
  assign \new_[35085]_  = ~A266 & ~A265;
  assign \new_[35086]_  = ~A235 & \new_[35085]_ ;
  assign \new_[35089]_  = ~A300 & ~A268;
  assign \new_[35092]_  = ~A302 & ~A301;
  assign \new_[35093]_  = \new_[35092]_  & \new_[35089]_ ;
  assign \new_[35094]_  = \new_[35093]_  & \new_[35086]_ ;
  assign \new_[35098]_  = ~A201 & A167;
  assign \new_[35099]_  = A168 & \new_[35098]_ ;
  assign \new_[35102]_  = ~A203 & ~A202;
  assign \new_[35105]_  = ~A233 & ~A232;
  assign \new_[35106]_  = \new_[35105]_  & \new_[35102]_ ;
  assign \new_[35107]_  = \new_[35106]_  & \new_[35099]_ ;
  assign \new_[35111]_  = ~A266 & ~A265;
  assign \new_[35112]_  = ~A235 & \new_[35111]_ ;
  assign \new_[35115]_  = ~A298 & ~A268;
  assign \new_[35118]_  = ~A301 & ~A299;
  assign \new_[35119]_  = \new_[35118]_  & \new_[35115]_ ;
  assign \new_[35120]_  = \new_[35119]_  & \new_[35112]_ ;
  assign \new_[35124]_  = ~A199 & A167;
  assign \new_[35125]_  = A168 & \new_[35124]_ ;
  assign \new_[35128]_  = ~A202 & ~A200;
  assign \new_[35131]_  = ~A235 & ~A234;
  assign \new_[35132]_  = \new_[35131]_  & \new_[35128]_ ;
  assign \new_[35133]_  = \new_[35132]_  & \new_[35125]_ ;
  assign \new_[35137]_  = ~A268 & ~A267;
  assign \new_[35138]_  = ~A236 & \new_[35137]_ ;
  assign \new_[35141]_  = ~A300 & ~A269;
  assign \new_[35144]_  = ~A302 & ~A301;
  assign \new_[35145]_  = \new_[35144]_  & \new_[35141]_ ;
  assign \new_[35146]_  = \new_[35145]_  & \new_[35138]_ ;
  assign \new_[35150]_  = ~A199 & A167;
  assign \new_[35151]_  = A168 & \new_[35150]_ ;
  assign \new_[35154]_  = ~A202 & ~A200;
  assign \new_[35157]_  = ~A235 & ~A234;
  assign \new_[35158]_  = \new_[35157]_  & \new_[35154]_ ;
  assign \new_[35159]_  = \new_[35158]_  & \new_[35151]_ ;
  assign \new_[35163]_  = ~A268 & ~A267;
  assign \new_[35164]_  = ~A236 & \new_[35163]_ ;
  assign \new_[35167]_  = ~A298 & ~A269;
  assign \new_[35170]_  = ~A301 & ~A299;
  assign \new_[35171]_  = \new_[35170]_  & \new_[35167]_ ;
  assign \new_[35172]_  = \new_[35171]_  & \new_[35164]_ ;
  assign \new_[35176]_  = ~A199 & A167;
  assign \new_[35177]_  = A168 & \new_[35176]_ ;
  assign \new_[35180]_  = ~A202 & ~A200;
  assign \new_[35183]_  = ~A235 & ~A234;
  assign \new_[35184]_  = \new_[35183]_  & \new_[35180]_ ;
  assign \new_[35185]_  = \new_[35184]_  & \new_[35177]_ ;
  assign \new_[35189]_  = ~A266 & ~A265;
  assign \new_[35190]_  = ~A236 & \new_[35189]_ ;
  assign \new_[35193]_  = ~A300 & ~A268;
  assign \new_[35196]_  = ~A302 & ~A301;
  assign \new_[35197]_  = \new_[35196]_  & \new_[35193]_ ;
  assign \new_[35198]_  = \new_[35197]_  & \new_[35190]_ ;
  assign \new_[35202]_  = ~A199 & A167;
  assign \new_[35203]_  = A168 & \new_[35202]_ ;
  assign \new_[35206]_  = ~A202 & ~A200;
  assign \new_[35209]_  = ~A235 & ~A234;
  assign \new_[35210]_  = \new_[35209]_  & \new_[35206]_ ;
  assign \new_[35211]_  = \new_[35210]_  & \new_[35203]_ ;
  assign \new_[35215]_  = ~A266 & ~A265;
  assign \new_[35216]_  = ~A236 & \new_[35215]_ ;
  assign \new_[35219]_  = ~A298 & ~A268;
  assign \new_[35222]_  = ~A301 & ~A299;
  assign \new_[35223]_  = \new_[35222]_  & \new_[35219]_ ;
  assign \new_[35224]_  = \new_[35223]_  & \new_[35216]_ ;
  assign \new_[35228]_  = ~A199 & A167;
  assign \new_[35229]_  = A168 & \new_[35228]_ ;
  assign \new_[35232]_  = ~A202 & ~A200;
  assign \new_[35235]_  = ~A233 & ~A232;
  assign \new_[35236]_  = \new_[35235]_  & \new_[35232]_ ;
  assign \new_[35237]_  = \new_[35236]_  & \new_[35229]_ ;
  assign \new_[35241]_  = ~A268 & ~A267;
  assign \new_[35242]_  = ~A235 & \new_[35241]_ ;
  assign \new_[35245]_  = ~A300 & ~A269;
  assign \new_[35248]_  = ~A302 & ~A301;
  assign \new_[35249]_  = \new_[35248]_  & \new_[35245]_ ;
  assign \new_[35250]_  = \new_[35249]_  & \new_[35242]_ ;
  assign \new_[35254]_  = ~A199 & A167;
  assign \new_[35255]_  = A168 & \new_[35254]_ ;
  assign \new_[35258]_  = ~A202 & ~A200;
  assign \new_[35261]_  = ~A233 & ~A232;
  assign \new_[35262]_  = \new_[35261]_  & \new_[35258]_ ;
  assign \new_[35263]_  = \new_[35262]_  & \new_[35255]_ ;
  assign \new_[35267]_  = ~A268 & ~A267;
  assign \new_[35268]_  = ~A235 & \new_[35267]_ ;
  assign \new_[35271]_  = ~A298 & ~A269;
  assign \new_[35274]_  = ~A301 & ~A299;
  assign \new_[35275]_  = \new_[35274]_  & \new_[35271]_ ;
  assign \new_[35276]_  = \new_[35275]_  & \new_[35268]_ ;
  assign \new_[35280]_  = ~A199 & A167;
  assign \new_[35281]_  = A168 & \new_[35280]_ ;
  assign \new_[35284]_  = ~A202 & ~A200;
  assign \new_[35287]_  = ~A233 & ~A232;
  assign \new_[35288]_  = \new_[35287]_  & \new_[35284]_ ;
  assign \new_[35289]_  = \new_[35288]_  & \new_[35281]_ ;
  assign \new_[35293]_  = ~A266 & ~A265;
  assign \new_[35294]_  = ~A235 & \new_[35293]_ ;
  assign \new_[35297]_  = ~A300 & ~A268;
  assign \new_[35300]_  = ~A302 & ~A301;
  assign \new_[35301]_  = \new_[35300]_  & \new_[35297]_ ;
  assign \new_[35302]_  = \new_[35301]_  & \new_[35294]_ ;
  assign \new_[35306]_  = ~A199 & A167;
  assign \new_[35307]_  = A168 & \new_[35306]_ ;
  assign \new_[35310]_  = ~A202 & ~A200;
  assign \new_[35313]_  = ~A233 & ~A232;
  assign \new_[35314]_  = \new_[35313]_  & \new_[35310]_ ;
  assign \new_[35315]_  = \new_[35314]_  & \new_[35307]_ ;
  assign \new_[35319]_  = ~A266 & ~A265;
  assign \new_[35320]_  = ~A235 & \new_[35319]_ ;
  assign \new_[35323]_  = ~A298 & ~A268;
  assign \new_[35326]_  = ~A301 & ~A299;
  assign \new_[35327]_  = \new_[35326]_  & \new_[35323]_ ;
  assign \new_[35328]_  = \new_[35327]_  & \new_[35320]_ ;
  assign \new_[35332]_  = ~A202 & ~A201;
  assign \new_[35333]_  = A169 & \new_[35332]_ ;
  assign \new_[35336]_  = ~A234 & ~A203;
  assign \new_[35339]_  = ~A236 & ~A235;
  assign \new_[35340]_  = \new_[35339]_  & \new_[35336]_ ;
  assign \new_[35341]_  = \new_[35340]_  & \new_[35333]_ ;
  assign \new_[35345]_  = ~A269 & ~A268;
  assign \new_[35346]_  = ~A267 & \new_[35345]_ ;
  assign \new_[35349]_  = A299 & A298;
  assign \new_[35352]_  = ~A301 & ~A300;
  assign \new_[35353]_  = \new_[35352]_  & \new_[35349]_ ;
  assign \new_[35354]_  = \new_[35353]_  & \new_[35346]_ ;
  assign \new_[35358]_  = ~A202 & ~A201;
  assign \new_[35359]_  = A169 & \new_[35358]_ ;
  assign \new_[35362]_  = ~A234 & ~A203;
  assign \new_[35365]_  = ~A236 & ~A235;
  assign \new_[35366]_  = \new_[35365]_  & \new_[35362]_ ;
  assign \new_[35367]_  = \new_[35366]_  & \new_[35359]_ ;
  assign \new_[35371]_  = ~A267 & A266;
  assign \new_[35372]_  = A265 & \new_[35371]_ ;
  assign \new_[35375]_  = ~A300 & ~A268;
  assign \new_[35378]_  = ~A302 & ~A301;
  assign \new_[35379]_  = \new_[35378]_  & \new_[35375]_ ;
  assign \new_[35380]_  = \new_[35379]_  & \new_[35372]_ ;
  assign \new_[35384]_  = ~A202 & ~A201;
  assign \new_[35385]_  = A169 & \new_[35384]_ ;
  assign \new_[35388]_  = ~A234 & ~A203;
  assign \new_[35391]_  = ~A236 & ~A235;
  assign \new_[35392]_  = \new_[35391]_  & \new_[35388]_ ;
  assign \new_[35393]_  = \new_[35392]_  & \new_[35385]_ ;
  assign \new_[35397]_  = ~A267 & A266;
  assign \new_[35398]_  = A265 & \new_[35397]_ ;
  assign \new_[35401]_  = ~A298 & ~A268;
  assign \new_[35404]_  = ~A301 & ~A299;
  assign \new_[35405]_  = \new_[35404]_  & \new_[35401]_ ;
  assign \new_[35406]_  = \new_[35405]_  & \new_[35398]_ ;
  assign \new_[35410]_  = ~A202 & ~A201;
  assign \new_[35411]_  = A169 & \new_[35410]_ ;
  assign \new_[35414]_  = ~A234 & ~A203;
  assign \new_[35417]_  = ~A236 & ~A235;
  assign \new_[35418]_  = \new_[35417]_  & \new_[35414]_ ;
  assign \new_[35419]_  = \new_[35418]_  & \new_[35411]_ ;
  assign \new_[35423]_  = ~A268 & ~A266;
  assign \new_[35424]_  = ~A265 & \new_[35423]_ ;
  assign \new_[35427]_  = A299 & A298;
  assign \new_[35430]_  = ~A301 & ~A300;
  assign \new_[35431]_  = \new_[35430]_  & \new_[35427]_ ;
  assign \new_[35432]_  = \new_[35431]_  & \new_[35424]_ ;
  assign \new_[35436]_  = ~A202 & ~A201;
  assign \new_[35437]_  = A169 & \new_[35436]_ ;
  assign \new_[35440]_  = A232 & ~A203;
  assign \new_[35443]_  = ~A234 & A233;
  assign \new_[35444]_  = \new_[35443]_  & \new_[35440]_ ;
  assign \new_[35445]_  = \new_[35444]_  & \new_[35437]_ ;
  assign \new_[35449]_  = ~A268 & ~A267;
  assign \new_[35450]_  = ~A235 & \new_[35449]_ ;
  assign \new_[35453]_  = ~A300 & ~A269;
  assign \new_[35456]_  = ~A302 & ~A301;
  assign \new_[35457]_  = \new_[35456]_  & \new_[35453]_ ;
  assign \new_[35458]_  = \new_[35457]_  & \new_[35450]_ ;
  assign \new_[35462]_  = ~A202 & ~A201;
  assign \new_[35463]_  = A169 & \new_[35462]_ ;
  assign \new_[35466]_  = A232 & ~A203;
  assign \new_[35469]_  = ~A234 & A233;
  assign \new_[35470]_  = \new_[35469]_  & \new_[35466]_ ;
  assign \new_[35471]_  = \new_[35470]_  & \new_[35463]_ ;
  assign \new_[35475]_  = ~A268 & ~A267;
  assign \new_[35476]_  = ~A235 & \new_[35475]_ ;
  assign \new_[35479]_  = ~A298 & ~A269;
  assign \new_[35482]_  = ~A301 & ~A299;
  assign \new_[35483]_  = \new_[35482]_  & \new_[35479]_ ;
  assign \new_[35484]_  = \new_[35483]_  & \new_[35476]_ ;
  assign \new_[35488]_  = ~A202 & ~A201;
  assign \new_[35489]_  = A169 & \new_[35488]_ ;
  assign \new_[35492]_  = A232 & ~A203;
  assign \new_[35495]_  = ~A234 & A233;
  assign \new_[35496]_  = \new_[35495]_  & \new_[35492]_ ;
  assign \new_[35497]_  = \new_[35496]_  & \new_[35489]_ ;
  assign \new_[35501]_  = ~A266 & ~A265;
  assign \new_[35502]_  = ~A235 & \new_[35501]_ ;
  assign \new_[35505]_  = ~A300 & ~A268;
  assign \new_[35508]_  = ~A302 & ~A301;
  assign \new_[35509]_  = \new_[35508]_  & \new_[35505]_ ;
  assign \new_[35510]_  = \new_[35509]_  & \new_[35502]_ ;
  assign \new_[35514]_  = ~A202 & ~A201;
  assign \new_[35515]_  = A169 & \new_[35514]_ ;
  assign \new_[35518]_  = A232 & ~A203;
  assign \new_[35521]_  = ~A234 & A233;
  assign \new_[35522]_  = \new_[35521]_  & \new_[35518]_ ;
  assign \new_[35523]_  = \new_[35522]_  & \new_[35515]_ ;
  assign \new_[35527]_  = ~A266 & ~A265;
  assign \new_[35528]_  = ~A235 & \new_[35527]_ ;
  assign \new_[35531]_  = ~A298 & ~A268;
  assign \new_[35534]_  = ~A301 & ~A299;
  assign \new_[35535]_  = \new_[35534]_  & \new_[35531]_ ;
  assign \new_[35536]_  = \new_[35535]_  & \new_[35528]_ ;
  assign \new_[35540]_  = ~A202 & ~A201;
  assign \new_[35541]_  = A169 & \new_[35540]_ ;
  assign \new_[35544]_  = ~A232 & ~A203;
  assign \new_[35547]_  = ~A235 & ~A233;
  assign \new_[35548]_  = \new_[35547]_  & \new_[35544]_ ;
  assign \new_[35549]_  = \new_[35548]_  & \new_[35541]_ ;
  assign \new_[35553]_  = ~A269 & ~A268;
  assign \new_[35554]_  = ~A267 & \new_[35553]_ ;
  assign \new_[35557]_  = A299 & A298;
  assign \new_[35560]_  = ~A301 & ~A300;
  assign \new_[35561]_  = \new_[35560]_  & \new_[35557]_ ;
  assign \new_[35562]_  = \new_[35561]_  & \new_[35554]_ ;
  assign \new_[35566]_  = ~A202 & ~A201;
  assign \new_[35567]_  = A169 & \new_[35566]_ ;
  assign \new_[35570]_  = ~A232 & ~A203;
  assign \new_[35573]_  = ~A235 & ~A233;
  assign \new_[35574]_  = \new_[35573]_  & \new_[35570]_ ;
  assign \new_[35575]_  = \new_[35574]_  & \new_[35567]_ ;
  assign \new_[35579]_  = ~A267 & A266;
  assign \new_[35580]_  = A265 & \new_[35579]_ ;
  assign \new_[35583]_  = ~A300 & ~A268;
  assign \new_[35586]_  = ~A302 & ~A301;
  assign \new_[35587]_  = \new_[35586]_  & \new_[35583]_ ;
  assign \new_[35588]_  = \new_[35587]_  & \new_[35580]_ ;
  assign \new_[35592]_  = ~A202 & ~A201;
  assign \new_[35593]_  = A169 & \new_[35592]_ ;
  assign \new_[35596]_  = ~A232 & ~A203;
  assign \new_[35599]_  = ~A235 & ~A233;
  assign \new_[35600]_  = \new_[35599]_  & \new_[35596]_ ;
  assign \new_[35601]_  = \new_[35600]_  & \new_[35593]_ ;
  assign \new_[35605]_  = ~A267 & A266;
  assign \new_[35606]_  = A265 & \new_[35605]_ ;
  assign \new_[35609]_  = ~A298 & ~A268;
  assign \new_[35612]_  = ~A301 & ~A299;
  assign \new_[35613]_  = \new_[35612]_  & \new_[35609]_ ;
  assign \new_[35614]_  = \new_[35613]_  & \new_[35606]_ ;
  assign \new_[35618]_  = ~A202 & ~A201;
  assign \new_[35619]_  = A169 & \new_[35618]_ ;
  assign \new_[35622]_  = ~A232 & ~A203;
  assign \new_[35625]_  = ~A235 & ~A233;
  assign \new_[35626]_  = \new_[35625]_  & \new_[35622]_ ;
  assign \new_[35627]_  = \new_[35626]_  & \new_[35619]_ ;
  assign \new_[35631]_  = ~A268 & ~A266;
  assign \new_[35632]_  = ~A265 & \new_[35631]_ ;
  assign \new_[35635]_  = A299 & A298;
  assign \new_[35638]_  = ~A301 & ~A300;
  assign \new_[35639]_  = \new_[35638]_  & \new_[35635]_ ;
  assign \new_[35640]_  = \new_[35639]_  & \new_[35632]_ ;
  assign \new_[35644]_  = A200 & A199;
  assign \new_[35645]_  = A169 & \new_[35644]_ ;
  assign \new_[35648]_  = ~A202 & ~A201;
  assign \new_[35651]_  = ~A235 & ~A234;
  assign \new_[35652]_  = \new_[35651]_  & \new_[35648]_ ;
  assign \new_[35653]_  = \new_[35652]_  & \new_[35645]_ ;
  assign \new_[35657]_  = ~A268 & ~A267;
  assign \new_[35658]_  = ~A236 & \new_[35657]_ ;
  assign \new_[35661]_  = ~A300 & ~A269;
  assign \new_[35664]_  = ~A302 & ~A301;
  assign \new_[35665]_  = \new_[35664]_  & \new_[35661]_ ;
  assign \new_[35666]_  = \new_[35665]_  & \new_[35658]_ ;
  assign \new_[35670]_  = A200 & A199;
  assign \new_[35671]_  = A169 & \new_[35670]_ ;
  assign \new_[35674]_  = ~A202 & ~A201;
  assign \new_[35677]_  = ~A235 & ~A234;
  assign \new_[35678]_  = \new_[35677]_  & \new_[35674]_ ;
  assign \new_[35679]_  = \new_[35678]_  & \new_[35671]_ ;
  assign \new_[35683]_  = ~A268 & ~A267;
  assign \new_[35684]_  = ~A236 & \new_[35683]_ ;
  assign \new_[35687]_  = ~A298 & ~A269;
  assign \new_[35690]_  = ~A301 & ~A299;
  assign \new_[35691]_  = \new_[35690]_  & \new_[35687]_ ;
  assign \new_[35692]_  = \new_[35691]_  & \new_[35684]_ ;
  assign \new_[35696]_  = A200 & A199;
  assign \new_[35697]_  = A169 & \new_[35696]_ ;
  assign \new_[35700]_  = ~A202 & ~A201;
  assign \new_[35703]_  = ~A235 & ~A234;
  assign \new_[35704]_  = \new_[35703]_  & \new_[35700]_ ;
  assign \new_[35705]_  = \new_[35704]_  & \new_[35697]_ ;
  assign \new_[35709]_  = ~A266 & ~A265;
  assign \new_[35710]_  = ~A236 & \new_[35709]_ ;
  assign \new_[35713]_  = ~A300 & ~A268;
  assign \new_[35716]_  = ~A302 & ~A301;
  assign \new_[35717]_  = \new_[35716]_  & \new_[35713]_ ;
  assign \new_[35718]_  = \new_[35717]_  & \new_[35710]_ ;
  assign \new_[35722]_  = A200 & A199;
  assign \new_[35723]_  = A169 & \new_[35722]_ ;
  assign \new_[35726]_  = ~A202 & ~A201;
  assign \new_[35729]_  = ~A235 & ~A234;
  assign \new_[35730]_  = \new_[35729]_  & \new_[35726]_ ;
  assign \new_[35731]_  = \new_[35730]_  & \new_[35723]_ ;
  assign \new_[35735]_  = ~A266 & ~A265;
  assign \new_[35736]_  = ~A236 & \new_[35735]_ ;
  assign \new_[35739]_  = ~A298 & ~A268;
  assign \new_[35742]_  = ~A301 & ~A299;
  assign \new_[35743]_  = \new_[35742]_  & \new_[35739]_ ;
  assign \new_[35744]_  = \new_[35743]_  & \new_[35736]_ ;
  assign \new_[35748]_  = A200 & A199;
  assign \new_[35749]_  = A169 & \new_[35748]_ ;
  assign \new_[35752]_  = ~A202 & ~A201;
  assign \new_[35755]_  = ~A233 & ~A232;
  assign \new_[35756]_  = \new_[35755]_  & \new_[35752]_ ;
  assign \new_[35757]_  = \new_[35756]_  & \new_[35749]_ ;
  assign \new_[35761]_  = ~A268 & ~A267;
  assign \new_[35762]_  = ~A235 & \new_[35761]_ ;
  assign \new_[35765]_  = ~A300 & ~A269;
  assign \new_[35768]_  = ~A302 & ~A301;
  assign \new_[35769]_  = \new_[35768]_  & \new_[35765]_ ;
  assign \new_[35770]_  = \new_[35769]_  & \new_[35762]_ ;
  assign \new_[35774]_  = A200 & A199;
  assign \new_[35775]_  = A169 & \new_[35774]_ ;
  assign \new_[35778]_  = ~A202 & ~A201;
  assign \new_[35781]_  = ~A233 & ~A232;
  assign \new_[35782]_  = \new_[35781]_  & \new_[35778]_ ;
  assign \new_[35783]_  = \new_[35782]_  & \new_[35775]_ ;
  assign \new_[35787]_  = ~A268 & ~A267;
  assign \new_[35788]_  = ~A235 & \new_[35787]_ ;
  assign \new_[35791]_  = ~A298 & ~A269;
  assign \new_[35794]_  = ~A301 & ~A299;
  assign \new_[35795]_  = \new_[35794]_  & \new_[35791]_ ;
  assign \new_[35796]_  = \new_[35795]_  & \new_[35788]_ ;
  assign \new_[35800]_  = A200 & A199;
  assign \new_[35801]_  = A169 & \new_[35800]_ ;
  assign \new_[35804]_  = ~A202 & ~A201;
  assign \new_[35807]_  = ~A233 & ~A232;
  assign \new_[35808]_  = \new_[35807]_  & \new_[35804]_ ;
  assign \new_[35809]_  = \new_[35808]_  & \new_[35801]_ ;
  assign \new_[35813]_  = ~A266 & ~A265;
  assign \new_[35814]_  = ~A235 & \new_[35813]_ ;
  assign \new_[35817]_  = ~A300 & ~A268;
  assign \new_[35820]_  = ~A302 & ~A301;
  assign \new_[35821]_  = \new_[35820]_  & \new_[35817]_ ;
  assign \new_[35822]_  = \new_[35821]_  & \new_[35814]_ ;
  assign \new_[35826]_  = A200 & A199;
  assign \new_[35827]_  = A169 & \new_[35826]_ ;
  assign \new_[35830]_  = ~A202 & ~A201;
  assign \new_[35833]_  = ~A233 & ~A232;
  assign \new_[35834]_  = \new_[35833]_  & \new_[35830]_ ;
  assign \new_[35835]_  = \new_[35834]_  & \new_[35827]_ ;
  assign \new_[35839]_  = ~A266 & ~A265;
  assign \new_[35840]_  = ~A235 & \new_[35839]_ ;
  assign \new_[35843]_  = ~A298 & ~A268;
  assign \new_[35846]_  = ~A301 & ~A299;
  assign \new_[35847]_  = \new_[35846]_  & \new_[35843]_ ;
  assign \new_[35848]_  = \new_[35847]_  & \new_[35840]_ ;
  assign \new_[35852]_  = ~A200 & ~A199;
  assign \new_[35853]_  = A169 & \new_[35852]_ ;
  assign \new_[35856]_  = ~A234 & ~A202;
  assign \new_[35859]_  = ~A236 & ~A235;
  assign \new_[35860]_  = \new_[35859]_  & \new_[35856]_ ;
  assign \new_[35861]_  = \new_[35860]_  & \new_[35853]_ ;
  assign \new_[35865]_  = ~A269 & ~A268;
  assign \new_[35866]_  = ~A267 & \new_[35865]_ ;
  assign \new_[35869]_  = A299 & A298;
  assign \new_[35872]_  = ~A301 & ~A300;
  assign \new_[35873]_  = \new_[35872]_  & \new_[35869]_ ;
  assign \new_[35874]_  = \new_[35873]_  & \new_[35866]_ ;
  assign \new_[35878]_  = ~A200 & ~A199;
  assign \new_[35879]_  = A169 & \new_[35878]_ ;
  assign \new_[35882]_  = ~A234 & ~A202;
  assign \new_[35885]_  = ~A236 & ~A235;
  assign \new_[35886]_  = \new_[35885]_  & \new_[35882]_ ;
  assign \new_[35887]_  = \new_[35886]_  & \new_[35879]_ ;
  assign \new_[35891]_  = ~A267 & A266;
  assign \new_[35892]_  = A265 & \new_[35891]_ ;
  assign \new_[35895]_  = ~A300 & ~A268;
  assign \new_[35898]_  = ~A302 & ~A301;
  assign \new_[35899]_  = \new_[35898]_  & \new_[35895]_ ;
  assign \new_[35900]_  = \new_[35899]_  & \new_[35892]_ ;
  assign \new_[35904]_  = ~A200 & ~A199;
  assign \new_[35905]_  = A169 & \new_[35904]_ ;
  assign \new_[35908]_  = ~A234 & ~A202;
  assign \new_[35911]_  = ~A236 & ~A235;
  assign \new_[35912]_  = \new_[35911]_  & \new_[35908]_ ;
  assign \new_[35913]_  = \new_[35912]_  & \new_[35905]_ ;
  assign \new_[35917]_  = ~A267 & A266;
  assign \new_[35918]_  = A265 & \new_[35917]_ ;
  assign \new_[35921]_  = ~A298 & ~A268;
  assign \new_[35924]_  = ~A301 & ~A299;
  assign \new_[35925]_  = \new_[35924]_  & \new_[35921]_ ;
  assign \new_[35926]_  = \new_[35925]_  & \new_[35918]_ ;
  assign \new_[35930]_  = ~A200 & ~A199;
  assign \new_[35931]_  = A169 & \new_[35930]_ ;
  assign \new_[35934]_  = ~A234 & ~A202;
  assign \new_[35937]_  = ~A236 & ~A235;
  assign \new_[35938]_  = \new_[35937]_  & \new_[35934]_ ;
  assign \new_[35939]_  = \new_[35938]_  & \new_[35931]_ ;
  assign \new_[35943]_  = ~A268 & ~A266;
  assign \new_[35944]_  = ~A265 & \new_[35943]_ ;
  assign \new_[35947]_  = A299 & A298;
  assign \new_[35950]_  = ~A301 & ~A300;
  assign \new_[35951]_  = \new_[35950]_  & \new_[35947]_ ;
  assign \new_[35952]_  = \new_[35951]_  & \new_[35944]_ ;
  assign \new_[35956]_  = ~A200 & ~A199;
  assign \new_[35957]_  = A169 & \new_[35956]_ ;
  assign \new_[35960]_  = A232 & ~A202;
  assign \new_[35963]_  = ~A234 & A233;
  assign \new_[35964]_  = \new_[35963]_  & \new_[35960]_ ;
  assign \new_[35965]_  = \new_[35964]_  & \new_[35957]_ ;
  assign \new_[35969]_  = ~A268 & ~A267;
  assign \new_[35970]_  = ~A235 & \new_[35969]_ ;
  assign \new_[35973]_  = ~A300 & ~A269;
  assign \new_[35976]_  = ~A302 & ~A301;
  assign \new_[35977]_  = \new_[35976]_  & \new_[35973]_ ;
  assign \new_[35978]_  = \new_[35977]_  & \new_[35970]_ ;
  assign \new_[35982]_  = ~A200 & ~A199;
  assign \new_[35983]_  = A169 & \new_[35982]_ ;
  assign \new_[35986]_  = A232 & ~A202;
  assign \new_[35989]_  = ~A234 & A233;
  assign \new_[35990]_  = \new_[35989]_  & \new_[35986]_ ;
  assign \new_[35991]_  = \new_[35990]_  & \new_[35983]_ ;
  assign \new_[35995]_  = ~A268 & ~A267;
  assign \new_[35996]_  = ~A235 & \new_[35995]_ ;
  assign \new_[35999]_  = ~A298 & ~A269;
  assign \new_[36002]_  = ~A301 & ~A299;
  assign \new_[36003]_  = \new_[36002]_  & \new_[35999]_ ;
  assign \new_[36004]_  = \new_[36003]_  & \new_[35996]_ ;
  assign \new_[36008]_  = ~A200 & ~A199;
  assign \new_[36009]_  = A169 & \new_[36008]_ ;
  assign \new_[36012]_  = A232 & ~A202;
  assign \new_[36015]_  = ~A234 & A233;
  assign \new_[36016]_  = \new_[36015]_  & \new_[36012]_ ;
  assign \new_[36017]_  = \new_[36016]_  & \new_[36009]_ ;
  assign \new_[36021]_  = ~A266 & ~A265;
  assign \new_[36022]_  = ~A235 & \new_[36021]_ ;
  assign \new_[36025]_  = ~A300 & ~A268;
  assign \new_[36028]_  = ~A302 & ~A301;
  assign \new_[36029]_  = \new_[36028]_  & \new_[36025]_ ;
  assign \new_[36030]_  = \new_[36029]_  & \new_[36022]_ ;
  assign \new_[36034]_  = ~A200 & ~A199;
  assign \new_[36035]_  = A169 & \new_[36034]_ ;
  assign \new_[36038]_  = A232 & ~A202;
  assign \new_[36041]_  = ~A234 & A233;
  assign \new_[36042]_  = \new_[36041]_  & \new_[36038]_ ;
  assign \new_[36043]_  = \new_[36042]_  & \new_[36035]_ ;
  assign \new_[36047]_  = ~A266 & ~A265;
  assign \new_[36048]_  = ~A235 & \new_[36047]_ ;
  assign \new_[36051]_  = ~A298 & ~A268;
  assign \new_[36054]_  = ~A301 & ~A299;
  assign \new_[36055]_  = \new_[36054]_  & \new_[36051]_ ;
  assign \new_[36056]_  = \new_[36055]_  & \new_[36048]_ ;
  assign \new_[36060]_  = ~A200 & ~A199;
  assign \new_[36061]_  = A169 & \new_[36060]_ ;
  assign \new_[36064]_  = ~A232 & ~A202;
  assign \new_[36067]_  = ~A235 & ~A233;
  assign \new_[36068]_  = \new_[36067]_  & \new_[36064]_ ;
  assign \new_[36069]_  = \new_[36068]_  & \new_[36061]_ ;
  assign \new_[36073]_  = ~A269 & ~A268;
  assign \new_[36074]_  = ~A267 & \new_[36073]_ ;
  assign \new_[36077]_  = A299 & A298;
  assign \new_[36080]_  = ~A301 & ~A300;
  assign \new_[36081]_  = \new_[36080]_  & \new_[36077]_ ;
  assign \new_[36082]_  = \new_[36081]_  & \new_[36074]_ ;
  assign \new_[36086]_  = ~A200 & ~A199;
  assign \new_[36087]_  = A169 & \new_[36086]_ ;
  assign \new_[36090]_  = ~A232 & ~A202;
  assign \new_[36093]_  = ~A235 & ~A233;
  assign \new_[36094]_  = \new_[36093]_  & \new_[36090]_ ;
  assign \new_[36095]_  = \new_[36094]_  & \new_[36087]_ ;
  assign \new_[36099]_  = ~A267 & A266;
  assign \new_[36100]_  = A265 & \new_[36099]_ ;
  assign \new_[36103]_  = ~A300 & ~A268;
  assign \new_[36106]_  = ~A302 & ~A301;
  assign \new_[36107]_  = \new_[36106]_  & \new_[36103]_ ;
  assign \new_[36108]_  = \new_[36107]_  & \new_[36100]_ ;
  assign \new_[36112]_  = ~A200 & ~A199;
  assign \new_[36113]_  = A169 & \new_[36112]_ ;
  assign \new_[36116]_  = ~A232 & ~A202;
  assign \new_[36119]_  = ~A235 & ~A233;
  assign \new_[36120]_  = \new_[36119]_  & \new_[36116]_ ;
  assign \new_[36121]_  = \new_[36120]_  & \new_[36113]_ ;
  assign \new_[36125]_  = ~A267 & A266;
  assign \new_[36126]_  = A265 & \new_[36125]_ ;
  assign \new_[36129]_  = ~A298 & ~A268;
  assign \new_[36132]_  = ~A301 & ~A299;
  assign \new_[36133]_  = \new_[36132]_  & \new_[36129]_ ;
  assign \new_[36134]_  = \new_[36133]_  & \new_[36126]_ ;
  assign \new_[36138]_  = ~A200 & ~A199;
  assign \new_[36139]_  = A169 & \new_[36138]_ ;
  assign \new_[36142]_  = ~A232 & ~A202;
  assign \new_[36145]_  = ~A235 & ~A233;
  assign \new_[36146]_  = \new_[36145]_  & \new_[36142]_ ;
  assign \new_[36147]_  = \new_[36146]_  & \new_[36139]_ ;
  assign \new_[36151]_  = ~A268 & ~A266;
  assign \new_[36152]_  = ~A265 & \new_[36151]_ ;
  assign \new_[36155]_  = A299 & A298;
  assign \new_[36158]_  = ~A301 & ~A300;
  assign \new_[36159]_  = \new_[36158]_  & \new_[36155]_ ;
  assign \new_[36160]_  = \new_[36159]_  & \new_[36152]_ ;
  assign \new_[36164]_  = ~A166 & ~A167;
  assign \new_[36165]_  = ~A169 & \new_[36164]_ ;
  assign \new_[36168]_  = ~A234 & A202;
  assign \new_[36171]_  = ~A236 & ~A235;
  assign \new_[36172]_  = \new_[36171]_  & \new_[36168]_ ;
  assign \new_[36173]_  = \new_[36172]_  & \new_[36165]_ ;
  assign \new_[36177]_  = ~A269 & ~A268;
  assign \new_[36178]_  = ~A267 & \new_[36177]_ ;
  assign \new_[36181]_  = A299 & A298;
  assign \new_[36184]_  = ~A301 & ~A300;
  assign \new_[36185]_  = \new_[36184]_  & \new_[36181]_ ;
  assign \new_[36186]_  = \new_[36185]_  & \new_[36178]_ ;
  assign \new_[36190]_  = ~A166 & ~A167;
  assign \new_[36191]_  = ~A169 & \new_[36190]_ ;
  assign \new_[36194]_  = ~A234 & A202;
  assign \new_[36197]_  = ~A236 & ~A235;
  assign \new_[36198]_  = \new_[36197]_  & \new_[36194]_ ;
  assign \new_[36199]_  = \new_[36198]_  & \new_[36191]_ ;
  assign \new_[36203]_  = ~A267 & A266;
  assign \new_[36204]_  = A265 & \new_[36203]_ ;
  assign \new_[36207]_  = ~A300 & ~A268;
  assign \new_[36210]_  = ~A302 & ~A301;
  assign \new_[36211]_  = \new_[36210]_  & \new_[36207]_ ;
  assign \new_[36212]_  = \new_[36211]_  & \new_[36204]_ ;
  assign \new_[36216]_  = ~A166 & ~A167;
  assign \new_[36217]_  = ~A169 & \new_[36216]_ ;
  assign \new_[36220]_  = ~A234 & A202;
  assign \new_[36223]_  = ~A236 & ~A235;
  assign \new_[36224]_  = \new_[36223]_  & \new_[36220]_ ;
  assign \new_[36225]_  = \new_[36224]_  & \new_[36217]_ ;
  assign \new_[36229]_  = ~A267 & A266;
  assign \new_[36230]_  = A265 & \new_[36229]_ ;
  assign \new_[36233]_  = ~A298 & ~A268;
  assign \new_[36236]_  = ~A301 & ~A299;
  assign \new_[36237]_  = \new_[36236]_  & \new_[36233]_ ;
  assign \new_[36238]_  = \new_[36237]_  & \new_[36230]_ ;
  assign \new_[36242]_  = ~A166 & ~A167;
  assign \new_[36243]_  = ~A169 & \new_[36242]_ ;
  assign \new_[36246]_  = ~A234 & A202;
  assign \new_[36249]_  = ~A236 & ~A235;
  assign \new_[36250]_  = \new_[36249]_  & \new_[36246]_ ;
  assign \new_[36251]_  = \new_[36250]_  & \new_[36243]_ ;
  assign \new_[36255]_  = ~A268 & ~A266;
  assign \new_[36256]_  = ~A265 & \new_[36255]_ ;
  assign \new_[36259]_  = A299 & A298;
  assign \new_[36262]_  = ~A301 & ~A300;
  assign \new_[36263]_  = \new_[36262]_  & \new_[36259]_ ;
  assign \new_[36264]_  = \new_[36263]_  & \new_[36256]_ ;
  assign \new_[36268]_  = ~A166 & ~A167;
  assign \new_[36269]_  = ~A169 & \new_[36268]_ ;
  assign \new_[36272]_  = A232 & A202;
  assign \new_[36275]_  = ~A234 & A233;
  assign \new_[36276]_  = \new_[36275]_  & \new_[36272]_ ;
  assign \new_[36277]_  = \new_[36276]_  & \new_[36269]_ ;
  assign \new_[36281]_  = ~A268 & ~A267;
  assign \new_[36282]_  = ~A235 & \new_[36281]_ ;
  assign \new_[36285]_  = ~A300 & ~A269;
  assign \new_[36288]_  = ~A302 & ~A301;
  assign \new_[36289]_  = \new_[36288]_  & \new_[36285]_ ;
  assign \new_[36290]_  = \new_[36289]_  & \new_[36282]_ ;
  assign \new_[36294]_  = ~A166 & ~A167;
  assign \new_[36295]_  = ~A169 & \new_[36294]_ ;
  assign \new_[36298]_  = A232 & A202;
  assign \new_[36301]_  = ~A234 & A233;
  assign \new_[36302]_  = \new_[36301]_  & \new_[36298]_ ;
  assign \new_[36303]_  = \new_[36302]_  & \new_[36295]_ ;
  assign \new_[36307]_  = ~A268 & ~A267;
  assign \new_[36308]_  = ~A235 & \new_[36307]_ ;
  assign \new_[36311]_  = ~A298 & ~A269;
  assign \new_[36314]_  = ~A301 & ~A299;
  assign \new_[36315]_  = \new_[36314]_  & \new_[36311]_ ;
  assign \new_[36316]_  = \new_[36315]_  & \new_[36308]_ ;
  assign \new_[36320]_  = ~A166 & ~A167;
  assign \new_[36321]_  = ~A169 & \new_[36320]_ ;
  assign \new_[36324]_  = A232 & A202;
  assign \new_[36327]_  = ~A234 & A233;
  assign \new_[36328]_  = \new_[36327]_  & \new_[36324]_ ;
  assign \new_[36329]_  = \new_[36328]_  & \new_[36321]_ ;
  assign \new_[36333]_  = ~A266 & ~A265;
  assign \new_[36334]_  = ~A235 & \new_[36333]_ ;
  assign \new_[36337]_  = ~A300 & ~A268;
  assign \new_[36340]_  = ~A302 & ~A301;
  assign \new_[36341]_  = \new_[36340]_  & \new_[36337]_ ;
  assign \new_[36342]_  = \new_[36341]_  & \new_[36334]_ ;
  assign \new_[36346]_  = ~A166 & ~A167;
  assign \new_[36347]_  = ~A169 & \new_[36346]_ ;
  assign \new_[36350]_  = A232 & A202;
  assign \new_[36353]_  = ~A234 & A233;
  assign \new_[36354]_  = \new_[36353]_  & \new_[36350]_ ;
  assign \new_[36355]_  = \new_[36354]_  & \new_[36347]_ ;
  assign \new_[36359]_  = ~A266 & ~A265;
  assign \new_[36360]_  = ~A235 & \new_[36359]_ ;
  assign \new_[36363]_  = ~A298 & ~A268;
  assign \new_[36366]_  = ~A301 & ~A299;
  assign \new_[36367]_  = \new_[36366]_  & \new_[36363]_ ;
  assign \new_[36368]_  = \new_[36367]_  & \new_[36360]_ ;
  assign \new_[36372]_  = ~A166 & ~A167;
  assign \new_[36373]_  = ~A169 & \new_[36372]_ ;
  assign \new_[36376]_  = ~A232 & A202;
  assign \new_[36379]_  = ~A235 & ~A233;
  assign \new_[36380]_  = \new_[36379]_  & \new_[36376]_ ;
  assign \new_[36381]_  = \new_[36380]_  & \new_[36373]_ ;
  assign \new_[36385]_  = ~A269 & ~A268;
  assign \new_[36386]_  = ~A267 & \new_[36385]_ ;
  assign \new_[36389]_  = A299 & A298;
  assign \new_[36392]_  = ~A301 & ~A300;
  assign \new_[36393]_  = \new_[36392]_  & \new_[36389]_ ;
  assign \new_[36394]_  = \new_[36393]_  & \new_[36386]_ ;
  assign \new_[36398]_  = ~A166 & ~A167;
  assign \new_[36399]_  = ~A169 & \new_[36398]_ ;
  assign \new_[36402]_  = ~A232 & A202;
  assign \new_[36405]_  = ~A235 & ~A233;
  assign \new_[36406]_  = \new_[36405]_  & \new_[36402]_ ;
  assign \new_[36407]_  = \new_[36406]_  & \new_[36399]_ ;
  assign \new_[36411]_  = ~A267 & A266;
  assign \new_[36412]_  = A265 & \new_[36411]_ ;
  assign \new_[36415]_  = ~A300 & ~A268;
  assign \new_[36418]_  = ~A302 & ~A301;
  assign \new_[36419]_  = \new_[36418]_  & \new_[36415]_ ;
  assign \new_[36420]_  = \new_[36419]_  & \new_[36412]_ ;
  assign \new_[36424]_  = ~A166 & ~A167;
  assign \new_[36425]_  = ~A169 & \new_[36424]_ ;
  assign \new_[36428]_  = ~A232 & A202;
  assign \new_[36431]_  = ~A235 & ~A233;
  assign \new_[36432]_  = \new_[36431]_  & \new_[36428]_ ;
  assign \new_[36433]_  = \new_[36432]_  & \new_[36425]_ ;
  assign \new_[36437]_  = ~A267 & A266;
  assign \new_[36438]_  = A265 & \new_[36437]_ ;
  assign \new_[36441]_  = ~A298 & ~A268;
  assign \new_[36444]_  = ~A301 & ~A299;
  assign \new_[36445]_  = \new_[36444]_  & \new_[36441]_ ;
  assign \new_[36446]_  = \new_[36445]_  & \new_[36438]_ ;
  assign \new_[36450]_  = ~A166 & ~A167;
  assign \new_[36451]_  = ~A169 & \new_[36450]_ ;
  assign \new_[36454]_  = ~A232 & A202;
  assign \new_[36457]_  = ~A235 & ~A233;
  assign \new_[36458]_  = \new_[36457]_  & \new_[36454]_ ;
  assign \new_[36459]_  = \new_[36458]_  & \new_[36451]_ ;
  assign \new_[36463]_  = ~A268 & ~A266;
  assign \new_[36464]_  = ~A265 & \new_[36463]_ ;
  assign \new_[36467]_  = A299 & A298;
  assign \new_[36470]_  = ~A301 & ~A300;
  assign \new_[36471]_  = \new_[36470]_  & \new_[36467]_ ;
  assign \new_[36472]_  = \new_[36471]_  & \new_[36464]_ ;
  assign \new_[36476]_  = ~A166 & ~A167;
  assign \new_[36477]_  = ~A169 & \new_[36476]_ ;
  assign \new_[36480]_  = A201 & A199;
  assign \new_[36483]_  = ~A235 & ~A234;
  assign \new_[36484]_  = \new_[36483]_  & \new_[36480]_ ;
  assign \new_[36485]_  = \new_[36484]_  & \new_[36477]_ ;
  assign \new_[36489]_  = ~A268 & ~A267;
  assign \new_[36490]_  = ~A236 & \new_[36489]_ ;
  assign \new_[36493]_  = ~A300 & ~A269;
  assign \new_[36496]_  = ~A302 & ~A301;
  assign \new_[36497]_  = \new_[36496]_  & \new_[36493]_ ;
  assign \new_[36498]_  = \new_[36497]_  & \new_[36490]_ ;
  assign \new_[36502]_  = ~A166 & ~A167;
  assign \new_[36503]_  = ~A169 & \new_[36502]_ ;
  assign \new_[36506]_  = A201 & A199;
  assign \new_[36509]_  = ~A235 & ~A234;
  assign \new_[36510]_  = \new_[36509]_  & \new_[36506]_ ;
  assign \new_[36511]_  = \new_[36510]_  & \new_[36503]_ ;
  assign \new_[36515]_  = ~A268 & ~A267;
  assign \new_[36516]_  = ~A236 & \new_[36515]_ ;
  assign \new_[36519]_  = ~A298 & ~A269;
  assign \new_[36522]_  = ~A301 & ~A299;
  assign \new_[36523]_  = \new_[36522]_  & \new_[36519]_ ;
  assign \new_[36524]_  = \new_[36523]_  & \new_[36516]_ ;
  assign \new_[36528]_  = ~A166 & ~A167;
  assign \new_[36529]_  = ~A169 & \new_[36528]_ ;
  assign \new_[36532]_  = A201 & A199;
  assign \new_[36535]_  = ~A235 & ~A234;
  assign \new_[36536]_  = \new_[36535]_  & \new_[36532]_ ;
  assign \new_[36537]_  = \new_[36536]_  & \new_[36529]_ ;
  assign \new_[36541]_  = ~A266 & ~A265;
  assign \new_[36542]_  = ~A236 & \new_[36541]_ ;
  assign \new_[36545]_  = ~A300 & ~A268;
  assign \new_[36548]_  = ~A302 & ~A301;
  assign \new_[36549]_  = \new_[36548]_  & \new_[36545]_ ;
  assign \new_[36550]_  = \new_[36549]_  & \new_[36542]_ ;
  assign \new_[36554]_  = ~A166 & ~A167;
  assign \new_[36555]_  = ~A169 & \new_[36554]_ ;
  assign \new_[36558]_  = A201 & A199;
  assign \new_[36561]_  = ~A235 & ~A234;
  assign \new_[36562]_  = \new_[36561]_  & \new_[36558]_ ;
  assign \new_[36563]_  = \new_[36562]_  & \new_[36555]_ ;
  assign \new_[36567]_  = ~A266 & ~A265;
  assign \new_[36568]_  = ~A236 & \new_[36567]_ ;
  assign \new_[36571]_  = ~A298 & ~A268;
  assign \new_[36574]_  = ~A301 & ~A299;
  assign \new_[36575]_  = \new_[36574]_  & \new_[36571]_ ;
  assign \new_[36576]_  = \new_[36575]_  & \new_[36568]_ ;
  assign \new_[36580]_  = ~A166 & ~A167;
  assign \new_[36581]_  = ~A169 & \new_[36580]_ ;
  assign \new_[36584]_  = A201 & A199;
  assign \new_[36587]_  = ~A233 & ~A232;
  assign \new_[36588]_  = \new_[36587]_  & \new_[36584]_ ;
  assign \new_[36589]_  = \new_[36588]_  & \new_[36581]_ ;
  assign \new_[36593]_  = ~A268 & ~A267;
  assign \new_[36594]_  = ~A235 & \new_[36593]_ ;
  assign \new_[36597]_  = ~A300 & ~A269;
  assign \new_[36600]_  = ~A302 & ~A301;
  assign \new_[36601]_  = \new_[36600]_  & \new_[36597]_ ;
  assign \new_[36602]_  = \new_[36601]_  & \new_[36594]_ ;
  assign \new_[36606]_  = ~A166 & ~A167;
  assign \new_[36607]_  = ~A169 & \new_[36606]_ ;
  assign \new_[36610]_  = A201 & A199;
  assign \new_[36613]_  = ~A233 & ~A232;
  assign \new_[36614]_  = \new_[36613]_  & \new_[36610]_ ;
  assign \new_[36615]_  = \new_[36614]_  & \new_[36607]_ ;
  assign \new_[36619]_  = ~A268 & ~A267;
  assign \new_[36620]_  = ~A235 & \new_[36619]_ ;
  assign \new_[36623]_  = ~A298 & ~A269;
  assign \new_[36626]_  = ~A301 & ~A299;
  assign \new_[36627]_  = \new_[36626]_  & \new_[36623]_ ;
  assign \new_[36628]_  = \new_[36627]_  & \new_[36620]_ ;
  assign \new_[36632]_  = ~A166 & ~A167;
  assign \new_[36633]_  = ~A169 & \new_[36632]_ ;
  assign \new_[36636]_  = A201 & A199;
  assign \new_[36639]_  = ~A233 & ~A232;
  assign \new_[36640]_  = \new_[36639]_  & \new_[36636]_ ;
  assign \new_[36641]_  = \new_[36640]_  & \new_[36633]_ ;
  assign \new_[36645]_  = ~A266 & ~A265;
  assign \new_[36646]_  = ~A235 & \new_[36645]_ ;
  assign \new_[36649]_  = ~A300 & ~A268;
  assign \new_[36652]_  = ~A302 & ~A301;
  assign \new_[36653]_  = \new_[36652]_  & \new_[36649]_ ;
  assign \new_[36654]_  = \new_[36653]_  & \new_[36646]_ ;
  assign \new_[36658]_  = ~A166 & ~A167;
  assign \new_[36659]_  = ~A169 & \new_[36658]_ ;
  assign \new_[36662]_  = A201 & A199;
  assign \new_[36665]_  = ~A233 & ~A232;
  assign \new_[36666]_  = \new_[36665]_  & \new_[36662]_ ;
  assign \new_[36667]_  = \new_[36666]_  & \new_[36659]_ ;
  assign \new_[36671]_  = ~A266 & ~A265;
  assign \new_[36672]_  = ~A235 & \new_[36671]_ ;
  assign \new_[36675]_  = ~A298 & ~A268;
  assign \new_[36678]_  = ~A301 & ~A299;
  assign \new_[36679]_  = \new_[36678]_  & \new_[36675]_ ;
  assign \new_[36680]_  = \new_[36679]_  & \new_[36672]_ ;
  assign \new_[36684]_  = ~A166 & ~A167;
  assign \new_[36685]_  = ~A169 & \new_[36684]_ ;
  assign \new_[36688]_  = A201 & A200;
  assign \new_[36691]_  = ~A235 & ~A234;
  assign \new_[36692]_  = \new_[36691]_  & \new_[36688]_ ;
  assign \new_[36693]_  = \new_[36692]_  & \new_[36685]_ ;
  assign \new_[36697]_  = ~A268 & ~A267;
  assign \new_[36698]_  = ~A236 & \new_[36697]_ ;
  assign \new_[36701]_  = ~A300 & ~A269;
  assign \new_[36704]_  = ~A302 & ~A301;
  assign \new_[36705]_  = \new_[36704]_  & \new_[36701]_ ;
  assign \new_[36706]_  = \new_[36705]_  & \new_[36698]_ ;
  assign \new_[36710]_  = ~A166 & ~A167;
  assign \new_[36711]_  = ~A169 & \new_[36710]_ ;
  assign \new_[36714]_  = A201 & A200;
  assign \new_[36717]_  = ~A235 & ~A234;
  assign \new_[36718]_  = \new_[36717]_  & \new_[36714]_ ;
  assign \new_[36719]_  = \new_[36718]_  & \new_[36711]_ ;
  assign \new_[36723]_  = ~A268 & ~A267;
  assign \new_[36724]_  = ~A236 & \new_[36723]_ ;
  assign \new_[36727]_  = ~A298 & ~A269;
  assign \new_[36730]_  = ~A301 & ~A299;
  assign \new_[36731]_  = \new_[36730]_  & \new_[36727]_ ;
  assign \new_[36732]_  = \new_[36731]_  & \new_[36724]_ ;
  assign \new_[36736]_  = ~A166 & ~A167;
  assign \new_[36737]_  = ~A169 & \new_[36736]_ ;
  assign \new_[36740]_  = A201 & A200;
  assign \new_[36743]_  = ~A235 & ~A234;
  assign \new_[36744]_  = \new_[36743]_  & \new_[36740]_ ;
  assign \new_[36745]_  = \new_[36744]_  & \new_[36737]_ ;
  assign \new_[36749]_  = ~A266 & ~A265;
  assign \new_[36750]_  = ~A236 & \new_[36749]_ ;
  assign \new_[36753]_  = ~A300 & ~A268;
  assign \new_[36756]_  = ~A302 & ~A301;
  assign \new_[36757]_  = \new_[36756]_  & \new_[36753]_ ;
  assign \new_[36758]_  = \new_[36757]_  & \new_[36750]_ ;
  assign \new_[36762]_  = ~A166 & ~A167;
  assign \new_[36763]_  = ~A169 & \new_[36762]_ ;
  assign \new_[36766]_  = A201 & A200;
  assign \new_[36769]_  = ~A235 & ~A234;
  assign \new_[36770]_  = \new_[36769]_  & \new_[36766]_ ;
  assign \new_[36771]_  = \new_[36770]_  & \new_[36763]_ ;
  assign \new_[36775]_  = ~A266 & ~A265;
  assign \new_[36776]_  = ~A236 & \new_[36775]_ ;
  assign \new_[36779]_  = ~A298 & ~A268;
  assign \new_[36782]_  = ~A301 & ~A299;
  assign \new_[36783]_  = \new_[36782]_  & \new_[36779]_ ;
  assign \new_[36784]_  = \new_[36783]_  & \new_[36776]_ ;
  assign \new_[36788]_  = ~A166 & ~A167;
  assign \new_[36789]_  = ~A169 & \new_[36788]_ ;
  assign \new_[36792]_  = A201 & A200;
  assign \new_[36795]_  = ~A233 & ~A232;
  assign \new_[36796]_  = \new_[36795]_  & \new_[36792]_ ;
  assign \new_[36797]_  = \new_[36796]_  & \new_[36789]_ ;
  assign \new_[36801]_  = ~A268 & ~A267;
  assign \new_[36802]_  = ~A235 & \new_[36801]_ ;
  assign \new_[36805]_  = ~A300 & ~A269;
  assign \new_[36808]_  = ~A302 & ~A301;
  assign \new_[36809]_  = \new_[36808]_  & \new_[36805]_ ;
  assign \new_[36810]_  = \new_[36809]_  & \new_[36802]_ ;
  assign \new_[36814]_  = ~A166 & ~A167;
  assign \new_[36815]_  = ~A169 & \new_[36814]_ ;
  assign \new_[36818]_  = A201 & A200;
  assign \new_[36821]_  = ~A233 & ~A232;
  assign \new_[36822]_  = \new_[36821]_  & \new_[36818]_ ;
  assign \new_[36823]_  = \new_[36822]_  & \new_[36815]_ ;
  assign \new_[36827]_  = ~A268 & ~A267;
  assign \new_[36828]_  = ~A235 & \new_[36827]_ ;
  assign \new_[36831]_  = ~A298 & ~A269;
  assign \new_[36834]_  = ~A301 & ~A299;
  assign \new_[36835]_  = \new_[36834]_  & \new_[36831]_ ;
  assign \new_[36836]_  = \new_[36835]_  & \new_[36828]_ ;
  assign \new_[36840]_  = ~A166 & ~A167;
  assign \new_[36841]_  = ~A169 & \new_[36840]_ ;
  assign \new_[36844]_  = A201 & A200;
  assign \new_[36847]_  = ~A233 & ~A232;
  assign \new_[36848]_  = \new_[36847]_  & \new_[36844]_ ;
  assign \new_[36849]_  = \new_[36848]_  & \new_[36841]_ ;
  assign \new_[36853]_  = ~A266 & ~A265;
  assign \new_[36854]_  = ~A235 & \new_[36853]_ ;
  assign \new_[36857]_  = ~A300 & ~A268;
  assign \new_[36860]_  = ~A302 & ~A301;
  assign \new_[36861]_  = \new_[36860]_  & \new_[36857]_ ;
  assign \new_[36862]_  = \new_[36861]_  & \new_[36854]_ ;
  assign \new_[36866]_  = ~A166 & ~A167;
  assign \new_[36867]_  = ~A169 & \new_[36866]_ ;
  assign \new_[36870]_  = A201 & A200;
  assign \new_[36873]_  = ~A233 & ~A232;
  assign \new_[36874]_  = \new_[36873]_  & \new_[36870]_ ;
  assign \new_[36875]_  = \new_[36874]_  & \new_[36867]_ ;
  assign \new_[36879]_  = ~A266 & ~A265;
  assign \new_[36880]_  = ~A235 & \new_[36879]_ ;
  assign \new_[36883]_  = ~A298 & ~A268;
  assign \new_[36886]_  = ~A301 & ~A299;
  assign \new_[36887]_  = \new_[36886]_  & \new_[36883]_ ;
  assign \new_[36888]_  = \new_[36887]_  & \new_[36880]_ ;
  assign \new_[36892]_  = A167 & ~A168;
  assign \new_[36893]_  = ~A169 & \new_[36892]_ ;
  assign \new_[36896]_  = A202 & A166;
  assign \new_[36899]_  = ~A235 & ~A234;
  assign \new_[36900]_  = \new_[36899]_  & \new_[36896]_ ;
  assign \new_[36901]_  = \new_[36900]_  & \new_[36893]_ ;
  assign \new_[36905]_  = ~A268 & ~A267;
  assign \new_[36906]_  = ~A236 & \new_[36905]_ ;
  assign \new_[36909]_  = ~A300 & ~A269;
  assign \new_[36912]_  = ~A302 & ~A301;
  assign \new_[36913]_  = \new_[36912]_  & \new_[36909]_ ;
  assign \new_[36914]_  = \new_[36913]_  & \new_[36906]_ ;
  assign \new_[36918]_  = A167 & ~A168;
  assign \new_[36919]_  = ~A169 & \new_[36918]_ ;
  assign \new_[36922]_  = A202 & A166;
  assign \new_[36925]_  = ~A235 & ~A234;
  assign \new_[36926]_  = \new_[36925]_  & \new_[36922]_ ;
  assign \new_[36927]_  = \new_[36926]_  & \new_[36919]_ ;
  assign \new_[36931]_  = ~A268 & ~A267;
  assign \new_[36932]_  = ~A236 & \new_[36931]_ ;
  assign \new_[36935]_  = ~A298 & ~A269;
  assign \new_[36938]_  = ~A301 & ~A299;
  assign \new_[36939]_  = \new_[36938]_  & \new_[36935]_ ;
  assign \new_[36940]_  = \new_[36939]_  & \new_[36932]_ ;
  assign \new_[36944]_  = A167 & ~A168;
  assign \new_[36945]_  = ~A169 & \new_[36944]_ ;
  assign \new_[36948]_  = A202 & A166;
  assign \new_[36951]_  = ~A235 & ~A234;
  assign \new_[36952]_  = \new_[36951]_  & \new_[36948]_ ;
  assign \new_[36953]_  = \new_[36952]_  & \new_[36945]_ ;
  assign \new_[36957]_  = ~A266 & ~A265;
  assign \new_[36958]_  = ~A236 & \new_[36957]_ ;
  assign \new_[36961]_  = ~A300 & ~A268;
  assign \new_[36964]_  = ~A302 & ~A301;
  assign \new_[36965]_  = \new_[36964]_  & \new_[36961]_ ;
  assign \new_[36966]_  = \new_[36965]_  & \new_[36958]_ ;
  assign \new_[36970]_  = A167 & ~A168;
  assign \new_[36971]_  = ~A169 & \new_[36970]_ ;
  assign \new_[36974]_  = A202 & A166;
  assign \new_[36977]_  = ~A235 & ~A234;
  assign \new_[36978]_  = \new_[36977]_  & \new_[36974]_ ;
  assign \new_[36979]_  = \new_[36978]_  & \new_[36971]_ ;
  assign \new_[36983]_  = ~A266 & ~A265;
  assign \new_[36984]_  = ~A236 & \new_[36983]_ ;
  assign \new_[36987]_  = ~A298 & ~A268;
  assign \new_[36990]_  = ~A301 & ~A299;
  assign \new_[36991]_  = \new_[36990]_  & \new_[36987]_ ;
  assign \new_[36992]_  = \new_[36991]_  & \new_[36984]_ ;
  assign \new_[36996]_  = A167 & ~A168;
  assign \new_[36997]_  = ~A169 & \new_[36996]_ ;
  assign \new_[37000]_  = A202 & A166;
  assign \new_[37003]_  = ~A233 & ~A232;
  assign \new_[37004]_  = \new_[37003]_  & \new_[37000]_ ;
  assign \new_[37005]_  = \new_[37004]_  & \new_[36997]_ ;
  assign \new_[37009]_  = ~A268 & ~A267;
  assign \new_[37010]_  = ~A235 & \new_[37009]_ ;
  assign \new_[37013]_  = ~A300 & ~A269;
  assign \new_[37016]_  = ~A302 & ~A301;
  assign \new_[37017]_  = \new_[37016]_  & \new_[37013]_ ;
  assign \new_[37018]_  = \new_[37017]_  & \new_[37010]_ ;
  assign \new_[37022]_  = A167 & ~A168;
  assign \new_[37023]_  = ~A169 & \new_[37022]_ ;
  assign \new_[37026]_  = A202 & A166;
  assign \new_[37029]_  = ~A233 & ~A232;
  assign \new_[37030]_  = \new_[37029]_  & \new_[37026]_ ;
  assign \new_[37031]_  = \new_[37030]_  & \new_[37023]_ ;
  assign \new_[37035]_  = ~A268 & ~A267;
  assign \new_[37036]_  = ~A235 & \new_[37035]_ ;
  assign \new_[37039]_  = ~A298 & ~A269;
  assign \new_[37042]_  = ~A301 & ~A299;
  assign \new_[37043]_  = \new_[37042]_  & \new_[37039]_ ;
  assign \new_[37044]_  = \new_[37043]_  & \new_[37036]_ ;
  assign \new_[37048]_  = A167 & ~A168;
  assign \new_[37049]_  = ~A169 & \new_[37048]_ ;
  assign \new_[37052]_  = A202 & A166;
  assign \new_[37055]_  = ~A233 & ~A232;
  assign \new_[37056]_  = \new_[37055]_  & \new_[37052]_ ;
  assign \new_[37057]_  = \new_[37056]_  & \new_[37049]_ ;
  assign \new_[37061]_  = ~A266 & ~A265;
  assign \new_[37062]_  = ~A235 & \new_[37061]_ ;
  assign \new_[37065]_  = ~A300 & ~A268;
  assign \new_[37068]_  = ~A302 & ~A301;
  assign \new_[37069]_  = \new_[37068]_  & \new_[37065]_ ;
  assign \new_[37070]_  = \new_[37069]_  & \new_[37062]_ ;
  assign \new_[37074]_  = A167 & ~A168;
  assign \new_[37075]_  = ~A169 & \new_[37074]_ ;
  assign \new_[37078]_  = A202 & A166;
  assign \new_[37081]_  = ~A233 & ~A232;
  assign \new_[37082]_  = \new_[37081]_  & \new_[37078]_ ;
  assign \new_[37083]_  = \new_[37082]_  & \new_[37075]_ ;
  assign \new_[37087]_  = ~A266 & ~A265;
  assign \new_[37088]_  = ~A235 & \new_[37087]_ ;
  assign \new_[37091]_  = ~A298 & ~A268;
  assign \new_[37094]_  = ~A301 & ~A299;
  assign \new_[37095]_  = \new_[37094]_  & \new_[37091]_ ;
  assign \new_[37096]_  = \new_[37095]_  & \new_[37088]_ ;
  assign \new_[37100]_  = ~A168 & ~A169;
  assign \new_[37101]_  = ~A170 & \new_[37100]_ ;
  assign \new_[37104]_  = ~A234 & A202;
  assign \new_[37107]_  = ~A236 & ~A235;
  assign \new_[37108]_  = \new_[37107]_  & \new_[37104]_ ;
  assign \new_[37109]_  = \new_[37108]_  & \new_[37101]_ ;
  assign \new_[37113]_  = ~A269 & ~A268;
  assign \new_[37114]_  = ~A267 & \new_[37113]_ ;
  assign \new_[37117]_  = A299 & A298;
  assign \new_[37120]_  = ~A301 & ~A300;
  assign \new_[37121]_  = \new_[37120]_  & \new_[37117]_ ;
  assign \new_[37122]_  = \new_[37121]_  & \new_[37114]_ ;
  assign \new_[37126]_  = ~A168 & ~A169;
  assign \new_[37127]_  = ~A170 & \new_[37126]_ ;
  assign \new_[37130]_  = ~A234 & A202;
  assign \new_[37133]_  = ~A236 & ~A235;
  assign \new_[37134]_  = \new_[37133]_  & \new_[37130]_ ;
  assign \new_[37135]_  = \new_[37134]_  & \new_[37127]_ ;
  assign \new_[37139]_  = ~A267 & A266;
  assign \new_[37140]_  = A265 & \new_[37139]_ ;
  assign \new_[37143]_  = ~A300 & ~A268;
  assign \new_[37146]_  = ~A302 & ~A301;
  assign \new_[37147]_  = \new_[37146]_  & \new_[37143]_ ;
  assign \new_[37148]_  = \new_[37147]_  & \new_[37140]_ ;
  assign \new_[37152]_  = ~A168 & ~A169;
  assign \new_[37153]_  = ~A170 & \new_[37152]_ ;
  assign \new_[37156]_  = ~A234 & A202;
  assign \new_[37159]_  = ~A236 & ~A235;
  assign \new_[37160]_  = \new_[37159]_  & \new_[37156]_ ;
  assign \new_[37161]_  = \new_[37160]_  & \new_[37153]_ ;
  assign \new_[37165]_  = ~A267 & A266;
  assign \new_[37166]_  = A265 & \new_[37165]_ ;
  assign \new_[37169]_  = ~A298 & ~A268;
  assign \new_[37172]_  = ~A301 & ~A299;
  assign \new_[37173]_  = \new_[37172]_  & \new_[37169]_ ;
  assign \new_[37174]_  = \new_[37173]_  & \new_[37166]_ ;
  assign \new_[37178]_  = ~A168 & ~A169;
  assign \new_[37179]_  = ~A170 & \new_[37178]_ ;
  assign \new_[37182]_  = ~A234 & A202;
  assign \new_[37185]_  = ~A236 & ~A235;
  assign \new_[37186]_  = \new_[37185]_  & \new_[37182]_ ;
  assign \new_[37187]_  = \new_[37186]_  & \new_[37179]_ ;
  assign \new_[37191]_  = ~A268 & ~A266;
  assign \new_[37192]_  = ~A265 & \new_[37191]_ ;
  assign \new_[37195]_  = A299 & A298;
  assign \new_[37198]_  = ~A301 & ~A300;
  assign \new_[37199]_  = \new_[37198]_  & \new_[37195]_ ;
  assign \new_[37200]_  = \new_[37199]_  & \new_[37192]_ ;
  assign \new_[37204]_  = ~A168 & ~A169;
  assign \new_[37205]_  = ~A170 & \new_[37204]_ ;
  assign \new_[37208]_  = A232 & A202;
  assign \new_[37211]_  = ~A234 & A233;
  assign \new_[37212]_  = \new_[37211]_  & \new_[37208]_ ;
  assign \new_[37213]_  = \new_[37212]_  & \new_[37205]_ ;
  assign \new_[37217]_  = ~A268 & ~A267;
  assign \new_[37218]_  = ~A235 & \new_[37217]_ ;
  assign \new_[37221]_  = ~A300 & ~A269;
  assign \new_[37224]_  = ~A302 & ~A301;
  assign \new_[37225]_  = \new_[37224]_  & \new_[37221]_ ;
  assign \new_[37226]_  = \new_[37225]_  & \new_[37218]_ ;
  assign \new_[37230]_  = ~A168 & ~A169;
  assign \new_[37231]_  = ~A170 & \new_[37230]_ ;
  assign \new_[37234]_  = A232 & A202;
  assign \new_[37237]_  = ~A234 & A233;
  assign \new_[37238]_  = \new_[37237]_  & \new_[37234]_ ;
  assign \new_[37239]_  = \new_[37238]_  & \new_[37231]_ ;
  assign \new_[37243]_  = ~A268 & ~A267;
  assign \new_[37244]_  = ~A235 & \new_[37243]_ ;
  assign \new_[37247]_  = ~A298 & ~A269;
  assign \new_[37250]_  = ~A301 & ~A299;
  assign \new_[37251]_  = \new_[37250]_  & \new_[37247]_ ;
  assign \new_[37252]_  = \new_[37251]_  & \new_[37244]_ ;
  assign \new_[37256]_  = ~A168 & ~A169;
  assign \new_[37257]_  = ~A170 & \new_[37256]_ ;
  assign \new_[37260]_  = A232 & A202;
  assign \new_[37263]_  = ~A234 & A233;
  assign \new_[37264]_  = \new_[37263]_  & \new_[37260]_ ;
  assign \new_[37265]_  = \new_[37264]_  & \new_[37257]_ ;
  assign \new_[37269]_  = ~A266 & ~A265;
  assign \new_[37270]_  = ~A235 & \new_[37269]_ ;
  assign \new_[37273]_  = ~A300 & ~A268;
  assign \new_[37276]_  = ~A302 & ~A301;
  assign \new_[37277]_  = \new_[37276]_  & \new_[37273]_ ;
  assign \new_[37278]_  = \new_[37277]_  & \new_[37270]_ ;
  assign \new_[37282]_  = ~A168 & ~A169;
  assign \new_[37283]_  = ~A170 & \new_[37282]_ ;
  assign \new_[37286]_  = A232 & A202;
  assign \new_[37289]_  = ~A234 & A233;
  assign \new_[37290]_  = \new_[37289]_  & \new_[37286]_ ;
  assign \new_[37291]_  = \new_[37290]_  & \new_[37283]_ ;
  assign \new_[37295]_  = ~A266 & ~A265;
  assign \new_[37296]_  = ~A235 & \new_[37295]_ ;
  assign \new_[37299]_  = ~A298 & ~A268;
  assign \new_[37302]_  = ~A301 & ~A299;
  assign \new_[37303]_  = \new_[37302]_  & \new_[37299]_ ;
  assign \new_[37304]_  = \new_[37303]_  & \new_[37296]_ ;
  assign \new_[37308]_  = ~A168 & ~A169;
  assign \new_[37309]_  = ~A170 & \new_[37308]_ ;
  assign \new_[37312]_  = ~A232 & A202;
  assign \new_[37315]_  = ~A235 & ~A233;
  assign \new_[37316]_  = \new_[37315]_  & \new_[37312]_ ;
  assign \new_[37317]_  = \new_[37316]_  & \new_[37309]_ ;
  assign \new_[37321]_  = ~A269 & ~A268;
  assign \new_[37322]_  = ~A267 & \new_[37321]_ ;
  assign \new_[37325]_  = A299 & A298;
  assign \new_[37328]_  = ~A301 & ~A300;
  assign \new_[37329]_  = \new_[37328]_  & \new_[37325]_ ;
  assign \new_[37330]_  = \new_[37329]_  & \new_[37322]_ ;
  assign \new_[37334]_  = ~A168 & ~A169;
  assign \new_[37335]_  = ~A170 & \new_[37334]_ ;
  assign \new_[37338]_  = ~A232 & A202;
  assign \new_[37341]_  = ~A235 & ~A233;
  assign \new_[37342]_  = \new_[37341]_  & \new_[37338]_ ;
  assign \new_[37343]_  = \new_[37342]_  & \new_[37335]_ ;
  assign \new_[37347]_  = ~A267 & A266;
  assign \new_[37348]_  = A265 & \new_[37347]_ ;
  assign \new_[37351]_  = ~A300 & ~A268;
  assign \new_[37354]_  = ~A302 & ~A301;
  assign \new_[37355]_  = \new_[37354]_  & \new_[37351]_ ;
  assign \new_[37356]_  = \new_[37355]_  & \new_[37348]_ ;
  assign \new_[37360]_  = ~A168 & ~A169;
  assign \new_[37361]_  = ~A170 & \new_[37360]_ ;
  assign \new_[37364]_  = ~A232 & A202;
  assign \new_[37367]_  = ~A235 & ~A233;
  assign \new_[37368]_  = \new_[37367]_  & \new_[37364]_ ;
  assign \new_[37369]_  = \new_[37368]_  & \new_[37361]_ ;
  assign \new_[37373]_  = ~A267 & A266;
  assign \new_[37374]_  = A265 & \new_[37373]_ ;
  assign \new_[37377]_  = ~A298 & ~A268;
  assign \new_[37380]_  = ~A301 & ~A299;
  assign \new_[37381]_  = \new_[37380]_  & \new_[37377]_ ;
  assign \new_[37382]_  = \new_[37381]_  & \new_[37374]_ ;
  assign \new_[37386]_  = ~A168 & ~A169;
  assign \new_[37387]_  = ~A170 & \new_[37386]_ ;
  assign \new_[37390]_  = ~A232 & A202;
  assign \new_[37393]_  = ~A235 & ~A233;
  assign \new_[37394]_  = \new_[37393]_  & \new_[37390]_ ;
  assign \new_[37395]_  = \new_[37394]_  & \new_[37387]_ ;
  assign \new_[37399]_  = ~A268 & ~A266;
  assign \new_[37400]_  = ~A265 & \new_[37399]_ ;
  assign \new_[37403]_  = A299 & A298;
  assign \new_[37406]_  = ~A301 & ~A300;
  assign \new_[37407]_  = \new_[37406]_  & \new_[37403]_ ;
  assign \new_[37408]_  = \new_[37407]_  & \new_[37400]_ ;
  assign \new_[37412]_  = ~A168 & ~A169;
  assign \new_[37413]_  = ~A170 & \new_[37412]_ ;
  assign \new_[37416]_  = A201 & A199;
  assign \new_[37419]_  = ~A235 & ~A234;
  assign \new_[37420]_  = \new_[37419]_  & \new_[37416]_ ;
  assign \new_[37421]_  = \new_[37420]_  & \new_[37413]_ ;
  assign \new_[37425]_  = ~A268 & ~A267;
  assign \new_[37426]_  = ~A236 & \new_[37425]_ ;
  assign \new_[37429]_  = ~A300 & ~A269;
  assign \new_[37432]_  = ~A302 & ~A301;
  assign \new_[37433]_  = \new_[37432]_  & \new_[37429]_ ;
  assign \new_[37434]_  = \new_[37433]_  & \new_[37426]_ ;
  assign \new_[37438]_  = ~A168 & ~A169;
  assign \new_[37439]_  = ~A170 & \new_[37438]_ ;
  assign \new_[37442]_  = A201 & A199;
  assign \new_[37445]_  = ~A235 & ~A234;
  assign \new_[37446]_  = \new_[37445]_  & \new_[37442]_ ;
  assign \new_[37447]_  = \new_[37446]_  & \new_[37439]_ ;
  assign \new_[37451]_  = ~A268 & ~A267;
  assign \new_[37452]_  = ~A236 & \new_[37451]_ ;
  assign \new_[37455]_  = ~A298 & ~A269;
  assign \new_[37458]_  = ~A301 & ~A299;
  assign \new_[37459]_  = \new_[37458]_  & \new_[37455]_ ;
  assign \new_[37460]_  = \new_[37459]_  & \new_[37452]_ ;
  assign \new_[37464]_  = ~A168 & ~A169;
  assign \new_[37465]_  = ~A170 & \new_[37464]_ ;
  assign \new_[37468]_  = A201 & A199;
  assign \new_[37471]_  = ~A235 & ~A234;
  assign \new_[37472]_  = \new_[37471]_  & \new_[37468]_ ;
  assign \new_[37473]_  = \new_[37472]_  & \new_[37465]_ ;
  assign \new_[37477]_  = ~A266 & ~A265;
  assign \new_[37478]_  = ~A236 & \new_[37477]_ ;
  assign \new_[37481]_  = ~A300 & ~A268;
  assign \new_[37484]_  = ~A302 & ~A301;
  assign \new_[37485]_  = \new_[37484]_  & \new_[37481]_ ;
  assign \new_[37486]_  = \new_[37485]_  & \new_[37478]_ ;
  assign \new_[37490]_  = ~A168 & ~A169;
  assign \new_[37491]_  = ~A170 & \new_[37490]_ ;
  assign \new_[37494]_  = A201 & A199;
  assign \new_[37497]_  = ~A235 & ~A234;
  assign \new_[37498]_  = \new_[37497]_  & \new_[37494]_ ;
  assign \new_[37499]_  = \new_[37498]_  & \new_[37491]_ ;
  assign \new_[37503]_  = ~A266 & ~A265;
  assign \new_[37504]_  = ~A236 & \new_[37503]_ ;
  assign \new_[37507]_  = ~A298 & ~A268;
  assign \new_[37510]_  = ~A301 & ~A299;
  assign \new_[37511]_  = \new_[37510]_  & \new_[37507]_ ;
  assign \new_[37512]_  = \new_[37511]_  & \new_[37504]_ ;
  assign \new_[37516]_  = ~A168 & ~A169;
  assign \new_[37517]_  = ~A170 & \new_[37516]_ ;
  assign \new_[37520]_  = A201 & A199;
  assign \new_[37523]_  = ~A233 & ~A232;
  assign \new_[37524]_  = \new_[37523]_  & \new_[37520]_ ;
  assign \new_[37525]_  = \new_[37524]_  & \new_[37517]_ ;
  assign \new_[37529]_  = ~A268 & ~A267;
  assign \new_[37530]_  = ~A235 & \new_[37529]_ ;
  assign \new_[37533]_  = ~A300 & ~A269;
  assign \new_[37536]_  = ~A302 & ~A301;
  assign \new_[37537]_  = \new_[37536]_  & \new_[37533]_ ;
  assign \new_[37538]_  = \new_[37537]_  & \new_[37530]_ ;
  assign \new_[37542]_  = ~A168 & ~A169;
  assign \new_[37543]_  = ~A170 & \new_[37542]_ ;
  assign \new_[37546]_  = A201 & A199;
  assign \new_[37549]_  = ~A233 & ~A232;
  assign \new_[37550]_  = \new_[37549]_  & \new_[37546]_ ;
  assign \new_[37551]_  = \new_[37550]_  & \new_[37543]_ ;
  assign \new_[37555]_  = ~A268 & ~A267;
  assign \new_[37556]_  = ~A235 & \new_[37555]_ ;
  assign \new_[37559]_  = ~A298 & ~A269;
  assign \new_[37562]_  = ~A301 & ~A299;
  assign \new_[37563]_  = \new_[37562]_  & \new_[37559]_ ;
  assign \new_[37564]_  = \new_[37563]_  & \new_[37556]_ ;
  assign \new_[37568]_  = ~A168 & ~A169;
  assign \new_[37569]_  = ~A170 & \new_[37568]_ ;
  assign \new_[37572]_  = A201 & A199;
  assign \new_[37575]_  = ~A233 & ~A232;
  assign \new_[37576]_  = \new_[37575]_  & \new_[37572]_ ;
  assign \new_[37577]_  = \new_[37576]_  & \new_[37569]_ ;
  assign \new_[37581]_  = ~A266 & ~A265;
  assign \new_[37582]_  = ~A235 & \new_[37581]_ ;
  assign \new_[37585]_  = ~A300 & ~A268;
  assign \new_[37588]_  = ~A302 & ~A301;
  assign \new_[37589]_  = \new_[37588]_  & \new_[37585]_ ;
  assign \new_[37590]_  = \new_[37589]_  & \new_[37582]_ ;
  assign \new_[37594]_  = ~A168 & ~A169;
  assign \new_[37595]_  = ~A170 & \new_[37594]_ ;
  assign \new_[37598]_  = A201 & A199;
  assign \new_[37601]_  = ~A233 & ~A232;
  assign \new_[37602]_  = \new_[37601]_  & \new_[37598]_ ;
  assign \new_[37603]_  = \new_[37602]_  & \new_[37595]_ ;
  assign \new_[37607]_  = ~A266 & ~A265;
  assign \new_[37608]_  = ~A235 & \new_[37607]_ ;
  assign \new_[37611]_  = ~A298 & ~A268;
  assign \new_[37614]_  = ~A301 & ~A299;
  assign \new_[37615]_  = \new_[37614]_  & \new_[37611]_ ;
  assign \new_[37616]_  = \new_[37615]_  & \new_[37608]_ ;
  assign \new_[37620]_  = ~A168 & ~A169;
  assign \new_[37621]_  = ~A170 & \new_[37620]_ ;
  assign \new_[37624]_  = A201 & A200;
  assign \new_[37627]_  = ~A235 & ~A234;
  assign \new_[37628]_  = \new_[37627]_  & \new_[37624]_ ;
  assign \new_[37629]_  = \new_[37628]_  & \new_[37621]_ ;
  assign \new_[37633]_  = ~A268 & ~A267;
  assign \new_[37634]_  = ~A236 & \new_[37633]_ ;
  assign \new_[37637]_  = ~A300 & ~A269;
  assign \new_[37640]_  = ~A302 & ~A301;
  assign \new_[37641]_  = \new_[37640]_  & \new_[37637]_ ;
  assign \new_[37642]_  = \new_[37641]_  & \new_[37634]_ ;
  assign \new_[37646]_  = ~A168 & ~A169;
  assign \new_[37647]_  = ~A170 & \new_[37646]_ ;
  assign \new_[37650]_  = A201 & A200;
  assign \new_[37653]_  = ~A235 & ~A234;
  assign \new_[37654]_  = \new_[37653]_  & \new_[37650]_ ;
  assign \new_[37655]_  = \new_[37654]_  & \new_[37647]_ ;
  assign \new_[37659]_  = ~A268 & ~A267;
  assign \new_[37660]_  = ~A236 & \new_[37659]_ ;
  assign \new_[37663]_  = ~A298 & ~A269;
  assign \new_[37666]_  = ~A301 & ~A299;
  assign \new_[37667]_  = \new_[37666]_  & \new_[37663]_ ;
  assign \new_[37668]_  = \new_[37667]_  & \new_[37660]_ ;
  assign \new_[37672]_  = ~A168 & ~A169;
  assign \new_[37673]_  = ~A170 & \new_[37672]_ ;
  assign \new_[37676]_  = A201 & A200;
  assign \new_[37679]_  = ~A235 & ~A234;
  assign \new_[37680]_  = \new_[37679]_  & \new_[37676]_ ;
  assign \new_[37681]_  = \new_[37680]_  & \new_[37673]_ ;
  assign \new_[37685]_  = ~A266 & ~A265;
  assign \new_[37686]_  = ~A236 & \new_[37685]_ ;
  assign \new_[37689]_  = ~A300 & ~A268;
  assign \new_[37692]_  = ~A302 & ~A301;
  assign \new_[37693]_  = \new_[37692]_  & \new_[37689]_ ;
  assign \new_[37694]_  = \new_[37693]_  & \new_[37686]_ ;
  assign \new_[37698]_  = ~A168 & ~A169;
  assign \new_[37699]_  = ~A170 & \new_[37698]_ ;
  assign \new_[37702]_  = A201 & A200;
  assign \new_[37705]_  = ~A235 & ~A234;
  assign \new_[37706]_  = \new_[37705]_  & \new_[37702]_ ;
  assign \new_[37707]_  = \new_[37706]_  & \new_[37699]_ ;
  assign \new_[37711]_  = ~A266 & ~A265;
  assign \new_[37712]_  = ~A236 & \new_[37711]_ ;
  assign \new_[37715]_  = ~A298 & ~A268;
  assign \new_[37718]_  = ~A301 & ~A299;
  assign \new_[37719]_  = \new_[37718]_  & \new_[37715]_ ;
  assign \new_[37720]_  = \new_[37719]_  & \new_[37712]_ ;
  assign \new_[37724]_  = ~A168 & ~A169;
  assign \new_[37725]_  = ~A170 & \new_[37724]_ ;
  assign \new_[37728]_  = A201 & A200;
  assign \new_[37731]_  = ~A233 & ~A232;
  assign \new_[37732]_  = \new_[37731]_  & \new_[37728]_ ;
  assign \new_[37733]_  = \new_[37732]_  & \new_[37725]_ ;
  assign \new_[37737]_  = ~A268 & ~A267;
  assign \new_[37738]_  = ~A235 & \new_[37737]_ ;
  assign \new_[37741]_  = ~A300 & ~A269;
  assign \new_[37744]_  = ~A302 & ~A301;
  assign \new_[37745]_  = \new_[37744]_  & \new_[37741]_ ;
  assign \new_[37746]_  = \new_[37745]_  & \new_[37738]_ ;
  assign \new_[37750]_  = ~A168 & ~A169;
  assign \new_[37751]_  = ~A170 & \new_[37750]_ ;
  assign \new_[37754]_  = A201 & A200;
  assign \new_[37757]_  = ~A233 & ~A232;
  assign \new_[37758]_  = \new_[37757]_  & \new_[37754]_ ;
  assign \new_[37759]_  = \new_[37758]_  & \new_[37751]_ ;
  assign \new_[37763]_  = ~A268 & ~A267;
  assign \new_[37764]_  = ~A235 & \new_[37763]_ ;
  assign \new_[37767]_  = ~A298 & ~A269;
  assign \new_[37770]_  = ~A301 & ~A299;
  assign \new_[37771]_  = \new_[37770]_  & \new_[37767]_ ;
  assign \new_[37772]_  = \new_[37771]_  & \new_[37764]_ ;
  assign \new_[37776]_  = ~A168 & ~A169;
  assign \new_[37777]_  = ~A170 & \new_[37776]_ ;
  assign \new_[37780]_  = A201 & A200;
  assign \new_[37783]_  = ~A233 & ~A232;
  assign \new_[37784]_  = \new_[37783]_  & \new_[37780]_ ;
  assign \new_[37785]_  = \new_[37784]_  & \new_[37777]_ ;
  assign \new_[37789]_  = ~A266 & ~A265;
  assign \new_[37790]_  = ~A235 & \new_[37789]_ ;
  assign \new_[37793]_  = ~A300 & ~A268;
  assign \new_[37796]_  = ~A302 & ~A301;
  assign \new_[37797]_  = \new_[37796]_  & \new_[37793]_ ;
  assign \new_[37798]_  = \new_[37797]_  & \new_[37790]_ ;
  assign \new_[37802]_  = ~A168 & ~A169;
  assign \new_[37803]_  = ~A170 & \new_[37802]_ ;
  assign \new_[37806]_  = A201 & A200;
  assign \new_[37809]_  = ~A233 & ~A232;
  assign \new_[37810]_  = \new_[37809]_  & \new_[37806]_ ;
  assign \new_[37811]_  = \new_[37810]_  & \new_[37803]_ ;
  assign \new_[37815]_  = ~A266 & ~A265;
  assign \new_[37816]_  = ~A235 & \new_[37815]_ ;
  assign \new_[37819]_  = ~A298 & ~A268;
  assign \new_[37822]_  = ~A301 & ~A299;
  assign \new_[37823]_  = \new_[37822]_  & \new_[37819]_ ;
  assign \new_[37824]_  = \new_[37823]_  & \new_[37816]_ ;
  assign \new_[37828]_  = ~A201 & A166;
  assign \new_[37829]_  = A168 & \new_[37828]_ ;
  assign \new_[37832]_  = ~A203 & ~A202;
  assign \new_[37835]_  = ~A235 & ~A234;
  assign \new_[37836]_  = \new_[37835]_  & \new_[37832]_ ;
  assign \new_[37837]_  = \new_[37836]_  & \new_[37829]_ ;
  assign \new_[37840]_  = ~A267 & ~A236;
  assign \new_[37843]_  = ~A269 & ~A268;
  assign \new_[37844]_  = \new_[37843]_  & \new_[37840]_ ;
  assign \new_[37847]_  = A299 & A298;
  assign \new_[37850]_  = ~A301 & ~A300;
  assign \new_[37851]_  = \new_[37850]_  & \new_[37847]_ ;
  assign \new_[37852]_  = \new_[37851]_  & \new_[37844]_ ;
  assign \new_[37856]_  = ~A201 & A166;
  assign \new_[37857]_  = A168 & \new_[37856]_ ;
  assign \new_[37860]_  = ~A203 & ~A202;
  assign \new_[37863]_  = ~A235 & ~A234;
  assign \new_[37864]_  = \new_[37863]_  & \new_[37860]_ ;
  assign \new_[37865]_  = \new_[37864]_  & \new_[37857]_ ;
  assign \new_[37868]_  = A265 & ~A236;
  assign \new_[37871]_  = ~A267 & A266;
  assign \new_[37872]_  = \new_[37871]_  & \new_[37868]_ ;
  assign \new_[37875]_  = ~A300 & ~A268;
  assign \new_[37878]_  = ~A302 & ~A301;
  assign \new_[37879]_  = \new_[37878]_  & \new_[37875]_ ;
  assign \new_[37880]_  = \new_[37879]_  & \new_[37872]_ ;
  assign \new_[37884]_  = ~A201 & A166;
  assign \new_[37885]_  = A168 & \new_[37884]_ ;
  assign \new_[37888]_  = ~A203 & ~A202;
  assign \new_[37891]_  = ~A235 & ~A234;
  assign \new_[37892]_  = \new_[37891]_  & \new_[37888]_ ;
  assign \new_[37893]_  = \new_[37892]_  & \new_[37885]_ ;
  assign \new_[37896]_  = A265 & ~A236;
  assign \new_[37899]_  = ~A267 & A266;
  assign \new_[37900]_  = \new_[37899]_  & \new_[37896]_ ;
  assign \new_[37903]_  = ~A298 & ~A268;
  assign \new_[37906]_  = ~A301 & ~A299;
  assign \new_[37907]_  = \new_[37906]_  & \new_[37903]_ ;
  assign \new_[37908]_  = \new_[37907]_  & \new_[37900]_ ;
  assign \new_[37912]_  = ~A201 & A166;
  assign \new_[37913]_  = A168 & \new_[37912]_ ;
  assign \new_[37916]_  = ~A203 & ~A202;
  assign \new_[37919]_  = ~A235 & ~A234;
  assign \new_[37920]_  = \new_[37919]_  & \new_[37916]_ ;
  assign \new_[37921]_  = \new_[37920]_  & \new_[37913]_ ;
  assign \new_[37924]_  = ~A265 & ~A236;
  assign \new_[37927]_  = ~A268 & ~A266;
  assign \new_[37928]_  = \new_[37927]_  & \new_[37924]_ ;
  assign \new_[37931]_  = A299 & A298;
  assign \new_[37934]_  = ~A301 & ~A300;
  assign \new_[37935]_  = \new_[37934]_  & \new_[37931]_ ;
  assign \new_[37936]_  = \new_[37935]_  & \new_[37928]_ ;
  assign \new_[37940]_  = ~A201 & A166;
  assign \new_[37941]_  = A168 & \new_[37940]_ ;
  assign \new_[37944]_  = ~A203 & ~A202;
  assign \new_[37947]_  = A233 & A232;
  assign \new_[37948]_  = \new_[37947]_  & \new_[37944]_ ;
  assign \new_[37949]_  = \new_[37948]_  & \new_[37941]_ ;
  assign \new_[37952]_  = ~A235 & ~A234;
  assign \new_[37955]_  = ~A268 & ~A267;
  assign \new_[37956]_  = \new_[37955]_  & \new_[37952]_ ;
  assign \new_[37959]_  = ~A300 & ~A269;
  assign \new_[37962]_  = ~A302 & ~A301;
  assign \new_[37963]_  = \new_[37962]_  & \new_[37959]_ ;
  assign \new_[37964]_  = \new_[37963]_  & \new_[37956]_ ;
  assign \new_[37968]_  = ~A201 & A166;
  assign \new_[37969]_  = A168 & \new_[37968]_ ;
  assign \new_[37972]_  = ~A203 & ~A202;
  assign \new_[37975]_  = A233 & A232;
  assign \new_[37976]_  = \new_[37975]_  & \new_[37972]_ ;
  assign \new_[37977]_  = \new_[37976]_  & \new_[37969]_ ;
  assign \new_[37980]_  = ~A235 & ~A234;
  assign \new_[37983]_  = ~A268 & ~A267;
  assign \new_[37984]_  = \new_[37983]_  & \new_[37980]_ ;
  assign \new_[37987]_  = ~A298 & ~A269;
  assign \new_[37990]_  = ~A301 & ~A299;
  assign \new_[37991]_  = \new_[37990]_  & \new_[37987]_ ;
  assign \new_[37992]_  = \new_[37991]_  & \new_[37984]_ ;
  assign \new_[37996]_  = ~A201 & A166;
  assign \new_[37997]_  = A168 & \new_[37996]_ ;
  assign \new_[38000]_  = ~A203 & ~A202;
  assign \new_[38003]_  = A233 & A232;
  assign \new_[38004]_  = \new_[38003]_  & \new_[38000]_ ;
  assign \new_[38005]_  = \new_[38004]_  & \new_[37997]_ ;
  assign \new_[38008]_  = ~A235 & ~A234;
  assign \new_[38011]_  = ~A266 & ~A265;
  assign \new_[38012]_  = \new_[38011]_  & \new_[38008]_ ;
  assign \new_[38015]_  = ~A300 & ~A268;
  assign \new_[38018]_  = ~A302 & ~A301;
  assign \new_[38019]_  = \new_[38018]_  & \new_[38015]_ ;
  assign \new_[38020]_  = \new_[38019]_  & \new_[38012]_ ;
  assign \new_[38024]_  = ~A201 & A166;
  assign \new_[38025]_  = A168 & \new_[38024]_ ;
  assign \new_[38028]_  = ~A203 & ~A202;
  assign \new_[38031]_  = A233 & A232;
  assign \new_[38032]_  = \new_[38031]_  & \new_[38028]_ ;
  assign \new_[38033]_  = \new_[38032]_  & \new_[38025]_ ;
  assign \new_[38036]_  = ~A235 & ~A234;
  assign \new_[38039]_  = ~A266 & ~A265;
  assign \new_[38040]_  = \new_[38039]_  & \new_[38036]_ ;
  assign \new_[38043]_  = ~A298 & ~A268;
  assign \new_[38046]_  = ~A301 & ~A299;
  assign \new_[38047]_  = \new_[38046]_  & \new_[38043]_ ;
  assign \new_[38048]_  = \new_[38047]_  & \new_[38040]_ ;
  assign \new_[38052]_  = ~A201 & A166;
  assign \new_[38053]_  = A168 & \new_[38052]_ ;
  assign \new_[38056]_  = ~A203 & ~A202;
  assign \new_[38059]_  = ~A233 & ~A232;
  assign \new_[38060]_  = \new_[38059]_  & \new_[38056]_ ;
  assign \new_[38061]_  = \new_[38060]_  & \new_[38053]_ ;
  assign \new_[38064]_  = ~A267 & ~A235;
  assign \new_[38067]_  = ~A269 & ~A268;
  assign \new_[38068]_  = \new_[38067]_  & \new_[38064]_ ;
  assign \new_[38071]_  = A299 & A298;
  assign \new_[38074]_  = ~A301 & ~A300;
  assign \new_[38075]_  = \new_[38074]_  & \new_[38071]_ ;
  assign \new_[38076]_  = \new_[38075]_  & \new_[38068]_ ;
  assign \new_[38080]_  = ~A201 & A166;
  assign \new_[38081]_  = A168 & \new_[38080]_ ;
  assign \new_[38084]_  = ~A203 & ~A202;
  assign \new_[38087]_  = ~A233 & ~A232;
  assign \new_[38088]_  = \new_[38087]_  & \new_[38084]_ ;
  assign \new_[38089]_  = \new_[38088]_  & \new_[38081]_ ;
  assign \new_[38092]_  = A265 & ~A235;
  assign \new_[38095]_  = ~A267 & A266;
  assign \new_[38096]_  = \new_[38095]_  & \new_[38092]_ ;
  assign \new_[38099]_  = ~A300 & ~A268;
  assign \new_[38102]_  = ~A302 & ~A301;
  assign \new_[38103]_  = \new_[38102]_  & \new_[38099]_ ;
  assign \new_[38104]_  = \new_[38103]_  & \new_[38096]_ ;
  assign \new_[38108]_  = ~A201 & A166;
  assign \new_[38109]_  = A168 & \new_[38108]_ ;
  assign \new_[38112]_  = ~A203 & ~A202;
  assign \new_[38115]_  = ~A233 & ~A232;
  assign \new_[38116]_  = \new_[38115]_  & \new_[38112]_ ;
  assign \new_[38117]_  = \new_[38116]_  & \new_[38109]_ ;
  assign \new_[38120]_  = A265 & ~A235;
  assign \new_[38123]_  = ~A267 & A266;
  assign \new_[38124]_  = \new_[38123]_  & \new_[38120]_ ;
  assign \new_[38127]_  = ~A298 & ~A268;
  assign \new_[38130]_  = ~A301 & ~A299;
  assign \new_[38131]_  = \new_[38130]_  & \new_[38127]_ ;
  assign \new_[38132]_  = \new_[38131]_  & \new_[38124]_ ;
  assign \new_[38136]_  = ~A201 & A166;
  assign \new_[38137]_  = A168 & \new_[38136]_ ;
  assign \new_[38140]_  = ~A203 & ~A202;
  assign \new_[38143]_  = ~A233 & ~A232;
  assign \new_[38144]_  = \new_[38143]_  & \new_[38140]_ ;
  assign \new_[38145]_  = \new_[38144]_  & \new_[38137]_ ;
  assign \new_[38148]_  = ~A265 & ~A235;
  assign \new_[38151]_  = ~A268 & ~A266;
  assign \new_[38152]_  = \new_[38151]_  & \new_[38148]_ ;
  assign \new_[38155]_  = A299 & A298;
  assign \new_[38158]_  = ~A301 & ~A300;
  assign \new_[38159]_  = \new_[38158]_  & \new_[38155]_ ;
  assign \new_[38160]_  = \new_[38159]_  & \new_[38152]_ ;
  assign \new_[38164]_  = A199 & A166;
  assign \new_[38165]_  = A168 & \new_[38164]_ ;
  assign \new_[38168]_  = ~A201 & A200;
  assign \new_[38171]_  = ~A234 & ~A202;
  assign \new_[38172]_  = \new_[38171]_  & \new_[38168]_ ;
  assign \new_[38173]_  = \new_[38172]_  & \new_[38165]_ ;
  assign \new_[38176]_  = ~A236 & ~A235;
  assign \new_[38179]_  = ~A268 & ~A267;
  assign \new_[38180]_  = \new_[38179]_  & \new_[38176]_ ;
  assign \new_[38183]_  = ~A300 & ~A269;
  assign \new_[38186]_  = ~A302 & ~A301;
  assign \new_[38187]_  = \new_[38186]_  & \new_[38183]_ ;
  assign \new_[38188]_  = \new_[38187]_  & \new_[38180]_ ;
  assign \new_[38192]_  = A199 & A166;
  assign \new_[38193]_  = A168 & \new_[38192]_ ;
  assign \new_[38196]_  = ~A201 & A200;
  assign \new_[38199]_  = ~A234 & ~A202;
  assign \new_[38200]_  = \new_[38199]_  & \new_[38196]_ ;
  assign \new_[38201]_  = \new_[38200]_  & \new_[38193]_ ;
  assign \new_[38204]_  = ~A236 & ~A235;
  assign \new_[38207]_  = ~A268 & ~A267;
  assign \new_[38208]_  = \new_[38207]_  & \new_[38204]_ ;
  assign \new_[38211]_  = ~A298 & ~A269;
  assign \new_[38214]_  = ~A301 & ~A299;
  assign \new_[38215]_  = \new_[38214]_  & \new_[38211]_ ;
  assign \new_[38216]_  = \new_[38215]_  & \new_[38208]_ ;
  assign \new_[38220]_  = A199 & A166;
  assign \new_[38221]_  = A168 & \new_[38220]_ ;
  assign \new_[38224]_  = ~A201 & A200;
  assign \new_[38227]_  = ~A234 & ~A202;
  assign \new_[38228]_  = \new_[38227]_  & \new_[38224]_ ;
  assign \new_[38229]_  = \new_[38228]_  & \new_[38221]_ ;
  assign \new_[38232]_  = ~A236 & ~A235;
  assign \new_[38235]_  = ~A266 & ~A265;
  assign \new_[38236]_  = \new_[38235]_  & \new_[38232]_ ;
  assign \new_[38239]_  = ~A300 & ~A268;
  assign \new_[38242]_  = ~A302 & ~A301;
  assign \new_[38243]_  = \new_[38242]_  & \new_[38239]_ ;
  assign \new_[38244]_  = \new_[38243]_  & \new_[38236]_ ;
  assign \new_[38248]_  = A199 & A166;
  assign \new_[38249]_  = A168 & \new_[38248]_ ;
  assign \new_[38252]_  = ~A201 & A200;
  assign \new_[38255]_  = ~A234 & ~A202;
  assign \new_[38256]_  = \new_[38255]_  & \new_[38252]_ ;
  assign \new_[38257]_  = \new_[38256]_  & \new_[38249]_ ;
  assign \new_[38260]_  = ~A236 & ~A235;
  assign \new_[38263]_  = ~A266 & ~A265;
  assign \new_[38264]_  = \new_[38263]_  & \new_[38260]_ ;
  assign \new_[38267]_  = ~A298 & ~A268;
  assign \new_[38270]_  = ~A301 & ~A299;
  assign \new_[38271]_  = \new_[38270]_  & \new_[38267]_ ;
  assign \new_[38272]_  = \new_[38271]_  & \new_[38264]_ ;
  assign \new_[38276]_  = A199 & A166;
  assign \new_[38277]_  = A168 & \new_[38276]_ ;
  assign \new_[38280]_  = ~A201 & A200;
  assign \new_[38283]_  = ~A232 & ~A202;
  assign \new_[38284]_  = \new_[38283]_  & \new_[38280]_ ;
  assign \new_[38285]_  = \new_[38284]_  & \new_[38277]_ ;
  assign \new_[38288]_  = ~A235 & ~A233;
  assign \new_[38291]_  = ~A268 & ~A267;
  assign \new_[38292]_  = \new_[38291]_  & \new_[38288]_ ;
  assign \new_[38295]_  = ~A300 & ~A269;
  assign \new_[38298]_  = ~A302 & ~A301;
  assign \new_[38299]_  = \new_[38298]_  & \new_[38295]_ ;
  assign \new_[38300]_  = \new_[38299]_  & \new_[38292]_ ;
  assign \new_[38304]_  = A199 & A166;
  assign \new_[38305]_  = A168 & \new_[38304]_ ;
  assign \new_[38308]_  = ~A201 & A200;
  assign \new_[38311]_  = ~A232 & ~A202;
  assign \new_[38312]_  = \new_[38311]_  & \new_[38308]_ ;
  assign \new_[38313]_  = \new_[38312]_  & \new_[38305]_ ;
  assign \new_[38316]_  = ~A235 & ~A233;
  assign \new_[38319]_  = ~A268 & ~A267;
  assign \new_[38320]_  = \new_[38319]_  & \new_[38316]_ ;
  assign \new_[38323]_  = ~A298 & ~A269;
  assign \new_[38326]_  = ~A301 & ~A299;
  assign \new_[38327]_  = \new_[38326]_  & \new_[38323]_ ;
  assign \new_[38328]_  = \new_[38327]_  & \new_[38320]_ ;
  assign \new_[38332]_  = A199 & A166;
  assign \new_[38333]_  = A168 & \new_[38332]_ ;
  assign \new_[38336]_  = ~A201 & A200;
  assign \new_[38339]_  = ~A232 & ~A202;
  assign \new_[38340]_  = \new_[38339]_  & \new_[38336]_ ;
  assign \new_[38341]_  = \new_[38340]_  & \new_[38333]_ ;
  assign \new_[38344]_  = ~A235 & ~A233;
  assign \new_[38347]_  = ~A266 & ~A265;
  assign \new_[38348]_  = \new_[38347]_  & \new_[38344]_ ;
  assign \new_[38351]_  = ~A300 & ~A268;
  assign \new_[38354]_  = ~A302 & ~A301;
  assign \new_[38355]_  = \new_[38354]_  & \new_[38351]_ ;
  assign \new_[38356]_  = \new_[38355]_  & \new_[38348]_ ;
  assign \new_[38360]_  = A199 & A166;
  assign \new_[38361]_  = A168 & \new_[38360]_ ;
  assign \new_[38364]_  = ~A201 & A200;
  assign \new_[38367]_  = ~A232 & ~A202;
  assign \new_[38368]_  = \new_[38367]_  & \new_[38364]_ ;
  assign \new_[38369]_  = \new_[38368]_  & \new_[38361]_ ;
  assign \new_[38372]_  = ~A235 & ~A233;
  assign \new_[38375]_  = ~A266 & ~A265;
  assign \new_[38376]_  = \new_[38375]_  & \new_[38372]_ ;
  assign \new_[38379]_  = ~A298 & ~A268;
  assign \new_[38382]_  = ~A301 & ~A299;
  assign \new_[38383]_  = \new_[38382]_  & \new_[38379]_ ;
  assign \new_[38384]_  = \new_[38383]_  & \new_[38376]_ ;
  assign \new_[38388]_  = ~A199 & A166;
  assign \new_[38389]_  = A168 & \new_[38388]_ ;
  assign \new_[38392]_  = ~A202 & ~A200;
  assign \new_[38395]_  = ~A235 & ~A234;
  assign \new_[38396]_  = \new_[38395]_  & \new_[38392]_ ;
  assign \new_[38397]_  = \new_[38396]_  & \new_[38389]_ ;
  assign \new_[38400]_  = ~A267 & ~A236;
  assign \new_[38403]_  = ~A269 & ~A268;
  assign \new_[38404]_  = \new_[38403]_  & \new_[38400]_ ;
  assign \new_[38407]_  = A299 & A298;
  assign \new_[38410]_  = ~A301 & ~A300;
  assign \new_[38411]_  = \new_[38410]_  & \new_[38407]_ ;
  assign \new_[38412]_  = \new_[38411]_  & \new_[38404]_ ;
  assign \new_[38416]_  = ~A199 & A166;
  assign \new_[38417]_  = A168 & \new_[38416]_ ;
  assign \new_[38420]_  = ~A202 & ~A200;
  assign \new_[38423]_  = ~A235 & ~A234;
  assign \new_[38424]_  = \new_[38423]_  & \new_[38420]_ ;
  assign \new_[38425]_  = \new_[38424]_  & \new_[38417]_ ;
  assign \new_[38428]_  = A265 & ~A236;
  assign \new_[38431]_  = ~A267 & A266;
  assign \new_[38432]_  = \new_[38431]_  & \new_[38428]_ ;
  assign \new_[38435]_  = ~A300 & ~A268;
  assign \new_[38438]_  = ~A302 & ~A301;
  assign \new_[38439]_  = \new_[38438]_  & \new_[38435]_ ;
  assign \new_[38440]_  = \new_[38439]_  & \new_[38432]_ ;
  assign \new_[38444]_  = ~A199 & A166;
  assign \new_[38445]_  = A168 & \new_[38444]_ ;
  assign \new_[38448]_  = ~A202 & ~A200;
  assign \new_[38451]_  = ~A235 & ~A234;
  assign \new_[38452]_  = \new_[38451]_  & \new_[38448]_ ;
  assign \new_[38453]_  = \new_[38452]_  & \new_[38445]_ ;
  assign \new_[38456]_  = A265 & ~A236;
  assign \new_[38459]_  = ~A267 & A266;
  assign \new_[38460]_  = \new_[38459]_  & \new_[38456]_ ;
  assign \new_[38463]_  = ~A298 & ~A268;
  assign \new_[38466]_  = ~A301 & ~A299;
  assign \new_[38467]_  = \new_[38466]_  & \new_[38463]_ ;
  assign \new_[38468]_  = \new_[38467]_  & \new_[38460]_ ;
  assign \new_[38472]_  = ~A199 & A166;
  assign \new_[38473]_  = A168 & \new_[38472]_ ;
  assign \new_[38476]_  = ~A202 & ~A200;
  assign \new_[38479]_  = ~A235 & ~A234;
  assign \new_[38480]_  = \new_[38479]_  & \new_[38476]_ ;
  assign \new_[38481]_  = \new_[38480]_  & \new_[38473]_ ;
  assign \new_[38484]_  = ~A265 & ~A236;
  assign \new_[38487]_  = ~A268 & ~A266;
  assign \new_[38488]_  = \new_[38487]_  & \new_[38484]_ ;
  assign \new_[38491]_  = A299 & A298;
  assign \new_[38494]_  = ~A301 & ~A300;
  assign \new_[38495]_  = \new_[38494]_  & \new_[38491]_ ;
  assign \new_[38496]_  = \new_[38495]_  & \new_[38488]_ ;
  assign \new_[38500]_  = ~A199 & A166;
  assign \new_[38501]_  = A168 & \new_[38500]_ ;
  assign \new_[38504]_  = ~A202 & ~A200;
  assign \new_[38507]_  = A233 & A232;
  assign \new_[38508]_  = \new_[38507]_  & \new_[38504]_ ;
  assign \new_[38509]_  = \new_[38508]_  & \new_[38501]_ ;
  assign \new_[38512]_  = ~A235 & ~A234;
  assign \new_[38515]_  = ~A268 & ~A267;
  assign \new_[38516]_  = \new_[38515]_  & \new_[38512]_ ;
  assign \new_[38519]_  = ~A300 & ~A269;
  assign \new_[38522]_  = ~A302 & ~A301;
  assign \new_[38523]_  = \new_[38522]_  & \new_[38519]_ ;
  assign \new_[38524]_  = \new_[38523]_  & \new_[38516]_ ;
  assign \new_[38528]_  = ~A199 & A166;
  assign \new_[38529]_  = A168 & \new_[38528]_ ;
  assign \new_[38532]_  = ~A202 & ~A200;
  assign \new_[38535]_  = A233 & A232;
  assign \new_[38536]_  = \new_[38535]_  & \new_[38532]_ ;
  assign \new_[38537]_  = \new_[38536]_  & \new_[38529]_ ;
  assign \new_[38540]_  = ~A235 & ~A234;
  assign \new_[38543]_  = ~A268 & ~A267;
  assign \new_[38544]_  = \new_[38543]_  & \new_[38540]_ ;
  assign \new_[38547]_  = ~A298 & ~A269;
  assign \new_[38550]_  = ~A301 & ~A299;
  assign \new_[38551]_  = \new_[38550]_  & \new_[38547]_ ;
  assign \new_[38552]_  = \new_[38551]_  & \new_[38544]_ ;
  assign \new_[38556]_  = ~A199 & A166;
  assign \new_[38557]_  = A168 & \new_[38556]_ ;
  assign \new_[38560]_  = ~A202 & ~A200;
  assign \new_[38563]_  = A233 & A232;
  assign \new_[38564]_  = \new_[38563]_  & \new_[38560]_ ;
  assign \new_[38565]_  = \new_[38564]_  & \new_[38557]_ ;
  assign \new_[38568]_  = ~A235 & ~A234;
  assign \new_[38571]_  = ~A266 & ~A265;
  assign \new_[38572]_  = \new_[38571]_  & \new_[38568]_ ;
  assign \new_[38575]_  = ~A300 & ~A268;
  assign \new_[38578]_  = ~A302 & ~A301;
  assign \new_[38579]_  = \new_[38578]_  & \new_[38575]_ ;
  assign \new_[38580]_  = \new_[38579]_  & \new_[38572]_ ;
  assign \new_[38584]_  = ~A199 & A166;
  assign \new_[38585]_  = A168 & \new_[38584]_ ;
  assign \new_[38588]_  = ~A202 & ~A200;
  assign \new_[38591]_  = A233 & A232;
  assign \new_[38592]_  = \new_[38591]_  & \new_[38588]_ ;
  assign \new_[38593]_  = \new_[38592]_  & \new_[38585]_ ;
  assign \new_[38596]_  = ~A235 & ~A234;
  assign \new_[38599]_  = ~A266 & ~A265;
  assign \new_[38600]_  = \new_[38599]_  & \new_[38596]_ ;
  assign \new_[38603]_  = ~A298 & ~A268;
  assign \new_[38606]_  = ~A301 & ~A299;
  assign \new_[38607]_  = \new_[38606]_  & \new_[38603]_ ;
  assign \new_[38608]_  = \new_[38607]_  & \new_[38600]_ ;
  assign \new_[38612]_  = ~A199 & A166;
  assign \new_[38613]_  = A168 & \new_[38612]_ ;
  assign \new_[38616]_  = ~A202 & ~A200;
  assign \new_[38619]_  = ~A233 & ~A232;
  assign \new_[38620]_  = \new_[38619]_  & \new_[38616]_ ;
  assign \new_[38621]_  = \new_[38620]_  & \new_[38613]_ ;
  assign \new_[38624]_  = ~A267 & ~A235;
  assign \new_[38627]_  = ~A269 & ~A268;
  assign \new_[38628]_  = \new_[38627]_  & \new_[38624]_ ;
  assign \new_[38631]_  = A299 & A298;
  assign \new_[38634]_  = ~A301 & ~A300;
  assign \new_[38635]_  = \new_[38634]_  & \new_[38631]_ ;
  assign \new_[38636]_  = \new_[38635]_  & \new_[38628]_ ;
  assign \new_[38640]_  = ~A199 & A166;
  assign \new_[38641]_  = A168 & \new_[38640]_ ;
  assign \new_[38644]_  = ~A202 & ~A200;
  assign \new_[38647]_  = ~A233 & ~A232;
  assign \new_[38648]_  = \new_[38647]_  & \new_[38644]_ ;
  assign \new_[38649]_  = \new_[38648]_  & \new_[38641]_ ;
  assign \new_[38652]_  = A265 & ~A235;
  assign \new_[38655]_  = ~A267 & A266;
  assign \new_[38656]_  = \new_[38655]_  & \new_[38652]_ ;
  assign \new_[38659]_  = ~A300 & ~A268;
  assign \new_[38662]_  = ~A302 & ~A301;
  assign \new_[38663]_  = \new_[38662]_  & \new_[38659]_ ;
  assign \new_[38664]_  = \new_[38663]_  & \new_[38656]_ ;
  assign \new_[38668]_  = ~A199 & A166;
  assign \new_[38669]_  = A168 & \new_[38668]_ ;
  assign \new_[38672]_  = ~A202 & ~A200;
  assign \new_[38675]_  = ~A233 & ~A232;
  assign \new_[38676]_  = \new_[38675]_  & \new_[38672]_ ;
  assign \new_[38677]_  = \new_[38676]_  & \new_[38669]_ ;
  assign \new_[38680]_  = A265 & ~A235;
  assign \new_[38683]_  = ~A267 & A266;
  assign \new_[38684]_  = \new_[38683]_  & \new_[38680]_ ;
  assign \new_[38687]_  = ~A298 & ~A268;
  assign \new_[38690]_  = ~A301 & ~A299;
  assign \new_[38691]_  = \new_[38690]_  & \new_[38687]_ ;
  assign \new_[38692]_  = \new_[38691]_  & \new_[38684]_ ;
  assign \new_[38696]_  = ~A199 & A166;
  assign \new_[38697]_  = A168 & \new_[38696]_ ;
  assign \new_[38700]_  = ~A202 & ~A200;
  assign \new_[38703]_  = ~A233 & ~A232;
  assign \new_[38704]_  = \new_[38703]_  & \new_[38700]_ ;
  assign \new_[38705]_  = \new_[38704]_  & \new_[38697]_ ;
  assign \new_[38708]_  = ~A265 & ~A235;
  assign \new_[38711]_  = ~A268 & ~A266;
  assign \new_[38712]_  = \new_[38711]_  & \new_[38708]_ ;
  assign \new_[38715]_  = A299 & A298;
  assign \new_[38718]_  = ~A301 & ~A300;
  assign \new_[38719]_  = \new_[38718]_  & \new_[38715]_ ;
  assign \new_[38720]_  = \new_[38719]_  & \new_[38712]_ ;
  assign \new_[38724]_  = ~A201 & A167;
  assign \new_[38725]_  = A168 & \new_[38724]_ ;
  assign \new_[38728]_  = ~A203 & ~A202;
  assign \new_[38731]_  = ~A235 & ~A234;
  assign \new_[38732]_  = \new_[38731]_  & \new_[38728]_ ;
  assign \new_[38733]_  = \new_[38732]_  & \new_[38725]_ ;
  assign \new_[38736]_  = ~A267 & ~A236;
  assign \new_[38739]_  = ~A269 & ~A268;
  assign \new_[38740]_  = \new_[38739]_  & \new_[38736]_ ;
  assign \new_[38743]_  = A299 & A298;
  assign \new_[38746]_  = ~A301 & ~A300;
  assign \new_[38747]_  = \new_[38746]_  & \new_[38743]_ ;
  assign \new_[38748]_  = \new_[38747]_  & \new_[38740]_ ;
  assign \new_[38752]_  = ~A201 & A167;
  assign \new_[38753]_  = A168 & \new_[38752]_ ;
  assign \new_[38756]_  = ~A203 & ~A202;
  assign \new_[38759]_  = ~A235 & ~A234;
  assign \new_[38760]_  = \new_[38759]_  & \new_[38756]_ ;
  assign \new_[38761]_  = \new_[38760]_  & \new_[38753]_ ;
  assign \new_[38764]_  = A265 & ~A236;
  assign \new_[38767]_  = ~A267 & A266;
  assign \new_[38768]_  = \new_[38767]_  & \new_[38764]_ ;
  assign \new_[38771]_  = ~A300 & ~A268;
  assign \new_[38774]_  = ~A302 & ~A301;
  assign \new_[38775]_  = \new_[38774]_  & \new_[38771]_ ;
  assign \new_[38776]_  = \new_[38775]_  & \new_[38768]_ ;
  assign \new_[38780]_  = ~A201 & A167;
  assign \new_[38781]_  = A168 & \new_[38780]_ ;
  assign \new_[38784]_  = ~A203 & ~A202;
  assign \new_[38787]_  = ~A235 & ~A234;
  assign \new_[38788]_  = \new_[38787]_  & \new_[38784]_ ;
  assign \new_[38789]_  = \new_[38788]_  & \new_[38781]_ ;
  assign \new_[38792]_  = A265 & ~A236;
  assign \new_[38795]_  = ~A267 & A266;
  assign \new_[38796]_  = \new_[38795]_  & \new_[38792]_ ;
  assign \new_[38799]_  = ~A298 & ~A268;
  assign \new_[38802]_  = ~A301 & ~A299;
  assign \new_[38803]_  = \new_[38802]_  & \new_[38799]_ ;
  assign \new_[38804]_  = \new_[38803]_  & \new_[38796]_ ;
  assign \new_[38808]_  = ~A201 & A167;
  assign \new_[38809]_  = A168 & \new_[38808]_ ;
  assign \new_[38812]_  = ~A203 & ~A202;
  assign \new_[38815]_  = ~A235 & ~A234;
  assign \new_[38816]_  = \new_[38815]_  & \new_[38812]_ ;
  assign \new_[38817]_  = \new_[38816]_  & \new_[38809]_ ;
  assign \new_[38820]_  = ~A265 & ~A236;
  assign \new_[38823]_  = ~A268 & ~A266;
  assign \new_[38824]_  = \new_[38823]_  & \new_[38820]_ ;
  assign \new_[38827]_  = A299 & A298;
  assign \new_[38830]_  = ~A301 & ~A300;
  assign \new_[38831]_  = \new_[38830]_  & \new_[38827]_ ;
  assign \new_[38832]_  = \new_[38831]_  & \new_[38824]_ ;
  assign \new_[38836]_  = ~A201 & A167;
  assign \new_[38837]_  = A168 & \new_[38836]_ ;
  assign \new_[38840]_  = ~A203 & ~A202;
  assign \new_[38843]_  = A233 & A232;
  assign \new_[38844]_  = \new_[38843]_  & \new_[38840]_ ;
  assign \new_[38845]_  = \new_[38844]_  & \new_[38837]_ ;
  assign \new_[38848]_  = ~A235 & ~A234;
  assign \new_[38851]_  = ~A268 & ~A267;
  assign \new_[38852]_  = \new_[38851]_  & \new_[38848]_ ;
  assign \new_[38855]_  = ~A300 & ~A269;
  assign \new_[38858]_  = ~A302 & ~A301;
  assign \new_[38859]_  = \new_[38858]_  & \new_[38855]_ ;
  assign \new_[38860]_  = \new_[38859]_  & \new_[38852]_ ;
  assign \new_[38864]_  = ~A201 & A167;
  assign \new_[38865]_  = A168 & \new_[38864]_ ;
  assign \new_[38868]_  = ~A203 & ~A202;
  assign \new_[38871]_  = A233 & A232;
  assign \new_[38872]_  = \new_[38871]_  & \new_[38868]_ ;
  assign \new_[38873]_  = \new_[38872]_  & \new_[38865]_ ;
  assign \new_[38876]_  = ~A235 & ~A234;
  assign \new_[38879]_  = ~A268 & ~A267;
  assign \new_[38880]_  = \new_[38879]_  & \new_[38876]_ ;
  assign \new_[38883]_  = ~A298 & ~A269;
  assign \new_[38886]_  = ~A301 & ~A299;
  assign \new_[38887]_  = \new_[38886]_  & \new_[38883]_ ;
  assign \new_[38888]_  = \new_[38887]_  & \new_[38880]_ ;
  assign \new_[38892]_  = ~A201 & A167;
  assign \new_[38893]_  = A168 & \new_[38892]_ ;
  assign \new_[38896]_  = ~A203 & ~A202;
  assign \new_[38899]_  = A233 & A232;
  assign \new_[38900]_  = \new_[38899]_  & \new_[38896]_ ;
  assign \new_[38901]_  = \new_[38900]_  & \new_[38893]_ ;
  assign \new_[38904]_  = ~A235 & ~A234;
  assign \new_[38907]_  = ~A266 & ~A265;
  assign \new_[38908]_  = \new_[38907]_  & \new_[38904]_ ;
  assign \new_[38911]_  = ~A300 & ~A268;
  assign \new_[38914]_  = ~A302 & ~A301;
  assign \new_[38915]_  = \new_[38914]_  & \new_[38911]_ ;
  assign \new_[38916]_  = \new_[38915]_  & \new_[38908]_ ;
  assign \new_[38920]_  = ~A201 & A167;
  assign \new_[38921]_  = A168 & \new_[38920]_ ;
  assign \new_[38924]_  = ~A203 & ~A202;
  assign \new_[38927]_  = A233 & A232;
  assign \new_[38928]_  = \new_[38927]_  & \new_[38924]_ ;
  assign \new_[38929]_  = \new_[38928]_  & \new_[38921]_ ;
  assign \new_[38932]_  = ~A235 & ~A234;
  assign \new_[38935]_  = ~A266 & ~A265;
  assign \new_[38936]_  = \new_[38935]_  & \new_[38932]_ ;
  assign \new_[38939]_  = ~A298 & ~A268;
  assign \new_[38942]_  = ~A301 & ~A299;
  assign \new_[38943]_  = \new_[38942]_  & \new_[38939]_ ;
  assign \new_[38944]_  = \new_[38943]_  & \new_[38936]_ ;
  assign \new_[38948]_  = ~A201 & A167;
  assign \new_[38949]_  = A168 & \new_[38948]_ ;
  assign \new_[38952]_  = ~A203 & ~A202;
  assign \new_[38955]_  = ~A233 & ~A232;
  assign \new_[38956]_  = \new_[38955]_  & \new_[38952]_ ;
  assign \new_[38957]_  = \new_[38956]_  & \new_[38949]_ ;
  assign \new_[38960]_  = ~A267 & ~A235;
  assign \new_[38963]_  = ~A269 & ~A268;
  assign \new_[38964]_  = \new_[38963]_  & \new_[38960]_ ;
  assign \new_[38967]_  = A299 & A298;
  assign \new_[38970]_  = ~A301 & ~A300;
  assign \new_[38971]_  = \new_[38970]_  & \new_[38967]_ ;
  assign \new_[38972]_  = \new_[38971]_  & \new_[38964]_ ;
  assign \new_[38976]_  = ~A201 & A167;
  assign \new_[38977]_  = A168 & \new_[38976]_ ;
  assign \new_[38980]_  = ~A203 & ~A202;
  assign \new_[38983]_  = ~A233 & ~A232;
  assign \new_[38984]_  = \new_[38983]_  & \new_[38980]_ ;
  assign \new_[38985]_  = \new_[38984]_  & \new_[38977]_ ;
  assign \new_[38988]_  = A265 & ~A235;
  assign \new_[38991]_  = ~A267 & A266;
  assign \new_[38992]_  = \new_[38991]_  & \new_[38988]_ ;
  assign \new_[38995]_  = ~A300 & ~A268;
  assign \new_[38998]_  = ~A302 & ~A301;
  assign \new_[38999]_  = \new_[38998]_  & \new_[38995]_ ;
  assign \new_[39000]_  = \new_[38999]_  & \new_[38992]_ ;
  assign \new_[39004]_  = ~A201 & A167;
  assign \new_[39005]_  = A168 & \new_[39004]_ ;
  assign \new_[39008]_  = ~A203 & ~A202;
  assign \new_[39011]_  = ~A233 & ~A232;
  assign \new_[39012]_  = \new_[39011]_  & \new_[39008]_ ;
  assign \new_[39013]_  = \new_[39012]_  & \new_[39005]_ ;
  assign \new_[39016]_  = A265 & ~A235;
  assign \new_[39019]_  = ~A267 & A266;
  assign \new_[39020]_  = \new_[39019]_  & \new_[39016]_ ;
  assign \new_[39023]_  = ~A298 & ~A268;
  assign \new_[39026]_  = ~A301 & ~A299;
  assign \new_[39027]_  = \new_[39026]_  & \new_[39023]_ ;
  assign \new_[39028]_  = \new_[39027]_  & \new_[39020]_ ;
  assign \new_[39032]_  = ~A201 & A167;
  assign \new_[39033]_  = A168 & \new_[39032]_ ;
  assign \new_[39036]_  = ~A203 & ~A202;
  assign \new_[39039]_  = ~A233 & ~A232;
  assign \new_[39040]_  = \new_[39039]_  & \new_[39036]_ ;
  assign \new_[39041]_  = \new_[39040]_  & \new_[39033]_ ;
  assign \new_[39044]_  = ~A265 & ~A235;
  assign \new_[39047]_  = ~A268 & ~A266;
  assign \new_[39048]_  = \new_[39047]_  & \new_[39044]_ ;
  assign \new_[39051]_  = A299 & A298;
  assign \new_[39054]_  = ~A301 & ~A300;
  assign \new_[39055]_  = \new_[39054]_  & \new_[39051]_ ;
  assign \new_[39056]_  = \new_[39055]_  & \new_[39048]_ ;
  assign \new_[39060]_  = A199 & A167;
  assign \new_[39061]_  = A168 & \new_[39060]_ ;
  assign \new_[39064]_  = ~A201 & A200;
  assign \new_[39067]_  = ~A234 & ~A202;
  assign \new_[39068]_  = \new_[39067]_  & \new_[39064]_ ;
  assign \new_[39069]_  = \new_[39068]_  & \new_[39061]_ ;
  assign \new_[39072]_  = ~A236 & ~A235;
  assign \new_[39075]_  = ~A268 & ~A267;
  assign \new_[39076]_  = \new_[39075]_  & \new_[39072]_ ;
  assign \new_[39079]_  = ~A300 & ~A269;
  assign \new_[39082]_  = ~A302 & ~A301;
  assign \new_[39083]_  = \new_[39082]_  & \new_[39079]_ ;
  assign \new_[39084]_  = \new_[39083]_  & \new_[39076]_ ;
  assign \new_[39088]_  = A199 & A167;
  assign \new_[39089]_  = A168 & \new_[39088]_ ;
  assign \new_[39092]_  = ~A201 & A200;
  assign \new_[39095]_  = ~A234 & ~A202;
  assign \new_[39096]_  = \new_[39095]_  & \new_[39092]_ ;
  assign \new_[39097]_  = \new_[39096]_  & \new_[39089]_ ;
  assign \new_[39100]_  = ~A236 & ~A235;
  assign \new_[39103]_  = ~A268 & ~A267;
  assign \new_[39104]_  = \new_[39103]_  & \new_[39100]_ ;
  assign \new_[39107]_  = ~A298 & ~A269;
  assign \new_[39110]_  = ~A301 & ~A299;
  assign \new_[39111]_  = \new_[39110]_  & \new_[39107]_ ;
  assign \new_[39112]_  = \new_[39111]_  & \new_[39104]_ ;
  assign \new_[39116]_  = A199 & A167;
  assign \new_[39117]_  = A168 & \new_[39116]_ ;
  assign \new_[39120]_  = ~A201 & A200;
  assign \new_[39123]_  = ~A234 & ~A202;
  assign \new_[39124]_  = \new_[39123]_  & \new_[39120]_ ;
  assign \new_[39125]_  = \new_[39124]_  & \new_[39117]_ ;
  assign \new_[39128]_  = ~A236 & ~A235;
  assign \new_[39131]_  = ~A266 & ~A265;
  assign \new_[39132]_  = \new_[39131]_  & \new_[39128]_ ;
  assign \new_[39135]_  = ~A300 & ~A268;
  assign \new_[39138]_  = ~A302 & ~A301;
  assign \new_[39139]_  = \new_[39138]_  & \new_[39135]_ ;
  assign \new_[39140]_  = \new_[39139]_  & \new_[39132]_ ;
  assign \new_[39144]_  = A199 & A167;
  assign \new_[39145]_  = A168 & \new_[39144]_ ;
  assign \new_[39148]_  = ~A201 & A200;
  assign \new_[39151]_  = ~A234 & ~A202;
  assign \new_[39152]_  = \new_[39151]_  & \new_[39148]_ ;
  assign \new_[39153]_  = \new_[39152]_  & \new_[39145]_ ;
  assign \new_[39156]_  = ~A236 & ~A235;
  assign \new_[39159]_  = ~A266 & ~A265;
  assign \new_[39160]_  = \new_[39159]_  & \new_[39156]_ ;
  assign \new_[39163]_  = ~A298 & ~A268;
  assign \new_[39166]_  = ~A301 & ~A299;
  assign \new_[39167]_  = \new_[39166]_  & \new_[39163]_ ;
  assign \new_[39168]_  = \new_[39167]_  & \new_[39160]_ ;
  assign \new_[39172]_  = A199 & A167;
  assign \new_[39173]_  = A168 & \new_[39172]_ ;
  assign \new_[39176]_  = ~A201 & A200;
  assign \new_[39179]_  = ~A232 & ~A202;
  assign \new_[39180]_  = \new_[39179]_  & \new_[39176]_ ;
  assign \new_[39181]_  = \new_[39180]_  & \new_[39173]_ ;
  assign \new_[39184]_  = ~A235 & ~A233;
  assign \new_[39187]_  = ~A268 & ~A267;
  assign \new_[39188]_  = \new_[39187]_  & \new_[39184]_ ;
  assign \new_[39191]_  = ~A300 & ~A269;
  assign \new_[39194]_  = ~A302 & ~A301;
  assign \new_[39195]_  = \new_[39194]_  & \new_[39191]_ ;
  assign \new_[39196]_  = \new_[39195]_  & \new_[39188]_ ;
  assign \new_[39200]_  = A199 & A167;
  assign \new_[39201]_  = A168 & \new_[39200]_ ;
  assign \new_[39204]_  = ~A201 & A200;
  assign \new_[39207]_  = ~A232 & ~A202;
  assign \new_[39208]_  = \new_[39207]_  & \new_[39204]_ ;
  assign \new_[39209]_  = \new_[39208]_  & \new_[39201]_ ;
  assign \new_[39212]_  = ~A235 & ~A233;
  assign \new_[39215]_  = ~A268 & ~A267;
  assign \new_[39216]_  = \new_[39215]_  & \new_[39212]_ ;
  assign \new_[39219]_  = ~A298 & ~A269;
  assign \new_[39222]_  = ~A301 & ~A299;
  assign \new_[39223]_  = \new_[39222]_  & \new_[39219]_ ;
  assign \new_[39224]_  = \new_[39223]_  & \new_[39216]_ ;
  assign \new_[39228]_  = A199 & A167;
  assign \new_[39229]_  = A168 & \new_[39228]_ ;
  assign \new_[39232]_  = ~A201 & A200;
  assign \new_[39235]_  = ~A232 & ~A202;
  assign \new_[39236]_  = \new_[39235]_  & \new_[39232]_ ;
  assign \new_[39237]_  = \new_[39236]_  & \new_[39229]_ ;
  assign \new_[39240]_  = ~A235 & ~A233;
  assign \new_[39243]_  = ~A266 & ~A265;
  assign \new_[39244]_  = \new_[39243]_  & \new_[39240]_ ;
  assign \new_[39247]_  = ~A300 & ~A268;
  assign \new_[39250]_  = ~A302 & ~A301;
  assign \new_[39251]_  = \new_[39250]_  & \new_[39247]_ ;
  assign \new_[39252]_  = \new_[39251]_  & \new_[39244]_ ;
  assign \new_[39256]_  = A199 & A167;
  assign \new_[39257]_  = A168 & \new_[39256]_ ;
  assign \new_[39260]_  = ~A201 & A200;
  assign \new_[39263]_  = ~A232 & ~A202;
  assign \new_[39264]_  = \new_[39263]_  & \new_[39260]_ ;
  assign \new_[39265]_  = \new_[39264]_  & \new_[39257]_ ;
  assign \new_[39268]_  = ~A235 & ~A233;
  assign \new_[39271]_  = ~A266 & ~A265;
  assign \new_[39272]_  = \new_[39271]_  & \new_[39268]_ ;
  assign \new_[39275]_  = ~A298 & ~A268;
  assign \new_[39278]_  = ~A301 & ~A299;
  assign \new_[39279]_  = \new_[39278]_  & \new_[39275]_ ;
  assign \new_[39280]_  = \new_[39279]_  & \new_[39272]_ ;
  assign \new_[39284]_  = ~A199 & A167;
  assign \new_[39285]_  = A168 & \new_[39284]_ ;
  assign \new_[39288]_  = ~A202 & ~A200;
  assign \new_[39291]_  = ~A235 & ~A234;
  assign \new_[39292]_  = \new_[39291]_  & \new_[39288]_ ;
  assign \new_[39293]_  = \new_[39292]_  & \new_[39285]_ ;
  assign \new_[39296]_  = ~A267 & ~A236;
  assign \new_[39299]_  = ~A269 & ~A268;
  assign \new_[39300]_  = \new_[39299]_  & \new_[39296]_ ;
  assign \new_[39303]_  = A299 & A298;
  assign \new_[39306]_  = ~A301 & ~A300;
  assign \new_[39307]_  = \new_[39306]_  & \new_[39303]_ ;
  assign \new_[39308]_  = \new_[39307]_  & \new_[39300]_ ;
  assign \new_[39312]_  = ~A199 & A167;
  assign \new_[39313]_  = A168 & \new_[39312]_ ;
  assign \new_[39316]_  = ~A202 & ~A200;
  assign \new_[39319]_  = ~A235 & ~A234;
  assign \new_[39320]_  = \new_[39319]_  & \new_[39316]_ ;
  assign \new_[39321]_  = \new_[39320]_  & \new_[39313]_ ;
  assign \new_[39324]_  = A265 & ~A236;
  assign \new_[39327]_  = ~A267 & A266;
  assign \new_[39328]_  = \new_[39327]_  & \new_[39324]_ ;
  assign \new_[39331]_  = ~A300 & ~A268;
  assign \new_[39334]_  = ~A302 & ~A301;
  assign \new_[39335]_  = \new_[39334]_  & \new_[39331]_ ;
  assign \new_[39336]_  = \new_[39335]_  & \new_[39328]_ ;
  assign \new_[39340]_  = ~A199 & A167;
  assign \new_[39341]_  = A168 & \new_[39340]_ ;
  assign \new_[39344]_  = ~A202 & ~A200;
  assign \new_[39347]_  = ~A235 & ~A234;
  assign \new_[39348]_  = \new_[39347]_  & \new_[39344]_ ;
  assign \new_[39349]_  = \new_[39348]_  & \new_[39341]_ ;
  assign \new_[39352]_  = A265 & ~A236;
  assign \new_[39355]_  = ~A267 & A266;
  assign \new_[39356]_  = \new_[39355]_  & \new_[39352]_ ;
  assign \new_[39359]_  = ~A298 & ~A268;
  assign \new_[39362]_  = ~A301 & ~A299;
  assign \new_[39363]_  = \new_[39362]_  & \new_[39359]_ ;
  assign \new_[39364]_  = \new_[39363]_  & \new_[39356]_ ;
  assign \new_[39368]_  = ~A199 & A167;
  assign \new_[39369]_  = A168 & \new_[39368]_ ;
  assign \new_[39372]_  = ~A202 & ~A200;
  assign \new_[39375]_  = ~A235 & ~A234;
  assign \new_[39376]_  = \new_[39375]_  & \new_[39372]_ ;
  assign \new_[39377]_  = \new_[39376]_  & \new_[39369]_ ;
  assign \new_[39380]_  = ~A265 & ~A236;
  assign \new_[39383]_  = ~A268 & ~A266;
  assign \new_[39384]_  = \new_[39383]_  & \new_[39380]_ ;
  assign \new_[39387]_  = A299 & A298;
  assign \new_[39390]_  = ~A301 & ~A300;
  assign \new_[39391]_  = \new_[39390]_  & \new_[39387]_ ;
  assign \new_[39392]_  = \new_[39391]_  & \new_[39384]_ ;
  assign \new_[39396]_  = ~A199 & A167;
  assign \new_[39397]_  = A168 & \new_[39396]_ ;
  assign \new_[39400]_  = ~A202 & ~A200;
  assign \new_[39403]_  = A233 & A232;
  assign \new_[39404]_  = \new_[39403]_  & \new_[39400]_ ;
  assign \new_[39405]_  = \new_[39404]_  & \new_[39397]_ ;
  assign \new_[39408]_  = ~A235 & ~A234;
  assign \new_[39411]_  = ~A268 & ~A267;
  assign \new_[39412]_  = \new_[39411]_  & \new_[39408]_ ;
  assign \new_[39415]_  = ~A300 & ~A269;
  assign \new_[39418]_  = ~A302 & ~A301;
  assign \new_[39419]_  = \new_[39418]_  & \new_[39415]_ ;
  assign \new_[39420]_  = \new_[39419]_  & \new_[39412]_ ;
  assign \new_[39424]_  = ~A199 & A167;
  assign \new_[39425]_  = A168 & \new_[39424]_ ;
  assign \new_[39428]_  = ~A202 & ~A200;
  assign \new_[39431]_  = A233 & A232;
  assign \new_[39432]_  = \new_[39431]_  & \new_[39428]_ ;
  assign \new_[39433]_  = \new_[39432]_  & \new_[39425]_ ;
  assign \new_[39436]_  = ~A235 & ~A234;
  assign \new_[39439]_  = ~A268 & ~A267;
  assign \new_[39440]_  = \new_[39439]_  & \new_[39436]_ ;
  assign \new_[39443]_  = ~A298 & ~A269;
  assign \new_[39446]_  = ~A301 & ~A299;
  assign \new_[39447]_  = \new_[39446]_  & \new_[39443]_ ;
  assign \new_[39448]_  = \new_[39447]_  & \new_[39440]_ ;
  assign \new_[39452]_  = ~A199 & A167;
  assign \new_[39453]_  = A168 & \new_[39452]_ ;
  assign \new_[39456]_  = ~A202 & ~A200;
  assign \new_[39459]_  = A233 & A232;
  assign \new_[39460]_  = \new_[39459]_  & \new_[39456]_ ;
  assign \new_[39461]_  = \new_[39460]_  & \new_[39453]_ ;
  assign \new_[39464]_  = ~A235 & ~A234;
  assign \new_[39467]_  = ~A266 & ~A265;
  assign \new_[39468]_  = \new_[39467]_  & \new_[39464]_ ;
  assign \new_[39471]_  = ~A300 & ~A268;
  assign \new_[39474]_  = ~A302 & ~A301;
  assign \new_[39475]_  = \new_[39474]_  & \new_[39471]_ ;
  assign \new_[39476]_  = \new_[39475]_  & \new_[39468]_ ;
  assign \new_[39480]_  = ~A199 & A167;
  assign \new_[39481]_  = A168 & \new_[39480]_ ;
  assign \new_[39484]_  = ~A202 & ~A200;
  assign \new_[39487]_  = A233 & A232;
  assign \new_[39488]_  = \new_[39487]_  & \new_[39484]_ ;
  assign \new_[39489]_  = \new_[39488]_  & \new_[39481]_ ;
  assign \new_[39492]_  = ~A235 & ~A234;
  assign \new_[39495]_  = ~A266 & ~A265;
  assign \new_[39496]_  = \new_[39495]_  & \new_[39492]_ ;
  assign \new_[39499]_  = ~A298 & ~A268;
  assign \new_[39502]_  = ~A301 & ~A299;
  assign \new_[39503]_  = \new_[39502]_  & \new_[39499]_ ;
  assign \new_[39504]_  = \new_[39503]_  & \new_[39496]_ ;
  assign \new_[39508]_  = ~A199 & A167;
  assign \new_[39509]_  = A168 & \new_[39508]_ ;
  assign \new_[39512]_  = ~A202 & ~A200;
  assign \new_[39515]_  = ~A233 & ~A232;
  assign \new_[39516]_  = \new_[39515]_  & \new_[39512]_ ;
  assign \new_[39517]_  = \new_[39516]_  & \new_[39509]_ ;
  assign \new_[39520]_  = ~A267 & ~A235;
  assign \new_[39523]_  = ~A269 & ~A268;
  assign \new_[39524]_  = \new_[39523]_  & \new_[39520]_ ;
  assign \new_[39527]_  = A299 & A298;
  assign \new_[39530]_  = ~A301 & ~A300;
  assign \new_[39531]_  = \new_[39530]_  & \new_[39527]_ ;
  assign \new_[39532]_  = \new_[39531]_  & \new_[39524]_ ;
  assign \new_[39536]_  = ~A199 & A167;
  assign \new_[39537]_  = A168 & \new_[39536]_ ;
  assign \new_[39540]_  = ~A202 & ~A200;
  assign \new_[39543]_  = ~A233 & ~A232;
  assign \new_[39544]_  = \new_[39543]_  & \new_[39540]_ ;
  assign \new_[39545]_  = \new_[39544]_  & \new_[39537]_ ;
  assign \new_[39548]_  = A265 & ~A235;
  assign \new_[39551]_  = ~A267 & A266;
  assign \new_[39552]_  = \new_[39551]_  & \new_[39548]_ ;
  assign \new_[39555]_  = ~A300 & ~A268;
  assign \new_[39558]_  = ~A302 & ~A301;
  assign \new_[39559]_  = \new_[39558]_  & \new_[39555]_ ;
  assign \new_[39560]_  = \new_[39559]_  & \new_[39552]_ ;
  assign \new_[39564]_  = ~A199 & A167;
  assign \new_[39565]_  = A168 & \new_[39564]_ ;
  assign \new_[39568]_  = ~A202 & ~A200;
  assign \new_[39571]_  = ~A233 & ~A232;
  assign \new_[39572]_  = \new_[39571]_  & \new_[39568]_ ;
  assign \new_[39573]_  = \new_[39572]_  & \new_[39565]_ ;
  assign \new_[39576]_  = A265 & ~A235;
  assign \new_[39579]_  = ~A267 & A266;
  assign \new_[39580]_  = \new_[39579]_  & \new_[39576]_ ;
  assign \new_[39583]_  = ~A298 & ~A268;
  assign \new_[39586]_  = ~A301 & ~A299;
  assign \new_[39587]_  = \new_[39586]_  & \new_[39583]_ ;
  assign \new_[39588]_  = \new_[39587]_  & \new_[39580]_ ;
  assign \new_[39592]_  = ~A199 & A167;
  assign \new_[39593]_  = A168 & \new_[39592]_ ;
  assign \new_[39596]_  = ~A202 & ~A200;
  assign \new_[39599]_  = ~A233 & ~A232;
  assign \new_[39600]_  = \new_[39599]_  & \new_[39596]_ ;
  assign \new_[39601]_  = \new_[39600]_  & \new_[39593]_ ;
  assign \new_[39604]_  = ~A265 & ~A235;
  assign \new_[39607]_  = ~A268 & ~A266;
  assign \new_[39608]_  = \new_[39607]_  & \new_[39604]_ ;
  assign \new_[39611]_  = A299 & A298;
  assign \new_[39614]_  = ~A301 & ~A300;
  assign \new_[39615]_  = \new_[39614]_  & \new_[39611]_ ;
  assign \new_[39616]_  = \new_[39615]_  & \new_[39608]_ ;
  assign \new_[39620]_  = ~A166 & A167;
  assign \new_[39621]_  = A170 & \new_[39620]_ ;
  assign \new_[39624]_  = ~A202 & ~A201;
  assign \new_[39627]_  = ~A234 & ~A203;
  assign \new_[39628]_  = \new_[39627]_  & \new_[39624]_ ;
  assign \new_[39629]_  = \new_[39628]_  & \new_[39621]_ ;
  assign \new_[39632]_  = ~A236 & ~A235;
  assign \new_[39635]_  = ~A268 & ~A267;
  assign \new_[39636]_  = \new_[39635]_  & \new_[39632]_ ;
  assign \new_[39639]_  = ~A300 & ~A269;
  assign \new_[39642]_  = ~A302 & ~A301;
  assign \new_[39643]_  = \new_[39642]_  & \new_[39639]_ ;
  assign \new_[39644]_  = \new_[39643]_  & \new_[39636]_ ;
  assign \new_[39648]_  = ~A166 & A167;
  assign \new_[39649]_  = A170 & \new_[39648]_ ;
  assign \new_[39652]_  = ~A202 & ~A201;
  assign \new_[39655]_  = ~A234 & ~A203;
  assign \new_[39656]_  = \new_[39655]_  & \new_[39652]_ ;
  assign \new_[39657]_  = \new_[39656]_  & \new_[39649]_ ;
  assign \new_[39660]_  = ~A236 & ~A235;
  assign \new_[39663]_  = ~A268 & ~A267;
  assign \new_[39664]_  = \new_[39663]_  & \new_[39660]_ ;
  assign \new_[39667]_  = ~A298 & ~A269;
  assign \new_[39670]_  = ~A301 & ~A299;
  assign \new_[39671]_  = \new_[39670]_  & \new_[39667]_ ;
  assign \new_[39672]_  = \new_[39671]_  & \new_[39664]_ ;
  assign \new_[39676]_  = ~A166 & A167;
  assign \new_[39677]_  = A170 & \new_[39676]_ ;
  assign \new_[39680]_  = ~A202 & ~A201;
  assign \new_[39683]_  = ~A234 & ~A203;
  assign \new_[39684]_  = \new_[39683]_  & \new_[39680]_ ;
  assign \new_[39685]_  = \new_[39684]_  & \new_[39677]_ ;
  assign \new_[39688]_  = ~A236 & ~A235;
  assign \new_[39691]_  = ~A266 & ~A265;
  assign \new_[39692]_  = \new_[39691]_  & \new_[39688]_ ;
  assign \new_[39695]_  = ~A300 & ~A268;
  assign \new_[39698]_  = ~A302 & ~A301;
  assign \new_[39699]_  = \new_[39698]_  & \new_[39695]_ ;
  assign \new_[39700]_  = \new_[39699]_  & \new_[39692]_ ;
  assign \new_[39704]_  = ~A166 & A167;
  assign \new_[39705]_  = A170 & \new_[39704]_ ;
  assign \new_[39708]_  = ~A202 & ~A201;
  assign \new_[39711]_  = ~A234 & ~A203;
  assign \new_[39712]_  = \new_[39711]_  & \new_[39708]_ ;
  assign \new_[39713]_  = \new_[39712]_  & \new_[39705]_ ;
  assign \new_[39716]_  = ~A236 & ~A235;
  assign \new_[39719]_  = ~A266 & ~A265;
  assign \new_[39720]_  = \new_[39719]_  & \new_[39716]_ ;
  assign \new_[39723]_  = ~A298 & ~A268;
  assign \new_[39726]_  = ~A301 & ~A299;
  assign \new_[39727]_  = \new_[39726]_  & \new_[39723]_ ;
  assign \new_[39728]_  = \new_[39727]_  & \new_[39720]_ ;
  assign \new_[39732]_  = ~A166 & A167;
  assign \new_[39733]_  = A170 & \new_[39732]_ ;
  assign \new_[39736]_  = ~A202 & ~A201;
  assign \new_[39739]_  = ~A232 & ~A203;
  assign \new_[39740]_  = \new_[39739]_  & \new_[39736]_ ;
  assign \new_[39741]_  = \new_[39740]_  & \new_[39733]_ ;
  assign \new_[39744]_  = ~A235 & ~A233;
  assign \new_[39747]_  = ~A268 & ~A267;
  assign \new_[39748]_  = \new_[39747]_  & \new_[39744]_ ;
  assign \new_[39751]_  = ~A300 & ~A269;
  assign \new_[39754]_  = ~A302 & ~A301;
  assign \new_[39755]_  = \new_[39754]_  & \new_[39751]_ ;
  assign \new_[39756]_  = \new_[39755]_  & \new_[39748]_ ;
  assign \new_[39760]_  = ~A166 & A167;
  assign \new_[39761]_  = A170 & \new_[39760]_ ;
  assign \new_[39764]_  = ~A202 & ~A201;
  assign \new_[39767]_  = ~A232 & ~A203;
  assign \new_[39768]_  = \new_[39767]_  & \new_[39764]_ ;
  assign \new_[39769]_  = \new_[39768]_  & \new_[39761]_ ;
  assign \new_[39772]_  = ~A235 & ~A233;
  assign \new_[39775]_  = ~A268 & ~A267;
  assign \new_[39776]_  = \new_[39775]_  & \new_[39772]_ ;
  assign \new_[39779]_  = ~A298 & ~A269;
  assign \new_[39782]_  = ~A301 & ~A299;
  assign \new_[39783]_  = \new_[39782]_  & \new_[39779]_ ;
  assign \new_[39784]_  = \new_[39783]_  & \new_[39776]_ ;
  assign \new_[39788]_  = ~A166 & A167;
  assign \new_[39789]_  = A170 & \new_[39788]_ ;
  assign \new_[39792]_  = ~A202 & ~A201;
  assign \new_[39795]_  = ~A232 & ~A203;
  assign \new_[39796]_  = \new_[39795]_  & \new_[39792]_ ;
  assign \new_[39797]_  = \new_[39796]_  & \new_[39789]_ ;
  assign \new_[39800]_  = ~A235 & ~A233;
  assign \new_[39803]_  = ~A266 & ~A265;
  assign \new_[39804]_  = \new_[39803]_  & \new_[39800]_ ;
  assign \new_[39807]_  = ~A300 & ~A268;
  assign \new_[39810]_  = ~A302 & ~A301;
  assign \new_[39811]_  = \new_[39810]_  & \new_[39807]_ ;
  assign \new_[39812]_  = \new_[39811]_  & \new_[39804]_ ;
  assign \new_[39816]_  = ~A166 & A167;
  assign \new_[39817]_  = A170 & \new_[39816]_ ;
  assign \new_[39820]_  = ~A202 & ~A201;
  assign \new_[39823]_  = ~A232 & ~A203;
  assign \new_[39824]_  = \new_[39823]_  & \new_[39820]_ ;
  assign \new_[39825]_  = \new_[39824]_  & \new_[39817]_ ;
  assign \new_[39828]_  = ~A235 & ~A233;
  assign \new_[39831]_  = ~A266 & ~A265;
  assign \new_[39832]_  = \new_[39831]_  & \new_[39828]_ ;
  assign \new_[39835]_  = ~A298 & ~A268;
  assign \new_[39838]_  = ~A301 & ~A299;
  assign \new_[39839]_  = \new_[39838]_  & \new_[39835]_ ;
  assign \new_[39840]_  = \new_[39839]_  & \new_[39832]_ ;
  assign \new_[39844]_  = ~A166 & A167;
  assign \new_[39845]_  = A170 & \new_[39844]_ ;
  assign \new_[39848]_  = ~A200 & ~A199;
  assign \new_[39851]_  = ~A234 & ~A202;
  assign \new_[39852]_  = \new_[39851]_  & \new_[39848]_ ;
  assign \new_[39853]_  = \new_[39852]_  & \new_[39845]_ ;
  assign \new_[39856]_  = ~A236 & ~A235;
  assign \new_[39859]_  = ~A268 & ~A267;
  assign \new_[39860]_  = \new_[39859]_  & \new_[39856]_ ;
  assign \new_[39863]_  = ~A300 & ~A269;
  assign \new_[39866]_  = ~A302 & ~A301;
  assign \new_[39867]_  = \new_[39866]_  & \new_[39863]_ ;
  assign \new_[39868]_  = \new_[39867]_  & \new_[39860]_ ;
  assign \new_[39872]_  = ~A166 & A167;
  assign \new_[39873]_  = A170 & \new_[39872]_ ;
  assign \new_[39876]_  = ~A200 & ~A199;
  assign \new_[39879]_  = ~A234 & ~A202;
  assign \new_[39880]_  = \new_[39879]_  & \new_[39876]_ ;
  assign \new_[39881]_  = \new_[39880]_  & \new_[39873]_ ;
  assign \new_[39884]_  = ~A236 & ~A235;
  assign \new_[39887]_  = ~A268 & ~A267;
  assign \new_[39888]_  = \new_[39887]_  & \new_[39884]_ ;
  assign \new_[39891]_  = ~A298 & ~A269;
  assign \new_[39894]_  = ~A301 & ~A299;
  assign \new_[39895]_  = \new_[39894]_  & \new_[39891]_ ;
  assign \new_[39896]_  = \new_[39895]_  & \new_[39888]_ ;
  assign \new_[39900]_  = ~A166 & A167;
  assign \new_[39901]_  = A170 & \new_[39900]_ ;
  assign \new_[39904]_  = ~A200 & ~A199;
  assign \new_[39907]_  = ~A234 & ~A202;
  assign \new_[39908]_  = \new_[39907]_  & \new_[39904]_ ;
  assign \new_[39909]_  = \new_[39908]_  & \new_[39901]_ ;
  assign \new_[39912]_  = ~A236 & ~A235;
  assign \new_[39915]_  = ~A266 & ~A265;
  assign \new_[39916]_  = \new_[39915]_  & \new_[39912]_ ;
  assign \new_[39919]_  = ~A300 & ~A268;
  assign \new_[39922]_  = ~A302 & ~A301;
  assign \new_[39923]_  = \new_[39922]_  & \new_[39919]_ ;
  assign \new_[39924]_  = \new_[39923]_  & \new_[39916]_ ;
  assign \new_[39928]_  = ~A166 & A167;
  assign \new_[39929]_  = A170 & \new_[39928]_ ;
  assign \new_[39932]_  = ~A200 & ~A199;
  assign \new_[39935]_  = ~A234 & ~A202;
  assign \new_[39936]_  = \new_[39935]_  & \new_[39932]_ ;
  assign \new_[39937]_  = \new_[39936]_  & \new_[39929]_ ;
  assign \new_[39940]_  = ~A236 & ~A235;
  assign \new_[39943]_  = ~A266 & ~A265;
  assign \new_[39944]_  = \new_[39943]_  & \new_[39940]_ ;
  assign \new_[39947]_  = ~A298 & ~A268;
  assign \new_[39950]_  = ~A301 & ~A299;
  assign \new_[39951]_  = \new_[39950]_  & \new_[39947]_ ;
  assign \new_[39952]_  = \new_[39951]_  & \new_[39944]_ ;
  assign \new_[39956]_  = ~A166 & A167;
  assign \new_[39957]_  = A170 & \new_[39956]_ ;
  assign \new_[39960]_  = ~A200 & ~A199;
  assign \new_[39963]_  = ~A232 & ~A202;
  assign \new_[39964]_  = \new_[39963]_  & \new_[39960]_ ;
  assign \new_[39965]_  = \new_[39964]_  & \new_[39957]_ ;
  assign \new_[39968]_  = ~A235 & ~A233;
  assign \new_[39971]_  = ~A268 & ~A267;
  assign \new_[39972]_  = \new_[39971]_  & \new_[39968]_ ;
  assign \new_[39975]_  = ~A300 & ~A269;
  assign \new_[39978]_  = ~A302 & ~A301;
  assign \new_[39979]_  = \new_[39978]_  & \new_[39975]_ ;
  assign \new_[39980]_  = \new_[39979]_  & \new_[39972]_ ;
  assign \new_[39984]_  = ~A166 & A167;
  assign \new_[39985]_  = A170 & \new_[39984]_ ;
  assign \new_[39988]_  = ~A200 & ~A199;
  assign \new_[39991]_  = ~A232 & ~A202;
  assign \new_[39992]_  = \new_[39991]_  & \new_[39988]_ ;
  assign \new_[39993]_  = \new_[39992]_  & \new_[39985]_ ;
  assign \new_[39996]_  = ~A235 & ~A233;
  assign \new_[39999]_  = ~A268 & ~A267;
  assign \new_[40000]_  = \new_[39999]_  & \new_[39996]_ ;
  assign \new_[40003]_  = ~A298 & ~A269;
  assign \new_[40006]_  = ~A301 & ~A299;
  assign \new_[40007]_  = \new_[40006]_  & \new_[40003]_ ;
  assign \new_[40008]_  = \new_[40007]_  & \new_[40000]_ ;
  assign \new_[40012]_  = ~A166 & A167;
  assign \new_[40013]_  = A170 & \new_[40012]_ ;
  assign \new_[40016]_  = ~A200 & ~A199;
  assign \new_[40019]_  = ~A232 & ~A202;
  assign \new_[40020]_  = \new_[40019]_  & \new_[40016]_ ;
  assign \new_[40021]_  = \new_[40020]_  & \new_[40013]_ ;
  assign \new_[40024]_  = ~A235 & ~A233;
  assign \new_[40027]_  = ~A266 & ~A265;
  assign \new_[40028]_  = \new_[40027]_  & \new_[40024]_ ;
  assign \new_[40031]_  = ~A300 & ~A268;
  assign \new_[40034]_  = ~A302 & ~A301;
  assign \new_[40035]_  = \new_[40034]_  & \new_[40031]_ ;
  assign \new_[40036]_  = \new_[40035]_  & \new_[40028]_ ;
  assign \new_[40040]_  = ~A166 & A167;
  assign \new_[40041]_  = A170 & \new_[40040]_ ;
  assign \new_[40044]_  = ~A200 & ~A199;
  assign \new_[40047]_  = ~A232 & ~A202;
  assign \new_[40048]_  = \new_[40047]_  & \new_[40044]_ ;
  assign \new_[40049]_  = \new_[40048]_  & \new_[40041]_ ;
  assign \new_[40052]_  = ~A235 & ~A233;
  assign \new_[40055]_  = ~A266 & ~A265;
  assign \new_[40056]_  = \new_[40055]_  & \new_[40052]_ ;
  assign \new_[40059]_  = ~A298 & ~A268;
  assign \new_[40062]_  = ~A301 & ~A299;
  assign \new_[40063]_  = \new_[40062]_  & \new_[40059]_ ;
  assign \new_[40064]_  = \new_[40063]_  & \new_[40056]_ ;
  assign \new_[40068]_  = A166 & ~A167;
  assign \new_[40069]_  = A170 & \new_[40068]_ ;
  assign \new_[40072]_  = ~A202 & ~A201;
  assign \new_[40075]_  = ~A234 & ~A203;
  assign \new_[40076]_  = \new_[40075]_  & \new_[40072]_ ;
  assign \new_[40077]_  = \new_[40076]_  & \new_[40069]_ ;
  assign \new_[40080]_  = ~A236 & ~A235;
  assign \new_[40083]_  = ~A268 & ~A267;
  assign \new_[40084]_  = \new_[40083]_  & \new_[40080]_ ;
  assign \new_[40087]_  = ~A300 & ~A269;
  assign \new_[40090]_  = ~A302 & ~A301;
  assign \new_[40091]_  = \new_[40090]_  & \new_[40087]_ ;
  assign \new_[40092]_  = \new_[40091]_  & \new_[40084]_ ;
  assign \new_[40096]_  = A166 & ~A167;
  assign \new_[40097]_  = A170 & \new_[40096]_ ;
  assign \new_[40100]_  = ~A202 & ~A201;
  assign \new_[40103]_  = ~A234 & ~A203;
  assign \new_[40104]_  = \new_[40103]_  & \new_[40100]_ ;
  assign \new_[40105]_  = \new_[40104]_  & \new_[40097]_ ;
  assign \new_[40108]_  = ~A236 & ~A235;
  assign \new_[40111]_  = ~A268 & ~A267;
  assign \new_[40112]_  = \new_[40111]_  & \new_[40108]_ ;
  assign \new_[40115]_  = ~A298 & ~A269;
  assign \new_[40118]_  = ~A301 & ~A299;
  assign \new_[40119]_  = \new_[40118]_  & \new_[40115]_ ;
  assign \new_[40120]_  = \new_[40119]_  & \new_[40112]_ ;
  assign \new_[40124]_  = A166 & ~A167;
  assign \new_[40125]_  = A170 & \new_[40124]_ ;
  assign \new_[40128]_  = ~A202 & ~A201;
  assign \new_[40131]_  = ~A234 & ~A203;
  assign \new_[40132]_  = \new_[40131]_  & \new_[40128]_ ;
  assign \new_[40133]_  = \new_[40132]_  & \new_[40125]_ ;
  assign \new_[40136]_  = ~A236 & ~A235;
  assign \new_[40139]_  = ~A266 & ~A265;
  assign \new_[40140]_  = \new_[40139]_  & \new_[40136]_ ;
  assign \new_[40143]_  = ~A300 & ~A268;
  assign \new_[40146]_  = ~A302 & ~A301;
  assign \new_[40147]_  = \new_[40146]_  & \new_[40143]_ ;
  assign \new_[40148]_  = \new_[40147]_  & \new_[40140]_ ;
  assign \new_[40152]_  = A166 & ~A167;
  assign \new_[40153]_  = A170 & \new_[40152]_ ;
  assign \new_[40156]_  = ~A202 & ~A201;
  assign \new_[40159]_  = ~A234 & ~A203;
  assign \new_[40160]_  = \new_[40159]_  & \new_[40156]_ ;
  assign \new_[40161]_  = \new_[40160]_  & \new_[40153]_ ;
  assign \new_[40164]_  = ~A236 & ~A235;
  assign \new_[40167]_  = ~A266 & ~A265;
  assign \new_[40168]_  = \new_[40167]_  & \new_[40164]_ ;
  assign \new_[40171]_  = ~A298 & ~A268;
  assign \new_[40174]_  = ~A301 & ~A299;
  assign \new_[40175]_  = \new_[40174]_  & \new_[40171]_ ;
  assign \new_[40176]_  = \new_[40175]_  & \new_[40168]_ ;
  assign \new_[40180]_  = A166 & ~A167;
  assign \new_[40181]_  = A170 & \new_[40180]_ ;
  assign \new_[40184]_  = ~A202 & ~A201;
  assign \new_[40187]_  = ~A232 & ~A203;
  assign \new_[40188]_  = \new_[40187]_  & \new_[40184]_ ;
  assign \new_[40189]_  = \new_[40188]_  & \new_[40181]_ ;
  assign \new_[40192]_  = ~A235 & ~A233;
  assign \new_[40195]_  = ~A268 & ~A267;
  assign \new_[40196]_  = \new_[40195]_  & \new_[40192]_ ;
  assign \new_[40199]_  = ~A300 & ~A269;
  assign \new_[40202]_  = ~A302 & ~A301;
  assign \new_[40203]_  = \new_[40202]_  & \new_[40199]_ ;
  assign \new_[40204]_  = \new_[40203]_  & \new_[40196]_ ;
  assign \new_[40208]_  = A166 & ~A167;
  assign \new_[40209]_  = A170 & \new_[40208]_ ;
  assign \new_[40212]_  = ~A202 & ~A201;
  assign \new_[40215]_  = ~A232 & ~A203;
  assign \new_[40216]_  = \new_[40215]_  & \new_[40212]_ ;
  assign \new_[40217]_  = \new_[40216]_  & \new_[40209]_ ;
  assign \new_[40220]_  = ~A235 & ~A233;
  assign \new_[40223]_  = ~A268 & ~A267;
  assign \new_[40224]_  = \new_[40223]_  & \new_[40220]_ ;
  assign \new_[40227]_  = ~A298 & ~A269;
  assign \new_[40230]_  = ~A301 & ~A299;
  assign \new_[40231]_  = \new_[40230]_  & \new_[40227]_ ;
  assign \new_[40232]_  = \new_[40231]_  & \new_[40224]_ ;
  assign \new_[40236]_  = A166 & ~A167;
  assign \new_[40237]_  = A170 & \new_[40236]_ ;
  assign \new_[40240]_  = ~A202 & ~A201;
  assign \new_[40243]_  = ~A232 & ~A203;
  assign \new_[40244]_  = \new_[40243]_  & \new_[40240]_ ;
  assign \new_[40245]_  = \new_[40244]_  & \new_[40237]_ ;
  assign \new_[40248]_  = ~A235 & ~A233;
  assign \new_[40251]_  = ~A266 & ~A265;
  assign \new_[40252]_  = \new_[40251]_  & \new_[40248]_ ;
  assign \new_[40255]_  = ~A300 & ~A268;
  assign \new_[40258]_  = ~A302 & ~A301;
  assign \new_[40259]_  = \new_[40258]_  & \new_[40255]_ ;
  assign \new_[40260]_  = \new_[40259]_  & \new_[40252]_ ;
  assign \new_[40264]_  = A166 & ~A167;
  assign \new_[40265]_  = A170 & \new_[40264]_ ;
  assign \new_[40268]_  = ~A202 & ~A201;
  assign \new_[40271]_  = ~A232 & ~A203;
  assign \new_[40272]_  = \new_[40271]_  & \new_[40268]_ ;
  assign \new_[40273]_  = \new_[40272]_  & \new_[40265]_ ;
  assign \new_[40276]_  = ~A235 & ~A233;
  assign \new_[40279]_  = ~A266 & ~A265;
  assign \new_[40280]_  = \new_[40279]_  & \new_[40276]_ ;
  assign \new_[40283]_  = ~A298 & ~A268;
  assign \new_[40286]_  = ~A301 & ~A299;
  assign \new_[40287]_  = \new_[40286]_  & \new_[40283]_ ;
  assign \new_[40288]_  = \new_[40287]_  & \new_[40280]_ ;
  assign \new_[40292]_  = A166 & ~A167;
  assign \new_[40293]_  = A170 & \new_[40292]_ ;
  assign \new_[40296]_  = ~A200 & ~A199;
  assign \new_[40299]_  = ~A234 & ~A202;
  assign \new_[40300]_  = \new_[40299]_  & \new_[40296]_ ;
  assign \new_[40301]_  = \new_[40300]_  & \new_[40293]_ ;
  assign \new_[40304]_  = ~A236 & ~A235;
  assign \new_[40307]_  = ~A268 & ~A267;
  assign \new_[40308]_  = \new_[40307]_  & \new_[40304]_ ;
  assign \new_[40311]_  = ~A300 & ~A269;
  assign \new_[40314]_  = ~A302 & ~A301;
  assign \new_[40315]_  = \new_[40314]_  & \new_[40311]_ ;
  assign \new_[40316]_  = \new_[40315]_  & \new_[40308]_ ;
  assign \new_[40320]_  = A166 & ~A167;
  assign \new_[40321]_  = A170 & \new_[40320]_ ;
  assign \new_[40324]_  = ~A200 & ~A199;
  assign \new_[40327]_  = ~A234 & ~A202;
  assign \new_[40328]_  = \new_[40327]_  & \new_[40324]_ ;
  assign \new_[40329]_  = \new_[40328]_  & \new_[40321]_ ;
  assign \new_[40332]_  = ~A236 & ~A235;
  assign \new_[40335]_  = ~A268 & ~A267;
  assign \new_[40336]_  = \new_[40335]_  & \new_[40332]_ ;
  assign \new_[40339]_  = ~A298 & ~A269;
  assign \new_[40342]_  = ~A301 & ~A299;
  assign \new_[40343]_  = \new_[40342]_  & \new_[40339]_ ;
  assign \new_[40344]_  = \new_[40343]_  & \new_[40336]_ ;
  assign \new_[40348]_  = A166 & ~A167;
  assign \new_[40349]_  = A170 & \new_[40348]_ ;
  assign \new_[40352]_  = ~A200 & ~A199;
  assign \new_[40355]_  = ~A234 & ~A202;
  assign \new_[40356]_  = \new_[40355]_  & \new_[40352]_ ;
  assign \new_[40357]_  = \new_[40356]_  & \new_[40349]_ ;
  assign \new_[40360]_  = ~A236 & ~A235;
  assign \new_[40363]_  = ~A266 & ~A265;
  assign \new_[40364]_  = \new_[40363]_  & \new_[40360]_ ;
  assign \new_[40367]_  = ~A300 & ~A268;
  assign \new_[40370]_  = ~A302 & ~A301;
  assign \new_[40371]_  = \new_[40370]_  & \new_[40367]_ ;
  assign \new_[40372]_  = \new_[40371]_  & \new_[40364]_ ;
  assign \new_[40376]_  = A166 & ~A167;
  assign \new_[40377]_  = A170 & \new_[40376]_ ;
  assign \new_[40380]_  = ~A200 & ~A199;
  assign \new_[40383]_  = ~A234 & ~A202;
  assign \new_[40384]_  = \new_[40383]_  & \new_[40380]_ ;
  assign \new_[40385]_  = \new_[40384]_  & \new_[40377]_ ;
  assign \new_[40388]_  = ~A236 & ~A235;
  assign \new_[40391]_  = ~A266 & ~A265;
  assign \new_[40392]_  = \new_[40391]_  & \new_[40388]_ ;
  assign \new_[40395]_  = ~A298 & ~A268;
  assign \new_[40398]_  = ~A301 & ~A299;
  assign \new_[40399]_  = \new_[40398]_  & \new_[40395]_ ;
  assign \new_[40400]_  = \new_[40399]_  & \new_[40392]_ ;
  assign \new_[40404]_  = A166 & ~A167;
  assign \new_[40405]_  = A170 & \new_[40404]_ ;
  assign \new_[40408]_  = ~A200 & ~A199;
  assign \new_[40411]_  = ~A232 & ~A202;
  assign \new_[40412]_  = \new_[40411]_  & \new_[40408]_ ;
  assign \new_[40413]_  = \new_[40412]_  & \new_[40405]_ ;
  assign \new_[40416]_  = ~A235 & ~A233;
  assign \new_[40419]_  = ~A268 & ~A267;
  assign \new_[40420]_  = \new_[40419]_  & \new_[40416]_ ;
  assign \new_[40423]_  = ~A300 & ~A269;
  assign \new_[40426]_  = ~A302 & ~A301;
  assign \new_[40427]_  = \new_[40426]_  & \new_[40423]_ ;
  assign \new_[40428]_  = \new_[40427]_  & \new_[40420]_ ;
  assign \new_[40432]_  = A166 & ~A167;
  assign \new_[40433]_  = A170 & \new_[40432]_ ;
  assign \new_[40436]_  = ~A200 & ~A199;
  assign \new_[40439]_  = ~A232 & ~A202;
  assign \new_[40440]_  = \new_[40439]_  & \new_[40436]_ ;
  assign \new_[40441]_  = \new_[40440]_  & \new_[40433]_ ;
  assign \new_[40444]_  = ~A235 & ~A233;
  assign \new_[40447]_  = ~A268 & ~A267;
  assign \new_[40448]_  = \new_[40447]_  & \new_[40444]_ ;
  assign \new_[40451]_  = ~A298 & ~A269;
  assign \new_[40454]_  = ~A301 & ~A299;
  assign \new_[40455]_  = \new_[40454]_  & \new_[40451]_ ;
  assign \new_[40456]_  = \new_[40455]_  & \new_[40448]_ ;
  assign \new_[40460]_  = A166 & ~A167;
  assign \new_[40461]_  = A170 & \new_[40460]_ ;
  assign \new_[40464]_  = ~A200 & ~A199;
  assign \new_[40467]_  = ~A232 & ~A202;
  assign \new_[40468]_  = \new_[40467]_  & \new_[40464]_ ;
  assign \new_[40469]_  = \new_[40468]_  & \new_[40461]_ ;
  assign \new_[40472]_  = ~A235 & ~A233;
  assign \new_[40475]_  = ~A266 & ~A265;
  assign \new_[40476]_  = \new_[40475]_  & \new_[40472]_ ;
  assign \new_[40479]_  = ~A300 & ~A268;
  assign \new_[40482]_  = ~A302 & ~A301;
  assign \new_[40483]_  = \new_[40482]_  & \new_[40479]_ ;
  assign \new_[40484]_  = \new_[40483]_  & \new_[40476]_ ;
  assign \new_[40488]_  = A166 & ~A167;
  assign \new_[40489]_  = A170 & \new_[40488]_ ;
  assign \new_[40492]_  = ~A200 & ~A199;
  assign \new_[40495]_  = ~A232 & ~A202;
  assign \new_[40496]_  = \new_[40495]_  & \new_[40492]_ ;
  assign \new_[40497]_  = \new_[40496]_  & \new_[40489]_ ;
  assign \new_[40500]_  = ~A235 & ~A233;
  assign \new_[40503]_  = ~A266 & ~A265;
  assign \new_[40504]_  = \new_[40503]_  & \new_[40500]_ ;
  assign \new_[40507]_  = ~A298 & ~A268;
  assign \new_[40510]_  = ~A301 & ~A299;
  assign \new_[40511]_  = \new_[40510]_  & \new_[40507]_ ;
  assign \new_[40512]_  = \new_[40511]_  & \new_[40504]_ ;
  assign \new_[40516]_  = ~A202 & ~A201;
  assign \new_[40517]_  = A169 & \new_[40516]_ ;
  assign \new_[40520]_  = ~A234 & ~A203;
  assign \new_[40523]_  = ~A236 & ~A235;
  assign \new_[40524]_  = \new_[40523]_  & \new_[40520]_ ;
  assign \new_[40525]_  = \new_[40524]_  & \new_[40517]_ ;
  assign \new_[40528]_  = A266 & A265;
  assign \new_[40531]_  = ~A268 & ~A267;
  assign \new_[40532]_  = \new_[40531]_  & \new_[40528]_ ;
  assign \new_[40535]_  = A299 & A298;
  assign \new_[40538]_  = ~A301 & ~A300;
  assign \new_[40539]_  = \new_[40538]_  & \new_[40535]_ ;
  assign \new_[40540]_  = \new_[40539]_  & \new_[40532]_ ;
  assign \new_[40544]_  = ~A202 & ~A201;
  assign \new_[40545]_  = A169 & \new_[40544]_ ;
  assign \new_[40548]_  = A232 & ~A203;
  assign \new_[40551]_  = ~A234 & A233;
  assign \new_[40552]_  = \new_[40551]_  & \new_[40548]_ ;
  assign \new_[40553]_  = \new_[40552]_  & \new_[40545]_ ;
  assign \new_[40556]_  = ~A267 & ~A235;
  assign \new_[40559]_  = ~A269 & ~A268;
  assign \new_[40560]_  = \new_[40559]_  & \new_[40556]_ ;
  assign \new_[40563]_  = A299 & A298;
  assign \new_[40566]_  = ~A301 & ~A300;
  assign \new_[40567]_  = \new_[40566]_  & \new_[40563]_ ;
  assign \new_[40568]_  = \new_[40567]_  & \new_[40560]_ ;
  assign \new_[40572]_  = ~A202 & ~A201;
  assign \new_[40573]_  = A169 & \new_[40572]_ ;
  assign \new_[40576]_  = A232 & ~A203;
  assign \new_[40579]_  = ~A234 & A233;
  assign \new_[40580]_  = \new_[40579]_  & \new_[40576]_ ;
  assign \new_[40581]_  = \new_[40580]_  & \new_[40573]_ ;
  assign \new_[40584]_  = A265 & ~A235;
  assign \new_[40587]_  = ~A267 & A266;
  assign \new_[40588]_  = \new_[40587]_  & \new_[40584]_ ;
  assign \new_[40591]_  = ~A300 & ~A268;
  assign \new_[40594]_  = ~A302 & ~A301;
  assign \new_[40595]_  = \new_[40594]_  & \new_[40591]_ ;
  assign \new_[40596]_  = \new_[40595]_  & \new_[40588]_ ;
  assign \new_[40600]_  = ~A202 & ~A201;
  assign \new_[40601]_  = A169 & \new_[40600]_ ;
  assign \new_[40604]_  = A232 & ~A203;
  assign \new_[40607]_  = ~A234 & A233;
  assign \new_[40608]_  = \new_[40607]_  & \new_[40604]_ ;
  assign \new_[40609]_  = \new_[40608]_  & \new_[40601]_ ;
  assign \new_[40612]_  = A265 & ~A235;
  assign \new_[40615]_  = ~A267 & A266;
  assign \new_[40616]_  = \new_[40615]_  & \new_[40612]_ ;
  assign \new_[40619]_  = ~A298 & ~A268;
  assign \new_[40622]_  = ~A301 & ~A299;
  assign \new_[40623]_  = \new_[40622]_  & \new_[40619]_ ;
  assign \new_[40624]_  = \new_[40623]_  & \new_[40616]_ ;
  assign \new_[40628]_  = ~A202 & ~A201;
  assign \new_[40629]_  = A169 & \new_[40628]_ ;
  assign \new_[40632]_  = A232 & ~A203;
  assign \new_[40635]_  = ~A234 & A233;
  assign \new_[40636]_  = \new_[40635]_  & \new_[40632]_ ;
  assign \new_[40637]_  = \new_[40636]_  & \new_[40629]_ ;
  assign \new_[40640]_  = ~A265 & ~A235;
  assign \new_[40643]_  = ~A268 & ~A266;
  assign \new_[40644]_  = \new_[40643]_  & \new_[40640]_ ;
  assign \new_[40647]_  = A299 & A298;
  assign \new_[40650]_  = ~A301 & ~A300;
  assign \new_[40651]_  = \new_[40650]_  & \new_[40647]_ ;
  assign \new_[40652]_  = \new_[40651]_  & \new_[40644]_ ;
  assign \new_[40656]_  = ~A202 & ~A201;
  assign \new_[40657]_  = A169 & \new_[40656]_ ;
  assign \new_[40660]_  = ~A232 & ~A203;
  assign \new_[40663]_  = ~A235 & ~A233;
  assign \new_[40664]_  = \new_[40663]_  & \new_[40660]_ ;
  assign \new_[40665]_  = \new_[40664]_  & \new_[40657]_ ;
  assign \new_[40668]_  = A266 & A265;
  assign \new_[40671]_  = ~A268 & ~A267;
  assign \new_[40672]_  = \new_[40671]_  & \new_[40668]_ ;
  assign \new_[40675]_  = A299 & A298;
  assign \new_[40678]_  = ~A301 & ~A300;
  assign \new_[40679]_  = \new_[40678]_  & \new_[40675]_ ;
  assign \new_[40680]_  = \new_[40679]_  & \new_[40672]_ ;
  assign \new_[40684]_  = A200 & A199;
  assign \new_[40685]_  = A169 & \new_[40684]_ ;
  assign \new_[40688]_  = ~A202 & ~A201;
  assign \new_[40691]_  = ~A235 & ~A234;
  assign \new_[40692]_  = \new_[40691]_  & \new_[40688]_ ;
  assign \new_[40693]_  = \new_[40692]_  & \new_[40685]_ ;
  assign \new_[40696]_  = ~A267 & ~A236;
  assign \new_[40699]_  = ~A269 & ~A268;
  assign \new_[40700]_  = \new_[40699]_  & \new_[40696]_ ;
  assign \new_[40703]_  = A299 & A298;
  assign \new_[40706]_  = ~A301 & ~A300;
  assign \new_[40707]_  = \new_[40706]_  & \new_[40703]_ ;
  assign \new_[40708]_  = \new_[40707]_  & \new_[40700]_ ;
  assign \new_[40712]_  = A200 & A199;
  assign \new_[40713]_  = A169 & \new_[40712]_ ;
  assign \new_[40716]_  = ~A202 & ~A201;
  assign \new_[40719]_  = ~A235 & ~A234;
  assign \new_[40720]_  = \new_[40719]_  & \new_[40716]_ ;
  assign \new_[40721]_  = \new_[40720]_  & \new_[40713]_ ;
  assign \new_[40724]_  = A265 & ~A236;
  assign \new_[40727]_  = ~A267 & A266;
  assign \new_[40728]_  = \new_[40727]_  & \new_[40724]_ ;
  assign \new_[40731]_  = ~A300 & ~A268;
  assign \new_[40734]_  = ~A302 & ~A301;
  assign \new_[40735]_  = \new_[40734]_  & \new_[40731]_ ;
  assign \new_[40736]_  = \new_[40735]_  & \new_[40728]_ ;
  assign \new_[40740]_  = A200 & A199;
  assign \new_[40741]_  = A169 & \new_[40740]_ ;
  assign \new_[40744]_  = ~A202 & ~A201;
  assign \new_[40747]_  = ~A235 & ~A234;
  assign \new_[40748]_  = \new_[40747]_  & \new_[40744]_ ;
  assign \new_[40749]_  = \new_[40748]_  & \new_[40741]_ ;
  assign \new_[40752]_  = A265 & ~A236;
  assign \new_[40755]_  = ~A267 & A266;
  assign \new_[40756]_  = \new_[40755]_  & \new_[40752]_ ;
  assign \new_[40759]_  = ~A298 & ~A268;
  assign \new_[40762]_  = ~A301 & ~A299;
  assign \new_[40763]_  = \new_[40762]_  & \new_[40759]_ ;
  assign \new_[40764]_  = \new_[40763]_  & \new_[40756]_ ;
  assign \new_[40768]_  = A200 & A199;
  assign \new_[40769]_  = A169 & \new_[40768]_ ;
  assign \new_[40772]_  = ~A202 & ~A201;
  assign \new_[40775]_  = ~A235 & ~A234;
  assign \new_[40776]_  = \new_[40775]_  & \new_[40772]_ ;
  assign \new_[40777]_  = \new_[40776]_  & \new_[40769]_ ;
  assign \new_[40780]_  = ~A265 & ~A236;
  assign \new_[40783]_  = ~A268 & ~A266;
  assign \new_[40784]_  = \new_[40783]_  & \new_[40780]_ ;
  assign \new_[40787]_  = A299 & A298;
  assign \new_[40790]_  = ~A301 & ~A300;
  assign \new_[40791]_  = \new_[40790]_  & \new_[40787]_ ;
  assign \new_[40792]_  = \new_[40791]_  & \new_[40784]_ ;
  assign \new_[40796]_  = A200 & A199;
  assign \new_[40797]_  = A169 & \new_[40796]_ ;
  assign \new_[40800]_  = ~A202 & ~A201;
  assign \new_[40803]_  = A233 & A232;
  assign \new_[40804]_  = \new_[40803]_  & \new_[40800]_ ;
  assign \new_[40805]_  = \new_[40804]_  & \new_[40797]_ ;
  assign \new_[40808]_  = ~A235 & ~A234;
  assign \new_[40811]_  = ~A268 & ~A267;
  assign \new_[40812]_  = \new_[40811]_  & \new_[40808]_ ;
  assign \new_[40815]_  = ~A300 & ~A269;
  assign \new_[40818]_  = ~A302 & ~A301;
  assign \new_[40819]_  = \new_[40818]_  & \new_[40815]_ ;
  assign \new_[40820]_  = \new_[40819]_  & \new_[40812]_ ;
  assign \new_[40824]_  = A200 & A199;
  assign \new_[40825]_  = A169 & \new_[40824]_ ;
  assign \new_[40828]_  = ~A202 & ~A201;
  assign \new_[40831]_  = A233 & A232;
  assign \new_[40832]_  = \new_[40831]_  & \new_[40828]_ ;
  assign \new_[40833]_  = \new_[40832]_  & \new_[40825]_ ;
  assign \new_[40836]_  = ~A235 & ~A234;
  assign \new_[40839]_  = ~A268 & ~A267;
  assign \new_[40840]_  = \new_[40839]_  & \new_[40836]_ ;
  assign \new_[40843]_  = ~A298 & ~A269;
  assign \new_[40846]_  = ~A301 & ~A299;
  assign \new_[40847]_  = \new_[40846]_  & \new_[40843]_ ;
  assign \new_[40848]_  = \new_[40847]_  & \new_[40840]_ ;
  assign \new_[40852]_  = A200 & A199;
  assign \new_[40853]_  = A169 & \new_[40852]_ ;
  assign \new_[40856]_  = ~A202 & ~A201;
  assign \new_[40859]_  = A233 & A232;
  assign \new_[40860]_  = \new_[40859]_  & \new_[40856]_ ;
  assign \new_[40861]_  = \new_[40860]_  & \new_[40853]_ ;
  assign \new_[40864]_  = ~A235 & ~A234;
  assign \new_[40867]_  = ~A266 & ~A265;
  assign \new_[40868]_  = \new_[40867]_  & \new_[40864]_ ;
  assign \new_[40871]_  = ~A300 & ~A268;
  assign \new_[40874]_  = ~A302 & ~A301;
  assign \new_[40875]_  = \new_[40874]_  & \new_[40871]_ ;
  assign \new_[40876]_  = \new_[40875]_  & \new_[40868]_ ;
  assign \new_[40880]_  = A200 & A199;
  assign \new_[40881]_  = A169 & \new_[40880]_ ;
  assign \new_[40884]_  = ~A202 & ~A201;
  assign \new_[40887]_  = A233 & A232;
  assign \new_[40888]_  = \new_[40887]_  & \new_[40884]_ ;
  assign \new_[40889]_  = \new_[40888]_  & \new_[40881]_ ;
  assign \new_[40892]_  = ~A235 & ~A234;
  assign \new_[40895]_  = ~A266 & ~A265;
  assign \new_[40896]_  = \new_[40895]_  & \new_[40892]_ ;
  assign \new_[40899]_  = ~A298 & ~A268;
  assign \new_[40902]_  = ~A301 & ~A299;
  assign \new_[40903]_  = \new_[40902]_  & \new_[40899]_ ;
  assign \new_[40904]_  = \new_[40903]_  & \new_[40896]_ ;
  assign \new_[40908]_  = A200 & A199;
  assign \new_[40909]_  = A169 & \new_[40908]_ ;
  assign \new_[40912]_  = ~A202 & ~A201;
  assign \new_[40915]_  = ~A233 & ~A232;
  assign \new_[40916]_  = \new_[40915]_  & \new_[40912]_ ;
  assign \new_[40917]_  = \new_[40916]_  & \new_[40909]_ ;
  assign \new_[40920]_  = ~A267 & ~A235;
  assign \new_[40923]_  = ~A269 & ~A268;
  assign \new_[40924]_  = \new_[40923]_  & \new_[40920]_ ;
  assign \new_[40927]_  = A299 & A298;
  assign \new_[40930]_  = ~A301 & ~A300;
  assign \new_[40931]_  = \new_[40930]_  & \new_[40927]_ ;
  assign \new_[40932]_  = \new_[40931]_  & \new_[40924]_ ;
  assign \new_[40936]_  = A200 & A199;
  assign \new_[40937]_  = A169 & \new_[40936]_ ;
  assign \new_[40940]_  = ~A202 & ~A201;
  assign \new_[40943]_  = ~A233 & ~A232;
  assign \new_[40944]_  = \new_[40943]_  & \new_[40940]_ ;
  assign \new_[40945]_  = \new_[40944]_  & \new_[40937]_ ;
  assign \new_[40948]_  = A265 & ~A235;
  assign \new_[40951]_  = ~A267 & A266;
  assign \new_[40952]_  = \new_[40951]_  & \new_[40948]_ ;
  assign \new_[40955]_  = ~A300 & ~A268;
  assign \new_[40958]_  = ~A302 & ~A301;
  assign \new_[40959]_  = \new_[40958]_  & \new_[40955]_ ;
  assign \new_[40960]_  = \new_[40959]_  & \new_[40952]_ ;
  assign \new_[40964]_  = A200 & A199;
  assign \new_[40965]_  = A169 & \new_[40964]_ ;
  assign \new_[40968]_  = ~A202 & ~A201;
  assign \new_[40971]_  = ~A233 & ~A232;
  assign \new_[40972]_  = \new_[40971]_  & \new_[40968]_ ;
  assign \new_[40973]_  = \new_[40972]_  & \new_[40965]_ ;
  assign \new_[40976]_  = A265 & ~A235;
  assign \new_[40979]_  = ~A267 & A266;
  assign \new_[40980]_  = \new_[40979]_  & \new_[40976]_ ;
  assign \new_[40983]_  = ~A298 & ~A268;
  assign \new_[40986]_  = ~A301 & ~A299;
  assign \new_[40987]_  = \new_[40986]_  & \new_[40983]_ ;
  assign \new_[40988]_  = \new_[40987]_  & \new_[40980]_ ;
  assign \new_[40992]_  = A200 & A199;
  assign \new_[40993]_  = A169 & \new_[40992]_ ;
  assign \new_[40996]_  = ~A202 & ~A201;
  assign \new_[40999]_  = ~A233 & ~A232;
  assign \new_[41000]_  = \new_[40999]_  & \new_[40996]_ ;
  assign \new_[41001]_  = \new_[41000]_  & \new_[40993]_ ;
  assign \new_[41004]_  = ~A265 & ~A235;
  assign \new_[41007]_  = ~A268 & ~A266;
  assign \new_[41008]_  = \new_[41007]_  & \new_[41004]_ ;
  assign \new_[41011]_  = A299 & A298;
  assign \new_[41014]_  = ~A301 & ~A300;
  assign \new_[41015]_  = \new_[41014]_  & \new_[41011]_ ;
  assign \new_[41016]_  = \new_[41015]_  & \new_[41008]_ ;
  assign \new_[41020]_  = ~A200 & ~A199;
  assign \new_[41021]_  = A169 & \new_[41020]_ ;
  assign \new_[41024]_  = ~A234 & ~A202;
  assign \new_[41027]_  = ~A236 & ~A235;
  assign \new_[41028]_  = \new_[41027]_  & \new_[41024]_ ;
  assign \new_[41029]_  = \new_[41028]_  & \new_[41021]_ ;
  assign \new_[41032]_  = A266 & A265;
  assign \new_[41035]_  = ~A268 & ~A267;
  assign \new_[41036]_  = \new_[41035]_  & \new_[41032]_ ;
  assign \new_[41039]_  = A299 & A298;
  assign \new_[41042]_  = ~A301 & ~A300;
  assign \new_[41043]_  = \new_[41042]_  & \new_[41039]_ ;
  assign \new_[41044]_  = \new_[41043]_  & \new_[41036]_ ;
  assign \new_[41048]_  = ~A200 & ~A199;
  assign \new_[41049]_  = A169 & \new_[41048]_ ;
  assign \new_[41052]_  = A232 & ~A202;
  assign \new_[41055]_  = ~A234 & A233;
  assign \new_[41056]_  = \new_[41055]_  & \new_[41052]_ ;
  assign \new_[41057]_  = \new_[41056]_  & \new_[41049]_ ;
  assign \new_[41060]_  = ~A267 & ~A235;
  assign \new_[41063]_  = ~A269 & ~A268;
  assign \new_[41064]_  = \new_[41063]_  & \new_[41060]_ ;
  assign \new_[41067]_  = A299 & A298;
  assign \new_[41070]_  = ~A301 & ~A300;
  assign \new_[41071]_  = \new_[41070]_  & \new_[41067]_ ;
  assign \new_[41072]_  = \new_[41071]_  & \new_[41064]_ ;
  assign \new_[41076]_  = ~A200 & ~A199;
  assign \new_[41077]_  = A169 & \new_[41076]_ ;
  assign \new_[41080]_  = A232 & ~A202;
  assign \new_[41083]_  = ~A234 & A233;
  assign \new_[41084]_  = \new_[41083]_  & \new_[41080]_ ;
  assign \new_[41085]_  = \new_[41084]_  & \new_[41077]_ ;
  assign \new_[41088]_  = A265 & ~A235;
  assign \new_[41091]_  = ~A267 & A266;
  assign \new_[41092]_  = \new_[41091]_  & \new_[41088]_ ;
  assign \new_[41095]_  = ~A300 & ~A268;
  assign \new_[41098]_  = ~A302 & ~A301;
  assign \new_[41099]_  = \new_[41098]_  & \new_[41095]_ ;
  assign \new_[41100]_  = \new_[41099]_  & \new_[41092]_ ;
  assign \new_[41104]_  = ~A200 & ~A199;
  assign \new_[41105]_  = A169 & \new_[41104]_ ;
  assign \new_[41108]_  = A232 & ~A202;
  assign \new_[41111]_  = ~A234 & A233;
  assign \new_[41112]_  = \new_[41111]_  & \new_[41108]_ ;
  assign \new_[41113]_  = \new_[41112]_  & \new_[41105]_ ;
  assign \new_[41116]_  = A265 & ~A235;
  assign \new_[41119]_  = ~A267 & A266;
  assign \new_[41120]_  = \new_[41119]_  & \new_[41116]_ ;
  assign \new_[41123]_  = ~A298 & ~A268;
  assign \new_[41126]_  = ~A301 & ~A299;
  assign \new_[41127]_  = \new_[41126]_  & \new_[41123]_ ;
  assign \new_[41128]_  = \new_[41127]_  & \new_[41120]_ ;
  assign \new_[41132]_  = ~A200 & ~A199;
  assign \new_[41133]_  = A169 & \new_[41132]_ ;
  assign \new_[41136]_  = A232 & ~A202;
  assign \new_[41139]_  = ~A234 & A233;
  assign \new_[41140]_  = \new_[41139]_  & \new_[41136]_ ;
  assign \new_[41141]_  = \new_[41140]_  & \new_[41133]_ ;
  assign \new_[41144]_  = ~A265 & ~A235;
  assign \new_[41147]_  = ~A268 & ~A266;
  assign \new_[41148]_  = \new_[41147]_  & \new_[41144]_ ;
  assign \new_[41151]_  = A299 & A298;
  assign \new_[41154]_  = ~A301 & ~A300;
  assign \new_[41155]_  = \new_[41154]_  & \new_[41151]_ ;
  assign \new_[41156]_  = \new_[41155]_  & \new_[41148]_ ;
  assign \new_[41160]_  = ~A200 & ~A199;
  assign \new_[41161]_  = A169 & \new_[41160]_ ;
  assign \new_[41164]_  = ~A232 & ~A202;
  assign \new_[41167]_  = ~A235 & ~A233;
  assign \new_[41168]_  = \new_[41167]_  & \new_[41164]_ ;
  assign \new_[41169]_  = \new_[41168]_  & \new_[41161]_ ;
  assign \new_[41172]_  = A266 & A265;
  assign \new_[41175]_  = ~A268 & ~A267;
  assign \new_[41176]_  = \new_[41175]_  & \new_[41172]_ ;
  assign \new_[41179]_  = A299 & A298;
  assign \new_[41182]_  = ~A301 & ~A300;
  assign \new_[41183]_  = \new_[41182]_  & \new_[41179]_ ;
  assign \new_[41184]_  = \new_[41183]_  & \new_[41176]_ ;
  assign \new_[41188]_  = ~A166 & ~A167;
  assign \new_[41189]_  = ~A169 & \new_[41188]_ ;
  assign \new_[41192]_  = ~A234 & A202;
  assign \new_[41195]_  = ~A236 & ~A235;
  assign \new_[41196]_  = \new_[41195]_  & \new_[41192]_ ;
  assign \new_[41197]_  = \new_[41196]_  & \new_[41189]_ ;
  assign \new_[41200]_  = A266 & A265;
  assign \new_[41203]_  = ~A268 & ~A267;
  assign \new_[41204]_  = \new_[41203]_  & \new_[41200]_ ;
  assign \new_[41207]_  = A299 & A298;
  assign \new_[41210]_  = ~A301 & ~A300;
  assign \new_[41211]_  = \new_[41210]_  & \new_[41207]_ ;
  assign \new_[41212]_  = \new_[41211]_  & \new_[41204]_ ;
  assign \new_[41216]_  = ~A166 & ~A167;
  assign \new_[41217]_  = ~A169 & \new_[41216]_ ;
  assign \new_[41220]_  = A232 & A202;
  assign \new_[41223]_  = ~A234 & A233;
  assign \new_[41224]_  = \new_[41223]_  & \new_[41220]_ ;
  assign \new_[41225]_  = \new_[41224]_  & \new_[41217]_ ;
  assign \new_[41228]_  = ~A267 & ~A235;
  assign \new_[41231]_  = ~A269 & ~A268;
  assign \new_[41232]_  = \new_[41231]_  & \new_[41228]_ ;
  assign \new_[41235]_  = A299 & A298;
  assign \new_[41238]_  = ~A301 & ~A300;
  assign \new_[41239]_  = \new_[41238]_  & \new_[41235]_ ;
  assign \new_[41240]_  = \new_[41239]_  & \new_[41232]_ ;
  assign \new_[41244]_  = ~A166 & ~A167;
  assign \new_[41245]_  = ~A169 & \new_[41244]_ ;
  assign \new_[41248]_  = A232 & A202;
  assign \new_[41251]_  = ~A234 & A233;
  assign \new_[41252]_  = \new_[41251]_  & \new_[41248]_ ;
  assign \new_[41253]_  = \new_[41252]_  & \new_[41245]_ ;
  assign \new_[41256]_  = A265 & ~A235;
  assign \new_[41259]_  = ~A267 & A266;
  assign \new_[41260]_  = \new_[41259]_  & \new_[41256]_ ;
  assign \new_[41263]_  = ~A300 & ~A268;
  assign \new_[41266]_  = ~A302 & ~A301;
  assign \new_[41267]_  = \new_[41266]_  & \new_[41263]_ ;
  assign \new_[41268]_  = \new_[41267]_  & \new_[41260]_ ;
  assign \new_[41272]_  = ~A166 & ~A167;
  assign \new_[41273]_  = ~A169 & \new_[41272]_ ;
  assign \new_[41276]_  = A232 & A202;
  assign \new_[41279]_  = ~A234 & A233;
  assign \new_[41280]_  = \new_[41279]_  & \new_[41276]_ ;
  assign \new_[41281]_  = \new_[41280]_  & \new_[41273]_ ;
  assign \new_[41284]_  = A265 & ~A235;
  assign \new_[41287]_  = ~A267 & A266;
  assign \new_[41288]_  = \new_[41287]_  & \new_[41284]_ ;
  assign \new_[41291]_  = ~A298 & ~A268;
  assign \new_[41294]_  = ~A301 & ~A299;
  assign \new_[41295]_  = \new_[41294]_  & \new_[41291]_ ;
  assign \new_[41296]_  = \new_[41295]_  & \new_[41288]_ ;
  assign \new_[41300]_  = ~A166 & ~A167;
  assign \new_[41301]_  = ~A169 & \new_[41300]_ ;
  assign \new_[41304]_  = A232 & A202;
  assign \new_[41307]_  = ~A234 & A233;
  assign \new_[41308]_  = \new_[41307]_  & \new_[41304]_ ;
  assign \new_[41309]_  = \new_[41308]_  & \new_[41301]_ ;
  assign \new_[41312]_  = ~A265 & ~A235;
  assign \new_[41315]_  = ~A268 & ~A266;
  assign \new_[41316]_  = \new_[41315]_  & \new_[41312]_ ;
  assign \new_[41319]_  = A299 & A298;
  assign \new_[41322]_  = ~A301 & ~A300;
  assign \new_[41323]_  = \new_[41322]_  & \new_[41319]_ ;
  assign \new_[41324]_  = \new_[41323]_  & \new_[41316]_ ;
  assign \new_[41328]_  = ~A166 & ~A167;
  assign \new_[41329]_  = ~A169 & \new_[41328]_ ;
  assign \new_[41332]_  = ~A232 & A202;
  assign \new_[41335]_  = ~A235 & ~A233;
  assign \new_[41336]_  = \new_[41335]_  & \new_[41332]_ ;
  assign \new_[41337]_  = \new_[41336]_  & \new_[41329]_ ;
  assign \new_[41340]_  = A266 & A265;
  assign \new_[41343]_  = ~A268 & ~A267;
  assign \new_[41344]_  = \new_[41343]_  & \new_[41340]_ ;
  assign \new_[41347]_  = A299 & A298;
  assign \new_[41350]_  = ~A301 & ~A300;
  assign \new_[41351]_  = \new_[41350]_  & \new_[41347]_ ;
  assign \new_[41352]_  = \new_[41351]_  & \new_[41344]_ ;
  assign \new_[41356]_  = ~A166 & ~A167;
  assign \new_[41357]_  = ~A169 & \new_[41356]_ ;
  assign \new_[41360]_  = A201 & A199;
  assign \new_[41363]_  = ~A235 & ~A234;
  assign \new_[41364]_  = \new_[41363]_  & \new_[41360]_ ;
  assign \new_[41365]_  = \new_[41364]_  & \new_[41357]_ ;
  assign \new_[41368]_  = ~A267 & ~A236;
  assign \new_[41371]_  = ~A269 & ~A268;
  assign \new_[41372]_  = \new_[41371]_  & \new_[41368]_ ;
  assign \new_[41375]_  = A299 & A298;
  assign \new_[41378]_  = ~A301 & ~A300;
  assign \new_[41379]_  = \new_[41378]_  & \new_[41375]_ ;
  assign \new_[41380]_  = \new_[41379]_  & \new_[41372]_ ;
  assign \new_[41384]_  = ~A166 & ~A167;
  assign \new_[41385]_  = ~A169 & \new_[41384]_ ;
  assign \new_[41388]_  = A201 & A199;
  assign \new_[41391]_  = ~A235 & ~A234;
  assign \new_[41392]_  = \new_[41391]_  & \new_[41388]_ ;
  assign \new_[41393]_  = \new_[41392]_  & \new_[41385]_ ;
  assign \new_[41396]_  = A265 & ~A236;
  assign \new_[41399]_  = ~A267 & A266;
  assign \new_[41400]_  = \new_[41399]_  & \new_[41396]_ ;
  assign \new_[41403]_  = ~A300 & ~A268;
  assign \new_[41406]_  = ~A302 & ~A301;
  assign \new_[41407]_  = \new_[41406]_  & \new_[41403]_ ;
  assign \new_[41408]_  = \new_[41407]_  & \new_[41400]_ ;
  assign \new_[41412]_  = ~A166 & ~A167;
  assign \new_[41413]_  = ~A169 & \new_[41412]_ ;
  assign \new_[41416]_  = A201 & A199;
  assign \new_[41419]_  = ~A235 & ~A234;
  assign \new_[41420]_  = \new_[41419]_  & \new_[41416]_ ;
  assign \new_[41421]_  = \new_[41420]_  & \new_[41413]_ ;
  assign \new_[41424]_  = A265 & ~A236;
  assign \new_[41427]_  = ~A267 & A266;
  assign \new_[41428]_  = \new_[41427]_  & \new_[41424]_ ;
  assign \new_[41431]_  = ~A298 & ~A268;
  assign \new_[41434]_  = ~A301 & ~A299;
  assign \new_[41435]_  = \new_[41434]_  & \new_[41431]_ ;
  assign \new_[41436]_  = \new_[41435]_  & \new_[41428]_ ;
  assign \new_[41440]_  = ~A166 & ~A167;
  assign \new_[41441]_  = ~A169 & \new_[41440]_ ;
  assign \new_[41444]_  = A201 & A199;
  assign \new_[41447]_  = ~A235 & ~A234;
  assign \new_[41448]_  = \new_[41447]_  & \new_[41444]_ ;
  assign \new_[41449]_  = \new_[41448]_  & \new_[41441]_ ;
  assign \new_[41452]_  = ~A265 & ~A236;
  assign \new_[41455]_  = ~A268 & ~A266;
  assign \new_[41456]_  = \new_[41455]_  & \new_[41452]_ ;
  assign \new_[41459]_  = A299 & A298;
  assign \new_[41462]_  = ~A301 & ~A300;
  assign \new_[41463]_  = \new_[41462]_  & \new_[41459]_ ;
  assign \new_[41464]_  = \new_[41463]_  & \new_[41456]_ ;
  assign \new_[41468]_  = ~A166 & ~A167;
  assign \new_[41469]_  = ~A169 & \new_[41468]_ ;
  assign \new_[41472]_  = A201 & A199;
  assign \new_[41475]_  = A233 & A232;
  assign \new_[41476]_  = \new_[41475]_  & \new_[41472]_ ;
  assign \new_[41477]_  = \new_[41476]_  & \new_[41469]_ ;
  assign \new_[41480]_  = ~A235 & ~A234;
  assign \new_[41483]_  = ~A268 & ~A267;
  assign \new_[41484]_  = \new_[41483]_  & \new_[41480]_ ;
  assign \new_[41487]_  = ~A300 & ~A269;
  assign \new_[41490]_  = ~A302 & ~A301;
  assign \new_[41491]_  = \new_[41490]_  & \new_[41487]_ ;
  assign \new_[41492]_  = \new_[41491]_  & \new_[41484]_ ;
  assign \new_[41496]_  = ~A166 & ~A167;
  assign \new_[41497]_  = ~A169 & \new_[41496]_ ;
  assign \new_[41500]_  = A201 & A199;
  assign \new_[41503]_  = A233 & A232;
  assign \new_[41504]_  = \new_[41503]_  & \new_[41500]_ ;
  assign \new_[41505]_  = \new_[41504]_  & \new_[41497]_ ;
  assign \new_[41508]_  = ~A235 & ~A234;
  assign \new_[41511]_  = ~A268 & ~A267;
  assign \new_[41512]_  = \new_[41511]_  & \new_[41508]_ ;
  assign \new_[41515]_  = ~A298 & ~A269;
  assign \new_[41518]_  = ~A301 & ~A299;
  assign \new_[41519]_  = \new_[41518]_  & \new_[41515]_ ;
  assign \new_[41520]_  = \new_[41519]_  & \new_[41512]_ ;
  assign \new_[41524]_  = ~A166 & ~A167;
  assign \new_[41525]_  = ~A169 & \new_[41524]_ ;
  assign \new_[41528]_  = A201 & A199;
  assign \new_[41531]_  = A233 & A232;
  assign \new_[41532]_  = \new_[41531]_  & \new_[41528]_ ;
  assign \new_[41533]_  = \new_[41532]_  & \new_[41525]_ ;
  assign \new_[41536]_  = ~A235 & ~A234;
  assign \new_[41539]_  = ~A266 & ~A265;
  assign \new_[41540]_  = \new_[41539]_  & \new_[41536]_ ;
  assign \new_[41543]_  = ~A300 & ~A268;
  assign \new_[41546]_  = ~A302 & ~A301;
  assign \new_[41547]_  = \new_[41546]_  & \new_[41543]_ ;
  assign \new_[41548]_  = \new_[41547]_  & \new_[41540]_ ;
  assign \new_[41552]_  = ~A166 & ~A167;
  assign \new_[41553]_  = ~A169 & \new_[41552]_ ;
  assign \new_[41556]_  = A201 & A199;
  assign \new_[41559]_  = A233 & A232;
  assign \new_[41560]_  = \new_[41559]_  & \new_[41556]_ ;
  assign \new_[41561]_  = \new_[41560]_  & \new_[41553]_ ;
  assign \new_[41564]_  = ~A235 & ~A234;
  assign \new_[41567]_  = ~A266 & ~A265;
  assign \new_[41568]_  = \new_[41567]_  & \new_[41564]_ ;
  assign \new_[41571]_  = ~A298 & ~A268;
  assign \new_[41574]_  = ~A301 & ~A299;
  assign \new_[41575]_  = \new_[41574]_  & \new_[41571]_ ;
  assign \new_[41576]_  = \new_[41575]_  & \new_[41568]_ ;
  assign \new_[41580]_  = ~A166 & ~A167;
  assign \new_[41581]_  = ~A169 & \new_[41580]_ ;
  assign \new_[41584]_  = A201 & A199;
  assign \new_[41587]_  = ~A233 & ~A232;
  assign \new_[41588]_  = \new_[41587]_  & \new_[41584]_ ;
  assign \new_[41589]_  = \new_[41588]_  & \new_[41581]_ ;
  assign \new_[41592]_  = ~A267 & ~A235;
  assign \new_[41595]_  = ~A269 & ~A268;
  assign \new_[41596]_  = \new_[41595]_  & \new_[41592]_ ;
  assign \new_[41599]_  = A299 & A298;
  assign \new_[41602]_  = ~A301 & ~A300;
  assign \new_[41603]_  = \new_[41602]_  & \new_[41599]_ ;
  assign \new_[41604]_  = \new_[41603]_  & \new_[41596]_ ;
  assign \new_[41608]_  = ~A166 & ~A167;
  assign \new_[41609]_  = ~A169 & \new_[41608]_ ;
  assign \new_[41612]_  = A201 & A199;
  assign \new_[41615]_  = ~A233 & ~A232;
  assign \new_[41616]_  = \new_[41615]_  & \new_[41612]_ ;
  assign \new_[41617]_  = \new_[41616]_  & \new_[41609]_ ;
  assign \new_[41620]_  = A265 & ~A235;
  assign \new_[41623]_  = ~A267 & A266;
  assign \new_[41624]_  = \new_[41623]_  & \new_[41620]_ ;
  assign \new_[41627]_  = ~A300 & ~A268;
  assign \new_[41630]_  = ~A302 & ~A301;
  assign \new_[41631]_  = \new_[41630]_  & \new_[41627]_ ;
  assign \new_[41632]_  = \new_[41631]_  & \new_[41624]_ ;
  assign \new_[41636]_  = ~A166 & ~A167;
  assign \new_[41637]_  = ~A169 & \new_[41636]_ ;
  assign \new_[41640]_  = A201 & A199;
  assign \new_[41643]_  = ~A233 & ~A232;
  assign \new_[41644]_  = \new_[41643]_  & \new_[41640]_ ;
  assign \new_[41645]_  = \new_[41644]_  & \new_[41637]_ ;
  assign \new_[41648]_  = A265 & ~A235;
  assign \new_[41651]_  = ~A267 & A266;
  assign \new_[41652]_  = \new_[41651]_  & \new_[41648]_ ;
  assign \new_[41655]_  = ~A298 & ~A268;
  assign \new_[41658]_  = ~A301 & ~A299;
  assign \new_[41659]_  = \new_[41658]_  & \new_[41655]_ ;
  assign \new_[41660]_  = \new_[41659]_  & \new_[41652]_ ;
  assign \new_[41664]_  = ~A166 & ~A167;
  assign \new_[41665]_  = ~A169 & \new_[41664]_ ;
  assign \new_[41668]_  = A201 & A199;
  assign \new_[41671]_  = ~A233 & ~A232;
  assign \new_[41672]_  = \new_[41671]_  & \new_[41668]_ ;
  assign \new_[41673]_  = \new_[41672]_  & \new_[41665]_ ;
  assign \new_[41676]_  = ~A265 & ~A235;
  assign \new_[41679]_  = ~A268 & ~A266;
  assign \new_[41680]_  = \new_[41679]_  & \new_[41676]_ ;
  assign \new_[41683]_  = A299 & A298;
  assign \new_[41686]_  = ~A301 & ~A300;
  assign \new_[41687]_  = \new_[41686]_  & \new_[41683]_ ;
  assign \new_[41688]_  = \new_[41687]_  & \new_[41680]_ ;
  assign \new_[41692]_  = ~A166 & ~A167;
  assign \new_[41693]_  = ~A169 & \new_[41692]_ ;
  assign \new_[41696]_  = A201 & A200;
  assign \new_[41699]_  = ~A235 & ~A234;
  assign \new_[41700]_  = \new_[41699]_  & \new_[41696]_ ;
  assign \new_[41701]_  = \new_[41700]_  & \new_[41693]_ ;
  assign \new_[41704]_  = ~A267 & ~A236;
  assign \new_[41707]_  = ~A269 & ~A268;
  assign \new_[41708]_  = \new_[41707]_  & \new_[41704]_ ;
  assign \new_[41711]_  = A299 & A298;
  assign \new_[41714]_  = ~A301 & ~A300;
  assign \new_[41715]_  = \new_[41714]_  & \new_[41711]_ ;
  assign \new_[41716]_  = \new_[41715]_  & \new_[41708]_ ;
  assign \new_[41720]_  = ~A166 & ~A167;
  assign \new_[41721]_  = ~A169 & \new_[41720]_ ;
  assign \new_[41724]_  = A201 & A200;
  assign \new_[41727]_  = ~A235 & ~A234;
  assign \new_[41728]_  = \new_[41727]_  & \new_[41724]_ ;
  assign \new_[41729]_  = \new_[41728]_  & \new_[41721]_ ;
  assign \new_[41732]_  = A265 & ~A236;
  assign \new_[41735]_  = ~A267 & A266;
  assign \new_[41736]_  = \new_[41735]_  & \new_[41732]_ ;
  assign \new_[41739]_  = ~A300 & ~A268;
  assign \new_[41742]_  = ~A302 & ~A301;
  assign \new_[41743]_  = \new_[41742]_  & \new_[41739]_ ;
  assign \new_[41744]_  = \new_[41743]_  & \new_[41736]_ ;
  assign \new_[41748]_  = ~A166 & ~A167;
  assign \new_[41749]_  = ~A169 & \new_[41748]_ ;
  assign \new_[41752]_  = A201 & A200;
  assign \new_[41755]_  = ~A235 & ~A234;
  assign \new_[41756]_  = \new_[41755]_  & \new_[41752]_ ;
  assign \new_[41757]_  = \new_[41756]_  & \new_[41749]_ ;
  assign \new_[41760]_  = A265 & ~A236;
  assign \new_[41763]_  = ~A267 & A266;
  assign \new_[41764]_  = \new_[41763]_  & \new_[41760]_ ;
  assign \new_[41767]_  = ~A298 & ~A268;
  assign \new_[41770]_  = ~A301 & ~A299;
  assign \new_[41771]_  = \new_[41770]_  & \new_[41767]_ ;
  assign \new_[41772]_  = \new_[41771]_  & \new_[41764]_ ;
  assign \new_[41776]_  = ~A166 & ~A167;
  assign \new_[41777]_  = ~A169 & \new_[41776]_ ;
  assign \new_[41780]_  = A201 & A200;
  assign \new_[41783]_  = ~A235 & ~A234;
  assign \new_[41784]_  = \new_[41783]_  & \new_[41780]_ ;
  assign \new_[41785]_  = \new_[41784]_  & \new_[41777]_ ;
  assign \new_[41788]_  = ~A265 & ~A236;
  assign \new_[41791]_  = ~A268 & ~A266;
  assign \new_[41792]_  = \new_[41791]_  & \new_[41788]_ ;
  assign \new_[41795]_  = A299 & A298;
  assign \new_[41798]_  = ~A301 & ~A300;
  assign \new_[41799]_  = \new_[41798]_  & \new_[41795]_ ;
  assign \new_[41800]_  = \new_[41799]_  & \new_[41792]_ ;
  assign \new_[41804]_  = ~A166 & ~A167;
  assign \new_[41805]_  = ~A169 & \new_[41804]_ ;
  assign \new_[41808]_  = A201 & A200;
  assign \new_[41811]_  = A233 & A232;
  assign \new_[41812]_  = \new_[41811]_  & \new_[41808]_ ;
  assign \new_[41813]_  = \new_[41812]_  & \new_[41805]_ ;
  assign \new_[41816]_  = ~A235 & ~A234;
  assign \new_[41819]_  = ~A268 & ~A267;
  assign \new_[41820]_  = \new_[41819]_  & \new_[41816]_ ;
  assign \new_[41823]_  = ~A300 & ~A269;
  assign \new_[41826]_  = ~A302 & ~A301;
  assign \new_[41827]_  = \new_[41826]_  & \new_[41823]_ ;
  assign \new_[41828]_  = \new_[41827]_  & \new_[41820]_ ;
  assign \new_[41832]_  = ~A166 & ~A167;
  assign \new_[41833]_  = ~A169 & \new_[41832]_ ;
  assign \new_[41836]_  = A201 & A200;
  assign \new_[41839]_  = A233 & A232;
  assign \new_[41840]_  = \new_[41839]_  & \new_[41836]_ ;
  assign \new_[41841]_  = \new_[41840]_  & \new_[41833]_ ;
  assign \new_[41844]_  = ~A235 & ~A234;
  assign \new_[41847]_  = ~A268 & ~A267;
  assign \new_[41848]_  = \new_[41847]_  & \new_[41844]_ ;
  assign \new_[41851]_  = ~A298 & ~A269;
  assign \new_[41854]_  = ~A301 & ~A299;
  assign \new_[41855]_  = \new_[41854]_  & \new_[41851]_ ;
  assign \new_[41856]_  = \new_[41855]_  & \new_[41848]_ ;
  assign \new_[41860]_  = ~A166 & ~A167;
  assign \new_[41861]_  = ~A169 & \new_[41860]_ ;
  assign \new_[41864]_  = A201 & A200;
  assign \new_[41867]_  = A233 & A232;
  assign \new_[41868]_  = \new_[41867]_  & \new_[41864]_ ;
  assign \new_[41869]_  = \new_[41868]_  & \new_[41861]_ ;
  assign \new_[41872]_  = ~A235 & ~A234;
  assign \new_[41875]_  = ~A266 & ~A265;
  assign \new_[41876]_  = \new_[41875]_  & \new_[41872]_ ;
  assign \new_[41879]_  = ~A300 & ~A268;
  assign \new_[41882]_  = ~A302 & ~A301;
  assign \new_[41883]_  = \new_[41882]_  & \new_[41879]_ ;
  assign \new_[41884]_  = \new_[41883]_  & \new_[41876]_ ;
  assign \new_[41888]_  = ~A166 & ~A167;
  assign \new_[41889]_  = ~A169 & \new_[41888]_ ;
  assign \new_[41892]_  = A201 & A200;
  assign \new_[41895]_  = A233 & A232;
  assign \new_[41896]_  = \new_[41895]_  & \new_[41892]_ ;
  assign \new_[41897]_  = \new_[41896]_  & \new_[41889]_ ;
  assign \new_[41900]_  = ~A235 & ~A234;
  assign \new_[41903]_  = ~A266 & ~A265;
  assign \new_[41904]_  = \new_[41903]_  & \new_[41900]_ ;
  assign \new_[41907]_  = ~A298 & ~A268;
  assign \new_[41910]_  = ~A301 & ~A299;
  assign \new_[41911]_  = \new_[41910]_  & \new_[41907]_ ;
  assign \new_[41912]_  = \new_[41911]_  & \new_[41904]_ ;
  assign \new_[41916]_  = ~A166 & ~A167;
  assign \new_[41917]_  = ~A169 & \new_[41916]_ ;
  assign \new_[41920]_  = A201 & A200;
  assign \new_[41923]_  = ~A233 & ~A232;
  assign \new_[41924]_  = \new_[41923]_  & \new_[41920]_ ;
  assign \new_[41925]_  = \new_[41924]_  & \new_[41917]_ ;
  assign \new_[41928]_  = ~A267 & ~A235;
  assign \new_[41931]_  = ~A269 & ~A268;
  assign \new_[41932]_  = \new_[41931]_  & \new_[41928]_ ;
  assign \new_[41935]_  = A299 & A298;
  assign \new_[41938]_  = ~A301 & ~A300;
  assign \new_[41939]_  = \new_[41938]_  & \new_[41935]_ ;
  assign \new_[41940]_  = \new_[41939]_  & \new_[41932]_ ;
  assign \new_[41944]_  = ~A166 & ~A167;
  assign \new_[41945]_  = ~A169 & \new_[41944]_ ;
  assign \new_[41948]_  = A201 & A200;
  assign \new_[41951]_  = ~A233 & ~A232;
  assign \new_[41952]_  = \new_[41951]_  & \new_[41948]_ ;
  assign \new_[41953]_  = \new_[41952]_  & \new_[41945]_ ;
  assign \new_[41956]_  = A265 & ~A235;
  assign \new_[41959]_  = ~A267 & A266;
  assign \new_[41960]_  = \new_[41959]_  & \new_[41956]_ ;
  assign \new_[41963]_  = ~A300 & ~A268;
  assign \new_[41966]_  = ~A302 & ~A301;
  assign \new_[41967]_  = \new_[41966]_  & \new_[41963]_ ;
  assign \new_[41968]_  = \new_[41967]_  & \new_[41960]_ ;
  assign \new_[41972]_  = ~A166 & ~A167;
  assign \new_[41973]_  = ~A169 & \new_[41972]_ ;
  assign \new_[41976]_  = A201 & A200;
  assign \new_[41979]_  = ~A233 & ~A232;
  assign \new_[41980]_  = \new_[41979]_  & \new_[41976]_ ;
  assign \new_[41981]_  = \new_[41980]_  & \new_[41973]_ ;
  assign \new_[41984]_  = A265 & ~A235;
  assign \new_[41987]_  = ~A267 & A266;
  assign \new_[41988]_  = \new_[41987]_  & \new_[41984]_ ;
  assign \new_[41991]_  = ~A298 & ~A268;
  assign \new_[41994]_  = ~A301 & ~A299;
  assign \new_[41995]_  = \new_[41994]_  & \new_[41991]_ ;
  assign \new_[41996]_  = \new_[41995]_  & \new_[41988]_ ;
  assign \new_[42000]_  = ~A166 & ~A167;
  assign \new_[42001]_  = ~A169 & \new_[42000]_ ;
  assign \new_[42004]_  = A201 & A200;
  assign \new_[42007]_  = ~A233 & ~A232;
  assign \new_[42008]_  = \new_[42007]_  & \new_[42004]_ ;
  assign \new_[42009]_  = \new_[42008]_  & \new_[42001]_ ;
  assign \new_[42012]_  = ~A265 & ~A235;
  assign \new_[42015]_  = ~A268 & ~A266;
  assign \new_[42016]_  = \new_[42015]_  & \new_[42012]_ ;
  assign \new_[42019]_  = A299 & A298;
  assign \new_[42022]_  = ~A301 & ~A300;
  assign \new_[42023]_  = \new_[42022]_  & \new_[42019]_ ;
  assign \new_[42024]_  = \new_[42023]_  & \new_[42016]_ ;
  assign \new_[42028]_  = ~A166 & ~A167;
  assign \new_[42029]_  = ~A169 & \new_[42028]_ ;
  assign \new_[42032]_  = A200 & ~A199;
  assign \new_[42035]_  = ~A234 & A203;
  assign \new_[42036]_  = \new_[42035]_  & \new_[42032]_ ;
  assign \new_[42037]_  = \new_[42036]_  & \new_[42029]_ ;
  assign \new_[42040]_  = ~A236 & ~A235;
  assign \new_[42043]_  = ~A268 & ~A267;
  assign \new_[42044]_  = \new_[42043]_  & \new_[42040]_ ;
  assign \new_[42047]_  = ~A300 & ~A269;
  assign \new_[42050]_  = ~A302 & ~A301;
  assign \new_[42051]_  = \new_[42050]_  & \new_[42047]_ ;
  assign \new_[42052]_  = \new_[42051]_  & \new_[42044]_ ;
  assign \new_[42056]_  = ~A166 & ~A167;
  assign \new_[42057]_  = ~A169 & \new_[42056]_ ;
  assign \new_[42060]_  = A200 & ~A199;
  assign \new_[42063]_  = ~A234 & A203;
  assign \new_[42064]_  = \new_[42063]_  & \new_[42060]_ ;
  assign \new_[42065]_  = \new_[42064]_  & \new_[42057]_ ;
  assign \new_[42068]_  = ~A236 & ~A235;
  assign \new_[42071]_  = ~A268 & ~A267;
  assign \new_[42072]_  = \new_[42071]_  & \new_[42068]_ ;
  assign \new_[42075]_  = ~A298 & ~A269;
  assign \new_[42078]_  = ~A301 & ~A299;
  assign \new_[42079]_  = \new_[42078]_  & \new_[42075]_ ;
  assign \new_[42080]_  = \new_[42079]_  & \new_[42072]_ ;
  assign \new_[42084]_  = ~A166 & ~A167;
  assign \new_[42085]_  = ~A169 & \new_[42084]_ ;
  assign \new_[42088]_  = A200 & ~A199;
  assign \new_[42091]_  = ~A234 & A203;
  assign \new_[42092]_  = \new_[42091]_  & \new_[42088]_ ;
  assign \new_[42093]_  = \new_[42092]_  & \new_[42085]_ ;
  assign \new_[42096]_  = ~A236 & ~A235;
  assign \new_[42099]_  = ~A266 & ~A265;
  assign \new_[42100]_  = \new_[42099]_  & \new_[42096]_ ;
  assign \new_[42103]_  = ~A300 & ~A268;
  assign \new_[42106]_  = ~A302 & ~A301;
  assign \new_[42107]_  = \new_[42106]_  & \new_[42103]_ ;
  assign \new_[42108]_  = \new_[42107]_  & \new_[42100]_ ;
  assign \new_[42112]_  = ~A166 & ~A167;
  assign \new_[42113]_  = ~A169 & \new_[42112]_ ;
  assign \new_[42116]_  = A200 & ~A199;
  assign \new_[42119]_  = ~A234 & A203;
  assign \new_[42120]_  = \new_[42119]_  & \new_[42116]_ ;
  assign \new_[42121]_  = \new_[42120]_  & \new_[42113]_ ;
  assign \new_[42124]_  = ~A236 & ~A235;
  assign \new_[42127]_  = ~A266 & ~A265;
  assign \new_[42128]_  = \new_[42127]_  & \new_[42124]_ ;
  assign \new_[42131]_  = ~A298 & ~A268;
  assign \new_[42134]_  = ~A301 & ~A299;
  assign \new_[42135]_  = \new_[42134]_  & \new_[42131]_ ;
  assign \new_[42136]_  = \new_[42135]_  & \new_[42128]_ ;
  assign \new_[42140]_  = ~A166 & ~A167;
  assign \new_[42141]_  = ~A169 & \new_[42140]_ ;
  assign \new_[42144]_  = A200 & ~A199;
  assign \new_[42147]_  = ~A232 & A203;
  assign \new_[42148]_  = \new_[42147]_  & \new_[42144]_ ;
  assign \new_[42149]_  = \new_[42148]_  & \new_[42141]_ ;
  assign \new_[42152]_  = ~A235 & ~A233;
  assign \new_[42155]_  = ~A268 & ~A267;
  assign \new_[42156]_  = \new_[42155]_  & \new_[42152]_ ;
  assign \new_[42159]_  = ~A300 & ~A269;
  assign \new_[42162]_  = ~A302 & ~A301;
  assign \new_[42163]_  = \new_[42162]_  & \new_[42159]_ ;
  assign \new_[42164]_  = \new_[42163]_  & \new_[42156]_ ;
  assign \new_[42168]_  = ~A166 & ~A167;
  assign \new_[42169]_  = ~A169 & \new_[42168]_ ;
  assign \new_[42172]_  = A200 & ~A199;
  assign \new_[42175]_  = ~A232 & A203;
  assign \new_[42176]_  = \new_[42175]_  & \new_[42172]_ ;
  assign \new_[42177]_  = \new_[42176]_  & \new_[42169]_ ;
  assign \new_[42180]_  = ~A235 & ~A233;
  assign \new_[42183]_  = ~A268 & ~A267;
  assign \new_[42184]_  = \new_[42183]_  & \new_[42180]_ ;
  assign \new_[42187]_  = ~A298 & ~A269;
  assign \new_[42190]_  = ~A301 & ~A299;
  assign \new_[42191]_  = \new_[42190]_  & \new_[42187]_ ;
  assign \new_[42192]_  = \new_[42191]_  & \new_[42184]_ ;
  assign \new_[42196]_  = ~A166 & ~A167;
  assign \new_[42197]_  = ~A169 & \new_[42196]_ ;
  assign \new_[42200]_  = A200 & ~A199;
  assign \new_[42203]_  = ~A232 & A203;
  assign \new_[42204]_  = \new_[42203]_  & \new_[42200]_ ;
  assign \new_[42205]_  = \new_[42204]_  & \new_[42197]_ ;
  assign \new_[42208]_  = ~A235 & ~A233;
  assign \new_[42211]_  = ~A266 & ~A265;
  assign \new_[42212]_  = \new_[42211]_  & \new_[42208]_ ;
  assign \new_[42215]_  = ~A300 & ~A268;
  assign \new_[42218]_  = ~A302 & ~A301;
  assign \new_[42219]_  = \new_[42218]_  & \new_[42215]_ ;
  assign \new_[42220]_  = \new_[42219]_  & \new_[42212]_ ;
  assign \new_[42224]_  = ~A166 & ~A167;
  assign \new_[42225]_  = ~A169 & \new_[42224]_ ;
  assign \new_[42228]_  = A200 & ~A199;
  assign \new_[42231]_  = ~A232 & A203;
  assign \new_[42232]_  = \new_[42231]_  & \new_[42228]_ ;
  assign \new_[42233]_  = \new_[42232]_  & \new_[42225]_ ;
  assign \new_[42236]_  = ~A235 & ~A233;
  assign \new_[42239]_  = ~A266 & ~A265;
  assign \new_[42240]_  = \new_[42239]_  & \new_[42236]_ ;
  assign \new_[42243]_  = ~A298 & ~A268;
  assign \new_[42246]_  = ~A301 & ~A299;
  assign \new_[42247]_  = \new_[42246]_  & \new_[42243]_ ;
  assign \new_[42248]_  = \new_[42247]_  & \new_[42240]_ ;
  assign \new_[42252]_  = ~A166 & ~A167;
  assign \new_[42253]_  = ~A169 & \new_[42252]_ ;
  assign \new_[42256]_  = ~A200 & A199;
  assign \new_[42259]_  = ~A234 & A203;
  assign \new_[42260]_  = \new_[42259]_  & \new_[42256]_ ;
  assign \new_[42261]_  = \new_[42260]_  & \new_[42253]_ ;
  assign \new_[42264]_  = ~A236 & ~A235;
  assign \new_[42267]_  = ~A268 & ~A267;
  assign \new_[42268]_  = \new_[42267]_  & \new_[42264]_ ;
  assign \new_[42271]_  = ~A300 & ~A269;
  assign \new_[42274]_  = ~A302 & ~A301;
  assign \new_[42275]_  = \new_[42274]_  & \new_[42271]_ ;
  assign \new_[42276]_  = \new_[42275]_  & \new_[42268]_ ;
  assign \new_[42280]_  = ~A166 & ~A167;
  assign \new_[42281]_  = ~A169 & \new_[42280]_ ;
  assign \new_[42284]_  = ~A200 & A199;
  assign \new_[42287]_  = ~A234 & A203;
  assign \new_[42288]_  = \new_[42287]_  & \new_[42284]_ ;
  assign \new_[42289]_  = \new_[42288]_  & \new_[42281]_ ;
  assign \new_[42292]_  = ~A236 & ~A235;
  assign \new_[42295]_  = ~A268 & ~A267;
  assign \new_[42296]_  = \new_[42295]_  & \new_[42292]_ ;
  assign \new_[42299]_  = ~A298 & ~A269;
  assign \new_[42302]_  = ~A301 & ~A299;
  assign \new_[42303]_  = \new_[42302]_  & \new_[42299]_ ;
  assign \new_[42304]_  = \new_[42303]_  & \new_[42296]_ ;
  assign \new_[42308]_  = ~A166 & ~A167;
  assign \new_[42309]_  = ~A169 & \new_[42308]_ ;
  assign \new_[42312]_  = ~A200 & A199;
  assign \new_[42315]_  = ~A234 & A203;
  assign \new_[42316]_  = \new_[42315]_  & \new_[42312]_ ;
  assign \new_[42317]_  = \new_[42316]_  & \new_[42309]_ ;
  assign \new_[42320]_  = ~A236 & ~A235;
  assign \new_[42323]_  = ~A266 & ~A265;
  assign \new_[42324]_  = \new_[42323]_  & \new_[42320]_ ;
  assign \new_[42327]_  = ~A300 & ~A268;
  assign \new_[42330]_  = ~A302 & ~A301;
  assign \new_[42331]_  = \new_[42330]_  & \new_[42327]_ ;
  assign \new_[42332]_  = \new_[42331]_  & \new_[42324]_ ;
  assign \new_[42336]_  = ~A166 & ~A167;
  assign \new_[42337]_  = ~A169 & \new_[42336]_ ;
  assign \new_[42340]_  = ~A200 & A199;
  assign \new_[42343]_  = ~A234 & A203;
  assign \new_[42344]_  = \new_[42343]_  & \new_[42340]_ ;
  assign \new_[42345]_  = \new_[42344]_  & \new_[42337]_ ;
  assign \new_[42348]_  = ~A236 & ~A235;
  assign \new_[42351]_  = ~A266 & ~A265;
  assign \new_[42352]_  = \new_[42351]_  & \new_[42348]_ ;
  assign \new_[42355]_  = ~A298 & ~A268;
  assign \new_[42358]_  = ~A301 & ~A299;
  assign \new_[42359]_  = \new_[42358]_  & \new_[42355]_ ;
  assign \new_[42360]_  = \new_[42359]_  & \new_[42352]_ ;
  assign \new_[42364]_  = ~A166 & ~A167;
  assign \new_[42365]_  = ~A169 & \new_[42364]_ ;
  assign \new_[42368]_  = ~A200 & A199;
  assign \new_[42371]_  = ~A232 & A203;
  assign \new_[42372]_  = \new_[42371]_  & \new_[42368]_ ;
  assign \new_[42373]_  = \new_[42372]_  & \new_[42365]_ ;
  assign \new_[42376]_  = ~A235 & ~A233;
  assign \new_[42379]_  = ~A268 & ~A267;
  assign \new_[42380]_  = \new_[42379]_  & \new_[42376]_ ;
  assign \new_[42383]_  = ~A300 & ~A269;
  assign \new_[42386]_  = ~A302 & ~A301;
  assign \new_[42387]_  = \new_[42386]_  & \new_[42383]_ ;
  assign \new_[42388]_  = \new_[42387]_  & \new_[42380]_ ;
  assign \new_[42392]_  = ~A166 & ~A167;
  assign \new_[42393]_  = ~A169 & \new_[42392]_ ;
  assign \new_[42396]_  = ~A200 & A199;
  assign \new_[42399]_  = ~A232 & A203;
  assign \new_[42400]_  = \new_[42399]_  & \new_[42396]_ ;
  assign \new_[42401]_  = \new_[42400]_  & \new_[42393]_ ;
  assign \new_[42404]_  = ~A235 & ~A233;
  assign \new_[42407]_  = ~A268 & ~A267;
  assign \new_[42408]_  = \new_[42407]_  & \new_[42404]_ ;
  assign \new_[42411]_  = ~A298 & ~A269;
  assign \new_[42414]_  = ~A301 & ~A299;
  assign \new_[42415]_  = \new_[42414]_  & \new_[42411]_ ;
  assign \new_[42416]_  = \new_[42415]_  & \new_[42408]_ ;
  assign \new_[42420]_  = ~A166 & ~A167;
  assign \new_[42421]_  = ~A169 & \new_[42420]_ ;
  assign \new_[42424]_  = ~A200 & A199;
  assign \new_[42427]_  = ~A232 & A203;
  assign \new_[42428]_  = \new_[42427]_  & \new_[42424]_ ;
  assign \new_[42429]_  = \new_[42428]_  & \new_[42421]_ ;
  assign \new_[42432]_  = ~A235 & ~A233;
  assign \new_[42435]_  = ~A266 & ~A265;
  assign \new_[42436]_  = \new_[42435]_  & \new_[42432]_ ;
  assign \new_[42439]_  = ~A300 & ~A268;
  assign \new_[42442]_  = ~A302 & ~A301;
  assign \new_[42443]_  = \new_[42442]_  & \new_[42439]_ ;
  assign \new_[42444]_  = \new_[42443]_  & \new_[42436]_ ;
  assign \new_[42448]_  = ~A166 & ~A167;
  assign \new_[42449]_  = ~A169 & \new_[42448]_ ;
  assign \new_[42452]_  = ~A200 & A199;
  assign \new_[42455]_  = ~A232 & A203;
  assign \new_[42456]_  = \new_[42455]_  & \new_[42452]_ ;
  assign \new_[42457]_  = \new_[42456]_  & \new_[42449]_ ;
  assign \new_[42460]_  = ~A235 & ~A233;
  assign \new_[42463]_  = ~A266 & ~A265;
  assign \new_[42464]_  = \new_[42463]_  & \new_[42460]_ ;
  assign \new_[42467]_  = ~A298 & ~A268;
  assign \new_[42470]_  = ~A301 & ~A299;
  assign \new_[42471]_  = \new_[42470]_  & \new_[42467]_ ;
  assign \new_[42472]_  = \new_[42471]_  & \new_[42464]_ ;
  assign \new_[42476]_  = A167 & ~A168;
  assign \new_[42477]_  = ~A169 & \new_[42476]_ ;
  assign \new_[42480]_  = A202 & A166;
  assign \new_[42483]_  = ~A235 & ~A234;
  assign \new_[42484]_  = \new_[42483]_  & \new_[42480]_ ;
  assign \new_[42485]_  = \new_[42484]_  & \new_[42477]_ ;
  assign \new_[42488]_  = ~A267 & ~A236;
  assign \new_[42491]_  = ~A269 & ~A268;
  assign \new_[42492]_  = \new_[42491]_  & \new_[42488]_ ;
  assign \new_[42495]_  = A299 & A298;
  assign \new_[42498]_  = ~A301 & ~A300;
  assign \new_[42499]_  = \new_[42498]_  & \new_[42495]_ ;
  assign \new_[42500]_  = \new_[42499]_  & \new_[42492]_ ;
  assign \new_[42504]_  = A167 & ~A168;
  assign \new_[42505]_  = ~A169 & \new_[42504]_ ;
  assign \new_[42508]_  = A202 & A166;
  assign \new_[42511]_  = ~A235 & ~A234;
  assign \new_[42512]_  = \new_[42511]_  & \new_[42508]_ ;
  assign \new_[42513]_  = \new_[42512]_  & \new_[42505]_ ;
  assign \new_[42516]_  = A265 & ~A236;
  assign \new_[42519]_  = ~A267 & A266;
  assign \new_[42520]_  = \new_[42519]_  & \new_[42516]_ ;
  assign \new_[42523]_  = ~A300 & ~A268;
  assign \new_[42526]_  = ~A302 & ~A301;
  assign \new_[42527]_  = \new_[42526]_  & \new_[42523]_ ;
  assign \new_[42528]_  = \new_[42527]_  & \new_[42520]_ ;
  assign \new_[42532]_  = A167 & ~A168;
  assign \new_[42533]_  = ~A169 & \new_[42532]_ ;
  assign \new_[42536]_  = A202 & A166;
  assign \new_[42539]_  = ~A235 & ~A234;
  assign \new_[42540]_  = \new_[42539]_  & \new_[42536]_ ;
  assign \new_[42541]_  = \new_[42540]_  & \new_[42533]_ ;
  assign \new_[42544]_  = A265 & ~A236;
  assign \new_[42547]_  = ~A267 & A266;
  assign \new_[42548]_  = \new_[42547]_  & \new_[42544]_ ;
  assign \new_[42551]_  = ~A298 & ~A268;
  assign \new_[42554]_  = ~A301 & ~A299;
  assign \new_[42555]_  = \new_[42554]_  & \new_[42551]_ ;
  assign \new_[42556]_  = \new_[42555]_  & \new_[42548]_ ;
  assign \new_[42560]_  = A167 & ~A168;
  assign \new_[42561]_  = ~A169 & \new_[42560]_ ;
  assign \new_[42564]_  = A202 & A166;
  assign \new_[42567]_  = ~A235 & ~A234;
  assign \new_[42568]_  = \new_[42567]_  & \new_[42564]_ ;
  assign \new_[42569]_  = \new_[42568]_  & \new_[42561]_ ;
  assign \new_[42572]_  = ~A265 & ~A236;
  assign \new_[42575]_  = ~A268 & ~A266;
  assign \new_[42576]_  = \new_[42575]_  & \new_[42572]_ ;
  assign \new_[42579]_  = A299 & A298;
  assign \new_[42582]_  = ~A301 & ~A300;
  assign \new_[42583]_  = \new_[42582]_  & \new_[42579]_ ;
  assign \new_[42584]_  = \new_[42583]_  & \new_[42576]_ ;
  assign \new_[42588]_  = A167 & ~A168;
  assign \new_[42589]_  = ~A169 & \new_[42588]_ ;
  assign \new_[42592]_  = A202 & A166;
  assign \new_[42595]_  = A233 & A232;
  assign \new_[42596]_  = \new_[42595]_  & \new_[42592]_ ;
  assign \new_[42597]_  = \new_[42596]_  & \new_[42589]_ ;
  assign \new_[42600]_  = ~A235 & ~A234;
  assign \new_[42603]_  = ~A268 & ~A267;
  assign \new_[42604]_  = \new_[42603]_  & \new_[42600]_ ;
  assign \new_[42607]_  = ~A300 & ~A269;
  assign \new_[42610]_  = ~A302 & ~A301;
  assign \new_[42611]_  = \new_[42610]_  & \new_[42607]_ ;
  assign \new_[42612]_  = \new_[42611]_  & \new_[42604]_ ;
  assign \new_[42616]_  = A167 & ~A168;
  assign \new_[42617]_  = ~A169 & \new_[42616]_ ;
  assign \new_[42620]_  = A202 & A166;
  assign \new_[42623]_  = A233 & A232;
  assign \new_[42624]_  = \new_[42623]_  & \new_[42620]_ ;
  assign \new_[42625]_  = \new_[42624]_  & \new_[42617]_ ;
  assign \new_[42628]_  = ~A235 & ~A234;
  assign \new_[42631]_  = ~A268 & ~A267;
  assign \new_[42632]_  = \new_[42631]_  & \new_[42628]_ ;
  assign \new_[42635]_  = ~A298 & ~A269;
  assign \new_[42638]_  = ~A301 & ~A299;
  assign \new_[42639]_  = \new_[42638]_  & \new_[42635]_ ;
  assign \new_[42640]_  = \new_[42639]_  & \new_[42632]_ ;
  assign \new_[42644]_  = A167 & ~A168;
  assign \new_[42645]_  = ~A169 & \new_[42644]_ ;
  assign \new_[42648]_  = A202 & A166;
  assign \new_[42651]_  = A233 & A232;
  assign \new_[42652]_  = \new_[42651]_  & \new_[42648]_ ;
  assign \new_[42653]_  = \new_[42652]_  & \new_[42645]_ ;
  assign \new_[42656]_  = ~A235 & ~A234;
  assign \new_[42659]_  = ~A266 & ~A265;
  assign \new_[42660]_  = \new_[42659]_  & \new_[42656]_ ;
  assign \new_[42663]_  = ~A300 & ~A268;
  assign \new_[42666]_  = ~A302 & ~A301;
  assign \new_[42667]_  = \new_[42666]_  & \new_[42663]_ ;
  assign \new_[42668]_  = \new_[42667]_  & \new_[42660]_ ;
  assign \new_[42672]_  = A167 & ~A168;
  assign \new_[42673]_  = ~A169 & \new_[42672]_ ;
  assign \new_[42676]_  = A202 & A166;
  assign \new_[42679]_  = A233 & A232;
  assign \new_[42680]_  = \new_[42679]_  & \new_[42676]_ ;
  assign \new_[42681]_  = \new_[42680]_  & \new_[42673]_ ;
  assign \new_[42684]_  = ~A235 & ~A234;
  assign \new_[42687]_  = ~A266 & ~A265;
  assign \new_[42688]_  = \new_[42687]_  & \new_[42684]_ ;
  assign \new_[42691]_  = ~A298 & ~A268;
  assign \new_[42694]_  = ~A301 & ~A299;
  assign \new_[42695]_  = \new_[42694]_  & \new_[42691]_ ;
  assign \new_[42696]_  = \new_[42695]_  & \new_[42688]_ ;
  assign \new_[42700]_  = A167 & ~A168;
  assign \new_[42701]_  = ~A169 & \new_[42700]_ ;
  assign \new_[42704]_  = A202 & A166;
  assign \new_[42707]_  = ~A233 & ~A232;
  assign \new_[42708]_  = \new_[42707]_  & \new_[42704]_ ;
  assign \new_[42709]_  = \new_[42708]_  & \new_[42701]_ ;
  assign \new_[42712]_  = ~A267 & ~A235;
  assign \new_[42715]_  = ~A269 & ~A268;
  assign \new_[42716]_  = \new_[42715]_  & \new_[42712]_ ;
  assign \new_[42719]_  = A299 & A298;
  assign \new_[42722]_  = ~A301 & ~A300;
  assign \new_[42723]_  = \new_[42722]_  & \new_[42719]_ ;
  assign \new_[42724]_  = \new_[42723]_  & \new_[42716]_ ;
  assign \new_[42728]_  = A167 & ~A168;
  assign \new_[42729]_  = ~A169 & \new_[42728]_ ;
  assign \new_[42732]_  = A202 & A166;
  assign \new_[42735]_  = ~A233 & ~A232;
  assign \new_[42736]_  = \new_[42735]_  & \new_[42732]_ ;
  assign \new_[42737]_  = \new_[42736]_  & \new_[42729]_ ;
  assign \new_[42740]_  = A265 & ~A235;
  assign \new_[42743]_  = ~A267 & A266;
  assign \new_[42744]_  = \new_[42743]_  & \new_[42740]_ ;
  assign \new_[42747]_  = ~A300 & ~A268;
  assign \new_[42750]_  = ~A302 & ~A301;
  assign \new_[42751]_  = \new_[42750]_  & \new_[42747]_ ;
  assign \new_[42752]_  = \new_[42751]_  & \new_[42744]_ ;
  assign \new_[42756]_  = A167 & ~A168;
  assign \new_[42757]_  = ~A169 & \new_[42756]_ ;
  assign \new_[42760]_  = A202 & A166;
  assign \new_[42763]_  = ~A233 & ~A232;
  assign \new_[42764]_  = \new_[42763]_  & \new_[42760]_ ;
  assign \new_[42765]_  = \new_[42764]_  & \new_[42757]_ ;
  assign \new_[42768]_  = A265 & ~A235;
  assign \new_[42771]_  = ~A267 & A266;
  assign \new_[42772]_  = \new_[42771]_  & \new_[42768]_ ;
  assign \new_[42775]_  = ~A298 & ~A268;
  assign \new_[42778]_  = ~A301 & ~A299;
  assign \new_[42779]_  = \new_[42778]_  & \new_[42775]_ ;
  assign \new_[42780]_  = \new_[42779]_  & \new_[42772]_ ;
  assign \new_[42784]_  = A167 & ~A168;
  assign \new_[42785]_  = ~A169 & \new_[42784]_ ;
  assign \new_[42788]_  = A202 & A166;
  assign \new_[42791]_  = ~A233 & ~A232;
  assign \new_[42792]_  = \new_[42791]_  & \new_[42788]_ ;
  assign \new_[42793]_  = \new_[42792]_  & \new_[42785]_ ;
  assign \new_[42796]_  = ~A265 & ~A235;
  assign \new_[42799]_  = ~A268 & ~A266;
  assign \new_[42800]_  = \new_[42799]_  & \new_[42796]_ ;
  assign \new_[42803]_  = A299 & A298;
  assign \new_[42806]_  = ~A301 & ~A300;
  assign \new_[42807]_  = \new_[42806]_  & \new_[42803]_ ;
  assign \new_[42808]_  = \new_[42807]_  & \new_[42800]_ ;
  assign \new_[42812]_  = A167 & ~A168;
  assign \new_[42813]_  = ~A169 & \new_[42812]_ ;
  assign \new_[42816]_  = A199 & A166;
  assign \new_[42819]_  = ~A234 & A201;
  assign \new_[42820]_  = \new_[42819]_  & \new_[42816]_ ;
  assign \new_[42821]_  = \new_[42820]_  & \new_[42813]_ ;
  assign \new_[42824]_  = ~A236 & ~A235;
  assign \new_[42827]_  = ~A268 & ~A267;
  assign \new_[42828]_  = \new_[42827]_  & \new_[42824]_ ;
  assign \new_[42831]_  = ~A300 & ~A269;
  assign \new_[42834]_  = ~A302 & ~A301;
  assign \new_[42835]_  = \new_[42834]_  & \new_[42831]_ ;
  assign \new_[42836]_  = \new_[42835]_  & \new_[42828]_ ;
  assign \new_[42840]_  = A167 & ~A168;
  assign \new_[42841]_  = ~A169 & \new_[42840]_ ;
  assign \new_[42844]_  = A199 & A166;
  assign \new_[42847]_  = ~A234 & A201;
  assign \new_[42848]_  = \new_[42847]_  & \new_[42844]_ ;
  assign \new_[42849]_  = \new_[42848]_  & \new_[42841]_ ;
  assign \new_[42852]_  = ~A236 & ~A235;
  assign \new_[42855]_  = ~A268 & ~A267;
  assign \new_[42856]_  = \new_[42855]_  & \new_[42852]_ ;
  assign \new_[42859]_  = ~A298 & ~A269;
  assign \new_[42862]_  = ~A301 & ~A299;
  assign \new_[42863]_  = \new_[42862]_  & \new_[42859]_ ;
  assign \new_[42864]_  = \new_[42863]_  & \new_[42856]_ ;
  assign \new_[42868]_  = A167 & ~A168;
  assign \new_[42869]_  = ~A169 & \new_[42868]_ ;
  assign \new_[42872]_  = A199 & A166;
  assign \new_[42875]_  = ~A234 & A201;
  assign \new_[42876]_  = \new_[42875]_  & \new_[42872]_ ;
  assign \new_[42877]_  = \new_[42876]_  & \new_[42869]_ ;
  assign \new_[42880]_  = ~A236 & ~A235;
  assign \new_[42883]_  = ~A266 & ~A265;
  assign \new_[42884]_  = \new_[42883]_  & \new_[42880]_ ;
  assign \new_[42887]_  = ~A300 & ~A268;
  assign \new_[42890]_  = ~A302 & ~A301;
  assign \new_[42891]_  = \new_[42890]_  & \new_[42887]_ ;
  assign \new_[42892]_  = \new_[42891]_  & \new_[42884]_ ;
  assign \new_[42896]_  = A167 & ~A168;
  assign \new_[42897]_  = ~A169 & \new_[42896]_ ;
  assign \new_[42900]_  = A199 & A166;
  assign \new_[42903]_  = ~A234 & A201;
  assign \new_[42904]_  = \new_[42903]_  & \new_[42900]_ ;
  assign \new_[42905]_  = \new_[42904]_  & \new_[42897]_ ;
  assign \new_[42908]_  = ~A236 & ~A235;
  assign \new_[42911]_  = ~A266 & ~A265;
  assign \new_[42912]_  = \new_[42911]_  & \new_[42908]_ ;
  assign \new_[42915]_  = ~A298 & ~A268;
  assign \new_[42918]_  = ~A301 & ~A299;
  assign \new_[42919]_  = \new_[42918]_  & \new_[42915]_ ;
  assign \new_[42920]_  = \new_[42919]_  & \new_[42912]_ ;
  assign \new_[42924]_  = A167 & ~A168;
  assign \new_[42925]_  = ~A169 & \new_[42924]_ ;
  assign \new_[42928]_  = A199 & A166;
  assign \new_[42931]_  = ~A232 & A201;
  assign \new_[42932]_  = \new_[42931]_  & \new_[42928]_ ;
  assign \new_[42933]_  = \new_[42932]_  & \new_[42925]_ ;
  assign \new_[42936]_  = ~A235 & ~A233;
  assign \new_[42939]_  = ~A268 & ~A267;
  assign \new_[42940]_  = \new_[42939]_  & \new_[42936]_ ;
  assign \new_[42943]_  = ~A300 & ~A269;
  assign \new_[42946]_  = ~A302 & ~A301;
  assign \new_[42947]_  = \new_[42946]_  & \new_[42943]_ ;
  assign \new_[42948]_  = \new_[42947]_  & \new_[42940]_ ;
  assign \new_[42952]_  = A167 & ~A168;
  assign \new_[42953]_  = ~A169 & \new_[42952]_ ;
  assign \new_[42956]_  = A199 & A166;
  assign \new_[42959]_  = ~A232 & A201;
  assign \new_[42960]_  = \new_[42959]_  & \new_[42956]_ ;
  assign \new_[42961]_  = \new_[42960]_  & \new_[42953]_ ;
  assign \new_[42964]_  = ~A235 & ~A233;
  assign \new_[42967]_  = ~A268 & ~A267;
  assign \new_[42968]_  = \new_[42967]_  & \new_[42964]_ ;
  assign \new_[42971]_  = ~A298 & ~A269;
  assign \new_[42974]_  = ~A301 & ~A299;
  assign \new_[42975]_  = \new_[42974]_  & \new_[42971]_ ;
  assign \new_[42976]_  = \new_[42975]_  & \new_[42968]_ ;
  assign \new_[42980]_  = A167 & ~A168;
  assign \new_[42981]_  = ~A169 & \new_[42980]_ ;
  assign \new_[42984]_  = A199 & A166;
  assign \new_[42987]_  = ~A232 & A201;
  assign \new_[42988]_  = \new_[42987]_  & \new_[42984]_ ;
  assign \new_[42989]_  = \new_[42988]_  & \new_[42981]_ ;
  assign \new_[42992]_  = ~A235 & ~A233;
  assign \new_[42995]_  = ~A266 & ~A265;
  assign \new_[42996]_  = \new_[42995]_  & \new_[42992]_ ;
  assign \new_[42999]_  = ~A300 & ~A268;
  assign \new_[43002]_  = ~A302 & ~A301;
  assign \new_[43003]_  = \new_[43002]_  & \new_[42999]_ ;
  assign \new_[43004]_  = \new_[43003]_  & \new_[42996]_ ;
  assign \new_[43008]_  = A167 & ~A168;
  assign \new_[43009]_  = ~A169 & \new_[43008]_ ;
  assign \new_[43012]_  = A199 & A166;
  assign \new_[43015]_  = ~A232 & A201;
  assign \new_[43016]_  = \new_[43015]_  & \new_[43012]_ ;
  assign \new_[43017]_  = \new_[43016]_  & \new_[43009]_ ;
  assign \new_[43020]_  = ~A235 & ~A233;
  assign \new_[43023]_  = ~A266 & ~A265;
  assign \new_[43024]_  = \new_[43023]_  & \new_[43020]_ ;
  assign \new_[43027]_  = ~A298 & ~A268;
  assign \new_[43030]_  = ~A301 & ~A299;
  assign \new_[43031]_  = \new_[43030]_  & \new_[43027]_ ;
  assign \new_[43032]_  = \new_[43031]_  & \new_[43024]_ ;
  assign \new_[43036]_  = A167 & ~A168;
  assign \new_[43037]_  = ~A169 & \new_[43036]_ ;
  assign \new_[43040]_  = A200 & A166;
  assign \new_[43043]_  = ~A234 & A201;
  assign \new_[43044]_  = \new_[43043]_  & \new_[43040]_ ;
  assign \new_[43045]_  = \new_[43044]_  & \new_[43037]_ ;
  assign \new_[43048]_  = ~A236 & ~A235;
  assign \new_[43051]_  = ~A268 & ~A267;
  assign \new_[43052]_  = \new_[43051]_  & \new_[43048]_ ;
  assign \new_[43055]_  = ~A300 & ~A269;
  assign \new_[43058]_  = ~A302 & ~A301;
  assign \new_[43059]_  = \new_[43058]_  & \new_[43055]_ ;
  assign \new_[43060]_  = \new_[43059]_  & \new_[43052]_ ;
  assign \new_[43064]_  = A167 & ~A168;
  assign \new_[43065]_  = ~A169 & \new_[43064]_ ;
  assign \new_[43068]_  = A200 & A166;
  assign \new_[43071]_  = ~A234 & A201;
  assign \new_[43072]_  = \new_[43071]_  & \new_[43068]_ ;
  assign \new_[43073]_  = \new_[43072]_  & \new_[43065]_ ;
  assign \new_[43076]_  = ~A236 & ~A235;
  assign \new_[43079]_  = ~A268 & ~A267;
  assign \new_[43080]_  = \new_[43079]_  & \new_[43076]_ ;
  assign \new_[43083]_  = ~A298 & ~A269;
  assign \new_[43086]_  = ~A301 & ~A299;
  assign \new_[43087]_  = \new_[43086]_  & \new_[43083]_ ;
  assign \new_[43088]_  = \new_[43087]_  & \new_[43080]_ ;
  assign \new_[43092]_  = A167 & ~A168;
  assign \new_[43093]_  = ~A169 & \new_[43092]_ ;
  assign \new_[43096]_  = A200 & A166;
  assign \new_[43099]_  = ~A234 & A201;
  assign \new_[43100]_  = \new_[43099]_  & \new_[43096]_ ;
  assign \new_[43101]_  = \new_[43100]_  & \new_[43093]_ ;
  assign \new_[43104]_  = ~A236 & ~A235;
  assign \new_[43107]_  = ~A266 & ~A265;
  assign \new_[43108]_  = \new_[43107]_  & \new_[43104]_ ;
  assign \new_[43111]_  = ~A300 & ~A268;
  assign \new_[43114]_  = ~A302 & ~A301;
  assign \new_[43115]_  = \new_[43114]_  & \new_[43111]_ ;
  assign \new_[43116]_  = \new_[43115]_  & \new_[43108]_ ;
  assign \new_[43120]_  = A167 & ~A168;
  assign \new_[43121]_  = ~A169 & \new_[43120]_ ;
  assign \new_[43124]_  = A200 & A166;
  assign \new_[43127]_  = ~A234 & A201;
  assign \new_[43128]_  = \new_[43127]_  & \new_[43124]_ ;
  assign \new_[43129]_  = \new_[43128]_  & \new_[43121]_ ;
  assign \new_[43132]_  = ~A236 & ~A235;
  assign \new_[43135]_  = ~A266 & ~A265;
  assign \new_[43136]_  = \new_[43135]_  & \new_[43132]_ ;
  assign \new_[43139]_  = ~A298 & ~A268;
  assign \new_[43142]_  = ~A301 & ~A299;
  assign \new_[43143]_  = \new_[43142]_  & \new_[43139]_ ;
  assign \new_[43144]_  = \new_[43143]_  & \new_[43136]_ ;
  assign \new_[43148]_  = A167 & ~A168;
  assign \new_[43149]_  = ~A169 & \new_[43148]_ ;
  assign \new_[43152]_  = A200 & A166;
  assign \new_[43155]_  = ~A232 & A201;
  assign \new_[43156]_  = \new_[43155]_  & \new_[43152]_ ;
  assign \new_[43157]_  = \new_[43156]_  & \new_[43149]_ ;
  assign \new_[43160]_  = ~A235 & ~A233;
  assign \new_[43163]_  = ~A268 & ~A267;
  assign \new_[43164]_  = \new_[43163]_  & \new_[43160]_ ;
  assign \new_[43167]_  = ~A300 & ~A269;
  assign \new_[43170]_  = ~A302 & ~A301;
  assign \new_[43171]_  = \new_[43170]_  & \new_[43167]_ ;
  assign \new_[43172]_  = \new_[43171]_  & \new_[43164]_ ;
  assign \new_[43176]_  = A167 & ~A168;
  assign \new_[43177]_  = ~A169 & \new_[43176]_ ;
  assign \new_[43180]_  = A200 & A166;
  assign \new_[43183]_  = ~A232 & A201;
  assign \new_[43184]_  = \new_[43183]_  & \new_[43180]_ ;
  assign \new_[43185]_  = \new_[43184]_  & \new_[43177]_ ;
  assign \new_[43188]_  = ~A235 & ~A233;
  assign \new_[43191]_  = ~A268 & ~A267;
  assign \new_[43192]_  = \new_[43191]_  & \new_[43188]_ ;
  assign \new_[43195]_  = ~A298 & ~A269;
  assign \new_[43198]_  = ~A301 & ~A299;
  assign \new_[43199]_  = \new_[43198]_  & \new_[43195]_ ;
  assign \new_[43200]_  = \new_[43199]_  & \new_[43192]_ ;
  assign \new_[43204]_  = A167 & ~A168;
  assign \new_[43205]_  = ~A169 & \new_[43204]_ ;
  assign \new_[43208]_  = A200 & A166;
  assign \new_[43211]_  = ~A232 & A201;
  assign \new_[43212]_  = \new_[43211]_  & \new_[43208]_ ;
  assign \new_[43213]_  = \new_[43212]_  & \new_[43205]_ ;
  assign \new_[43216]_  = ~A235 & ~A233;
  assign \new_[43219]_  = ~A266 & ~A265;
  assign \new_[43220]_  = \new_[43219]_  & \new_[43216]_ ;
  assign \new_[43223]_  = ~A300 & ~A268;
  assign \new_[43226]_  = ~A302 & ~A301;
  assign \new_[43227]_  = \new_[43226]_  & \new_[43223]_ ;
  assign \new_[43228]_  = \new_[43227]_  & \new_[43220]_ ;
  assign \new_[43232]_  = A167 & ~A168;
  assign \new_[43233]_  = ~A169 & \new_[43232]_ ;
  assign \new_[43236]_  = A200 & A166;
  assign \new_[43239]_  = ~A232 & A201;
  assign \new_[43240]_  = \new_[43239]_  & \new_[43236]_ ;
  assign \new_[43241]_  = \new_[43240]_  & \new_[43233]_ ;
  assign \new_[43244]_  = ~A235 & ~A233;
  assign \new_[43247]_  = ~A266 & ~A265;
  assign \new_[43248]_  = \new_[43247]_  & \new_[43244]_ ;
  assign \new_[43251]_  = ~A298 & ~A268;
  assign \new_[43254]_  = ~A301 & ~A299;
  assign \new_[43255]_  = \new_[43254]_  & \new_[43251]_ ;
  assign \new_[43256]_  = \new_[43255]_  & \new_[43248]_ ;
  assign \new_[43260]_  = ~A168 & ~A169;
  assign \new_[43261]_  = ~A170 & \new_[43260]_ ;
  assign \new_[43264]_  = ~A234 & A202;
  assign \new_[43267]_  = ~A236 & ~A235;
  assign \new_[43268]_  = \new_[43267]_  & \new_[43264]_ ;
  assign \new_[43269]_  = \new_[43268]_  & \new_[43261]_ ;
  assign \new_[43272]_  = A266 & A265;
  assign \new_[43275]_  = ~A268 & ~A267;
  assign \new_[43276]_  = \new_[43275]_  & \new_[43272]_ ;
  assign \new_[43279]_  = A299 & A298;
  assign \new_[43282]_  = ~A301 & ~A300;
  assign \new_[43283]_  = \new_[43282]_  & \new_[43279]_ ;
  assign \new_[43284]_  = \new_[43283]_  & \new_[43276]_ ;
  assign \new_[43288]_  = ~A168 & ~A169;
  assign \new_[43289]_  = ~A170 & \new_[43288]_ ;
  assign \new_[43292]_  = A232 & A202;
  assign \new_[43295]_  = ~A234 & A233;
  assign \new_[43296]_  = \new_[43295]_  & \new_[43292]_ ;
  assign \new_[43297]_  = \new_[43296]_  & \new_[43289]_ ;
  assign \new_[43300]_  = ~A267 & ~A235;
  assign \new_[43303]_  = ~A269 & ~A268;
  assign \new_[43304]_  = \new_[43303]_  & \new_[43300]_ ;
  assign \new_[43307]_  = A299 & A298;
  assign \new_[43310]_  = ~A301 & ~A300;
  assign \new_[43311]_  = \new_[43310]_  & \new_[43307]_ ;
  assign \new_[43312]_  = \new_[43311]_  & \new_[43304]_ ;
  assign \new_[43316]_  = ~A168 & ~A169;
  assign \new_[43317]_  = ~A170 & \new_[43316]_ ;
  assign \new_[43320]_  = A232 & A202;
  assign \new_[43323]_  = ~A234 & A233;
  assign \new_[43324]_  = \new_[43323]_  & \new_[43320]_ ;
  assign \new_[43325]_  = \new_[43324]_  & \new_[43317]_ ;
  assign \new_[43328]_  = A265 & ~A235;
  assign \new_[43331]_  = ~A267 & A266;
  assign \new_[43332]_  = \new_[43331]_  & \new_[43328]_ ;
  assign \new_[43335]_  = ~A300 & ~A268;
  assign \new_[43338]_  = ~A302 & ~A301;
  assign \new_[43339]_  = \new_[43338]_  & \new_[43335]_ ;
  assign \new_[43340]_  = \new_[43339]_  & \new_[43332]_ ;
  assign \new_[43344]_  = ~A168 & ~A169;
  assign \new_[43345]_  = ~A170 & \new_[43344]_ ;
  assign \new_[43348]_  = A232 & A202;
  assign \new_[43351]_  = ~A234 & A233;
  assign \new_[43352]_  = \new_[43351]_  & \new_[43348]_ ;
  assign \new_[43353]_  = \new_[43352]_  & \new_[43345]_ ;
  assign \new_[43356]_  = A265 & ~A235;
  assign \new_[43359]_  = ~A267 & A266;
  assign \new_[43360]_  = \new_[43359]_  & \new_[43356]_ ;
  assign \new_[43363]_  = ~A298 & ~A268;
  assign \new_[43366]_  = ~A301 & ~A299;
  assign \new_[43367]_  = \new_[43366]_  & \new_[43363]_ ;
  assign \new_[43368]_  = \new_[43367]_  & \new_[43360]_ ;
  assign \new_[43372]_  = ~A168 & ~A169;
  assign \new_[43373]_  = ~A170 & \new_[43372]_ ;
  assign \new_[43376]_  = A232 & A202;
  assign \new_[43379]_  = ~A234 & A233;
  assign \new_[43380]_  = \new_[43379]_  & \new_[43376]_ ;
  assign \new_[43381]_  = \new_[43380]_  & \new_[43373]_ ;
  assign \new_[43384]_  = ~A265 & ~A235;
  assign \new_[43387]_  = ~A268 & ~A266;
  assign \new_[43388]_  = \new_[43387]_  & \new_[43384]_ ;
  assign \new_[43391]_  = A299 & A298;
  assign \new_[43394]_  = ~A301 & ~A300;
  assign \new_[43395]_  = \new_[43394]_  & \new_[43391]_ ;
  assign \new_[43396]_  = \new_[43395]_  & \new_[43388]_ ;
  assign \new_[43400]_  = ~A168 & ~A169;
  assign \new_[43401]_  = ~A170 & \new_[43400]_ ;
  assign \new_[43404]_  = ~A232 & A202;
  assign \new_[43407]_  = ~A235 & ~A233;
  assign \new_[43408]_  = \new_[43407]_  & \new_[43404]_ ;
  assign \new_[43409]_  = \new_[43408]_  & \new_[43401]_ ;
  assign \new_[43412]_  = A266 & A265;
  assign \new_[43415]_  = ~A268 & ~A267;
  assign \new_[43416]_  = \new_[43415]_  & \new_[43412]_ ;
  assign \new_[43419]_  = A299 & A298;
  assign \new_[43422]_  = ~A301 & ~A300;
  assign \new_[43423]_  = \new_[43422]_  & \new_[43419]_ ;
  assign \new_[43424]_  = \new_[43423]_  & \new_[43416]_ ;
  assign \new_[43428]_  = ~A168 & ~A169;
  assign \new_[43429]_  = ~A170 & \new_[43428]_ ;
  assign \new_[43432]_  = A201 & A199;
  assign \new_[43435]_  = ~A235 & ~A234;
  assign \new_[43436]_  = \new_[43435]_  & \new_[43432]_ ;
  assign \new_[43437]_  = \new_[43436]_  & \new_[43429]_ ;
  assign \new_[43440]_  = ~A267 & ~A236;
  assign \new_[43443]_  = ~A269 & ~A268;
  assign \new_[43444]_  = \new_[43443]_  & \new_[43440]_ ;
  assign \new_[43447]_  = A299 & A298;
  assign \new_[43450]_  = ~A301 & ~A300;
  assign \new_[43451]_  = \new_[43450]_  & \new_[43447]_ ;
  assign \new_[43452]_  = \new_[43451]_  & \new_[43444]_ ;
  assign \new_[43456]_  = ~A168 & ~A169;
  assign \new_[43457]_  = ~A170 & \new_[43456]_ ;
  assign \new_[43460]_  = A201 & A199;
  assign \new_[43463]_  = ~A235 & ~A234;
  assign \new_[43464]_  = \new_[43463]_  & \new_[43460]_ ;
  assign \new_[43465]_  = \new_[43464]_  & \new_[43457]_ ;
  assign \new_[43468]_  = A265 & ~A236;
  assign \new_[43471]_  = ~A267 & A266;
  assign \new_[43472]_  = \new_[43471]_  & \new_[43468]_ ;
  assign \new_[43475]_  = ~A300 & ~A268;
  assign \new_[43478]_  = ~A302 & ~A301;
  assign \new_[43479]_  = \new_[43478]_  & \new_[43475]_ ;
  assign \new_[43480]_  = \new_[43479]_  & \new_[43472]_ ;
  assign \new_[43484]_  = ~A168 & ~A169;
  assign \new_[43485]_  = ~A170 & \new_[43484]_ ;
  assign \new_[43488]_  = A201 & A199;
  assign \new_[43491]_  = ~A235 & ~A234;
  assign \new_[43492]_  = \new_[43491]_  & \new_[43488]_ ;
  assign \new_[43493]_  = \new_[43492]_  & \new_[43485]_ ;
  assign \new_[43496]_  = A265 & ~A236;
  assign \new_[43499]_  = ~A267 & A266;
  assign \new_[43500]_  = \new_[43499]_  & \new_[43496]_ ;
  assign \new_[43503]_  = ~A298 & ~A268;
  assign \new_[43506]_  = ~A301 & ~A299;
  assign \new_[43507]_  = \new_[43506]_  & \new_[43503]_ ;
  assign \new_[43508]_  = \new_[43507]_  & \new_[43500]_ ;
  assign \new_[43512]_  = ~A168 & ~A169;
  assign \new_[43513]_  = ~A170 & \new_[43512]_ ;
  assign \new_[43516]_  = A201 & A199;
  assign \new_[43519]_  = ~A235 & ~A234;
  assign \new_[43520]_  = \new_[43519]_  & \new_[43516]_ ;
  assign \new_[43521]_  = \new_[43520]_  & \new_[43513]_ ;
  assign \new_[43524]_  = ~A265 & ~A236;
  assign \new_[43527]_  = ~A268 & ~A266;
  assign \new_[43528]_  = \new_[43527]_  & \new_[43524]_ ;
  assign \new_[43531]_  = A299 & A298;
  assign \new_[43534]_  = ~A301 & ~A300;
  assign \new_[43535]_  = \new_[43534]_  & \new_[43531]_ ;
  assign \new_[43536]_  = \new_[43535]_  & \new_[43528]_ ;
  assign \new_[43540]_  = ~A168 & ~A169;
  assign \new_[43541]_  = ~A170 & \new_[43540]_ ;
  assign \new_[43544]_  = A201 & A199;
  assign \new_[43547]_  = A233 & A232;
  assign \new_[43548]_  = \new_[43547]_  & \new_[43544]_ ;
  assign \new_[43549]_  = \new_[43548]_  & \new_[43541]_ ;
  assign \new_[43552]_  = ~A235 & ~A234;
  assign \new_[43555]_  = ~A268 & ~A267;
  assign \new_[43556]_  = \new_[43555]_  & \new_[43552]_ ;
  assign \new_[43559]_  = ~A300 & ~A269;
  assign \new_[43562]_  = ~A302 & ~A301;
  assign \new_[43563]_  = \new_[43562]_  & \new_[43559]_ ;
  assign \new_[43564]_  = \new_[43563]_  & \new_[43556]_ ;
  assign \new_[43568]_  = ~A168 & ~A169;
  assign \new_[43569]_  = ~A170 & \new_[43568]_ ;
  assign \new_[43572]_  = A201 & A199;
  assign \new_[43575]_  = A233 & A232;
  assign \new_[43576]_  = \new_[43575]_  & \new_[43572]_ ;
  assign \new_[43577]_  = \new_[43576]_  & \new_[43569]_ ;
  assign \new_[43580]_  = ~A235 & ~A234;
  assign \new_[43583]_  = ~A268 & ~A267;
  assign \new_[43584]_  = \new_[43583]_  & \new_[43580]_ ;
  assign \new_[43587]_  = ~A298 & ~A269;
  assign \new_[43590]_  = ~A301 & ~A299;
  assign \new_[43591]_  = \new_[43590]_  & \new_[43587]_ ;
  assign \new_[43592]_  = \new_[43591]_  & \new_[43584]_ ;
  assign \new_[43596]_  = ~A168 & ~A169;
  assign \new_[43597]_  = ~A170 & \new_[43596]_ ;
  assign \new_[43600]_  = A201 & A199;
  assign \new_[43603]_  = A233 & A232;
  assign \new_[43604]_  = \new_[43603]_  & \new_[43600]_ ;
  assign \new_[43605]_  = \new_[43604]_  & \new_[43597]_ ;
  assign \new_[43608]_  = ~A235 & ~A234;
  assign \new_[43611]_  = ~A266 & ~A265;
  assign \new_[43612]_  = \new_[43611]_  & \new_[43608]_ ;
  assign \new_[43615]_  = ~A300 & ~A268;
  assign \new_[43618]_  = ~A302 & ~A301;
  assign \new_[43619]_  = \new_[43618]_  & \new_[43615]_ ;
  assign \new_[43620]_  = \new_[43619]_  & \new_[43612]_ ;
  assign \new_[43624]_  = ~A168 & ~A169;
  assign \new_[43625]_  = ~A170 & \new_[43624]_ ;
  assign \new_[43628]_  = A201 & A199;
  assign \new_[43631]_  = A233 & A232;
  assign \new_[43632]_  = \new_[43631]_  & \new_[43628]_ ;
  assign \new_[43633]_  = \new_[43632]_  & \new_[43625]_ ;
  assign \new_[43636]_  = ~A235 & ~A234;
  assign \new_[43639]_  = ~A266 & ~A265;
  assign \new_[43640]_  = \new_[43639]_  & \new_[43636]_ ;
  assign \new_[43643]_  = ~A298 & ~A268;
  assign \new_[43646]_  = ~A301 & ~A299;
  assign \new_[43647]_  = \new_[43646]_  & \new_[43643]_ ;
  assign \new_[43648]_  = \new_[43647]_  & \new_[43640]_ ;
  assign \new_[43652]_  = ~A168 & ~A169;
  assign \new_[43653]_  = ~A170 & \new_[43652]_ ;
  assign \new_[43656]_  = A201 & A199;
  assign \new_[43659]_  = ~A233 & ~A232;
  assign \new_[43660]_  = \new_[43659]_  & \new_[43656]_ ;
  assign \new_[43661]_  = \new_[43660]_  & \new_[43653]_ ;
  assign \new_[43664]_  = ~A267 & ~A235;
  assign \new_[43667]_  = ~A269 & ~A268;
  assign \new_[43668]_  = \new_[43667]_  & \new_[43664]_ ;
  assign \new_[43671]_  = A299 & A298;
  assign \new_[43674]_  = ~A301 & ~A300;
  assign \new_[43675]_  = \new_[43674]_  & \new_[43671]_ ;
  assign \new_[43676]_  = \new_[43675]_  & \new_[43668]_ ;
  assign \new_[43680]_  = ~A168 & ~A169;
  assign \new_[43681]_  = ~A170 & \new_[43680]_ ;
  assign \new_[43684]_  = A201 & A199;
  assign \new_[43687]_  = ~A233 & ~A232;
  assign \new_[43688]_  = \new_[43687]_  & \new_[43684]_ ;
  assign \new_[43689]_  = \new_[43688]_  & \new_[43681]_ ;
  assign \new_[43692]_  = A265 & ~A235;
  assign \new_[43695]_  = ~A267 & A266;
  assign \new_[43696]_  = \new_[43695]_  & \new_[43692]_ ;
  assign \new_[43699]_  = ~A300 & ~A268;
  assign \new_[43702]_  = ~A302 & ~A301;
  assign \new_[43703]_  = \new_[43702]_  & \new_[43699]_ ;
  assign \new_[43704]_  = \new_[43703]_  & \new_[43696]_ ;
  assign \new_[43708]_  = ~A168 & ~A169;
  assign \new_[43709]_  = ~A170 & \new_[43708]_ ;
  assign \new_[43712]_  = A201 & A199;
  assign \new_[43715]_  = ~A233 & ~A232;
  assign \new_[43716]_  = \new_[43715]_  & \new_[43712]_ ;
  assign \new_[43717]_  = \new_[43716]_  & \new_[43709]_ ;
  assign \new_[43720]_  = A265 & ~A235;
  assign \new_[43723]_  = ~A267 & A266;
  assign \new_[43724]_  = \new_[43723]_  & \new_[43720]_ ;
  assign \new_[43727]_  = ~A298 & ~A268;
  assign \new_[43730]_  = ~A301 & ~A299;
  assign \new_[43731]_  = \new_[43730]_  & \new_[43727]_ ;
  assign \new_[43732]_  = \new_[43731]_  & \new_[43724]_ ;
  assign \new_[43736]_  = ~A168 & ~A169;
  assign \new_[43737]_  = ~A170 & \new_[43736]_ ;
  assign \new_[43740]_  = A201 & A199;
  assign \new_[43743]_  = ~A233 & ~A232;
  assign \new_[43744]_  = \new_[43743]_  & \new_[43740]_ ;
  assign \new_[43745]_  = \new_[43744]_  & \new_[43737]_ ;
  assign \new_[43748]_  = ~A265 & ~A235;
  assign \new_[43751]_  = ~A268 & ~A266;
  assign \new_[43752]_  = \new_[43751]_  & \new_[43748]_ ;
  assign \new_[43755]_  = A299 & A298;
  assign \new_[43758]_  = ~A301 & ~A300;
  assign \new_[43759]_  = \new_[43758]_  & \new_[43755]_ ;
  assign \new_[43760]_  = \new_[43759]_  & \new_[43752]_ ;
  assign \new_[43764]_  = ~A168 & ~A169;
  assign \new_[43765]_  = ~A170 & \new_[43764]_ ;
  assign \new_[43768]_  = A201 & A200;
  assign \new_[43771]_  = ~A235 & ~A234;
  assign \new_[43772]_  = \new_[43771]_  & \new_[43768]_ ;
  assign \new_[43773]_  = \new_[43772]_  & \new_[43765]_ ;
  assign \new_[43776]_  = ~A267 & ~A236;
  assign \new_[43779]_  = ~A269 & ~A268;
  assign \new_[43780]_  = \new_[43779]_  & \new_[43776]_ ;
  assign \new_[43783]_  = A299 & A298;
  assign \new_[43786]_  = ~A301 & ~A300;
  assign \new_[43787]_  = \new_[43786]_  & \new_[43783]_ ;
  assign \new_[43788]_  = \new_[43787]_  & \new_[43780]_ ;
  assign \new_[43792]_  = ~A168 & ~A169;
  assign \new_[43793]_  = ~A170 & \new_[43792]_ ;
  assign \new_[43796]_  = A201 & A200;
  assign \new_[43799]_  = ~A235 & ~A234;
  assign \new_[43800]_  = \new_[43799]_  & \new_[43796]_ ;
  assign \new_[43801]_  = \new_[43800]_  & \new_[43793]_ ;
  assign \new_[43804]_  = A265 & ~A236;
  assign \new_[43807]_  = ~A267 & A266;
  assign \new_[43808]_  = \new_[43807]_  & \new_[43804]_ ;
  assign \new_[43811]_  = ~A300 & ~A268;
  assign \new_[43814]_  = ~A302 & ~A301;
  assign \new_[43815]_  = \new_[43814]_  & \new_[43811]_ ;
  assign \new_[43816]_  = \new_[43815]_  & \new_[43808]_ ;
  assign \new_[43820]_  = ~A168 & ~A169;
  assign \new_[43821]_  = ~A170 & \new_[43820]_ ;
  assign \new_[43824]_  = A201 & A200;
  assign \new_[43827]_  = ~A235 & ~A234;
  assign \new_[43828]_  = \new_[43827]_  & \new_[43824]_ ;
  assign \new_[43829]_  = \new_[43828]_  & \new_[43821]_ ;
  assign \new_[43832]_  = A265 & ~A236;
  assign \new_[43835]_  = ~A267 & A266;
  assign \new_[43836]_  = \new_[43835]_  & \new_[43832]_ ;
  assign \new_[43839]_  = ~A298 & ~A268;
  assign \new_[43842]_  = ~A301 & ~A299;
  assign \new_[43843]_  = \new_[43842]_  & \new_[43839]_ ;
  assign \new_[43844]_  = \new_[43843]_  & \new_[43836]_ ;
  assign \new_[43848]_  = ~A168 & ~A169;
  assign \new_[43849]_  = ~A170 & \new_[43848]_ ;
  assign \new_[43852]_  = A201 & A200;
  assign \new_[43855]_  = ~A235 & ~A234;
  assign \new_[43856]_  = \new_[43855]_  & \new_[43852]_ ;
  assign \new_[43857]_  = \new_[43856]_  & \new_[43849]_ ;
  assign \new_[43860]_  = ~A265 & ~A236;
  assign \new_[43863]_  = ~A268 & ~A266;
  assign \new_[43864]_  = \new_[43863]_  & \new_[43860]_ ;
  assign \new_[43867]_  = A299 & A298;
  assign \new_[43870]_  = ~A301 & ~A300;
  assign \new_[43871]_  = \new_[43870]_  & \new_[43867]_ ;
  assign \new_[43872]_  = \new_[43871]_  & \new_[43864]_ ;
  assign \new_[43876]_  = ~A168 & ~A169;
  assign \new_[43877]_  = ~A170 & \new_[43876]_ ;
  assign \new_[43880]_  = A201 & A200;
  assign \new_[43883]_  = A233 & A232;
  assign \new_[43884]_  = \new_[43883]_  & \new_[43880]_ ;
  assign \new_[43885]_  = \new_[43884]_  & \new_[43877]_ ;
  assign \new_[43888]_  = ~A235 & ~A234;
  assign \new_[43891]_  = ~A268 & ~A267;
  assign \new_[43892]_  = \new_[43891]_  & \new_[43888]_ ;
  assign \new_[43895]_  = ~A300 & ~A269;
  assign \new_[43898]_  = ~A302 & ~A301;
  assign \new_[43899]_  = \new_[43898]_  & \new_[43895]_ ;
  assign \new_[43900]_  = \new_[43899]_  & \new_[43892]_ ;
  assign \new_[43904]_  = ~A168 & ~A169;
  assign \new_[43905]_  = ~A170 & \new_[43904]_ ;
  assign \new_[43908]_  = A201 & A200;
  assign \new_[43911]_  = A233 & A232;
  assign \new_[43912]_  = \new_[43911]_  & \new_[43908]_ ;
  assign \new_[43913]_  = \new_[43912]_  & \new_[43905]_ ;
  assign \new_[43916]_  = ~A235 & ~A234;
  assign \new_[43919]_  = ~A268 & ~A267;
  assign \new_[43920]_  = \new_[43919]_  & \new_[43916]_ ;
  assign \new_[43923]_  = ~A298 & ~A269;
  assign \new_[43926]_  = ~A301 & ~A299;
  assign \new_[43927]_  = \new_[43926]_  & \new_[43923]_ ;
  assign \new_[43928]_  = \new_[43927]_  & \new_[43920]_ ;
  assign \new_[43932]_  = ~A168 & ~A169;
  assign \new_[43933]_  = ~A170 & \new_[43932]_ ;
  assign \new_[43936]_  = A201 & A200;
  assign \new_[43939]_  = A233 & A232;
  assign \new_[43940]_  = \new_[43939]_  & \new_[43936]_ ;
  assign \new_[43941]_  = \new_[43940]_  & \new_[43933]_ ;
  assign \new_[43944]_  = ~A235 & ~A234;
  assign \new_[43947]_  = ~A266 & ~A265;
  assign \new_[43948]_  = \new_[43947]_  & \new_[43944]_ ;
  assign \new_[43951]_  = ~A300 & ~A268;
  assign \new_[43954]_  = ~A302 & ~A301;
  assign \new_[43955]_  = \new_[43954]_  & \new_[43951]_ ;
  assign \new_[43956]_  = \new_[43955]_  & \new_[43948]_ ;
  assign \new_[43960]_  = ~A168 & ~A169;
  assign \new_[43961]_  = ~A170 & \new_[43960]_ ;
  assign \new_[43964]_  = A201 & A200;
  assign \new_[43967]_  = A233 & A232;
  assign \new_[43968]_  = \new_[43967]_  & \new_[43964]_ ;
  assign \new_[43969]_  = \new_[43968]_  & \new_[43961]_ ;
  assign \new_[43972]_  = ~A235 & ~A234;
  assign \new_[43975]_  = ~A266 & ~A265;
  assign \new_[43976]_  = \new_[43975]_  & \new_[43972]_ ;
  assign \new_[43979]_  = ~A298 & ~A268;
  assign \new_[43982]_  = ~A301 & ~A299;
  assign \new_[43983]_  = \new_[43982]_  & \new_[43979]_ ;
  assign \new_[43984]_  = \new_[43983]_  & \new_[43976]_ ;
  assign \new_[43988]_  = ~A168 & ~A169;
  assign \new_[43989]_  = ~A170 & \new_[43988]_ ;
  assign \new_[43992]_  = A201 & A200;
  assign \new_[43995]_  = ~A233 & ~A232;
  assign \new_[43996]_  = \new_[43995]_  & \new_[43992]_ ;
  assign \new_[43997]_  = \new_[43996]_  & \new_[43989]_ ;
  assign \new_[44000]_  = ~A267 & ~A235;
  assign \new_[44003]_  = ~A269 & ~A268;
  assign \new_[44004]_  = \new_[44003]_  & \new_[44000]_ ;
  assign \new_[44007]_  = A299 & A298;
  assign \new_[44010]_  = ~A301 & ~A300;
  assign \new_[44011]_  = \new_[44010]_  & \new_[44007]_ ;
  assign \new_[44012]_  = \new_[44011]_  & \new_[44004]_ ;
  assign \new_[44016]_  = ~A168 & ~A169;
  assign \new_[44017]_  = ~A170 & \new_[44016]_ ;
  assign \new_[44020]_  = A201 & A200;
  assign \new_[44023]_  = ~A233 & ~A232;
  assign \new_[44024]_  = \new_[44023]_  & \new_[44020]_ ;
  assign \new_[44025]_  = \new_[44024]_  & \new_[44017]_ ;
  assign \new_[44028]_  = A265 & ~A235;
  assign \new_[44031]_  = ~A267 & A266;
  assign \new_[44032]_  = \new_[44031]_  & \new_[44028]_ ;
  assign \new_[44035]_  = ~A300 & ~A268;
  assign \new_[44038]_  = ~A302 & ~A301;
  assign \new_[44039]_  = \new_[44038]_  & \new_[44035]_ ;
  assign \new_[44040]_  = \new_[44039]_  & \new_[44032]_ ;
  assign \new_[44044]_  = ~A168 & ~A169;
  assign \new_[44045]_  = ~A170 & \new_[44044]_ ;
  assign \new_[44048]_  = A201 & A200;
  assign \new_[44051]_  = ~A233 & ~A232;
  assign \new_[44052]_  = \new_[44051]_  & \new_[44048]_ ;
  assign \new_[44053]_  = \new_[44052]_  & \new_[44045]_ ;
  assign \new_[44056]_  = A265 & ~A235;
  assign \new_[44059]_  = ~A267 & A266;
  assign \new_[44060]_  = \new_[44059]_  & \new_[44056]_ ;
  assign \new_[44063]_  = ~A298 & ~A268;
  assign \new_[44066]_  = ~A301 & ~A299;
  assign \new_[44067]_  = \new_[44066]_  & \new_[44063]_ ;
  assign \new_[44068]_  = \new_[44067]_  & \new_[44060]_ ;
  assign \new_[44072]_  = ~A168 & ~A169;
  assign \new_[44073]_  = ~A170 & \new_[44072]_ ;
  assign \new_[44076]_  = A201 & A200;
  assign \new_[44079]_  = ~A233 & ~A232;
  assign \new_[44080]_  = \new_[44079]_  & \new_[44076]_ ;
  assign \new_[44081]_  = \new_[44080]_  & \new_[44073]_ ;
  assign \new_[44084]_  = ~A265 & ~A235;
  assign \new_[44087]_  = ~A268 & ~A266;
  assign \new_[44088]_  = \new_[44087]_  & \new_[44084]_ ;
  assign \new_[44091]_  = A299 & A298;
  assign \new_[44094]_  = ~A301 & ~A300;
  assign \new_[44095]_  = \new_[44094]_  & \new_[44091]_ ;
  assign \new_[44096]_  = \new_[44095]_  & \new_[44088]_ ;
  assign \new_[44100]_  = ~A168 & ~A169;
  assign \new_[44101]_  = ~A170 & \new_[44100]_ ;
  assign \new_[44104]_  = A200 & ~A199;
  assign \new_[44107]_  = ~A234 & A203;
  assign \new_[44108]_  = \new_[44107]_  & \new_[44104]_ ;
  assign \new_[44109]_  = \new_[44108]_  & \new_[44101]_ ;
  assign \new_[44112]_  = ~A236 & ~A235;
  assign \new_[44115]_  = ~A268 & ~A267;
  assign \new_[44116]_  = \new_[44115]_  & \new_[44112]_ ;
  assign \new_[44119]_  = ~A300 & ~A269;
  assign \new_[44122]_  = ~A302 & ~A301;
  assign \new_[44123]_  = \new_[44122]_  & \new_[44119]_ ;
  assign \new_[44124]_  = \new_[44123]_  & \new_[44116]_ ;
  assign \new_[44128]_  = ~A168 & ~A169;
  assign \new_[44129]_  = ~A170 & \new_[44128]_ ;
  assign \new_[44132]_  = A200 & ~A199;
  assign \new_[44135]_  = ~A234 & A203;
  assign \new_[44136]_  = \new_[44135]_  & \new_[44132]_ ;
  assign \new_[44137]_  = \new_[44136]_  & \new_[44129]_ ;
  assign \new_[44140]_  = ~A236 & ~A235;
  assign \new_[44143]_  = ~A268 & ~A267;
  assign \new_[44144]_  = \new_[44143]_  & \new_[44140]_ ;
  assign \new_[44147]_  = ~A298 & ~A269;
  assign \new_[44150]_  = ~A301 & ~A299;
  assign \new_[44151]_  = \new_[44150]_  & \new_[44147]_ ;
  assign \new_[44152]_  = \new_[44151]_  & \new_[44144]_ ;
  assign \new_[44156]_  = ~A168 & ~A169;
  assign \new_[44157]_  = ~A170 & \new_[44156]_ ;
  assign \new_[44160]_  = A200 & ~A199;
  assign \new_[44163]_  = ~A234 & A203;
  assign \new_[44164]_  = \new_[44163]_  & \new_[44160]_ ;
  assign \new_[44165]_  = \new_[44164]_  & \new_[44157]_ ;
  assign \new_[44168]_  = ~A236 & ~A235;
  assign \new_[44171]_  = ~A266 & ~A265;
  assign \new_[44172]_  = \new_[44171]_  & \new_[44168]_ ;
  assign \new_[44175]_  = ~A300 & ~A268;
  assign \new_[44178]_  = ~A302 & ~A301;
  assign \new_[44179]_  = \new_[44178]_  & \new_[44175]_ ;
  assign \new_[44180]_  = \new_[44179]_  & \new_[44172]_ ;
  assign \new_[44184]_  = ~A168 & ~A169;
  assign \new_[44185]_  = ~A170 & \new_[44184]_ ;
  assign \new_[44188]_  = A200 & ~A199;
  assign \new_[44191]_  = ~A234 & A203;
  assign \new_[44192]_  = \new_[44191]_  & \new_[44188]_ ;
  assign \new_[44193]_  = \new_[44192]_  & \new_[44185]_ ;
  assign \new_[44196]_  = ~A236 & ~A235;
  assign \new_[44199]_  = ~A266 & ~A265;
  assign \new_[44200]_  = \new_[44199]_  & \new_[44196]_ ;
  assign \new_[44203]_  = ~A298 & ~A268;
  assign \new_[44206]_  = ~A301 & ~A299;
  assign \new_[44207]_  = \new_[44206]_  & \new_[44203]_ ;
  assign \new_[44208]_  = \new_[44207]_  & \new_[44200]_ ;
  assign \new_[44212]_  = ~A168 & ~A169;
  assign \new_[44213]_  = ~A170 & \new_[44212]_ ;
  assign \new_[44216]_  = A200 & ~A199;
  assign \new_[44219]_  = ~A232 & A203;
  assign \new_[44220]_  = \new_[44219]_  & \new_[44216]_ ;
  assign \new_[44221]_  = \new_[44220]_  & \new_[44213]_ ;
  assign \new_[44224]_  = ~A235 & ~A233;
  assign \new_[44227]_  = ~A268 & ~A267;
  assign \new_[44228]_  = \new_[44227]_  & \new_[44224]_ ;
  assign \new_[44231]_  = ~A300 & ~A269;
  assign \new_[44234]_  = ~A302 & ~A301;
  assign \new_[44235]_  = \new_[44234]_  & \new_[44231]_ ;
  assign \new_[44236]_  = \new_[44235]_  & \new_[44228]_ ;
  assign \new_[44240]_  = ~A168 & ~A169;
  assign \new_[44241]_  = ~A170 & \new_[44240]_ ;
  assign \new_[44244]_  = A200 & ~A199;
  assign \new_[44247]_  = ~A232 & A203;
  assign \new_[44248]_  = \new_[44247]_  & \new_[44244]_ ;
  assign \new_[44249]_  = \new_[44248]_  & \new_[44241]_ ;
  assign \new_[44252]_  = ~A235 & ~A233;
  assign \new_[44255]_  = ~A268 & ~A267;
  assign \new_[44256]_  = \new_[44255]_  & \new_[44252]_ ;
  assign \new_[44259]_  = ~A298 & ~A269;
  assign \new_[44262]_  = ~A301 & ~A299;
  assign \new_[44263]_  = \new_[44262]_  & \new_[44259]_ ;
  assign \new_[44264]_  = \new_[44263]_  & \new_[44256]_ ;
  assign \new_[44268]_  = ~A168 & ~A169;
  assign \new_[44269]_  = ~A170 & \new_[44268]_ ;
  assign \new_[44272]_  = A200 & ~A199;
  assign \new_[44275]_  = ~A232 & A203;
  assign \new_[44276]_  = \new_[44275]_  & \new_[44272]_ ;
  assign \new_[44277]_  = \new_[44276]_  & \new_[44269]_ ;
  assign \new_[44280]_  = ~A235 & ~A233;
  assign \new_[44283]_  = ~A266 & ~A265;
  assign \new_[44284]_  = \new_[44283]_  & \new_[44280]_ ;
  assign \new_[44287]_  = ~A300 & ~A268;
  assign \new_[44290]_  = ~A302 & ~A301;
  assign \new_[44291]_  = \new_[44290]_  & \new_[44287]_ ;
  assign \new_[44292]_  = \new_[44291]_  & \new_[44284]_ ;
  assign \new_[44296]_  = ~A168 & ~A169;
  assign \new_[44297]_  = ~A170 & \new_[44296]_ ;
  assign \new_[44300]_  = A200 & ~A199;
  assign \new_[44303]_  = ~A232 & A203;
  assign \new_[44304]_  = \new_[44303]_  & \new_[44300]_ ;
  assign \new_[44305]_  = \new_[44304]_  & \new_[44297]_ ;
  assign \new_[44308]_  = ~A235 & ~A233;
  assign \new_[44311]_  = ~A266 & ~A265;
  assign \new_[44312]_  = \new_[44311]_  & \new_[44308]_ ;
  assign \new_[44315]_  = ~A298 & ~A268;
  assign \new_[44318]_  = ~A301 & ~A299;
  assign \new_[44319]_  = \new_[44318]_  & \new_[44315]_ ;
  assign \new_[44320]_  = \new_[44319]_  & \new_[44312]_ ;
  assign \new_[44324]_  = ~A168 & ~A169;
  assign \new_[44325]_  = ~A170 & \new_[44324]_ ;
  assign \new_[44328]_  = ~A200 & A199;
  assign \new_[44331]_  = ~A234 & A203;
  assign \new_[44332]_  = \new_[44331]_  & \new_[44328]_ ;
  assign \new_[44333]_  = \new_[44332]_  & \new_[44325]_ ;
  assign \new_[44336]_  = ~A236 & ~A235;
  assign \new_[44339]_  = ~A268 & ~A267;
  assign \new_[44340]_  = \new_[44339]_  & \new_[44336]_ ;
  assign \new_[44343]_  = ~A300 & ~A269;
  assign \new_[44346]_  = ~A302 & ~A301;
  assign \new_[44347]_  = \new_[44346]_  & \new_[44343]_ ;
  assign \new_[44348]_  = \new_[44347]_  & \new_[44340]_ ;
  assign \new_[44352]_  = ~A168 & ~A169;
  assign \new_[44353]_  = ~A170 & \new_[44352]_ ;
  assign \new_[44356]_  = ~A200 & A199;
  assign \new_[44359]_  = ~A234 & A203;
  assign \new_[44360]_  = \new_[44359]_  & \new_[44356]_ ;
  assign \new_[44361]_  = \new_[44360]_  & \new_[44353]_ ;
  assign \new_[44364]_  = ~A236 & ~A235;
  assign \new_[44367]_  = ~A268 & ~A267;
  assign \new_[44368]_  = \new_[44367]_  & \new_[44364]_ ;
  assign \new_[44371]_  = ~A298 & ~A269;
  assign \new_[44374]_  = ~A301 & ~A299;
  assign \new_[44375]_  = \new_[44374]_  & \new_[44371]_ ;
  assign \new_[44376]_  = \new_[44375]_  & \new_[44368]_ ;
  assign \new_[44380]_  = ~A168 & ~A169;
  assign \new_[44381]_  = ~A170 & \new_[44380]_ ;
  assign \new_[44384]_  = ~A200 & A199;
  assign \new_[44387]_  = ~A234 & A203;
  assign \new_[44388]_  = \new_[44387]_  & \new_[44384]_ ;
  assign \new_[44389]_  = \new_[44388]_  & \new_[44381]_ ;
  assign \new_[44392]_  = ~A236 & ~A235;
  assign \new_[44395]_  = ~A266 & ~A265;
  assign \new_[44396]_  = \new_[44395]_  & \new_[44392]_ ;
  assign \new_[44399]_  = ~A300 & ~A268;
  assign \new_[44402]_  = ~A302 & ~A301;
  assign \new_[44403]_  = \new_[44402]_  & \new_[44399]_ ;
  assign \new_[44404]_  = \new_[44403]_  & \new_[44396]_ ;
  assign \new_[44408]_  = ~A168 & ~A169;
  assign \new_[44409]_  = ~A170 & \new_[44408]_ ;
  assign \new_[44412]_  = ~A200 & A199;
  assign \new_[44415]_  = ~A234 & A203;
  assign \new_[44416]_  = \new_[44415]_  & \new_[44412]_ ;
  assign \new_[44417]_  = \new_[44416]_  & \new_[44409]_ ;
  assign \new_[44420]_  = ~A236 & ~A235;
  assign \new_[44423]_  = ~A266 & ~A265;
  assign \new_[44424]_  = \new_[44423]_  & \new_[44420]_ ;
  assign \new_[44427]_  = ~A298 & ~A268;
  assign \new_[44430]_  = ~A301 & ~A299;
  assign \new_[44431]_  = \new_[44430]_  & \new_[44427]_ ;
  assign \new_[44432]_  = \new_[44431]_  & \new_[44424]_ ;
  assign \new_[44436]_  = ~A168 & ~A169;
  assign \new_[44437]_  = ~A170 & \new_[44436]_ ;
  assign \new_[44440]_  = ~A200 & A199;
  assign \new_[44443]_  = ~A232 & A203;
  assign \new_[44444]_  = \new_[44443]_  & \new_[44440]_ ;
  assign \new_[44445]_  = \new_[44444]_  & \new_[44437]_ ;
  assign \new_[44448]_  = ~A235 & ~A233;
  assign \new_[44451]_  = ~A268 & ~A267;
  assign \new_[44452]_  = \new_[44451]_  & \new_[44448]_ ;
  assign \new_[44455]_  = ~A300 & ~A269;
  assign \new_[44458]_  = ~A302 & ~A301;
  assign \new_[44459]_  = \new_[44458]_  & \new_[44455]_ ;
  assign \new_[44460]_  = \new_[44459]_  & \new_[44452]_ ;
  assign \new_[44464]_  = ~A168 & ~A169;
  assign \new_[44465]_  = ~A170 & \new_[44464]_ ;
  assign \new_[44468]_  = ~A200 & A199;
  assign \new_[44471]_  = ~A232 & A203;
  assign \new_[44472]_  = \new_[44471]_  & \new_[44468]_ ;
  assign \new_[44473]_  = \new_[44472]_  & \new_[44465]_ ;
  assign \new_[44476]_  = ~A235 & ~A233;
  assign \new_[44479]_  = ~A268 & ~A267;
  assign \new_[44480]_  = \new_[44479]_  & \new_[44476]_ ;
  assign \new_[44483]_  = ~A298 & ~A269;
  assign \new_[44486]_  = ~A301 & ~A299;
  assign \new_[44487]_  = \new_[44486]_  & \new_[44483]_ ;
  assign \new_[44488]_  = \new_[44487]_  & \new_[44480]_ ;
  assign \new_[44492]_  = ~A168 & ~A169;
  assign \new_[44493]_  = ~A170 & \new_[44492]_ ;
  assign \new_[44496]_  = ~A200 & A199;
  assign \new_[44499]_  = ~A232 & A203;
  assign \new_[44500]_  = \new_[44499]_  & \new_[44496]_ ;
  assign \new_[44501]_  = \new_[44500]_  & \new_[44493]_ ;
  assign \new_[44504]_  = ~A235 & ~A233;
  assign \new_[44507]_  = ~A266 & ~A265;
  assign \new_[44508]_  = \new_[44507]_  & \new_[44504]_ ;
  assign \new_[44511]_  = ~A300 & ~A268;
  assign \new_[44514]_  = ~A302 & ~A301;
  assign \new_[44515]_  = \new_[44514]_  & \new_[44511]_ ;
  assign \new_[44516]_  = \new_[44515]_  & \new_[44508]_ ;
  assign \new_[44520]_  = ~A168 & ~A169;
  assign \new_[44521]_  = ~A170 & \new_[44520]_ ;
  assign \new_[44524]_  = ~A200 & A199;
  assign \new_[44527]_  = ~A232 & A203;
  assign \new_[44528]_  = \new_[44527]_  & \new_[44524]_ ;
  assign \new_[44529]_  = \new_[44528]_  & \new_[44521]_ ;
  assign \new_[44532]_  = ~A235 & ~A233;
  assign \new_[44535]_  = ~A266 & ~A265;
  assign \new_[44536]_  = \new_[44535]_  & \new_[44532]_ ;
  assign \new_[44539]_  = ~A298 & ~A268;
  assign \new_[44542]_  = ~A301 & ~A299;
  assign \new_[44543]_  = \new_[44542]_  & \new_[44539]_ ;
  assign \new_[44544]_  = \new_[44543]_  & \new_[44536]_ ;
  assign \new_[44547]_  = A166 & A168;
  assign \new_[44550]_  = ~A202 & ~A201;
  assign \new_[44551]_  = \new_[44550]_  & \new_[44547]_ ;
  assign \new_[44554]_  = ~A234 & ~A203;
  assign \new_[44557]_  = ~A236 & ~A235;
  assign \new_[44558]_  = \new_[44557]_  & \new_[44554]_ ;
  assign \new_[44559]_  = \new_[44558]_  & \new_[44551]_ ;
  assign \new_[44562]_  = A266 & A265;
  assign \new_[44565]_  = ~A268 & ~A267;
  assign \new_[44566]_  = \new_[44565]_  & \new_[44562]_ ;
  assign \new_[44569]_  = A299 & A298;
  assign \new_[44572]_  = ~A301 & ~A300;
  assign \new_[44573]_  = \new_[44572]_  & \new_[44569]_ ;
  assign \new_[44574]_  = \new_[44573]_  & \new_[44566]_ ;
  assign \new_[44577]_  = A166 & A168;
  assign \new_[44580]_  = ~A202 & ~A201;
  assign \new_[44581]_  = \new_[44580]_  & \new_[44577]_ ;
  assign \new_[44584]_  = A232 & ~A203;
  assign \new_[44587]_  = ~A234 & A233;
  assign \new_[44588]_  = \new_[44587]_  & \new_[44584]_ ;
  assign \new_[44589]_  = \new_[44588]_  & \new_[44581]_ ;
  assign \new_[44592]_  = ~A267 & ~A235;
  assign \new_[44595]_  = ~A269 & ~A268;
  assign \new_[44596]_  = \new_[44595]_  & \new_[44592]_ ;
  assign \new_[44599]_  = A299 & A298;
  assign \new_[44602]_  = ~A301 & ~A300;
  assign \new_[44603]_  = \new_[44602]_  & \new_[44599]_ ;
  assign \new_[44604]_  = \new_[44603]_  & \new_[44596]_ ;
  assign \new_[44607]_  = A166 & A168;
  assign \new_[44610]_  = ~A202 & ~A201;
  assign \new_[44611]_  = \new_[44610]_  & \new_[44607]_ ;
  assign \new_[44614]_  = A232 & ~A203;
  assign \new_[44617]_  = ~A234 & A233;
  assign \new_[44618]_  = \new_[44617]_  & \new_[44614]_ ;
  assign \new_[44619]_  = \new_[44618]_  & \new_[44611]_ ;
  assign \new_[44622]_  = A265 & ~A235;
  assign \new_[44625]_  = ~A267 & A266;
  assign \new_[44626]_  = \new_[44625]_  & \new_[44622]_ ;
  assign \new_[44629]_  = ~A300 & ~A268;
  assign \new_[44632]_  = ~A302 & ~A301;
  assign \new_[44633]_  = \new_[44632]_  & \new_[44629]_ ;
  assign \new_[44634]_  = \new_[44633]_  & \new_[44626]_ ;
  assign \new_[44637]_  = A166 & A168;
  assign \new_[44640]_  = ~A202 & ~A201;
  assign \new_[44641]_  = \new_[44640]_  & \new_[44637]_ ;
  assign \new_[44644]_  = A232 & ~A203;
  assign \new_[44647]_  = ~A234 & A233;
  assign \new_[44648]_  = \new_[44647]_  & \new_[44644]_ ;
  assign \new_[44649]_  = \new_[44648]_  & \new_[44641]_ ;
  assign \new_[44652]_  = A265 & ~A235;
  assign \new_[44655]_  = ~A267 & A266;
  assign \new_[44656]_  = \new_[44655]_  & \new_[44652]_ ;
  assign \new_[44659]_  = ~A298 & ~A268;
  assign \new_[44662]_  = ~A301 & ~A299;
  assign \new_[44663]_  = \new_[44662]_  & \new_[44659]_ ;
  assign \new_[44664]_  = \new_[44663]_  & \new_[44656]_ ;
  assign \new_[44667]_  = A166 & A168;
  assign \new_[44670]_  = ~A202 & ~A201;
  assign \new_[44671]_  = \new_[44670]_  & \new_[44667]_ ;
  assign \new_[44674]_  = A232 & ~A203;
  assign \new_[44677]_  = ~A234 & A233;
  assign \new_[44678]_  = \new_[44677]_  & \new_[44674]_ ;
  assign \new_[44679]_  = \new_[44678]_  & \new_[44671]_ ;
  assign \new_[44682]_  = ~A265 & ~A235;
  assign \new_[44685]_  = ~A268 & ~A266;
  assign \new_[44686]_  = \new_[44685]_  & \new_[44682]_ ;
  assign \new_[44689]_  = A299 & A298;
  assign \new_[44692]_  = ~A301 & ~A300;
  assign \new_[44693]_  = \new_[44692]_  & \new_[44689]_ ;
  assign \new_[44694]_  = \new_[44693]_  & \new_[44686]_ ;
  assign \new_[44697]_  = A166 & A168;
  assign \new_[44700]_  = ~A202 & ~A201;
  assign \new_[44701]_  = \new_[44700]_  & \new_[44697]_ ;
  assign \new_[44704]_  = ~A232 & ~A203;
  assign \new_[44707]_  = ~A235 & ~A233;
  assign \new_[44708]_  = \new_[44707]_  & \new_[44704]_ ;
  assign \new_[44709]_  = \new_[44708]_  & \new_[44701]_ ;
  assign \new_[44712]_  = A266 & A265;
  assign \new_[44715]_  = ~A268 & ~A267;
  assign \new_[44716]_  = \new_[44715]_  & \new_[44712]_ ;
  assign \new_[44719]_  = A299 & A298;
  assign \new_[44722]_  = ~A301 & ~A300;
  assign \new_[44723]_  = \new_[44722]_  & \new_[44719]_ ;
  assign \new_[44724]_  = \new_[44723]_  & \new_[44716]_ ;
  assign \new_[44727]_  = A166 & A168;
  assign \new_[44730]_  = A200 & A199;
  assign \new_[44731]_  = \new_[44730]_  & \new_[44727]_ ;
  assign \new_[44734]_  = ~A202 & ~A201;
  assign \new_[44737]_  = ~A235 & ~A234;
  assign \new_[44738]_  = \new_[44737]_  & \new_[44734]_ ;
  assign \new_[44739]_  = \new_[44738]_  & \new_[44731]_ ;
  assign \new_[44742]_  = ~A267 & ~A236;
  assign \new_[44745]_  = ~A269 & ~A268;
  assign \new_[44746]_  = \new_[44745]_  & \new_[44742]_ ;
  assign \new_[44749]_  = A299 & A298;
  assign \new_[44752]_  = ~A301 & ~A300;
  assign \new_[44753]_  = \new_[44752]_  & \new_[44749]_ ;
  assign \new_[44754]_  = \new_[44753]_  & \new_[44746]_ ;
  assign \new_[44757]_  = A166 & A168;
  assign \new_[44760]_  = A200 & A199;
  assign \new_[44761]_  = \new_[44760]_  & \new_[44757]_ ;
  assign \new_[44764]_  = ~A202 & ~A201;
  assign \new_[44767]_  = ~A235 & ~A234;
  assign \new_[44768]_  = \new_[44767]_  & \new_[44764]_ ;
  assign \new_[44769]_  = \new_[44768]_  & \new_[44761]_ ;
  assign \new_[44772]_  = A265 & ~A236;
  assign \new_[44775]_  = ~A267 & A266;
  assign \new_[44776]_  = \new_[44775]_  & \new_[44772]_ ;
  assign \new_[44779]_  = ~A300 & ~A268;
  assign \new_[44782]_  = ~A302 & ~A301;
  assign \new_[44783]_  = \new_[44782]_  & \new_[44779]_ ;
  assign \new_[44784]_  = \new_[44783]_  & \new_[44776]_ ;
  assign \new_[44787]_  = A166 & A168;
  assign \new_[44790]_  = A200 & A199;
  assign \new_[44791]_  = \new_[44790]_  & \new_[44787]_ ;
  assign \new_[44794]_  = ~A202 & ~A201;
  assign \new_[44797]_  = ~A235 & ~A234;
  assign \new_[44798]_  = \new_[44797]_  & \new_[44794]_ ;
  assign \new_[44799]_  = \new_[44798]_  & \new_[44791]_ ;
  assign \new_[44802]_  = A265 & ~A236;
  assign \new_[44805]_  = ~A267 & A266;
  assign \new_[44806]_  = \new_[44805]_  & \new_[44802]_ ;
  assign \new_[44809]_  = ~A298 & ~A268;
  assign \new_[44812]_  = ~A301 & ~A299;
  assign \new_[44813]_  = \new_[44812]_  & \new_[44809]_ ;
  assign \new_[44814]_  = \new_[44813]_  & \new_[44806]_ ;
  assign \new_[44817]_  = A166 & A168;
  assign \new_[44820]_  = A200 & A199;
  assign \new_[44821]_  = \new_[44820]_  & \new_[44817]_ ;
  assign \new_[44824]_  = ~A202 & ~A201;
  assign \new_[44827]_  = ~A235 & ~A234;
  assign \new_[44828]_  = \new_[44827]_  & \new_[44824]_ ;
  assign \new_[44829]_  = \new_[44828]_  & \new_[44821]_ ;
  assign \new_[44832]_  = ~A265 & ~A236;
  assign \new_[44835]_  = ~A268 & ~A266;
  assign \new_[44836]_  = \new_[44835]_  & \new_[44832]_ ;
  assign \new_[44839]_  = A299 & A298;
  assign \new_[44842]_  = ~A301 & ~A300;
  assign \new_[44843]_  = \new_[44842]_  & \new_[44839]_ ;
  assign \new_[44844]_  = \new_[44843]_  & \new_[44836]_ ;
  assign \new_[44847]_  = A166 & A168;
  assign \new_[44850]_  = A200 & A199;
  assign \new_[44851]_  = \new_[44850]_  & \new_[44847]_ ;
  assign \new_[44854]_  = ~A202 & ~A201;
  assign \new_[44857]_  = A233 & A232;
  assign \new_[44858]_  = \new_[44857]_  & \new_[44854]_ ;
  assign \new_[44859]_  = \new_[44858]_  & \new_[44851]_ ;
  assign \new_[44862]_  = ~A235 & ~A234;
  assign \new_[44865]_  = ~A268 & ~A267;
  assign \new_[44866]_  = \new_[44865]_  & \new_[44862]_ ;
  assign \new_[44869]_  = ~A300 & ~A269;
  assign \new_[44872]_  = ~A302 & ~A301;
  assign \new_[44873]_  = \new_[44872]_  & \new_[44869]_ ;
  assign \new_[44874]_  = \new_[44873]_  & \new_[44866]_ ;
  assign \new_[44877]_  = A166 & A168;
  assign \new_[44880]_  = A200 & A199;
  assign \new_[44881]_  = \new_[44880]_  & \new_[44877]_ ;
  assign \new_[44884]_  = ~A202 & ~A201;
  assign \new_[44887]_  = A233 & A232;
  assign \new_[44888]_  = \new_[44887]_  & \new_[44884]_ ;
  assign \new_[44889]_  = \new_[44888]_  & \new_[44881]_ ;
  assign \new_[44892]_  = ~A235 & ~A234;
  assign \new_[44895]_  = ~A268 & ~A267;
  assign \new_[44896]_  = \new_[44895]_  & \new_[44892]_ ;
  assign \new_[44899]_  = ~A298 & ~A269;
  assign \new_[44902]_  = ~A301 & ~A299;
  assign \new_[44903]_  = \new_[44902]_  & \new_[44899]_ ;
  assign \new_[44904]_  = \new_[44903]_  & \new_[44896]_ ;
  assign \new_[44907]_  = A166 & A168;
  assign \new_[44910]_  = A200 & A199;
  assign \new_[44911]_  = \new_[44910]_  & \new_[44907]_ ;
  assign \new_[44914]_  = ~A202 & ~A201;
  assign \new_[44917]_  = A233 & A232;
  assign \new_[44918]_  = \new_[44917]_  & \new_[44914]_ ;
  assign \new_[44919]_  = \new_[44918]_  & \new_[44911]_ ;
  assign \new_[44922]_  = ~A235 & ~A234;
  assign \new_[44925]_  = ~A266 & ~A265;
  assign \new_[44926]_  = \new_[44925]_  & \new_[44922]_ ;
  assign \new_[44929]_  = ~A300 & ~A268;
  assign \new_[44932]_  = ~A302 & ~A301;
  assign \new_[44933]_  = \new_[44932]_  & \new_[44929]_ ;
  assign \new_[44934]_  = \new_[44933]_  & \new_[44926]_ ;
  assign \new_[44937]_  = A166 & A168;
  assign \new_[44940]_  = A200 & A199;
  assign \new_[44941]_  = \new_[44940]_  & \new_[44937]_ ;
  assign \new_[44944]_  = ~A202 & ~A201;
  assign \new_[44947]_  = A233 & A232;
  assign \new_[44948]_  = \new_[44947]_  & \new_[44944]_ ;
  assign \new_[44949]_  = \new_[44948]_  & \new_[44941]_ ;
  assign \new_[44952]_  = ~A235 & ~A234;
  assign \new_[44955]_  = ~A266 & ~A265;
  assign \new_[44956]_  = \new_[44955]_  & \new_[44952]_ ;
  assign \new_[44959]_  = ~A298 & ~A268;
  assign \new_[44962]_  = ~A301 & ~A299;
  assign \new_[44963]_  = \new_[44962]_  & \new_[44959]_ ;
  assign \new_[44964]_  = \new_[44963]_  & \new_[44956]_ ;
  assign \new_[44967]_  = A166 & A168;
  assign \new_[44970]_  = A200 & A199;
  assign \new_[44971]_  = \new_[44970]_  & \new_[44967]_ ;
  assign \new_[44974]_  = ~A202 & ~A201;
  assign \new_[44977]_  = ~A233 & ~A232;
  assign \new_[44978]_  = \new_[44977]_  & \new_[44974]_ ;
  assign \new_[44979]_  = \new_[44978]_  & \new_[44971]_ ;
  assign \new_[44982]_  = ~A267 & ~A235;
  assign \new_[44985]_  = ~A269 & ~A268;
  assign \new_[44986]_  = \new_[44985]_  & \new_[44982]_ ;
  assign \new_[44989]_  = A299 & A298;
  assign \new_[44992]_  = ~A301 & ~A300;
  assign \new_[44993]_  = \new_[44992]_  & \new_[44989]_ ;
  assign \new_[44994]_  = \new_[44993]_  & \new_[44986]_ ;
  assign \new_[44997]_  = A166 & A168;
  assign \new_[45000]_  = A200 & A199;
  assign \new_[45001]_  = \new_[45000]_  & \new_[44997]_ ;
  assign \new_[45004]_  = ~A202 & ~A201;
  assign \new_[45007]_  = ~A233 & ~A232;
  assign \new_[45008]_  = \new_[45007]_  & \new_[45004]_ ;
  assign \new_[45009]_  = \new_[45008]_  & \new_[45001]_ ;
  assign \new_[45012]_  = A265 & ~A235;
  assign \new_[45015]_  = ~A267 & A266;
  assign \new_[45016]_  = \new_[45015]_  & \new_[45012]_ ;
  assign \new_[45019]_  = ~A300 & ~A268;
  assign \new_[45022]_  = ~A302 & ~A301;
  assign \new_[45023]_  = \new_[45022]_  & \new_[45019]_ ;
  assign \new_[45024]_  = \new_[45023]_  & \new_[45016]_ ;
  assign \new_[45027]_  = A166 & A168;
  assign \new_[45030]_  = A200 & A199;
  assign \new_[45031]_  = \new_[45030]_  & \new_[45027]_ ;
  assign \new_[45034]_  = ~A202 & ~A201;
  assign \new_[45037]_  = ~A233 & ~A232;
  assign \new_[45038]_  = \new_[45037]_  & \new_[45034]_ ;
  assign \new_[45039]_  = \new_[45038]_  & \new_[45031]_ ;
  assign \new_[45042]_  = A265 & ~A235;
  assign \new_[45045]_  = ~A267 & A266;
  assign \new_[45046]_  = \new_[45045]_  & \new_[45042]_ ;
  assign \new_[45049]_  = ~A298 & ~A268;
  assign \new_[45052]_  = ~A301 & ~A299;
  assign \new_[45053]_  = \new_[45052]_  & \new_[45049]_ ;
  assign \new_[45054]_  = \new_[45053]_  & \new_[45046]_ ;
  assign \new_[45057]_  = A166 & A168;
  assign \new_[45060]_  = A200 & A199;
  assign \new_[45061]_  = \new_[45060]_  & \new_[45057]_ ;
  assign \new_[45064]_  = ~A202 & ~A201;
  assign \new_[45067]_  = ~A233 & ~A232;
  assign \new_[45068]_  = \new_[45067]_  & \new_[45064]_ ;
  assign \new_[45069]_  = \new_[45068]_  & \new_[45061]_ ;
  assign \new_[45072]_  = ~A265 & ~A235;
  assign \new_[45075]_  = ~A268 & ~A266;
  assign \new_[45076]_  = \new_[45075]_  & \new_[45072]_ ;
  assign \new_[45079]_  = A299 & A298;
  assign \new_[45082]_  = ~A301 & ~A300;
  assign \new_[45083]_  = \new_[45082]_  & \new_[45079]_ ;
  assign \new_[45084]_  = \new_[45083]_  & \new_[45076]_ ;
  assign \new_[45087]_  = A166 & A168;
  assign \new_[45090]_  = ~A200 & ~A199;
  assign \new_[45091]_  = \new_[45090]_  & \new_[45087]_ ;
  assign \new_[45094]_  = ~A234 & ~A202;
  assign \new_[45097]_  = ~A236 & ~A235;
  assign \new_[45098]_  = \new_[45097]_  & \new_[45094]_ ;
  assign \new_[45099]_  = \new_[45098]_  & \new_[45091]_ ;
  assign \new_[45102]_  = A266 & A265;
  assign \new_[45105]_  = ~A268 & ~A267;
  assign \new_[45106]_  = \new_[45105]_  & \new_[45102]_ ;
  assign \new_[45109]_  = A299 & A298;
  assign \new_[45112]_  = ~A301 & ~A300;
  assign \new_[45113]_  = \new_[45112]_  & \new_[45109]_ ;
  assign \new_[45114]_  = \new_[45113]_  & \new_[45106]_ ;
  assign \new_[45117]_  = A166 & A168;
  assign \new_[45120]_  = ~A200 & ~A199;
  assign \new_[45121]_  = \new_[45120]_  & \new_[45117]_ ;
  assign \new_[45124]_  = A232 & ~A202;
  assign \new_[45127]_  = ~A234 & A233;
  assign \new_[45128]_  = \new_[45127]_  & \new_[45124]_ ;
  assign \new_[45129]_  = \new_[45128]_  & \new_[45121]_ ;
  assign \new_[45132]_  = ~A267 & ~A235;
  assign \new_[45135]_  = ~A269 & ~A268;
  assign \new_[45136]_  = \new_[45135]_  & \new_[45132]_ ;
  assign \new_[45139]_  = A299 & A298;
  assign \new_[45142]_  = ~A301 & ~A300;
  assign \new_[45143]_  = \new_[45142]_  & \new_[45139]_ ;
  assign \new_[45144]_  = \new_[45143]_  & \new_[45136]_ ;
  assign \new_[45147]_  = A166 & A168;
  assign \new_[45150]_  = ~A200 & ~A199;
  assign \new_[45151]_  = \new_[45150]_  & \new_[45147]_ ;
  assign \new_[45154]_  = A232 & ~A202;
  assign \new_[45157]_  = ~A234 & A233;
  assign \new_[45158]_  = \new_[45157]_  & \new_[45154]_ ;
  assign \new_[45159]_  = \new_[45158]_  & \new_[45151]_ ;
  assign \new_[45162]_  = A265 & ~A235;
  assign \new_[45165]_  = ~A267 & A266;
  assign \new_[45166]_  = \new_[45165]_  & \new_[45162]_ ;
  assign \new_[45169]_  = ~A300 & ~A268;
  assign \new_[45172]_  = ~A302 & ~A301;
  assign \new_[45173]_  = \new_[45172]_  & \new_[45169]_ ;
  assign \new_[45174]_  = \new_[45173]_  & \new_[45166]_ ;
  assign \new_[45177]_  = A166 & A168;
  assign \new_[45180]_  = ~A200 & ~A199;
  assign \new_[45181]_  = \new_[45180]_  & \new_[45177]_ ;
  assign \new_[45184]_  = A232 & ~A202;
  assign \new_[45187]_  = ~A234 & A233;
  assign \new_[45188]_  = \new_[45187]_  & \new_[45184]_ ;
  assign \new_[45189]_  = \new_[45188]_  & \new_[45181]_ ;
  assign \new_[45192]_  = A265 & ~A235;
  assign \new_[45195]_  = ~A267 & A266;
  assign \new_[45196]_  = \new_[45195]_  & \new_[45192]_ ;
  assign \new_[45199]_  = ~A298 & ~A268;
  assign \new_[45202]_  = ~A301 & ~A299;
  assign \new_[45203]_  = \new_[45202]_  & \new_[45199]_ ;
  assign \new_[45204]_  = \new_[45203]_  & \new_[45196]_ ;
  assign \new_[45207]_  = A166 & A168;
  assign \new_[45210]_  = ~A200 & ~A199;
  assign \new_[45211]_  = \new_[45210]_  & \new_[45207]_ ;
  assign \new_[45214]_  = A232 & ~A202;
  assign \new_[45217]_  = ~A234 & A233;
  assign \new_[45218]_  = \new_[45217]_  & \new_[45214]_ ;
  assign \new_[45219]_  = \new_[45218]_  & \new_[45211]_ ;
  assign \new_[45222]_  = ~A265 & ~A235;
  assign \new_[45225]_  = ~A268 & ~A266;
  assign \new_[45226]_  = \new_[45225]_  & \new_[45222]_ ;
  assign \new_[45229]_  = A299 & A298;
  assign \new_[45232]_  = ~A301 & ~A300;
  assign \new_[45233]_  = \new_[45232]_  & \new_[45229]_ ;
  assign \new_[45234]_  = \new_[45233]_  & \new_[45226]_ ;
  assign \new_[45237]_  = A166 & A168;
  assign \new_[45240]_  = ~A200 & ~A199;
  assign \new_[45241]_  = \new_[45240]_  & \new_[45237]_ ;
  assign \new_[45244]_  = ~A232 & ~A202;
  assign \new_[45247]_  = ~A235 & ~A233;
  assign \new_[45248]_  = \new_[45247]_  & \new_[45244]_ ;
  assign \new_[45249]_  = \new_[45248]_  & \new_[45241]_ ;
  assign \new_[45252]_  = A266 & A265;
  assign \new_[45255]_  = ~A268 & ~A267;
  assign \new_[45256]_  = \new_[45255]_  & \new_[45252]_ ;
  assign \new_[45259]_  = A299 & A298;
  assign \new_[45262]_  = ~A301 & ~A300;
  assign \new_[45263]_  = \new_[45262]_  & \new_[45259]_ ;
  assign \new_[45264]_  = \new_[45263]_  & \new_[45256]_ ;
  assign \new_[45267]_  = A167 & A168;
  assign \new_[45270]_  = ~A202 & ~A201;
  assign \new_[45271]_  = \new_[45270]_  & \new_[45267]_ ;
  assign \new_[45274]_  = ~A234 & ~A203;
  assign \new_[45277]_  = ~A236 & ~A235;
  assign \new_[45278]_  = \new_[45277]_  & \new_[45274]_ ;
  assign \new_[45279]_  = \new_[45278]_  & \new_[45271]_ ;
  assign \new_[45282]_  = A266 & A265;
  assign \new_[45285]_  = ~A268 & ~A267;
  assign \new_[45286]_  = \new_[45285]_  & \new_[45282]_ ;
  assign \new_[45289]_  = A299 & A298;
  assign \new_[45292]_  = ~A301 & ~A300;
  assign \new_[45293]_  = \new_[45292]_  & \new_[45289]_ ;
  assign \new_[45294]_  = \new_[45293]_  & \new_[45286]_ ;
  assign \new_[45297]_  = A167 & A168;
  assign \new_[45300]_  = ~A202 & ~A201;
  assign \new_[45301]_  = \new_[45300]_  & \new_[45297]_ ;
  assign \new_[45304]_  = A232 & ~A203;
  assign \new_[45307]_  = ~A234 & A233;
  assign \new_[45308]_  = \new_[45307]_  & \new_[45304]_ ;
  assign \new_[45309]_  = \new_[45308]_  & \new_[45301]_ ;
  assign \new_[45312]_  = ~A267 & ~A235;
  assign \new_[45315]_  = ~A269 & ~A268;
  assign \new_[45316]_  = \new_[45315]_  & \new_[45312]_ ;
  assign \new_[45319]_  = A299 & A298;
  assign \new_[45322]_  = ~A301 & ~A300;
  assign \new_[45323]_  = \new_[45322]_  & \new_[45319]_ ;
  assign \new_[45324]_  = \new_[45323]_  & \new_[45316]_ ;
  assign \new_[45327]_  = A167 & A168;
  assign \new_[45330]_  = ~A202 & ~A201;
  assign \new_[45331]_  = \new_[45330]_  & \new_[45327]_ ;
  assign \new_[45334]_  = A232 & ~A203;
  assign \new_[45337]_  = ~A234 & A233;
  assign \new_[45338]_  = \new_[45337]_  & \new_[45334]_ ;
  assign \new_[45339]_  = \new_[45338]_  & \new_[45331]_ ;
  assign \new_[45342]_  = A265 & ~A235;
  assign \new_[45345]_  = ~A267 & A266;
  assign \new_[45346]_  = \new_[45345]_  & \new_[45342]_ ;
  assign \new_[45349]_  = ~A300 & ~A268;
  assign \new_[45352]_  = ~A302 & ~A301;
  assign \new_[45353]_  = \new_[45352]_  & \new_[45349]_ ;
  assign \new_[45354]_  = \new_[45353]_  & \new_[45346]_ ;
  assign \new_[45357]_  = A167 & A168;
  assign \new_[45360]_  = ~A202 & ~A201;
  assign \new_[45361]_  = \new_[45360]_  & \new_[45357]_ ;
  assign \new_[45364]_  = A232 & ~A203;
  assign \new_[45367]_  = ~A234 & A233;
  assign \new_[45368]_  = \new_[45367]_  & \new_[45364]_ ;
  assign \new_[45369]_  = \new_[45368]_  & \new_[45361]_ ;
  assign \new_[45372]_  = A265 & ~A235;
  assign \new_[45375]_  = ~A267 & A266;
  assign \new_[45376]_  = \new_[45375]_  & \new_[45372]_ ;
  assign \new_[45379]_  = ~A298 & ~A268;
  assign \new_[45382]_  = ~A301 & ~A299;
  assign \new_[45383]_  = \new_[45382]_  & \new_[45379]_ ;
  assign \new_[45384]_  = \new_[45383]_  & \new_[45376]_ ;
  assign \new_[45387]_  = A167 & A168;
  assign \new_[45390]_  = ~A202 & ~A201;
  assign \new_[45391]_  = \new_[45390]_  & \new_[45387]_ ;
  assign \new_[45394]_  = A232 & ~A203;
  assign \new_[45397]_  = ~A234 & A233;
  assign \new_[45398]_  = \new_[45397]_  & \new_[45394]_ ;
  assign \new_[45399]_  = \new_[45398]_  & \new_[45391]_ ;
  assign \new_[45402]_  = ~A265 & ~A235;
  assign \new_[45405]_  = ~A268 & ~A266;
  assign \new_[45406]_  = \new_[45405]_  & \new_[45402]_ ;
  assign \new_[45409]_  = A299 & A298;
  assign \new_[45412]_  = ~A301 & ~A300;
  assign \new_[45413]_  = \new_[45412]_  & \new_[45409]_ ;
  assign \new_[45414]_  = \new_[45413]_  & \new_[45406]_ ;
  assign \new_[45417]_  = A167 & A168;
  assign \new_[45420]_  = ~A202 & ~A201;
  assign \new_[45421]_  = \new_[45420]_  & \new_[45417]_ ;
  assign \new_[45424]_  = ~A232 & ~A203;
  assign \new_[45427]_  = ~A235 & ~A233;
  assign \new_[45428]_  = \new_[45427]_  & \new_[45424]_ ;
  assign \new_[45429]_  = \new_[45428]_  & \new_[45421]_ ;
  assign \new_[45432]_  = A266 & A265;
  assign \new_[45435]_  = ~A268 & ~A267;
  assign \new_[45436]_  = \new_[45435]_  & \new_[45432]_ ;
  assign \new_[45439]_  = A299 & A298;
  assign \new_[45442]_  = ~A301 & ~A300;
  assign \new_[45443]_  = \new_[45442]_  & \new_[45439]_ ;
  assign \new_[45444]_  = \new_[45443]_  & \new_[45436]_ ;
  assign \new_[45447]_  = A167 & A168;
  assign \new_[45450]_  = A200 & A199;
  assign \new_[45451]_  = \new_[45450]_  & \new_[45447]_ ;
  assign \new_[45454]_  = ~A202 & ~A201;
  assign \new_[45457]_  = ~A235 & ~A234;
  assign \new_[45458]_  = \new_[45457]_  & \new_[45454]_ ;
  assign \new_[45459]_  = \new_[45458]_  & \new_[45451]_ ;
  assign \new_[45462]_  = ~A267 & ~A236;
  assign \new_[45465]_  = ~A269 & ~A268;
  assign \new_[45466]_  = \new_[45465]_  & \new_[45462]_ ;
  assign \new_[45469]_  = A299 & A298;
  assign \new_[45472]_  = ~A301 & ~A300;
  assign \new_[45473]_  = \new_[45472]_  & \new_[45469]_ ;
  assign \new_[45474]_  = \new_[45473]_  & \new_[45466]_ ;
  assign \new_[45477]_  = A167 & A168;
  assign \new_[45480]_  = A200 & A199;
  assign \new_[45481]_  = \new_[45480]_  & \new_[45477]_ ;
  assign \new_[45484]_  = ~A202 & ~A201;
  assign \new_[45487]_  = ~A235 & ~A234;
  assign \new_[45488]_  = \new_[45487]_  & \new_[45484]_ ;
  assign \new_[45489]_  = \new_[45488]_  & \new_[45481]_ ;
  assign \new_[45492]_  = A265 & ~A236;
  assign \new_[45495]_  = ~A267 & A266;
  assign \new_[45496]_  = \new_[45495]_  & \new_[45492]_ ;
  assign \new_[45499]_  = ~A300 & ~A268;
  assign \new_[45502]_  = ~A302 & ~A301;
  assign \new_[45503]_  = \new_[45502]_  & \new_[45499]_ ;
  assign \new_[45504]_  = \new_[45503]_  & \new_[45496]_ ;
  assign \new_[45507]_  = A167 & A168;
  assign \new_[45510]_  = A200 & A199;
  assign \new_[45511]_  = \new_[45510]_  & \new_[45507]_ ;
  assign \new_[45514]_  = ~A202 & ~A201;
  assign \new_[45517]_  = ~A235 & ~A234;
  assign \new_[45518]_  = \new_[45517]_  & \new_[45514]_ ;
  assign \new_[45519]_  = \new_[45518]_  & \new_[45511]_ ;
  assign \new_[45522]_  = A265 & ~A236;
  assign \new_[45525]_  = ~A267 & A266;
  assign \new_[45526]_  = \new_[45525]_  & \new_[45522]_ ;
  assign \new_[45529]_  = ~A298 & ~A268;
  assign \new_[45532]_  = ~A301 & ~A299;
  assign \new_[45533]_  = \new_[45532]_  & \new_[45529]_ ;
  assign \new_[45534]_  = \new_[45533]_  & \new_[45526]_ ;
  assign \new_[45537]_  = A167 & A168;
  assign \new_[45540]_  = A200 & A199;
  assign \new_[45541]_  = \new_[45540]_  & \new_[45537]_ ;
  assign \new_[45544]_  = ~A202 & ~A201;
  assign \new_[45547]_  = ~A235 & ~A234;
  assign \new_[45548]_  = \new_[45547]_  & \new_[45544]_ ;
  assign \new_[45549]_  = \new_[45548]_  & \new_[45541]_ ;
  assign \new_[45552]_  = ~A265 & ~A236;
  assign \new_[45555]_  = ~A268 & ~A266;
  assign \new_[45556]_  = \new_[45555]_  & \new_[45552]_ ;
  assign \new_[45559]_  = A299 & A298;
  assign \new_[45562]_  = ~A301 & ~A300;
  assign \new_[45563]_  = \new_[45562]_  & \new_[45559]_ ;
  assign \new_[45564]_  = \new_[45563]_  & \new_[45556]_ ;
  assign \new_[45567]_  = A167 & A168;
  assign \new_[45570]_  = A200 & A199;
  assign \new_[45571]_  = \new_[45570]_  & \new_[45567]_ ;
  assign \new_[45574]_  = ~A202 & ~A201;
  assign \new_[45577]_  = A233 & A232;
  assign \new_[45578]_  = \new_[45577]_  & \new_[45574]_ ;
  assign \new_[45579]_  = \new_[45578]_  & \new_[45571]_ ;
  assign \new_[45582]_  = ~A235 & ~A234;
  assign \new_[45585]_  = ~A268 & ~A267;
  assign \new_[45586]_  = \new_[45585]_  & \new_[45582]_ ;
  assign \new_[45589]_  = ~A300 & ~A269;
  assign \new_[45592]_  = ~A302 & ~A301;
  assign \new_[45593]_  = \new_[45592]_  & \new_[45589]_ ;
  assign \new_[45594]_  = \new_[45593]_  & \new_[45586]_ ;
  assign \new_[45597]_  = A167 & A168;
  assign \new_[45600]_  = A200 & A199;
  assign \new_[45601]_  = \new_[45600]_  & \new_[45597]_ ;
  assign \new_[45604]_  = ~A202 & ~A201;
  assign \new_[45607]_  = A233 & A232;
  assign \new_[45608]_  = \new_[45607]_  & \new_[45604]_ ;
  assign \new_[45609]_  = \new_[45608]_  & \new_[45601]_ ;
  assign \new_[45612]_  = ~A235 & ~A234;
  assign \new_[45615]_  = ~A268 & ~A267;
  assign \new_[45616]_  = \new_[45615]_  & \new_[45612]_ ;
  assign \new_[45619]_  = ~A298 & ~A269;
  assign \new_[45622]_  = ~A301 & ~A299;
  assign \new_[45623]_  = \new_[45622]_  & \new_[45619]_ ;
  assign \new_[45624]_  = \new_[45623]_  & \new_[45616]_ ;
  assign \new_[45627]_  = A167 & A168;
  assign \new_[45630]_  = A200 & A199;
  assign \new_[45631]_  = \new_[45630]_  & \new_[45627]_ ;
  assign \new_[45634]_  = ~A202 & ~A201;
  assign \new_[45637]_  = A233 & A232;
  assign \new_[45638]_  = \new_[45637]_  & \new_[45634]_ ;
  assign \new_[45639]_  = \new_[45638]_  & \new_[45631]_ ;
  assign \new_[45642]_  = ~A235 & ~A234;
  assign \new_[45645]_  = ~A266 & ~A265;
  assign \new_[45646]_  = \new_[45645]_  & \new_[45642]_ ;
  assign \new_[45649]_  = ~A300 & ~A268;
  assign \new_[45652]_  = ~A302 & ~A301;
  assign \new_[45653]_  = \new_[45652]_  & \new_[45649]_ ;
  assign \new_[45654]_  = \new_[45653]_  & \new_[45646]_ ;
  assign \new_[45657]_  = A167 & A168;
  assign \new_[45660]_  = A200 & A199;
  assign \new_[45661]_  = \new_[45660]_  & \new_[45657]_ ;
  assign \new_[45664]_  = ~A202 & ~A201;
  assign \new_[45667]_  = A233 & A232;
  assign \new_[45668]_  = \new_[45667]_  & \new_[45664]_ ;
  assign \new_[45669]_  = \new_[45668]_  & \new_[45661]_ ;
  assign \new_[45672]_  = ~A235 & ~A234;
  assign \new_[45675]_  = ~A266 & ~A265;
  assign \new_[45676]_  = \new_[45675]_  & \new_[45672]_ ;
  assign \new_[45679]_  = ~A298 & ~A268;
  assign \new_[45682]_  = ~A301 & ~A299;
  assign \new_[45683]_  = \new_[45682]_  & \new_[45679]_ ;
  assign \new_[45684]_  = \new_[45683]_  & \new_[45676]_ ;
  assign \new_[45687]_  = A167 & A168;
  assign \new_[45690]_  = A200 & A199;
  assign \new_[45691]_  = \new_[45690]_  & \new_[45687]_ ;
  assign \new_[45694]_  = ~A202 & ~A201;
  assign \new_[45697]_  = ~A233 & ~A232;
  assign \new_[45698]_  = \new_[45697]_  & \new_[45694]_ ;
  assign \new_[45699]_  = \new_[45698]_  & \new_[45691]_ ;
  assign \new_[45702]_  = ~A267 & ~A235;
  assign \new_[45705]_  = ~A269 & ~A268;
  assign \new_[45706]_  = \new_[45705]_  & \new_[45702]_ ;
  assign \new_[45709]_  = A299 & A298;
  assign \new_[45712]_  = ~A301 & ~A300;
  assign \new_[45713]_  = \new_[45712]_  & \new_[45709]_ ;
  assign \new_[45714]_  = \new_[45713]_  & \new_[45706]_ ;
  assign \new_[45717]_  = A167 & A168;
  assign \new_[45720]_  = A200 & A199;
  assign \new_[45721]_  = \new_[45720]_  & \new_[45717]_ ;
  assign \new_[45724]_  = ~A202 & ~A201;
  assign \new_[45727]_  = ~A233 & ~A232;
  assign \new_[45728]_  = \new_[45727]_  & \new_[45724]_ ;
  assign \new_[45729]_  = \new_[45728]_  & \new_[45721]_ ;
  assign \new_[45732]_  = A265 & ~A235;
  assign \new_[45735]_  = ~A267 & A266;
  assign \new_[45736]_  = \new_[45735]_  & \new_[45732]_ ;
  assign \new_[45739]_  = ~A300 & ~A268;
  assign \new_[45742]_  = ~A302 & ~A301;
  assign \new_[45743]_  = \new_[45742]_  & \new_[45739]_ ;
  assign \new_[45744]_  = \new_[45743]_  & \new_[45736]_ ;
  assign \new_[45747]_  = A167 & A168;
  assign \new_[45750]_  = A200 & A199;
  assign \new_[45751]_  = \new_[45750]_  & \new_[45747]_ ;
  assign \new_[45754]_  = ~A202 & ~A201;
  assign \new_[45757]_  = ~A233 & ~A232;
  assign \new_[45758]_  = \new_[45757]_  & \new_[45754]_ ;
  assign \new_[45759]_  = \new_[45758]_  & \new_[45751]_ ;
  assign \new_[45762]_  = A265 & ~A235;
  assign \new_[45765]_  = ~A267 & A266;
  assign \new_[45766]_  = \new_[45765]_  & \new_[45762]_ ;
  assign \new_[45769]_  = ~A298 & ~A268;
  assign \new_[45772]_  = ~A301 & ~A299;
  assign \new_[45773]_  = \new_[45772]_  & \new_[45769]_ ;
  assign \new_[45774]_  = \new_[45773]_  & \new_[45766]_ ;
  assign \new_[45777]_  = A167 & A168;
  assign \new_[45780]_  = A200 & A199;
  assign \new_[45781]_  = \new_[45780]_  & \new_[45777]_ ;
  assign \new_[45784]_  = ~A202 & ~A201;
  assign \new_[45787]_  = ~A233 & ~A232;
  assign \new_[45788]_  = \new_[45787]_  & \new_[45784]_ ;
  assign \new_[45789]_  = \new_[45788]_  & \new_[45781]_ ;
  assign \new_[45792]_  = ~A265 & ~A235;
  assign \new_[45795]_  = ~A268 & ~A266;
  assign \new_[45796]_  = \new_[45795]_  & \new_[45792]_ ;
  assign \new_[45799]_  = A299 & A298;
  assign \new_[45802]_  = ~A301 & ~A300;
  assign \new_[45803]_  = \new_[45802]_  & \new_[45799]_ ;
  assign \new_[45804]_  = \new_[45803]_  & \new_[45796]_ ;
  assign \new_[45807]_  = A167 & A168;
  assign \new_[45810]_  = ~A200 & ~A199;
  assign \new_[45811]_  = \new_[45810]_  & \new_[45807]_ ;
  assign \new_[45814]_  = ~A234 & ~A202;
  assign \new_[45817]_  = ~A236 & ~A235;
  assign \new_[45818]_  = \new_[45817]_  & \new_[45814]_ ;
  assign \new_[45819]_  = \new_[45818]_  & \new_[45811]_ ;
  assign \new_[45822]_  = A266 & A265;
  assign \new_[45825]_  = ~A268 & ~A267;
  assign \new_[45826]_  = \new_[45825]_  & \new_[45822]_ ;
  assign \new_[45829]_  = A299 & A298;
  assign \new_[45832]_  = ~A301 & ~A300;
  assign \new_[45833]_  = \new_[45832]_  & \new_[45829]_ ;
  assign \new_[45834]_  = \new_[45833]_  & \new_[45826]_ ;
  assign \new_[45837]_  = A167 & A168;
  assign \new_[45840]_  = ~A200 & ~A199;
  assign \new_[45841]_  = \new_[45840]_  & \new_[45837]_ ;
  assign \new_[45844]_  = A232 & ~A202;
  assign \new_[45847]_  = ~A234 & A233;
  assign \new_[45848]_  = \new_[45847]_  & \new_[45844]_ ;
  assign \new_[45849]_  = \new_[45848]_  & \new_[45841]_ ;
  assign \new_[45852]_  = ~A267 & ~A235;
  assign \new_[45855]_  = ~A269 & ~A268;
  assign \new_[45856]_  = \new_[45855]_  & \new_[45852]_ ;
  assign \new_[45859]_  = A299 & A298;
  assign \new_[45862]_  = ~A301 & ~A300;
  assign \new_[45863]_  = \new_[45862]_  & \new_[45859]_ ;
  assign \new_[45864]_  = \new_[45863]_  & \new_[45856]_ ;
  assign \new_[45867]_  = A167 & A168;
  assign \new_[45870]_  = ~A200 & ~A199;
  assign \new_[45871]_  = \new_[45870]_  & \new_[45867]_ ;
  assign \new_[45874]_  = A232 & ~A202;
  assign \new_[45877]_  = ~A234 & A233;
  assign \new_[45878]_  = \new_[45877]_  & \new_[45874]_ ;
  assign \new_[45879]_  = \new_[45878]_  & \new_[45871]_ ;
  assign \new_[45882]_  = A265 & ~A235;
  assign \new_[45885]_  = ~A267 & A266;
  assign \new_[45886]_  = \new_[45885]_  & \new_[45882]_ ;
  assign \new_[45889]_  = ~A300 & ~A268;
  assign \new_[45892]_  = ~A302 & ~A301;
  assign \new_[45893]_  = \new_[45892]_  & \new_[45889]_ ;
  assign \new_[45894]_  = \new_[45893]_  & \new_[45886]_ ;
  assign \new_[45897]_  = A167 & A168;
  assign \new_[45900]_  = ~A200 & ~A199;
  assign \new_[45901]_  = \new_[45900]_  & \new_[45897]_ ;
  assign \new_[45904]_  = A232 & ~A202;
  assign \new_[45907]_  = ~A234 & A233;
  assign \new_[45908]_  = \new_[45907]_  & \new_[45904]_ ;
  assign \new_[45909]_  = \new_[45908]_  & \new_[45901]_ ;
  assign \new_[45912]_  = A265 & ~A235;
  assign \new_[45915]_  = ~A267 & A266;
  assign \new_[45916]_  = \new_[45915]_  & \new_[45912]_ ;
  assign \new_[45919]_  = ~A298 & ~A268;
  assign \new_[45922]_  = ~A301 & ~A299;
  assign \new_[45923]_  = \new_[45922]_  & \new_[45919]_ ;
  assign \new_[45924]_  = \new_[45923]_  & \new_[45916]_ ;
  assign \new_[45927]_  = A167 & A168;
  assign \new_[45930]_  = ~A200 & ~A199;
  assign \new_[45931]_  = \new_[45930]_  & \new_[45927]_ ;
  assign \new_[45934]_  = A232 & ~A202;
  assign \new_[45937]_  = ~A234 & A233;
  assign \new_[45938]_  = \new_[45937]_  & \new_[45934]_ ;
  assign \new_[45939]_  = \new_[45938]_  & \new_[45931]_ ;
  assign \new_[45942]_  = ~A265 & ~A235;
  assign \new_[45945]_  = ~A268 & ~A266;
  assign \new_[45946]_  = \new_[45945]_  & \new_[45942]_ ;
  assign \new_[45949]_  = A299 & A298;
  assign \new_[45952]_  = ~A301 & ~A300;
  assign \new_[45953]_  = \new_[45952]_  & \new_[45949]_ ;
  assign \new_[45954]_  = \new_[45953]_  & \new_[45946]_ ;
  assign \new_[45957]_  = A167 & A168;
  assign \new_[45960]_  = ~A200 & ~A199;
  assign \new_[45961]_  = \new_[45960]_  & \new_[45957]_ ;
  assign \new_[45964]_  = ~A232 & ~A202;
  assign \new_[45967]_  = ~A235 & ~A233;
  assign \new_[45968]_  = \new_[45967]_  & \new_[45964]_ ;
  assign \new_[45969]_  = \new_[45968]_  & \new_[45961]_ ;
  assign \new_[45972]_  = A266 & A265;
  assign \new_[45975]_  = ~A268 & ~A267;
  assign \new_[45976]_  = \new_[45975]_  & \new_[45972]_ ;
  assign \new_[45979]_  = A299 & A298;
  assign \new_[45982]_  = ~A301 & ~A300;
  assign \new_[45983]_  = \new_[45982]_  & \new_[45979]_ ;
  assign \new_[45984]_  = \new_[45983]_  & \new_[45976]_ ;
  assign \new_[45987]_  = A167 & A170;
  assign \new_[45990]_  = ~A201 & ~A166;
  assign \new_[45991]_  = \new_[45990]_  & \new_[45987]_ ;
  assign \new_[45994]_  = ~A203 & ~A202;
  assign \new_[45997]_  = ~A235 & ~A234;
  assign \new_[45998]_  = \new_[45997]_  & \new_[45994]_ ;
  assign \new_[45999]_  = \new_[45998]_  & \new_[45991]_ ;
  assign \new_[46002]_  = ~A267 & ~A236;
  assign \new_[46005]_  = ~A269 & ~A268;
  assign \new_[46006]_  = \new_[46005]_  & \new_[46002]_ ;
  assign \new_[46009]_  = A299 & A298;
  assign \new_[46012]_  = ~A301 & ~A300;
  assign \new_[46013]_  = \new_[46012]_  & \new_[46009]_ ;
  assign \new_[46014]_  = \new_[46013]_  & \new_[46006]_ ;
  assign \new_[46017]_  = A167 & A170;
  assign \new_[46020]_  = ~A201 & ~A166;
  assign \new_[46021]_  = \new_[46020]_  & \new_[46017]_ ;
  assign \new_[46024]_  = ~A203 & ~A202;
  assign \new_[46027]_  = ~A235 & ~A234;
  assign \new_[46028]_  = \new_[46027]_  & \new_[46024]_ ;
  assign \new_[46029]_  = \new_[46028]_  & \new_[46021]_ ;
  assign \new_[46032]_  = A265 & ~A236;
  assign \new_[46035]_  = ~A267 & A266;
  assign \new_[46036]_  = \new_[46035]_  & \new_[46032]_ ;
  assign \new_[46039]_  = ~A300 & ~A268;
  assign \new_[46042]_  = ~A302 & ~A301;
  assign \new_[46043]_  = \new_[46042]_  & \new_[46039]_ ;
  assign \new_[46044]_  = \new_[46043]_  & \new_[46036]_ ;
  assign \new_[46047]_  = A167 & A170;
  assign \new_[46050]_  = ~A201 & ~A166;
  assign \new_[46051]_  = \new_[46050]_  & \new_[46047]_ ;
  assign \new_[46054]_  = ~A203 & ~A202;
  assign \new_[46057]_  = ~A235 & ~A234;
  assign \new_[46058]_  = \new_[46057]_  & \new_[46054]_ ;
  assign \new_[46059]_  = \new_[46058]_  & \new_[46051]_ ;
  assign \new_[46062]_  = A265 & ~A236;
  assign \new_[46065]_  = ~A267 & A266;
  assign \new_[46066]_  = \new_[46065]_  & \new_[46062]_ ;
  assign \new_[46069]_  = ~A298 & ~A268;
  assign \new_[46072]_  = ~A301 & ~A299;
  assign \new_[46073]_  = \new_[46072]_  & \new_[46069]_ ;
  assign \new_[46074]_  = \new_[46073]_  & \new_[46066]_ ;
  assign \new_[46077]_  = A167 & A170;
  assign \new_[46080]_  = ~A201 & ~A166;
  assign \new_[46081]_  = \new_[46080]_  & \new_[46077]_ ;
  assign \new_[46084]_  = ~A203 & ~A202;
  assign \new_[46087]_  = ~A235 & ~A234;
  assign \new_[46088]_  = \new_[46087]_  & \new_[46084]_ ;
  assign \new_[46089]_  = \new_[46088]_  & \new_[46081]_ ;
  assign \new_[46092]_  = ~A265 & ~A236;
  assign \new_[46095]_  = ~A268 & ~A266;
  assign \new_[46096]_  = \new_[46095]_  & \new_[46092]_ ;
  assign \new_[46099]_  = A299 & A298;
  assign \new_[46102]_  = ~A301 & ~A300;
  assign \new_[46103]_  = \new_[46102]_  & \new_[46099]_ ;
  assign \new_[46104]_  = \new_[46103]_  & \new_[46096]_ ;
  assign \new_[46107]_  = A167 & A170;
  assign \new_[46110]_  = ~A201 & ~A166;
  assign \new_[46111]_  = \new_[46110]_  & \new_[46107]_ ;
  assign \new_[46114]_  = ~A203 & ~A202;
  assign \new_[46117]_  = A233 & A232;
  assign \new_[46118]_  = \new_[46117]_  & \new_[46114]_ ;
  assign \new_[46119]_  = \new_[46118]_  & \new_[46111]_ ;
  assign \new_[46122]_  = ~A235 & ~A234;
  assign \new_[46125]_  = ~A268 & ~A267;
  assign \new_[46126]_  = \new_[46125]_  & \new_[46122]_ ;
  assign \new_[46129]_  = ~A300 & ~A269;
  assign \new_[46132]_  = ~A302 & ~A301;
  assign \new_[46133]_  = \new_[46132]_  & \new_[46129]_ ;
  assign \new_[46134]_  = \new_[46133]_  & \new_[46126]_ ;
  assign \new_[46137]_  = A167 & A170;
  assign \new_[46140]_  = ~A201 & ~A166;
  assign \new_[46141]_  = \new_[46140]_  & \new_[46137]_ ;
  assign \new_[46144]_  = ~A203 & ~A202;
  assign \new_[46147]_  = A233 & A232;
  assign \new_[46148]_  = \new_[46147]_  & \new_[46144]_ ;
  assign \new_[46149]_  = \new_[46148]_  & \new_[46141]_ ;
  assign \new_[46152]_  = ~A235 & ~A234;
  assign \new_[46155]_  = ~A268 & ~A267;
  assign \new_[46156]_  = \new_[46155]_  & \new_[46152]_ ;
  assign \new_[46159]_  = ~A298 & ~A269;
  assign \new_[46162]_  = ~A301 & ~A299;
  assign \new_[46163]_  = \new_[46162]_  & \new_[46159]_ ;
  assign \new_[46164]_  = \new_[46163]_  & \new_[46156]_ ;
  assign \new_[46167]_  = A167 & A170;
  assign \new_[46170]_  = ~A201 & ~A166;
  assign \new_[46171]_  = \new_[46170]_  & \new_[46167]_ ;
  assign \new_[46174]_  = ~A203 & ~A202;
  assign \new_[46177]_  = A233 & A232;
  assign \new_[46178]_  = \new_[46177]_  & \new_[46174]_ ;
  assign \new_[46179]_  = \new_[46178]_  & \new_[46171]_ ;
  assign \new_[46182]_  = ~A235 & ~A234;
  assign \new_[46185]_  = ~A266 & ~A265;
  assign \new_[46186]_  = \new_[46185]_  & \new_[46182]_ ;
  assign \new_[46189]_  = ~A300 & ~A268;
  assign \new_[46192]_  = ~A302 & ~A301;
  assign \new_[46193]_  = \new_[46192]_  & \new_[46189]_ ;
  assign \new_[46194]_  = \new_[46193]_  & \new_[46186]_ ;
  assign \new_[46197]_  = A167 & A170;
  assign \new_[46200]_  = ~A201 & ~A166;
  assign \new_[46201]_  = \new_[46200]_  & \new_[46197]_ ;
  assign \new_[46204]_  = ~A203 & ~A202;
  assign \new_[46207]_  = A233 & A232;
  assign \new_[46208]_  = \new_[46207]_  & \new_[46204]_ ;
  assign \new_[46209]_  = \new_[46208]_  & \new_[46201]_ ;
  assign \new_[46212]_  = ~A235 & ~A234;
  assign \new_[46215]_  = ~A266 & ~A265;
  assign \new_[46216]_  = \new_[46215]_  & \new_[46212]_ ;
  assign \new_[46219]_  = ~A298 & ~A268;
  assign \new_[46222]_  = ~A301 & ~A299;
  assign \new_[46223]_  = \new_[46222]_  & \new_[46219]_ ;
  assign \new_[46224]_  = \new_[46223]_  & \new_[46216]_ ;
  assign \new_[46227]_  = A167 & A170;
  assign \new_[46230]_  = ~A201 & ~A166;
  assign \new_[46231]_  = \new_[46230]_  & \new_[46227]_ ;
  assign \new_[46234]_  = ~A203 & ~A202;
  assign \new_[46237]_  = ~A233 & ~A232;
  assign \new_[46238]_  = \new_[46237]_  & \new_[46234]_ ;
  assign \new_[46239]_  = \new_[46238]_  & \new_[46231]_ ;
  assign \new_[46242]_  = ~A267 & ~A235;
  assign \new_[46245]_  = ~A269 & ~A268;
  assign \new_[46246]_  = \new_[46245]_  & \new_[46242]_ ;
  assign \new_[46249]_  = A299 & A298;
  assign \new_[46252]_  = ~A301 & ~A300;
  assign \new_[46253]_  = \new_[46252]_  & \new_[46249]_ ;
  assign \new_[46254]_  = \new_[46253]_  & \new_[46246]_ ;
  assign \new_[46257]_  = A167 & A170;
  assign \new_[46260]_  = ~A201 & ~A166;
  assign \new_[46261]_  = \new_[46260]_  & \new_[46257]_ ;
  assign \new_[46264]_  = ~A203 & ~A202;
  assign \new_[46267]_  = ~A233 & ~A232;
  assign \new_[46268]_  = \new_[46267]_  & \new_[46264]_ ;
  assign \new_[46269]_  = \new_[46268]_  & \new_[46261]_ ;
  assign \new_[46272]_  = A265 & ~A235;
  assign \new_[46275]_  = ~A267 & A266;
  assign \new_[46276]_  = \new_[46275]_  & \new_[46272]_ ;
  assign \new_[46279]_  = ~A300 & ~A268;
  assign \new_[46282]_  = ~A302 & ~A301;
  assign \new_[46283]_  = \new_[46282]_  & \new_[46279]_ ;
  assign \new_[46284]_  = \new_[46283]_  & \new_[46276]_ ;
  assign \new_[46287]_  = A167 & A170;
  assign \new_[46290]_  = ~A201 & ~A166;
  assign \new_[46291]_  = \new_[46290]_  & \new_[46287]_ ;
  assign \new_[46294]_  = ~A203 & ~A202;
  assign \new_[46297]_  = ~A233 & ~A232;
  assign \new_[46298]_  = \new_[46297]_  & \new_[46294]_ ;
  assign \new_[46299]_  = \new_[46298]_  & \new_[46291]_ ;
  assign \new_[46302]_  = A265 & ~A235;
  assign \new_[46305]_  = ~A267 & A266;
  assign \new_[46306]_  = \new_[46305]_  & \new_[46302]_ ;
  assign \new_[46309]_  = ~A298 & ~A268;
  assign \new_[46312]_  = ~A301 & ~A299;
  assign \new_[46313]_  = \new_[46312]_  & \new_[46309]_ ;
  assign \new_[46314]_  = \new_[46313]_  & \new_[46306]_ ;
  assign \new_[46317]_  = A167 & A170;
  assign \new_[46320]_  = ~A201 & ~A166;
  assign \new_[46321]_  = \new_[46320]_  & \new_[46317]_ ;
  assign \new_[46324]_  = ~A203 & ~A202;
  assign \new_[46327]_  = ~A233 & ~A232;
  assign \new_[46328]_  = \new_[46327]_  & \new_[46324]_ ;
  assign \new_[46329]_  = \new_[46328]_  & \new_[46321]_ ;
  assign \new_[46332]_  = ~A265 & ~A235;
  assign \new_[46335]_  = ~A268 & ~A266;
  assign \new_[46336]_  = \new_[46335]_  & \new_[46332]_ ;
  assign \new_[46339]_  = A299 & A298;
  assign \new_[46342]_  = ~A301 & ~A300;
  assign \new_[46343]_  = \new_[46342]_  & \new_[46339]_ ;
  assign \new_[46344]_  = \new_[46343]_  & \new_[46336]_ ;
  assign \new_[46347]_  = A167 & A170;
  assign \new_[46350]_  = A199 & ~A166;
  assign \new_[46351]_  = \new_[46350]_  & \new_[46347]_ ;
  assign \new_[46354]_  = ~A201 & A200;
  assign \new_[46357]_  = ~A234 & ~A202;
  assign \new_[46358]_  = \new_[46357]_  & \new_[46354]_ ;
  assign \new_[46359]_  = \new_[46358]_  & \new_[46351]_ ;
  assign \new_[46362]_  = ~A236 & ~A235;
  assign \new_[46365]_  = ~A268 & ~A267;
  assign \new_[46366]_  = \new_[46365]_  & \new_[46362]_ ;
  assign \new_[46369]_  = ~A300 & ~A269;
  assign \new_[46372]_  = ~A302 & ~A301;
  assign \new_[46373]_  = \new_[46372]_  & \new_[46369]_ ;
  assign \new_[46374]_  = \new_[46373]_  & \new_[46366]_ ;
  assign \new_[46377]_  = A167 & A170;
  assign \new_[46380]_  = A199 & ~A166;
  assign \new_[46381]_  = \new_[46380]_  & \new_[46377]_ ;
  assign \new_[46384]_  = ~A201 & A200;
  assign \new_[46387]_  = ~A234 & ~A202;
  assign \new_[46388]_  = \new_[46387]_  & \new_[46384]_ ;
  assign \new_[46389]_  = \new_[46388]_  & \new_[46381]_ ;
  assign \new_[46392]_  = ~A236 & ~A235;
  assign \new_[46395]_  = ~A268 & ~A267;
  assign \new_[46396]_  = \new_[46395]_  & \new_[46392]_ ;
  assign \new_[46399]_  = ~A298 & ~A269;
  assign \new_[46402]_  = ~A301 & ~A299;
  assign \new_[46403]_  = \new_[46402]_  & \new_[46399]_ ;
  assign \new_[46404]_  = \new_[46403]_  & \new_[46396]_ ;
  assign \new_[46407]_  = A167 & A170;
  assign \new_[46410]_  = A199 & ~A166;
  assign \new_[46411]_  = \new_[46410]_  & \new_[46407]_ ;
  assign \new_[46414]_  = ~A201 & A200;
  assign \new_[46417]_  = ~A234 & ~A202;
  assign \new_[46418]_  = \new_[46417]_  & \new_[46414]_ ;
  assign \new_[46419]_  = \new_[46418]_  & \new_[46411]_ ;
  assign \new_[46422]_  = ~A236 & ~A235;
  assign \new_[46425]_  = ~A266 & ~A265;
  assign \new_[46426]_  = \new_[46425]_  & \new_[46422]_ ;
  assign \new_[46429]_  = ~A300 & ~A268;
  assign \new_[46432]_  = ~A302 & ~A301;
  assign \new_[46433]_  = \new_[46432]_  & \new_[46429]_ ;
  assign \new_[46434]_  = \new_[46433]_  & \new_[46426]_ ;
  assign \new_[46437]_  = A167 & A170;
  assign \new_[46440]_  = A199 & ~A166;
  assign \new_[46441]_  = \new_[46440]_  & \new_[46437]_ ;
  assign \new_[46444]_  = ~A201 & A200;
  assign \new_[46447]_  = ~A234 & ~A202;
  assign \new_[46448]_  = \new_[46447]_  & \new_[46444]_ ;
  assign \new_[46449]_  = \new_[46448]_  & \new_[46441]_ ;
  assign \new_[46452]_  = ~A236 & ~A235;
  assign \new_[46455]_  = ~A266 & ~A265;
  assign \new_[46456]_  = \new_[46455]_  & \new_[46452]_ ;
  assign \new_[46459]_  = ~A298 & ~A268;
  assign \new_[46462]_  = ~A301 & ~A299;
  assign \new_[46463]_  = \new_[46462]_  & \new_[46459]_ ;
  assign \new_[46464]_  = \new_[46463]_  & \new_[46456]_ ;
  assign \new_[46467]_  = A167 & A170;
  assign \new_[46470]_  = A199 & ~A166;
  assign \new_[46471]_  = \new_[46470]_  & \new_[46467]_ ;
  assign \new_[46474]_  = ~A201 & A200;
  assign \new_[46477]_  = ~A232 & ~A202;
  assign \new_[46478]_  = \new_[46477]_  & \new_[46474]_ ;
  assign \new_[46479]_  = \new_[46478]_  & \new_[46471]_ ;
  assign \new_[46482]_  = ~A235 & ~A233;
  assign \new_[46485]_  = ~A268 & ~A267;
  assign \new_[46486]_  = \new_[46485]_  & \new_[46482]_ ;
  assign \new_[46489]_  = ~A300 & ~A269;
  assign \new_[46492]_  = ~A302 & ~A301;
  assign \new_[46493]_  = \new_[46492]_  & \new_[46489]_ ;
  assign \new_[46494]_  = \new_[46493]_  & \new_[46486]_ ;
  assign \new_[46497]_  = A167 & A170;
  assign \new_[46500]_  = A199 & ~A166;
  assign \new_[46501]_  = \new_[46500]_  & \new_[46497]_ ;
  assign \new_[46504]_  = ~A201 & A200;
  assign \new_[46507]_  = ~A232 & ~A202;
  assign \new_[46508]_  = \new_[46507]_  & \new_[46504]_ ;
  assign \new_[46509]_  = \new_[46508]_  & \new_[46501]_ ;
  assign \new_[46512]_  = ~A235 & ~A233;
  assign \new_[46515]_  = ~A268 & ~A267;
  assign \new_[46516]_  = \new_[46515]_  & \new_[46512]_ ;
  assign \new_[46519]_  = ~A298 & ~A269;
  assign \new_[46522]_  = ~A301 & ~A299;
  assign \new_[46523]_  = \new_[46522]_  & \new_[46519]_ ;
  assign \new_[46524]_  = \new_[46523]_  & \new_[46516]_ ;
  assign \new_[46527]_  = A167 & A170;
  assign \new_[46530]_  = A199 & ~A166;
  assign \new_[46531]_  = \new_[46530]_  & \new_[46527]_ ;
  assign \new_[46534]_  = ~A201 & A200;
  assign \new_[46537]_  = ~A232 & ~A202;
  assign \new_[46538]_  = \new_[46537]_  & \new_[46534]_ ;
  assign \new_[46539]_  = \new_[46538]_  & \new_[46531]_ ;
  assign \new_[46542]_  = ~A235 & ~A233;
  assign \new_[46545]_  = ~A266 & ~A265;
  assign \new_[46546]_  = \new_[46545]_  & \new_[46542]_ ;
  assign \new_[46549]_  = ~A300 & ~A268;
  assign \new_[46552]_  = ~A302 & ~A301;
  assign \new_[46553]_  = \new_[46552]_  & \new_[46549]_ ;
  assign \new_[46554]_  = \new_[46553]_  & \new_[46546]_ ;
  assign \new_[46557]_  = A167 & A170;
  assign \new_[46560]_  = A199 & ~A166;
  assign \new_[46561]_  = \new_[46560]_  & \new_[46557]_ ;
  assign \new_[46564]_  = ~A201 & A200;
  assign \new_[46567]_  = ~A232 & ~A202;
  assign \new_[46568]_  = \new_[46567]_  & \new_[46564]_ ;
  assign \new_[46569]_  = \new_[46568]_  & \new_[46561]_ ;
  assign \new_[46572]_  = ~A235 & ~A233;
  assign \new_[46575]_  = ~A266 & ~A265;
  assign \new_[46576]_  = \new_[46575]_  & \new_[46572]_ ;
  assign \new_[46579]_  = ~A298 & ~A268;
  assign \new_[46582]_  = ~A301 & ~A299;
  assign \new_[46583]_  = \new_[46582]_  & \new_[46579]_ ;
  assign \new_[46584]_  = \new_[46583]_  & \new_[46576]_ ;
  assign \new_[46587]_  = A167 & A170;
  assign \new_[46590]_  = ~A199 & ~A166;
  assign \new_[46591]_  = \new_[46590]_  & \new_[46587]_ ;
  assign \new_[46594]_  = ~A202 & ~A200;
  assign \new_[46597]_  = ~A235 & ~A234;
  assign \new_[46598]_  = \new_[46597]_  & \new_[46594]_ ;
  assign \new_[46599]_  = \new_[46598]_  & \new_[46591]_ ;
  assign \new_[46602]_  = ~A267 & ~A236;
  assign \new_[46605]_  = ~A269 & ~A268;
  assign \new_[46606]_  = \new_[46605]_  & \new_[46602]_ ;
  assign \new_[46609]_  = A299 & A298;
  assign \new_[46612]_  = ~A301 & ~A300;
  assign \new_[46613]_  = \new_[46612]_  & \new_[46609]_ ;
  assign \new_[46614]_  = \new_[46613]_  & \new_[46606]_ ;
  assign \new_[46617]_  = A167 & A170;
  assign \new_[46620]_  = ~A199 & ~A166;
  assign \new_[46621]_  = \new_[46620]_  & \new_[46617]_ ;
  assign \new_[46624]_  = ~A202 & ~A200;
  assign \new_[46627]_  = ~A235 & ~A234;
  assign \new_[46628]_  = \new_[46627]_  & \new_[46624]_ ;
  assign \new_[46629]_  = \new_[46628]_  & \new_[46621]_ ;
  assign \new_[46632]_  = A265 & ~A236;
  assign \new_[46635]_  = ~A267 & A266;
  assign \new_[46636]_  = \new_[46635]_  & \new_[46632]_ ;
  assign \new_[46639]_  = ~A300 & ~A268;
  assign \new_[46642]_  = ~A302 & ~A301;
  assign \new_[46643]_  = \new_[46642]_  & \new_[46639]_ ;
  assign \new_[46644]_  = \new_[46643]_  & \new_[46636]_ ;
  assign \new_[46647]_  = A167 & A170;
  assign \new_[46650]_  = ~A199 & ~A166;
  assign \new_[46651]_  = \new_[46650]_  & \new_[46647]_ ;
  assign \new_[46654]_  = ~A202 & ~A200;
  assign \new_[46657]_  = ~A235 & ~A234;
  assign \new_[46658]_  = \new_[46657]_  & \new_[46654]_ ;
  assign \new_[46659]_  = \new_[46658]_  & \new_[46651]_ ;
  assign \new_[46662]_  = A265 & ~A236;
  assign \new_[46665]_  = ~A267 & A266;
  assign \new_[46666]_  = \new_[46665]_  & \new_[46662]_ ;
  assign \new_[46669]_  = ~A298 & ~A268;
  assign \new_[46672]_  = ~A301 & ~A299;
  assign \new_[46673]_  = \new_[46672]_  & \new_[46669]_ ;
  assign \new_[46674]_  = \new_[46673]_  & \new_[46666]_ ;
  assign \new_[46677]_  = A167 & A170;
  assign \new_[46680]_  = ~A199 & ~A166;
  assign \new_[46681]_  = \new_[46680]_  & \new_[46677]_ ;
  assign \new_[46684]_  = ~A202 & ~A200;
  assign \new_[46687]_  = ~A235 & ~A234;
  assign \new_[46688]_  = \new_[46687]_  & \new_[46684]_ ;
  assign \new_[46689]_  = \new_[46688]_  & \new_[46681]_ ;
  assign \new_[46692]_  = ~A265 & ~A236;
  assign \new_[46695]_  = ~A268 & ~A266;
  assign \new_[46696]_  = \new_[46695]_  & \new_[46692]_ ;
  assign \new_[46699]_  = A299 & A298;
  assign \new_[46702]_  = ~A301 & ~A300;
  assign \new_[46703]_  = \new_[46702]_  & \new_[46699]_ ;
  assign \new_[46704]_  = \new_[46703]_  & \new_[46696]_ ;
  assign \new_[46707]_  = A167 & A170;
  assign \new_[46710]_  = ~A199 & ~A166;
  assign \new_[46711]_  = \new_[46710]_  & \new_[46707]_ ;
  assign \new_[46714]_  = ~A202 & ~A200;
  assign \new_[46717]_  = A233 & A232;
  assign \new_[46718]_  = \new_[46717]_  & \new_[46714]_ ;
  assign \new_[46719]_  = \new_[46718]_  & \new_[46711]_ ;
  assign \new_[46722]_  = ~A235 & ~A234;
  assign \new_[46725]_  = ~A268 & ~A267;
  assign \new_[46726]_  = \new_[46725]_  & \new_[46722]_ ;
  assign \new_[46729]_  = ~A300 & ~A269;
  assign \new_[46732]_  = ~A302 & ~A301;
  assign \new_[46733]_  = \new_[46732]_  & \new_[46729]_ ;
  assign \new_[46734]_  = \new_[46733]_  & \new_[46726]_ ;
  assign \new_[46737]_  = A167 & A170;
  assign \new_[46740]_  = ~A199 & ~A166;
  assign \new_[46741]_  = \new_[46740]_  & \new_[46737]_ ;
  assign \new_[46744]_  = ~A202 & ~A200;
  assign \new_[46747]_  = A233 & A232;
  assign \new_[46748]_  = \new_[46747]_  & \new_[46744]_ ;
  assign \new_[46749]_  = \new_[46748]_  & \new_[46741]_ ;
  assign \new_[46752]_  = ~A235 & ~A234;
  assign \new_[46755]_  = ~A268 & ~A267;
  assign \new_[46756]_  = \new_[46755]_  & \new_[46752]_ ;
  assign \new_[46759]_  = ~A298 & ~A269;
  assign \new_[46762]_  = ~A301 & ~A299;
  assign \new_[46763]_  = \new_[46762]_  & \new_[46759]_ ;
  assign \new_[46764]_  = \new_[46763]_  & \new_[46756]_ ;
  assign \new_[46767]_  = A167 & A170;
  assign \new_[46770]_  = ~A199 & ~A166;
  assign \new_[46771]_  = \new_[46770]_  & \new_[46767]_ ;
  assign \new_[46774]_  = ~A202 & ~A200;
  assign \new_[46777]_  = A233 & A232;
  assign \new_[46778]_  = \new_[46777]_  & \new_[46774]_ ;
  assign \new_[46779]_  = \new_[46778]_  & \new_[46771]_ ;
  assign \new_[46782]_  = ~A235 & ~A234;
  assign \new_[46785]_  = ~A266 & ~A265;
  assign \new_[46786]_  = \new_[46785]_  & \new_[46782]_ ;
  assign \new_[46789]_  = ~A300 & ~A268;
  assign \new_[46792]_  = ~A302 & ~A301;
  assign \new_[46793]_  = \new_[46792]_  & \new_[46789]_ ;
  assign \new_[46794]_  = \new_[46793]_  & \new_[46786]_ ;
  assign \new_[46797]_  = A167 & A170;
  assign \new_[46800]_  = ~A199 & ~A166;
  assign \new_[46801]_  = \new_[46800]_  & \new_[46797]_ ;
  assign \new_[46804]_  = ~A202 & ~A200;
  assign \new_[46807]_  = A233 & A232;
  assign \new_[46808]_  = \new_[46807]_  & \new_[46804]_ ;
  assign \new_[46809]_  = \new_[46808]_  & \new_[46801]_ ;
  assign \new_[46812]_  = ~A235 & ~A234;
  assign \new_[46815]_  = ~A266 & ~A265;
  assign \new_[46816]_  = \new_[46815]_  & \new_[46812]_ ;
  assign \new_[46819]_  = ~A298 & ~A268;
  assign \new_[46822]_  = ~A301 & ~A299;
  assign \new_[46823]_  = \new_[46822]_  & \new_[46819]_ ;
  assign \new_[46824]_  = \new_[46823]_  & \new_[46816]_ ;
  assign \new_[46827]_  = A167 & A170;
  assign \new_[46830]_  = ~A199 & ~A166;
  assign \new_[46831]_  = \new_[46830]_  & \new_[46827]_ ;
  assign \new_[46834]_  = ~A202 & ~A200;
  assign \new_[46837]_  = ~A233 & ~A232;
  assign \new_[46838]_  = \new_[46837]_  & \new_[46834]_ ;
  assign \new_[46839]_  = \new_[46838]_  & \new_[46831]_ ;
  assign \new_[46842]_  = ~A267 & ~A235;
  assign \new_[46845]_  = ~A269 & ~A268;
  assign \new_[46846]_  = \new_[46845]_  & \new_[46842]_ ;
  assign \new_[46849]_  = A299 & A298;
  assign \new_[46852]_  = ~A301 & ~A300;
  assign \new_[46853]_  = \new_[46852]_  & \new_[46849]_ ;
  assign \new_[46854]_  = \new_[46853]_  & \new_[46846]_ ;
  assign \new_[46857]_  = A167 & A170;
  assign \new_[46860]_  = ~A199 & ~A166;
  assign \new_[46861]_  = \new_[46860]_  & \new_[46857]_ ;
  assign \new_[46864]_  = ~A202 & ~A200;
  assign \new_[46867]_  = ~A233 & ~A232;
  assign \new_[46868]_  = \new_[46867]_  & \new_[46864]_ ;
  assign \new_[46869]_  = \new_[46868]_  & \new_[46861]_ ;
  assign \new_[46872]_  = A265 & ~A235;
  assign \new_[46875]_  = ~A267 & A266;
  assign \new_[46876]_  = \new_[46875]_  & \new_[46872]_ ;
  assign \new_[46879]_  = ~A300 & ~A268;
  assign \new_[46882]_  = ~A302 & ~A301;
  assign \new_[46883]_  = \new_[46882]_  & \new_[46879]_ ;
  assign \new_[46884]_  = \new_[46883]_  & \new_[46876]_ ;
  assign \new_[46887]_  = A167 & A170;
  assign \new_[46890]_  = ~A199 & ~A166;
  assign \new_[46891]_  = \new_[46890]_  & \new_[46887]_ ;
  assign \new_[46894]_  = ~A202 & ~A200;
  assign \new_[46897]_  = ~A233 & ~A232;
  assign \new_[46898]_  = \new_[46897]_  & \new_[46894]_ ;
  assign \new_[46899]_  = \new_[46898]_  & \new_[46891]_ ;
  assign \new_[46902]_  = A265 & ~A235;
  assign \new_[46905]_  = ~A267 & A266;
  assign \new_[46906]_  = \new_[46905]_  & \new_[46902]_ ;
  assign \new_[46909]_  = ~A298 & ~A268;
  assign \new_[46912]_  = ~A301 & ~A299;
  assign \new_[46913]_  = \new_[46912]_  & \new_[46909]_ ;
  assign \new_[46914]_  = \new_[46913]_  & \new_[46906]_ ;
  assign \new_[46917]_  = A167 & A170;
  assign \new_[46920]_  = ~A199 & ~A166;
  assign \new_[46921]_  = \new_[46920]_  & \new_[46917]_ ;
  assign \new_[46924]_  = ~A202 & ~A200;
  assign \new_[46927]_  = ~A233 & ~A232;
  assign \new_[46928]_  = \new_[46927]_  & \new_[46924]_ ;
  assign \new_[46929]_  = \new_[46928]_  & \new_[46921]_ ;
  assign \new_[46932]_  = ~A265 & ~A235;
  assign \new_[46935]_  = ~A268 & ~A266;
  assign \new_[46936]_  = \new_[46935]_  & \new_[46932]_ ;
  assign \new_[46939]_  = A299 & A298;
  assign \new_[46942]_  = ~A301 & ~A300;
  assign \new_[46943]_  = \new_[46942]_  & \new_[46939]_ ;
  assign \new_[46944]_  = \new_[46943]_  & \new_[46936]_ ;
  assign \new_[46947]_  = ~A167 & A170;
  assign \new_[46950]_  = ~A201 & A166;
  assign \new_[46951]_  = \new_[46950]_  & \new_[46947]_ ;
  assign \new_[46954]_  = ~A203 & ~A202;
  assign \new_[46957]_  = ~A235 & ~A234;
  assign \new_[46958]_  = \new_[46957]_  & \new_[46954]_ ;
  assign \new_[46959]_  = \new_[46958]_  & \new_[46951]_ ;
  assign \new_[46962]_  = ~A267 & ~A236;
  assign \new_[46965]_  = ~A269 & ~A268;
  assign \new_[46966]_  = \new_[46965]_  & \new_[46962]_ ;
  assign \new_[46969]_  = A299 & A298;
  assign \new_[46972]_  = ~A301 & ~A300;
  assign \new_[46973]_  = \new_[46972]_  & \new_[46969]_ ;
  assign \new_[46974]_  = \new_[46973]_  & \new_[46966]_ ;
  assign \new_[46977]_  = ~A167 & A170;
  assign \new_[46980]_  = ~A201 & A166;
  assign \new_[46981]_  = \new_[46980]_  & \new_[46977]_ ;
  assign \new_[46984]_  = ~A203 & ~A202;
  assign \new_[46987]_  = ~A235 & ~A234;
  assign \new_[46988]_  = \new_[46987]_  & \new_[46984]_ ;
  assign \new_[46989]_  = \new_[46988]_  & \new_[46981]_ ;
  assign \new_[46992]_  = A265 & ~A236;
  assign \new_[46995]_  = ~A267 & A266;
  assign \new_[46996]_  = \new_[46995]_  & \new_[46992]_ ;
  assign \new_[46999]_  = ~A300 & ~A268;
  assign \new_[47002]_  = ~A302 & ~A301;
  assign \new_[47003]_  = \new_[47002]_  & \new_[46999]_ ;
  assign \new_[47004]_  = \new_[47003]_  & \new_[46996]_ ;
  assign \new_[47007]_  = ~A167 & A170;
  assign \new_[47010]_  = ~A201 & A166;
  assign \new_[47011]_  = \new_[47010]_  & \new_[47007]_ ;
  assign \new_[47014]_  = ~A203 & ~A202;
  assign \new_[47017]_  = ~A235 & ~A234;
  assign \new_[47018]_  = \new_[47017]_  & \new_[47014]_ ;
  assign \new_[47019]_  = \new_[47018]_  & \new_[47011]_ ;
  assign \new_[47022]_  = A265 & ~A236;
  assign \new_[47025]_  = ~A267 & A266;
  assign \new_[47026]_  = \new_[47025]_  & \new_[47022]_ ;
  assign \new_[47029]_  = ~A298 & ~A268;
  assign \new_[47032]_  = ~A301 & ~A299;
  assign \new_[47033]_  = \new_[47032]_  & \new_[47029]_ ;
  assign \new_[47034]_  = \new_[47033]_  & \new_[47026]_ ;
  assign \new_[47037]_  = ~A167 & A170;
  assign \new_[47040]_  = ~A201 & A166;
  assign \new_[47041]_  = \new_[47040]_  & \new_[47037]_ ;
  assign \new_[47044]_  = ~A203 & ~A202;
  assign \new_[47047]_  = ~A235 & ~A234;
  assign \new_[47048]_  = \new_[47047]_  & \new_[47044]_ ;
  assign \new_[47049]_  = \new_[47048]_  & \new_[47041]_ ;
  assign \new_[47052]_  = ~A265 & ~A236;
  assign \new_[47055]_  = ~A268 & ~A266;
  assign \new_[47056]_  = \new_[47055]_  & \new_[47052]_ ;
  assign \new_[47059]_  = A299 & A298;
  assign \new_[47062]_  = ~A301 & ~A300;
  assign \new_[47063]_  = \new_[47062]_  & \new_[47059]_ ;
  assign \new_[47064]_  = \new_[47063]_  & \new_[47056]_ ;
  assign \new_[47067]_  = ~A167 & A170;
  assign \new_[47070]_  = ~A201 & A166;
  assign \new_[47071]_  = \new_[47070]_  & \new_[47067]_ ;
  assign \new_[47074]_  = ~A203 & ~A202;
  assign \new_[47077]_  = A233 & A232;
  assign \new_[47078]_  = \new_[47077]_  & \new_[47074]_ ;
  assign \new_[47079]_  = \new_[47078]_  & \new_[47071]_ ;
  assign \new_[47082]_  = ~A235 & ~A234;
  assign \new_[47085]_  = ~A268 & ~A267;
  assign \new_[47086]_  = \new_[47085]_  & \new_[47082]_ ;
  assign \new_[47089]_  = ~A300 & ~A269;
  assign \new_[47092]_  = ~A302 & ~A301;
  assign \new_[47093]_  = \new_[47092]_  & \new_[47089]_ ;
  assign \new_[47094]_  = \new_[47093]_  & \new_[47086]_ ;
  assign \new_[47097]_  = ~A167 & A170;
  assign \new_[47100]_  = ~A201 & A166;
  assign \new_[47101]_  = \new_[47100]_  & \new_[47097]_ ;
  assign \new_[47104]_  = ~A203 & ~A202;
  assign \new_[47107]_  = A233 & A232;
  assign \new_[47108]_  = \new_[47107]_  & \new_[47104]_ ;
  assign \new_[47109]_  = \new_[47108]_  & \new_[47101]_ ;
  assign \new_[47112]_  = ~A235 & ~A234;
  assign \new_[47115]_  = ~A268 & ~A267;
  assign \new_[47116]_  = \new_[47115]_  & \new_[47112]_ ;
  assign \new_[47119]_  = ~A298 & ~A269;
  assign \new_[47122]_  = ~A301 & ~A299;
  assign \new_[47123]_  = \new_[47122]_  & \new_[47119]_ ;
  assign \new_[47124]_  = \new_[47123]_  & \new_[47116]_ ;
  assign \new_[47127]_  = ~A167 & A170;
  assign \new_[47130]_  = ~A201 & A166;
  assign \new_[47131]_  = \new_[47130]_  & \new_[47127]_ ;
  assign \new_[47134]_  = ~A203 & ~A202;
  assign \new_[47137]_  = A233 & A232;
  assign \new_[47138]_  = \new_[47137]_  & \new_[47134]_ ;
  assign \new_[47139]_  = \new_[47138]_  & \new_[47131]_ ;
  assign \new_[47142]_  = ~A235 & ~A234;
  assign \new_[47145]_  = ~A266 & ~A265;
  assign \new_[47146]_  = \new_[47145]_  & \new_[47142]_ ;
  assign \new_[47149]_  = ~A300 & ~A268;
  assign \new_[47152]_  = ~A302 & ~A301;
  assign \new_[47153]_  = \new_[47152]_  & \new_[47149]_ ;
  assign \new_[47154]_  = \new_[47153]_  & \new_[47146]_ ;
  assign \new_[47157]_  = ~A167 & A170;
  assign \new_[47160]_  = ~A201 & A166;
  assign \new_[47161]_  = \new_[47160]_  & \new_[47157]_ ;
  assign \new_[47164]_  = ~A203 & ~A202;
  assign \new_[47167]_  = A233 & A232;
  assign \new_[47168]_  = \new_[47167]_  & \new_[47164]_ ;
  assign \new_[47169]_  = \new_[47168]_  & \new_[47161]_ ;
  assign \new_[47172]_  = ~A235 & ~A234;
  assign \new_[47175]_  = ~A266 & ~A265;
  assign \new_[47176]_  = \new_[47175]_  & \new_[47172]_ ;
  assign \new_[47179]_  = ~A298 & ~A268;
  assign \new_[47182]_  = ~A301 & ~A299;
  assign \new_[47183]_  = \new_[47182]_  & \new_[47179]_ ;
  assign \new_[47184]_  = \new_[47183]_  & \new_[47176]_ ;
  assign \new_[47187]_  = ~A167 & A170;
  assign \new_[47190]_  = ~A201 & A166;
  assign \new_[47191]_  = \new_[47190]_  & \new_[47187]_ ;
  assign \new_[47194]_  = ~A203 & ~A202;
  assign \new_[47197]_  = ~A233 & ~A232;
  assign \new_[47198]_  = \new_[47197]_  & \new_[47194]_ ;
  assign \new_[47199]_  = \new_[47198]_  & \new_[47191]_ ;
  assign \new_[47202]_  = ~A267 & ~A235;
  assign \new_[47205]_  = ~A269 & ~A268;
  assign \new_[47206]_  = \new_[47205]_  & \new_[47202]_ ;
  assign \new_[47209]_  = A299 & A298;
  assign \new_[47212]_  = ~A301 & ~A300;
  assign \new_[47213]_  = \new_[47212]_  & \new_[47209]_ ;
  assign \new_[47214]_  = \new_[47213]_  & \new_[47206]_ ;
  assign \new_[47217]_  = ~A167 & A170;
  assign \new_[47220]_  = ~A201 & A166;
  assign \new_[47221]_  = \new_[47220]_  & \new_[47217]_ ;
  assign \new_[47224]_  = ~A203 & ~A202;
  assign \new_[47227]_  = ~A233 & ~A232;
  assign \new_[47228]_  = \new_[47227]_  & \new_[47224]_ ;
  assign \new_[47229]_  = \new_[47228]_  & \new_[47221]_ ;
  assign \new_[47232]_  = A265 & ~A235;
  assign \new_[47235]_  = ~A267 & A266;
  assign \new_[47236]_  = \new_[47235]_  & \new_[47232]_ ;
  assign \new_[47239]_  = ~A300 & ~A268;
  assign \new_[47242]_  = ~A302 & ~A301;
  assign \new_[47243]_  = \new_[47242]_  & \new_[47239]_ ;
  assign \new_[47244]_  = \new_[47243]_  & \new_[47236]_ ;
  assign \new_[47247]_  = ~A167 & A170;
  assign \new_[47250]_  = ~A201 & A166;
  assign \new_[47251]_  = \new_[47250]_  & \new_[47247]_ ;
  assign \new_[47254]_  = ~A203 & ~A202;
  assign \new_[47257]_  = ~A233 & ~A232;
  assign \new_[47258]_  = \new_[47257]_  & \new_[47254]_ ;
  assign \new_[47259]_  = \new_[47258]_  & \new_[47251]_ ;
  assign \new_[47262]_  = A265 & ~A235;
  assign \new_[47265]_  = ~A267 & A266;
  assign \new_[47266]_  = \new_[47265]_  & \new_[47262]_ ;
  assign \new_[47269]_  = ~A298 & ~A268;
  assign \new_[47272]_  = ~A301 & ~A299;
  assign \new_[47273]_  = \new_[47272]_  & \new_[47269]_ ;
  assign \new_[47274]_  = \new_[47273]_  & \new_[47266]_ ;
  assign \new_[47277]_  = ~A167 & A170;
  assign \new_[47280]_  = ~A201 & A166;
  assign \new_[47281]_  = \new_[47280]_  & \new_[47277]_ ;
  assign \new_[47284]_  = ~A203 & ~A202;
  assign \new_[47287]_  = ~A233 & ~A232;
  assign \new_[47288]_  = \new_[47287]_  & \new_[47284]_ ;
  assign \new_[47289]_  = \new_[47288]_  & \new_[47281]_ ;
  assign \new_[47292]_  = ~A265 & ~A235;
  assign \new_[47295]_  = ~A268 & ~A266;
  assign \new_[47296]_  = \new_[47295]_  & \new_[47292]_ ;
  assign \new_[47299]_  = A299 & A298;
  assign \new_[47302]_  = ~A301 & ~A300;
  assign \new_[47303]_  = \new_[47302]_  & \new_[47299]_ ;
  assign \new_[47304]_  = \new_[47303]_  & \new_[47296]_ ;
  assign \new_[47307]_  = ~A167 & A170;
  assign \new_[47310]_  = A199 & A166;
  assign \new_[47311]_  = \new_[47310]_  & \new_[47307]_ ;
  assign \new_[47314]_  = ~A201 & A200;
  assign \new_[47317]_  = ~A234 & ~A202;
  assign \new_[47318]_  = \new_[47317]_  & \new_[47314]_ ;
  assign \new_[47319]_  = \new_[47318]_  & \new_[47311]_ ;
  assign \new_[47322]_  = ~A236 & ~A235;
  assign \new_[47325]_  = ~A268 & ~A267;
  assign \new_[47326]_  = \new_[47325]_  & \new_[47322]_ ;
  assign \new_[47329]_  = ~A300 & ~A269;
  assign \new_[47332]_  = ~A302 & ~A301;
  assign \new_[47333]_  = \new_[47332]_  & \new_[47329]_ ;
  assign \new_[47334]_  = \new_[47333]_  & \new_[47326]_ ;
  assign \new_[47337]_  = ~A167 & A170;
  assign \new_[47340]_  = A199 & A166;
  assign \new_[47341]_  = \new_[47340]_  & \new_[47337]_ ;
  assign \new_[47344]_  = ~A201 & A200;
  assign \new_[47347]_  = ~A234 & ~A202;
  assign \new_[47348]_  = \new_[47347]_  & \new_[47344]_ ;
  assign \new_[47349]_  = \new_[47348]_  & \new_[47341]_ ;
  assign \new_[47352]_  = ~A236 & ~A235;
  assign \new_[47355]_  = ~A268 & ~A267;
  assign \new_[47356]_  = \new_[47355]_  & \new_[47352]_ ;
  assign \new_[47359]_  = ~A298 & ~A269;
  assign \new_[47362]_  = ~A301 & ~A299;
  assign \new_[47363]_  = \new_[47362]_  & \new_[47359]_ ;
  assign \new_[47364]_  = \new_[47363]_  & \new_[47356]_ ;
  assign \new_[47367]_  = ~A167 & A170;
  assign \new_[47370]_  = A199 & A166;
  assign \new_[47371]_  = \new_[47370]_  & \new_[47367]_ ;
  assign \new_[47374]_  = ~A201 & A200;
  assign \new_[47377]_  = ~A234 & ~A202;
  assign \new_[47378]_  = \new_[47377]_  & \new_[47374]_ ;
  assign \new_[47379]_  = \new_[47378]_  & \new_[47371]_ ;
  assign \new_[47382]_  = ~A236 & ~A235;
  assign \new_[47385]_  = ~A266 & ~A265;
  assign \new_[47386]_  = \new_[47385]_  & \new_[47382]_ ;
  assign \new_[47389]_  = ~A300 & ~A268;
  assign \new_[47392]_  = ~A302 & ~A301;
  assign \new_[47393]_  = \new_[47392]_  & \new_[47389]_ ;
  assign \new_[47394]_  = \new_[47393]_  & \new_[47386]_ ;
  assign \new_[47397]_  = ~A167 & A170;
  assign \new_[47400]_  = A199 & A166;
  assign \new_[47401]_  = \new_[47400]_  & \new_[47397]_ ;
  assign \new_[47404]_  = ~A201 & A200;
  assign \new_[47407]_  = ~A234 & ~A202;
  assign \new_[47408]_  = \new_[47407]_  & \new_[47404]_ ;
  assign \new_[47409]_  = \new_[47408]_  & \new_[47401]_ ;
  assign \new_[47412]_  = ~A236 & ~A235;
  assign \new_[47415]_  = ~A266 & ~A265;
  assign \new_[47416]_  = \new_[47415]_  & \new_[47412]_ ;
  assign \new_[47419]_  = ~A298 & ~A268;
  assign \new_[47422]_  = ~A301 & ~A299;
  assign \new_[47423]_  = \new_[47422]_  & \new_[47419]_ ;
  assign \new_[47424]_  = \new_[47423]_  & \new_[47416]_ ;
  assign \new_[47427]_  = ~A167 & A170;
  assign \new_[47430]_  = A199 & A166;
  assign \new_[47431]_  = \new_[47430]_  & \new_[47427]_ ;
  assign \new_[47434]_  = ~A201 & A200;
  assign \new_[47437]_  = ~A232 & ~A202;
  assign \new_[47438]_  = \new_[47437]_  & \new_[47434]_ ;
  assign \new_[47439]_  = \new_[47438]_  & \new_[47431]_ ;
  assign \new_[47442]_  = ~A235 & ~A233;
  assign \new_[47445]_  = ~A268 & ~A267;
  assign \new_[47446]_  = \new_[47445]_  & \new_[47442]_ ;
  assign \new_[47449]_  = ~A300 & ~A269;
  assign \new_[47452]_  = ~A302 & ~A301;
  assign \new_[47453]_  = \new_[47452]_  & \new_[47449]_ ;
  assign \new_[47454]_  = \new_[47453]_  & \new_[47446]_ ;
  assign \new_[47457]_  = ~A167 & A170;
  assign \new_[47460]_  = A199 & A166;
  assign \new_[47461]_  = \new_[47460]_  & \new_[47457]_ ;
  assign \new_[47464]_  = ~A201 & A200;
  assign \new_[47467]_  = ~A232 & ~A202;
  assign \new_[47468]_  = \new_[47467]_  & \new_[47464]_ ;
  assign \new_[47469]_  = \new_[47468]_  & \new_[47461]_ ;
  assign \new_[47472]_  = ~A235 & ~A233;
  assign \new_[47475]_  = ~A268 & ~A267;
  assign \new_[47476]_  = \new_[47475]_  & \new_[47472]_ ;
  assign \new_[47479]_  = ~A298 & ~A269;
  assign \new_[47482]_  = ~A301 & ~A299;
  assign \new_[47483]_  = \new_[47482]_  & \new_[47479]_ ;
  assign \new_[47484]_  = \new_[47483]_  & \new_[47476]_ ;
  assign \new_[47487]_  = ~A167 & A170;
  assign \new_[47490]_  = A199 & A166;
  assign \new_[47491]_  = \new_[47490]_  & \new_[47487]_ ;
  assign \new_[47494]_  = ~A201 & A200;
  assign \new_[47497]_  = ~A232 & ~A202;
  assign \new_[47498]_  = \new_[47497]_  & \new_[47494]_ ;
  assign \new_[47499]_  = \new_[47498]_  & \new_[47491]_ ;
  assign \new_[47502]_  = ~A235 & ~A233;
  assign \new_[47505]_  = ~A266 & ~A265;
  assign \new_[47506]_  = \new_[47505]_  & \new_[47502]_ ;
  assign \new_[47509]_  = ~A300 & ~A268;
  assign \new_[47512]_  = ~A302 & ~A301;
  assign \new_[47513]_  = \new_[47512]_  & \new_[47509]_ ;
  assign \new_[47514]_  = \new_[47513]_  & \new_[47506]_ ;
  assign \new_[47517]_  = ~A167 & A170;
  assign \new_[47520]_  = A199 & A166;
  assign \new_[47521]_  = \new_[47520]_  & \new_[47517]_ ;
  assign \new_[47524]_  = ~A201 & A200;
  assign \new_[47527]_  = ~A232 & ~A202;
  assign \new_[47528]_  = \new_[47527]_  & \new_[47524]_ ;
  assign \new_[47529]_  = \new_[47528]_  & \new_[47521]_ ;
  assign \new_[47532]_  = ~A235 & ~A233;
  assign \new_[47535]_  = ~A266 & ~A265;
  assign \new_[47536]_  = \new_[47535]_  & \new_[47532]_ ;
  assign \new_[47539]_  = ~A298 & ~A268;
  assign \new_[47542]_  = ~A301 & ~A299;
  assign \new_[47543]_  = \new_[47542]_  & \new_[47539]_ ;
  assign \new_[47544]_  = \new_[47543]_  & \new_[47536]_ ;
  assign \new_[47547]_  = ~A167 & A170;
  assign \new_[47550]_  = ~A199 & A166;
  assign \new_[47551]_  = \new_[47550]_  & \new_[47547]_ ;
  assign \new_[47554]_  = ~A202 & ~A200;
  assign \new_[47557]_  = ~A235 & ~A234;
  assign \new_[47558]_  = \new_[47557]_  & \new_[47554]_ ;
  assign \new_[47559]_  = \new_[47558]_  & \new_[47551]_ ;
  assign \new_[47562]_  = ~A267 & ~A236;
  assign \new_[47565]_  = ~A269 & ~A268;
  assign \new_[47566]_  = \new_[47565]_  & \new_[47562]_ ;
  assign \new_[47569]_  = A299 & A298;
  assign \new_[47572]_  = ~A301 & ~A300;
  assign \new_[47573]_  = \new_[47572]_  & \new_[47569]_ ;
  assign \new_[47574]_  = \new_[47573]_  & \new_[47566]_ ;
  assign \new_[47577]_  = ~A167 & A170;
  assign \new_[47580]_  = ~A199 & A166;
  assign \new_[47581]_  = \new_[47580]_  & \new_[47577]_ ;
  assign \new_[47584]_  = ~A202 & ~A200;
  assign \new_[47587]_  = ~A235 & ~A234;
  assign \new_[47588]_  = \new_[47587]_  & \new_[47584]_ ;
  assign \new_[47589]_  = \new_[47588]_  & \new_[47581]_ ;
  assign \new_[47592]_  = A265 & ~A236;
  assign \new_[47595]_  = ~A267 & A266;
  assign \new_[47596]_  = \new_[47595]_  & \new_[47592]_ ;
  assign \new_[47599]_  = ~A300 & ~A268;
  assign \new_[47602]_  = ~A302 & ~A301;
  assign \new_[47603]_  = \new_[47602]_  & \new_[47599]_ ;
  assign \new_[47604]_  = \new_[47603]_  & \new_[47596]_ ;
  assign \new_[47607]_  = ~A167 & A170;
  assign \new_[47610]_  = ~A199 & A166;
  assign \new_[47611]_  = \new_[47610]_  & \new_[47607]_ ;
  assign \new_[47614]_  = ~A202 & ~A200;
  assign \new_[47617]_  = ~A235 & ~A234;
  assign \new_[47618]_  = \new_[47617]_  & \new_[47614]_ ;
  assign \new_[47619]_  = \new_[47618]_  & \new_[47611]_ ;
  assign \new_[47622]_  = A265 & ~A236;
  assign \new_[47625]_  = ~A267 & A266;
  assign \new_[47626]_  = \new_[47625]_  & \new_[47622]_ ;
  assign \new_[47629]_  = ~A298 & ~A268;
  assign \new_[47632]_  = ~A301 & ~A299;
  assign \new_[47633]_  = \new_[47632]_  & \new_[47629]_ ;
  assign \new_[47634]_  = \new_[47633]_  & \new_[47626]_ ;
  assign \new_[47637]_  = ~A167 & A170;
  assign \new_[47640]_  = ~A199 & A166;
  assign \new_[47641]_  = \new_[47640]_  & \new_[47637]_ ;
  assign \new_[47644]_  = ~A202 & ~A200;
  assign \new_[47647]_  = ~A235 & ~A234;
  assign \new_[47648]_  = \new_[47647]_  & \new_[47644]_ ;
  assign \new_[47649]_  = \new_[47648]_  & \new_[47641]_ ;
  assign \new_[47652]_  = ~A265 & ~A236;
  assign \new_[47655]_  = ~A268 & ~A266;
  assign \new_[47656]_  = \new_[47655]_  & \new_[47652]_ ;
  assign \new_[47659]_  = A299 & A298;
  assign \new_[47662]_  = ~A301 & ~A300;
  assign \new_[47663]_  = \new_[47662]_  & \new_[47659]_ ;
  assign \new_[47664]_  = \new_[47663]_  & \new_[47656]_ ;
  assign \new_[47667]_  = ~A167 & A170;
  assign \new_[47670]_  = ~A199 & A166;
  assign \new_[47671]_  = \new_[47670]_  & \new_[47667]_ ;
  assign \new_[47674]_  = ~A202 & ~A200;
  assign \new_[47677]_  = A233 & A232;
  assign \new_[47678]_  = \new_[47677]_  & \new_[47674]_ ;
  assign \new_[47679]_  = \new_[47678]_  & \new_[47671]_ ;
  assign \new_[47682]_  = ~A235 & ~A234;
  assign \new_[47685]_  = ~A268 & ~A267;
  assign \new_[47686]_  = \new_[47685]_  & \new_[47682]_ ;
  assign \new_[47689]_  = ~A300 & ~A269;
  assign \new_[47692]_  = ~A302 & ~A301;
  assign \new_[47693]_  = \new_[47692]_  & \new_[47689]_ ;
  assign \new_[47694]_  = \new_[47693]_  & \new_[47686]_ ;
  assign \new_[47697]_  = ~A167 & A170;
  assign \new_[47700]_  = ~A199 & A166;
  assign \new_[47701]_  = \new_[47700]_  & \new_[47697]_ ;
  assign \new_[47704]_  = ~A202 & ~A200;
  assign \new_[47707]_  = A233 & A232;
  assign \new_[47708]_  = \new_[47707]_  & \new_[47704]_ ;
  assign \new_[47709]_  = \new_[47708]_  & \new_[47701]_ ;
  assign \new_[47712]_  = ~A235 & ~A234;
  assign \new_[47715]_  = ~A268 & ~A267;
  assign \new_[47716]_  = \new_[47715]_  & \new_[47712]_ ;
  assign \new_[47719]_  = ~A298 & ~A269;
  assign \new_[47722]_  = ~A301 & ~A299;
  assign \new_[47723]_  = \new_[47722]_  & \new_[47719]_ ;
  assign \new_[47724]_  = \new_[47723]_  & \new_[47716]_ ;
  assign \new_[47727]_  = ~A167 & A170;
  assign \new_[47730]_  = ~A199 & A166;
  assign \new_[47731]_  = \new_[47730]_  & \new_[47727]_ ;
  assign \new_[47734]_  = ~A202 & ~A200;
  assign \new_[47737]_  = A233 & A232;
  assign \new_[47738]_  = \new_[47737]_  & \new_[47734]_ ;
  assign \new_[47739]_  = \new_[47738]_  & \new_[47731]_ ;
  assign \new_[47742]_  = ~A235 & ~A234;
  assign \new_[47745]_  = ~A266 & ~A265;
  assign \new_[47746]_  = \new_[47745]_  & \new_[47742]_ ;
  assign \new_[47749]_  = ~A300 & ~A268;
  assign \new_[47752]_  = ~A302 & ~A301;
  assign \new_[47753]_  = \new_[47752]_  & \new_[47749]_ ;
  assign \new_[47754]_  = \new_[47753]_  & \new_[47746]_ ;
  assign \new_[47757]_  = ~A167 & A170;
  assign \new_[47760]_  = ~A199 & A166;
  assign \new_[47761]_  = \new_[47760]_  & \new_[47757]_ ;
  assign \new_[47764]_  = ~A202 & ~A200;
  assign \new_[47767]_  = A233 & A232;
  assign \new_[47768]_  = \new_[47767]_  & \new_[47764]_ ;
  assign \new_[47769]_  = \new_[47768]_  & \new_[47761]_ ;
  assign \new_[47772]_  = ~A235 & ~A234;
  assign \new_[47775]_  = ~A266 & ~A265;
  assign \new_[47776]_  = \new_[47775]_  & \new_[47772]_ ;
  assign \new_[47779]_  = ~A298 & ~A268;
  assign \new_[47782]_  = ~A301 & ~A299;
  assign \new_[47783]_  = \new_[47782]_  & \new_[47779]_ ;
  assign \new_[47784]_  = \new_[47783]_  & \new_[47776]_ ;
  assign \new_[47787]_  = ~A167 & A170;
  assign \new_[47790]_  = ~A199 & A166;
  assign \new_[47791]_  = \new_[47790]_  & \new_[47787]_ ;
  assign \new_[47794]_  = ~A202 & ~A200;
  assign \new_[47797]_  = ~A233 & ~A232;
  assign \new_[47798]_  = \new_[47797]_  & \new_[47794]_ ;
  assign \new_[47799]_  = \new_[47798]_  & \new_[47791]_ ;
  assign \new_[47802]_  = ~A267 & ~A235;
  assign \new_[47805]_  = ~A269 & ~A268;
  assign \new_[47806]_  = \new_[47805]_  & \new_[47802]_ ;
  assign \new_[47809]_  = A299 & A298;
  assign \new_[47812]_  = ~A301 & ~A300;
  assign \new_[47813]_  = \new_[47812]_  & \new_[47809]_ ;
  assign \new_[47814]_  = \new_[47813]_  & \new_[47806]_ ;
  assign \new_[47817]_  = ~A167 & A170;
  assign \new_[47820]_  = ~A199 & A166;
  assign \new_[47821]_  = \new_[47820]_  & \new_[47817]_ ;
  assign \new_[47824]_  = ~A202 & ~A200;
  assign \new_[47827]_  = ~A233 & ~A232;
  assign \new_[47828]_  = \new_[47827]_  & \new_[47824]_ ;
  assign \new_[47829]_  = \new_[47828]_  & \new_[47821]_ ;
  assign \new_[47832]_  = A265 & ~A235;
  assign \new_[47835]_  = ~A267 & A266;
  assign \new_[47836]_  = \new_[47835]_  & \new_[47832]_ ;
  assign \new_[47839]_  = ~A300 & ~A268;
  assign \new_[47842]_  = ~A302 & ~A301;
  assign \new_[47843]_  = \new_[47842]_  & \new_[47839]_ ;
  assign \new_[47844]_  = \new_[47843]_  & \new_[47836]_ ;
  assign \new_[47847]_  = ~A167 & A170;
  assign \new_[47850]_  = ~A199 & A166;
  assign \new_[47851]_  = \new_[47850]_  & \new_[47847]_ ;
  assign \new_[47854]_  = ~A202 & ~A200;
  assign \new_[47857]_  = ~A233 & ~A232;
  assign \new_[47858]_  = \new_[47857]_  & \new_[47854]_ ;
  assign \new_[47859]_  = \new_[47858]_  & \new_[47851]_ ;
  assign \new_[47862]_  = A265 & ~A235;
  assign \new_[47865]_  = ~A267 & A266;
  assign \new_[47866]_  = \new_[47865]_  & \new_[47862]_ ;
  assign \new_[47869]_  = ~A298 & ~A268;
  assign \new_[47872]_  = ~A301 & ~A299;
  assign \new_[47873]_  = \new_[47872]_  & \new_[47869]_ ;
  assign \new_[47874]_  = \new_[47873]_  & \new_[47866]_ ;
  assign \new_[47877]_  = ~A167 & A170;
  assign \new_[47880]_  = ~A199 & A166;
  assign \new_[47881]_  = \new_[47880]_  & \new_[47877]_ ;
  assign \new_[47884]_  = ~A202 & ~A200;
  assign \new_[47887]_  = ~A233 & ~A232;
  assign \new_[47888]_  = \new_[47887]_  & \new_[47884]_ ;
  assign \new_[47889]_  = \new_[47888]_  & \new_[47881]_ ;
  assign \new_[47892]_  = ~A265 & ~A235;
  assign \new_[47895]_  = ~A268 & ~A266;
  assign \new_[47896]_  = \new_[47895]_  & \new_[47892]_ ;
  assign \new_[47899]_  = A299 & A298;
  assign \new_[47902]_  = ~A301 & ~A300;
  assign \new_[47903]_  = \new_[47902]_  & \new_[47899]_ ;
  assign \new_[47904]_  = \new_[47903]_  & \new_[47896]_ ;
  assign \new_[47907]_  = ~A201 & A169;
  assign \new_[47910]_  = ~A203 & ~A202;
  assign \new_[47911]_  = \new_[47910]_  & \new_[47907]_ ;
  assign \new_[47914]_  = A233 & A232;
  assign \new_[47917]_  = ~A235 & ~A234;
  assign \new_[47918]_  = \new_[47917]_  & \new_[47914]_ ;
  assign \new_[47919]_  = \new_[47918]_  & \new_[47911]_ ;
  assign \new_[47922]_  = A266 & A265;
  assign \new_[47925]_  = ~A268 & ~A267;
  assign \new_[47926]_  = \new_[47925]_  & \new_[47922]_ ;
  assign \new_[47929]_  = A299 & A298;
  assign \new_[47932]_  = ~A301 & ~A300;
  assign \new_[47933]_  = \new_[47932]_  & \new_[47929]_ ;
  assign \new_[47934]_  = \new_[47933]_  & \new_[47926]_ ;
  assign \new_[47937]_  = A199 & A169;
  assign \new_[47940]_  = ~A201 & A200;
  assign \new_[47941]_  = \new_[47940]_  & \new_[47937]_ ;
  assign \new_[47944]_  = ~A234 & ~A202;
  assign \new_[47947]_  = ~A236 & ~A235;
  assign \new_[47948]_  = \new_[47947]_  & \new_[47944]_ ;
  assign \new_[47949]_  = \new_[47948]_  & \new_[47941]_ ;
  assign \new_[47952]_  = A266 & A265;
  assign \new_[47955]_  = ~A268 & ~A267;
  assign \new_[47956]_  = \new_[47955]_  & \new_[47952]_ ;
  assign \new_[47959]_  = A299 & A298;
  assign \new_[47962]_  = ~A301 & ~A300;
  assign \new_[47963]_  = \new_[47962]_  & \new_[47959]_ ;
  assign \new_[47964]_  = \new_[47963]_  & \new_[47956]_ ;
  assign \new_[47967]_  = A199 & A169;
  assign \new_[47970]_  = ~A201 & A200;
  assign \new_[47971]_  = \new_[47970]_  & \new_[47967]_ ;
  assign \new_[47974]_  = A232 & ~A202;
  assign \new_[47977]_  = ~A234 & A233;
  assign \new_[47978]_  = \new_[47977]_  & \new_[47974]_ ;
  assign \new_[47979]_  = \new_[47978]_  & \new_[47971]_ ;
  assign \new_[47982]_  = ~A267 & ~A235;
  assign \new_[47985]_  = ~A269 & ~A268;
  assign \new_[47986]_  = \new_[47985]_  & \new_[47982]_ ;
  assign \new_[47989]_  = A299 & A298;
  assign \new_[47992]_  = ~A301 & ~A300;
  assign \new_[47993]_  = \new_[47992]_  & \new_[47989]_ ;
  assign \new_[47994]_  = \new_[47993]_  & \new_[47986]_ ;
  assign \new_[47997]_  = A199 & A169;
  assign \new_[48000]_  = ~A201 & A200;
  assign \new_[48001]_  = \new_[48000]_  & \new_[47997]_ ;
  assign \new_[48004]_  = A232 & ~A202;
  assign \new_[48007]_  = ~A234 & A233;
  assign \new_[48008]_  = \new_[48007]_  & \new_[48004]_ ;
  assign \new_[48009]_  = \new_[48008]_  & \new_[48001]_ ;
  assign \new_[48012]_  = A265 & ~A235;
  assign \new_[48015]_  = ~A267 & A266;
  assign \new_[48016]_  = \new_[48015]_  & \new_[48012]_ ;
  assign \new_[48019]_  = ~A300 & ~A268;
  assign \new_[48022]_  = ~A302 & ~A301;
  assign \new_[48023]_  = \new_[48022]_  & \new_[48019]_ ;
  assign \new_[48024]_  = \new_[48023]_  & \new_[48016]_ ;
  assign \new_[48027]_  = A199 & A169;
  assign \new_[48030]_  = ~A201 & A200;
  assign \new_[48031]_  = \new_[48030]_  & \new_[48027]_ ;
  assign \new_[48034]_  = A232 & ~A202;
  assign \new_[48037]_  = ~A234 & A233;
  assign \new_[48038]_  = \new_[48037]_  & \new_[48034]_ ;
  assign \new_[48039]_  = \new_[48038]_  & \new_[48031]_ ;
  assign \new_[48042]_  = A265 & ~A235;
  assign \new_[48045]_  = ~A267 & A266;
  assign \new_[48046]_  = \new_[48045]_  & \new_[48042]_ ;
  assign \new_[48049]_  = ~A298 & ~A268;
  assign \new_[48052]_  = ~A301 & ~A299;
  assign \new_[48053]_  = \new_[48052]_  & \new_[48049]_ ;
  assign \new_[48054]_  = \new_[48053]_  & \new_[48046]_ ;
  assign \new_[48057]_  = A199 & A169;
  assign \new_[48060]_  = ~A201 & A200;
  assign \new_[48061]_  = \new_[48060]_  & \new_[48057]_ ;
  assign \new_[48064]_  = A232 & ~A202;
  assign \new_[48067]_  = ~A234 & A233;
  assign \new_[48068]_  = \new_[48067]_  & \new_[48064]_ ;
  assign \new_[48069]_  = \new_[48068]_  & \new_[48061]_ ;
  assign \new_[48072]_  = ~A265 & ~A235;
  assign \new_[48075]_  = ~A268 & ~A266;
  assign \new_[48076]_  = \new_[48075]_  & \new_[48072]_ ;
  assign \new_[48079]_  = A299 & A298;
  assign \new_[48082]_  = ~A301 & ~A300;
  assign \new_[48083]_  = \new_[48082]_  & \new_[48079]_ ;
  assign \new_[48084]_  = \new_[48083]_  & \new_[48076]_ ;
  assign \new_[48087]_  = A199 & A169;
  assign \new_[48090]_  = ~A201 & A200;
  assign \new_[48091]_  = \new_[48090]_  & \new_[48087]_ ;
  assign \new_[48094]_  = ~A232 & ~A202;
  assign \new_[48097]_  = ~A235 & ~A233;
  assign \new_[48098]_  = \new_[48097]_  & \new_[48094]_ ;
  assign \new_[48099]_  = \new_[48098]_  & \new_[48091]_ ;
  assign \new_[48102]_  = A266 & A265;
  assign \new_[48105]_  = ~A268 & ~A267;
  assign \new_[48106]_  = \new_[48105]_  & \new_[48102]_ ;
  assign \new_[48109]_  = A299 & A298;
  assign \new_[48112]_  = ~A301 & ~A300;
  assign \new_[48113]_  = \new_[48112]_  & \new_[48109]_ ;
  assign \new_[48114]_  = \new_[48113]_  & \new_[48106]_ ;
  assign \new_[48117]_  = ~A199 & A169;
  assign \new_[48120]_  = ~A202 & ~A200;
  assign \new_[48121]_  = \new_[48120]_  & \new_[48117]_ ;
  assign \new_[48124]_  = A233 & A232;
  assign \new_[48127]_  = ~A235 & ~A234;
  assign \new_[48128]_  = \new_[48127]_  & \new_[48124]_ ;
  assign \new_[48129]_  = \new_[48128]_  & \new_[48121]_ ;
  assign \new_[48132]_  = A266 & A265;
  assign \new_[48135]_  = ~A268 & ~A267;
  assign \new_[48136]_  = \new_[48135]_  & \new_[48132]_ ;
  assign \new_[48139]_  = A299 & A298;
  assign \new_[48142]_  = ~A301 & ~A300;
  assign \new_[48143]_  = \new_[48142]_  & \new_[48139]_ ;
  assign \new_[48144]_  = \new_[48143]_  & \new_[48136]_ ;
  assign \new_[48147]_  = ~A167 & ~A169;
  assign \new_[48150]_  = A202 & ~A166;
  assign \new_[48151]_  = \new_[48150]_  & \new_[48147]_ ;
  assign \new_[48154]_  = A233 & A232;
  assign \new_[48157]_  = ~A235 & ~A234;
  assign \new_[48158]_  = \new_[48157]_  & \new_[48154]_ ;
  assign \new_[48159]_  = \new_[48158]_  & \new_[48151]_ ;
  assign \new_[48162]_  = A266 & A265;
  assign \new_[48165]_  = ~A268 & ~A267;
  assign \new_[48166]_  = \new_[48165]_  & \new_[48162]_ ;
  assign \new_[48169]_  = A299 & A298;
  assign \new_[48172]_  = ~A301 & ~A300;
  assign \new_[48173]_  = \new_[48172]_  & \new_[48169]_ ;
  assign \new_[48174]_  = \new_[48173]_  & \new_[48166]_ ;
  assign \new_[48177]_  = ~A167 & ~A169;
  assign \new_[48180]_  = A199 & ~A166;
  assign \new_[48181]_  = \new_[48180]_  & \new_[48177]_ ;
  assign \new_[48184]_  = ~A234 & A201;
  assign \new_[48187]_  = ~A236 & ~A235;
  assign \new_[48188]_  = \new_[48187]_  & \new_[48184]_ ;
  assign \new_[48189]_  = \new_[48188]_  & \new_[48181]_ ;
  assign \new_[48192]_  = A266 & A265;
  assign \new_[48195]_  = ~A268 & ~A267;
  assign \new_[48196]_  = \new_[48195]_  & \new_[48192]_ ;
  assign \new_[48199]_  = A299 & A298;
  assign \new_[48202]_  = ~A301 & ~A300;
  assign \new_[48203]_  = \new_[48202]_  & \new_[48199]_ ;
  assign \new_[48204]_  = \new_[48203]_  & \new_[48196]_ ;
  assign \new_[48207]_  = ~A167 & ~A169;
  assign \new_[48210]_  = A199 & ~A166;
  assign \new_[48211]_  = \new_[48210]_  & \new_[48207]_ ;
  assign \new_[48214]_  = A232 & A201;
  assign \new_[48217]_  = ~A234 & A233;
  assign \new_[48218]_  = \new_[48217]_  & \new_[48214]_ ;
  assign \new_[48219]_  = \new_[48218]_  & \new_[48211]_ ;
  assign \new_[48222]_  = ~A267 & ~A235;
  assign \new_[48225]_  = ~A269 & ~A268;
  assign \new_[48226]_  = \new_[48225]_  & \new_[48222]_ ;
  assign \new_[48229]_  = A299 & A298;
  assign \new_[48232]_  = ~A301 & ~A300;
  assign \new_[48233]_  = \new_[48232]_  & \new_[48229]_ ;
  assign \new_[48234]_  = \new_[48233]_  & \new_[48226]_ ;
  assign \new_[48237]_  = ~A167 & ~A169;
  assign \new_[48240]_  = A199 & ~A166;
  assign \new_[48241]_  = \new_[48240]_  & \new_[48237]_ ;
  assign \new_[48244]_  = A232 & A201;
  assign \new_[48247]_  = ~A234 & A233;
  assign \new_[48248]_  = \new_[48247]_  & \new_[48244]_ ;
  assign \new_[48249]_  = \new_[48248]_  & \new_[48241]_ ;
  assign \new_[48252]_  = A265 & ~A235;
  assign \new_[48255]_  = ~A267 & A266;
  assign \new_[48256]_  = \new_[48255]_  & \new_[48252]_ ;
  assign \new_[48259]_  = ~A300 & ~A268;
  assign \new_[48262]_  = ~A302 & ~A301;
  assign \new_[48263]_  = \new_[48262]_  & \new_[48259]_ ;
  assign \new_[48264]_  = \new_[48263]_  & \new_[48256]_ ;
  assign \new_[48267]_  = ~A167 & ~A169;
  assign \new_[48270]_  = A199 & ~A166;
  assign \new_[48271]_  = \new_[48270]_  & \new_[48267]_ ;
  assign \new_[48274]_  = A232 & A201;
  assign \new_[48277]_  = ~A234 & A233;
  assign \new_[48278]_  = \new_[48277]_  & \new_[48274]_ ;
  assign \new_[48279]_  = \new_[48278]_  & \new_[48271]_ ;
  assign \new_[48282]_  = A265 & ~A235;
  assign \new_[48285]_  = ~A267 & A266;
  assign \new_[48286]_  = \new_[48285]_  & \new_[48282]_ ;
  assign \new_[48289]_  = ~A298 & ~A268;
  assign \new_[48292]_  = ~A301 & ~A299;
  assign \new_[48293]_  = \new_[48292]_  & \new_[48289]_ ;
  assign \new_[48294]_  = \new_[48293]_  & \new_[48286]_ ;
  assign \new_[48297]_  = ~A167 & ~A169;
  assign \new_[48300]_  = A199 & ~A166;
  assign \new_[48301]_  = \new_[48300]_  & \new_[48297]_ ;
  assign \new_[48304]_  = A232 & A201;
  assign \new_[48307]_  = ~A234 & A233;
  assign \new_[48308]_  = \new_[48307]_  & \new_[48304]_ ;
  assign \new_[48309]_  = \new_[48308]_  & \new_[48301]_ ;
  assign \new_[48312]_  = ~A265 & ~A235;
  assign \new_[48315]_  = ~A268 & ~A266;
  assign \new_[48316]_  = \new_[48315]_  & \new_[48312]_ ;
  assign \new_[48319]_  = A299 & A298;
  assign \new_[48322]_  = ~A301 & ~A300;
  assign \new_[48323]_  = \new_[48322]_  & \new_[48319]_ ;
  assign \new_[48324]_  = \new_[48323]_  & \new_[48316]_ ;
  assign \new_[48327]_  = ~A167 & ~A169;
  assign \new_[48330]_  = A199 & ~A166;
  assign \new_[48331]_  = \new_[48330]_  & \new_[48327]_ ;
  assign \new_[48334]_  = ~A232 & A201;
  assign \new_[48337]_  = ~A235 & ~A233;
  assign \new_[48338]_  = \new_[48337]_  & \new_[48334]_ ;
  assign \new_[48339]_  = \new_[48338]_  & \new_[48331]_ ;
  assign \new_[48342]_  = A266 & A265;
  assign \new_[48345]_  = ~A268 & ~A267;
  assign \new_[48346]_  = \new_[48345]_  & \new_[48342]_ ;
  assign \new_[48349]_  = A299 & A298;
  assign \new_[48352]_  = ~A301 & ~A300;
  assign \new_[48353]_  = \new_[48352]_  & \new_[48349]_ ;
  assign \new_[48354]_  = \new_[48353]_  & \new_[48346]_ ;
  assign \new_[48357]_  = ~A167 & ~A169;
  assign \new_[48360]_  = A200 & ~A166;
  assign \new_[48361]_  = \new_[48360]_  & \new_[48357]_ ;
  assign \new_[48364]_  = ~A234 & A201;
  assign \new_[48367]_  = ~A236 & ~A235;
  assign \new_[48368]_  = \new_[48367]_  & \new_[48364]_ ;
  assign \new_[48369]_  = \new_[48368]_  & \new_[48361]_ ;
  assign \new_[48372]_  = A266 & A265;
  assign \new_[48375]_  = ~A268 & ~A267;
  assign \new_[48376]_  = \new_[48375]_  & \new_[48372]_ ;
  assign \new_[48379]_  = A299 & A298;
  assign \new_[48382]_  = ~A301 & ~A300;
  assign \new_[48383]_  = \new_[48382]_  & \new_[48379]_ ;
  assign \new_[48384]_  = \new_[48383]_  & \new_[48376]_ ;
  assign \new_[48387]_  = ~A167 & ~A169;
  assign \new_[48390]_  = A200 & ~A166;
  assign \new_[48391]_  = \new_[48390]_  & \new_[48387]_ ;
  assign \new_[48394]_  = A232 & A201;
  assign \new_[48397]_  = ~A234 & A233;
  assign \new_[48398]_  = \new_[48397]_  & \new_[48394]_ ;
  assign \new_[48399]_  = \new_[48398]_  & \new_[48391]_ ;
  assign \new_[48402]_  = ~A267 & ~A235;
  assign \new_[48405]_  = ~A269 & ~A268;
  assign \new_[48406]_  = \new_[48405]_  & \new_[48402]_ ;
  assign \new_[48409]_  = A299 & A298;
  assign \new_[48412]_  = ~A301 & ~A300;
  assign \new_[48413]_  = \new_[48412]_  & \new_[48409]_ ;
  assign \new_[48414]_  = \new_[48413]_  & \new_[48406]_ ;
  assign \new_[48417]_  = ~A167 & ~A169;
  assign \new_[48420]_  = A200 & ~A166;
  assign \new_[48421]_  = \new_[48420]_  & \new_[48417]_ ;
  assign \new_[48424]_  = A232 & A201;
  assign \new_[48427]_  = ~A234 & A233;
  assign \new_[48428]_  = \new_[48427]_  & \new_[48424]_ ;
  assign \new_[48429]_  = \new_[48428]_  & \new_[48421]_ ;
  assign \new_[48432]_  = A265 & ~A235;
  assign \new_[48435]_  = ~A267 & A266;
  assign \new_[48436]_  = \new_[48435]_  & \new_[48432]_ ;
  assign \new_[48439]_  = ~A300 & ~A268;
  assign \new_[48442]_  = ~A302 & ~A301;
  assign \new_[48443]_  = \new_[48442]_  & \new_[48439]_ ;
  assign \new_[48444]_  = \new_[48443]_  & \new_[48436]_ ;
  assign \new_[48447]_  = ~A167 & ~A169;
  assign \new_[48450]_  = A200 & ~A166;
  assign \new_[48451]_  = \new_[48450]_  & \new_[48447]_ ;
  assign \new_[48454]_  = A232 & A201;
  assign \new_[48457]_  = ~A234 & A233;
  assign \new_[48458]_  = \new_[48457]_  & \new_[48454]_ ;
  assign \new_[48459]_  = \new_[48458]_  & \new_[48451]_ ;
  assign \new_[48462]_  = A265 & ~A235;
  assign \new_[48465]_  = ~A267 & A266;
  assign \new_[48466]_  = \new_[48465]_  & \new_[48462]_ ;
  assign \new_[48469]_  = ~A298 & ~A268;
  assign \new_[48472]_  = ~A301 & ~A299;
  assign \new_[48473]_  = \new_[48472]_  & \new_[48469]_ ;
  assign \new_[48474]_  = \new_[48473]_  & \new_[48466]_ ;
  assign \new_[48477]_  = ~A167 & ~A169;
  assign \new_[48480]_  = A200 & ~A166;
  assign \new_[48481]_  = \new_[48480]_  & \new_[48477]_ ;
  assign \new_[48484]_  = A232 & A201;
  assign \new_[48487]_  = ~A234 & A233;
  assign \new_[48488]_  = \new_[48487]_  & \new_[48484]_ ;
  assign \new_[48489]_  = \new_[48488]_  & \new_[48481]_ ;
  assign \new_[48492]_  = ~A265 & ~A235;
  assign \new_[48495]_  = ~A268 & ~A266;
  assign \new_[48496]_  = \new_[48495]_  & \new_[48492]_ ;
  assign \new_[48499]_  = A299 & A298;
  assign \new_[48502]_  = ~A301 & ~A300;
  assign \new_[48503]_  = \new_[48502]_  & \new_[48499]_ ;
  assign \new_[48504]_  = \new_[48503]_  & \new_[48496]_ ;
  assign \new_[48507]_  = ~A167 & ~A169;
  assign \new_[48510]_  = A200 & ~A166;
  assign \new_[48511]_  = \new_[48510]_  & \new_[48507]_ ;
  assign \new_[48514]_  = ~A232 & A201;
  assign \new_[48517]_  = ~A235 & ~A233;
  assign \new_[48518]_  = \new_[48517]_  & \new_[48514]_ ;
  assign \new_[48519]_  = \new_[48518]_  & \new_[48511]_ ;
  assign \new_[48522]_  = A266 & A265;
  assign \new_[48525]_  = ~A268 & ~A267;
  assign \new_[48526]_  = \new_[48525]_  & \new_[48522]_ ;
  assign \new_[48529]_  = A299 & A298;
  assign \new_[48532]_  = ~A301 & ~A300;
  assign \new_[48533]_  = \new_[48532]_  & \new_[48529]_ ;
  assign \new_[48534]_  = \new_[48533]_  & \new_[48526]_ ;
  assign \new_[48537]_  = ~A167 & ~A169;
  assign \new_[48540]_  = ~A199 & ~A166;
  assign \new_[48541]_  = \new_[48540]_  & \new_[48537]_ ;
  assign \new_[48544]_  = A203 & A200;
  assign \new_[48547]_  = ~A235 & ~A234;
  assign \new_[48548]_  = \new_[48547]_  & \new_[48544]_ ;
  assign \new_[48549]_  = \new_[48548]_  & \new_[48541]_ ;
  assign \new_[48552]_  = ~A267 & ~A236;
  assign \new_[48555]_  = ~A269 & ~A268;
  assign \new_[48556]_  = \new_[48555]_  & \new_[48552]_ ;
  assign \new_[48559]_  = A299 & A298;
  assign \new_[48562]_  = ~A301 & ~A300;
  assign \new_[48563]_  = \new_[48562]_  & \new_[48559]_ ;
  assign \new_[48564]_  = \new_[48563]_  & \new_[48556]_ ;
  assign \new_[48567]_  = ~A167 & ~A169;
  assign \new_[48570]_  = ~A199 & ~A166;
  assign \new_[48571]_  = \new_[48570]_  & \new_[48567]_ ;
  assign \new_[48574]_  = A203 & A200;
  assign \new_[48577]_  = ~A235 & ~A234;
  assign \new_[48578]_  = \new_[48577]_  & \new_[48574]_ ;
  assign \new_[48579]_  = \new_[48578]_  & \new_[48571]_ ;
  assign \new_[48582]_  = A265 & ~A236;
  assign \new_[48585]_  = ~A267 & A266;
  assign \new_[48586]_  = \new_[48585]_  & \new_[48582]_ ;
  assign \new_[48589]_  = ~A300 & ~A268;
  assign \new_[48592]_  = ~A302 & ~A301;
  assign \new_[48593]_  = \new_[48592]_  & \new_[48589]_ ;
  assign \new_[48594]_  = \new_[48593]_  & \new_[48586]_ ;
  assign \new_[48597]_  = ~A167 & ~A169;
  assign \new_[48600]_  = ~A199 & ~A166;
  assign \new_[48601]_  = \new_[48600]_  & \new_[48597]_ ;
  assign \new_[48604]_  = A203 & A200;
  assign \new_[48607]_  = ~A235 & ~A234;
  assign \new_[48608]_  = \new_[48607]_  & \new_[48604]_ ;
  assign \new_[48609]_  = \new_[48608]_  & \new_[48601]_ ;
  assign \new_[48612]_  = A265 & ~A236;
  assign \new_[48615]_  = ~A267 & A266;
  assign \new_[48616]_  = \new_[48615]_  & \new_[48612]_ ;
  assign \new_[48619]_  = ~A298 & ~A268;
  assign \new_[48622]_  = ~A301 & ~A299;
  assign \new_[48623]_  = \new_[48622]_  & \new_[48619]_ ;
  assign \new_[48624]_  = \new_[48623]_  & \new_[48616]_ ;
  assign \new_[48627]_  = ~A167 & ~A169;
  assign \new_[48630]_  = ~A199 & ~A166;
  assign \new_[48631]_  = \new_[48630]_  & \new_[48627]_ ;
  assign \new_[48634]_  = A203 & A200;
  assign \new_[48637]_  = ~A235 & ~A234;
  assign \new_[48638]_  = \new_[48637]_  & \new_[48634]_ ;
  assign \new_[48639]_  = \new_[48638]_  & \new_[48631]_ ;
  assign \new_[48642]_  = ~A265 & ~A236;
  assign \new_[48645]_  = ~A268 & ~A266;
  assign \new_[48646]_  = \new_[48645]_  & \new_[48642]_ ;
  assign \new_[48649]_  = A299 & A298;
  assign \new_[48652]_  = ~A301 & ~A300;
  assign \new_[48653]_  = \new_[48652]_  & \new_[48649]_ ;
  assign \new_[48654]_  = \new_[48653]_  & \new_[48646]_ ;
  assign \new_[48657]_  = ~A167 & ~A169;
  assign \new_[48660]_  = ~A199 & ~A166;
  assign \new_[48661]_  = \new_[48660]_  & \new_[48657]_ ;
  assign \new_[48664]_  = A203 & A200;
  assign \new_[48667]_  = A233 & A232;
  assign \new_[48668]_  = \new_[48667]_  & \new_[48664]_ ;
  assign \new_[48669]_  = \new_[48668]_  & \new_[48661]_ ;
  assign \new_[48672]_  = ~A235 & ~A234;
  assign \new_[48675]_  = ~A268 & ~A267;
  assign \new_[48676]_  = \new_[48675]_  & \new_[48672]_ ;
  assign \new_[48679]_  = ~A300 & ~A269;
  assign \new_[48682]_  = ~A302 & ~A301;
  assign \new_[48683]_  = \new_[48682]_  & \new_[48679]_ ;
  assign \new_[48684]_  = \new_[48683]_  & \new_[48676]_ ;
  assign \new_[48687]_  = ~A167 & ~A169;
  assign \new_[48690]_  = ~A199 & ~A166;
  assign \new_[48691]_  = \new_[48690]_  & \new_[48687]_ ;
  assign \new_[48694]_  = A203 & A200;
  assign \new_[48697]_  = A233 & A232;
  assign \new_[48698]_  = \new_[48697]_  & \new_[48694]_ ;
  assign \new_[48699]_  = \new_[48698]_  & \new_[48691]_ ;
  assign \new_[48702]_  = ~A235 & ~A234;
  assign \new_[48705]_  = ~A268 & ~A267;
  assign \new_[48706]_  = \new_[48705]_  & \new_[48702]_ ;
  assign \new_[48709]_  = ~A298 & ~A269;
  assign \new_[48712]_  = ~A301 & ~A299;
  assign \new_[48713]_  = \new_[48712]_  & \new_[48709]_ ;
  assign \new_[48714]_  = \new_[48713]_  & \new_[48706]_ ;
  assign \new_[48717]_  = ~A167 & ~A169;
  assign \new_[48720]_  = ~A199 & ~A166;
  assign \new_[48721]_  = \new_[48720]_  & \new_[48717]_ ;
  assign \new_[48724]_  = A203 & A200;
  assign \new_[48727]_  = A233 & A232;
  assign \new_[48728]_  = \new_[48727]_  & \new_[48724]_ ;
  assign \new_[48729]_  = \new_[48728]_  & \new_[48721]_ ;
  assign \new_[48732]_  = ~A235 & ~A234;
  assign \new_[48735]_  = ~A266 & ~A265;
  assign \new_[48736]_  = \new_[48735]_  & \new_[48732]_ ;
  assign \new_[48739]_  = ~A300 & ~A268;
  assign \new_[48742]_  = ~A302 & ~A301;
  assign \new_[48743]_  = \new_[48742]_  & \new_[48739]_ ;
  assign \new_[48744]_  = \new_[48743]_  & \new_[48736]_ ;
  assign \new_[48747]_  = ~A167 & ~A169;
  assign \new_[48750]_  = ~A199 & ~A166;
  assign \new_[48751]_  = \new_[48750]_  & \new_[48747]_ ;
  assign \new_[48754]_  = A203 & A200;
  assign \new_[48757]_  = A233 & A232;
  assign \new_[48758]_  = \new_[48757]_  & \new_[48754]_ ;
  assign \new_[48759]_  = \new_[48758]_  & \new_[48751]_ ;
  assign \new_[48762]_  = ~A235 & ~A234;
  assign \new_[48765]_  = ~A266 & ~A265;
  assign \new_[48766]_  = \new_[48765]_  & \new_[48762]_ ;
  assign \new_[48769]_  = ~A298 & ~A268;
  assign \new_[48772]_  = ~A301 & ~A299;
  assign \new_[48773]_  = \new_[48772]_  & \new_[48769]_ ;
  assign \new_[48774]_  = \new_[48773]_  & \new_[48766]_ ;
  assign \new_[48777]_  = ~A167 & ~A169;
  assign \new_[48780]_  = ~A199 & ~A166;
  assign \new_[48781]_  = \new_[48780]_  & \new_[48777]_ ;
  assign \new_[48784]_  = A203 & A200;
  assign \new_[48787]_  = ~A233 & ~A232;
  assign \new_[48788]_  = \new_[48787]_  & \new_[48784]_ ;
  assign \new_[48789]_  = \new_[48788]_  & \new_[48781]_ ;
  assign \new_[48792]_  = ~A267 & ~A235;
  assign \new_[48795]_  = ~A269 & ~A268;
  assign \new_[48796]_  = \new_[48795]_  & \new_[48792]_ ;
  assign \new_[48799]_  = A299 & A298;
  assign \new_[48802]_  = ~A301 & ~A300;
  assign \new_[48803]_  = \new_[48802]_  & \new_[48799]_ ;
  assign \new_[48804]_  = \new_[48803]_  & \new_[48796]_ ;
  assign \new_[48807]_  = ~A167 & ~A169;
  assign \new_[48810]_  = ~A199 & ~A166;
  assign \new_[48811]_  = \new_[48810]_  & \new_[48807]_ ;
  assign \new_[48814]_  = A203 & A200;
  assign \new_[48817]_  = ~A233 & ~A232;
  assign \new_[48818]_  = \new_[48817]_  & \new_[48814]_ ;
  assign \new_[48819]_  = \new_[48818]_  & \new_[48811]_ ;
  assign \new_[48822]_  = A265 & ~A235;
  assign \new_[48825]_  = ~A267 & A266;
  assign \new_[48826]_  = \new_[48825]_  & \new_[48822]_ ;
  assign \new_[48829]_  = ~A300 & ~A268;
  assign \new_[48832]_  = ~A302 & ~A301;
  assign \new_[48833]_  = \new_[48832]_  & \new_[48829]_ ;
  assign \new_[48834]_  = \new_[48833]_  & \new_[48826]_ ;
  assign \new_[48837]_  = ~A167 & ~A169;
  assign \new_[48840]_  = ~A199 & ~A166;
  assign \new_[48841]_  = \new_[48840]_  & \new_[48837]_ ;
  assign \new_[48844]_  = A203 & A200;
  assign \new_[48847]_  = ~A233 & ~A232;
  assign \new_[48848]_  = \new_[48847]_  & \new_[48844]_ ;
  assign \new_[48849]_  = \new_[48848]_  & \new_[48841]_ ;
  assign \new_[48852]_  = A265 & ~A235;
  assign \new_[48855]_  = ~A267 & A266;
  assign \new_[48856]_  = \new_[48855]_  & \new_[48852]_ ;
  assign \new_[48859]_  = ~A298 & ~A268;
  assign \new_[48862]_  = ~A301 & ~A299;
  assign \new_[48863]_  = \new_[48862]_  & \new_[48859]_ ;
  assign \new_[48864]_  = \new_[48863]_  & \new_[48856]_ ;
  assign \new_[48867]_  = ~A167 & ~A169;
  assign \new_[48870]_  = ~A199 & ~A166;
  assign \new_[48871]_  = \new_[48870]_  & \new_[48867]_ ;
  assign \new_[48874]_  = A203 & A200;
  assign \new_[48877]_  = ~A233 & ~A232;
  assign \new_[48878]_  = \new_[48877]_  & \new_[48874]_ ;
  assign \new_[48879]_  = \new_[48878]_  & \new_[48871]_ ;
  assign \new_[48882]_  = ~A265 & ~A235;
  assign \new_[48885]_  = ~A268 & ~A266;
  assign \new_[48886]_  = \new_[48885]_  & \new_[48882]_ ;
  assign \new_[48889]_  = A299 & A298;
  assign \new_[48892]_  = ~A301 & ~A300;
  assign \new_[48893]_  = \new_[48892]_  & \new_[48889]_ ;
  assign \new_[48894]_  = \new_[48893]_  & \new_[48886]_ ;
  assign \new_[48897]_  = ~A167 & ~A169;
  assign \new_[48900]_  = A199 & ~A166;
  assign \new_[48901]_  = \new_[48900]_  & \new_[48897]_ ;
  assign \new_[48904]_  = A203 & ~A200;
  assign \new_[48907]_  = ~A235 & ~A234;
  assign \new_[48908]_  = \new_[48907]_  & \new_[48904]_ ;
  assign \new_[48909]_  = \new_[48908]_  & \new_[48901]_ ;
  assign \new_[48912]_  = ~A267 & ~A236;
  assign \new_[48915]_  = ~A269 & ~A268;
  assign \new_[48916]_  = \new_[48915]_  & \new_[48912]_ ;
  assign \new_[48919]_  = A299 & A298;
  assign \new_[48922]_  = ~A301 & ~A300;
  assign \new_[48923]_  = \new_[48922]_  & \new_[48919]_ ;
  assign \new_[48924]_  = \new_[48923]_  & \new_[48916]_ ;
  assign \new_[48927]_  = ~A167 & ~A169;
  assign \new_[48930]_  = A199 & ~A166;
  assign \new_[48931]_  = \new_[48930]_  & \new_[48927]_ ;
  assign \new_[48934]_  = A203 & ~A200;
  assign \new_[48937]_  = ~A235 & ~A234;
  assign \new_[48938]_  = \new_[48937]_  & \new_[48934]_ ;
  assign \new_[48939]_  = \new_[48938]_  & \new_[48931]_ ;
  assign \new_[48942]_  = A265 & ~A236;
  assign \new_[48945]_  = ~A267 & A266;
  assign \new_[48946]_  = \new_[48945]_  & \new_[48942]_ ;
  assign \new_[48949]_  = ~A300 & ~A268;
  assign \new_[48952]_  = ~A302 & ~A301;
  assign \new_[48953]_  = \new_[48952]_  & \new_[48949]_ ;
  assign \new_[48954]_  = \new_[48953]_  & \new_[48946]_ ;
  assign \new_[48957]_  = ~A167 & ~A169;
  assign \new_[48960]_  = A199 & ~A166;
  assign \new_[48961]_  = \new_[48960]_  & \new_[48957]_ ;
  assign \new_[48964]_  = A203 & ~A200;
  assign \new_[48967]_  = ~A235 & ~A234;
  assign \new_[48968]_  = \new_[48967]_  & \new_[48964]_ ;
  assign \new_[48969]_  = \new_[48968]_  & \new_[48961]_ ;
  assign \new_[48972]_  = A265 & ~A236;
  assign \new_[48975]_  = ~A267 & A266;
  assign \new_[48976]_  = \new_[48975]_  & \new_[48972]_ ;
  assign \new_[48979]_  = ~A298 & ~A268;
  assign \new_[48982]_  = ~A301 & ~A299;
  assign \new_[48983]_  = \new_[48982]_  & \new_[48979]_ ;
  assign \new_[48984]_  = \new_[48983]_  & \new_[48976]_ ;
  assign \new_[48987]_  = ~A167 & ~A169;
  assign \new_[48990]_  = A199 & ~A166;
  assign \new_[48991]_  = \new_[48990]_  & \new_[48987]_ ;
  assign \new_[48994]_  = A203 & ~A200;
  assign \new_[48997]_  = ~A235 & ~A234;
  assign \new_[48998]_  = \new_[48997]_  & \new_[48994]_ ;
  assign \new_[48999]_  = \new_[48998]_  & \new_[48991]_ ;
  assign \new_[49002]_  = ~A265 & ~A236;
  assign \new_[49005]_  = ~A268 & ~A266;
  assign \new_[49006]_  = \new_[49005]_  & \new_[49002]_ ;
  assign \new_[49009]_  = A299 & A298;
  assign \new_[49012]_  = ~A301 & ~A300;
  assign \new_[49013]_  = \new_[49012]_  & \new_[49009]_ ;
  assign \new_[49014]_  = \new_[49013]_  & \new_[49006]_ ;
  assign \new_[49017]_  = ~A167 & ~A169;
  assign \new_[49020]_  = A199 & ~A166;
  assign \new_[49021]_  = \new_[49020]_  & \new_[49017]_ ;
  assign \new_[49024]_  = A203 & ~A200;
  assign \new_[49027]_  = A233 & A232;
  assign \new_[49028]_  = \new_[49027]_  & \new_[49024]_ ;
  assign \new_[49029]_  = \new_[49028]_  & \new_[49021]_ ;
  assign \new_[49032]_  = ~A235 & ~A234;
  assign \new_[49035]_  = ~A268 & ~A267;
  assign \new_[49036]_  = \new_[49035]_  & \new_[49032]_ ;
  assign \new_[49039]_  = ~A300 & ~A269;
  assign \new_[49042]_  = ~A302 & ~A301;
  assign \new_[49043]_  = \new_[49042]_  & \new_[49039]_ ;
  assign \new_[49044]_  = \new_[49043]_  & \new_[49036]_ ;
  assign \new_[49047]_  = ~A167 & ~A169;
  assign \new_[49050]_  = A199 & ~A166;
  assign \new_[49051]_  = \new_[49050]_  & \new_[49047]_ ;
  assign \new_[49054]_  = A203 & ~A200;
  assign \new_[49057]_  = A233 & A232;
  assign \new_[49058]_  = \new_[49057]_  & \new_[49054]_ ;
  assign \new_[49059]_  = \new_[49058]_  & \new_[49051]_ ;
  assign \new_[49062]_  = ~A235 & ~A234;
  assign \new_[49065]_  = ~A268 & ~A267;
  assign \new_[49066]_  = \new_[49065]_  & \new_[49062]_ ;
  assign \new_[49069]_  = ~A298 & ~A269;
  assign \new_[49072]_  = ~A301 & ~A299;
  assign \new_[49073]_  = \new_[49072]_  & \new_[49069]_ ;
  assign \new_[49074]_  = \new_[49073]_  & \new_[49066]_ ;
  assign \new_[49077]_  = ~A167 & ~A169;
  assign \new_[49080]_  = A199 & ~A166;
  assign \new_[49081]_  = \new_[49080]_  & \new_[49077]_ ;
  assign \new_[49084]_  = A203 & ~A200;
  assign \new_[49087]_  = A233 & A232;
  assign \new_[49088]_  = \new_[49087]_  & \new_[49084]_ ;
  assign \new_[49089]_  = \new_[49088]_  & \new_[49081]_ ;
  assign \new_[49092]_  = ~A235 & ~A234;
  assign \new_[49095]_  = ~A266 & ~A265;
  assign \new_[49096]_  = \new_[49095]_  & \new_[49092]_ ;
  assign \new_[49099]_  = ~A300 & ~A268;
  assign \new_[49102]_  = ~A302 & ~A301;
  assign \new_[49103]_  = \new_[49102]_  & \new_[49099]_ ;
  assign \new_[49104]_  = \new_[49103]_  & \new_[49096]_ ;
  assign \new_[49107]_  = ~A167 & ~A169;
  assign \new_[49110]_  = A199 & ~A166;
  assign \new_[49111]_  = \new_[49110]_  & \new_[49107]_ ;
  assign \new_[49114]_  = A203 & ~A200;
  assign \new_[49117]_  = A233 & A232;
  assign \new_[49118]_  = \new_[49117]_  & \new_[49114]_ ;
  assign \new_[49119]_  = \new_[49118]_  & \new_[49111]_ ;
  assign \new_[49122]_  = ~A235 & ~A234;
  assign \new_[49125]_  = ~A266 & ~A265;
  assign \new_[49126]_  = \new_[49125]_  & \new_[49122]_ ;
  assign \new_[49129]_  = ~A298 & ~A268;
  assign \new_[49132]_  = ~A301 & ~A299;
  assign \new_[49133]_  = \new_[49132]_  & \new_[49129]_ ;
  assign \new_[49134]_  = \new_[49133]_  & \new_[49126]_ ;
  assign \new_[49137]_  = ~A167 & ~A169;
  assign \new_[49140]_  = A199 & ~A166;
  assign \new_[49141]_  = \new_[49140]_  & \new_[49137]_ ;
  assign \new_[49144]_  = A203 & ~A200;
  assign \new_[49147]_  = ~A233 & ~A232;
  assign \new_[49148]_  = \new_[49147]_  & \new_[49144]_ ;
  assign \new_[49149]_  = \new_[49148]_  & \new_[49141]_ ;
  assign \new_[49152]_  = ~A267 & ~A235;
  assign \new_[49155]_  = ~A269 & ~A268;
  assign \new_[49156]_  = \new_[49155]_  & \new_[49152]_ ;
  assign \new_[49159]_  = A299 & A298;
  assign \new_[49162]_  = ~A301 & ~A300;
  assign \new_[49163]_  = \new_[49162]_  & \new_[49159]_ ;
  assign \new_[49164]_  = \new_[49163]_  & \new_[49156]_ ;
  assign \new_[49167]_  = ~A167 & ~A169;
  assign \new_[49170]_  = A199 & ~A166;
  assign \new_[49171]_  = \new_[49170]_  & \new_[49167]_ ;
  assign \new_[49174]_  = A203 & ~A200;
  assign \new_[49177]_  = ~A233 & ~A232;
  assign \new_[49178]_  = \new_[49177]_  & \new_[49174]_ ;
  assign \new_[49179]_  = \new_[49178]_  & \new_[49171]_ ;
  assign \new_[49182]_  = A265 & ~A235;
  assign \new_[49185]_  = ~A267 & A266;
  assign \new_[49186]_  = \new_[49185]_  & \new_[49182]_ ;
  assign \new_[49189]_  = ~A300 & ~A268;
  assign \new_[49192]_  = ~A302 & ~A301;
  assign \new_[49193]_  = \new_[49192]_  & \new_[49189]_ ;
  assign \new_[49194]_  = \new_[49193]_  & \new_[49186]_ ;
  assign \new_[49197]_  = ~A167 & ~A169;
  assign \new_[49200]_  = A199 & ~A166;
  assign \new_[49201]_  = \new_[49200]_  & \new_[49197]_ ;
  assign \new_[49204]_  = A203 & ~A200;
  assign \new_[49207]_  = ~A233 & ~A232;
  assign \new_[49208]_  = \new_[49207]_  & \new_[49204]_ ;
  assign \new_[49209]_  = \new_[49208]_  & \new_[49201]_ ;
  assign \new_[49212]_  = A265 & ~A235;
  assign \new_[49215]_  = ~A267 & A266;
  assign \new_[49216]_  = \new_[49215]_  & \new_[49212]_ ;
  assign \new_[49219]_  = ~A298 & ~A268;
  assign \new_[49222]_  = ~A301 & ~A299;
  assign \new_[49223]_  = \new_[49222]_  & \new_[49219]_ ;
  assign \new_[49224]_  = \new_[49223]_  & \new_[49216]_ ;
  assign \new_[49227]_  = ~A167 & ~A169;
  assign \new_[49230]_  = A199 & ~A166;
  assign \new_[49231]_  = \new_[49230]_  & \new_[49227]_ ;
  assign \new_[49234]_  = A203 & ~A200;
  assign \new_[49237]_  = ~A233 & ~A232;
  assign \new_[49238]_  = \new_[49237]_  & \new_[49234]_ ;
  assign \new_[49239]_  = \new_[49238]_  & \new_[49231]_ ;
  assign \new_[49242]_  = ~A265 & ~A235;
  assign \new_[49245]_  = ~A268 & ~A266;
  assign \new_[49246]_  = \new_[49245]_  & \new_[49242]_ ;
  assign \new_[49249]_  = A299 & A298;
  assign \new_[49252]_  = ~A301 & ~A300;
  assign \new_[49253]_  = \new_[49252]_  & \new_[49249]_ ;
  assign \new_[49254]_  = \new_[49253]_  & \new_[49246]_ ;
  assign \new_[49257]_  = ~A168 & ~A169;
  assign \new_[49260]_  = A166 & A167;
  assign \new_[49261]_  = \new_[49260]_  & \new_[49257]_ ;
  assign \new_[49264]_  = ~A234 & A202;
  assign \new_[49267]_  = ~A236 & ~A235;
  assign \new_[49268]_  = \new_[49267]_  & \new_[49264]_ ;
  assign \new_[49269]_  = \new_[49268]_  & \new_[49261]_ ;
  assign \new_[49272]_  = A266 & A265;
  assign \new_[49275]_  = ~A268 & ~A267;
  assign \new_[49276]_  = \new_[49275]_  & \new_[49272]_ ;
  assign \new_[49279]_  = A299 & A298;
  assign \new_[49282]_  = ~A301 & ~A300;
  assign \new_[49283]_  = \new_[49282]_  & \new_[49279]_ ;
  assign \new_[49284]_  = \new_[49283]_  & \new_[49276]_ ;
  assign \new_[49287]_  = ~A168 & ~A169;
  assign \new_[49290]_  = A166 & A167;
  assign \new_[49291]_  = \new_[49290]_  & \new_[49287]_ ;
  assign \new_[49294]_  = A232 & A202;
  assign \new_[49297]_  = ~A234 & A233;
  assign \new_[49298]_  = \new_[49297]_  & \new_[49294]_ ;
  assign \new_[49299]_  = \new_[49298]_  & \new_[49291]_ ;
  assign \new_[49302]_  = ~A267 & ~A235;
  assign \new_[49305]_  = ~A269 & ~A268;
  assign \new_[49306]_  = \new_[49305]_  & \new_[49302]_ ;
  assign \new_[49309]_  = A299 & A298;
  assign \new_[49312]_  = ~A301 & ~A300;
  assign \new_[49313]_  = \new_[49312]_  & \new_[49309]_ ;
  assign \new_[49314]_  = \new_[49313]_  & \new_[49306]_ ;
  assign \new_[49317]_  = ~A168 & ~A169;
  assign \new_[49320]_  = A166 & A167;
  assign \new_[49321]_  = \new_[49320]_  & \new_[49317]_ ;
  assign \new_[49324]_  = A232 & A202;
  assign \new_[49327]_  = ~A234 & A233;
  assign \new_[49328]_  = \new_[49327]_  & \new_[49324]_ ;
  assign \new_[49329]_  = \new_[49328]_  & \new_[49321]_ ;
  assign \new_[49332]_  = A265 & ~A235;
  assign \new_[49335]_  = ~A267 & A266;
  assign \new_[49336]_  = \new_[49335]_  & \new_[49332]_ ;
  assign \new_[49339]_  = ~A300 & ~A268;
  assign \new_[49342]_  = ~A302 & ~A301;
  assign \new_[49343]_  = \new_[49342]_  & \new_[49339]_ ;
  assign \new_[49344]_  = \new_[49343]_  & \new_[49336]_ ;
  assign \new_[49347]_  = ~A168 & ~A169;
  assign \new_[49350]_  = A166 & A167;
  assign \new_[49351]_  = \new_[49350]_  & \new_[49347]_ ;
  assign \new_[49354]_  = A232 & A202;
  assign \new_[49357]_  = ~A234 & A233;
  assign \new_[49358]_  = \new_[49357]_  & \new_[49354]_ ;
  assign \new_[49359]_  = \new_[49358]_  & \new_[49351]_ ;
  assign \new_[49362]_  = A265 & ~A235;
  assign \new_[49365]_  = ~A267 & A266;
  assign \new_[49366]_  = \new_[49365]_  & \new_[49362]_ ;
  assign \new_[49369]_  = ~A298 & ~A268;
  assign \new_[49372]_  = ~A301 & ~A299;
  assign \new_[49373]_  = \new_[49372]_  & \new_[49369]_ ;
  assign \new_[49374]_  = \new_[49373]_  & \new_[49366]_ ;
  assign \new_[49377]_  = ~A168 & ~A169;
  assign \new_[49380]_  = A166 & A167;
  assign \new_[49381]_  = \new_[49380]_  & \new_[49377]_ ;
  assign \new_[49384]_  = A232 & A202;
  assign \new_[49387]_  = ~A234 & A233;
  assign \new_[49388]_  = \new_[49387]_  & \new_[49384]_ ;
  assign \new_[49389]_  = \new_[49388]_  & \new_[49381]_ ;
  assign \new_[49392]_  = ~A265 & ~A235;
  assign \new_[49395]_  = ~A268 & ~A266;
  assign \new_[49396]_  = \new_[49395]_  & \new_[49392]_ ;
  assign \new_[49399]_  = A299 & A298;
  assign \new_[49402]_  = ~A301 & ~A300;
  assign \new_[49403]_  = \new_[49402]_  & \new_[49399]_ ;
  assign \new_[49404]_  = \new_[49403]_  & \new_[49396]_ ;
  assign \new_[49407]_  = ~A168 & ~A169;
  assign \new_[49410]_  = A166 & A167;
  assign \new_[49411]_  = \new_[49410]_  & \new_[49407]_ ;
  assign \new_[49414]_  = ~A232 & A202;
  assign \new_[49417]_  = ~A235 & ~A233;
  assign \new_[49418]_  = \new_[49417]_  & \new_[49414]_ ;
  assign \new_[49419]_  = \new_[49418]_  & \new_[49411]_ ;
  assign \new_[49422]_  = A266 & A265;
  assign \new_[49425]_  = ~A268 & ~A267;
  assign \new_[49426]_  = \new_[49425]_  & \new_[49422]_ ;
  assign \new_[49429]_  = A299 & A298;
  assign \new_[49432]_  = ~A301 & ~A300;
  assign \new_[49433]_  = \new_[49432]_  & \new_[49429]_ ;
  assign \new_[49434]_  = \new_[49433]_  & \new_[49426]_ ;
  assign \new_[49437]_  = ~A168 & ~A169;
  assign \new_[49440]_  = A166 & A167;
  assign \new_[49441]_  = \new_[49440]_  & \new_[49437]_ ;
  assign \new_[49444]_  = A201 & A199;
  assign \new_[49447]_  = ~A235 & ~A234;
  assign \new_[49448]_  = \new_[49447]_  & \new_[49444]_ ;
  assign \new_[49449]_  = \new_[49448]_  & \new_[49441]_ ;
  assign \new_[49452]_  = ~A267 & ~A236;
  assign \new_[49455]_  = ~A269 & ~A268;
  assign \new_[49456]_  = \new_[49455]_  & \new_[49452]_ ;
  assign \new_[49459]_  = A299 & A298;
  assign \new_[49462]_  = ~A301 & ~A300;
  assign \new_[49463]_  = \new_[49462]_  & \new_[49459]_ ;
  assign \new_[49464]_  = \new_[49463]_  & \new_[49456]_ ;
  assign \new_[49467]_  = ~A168 & ~A169;
  assign \new_[49470]_  = A166 & A167;
  assign \new_[49471]_  = \new_[49470]_  & \new_[49467]_ ;
  assign \new_[49474]_  = A201 & A199;
  assign \new_[49477]_  = ~A235 & ~A234;
  assign \new_[49478]_  = \new_[49477]_  & \new_[49474]_ ;
  assign \new_[49479]_  = \new_[49478]_  & \new_[49471]_ ;
  assign \new_[49482]_  = A265 & ~A236;
  assign \new_[49485]_  = ~A267 & A266;
  assign \new_[49486]_  = \new_[49485]_  & \new_[49482]_ ;
  assign \new_[49489]_  = ~A300 & ~A268;
  assign \new_[49492]_  = ~A302 & ~A301;
  assign \new_[49493]_  = \new_[49492]_  & \new_[49489]_ ;
  assign \new_[49494]_  = \new_[49493]_  & \new_[49486]_ ;
  assign \new_[49497]_  = ~A168 & ~A169;
  assign \new_[49500]_  = A166 & A167;
  assign \new_[49501]_  = \new_[49500]_  & \new_[49497]_ ;
  assign \new_[49504]_  = A201 & A199;
  assign \new_[49507]_  = ~A235 & ~A234;
  assign \new_[49508]_  = \new_[49507]_  & \new_[49504]_ ;
  assign \new_[49509]_  = \new_[49508]_  & \new_[49501]_ ;
  assign \new_[49512]_  = A265 & ~A236;
  assign \new_[49515]_  = ~A267 & A266;
  assign \new_[49516]_  = \new_[49515]_  & \new_[49512]_ ;
  assign \new_[49519]_  = ~A298 & ~A268;
  assign \new_[49522]_  = ~A301 & ~A299;
  assign \new_[49523]_  = \new_[49522]_  & \new_[49519]_ ;
  assign \new_[49524]_  = \new_[49523]_  & \new_[49516]_ ;
  assign \new_[49527]_  = ~A168 & ~A169;
  assign \new_[49530]_  = A166 & A167;
  assign \new_[49531]_  = \new_[49530]_  & \new_[49527]_ ;
  assign \new_[49534]_  = A201 & A199;
  assign \new_[49537]_  = ~A235 & ~A234;
  assign \new_[49538]_  = \new_[49537]_  & \new_[49534]_ ;
  assign \new_[49539]_  = \new_[49538]_  & \new_[49531]_ ;
  assign \new_[49542]_  = ~A265 & ~A236;
  assign \new_[49545]_  = ~A268 & ~A266;
  assign \new_[49546]_  = \new_[49545]_  & \new_[49542]_ ;
  assign \new_[49549]_  = A299 & A298;
  assign \new_[49552]_  = ~A301 & ~A300;
  assign \new_[49553]_  = \new_[49552]_  & \new_[49549]_ ;
  assign \new_[49554]_  = \new_[49553]_  & \new_[49546]_ ;
  assign \new_[49557]_  = ~A168 & ~A169;
  assign \new_[49560]_  = A166 & A167;
  assign \new_[49561]_  = \new_[49560]_  & \new_[49557]_ ;
  assign \new_[49564]_  = A201 & A199;
  assign \new_[49567]_  = A233 & A232;
  assign \new_[49568]_  = \new_[49567]_  & \new_[49564]_ ;
  assign \new_[49569]_  = \new_[49568]_  & \new_[49561]_ ;
  assign \new_[49572]_  = ~A235 & ~A234;
  assign \new_[49575]_  = ~A268 & ~A267;
  assign \new_[49576]_  = \new_[49575]_  & \new_[49572]_ ;
  assign \new_[49579]_  = ~A300 & ~A269;
  assign \new_[49582]_  = ~A302 & ~A301;
  assign \new_[49583]_  = \new_[49582]_  & \new_[49579]_ ;
  assign \new_[49584]_  = \new_[49583]_  & \new_[49576]_ ;
  assign \new_[49587]_  = ~A168 & ~A169;
  assign \new_[49590]_  = A166 & A167;
  assign \new_[49591]_  = \new_[49590]_  & \new_[49587]_ ;
  assign \new_[49594]_  = A201 & A199;
  assign \new_[49597]_  = A233 & A232;
  assign \new_[49598]_  = \new_[49597]_  & \new_[49594]_ ;
  assign \new_[49599]_  = \new_[49598]_  & \new_[49591]_ ;
  assign \new_[49602]_  = ~A235 & ~A234;
  assign \new_[49605]_  = ~A268 & ~A267;
  assign \new_[49606]_  = \new_[49605]_  & \new_[49602]_ ;
  assign \new_[49609]_  = ~A298 & ~A269;
  assign \new_[49612]_  = ~A301 & ~A299;
  assign \new_[49613]_  = \new_[49612]_  & \new_[49609]_ ;
  assign \new_[49614]_  = \new_[49613]_  & \new_[49606]_ ;
  assign \new_[49617]_  = ~A168 & ~A169;
  assign \new_[49620]_  = A166 & A167;
  assign \new_[49621]_  = \new_[49620]_  & \new_[49617]_ ;
  assign \new_[49624]_  = A201 & A199;
  assign \new_[49627]_  = A233 & A232;
  assign \new_[49628]_  = \new_[49627]_  & \new_[49624]_ ;
  assign \new_[49629]_  = \new_[49628]_  & \new_[49621]_ ;
  assign \new_[49632]_  = ~A235 & ~A234;
  assign \new_[49635]_  = ~A266 & ~A265;
  assign \new_[49636]_  = \new_[49635]_  & \new_[49632]_ ;
  assign \new_[49639]_  = ~A300 & ~A268;
  assign \new_[49642]_  = ~A302 & ~A301;
  assign \new_[49643]_  = \new_[49642]_  & \new_[49639]_ ;
  assign \new_[49644]_  = \new_[49643]_  & \new_[49636]_ ;
  assign \new_[49647]_  = ~A168 & ~A169;
  assign \new_[49650]_  = A166 & A167;
  assign \new_[49651]_  = \new_[49650]_  & \new_[49647]_ ;
  assign \new_[49654]_  = A201 & A199;
  assign \new_[49657]_  = A233 & A232;
  assign \new_[49658]_  = \new_[49657]_  & \new_[49654]_ ;
  assign \new_[49659]_  = \new_[49658]_  & \new_[49651]_ ;
  assign \new_[49662]_  = ~A235 & ~A234;
  assign \new_[49665]_  = ~A266 & ~A265;
  assign \new_[49666]_  = \new_[49665]_  & \new_[49662]_ ;
  assign \new_[49669]_  = ~A298 & ~A268;
  assign \new_[49672]_  = ~A301 & ~A299;
  assign \new_[49673]_  = \new_[49672]_  & \new_[49669]_ ;
  assign \new_[49674]_  = \new_[49673]_  & \new_[49666]_ ;
  assign \new_[49677]_  = ~A168 & ~A169;
  assign \new_[49680]_  = A166 & A167;
  assign \new_[49681]_  = \new_[49680]_  & \new_[49677]_ ;
  assign \new_[49684]_  = A201 & A199;
  assign \new_[49687]_  = ~A233 & ~A232;
  assign \new_[49688]_  = \new_[49687]_  & \new_[49684]_ ;
  assign \new_[49689]_  = \new_[49688]_  & \new_[49681]_ ;
  assign \new_[49692]_  = ~A267 & ~A235;
  assign \new_[49695]_  = ~A269 & ~A268;
  assign \new_[49696]_  = \new_[49695]_  & \new_[49692]_ ;
  assign \new_[49699]_  = A299 & A298;
  assign \new_[49702]_  = ~A301 & ~A300;
  assign \new_[49703]_  = \new_[49702]_  & \new_[49699]_ ;
  assign \new_[49704]_  = \new_[49703]_  & \new_[49696]_ ;
  assign \new_[49707]_  = ~A168 & ~A169;
  assign \new_[49710]_  = A166 & A167;
  assign \new_[49711]_  = \new_[49710]_  & \new_[49707]_ ;
  assign \new_[49714]_  = A201 & A199;
  assign \new_[49717]_  = ~A233 & ~A232;
  assign \new_[49718]_  = \new_[49717]_  & \new_[49714]_ ;
  assign \new_[49719]_  = \new_[49718]_  & \new_[49711]_ ;
  assign \new_[49722]_  = A265 & ~A235;
  assign \new_[49725]_  = ~A267 & A266;
  assign \new_[49726]_  = \new_[49725]_  & \new_[49722]_ ;
  assign \new_[49729]_  = ~A300 & ~A268;
  assign \new_[49732]_  = ~A302 & ~A301;
  assign \new_[49733]_  = \new_[49732]_  & \new_[49729]_ ;
  assign \new_[49734]_  = \new_[49733]_  & \new_[49726]_ ;
  assign \new_[49737]_  = ~A168 & ~A169;
  assign \new_[49740]_  = A166 & A167;
  assign \new_[49741]_  = \new_[49740]_  & \new_[49737]_ ;
  assign \new_[49744]_  = A201 & A199;
  assign \new_[49747]_  = ~A233 & ~A232;
  assign \new_[49748]_  = \new_[49747]_  & \new_[49744]_ ;
  assign \new_[49749]_  = \new_[49748]_  & \new_[49741]_ ;
  assign \new_[49752]_  = A265 & ~A235;
  assign \new_[49755]_  = ~A267 & A266;
  assign \new_[49756]_  = \new_[49755]_  & \new_[49752]_ ;
  assign \new_[49759]_  = ~A298 & ~A268;
  assign \new_[49762]_  = ~A301 & ~A299;
  assign \new_[49763]_  = \new_[49762]_  & \new_[49759]_ ;
  assign \new_[49764]_  = \new_[49763]_  & \new_[49756]_ ;
  assign \new_[49767]_  = ~A168 & ~A169;
  assign \new_[49770]_  = A166 & A167;
  assign \new_[49771]_  = \new_[49770]_  & \new_[49767]_ ;
  assign \new_[49774]_  = A201 & A199;
  assign \new_[49777]_  = ~A233 & ~A232;
  assign \new_[49778]_  = \new_[49777]_  & \new_[49774]_ ;
  assign \new_[49779]_  = \new_[49778]_  & \new_[49771]_ ;
  assign \new_[49782]_  = ~A265 & ~A235;
  assign \new_[49785]_  = ~A268 & ~A266;
  assign \new_[49786]_  = \new_[49785]_  & \new_[49782]_ ;
  assign \new_[49789]_  = A299 & A298;
  assign \new_[49792]_  = ~A301 & ~A300;
  assign \new_[49793]_  = \new_[49792]_  & \new_[49789]_ ;
  assign \new_[49794]_  = \new_[49793]_  & \new_[49786]_ ;
  assign \new_[49797]_  = ~A168 & ~A169;
  assign \new_[49800]_  = A166 & A167;
  assign \new_[49801]_  = \new_[49800]_  & \new_[49797]_ ;
  assign \new_[49804]_  = A201 & A200;
  assign \new_[49807]_  = ~A235 & ~A234;
  assign \new_[49808]_  = \new_[49807]_  & \new_[49804]_ ;
  assign \new_[49809]_  = \new_[49808]_  & \new_[49801]_ ;
  assign \new_[49812]_  = ~A267 & ~A236;
  assign \new_[49815]_  = ~A269 & ~A268;
  assign \new_[49816]_  = \new_[49815]_  & \new_[49812]_ ;
  assign \new_[49819]_  = A299 & A298;
  assign \new_[49822]_  = ~A301 & ~A300;
  assign \new_[49823]_  = \new_[49822]_  & \new_[49819]_ ;
  assign \new_[49824]_  = \new_[49823]_  & \new_[49816]_ ;
  assign \new_[49827]_  = ~A168 & ~A169;
  assign \new_[49830]_  = A166 & A167;
  assign \new_[49831]_  = \new_[49830]_  & \new_[49827]_ ;
  assign \new_[49834]_  = A201 & A200;
  assign \new_[49837]_  = ~A235 & ~A234;
  assign \new_[49838]_  = \new_[49837]_  & \new_[49834]_ ;
  assign \new_[49839]_  = \new_[49838]_  & \new_[49831]_ ;
  assign \new_[49842]_  = A265 & ~A236;
  assign \new_[49845]_  = ~A267 & A266;
  assign \new_[49846]_  = \new_[49845]_  & \new_[49842]_ ;
  assign \new_[49849]_  = ~A300 & ~A268;
  assign \new_[49852]_  = ~A302 & ~A301;
  assign \new_[49853]_  = \new_[49852]_  & \new_[49849]_ ;
  assign \new_[49854]_  = \new_[49853]_  & \new_[49846]_ ;
  assign \new_[49857]_  = ~A168 & ~A169;
  assign \new_[49860]_  = A166 & A167;
  assign \new_[49861]_  = \new_[49860]_  & \new_[49857]_ ;
  assign \new_[49864]_  = A201 & A200;
  assign \new_[49867]_  = ~A235 & ~A234;
  assign \new_[49868]_  = \new_[49867]_  & \new_[49864]_ ;
  assign \new_[49869]_  = \new_[49868]_  & \new_[49861]_ ;
  assign \new_[49872]_  = A265 & ~A236;
  assign \new_[49875]_  = ~A267 & A266;
  assign \new_[49876]_  = \new_[49875]_  & \new_[49872]_ ;
  assign \new_[49879]_  = ~A298 & ~A268;
  assign \new_[49882]_  = ~A301 & ~A299;
  assign \new_[49883]_  = \new_[49882]_  & \new_[49879]_ ;
  assign \new_[49884]_  = \new_[49883]_  & \new_[49876]_ ;
  assign \new_[49887]_  = ~A168 & ~A169;
  assign \new_[49890]_  = A166 & A167;
  assign \new_[49891]_  = \new_[49890]_  & \new_[49887]_ ;
  assign \new_[49894]_  = A201 & A200;
  assign \new_[49897]_  = ~A235 & ~A234;
  assign \new_[49898]_  = \new_[49897]_  & \new_[49894]_ ;
  assign \new_[49899]_  = \new_[49898]_  & \new_[49891]_ ;
  assign \new_[49902]_  = ~A265 & ~A236;
  assign \new_[49905]_  = ~A268 & ~A266;
  assign \new_[49906]_  = \new_[49905]_  & \new_[49902]_ ;
  assign \new_[49909]_  = A299 & A298;
  assign \new_[49912]_  = ~A301 & ~A300;
  assign \new_[49913]_  = \new_[49912]_  & \new_[49909]_ ;
  assign \new_[49914]_  = \new_[49913]_  & \new_[49906]_ ;
  assign \new_[49917]_  = ~A168 & ~A169;
  assign \new_[49920]_  = A166 & A167;
  assign \new_[49921]_  = \new_[49920]_  & \new_[49917]_ ;
  assign \new_[49924]_  = A201 & A200;
  assign \new_[49927]_  = A233 & A232;
  assign \new_[49928]_  = \new_[49927]_  & \new_[49924]_ ;
  assign \new_[49929]_  = \new_[49928]_  & \new_[49921]_ ;
  assign \new_[49932]_  = ~A235 & ~A234;
  assign \new_[49935]_  = ~A268 & ~A267;
  assign \new_[49936]_  = \new_[49935]_  & \new_[49932]_ ;
  assign \new_[49939]_  = ~A300 & ~A269;
  assign \new_[49942]_  = ~A302 & ~A301;
  assign \new_[49943]_  = \new_[49942]_  & \new_[49939]_ ;
  assign \new_[49944]_  = \new_[49943]_  & \new_[49936]_ ;
  assign \new_[49947]_  = ~A168 & ~A169;
  assign \new_[49950]_  = A166 & A167;
  assign \new_[49951]_  = \new_[49950]_  & \new_[49947]_ ;
  assign \new_[49954]_  = A201 & A200;
  assign \new_[49957]_  = A233 & A232;
  assign \new_[49958]_  = \new_[49957]_  & \new_[49954]_ ;
  assign \new_[49959]_  = \new_[49958]_  & \new_[49951]_ ;
  assign \new_[49962]_  = ~A235 & ~A234;
  assign \new_[49965]_  = ~A268 & ~A267;
  assign \new_[49966]_  = \new_[49965]_  & \new_[49962]_ ;
  assign \new_[49969]_  = ~A298 & ~A269;
  assign \new_[49972]_  = ~A301 & ~A299;
  assign \new_[49973]_  = \new_[49972]_  & \new_[49969]_ ;
  assign \new_[49974]_  = \new_[49973]_  & \new_[49966]_ ;
  assign \new_[49977]_  = ~A168 & ~A169;
  assign \new_[49980]_  = A166 & A167;
  assign \new_[49981]_  = \new_[49980]_  & \new_[49977]_ ;
  assign \new_[49984]_  = A201 & A200;
  assign \new_[49987]_  = A233 & A232;
  assign \new_[49988]_  = \new_[49987]_  & \new_[49984]_ ;
  assign \new_[49989]_  = \new_[49988]_  & \new_[49981]_ ;
  assign \new_[49992]_  = ~A235 & ~A234;
  assign \new_[49995]_  = ~A266 & ~A265;
  assign \new_[49996]_  = \new_[49995]_  & \new_[49992]_ ;
  assign \new_[49999]_  = ~A300 & ~A268;
  assign \new_[50002]_  = ~A302 & ~A301;
  assign \new_[50003]_  = \new_[50002]_  & \new_[49999]_ ;
  assign \new_[50004]_  = \new_[50003]_  & \new_[49996]_ ;
  assign \new_[50007]_  = ~A168 & ~A169;
  assign \new_[50010]_  = A166 & A167;
  assign \new_[50011]_  = \new_[50010]_  & \new_[50007]_ ;
  assign \new_[50014]_  = A201 & A200;
  assign \new_[50017]_  = A233 & A232;
  assign \new_[50018]_  = \new_[50017]_  & \new_[50014]_ ;
  assign \new_[50019]_  = \new_[50018]_  & \new_[50011]_ ;
  assign \new_[50022]_  = ~A235 & ~A234;
  assign \new_[50025]_  = ~A266 & ~A265;
  assign \new_[50026]_  = \new_[50025]_  & \new_[50022]_ ;
  assign \new_[50029]_  = ~A298 & ~A268;
  assign \new_[50032]_  = ~A301 & ~A299;
  assign \new_[50033]_  = \new_[50032]_  & \new_[50029]_ ;
  assign \new_[50034]_  = \new_[50033]_  & \new_[50026]_ ;
  assign \new_[50037]_  = ~A168 & ~A169;
  assign \new_[50040]_  = A166 & A167;
  assign \new_[50041]_  = \new_[50040]_  & \new_[50037]_ ;
  assign \new_[50044]_  = A201 & A200;
  assign \new_[50047]_  = ~A233 & ~A232;
  assign \new_[50048]_  = \new_[50047]_  & \new_[50044]_ ;
  assign \new_[50049]_  = \new_[50048]_  & \new_[50041]_ ;
  assign \new_[50052]_  = ~A267 & ~A235;
  assign \new_[50055]_  = ~A269 & ~A268;
  assign \new_[50056]_  = \new_[50055]_  & \new_[50052]_ ;
  assign \new_[50059]_  = A299 & A298;
  assign \new_[50062]_  = ~A301 & ~A300;
  assign \new_[50063]_  = \new_[50062]_  & \new_[50059]_ ;
  assign \new_[50064]_  = \new_[50063]_  & \new_[50056]_ ;
  assign \new_[50067]_  = ~A168 & ~A169;
  assign \new_[50070]_  = A166 & A167;
  assign \new_[50071]_  = \new_[50070]_  & \new_[50067]_ ;
  assign \new_[50074]_  = A201 & A200;
  assign \new_[50077]_  = ~A233 & ~A232;
  assign \new_[50078]_  = \new_[50077]_  & \new_[50074]_ ;
  assign \new_[50079]_  = \new_[50078]_  & \new_[50071]_ ;
  assign \new_[50082]_  = A265 & ~A235;
  assign \new_[50085]_  = ~A267 & A266;
  assign \new_[50086]_  = \new_[50085]_  & \new_[50082]_ ;
  assign \new_[50089]_  = ~A300 & ~A268;
  assign \new_[50092]_  = ~A302 & ~A301;
  assign \new_[50093]_  = \new_[50092]_  & \new_[50089]_ ;
  assign \new_[50094]_  = \new_[50093]_  & \new_[50086]_ ;
  assign \new_[50097]_  = ~A168 & ~A169;
  assign \new_[50100]_  = A166 & A167;
  assign \new_[50101]_  = \new_[50100]_  & \new_[50097]_ ;
  assign \new_[50104]_  = A201 & A200;
  assign \new_[50107]_  = ~A233 & ~A232;
  assign \new_[50108]_  = \new_[50107]_  & \new_[50104]_ ;
  assign \new_[50109]_  = \new_[50108]_  & \new_[50101]_ ;
  assign \new_[50112]_  = A265 & ~A235;
  assign \new_[50115]_  = ~A267 & A266;
  assign \new_[50116]_  = \new_[50115]_  & \new_[50112]_ ;
  assign \new_[50119]_  = ~A298 & ~A268;
  assign \new_[50122]_  = ~A301 & ~A299;
  assign \new_[50123]_  = \new_[50122]_  & \new_[50119]_ ;
  assign \new_[50124]_  = \new_[50123]_  & \new_[50116]_ ;
  assign \new_[50127]_  = ~A168 & ~A169;
  assign \new_[50130]_  = A166 & A167;
  assign \new_[50131]_  = \new_[50130]_  & \new_[50127]_ ;
  assign \new_[50134]_  = A201 & A200;
  assign \new_[50137]_  = ~A233 & ~A232;
  assign \new_[50138]_  = \new_[50137]_  & \new_[50134]_ ;
  assign \new_[50139]_  = \new_[50138]_  & \new_[50131]_ ;
  assign \new_[50142]_  = ~A265 & ~A235;
  assign \new_[50145]_  = ~A268 & ~A266;
  assign \new_[50146]_  = \new_[50145]_  & \new_[50142]_ ;
  assign \new_[50149]_  = A299 & A298;
  assign \new_[50152]_  = ~A301 & ~A300;
  assign \new_[50153]_  = \new_[50152]_  & \new_[50149]_ ;
  assign \new_[50154]_  = \new_[50153]_  & \new_[50146]_ ;
  assign \new_[50157]_  = ~A168 & ~A169;
  assign \new_[50160]_  = A166 & A167;
  assign \new_[50161]_  = \new_[50160]_  & \new_[50157]_ ;
  assign \new_[50164]_  = A200 & ~A199;
  assign \new_[50167]_  = ~A234 & A203;
  assign \new_[50168]_  = \new_[50167]_  & \new_[50164]_ ;
  assign \new_[50169]_  = \new_[50168]_  & \new_[50161]_ ;
  assign \new_[50172]_  = ~A236 & ~A235;
  assign \new_[50175]_  = ~A268 & ~A267;
  assign \new_[50176]_  = \new_[50175]_  & \new_[50172]_ ;
  assign \new_[50179]_  = ~A300 & ~A269;
  assign \new_[50182]_  = ~A302 & ~A301;
  assign \new_[50183]_  = \new_[50182]_  & \new_[50179]_ ;
  assign \new_[50184]_  = \new_[50183]_  & \new_[50176]_ ;
  assign \new_[50187]_  = ~A168 & ~A169;
  assign \new_[50190]_  = A166 & A167;
  assign \new_[50191]_  = \new_[50190]_  & \new_[50187]_ ;
  assign \new_[50194]_  = A200 & ~A199;
  assign \new_[50197]_  = ~A234 & A203;
  assign \new_[50198]_  = \new_[50197]_  & \new_[50194]_ ;
  assign \new_[50199]_  = \new_[50198]_  & \new_[50191]_ ;
  assign \new_[50202]_  = ~A236 & ~A235;
  assign \new_[50205]_  = ~A268 & ~A267;
  assign \new_[50206]_  = \new_[50205]_  & \new_[50202]_ ;
  assign \new_[50209]_  = ~A298 & ~A269;
  assign \new_[50212]_  = ~A301 & ~A299;
  assign \new_[50213]_  = \new_[50212]_  & \new_[50209]_ ;
  assign \new_[50214]_  = \new_[50213]_  & \new_[50206]_ ;
  assign \new_[50217]_  = ~A168 & ~A169;
  assign \new_[50220]_  = A166 & A167;
  assign \new_[50221]_  = \new_[50220]_  & \new_[50217]_ ;
  assign \new_[50224]_  = A200 & ~A199;
  assign \new_[50227]_  = ~A234 & A203;
  assign \new_[50228]_  = \new_[50227]_  & \new_[50224]_ ;
  assign \new_[50229]_  = \new_[50228]_  & \new_[50221]_ ;
  assign \new_[50232]_  = ~A236 & ~A235;
  assign \new_[50235]_  = ~A266 & ~A265;
  assign \new_[50236]_  = \new_[50235]_  & \new_[50232]_ ;
  assign \new_[50239]_  = ~A300 & ~A268;
  assign \new_[50242]_  = ~A302 & ~A301;
  assign \new_[50243]_  = \new_[50242]_  & \new_[50239]_ ;
  assign \new_[50244]_  = \new_[50243]_  & \new_[50236]_ ;
  assign \new_[50247]_  = ~A168 & ~A169;
  assign \new_[50250]_  = A166 & A167;
  assign \new_[50251]_  = \new_[50250]_  & \new_[50247]_ ;
  assign \new_[50254]_  = A200 & ~A199;
  assign \new_[50257]_  = ~A234 & A203;
  assign \new_[50258]_  = \new_[50257]_  & \new_[50254]_ ;
  assign \new_[50259]_  = \new_[50258]_  & \new_[50251]_ ;
  assign \new_[50262]_  = ~A236 & ~A235;
  assign \new_[50265]_  = ~A266 & ~A265;
  assign \new_[50266]_  = \new_[50265]_  & \new_[50262]_ ;
  assign \new_[50269]_  = ~A298 & ~A268;
  assign \new_[50272]_  = ~A301 & ~A299;
  assign \new_[50273]_  = \new_[50272]_  & \new_[50269]_ ;
  assign \new_[50274]_  = \new_[50273]_  & \new_[50266]_ ;
  assign \new_[50277]_  = ~A168 & ~A169;
  assign \new_[50280]_  = A166 & A167;
  assign \new_[50281]_  = \new_[50280]_  & \new_[50277]_ ;
  assign \new_[50284]_  = A200 & ~A199;
  assign \new_[50287]_  = ~A232 & A203;
  assign \new_[50288]_  = \new_[50287]_  & \new_[50284]_ ;
  assign \new_[50289]_  = \new_[50288]_  & \new_[50281]_ ;
  assign \new_[50292]_  = ~A235 & ~A233;
  assign \new_[50295]_  = ~A268 & ~A267;
  assign \new_[50296]_  = \new_[50295]_  & \new_[50292]_ ;
  assign \new_[50299]_  = ~A300 & ~A269;
  assign \new_[50302]_  = ~A302 & ~A301;
  assign \new_[50303]_  = \new_[50302]_  & \new_[50299]_ ;
  assign \new_[50304]_  = \new_[50303]_  & \new_[50296]_ ;
  assign \new_[50307]_  = ~A168 & ~A169;
  assign \new_[50310]_  = A166 & A167;
  assign \new_[50311]_  = \new_[50310]_  & \new_[50307]_ ;
  assign \new_[50314]_  = A200 & ~A199;
  assign \new_[50317]_  = ~A232 & A203;
  assign \new_[50318]_  = \new_[50317]_  & \new_[50314]_ ;
  assign \new_[50319]_  = \new_[50318]_  & \new_[50311]_ ;
  assign \new_[50322]_  = ~A235 & ~A233;
  assign \new_[50325]_  = ~A268 & ~A267;
  assign \new_[50326]_  = \new_[50325]_  & \new_[50322]_ ;
  assign \new_[50329]_  = ~A298 & ~A269;
  assign \new_[50332]_  = ~A301 & ~A299;
  assign \new_[50333]_  = \new_[50332]_  & \new_[50329]_ ;
  assign \new_[50334]_  = \new_[50333]_  & \new_[50326]_ ;
  assign \new_[50337]_  = ~A168 & ~A169;
  assign \new_[50340]_  = A166 & A167;
  assign \new_[50341]_  = \new_[50340]_  & \new_[50337]_ ;
  assign \new_[50344]_  = A200 & ~A199;
  assign \new_[50347]_  = ~A232 & A203;
  assign \new_[50348]_  = \new_[50347]_  & \new_[50344]_ ;
  assign \new_[50349]_  = \new_[50348]_  & \new_[50341]_ ;
  assign \new_[50352]_  = ~A235 & ~A233;
  assign \new_[50355]_  = ~A266 & ~A265;
  assign \new_[50356]_  = \new_[50355]_  & \new_[50352]_ ;
  assign \new_[50359]_  = ~A300 & ~A268;
  assign \new_[50362]_  = ~A302 & ~A301;
  assign \new_[50363]_  = \new_[50362]_  & \new_[50359]_ ;
  assign \new_[50364]_  = \new_[50363]_  & \new_[50356]_ ;
  assign \new_[50367]_  = ~A168 & ~A169;
  assign \new_[50370]_  = A166 & A167;
  assign \new_[50371]_  = \new_[50370]_  & \new_[50367]_ ;
  assign \new_[50374]_  = A200 & ~A199;
  assign \new_[50377]_  = ~A232 & A203;
  assign \new_[50378]_  = \new_[50377]_  & \new_[50374]_ ;
  assign \new_[50379]_  = \new_[50378]_  & \new_[50371]_ ;
  assign \new_[50382]_  = ~A235 & ~A233;
  assign \new_[50385]_  = ~A266 & ~A265;
  assign \new_[50386]_  = \new_[50385]_  & \new_[50382]_ ;
  assign \new_[50389]_  = ~A298 & ~A268;
  assign \new_[50392]_  = ~A301 & ~A299;
  assign \new_[50393]_  = \new_[50392]_  & \new_[50389]_ ;
  assign \new_[50394]_  = \new_[50393]_  & \new_[50386]_ ;
  assign \new_[50397]_  = ~A168 & ~A169;
  assign \new_[50400]_  = A166 & A167;
  assign \new_[50401]_  = \new_[50400]_  & \new_[50397]_ ;
  assign \new_[50404]_  = ~A200 & A199;
  assign \new_[50407]_  = ~A234 & A203;
  assign \new_[50408]_  = \new_[50407]_  & \new_[50404]_ ;
  assign \new_[50409]_  = \new_[50408]_  & \new_[50401]_ ;
  assign \new_[50412]_  = ~A236 & ~A235;
  assign \new_[50415]_  = ~A268 & ~A267;
  assign \new_[50416]_  = \new_[50415]_  & \new_[50412]_ ;
  assign \new_[50419]_  = ~A300 & ~A269;
  assign \new_[50422]_  = ~A302 & ~A301;
  assign \new_[50423]_  = \new_[50422]_  & \new_[50419]_ ;
  assign \new_[50424]_  = \new_[50423]_  & \new_[50416]_ ;
  assign \new_[50427]_  = ~A168 & ~A169;
  assign \new_[50430]_  = A166 & A167;
  assign \new_[50431]_  = \new_[50430]_  & \new_[50427]_ ;
  assign \new_[50434]_  = ~A200 & A199;
  assign \new_[50437]_  = ~A234 & A203;
  assign \new_[50438]_  = \new_[50437]_  & \new_[50434]_ ;
  assign \new_[50439]_  = \new_[50438]_  & \new_[50431]_ ;
  assign \new_[50442]_  = ~A236 & ~A235;
  assign \new_[50445]_  = ~A268 & ~A267;
  assign \new_[50446]_  = \new_[50445]_  & \new_[50442]_ ;
  assign \new_[50449]_  = ~A298 & ~A269;
  assign \new_[50452]_  = ~A301 & ~A299;
  assign \new_[50453]_  = \new_[50452]_  & \new_[50449]_ ;
  assign \new_[50454]_  = \new_[50453]_  & \new_[50446]_ ;
  assign \new_[50457]_  = ~A168 & ~A169;
  assign \new_[50460]_  = A166 & A167;
  assign \new_[50461]_  = \new_[50460]_  & \new_[50457]_ ;
  assign \new_[50464]_  = ~A200 & A199;
  assign \new_[50467]_  = ~A234 & A203;
  assign \new_[50468]_  = \new_[50467]_  & \new_[50464]_ ;
  assign \new_[50469]_  = \new_[50468]_  & \new_[50461]_ ;
  assign \new_[50472]_  = ~A236 & ~A235;
  assign \new_[50475]_  = ~A266 & ~A265;
  assign \new_[50476]_  = \new_[50475]_  & \new_[50472]_ ;
  assign \new_[50479]_  = ~A300 & ~A268;
  assign \new_[50482]_  = ~A302 & ~A301;
  assign \new_[50483]_  = \new_[50482]_  & \new_[50479]_ ;
  assign \new_[50484]_  = \new_[50483]_  & \new_[50476]_ ;
  assign \new_[50487]_  = ~A168 & ~A169;
  assign \new_[50490]_  = A166 & A167;
  assign \new_[50491]_  = \new_[50490]_  & \new_[50487]_ ;
  assign \new_[50494]_  = ~A200 & A199;
  assign \new_[50497]_  = ~A234 & A203;
  assign \new_[50498]_  = \new_[50497]_  & \new_[50494]_ ;
  assign \new_[50499]_  = \new_[50498]_  & \new_[50491]_ ;
  assign \new_[50502]_  = ~A236 & ~A235;
  assign \new_[50505]_  = ~A266 & ~A265;
  assign \new_[50506]_  = \new_[50505]_  & \new_[50502]_ ;
  assign \new_[50509]_  = ~A298 & ~A268;
  assign \new_[50512]_  = ~A301 & ~A299;
  assign \new_[50513]_  = \new_[50512]_  & \new_[50509]_ ;
  assign \new_[50514]_  = \new_[50513]_  & \new_[50506]_ ;
  assign \new_[50517]_  = ~A168 & ~A169;
  assign \new_[50520]_  = A166 & A167;
  assign \new_[50521]_  = \new_[50520]_  & \new_[50517]_ ;
  assign \new_[50524]_  = ~A200 & A199;
  assign \new_[50527]_  = ~A232 & A203;
  assign \new_[50528]_  = \new_[50527]_  & \new_[50524]_ ;
  assign \new_[50529]_  = \new_[50528]_  & \new_[50521]_ ;
  assign \new_[50532]_  = ~A235 & ~A233;
  assign \new_[50535]_  = ~A268 & ~A267;
  assign \new_[50536]_  = \new_[50535]_  & \new_[50532]_ ;
  assign \new_[50539]_  = ~A300 & ~A269;
  assign \new_[50542]_  = ~A302 & ~A301;
  assign \new_[50543]_  = \new_[50542]_  & \new_[50539]_ ;
  assign \new_[50544]_  = \new_[50543]_  & \new_[50536]_ ;
  assign \new_[50547]_  = ~A168 & ~A169;
  assign \new_[50550]_  = A166 & A167;
  assign \new_[50551]_  = \new_[50550]_  & \new_[50547]_ ;
  assign \new_[50554]_  = ~A200 & A199;
  assign \new_[50557]_  = ~A232 & A203;
  assign \new_[50558]_  = \new_[50557]_  & \new_[50554]_ ;
  assign \new_[50559]_  = \new_[50558]_  & \new_[50551]_ ;
  assign \new_[50562]_  = ~A235 & ~A233;
  assign \new_[50565]_  = ~A268 & ~A267;
  assign \new_[50566]_  = \new_[50565]_  & \new_[50562]_ ;
  assign \new_[50569]_  = ~A298 & ~A269;
  assign \new_[50572]_  = ~A301 & ~A299;
  assign \new_[50573]_  = \new_[50572]_  & \new_[50569]_ ;
  assign \new_[50574]_  = \new_[50573]_  & \new_[50566]_ ;
  assign \new_[50577]_  = ~A168 & ~A169;
  assign \new_[50580]_  = A166 & A167;
  assign \new_[50581]_  = \new_[50580]_  & \new_[50577]_ ;
  assign \new_[50584]_  = ~A200 & A199;
  assign \new_[50587]_  = ~A232 & A203;
  assign \new_[50588]_  = \new_[50587]_  & \new_[50584]_ ;
  assign \new_[50589]_  = \new_[50588]_  & \new_[50581]_ ;
  assign \new_[50592]_  = ~A235 & ~A233;
  assign \new_[50595]_  = ~A266 & ~A265;
  assign \new_[50596]_  = \new_[50595]_  & \new_[50592]_ ;
  assign \new_[50599]_  = ~A300 & ~A268;
  assign \new_[50602]_  = ~A302 & ~A301;
  assign \new_[50603]_  = \new_[50602]_  & \new_[50599]_ ;
  assign \new_[50604]_  = \new_[50603]_  & \new_[50596]_ ;
  assign \new_[50607]_  = ~A168 & ~A169;
  assign \new_[50610]_  = A166 & A167;
  assign \new_[50611]_  = \new_[50610]_  & \new_[50607]_ ;
  assign \new_[50614]_  = ~A200 & A199;
  assign \new_[50617]_  = ~A232 & A203;
  assign \new_[50618]_  = \new_[50617]_  & \new_[50614]_ ;
  assign \new_[50619]_  = \new_[50618]_  & \new_[50611]_ ;
  assign \new_[50622]_  = ~A235 & ~A233;
  assign \new_[50625]_  = ~A266 & ~A265;
  assign \new_[50626]_  = \new_[50625]_  & \new_[50622]_ ;
  assign \new_[50629]_  = ~A298 & ~A268;
  assign \new_[50632]_  = ~A301 & ~A299;
  assign \new_[50633]_  = \new_[50632]_  & \new_[50629]_ ;
  assign \new_[50634]_  = \new_[50633]_  & \new_[50626]_ ;
  assign \new_[50637]_  = ~A169 & ~A170;
  assign \new_[50640]_  = A202 & ~A168;
  assign \new_[50641]_  = \new_[50640]_  & \new_[50637]_ ;
  assign \new_[50644]_  = A233 & A232;
  assign \new_[50647]_  = ~A235 & ~A234;
  assign \new_[50648]_  = \new_[50647]_  & \new_[50644]_ ;
  assign \new_[50649]_  = \new_[50648]_  & \new_[50641]_ ;
  assign \new_[50652]_  = A266 & A265;
  assign \new_[50655]_  = ~A268 & ~A267;
  assign \new_[50656]_  = \new_[50655]_  & \new_[50652]_ ;
  assign \new_[50659]_  = A299 & A298;
  assign \new_[50662]_  = ~A301 & ~A300;
  assign \new_[50663]_  = \new_[50662]_  & \new_[50659]_ ;
  assign \new_[50664]_  = \new_[50663]_  & \new_[50656]_ ;
  assign \new_[50667]_  = ~A169 & ~A170;
  assign \new_[50670]_  = A199 & ~A168;
  assign \new_[50671]_  = \new_[50670]_  & \new_[50667]_ ;
  assign \new_[50674]_  = ~A234 & A201;
  assign \new_[50677]_  = ~A236 & ~A235;
  assign \new_[50678]_  = \new_[50677]_  & \new_[50674]_ ;
  assign \new_[50679]_  = \new_[50678]_  & \new_[50671]_ ;
  assign \new_[50682]_  = A266 & A265;
  assign \new_[50685]_  = ~A268 & ~A267;
  assign \new_[50686]_  = \new_[50685]_  & \new_[50682]_ ;
  assign \new_[50689]_  = A299 & A298;
  assign \new_[50692]_  = ~A301 & ~A300;
  assign \new_[50693]_  = \new_[50692]_  & \new_[50689]_ ;
  assign \new_[50694]_  = \new_[50693]_  & \new_[50686]_ ;
  assign \new_[50697]_  = ~A169 & ~A170;
  assign \new_[50700]_  = A199 & ~A168;
  assign \new_[50701]_  = \new_[50700]_  & \new_[50697]_ ;
  assign \new_[50704]_  = A232 & A201;
  assign \new_[50707]_  = ~A234 & A233;
  assign \new_[50708]_  = \new_[50707]_  & \new_[50704]_ ;
  assign \new_[50709]_  = \new_[50708]_  & \new_[50701]_ ;
  assign \new_[50712]_  = ~A267 & ~A235;
  assign \new_[50715]_  = ~A269 & ~A268;
  assign \new_[50716]_  = \new_[50715]_  & \new_[50712]_ ;
  assign \new_[50719]_  = A299 & A298;
  assign \new_[50722]_  = ~A301 & ~A300;
  assign \new_[50723]_  = \new_[50722]_  & \new_[50719]_ ;
  assign \new_[50724]_  = \new_[50723]_  & \new_[50716]_ ;
  assign \new_[50727]_  = ~A169 & ~A170;
  assign \new_[50730]_  = A199 & ~A168;
  assign \new_[50731]_  = \new_[50730]_  & \new_[50727]_ ;
  assign \new_[50734]_  = A232 & A201;
  assign \new_[50737]_  = ~A234 & A233;
  assign \new_[50738]_  = \new_[50737]_  & \new_[50734]_ ;
  assign \new_[50739]_  = \new_[50738]_  & \new_[50731]_ ;
  assign \new_[50742]_  = A265 & ~A235;
  assign \new_[50745]_  = ~A267 & A266;
  assign \new_[50746]_  = \new_[50745]_  & \new_[50742]_ ;
  assign \new_[50749]_  = ~A300 & ~A268;
  assign \new_[50752]_  = ~A302 & ~A301;
  assign \new_[50753]_  = \new_[50752]_  & \new_[50749]_ ;
  assign \new_[50754]_  = \new_[50753]_  & \new_[50746]_ ;
  assign \new_[50757]_  = ~A169 & ~A170;
  assign \new_[50760]_  = A199 & ~A168;
  assign \new_[50761]_  = \new_[50760]_  & \new_[50757]_ ;
  assign \new_[50764]_  = A232 & A201;
  assign \new_[50767]_  = ~A234 & A233;
  assign \new_[50768]_  = \new_[50767]_  & \new_[50764]_ ;
  assign \new_[50769]_  = \new_[50768]_  & \new_[50761]_ ;
  assign \new_[50772]_  = A265 & ~A235;
  assign \new_[50775]_  = ~A267 & A266;
  assign \new_[50776]_  = \new_[50775]_  & \new_[50772]_ ;
  assign \new_[50779]_  = ~A298 & ~A268;
  assign \new_[50782]_  = ~A301 & ~A299;
  assign \new_[50783]_  = \new_[50782]_  & \new_[50779]_ ;
  assign \new_[50784]_  = \new_[50783]_  & \new_[50776]_ ;
  assign \new_[50787]_  = ~A169 & ~A170;
  assign \new_[50790]_  = A199 & ~A168;
  assign \new_[50791]_  = \new_[50790]_  & \new_[50787]_ ;
  assign \new_[50794]_  = A232 & A201;
  assign \new_[50797]_  = ~A234 & A233;
  assign \new_[50798]_  = \new_[50797]_  & \new_[50794]_ ;
  assign \new_[50799]_  = \new_[50798]_  & \new_[50791]_ ;
  assign \new_[50802]_  = ~A265 & ~A235;
  assign \new_[50805]_  = ~A268 & ~A266;
  assign \new_[50806]_  = \new_[50805]_  & \new_[50802]_ ;
  assign \new_[50809]_  = A299 & A298;
  assign \new_[50812]_  = ~A301 & ~A300;
  assign \new_[50813]_  = \new_[50812]_  & \new_[50809]_ ;
  assign \new_[50814]_  = \new_[50813]_  & \new_[50806]_ ;
  assign \new_[50817]_  = ~A169 & ~A170;
  assign \new_[50820]_  = A199 & ~A168;
  assign \new_[50821]_  = \new_[50820]_  & \new_[50817]_ ;
  assign \new_[50824]_  = ~A232 & A201;
  assign \new_[50827]_  = ~A235 & ~A233;
  assign \new_[50828]_  = \new_[50827]_  & \new_[50824]_ ;
  assign \new_[50829]_  = \new_[50828]_  & \new_[50821]_ ;
  assign \new_[50832]_  = A266 & A265;
  assign \new_[50835]_  = ~A268 & ~A267;
  assign \new_[50836]_  = \new_[50835]_  & \new_[50832]_ ;
  assign \new_[50839]_  = A299 & A298;
  assign \new_[50842]_  = ~A301 & ~A300;
  assign \new_[50843]_  = \new_[50842]_  & \new_[50839]_ ;
  assign \new_[50844]_  = \new_[50843]_  & \new_[50836]_ ;
  assign \new_[50847]_  = ~A169 & ~A170;
  assign \new_[50850]_  = A200 & ~A168;
  assign \new_[50851]_  = \new_[50850]_  & \new_[50847]_ ;
  assign \new_[50854]_  = ~A234 & A201;
  assign \new_[50857]_  = ~A236 & ~A235;
  assign \new_[50858]_  = \new_[50857]_  & \new_[50854]_ ;
  assign \new_[50859]_  = \new_[50858]_  & \new_[50851]_ ;
  assign \new_[50862]_  = A266 & A265;
  assign \new_[50865]_  = ~A268 & ~A267;
  assign \new_[50866]_  = \new_[50865]_  & \new_[50862]_ ;
  assign \new_[50869]_  = A299 & A298;
  assign \new_[50872]_  = ~A301 & ~A300;
  assign \new_[50873]_  = \new_[50872]_  & \new_[50869]_ ;
  assign \new_[50874]_  = \new_[50873]_  & \new_[50866]_ ;
  assign \new_[50877]_  = ~A169 & ~A170;
  assign \new_[50880]_  = A200 & ~A168;
  assign \new_[50881]_  = \new_[50880]_  & \new_[50877]_ ;
  assign \new_[50884]_  = A232 & A201;
  assign \new_[50887]_  = ~A234 & A233;
  assign \new_[50888]_  = \new_[50887]_  & \new_[50884]_ ;
  assign \new_[50889]_  = \new_[50888]_  & \new_[50881]_ ;
  assign \new_[50892]_  = ~A267 & ~A235;
  assign \new_[50895]_  = ~A269 & ~A268;
  assign \new_[50896]_  = \new_[50895]_  & \new_[50892]_ ;
  assign \new_[50899]_  = A299 & A298;
  assign \new_[50902]_  = ~A301 & ~A300;
  assign \new_[50903]_  = \new_[50902]_  & \new_[50899]_ ;
  assign \new_[50904]_  = \new_[50903]_  & \new_[50896]_ ;
  assign \new_[50907]_  = ~A169 & ~A170;
  assign \new_[50910]_  = A200 & ~A168;
  assign \new_[50911]_  = \new_[50910]_  & \new_[50907]_ ;
  assign \new_[50914]_  = A232 & A201;
  assign \new_[50917]_  = ~A234 & A233;
  assign \new_[50918]_  = \new_[50917]_  & \new_[50914]_ ;
  assign \new_[50919]_  = \new_[50918]_  & \new_[50911]_ ;
  assign \new_[50922]_  = A265 & ~A235;
  assign \new_[50925]_  = ~A267 & A266;
  assign \new_[50926]_  = \new_[50925]_  & \new_[50922]_ ;
  assign \new_[50929]_  = ~A300 & ~A268;
  assign \new_[50932]_  = ~A302 & ~A301;
  assign \new_[50933]_  = \new_[50932]_  & \new_[50929]_ ;
  assign \new_[50934]_  = \new_[50933]_  & \new_[50926]_ ;
  assign \new_[50937]_  = ~A169 & ~A170;
  assign \new_[50940]_  = A200 & ~A168;
  assign \new_[50941]_  = \new_[50940]_  & \new_[50937]_ ;
  assign \new_[50944]_  = A232 & A201;
  assign \new_[50947]_  = ~A234 & A233;
  assign \new_[50948]_  = \new_[50947]_  & \new_[50944]_ ;
  assign \new_[50949]_  = \new_[50948]_  & \new_[50941]_ ;
  assign \new_[50952]_  = A265 & ~A235;
  assign \new_[50955]_  = ~A267 & A266;
  assign \new_[50956]_  = \new_[50955]_  & \new_[50952]_ ;
  assign \new_[50959]_  = ~A298 & ~A268;
  assign \new_[50962]_  = ~A301 & ~A299;
  assign \new_[50963]_  = \new_[50962]_  & \new_[50959]_ ;
  assign \new_[50964]_  = \new_[50963]_  & \new_[50956]_ ;
  assign \new_[50967]_  = ~A169 & ~A170;
  assign \new_[50970]_  = A200 & ~A168;
  assign \new_[50971]_  = \new_[50970]_  & \new_[50967]_ ;
  assign \new_[50974]_  = A232 & A201;
  assign \new_[50977]_  = ~A234 & A233;
  assign \new_[50978]_  = \new_[50977]_  & \new_[50974]_ ;
  assign \new_[50979]_  = \new_[50978]_  & \new_[50971]_ ;
  assign \new_[50982]_  = ~A265 & ~A235;
  assign \new_[50985]_  = ~A268 & ~A266;
  assign \new_[50986]_  = \new_[50985]_  & \new_[50982]_ ;
  assign \new_[50989]_  = A299 & A298;
  assign \new_[50992]_  = ~A301 & ~A300;
  assign \new_[50993]_  = \new_[50992]_  & \new_[50989]_ ;
  assign \new_[50994]_  = \new_[50993]_  & \new_[50986]_ ;
  assign \new_[50997]_  = ~A169 & ~A170;
  assign \new_[51000]_  = A200 & ~A168;
  assign \new_[51001]_  = \new_[51000]_  & \new_[50997]_ ;
  assign \new_[51004]_  = ~A232 & A201;
  assign \new_[51007]_  = ~A235 & ~A233;
  assign \new_[51008]_  = \new_[51007]_  & \new_[51004]_ ;
  assign \new_[51009]_  = \new_[51008]_  & \new_[51001]_ ;
  assign \new_[51012]_  = A266 & A265;
  assign \new_[51015]_  = ~A268 & ~A267;
  assign \new_[51016]_  = \new_[51015]_  & \new_[51012]_ ;
  assign \new_[51019]_  = A299 & A298;
  assign \new_[51022]_  = ~A301 & ~A300;
  assign \new_[51023]_  = \new_[51022]_  & \new_[51019]_ ;
  assign \new_[51024]_  = \new_[51023]_  & \new_[51016]_ ;
  assign \new_[51027]_  = ~A169 & ~A170;
  assign \new_[51030]_  = ~A199 & ~A168;
  assign \new_[51031]_  = \new_[51030]_  & \new_[51027]_ ;
  assign \new_[51034]_  = A203 & A200;
  assign \new_[51037]_  = ~A235 & ~A234;
  assign \new_[51038]_  = \new_[51037]_  & \new_[51034]_ ;
  assign \new_[51039]_  = \new_[51038]_  & \new_[51031]_ ;
  assign \new_[51042]_  = ~A267 & ~A236;
  assign \new_[51045]_  = ~A269 & ~A268;
  assign \new_[51046]_  = \new_[51045]_  & \new_[51042]_ ;
  assign \new_[51049]_  = A299 & A298;
  assign \new_[51052]_  = ~A301 & ~A300;
  assign \new_[51053]_  = \new_[51052]_  & \new_[51049]_ ;
  assign \new_[51054]_  = \new_[51053]_  & \new_[51046]_ ;
  assign \new_[51057]_  = ~A169 & ~A170;
  assign \new_[51060]_  = ~A199 & ~A168;
  assign \new_[51061]_  = \new_[51060]_  & \new_[51057]_ ;
  assign \new_[51064]_  = A203 & A200;
  assign \new_[51067]_  = ~A235 & ~A234;
  assign \new_[51068]_  = \new_[51067]_  & \new_[51064]_ ;
  assign \new_[51069]_  = \new_[51068]_  & \new_[51061]_ ;
  assign \new_[51072]_  = A265 & ~A236;
  assign \new_[51075]_  = ~A267 & A266;
  assign \new_[51076]_  = \new_[51075]_  & \new_[51072]_ ;
  assign \new_[51079]_  = ~A300 & ~A268;
  assign \new_[51082]_  = ~A302 & ~A301;
  assign \new_[51083]_  = \new_[51082]_  & \new_[51079]_ ;
  assign \new_[51084]_  = \new_[51083]_  & \new_[51076]_ ;
  assign \new_[51087]_  = ~A169 & ~A170;
  assign \new_[51090]_  = ~A199 & ~A168;
  assign \new_[51091]_  = \new_[51090]_  & \new_[51087]_ ;
  assign \new_[51094]_  = A203 & A200;
  assign \new_[51097]_  = ~A235 & ~A234;
  assign \new_[51098]_  = \new_[51097]_  & \new_[51094]_ ;
  assign \new_[51099]_  = \new_[51098]_  & \new_[51091]_ ;
  assign \new_[51102]_  = A265 & ~A236;
  assign \new_[51105]_  = ~A267 & A266;
  assign \new_[51106]_  = \new_[51105]_  & \new_[51102]_ ;
  assign \new_[51109]_  = ~A298 & ~A268;
  assign \new_[51112]_  = ~A301 & ~A299;
  assign \new_[51113]_  = \new_[51112]_  & \new_[51109]_ ;
  assign \new_[51114]_  = \new_[51113]_  & \new_[51106]_ ;
  assign \new_[51117]_  = ~A169 & ~A170;
  assign \new_[51120]_  = ~A199 & ~A168;
  assign \new_[51121]_  = \new_[51120]_  & \new_[51117]_ ;
  assign \new_[51124]_  = A203 & A200;
  assign \new_[51127]_  = ~A235 & ~A234;
  assign \new_[51128]_  = \new_[51127]_  & \new_[51124]_ ;
  assign \new_[51129]_  = \new_[51128]_  & \new_[51121]_ ;
  assign \new_[51132]_  = ~A265 & ~A236;
  assign \new_[51135]_  = ~A268 & ~A266;
  assign \new_[51136]_  = \new_[51135]_  & \new_[51132]_ ;
  assign \new_[51139]_  = A299 & A298;
  assign \new_[51142]_  = ~A301 & ~A300;
  assign \new_[51143]_  = \new_[51142]_  & \new_[51139]_ ;
  assign \new_[51144]_  = \new_[51143]_  & \new_[51136]_ ;
  assign \new_[51147]_  = ~A169 & ~A170;
  assign \new_[51150]_  = ~A199 & ~A168;
  assign \new_[51151]_  = \new_[51150]_  & \new_[51147]_ ;
  assign \new_[51154]_  = A203 & A200;
  assign \new_[51157]_  = A233 & A232;
  assign \new_[51158]_  = \new_[51157]_  & \new_[51154]_ ;
  assign \new_[51159]_  = \new_[51158]_  & \new_[51151]_ ;
  assign \new_[51162]_  = ~A235 & ~A234;
  assign \new_[51165]_  = ~A268 & ~A267;
  assign \new_[51166]_  = \new_[51165]_  & \new_[51162]_ ;
  assign \new_[51169]_  = ~A300 & ~A269;
  assign \new_[51172]_  = ~A302 & ~A301;
  assign \new_[51173]_  = \new_[51172]_  & \new_[51169]_ ;
  assign \new_[51174]_  = \new_[51173]_  & \new_[51166]_ ;
  assign \new_[51177]_  = ~A169 & ~A170;
  assign \new_[51180]_  = ~A199 & ~A168;
  assign \new_[51181]_  = \new_[51180]_  & \new_[51177]_ ;
  assign \new_[51184]_  = A203 & A200;
  assign \new_[51187]_  = A233 & A232;
  assign \new_[51188]_  = \new_[51187]_  & \new_[51184]_ ;
  assign \new_[51189]_  = \new_[51188]_  & \new_[51181]_ ;
  assign \new_[51192]_  = ~A235 & ~A234;
  assign \new_[51195]_  = ~A268 & ~A267;
  assign \new_[51196]_  = \new_[51195]_  & \new_[51192]_ ;
  assign \new_[51199]_  = ~A298 & ~A269;
  assign \new_[51202]_  = ~A301 & ~A299;
  assign \new_[51203]_  = \new_[51202]_  & \new_[51199]_ ;
  assign \new_[51204]_  = \new_[51203]_  & \new_[51196]_ ;
  assign \new_[51207]_  = ~A169 & ~A170;
  assign \new_[51210]_  = ~A199 & ~A168;
  assign \new_[51211]_  = \new_[51210]_  & \new_[51207]_ ;
  assign \new_[51214]_  = A203 & A200;
  assign \new_[51217]_  = A233 & A232;
  assign \new_[51218]_  = \new_[51217]_  & \new_[51214]_ ;
  assign \new_[51219]_  = \new_[51218]_  & \new_[51211]_ ;
  assign \new_[51222]_  = ~A235 & ~A234;
  assign \new_[51225]_  = ~A266 & ~A265;
  assign \new_[51226]_  = \new_[51225]_  & \new_[51222]_ ;
  assign \new_[51229]_  = ~A300 & ~A268;
  assign \new_[51232]_  = ~A302 & ~A301;
  assign \new_[51233]_  = \new_[51232]_  & \new_[51229]_ ;
  assign \new_[51234]_  = \new_[51233]_  & \new_[51226]_ ;
  assign \new_[51237]_  = ~A169 & ~A170;
  assign \new_[51240]_  = ~A199 & ~A168;
  assign \new_[51241]_  = \new_[51240]_  & \new_[51237]_ ;
  assign \new_[51244]_  = A203 & A200;
  assign \new_[51247]_  = A233 & A232;
  assign \new_[51248]_  = \new_[51247]_  & \new_[51244]_ ;
  assign \new_[51249]_  = \new_[51248]_  & \new_[51241]_ ;
  assign \new_[51252]_  = ~A235 & ~A234;
  assign \new_[51255]_  = ~A266 & ~A265;
  assign \new_[51256]_  = \new_[51255]_  & \new_[51252]_ ;
  assign \new_[51259]_  = ~A298 & ~A268;
  assign \new_[51262]_  = ~A301 & ~A299;
  assign \new_[51263]_  = \new_[51262]_  & \new_[51259]_ ;
  assign \new_[51264]_  = \new_[51263]_  & \new_[51256]_ ;
  assign \new_[51267]_  = ~A169 & ~A170;
  assign \new_[51270]_  = ~A199 & ~A168;
  assign \new_[51271]_  = \new_[51270]_  & \new_[51267]_ ;
  assign \new_[51274]_  = A203 & A200;
  assign \new_[51277]_  = ~A233 & ~A232;
  assign \new_[51278]_  = \new_[51277]_  & \new_[51274]_ ;
  assign \new_[51279]_  = \new_[51278]_  & \new_[51271]_ ;
  assign \new_[51282]_  = ~A267 & ~A235;
  assign \new_[51285]_  = ~A269 & ~A268;
  assign \new_[51286]_  = \new_[51285]_  & \new_[51282]_ ;
  assign \new_[51289]_  = A299 & A298;
  assign \new_[51292]_  = ~A301 & ~A300;
  assign \new_[51293]_  = \new_[51292]_  & \new_[51289]_ ;
  assign \new_[51294]_  = \new_[51293]_  & \new_[51286]_ ;
  assign \new_[51297]_  = ~A169 & ~A170;
  assign \new_[51300]_  = ~A199 & ~A168;
  assign \new_[51301]_  = \new_[51300]_  & \new_[51297]_ ;
  assign \new_[51304]_  = A203 & A200;
  assign \new_[51307]_  = ~A233 & ~A232;
  assign \new_[51308]_  = \new_[51307]_  & \new_[51304]_ ;
  assign \new_[51309]_  = \new_[51308]_  & \new_[51301]_ ;
  assign \new_[51312]_  = A265 & ~A235;
  assign \new_[51315]_  = ~A267 & A266;
  assign \new_[51316]_  = \new_[51315]_  & \new_[51312]_ ;
  assign \new_[51319]_  = ~A300 & ~A268;
  assign \new_[51322]_  = ~A302 & ~A301;
  assign \new_[51323]_  = \new_[51322]_  & \new_[51319]_ ;
  assign \new_[51324]_  = \new_[51323]_  & \new_[51316]_ ;
  assign \new_[51327]_  = ~A169 & ~A170;
  assign \new_[51330]_  = ~A199 & ~A168;
  assign \new_[51331]_  = \new_[51330]_  & \new_[51327]_ ;
  assign \new_[51334]_  = A203 & A200;
  assign \new_[51337]_  = ~A233 & ~A232;
  assign \new_[51338]_  = \new_[51337]_  & \new_[51334]_ ;
  assign \new_[51339]_  = \new_[51338]_  & \new_[51331]_ ;
  assign \new_[51342]_  = A265 & ~A235;
  assign \new_[51345]_  = ~A267 & A266;
  assign \new_[51346]_  = \new_[51345]_  & \new_[51342]_ ;
  assign \new_[51349]_  = ~A298 & ~A268;
  assign \new_[51352]_  = ~A301 & ~A299;
  assign \new_[51353]_  = \new_[51352]_  & \new_[51349]_ ;
  assign \new_[51354]_  = \new_[51353]_  & \new_[51346]_ ;
  assign \new_[51357]_  = ~A169 & ~A170;
  assign \new_[51360]_  = ~A199 & ~A168;
  assign \new_[51361]_  = \new_[51360]_  & \new_[51357]_ ;
  assign \new_[51364]_  = A203 & A200;
  assign \new_[51367]_  = ~A233 & ~A232;
  assign \new_[51368]_  = \new_[51367]_  & \new_[51364]_ ;
  assign \new_[51369]_  = \new_[51368]_  & \new_[51361]_ ;
  assign \new_[51372]_  = ~A265 & ~A235;
  assign \new_[51375]_  = ~A268 & ~A266;
  assign \new_[51376]_  = \new_[51375]_  & \new_[51372]_ ;
  assign \new_[51379]_  = A299 & A298;
  assign \new_[51382]_  = ~A301 & ~A300;
  assign \new_[51383]_  = \new_[51382]_  & \new_[51379]_ ;
  assign \new_[51384]_  = \new_[51383]_  & \new_[51376]_ ;
  assign \new_[51387]_  = ~A169 & ~A170;
  assign \new_[51390]_  = A199 & ~A168;
  assign \new_[51391]_  = \new_[51390]_  & \new_[51387]_ ;
  assign \new_[51394]_  = A203 & ~A200;
  assign \new_[51397]_  = ~A235 & ~A234;
  assign \new_[51398]_  = \new_[51397]_  & \new_[51394]_ ;
  assign \new_[51399]_  = \new_[51398]_  & \new_[51391]_ ;
  assign \new_[51402]_  = ~A267 & ~A236;
  assign \new_[51405]_  = ~A269 & ~A268;
  assign \new_[51406]_  = \new_[51405]_  & \new_[51402]_ ;
  assign \new_[51409]_  = A299 & A298;
  assign \new_[51412]_  = ~A301 & ~A300;
  assign \new_[51413]_  = \new_[51412]_  & \new_[51409]_ ;
  assign \new_[51414]_  = \new_[51413]_  & \new_[51406]_ ;
  assign \new_[51417]_  = ~A169 & ~A170;
  assign \new_[51420]_  = A199 & ~A168;
  assign \new_[51421]_  = \new_[51420]_  & \new_[51417]_ ;
  assign \new_[51424]_  = A203 & ~A200;
  assign \new_[51427]_  = ~A235 & ~A234;
  assign \new_[51428]_  = \new_[51427]_  & \new_[51424]_ ;
  assign \new_[51429]_  = \new_[51428]_  & \new_[51421]_ ;
  assign \new_[51432]_  = A265 & ~A236;
  assign \new_[51435]_  = ~A267 & A266;
  assign \new_[51436]_  = \new_[51435]_  & \new_[51432]_ ;
  assign \new_[51439]_  = ~A300 & ~A268;
  assign \new_[51442]_  = ~A302 & ~A301;
  assign \new_[51443]_  = \new_[51442]_  & \new_[51439]_ ;
  assign \new_[51444]_  = \new_[51443]_  & \new_[51436]_ ;
  assign \new_[51447]_  = ~A169 & ~A170;
  assign \new_[51450]_  = A199 & ~A168;
  assign \new_[51451]_  = \new_[51450]_  & \new_[51447]_ ;
  assign \new_[51454]_  = A203 & ~A200;
  assign \new_[51457]_  = ~A235 & ~A234;
  assign \new_[51458]_  = \new_[51457]_  & \new_[51454]_ ;
  assign \new_[51459]_  = \new_[51458]_  & \new_[51451]_ ;
  assign \new_[51462]_  = A265 & ~A236;
  assign \new_[51465]_  = ~A267 & A266;
  assign \new_[51466]_  = \new_[51465]_  & \new_[51462]_ ;
  assign \new_[51469]_  = ~A298 & ~A268;
  assign \new_[51472]_  = ~A301 & ~A299;
  assign \new_[51473]_  = \new_[51472]_  & \new_[51469]_ ;
  assign \new_[51474]_  = \new_[51473]_  & \new_[51466]_ ;
  assign \new_[51477]_  = ~A169 & ~A170;
  assign \new_[51480]_  = A199 & ~A168;
  assign \new_[51481]_  = \new_[51480]_  & \new_[51477]_ ;
  assign \new_[51484]_  = A203 & ~A200;
  assign \new_[51487]_  = ~A235 & ~A234;
  assign \new_[51488]_  = \new_[51487]_  & \new_[51484]_ ;
  assign \new_[51489]_  = \new_[51488]_  & \new_[51481]_ ;
  assign \new_[51492]_  = ~A265 & ~A236;
  assign \new_[51495]_  = ~A268 & ~A266;
  assign \new_[51496]_  = \new_[51495]_  & \new_[51492]_ ;
  assign \new_[51499]_  = A299 & A298;
  assign \new_[51502]_  = ~A301 & ~A300;
  assign \new_[51503]_  = \new_[51502]_  & \new_[51499]_ ;
  assign \new_[51504]_  = \new_[51503]_  & \new_[51496]_ ;
  assign \new_[51507]_  = ~A169 & ~A170;
  assign \new_[51510]_  = A199 & ~A168;
  assign \new_[51511]_  = \new_[51510]_  & \new_[51507]_ ;
  assign \new_[51514]_  = A203 & ~A200;
  assign \new_[51517]_  = A233 & A232;
  assign \new_[51518]_  = \new_[51517]_  & \new_[51514]_ ;
  assign \new_[51519]_  = \new_[51518]_  & \new_[51511]_ ;
  assign \new_[51522]_  = ~A235 & ~A234;
  assign \new_[51525]_  = ~A268 & ~A267;
  assign \new_[51526]_  = \new_[51525]_  & \new_[51522]_ ;
  assign \new_[51529]_  = ~A300 & ~A269;
  assign \new_[51532]_  = ~A302 & ~A301;
  assign \new_[51533]_  = \new_[51532]_  & \new_[51529]_ ;
  assign \new_[51534]_  = \new_[51533]_  & \new_[51526]_ ;
  assign \new_[51537]_  = ~A169 & ~A170;
  assign \new_[51540]_  = A199 & ~A168;
  assign \new_[51541]_  = \new_[51540]_  & \new_[51537]_ ;
  assign \new_[51544]_  = A203 & ~A200;
  assign \new_[51547]_  = A233 & A232;
  assign \new_[51548]_  = \new_[51547]_  & \new_[51544]_ ;
  assign \new_[51549]_  = \new_[51548]_  & \new_[51541]_ ;
  assign \new_[51552]_  = ~A235 & ~A234;
  assign \new_[51555]_  = ~A268 & ~A267;
  assign \new_[51556]_  = \new_[51555]_  & \new_[51552]_ ;
  assign \new_[51559]_  = ~A298 & ~A269;
  assign \new_[51562]_  = ~A301 & ~A299;
  assign \new_[51563]_  = \new_[51562]_  & \new_[51559]_ ;
  assign \new_[51564]_  = \new_[51563]_  & \new_[51556]_ ;
  assign \new_[51567]_  = ~A169 & ~A170;
  assign \new_[51570]_  = A199 & ~A168;
  assign \new_[51571]_  = \new_[51570]_  & \new_[51567]_ ;
  assign \new_[51574]_  = A203 & ~A200;
  assign \new_[51577]_  = A233 & A232;
  assign \new_[51578]_  = \new_[51577]_  & \new_[51574]_ ;
  assign \new_[51579]_  = \new_[51578]_  & \new_[51571]_ ;
  assign \new_[51582]_  = ~A235 & ~A234;
  assign \new_[51585]_  = ~A266 & ~A265;
  assign \new_[51586]_  = \new_[51585]_  & \new_[51582]_ ;
  assign \new_[51589]_  = ~A300 & ~A268;
  assign \new_[51592]_  = ~A302 & ~A301;
  assign \new_[51593]_  = \new_[51592]_  & \new_[51589]_ ;
  assign \new_[51594]_  = \new_[51593]_  & \new_[51586]_ ;
  assign \new_[51597]_  = ~A169 & ~A170;
  assign \new_[51600]_  = A199 & ~A168;
  assign \new_[51601]_  = \new_[51600]_  & \new_[51597]_ ;
  assign \new_[51604]_  = A203 & ~A200;
  assign \new_[51607]_  = A233 & A232;
  assign \new_[51608]_  = \new_[51607]_  & \new_[51604]_ ;
  assign \new_[51609]_  = \new_[51608]_  & \new_[51601]_ ;
  assign \new_[51612]_  = ~A235 & ~A234;
  assign \new_[51615]_  = ~A266 & ~A265;
  assign \new_[51616]_  = \new_[51615]_  & \new_[51612]_ ;
  assign \new_[51619]_  = ~A298 & ~A268;
  assign \new_[51622]_  = ~A301 & ~A299;
  assign \new_[51623]_  = \new_[51622]_  & \new_[51619]_ ;
  assign \new_[51624]_  = \new_[51623]_  & \new_[51616]_ ;
  assign \new_[51627]_  = ~A169 & ~A170;
  assign \new_[51630]_  = A199 & ~A168;
  assign \new_[51631]_  = \new_[51630]_  & \new_[51627]_ ;
  assign \new_[51634]_  = A203 & ~A200;
  assign \new_[51637]_  = ~A233 & ~A232;
  assign \new_[51638]_  = \new_[51637]_  & \new_[51634]_ ;
  assign \new_[51639]_  = \new_[51638]_  & \new_[51631]_ ;
  assign \new_[51642]_  = ~A267 & ~A235;
  assign \new_[51645]_  = ~A269 & ~A268;
  assign \new_[51646]_  = \new_[51645]_  & \new_[51642]_ ;
  assign \new_[51649]_  = A299 & A298;
  assign \new_[51652]_  = ~A301 & ~A300;
  assign \new_[51653]_  = \new_[51652]_  & \new_[51649]_ ;
  assign \new_[51654]_  = \new_[51653]_  & \new_[51646]_ ;
  assign \new_[51657]_  = ~A169 & ~A170;
  assign \new_[51660]_  = A199 & ~A168;
  assign \new_[51661]_  = \new_[51660]_  & \new_[51657]_ ;
  assign \new_[51664]_  = A203 & ~A200;
  assign \new_[51667]_  = ~A233 & ~A232;
  assign \new_[51668]_  = \new_[51667]_  & \new_[51664]_ ;
  assign \new_[51669]_  = \new_[51668]_  & \new_[51661]_ ;
  assign \new_[51672]_  = A265 & ~A235;
  assign \new_[51675]_  = ~A267 & A266;
  assign \new_[51676]_  = \new_[51675]_  & \new_[51672]_ ;
  assign \new_[51679]_  = ~A300 & ~A268;
  assign \new_[51682]_  = ~A302 & ~A301;
  assign \new_[51683]_  = \new_[51682]_  & \new_[51679]_ ;
  assign \new_[51684]_  = \new_[51683]_  & \new_[51676]_ ;
  assign \new_[51687]_  = ~A169 & ~A170;
  assign \new_[51690]_  = A199 & ~A168;
  assign \new_[51691]_  = \new_[51690]_  & \new_[51687]_ ;
  assign \new_[51694]_  = A203 & ~A200;
  assign \new_[51697]_  = ~A233 & ~A232;
  assign \new_[51698]_  = \new_[51697]_  & \new_[51694]_ ;
  assign \new_[51699]_  = \new_[51698]_  & \new_[51691]_ ;
  assign \new_[51702]_  = A265 & ~A235;
  assign \new_[51705]_  = ~A267 & A266;
  assign \new_[51706]_  = \new_[51705]_  & \new_[51702]_ ;
  assign \new_[51709]_  = ~A298 & ~A268;
  assign \new_[51712]_  = ~A301 & ~A299;
  assign \new_[51713]_  = \new_[51712]_  & \new_[51709]_ ;
  assign \new_[51714]_  = \new_[51713]_  & \new_[51706]_ ;
  assign \new_[51717]_  = ~A169 & ~A170;
  assign \new_[51720]_  = A199 & ~A168;
  assign \new_[51721]_  = \new_[51720]_  & \new_[51717]_ ;
  assign \new_[51724]_  = A203 & ~A200;
  assign \new_[51727]_  = ~A233 & ~A232;
  assign \new_[51728]_  = \new_[51727]_  & \new_[51724]_ ;
  assign \new_[51729]_  = \new_[51728]_  & \new_[51721]_ ;
  assign \new_[51732]_  = ~A265 & ~A235;
  assign \new_[51735]_  = ~A268 & ~A266;
  assign \new_[51736]_  = \new_[51735]_  & \new_[51732]_ ;
  assign \new_[51739]_  = A299 & A298;
  assign \new_[51742]_  = ~A301 & ~A300;
  assign \new_[51743]_  = \new_[51742]_  & \new_[51739]_ ;
  assign \new_[51744]_  = \new_[51743]_  & \new_[51736]_ ;
  assign \new_[51747]_  = A166 & A168;
  assign \new_[51750]_  = ~A202 & ~A201;
  assign \new_[51751]_  = \new_[51750]_  & \new_[51747]_ ;
  assign \new_[51754]_  = A232 & ~A203;
  assign \new_[51757]_  = ~A234 & A233;
  assign \new_[51758]_  = \new_[51757]_  & \new_[51754]_ ;
  assign \new_[51759]_  = \new_[51758]_  & \new_[51751]_ ;
  assign \new_[51762]_  = A265 & ~A235;
  assign \new_[51765]_  = ~A267 & A266;
  assign \new_[51766]_  = \new_[51765]_  & \new_[51762]_ ;
  assign \new_[51769]_  = A298 & ~A268;
  assign \new_[51773]_  = ~A301 & ~A300;
  assign \new_[51774]_  = A299 & \new_[51773]_ ;
  assign \new_[51775]_  = \new_[51774]_  & \new_[51769]_ ;
  assign \new_[51776]_  = \new_[51775]_  & \new_[51766]_ ;
  assign \new_[51779]_  = A166 & A168;
  assign \new_[51782]_  = A200 & A199;
  assign \new_[51783]_  = \new_[51782]_  & \new_[51779]_ ;
  assign \new_[51786]_  = ~A202 & ~A201;
  assign \new_[51789]_  = ~A235 & ~A234;
  assign \new_[51790]_  = \new_[51789]_  & \new_[51786]_ ;
  assign \new_[51791]_  = \new_[51790]_  & \new_[51783]_ ;
  assign \new_[51794]_  = A265 & ~A236;
  assign \new_[51797]_  = ~A267 & A266;
  assign \new_[51798]_  = \new_[51797]_  & \new_[51794]_ ;
  assign \new_[51801]_  = A298 & ~A268;
  assign \new_[51805]_  = ~A301 & ~A300;
  assign \new_[51806]_  = A299 & \new_[51805]_ ;
  assign \new_[51807]_  = \new_[51806]_  & \new_[51801]_ ;
  assign \new_[51808]_  = \new_[51807]_  & \new_[51798]_ ;
  assign \new_[51811]_  = A166 & A168;
  assign \new_[51814]_  = A200 & A199;
  assign \new_[51815]_  = \new_[51814]_  & \new_[51811]_ ;
  assign \new_[51818]_  = ~A202 & ~A201;
  assign \new_[51821]_  = A233 & A232;
  assign \new_[51822]_  = \new_[51821]_  & \new_[51818]_ ;
  assign \new_[51823]_  = \new_[51822]_  & \new_[51815]_ ;
  assign \new_[51826]_  = ~A235 & ~A234;
  assign \new_[51829]_  = ~A268 & ~A267;
  assign \new_[51830]_  = \new_[51829]_  & \new_[51826]_ ;
  assign \new_[51833]_  = A298 & ~A269;
  assign \new_[51837]_  = ~A301 & ~A300;
  assign \new_[51838]_  = A299 & \new_[51837]_ ;
  assign \new_[51839]_  = \new_[51838]_  & \new_[51833]_ ;
  assign \new_[51840]_  = \new_[51839]_  & \new_[51830]_ ;
  assign \new_[51843]_  = A166 & A168;
  assign \new_[51846]_  = A200 & A199;
  assign \new_[51847]_  = \new_[51846]_  & \new_[51843]_ ;
  assign \new_[51850]_  = ~A202 & ~A201;
  assign \new_[51853]_  = A233 & A232;
  assign \new_[51854]_  = \new_[51853]_  & \new_[51850]_ ;
  assign \new_[51855]_  = \new_[51854]_  & \new_[51847]_ ;
  assign \new_[51858]_  = ~A235 & ~A234;
  assign \new_[51861]_  = A266 & A265;
  assign \new_[51862]_  = \new_[51861]_  & \new_[51858]_ ;
  assign \new_[51865]_  = ~A268 & ~A267;
  assign \new_[51869]_  = ~A302 & ~A301;
  assign \new_[51870]_  = ~A300 & \new_[51869]_ ;
  assign \new_[51871]_  = \new_[51870]_  & \new_[51865]_ ;
  assign \new_[51872]_  = \new_[51871]_  & \new_[51862]_ ;
  assign \new_[51875]_  = A166 & A168;
  assign \new_[51878]_  = A200 & A199;
  assign \new_[51879]_  = \new_[51878]_  & \new_[51875]_ ;
  assign \new_[51882]_  = ~A202 & ~A201;
  assign \new_[51885]_  = A233 & A232;
  assign \new_[51886]_  = \new_[51885]_  & \new_[51882]_ ;
  assign \new_[51887]_  = \new_[51886]_  & \new_[51879]_ ;
  assign \new_[51890]_  = ~A235 & ~A234;
  assign \new_[51893]_  = A266 & A265;
  assign \new_[51894]_  = \new_[51893]_  & \new_[51890]_ ;
  assign \new_[51897]_  = ~A268 & ~A267;
  assign \new_[51901]_  = ~A301 & ~A299;
  assign \new_[51902]_  = ~A298 & \new_[51901]_ ;
  assign \new_[51903]_  = \new_[51902]_  & \new_[51897]_ ;
  assign \new_[51904]_  = \new_[51903]_  & \new_[51894]_ ;
  assign \new_[51907]_  = A166 & A168;
  assign \new_[51910]_  = A200 & A199;
  assign \new_[51911]_  = \new_[51910]_  & \new_[51907]_ ;
  assign \new_[51914]_  = ~A202 & ~A201;
  assign \new_[51917]_  = A233 & A232;
  assign \new_[51918]_  = \new_[51917]_  & \new_[51914]_ ;
  assign \new_[51919]_  = \new_[51918]_  & \new_[51911]_ ;
  assign \new_[51922]_  = ~A235 & ~A234;
  assign \new_[51925]_  = ~A266 & ~A265;
  assign \new_[51926]_  = \new_[51925]_  & \new_[51922]_ ;
  assign \new_[51929]_  = A298 & ~A268;
  assign \new_[51933]_  = ~A301 & ~A300;
  assign \new_[51934]_  = A299 & \new_[51933]_ ;
  assign \new_[51935]_  = \new_[51934]_  & \new_[51929]_ ;
  assign \new_[51936]_  = \new_[51935]_  & \new_[51926]_ ;
  assign \new_[51939]_  = A166 & A168;
  assign \new_[51942]_  = A200 & A199;
  assign \new_[51943]_  = \new_[51942]_  & \new_[51939]_ ;
  assign \new_[51946]_  = ~A202 & ~A201;
  assign \new_[51949]_  = ~A233 & ~A232;
  assign \new_[51950]_  = \new_[51949]_  & \new_[51946]_ ;
  assign \new_[51951]_  = \new_[51950]_  & \new_[51943]_ ;
  assign \new_[51954]_  = A265 & ~A235;
  assign \new_[51957]_  = ~A267 & A266;
  assign \new_[51958]_  = \new_[51957]_  & \new_[51954]_ ;
  assign \new_[51961]_  = A298 & ~A268;
  assign \new_[51965]_  = ~A301 & ~A300;
  assign \new_[51966]_  = A299 & \new_[51965]_ ;
  assign \new_[51967]_  = \new_[51966]_  & \new_[51961]_ ;
  assign \new_[51968]_  = \new_[51967]_  & \new_[51958]_ ;
  assign \new_[51971]_  = A166 & A168;
  assign \new_[51974]_  = ~A200 & ~A199;
  assign \new_[51975]_  = \new_[51974]_  & \new_[51971]_ ;
  assign \new_[51978]_  = A232 & ~A202;
  assign \new_[51981]_  = ~A234 & A233;
  assign \new_[51982]_  = \new_[51981]_  & \new_[51978]_ ;
  assign \new_[51983]_  = \new_[51982]_  & \new_[51975]_ ;
  assign \new_[51986]_  = A265 & ~A235;
  assign \new_[51989]_  = ~A267 & A266;
  assign \new_[51990]_  = \new_[51989]_  & \new_[51986]_ ;
  assign \new_[51993]_  = A298 & ~A268;
  assign \new_[51997]_  = ~A301 & ~A300;
  assign \new_[51998]_  = A299 & \new_[51997]_ ;
  assign \new_[51999]_  = \new_[51998]_  & \new_[51993]_ ;
  assign \new_[52000]_  = \new_[51999]_  & \new_[51990]_ ;
  assign \new_[52003]_  = A167 & A168;
  assign \new_[52006]_  = ~A202 & ~A201;
  assign \new_[52007]_  = \new_[52006]_  & \new_[52003]_ ;
  assign \new_[52010]_  = A232 & ~A203;
  assign \new_[52013]_  = ~A234 & A233;
  assign \new_[52014]_  = \new_[52013]_  & \new_[52010]_ ;
  assign \new_[52015]_  = \new_[52014]_  & \new_[52007]_ ;
  assign \new_[52018]_  = A265 & ~A235;
  assign \new_[52021]_  = ~A267 & A266;
  assign \new_[52022]_  = \new_[52021]_  & \new_[52018]_ ;
  assign \new_[52025]_  = A298 & ~A268;
  assign \new_[52029]_  = ~A301 & ~A300;
  assign \new_[52030]_  = A299 & \new_[52029]_ ;
  assign \new_[52031]_  = \new_[52030]_  & \new_[52025]_ ;
  assign \new_[52032]_  = \new_[52031]_  & \new_[52022]_ ;
  assign \new_[52035]_  = A167 & A168;
  assign \new_[52038]_  = A200 & A199;
  assign \new_[52039]_  = \new_[52038]_  & \new_[52035]_ ;
  assign \new_[52042]_  = ~A202 & ~A201;
  assign \new_[52045]_  = ~A235 & ~A234;
  assign \new_[52046]_  = \new_[52045]_  & \new_[52042]_ ;
  assign \new_[52047]_  = \new_[52046]_  & \new_[52039]_ ;
  assign \new_[52050]_  = A265 & ~A236;
  assign \new_[52053]_  = ~A267 & A266;
  assign \new_[52054]_  = \new_[52053]_  & \new_[52050]_ ;
  assign \new_[52057]_  = A298 & ~A268;
  assign \new_[52061]_  = ~A301 & ~A300;
  assign \new_[52062]_  = A299 & \new_[52061]_ ;
  assign \new_[52063]_  = \new_[52062]_  & \new_[52057]_ ;
  assign \new_[52064]_  = \new_[52063]_  & \new_[52054]_ ;
  assign \new_[52067]_  = A167 & A168;
  assign \new_[52070]_  = A200 & A199;
  assign \new_[52071]_  = \new_[52070]_  & \new_[52067]_ ;
  assign \new_[52074]_  = ~A202 & ~A201;
  assign \new_[52077]_  = A233 & A232;
  assign \new_[52078]_  = \new_[52077]_  & \new_[52074]_ ;
  assign \new_[52079]_  = \new_[52078]_  & \new_[52071]_ ;
  assign \new_[52082]_  = ~A235 & ~A234;
  assign \new_[52085]_  = ~A268 & ~A267;
  assign \new_[52086]_  = \new_[52085]_  & \new_[52082]_ ;
  assign \new_[52089]_  = A298 & ~A269;
  assign \new_[52093]_  = ~A301 & ~A300;
  assign \new_[52094]_  = A299 & \new_[52093]_ ;
  assign \new_[52095]_  = \new_[52094]_  & \new_[52089]_ ;
  assign \new_[52096]_  = \new_[52095]_  & \new_[52086]_ ;
  assign \new_[52099]_  = A167 & A168;
  assign \new_[52102]_  = A200 & A199;
  assign \new_[52103]_  = \new_[52102]_  & \new_[52099]_ ;
  assign \new_[52106]_  = ~A202 & ~A201;
  assign \new_[52109]_  = A233 & A232;
  assign \new_[52110]_  = \new_[52109]_  & \new_[52106]_ ;
  assign \new_[52111]_  = \new_[52110]_  & \new_[52103]_ ;
  assign \new_[52114]_  = ~A235 & ~A234;
  assign \new_[52117]_  = A266 & A265;
  assign \new_[52118]_  = \new_[52117]_  & \new_[52114]_ ;
  assign \new_[52121]_  = ~A268 & ~A267;
  assign \new_[52125]_  = ~A302 & ~A301;
  assign \new_[52126]_  = ~A300 & \new_[52125]_ ;
  assign \new_[52127]_  = \new_[52126]_  & \new_[52121]_ ;
  assign \new_[52128]_  = \new_[52127]_  & \new_[52118]_ ;
  assign \new_[52131]_  = A167 & A168;
  assign \new_[52134]_  = A200 & A199;
  assign \new_[52135]_  = \new_[52134]_  & \new_[52131]_ ;
  assign \new_[52138]_  = ~A202 & ~A201;
  assign \new_[52141]_  = A233 & A232;
  assign \new_[52142]_  = \new_[52141]_  & \new_[52138]_ ;
  assign \new_[52143]_  = \new_[52142]_  & \new_[52135]_ ;
  assign \new_[52146]_  = ~A235 & ~A234;
  assign \new_[52149]_  = A266 & A265;
  assign \new_[52150]_  = \new_[52149]_  & \new_[52146]_ ;
  assign \new_[52153]_  = ~A268 & ~A267;
  assign \new_[52157]_  = ~A301 & ~A299;
  assign \new_[52158]_  = ~A298 & \new_[52157]_ ;
  assign \new_[52159]_  = \new_[52158]_  & \new_[52153]_ ;
  assign \new_[52160]_  = \new_[52159]_  & \new_[52150]_ ;
  assign \new_[52163]_  = A167 & A168;
  assign \new_[52166]_  = A200 & A199;
  assign \new_[52167]_  = \new_[52166]_  & \new_[52163]_ ;
  assign \new_[52170]_  = ~A202 & ~A201;
  assign \new_[52173]_  = A233 & A232;
  assign \new_[52174]_  = \new_[52173]_  & \new_[52170]_ ;
  assign \new_[52175]_  = \new_[52174]_  & \new_[52167]_ ;
  assign \new_[52178]_  = ~A235 & ~A234;
  assign \new_[52181]_  = ~A266 & ~A265;
  assign \new_[52182]_  = \new_[52181]_  & \new_[52178]_ ;
  assign \new_[52185]_  = A298 & ~A268;
  assign \new_[52189]_  = ~A301 & ~A300;
  assign \new_[52190]_  = A299 & \new_[52189]_ ;
  assign \new_[52191]_  = \new_[52190]_  & \new_[52185]_ ;
  assign \new_[52192]_  = \new_[52191]_  & \new_[52182]_ ;
  assign \new_[52195]_  = A167 & A168;
  assign \new_[52198]_  = A200 & A199;
  assign \new_[52199]_  = \new_[52198]_  & \new_[52195]_ ;
  assign \new_[52202]_  = ~A202 & ~A201;
  assign \new_[52205]_  = ~A233 & ~A232;
  assign \new_[52206]_  = \new_[52205]_  & \new_[52202]_ ;
  assign \new_[52207]_  = \new_[52206]_  & \new_[52199]_ ;
  assign \new_[52210]_  = A265 & ~A235;
  assign \new_[52213]_  = ~A267 & A266;
  assign \new_[52214]_  = \new_[52213]_  & \new_[52210]_ ;
  assign \new_[52217]_  = A298 & ~A268;
  assign \new_[52221]_  = ~A301 & ~A300;
  assign \new_[52222]_  = A299 & \new_[52221]_ ;
  assign \new_[52223]_  = \new_[52222]_  & \new_[52217]_ ;
  assign \new_[52224]_  = \new_[52223]_  & \new_[52214]_ ;
  assign \new_[52227]_  = A167 & A168;
  assign \new_[52230]_  = ~A200 & ~A199;
  assign \new_[52231]_  = \new_[52230]_  & \new_[52227]_ ;
  assign \new_[52234]_  = A232 & ~A202;
  assign \new_[52237]_  = ~A234 & A233;
  assign \new_[52238]_  = \new_[52237]_  & \new_[52234]_ ;
  assign \new_[52239]_  = \new_[52238]_  & \new_[52231]_ ;
  assign \new_[52242]_  = A265 & ~A235;
  assign \new_[52245]_  = ~A267 & A266;
  assign \new_[52246]_  = \new_[52245]_  & \new_[52242]_ ;
  assign \new_[52249]_  = A298 & ~A268;
  assign \new_[52253]_  = ~A301 & ~A300;
  assign \new_[52254]_  = A299 & \new_[52253]_ ;
  assign \new_[52255]_  = \new_[52254]_  & \new_[52249]_ ;
  assign \new_[52256]_  = \new_[52255]_  & \new_[52246]_ ;
  assign \new_[52259]_  = A167 & A170;
  assign \new_[52262]_  = ~A201 & ~A166;
  assign \new_[52263]_  = \new_[52262]_  & \new_[52259]_ ;
  assign \new_[52266]_  = ~A203 & ~A202;
  assign \new_[52269]_  = ~A235 & ~A234;
  assign \new_[52270]_  = \new_[52269]_  & \new_[52266]_ ;
  assign \new_[52271]_  = \new_[52270]_  & \new_[52263]_ ;
  assign \new_[52274]_  = A265 & ~A236;
  assign \new_[52277]_  = ~A267 & A266;
  assign \new_[52278]_  = \new_[52277]_  & \new_[52274]_ ;
  assign \new_[52281]_  = A298 & ~A268;
  assign \new_[52285]_  = ~A301 & ~A300;
  assign \new_[52286]_  = A299 & \new_[52285]_ ;
  assign \new_[52287]_  = \new_[52286]_  & \new_[52281]_ ;
  assign \new_[52288]_  = \new_[52287]_  & \new_[52278]_ ;
  assign \new_[52291]_  = A167 & A170;
  assign \new_[52294]_  = ~A201 & ~A166;
  assign \new_[52295]_  = \new_[52294]_  & \new_[52291]_ ;
  assign \new_[52298]_  = ~A203 & ~A202;
  assign \new_[52301]_  = A233 & A232;
  assign \new_[52302]_  = \new_[52301]_  & \new_[52298]_ ;
  assign \new_[52303]_  = \new_[52302]_  & \new_[52295]_ ;
  assign \new_[52306]_  = ~A235 & ~A234;
  assign \new_[52309]_  = ~A268 & ~A267;
  assign \new_[52310]_  = \new_[52309]_  & \new_[52306]_ ;
  assign \new_[52313]_  = A298 & ~A269;
  assign \new_[52317]_  = ~A301 & ~A300;
  assign \new_[52318]_  = A299 & \new_[52317]_ ;
  assign \new_[52319]_  = \new_[52318]_  & \new_[52313]_ ;
  assign \new_[52320]_  = \new_[52319]_  & \new_[52310]_ ;
  assign \new_[52323]_  = A167 & A170;
  assign \new_[52326]_  = ~A201 & ~A166;
  assign \new_[52327]_  = \new_[52326]_  & \new_[52323]_ ;
  assign \new_[52330]_  = ~A203 & ~A202;
  assign \new_[52333]_  = A233 & A232;
  assign \new_[52334]_  = \new_[52333]_  & \new_[52330]_ ;
  assign \new_[52335]_  = \new_[52334]_  & \new_[52327]_ ;
  assign \new_[52338]_  = ~A235 & ~A234;
  assign \new_[52341]_  = A266 & A265;
  assign \new_[52342]_  = \new_[52341]_  & \new_[52338]_ ;
  assign \new_[52345]_  = ~A268 & ~A267;
  assign \new_[52349]_  = ~A302 & ~A301;
  assign \new_[52350]_  = ~A300 & \new_[52349]_ ;
  assign \new_[52351]_  = \new_[52350]_  & \new_[52345]_ ;
  assign \new_[52352]_  = \new_[52351]_  & \new_[52342]_ ;
  assign \new_[52355]_  = A167 & A170;
  assign \new_[52358]_  = ~A201 & ~A166;
  assign \new_[52359]_  = \new_[52358]_  & \new_[52355]_ ;
  assign \new_[52362]_  = ~A203 & ~A202;
  assign \new_[52365]_  = A233 & A232;
  assign \new_[52366]_  = \new_[52365]_  & \new_[52362]_ ;
  assign \new_[52367]_  = \new_[52366]_  & \new_[52359]_ ;
  assign \new_[52370]_  = ~A235 & ~A234;
  assign \new_[52373]_  = A266 & A265;
  assign \new_[52374]_  = \new_[52373]_  & \new_[52370]_ ;
  assign \new_[52377]_  = ~A268 & ~A267;
  assign \new_[52381]_  = ~A301 & ~A299;
  assign \new_[52382]_  = ~A298 & \new_[52381]_ ;
  assign \new_[52383]_  = \new_[52382]_  & \new_[52377]_ ;
  assign \new_[52384]_  = \new_[52383]_  & \new_[52374]_ ;
  assign \new_[52387]_  = A167 & A170;
  assign \new_[52390]_  = ~A201 & ~A166;
  assign \new_[52391]_  = \new_[52390]_  & \new_[52387]_ ;
  assign \new_[52394]_  = ~A203 & ~A202;
  assign \new_[52397]_  = A233 & A232;
  assign \new_[52398]_  = \new_[52397]_  & \new_[52394]_ ;
  assign \new_[52399]_  = \new_[52398]_  & \new_[52391]_ ;
  assign \new_[52402]_  = ~A235 & ~A234;
  assign \new_[52405]_  = ~A266 & ~A265;
  assign \new_[52406]_  = \new_[52405]_  & \new_[52402]_ ;
  assign \new_[52409]_  = A298 & ~A268;
  assign \new_[52413]_  = ~A301 & ~A300;
  assign \new_[52414]_  = A299 & \new_[52413]_ ;
  assign \new_[52415]_  = \new_[52414]_  & \new_[52409]_ ;
  assign \new_[52416]_  = \new_[52415]_  & \new_[52406]_ ;
  assign \new_[52419]_  = A167 & A170;
  assign \new_[52422]_  = ~A201 & ~A166;
  assign \new_[52423]_  = \new_[52422]_  & \new_[52419]_ ;
  assign \new_[52426]_  = ~A203 & ~A202;
  assign \new_[52429]_  = ~A233 & ~A232;
  assign \new_[52430]_  = \new_[52429]_  & \new_[52426]_ ;
  assign \new_[52431]_  = \new_[52430]_  & \new_[52423]_ ;
  assign \new_[52434]_  = A265 & ~A235;
  assign \new_[52437]_  = ~A267 & A266;
  assign \new_[52438]_  = \new_[52437]_  & \new_[52434]_ ;
  assign \new_[52441]_  = A298 & ~A268;
  assign \new_[52445]_  = ~A301 & ~A300;
  assign \new_[52446]_  = A299 & \new_[52445]_ ;
  assign \new_[52447]_  = \new_[52446]_  & \new_[52441]_ ;
  assign \new_[52448]_  = \new_[52447]_  & \new_[52438]_ ;
  assign \new_[52451]_  = A167 & A170;
  assign \new_[52454]_  = A199 & ~A166;
  assign \new_[52455]_  = \new_[52454]_  & \new_[52451]_ ;
  assign \new_[52458]_  = ~A201 & A200;
  assign \new_[52461]_  = ~A234 & ~A202;
  assign \new_[52462]_  = \new_[52461]_  & \new_[52458]_ ;
  assign \new_[52463]_  = \new_[52462]_  & \new_[52455]_ ;
  assign \new_[52466]_  = ~A236 & ~A235;
  assign \new_[52469]_  = ~A268 & ~A267;
  assign \new_[52470]_  = \new_[52469]_  & \new_[52466]_ ;
  assign \new_[52473]_  = A298 & ~A269;
  assign \new_[52477]_  = ~A301 & ~A300;
  assign \new_[52478]_  = A299 & \new_[52477]_ ;
  assign \new_[52479]_  = \new_[52478]_  & \new_[52473]_ ;
  assign \new_[52480]_  = \new_[52479]_  & \new_[52470]_ ;
  assign \new_[52483]_  = A167 & A170;
  assign \new_[52486]_  = A199 & ~A166;
  assign \new_[52487]_  = \new_[52486]_  & \new_[52483]_ ;
  assign \new_[52490]_  = ~A201 & A200;
  assign \new_[52493]_  = ~A234 & ~A202;
  assign \new_[52494]_  = \new_[52493]_  & \new_[52490]_ ;
  assign \new_[52495]_  = \new_[52494]_  & \new_[52487]_ ;
  assign \new_[52498]_  = ~A236 & ~A235;
  assign \new_[52501]_  = A266 & A265;
  assign \new_[52502]_  = \new_[52501]_  & \new_[52498]_ ;
  assign \new_[52505]_  = ~A268 & ~A267;
  assign \new_[52509]_  = ~A302 & ~A301;
  assign \new_[52510]_  = ~A300 & \new_[52509]_ ;
  assign \new_[52511]_  = \new_[52510]_  & \new_[52505]_ ;
  assign \new_[52512]_  = \new_[52511]_  & \new_[52502]_ ;
  assign \new_[52515]_  = A167 & A170;
  assign \new_[52518]_  = A199 & ~A166;
  assign \new_[52519]_  = \new_[52518]_  & \new_[52515]_ ;
  assign \new_[52522]_  = ~A201 & A200;
  assign \new_[52525]_  = ~A234 & ~A202;
  assign \new_[52526]_  = \new_[52525]_  & \new_[52522]_ ;
  assign \new_[52527]_  = \new_[52526]_  & \new_[52519]_ ;
  assign \new_[52530]_  = ~A236 & ~A235;
  assign \new_[52533]_  = A266 & A265;
  assign \new_[52534]_  = \new_[52533]_  & \new_[52530]_ ;
  assign \new_[52537]_  = ~A268 & ~A267;
  assign \new_[52541]_  = ~A301 & ~A299;
  assign \new_[52542]_  = ~A298 & \new_[52541]_ ;
  assign \new_[52543]_  = \new_[52542]_  & \new_[52537]_ ;
  assign \new_[52544]_  = \new_[52543]_  & \new_[52534]_ ;
  assign \new_[52547]_  = A167 & A170;
  assign \new_[52550]_  = A199 & ~A166;
  assign \new_[52551]_  = \new_[52550]_  & \new_[52547]_ ;
  assign \new_[52554]_  = ~A201 & A200;
  assign \new_[52557]_  = ~A234 & ~A202;
  assign \new_[52558]_  = \new_[52557]_  & \new_[52554]_ ;
  assign \new_[52559]_  = \new_[52558]_  & \new_[52551]_ ;
  assign \new_[52562]_  = ~A236 & ~A235;
  assign \new_[52565]_  = ~A266 & ~A265;
  assign \new_[52566]_  = \new_[52565]_  & \new_[52562]_ ;
  assign \new_[52569]_  = A298 & ~A268;
  assign \new_[52573]_  = ~A301 & ~A300;
  assign \new_[52574]_  = A299 & \new_[52573]_ ;
  assign \new_[52575]_  = \new_[52574]_  & \new_[52569]_ ;
  assign \new_[52576]_  = \new_[52575]_  & \new_[52566]_ ;
  assign \new_[52579]_  = A167 & A170;
  assign \new_[52582]_  = A199 & ~A166;
  assign \new_[52583]_  = \new_[52582]_  & \new_[52579]_ ;
  assign \new_[52586]_  = ~A201 & A200;
  assign \new_[52589]_  = A232 & ~A202;
  assign \new_[52590]_  = \new_[52589]_  & \new_[52586]_ ;
  assign \new_[52591]_  = \new_[52590]_  & \new_[52583]_ ;
  assign \new_[52594]_  = ~A234 & A233;
  assign \new_[52597]_  = ~A267 & ~A235;
  assign \new_[52598]_  = \new_[52597]_  & \new_[52594]_ ;
  assign \new_[52601]_  = ~A269 & ~A268;
  assign \new_[52605]_  = ~A302 & ~A301;
  assign \new_[52606]_  = ~A300 & \new_[52605]_ ;
  assign \new_[52607]_  = \new_[52606]_  & \new_[52601]_ ;
  assign \new_[52608]_  = \new_[52607]_  & \new_[52598]_ ;
  assign \new_[52611]_  = A167 & A170;
  assign \new_[52614]_  = A199 & ~A166;
  assign \new_[52615]_  = \new_[52614]_  & \new_[52611]_ ;
  assign \new_[52618]_  = ~A201 & A200;
  assign \new_[52621]_  = A232 & ~A202;
  assign \new_[52622]_  = \new_[52621]_  & \new_[52618]_ ;
  assign \new_[52623]_  = \new_[52622]_  & \new_[52615]_ ;
  assign \new_[52626]_  = ~A234 & A233;
  assign \new_[52629]_  = ~A267 & ~A235;
  assign \new_[52630]_  = \new_[52629]_  & \new_[52626]_ ;
  assign \new_[52633]_  = ~A269 & ~A268;
  assign \new_[52637]_  = ~A301 & ~A299;
  assign \new_[52638]_  = ~A298 & \new_[52637]_ ;
  assign \new_[52639]_  = \new_[52638]_  & \new_[52633]_ ;
  assign \new_[52640]_  = \new_[52639]_  & \new_[52630]_ ;
  assign \new_[52643]_  = A167 & A170;
  assign \new_[52646]_  = A199 & ~A166;
  assign \new_[52647]_  = \new_[52646]_  & \new_[52643]_ ;
  assign \new_[52650]_  = ~A201 & A200;
  assign \new_[52653]_  = A232 & ~A202;
  assign \new_[52654]_  = \new_[52653]_  & \new_[52650]_ ;
  assign \new_[52655]_  = \new_[52654]_  & \new_[52647]_ ;
  assign \new_[52658]_  = ~A234 & A233;
  assign \new_[52661]_  = ~A265 & ~A235;
  assign \new_[52662]_  = \new_[52661]_  & \new_[52658]_ ;
  assign \new_[52665]_  = ~A268 & ~A266;
  assign \new_[52669]_  = ~A302 & ~A301;
  assign \new_[52670]_  = ~A300 & \new_[52669]_ ;
  assign \new_[52671]_  = \new_[52670]_  & \new_[52665]_ ;
  assign \new_[52672]_  = \new_[52671]_  & \new_[52662]_ ;
  assign \new_[52675]_  = A167 & A170;
  assign \new_[52678]_  = A199 & ~A166;
  assign \new_[52679]_  = \new_[52678]_  & \new_[52675]_ ;
  assign \new_[52682]_  = ~A201 & A200;
  assign \new_[52685]_  = A232 & ~A202;
  assign \new_[52686]_  = \new_[52685]_  & \new_[52682]_ ;
  assign \new_[52687]_  = \new_[52686]_  & \new_[52679]_ ;
  assign \new_[52690]_  = ~A234 & A233;
  assign \new_[52693]_  = ~A265 & ~A235;
  assign \new_[52694]_  = \new_[52693]_  & \new_[52690]_ ;
  assign \new_[52697]_  = ~A268 & ~A266;
  assign \new_[52701]_  = ~A301 & ~A299;
  assign \new_[52702]_  = ~A298 & \new_[52701]_ ;
  assign \new_[52703]_  = \new_[52702]_  & \new_[52697]_ ;
  assign \new_[52704]_  = \new_[52703]_  & \new_[52694]_ ;
  assign \new_[52707]_  = A167 & A170;
  assign \new_[52710]_  = A199 & ~A166;
  assign \new_[52711]_  = \new_[52710]_  & \new_[52707]_ ;
  assign \new_[52714]_  = ~A201 & A200;
  assign \new_[52717]_  = ~A232 & ~A202;
  assign \new_[52718]_  = \new_[52717]_  & \new_[52714]_ ;
  assign \new_[52719]_  = \new_[52718]_  & \new_[52711]_ ;
  assign \new_[52722]_  = ~A235 & ~A233;
  assign \new_[52725]_  = ~A268 & ~A267;
  assign \new_[52726]_  = \new_[52725]_  & \new_[52722]_ ;
  assign \new_[52729]_  = A298 & ~A269;
  assign \new_[52733]_  = ~A301 & ~A300;
  assign \new_[52734]_  = A299 & \new_[52733]_ ;
  assign \new_[52735]_  = \new_[52734]_  & \new_[52729]_ ;
  assign \new_[52736]_  = \new_[52735]_  & \new_[52726]_ ;
  assign \new_[52739]_  = A167 & A170;
  assign \new_[52742]_  = A199 & ~A166;
  assign \new_[52743]_  = \new_[52742]_  & \new_[52739]_ ;
  assign \new_[52746]_  = ~A201 & A200;
  assign \new_[52749]_  = ~A232 & ~A202;
  assign \new_[52750]_  = \new_[52749]_  & \new_[52746]_ ;
  assign \new_[52751]_  = \new_[52750]_  & \new_[52743]_ ;
  assign \new_[52754]_  = ~A235 & ~A233;
  assign \new_[52757]_  = A266 & A265;
  assign \new_[52758]_  = \new_[52757]_  & \new_[52754]_ ;
  assign \new_[52761]_  = ~A268 & ~A267;
  assign \new_[52765]_  = ~A302 & ~A301;
  assign \new_[52766]_  = ~A300 & \new_[52765]_ ;
  assign \new_[52767]_  = \new_[52766]_  & \new_[52761]_ ;
  assign \new_[52768]_  = \new_[52767]_  & \new_[52758]_ ;
  assign \new_[52771]_  = A167 & A170;
  assign \new_[52774]_  = A199 & ~A166;
  assign \new_[52775]_  = \new_[52774]_  & \new_[52771]_ ;
  assign \new_[52778]_  = ~A201 & A200;
  assign \new_[52781]_  = ~A232 & ~A202;
  assign \new_[52782]_  = \new_[52781]_  & \new_[52778]_ ;
  assign \new_[52783]_  = \new_[52782]_  & \new_[52775]_ ;
  assign \new_[52786]_  = ~A235 & ~A233;
  assign \new_[52789]_  = A266 & A265;
  assign \new_[52790]_  = \new_[52789]_  & \new_[52786]_ ;
  assign \new_[52793]_  = ~A268 & ~A267;
  assign \new_[52797]_  = ~A301 & ~A299;
  assign \new_[52798]_  = ~A298 & \new_[52797]_ ;
  assign \new_[52799]_  = \new_[52798]_  & \new_[52793]_ ;
  assign \new_[52800]_  = \new_[52799]_  & \new_[52790]_ ;
  assign \new_[52803]_  = A167 & A170;
  assign \new_[52806]_  = A199 & ~A166;
  assign \new_[52807]_  = \new_[52806]_  & \new_[52803]_ ;
  assign \new_[52810]_  = ~A201 & A200;
  assign \new_[52813]_  = ~A232 & ~A202;
  assign \new_[52814]_  = \new_[52813]_  & \new_[52810]_ ;
  assign \new_[52815]_  = \new_[52814]_  & \new_[52807]_ ;
  assign \new_[52818]_  = ~A235 & ~A233;
  assign \new_[52821]_  = ~A266 & ~A265;
  assign \new_[52822]_  = \new_[52821]_  & \new_[52818]_ ;
  assign \new_[52825]_  = A298 & ~A268;
  assign \new_[52829]_  = ~A301 & ~A300;
  assign \new_[52830]_  = A299 & \new_[52829]_ ;
  assign \new_[52831]_  = \new_[52830]_  & \new_[52825]_ ;
  assign \new_[52832]_  = \new_[52831]_  & \new_[52822]_ ;
  assign \new_[52835]_  = A167 & A170;
  assign \new_[52838]_  = ~A199 & ~A166;
  assign \new_[52839]_  = \new_[52838]_  & \new_[52835]_ ;
  assign \new_[52842]_  = ~A202 & ~A200;
  assign \new_[52845]_  = ~A235 & ~A234;
  assign \new_[52846]_  = \new_[52845]_  & \new_[52842]_ ;
  assign \new_[52847]_  = \new_[52846]_  & \new_[52839]_ ;
  assign \new_[52850]_  = A265 & ~A236;
  assign \new_[52853]_  = ~A267 & A266;
  assign \new_[52854]_  = \new_[52853]_  & \new_[52850]_ ;
  assign \new_[52857]_  = A298 & ~A268;
  assign \new_[52861]_  = ~A301 & ~A300;
  assign \new_[52862]_  = A299 & \new_[52861]_ ;
  assign \new_[52863]_  = \new_[52862]_  & \new_[52857]_ ;
  assign \new_[52864]_  = \new_[52863]_  & \new_[52854]_ ;
  assign \new_[52867]_  = A167 & A170;
  assign \new_[52870]_  = ~A199 & ~A166;
  assign \new_[52871]_  = \new_[52870]_  & \new_[52867]_ ;
  assign \new_[52874]_  = ~A202 & ~A200;
  assign \new_[52877]_  = A233 & A232;
  assign \new_[52878]_  = \new_[52877]_  & \new_[52874]_ ;
  assign \new_[52879]_  = \new_[52878]_  & \new_[52871]_ ;
  assign \new_[52882]_  = ~A235 & ~A234;
  assign \new_[52885]_  = ~A268 & ~A267;
  assign \new_[52886]_  = \new_[52885]_  & \new_[52882]_ ;
  assign \new_[52889]_  = A298 & ~A269;
  assign \new_[52893]_  = ~A301 & ~A300;
  assign \new_[52894]_  = A299 & \new_[52893]_ ;
  assign \new_[52895]_  = \new_[52894]_  & \new_[52889]_ ;
  assign \new_[52896]_  = \new_[52895]_  & \new_[52886]_ ;
  assign \new_[52899]_  = A167 & A170;
  assign \new_[52902]_  = ~A199 & ~A166;
  assign \new_[52903]_  = \new_[52902]_  & \new_[52899]_ ;
  assign \new_[52906]_  = ~A202 & ~A200;
  assign \new_[52909]_  = A233 & A232;
  assign \new_[52910]_  = \new_[52909]_  & \new_[52906]_ ;
  assign \new_[52911]_  = \new_[52910]_  & \new_[52903]_ ;
  assign \new_[52914]_  = ~A235 & ~A234;
  assign \new_[52917]_  = A266 & A265;
  assign \new_[52918]_  = \new_[52917]_  & \new_[52914]_ ;
  assign \new_[52921]_  = ~A268 & ~A267;
  assign \new_[52925]_  = ~A302 & ~A301;
  assign \new_[52926]_  = ~A300 & \new_[52925]_ ;
  assign \new_[52927]_  = \new_[52926]_  & \new_[52921]_ ;
  assign \new_[52928]_  = \new_[52927]_  & \new_[52918]_ ;
  assign \new_[52931]_  = A167 & A170;
  assign \new_[52934]_  = ~A199 & ~A166;
  assign \new_[52935]_  = \new_[52934]_  & \new_[52931]_ ;
  assign \new_[52938]_  = ~A202 & ~A200;
  assign \new_[52941]_  = A233 & A232;
  assign \new_[52942]_  = \new_[52941]_  & \new_[52938]_ ;
  assign \new_[52943]_  = \new_[52942]_  & \new_[52935]_ ;
  assign \new_[52946]_  = ~A235 & ~A234;
  assign \new_[52949]_  = A266 & A265;
  assign \new_[52950]_  = \new_[52949]_  & \new_[52946]_ ;
  assign \new_[52953]_  = ~A268 & ~A267;
  assign \new_[52957]_  = ~A301 & ~A299;
  assign \new_[52958]_  = ~A298 & \new_[52957]_ ;
  assign \new_[52959]_  = \new_[52958]_  & \new_[52953]_ ;
  assign \new_[52960]_  = \new_[52959]_  & \new_[52950]_ ;
  assign \new_[52963]_  = A167 & A170;
  assign \new_[52966]_  = ~A199 & ~A166;
  assign \new_[52967]_  = \new_[52966]_  & \new_[52963]_ ;
  assign \new_[52970]_  = ~A202 & ~A200;
  assign \new_[52973]_  = A233 & A232;
  assign \new_[52974]_  = \new_[52973]_  & \new_[52970]_ ;
  assign \new_[52975]_  = \new_[52974]_  & \new_[52967]_ ;
  assign \new_[52978]_  = ~A235 & ~A234;
  assign \new_[52981]_  = ~A266 & ~A265;
  assign \new_[52982]_  = \new_[52981]_  & \new_[52978]_ ;
  assign \new_[52985]_  = A298 & ~A268;
  assign \new_[52989]_  = ~A301 & ~A300;
  assign \new_[52990]_  = A299 & \new_[52989]_ ;
  assign \new_[52991]_  = \new_[52990]_  & \new_[52985]_ ;
  assign \new_[52992]_  = \new_[52991]_  & \new_[52982]_ ;
  assign \new_[52995]_  = A167 & A170;
  assign \new_[52998]_  = ~A199 & ~A166;
  assign \new_[52999]_  = \new_[52998]_  & \new_[52995]_ ;
  assign \new_[53002]_  = ~A202 & ~A200;
  assign \new_[53005]_  = ~A233 & ~A232;
  assign \new_[53006]_  = \new_[53005]_  & \new_[53002]_ ;
  assign \new_[53007]_  = \new_[53006]_  & \new_[52999]_ ;
  assign \new_[53010]_  = A265 & ~A235;
  assign \new_[53013]_  = ~A267 & A266;
  assign \new_[53014]_  = \new_[53013]_  & \new_[53010]_ ;
  assign \new_[53017]_  = A298 & ~A268;
  assign \new_[53021]_  = ~A301 & ~A300;
  assign \new_[53022]_  = A299 & \new_[53021]_ ;
  assign \new_[53023]_  = \new_[53022]_  & \new_[53017]_ ;
  assign \new_[53024]_  = \new_[53023]_  & \new_[53014]_ ;
  assign \new_[53027]_  = ~A167 & A170;
  assign \new_[53030]_  = ~A201 & A166;
  assign \new_[53031]_  = \new_[53030]_  & \new_[53027]_ ;
  assign \new_[53034]_  = ~A203 & ~A202;
  assign \new_[53037]_  = ~A235 & ~A234;
  assign \new_[53038]_  = \new_[53037]_  & \new_[53034]_ ;
  assign \new_[53039]_  = \new_[53038]_  & \new_[53031]_ ;
  assign \new_[53042]_  = A265 & ~A236;
  assign \new_[53045]_  = ~A267 & A266;
  assign \new_[53046]_  = \new_[53045]_  & \new_[53042]_ ;
  assign \new_[53049]_  = A298 & ~A268;
  assign \new_[53053]_  = ~A301 & ~A300;
  assign \new_[53054]_  = A299 & \new_[53053]_ ;
  assign \new_[53055]_  = \new_[53054]_  & \new_[53049]_ ;
  assign \new_[53056]_  = \new_[53055]_  & \new_[53046]_ ;
  assign \new_[53059]_  = ~A167 & A170;
  assign \new_[53062]_  = ~A201 & A166;
  assign \new_[53063]_  = \new_[53062]_  & \new_[53059]_ ;
  assign \new_[53066]_  = ~A203 & ~A202;
  assign \new_[53069]_  = A233 & A232;
  assign \new_[53070]_  = \new_[53069]_  & \new_[53066]_ ;
  assign \new_[53071]_  = \new_[53070]_  & \new_[53063]_ ;
  assign \new_[53074]_  = ~A235 & ~A234;
  assign \new_[53077]_  = ~A268 & ~A267;
  assign \new_[53078]_  = \new_[53077]_  & \new_[53074]_ ;
  assign \new_[53081]_  = A298 & ~A269;
  assign \new_[53085]_  = ~A301 & ~A300;
  assign \new_[53086]_  = A299 & \new_[53085]_ ;
  assign \new_[53087]_  = \new_[53086]_  & \new_[53081]_ ;
  assign \new_[53088]_  = \new_[53087]_  & \new_[53078]_ ;
  assign \new_[53091]_  = ~A167 & A170;
  assign \new_[53094]_  = ~A201 & A166;
  assign \new_[53095]_  = \new_[53094]_  & \new_[53091]_ ;
  assign \new_[53098]_  = ~A203 & ~A202;
  assign \new_[53101]_  = A233 & A232;
  assign \new_[53102]_  = \new_[53101]_  & \new_[53098]_ ;
  assign \new_[53103]_  = \new_[53102]_  & \new_[53095]_ ;
  assign \new_[53106]_  = ~A235 & ~A234;
  assign \new_[53109]_  = A266 & A265;
  assign \new_[53110]_  = \new_[53109]_  & \new_[53106]_ ;
  assign \new_[53113]_  = ~A268 & ~A267;
  assign \new_[53117]_  = ~A302 & ~A301;
  assign \new_[53118]_  = ~A300 & \new_[53117]_ ;
  assign \new_[53119]_  = \new_[53118]_  & \new_[53113]_ ;
  assign \new_[53120]_  = \new_[53119]_  & \new_[53110]_ ;
  assign \new_[53123]_  = ~A167 & A170;
  assign \new_[53126]_  = ~A201 & A166;
  assign \new_[53127]_  = \new_[53126]_  & \new_[53123]_ ;
  assign \new_[53130]_  = ~A203 & ~A202;
  assign \new_[53133]_  = A233 & A232;
  assign \new_[53134]_  = \new_[53133]_  & \new_[53130]_ ;
  assign \new_[53135]_  = \new_[53134]_  & \new_[53127]_ ;
  assign \new_[53138]_  = ~A235 & ~A234;
  assign \new_[53141]_  = A266 & A265;
  assign \new_[53142]_  = \new_[53141]_  & \new_[53138]_ ;
  assign \new_[53145]_  = ~A268 & ~A267;
  assign \new_[53149]_  = ~A301 & ~A299;
  assign \new_[53150]_  = ~A298 & \new_[53149]_ ;
  assign \new_[53151]_  = \new_[53150]_  & \new_[53145]_ ;
  assign \new_[53152]_  = \new_[53151]_  & \new_[53142]_ ;
  assign \new_[53155]_  = ~A167 & A170;
  assign \new_[53158]_  = ~A201 & A166;
  assign \new_[53159]_  = \new_[53158]_  & \new_[53155]_ ;
  assign \new_[53162]_  = ~A203 & ~A202;
  assign \new_[53165]_  = A233 & A232;
  assign \new_[53166]_  = \new_[53165]_  & \new_[53162]_ ;
  assign \new_[53167]_  = \new_[53166]_  & \new_[53159]_ ;
  assign \new_[53170]_  = ~A235 & ~A234;
  assign \new_[53173]_  = ~A266 & ~A265;
  assign \new_[53174]_  = \new_[53173]_  & \new_[53170]_ ;
  assign \new_[53177]_  = A298 & ~A268;
  assign \new_[53181]_  = ~A301 & ~A300;
  assign \new_[53182]_  = A299 & \new_[53181]_ ;
  assign \new_[53183]_  = \new_[53182]_  & \new_[53177]_ ;
  assign \new_[53184]_  = \new_[53183]_  & \new_[53174]_ ;
  assign \new_[53187]_  = ~A167 & A170;
  assign \new_[53190]_  = ~A201 & A166;
  assign \new_[53191]_  = \new_[53190]_  & \new_[53187]_ ;
  assign \new_[53194]_  = ~A203 & ~A202;
  assign \new_[53197]_  = ~A233 & ~A232;
  assign \new_[53198]_  = \new_[53197]_  & \new_[53194]_ ;
  assign \new_[53199]_  = \new_[53198]_  & \new_[53191]_ ;
  assign \new_[53202]_  = A265 & ~A235;
  assign \new_[53205]_  = ~A267 & A266;
  assign \new_[53206]_  = \new_[53205]_  & \new_[53202]_ ;
  assign \new_[53209]_  = A298 & ~A268;
  assign \new_[53213]_  = ~A301 & ~A300;
  assign \new_[53214]_  = A299 & \new_[53213]_ ;
  assign \new_[53215]_  = \new_[53214]_  & \new_[53209]_ ;
  assign \new_[53216]_  = \new_[53215]_  & \new_[53206]_ ;
  assign \new_[53219]_  = ~A167 & A170;
  assign \new_[53222]_  = A199 & A166;
  assign \new_[53223]_  = \new_[53222]_  & \new_[53219]_ ;
  assign \new_[53226]_  = ~A201 & A200;
  assign \new_[53229]_  = ~A234 & ~A202;
  assign \new_[53230]_  = \new_[53229]_  & \new_[53226]_ ;
  assign \new_[53231]_  = \new_[53230]_  & \new_[53223]_ ;
  assign \new_[53234]_  = ~A236 & ~A235;
  assign \new_[53237]_  = ~A268 & ~A267;
  assign \new_[53238]_  = \new_[53237]_  & \new_[53234]_ ;
  assign \new_[53241]_  = A298 & ~A269;
  assign \new_[53245]_  = ~A301 & ~A300;
  assign \new_[53246]_  = A299 & \new_[53245]_ ;
  assign \new_[53247]_  = \new_[53246]_  & \new_[53241]_ ;
  assign \new_[53248]_  = \new_[53247]_  & \new_[53238]_ ;
  assign \new_[53251]_  = ~A167 & A170;
  assign \new_[53254]_  = A199 & A166;
  assign \new_[53255]_  = \new_[53254]_  & \new_[53251]_ ;
  assign \new_[53258]_  = ~A201 & A200;
  assign \new_[53261]_  = ~A234 & ~A202;
  assign \new_[53262]_  = \new_[53261]_  & \new_[53258]_ ;
  assign \new_[53263]_  = \new_[53262]_  & \new_[53255]_ ;
  assign \new_[53266]_  = ~A236 & ~A235;
  assign \new_[53269]_  = A266 & A265;
  assign \new_[53270]_  = \new_[53269]_  & \new_[53266]_ ;
  assign \new_[53273]_  = ~A268 & ~A267;
  assign \new_[53277]_  = ~A302 & ~A301;
  assign \new_[53278]_  = ~A300 & \new_[53277]_ ;
  assign \new_[53279]_  = \new_[53278]_  & \new_[53273]_ ;
  assign \new_[53280]_  = \new_[53279]_  & \new_[53270]_ ;
  assign \new_[53283]_  = ~A167 & A170;
  assign \new_[53286]_  = A199 & A166;
  assign \new_[53287]_  = \new_[53286]_  & \new_[53283]_ ;
  assign \new_[53290]_  = ~A201 & A200;
  assign \new_[53293]_  = ~A234 & ~A202;
  assign \new_[53294]_  = \new_[53293]_  & \new_[53290]_ ;
  assign \new_[53295]_  = \new_[53294]_  & \new_[53287]_ ;
  assign \new_[53298]_  = ~A236 & ~A235;
  assign \new_[53301]_  = A266 & A265;
  assign \new_[53302]_  = \new_[53301]_  & \new_[53298]_ ;
  assign \new_[53305]_  = ~A268 & ~A267;
  assign \new_[53309]_  = ~A301 & ~A299;
  assign \new_[53310]_  = ~A298 & \new_[53309]_ ;
  assign \new_[53311]_  = \new_[53310]_  & \new_[53305]_ ;
  assign \new_[53312]_  = \new_[53311]_  & \new_[53302]_ ;
  assign \new_[53315]_  = ~A167 & A170;
  assign \new_[53318]_  = A199 & A166;
  assign \new_[53319]_  = \new_[53318]_  & \new_[53315]_ ;
  assign \new_[53322]_  = ~A201 & A200;
  assign \new_[53325]_  = ~A234 & ~A202;
  assign \new_[53326]_  = \new_[53325]_  & \new_[53322]_ ;
  assign \new_[53327]_  = \new_[53326]_  & \new_[53319]_ ;
  assign \new_[53330]_  = ~A236 & ~A235;
  assign \new_[53333]_  = ~A266 & ~A265;
  assign \new_[53334]_  = \new_[53333]_  & \new_[53330]_ ;
  assign \new_[53337]_  = A298 & ~A268;
  assign \new_[53341]_  = ~A301 & ~A300;
  assign \new_[53342]_  = A299 & \new_[53341]_ ;
  assign \new_[53343]_  = \new_[53342]_  & \new_[53337]_ ;
  assign \new_[53344]_  = \new_[53343]_  & \new_[53334]_ ;
  assign \new_[53347]_  = ~A167 & A170;
  assign \new_[53350]_  = A199 & A166;
  assign \new_[53351]_  = \new_[53350]_  & \new_[53347]_ ;
  assign \new_[53354]_  = ~A201 & A200;
  assign \new_[53357]_  = A232 & ~A202;
  assign \new_[53358]_  = \new_[53357]_  & \new_[53354]_ ;
  assign \new_[53359]_  = \new_[53358]_  & \new_[53351]_ ;
  assign \new_[53362]_  = ~A234 & A233;
  assign \new_[53365]_  = ~A267 & ~A235;
  assign \new_[53366]_  = \new_[53365]_  & \new_[53362]_ ;
  assign \new_[53369]_  = ~A269 & ~A268;
  assign \new_[53373]_  = ~A302 & ~A301;
  assign \new_[53374]_  = ~A300 & \new_[53373]_ ;
  assign \new_[53375]_  = \new_[53374]_  & \new_[53369]_ ;
  assign \new_[53376]_  = \new_[53375]_  & \new_[53366]_ ;
  assign \new_[53379]_  = ~A167 & A170;
  assign \new_[53382]_  = A199 & A166;
  assign \new_[53383]_  = \new_[53382]_  & \new_[53379]_ ;
  assign \new_[53386]_  = ~A201 & A200;
  assign \new_[53389]_  = A232 & ~A202;
  assign \new_[53390]_  = \new_[53389]_  & \new_[53386]_ ;
  assign \new_[53391]_  = \new_[53390]_  & \new_[53383]_ ;
  assign \new_[53394]_  = ~A234 & A233;
  assign \new_[53397]_  = ~A267 & ~A235;
  assign \new_[53398]_  = \new_[53397]_  & \new_[53394]_ ;
  assign \new_[53401]_  = ~A269 & ~A268;
  assign \new_[53405]_  = ~A301 & ~A299;
  assign \new_[53406]_  = ~A298 & \new_[53405]_ ;
  assign \new_[53407]_  = \new_[53406]_  & \new_[53401]_ ;
  assign \new_[53408]_  = \new_[53407]_  & \new_[53398]_ ;
  assign \new_[53411]_  = ~A167 & A170;
  assign \new_[53414]_  = A199 & A166;
  assign \new_[53415]_  = \new_[53414]_  & \new_[53411]_ ;
  assign \new_[53418]_  = ~A201 & A200;
  assign \new_[53421]_  = A232 & ~A202;
  assign \new_[53422]_  = \new_[53421]_  & \new_[53418]_ ;
  assign \new_[53423]_  = \new_[53422]_  & \new_[53415]_ ;
  assign \new_[53426]_  = ~A234 & A233;
  assign \new_[53429]_  = ~A265 & ~A235;
  assign \new_[53430]_  = \new_[53429]_  & \new_[53426]_ ;
  assign \new_[53433]_  = ~A268 & ~A266;
  assign \new_[53437]_  = ~A302 & ~A301;
  assign \new_[53438]_  = ~A300 & \new_[53437]_ ;
  assign \new_[53439]_  = \new_[53438]_  & \new_[53433]_ ;
  assign \new_[53440]_  = \new_[53439]_  & \new_[53430]_ ;
  assign \new_[53443]_  = ~A167 & A170;
  assign \new_[53446]_  = A199 & A166;
  assign \new_[53447]_  = \new_[53446]_  & \new_[53443]_ ;
  assign \new_[53450]_  = ~A201 & A200;
  assign \new_[53453]_  = A232 & ~A202;
  assign \new_[53454]_  = \new_[53453]_  & \new_[53450]_ ;
  assign \new_[53455]_  = \new_[53454]_  & \new_[53447]_ ;
  assign \new_[53458]_  = ~A234 & A233;
  assign \new_[53461]_  = ~A265 & ~A235;
  assign \new_[53462]_  = \new_[53461]_  & \new_[53458]_ ;
  assign \new_[53465]_  = ~A268 & ~A266;
  assign \new_[53469]_  = ~A301 & ~A299;
  assign \new_[53470]_  = ~A298 & \new_[53469]_ ;
  assign \new_[53471]_  = \new_[53470]_  & \new_[53465]_ ;
  assign \new_[53472]_  = \new_[53471]_  & \new_[53462]_ ;
  assign \new_[53475]_  = ~A167 & A170;
  assign \new_[53478]_  = A199 & A166;
  assign \new_[53479]_  = \new_[53478]_  & \new_[53475]_ ;
  assign \new_[53482]_  = ~A201 & A200;
  assign \new_[53485]_  = ~A232 & ~A202;
  assign \new_[53486]_  = \new_[53485]_  & \new_[53482]_ ;
  assign \new_[53487]_  = \new_[53486]_  & \new_[53479]_ ;
  assign \new_[53490]_  = ~A235 & ~A233;
  assign \new_[53493]_  = ~A268 & ~A267;
  assign \new_[53494]_  = \new_[53493]_  & \new_[53490]_ ;
  assign \new_[53497]_  = A298 & ~A269;
  assign \new_[53501]_  = ~A301 & ~A300;
  assign \new_[53502]_  = A299 & \new_[53501]_ ;
  assign \new_[53503]_  = \new_[53502]_  & \new_[53497]_ ;
  assign \new_[53504]_  = \new_[53503]_  & \new_[53494]_ ;
  assign \new_[53507]_  = ~A167 & A170;
  assign \new_[53510]_  = A199 & A166;
  assign \new_[53511]_  = \new_[53510]_  & \new_[53507]_ ;
  assign \new_[53514]_  = ~A201 & A200;
  assign \new_[53517]_  = ~A232 & ~A202;
  assign \new_[53518]_  = \new_[53517]_  & \new_[53514]_ ;
  assign \new_[53519]_  = \new_[53518]_  & \new_[53511]_ ;
  assign \new_[53522]_  = ~A235 & ~A233;
  assign \new_[53525]_  = A266 & A265;
  assign \new_[53526]_  = \new_[53525]_  & \new_[53522]_ ;
  assign \new_[53529]_  = ~A268 & ~A267;
  assign \new_[53533]_  = ~A302 & ~A301;
  assign \new_[53534]_  = ~A300 & \new_[53533]_ ;
  assign \new_[53535]_  = \new_[53534]_  & \new_[53529]_ ;
  assign \new_[53536]_  = \new_[53535]_  & \new_[53526]_ ;
  assign \new_[53539]_  = ~A167 & A170;
  assign \new_[53542]_  = A199 & A166;
  assign \new_[53543]_  = \new_[53542]_  & \new_[53539]_ ;
  assign \new_[53546]_  = ~A201 & A200;
  assign \new_[53549]_  = ~A232 & ~A202;
  assign \new_[53550]_  = \new_[53549]_  & \new_[53546]_ ;
  assign \new_[53551]_  = \new_[53550]_  & \new_[53543]_ ;
  assign \new_[53554]_  = ~A235 & ~A233;
  assign \new_[53557]_  = A266 & A265;
  assign \new_[53558]_  = \new_[53557]_  & \new_[53554]_ ;
  assign \new_[53561]_  = ~A268 & ~A267;
  assign \new_[53565]_  = ~A301 & ~A299;
  assign \new_[53566]_  = ~A298 & \new_[53565]_ ;
  assign \new_[53567]_  = \new_[53566]_  & \new_[53561]_ ;
  assign \new_[53568]_  = \new_[53567]_  & \new_[53558]_ ;
  assign \new_[53571]_  = ~A167 & A170;
  assign \new_[53574]_  = A199 & A166;
  assign \new_[53575]_  = \new_[53574]_  & \new_[53571]_ ;
  assign \new_[53578]_  = ~A201 & A200;
  assign \new_[53581]_  = ~A232 & ~A202;
  assign \new_[53582]_  = \new_[53581]_  & \new_[53578]_ ;
  assign \new_[53583]_  = \new_[53582]_  & \new_[53575]_ ;
  assign \new_[53586]_  = ~A235 & ~A233;
  assign \new_[53589]_  = ~A266 & ~A265;
  assign \new_[53590]_  = \new_[53589]_  & \new_[53586]_ ;
  assign \new_[53593]_  = A298 & ~A268;
  assign \new_[53597]_  = ~A301 & ~A300;
  assign \new_[53598]_  = A299 & \new_[53597]_ ;
  assign \new_[53599]_  = \new_[53598]_  & \new_[53593]_ ;
  assign \new_[53600]_  = \new_[53599]_  & \new_[53590]_ ;
  assign \new_[53603]_  = ~A167 & A170;
  assign \new_[53606]_  = ~A199 & A166;
  assign \new_[53607]_  = \new_[53606]_  & \new_[53603]_ ;
  assign \new_[53610]_  = ~A202 & ~A200;
  assign \new_[53613]_  = ~A235 & ~A234;
  assign \new_[53614]_  = \new_[53613]_  & \new_[53610]_ ;
  assign \new_[53615]_  = \new_[53614]_  & \new_[53607]_ ;
  assign \new_[53618]_  = A265 & ~A236;
  assign \new_[53621]_  = ~A267 & A266;
  assign \new_[53622]_  = \new_[53621]_  & \new_[53618]_ ;
  assign \new_[53625]_  = A298 & ~A268;
  assign \new_[53629]_  = ~A301 & ~A300;
  assign \new_[53630]_  = A299 & \new_[53629]_ ;
  assign \new_[53631]_  = \new_[53630]_  & \new_[53625]_ ;
  assign \new_[53632]_  = \new_[53631]_  & \new_[53622]_ ;
  assign \new_[53635]_  = ~A167 & A170;
  assign \new_[53638]_  = ~A199 & A166;
  assign \new_[53639]_  = \new_[53638]_  & \new_[53635]_ ;
  assign \new_[53642]_  = ~A202 & ~A200;
  assign \new_[53645]_  = A233 & A232;
  assign \new_[53646]_  = \new_[53645]_  & \new_[53642]_ ;
  assign \new_[53647]_  = \new_[53646]_  & \new_[53639]_ ;
  assign \new_[53650]_  = ~A235 & ~A234;
  assign \new_[53653]_  = ~A268 & ~A267;
  assign \new_[53654]_  = \new_[53653]_  & \new_[53650]_ ;
  assign \new_[53657]_  = A298 & ~A269;
  assign \new_[53661]_  = ~A301 & ~A300;
  assign \new_[53662]_  = A299 & \new_[53661]_ ;
  assign \new_[53663]_  = \new_[53662]_  & \new_[53657]_ ;
  assign \new_[53664]_  = \new_[53663]_  & \new_[53654]_ ;
  assign \new_[53667]_  = ~A167 & A170;
  assign \new_[53670]_  = ~A199 & A166;
  assign \new_[53671]_  = \new_[53670]_  & \new_[53667]_ ;
  assign \new_[53674]_  = ~A202 & ~A200;
  assign \new_[53677]_  = A233 & A232;
  assign \new_[53678]_  = \new_[53677]_  & \new_[53674]_ ;
  assign \new_[53679]_  = \new_[53678]_  & \new_[53671]_ ;
  assign \new_[53682]_  = ~A235 & ~A234;
  assign \new_[53685]_  = A266 & A265;
  assign \new_[53686]_  = \new_[53685]_  & \new_[53682]_ ;
  assign \new_[53689]_  = ~A268 & ~A267;
  assign \new_[53693]_  = ~A302 & ~A301;
  assign \new_[53694]_  = ~A300 & \new_[53693]_ ;
  assign \new_[53695]_  = \new_[53694]_  & \new_[53689]_ ;
  assign \new_[53696]_  = \new_[53695]_  & \new_[53686]_ ;
  assign \new_[53699]_  = ~A167 & A170;
  assign \new_[53702]_  = ~A199 & A166;
  assign \new_[53703]_  = \new_[53702]_  & \new_[53699]_ ;
  assign \new_[53706]_  = ~A202 & ~A200;
  assign \new_[53709]_  = A233 & A232;
  assign \new_[53710]_  = \new_[53709]_  & \new_[53706]_ ;
  assign \new_[53711]_  = \new_[53710]_  & \new_[53703]_ ;
  assign \new_[53714]_  = ~A235 & ~A234;
  assign \new_[53717]_  = A266 & A265;
  assign \new_[53718]_  = \new_[53717]_  & \new_[53714]_ ;
  assign \new_[53721]_  = ~A268 & ~A267;
  assign \new_[53725]_  = ~A301 & ~A299;
  assign \new_[53726]_  = ~A298 & \new_[53725]_ ;
  assign \new_[53727]_  = \new_[53726]_  & \new_[53721]_ ;
  assign \new_[53728]_  = \new_[53727]_  & \new_[53718]_ ;
  assign \new_[53731]_  = ~A167 & A170;
  assign \new_[53734]_  = ~A199 & A166;
  assign \new_[53735]_  = \new_[53734]_  & \new_[53731]_ ;
  assign \new_[53738]_  = ~A202 & ~A200;
  assign \new_[53741]_  = A233 & A232;
  assign \new_[53742]_  = \new_[53741]_  & \new_[53738]_ ;
  assign \new_[53743]_  = \new_[53742]_  & \new_[53735]_ ;
  assign \new_[53746]_  = ~A235 & ~A234;
  assign \new_[53749]_  = ~A266 & ~A265;
  assign \new_[53750]_  = \new_[53749]_  & \new_[53746]_ ;
  assign \new_[53753]_  = A298 & ~A268;
  assign \new_[53757]_  = ~A301 & ~A300;
  assign \new_[53758]_  = A299 & \new_[53757]_ ;
  assign \new_[53759]_  = \new_[53758]_  & \new_[53753]_ ;
  assign \new_[53760]_  = \new_[53759]_  & \new_[53750]_ ;
  assign \new_[53763]_  = ~A167 & A170;
  assign \new_[53766]_  = ~A199 & A166;
  assign \new_[53767]_  = \new_[53766]_  & \new_[53763]_ ;
  assign \new_[53770]_  = ~A202 & ~A200;
  assign \new_[53773]_  = ~A233 & ~A232;
  assign \new_[53774]_  = \new_[53773]_  & \new_[53770]_ ;
  assign \new_[53775]_  = \new_[53774]_  & \new_[53767]_ ;
  assign \new_[53778]_  = A265 & ~A235;
  assign \new_[53781]_  = ~A267 & A266;
  assign \new_[53782]_  = \new_[53781]_  & \new_[53778]_ ;
  assign \new_[53785]_  = A298 & ~A268;
  assign \new_[53789]_  = ~A301 & ~A300;
  assign \new_[53790]_  = A299 & \new_[53789]_ ;
  assign \new_[53791]_  = \new_[53790]_  & \new_[53785]_ ;
  assign \new_[53792]_  = \new_[53791]_  & \new_[53782]_ ;
  assign \new_[53795]_  = A199 & A169;
  assign \new_[53798]_  = ~A201 & A200;
  assign \new_[53799]_  = \new_[53798]_  & \new_[53795]_ ;
  assign \new_[53802]_  = A232 & ~A202;
  assign \new_[53805]_  = ~A234 & A233;
  assign \new_[53806]_  = \new_[53805]_  & \new_[53802]_ ;
  assign \new_[53807]_  = \new_[53806]_  & \new_[53799]_ ;
  assign \new_[53810]_  = A265 & ~A235;
  assign \new_[53813]_  = ~A267 & A266;
  assign \new_[53814]_  = \new_[53813]_  & \new_[53810]_ ;
  assign \new_[53817]_  = A298 & ~A268;
  assign \new_[53821]_  = ~A301 & ~A300;
  assign \new_[53822]_  = A299 & \new_[53821]_ ;
  assign \new_[53823]_  = \new_[53822]_  & \new_[53817]_ ;
  assign \new_[53824]_  = \new_[53823]_  & \new_[53814]_ ;
  assign \new_[53827]_  = ~A167 & ~A169;
  assign \new_[53830]_  = A199 & ~A166;
  assign \new_[53831]_  = \new_[53830]_  & \new_[53827]_ ;
  assign \new_[53834]_  = A232 & A201;
  assign \new_[53837]_  = ~A234 & A233;
  assign \new_[53838]_  = \new_[53837]_  & \new_[53834]_ ;
  assign \new_[53839]_  = \new_[53838]_  & \new_[53831]_ ;
  assign \new_[53842]_  = A265 & ~A235;
  assign \new_[53845]_  = ~A267 & A266;
  assign \new_[53846]_  = \new_[53845]_  & \new_[53842]_ ;
  assign \new_[53849]_  = A298 & ~A268;
  assign \new_[53853]_  = ~A301 & ~A300;
  assign \new_[53854]_  = A299 & \new_[53853]_ ;
  assign \new_[53855]_  = \new_[53854]_  & \new_[53849]_ ;
  assign \new_[53856]_  = \new_[53855]_  & \new_[53846]_ ;
  assign \new_[53859]_  = ~A167 & ~A169;
  assign \new_[53862]_  = A200 & ~A166;
  assign \new_[53863]_  = \new_[53862]_  & \new_[53859]_ ;
  assign \new_[53866]_  = A232 & A201;
  assign \new_[53869]_  = ~A234 & A233;
  assign \new_[53870]_  = \new_[53869]_  & \new_[53866]_ ;
  assign \new_[53871]_  = \new_[53870]_  & \new_[53863]_ ;
  assign \new_[53874]_  = A265 & ~A235;
  assign \new_[53877]_  = ~A267 & A266;
  assign \new_[53878]_  = \new_[53877]_  & \new_[53874]_ ;
  assign \new_[53881]_  = A298 & ~A268;
  assign \new_[53885]_  = ~A301 & ~A300;
  assign \new_[53886]_  = A299 & \new_[53885]_ ;
  assign \new_[53887]_  = \new_[53886]_  & \new_[53881]_ ;
  assign \new_[53888]_  = \new_[53887]_  & \new_[53878]_ ;
  assign \new_[53891]_  = ~A167 & ~A169;
  assign \new_[53894]_  = ~A199 & ~A166;
  assign \new_[53895]_  = \new_[53894]_  & \new_[53891]_ ;
  assign \new_[53898]_  = A203 & A200;
  assign \new_[53901]_  = ~A235 & ~A234;
  assign \new_[53902]_  = \new_[53901]_  & \new_[53898]_ ;
  assign \new_[53903]_  = \new_[53902]_  & \new_[53895]_ ;
  assign \new_[53906]_  = A265 & ~A236;
  assign \new_[53909]_  = ~A267 & A266;
  assign \new_[53910]_  = \new_[53909]_  & \new_[53906]_ ;
  assign \new_[53913]_  = A298 & ~A268;
  assign \new_[53917]_  = ~A301 & ~A300;
  assign \new_[53918]_  = A299 & \new_[53917]_ ;
  assign \new_[53919]_  = \new_[53918]_  & \new_[53913]_ ;
  assign \new_[53920]_  = \new_[53919]_  & \new_[53910]_ ;
  assign \new_[53923]_  = ~A167 & ~A169;
  assign \new_[53926]_  = ~A199 & ~A166;
  assign \new_[53927]_  = \new_[53926]_  & \new_[53923]_ ;
  assign \new_[53930]_  = A203 & A200;
  assign \new_[53933]_  = A233 & A232;
  assign \new_[53934]_  = \new_[53933]_  & \new_[53930]_ ;
  assign \new_[53935]_  = \new_[53934]_  & \new_[53927]_ ;
  assign \new_[53938]_  = ~A235 & ~A234;
  assign \new_[53941]_  = ~A268 & ~A267;
  assign \new_[53942]_  = \new_[53941]_  & \new_[53938]_ ;
  assign \new_[53945]_  = A298 & ~A269;
  assign \new_[53949]_  = ~A301 & ~A300;
  assign \new_[53950]_  = A299 & \new_[53949]_ ;
  assign \new_[53951]_  = \new_[53950]_  & \new_[53945]_ ;
  assign \new_[53952]_  = \new_[53951]_  & \new_[53942]_ ;
  assign \new_[53955]_  = ~A167 & ~A169;
  assign \new_[53958]_  = ~A199 & ~A166;
  assign \new_[53959]_  = \new_[53958]_  & \new_[53955]_ ;
  assign \new_[53962]_  = A203 & A200;
  assign \new_[53965]_  = A233 & A232;
  assign \new_[53966]_  = \new_[53965]_  & \new_[53962]_ ;
  assign \new_[53967]_  = \new_[53966]_  & \new_[53959]_ ;
  assign \new_[53970]_  = ~A235 & ~A234;
  assign \new_[53973]_  = A266 & A265;
  assign \new_[53974]_  = \new_[53973]_  & \new_[53970]_ ;
  assign \new_[53977]_  = ~A268 & ~A267;
  assign \new_[53981]_  = ~A302 & ~A301;
  assign \new_[53982]_  = ~A300 & \new_[53981]_ ;
  assign \new_[53983]_  = \new_[53982]_  & \new_[53977]_ ;
  assign \new_[53984]_  = \new_[53983]_  & \new_[53974]_ ;
  assign \new_[53987]_  = ~A167 & ~A169;
  assign \new_[53990]_  = ~A199 & ~A166;
  assign \new_[53991]_  = \new_[53990]_  & \new_[53987]_ ;
  assign \new_[53994]_  = A203 & A200;
  assign \new_[53997]_  = A233 & A232;
  assign \new_[53998]_  = \new_[53997]_  & \new_[53994]_ ;
  assign \new_[53999]_  = \new_[53998]_  & \new_[53991]_ ;
  assign \new_[54002]_  = ~A235 & ~A234;
  assign \new_[54005]_  = A266 & A265;
  assign \new_[54006]_  = \new_[54005]_  & \new_[54002]_ ;
  assign \new_[54009]_  = ~A268 & ~A267;
  assign \new_[54013]_  = ~A301 & ~A299;
  assign \new_[54014]_  = ~A298 & \new_[54013]_ ;
  assign \new_[54015]_  = \new_[54014]_  & \new_[54009]_ ;
  assign \new_[54016]_  = \new_[54015]_  & \new_[54006]_ ;
  assign \new_[54019]_  = ~A167 & ~A169;
  assign \new_[54022]_  = ~A199 & ~A166;
  assign \new_[54023]_  = \new_[54022]_  & \new_[54019]_ ;
  assign \new_[54026]_  = A203 & A200;
  assign \new_[54029]_  = A233 & A232;
  assign \new_[54030]_  = \new_[54029]_  & \new_[54026]_ ;
  assign \new_[54031]_  = \new_[54030]_  & \new_[54023]_ ;
  assign \new_[54034]_  = ~A235 & ~A234;
  assign \new_[54037]_  = ~A266 & ~A265;
  assign \new_[54038]_  = \new_[54037]_  & \new_[54034]_ ;
  assign \new_[54041]_  = A298 & ~A268;
  assign \new_[54045]_  = ~A301 & ~A300;
  assign \new_[54046]_  = A299 & \new_[54045]_ ;
  assign \new_[54047]_  = \new_[54046]_  & \new_[54041]_ ;
  assign \new_[54048]_  = \new_[54047]_  & \new_[54038]_ ;
  assign \new_[54051]_  = ~A167 & ~A169;
  assign \new_[54054]_  = ~A199 & ~A166;
  assign \new_[54055]_  = \new_[54054]_  & \new_[54051]_ ;
  assign \new_[54058]_  = A203 & A200;
  assign \new_[54061]_  = ~A233 & ~A232;
  assign \new_[54062]_  = \new_[54061]_  & \new_[54058]_ ;
  assign \new_[54063]_  = \new_[54062]_  & \new_[54055]_ ;
  assign \new_[54066]_  = A265 & ~A235;
  assign \new_[54069]_  = ~A267 & A266;
  assign \new_[54070]_  = \new_[54069]_  & \new_[54066]_ ;
  assign \new_[54073]_  = A298 & ~A268;
  assign \new_[54077]_  = ~A301 & ~A300;
  assign \new_[54078]_  = A299 & \new_[54077]_ ;
  assign \new_[54079]_  = \new_[54078]_  & \new_[54073]_ ;
  assign \new_[54080]_  = \new_[54079]_  & \new_[54070]_ ;
  assign \new_[54083]_  = ~A167 & ~A169;
  assign \new_[54086]_  = A199 & ~A166;
  assign \new_[54087]_  = \new_[54086]_  & \new_[54083]_ ;
  assign \new_[54090]_  = A203 & ~A200;
  assign \new_[54093]_  = ~A235 & ~A234;
  assign \new_[54094]_  = \new_[54093]_  & \new_[54090]_ ;
  assign \new_[54095]_  = \new_[54094]_  & \new_[54087]_ ;
  assign \new_[54098]_  = A265 & ~A236;
  assign \new_[54101]_  = ~A267 & A266;
  assign \new_[54102]_  = \new_[54101]_  & \new_[54098]_ ;
  assign \new_[54105]_  = A298 & ~A268;
  assign \new_[54109]_  = ~A301 & ~A300;
  assign \new_[54110]_  = A299 & \new_[54109]_ ;
  assign \new_[54111]_  = \new_[54110]_  & \new_[54105]_ ;
  assign \new_[54112]_  = \new_[54111]_  & \new_[54102]_ ;
  assign \new_[54115]_  = ~A167 & ~A169;
  assign \new_[54118]_  = A199 & ~A166;
  assign \new_[54119]_  = \new_[54118]_  & \new_[54115]_ ;
  assign \new_[54122]_  = A203 & ~A200;
  assign \new_[54125]_  = A233 & A232;
  assign \new_[54126]_  = \new_[54125]_  & \new_[54122]_ ;
  assign \new_[54127]_  = \new_[54126]_  & \new_[54119]_ ;
  assign \new_[54130]_  = ~A235 & ~A234;
  assign \new_[54133]_  = ~A268 & ~A267;
  assign \new_[54134]_  = \new_[54133]_  & \new_[54130]_ ;
  assign \new_[54137]_  = A298 & ~A269;
  assign \new_[54141]_  = ~A301 & ~A300;
  assign \new_[54142]_  = A299 & \new_[54141]_ ;
  assign \new_[54143]_  = \new_[54142]_  & \new_[54137]_ ;
  assign \new_[54144]_  = \new_[54143]_  & \new_[54134]_ ;
  assign \new_[54147]_  = ~A167 & ~A169;
  assign \new_[54150]_  = A199 & ~A166;
  assign \new_[54151]_  = \new_[54150]_  & \new_[54147]_ ;
  assign \new_[54154]_  = A203 & ~A200;
  assign \new_[54157]_  = A233 & A232;
  assign \new_[54158]_  = \new_[54157]_  & \new_[54154]_ ;
  assign \new_[54159]_  = \new_[54158]_  & \new_[54151]_ ;
  assign \new_[54162]_  = ~A235 & ~A234;
  assign \new_[54165]_  = A266 & A265;
  assign \new_[54166]_  = \new_[54165]_  & \new_[54162]_ ;
  assign \new_[54169]_  = ~A268 & ~A267;
  assign \new_[54173]_  = ~A302 & ~A301;
  assign \new_[54174]_  = ~A300 & \new_[54173]_ ;
  assign \new_[54175]_  = \new_[54174]_  & \new_[54169]_ ;
  assign \new_[54176]_  = \new_[54175]_  & \new_[54166]_ ;
  assign \new_[54179]_  = ~A167 & ~A169;
  assign \new_[54182]_  = A199 & ~A166;
  assign \new_[54183]_  = \new_[54182]_  & \new_[54179]_ ;
  assign \new_[54186]_  = A203 & ~A200;
  assign \new_[54189]_  = A233 & A232;
  assign \new_[54190]_  = \new_[54189]_  & \new_[54186]_ ;
  assign \new_[54191]_  = \new_[54190]_  & \new_[54183]_ ;
  assign \new_[54194]_  = ~A235 & ~A234;
  assign \new_[54197]_  = A266 & A265;
  assign \new_[54198]_  = \new_[54197]_  & \new_[54194]_ ;
  assign \new_[54201]_  = ~A268 & ~A267;
  assign \new_[54205]_  = ~A301 & ~A299;
  assign \new_[54206]_  = ~A298 & \new_[54205]_ ;
  assign \new_[54207]_  = \new_[54206]_  & \new_[54201]_ ;
  assign \new_[54208]_  = \new_[54207]_  & \new_[54198]_ ;
  assign \new_[54211]_  = ~A167 & ~A169;
  assign \new_[54214]_  = A199 & ~A166;
  assign \new_[54215]_  = \new_[54214]_  & \new_[54211]_ ;
  assign \new_[54218]_  = A203 & ~A200;
  assign \new_[54221]_  = A233 & A232;
  assign \new_[54222]_  = \new_[54221]_  & \new_[54218]_ ;
  assign \new_[54223]_  = \new_[54222]_  & \new_[54215]_ ;
  assign \new_[54226]_  = ~A235 & ~A234;
  assign \new_[54229]_  = ~A266 & ~A265;
  assign \new_[54230]_  = \new_[54229]_  & \new_[54226]_ ;
  assign \new_[54233]_  = A298 & ~A268;
  assign \new_[54237]_  = ~A301 & ~A300;
  assign \new_[54238]_  = A299 & \new_[54237]_ ;
  assign \new_[54239]_  = \new_[54238]_  & \new_[54233]_ ;
  assign \new_[54240]_  = \new_[54239]_  & \new_[54230]_ ;
  assign \new_[54243]_  = ~A167 & ~A169;
  assign \new_[54246]_  = A199 & ~A166;
  assign \new_[54247]_  = \new_[54246]_  & \new_[54243]_ ;
  assign \new_[54250]_  = A203 & ~A200;
  assign \new_[54253]_  = ~A233 & ~A232;
  assign \new_[54254]_  = \new_[54253]_  & \new_[54250]_ ;
  assign \new_[54255]_  = \new_[54254]_  & \new_[54247]_ ;
  assign \new_[54258]_  = A265 & ~A235;
  assign \new_[54261]_  = ~A267 & A266;
  assign \new_[54262]_  = \new_[54261]_  & \new_[54258]_ ;
  assign \new_[54265]_  = A298 & ~A268;
  assign \new_[54269]_  = ~A301 & ~A300;
  assign \new_[54270]_  = A299 & \new_[54269]_ ;
  assign \new_[54271]_  = \new_[54270]_  & \new_[54265]_ ;
  assign \new_[54272]_  = \new_[54271]_  & \new_[54262]_ ;
  assign \new_[54275]_  = ~A168 & ~A169;
  assign \new_[54278]_  = A166 & A167;
  assign \new_[54279]_  = \new_[54278]_  & \new_[54275]_ ;
  assign \new_[54282]_  = A232 & A202;
  assign \new_[54285]_  = ~A234 & A233;
  assign \new_[54286]_  = \new_[54285]_  & \new_[54282]_ ;
  assign \new_[54287]_  = \new_[54286]_  & \new_[54279]_ ;
  assign \new_[54290]_  = A265 & ~A235;
  assign \new_[54293]_  = ~A267 & A266;
  assign \new_[54294]_  = \new_[54293]_  & \new_[54290]_ ;
  assign \new_[54297]_  = A298 & ~A268;
  assign \new_[54301]_  = ~A301 & ~A300;
  assign \new_[54302]_  = A299 & \new_[54301]_ ;
  assign \new_[54303]_  = \new_[54302]_  & \new_[54297]_ ;
  assign \new_[54304]_  = \new_[54303]_  & \new_[54294]_ ;
  assign \new_[54307]_  = ~A168 & ~A169;
  assign \new_[54310]_  = A166 & A167;
  assign \new_[54311]_  = \new_[54310]_  & \new_[54307]_ ;
  assign \new_[54314]_  = A201 & A199;
  assign \new_[54317]_  = ~A235 & ~A234;
  assign \new_[54318]_  = \new_[54317]_  & \new_[54314]_ ;
  assign \new_[54319]_  = \new_[54318]_  & \new_[54311]_ ;
  assign \new_[54322]_  = A265 & ~A236;
  assign \new_[54325]_  = ~A267 & A266;
  assign \new_[54326]_  = \new_[54325]_  & \new_[54322]_ ;
  assign \new_[54329]_  = A298 & ~A268;
  assign \new_[54333]_  = ~A301 & ~A300;
  assign \new_[54334]_  = A299 & \new_[54333]_ ;
  assign \new_[54335]_  = \new_[54334]_  & \new_[54329]_ ;
  assign \new_[54336]_  = \new_[54335]_  & \new_[54326]_ ;
  assign \new_[54339]_  = ~A168 & ~A169;
  assign \new_[54342]_  = A166 & A167;
  assign \new_[54343]_  = \new_[54342]_  & \new_[54339]_ ;
  assign \new_[54346]_  = A201 & A199;
  assign \new_[54349]_  = A233 & A232;
  assign \new_[54350]_  = \new_[54349]_  & \new_[54346]_ ;
  assign \new_[54351]_  = \new_[54350]_  & \new_[54343]_ ;
  assign \new_[54354]_  = ~A235 & ~A234;
  assign \new_[54357]_  = ~A268 & ~A267;
  assign \new_[54358]_  = \new_[54357]_  & \new_[54354]_ ;
  assign \new_[54361]_  = A298 & ~A269;
  assign \new_[54365]_  = ~A301 & ~A300;
  assign \new_[54366]_  = A299 & \new_[54365]_ ;
  assign \new_[54367]_  = \new_[54366]_  & \new_[54361]_ ;
  assign \new_[54368]_  = \new_[54367]_  & \new_[54358]_ ;
  assign \new_[54371]_  = ~A168 & ~A169;
  assign \new_[54374]_  = A166 & A167;
  assign \new_[54375]_  = \new_[54374]_  & \new_[54371]_ ;
  assign \new_[54378]_  = A201 & A199;
  assign \new_[54381]_  = A233 & A232;
  assign \new_[54382]_  = \new_[54381]_  & \new_[54378]_ ;
  assign \new_[54383]_  = \new_[54382]_  & \new_[54375]_ ;
  assign \new_[54386]_  = ~A235 & ~A234;
  assign \new_[54389]_  = A266 & A265;
  assign \new_[54390]_  = \new_[54389]_  & \new_[54386]_ ;
  assign \new_[54393]_  = ~A268 & ~A267;
  assign \new_[54397]_  = ~A302 & ~A301;
  assign \new_[54398]_  = ~A300 & \new_[54397]_ ;
  assign \new_[54399]_  = \new_[54398]_  & \new_[54393]_ ;
  assign \new_[54400]_  = \new_[54399]_  & \new_[54390]_ ;
  assign \new_[54403]_  = ~A168 & ~A169;
  assign \new_[54406]_  = A166 & A167;
  assign \new_[54407]_  = \new_[54406]_  & \new_[54403]_ ;
  assign \new_[54410]_  = A201 & A199;
  assign \new_[54413]_  = A233 & A232;
  assign \new_[54414]_  = \new_[54413]_  & \new_[54410]_ ;
  assign \new_[54415]_  = \new_[54414]_  & \new_[54407]_ ;
  assign \new_[54418]_  = ~A235 & ~A234;
  assign \new_[54421]_  = A266 & A265;
  assign \new_[54422]_  = \new_[54421]_  & \new_[54418]_ ;
  assign \new_[54425]_  = ~A268 & ~A267;
  assign \new_[54429]_  = ~A301 & ~A299;
  assign \new_[54430]_  = ~A298 & \new_[54429]_ ;
  assign \new_[54431]_  = \new_[54430]_  & \new_[54425]_ ;
  assign \new_[54432]_  = \new_[54431]_  & \new_[54422]_ ;
  assign \new_[54435]_  = ~A168 & ~A169;
  assign \new_[54438]_  = A166 & A167;
  assign \new_[54439]_  = \new_[54438]_  & \new_[54435]_ ;
  assign \new_[54442]_  = A201 & A199;
  assign \new_[54445]_  = A233 & A232;
  assign \new_[54446]_  = \new_[54445]_  & \new_[54442]_ ;
  assign \new_[54447]_  = \new_[54446]_  & \new_[54439]_ ;
  assign \new_[54450]_  = ~A235 & ~A234;
  assign \new_[54453]_  = ~A266 & ~A265;
  assign \new_[54454]_  = \new_[54453]_  & \new_[54450]_ ;
  assign \new_[54457]_  = A298 & ~A268;
  assign \new_[54461]_  = ~A301 & ~A300;
  assign \new_[54462]_  = A299 & \new_[54461]_ ;
  assign \new_[54463]_  = \new_[54462]_  & \new_[54457]_ ;
  assign \new_[54464]_  = \new_[54463]_  & \new_[54454]_ ;
  assign \new_[54467]_  = ~A168 & ~A169;
  assign \new_[54470]_  = A166 & A167;
  assign \new_[54471]_  = \new_[54470]_  & \new_[54467]_ ;
  assign \new_[54474]_  = A201 & A199;
  assign \new_[54477]_  = ~A233 & ~A232;
  assign \new_[54478]_  = \new_[54477]_  & \new_[54474]_ ;
  assign \new_[54479]_  = \new_[54478]_  & \new_[54471]_ ;
  assign \new_[54482]_  = A265 & ~A235;
  assign \new_[54485]_  = ~A267 & A266;
  assign \new_[54486]_  = \new_[54485]_  & \new_[54482]_ ;
  assign \new_[54489]_  = A298 & ~A268;
  assign \new_[54493]_  = ~A301 & ~A300;
  assign \new_[54494]_  = A299 & \new_[54493]_ ;
  assign \new_[54495]_  = \new_[54494]_  & \new_[54489]_ ;
  assign \new_[54496]_  = \new_[54495]_  & \new_[54486]_ ;
  assign \new_[54499]_  = ~A168 & ~A169;
  assign \new_[54502]_  = A166 & A167;
  assign \new_[54503]_  = \new_[54502]_  & \new_[54499]_ ;
  assign \new_[54506]_  = A201 & A200;
  assign \new_[54509]_  = ~A235 & ~A234;
  assign \new_[54510]_  = \new_[54509]_  & \new_[54506]_ ;
  assign \new_[54511]_  = \new_[54510]_  & \new_[54503]_ ;
  assign \new_[54514]_  = A265 & ~A236;
  assign \new_[54517]_  = ~A267 & A266;
  assign \new_[54518]_  = \new_[54517]_  & \new_[54514]_ ;
  assign \new_[54521]_  = A298 & ~A268;
  assign \new_[54525]_  = ~A301 & ~A300;
  assign \new_[54526]_  = A299 & \new_[54525]_ ;
  assign \new_[54527]_  = \new_[54526]_  & \new_[54521]_ ;
  assign \new_[54528]_  = \new_[54527]_  & \new_[54518]_ ;
  assign \new_[54531]_  = ~A168 & ~A169;
  assign \new_[54534]_  = A166 & A167;
  assign \new_[54535]_  = \new_[54534]_  & \new_[54531]_ ;
  assign \new_[54538]_  = A201 & A200;
  assign \new_[54541]_  = A233 & A232;
  assign \new_[54542]_  = \new_[54541]_  & \new_[54538]_ ;
  assign \new_[54543]_  = \new_[54542]_  & \new_[54535]_ ;
  assign \new_[54546]_  = ~A235 & ~A234;
  assign \new_[54549]_  = ~A268 & ~A267;
  assign \new_[54550]_  = \new_[54549]_  & \new_[54546]_ ;
  assign \new_[54553]_  = A298 & ~A269;
  assign \new_[54557]_  = ~A301 & ~A300;
  assign \new_[54558]_  = A299 & \new_[54557]_ ;
  assign \new_[54559]_  = \new_[54558]_  & \new_[54553]_ ;
  assign \new_[54560]_  = \new_[54559]_  & \new_[54550]_ ;
  assign \new_[54563]_  = ~A168 & ~A169;
  assign \new_[54566]_  = A166 & A167;
  assign \new_[54567]_  = \new_[54566]_  & \new_[54563]_ ;
  assign \new_[54570]_  = A201 & A200;
  assign \new_[54573]_  = A233 & A232;
  assign \new_[54574]_  = \new_[54573]_  & \new_[54570]_ ;
  assign \new_[54575]_  = \new_[54574]_  & \new_[54567]_ ;
  assign \new_[54578]_  = ~A235 & ~A234;
  assign \new_[54581]_  = A266 & A265;
  assign \new_[54582]_  = \new_[54581]_  & \new_[54578]_ ;
  assign \new_[54585]_  = ~A268 & ~A267;
  assign \new_[54589]_  = ~A302 & ~A301;
  assign \new_[54590]_  = ~A300 & \new_[54589]_ ;
  assign \new_[54591]_  = \new_[54590]_  & \new_[54585]_ ;
  assign \new_[54592]_  = \new_[54591]_  & \new_[54582]_ ;
  assign \new_[54595]_  = ~A168 & ~A169;
  assign \new_[54598]_  = A166 & A167;
  assign \new_[54599]_  = \new_[54598]_  & \new_[54595]_ ;
  assign \new_[54602]_  = A201 & A200;
  assign \new_[54605]_  = A233 & A232;
  assign \new_[54606]_  = \new_[54605]_  & \new_[54602]_ ;
  assign \new_[54607]_  = \new_[54606]_  & \new_[54599]_ ;
  assign \new_[54610]_  = ~A235 & ~A234;
  assign \new_[54613]_  = A266 & A265;
  assign \new_[54614]_  = \new_[54613]_  & \new_[54610]_ ;
  assign \new_[54617]_  = ~A268 & ~A267;
  assign \new_[54621]_  = ~A301 & ~A299;
  assign \new_[54622]_  = ~A298 & \new_[54621]_ ;
  assign \new_[54623]_  = \new_[54622]_  & \new_[54617]_ ;
  assign \new_[54624]_  = \new_[54623]_  & \new_[54614]_ ;
  assign \new_[54627]_  = ~A168 & ~A169;
  assign \new_[54630]_  = A166 & A167;
  assign \new_[54631]_  = \new_[54630]_  & \new_[54627]_ ;
  assign \new_[54634]_  = A201 & A200;
  assign \new_[54637]_  = A233 & A232;
  assign \new_[54638]_  = \new_[54637]_  & \new_[54634]_ ;
  assign \new_[54639]_  = \new_[54638]_  & \new_[54631]_ ;
  assign \new_[54642]_  = ~A235 & ~A234;
  assign \new_[54645]_  = ~A266 & ~A265;
  assign \new_[54646]_  = \new_[54645]_  & \new_[54642]_ ;
  assign \new_[54649]_  = A298 & ~A268;
  assign \new_[54653]_  = ~A301 & ~A300;
  assign \new_[54654]_  = A299 & \new_[54653]_ ;
  assign \new_[54655]_  = \new_[54654]_  & \new_[54649]_ ;
  assign \new_[54656]_  = \new_[54655]_  & \new_[54646]_ ;
  assign \new_[54659]_  = ~A168 & ~A169;
  assign \new_[54662]_  = A166 & A167;
  assign \new_[54663]_  = \new_[54662]_  & \new_[54659]_ ;
  assign \new_[54666]_  = A201 & A200;
  assign \new_[54669]_  = ~A233 & ~A232;
  assign \new_[54670]_  = \new_[54669]_  & \new_[54666]_ ;
  assign \new_[54671]_  = \new_[54670]_  & \new_[54663]_ ;
  assign \new_[54674]_  = A265 & ~A235;
  assign \new_[54677]_  = ~A267 & A266;
  assign \new_[54678]_  = \new_[54677]_  & \new_[54674]_ ;
  assign \new_[54681]_  = A298 & ~A268;
  assign \new_[54685]_  = ~A301 & ~A300;
  assign \new_[54686]_  = A299 & \new_[54685]_ ;
  assign \new_[54687]_  = \new_[54686]_  & \new_[54681]_ ;
  assign \new_[54688]_  = \new_[54687]_  & \new_[54678]_ ;
  assign \new_[54691]_  = ~A168 & ~A169;
  assign \new_[54694]_  = A166 & A167;
  assign \new_[54695]_  = \new_[54694]_  & \new_[54691]_ ;
  assign \new_[54698]_  = A200 & ~A199;
  assign \new_[54701]_  = ~A234 & A203;
  assign \new_[54702]_  = \new_[54701]_  & \new_[54698]_ ;
  assign \new_[54703]_  = \new_[54702]_  & \new_[54695]_ ;
  assign \new_[54706]_  = ~A236 & ~A235;
  assign \new_[54709]_  = ~A268 & ~A267;
  assign \new_[54710]_  = \new_[54709]_  & \new_[54706]_ ;
  assign \new_[54713]_  = A298 & ~A269;
  assign \new_[54717]_  = ~A301 & ~A300;
  assign \new_[54718]_  = A299 & \new_[54717]_ ;
  assign \new_[54719]_  = \new_[54718]_  & \new_[54713]_ ;
  assign \new_[54720]_  = \new_[54719]_  & \new_[54710]_ ;
  assign \new_[54723]_  = ~A168 & ~A169;
  assign \new_[54726]_  = A166 & A167;
  assign \new_[54727]_  = \new_[54726]_  & \new_[54723]_ ;
  assign \new_[54730]_  = A200 & ~A199;
  assign \new_[54733]_  = ~A234 & A203;
  assign \new_[54734]_  = \new_[54733]_  & \new_[54730]_ ;
  assign \new_[54735]_  = \new_[54734]_  & \new_[54727]_ ;
  assign \new_[54738]_  = ~A236 & ~A235;
  assign \new_[54741]_  = A266 & A265;
  assign \new_[54742]_  = \new_[54741]_  & \new_[54738]_ ;
  assign \new_[54745]_  = ~A268 & ~A267;
  assign \new_[54749]_  = ~A302 & ~A301;
  assign \new_[54750]_  = ~A300 & \new_[54749]_ ;
  assign \new_[54751]_  = \new_[54750]_  & \new_[54745]_ ;
  assign \new_[54752]_  = \new_[54751]_  & \new_[54742]_ ;
  assign \new_[54755]_  = ~A168 & ~A169;
  assign \new_[54758]_  = A166 & A167;
  assign \new_[54759]_  = \new_[54758]_  & \new_[54755]_ ;
  assign \new_[54762]_  = A200 & ~A199;
  assign \new_[54765]_  = ~A234 & A203;
  assign \new_[54766]_  = \new_[54765]_  & \new_[54762]_ ;
  assign \new_[54767]_  = \new_[54766]_  & \new_[54759]_ ;
  assign \new_[54770]_  = ~A236 & ~A235;
  assign \new_[54773]_  = A266 & A265;
  assign \new_[54774]_  = \new_[54773]_  & \new_[54770]_ ;
  assign \new_[54777]_  = ~A268 & ~A267;
  assign \new_[54781]_  = ~A301 & ~A299;
  assign \new_[54782]_  = ~A298 & \new_[54781]_ ;
  assign \new_[54783]_  = \new_[54782]_  & \new_[54777]_ ;
  assign \new_[54784]_  = \new_[54783]_  & \new_[54774]_ ;
  assign \new_[54787]_  = ~A168 & ~A169;
  assign \new_[54790]_  = A166 & A167;
  assign \new_[54791]_  = \new_[54790]_  & \new_[54787]_ ;
  assign \new_[54794]_  = A200 & ~A199;
  assign \new_[54797]_  = ~A234 & A203;
  assign \new_[54798]_  = \new_[54797]_  & \new_[54794]_ ;
  assign \new_[54799]_  = \new_[54798]_  & \new_[54791]_ ;
  assign \new_[54802]_  = ~A236 & ~A235;
  assign \new_[54805]_  = ~A266 & ~A265;
  assign \new_[54806]_  = \new_[54805]_  & \new_[54802]_ ;
  assign \new_[54809]_  = A298 & ~A268;
  assign \new_[54813]_  = ~A301 & ~A300;
  assign \new_[54814]_  = A299 & \new_[54813]_ ;
  assign \new_[54815]_  = \new_[54814]_  & \new_[54809]_ ;
  assign \new_[54816]_  = \new_[54815]_  & \new_[54806]_ ;
  assign \new_[54819]_  = ~A168 & ~A169;
  assign \new_[54822]_  = A166 & A167;
  assign \new_[54823]_  = \new_[54822]_  & \new_[54819]_ ;
  assign \new_[54826]_  = A200 & ~A199;
  assign \new_[54829]_  = A232 & A203;
  assign \new_[54830]_  = \new_[54829]_  & \new_[54826]_ ;
  assign \new_[54831]_  = \new_[54830]_  & \new_[54823]_ ;
  assign \new_[54834]_  = ~A234 & A233;
  assign \new_[54837]_  = ~A267 & ~A235;
  assign \new_[54838]_  = \new_[54837]_  & \new_[54834]_ ;
  assign \new_[54841]_  = ~A269 & ~A268;
  assign \new_[54845]_  = ~A302 & ~A301;
  assign \new_[54846]_  = ~A300 & \new_[54845]_ ;
  assign \new_[54847]_  = \new_[54846]_  & \new_[54841]_ ;
  assign \new_[54848]_  = \new_[54847]_  & \new_[54838]_ ;
  assign \new_[54851]_  = ~A168 & ~A169;
  assign \new_[54854]_  = A166 & A167;
  assign \new_[54855]_  = \new_[54854]_  & \new_[54851]_ ;
  assign \new_[54858]_  = A200 & ~A199;
  assign \new_[54861]_  = A232 & A203;
  assign \new_[54862]_  = \new_[54861]_  & \new_[54858]_ ;
  assign \new_[54863]_  = \new_[54862]_  & \new_[54855]_ ;
  assign \new_[54866]_  = ~A234 & A233;
  assign \new_[54869]_  = ~A267 & ~A235;
  assign \new_[54870]_  = \new_[54869]_  & \new_[54866]_ ;
  assign \new_[54873]_  = ~A269 & ~A268;
  assign \new_[54877]_  = ~A301 & ~A299;
  assign \new_[54878]_  = ~A298 & \new_[54877]_ ;
  assign \new_[54879]_  = \new_[54878]_  & \new_[54873]_ ;
  assign \new_[54880]_  = \new_[54879]_  & \new_[54870]_ ;
  assign \new_[54883]_  = ~A168 & ~A169;
  assign \new_[54886]_  = A166 & A167;
  assign \new_[54887]_  = \new_[54886]_  & \new_[54883]_ ;
  assign \new_[54890]_  = A200 & ~A199;
  assign \new_[54893]_  = A232 & A203;
  assign \new_[54894]_  = \new_[54893]_  & \new_[54890]_ ;
  assign \new_[54895]_  = \new_[54894]_  & \new_[54887]_ ;
  assign \new_[54898]_  = ~A234 & A233;
  assign \new_[54901]_  = ~A265 & ~A235;
  assign \new_[54902]_  = \new_[54901]_  & \new_[54898]_ ;
  assign \new_[54905]_  = ~A268 & ~A266;
  assign \new_[54909]_  = ~A302 & ~A301;
  assign \new_[54910]_  = ~A300 & \new_[54909]_ ;
  assign \new_[54911]_  = \new_[54910]_  & \new_[54905]_ ;
  assign \new_[54912]_  = \new_[54911]_  & \new_[54902]_ ;
  assign \new_[54915]_  = ~A168 & ~A169;
  assign \new_[54918]_  = A166 & A167;
  assign \new_[54919]_  = \new_[54918]_  & \new_[54915]_ ;
  assign \new_[54922]_  = A200 & ~A199;
  assign \new_[54925]_  = A232 & A203;
  assign \new_[54926]_  = \new_[54925]_  & \new_[54922]_ ;
  assign \new_[54927]_  = \new_[54926]_  & \new_[54919]_ ;
  assign \new_[54930]_  = ~A234 & A233;
  assign \new_[54933]_  = ~A265 & ~A235;
  assign \new_[54934]_  = \new_[54933]_  & \new_[54930]_ ;
  assign \new_[54937]_  = ~A268 & ~A266;
  assign \new_[54941]_  = ~A301 & ~A299;
  assign \new_[54942]_  = ~A298 & \new_[54941]_ ;
  assign \new_[54943]_  = \new_[54942]_  & \new_[54937]_ ;
  assign \new_[54944]_  = \new_[54943]_  & \new_[54934]_ ;
  assign \new_[54947]_  = ~A168 & ~A169;
  assign \new_[54950]_  = A166 & A167;
  assign \new_[54951]_  = \new_[54950]_  & \new_[54947]_ ;
  assign \new_[54954]_  = A200 & ~A199;
  assign \new_[54957]_  = ~A232 & A203;
  assign \new_[54958]_  = \new_[54957]_  & \new_[54954]_ ;
  assign \new_[54959]_  = \new_[54958]_  & \new_[54951]_ ;
  assign \new_[54962]_  = ~A235 & ~A233;
  assign \new_[54965]_  = ~A268 & ~A267;
  assign \new_[54966]_  = \new_[54965]_  & \new_[54962]_ ;
  assign \new_[54969]_  = A298 & ~A269;
  assign \new_[54973]_  = ~A301 & ~A300;
  assign \new_[54974]_  = A299 & \new_[54973]_ ;
  assign \new_[54975]_  = \new_[54974]_  & \new_[54969]_ ;
  assign \new_[54976]_  = \new_[54975]_  & \new_[54966]_ ;
  assign \new_[54979]_  = ~A168 & ~A169;
  assign \new_[54982]_  = A166 & A167;
  assign \new_[54983]_  = \new_[54982]_  & \new_[54979]_ ;
  assign \new_[54986]_  = A200 & ~A199;
  assign \new_[54989]_  = ~A232 & A203;
  assign \new_[54990]_  = \new_[54989]_  & \new_[54986]_ ;
  assign \new_[54991]_  = \new_[54990]_  & \new_[54983]_ ;
  assign \new_[54994]_  = ~A235 & ~A233;
  assign \new_[54997]_  = A266 & A265;
  assign \new_[54998]_  = \new_[54997]_  & \new_[54994]_ ;
  assign \new_[55001]_  = ~A268 & ~A267;
  assign \new_[55005]_  = ~A302 & ~A301;
  assign \new_[55006]_  = ~A300 & \new_[55005]_ ;
  assign \new_[55007]_  = \new_[55006]_  & \new_[55001]_ ;
  assign \new_[55008]_  = \new_[55007]_  & \new_[54998]_ ;
  assign \new_[55011]_  = ~A168 & ~A169;
  assign \new_[55014]_  = A166 & A167;
  assign \new_[55015]_  = \new_[55014]_  & \new_[55011]_ ;
  assign \new_[55018]_  = A200 & ~A199;
  assign \new_[55021]_  = ~A232 & A203;
  assign \new_[55022]_  = \new_[55021]_  & \new_[55018]_ ;
  assign \new_[55023]_  = \new_[55022]_  & \new_[55015]_ ;
  assign \new_[55026]_  = ~A235 & ~A233;
  assign \new_[55029]_  = A266 & A265;
  assign \new_[55030]_  = \new_[55029]_  & \new_[55026]_ ;
  assign \new_[55033]_  = ~A268 & ~A267;
  assign \new_[55037]_  = ~A301 & ~A299;
  assign \new_[55038]_  = ~A298 & \new_[55037]_ ;
  assign \new_[55039]_  = \new_[55038]_  & \new_[55033]_ ;
  assign \new_[55040]_  = \new_[55039]_  & \new_[55030]_ ;
  assign \new_[55043]_  = ~A168 & ~A169;
  assign \new_[55046]_  = A166 & A167;
  assign \new_[55047]_  = \new_[55046]_  & \new_[55043]_ ;
  assign \new_[55050]_  = A200 & ~A199;
  assign \new_[55053]_  = ~A232 & A203;
  assign \new_[55054]_  = \new_[55053]_  & \new_[55050]_ ;
  assign \new_[55055]_  = \new_[55054]_  & \new_[55047]_ ;
  assign \new_[55058]_  = ~A235 & ~A233;
  assign \new_[55061]_  = ~A266 & ~A265;
  assign \new_[55062]_  = \new_[55061]_  & \new_[55058]_ ;
  assign \new_[55065]_  = A298 & ~A268;
  assign \new_[55069]_  = ~A301 & ~A300;
  assign \new_[55070]_  = A299 & \new_[55069]_ ;
  assign \new_[55071]_  = \new_[55070]_  & \new_[55065]_ ;
  assign \new_[55072]_  = \new_[55071]_  & \new_[55062]_ ;
  assign \new_[55075]_  = ~A168 & ~A169;
  assign \new_[55078]_  = A166 & A167;
  assign \new_[55079]_  = \new_[55078]_  & \new_[55075]_ ;
  assign \new_[55082]_  = ~A200 & A199;
  assign \new_[55085]_  = ~A234 & A203;
  assign \new_[55086]_  = \new_[55085]_  & \new_[55082]_ ;
  assign \new_[55087]_  = \new_[55086]_  & \new_[55079]_ ;
  assign \new_[55090]_  = ~A236 & ~A235;
  assign \new_[55093]_  = ~A268 & ~A267;
  assign \new_[55094]_  = \new_[55093]_  & \new_[55090]_ ;
  assign \new_[55097]_  = A298 & ~A269;
  assign \new_[55101]_  = ~A301 & ~A300;
  assign \new_[55102]_  = A299 & \new_[55101]_ ;
  assign \new_[55103]_  = \new_[55102]_  & \new_[55097]_ ;
  assign \new_[55104]_  = \new_[55103]_  & \new_[55094]_ ;
  assign \new_[55107]_  = ~A168 & ~A169;
  assign \new_[55110]_  = A166 & A167;
  assign \new_[55111]_  = \new_[55110]_  & \new_[55107]_ ;
  assign \new_[55114]_  = ~A200 & A199;
  assign \new_[55117]_  = ~A234 & A203;
  assign \new_[55118]_  = \new_[55117]_  & \new_[55114]_ ;
  assign \new_[55119]_  = \new_[55118]_  & \new_[55111]_ ;
  assign \new_[55122]_  = ~A236 & ~A235;
  assign \new_[55125]_  = A266 & A265;
  assign \new_[55126]_  = \new_[55125]_  & \new_[55122]_ ;
  assign \new_[55129]_  = ~A268 & ~A267;
  assign \new_[55133]_  = ~A302 & ~A301;
  assign \new_[55134]_  = ~A300 & \new_[55133]_ ;
  assign \new_[55135]_  = \new_[55134]_  & \new_[55129]_ ;
  assign \new_[55136]_  = \new_[55135]_  & \new_[55126]_ ;
  assign \new_[55139]_  = ~A168 & ~A169;
  assign \new_[55142]_  = A166 & A167;
  assign \new_[55143]_  = \new_[55142]_  & \new_[55139]_ ;
  assign \new_[55146]_  = ~A200 & A199;
  assign \new_[55149]_  = ~A234 & A203;
  assign \new_[55150]_  = \new_[55149]_  & \new_[55146]_ ;
  assign \new_[55151]_  = \new_[55150]_  & \new_[55143]_ ;
  assign \new_[55154]_  = ~A236 & ~A235;
  assign \new_[55157]_  = A266 & A265;
  assign \new_[55158]_  = \new_[55157]_  & \new_[55154]_ ;
  assign \new_[55161]_  = ~A268 & ~A267;
  assign \new_[55165]_  = ~A301 & ~A299;
  assign \new_[55166]_  = ~A298 & \new_[55165]_ ;
  assign \new_[55167]_  = \new_[55166]_  & \new_[55161]_ ;
  assign \new_[55168]_  = \new_[55167]_  & \new_[55158]_ ;
  assign \new_[55171]_  = ~A168 & ~A169;
  assign \new_[55174]_  = A166 & A167;
  assign \new_[55175]_  = \new_[55174]_  & \new_[55171]_ ;
  assign \new_[55178]_  = ~A200 & A199;
  assign \new_[55181]_  = ~A234 & A203;
  assign \new_[55182]_  = \new_[55181]_  & \new_[55178]_ ;
  assign \new_[55183]_  = \new_[55182]_  & \new_[55175]_ ;
  assign \new_[55186]_  = ~A236 & ~A235;
  assign \new_[55189]_  = ~A266 & ~A265;
  assign \new_[55190]_  = \new_[55189]_  & \new_[55186]_ ;
  assign \new_[55193]_  = A298 & ~A268;
  assign \new_[55197]_  = ~A301 & ~A300;
  assign \new_[55198]_  = A299 & \new_[55197]_ ;
  assign \new_[55199]_  = \new_[55198]_  & \new_[55193]_ ;
  assign \new_[55200]_  = \new_[55199]_  & \new_[55190]_ ;
  assign \new_[55203]_  = ~A168 & ~A169;
  assign \new_[55206]_  = A166 & A167;
  assign \new_[55207]_  = \new_[55206]_  & \new_[55203]_ ;
  assign \new_[55210]_  = ~A200 & A199;
  assign \new_[55213]_  = A232 & A203;
  assign \new_[55214]_  = \new_[55213]_  & \new_[55210]_ ;
  assign \new_[55215]_  = \new_[55214]_  & \new_[55207]_ ;
  assign \new_[55218]_  = ~A234 & A233;
  assign \new_[55221]_  = ~A267 & ~A235;
  assign \new_[55222]_  = \new_[55221]_  & \new_[55218]_ ;
  assign \new_[55225]_  = ~A269 & ~A268;
  assign \new_[55229]_  = ~A302 & ~A301;
  assign \new_[55230]_  = ~A300 & \new_[55229]_ ;
  assign \new_[55231]_  = \new_[55230]_  & \new_[55225]_ ;
  assign \new_[55232]_  = \new_[55231]_  & \new_[55222]_ ;
  assign \new_[55235]_  = ~A168 & ~A169;
  assign \new_[55238]_  = A166 & A167;
  assign \new_[55239]_  = \new_[55238]_  & \new_[55235]_ ;
  assign \new_[55242]_  = ~A200 & A199;
  assign \new_[55245]_  = A232 & A203;
  assign \new_[55246]_  = \new_[55245]_  & \new_[55242]_ ;
  assign \new_[55247]_  = \new_[55246]_  & \new_[55239]_ ;
  assign \new_[55250]_  = ~A234 & A233;
  assign \new_[55253]_  = ~A267 & ~A235;
  assign \new_[55254]_  = \new_[55253]_  & \new_[55250]_ ;
  assign \new_[55257]_  = ~A269 & ~A268;
  assign \new_[55261]_  = ~A301 & ~A299;
  assign \new_[55262]_  = ~A298 & \new_[55261]_ ;
  assign \new_[55263]_  = \new_[55262]_  & \new_[55257]_ ;
  assign \new_[55264]_  = \new_[55263]_  & \new_[55254]_ ;
  assign \new_[55267]_  = ~A168 & ~A169;
  assign \new_[55270]_  = A166 & A167;
  assign \new_[55271]_  = \new_[55270]_  & \new_[55267]_ ;
  assign \new_[55274]_  = ~A200 & A199;
  assign \new_[55277]_  = A232 & A203;
  assign \new_[55278]_  = \new_[55277]_  & \new_[55274]_ ;
  assign \new_[55279]_  = \new_[55278]_  & \new_[55271]_ ;
  assign \new_[55282]_  = ~A234 & A233;
  assign \new_[55285]_  = ~A265 & ~A235;
  assign \new_[55286]_  = \new_[55285]_  & \new_[55282]_ ;
  assign \new_[55289]_  = ~A268 & ~A266;
  assign \new_[55293]_  = ~A302 & ~A301;
  assign \new_[55294]_  = ~A300 & \new_[55293]_ ;
  assign \new_[55295]_  = \new_[55294]_  & \new_[55289]_ ;
  assign \new_[55296]_  = \new_[55295]_  & \new_[55286]_ ;
  assign \new_[55299]_  = ~A168 & ~A169;
  assign \new_[55302]_  = A166 & A167;
  assign \new_[55303]_  = \new_[55302]_  & \new_[55299]_ ;
  assign \new_[55306]_  = ~A200 & A199;
  assign \new_[55309]_  = A232 & A203;
  assign \new_[55310]_  = \new_[55309]_  & \new_[55306]_ ;
  assign \new_[55311]_  = \new_[55310]_  & \new_[55303]_ ;
  assign \new_[55314]_  = ~A234 & A233;
  assign \new_[55317]_  = ~A265 & ~A235;
  assign \new_[55318]_  = \new_[55317]_  & \new_[55314]_ ;
  assign \new_[55321]_  = ~A268 & ~A266;
  assign \new_[55325]_  = ~A301 & ~A299;
  assign \new_[55326]_  = ~A298 & \new_[55325]_ ;
  assign \new_[55327]_  = \new_[55326]_  & \new_[55321]_ ;
  assign \new_[55328]_  = \new_[55327]_  & \new_[55318]_ ;
  assign \new_[55331]_  = ~A168 & ~A169;
  assign \new_[55334]_  = A166 & A167;
  assign \new_[55335]_  = \new_[55334]_  & \new_[55331]_ ;
  assign \new_[55338]_  = ~A200 & A199;
  assign \new_[55341]_  = ~A232 & A203;
  assign \new_[55342]_  = \new_[55341]_  & \new_[55338]_ ;
  assign \new_[55343]_  = \new_[55342]_  & \new_[55335]_ ;
  assign \new_[55346]_  = ~A235 & ~A233;
  assign \new_[55349]_  = ~A268 & ~A267;
  assign \new_[55350]_  = \new_[55349]_  & \new_[55346]_ ;
  assign \new_[55353]_  = A298 & ~A269;
  assign \new_[55357]_  = ~A301 & ~A300;
  assign \new_[55358]_  = A299 & \new_[55357]_ ;
  assign \new_[55359]_  = \new_[55358]_  & \new_[55353]_ ;
  assign \new_[55360]_  = \new_[55359]_  & \new_[55350]_ ;
  assign \new_[55363]_  = ~A168 & ~A169;
  assign \new_[55366]_  = A166 & A167;
  assign \new_[55367]_  = \new_[55366]_  & \new_[55363]_ ;
  assign \new_[55370]_  = ~A200 & A199;
  assign \new_[55373]_  = ~A232 & A203;
  assign \new_[55374]_  = \new_[55373]_  & \new_[55370]_ ;
  assign \new_[55375]_  = \new_[55374]_  & \new_[55367]_ ;
  assign \new_[55378]_  = ~A235 & ~A233;
  assign \new_[55381]_  = A266 & A265;
  assign \new_[55382]_  = \new_[55381]_  & \new_[55378]_ ;
  assign \new_[55385]_  = ~A268 & ~A267;
  assign \new_[55389]_  = ~A302 & ~A301;
  assign \new_[55390]_  = ~A300 & \new_[55389]_ ;
  assign \new_[55391]_  = \new_[55390]_  & \new_[55385]_ ;
  assign \new_[55392]_  = \new_[55391]_  & \new_[55382]_ ;
  assign \new_[55395]_  = ~A168 & ~A169;
  assign \new_[55398]_  = A166 & A167;
  assign \new_[55399]_  = \new_[55398]_  & \new_[55395]_ ;
  assign \new_[55402]_  = ~A200 & A199;
  assign \new_[55405]_  = ~A232 & A203;
  assign \new_[55406]_  = \new_[55405]_  & \new_[55402]_ ;
  assign \new_[55407]_  = \new_[55406]_  & \new_[55399]_ ;
  assign \new_[55410]_  = ~A235 & ~A233;
  assign \new_[55413]_  = A266 & A265;
  assign \new_[55414]_  = \new_[55413]_  & \new_[55410]_ ;
  assign \new_[55417]_  = ~A268 & ~A267;
  assign \new_[55421]_  = ~A301 & ~A299;
  assign \new_[55422]_  = ~A298 & \new_[55421]_ ;
  assign \new_[55423]_  = \new_[55422]_  & \new_[55417]_ ;
  assign \new_[55424]_  = \new_[55423]_  & \new_[55414]_ ;
  assign \new_[55427]_  = ~A168 & ~A169;
  assign \new_[55430]_  = A166 & A167;
  assign \new_[55431]_  = \new_[55430]_  & \new_[55427]_ ;
  assign \new_[55434]_  = ~A200 & A199;
  assign \new_[55437]_  = ~A232 & A203;
  assign \new_[55438]_  = \new_[55437]_  & \new_[55434]_ ;
  assign \new_[55439]_  = \new_[55438]_  & \new_[55431]_ ;
  assign \new_[55442]_  = ~A235 & ~A233;
  assign \new_[55445]_  = ~A266 & ~A265;
  assign \new_[55446]_  = \new_[55445]_  & \new_[55442]_ ;
  assign \new_[55449]_  = A298 & ~A268;
  assign \new_[55453]_  = ~A301 & ~A300;
  assign \new_[55454]_  = A299 & \new_[55453]_ ;
  assign \new_[55455]_  = \new_[55454]_  & \new_[55449]_ ;
  assign \new_[55456]_  = \new_[55455]_  & \new_[55446]_ ;
  assign \new_[55459]_  = ~A169 & ~A170;
  assign \new_[55462]_  = A199 & ~A168;
  assign \new_[55463]_  = \new_[55462]_  & \new_[55459]_ ;
  assign \new_[55466]_  = A232 & A201;
  assign \new_[55469]_  = ~A234 & A233;
  assign \new_[55470]_  = \new_[55469]_  & \new_[55466]_ ;
  assign \new_[55471]_  = \new_[55470]_  & \new_[55463]_ ;
  assign \new_[55474]_  = A265 & ~A235;
  assign \new_[55477]_  = ~A267 & A266;
  assign \new_[55478]_  = \new_[55477]_  & \new_[55474]_ ;
  assign \new_[55481]_  = A298 & ~A268;
  assign \new_[55485]_  = ~A301 & ~A300;
  assign \new_[55486]_  = A299 & \new_[55485]_ ;
  assign \new_[55487]_  = \new_[55486]_  & \new_[55481]_ ;
  assign \new_[55488]_  = \new_[55487]_  & \new_[55478]_ ;
  assign \new_[55491]_  = ~A169 & ~A170;
  assign \new_[55494]_  = A200 & ~A168;
  assign \new_[55495]_  = \new_[55494]_  & \new_[55491]_ ;
  assign \new_[55498]_  = A232 & A201;
  assign \new_[55501]_  = ~A234 & A233;
  assign \new_[55502]_  = \new_[55501]_  & \new_[55498]_ ;
  assign \new_[55503]_  = \new_[55502]_  & \new_[55495]_ ;
  assign \new_[55506]_  = A265 & ~A235;
  assign \new_[55509]_  = ~A267 & A266;
  assign \new_[55510]_  = \new_[55509]_  & \new_[55506]_ ;
  assign \new_[55513]_  = A298 & ~A268;
  assign \new_[55517]_  = ~A301 & ~A300;
  assign \new_[55518]_  = A299 & \new_[55517]_ ;
  assign \new_[55519]_  = \new_[55518]_  & \new_[55513]_ ;
  assign \new_[55520]_  = \new_[55519]_  & \new_[55510]_ ;
  assign \new_[55523]_  = ~A169 & ~A170;
  assign \new_[55526]_  = ~A199 & ~A168;
  assign \new_[55527]_  = \new_[55526]_  & \new_[55523]_ ;
  assign \new_[55530]_  = A203 & A200;
  assign \new_[55533]_  = ~A235 & ~A234;
  assign \new_[55534]_  = \new_[55533]_  & \new_[55530]_ ;
  assign \new_[55535]_  = \new_[55534]_  & \new_[55527]_ ;
  assign \new_[55538]_  = A265 & ~A236;
  assign \new_[55541]_  = ~A267 & A266;
  assign \new_[55542]_  = \new_[55541]_  & \new_[55538]_ ;
  assign \new_[55545]_  = A298 & ~A268;
  assign \new_[55549]_  = ~A301 & ~A300;
  assign \new_[55550]_  = A299 & \new_[55549]_ ;
  assign \new_[55551]_  = \new_[55550]_  & \new_[55545]_ ;
  assign \new_[55552]_  = \new_[55551]_  & \new_[55542]_ ;
  assign \new_[55555]_  = ~A169 & ~A170;
  assign \new_[55558]_  = ~A199 & ~A168;
  assign \new_[55559]_  = \new_[55558]_  & \new_[55555]_ ;
  assign \new_[55562]_  = A203 & A200;
  assign \new_[55565]_  = A233 & A232;
  assign \new_[55566]_  = \new_[55565]_  & \new_[55562]_ ;
  assign \new_[55567]_  = \new_[55566]_  & \new_[55559]_ ;
  assign \new_[55570]_  = ~A235 & ~A234;
  assign \new_[55573]_  = ~A268 & ~A267;
  assign \new_[55574]_  = \new_[55573]_  & \new_[55570]_ ;
  assign \new_[55577]_  = A298 & ~A269;
  assign \new_[55581]_  = ~A301 & ~A300;
  assign \new_[55582]_  = A299 & \new_[55581]_ ;
  assign \new_[55583]_  = \new_[55582]_  & \new_[55577]_ ;
  assign \new_[55584]_  = \new_[55583]_  & \new_[55574]_ ;
  assign \new_[55587]_  = ~A169 & ~A170;
  assign \new_[55590]_  = ~A199 & ~A168;
  assign \new_[55591]_  = \new_[55590]_  & \new_[55587]_ ;
  assign \new_[55594]_  = A203 & A200;
  assign \new_[55597]_  = A233 & A232;
  assign \new_[55598]_  = \new_[55597]_  & \new_[55594]_ ;
  assign \new_[55599]_  = \new_[55598]_  & \new_[55591]_ ;
  assign \new_[55602]_  = ~A235 & ~A234;
  assign \new_[55605]_  = A266 & A265;
  assign \new_[55606]_  = \new_[55605]_  & \new_[55602]_ ;
  assign \new_[55609]_  = ~A268 & ~A267;
  assign \new_[55613]_  = ~A302 & ~A301;
  assign \new_[55614]_  = ~A300 & \new_[55613]_ ;
  assign \new_[55615]_  = \new_[55614]_  & \new_[55609]_ ;
  assign \new_[55616]_  = \new_[55615]_  & \new_[55606]_ ;
  assign \new_[55619]_  = ~A169 & ~A170;
  assign \new_[55622]_  = ~A199 & ~A168;
  assign \new_[55623]_  = \new_[55622]_  & \new_[55619]_ ;
  assign \new_[55626]_  = A203 & A200;
  assign \new_[55629]_  = A233 & A232;
  assign \new_[55630]_  = \new_[55629]_  & \new_[55626]_ ;
  assign \new_[55631]_  = \new_[55630]_  & \new_[55623]_ ;
  assign \new_[55634]_  = ~A235 & ~A234;
  assign \new_[55637]_  = A266 & A265;
  assign \new_[55638]_  = \new_[55637]_  & \new_[55634]_ ;
  assign \new_[55641]_  = ~A268 & ~A267;
  assign \new_[55645]_  = ~A301 & ~A299;
  assign \new_[55646]_  = ~A298 & \new_[55645]_ ;
  assign \new_[55647]_  = \new_[55646]_  & \new_[55641]_ ;
  assign \new_[55648]_  = \new_[55647]_  & \new_[55638]_ ;
  assign \new_[55651]_  = ~A169 & ~A170;
  assign \new_[55654]_  = ~A199 & ~A168;
  assign \new_[55655]_  = \new_[55654]_  & \new_[55651]_ ;
  assign \new_[55658]_  = A203 & A200;
  assign \new_[55661]_  = A233 & A232;
  assign \new_[55662]_  = \new_[55661]_  & \new_[55658]_ ;
  assign \new_[55663]_  = \new_[55662]_  & \new_[55655]_ ;
  assign \new_[55666]_  = ~A235 & ~A234;
  assign \new_[55669]_  = ~A266 & ~A265;
  assign \new_[55670]_  = \new_[55669]_  & \new_[55666]_ ;
  assign \new_[55673]_  = A298 & ~A268;
  assign \new_[55677]_  = ~A301 & ~A300;
  assign \new_[55678]_  = A299 & \new_[55677]_ ;
  assign \new_[55679]_  = \new_[55678]_  & \new_[55673]_ ;
  assign \new_[55680]_  = \new_[55679]_  & \new_[55670]_ ;
  assign \new_[55683]_  = ~A169 & ~A170;
  assign \new_[55686]_  = ~A199 & ~A168;
  assign \new_[55687]_  = \new_[55686]_  & \new_[55683]_ ;
  assign \new_[55690]_  = A203 & A200;
  assign \new_[55693]_  = ~A233 & ~A232;
  assign \new_[55694]_  = \new_[55693]_  & \new_[55690]_ ;
  assign \new_[55695]_  = \new_[55694]_  & \new_[55687]_ ;
  assign \new_[55698]_  = A265 & ~A235;
  assign \new_[55701]_  = ~A267 & A266;
  assign \new_[55702]_  = \new_[55701]_  & \new_[55698]_ ;
  assign \new_[55705]_  = A298 & ~A268;
  assign \new_[55709]_  = ~A301 & ~A300;
  assign \new_[55710]_  = A299 & \new_[55709]_ ;
  assign \new_[55711]_  = \new_[55710]_  & \new_[55705]_ ;
  assign \new_[55712]_  = \new_[55711]_  & \new_[55702]_ ;
  assign \new_[55715]_  = ~A169 & ~A170;
  assign \new_[55718]_  = A199 & ~A168;
  assign \new_[55719]_  = \new_[55718]_  & \new_[55715]_ ;
  assign \new_[55722]_  = A203 & ~A200;
  assign \new_[55725]_  = ~A235 & ~A234;
  assign \new_[55726]_  = \new_[55725]_  & \new_[55722]_ ;
  assign \new_[55727]_  = \new_[55726]_  & \new_[55719]_ ;
  assign \new_[55730]_  = A265 & ~A236;
  assign \new_[55733]_  = ~A267 & A266;
  assign \new_[55734]_  = \new_[55733]_  & \new_[55730]_ ;
  assign \new_[55737]_  = A298 & ~A268;
  assign \new_[55741]_  = ~A301 & ~A300;
  assign \new_[55742]_  = A299 & \new_[55741]_ ;
  assign \new_[55743]_  = \new_[55742]_  & \new_[55737]_ ;
  assign \new_[55744]_  = \new_[55743]_  & \new_[55734]_ ;
  assign \new_[55747]_  = ~A169 & ~A170;
  assign \new_[55750]_  = A199 & ~A168;
  assign \new_[55751]_  = \new_[55750]_  & \new_[55747]_ ;
  assign \new_[55754]_  = A203 & ~A200;
  assign \new_[55757]_  = A233 & A232;
  assign \new_[55758]_  = \new_[55757]_  & \new_[55754]_ ;
  assign \new_[55759]_  = \new_[55758]_  & \new_[55751]_ ;
  assign \new_[55762]_  = ~A235 & ~A234;
  assign \new_[55765]_  = ~A268 & ~A267;
  assign \new_[55766]_  = \new_[55765]_  & \new_[55762]_ ;
  assign \new_[55769]_  = A298 & ~A269;
  assign \new_[55773]_  = ~A301 & ~A300;
  assign \new_[55774]_  = A299 & \new_[55773]_ ;
  assign \new_[55775]_  = \new_[55774]_  & \new_[55769]_ ;
  assign \new_[55776]_  = \new_[55775]_  & \new_[55766]_ ;
  assign \new_[55779]_  = ~A169 & ~A170;
  assign \new_[55782]_  = A199 & ~A168;
  assign \new_[55783]_  = \new_[55782]_  & \new_[55779]_ ;
  assign \new_[55786]_  = A203 & ~A200;
  assign \new_[55789]_  = A233 & A232;
  assign \new_[55790]_  = \new_[55789]_  & \new_[55786]_ ;
  assign \new_[55791]_  = \new_[55790]_  & \new_[55783]_ ;
  assign \new_[55794]_  = ~A235 & ~A234;
  assign \new_[55797]_  = A266 & A265;
  assign \new_[55798]_  = \new_[55797]_  & \new_[55794]_ ;
  assign \new_[55801]_  = ~A268 & ~A267;
  assign \new_[55805]_  = ~A302 & ~A301;
  assign \new_[55806]_  = ~A300 & \new_[55805]_ ;
  assign \new_[55807]_  = \new_[55806]_  & \new_[55801]_ ;
  assign \new_[55808]_  = \new_[55807]_  & \new_[55798]_ ;
  assign \new_[55811]_  = ~A169 & ~A170;
  assign \new_[55814]_  = A199 & ~A168;
  assign \new_[55815]_  = \new_[55814]_  & \new_[55811]_ ;
  assign \new_[55818]_  = A203 & ~A200;
  assign \new_[55821]_  = A233 & A232;
  assign \new_[55822]_  = \new_[55821]_  & \new_[55818]_ ;
  assign \new_[55823]_  = \new_[55822]_  & \new_[55815]_ ;
  assign \new_[55826]_  = ~A235 & ~A234;
  assign \new_[55829]_  = A266 & A265;
  assign \new_[55830]_  = \new_[55829]_  & \new_[55826]_ ;
  assign \new_[55833]_  = ~A268 & ~A267;
  assign \new_[55837]_  = ~A301 & ~A299;
  assign \new_[55838]_  = ~A298 & \new_[55837]_ ;
  assign \new_[55839]_  = \new_[55838]_  & \new_[55833]_ ;
  assign \new_[55840]_  = \new_[55839]_  & \new_[55830]_ ;
  assign \new_[55843]_  = ~A169 & ~A170;
  assign \new_[55846]_  = A199 & ~A168;
  assign \new_[55847]_  = \new_[55846]_  & \new_[55843]_ ;
  assign \new_[55850]_  = A203 & ~A200;
  assign \new_[55853]_  = A233 & A232;
  assign \new_[55854]_  = \new_[55853]_  & \new_[55850]_ ;
  assign \new_[55855]_  = \new_[55854]_  & \new_[55847]_ ;
  assign \new_[55858]_  = ~A235 & ~A234;
  assign \new_[55861]_  = ~A266 & ~A265;
  assign \new_[55862]_  = \new_[55861]_  & \new_[55858]_ ;
  assign \new_[55865]_  = A298 & ~A268;
  assign \new_[55869]_  = ~A301 & ~A300;
  assign \new_[55870]_  = A299 & \new_[55869]_ ;
  assign \new_[55871]_  = \new_[55870]_  & \new_[55865]_ ;
  assign \new_[55872]_  = \new_[55871]_  & \new_[55862]_ ;
  assign \new_[55875]_  = ~A169 & ~A170;
  assign \new_[55878]_  = A199 & ~A168;
  assign \new_[55879]_  = \new_[55878]_  & \new_[55875]_ ;
  assign \new_[55882]_  = A203 & ~A200;
  assign \new_[55885]_  = ~A233 & ~A232;
  assign \new_[55886]_  = \new_[55885]_  & \new_[55882]_ ;
  assign \new_[55887]_  = \new_[55886]_  & \new_[55879]_ ;
  assign \new_[55890]_  = A265 & ~A235;
  assign \new_[55893]_  = ~A267 & A266;
  assign \new_[55894]_  = \new_[55893]_  & \new_[55890]_ ;
  assign \new_[55897]_  = A298 & ~A268;
  assign \new_[55901]_  = ~A301 & ~A300;
  assign \new_[55902]_  = A299 & \new_[55901]_ ;
  assign \new_[55903]_  = \new_[55902]_  & \new_[55897]_ ;
  assign \new_[55904]_  = \new_[55903]_  & \new_[55894]_ ;
  assign \new_[55907]_  = A166 & A168;
  assign \new_[55910]_  = A200 & A199;
  assign \new_[55911]_  = \new_[55910]_  & \new_[55907]_ ;
  assign \new_[55914]_  = ~A202 & ~A201;
  assign \new_[55918]_  = ~A234 & A233;
  assign \new_[55919]_  = A232 & \new_[55918]_ ;
  assign \new_[55920]_  = \new_[55919]_  & \new_[55914]_ ;
  assign \new_[55921]_  = \new_[55920]_  & \new_[55911]_ ;
  assign \new_[55924]_  = A265 & ~A235;
  assign \new_[55927]_  = ~A267 & A266;
  assign \new_[55928]_  = \new_[55927]_  & \new_[55924]_ ;
  assign \new_[55931]_  = A298 & ~A268;
  assign \new_[55935]_  = ~A301 & ~A300;
  assign \new_[55936]_  = A299 & \new_[55935]_ ;
  assign \new_[55937]_  = \new_[55936]_  & \new_[55931]_ ;
  assign \new_[55938]_  = \new_[55937]_  & \new_[55928]_ ;
  assign \new_[55941]_  = A167 & A168;
  assign \new_[55944]_  = A200 & A199;
  assign \new_[55945]_  = \new_[55944]_  & \new_[55941]_ ;
  assign \new_[55948]_  = ~A202 & ~A201;
  assign \new_[55952]_  = ~A234 & A233;
  assign \new_[55953]_  = A232 & \new_[55952]_ ;
  assign \new_[55954]_  = \new_[55953]_  & \new_[55948]_ ;
  assign \new_[55955]_  = \new_[55954]_  & \new_[55945]_ ;
  assign \new_[55958]_  = A265 & ~A235;
  assign \new_[55961]_  = ~A267 & A266;
  assign \new_[55962]_  = \new_[55961]_  & \new_[55958]_ ;
  assign \new_[55965]_  = A298 & ~A268;
  assign \new_[55969]_  = ~A301 & ~A300;
  assign \new_[55970]_  = A299 & \new_[55969]_ ;
  assign \new_[55971]_  = \new_[55970]_  & \new_[55965]_ ;
  assign \new_[55972]_  = \new_[55971]_  & \new_[55962]_ ;
  assign \new_[55975]_  = A167 & A170;
  assign \new_[55978]_  = ~A201 & ~A166;
  assign \new_[55979]_  = \new_[55978]_  & \new_[55975]_ ;
  assign \new_[55982]_  = ~A203 & ~A202;
  assign \new_[55986]_  = ~A234 & A233;
  assign \new_[55987]_  = A232 & \new_[55986]_ ;
  assign \new_[55988]_  = \new_[55987]_  & \new_[55982]_ ;
  assign \new_[55989]_  = \new_[55988]_  & \new_[55979]_ ;
  assign \new_[55992]_  = A265 & ~A235;
  assign \new_[55995]_  = ~A267 & A266;
  assign \new_[55996]_  = \new_[55995]_  & \new_[55992]_ ;
  assign \new_[55999]_  = A298 & ~A268;
  assign \new_[56003]_  = ~A301 & ~A300;
  assign \new_[56004]_  = A299 & \new_[56003]_ ;
  assign \new_[56005]_  = \new_[56004]_  & \new_[55999]_ ;
  assign \new_[56006]_  = \new_[56005]_  & \new_[55996]_ ;
  assign \new_[56009]_  = A167 & A170;
  assign \new_[56012]_  = A199 & ~A166;
  assign \new_[56013]_  = \new_[56012]_  & \new_[56009]_ ;
  assign \new_[56016]_  = ~A201 & A200;
  assign \new_[56020]_  = ~A235 & ~A234;
  assign \new_[56021]_  = ~A202 & \new_[56020]_ ;
  assign \new_[56022]_  = \new_[56021]_  & \new_[56016]_ ;
  assign \new_[56023]_  = \new_[56022]_  & \new_[56013]_ ;
  assign \new_[56026]_  = A265 & ~A236;
  assign \new_[56029]_  = ~A267 & A266;
  assign \new_[56030]_  = \new_[56029]_  & \new_[56026]_ ;
  assign \new_[56033]_  = A298 & ~A268;
  assign \new_[56037]_  = ~A301 & ~A300;
  assign \new_[56038]_  = A299 & \new_[56037]_ ;
  assign \new_[56039]_  = \new_[56038]_  & \new_[56033]_ ;
  assign \new_[56040]_  = \new_[56039]_  & \new_[56030]_ ;
  assign \new_[56043]_  = A167 & A170;
  assign \new_[56046]_  = A199 & ~A166;
  assign \new_[56047]_  = \new_[56046]_  & \new_[56043]_ ;
  assign \new_[56050]_  = ~A201 & A200;
  assign \new_[56054]_  = A233 & A232;
  assign \new_[56055]_  = ~A202 & \new_[56054]_ ;
  assign \new_[56056]_  = \new_[56055]_  & \new_[56050]_ ;
  assign \new_[56057]_  = \new_[56056]_  & \new_[56047]_ ;
  assign \new_[56060]_  = ~A235 & ~A234;
  assign \new_[56063]_  = ~A268 & ~A267;
  assign \new_[56064]_  = \new_[56063]_  & \new_[56060]_ ;
  assign \new_[56067]_  = A298 & ~A269;
  assign \new_[56071]_  = ~A301 & ~A300;
  assign \new_[56072]_  = A299 & \new_[56071]_ ;
  assign \new_[56073]_  = \new_[56072]_  & \new_[56067]_ ;
  assign \new_[56074]_  = \new_[56073]_  & \new_[56064]_ ;
  assign \new_[56077]_  = A167 & A170;
  assign \new_[56080]_  = A199 & ~A166;
  assign \new_[56081]_  = \new_[56080]_  & \new_[56077]_ ;
  assign \new_[56084]_  = ~A201 & A200;
  assign \new_[56088]_  = A233 & A232;
  assign \new_[56089]_  = ~A202 & \new_[56088]_ ;
  assign \new_[56090]_  = \new_[56089]_  & \new_[56084]_ ;
  assign \new_[56091]_  = \new_[56090]_  & \new_[56081]_ ;
  assign \new_[56094]_  = ~A235 & ~A234;
  assign \new_[56097]_  = A266 & A265;
  assign \new_[56098]_  = \new_[56097]_  & \new_[56094]_ ;
  assign \new_[56101]_  = ~A268 & ~A267;
  assign \new_[56105]_  = ~A302 & ~A301;
  assign \new_[56106]_  = ~A300 & \new_[56105]_ ;
  assign \new_[56107]_  = \new_[56106]_  & \new_[56101]_ ;
  assign \new_[56108]_  = \new_[56107]_  & \new_[56098]_ ;
  assign \new_[56111]_  = A167 & A170;
  assign \new_[56114]_  = A199 & ~A166;
  assign \new_[56115]_  = \new_[56114]_  & \new_[56111]_ ;
  assign \new_[56118]_  = ~A201 & A200;
  assign \new_[56122]_  = A233 & A232;
  assign \new_[56123]_  = ~A202 & \new_[56122]_ ;
  assign \new_[56124]_  = \new_[56123]_  & \new_[56118]_ ;
  assign \new_[56125]_  = \new_[56124]_  & \new_[56115]_ ;
  assign \new_[56128]_  = ~A235 & ~A234;
  assign \new_[56131]_  = A266 & A265;
  assign \new_[56132]_  = \new_[56131]_  & \new_[56128]_ ;
  assign \new_[56135]_  = ~A268 & ~A267;
  assign \new_[56139]_  = ~A301 & ~A299;
  assign \new_[56140]_  = ~A298 & \new_[56139]_ ;
  assign \new_[56141]_  = \new_[56140]_  & \new_[56135]_ ;
  assign \new_[56142]_  = \new_[56141]_  & \new_[56132]_ ;
  assign \new_[56145]_  = A167 & A170;
  assign \new_[56148]_  = A199 & ~A166;
  assign \new_[56149]_  = \new_[56148]_  & \new_[56145]_ ;
  assign \new_[56152]_  = ~A201 & A200;
  assign \new_[56156]_  = A233 & A232;
  assign \new_[56157]_  = ~A202 & \new_[56156]_ ;
  assign \new_[56158]_  = \new_[56157]_  & \new_[56152]_ ;
  assign \new_[56159]_  = \new_[56158]_  & \new_[56149]_ ;
  assign \new_[56162]_  = ~A235 & ~A234;
  assign \new_[56165]_  = ~A266 & ~A265;
  assign \new_[56166]_  = \new_[56165]_  & \new_[56162]_ ;
  assign \new_[56169]_  = A298 & ~A268;
  assign \new_[56173]_  = ~A301 & ~A300;
  assign \new_[56174]_  = A299 & \new_[56173]_ ;
  assign \new_[56175]_  = \new_[56174]_  & \new_[56169]_ ;
  assign \new_[56176]_  = \new_[56175]_  & \new_[56166]_ ;
  assign \new_[56179]_  = A167 & A170;
  assign \new_[56182]_  = A199 & ~A166;
  assign \new_[56183]_  = \new_[56182]_  & \new_[56179]_ ;
  assign \new_[56186]_  = ~A201 & A200;
  assign \new_[56190]_  = ~A233 & ~A232;
  assign \new_[56191]_  = ~A202 & \new_[56190]_ ;
  assign \new_[56192]_  = \new_[56191]_  & \new_[56186]_ ;
  assign \new_[56193]_  = \new_[56192]_  & \new_[56183]_ ;
  assign \new_[56196]_  = A265 & ~A235;
  assign \new_[56199]_  = ~A267 & A266;
  assign \new_[56200]_  = \new_[56199]_  & \new_[56196]_ ;
  assign \new_[56203]_  = A298 & ~A268;
  assign \new_[56207]_  = ~A301 & ~A300;
  assign \new_[56208]_  = A299 & \new_[56207]_ ;
  assign \new_[56209]_  = \new_[56208]_  & \new_[56203]_ ;
  assign \new_[56210]_  = \new_[56209]_  & \new_[56200]_ ;
  assign \new_[56213]_  = A167 & A170;
  assign \new_[56216]_  = ~A199 & ~A166;
  assign \new_[56217]_  = \new_[56216]_  & \new_[56213]_ ;
  assign \new_[56220]_  = ~A202 & ~A200;
  assign \new_[56224]_  = ~A234 & A233;
  assign \new_[56225]_  = A232 & \new_[56224]_ ;
  assign \new_[56226]_  = \new_[56225]_  & \new_[56220]_ ;
  assign \new_[56227]_  = \new_[56226]_  & \new_[56217]_ ;
  assign \new_[56230]_  = A265 & ~A235;
  assign \new_[56233]_  = ~A267 & A266;
  assign \new_[56234]_  = \new_[56233]_  & \new_[56230]_ ;
  assign \new_[56237]_  = A298 & ~A268;
  assign \new_[56241]_  = ~A301 & ~A300;
  assign \new_[56242]_  = A299 & \new_[56241]_ ;
  assign \new_[56243]_  = \new_[56242]_  & \new_[56237]_ ;
  assign \new_[56244]_  = \new_[56243]_  & \new_[56234]_ ;
  assign \new_[56247]_  = ~A167 & A170;
  assign \new_[56250]_  = ~A201 & A166;
  assign \new_[56251]_  = \new_[56250]_  & \new_[56247]_ ;
  assign \new_[56254]_  = ~A203 & ~A202;
  assign \new_[56258]_  = ~A234 & A233;
  assign \new_[56259]_  = A232 & \new_[56258]_ ;
  assign \new_[56260]_  = \new_[56259]_  & \new_[56254]_ ;
  assign \new_[56261]_  = \new_[56260]_  & \new_[56251]_ ;
  assign \new_[56264]_  = A265 & ~A235;
  assign \new_[56267]_  = ~A267 & A266;
  assign \new_[56268]_  = \new_[56267]_  & \new_[56264]_ ;
  assign \new_[56271]_  = A298 & ~A268;
  assign \new_[56275]_  = ~A301 & ~A300;
  assign \new_[56276]_  = A299 & \new_[56275]_ ;
  assign \new_[56277]_  = \new_[56276]_  & \new_[56271]_ ;
  assign \new_[56278]_  = \new_[56277]_  & \new_[56268]_ ;
  assign \new_[56281]_  = ~A167 & A170;
  assign \new_[56284]_  = A199 & A166;
  assign \new_[56285]_  = \new_[56284]_  & \new_[56281]_ ;
  assign \new_[56288]_  = ~A201 & A200;
  assign \new_[56292]_  = ~A235 & ~A234;
  assign \new_[56293]_  = ~A202 & \new_[56292]_ ;
  assign \new_[56294]_  = \new_[56293]_  & \new_[56288]_ ;
  assign \new_[56295]_  = \new_[56294]_  & \new_[56285]_ ;
  assign \new_[56298]_  = A265 & ~A236;
  assign \new_[56301]_  = ~A267 & A266;
  assign \new_[56302]_  = \new_[56301]_  & \new_[56298]_ ;
  assign \new_[56305]_  = A298 & ~A268;
  assign \new_[56309]_  = ~A301 & ~A300;
  assign \new_[56310]_  = A299 & \new_[56309]_ ;
  assign \new_[56311]_  = \new_[56310]_  & \new_[56305]_ ;
  assign \new_[56312]_  = \new_[56311]_  & \new_[56302]_ ;
  assign \new_[56315]_  = ~A167 & A170;
  assign \new_[56318]_  = A199 & A166;
  assign \new_[56319]_  = \new_[56318]_  & \new_[56315]_ ;
  assign \new_[56322]_  = ~A201 & A200;
  assign \new_[56326]_  = A233 & A232;
  assign \new_[56327]_  = ~A202 & \new_[56326]_ ;
  assign \new_[56328]_  = \new_[56327]_  & \new_[56322]_ ;
  assign \new_[56329]_  = \new_[56328]_  & \new_[56319]_ ;
  assign \new_[56332]_  = ~A235 & ~A234;
  assign \new_[56335]_  = ~A268 & ~A267;
  assign \new_[56336]_  = \new_[56335]_  & \new_[56332]_ ;
  assign \new_[56339]_  = A298 & ~A269;
  assign \new_[56343]_  = ~A301 & ~A300;
  assign \new_[56344]_  = A299 & \new_[56343]_ ;
  assign \new_[56345]_  = \new_[56344]_  & \new_[56339]_ ;
  assign \new_[56346]_  = \new_[56345]_  & \new_[56336]_ ;
  assign \new_[56349]_  = ~A167 & A170;
  assign \new_[56352]_  = A199 & A166;
  assign \new_[56353]_  = \new_[56352]_  & \new_[56349]_ ;
  assign \new_[56356]_  = ~A201 & A200;
  assign \new_[56360]_  = A233 & A232;
  assign \new_[56361]_  = ~A202 & \new_[56360]_ ;
  assign \new_[56362]_  = \new_[56361]_  & \new_[56356]_ ;
  assign \new_[56363]_  = \new_[56362]_  & \new_[56353]_ ;
  assign \new_[56366]_  = ~A235 & ~A234;
  assign \new_[56369]_  = A266 & A265;
  assign \new_[56370]_  = \new_[56369]_  & \new_[56366]_ ;
  assign \new_[56373]_  = ~A268 & ~A267;
  assign \new_[56377]_  = ~A302 & ~A301;
  assign \new_[56378]_  = ~A300 & \new_[56377]_ ;
  assign \new_[56379]_  = \new_[56378]_  & \new_[56373]_ ;
  assign \new_[56380]_  = \new_[56379]_  & \new_[56370]_ ;
  assign \new_[56383]_  = ~A167 & A170;
  assign \new_[56386]_  = A199 & A166;
  assign \new_[56387]_  = \new_[56386]_  & \new_[56383]_ ;
  assign \new_[56390]_  = ~A201 & A200;
  assign \new_[56394]_  = A233 & A232;
  assign \new_[56395]_  = ~A202 & \new_[56394]_ ;
  assign \new_[56396]_  = \new_[56395]_  & \new_[56390]_ ;
  assign \new_[56397]_  = \new_[56396]_  & \new_[56387]_ ;
  assign \new_[56400]_  = ~A235 & ~A234;
  assign \new_[56403]_  = A266 & A265;
  assign \new_[56404]_  = \new_[56403]_  & \new_[56400]_ ;
  assign \new_[56407]_  = ~A268 & ~A267;
  assign \new_[56411]_  = ~A301 & ~A299;
  assign \new_[56412]_  = ~A298 & \new_[56411]_ ;
  assign \new_[56413]_  = \new_[56412]_  & \new_[56407]_ ;
  assign \new_[56414]_  = \new_[56413]_  & \new_[56404]_ ;
  assign \new_[56417]_  = ~A167 & A170;
  assign \new_[56420]_  = A199 & A166;
  assign \new_[56421]_  = \new_[56420]_  & \new_[56417]_ ;
  assign \new_[56424]_  = ~A201 & A200;
  assign \new_[56428]_  = A233 & A232;
  assign \new_[56429]_  = ~A202 & \new_[56428]_ ;
  assign \new_[56430]_  = \new_[56429]_  & \new_[56424]_ ;
  assign \new_[56431]_  = \new_[56430]_  & \new_[56421]_ ;
  assign \new_[56434]_  = ~A235 & ~A234;
  assign \new_[56437]_  = ~A266 & ~A265;
  assign \new_[56438]_  = \new_[56437]_  & \new_[56434]_ ;
  assign \new_[56441]_  = A298 & ~A268;
  assign \new_[56445]_  = ~A301 & ~A300;
  assign \new_[56446]_  = A299 & \new_[56445]_ ;
  assign \new_[56447]_  = \new_[56446]_  & \new_[56441]_ ;
  assign \new_[56448]_  = \new_[56447]_  & \new_[56438]_ ;
  assign \new_[56451]_  = ~A167 & A170;
  assign \new_[56454]_  = A199 & A166;
  assign \new_[56455]_  = \new_[56454]_  & \new_[56451]_ ;
  assign \new_[56458]_  = ~A201 & A200;
  assign \new_[56462]_  = ~A233 & ~A232;
  assign \new_[56463]_  = ~A202 & \new_[56462]_ ;
  assign \new_[56464]_  = \new_[56463]_  & \new_[56458]_ ;
  assign \new_[56465]_  = \new_[56464]_  & \new_[56455]_ ;
  assign \new_[56468]_  = A265 & ~A235;
  assign \new_[56471]_  = ~A267 & A266;
  assign \new_[56472]_  = \new_[56471]_  & \new_[56468]_ ;
  assign \new_[56475]_  = A298 & ~A268;
  assign \new_[56479]_  = ~A301 & ~A300;
  assign \new_[56480]_  = A299 & \new_[56479]_ ;
  assign \new_[56481]_  = \new_[56480]_  & \new_[56475]_ ;
  assign \new_[56482]_  = \new_[56481]_  & \new_[56472]_ ;
  assign \new_[56485]_  = ~A167 & A170;
  assign \new_[56488]_  = ~A199 & A166;
  assign \new_[56489]_  = \new_[56488]_  & \new_[56485]_ ;
  assign \new_[56492]_  = ~A202 & ~A200;
  assign \new_[56496]_  = ~A234 & A233;
  assign \new_[56497]_  = A232 & \new_[56496]_ ;
  assign \new_[56498]_  = \new_[56497]_  & \new_[56492]_ ;
  assign \new_[56499]_  = \new_[56498]_  & \new_[56489]_ ;
  assign \new_[56502]_  = A265 & ~A235;
  assign \new_[56505]_  = ~A267 & A266;
  assign \new_[56506]_  = \new_[56505]_  & \new_[56502]_ ;
  assign \new_[56509]_  = A298 & ~A268;
  assign \new_[56513]_  = ~A301 & ~A300;
  assign \new_[56514]_  = A299 & \new_[56513]_ ;
  assign \new_[56515]_  = \new_[56514]_  & \new_[56509]_ ;
  assign \new_[56516]_  = \new_[56515]_  & \new_[56506]_ ;
  assign \new_[56519]_  = ~A167 & ~A169;
  assign \new_[56522]_  = ~A199 & ~A166;
  assign \new_[56523]_  = \new_[56522]_  & \new_[56519]_ ;
  assign \new_[56526]_  = A203 & A200;
  assign \new_[56530]_  = ~A234 & A233;
  assign \new_[56531]_  = A232 & \new_[56530]_ ;
  assign \new_[56532]_  = \new_[56531]_  & \new_[56526]_ ;
  assign \new_[56533]_  = \new_[56532]_  & \new_[56523]_ ;
  assign \new_[56536]_  = A265 & ~A235;
  assign \new_[56539]_  = ~A267 & A266;
  assign \new_[56540]_  = \new_[56539]_  & \new_[56536]_ ;
  assign \new_[56543]_  = A298 & ~A268;
  assign \new_[56547]_  = ~A301 & ~A300;
  assign \new_[56548]_  = A299 & \new_[56547]_ ;
  assign \new_[56549]_  = \new_[56548]_  & \new_[56543]_ ;
  assign \new_[56550]_  = \new_[56549]_  & \new_[56540]_ ;
  assign \new_[56553]_  = ~A167 & ~A169;
  assign \new_[56556]_  = A199 & ~A166;
  assign \new_[56557]_  = \new_[56556]_  & \new_[56553]_ ;
  assign \new_[56560]_  = A203 & ~A200;
  assign \new_[56564]_  = ~A234 & A233;
  assign \new_[56565]_  = A232 & \new_[56564]_ ;
  assign \new_[56566]_  = \new_[56565]_  & \new_[56560]_ ;
  assign \new_[56567]_  = \new_[56566]_  & \new_[56557]_ ;
  assign \new_[56570]_  = A265 & ~A235;
  assign \new_[56573]_  = ~A267 & A266;
  assign \new_[56574]_  = \new_[56573]_  & \new_[56570]_ ;
  assign \new_[56577]_  = A298 & ~A268;
  assign \new_[56581]_  = ~A301 & ~A300;
  assign \new_[56582]_  = A299 & \new_[56581]_ ;
  assign \new_[56583]_  = \new_[56582]_  & \new_[56577]_ ;
  assign \new_[56584]_  = \new_[56583]_  & \new_[56574]_ ;
  assign \new_[56587]_  = ~A168 & ~A169;
  assign \new_[56590]_  = A166 & A167;
  assign \new_[56591]_  = \new_[56590]_  & \new_[56587]_ ;
  assign \new_[56594]_  = A201 & A199;
  assign \new_[56598]_  = ~A234 & A233;
  assign \new_[56599]_  = A232 & \new_[56598]_ ;
  assign \new_[56600]_  = \new_[56599]_  & \new_[56594]_ ;
  assign \new_[56601]_  = \new_[56600]_  & \new_[56591]_ ;
  assign \new_[56604]_  = A265 & ~A235;
  assign \new_[56607]_  = ~A267 & A266;
  assign \new_[56608]_  = \new_[56607]_  & \new_[56604]_ ;
  assign \new_[56611]_  = A298 & ~A268;
  assign \new_[56615]_  = ~A301 & ~A300;
  assign \new_[56616]_  = A299 & \new_[56615]_ ;
  assign \new_[56617]_  = \new_[56616]_  & \new_[56611]_ ;
  assign \new_[56618]_  = \new_[56617]_  & \new_[56608]_ ;
  assign \new_[56621]_  = ~A168 & ~A169;
  assign \new_[56624]_  = A166 & A167;
  assign \new_[56625]_  = \new_[56624]_  & \new_[56621]_ ;
  assign \new_[56628]_  = A201 & A200;
  assign \new_[56632]_  = ~A234 & A233;
  assign \new_[56633]_  = A232 & \new_[56632]_ ;
  assign \new_[56634]_  = \new_[56633]_  & \new_[56628]_ ;
  assign \new_[56635]_  = \new_[56634]_  & \new_[56625]_ ;
  assign \new_[56638]_  = A265 & ~A235;
  assign \new_[56641]_  = ~A267 & A266;
  assign \new_[56642]_  = \new_[56641]_  & \new_[56638]_ ;
  assign \new_[56645]_  = A298 & ~A268;
  assign \new_[56649]_  = ~A301 & ~A300;
  assign \new_[56650]_  = A299 & \new_[56649]_ ;
  assign \new_[56651]_  = \new_[56650]_  & \new_[56645]_ ;
  assign \new_[56652]_  = \new_[56651]_  & \new_[56642]_ ;
  assign \new_[56655]_  = ~A168 & ~A169;
  assign \new_[56658]_  = A166 & A167;
  assign \new_[56659]_  = \new_[56658]_  & \new_[56655]_ ;
  assign \new_[56662]_  = A200 & ~A199;
  assign \new_[56666]_  = ~A235 & ~A234;
  assign \new_[56667]_  = A203 & \new_[56666]_ ;
  assign \new_[56668]_  = \new_[56667]_  & \new_[56662]_ ;
  assign \new_[56669]_  = \new_[56668]_  & \new_[56659]_ ;
  assign \new_[56672]_  = A265 & ~A236;
  assign \new_[56675]_  = ~A267 & A266;
  assign \new_[56676]_  = \new_[56675]_  & \new_[56672]_ ;
  assign \new_[56679]_  = A298 & ~A268;
  assign \new_[56683]_  = ~A301 & ~A300;
  assign \new_[56684]_  = A299 & \new_[56683]_ ;
  assign \new_[56685]_  = \new_[56684]_  & \new_[56679]_ ;
  assign \new_[56686]_  = \new_[56685]_  & \new_[56676]_ ;
  assign \new_[56689]_  = ~A168 & ~A169;
  assign \new_[56692]_  = A166 & A167;
  assign \new_[56693]_  = \new_[56692]_  & \new_[56689]_ ;
  assign \new_[56696]_  = A200 & ~A199;
  assign \new_[56700]_  = A233 & A232;
  assign \new_[56701]_  = A203 & \new_[56700]_ ;
  assign \new_[56702]_  = \new_[56701]_  & \new_[56696]_ ;
  assign \new_[56703]_  = \new_[56702]_  & \new_[56693]_ ;
  assign \new_[56706]_  = ~A235 & ~A234;
  assign \new_[56709]_  = ~A268 & ~A267;
  assign \new_[56710]_  = \new_[56709]_  & \new_[56706]_ ;
  assign \new_[56713]_  = A298 & ~A269;
  assign \new_[56717]_  = ~A301 & ~A300;
  assign \new_[56718]_  = A299 & \new_[56717]_ ;
  assign \new_[56719]_  = \new_[56718]_  & \new_[56713]_ ;
  assign \new_[56720]_  = \new_[56719]_  & \new_[56710]_ ;
  assign \new_[56723]_  = ~A168 & ~A169;
  assign \new_[56726]_  = A166 & A167;
  assign \new_[56727]_  = \new_[56726]_  & \new_[56723]_ ;
  assign \new_[56730]_  = A200 & ~A199;
  assign \new_[56734]_  = A233 & A232;
  assign \new_[56735]_  = A203 & \new_[56734]_ ;
  assign \new_[56736]_  = \new_[56735]_  & \new_[56730]_ ;
  assign \new_[56737]_  = \new_[56736]_  & \new_[56727]_ ;
  assign \new_[56740]_  = ~A235 & ~A234;
  assign \new_[56743]_  = A266 & A265;
  assign \new_[56744]_  = \new_[56743]_  & \new_[56740]_ ;
  assign \new_[56747]_  = ~A268 & ~A267;
  assign \new_[56751]_  = ~A302 & ~A301;
  assign \new_[56752]_  = ~A300 & \new_[56751]_ ;
  assign \new_[56753]_  = \new_[56752]_  & \new_[56747]_ ;
  assign \new_[56754]_  = \new_[56753]_  & \new_[56744]_ ;
  assign \new_[56757]_  = ~A168 & ~A169;
  assign \new_[56760]_  = A166 & A167;
  assign \new_[56761]_  = \new_[56760]_  & \new_[56757]_ ;
  assign \new_[56764]_  = A200 & ~A199;
  assign \new_[56768]_  = A233 & A232;
  assign \new_[56769]_  = A203 & \new_[56768]_ ;
  assign \new_[56770]_  = \new_[56769]_  & \new_[56764]_ ;
  assign \new_[56771]_  = \new_[56770]_  & \new_[56761]_ ;
  assign \new_[56774]_  = ~A235 & ~A234;
  assign \new_[56777]_  = A266 & A265;
  assign \new_[56778]_  = \new_[56777]_  & \new_[56774]_ ;
  assign \new_[56781]_  = ~A268 & ~A267;
  assign \new_[56785]_  = ~A301 & ~A299;
  assign \new_[56786]_  = ~A298 & \new_[56785]_ ;
  assign \new_[56787]_  = \new_[56786]_  & \new_[56781]_ ;
  assign \new_[56788]_  = \new_[56787]_  & \new_[56778]_ ;
  assign \new_[56791]_  = ~A168 & ~A169;
  assign \new_[56794]_  = A166 & A167;
  assign \new_[56795]_  = \new_[56794]_  & \new_[56791]_ ;
  assign \new_[56798]_  = A200 & ~A199;
  assign \new_[56802]_  = A233 & A232;
  assign \new_[56803]_  = A203 & \new_[56802]_ ;
  assign \new_[56804]_  = \new_[56803]_  & \new_[56798]_ ;
  assign \new_[56805]_  = \new_[56804]_  & \new_[56795]_ ;
  assign \new_[56808]_  = ~A235 & ~A234;
  assign \new_[56811]_  = ~A266 & ~A265;
  assign \new_[56812]_  = \new_[56811]_  & \new_[56808]_ ;
  assign \new_[56815]_  = A298 & ~A268;
  assign \new_[56819]_  = ~A301 & ~A300;
  assign \new_[56820]_  = A299 & \new_[56819]_ ;
  assign \new_[56821]_  = \new_[56820]_  & \new_[56815]_ ;
  assign \new_[56822]_  = \new_[56821]_  & \new_[56812]_ ;
  assign \new_[56825]_  = ~A168 & ~A169;
  assign \new_[56828]_  = A166 & A167;
  assign \new_[56829]_  = \new_[56828]_  & \new_[56825]_ ;
  assign \new_[56832]_  = A200 & ~A199;
  assign \new_[56836]_  = ~A233 & ~A232;
  assign \new_[56837]_  = A203 & \new_[56836]_ ;
  assign \new_[56838]_  = \new_[56837]_  & \new_[56832]_ ;
  assign \new_[56839]_  = \new_[56838]_  & \new_[56829]_ ;
  assign \new_[56842]_  = A265 & ~A235;
  assign \new_[56845]_  = ~A267 & A266;
  assign \new_[56846]_  = \new_[56845]_  & \new_[56842]_ ;
  assign \new_[56849]_  = A298 & ~A268;
  assign \new_[56853]_  = ~A301 & ~A300;
  assign \new_[56854]_  = A299 & \new_[56853]_ ;
  assign \new_[56855]_  = \new_[56854]_  & \new_[56849]_ ;
  assign \new_[56856]_  = \new_[56855]_  & \new_[56846]_ ;
  assign \new_[56859]_  = ~A168 & ~A169;
  assign \new_[56862]_  = A166 & A167;
  assign \new_[56863]_  = \new_[56862]_  & \new_[56859]_ ;
  assign \new_[56866]_  = ~A200 & A199;
  assign \new_[56870]_  = ~A235 & ~A234;
  assign \new_[56871]_  = A203 & \new_[56870]_ ;
  assign \new_[56872]_  = \new_[56871]_  & \new_[56866]_ ;
  assign \new_[56873]_  = \new_[56872]_  & \new_[56863]_ ;
  assign \new_[56876]_  = A265 & ~A236;
  assign \new_[56879]_  = ~A267 & A266;
  assign \new_[56880]_  = \new_[56879]_  & \new_[56876]_ ;
  assign \new_[56883]_  = A298 & ~A268;
  assign \new_[56887]_  = ~A301 & ~A300;
  assign \new_[56888]_  = A299 & \new_[56887]_ ;
  assign \new_[56889]_  = \new_[56888]_  & \new_[56883]_ ;
  assign \new_[56890]_  = \new_[56889]_  & \new_[56880]_ ;
  assign \new_[56893]_  = ~A168 & ~A169;
  assign \new_[56896]_  = A166 & A167;
  assign \new_[56897]_  = \new_[56896]_  & \new_[56893]_ ;
  assign \new_[56900]_  = ~A200 & A199;
  assign \new_[56904]_  = A233 & A232;
  assign \new_[56905]_  = A203 & \new_[56904]_ ;
  assign \new_[56906]_  = \new_[56905]_  & \new_[56900]_ ;
  assign \new_[56907]_  = \new_[56906]_  & \new_[56897]_ ;
  assign \new_[56910]_  = ~A235 & ~A234;
  assign \new_[56913]_  = ~A268 & ~A267;
  assign \new_[56914]_  = \new_[56913]_  & \new_[56910]_ ;
  assign \new_[56917]_  = A298 & ~A269;
  assign \new_[56921]_  = ~A301 & ~A300;
  assign \new_[56922]_  = A299 & \new_[56921]_ ;
  assign \new_[56923]_  = \new_[56922]_  & \new_[56917]_ ;
  assign \new_[56924]_  = \new_[56923]_  & \new_[56914]_ ;
  assign \new_[56927]_  = ~A168 & ~A169;
  assign \new_[56930]_  = A166 & A167;
  assign \new_[56931]_  = \new_[56930]_  & \new_[56927]_ ;
  assign \new_[56934]_  = ~A200 & A199;
  assign \new_[56938]_  = A233 & A232;
  assign \new_[56939]_  = A203 & \new_[56938]_ ;
  assign \new_[56940]_  = \new_[56939]_  & \new_[56934]_ ;
  assign \new_[56941]_  = \new_[56940]_  & \new_[56931]_ ;
  assign \new_[56944]_  = ~A235 & ~A234;
  assign \new_[56947]_  = A266 & A265;
  assign \new_[56948]_  = \new_[56947]_  & \new_[56944]_ ;
  assign \new_[56951]_  = ~A268 & ~A267;
  assign \new_[56955]_  = ~A302 & ~A301;
  assign \new_[56956]_  = ~A300 & \new_[56955]_ ;
  assign \new_[56957]_  = \new_[56956]_  & \new_[56951]_ ;
  assign \new_[56958]_  = \new_[56957]_  & \new_[56948]_ ;
  assign \new_[56961]_  = ~A168 & ~A169;
  assign \new_[56964]_  = A166 & A167;
  assign \new_[56965]_  = \new_[56964]_  & \new_[56961]_ ;
  assign \new_[56968]_  = ~A200 & A199;
  assign \new_[56972]_  = A233 & A232;
  assign \new_[56973]_  = A203 & \new_[56972]_ ;
  assign \new_[56974]_  = \new_[56973]_  & \new_[56968]_ ;
  assign \new_[56975]_  = \new_[56974]_  & \new_[56965]_ ;
  assign \new_[56978]_  = ~A235 & ~A234;
  assign \new_[56981]_  = A266 & A265;
  assign \new_[56982]_  = \new_[56981]_  & \new_[56978]_ ;
  assign \new_[56985]_  = ~A268 & ~A267;
  assign \new_[56989]_  = ~A301 & ~A299;
  assign \new_[56990]_  = ~A298 & \new_[56989]_ ;
  assign \new_[56991]_  = \new_[56990]_  & \new_[56985]_ ;
  assign \new_[56992]_  = \new_[56991]_  & \new_[56982]_ ;
  assign \new_[56995]_  = ~A168 & ~A169;
  assign \new_[56998]_  = A166 & A167;
  assign \new_[56999]_  = \new_[56998]_  & \new_[56995]_ ;
  assign \new_[57002]_  = ~A200 & A199;
  assign \new_[57006]_  = A233 & A232;
  assign \new_[57007]_  = A203 & \new_[57006]_ ;
  assign \new_[57008]_  = \new_[57007]_  & \new_[57002]_ ;
  assign \new_[57009]_  = \new_[57008]_  & \new_[56999]_ ;
  assign \new_[57012]_  = ~A235 & ~A234;
  assign \new_[57015]_  = ~A266 & ~A265;
  assign \new_[57016]_  = \new_[57015]_  & \new_[57012]_ ;
  assign \new_[57019]_  = A298 & ~A268;
  assign \new_[57023]_  = ~A301 & ~A300;
  assign \new_[57024]_  = A299 & \new_[57023]_ ;
  assign \new_[57025]_  = \new_[57024]_  & \new_[57019]_ ;
  assign \new_[57026]_  = \new_[57025]_  & \new_[57016]_ ;
  assign \new_[57029]_  = ~A168 & ~A169;
  assign \new_[57032]_  = A166 & A167;
  assign \new_[57033]_  = \new_[57032]_  & \new_[57029]_ ;
  assign \new_[57036]_  = ~A200 & A199;
  assign \new_[57040]_  = ~A233 & ~A232;
  assign \new_[57041]_  = A203 & \new_[57040]_ ;
  assign \new_[57042]_  = \new_[57041]_  & \new_[57036]_ ;
  assign \new_[57043]_  = \new_[57042]_  & \new_[57033]_ ;
  assign \new_[57046]_  = A265 & ~A235;
  assign \new_[57049]_  = ~A267 & A266;
  assign \new_[57050]_  = \new_[57049]_  & \new_[57046]_ ;
  assign \new_[57053]_  = A298 & ~A268;
  assign \new_[57057]_  = ~A301 & ~A300;
  assign \new_[57058]_  = A299 & \new_[57057]_ ;
  assign \new_[57059]_  = \new_[57058]_  & \new_[57053]_ ;
  assign \new_[57060]_  = \new_[57059]_  & \new_[57050]_ ;
  assign \new_[57063]_  = ~A169 & ~A170;
  assign \new_[57066]_  = ~A199 & ~A168;
  assign \new_[57067]_  = \new_[57066]_  & \new_[57063]_ ;
  assign \new_[57070]_  = A203 & A200;
  assign \new_[57074]_  = ~A234 & A233;
  assign \new_[57075]_  = A232 & \new_[57074]_ ;
  assign \new_[57076]_  = \new_[57075]_  & \new_[57070]_ ;
  assign \new_[57077]_  = \new_[57076]_  & \new_[57067]_ ;
  assign \new_[57080]_  = A265 & ~A235;
  assign \new_[57083]_  = ~A267 & A266;
  assign \new_[57084]_  = \new_[57083]_  & \new_[57080]_ ;
  assign \new_[57087]_  = A298 & ~A268;
  assign \new_[57091]_  = ~A301 & ~A300;
  assign \new_[57092]_  = A299 & \new_[57091]_ ;
  assign \new_[57093]_  = \new_[57092]_  & \new_[57087]_ ;
  assign \new_[57094]_  = \new_[57093]_  & \new_[57084]_ ;
  assign \new_[57097]_  = ~A169 & ~A170;
  assign \new_[57100]_  = A199 & ~A168;
  assign \new_[57101]_  = \new_[57100]_  & \new_[57097]_ ;
  assign \new_[57104]_  = A203 & ~A200;
  assign \new_[57108]_  = ~A234 & A233;
  assign \new_[57109]_  = A232 & \new_[57108]_ ;
  assign \new_[57110]_  = \new_[57109]_  & \new_[57104]_ ;
  assign \new_[57111]_  = \new_[57110]_  & \new_[57101]_ ;
  assign \new_[57114]_  = A265 & ~A235;
  assign \new_[57117]_  = ~A267 & A266;
  assign \new_[57118]_  = \new_[57117]_  & \new_[57114]_ ;
  assign \new_[57121]_  = A298 & ~A268;
  assign \new_[57125]_  = ~A301 & ~A300;
  assign \new_[57126]_  = A299 & \new_[57125]_ ;
  assign \new_[57127]_  = \new_[57126]_  & \new_[57121]_ ;
  assign \new_[57128]_  = \new_[57127]_  & \new_[57118]_ ;
  assign \new_[57131]_  = A167 & A170;
  assign \new_[57134]_  = A199 & ~A166;
  assign \new_[57135]_  = \new_[57134]_  & \new_[57131]_ ;
  assign \new_[57138]_  = ~A201 & A200;
  assign \new_[57142]_  = A233 & A232;
  assign \new_[57143]_  = ~A202 & \new_[57142]_ ;
  assign \new_[57144]_  = \new_[57143]_  & \new_[57138]_ ;
  assign \new_[57145]_  = \new_[57144]_  & \new_[57135]_ ;
  assign \new_[57148]_  = ~A235 & ~A234;
  assign \new_[57152]_  = ~A267 & A266;
  assign \new_[57153]_  = A265 & \new_[57152]_ ;
  assign \new_[57154]_  = \new_[57153]_  & \new_[57148]_ ;
  assign \new_[57157]_  = A298 & ~A268;
  assign \new_[57161]_  = ~A301 & ~A300;
  assign \new_[57162]_  = A299 & \new_[57161]_ ;
  assign \new_[57163]_  = \new_[57162]_  & \new_[57157]_ ;
  assign \new_[57164]_  = \new_[57163]_  & \new_[57154]_ ;
  assign \new_[57167]_  = ~A167 & A170;
  assign \new_[57170]_  = A199 & A166;
  assign \new_[57171]_  = \new_[57170]_  & \new_[57167]_ ;
  assign \new_[57174]_  = ~A201 & A200;
  assign \new_[57178]_  = A233 & A232;
  assign \new_[57179]_  = ~A202 & \new_[57178]_ ;
  assign \new_[57180]_  = \new_[57179]_  & \new_[57174]_ ;
  assign \new_[57181]_  = \new_[57180]_  & \new_[57171]_ ;
  assign \new_[57184]_  = ~A235 & ~A234;
  assign \new_[57188]_  = ~A267 & A266;
  assign \new_[57189]_  = A265 & \new_[57188]_ ;
  assign \new_[57190]_  = \new_[57189]_  & \new_[57184]_ ;
  assign \new_[57193]_  = A298 & ~A268;
  assign \new_[57197]_  = ~A301 & ~A300;
  assign \new_[57198]_  = A299 & \new_[57197]_ ;
  assign \new_[57199]_  = \new_[57198]_  & \new_[57193]_ ;
  assign \new_[57200]_  = \new_[57199]_  & \new_[57190]_ ;
  assign \new_[57203]_  = ~A168 & ~A169;
  assign \new_[57206]_  = A166 & A167;
  assign \new_[57207]_  = \new_[57206]_  & \new_[57203]_ ;
  assign \new_[57210]_  = A200 & ~A199;
  assign \new_[57214]_  = A233 & A232;
  assign \new_[57215]_  = A203 & \new_[57214]_ ;
  assign \new_[57216]_  = \new_[57215]_  & \new_[57210]_ ;
  assign \new_[57217]_  = \new_[57216]_  & \new_[57207]_ ;
  assign \new_[57220]_  = ~A235 & ~A234;
  assign \new_[57224]_  = ~A267 & A266;
  assign \new_[57225]_  = A265 & \new_[57224]_ ;
  assign \new_[57226]_  = \new_[57225]_  & \new_[57220]_ ;
  assign \new_[57229]_  = A298 & ~A268;
  assign \new_[57233]_  = ~A301 & ~A300;
  assign \new_[57234]_  = A299 & \new_[57233]_ ;
  assign \new_[57235]_  = \new_[57234]_  & \new_[57229]_ ;
  assign \new_[57236]_  = \new_[57235]_  & \new_[57226]_ ;
  assign \new_[57239]_  = ~A168 & ~A169;
  assign \new_[57242]_  = A166 & A167;
  assign \new_[57243]_  = \new_[57242]_  & \new_[57239]_ ;
  assign \new_[57246]_  = ~A200 & A199;
  assign \new_[57250]_  = A233 & A232;
  assign \new_[57251]_  = A203 & \new_[57250]_ ;
  assign \new_[57252]_  = \new_[57251]_  & \new_[57246]_ ;
  assign \new_[57253]_  = \new_[57252]_  & \new_[57243]_ ;
  assign \new_[57256]_  = ~A235 & ~A234;
  assign \new_[57260]_  = ~A267 & A266;
  assign \new_[57261]_  = A265 & \new_[57260]_ ;
  assign \new_[57262]_  = \new_[57261]_  & \new_[57256]_ ;
  assign \new_[57265]_  = A298 & ~A268;
  assign \new_[57269]_  = ~A301 & ~A300;
  assign \new_[57270]_  = A299 & \new_[57269]_ ;
  assign \new_[57271]_  = \new_[57270]_  & \new_[57265]_ ;
  assign \new_[57272]_  = \new_[57271]_  & \new_[57262]_ ;
endmodule


