module top ( 
    pp, pq, pr, ps, pt, pu, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk, pl,
    pm, pn, po,
    pv  );
  input  pp, pq, pr, ps, pt, pu, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj,
    pk, pl, pm, pn, po;
  output pv;
  wire new_n23_, new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_,
    new_n30_, new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_,
    new_n37_, new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_,
    new_n44_, new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_,
    new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_,
    new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_,
    new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_,
    new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_,
    new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_, new_n114_, new_n115_, new_n116_, new_n117_,
    new_n118_, new_n119_, new_n120_, new_n121_, new_n122_, new_n123_,
    new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_,
    new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_,
    new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_,
    new_n142_, new_n143_, new_n144_;
  assign new_n23_ = ps & pt;
  assign new_n24_ = ~pe & new_n23_;
  assign new_n25_ = ~ps & pt;
  assign new_n26_ = ~pg & new_n25_;
  assign new_n27_ = ~ps & ~ph;
  assign new_n28_ = ~pg & new_n27_;
  assign new_n29_ = pt & ~pg;
  assign new_n30_ = ~pe & new_n29_;
  assign new_n31_ = ps & ~pf;
  assign new_n32_ = ~pe & new_n31_;
  assign new_n33_ = ~ps & ~pt;
  assign new_n34_ = ~ph & new_n33_;
  assign new_n35_ = ~pf & ~ph;
  assign new_n36_ = ~pg & new_n35_;
  assign new_n37_ = ~pe & new_n36_;
  assign new_n38_ = ~pt & ~ph;
  assign new_n39_ = ~pf & new_n38_;
  assign new_n40_ = ps & ~pt;
  assign new_n41_ = ~pf & new_n40_;
  assign new_n42_ = ~new_n39_ & ~new_n41_;
  assign new_n43_ = ~new_n34_ & ~new_n37_;
  assign new_n44_ = new_n42_ & new_n43_;
  assign new_n45_ = ~new_n30_ & ~new_n32_;
  assign new_n46_ = ~new_n24_ & ~new_n26_;
  assign new_n47_ = ~new_n28_ & new_n46_;
  assign new_n48_ = new_n45_ & new_n47_;
  assign new_n49_ = new_n44_ & new_n48_;
  assign new_n50_ = ~pr & new_n49_;
  assign new_n51_ = pq & new_n50_;
  assign new_n52_ = ~pm & new_n23_;
  assign new_n53_ = ~po & new_n25_;
  assign new_n54_ = ~pp & ~ps;
  assign new_n55_ = ~po & new_n54_;
  assign new_n56_ = pt & ~po;
  assign new_n57_ = ~pm & new_n56_;
  assign new_n58_ = ps & ~pn;
  assign new_n59_ = ~pm & new_n58_;
  assign new_n60_ = ~pp & new_n33_;
  assign new_n61_ = ~pp & ~pn;
  assign new_n62_ = ~po & new_n61_;
  assign new_n63_ = ~pm & new_n62_;
  assign new_n64_ = ~pp & ~pt;
  assign new_n65_ = ~pn & new_n64_;
  assign new_n66_ = ~pn & new_n40_;
  assign new_n67_ = ~new_n65_ & ~new_n66_;
  assign new_n68_ = ~new_n60_ & ~new_n63_;
  assign new_n69_ = new_n67_ & new_n68_;
  assign new_n70_ = ~new_n57_ & ~new_n59_;
  assign new_n71_ = ~new_n52_ & ~new_n53_;
  assign new_n72_ = ~new_n55_ & new_n71_;
  assign new_n73_ = new_n70_ & new_n72_;
  assign new_n74_ = new_n69_ & new_n73_;
  assign new_n75_ = new_n49_ & new_n74_;
  assign new_n76_ = ~pr & new_n75_;
  assign new_n77_ = ~pi & new_n23_;
  assign new_n78_ = ~pk & new_n25_;
  assign new_n79_ = ~ps & ~pl;
  assign new_n80_ = ~pk & new_n79_;
  assign new_n81_ = pt & ~pk;
  assign new_n82_ = ~pi & new_n81_;
  assign new_n83_ = ps & ~pj;
  assign new_n84_ = ~pi & new_n83_;
  assign new_n85_ = ~pl & new_n33_;
  assign new_n86_ = ~pj & ~pl;
  assign new_n87_ = ~pk & new_n86_;
  assign new_n88_ = ~pi & new_n87_;
  assign new_n89_ = ~pt & ~pl;
  assign new_n90_ = ~pj & new_n89_;
  assign new_n91_ = ~pj & new_n40_;
  assign new_n92_ = ~new_n90_ & ~new_n91_;
  assign new_n93_ = ~new_n85_ & ~new_n88_;
  assign new_n94_ = new_n92_ & new_n93_;
  assign new_n95_ = ~new_n82_ & ~new_n84_;
  assign new_n96_ = ~new_n77_ & ~new_n78_;
  assign new_n97_ = ~new_n80_ & new_n96_;
  assign new_n98_ = new_n95_ & new_n97_;
  assign new_n99_ = new_n94_ & new_n98_;
  assign new_n100_ = pr & new_n99_;
  assign new_n101_ = ~pq & new_n100_;
  assign new_n102_ = new_n74_ & new_n99_;
  assign new_n103_ = ~pq & new_n102_;
  assign new_n104_ = ~pr & new_n74_;
  assign new_n105_ = ~pq & new_n104_;
  assign new_n106_ = ~pa & new_n23_;
  assign new_n107_ = ~pc & new_n25_;
  assign new_n108_ = ~ps & ~pd;
  assign new_n109_ = ~pc & new_n108_;
  assign new_n110_ = pt & ~pc;
  assign new_n111_ = ~pa & new_n110_;
  assign new_n112_ = ps & ~pb;
  assign new_n113_ = ~pa & new_n112_;
  assign new_n114_ = ~pd & new_n33_;
  assign new_n115_ = ~pb & ~pd;
  assign new_n116_ = ~pc & new_n115_;
  assign new_n117_ = ~pa & new_n116_;
  assign new_n118_ = ~pt & ~pd;
  assign new_n119_ = ~pb & new_n118_;
  assign new_n120_ = ~pb & new_n40_;
  assign new_n121_ = ~new_n119_ & ~new_n120_;
  assign new_n122_ = ~new_n114_ & ~new_n117_;
  assign new_n123_ = new_n121_ & new_n122_;
  assign new_n124_ = ~new_n111_ & ~new_n113_;
  assign new_n125_ = ~new_n106_ & ~new_n107_;
  assign new_n126_ = ~new_n109_ & new_n125_;
  assign new_n127_ = new_n124_ & new_n126_;
  assign new_n128_ = new_n123_ & new_n127_;
  assign new_n129_ = new_n49_ & new_n128_;
  assign new_n130_ = pq & new_n129_;
  assign new_n131_ = new_n99_ & new_n128_;
  assign new_n132_ = new_n49_ & new_n131_;
  assign new_n133_ = new_n74_ & new_n132_;
  assign new_n134_ = pr & new_n128_;
  assign new_n135_ = pq & new_n134_;
  assign new_n136_ = pr & new_n131_;
  assign new_n137_ = ~new_n135_ & ~new_n136_;
  assign new_n138_ = ~new_n130_ & ~new_n133_;
  assign new_n139_ = new_n137_ & new_n138_;
  assign new_n140_ = ~new_n103_ & ~new_n105_;
  assign new_n141_ = ~new_n51_ & ~new_n76_;
  assign new_n142_ = ~new_n101_ & new_n141_;
  assign new_n143_ = new_n140_ & new_n142_;
  assign new_n144_ = new_n139_ & new_n143_;
  assign pv = pu & ~new_n144_;
endmodule

