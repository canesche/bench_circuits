module top ( clock, 
    p_10, p_12, p_11, pclk, p_14, p_13, p_16, p_15, p_9, p_18, p_8, p_17,
    p_7, p_6, p_5, p_4, p_3, p_1,
    p_36  );
  input  clock;
  input  p_10, p_12, p_11, pclk, p_14, p_13, p_16, p_15, p_9, p_18, p_8,
    p_17, p_7, p_6, p_5, p_4, p_3, p_1;
  output p_36;
  reg n_28, n_24, n_25, n_26, n_27, n_20, n_21, n_22, n_23, n_2, n_29, n_30,
    n_31, n_32, n_33, n_34;
  wire new_n68_, new_n69_, new_n70_1_, new_n72_, new_n73_, new_n74_,
    new_n75_1_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_1_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_1_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_1_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_1_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_1_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_1_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_1_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_1_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, n40, n45, n50,
    n55, n60, n65, n70, n75, n80, n85, n90, n95, n100, n105, n110, n115;
  assign new_n68_ = p_3 & p_1;
  assign new_n69_ = ~n_20 & new_n68_;
  assign new_n70_1_ = n_20 & ~new_n68_;
  assign p_36 = new_n69_ | new_n70_1_;
  assign new_n72_ = p_11 & p_1;
  assign new_n73_ = n_28 & new_n72_;
  assign new_n74_ = p_10 & p_1;
  assign new_n75_1_ = n_27 & new_n74_;
  assign new_n76_ = p_9 & p_1;
  assign new_n77_ = n_26 & new_n76_;
  assign new_n78_ = p_8 & p_1;
  assign new_n79_ = n_25 & new_n78_;
  assign new_n80_1_ = p_7 & p_1;
  assign new_n81_ = n_24 & new_n80_1_;
  assign new_n82_ = p_6 & p_1;
  assign new_n83_ = n_23 & new_n82_;
  assign new_n84_ = p_5 & p_1;
  assign new_n85_1_ = n_22 & new_n84_;
  assign new_n86_ = p_4 & p_1;
  assign new_n87_ = n_21 & new_n86_;
  assign new_n88_ = n_20 & new_n68_;
  assign new_n89_ = n_21 & new_n88_;
  assign new_n90_1_ = new_n86_ & new_n88_;
  assign new_n91_ = ~new_n87_ & ~new_n89_;
  assign new_n92_ = ~new_n90_1_ & new_n91_;
  assign new_n93_ = n_22 & ~new_n92_;
  assign new_n94_ = new_n84_ & ~new_n92_;
  assign new_n95_1_ = ~new_n85_1_ & ~new_n93_;
  assign new_n96_ = ~new_n94_ & new_n95_1_;
  assign new_n97_ = n_23 & ~new_n96_;
  assign new_n98_ = new_n82_ & ~new_n96_;
  assign new_n99_ = ~new_n83_ & ~new_n97_;
  assign new_n100_1_ = ~new_n98_ & new_n99_;
  assign new_n101_ = n_24 & ~new_n100_1_;
  assign new_n102_ = new_n80_1_ & ~new_n100_1_;
  assign new_n103_ = ~new_n81_ & ~new_n101_;
  assign new_n104_ = ~new_n102_ & new_n103_;
  assign new_n105_1_ = n_25 & ~new_n104_;
  assign new_n106_ = new_n78_ & ~new_n104_;
  assign new_n107_ = ~new_n79_ & ~new_n105_1_;
  assign new_n108_ = ~new_n106_ & new_n107_;
  assign new_n109_ = n_26 & ~new_n108_;
  assign new_n110_1_ = new_n76_ & ~new_n108_;
  assign new_n111_ = ~new_n77_ & ~new_n109_;
  assign new_n112_ = ~new_n110_1_ & new_n111_;
  assign new_n113_ = n_27 & ~new_n112_;
  assign new_n114_ = new_n74_ & ~new_n112_;
  assign new_n115_1_ = ~new_n75_1_ & ~new_n113_;
  assign new_n116_ = ~new_n114_ & new_n115_1_;
  assign new_n117_ = n_28 & ~new_n116_;
  assign new_n118_ = new_n72_ & ~new_n116_;
  assign new_n119_ = ~new_n73_ & ~new_n117_;
  assign new_n120_ = ~new_n118_ & new_n119_;
  assign new_n121_ = p_12 & p_1;
  assign new_n122_ = ~new_n120_ & new_n121_;
  assign new_n123_ = n_29 & new_n122_;
  assign new_n124_ = new_n120_ & new_n121_;
  assign new_n125_ = ~n_29 & new_n124_;
  assign new_n126_ = new_n120_ & ~new_n121_;
  assign new_n127_ = n_29 & new_n126_;
  assign new_n128_ = ~new_n120_ & ~new_n121_;
  assign new_n129_ = ~n_29 & new_n128_;
  assign new_n130_ = ~new_n123_ & ~new_n125_;
  assign new_n131_ = ~new_n127_ & ~new_n129_;
  assign n40 = ~new_n130_ | ~new_n131_;
  assign new_n133_ = n_25 & new_n106_;
  assign new_n134_ = new_n78_ & new_n104_;
  assign new_n135_ = ~n_25 & new_n134_;
  assign new_n136_ = ~new_n78_ & new_n104_;
  assign new_n137_ = n_25 & new_n136_;
  assign new_n138_ = ~new_n78_ & ~new_n104_;
  assign new_n139_ = ~n_25 & new_n138_;
  assign new_n140_ = ~new_n133_ & ~new_n135_;
  assign new_n141_ = ~new_n137_ & ~new_n139_;
  assign n45 = ~new_n140_ | ~new_n141_;
  assign new_n143_ = n_26 & new_n110_1_;
  assign new_n144_ = new_n76_ & new_n108_;
  assign new_n145_ = ~n_26 & new_n144_;
  assign new_n146_ = ~new_n76_ & new_n108_;
  assign new_n147_ = n_26 & new_n146_;
  assign new_n148_ = ~new_n76_ & ~new_n108_;
  assign new_n149_ = ~n_26 & new_n148_;
  assign new_n150_ = ~new_n143_ & ~new_n145_;
  assign new_n151_ = ~new_n147_ & ~new_n149_;
  assign n50 = ~new_n150_ | ~new_n151_;
  assign new_n153_ = n_27 & new_n114_;
  assign new_n154_ = new_n74_ & new_n112_;
  assign new_n155_ = ~n_27 & new_n154_;
  assign new_n156_ = ~new_n74_ & new_n112_;
  assign new_n157_ = n_27 & new_n156_;
  assign new_n158_ = ~new_n74_ & ~new_n112_;
  assign new_n159_ = ~n_27 & new_n158_;
  assign new_n160_ = ~new_n153_ & ~new_n155_;
  assign new_n161_ = ~new_n157_ & ~new_n159_;
  assign n55 = ~new_n160_ | ~new_n161_;
  assign new_n163_ = n_28 & new_n118_;
  assign new_n164_ = new_n72_ & new_n116_;
  assign new_n165_ = ~n_28 & new_n164_;
  assign new_n166_ = ~new_n72_ & new_n116_;
  assign new_n167_ = n_28 & new_n166_;
  assign new_n168_ = ~new_n72_ & ~new_n116_;
  assign new_n169_ = ~n_28 & new_n168_;
  assign new_n170_ = ~new_n163_ & ~new_n165_;
  assign new_n171_ = ~new_n167_ & ~new_n169_;
  assign n60 = ~new_n170_ | ~new_n171_;
  assign new_n173_ = n_21 & new_n90_1_;
  assign new_n174_ = new_n86_ & ~new_n88_;
  assign new_n175_ = ~n_21 & new_n174_;
  assign new_n176_ = ~new_n86_ & ~new_n88_;
  assign new_n177_ = n_21 & new_n176_;
  assign new_n178_ = ~new_n86_ & new_n88_;
  assign new_n179_ = ~n_21 & new_n178_;
  assign new_n180_ = ~new_n173_ & ~new_n175_;
  assign new_n181_ = ~new_n177_ & ~new_n179_;
  assign n65 = ~new_n180_ | ~new_n181_;
  assign new_n183_ = n_22 & new_n94_;
  assign new_n184_ = new_n84_ & new_n92_;
  assign new_n185_ = ~n_22 & new_n184_;
  assign new_n186_ = ~new_n84_ & new_n92_;
  assign new_n187_ = n_22 & new_n186_;
  assign new_n188_ = ~new_n84_ & ~new_n92_;
  assign new_n189_ = ~n_22 & new_n188_;
  assign new_n190_ = ~new_n183_ & ~new_n185_;
  assign new_n191_ = ~new_n187_ & ~new_n189_;
  assign n70 = ~new_n190_ | ~new_n191_;
  assign new_n193_ = n_23 & new_n98_;
  assign new_n194_ = new_n82_ & new_n96_;
  assign new_n195_ = ~n_23 & new_n194_;
  assign new_n196_ = ~new_n82_ & new_n96_;
  assign new_n197_ = n_23 & new_n196_;
  assign new_n198_ = ~new_n82_ & ~new_n96_;
  assign new_n199_ = ~n_23 & new_n198_;
  assign new_n200_ = ~new_n193_ & ~new_n195_;
  assign new_n201_ = ~new_n197_ & ~new_n199_;
  assign n75 = ~new_n200_ | ~new_n201_;
  assign new_n203_ = n_24 & new_n102_;
  assign new_n204_ = new_n80_1_ & new_n100_1_;
  assign new_n205_ = ~n_24 & new_n204_;
  assign new_n206_ = ~new_n80_1_ & new_n100_1_;
  assign new_n207_ = n_24 & new_n206_;
  assign new_n208_ = ~new_n80_1_ & ~new_n100_1_;
  assign new_n209_ = ~n_24 & new_n208_;
  assign new_n210_ = ~new_n203_ & ~new_n205_;
  assign new_n211_ = ~new_n207_ & ~new_n209_;
  assign n80 = ~new_n210_ | ~new_n211_;
  assign new_n213_ = p_17 & p_1;
  assign new_n214_ = n_34 & new_n213_;
  assign new_n215_ = p_16 & p_1;
  assign new_n216_ = n_33 & new_n215_;
  assign new_n217_ = p_15 & p_1;
  assign new_n218_ = n_32 & new_n217_;
  assign new_n219_ = p_14 & p_1;
  assign new_n220_ = n_31 & new_n219_;
  assign new_n221_ = p_13 & p_1;
  assign new_n222_ = n_30 & new_n221_;
  assign new_n223_ = n_29 & new_n121_;
  assign new_n224_ = n_29 & ~new_n120_;
  assign new_n225_ = ~new_n223_ & ~new_n224_;
  assign new_n226_ = ~new_n122_ & new_n225_;
  assign new_n227_ = n_30 & ~new_n226_;
  assign new_n228_ = new_n221_ & ~new_n226_;
  assign new_n229_ = ~new_n222_ & ~new_n227_;
  assign new_n230_ = ~new_n228_ & new_n229_;
  assign new_n231_ = n_31 & ~new_n230_;
  assign new_n232_ = new_n219_ & ~new_n230_;
  assign new_n233_ = ~new_n220_ & ~new_n231_;
  assign new_n234_ = ~new_n232_ & new_n233_;
  assign new_n235_ = n_32 & ~new_n234_;
  assign new_n236_ = new_n217_ & ~new_n234_;
  assign new_n237_ = ~new_n218_ & ~new_n235_;
  assign new_n238_ = ~new_n236_ & new_n237_;
  assign new_n239_ = n_33 & ~new_n238_;
  assign new_n240_ = new_n215_ & ~new_n238_;
  assign new_n241_ = ~new_n216_ & ~new_n239_;
  assign new_n242_ = ~new_n240_ & new_n241_;
  assign new_n243_ = n_34 & ~new_n242_;
  assign new_n244_ = new_n213_ & ~new_n242_;
  assign new_n245_ = ~new_n214_ & ~new_n243_;
  assign new_n246_ = ~new_n244_ & new_n245_;
  assign new_n247_ = p_18 & p_1;
  assign new_n248_ = n_2 & new_n247_;
  assign new_n249_ = new_n246_ & new_n248_;
  assign new_n250_ = n_2 & ~new_n247_;
  assign new_n251_ = ~new_n246_ & new_n250_;
  assign new_n252_ = ~new_n249_ & ~new_n251_;
  assign new_n253_ = ~n_2 & new_n247_;
  assign new_n254_ = ~new_n246_ & new_n253_;
  assign new_n255_ = ~new_n246_ & new_n248_;
  assign new_n256_ = ~new_n254_ & ~new_n255_;
  assign n85 = ~new_n252_ | ~new_n256_;
  assign new_n258_ = n_30 & new_n228_;
  assign new_n259_ = new_n221_ & new_n226_;
  assign new_n260_ = ~n_30 & new_n259_;
  assign new_n261_ = ~new_n221_ & new_n226_;
  assign new_n262_ = n_30 & new_n261_;
  assign new_n263_ = ~new_n221_ & ~new_n226_;
  assign new_n264_ = ~n_30 & new_n263_;
  assign new_n265_ = ~new_n258_ & ~new_n260_;
  assign new_n266_ = ~new_n262_ & ~new_n264_;
  assign n90 = ~new_n265_ | ~new_n266_;
  assign new_n268_ = n_31 & new_n232_;
  assign new_n269_ = new_n219_ & new_n230_;
  assign new_n270_ = ~n_31 & new_n269_;
  assign new_n271_ = ~new_n219_ & new_n230_;
  assign new_n272_ = n_31 & new_n271_;
  assign new_n273_ = ~new_n219_ & ~new_n230_;
  assign new_n274_ = ~n_31 & new_n273_;
  assign new_n275_ = ~new_n268_ & ~new_n270_;
  assign new_n276_ = ~new_n272_ & ~new_n274_;
  assign n95 = ~new_n275_ | ~new_n276_;
  assign new_n278_ = n_32 & new_n236_;
  assign new_n279_ = new_n217_ & new_n234_;
  assign new_n280_ = ~n_32 & new_n279_;
  assign new_n281_ = ~new_n217_ & new_n234_;
  assign new_n282_ = n_32 & new_n281_;
  assign new_n283_ = ~new_n217_ & ~new_n234_;
  assign new_n284_ = ~n_32 & new_n283_;
  assign new_n285_ = ~new_n278_ & ~new_n280_;
  assign new_n286_ = ~new_n282_ & ~new_n284_;
  assign n100 = ~new_n285_ | ~new_n286_;
  assign new_n288_ = n_33 & new_n240_;
  assign new_n289_ = new_n215_ & new_n238_;
  assign new_n290_ = ~n_33 & new_n289_;
  assign new_n291_ = ~new_n215_ & new_n238_;
  assign new_n292_ = n_33 & new_n291_;
  assign new_n293_ = ~new_n215_ & ~new_n238_;
  assign new_n294_ = ~n_33 & new_n293_;
  assign new_n295_ = ~new_n288_ & ~new_n290_;
  assign new_n296_ = ~new_n292_ & ~new_n294_;
  assign n105 = ~new_n295_ | ~new_n296_;
  assign new_n298_ = n_34 & new_n244_;
  assign new_n299_ = new_n213_ & new_n242_;
  assign new_n300_ = ~n_34 & new_n299_;
  assign new_n301_ = ~new_n213_ & new_n242_;
  assign new_n302_ = n_34 & new_n301_;
  assign new_n303_ = ~new_n213_ & ~new_n242_;
  assign new_n304_ = ~n_34 & new_n303_;
  assign new_n305_ = ~new_n298_ & ~new_n300_;
  assign new_n306_ = ~new_n302_ & ~new_n304_;
  assign n110 = ~new_n305_ | ~new_n306_;
  assign new_n308_ = ~new_n246_ & ~new_n247_;
  assign new_n309_ = new_n246_ & new_n247_;
  assign new_n310_ = ~new_n308_ & ~new_n309_;
  assign new_n311_ = ~n_2 & ~new_n310_;
  assign new_n312_ = n_2 & new_n310_;
  assign n115 = new_n311_ | new_n312_;
  always @ (posedge clock) begin
    n_28 <= n40;
    n_24 <= n45;
    n_25 <= n50;
    n_26 <= n55;
    n_27 <= n60;
    n_20 <= n65;
    n_21 <= n70;
    n_22 <= n75;
    n_23 <= n80;
    n_2 <= n85;
    n_29 <= n90;
    n_30 <= n95;
    n_31 <= n100;
    n_32 <= n105;
    n_33 <= n110;
    n_34 <= n115;
  end
endmodule

