// Benchmark "testing" written by ABC on Thu Oct  8 22:16:45 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A108  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A108;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ , \new_[350]_ ,
    \new_[351]_ , \new_[352]_ , \new_[353]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[405]_ ,
    \new_[406]_ , \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ ,
    \new_[411]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[436]_ , \new_[437]_ , \new_[438]_ , \new_[439]_ , \new_[440]_ ,
    \new_[441]_ , \new_[442]_ , \new_[443]_ , \new_[444]_ , \new_[445]_ ,
    \new_[446]_ , \new_[447]_ , \new_[448]_ , \new_[449]_ , \new_[450]_ ,
    \new_[451]_ , \new_[452]_ , \new_[453]_ , \new_[454]_ , \new_[455]_ ,
    \new_[456]_ , \new_[460]_ , \new_[461]_ , \new_[464]_ , \new_[467]_ ,
    \new_[468]_ , \new_[469]_ , \new_[473]_ , \new_[474]_ , \new_[477]_ ,
    \new_[480]_ , \new_[481]_ , \new_[482]_ , \new_[483]_ , \new_[487]_ ,
    \new_[488]_ , \new_[491]_ , \new_[494]_ , \new_[495]_ , \new_[496]_ ,
    \new_[500]_ , \new_[501]_ , \new_[504]_ , \new_[507]_ , \new_[508]_ ,
    \new_[509]_ , \new_[510]_ , \new_[511]_ , \new_[515]_ , \new_[516]_ ,
    \new_[519]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[528]_ ,
    \new_[529]_ , \new_[532]_ , \new_[535]_ , \new_[536]_ , \new_[537]_ ,
    \new_[538]_ , \new_[542]_ , \new_[543]_ , \new_[546]_ , \new_[549]_ ,
    \new_[550]_ , \new_[551]_ , \new_[554]_ , \new_[557]_ , \new_[558]_ ,
    \new_[561]_ , \new_[564]_ , \new_[565]_ , \new_[566]_ , \new_[567]_ ,
    \new_[568]_ , \new_[569]_ , \new_[573]_ , \new_[574]_ , \new_[577]_ ,
    \new_[580]_ , \new_[581]_ , \new_[582]_ , \new_[586]_ , \new_[587]_ ,
    \new_[590]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ , \new_[596]_ ,
    \new_[600]_ , \new_[601]_ , \new_[604]_ , \new_[607]_ , \new_[608]_ ,
    \new_[609]_ , \new_[613]_ , \new_[614]_ , \new_[617]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[628]_ ,
    \new_[629]_ , \new_[632]_ , \new_[635]_ , \new_[636]_ , \new_[637]_ ,
    \new_[641]_ , \new_[642]_ , \new_[645]_ , \new_[648]_ , \new_[649]_ ,
    \new_[650]_ , \new_[651]_ , \new_[655]_ , \new_[656]_ , \new_[659]_ ,
    \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[667]_ , \new_[670]_ ,
    \new_[671]_ , \new_[674]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ ,
    \new_[680]_ , \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[687]_ ,
    \new_[688]_ , \new_[691]_ , \new_[694]_ , \new_[695]_ , \new_[696]_ ,
    \new_[700]_ , \new_[701]_ , \new_[704]_ , \new_[707]_ , \new_[708]_ ,
    \new_[709]_ , \new_[710]_ , \new_[714]_ , \new_[715]_ , \new_[718]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[727]_ , \new_[728]_ ,
    \new_[731]_ , \new_[734]_ , \new_[735]_ , \new_[736]_ , \new_[737]_ ,
    \new_[738]_ , \new_[742]_ , \new_[743]_ , \new_[746]_ , \new_[749]_ ,
    \new_[750]_ , \new_[751]_ , \new_[755]_ , \new_[756]_ , \new_[759]_ ,
    \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ , \new_[769]_ ,
    \new_[770]_ , \new_[773]_ , \new_[776]_ , \new_[777]_ , \new_[778]_ ,
    \new_[781]_ , \new_[784]_ , \new_[785]_ , \new_[788]_ , \new_[791]_ ,
    \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ , \new_[796]_ ,
    \new_[800]_ , \new_[801]_ , \new_[804]_ , \new_[807]_ , \new_[808]_ ,
    \new_[809]_ , \new_[813]_ , \new_[814]_ , \new_[817]_ , \new_[820]_ ,
    \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[827]_ , \new_[828]_ ,
    \new_[831]_ , \new_[834]_ , \new_[835]_ , \new_[836]_ , \new_[840]_ ,
    \new_[841]_ , \new_[844]_ , \new_[847]_ , \new_[848]_ , \new_[849]_ ,
    \new_[850]_ , \new_[851]_ , \new_[855]_ , \new_[856]_ , \new_[859]_ ,
    \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[868]_ , \new_[869]_ ,
    \new_[872]_ , \new_[875]_ , \new_[876]_ , \new_[877]_ , \new_[878]_ ,
    \new_[882]_ , \new_[883]_ , \new_[886]_ , \new_[889]_ , \new_[890]_ ,
    \new_[891]_ , \new_[894]_ , \new_[897]_ , \new_[898]_ , \new_[901]_ ,
    \new_[904]_ , \new_[905]_ , \new_[906]_ , \new_[907]_ , \new_[908]_ ,
    \new_[909]_ , \new_[910]_ , \new_[911]_ , \new_[915]_ , \new_[916]_ ,
    \new_[919]_ , \new_[922]_ , \new_[923]_ , \new_[924]_ , \new_[928]_ ,
    \new_[929]_ , \new_[932]_ , \new_[935]_ , \new_[936]_ , \new_[937]_ ,
    \new_[938]_ , \new_[942]_ , \new_[943]_ , \new_[946]_ , \new_[949]_ ,
    \new_[950]_ , \new_[951]_ , \new_[955]_ , \new_[956]_ , \new_[959]_ ,
    \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ , \new_[966]_ ,
    \new_[970]_ , \new_[971]_ , \new_[974]_ , \new_[977]_ , \new_[978]_ ,
    \new_[979]_ , \new_[983]_ , \new_[984]_ , \new_[987]_ , \new_[990]_ ,
    \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[997]_ , \new_[998]_ ,
    \new_[1001]_ , \new_[1004]_ , \new_[1005]_ , \new_[1006]_ ,
    \new_[1009]_ , \new_[1012]_ , \new_[1013]_ , \new_[1016]_ ,
    \new_[1019]_ , \new_[1020]_ , \new_[1021]_ , \new_[1022]_ ,
    \new_[1023]_ , \new_[1024]_ , \new_[1028]_ , \new_[1029]_ ,
    \new_[1032]_ , \new_[1035]_ , \new_[1036]_ , \new_[1037]_ ,
    \new_[1041]_ , \new_[1042]_ , \new_[1045]_ , \new_[1048]_ ,
    \new_[1049]_ , \new_[1050]_ , \new_[1051]_ , \new_[1055]_ ,
    \new_[1056]_ , \new_[1059]_ , \new_[1062]_ , \new_[1063]_ ,
    \new_[1064]_ , \new_[1068]_ , \new_[1069]_ , \new_[1072]_ ,
    \new_[1075]_ , \new_[1076]_ , \new_[1077]_ , \new_[1078]_ ,
    \new_[1079]_ , \new_[1083]_ , \new_[1084]_ , \new_[1087]_ ,
    \new_[1090]_ , \new_[1091]_ , \new_[1092]_ , \new_[1096]_ ,
    \new_[1097]_ , \new_[1100]_ , \new_[1103]_ , \new_[1104]_ ,
    \new_[1105]_ , \new_[1106]_ , \new_[1110]_ , \new_[1111]_ ,
    \new_[1114]_ , \new_[1117]_ , \new_[1118]_ , \new_[1119]_ ,
    \new_[1122]_ , \new_[1125]_ , \new_[1126]_ , \new_[1129]_ ,
    \new_[1132]_ , \new_[1133]_ , \new_[1134]_ , \new_[1135]_ ,
    \new_[1136]_ , \new_[1137]_ , \new_[1138]_ , \new_[1142]_ ,
    \new_[1143]_ , \new_[1146]_ , \new_[1149]_ , \new_[1150]_ ,
    \new_[1151]_ , \new_[1155]_ , \new_[1156]_ , \new_[1159]_ ,
    \new_[1162]_ , \new_[1163]_ , \new_[1164]_ , \new_[1165]_ ,
    \new_[1169]_ , \new_[1170]_ , \new_[1173]_ , \new_[1176]_ ,
    \new_[1177]_ , \new_[1178]_ , \new_[1182]_ , \new_[1183]_ ,
    \new_[1186]_ , \new_[1189]_ , \new_[1190]_ , \new_[1191]_ ,
    \new_[1192]_ , \new_[1193]_ , \new_[1197]_ , \new_[1198]_ ,
    \new_[1201]_ , \new_[1204]_ , \new_[1205]_ , \new_[1206]_ ,
    \new_[1210]_ , \new_[1211]_ , \new_[1214]_ , \new_[1217]_ ,
    \new_[1218]_ , \new_[1219]_ , \new_[1220]_ , \new_[1224]_ ,
    \new_[1225]_ , \new_[1228]_ , \new_[1231]_ , \new_[1232]_ ,
    \new_[1233]_ , \new_[1236]_ , \new_[1239]_ , \new_[1240]_ ,
    \new_[1243]_ , \new_[1246]_ , \new_[1247]_ , \new_[1248]_ ,
    \new_[1249]_ , \new_[1250]_ , \new_[1251]_ , \new_[1255]_ ,
    \new_[1256]_ , \new_[1259]_ , \new_[1262]_ , \new_[1263]_ ,
    \new_[1264]_ , \new_[1268]_ , \new_[1269]_ , \new_[1272]_ ,
    \new_[1275]_ , \new_[1276]_ , \new_[1277]_ , \new_[1278]_ ,
    \new_[1282]_ , \new_[1283]_ , \new_[1286]_ , \new_[1289]_ ,
    \new_[1290]_ , \new_[1291]_ , \new_[1295]_ , \new_[1296]_ ,
    \new_[1299]_ , \new_[1302]_ , \new_[1303]_ , \new_[1304]_ ,
    \new_[1305]_ , \new_[1306]_ , \new_[1310]_ , \new_[1311]_ ,
    \new_[1314]_ , \new_[1317]_ , \new_[1318]_ , \new_[1319]_ ,
    \new_[1323]_ , \new_[1324]_ , \new_[1327]_ , \new_[1330]_ ,
    \new_[1331]_ , \new_[1332]_ , \new_[1333]_ , \new_[1337]_ ,
    \new_[1338]_ , \new_[1341]_ , \new_[1344]_ , \new_[1345]_ ,
    \new_[1346]_ , \new_[1349]_ , \new_[1352]_ , \new_[1353]_ ,
    \new_[1356]_ , \new_[1359]_ , \new_[1360]_ , \new_[1361]_ ,
    \new_[1362]_ , \new_[1363]_ , \new_[1364]_ , \new_[1365]_ ,
    \new_[1366]_ , \new_[1369]_ , \new_[1373]_ , \new_[1374]_ ,
    \new_[1377]_ , \new_[1381]_ , \new_[1382]_ , \new_[1386]_ ,
    \new_[1387]_ , \new_[1391]_ , \new_[1392]_ , \new_[1396]_ ,
    \new_[1397]_ , \new_[1401]_ , \new_[1402]_ , \new_[1406]_ ,
    \new_[1407]_ , \new_[1411]_ , \new_[1412]_ , \new_[1416]_ ,
    \new_[1417]_ , \new_[1421]_ , \new_[1422]_ , \new_[1426]_ ,
    \new_[1427]_ , \new_[1431]_ , \new_[1432]_ , \new_[1436]_ ,
    \new_[1437]_ , \new_[1441]_ , \new_[1442]_ , \new_[1446]_ ,
    \new_[1447]_ , \new_[1450]_ , \new_[1453]_ , \new_[1454]_ ,
    \new_[1458]_ , \new_[1459]_ , \new_[1462]_ , \new_[1465]_ ,
    \new_[1466]_ , \new_[1470]_ , \new_[1471]_ , \new_[1474]_ ,
    \new_[1477]_ , \new_[1478]_ , \new_[1482]_ , \new_[1483]_ ,
    \new_[1486]_ , \new_[1489]_ , \new_[1490]_ , \new_[1493]_ ,
    \new_[1496]_ , \new_[1497]_ , \new_[1500]_ , \new_[1503]_ ,
    \new_[1504]_ , \new_[1507]_ , \new_[1510]_ , \new_[1511]_ ,
    \new_[1514]_ , \new_[1517]_ , \new_[1518]_ , \new_[1521]_ ,
    \new_[1524]_ , \new_[1525]_ , \new_[1528]_ , \new_[1531]_ ,
    \new_[1532]_ , \new_[1535]_ , \new_[1538]_ , \new_[1539]_ ,
    \new_[1542]_ , \new_[1545]_ , \new_[1546]_ , \new_[1549]_ ,
    \new_[1552]_ , \new_[1553]_ , \new_[1556]_ , \new_[1559]_ ,
    \new_[1560]_ , \new_[1563]_ , \new_[1566]_ , \new_[1567]_ ,
    \new_[1570]_ , \new_[1573]_ , \new_[1574]_ , \new_[1577]_ ,
    \new_[1580]_ , \new_[1581]_ , \new_[1584]_ , \new_[1587]_ ,
    \new_[1588]_ , \new_[1591]_ , \new_[1594]_ , \new_[1595]_ ,
    \new_[1598]_ , \new_[1601]_ , \new_[1602]_ , \new_[1605]_ ,
    \new_[1608]_ , \new_[1609]_ , \new_[1612]_ , \new_[1615]_ ,
    \new_[1616]_ , \new_[1619]_ , \new_[1622]_ , \new_[1623]_ ,
    \new_[1626]_ , \new_[1629]_ , \new_[1630]_ , \new_[1633]_ ,
    \new_[1636]_ , \new_[1637]_ , \new_[1640]_ , \new_[1643]_ ,
    \new_[1644]_ , \new_[1647]_ , \new_[1650]_ , \new_[1651]_ ,
    \new_[1654]_ , \new_[1657]_ , \new_[1658]_ , \new_[1661]_ ,
    \new_[1664]_ , \new_[1665]_ , \new_[1668]_ , \new_[1671]_ ,
    \new_[1672]_ , \new_[1675]_ , \new_[1678]_ , \new_[1679]_ ,
    \new_[1682]_ , \new_[1685]_ , \new_[1686]_ , \new_[1689]_ ,
    \new_[1692]_ , \new_[1693]_ , \new_[1696]_ , \new_[1699]_ ,
    \new_[1700]_ , \new_[1703]_ , \new_[1706]_ , \new_[1707]_ ,
    \new_[1710]_ , \new_[1713]_ , \new_[1714]_ , \new_[1717]_ ,
    \new_[1720]_ , \new_[1721]_ , \new_[1724]_ , \new_[1727]_ ,
    \new_[1728]_ , \new_[1731]_ , \new_[1734]_ , \new_[1735]_ ,
    \new_[1738]_ , \new_[1741]_ , \new_[1742]_ , \new_[1745]_ ,
    \new_[1748]_ , \new_[1749]_ , \new_[1752]_ , \new_[1755]_ ,
    \new_[1756]_ , \new_[1759]_ , \new_[1762]_ , \new_[1763]_ ,
    \new_[1766]_ , \new_[1769]_ , \new_[1770]_ , \new_[1773]_ ,
    \new_[1776]_ , \new_[1777]_ , \new_[1780]_ , \new_[1783]_ ,
    \new_[1784]_ , \new_[1787]_ , \new_[1790]_ , \new_[1791]_ ,
    \new_[1794]_ , \new_[1797]_ , \new_[1798]_ , \new_[1801]_ ,
    \new_[1804]_ , \new_[1805]_ , \new_[1808]_ , \new_[1811]_ ,
    \new_[1812]_ , \new_[1815]_ , \new_[1818]_ , \new_[1819]_ ,
    \new_[1822]_ , \new_[1825]_ , \new_[1826]_ , \new_[1829]_ ,
    \new_[1832]_ , \new_[1833]_ , \new_[1836]_ , \new_[1840]_ ,
    \new_[1841]_ , \new_[1842]_ , \new_[1845]_ , \new_[1848]_ ,
    \new_[1849]_ , \new_[1852]_ , \new_[1856]_ , \new_[1857]_ ,
    \new_[1858]_ , \new_[1861]_ , \new_[1864]_ , \new_[1865]_ ,
    \new_[1868]_ , \new_[1872]_ , \new_[1873]_ , \new_[1874]_ ,
    \new_[1877]_ , \new_[1880]_ , \new_[1881]_ , \new_[1884]_ ,
    \new_[1888]_ , \new_[1889]_ , \new_[1890]_ , \new_[1893]_ ,
    \new_[1897]_ , \new_[1898]_ , \new_[1899]_ , \new_[1902]_ ,
    \new_[1906]_ , \new_[1907]_ , \new_[1908]_ , \new_[1911]_ ,
    \new_[1915]_ , \new_[1916]_ , \new_[1917]_ , \new_[1920]_ ,
    \new_[1924]_ , \new_[1925]_ , \new_[1926]_ , \new_[1929]_ ,
    \new_[1933]_ , \new_[1934]_ , \new_[1935]_ , \new_[1938]_ ,
    \new_[1942]_ , \new_[1943]_ , \new_[1944]_ , \new_[1947]_ ,
    \new_[1951]_ , \new_[1952]_ , \new_[1953]_ , \new_[1956]_ ,
    \new_[1960]_ , \new_[1961]_ , \new_[1962]_ , \new_[1965]_ ,
    \new_[1969]_ , \new_[1970]_ , \new_[1971]_ , \new_[1974]_ ,
    \new_[1978]_ , \new_[1979]_ , \new_[1980]_ , \new_[1983]_ ,
    \new_[1987]_ , \new_[1988]_ , \new_[1989]_ , \new_[1992]_ ,
    \new_[1996]_ , \new_[1997]_ , \new_[1998]_ , \new_[2001]_ ,
    \new_[2005]_ , \new_[2006]_ , \new_[2007]_ , \new_[2010]_ ,
    \new_[2014]_ , \new_[2015]_ , \new_[2016]_ , \new_[2019]_ ,
    \new_[2023]_ , \new_[2024]_ , \new_[2025]_ , \new_[2028]_ ,
    \new_[2032]_ , \new_[2033]_ , \new_[2034]_ , \new_[2037]_ ,
    \new_[2041]_ , \new_[2042]_ , \new_[2043]_ , \new_[2046]_ ,
    \new_[2050]_ , \new_[2051]_ , \new_[2052]_ , \new_[2055]_ ,
    \new_[2059]_ , \new_[2060]_ , \new_[2061]_ , \new_[2064]_ ,
    \new_[2068]_ , \new_[2069]_ , \new_[2070]_ , \new_[2073]_ ,
    \new_[2077]_ , \new_[2078]_ , \new_[2079]_ , \new_[2082]_ ,
    \new_[2086]_ , \new_[2087]_ , \new_[2088]_ , \new_[2091]_ ,
    \new_[2095]_ , \new_[2096]_ , \new_[2097]_ , \new_[2100]_ ,
    \new_[2104]_ , \new_[2105]_ , \new_[2106]_ , \new_[2109]_ ,
    \new_[2113]_ , \new_[2114]_ , \new_[2115]_ , \new_[2118]_ ,
    \new_[2122]_ , \new_[2123]_ , \new_[2124]_ , \new_[2127]_ ,
    \new_[2131]_ , \new_[2132]_ , \new_[2133]_ , \new_[2136]_ ,
    \new_[2140]_ , \new_[2141]_ , \new_[2142]_ , \new_[2145]_ ,
    \new_[2149]_ , \new_[2150]_ , \new_[2151]_ , \new_[2154]_ ,
    \new_[2158]_ , \new_[2159]_ , \new_[2160]_ , \new_[2163]_ ,
    \new_[2167]_ , \new_[2168]_ , \new_[2169]_ , \new_[2172]_ ,
    \new_[2176]_ , \new_[2177]_ , \new_[2178]_ , \new_[2181]_ ,
    \new_[2185]_ , \new_[2186]_ , \new_[2187]_ , \new_[2190]_ ,
    \new_[2194]_ , \new_[2195]_ , \new_[2196]_ , \new_[2199]_ ,
    \new_[2203]_ , \new_[2204]_ , \new_[2205]_ , \new_[2208]_ ,
    \new_[2212]_ , \new_[2213]_ , \new_[2214]_ , \new_[2217]_ ,
    \new_[2221]_ , \new_[2222]_ , \new_[2223]_ , \new_[2226]_ ,
    \new_[2230]_ , \new_[2231]_ , \new_[2232]_ , \new_[2235]_ ,
    \new_[2239]_ , \new_[2240]_ , \new_[2241]_ , \new_[2244]_ ,
    \new_[2248]_ , \new_[2249]_ , \new_[2250]_ , \new_[2253]_ ,
    \new_[2257]_ , \new_[2258]_ , \new_[2259]_ , \new_[2262]_ ,
    \new_[2266]_ , \new_[2267]_ , \new_[2268]_ , \new_[2271]_ ,
    \new_[2275]_ , \new_[2276]_ , \new_[2277]_ , \new_[2280]_ ,
    \new_[2284]_ , \new_[2285]_ , \new_[2286]_ , \new_[2289]_ ,
    \new_[2293]_ , \new_[2294]_ , \new_[2295]_ , \new_[2298]_ ,
    \new_[2302]_ , \new_[2303]_ , \new_[2304]_ , \new_[2307]_ ,
    \new_[2311]_ , \new_[2312]_ , \new_[2313]_ , \new_[2316]_ ,
    \new_[2320]_ , \new_[2321]_ , \new_[2322]_ , \new_[2325]_ ,
    \new_[2329]_ , \new_[2330]_ , \new_[2331]_ , \new_[2334]_ ,
    \new_[2338]_ , \new_[2339]_ , \new_[2340]_ , \new_[2343]_ ,
    \new_[2347]_ , \new_[2348]_ , \new_[2349]_ , \new_[2352]_ ,
    \new_[2356]_ , \new_[2357]_ , \new_[2358]_ , \new_[2361]_ ,
    \new_[2365]_ , \new_[2366]_ , \new_[2367]_ , \new_[2370]_ ,
    \new_[2374]_ , \new_[2375]_ , \new_[2376]_ , \new_[2379]_ ,
    \new_[2383]_ , \new_[2384]_ , \new_[2385]_ , \new_[2388]_ ,
    \new_[2392]_ , \new_[2393]_ , \new_[2394]_ , \new_[2397]_ ,
    \new_[2401]_ , \new_[2402]_ , \new_[2403]_ , \new_[2406]_ ,
    \new_[2410]_ , \new_[2411]_ , \new_[2412]_ , \new_[2415]_ ,
    \new_[2419]_ , \new_[2420]_ , \new_[2421]_ , \new_[2424]_ ,
    \new_[2428]_ , \new_[2429]_ , \new_[2430]_ , \new_[2433]_ ,
    \new_[2437]_ , \new_[2438]_ , \new_[2439]_ , \new_[2442]_ ,
    \new_[2446]_ , \new_[2447]_ , \new_[2448]_ , \new_[2451]_ ,
    \new_[2455]_ , \new_[2456]_ , \new_[2457]_ , \new_[2460]_ ,
    \new_[2464]_ , \new_[2465]_ , \new_[2466]_ , \new_[2469]_ ,
    \new_[2473]_ , \new_[2474]_ , \new_[2475]_ , \new_[2478]_ ,
    \new_[2482]_ , \new_[2483]_ , \new_[2484]_ , \new_[2487]_ ,
    \new_[2491]_ , \new_[2492]_ , \new_[2493]_ , \new_[2496]_ ,
    \new_[2500]_ , \new_[2501]_ , \new_[2502]_ , \new_[2505]_ ,
    \new_[2509]_ , \new_[2510]_ , \new_[2511]_ , \new_[2514]_ ,
    \new_[2518]_ , \new_[2519]_ , \new_[2520]_ , \new_[2523]_ ,
    \new_[2527]_ , \new_[2528]_ , \new_[2529]_ , \new_[2532]_ ,
    \new_[2536]_ , \new_[2537]_ , \new_[2538]_ , \new_[2541]_ ,
    \new_[2545]_ , \new_[2546]_ , \new_[2547]_ , \new_[2550]_ ,
    \new_[2554]_ , \new_[2555]_ , \new_[2556]_ , \new_[2559]_ ,
    \new_[2563]_ , \new_[2564]_ , \new_[2565]_ , \new_[2568]_ ,
    \new_[2572]_ , \new_[2573]_ , \new_[2574]_ , \new_[2577]_ ,
    \new_[2581]_ , \new_[2582]_ , \new_[2583]_ , \new_[2586]_ ,
    \new_[2590]_ , \new_[2591]_ , \new_[2592]_ , \new_[2595]_ ,
    \new_[2599]_ , \new_[2600]_ , \new_[2601]_ , \new_[2604]_ ,
    \new_[2608]_ , \new_[2609]_ , \new_[2610]_ , \new_[2613]_ ,
    \new_[2617]_ , \new_[2618]_ , \new_[2619]_ , \new_[2622]_ ,
    \new_[2626]_ , \new_[2627]_ , \new_[2628]_ , \new_[2631]_ ,
    \new_[2635]_ , \new_[2636]_ , \new_[2637]_ , \new_[2640]_ ,
    \new_[2644]_ , \new_[2645]_ , \new_[2646]_ , \new_[2649]_ ,
    \new_[2653]_ , \new_[2654]_ , \new_[2655]_ , \new_[2658]_ ,
    \new_[2662]_ , \new_[2663]_ , \new_[2664]_ , \new_[2667]_ ,
    \new_[2671]_ , \new_[2672]_ , \new_[2673]_ , \new_[2676]_ ,
    \new_[2680]_ , \new_[2681]_ , \new_[2682]_ , \new_[2685]_ ,
    \new_[2689]_ , \new_[2690]_ , \new_[2691]_ , \new_[2694]_ ,
    \new_[2698]_ , \new_[2699]_ , \new_[2700]_ , \new_[2703]_ ,
    \new_[2707]_ , \new_[2708]_ , \new_[2709]_ , \new_[2712]_ ,
    \new_[2716]_ , \new_[2717]_ , \new_[2718]_ , \new_[2721]_ ,
    \new_[2725]_ , \new_[2726]_ , \new_[2727]_ , \new_[2730]_ ,
    \new_[2734]_ , \new_[2735]_ , \new_[2736]_ , \new_[2739]_ ,
    \new_[2743]_ , \new_[2744]_ , \new_[2745]_ , \new_[2748]_ ,
    \new_[2752]_ , \new_[2753]_ , \new_[2754]_ , \new_[2757]_ ,
    \new_[2761]_ , \new_[2762]_ , \new_[2763]_ , \new_[2766]_ ,
    \new_[2770]_ , \new_[2771]_ , \new_[2772]_ , \new_[2775]_ ,
    \new_[2779]_ , \new_[2780]_ , \new_[2781]_ , \new_[2784]_ ,
    \new_[2788]_ , \new_[2789]_ , \new_[2790]_ , \new_[2793]_ ,
    \new_[2797]_ , \new_[2798]_ , \new_[2799]_ , \new_[2802]_ ,
    \new_[2806]_ , \new_[2807]_ , \new_[2808]_ , \new_[2811]_ ,
    \new_[2815]_ , \new_[2816]_ , \new_[2817]_ , \new_[2820]_ ,
    \new_[2824]_ , \new_[2825]_ , \new_[2826]_ , \new_[2829]_ ,
    \new_[2833]_ , \new_[2834]_ , \new_[2835]_ , \new_[2838]_ ,
    \new_[2842]_ , \new_[2843]_ , \new_[2844]_ , \new_[2847]_ ,
    \new_[2851]_ , \new_[2852]_ , \new_[2853]_ , \new_[2856]_ ,
    \new_[2860]_ , \new_[2861]_ , \new_[2862]_ , \new_[2865]_ ,
    \new_[2869]_ , \new_[2870]_ , \new_[2871]_ , \new_[2874]_ ,
    \new_[2878]_ , \new_[2879]_ , \new_[2880]_ , \new_[2883]_ ,
    \new_[2887]_ , \new_[2888]_ , \new_[2889]_ , \new_[2892]_ ,
    \new_[2896]_ , \new_[2897]_ , \new_[2898]_ , \new_[2901]_ ,
    \new_[2905]_ , \new_[2906]_ , \new_[2907]_ , \new_[2910]_ ,
    \new_[2914]_ , \new_[2915]_ , \new_[2916]_ , \new_[2919]_ ,
    \new_[2923]_ , \new_[2924]_ , \new_[2925]_ , \new_[2928]_ ,
    \new_[2932]_ , \new_[2933]_ , \new_[2934]_ , \new_[2937]_ ,
    \new_[2941]_ , \new_[2942]_ , \new_[2943]_ , \new_[2946]_ ,
    \new_[2950]_ , \new_[2951]_ , \new_[2952]_ , \new_[2955]_ ,
    \new_[2959]_ , \new_[2960]_ , \new_[2961]_ , \new_[2964]_ ,
    \new_[2968]_ , \new_[2969]_ , \new_[2970]_ , \new_[2973]_ ,
    \new_[2977]_ , \new_[2978]_ , \new_[2979]_ , \new_[2982]_ ,
    \new_[2986]_ , \new_[2987]_ , \new_[2988]_ , \new_[2991]_ ,
    \new_[2995]_ , \new_[2996]_ , \new_[2997]_ , \new_[3000]_ ,
    \new_[3004]_ , \new_[3005]_ , \new_[3006]_ , \new_[3009]_ ,
    \new_[3013]_ , \new_[3014]_ , \new_[3015]_ , \new_[3018]_ ,
    \new_[3022]_ , \new_[3023]_ , \new_[3024]_ , \new_[3027]_ ,
    \new_[3031]_ , \new_[3032]_ , \new_[3033]_ , \new_[3036]_ ,
    \new_[3040]_ , \new_[3041]_ , \new_[3042]_ , \new_[3045]_ ,
    \new_[3049]_ , \new_[3050]_ , \new_[3051]_ , \new_[3054]_ ,
    \new_[3058]_ , \new_[3059]_ , \new_[3060]_ , \new_[3063]_ ,
    \new_[3067]_ , \new_[3068]_ , \new_[3069]_ , \new_[3072]_ ,
    \new_[3076]_ , \new_[3077]_ , \new_[3078]_ , \new_[3081]_ ,
    \new_[3085]_ , \new_[3086]_ , \new_[3087]_ , \new_[3090]_ ,
    \new_[3094]_ , \new_[3095]_ , \new_[3096]_ , \new_[3099]_ ,
    \new_[3103]_ , \new_[3104]_ , \new_[3105]_ , \new_[3108]_ ,
    \new_[3112]_ , \new_[3113]_ , \new_[3114]_ , \new_[3117]_ ,
    \new_[3121]_ , \new_[3122]_ , \new_[3123]_ , \new_[3126]_ ,
    \new_[3130]_ , \new_[3131]_ , \new_[3132]_ , \new_[3135]_ ,
    \new_[3139]_ , \new_[3140]_ , \new_[3141]_ , \new_[3144]_ ,
    \new_[3148]_ , \new_[3149]_ , \new_[3150]_ , \new_[3153]_ ,
    \new_[3157]_ , \new_[3158]_ , \new_[3159]_ , \new_[3162]_ ,
    \new_[3166]_ , \new_[3167]_ , \new_[3168]_ , \new_[3171]_ ,
    \new_[3175]_ , \new_[3176]_ , \new_[3177]_ , \new_[3180]_ ,
    \new_[3184]_ , \new_[3185]_ , \new_[3186]_ , \new_[3189]_ ,
    \new_[3193]_ , \new_[3194]_ , \new_[3195]_ , \new_[3199]_ ,
    \new_[3200]_ , \new_[3204]_ , \new_[3205]_ , \new_[3206]_ ,
    \new_[3209]_ , \new_[3213]_ , \new_[3214]_ , \new_[3215]_ ,
    \new_[3219]_ , \new_[3220]_ , \new_[3224]_ , \new_[3225]_ ,
    \new_[3226]_ , \new_[3229]_ , \new_[3233]_ , \new_[3234]_ ,
    \new_[3235]_ , \new_[3239]_ , \new_[3240]_ , \new_[3244]_ ,
    \new_[3245]_ , \new_[3246]_ , \new_[3249]_ , \new_[3253]_ ,
    \new_[3254]_ , \new_[3255]_ , \new_[3259]_ , \new_[3260]_ ,
    \new_[3264]_ , \new_[3265]_ , \new_[3266]_ , \new_[3269]_ ,
    \new_[3273]_ , \new_[3274]_ , \new_[3275]_ , \new_[3279]_ ,
    \new_[3280]_ , \new_[3284]_ , \new_[3285]_ , \new_[3286]_ ,
    \new_[3289]_ , \new_[3293]_ , \new_[3294]_ , \new_[3295]_ ,
    \new_[3299]_ , \new_[3300]_ , \new_[3304]_ , \new_[3305]_ ,
    \new_[3306]_ , \new_[3309]_ , \new_[3313]_ , \new_[3314]_ ,
    \new_[3315]_ , \new_[3319]_ , \new_[3320]_ , \new_[3324]_ ,
    \new_[3325]_ , \new_[3326]_ , \new_[3329]_ , \new_[3333]_ ,
    \new_[3334]_ , \new_[3335]_ , \new_[3339]_ , \new_[3340]_ ,
    \new_[3344]_ , \new_[3345]_ , \new_[3346]_ , \new_[3349]_ ,
    \new_[3353]_ , \new_[3354]_ , \new_[3355]_ , \new_[3359]_ ,
    \new_[3360]_ , \new_[3364]_ , \new_[3365]_ , \new_[3366]_ ,
    \new_[3369]_ , \new_[3373]_ , \new_[3374]_ , \new_[3375]_ ,
    \new_[3379]_ , \new_[3380]_ , \new_[3384]_ , \new_[3385]_ ,
    \new_[3386]_ , \new_[3389]_ , \new_[3393]_ , \new_[3394]_ ,
    \new_[3395]_ , \new_[3399]_ , \new_[3400]_ , \new_[3404]_ ,
    \new_[3405]_ , \new_[3406]_ , \new_[3409]_ , \new_[3413]_ ,
    \new_[3414]_ , \new_[3415]_ , \new_[3419]_ , \new_[3420]_ ,
    \new_[3424]_ , \new_[3425]_ , \new_[3426]_ , \new_[3429]_ ,
    \new_[3433]_ , \new_[3434]_ , \new_[3435]_ , \new_[3439]_ ,
    \new_[3440]_ , \new_[3444]_ , \new_[3445]_ , \new_[3446]_ ,
    \new_[3449]_ , \new_[3453]_ , \new_[3454]_ , \new_[3455]_ ,
    \new_[3459]_ , \new_[3460]_ , \new_[3464]_ , \new_[3465]_ ,
    \new_[3466]_ , \new_[3469]_ , \new_[3473]_ , \new_[3474]_ ,
    \new_[3475]_ , \new_[3479]_ , \new_[3480]_ , \new_[3484]_ ,
    \new_[3485]_ , \new_[3486]_ , \new_[3489]_ , \new_[3493]_ ,
    \new_[3494]_ , \new_[3495]_ , \new_[3499]_ , \new_[3500]_ ,
    \new_[3504]_ , \new_[3505]_ , \new_[3506]_ , \new_[3509]_ ,
    \new_[3513]_ , \new_[3514]_ , \new_[3515]_ , \new_[3519]_ ,
    \new_[3520]_ , \new_[3524]_ , \new_[3525]_ , \new_[3526]_ ,
    \new_[3529]_ , \new_[3533]_ , \new_[3534]_ , \new_[3535]_ ,
    \new_[3539]_ , \new_[3540]_ , \new_[3544]_ , \new_[3545]_ ,
    \new_[3546]_ , \new_[3549]_ , \new_[3553]_ , \new_[3554]_ ,
    \new_[3555]_ , \new_[3559]_ , \new_[3560]_ , \new_[3564]_ ,
    \new_[3565]_ , \new_[3566]_ , \new_[3569]_ , \new_[3573]_ ,
    \new_[3574]_ , \new_[3575]_ , \new_[3579]_ , \new_[3580]_ ,
    \new_[3584]_ , \new_[3585]_ , \new_[3586]_ , \new_[3589]_ ,
    \new_[3593]_ , \new_[3594]_ , \new_[3595]_ , \new_[3599]_ ,
    \new_[3600]_ , \new_[3604]_ , \new_[3605]_ , \new_[3606]_ ,
    \new_[3609]_ , \new_[3613]_ , \new_[3614]_ , \new_[3615]_ ,
    \new_[3619]_ , \new_[3620]_ , \new_[3624]_ , \new_[3625]_ ,
    \new_[3626]_ , \new_[3629]_ , \new_[3633]_ , \new_[3634]_ ,
    \new_[3635]_ , \new_[3639]_ , \new_[3640]_ , \new_[3644]_ ,
    \new_[3645]_ , \new_[3646]_ , \new_[3649]_ , \new_[3653]_ ,
    \new_[3654]_ , \new_[3655]_ , \new_[3659]_ , \new_[3660]_ ,
    \new_[3664]_ , \new_[3665]_ , \new_[3666]_ , \new_[3670]_ ,
    \new_[3671]_ , \new_[3675]_ , \new_[3676]_ , \new_[3677]_ ,
    \new_[3681]_ , \new_[3682]_ , \new_[3686]_ , \new_[3687]_ ,
    \new_[3688]_ , \new_[3692]_ , \new_[3693]_ , \new_[3697]_ ,
    \new_[3698]_ , \new_[3699]_ , \new_[3703]_ , \new_[3704]_ ,
    \new_[3708]_ , \new_[3709]_ , \new_[3710]_ , \new_[3714]_ ,
    \new_[3715]_ , \new_[3719]_ , \new_[3720]_ , \new_[3721]_ ,
    \new_[3725]_ , \new_[3726]_ , \new_[3730]_ , \new_[3731]_ ,
    \new_[3732]_ , \new_[3736]_ , \new_[3737]_ , \new_[3741]_ ,
    \new_[3742]_ , \new_[3743]_ , \new_[3747]_ , \new_[3748]_ ,
    \new_[3752]_ , \new_[3753]_ , \new_[3754]_ , \new_[3758]_ ,
    \new_[3759]_ , \new_[3763]_ , \new_[3764]_ , \new_[3765]_ ,
    \new_[3769]_ , \new_[3770]_ , \new_[3774]_ , \new_[3775]_ ,
    \new_[3776]_ , \new_[3780]_ , \new_[3781]_ , \new_[3785]_ ,
    \new_[3786]_ , \new_[3787]_ , \new_[3791]_ , \new_[3792]_ ,
    \new_[3796]_ , \new_[3797]_ , \new_[3798]_ , \new_[3802]_ ,
    \new_[3803]_ , \new_[3807]_ , \new_[3808]_ , \new_[3809]_ ,
    \new_[3813]_ , \new_[3814]_ , \new_[3818]_ , \new_[3819]_ ,
    \new_[3820]_ , \new_[3824]_ , \new_[3825]_ , \new_[3829]_ ,
    \new_[3830]_ , \new_[3831]_ , \new_[3835]_ , \new_[3836]_ ,
    \new_[3840]_ , \new_[3841]_ , \new_[3842]_ , \new_[3846]_ ,
    \new_[3847]_ , \new_[3851]_ , \new_[3852]_ , \new_[3853]_ ,
    \new_[3857]_ , \new_[3858]_ , \new_[3862]_ , \new_[3863]_ ,
    \new_[3864]_ , \new_[3868]_ , \new_[3869]_ , \new_[3873]_ ,
    \new_[3874]_ , \new_[3875]_ , \new_[3879]_ , \new_[3880]_ ,
    \new_[3884]_ , \new_[3885]_ , \new_[3886]_ , \new_[3890]_ ,
    \new_[3891]_ , \new_[3895]_ , \new_[3896]_ , \new_[3897]_ ,
    \new_[3901]_ , \new_[3902]_ , \new_[3906]_ , \new_[3907]_ ,
    \new_[3908]_ , \new_[3912]_ , \new_[3913]_ , \new_[3917]_ ,
    \new_[3918]_ , \new_[3919]_ , \new_[3923]_ , \new_[3924]_ ,
    \new_[3928]_ , \new_[3929]_ , \new_[3930]_ , \new_[3934]_ ,
    \new_[3935]_ , \new_[3939]_ , \new_[3940]_ , \new_[3941]_ ,
    \new_[3945]_ , \new_[3946]_ , \new_[3950]_ , \new_[3951]_ ,
    \new_[3952]_ , \new_[3956]_ , \new_[3957]_ , \new_[3961]_ ,
    \new_[3962]_ , \new_[3963]_ , \new_[3967]_ , \new_[3968]_ ,
    \new_[3972]_ , \new_[3973]_ , \new_[3974]_ , \new_[3978]_ ,
    \new_[3979]_ , \new_[3983]_ , \new_[3984]_ , \new_[3985]_ ,
    \new_[3989]_ , \new_[3990]_ , \new_[3994]_ , \new_[3995]_ ,
    \new_[3996]_ , \new_[4000]_ , \new_[4001]_ , \new_[4005]_ ,
    \new_[4006]_ , \new_[4007]_ , \new_[4011]_ , \new_[4012]_ ,
    \new_[4016]_ , \new_[4017]_ , \new_[4018]_ , \new_[4022]_ ,
    \new_[4023]_ , \new_[4027]_ , \new_[4028]_ , \new_[4029]_ ,
    \new_[4033]_ , \new_[4034]_ , \new_[4038]_ , \new_[4039]_ ,
    \new_[4040]_ , \new_[4044]_ , \new_[4045]_ , \new_[4049]_ ,
    \new_[4050]_ , \new_[4051]_ , \new_[4055]_ , \new_[4056]_ ,
    \new_[4060]_ , \new_[4061]_ , \new_[4062]_ , \new_[4066]_ ,
    \new_[4067]_ , \new_[4071]_ , \new_[4072]_ , \new_[4073]_ ,
    \new_[4077]_ , \new_[4078]_ , \new_[4082]_ , \new_[4083]_ ,
    \new_[4084]_ , \new_[4088]_ , \new_[4089]_ , \new_[4093]_ ,
    \new_[4094]_ , \new_[4095]_ , \new_[4099]_ , \new_[4100]_ ,
    \new_[4104]_ , \new_[4105]_ , \new_[4106]_ , \new_[4110]_ ,
    \new_[4111]_ , \new_[4115]_ , \new_[4116]_ , \new_[4117]_ ,
    \new_[4121]_ , \new_[4122]_ , \new_[4126]_ , \new_[4127]_ ,
    \new_[4128]_ , \new_[4132]_ , \new_[4133]_ , \new_[4137]_ ,
    \new_[4138]_ , \new_[4139]_ , \new_[4143]_ , \new_[4144]_ ,
    \new_[4148]_ , \new_[4149]_ , \new_[4150]_ , \new_[4154]_ ,
    \new_[4155]_ , \new_[4159]_ , \new_[4160]_ , \new_[4161]_ ,
    \new_[4165]_ , \new_[4166]_ , \new_[4170]_ , \new_[4171]_ ,
    \new_[4172]_ , \new_[4176]_ , \new_[4177]_ , \new_[4181]_ ,
    \new_[4182]_ , \new_[4183]_ , \new_[4187]_ , \new_[4188]_ ,
    \new_[4192]_ , \new_[4193]_ , \new_[4194]_ , \new_[4198]_ ,
    \new_[4199]_ , \new_[4203]_ , \new_[4204]_ , \new_[4205]_ ,
    \new_[4209]_ , \new_[4210]_ , \new_[4214]_ , \new_[4215]_ ,
    \new_[4216]_ , \new_[4220]_ , \new_[4221]_ , \new_[4225]_ ,
    \new_[4226]_ , \new_[4227]_ , \new_[4231]_ , \new_[4232]_ ,
    \new_[4236]_ , \new_[4237]_ , \new_[4238]_ , \new_[4242]_ ,
    \new_[4243]_ , \new_[4247]_ , \new_[4248]_ , \new_[4249]_ ,
    \new_[4253]_ , \new_[4254]_ , \new_[4258]_ , \new_[4259]_ ,
    \new_[4260]_ , \new_[4264]_ , \new_[4265]_ , \new_[4269]_ ,
    \new_[4270]_ , \new_[4271]_ , \new_[4275]_ , \new_[4276]_ ,
    \new_[4280]_ , \new_[4281]_ , \new_[4282]_ , \new_[4286]_ ,
    \new_[4287]_ , \new_[4291]_ , \new_[4292]_ , \new_[4293]_ ,
    \new_[4297]_ , \new_[4298]_ , \new_[4302]_ , \new_[4303]_ ,
    \new_[4304]_ , \new_[4308]_ , \new_[4309]_ , \new_[4313]_ ,
    \new_[4314]_ , \new_[4315]_ , \new_[4319]_ , \new_[4320]_ ,
    \new_[4324]_ , \new_[4325]_ , \new_[4326]_ , \new_[4330]_ ,
    \new_[4331]_ , \new_[4335]_ , \new_[4336]_ , \new_[4337]_ ,
    \new_[4341]_ , \new_[4342]_ , \new_[4346]_ , \new_[4347]_ ,
    \new_[4348]_ , \new_[4352]_ , \new_[4353]_ , \new_[4357]_ ,
    \new_[4358]_ , \new_[4359]_ , \new_[4363]_ , \new_[4364]_ ,
    \new_[4368]_ , \new_[4369]_ , \new_[4370]_ , \new_[4374]_ ,
    \new_[4375]_ , \new_[4379]_ , \new_[4380]_ , \new_[4381]_ ,
    \new_[4385]_ , \new_[4386]_ , \new_[4390]_ , \new_[4391]_ ,
    \new_[4392]_ , \new_[4396]_ , \new_[4397]_ , \new_[4401]_ ,
    \new_[4402]_ , \new_[4403]_ , \new_[4407]_ , \new_[4408]_ ,
    \new_[4412]_ , \new_[4413]_ , \new_[4414]_ , \new_[4418]_ ,
    \new_[4419]_ , \new_[4423]_ , \new_[4424]_ , \new_[4425]_ ,
    \new_[4429]_ , \new_[4430]_ , \new_[4434]_ , \new_[4435]_ ,
    \new_[4436]_ , \new_[4440]_ , \new_[4441]_ , \new_[4445]_ ,
    \new_[4446]_ , \new_[4447]_ , \new_[4451]_ , \new_[4452]_ ,
    \new_[4456]_ , \new_[4457]_ , \new_[4458]_ , \new_[4462]_ ,
    \new_[4463]_ , \new_[4467]_ , \new_[4468]_ , \new_[4469]_ ,
    \new_[4473]_ , \new_[4474]_ , \new_[4478]_ , \new_[4479]_ ,
    \new_[4480]_ , \new_[4484]_ , \new_[4485]_ , \new_[4489]_ ,
    \new_[4490]_ , \new_[4491]_ , \new_[4495]_ , \new_[4496]_ ,
    \new_[4500]_ , \new_[4501]_ , \new_[4502]_ , \new_[4506]_ ,
    \new_[4507]_ , \new_[4511]_ , \new_[4512]_ , \new_[4513]_ ,
    \new_[4517]_ , \new_[4518]_ , \new_[4522]_ , \new_[4523]_ ,
    \new_[4524]_ , \new_[4528]_ , \new_[4529]_ , \new_[4533]_ ,
    \new_[4534]_ , \new_[4535]_ , \new_[4539]_ , \new_[4540]_ ,
    \new_[4544]_ , \new_[4545]_ , \new_[4546]_ , \new_[4550]_ ,
    \new_[4551]_ , \new_[4555]_ , \new_[4556]_ , \new_[4557]_ ,
    \new_[4561]_ , \new_[4562]_ , \new_[4566]_ , \new_[4567]_ ,
    \new_[4568]_ , \new_[4572]_ , \new_[4573]_ , \new_[4577]_ ,
    \new_[4578]_ , \new_[4579]_ , \new_[4583]_ , \new_[4584]_ ,
    \new_[4588]_ , \new_[4589]_ , \new_[4590]_ , \new_[4594]_ ,
    \new_[4595]_ , \new_[4599]_ , \new_[4600]_ , \new_[4601]_ ,
    \new_[4605]_ , \new_[4606]_ , \new_[4610]_ , \new_[4611]_ ,
    \new_[4612]_ , \new_[4616]_ , \new_[4617]_ , \new_[4621]_ ,
    \new_[4622]_ , \new_[4623]_ , \new_[4627]_ , \new_[4628]_ ,
    \new_[4632]_ , \new_[4633]_ , \new_[4634]_ , \new_[4638]_ ,
    \new_[4639]_ , \new_[4643]_ , \new_[4644]_ , \new_[4645]_ ,
    \new_[4649]_ , \new_[4650]_ , \new_[4654]_ , \new_[4655]_ ,
    \new_[4656]_ , \new_[4660]_ , \new_[4661]_ , \new_[4665]_ ,
    \new_[4666]_ , \new_[4667]_ , \new_[4671]_ , \new_[4672]_ ,
    \new_[4676]_ , \new_[4677]_ , \new_[4678]_ , \new_[4682]_ ,
    \new_[4683]_ , \new_[4687]_ , \new_[4688]_ , \new_[4689]_ ,
    \new_[4693]_ , \new_[4694]_ , \new_[4698]_ , \new_[4699]_ ,
    \new_[4700]_ , \new_[4704]_ , \new_[4705]_ , \new_[4709]_ ,
    \new_[4710]_ , \new_[4711]_ , \new_[4715]_ , \new_[4716]_ ,
    \new_[4720]_ , \new_[4721]_ , \new_[4722]_ , \new_[4726]_ ,
    \new_[4727]_ , \new_[4731]_ , \new_[4732]_ , \new_[4733]_ ,
    \new_[4737]_ , \new_[4738]_ , \new_[4742]_ , \new_[4743]_ ,
    \new_[4744]_ , \new_[4748]_ , \new_[4749]_ , \new_[4753]_ ,
    \new_[4754]_ , \new_[4755]_ , \new_[4759]_ , \new_[4760]_ ,
    \new_[4764]_ , \new_[4765]_ , \new_[4766]_ , \new_[4770]_ ,
    \new_[4771]_ , \new_[4775]_ , \new_[4776]_ , \new_[4777]_ ,
    \new_[4781]_ , \new_[4782]_ , \new_[4786]_ , \new_[4787]_ ,
    \new_[4788]_ , \new_[4792]_ , \new_[4793]_ , \new_[4797]_ ,
    \new_[4798]_ , \new_[4799]_ , \new_[4803]_ , \new_[4804]_ ,
    \new_[4808]_ , \new_[4809]_ , \new_[4810]_ , \new_[4814]_ ,
    \new_[4815]_ , \new_[4819]_ , \new_[4820]_ , \new_[4821]_ ,
    \new_[4825]_ , \new_[4826]_ , \new_[4830]_ , \new_[4831]_ ,
    \new_[4832]_ , \new_[4836]_ , \new_[4837]_ , \new_[4841]_ ,
    \new_[4842]_ , \new_[4843]_ , \new_[4847]_ , \new_[4848]_ ,
    \new_[4852]_ , \new_[4853]_ , \new_[4854]_ , \new_[4858]_ ,
    \new_[4859]_ , \new_[4863]_ , \new_[4864]_ , \new_[4865]_ ,
    \new_[4869]_ , \new_[4870]_ , \new_[4874]_ , \new_[4875]_ ,
    \new_[4876]_ , \new_[4880]_ , \new_[4881]_ , \new_[4885]_ ,
    \new_[4886]_ , \new_[4887]_ , \new_[4891]_ , \new_[4892]_ ,
    \new_[4896]_ , \new_[4897]_ , \new_[4898]_ , \new_[4902]_ ,
    \new_[4903]_ , \new_[4907]_ , \new_[4908]_ , \new_[4909]_ ,
    \new_[4913]_ , \new_[4914]_ , \new_[4918]_ , \new_[4919]_ ,
    \new_[4920]_ , \new_[4924]_ , \new_[4925]_ , \new_[4929]_ ,
    \new_[4930]_ , \new_[4931]_ , \new_[4935]_ , \new_[4936]_ ,
    \new_[4940]_ , \new_[4941]_ , \new_[4942]_ , \new_[4946]_ ,
    \new_[4947]_ , \new_[4951]_ , \new_[4952]_ , \new_[4953]_ ,
    \new_[4957]_ , \new_[4958]_ , \new_[4962]_ , \new_[4963]_ ,
    \new_[4964]_ , \new_[4968]_ , \new_[4969]_ , \new_[4973]_ ,
    \new_[4974]_ , \new_[4975]_ , \new_[4979]_ , \new_[4980]_ ,
    \new_[4984]_ , \new_[4985]_ , \new_[4986]_ , \new_[4990]_ ,
    \new_[4991]_ , \new_[4995]_ , \new_[4996]_ , \new_[4997]_ ,
    \new_[5001]_ , \new_[5002]_ , \new_[5006]_ , \new_[5007]_ ,
    \new_[5008]_ , \new_[5012]_ , \new_[5013]_ , \new_[5017]_ ,
    \new_[5018]_ , \new_[5019]_ , \new_[5023]_ , \new_[5024]_ ,
    \new_[5028]_ , \new_[5029]_ , \new_[5030]_ , \new_[5034]_ ,
    \new_[5035]_ , \new_[5039]_ , \new_[5040]_ , \new_[5041]_ ,
    \new_[5045]_ , \new_[5046]_ , \new_[5050]_ , \new_[5051]_ ,
    \new_[5052]_ , \new_[5056]_ , \new_[5057]_ , \new_[5061]_ ,
    \new_[5062]_ , \new_[5063]_ , \new_[5067]_ , \new_[5068]_ ,
    \new_[5072]_ , \new_[5073]_ , \new_[5074]_ , \new_[5078]_ ,
    \new_[5079]_ , \new_[5083]_ , \new_[5084]_ , \new_[5085]_ ,
    \new_[5089]_ , \new_[5090]_ , \new_[5094]_ , \new_[5095]_ ,
    \new_[5096]_ , \new_[5100]_ , \new_[5101]_ , \new_[5105]_ ,
    \new_[5106]_ , \new_[5107]_ , \new_[5111]_ , \new_[5112]_ ,
    \new_[5116]_ , \new_[5117]_ , \new_[5118]_ , \new_[5122]_ ,
    \new_[5123]_ , \new_[5127]_ , \new_[5128]_ , \new_[5129]_ ,
    \new_[5133]_ , \new_[5134]_ , \new_[5138]_ , \new_[5139]_ ,
    \new_[5140]_ , \new_[5144]_ , \new_[5145]_ , \new_[5149]_ ,
    \new_[5150]_ , \new_[5151]_ , \new_[5155]_ , \new_[5156]_ ,
    \new_[5160]_ , \new_[5161]_ , \new_[5162]_ , \new_[5166]_ ,
    \new_[5167]_ , \new_[5171]_ , \new_[5172]_ , \new_[5173]_ ,
    \new_[5177]_ , \new_[5178]_ , \new_[5182]_ , \new_[5183]_ ,
    \new_[5184]_ , \new_[5188]_ , \new_[5189]_ , \new_[5193]_ ,
    \new_[5194]_ , \new_[5195]_ , \new_[5199]_ , \new_[5200]_ ,
    \new_[5204]_ , \new_[5205]_ , \new_[5206]_ , \new_[5210]_ ,
    \new_[5211]_ , \new_[5215]_ , \new_[5216]_ , \new_[5217]_ ,
    \new_[5221]_ , \new_[5222]_ , \new_[5226]_ , \new_[5227]_ ,
    \new_[5228]_ , \new_[5232]_ , \new_[5233]_ , \new_[5237]_ ,
    \new_[5238]_ , \new_[5239]_ , \new_[5243]_ , \new_[5244]_ ,
    \new_[5248]_ , \new_[5249]_ , \new_[5250]_ , \new_[5254]_ ,
    \new_[5255]_ , \new_[5259]_ , \new_[5260]_ , \new_[5261]_ ,
    \new_[5265]_ , \new_[5266]_ , \new_[5270]_ , \new_[5271]_ ,
    \new_[5272]_ , \new_[5276]_ , \new_[5277]_ , \new_[5281]_ ,
    \new_[5282]_ , \new_[5283]_ , \new_[5287]_ , \new_[5288]_ ,
    \new_[5292]_ , \new_[5293]_ , \new_[5294]_ , \new_[5298]_ ,
    \new_[5299]_ , \new_[5303]_ , \new_[5304]_ , \new_[5305]_ ,
    \new_[5309]_ , \new_[5310]_ , \new_[5314]_ , \new_[5315]_ ,
    \new_[5316]_ , \new_[5320]_ , \new_[5321]_ , \new_[5325]_ ,
    \new_[5326]_ , \new_[5327]_ , \new_[5331]_ , \new_[5332]_ ,
    \new_[5336]_ , \new_[5337]_ , \new_[5338]_ , \new_[5342]_ ,
    \new_[5343]_ , \new_[5347]_ , \new_[5348]_ , \new_[5349]_ ,
    \new_[5353]_ , \new_[5354]_ , \new_[5358]_ , \new_[5359]_ ,
    \new_[5360]_ , \new_[5364]_ , \new_[5365]_ , \new_[5369]_ ,
    \new_[5370]_ , \new_[5371]_ , \new_[5375]_ , \new_[5376]_ ,
    \new_[5380]_ , \new_[5381]_ , \new_[5382]_ , \new_[5386]_ ,
    \new_[5387]_ , \new_[5391]_ , \new_[5392]_ , \new_[5393]_ ,
    \new_[5397]_ , \new_[5398]_ , \new_[5402]_ , \new_[5403]_ ,
    \new_[5404]_ , \new_[5408]_ , \new_[5409]_ , \new_[5413]_ ,
    \new_[5414]_ , \new_[5415]_ , \new_[5419]_ , \new_[5420]_ ,
    \new_[5424]_ , \new_[5425]_ , \new_[5426]_ , \new_[5430]_ ,
    \new_[5431]_ , \new_[5435]_ , \new_[5436]_ , \new_[5437]_ ,
    \new_[5441]_ , \new_[5442]_ , \new_[5446]_ , \new_[5447]_ ,
    \new_[5448]_ , \new_[5452]_ , \new_[5453]_ , \new_[5457]_ ,
    \new_[5458]_ , \new_[5459]_ , \new_[5463]_ , \new_[5464]_ ,
    \new_[5468]_ , \new_[5469]_ , \new_[5470]_ , \new_[5474]_ ,
    \new_[5475]_ , \new_[5479]_ , \new_[5480]_ , \new_[5481]_ ,
    \new_[5485]_ , \new_[5486]_ , \new_[5490]_ , \new_[5491]_ ,
    \new_[5492]_ , \new_[5496]_ , \new_[5497]_ , \new_[5501]_ ,
    \new_[5502]_ , \new_[5503]_ , \new_[5507]_ , \new_[5508]_ ,
    \new_[5512]_ , \new_[5513]_ , \new_[5514]_ , \new_[5518]_ ,
    \new_[5519]_ , \new_[5523]_ , \new_[5524]_ , \new_[5525]_ ,
    \new_[5529]_ , \new_[5530]_ , \new_[5534]_ , \new_[5535]_ ,
    \new_[5536]_ , \new_[5540]_ , \new_[5541]_ , \new_[5545]_ ,
    \new_[5546]_ , \new_[5547]_ , \new_[5551]_ , \new_[5552]_ ,
    \new_[5556]_ , \new_[5557]_ , \new_[5558]_ , \new_[5562]_ ,
    \new_[5563]_ , \new_[5567]_ , \new_[5568]_ , \new_[5569]_ ,
    \new_[5573]_ , \new_[5574]_ , \new_[5578]_ , \new_[5579]_ ,
    \new_[5580]_ , \new_[5584]_ , \new_[5585]_ , \new_[5589]_ ,
    \new_[5590]_ , \new_[5591]_ , \new_[5595]_ , \new_[5596]_ ,
    \new_[5600]_ , \new_[5601]_ , \new_[5602]_ , \new_[5606]_ ,
    \new_[5607]_ , \new_[5611]_ , \new_[5612]_ , \new_[5613]_ ,
    \new_[5617]_ , \new_[5618]_ , \new_[5622]_ , \new_[5623]_ ,
    \new_[5624]_ , \new_[5628]_ , \new_[5629]_ , \new_[5633]_ ,
    \new_[5634]_ , \new_[5635]_ , \new_[5639]_ , \new_[5640]_ ,
    \new_[5644]_ , \new_[5645]_ , \new_[5646]_ , \new_[5650]_ ,
    \new_[5651]_ , \new_[5655]_ , \new_[5656]_ , \new_[5657]_ ,
    \new_[5661]_ , \new_[5662]_ , \new_[5666]_ , \new_[5667]_ ,
    \new_[5668]_ , \new_[5672]_ , \new_[5673]_ , \new_[5677]_ ,
    \new_[5678]_ , \new_[5679]_ , \new_[5683]_ , \new_[5684]_ ,
    \new_[5688]_ , \new_[5689]_ , \new_[5690]_ , \new_[5694]_ ,
    \new_[5695]_ , \new_[5699]_ , \new_[5700]_ , \new_[5701]_ ,
    \new_[5705]_ , \new_[5706]_ , \new_[5710]_ , \new_[5711]_ ,
    \new_[5712]_ , \new_[5716]_ , \new_[5717]_ , \new_[5721]_ ,
    \new_[5722]_ , \new_[5723]_ , \new_[5727]_ , \new_[5728]_ ,
    \new_[5732]_ , \new_[5733]_ , \new_[5734]_ , \new_[5738]_ ,
    \new_[5739]_ , \new_[5743]_ , \new_[5744]_ , \new_[5745]_ ,
    \new_[5749]_ , \new_[5750]_ , \new_[5754]_ , \new_[5755]_ ,
    \new_[5756]_ , \new_[5760]_ , \new_[5761]_ , \new_[5765]_ ,
    \new_[5766]_ , \new_[5767]_ , \new_[5771]_ , \new_[5772]_ ,
    \new_[5776]_ , \new_[5777]_ , \new_[5778]_ , \new_[5782]_ ,
    \new_[5783]_ , \new_[5787]_ , \new_[5788]_ , \new_[5789]_ ,
    \new_[5793]_ , \new_[5794]_ , \new_[5798]_ , \new_[5799]_ ,
    \new_[5800]_ , \new_[5804]_ , \new_[5805]_ , \new_[5809]_ ,
    \new_[5810]_ , \new_[5811]_ , \new_[5815]_ , \new_[5816]_ ,
    \new_[5820]_ , \new_[5821]_ , \new_[5822]_ , \new_[5826]_ ,
    \new_[5827]_ , \new_[5831]_ , \new_[5832]_ , \new_[5833]_ ,
    \new_[5837]_ , \new_[5838]_ , \new_[5842]_ , \new_[5843]_ ,
    \new_[5844]_ , \new_[5848]_ , \new_[5849]_ , \new_[5853]_ ,
    \new_[5854]_ , \new_[5855]_ , \new_[5859]_ , \new_[5860]_ ,
    \new_[5864]_ , \new_[5865]_ , \new_[5866]_ , \new_[5870]_ ,
    \new_[5871]_ , \new_[5875]_ , \new_[5876]_ , \new_[5877]_ ,
    \new_[5881]_ , \new_[5882]_ , \new_[5886]_ , \new_[5887]_ ,
    \new_[5888]_ , \new_[5892]_ , \new_[5893]_ , \new_[5897]_ ,
    \new_[5898]_ , \new_[5899]_ , \new_[5903]_ , \new_[5904]_ ,
    \new_[5908]_ , \new_[5909]_ , \new_[5910]_ , \new_[5914]_ ,
    \new_[5915]_ , \new_[5919]_ , \new_[5920]_ , \new_[5921]_ ,
    \new_[5925]_ , \new_[5926]_ , \new_[5930]_ , \new_[5931]_ ,
    \new_[5932]_ , \new_[5936]_ , \new_[5937]_ , \new_[5941]_ ,
    \new_[5942]_ , \new_[5943]_ , \new_[5947]_ , \new_[5948]_ ,
    \new_[5952]_ , \new_[5953]_ , \new_[5954]_ , \new_[5958]_ ,
    \new_[5959]_ , \new_[5963]_ , \new_[5964]_ , \new_[5965]_ ,
    \new_[5969]_ , \new_[5970]_ , \new_[5974]_ , \new_[5975]_ ,
    \new_[5976]_ , \new_[5980]_ , \new_[5981]_ , \new_[5985]_ ,
    \new_[5986]_ , \new_[5987]_ , \new_[5991]_ , \new_[5992]_ ,
    \new_[5996]_ , \new_[5997]_ , \new_[5998]_ , \new_[6002]_ ,
    \new_[6003]_ , \new_[6007]_ , \new_[6008]_ , \new_[6009]_ ,
    \new_[6013]_ , \new_[6014]_ , \new_[6018]_ , \new_[6019]_ ,
    \new_[6020]_ , \new_[6024]_ , \new_[6025]_ , \new_[6029]_ ,
    \new_[6030]_ , \new_[6031]_ , \new_[6035]_ , \new_[6036]_ ,
    \new_[6040]_ , \new_[6041]_ , \new_[6042]_ , \new_[6046]_ ,
    \new_[6047]_ , \new_[6051]_ , \new_[6052]_ , \new_[6053]_ ,
    \new_[6057]_ , \new_[6058]_ , \new_[6062]_ , \new_[6063]_ ,
    \new_[6064]_ , \new_[6068]_ , \new_[6069]_ , \new_[6073]_ ,
    \new_[6074]_ , \new_[6075]_ , \new_[6079]_ , \new_[6080]_ ,
    \new_[6084]_ , \new_[6085]_ , \new_[6086]_ , \new_[6090]_ ,
    \new_[6091]_ , \new_[6095]_ , \new_[6096]_ , \new_[6097]_ ,
    \new_[6101]_ , \new_[6102]_ , \new_[6106]_ , \new_[6107]_ ,
    \new_[6108]_ , \new_[6112]_ , \new_[6113]_ , \new_[6117]_ ,
    \new_[6118]_ , \new_[6119]_ , \new_[6123]_ , \new_[6124]_ ,
    \new_[6128]_ , \new_[6129]_ , \new_[6130]_ , \new_[6134]_ ,
    \new_[6135]_ , \new_[6139]_ , \new_[6140]_ , \new_[6141]_ ,
    \new_[6145]_ , \new_[6146]_ , \new_[6150]_ , \new_[6151]_ ,
    \new_[6152]_ , \new_[6156]_ , \new_[6157]_ , \new_[6161]_ ,
    \new_[6162]_ , \new_[6163]_ , \new_[6167]_ , \new_[6168]_ ,
    \new_[6172]_ , \new_[6173]_ , \new_[6174]_ , \new_[6178]_ ,
    \new_[6179]_ , \new_[6183]_ , \new_[6184]_ , \new_[6185]_ ,
    \new_[6189]_ , \new_[6190]_ , \new_[6194]_ , \new_[6195]_ ,
    \new_[6196]_ , \new_[6200]_ , \new_[6201]_ , \new_[6205]_ ,
    \new_[6206]_ , \new_[6207]_ , \new_[6211]_ , \new_[6212]_ ,
    \new_[6216]_ , \new_[6217]_ , \new_[6218]_ , \new_[6222]_ ,
    \new_[6223]_ , \new_[6227]_ , \new_[6228]_ , \new_[6229]_ ,
    \new_[6233]_ , \new_[6234]_ , \new_[6238]_ , \new_[6239]_ ,
    \new_[6240]_ , \new_[6244]_ , \new_[6245]_ , \new_[6249]_ ,
    \new_[6250]_ , \new_[6251]_ , \new_[6255]_ , \new_[6256]_ ,
    \new_[6260]_ , \new_[6261]_ , \new_[6262]_ , \new_[6266]_ ,
    \new_[6267]_ , \new_[6271]_ , \new_[6272]_ , \new_[6273]_ ,
    \new_[6277]_ , \new_[6278]_ , \new_[6282]_ , \new_[6283]_ ,
    \new_[6284]_ , \new_[6288]_ , \new_[6289]_ , \new_[6293]_ ,
    \new_[6294]_ , \new_[6295]_ , \new_[6299]_ , \new_[6300]_ ,
    \new_[6304]_ , \new_[6305]_ , \new_[6306]_ , \new_[6310]_ ,
    \new_[6311]_ , \new_[6315]_ , \new_[6316]_ , \new_[6317]_ ,
    \new_[6321]_ , \new_[6322]_ , \new_[6326]_ , \new_[6327]_ ,
    \new_[6328]_ , \new_[6332]_ , \new_[6333]_ , \new_[6337]_ ,
    \new_[6338]_ , \new_[6339]_ , \new_[6343]_ , \new_[6344]_ ,
    \new_[6348]_ , \new_[6349]_ , \new_[6350]_ , \new_[6354]_ ,
    \new_[6355]_ , \new_[6359]_ , \new_[6360]_ , \new_[6361]_ ,
    \new_[6365]_ , \new_[6366]_ , \new_[6370]_ , \new_[6371]_ ,
    \new_[6372]_ , \new_[6376]_ , \new_[6377]_ , \new_[6381]_ ,
    \new_[6382]_ , \new_[6383]_ , \new_[6387]_ , \new_[6388]_ ,
    \new_[6392]_ , \new_[6393]_ , \new_[6394]_ , \new_[6398]_ ,
    \new_[6399]_ , \new_[6403]_ , \new_[6404]_ , \new_[6405]_ ,
    \new_[6409]_ , \new_[6410]_ , \new_[6414]_ , \new_[6415]_ ,
    \new_[6416]_ , \new_[6420]_ , \new_[6421]_ , \new_[6425]_ ,
    \new_[6426]_ , \new_[6427]_ , \new_[6431]_ , \new_[6432]_ ,
    \new_[6436]_ , \new_[6437]_ , \new_[6438]_ , \new_[6442]_ ,
    \new_[6443]_ , \new_[6447]_ , \new_[6448]_ , \new_[6449]_ ,
    \new_[6453]_ , \new_[6454]_ , \new_[6458]_ , \new_[6459]_ ,
    \new_[6460]_ , \new_[6464]_ , \new_[6465]_ , \new_[6469]_ ,
    \new_[6470]_ , \new_[6471]_ , \new_[6475]_ , \new_[6476]_ ,
    \new_[6480]_ , \new_[6481]_ , \new_[6482]_ , \new_[6486]_ ,
    \new_[6487]_ , \new_[6491]_ , \new_[6492]_ , \new_[6493]_ ,
    \new_[6497]_ , \new_[6498]_ , \new_[6502]_ , \new_[6503]_ ,
    \new_[6504]_ , \new_[6508]_ , \new_[6509]_ , \new_[6513]_ ,
    \new_[6514]_ , \new_[6515]_ , \new_[6519]_ , \new_[6520]_ ,
    \new_[6524]_ , \new_[6525]_ , \new_[6526]_ , \new_[6530]_ ,
    \new_[6531]_ , \new_[6535]_ , \new_[6536]_ , \new_[6537]_ ,
    \new_[6541]_ , \new_[6542]_ , \new_[6546]_ , \new_[6547]_ ,
    \new_[6548]_ , \new_[6552]_ , \new_[6553]_ , \new_[6557]_ ,
    \new_[6558]_ , \new_[6559]_ , \new_[6563]_ , \new_[6564]_ ,
    \new_[6568]_ , \new_[6569]_ , \new_[6570]_ , \new_[6574]_ ,
    \new_[6575]_ , \new_[6579]_ , \new_[6580]_ , \new_[6581]_ ,
    \new_[6585]_ , \new_[6586]_ , \new_[6590]_ , \new_[6591]_ ,
    \new_[6592]_ , \new_[6596]_ , \new_[6597]_ , \new_[6601]_ ,
    \new_[6602]_ , \new_[6603]_ , \new_[6607]_ , \new_[6608]_ ,
    \new_[6612]_ , \new_[6613]_ , \new_[6614]_ , \new_[6618]_ ,
    \new_[6619]_ , \new_[6623]_ , \new_[6624]_ , \new_[6625]_ ,
    \new_[6629]_ , \new_[6630]_ , \new_[6634]_ , \new_[6635]_ ,
    \new_[6636]_ , \new_[6640]_ , \new_[6641]_ , \new_[6645]_ ,
    \new_[6646]_ , \new_[6647]_ , \new_[6651]_ , \new_[6652]_ ,
    \new_[6656]_ , \new_[6657]_ , \new_[6658]_ , \new_[6662]_ ,
    \new_[6663]_ , \new_[6667]_ , \new_[6668]_ , \new_[6669]_ ,
    \new_[6673]_ , \new_[6674]_ , \new_[6678]_ , \new_[6679]_ ,
    \new_[6680]_ , \new_[6684]_ , \new_[6685]_ , \new_[6689]_ ,
    \new_[6690]_ , \new_[6691]_ , \new_[6695]_ , \new_[6696]_ ,
    \new_[6700]_ , \new_[6701]_ , \new_[6702]_ , \new_[6706]_ ,
    \new_[6707]_ , \new_[6711]_ , \new_[6712]_ , \new_[6713]_ ,
    \new_[6717]_ , \new_[6718]_ , \new_[6722]_ , \new_[6723]_ ,
    \new_[6724]_ , \new_[6728]_ , \new_[6729]_ , \new_[6733]_ ,
    \new_[6734]_ , \new_[6735]_ , \new_[6739]_ , \new_[6740]_ ,
    \new_[6744]_ , \new_[6745]_ , \new_[6746]_ , \new_[6750]_ ,
    \new_[6751]_ , \new_[6755]_ , \new_[6756]_ , \new_[6757]_ ,
    \new_[6761]_ , \new_[6762]_ , \new_[6766]_ , \new_[6767]_ ,
    \new_[6768]_ , \new_[6772]_ , \new_[6773]_ , \new_[6777]_ ,
    \new_[6778]_ , \new_[6779]_ , \new_[6783]_ , \new_[6784]_ ,
    \new_[6788]_ , \new_[6789]_ , \new_[6790]_ , \new_[6794]_ ,
    \new_[6795]_ , \new_[6799]_ , \new_[6800]_ , \new_[6801]_ ,
    \new_[6805]_ , \new_[6806]_ , \new_[6810]_ , \new_[6811]_ ,
    \new_[6812]_ , \new_[6816]_ , \new_[6817]_ , \new_[6821]_ ,
    \new_[6822]_ , \new_[6823]_ , \new_[6827]_ , \new_[6828]_ ,
    \new_[6832]_ , \new_[6833]_ , \new_[6834]_ , \new_[6838]_ ,
    \new_[6839]_ , \new_[6843]_ , \new_[6844]_ , \new_[6845]_ ,
    \new_[6849]_ , \new_[6850]_ , \new_[6853]_ , \new_[6856]_ ,
    \new_[6857]_ , \new_[6858]_ , \new_[6862]_ , \new_[6863]_ ,
    \new_[6867]_ , \new_[6868]_ , \new_[6869]_ , \new_[6873]_ ,
    \new_[6874]_ , \new_[6877]_ , \new_[6880]_ , \new_[6881]_ ,
    \new_[6882]_ , \new_[6886]_ , \new_[6887]_ , \new_[6891]_ ,
    \new_[6892]_ , \new_[6893]_ , \new_[6897]_ , \new_[6898]_ ,
    \new_[6901]_ , \new_[6904]_ , \new_[6905]_ , \new_[6906]_ ,
    \new_[6910]_ , \new_[6911]_ , \new_[6915]_ , \new_[6916]_ ,
    \new_[6917]_ , \new_[6921]_ , \new_[6922]_ , \new_[6925]_ ,
    \new_[6928]_ , \new_[6929]_ , \new_[6930]_ , \new_[6934]_ ,
    \new_[6935]_ , \new_[6939]_ , \new_[6940]_ , \new_[6941]_ ,
    \new_[6945]_ , \new_[6946]_ , \new_[6949]_ , \new_[6952]_ ,
    \new_[6953]_ , \new_[6954]_ , \new_[6958]_ , \new_[6959]_ ,
    \new_[6963]_ , \new_[6964]_ , \new_[6965]_ , \new_[6969]_ ,
    \new_[6970]_ , \new_[6973]_ , \new_[6976]_ , \new_[6977]_ ,
    \new_[6978]_ , \new_[6982]_ , \new_[6983]_ , \new_[6987]_ ,
    \new_[6988]_ , \new_[6989]_ , \new_[6993]_ , \new_[6994]_ ,
    \new_[6997]_ , \new_[7000]_ , \new_[7001]_ , \new_[7002]_ ,
    \new_[7006]_ , \new_[7007]_ , \new_[7011]_ , \new_[7012]_ ,
    \new_[7013]_ , \new_[7017]_ , \new_[7018]_ , \new_[7021]_ ,
    \new_[7024]_ , \new_[7025]_ , \new_[7026]_ , \new_[7030]_ ,
    \new_[7031]_ , \new_[7035]_ , \new_[7036]_ , \new_[7037]_ ,
    \new_[7041]_ , \new_[7042]_ , \new_[7045]_ , \new_[7048]_ ,
    \new_[7049]_ , \new_[7050]_ , \new_[7054]_ , \new_[7055]_ ,
    \new_[7059]_ , \new_[7060]_ , \new_[7061]_ , \new_[7065]_ ,
    \new_[7066]_ , \new_[7069]_ , \new_[7072]_ , \new_[7073]_ ,
    \new_[7074]_ , \new_[7078]_ , \new_[7079]_ , \new_[7083]_ ,
    \new_[7084]_ , \new_[7085]_ , \new_[7089]_ , \new_[7090]_ ,
    \new_[7093]_ , \new_[7096]_ , \new_[7097]_ , \new_[7098]_ ,
    \new_[7102]_ , \new_[7103]_ , \new_[7107]_ , \new_[7108]_ ,
    \new_[7109]_ , \new_[7113]_ , \new_[7114]_ , \new_[7117]_ ,
    \new_[7120]_ , \new_[7121]_ , \new_[7122]_ , \new_[7126]_ ,
    \new_[7127]_ , \new_[7131]_ , \new_[7132]_ , \new_[7133]_ ,
    \new_[7137]_ , \new_[7138]_ , \new_[7141]_ , \new_[7144]_ ,
    \new_[7145]_ , \new_[7146]_ , \new_[7150]_ , \new_[7151]_ ,
    \new_[7155]_ , \new_[7156]_ , \new_[7157]_ , \new_[7161]_ ,
    \new_[7162]_ , \new_[7165]_ , \new_[7168]_ , \new_[7169]_ ,
    \new_[7170]_ , \new_[7174]_ , \new_[7175]_ , \new_[7179]_ ,
    \new_[7180]_ , \new_[7181]_ , \new_[7185]_ , \new_[7186]_ ,
    \new_[7189]_ , \new_[7192]_ , \new_[7193]_ , \new_[7194]_ ,
    \new_[7198]_ , \new_[7199]_ , \new_[7203]_ , \new_[7204]_ ,
    \new_[7205]_ , \new_[7209]_ , \new_[7210]_ , \new_[7213]_ ,
    \new_[7216]_ , \new_[7217]_ , \new_[7218]_ , \new_[7222]_ ,
    \new_[7223]_ , \new_[7227]_ , \new_[7228]_ , \new_[7229]_ ,
    \new_[7233]_ , \new_[7234]_ , \new_[7237]_ , \new_[7240]_ ,
    \new_[7241]_ , \new_[7242]_ , \new_[7246]_ , \new_[7247]_ ,
    \new_[7251]_ , \new_[7252]_ , \new_[7253]_ , \new_[7257]_ ,
    \new_[7258]_ , \new_[7261]_ , \new_[7264]_ , \new_[7265]_ ,
    \new_[7266]_ , \new_[7270]_ , \new_[7271]_ , \new_[7275]_ ,
    \new_[7276]_ , \new_[7277]_ , \new_[7281]_ , \new_[7282]_ ,
    \new_[7285]_ , \new_[7288]_ , \new_[7289]_ , \new_[7290]_ ,
    \new_[7294]_ , \new_[7295]_ , \new_[7299]_ , \new_[7300]_ ,
    \new_[7301]_ , \new_[7305]_ , \new_[7306]_ , \new_[7309]_ ,
    \new_[7312]_ , \new_[7313]_ , \new_[7314]_ , \new_[7318]_ ,
    \new_[7319]_ , \new_[7323]_ , \new_[7324]_ , \new_[7325]_ ,
    \new_[7329]_ , \new_[7330]_ , \new_[7333]_ , \new_[7336]_ ,
    \new_[7337]_ , \new_[7338]_ , \new_[7342]_ , \new_[7343]_ ,
    \new_[7347]_ , \new_[7348]_ , \new_[7349]_ , \new_[7353]_ ,
    \new_[7354]_ , \new_[7357]_ , \new_[7360]_ , \new_[7361]_ ,
    \new_[7362]_ , \new_[7366]_ , \new_[7367]_ , \new_[7371]_ ,
    \new_[7372]_ , \new_[7373]_ , \new_[7377]_ , \new_[7378]_ ,
    \new_[7381]_ , \new_[7384]_ , \new_[7385]_ , \new_[7386]_ ,
    \new_[7390]_ , \new_[7391]_ , \new_[7395]_ , \new_[7396]_ ,
    \new_[7397]_ , \new_[7401]_ , \new_[7402]_ , \new_[7405]_ ,
    \new_[7408]_ , \new_[7409]_ , \new_[7410]_ , \new_[7414]_ ,
    \new_[7415]_ , \new_[7419]_ , \new_[7420]_ , \new_[7421]_ ,
    \new_[7425]_ , \new_[7426]_ , \new_[7429]_ , \new_[7432]_ ,
    \new_[7433]_ , \new_[7434]_ , \new_[7438]_ , \new_[7439]_ ,
    \new_[7443]_ , \new_[7444]_ , \new_[7445]_ , \new_[7449]_ ,
    \new_[7450]_ , \new_[7453]_ , \new_[7456]_ , \new_[7457]_ ,
    \new_[7458]_ , \new_[7462]_ , \new_[7463]_ , \new_[7467]_ ,
    \new_[7468]_ , \new_[7469]_ , \new_[7473]_ , \new_[7474]_ ,
    \new_[7477]_ , \new_[7480]_ , \new_[7481]_ , \new_[7482]_ ,
    \new_[7486]_ , \new_[7487]_ , \new_[7491]_ , \new_[7492]_ ,
    \new_[7493]_ , \new_[7497]_ , \new_[7498]_ , \new_[7501]_ ,
    \new_[7504]_ , \new_[7505]_ , \new_[7506]_ , \new_[7510]_ ,
    \new_[7511]_ , \new_[7515]_ , \new_[7516]_ , \new_[7517]_ ,
    \new_[7521]_ , \new_[7522]_ , \new_[7525]_ , \new_[7528]_ ,
    \new_[7529]_ , \new_[7530]_ , \new_[7534]_ , \new_[7535]_ ,
    \new_[7539]_ , \new_[7540]_ , \new_[7541]_ , \new_[7545]_ ,
    \new_[7546]_ , \new_[7549]_ , \new_[7552]_ , \new_[7553]_ ,
    \new_[7554]_ , \new_[7558]_ , \new_[7559]_ , \new_[7563]_ ,
    \new_[7564]_ , \new_[7565]_ , \new_[7569]_ , \new_[7570]_ ,
    \new_[7573]_ , \new_[7576]_ , \new_[7577]_ , \new_[7578]_ ,
    \new_[7582]_ , \new_[7583]_ , \new_[7587]_ , \new_[7588]_ ,
    \new_[7589]_ , \new_[7593]_ , \new_[7594]_ , \new_[7597]_ ,
    \new_[7600]_ , \new_[7601]_ , \new_[7602]_ , \new_[7606]_ ,
    \new_[7607]_ , \new_[7611]_ , \new_[7612]_ , \new_[7613]_ ,
    \new_[7617]_ , \new_[7618]_ , \new_[7621]_ , \new_[7624]_ ,
    \new_[7625]_ , \new_[7626]_ , \new_[7630]_ , \new_[7631]_ ,
    \new_[7635]_ , \new_[7636]_ , \new_[7637]_ , \new_[7641]_ ,
    \new_[7642]_ , \new_[7645]_ , \new_[7648]_ , \new_[7649]_ ,
    \new_[7650]_ , \new_[7654]_ , \new_[7655]_ , \new_[7659]_ ,
    \new_[7660]_ , \new_[7661]_ , \new_[7665]_ , \new_[7666]_ ,
    \new_[7669]_ , \new_[7672]_ , \new_[7673]_ , \new_[7674]_ ,
    \new_[7678]_ , \new_[7679]_ , \new_[7683]_ , \new_[7684]_ ,
    \new_[7685]_ , \new_[7689]_ , \new_[7690]_ , \new_[7693]_ ,
    \new_[7696]_ , \new_[7697]_ , \new_[7698]_ , \new_[7702]_ ,
    \new_[7703]_ , \new_[7707]_ , \new_[7708]_ , \new_[7709]_ ,
    \new_[7713]_ , \new_[7714]_ , \new_[7717]_ , \new_[7720]_ ,
    \new_[7721]_ , \new_[7722]_ , \new_[7726]_ , \new_[7727]_ ,
    \new_[7731]_ , \new_[7732]_ , \new_[7733]_ , \new_[7737]_ ,
    \new_[7738]_ , \new_[7741]_ , \new_[7744]_ , \new_[7745]_ ,
    \new_[7746]_ , \new_[7750]_ , \new_[7751]_ , \new_[7755]_ ,
    \new_[7756]_ , \new_[7757]_ , \new_[7761]_ , \new_[7762]_ ,
    \new_[7765]_ , \new_[7768]_ , \new_[7769]_ , \new_[7770]_ ,
    \new_[7774]_ , \new_[7775]_ , \new_[7779]_ , \new_[7780]_ ,
    \new_[7781]_ , \new_[7785]_ , \new_[7786]_ , \new_[7789]_ ,
    \new_[7792]_ , \new_[7793]_ , \new_[7794]_ , \new_[7798]_ ,
    \new_[7799]_ , \new_[7803]_ , \new_[7804]_ , \new_[7805]_ ,
    \new_[7809]_ , \new_[7810]_ , \new_[7813]_ , \new_[7816]_ ,
    \new_[7817]_ , \new_[7818]_ , \new_[7822]_ , \new_[7823]_ ,
    \new_[7827]_ , \new_[7828]_ , \new_[7829]_ , \new_[7833]_ ,
    \new_[7834]_ , \new_[7837]_ , \new_[7840]_ , \new_[7841]_ ,
    \new_[7842]_ , \new_[7846]_ , \new_[7847]_ , \new_[7851]_ ,
    \new_[7852]_ , \new_[7853]_ , \new_[7857]_ , \new_[7858]_ ,
    \new_[7861]_ , \new_[7864]_ , \new_[7865]_ , \new_[7866]_ ,
    \new_[7870]_ , \new_[7871]_ , \new_[7875]_ , \new_[7876]_ ,
    \new_[7877]_ , \new_[7881]_ , \new_[7882]_ , \new_[7885]_ ,
    \new_[7888]_ , \new_[7889]_ , \new_[7890]_ , \new_[7894]_ ,
    \new_[7895]_ , \new_[7899]_ , \new_[7900]_ , \new_[7901]_ ,
    \new_[7905]_ , \new_[7906]_ , \new_[7909]_ , \new_[7912]_ ,
    \new_[7913]_ , \new_[7914]_ , \new_[7918]_ , \new_[7919]_ ,
    \new_[7923]_ , \new_[7924]_ , \new_[7925]_ , \new_[7929]_ ,
    \new_[7930]_ , \new_[7933]_ , \new_[7936]_ , \new_[7937]_ ,
    \new_[7938]_ , \new_[7942]_ , \new_[7943]_ , \new_[7947]_ ,
    \new_[7948]_ , \new_[7949]_ , \new_[7953]_ , \new_[7954]_ ,
    \new_[7957]_ , \new_[7960]_ , \new_[7961]_ , \new_[7962]_ ,
    \new_[7966]_ , \new_[7967]_ , \new_[7971]_ , \new_[7972]_ ,
    \new_[7973]_ , \new_[7977]_ , \new_[7978]_ , \new_[7981]_ ,
    \new_[7984]_ , \new_[7985]_ , \new_[7986]_ , \new_[7990]_ ,
    \new_[7991]_ , \new_[7994]_ , \new_[7997]_ , \new_[7998]_ ,
    \new_[7999]_ , \new_[8003]_ , \new_[8004]_ , \new_[8007]_ ,
    \new_[8010]_ , \new_[8011]_ , \new_[8012]_ , \new_[8016]_ ,
    \new_[8017]_ , \new_[8020]_ , \new_[8023]_ , \new_[8024]_ ,
    \new_[8025]_ , \new_[8029]_ , \new_[8030]_ , \new_[8033]_ ,
    \new_[8036]_ , \new_[8037]_ , \new_[8038]_ , \new_[8042]_ ,
    \new_[8043]_ , \new_[8046]_ , \new_[8049]_ , \new_[8050]_ ,
    \new_[8051]_ , \new_[8055]_ , \new_[8056]_ , \new_[8059]_ ,
    \new_[8062]_ , \new_[8063]_ , \new_[8064]_ , \new_[8068]_ ,
    \new_[8069]_ , \new_[8072]_ , \new_[8075]_ , \new_[8076]_ ,
    \new_[8077]_ , \new_[8081]_ , \new_[8082]_ , \new_[8085]_ ,
    \new_[8088]_ , \new_[8089]_ , \new_[8090]_ , \new_[8094]_ ,
    \new_[8095]_ , \new_[8098]_ , \new_[8101]_ , \new_[8102]_ ,
    \new_[8103]_ , \new_[8107]_ , \new_[8108]_ , \new_[8111]_ ,
    \new_[8114]_ , \new_[8115]_ , \new_[8116]_ , \new_[8120]_ ,
    \new_[8121]_ , \new_[8124]_ , \new_[8127]_ , \new_[8128]_ ,
    \new_[8129]_ , \new_[8133]_ , \new_[8134]_ , \new_[8137]_ ,
    \new_[8140]_ , \new_[8141]_ , \new_[8142]_ , \new_[8146]_ ,
    \new_[8147]_ , \new_[8150]_ , \new_[8153]_ , \new_[8154]_ ,
    \new_[8155]_ , \new_[8159]_ , \new_[8160]_ , \new_[8163]_ ,
    \new_[8166]_ , \new_[8167]_ , \new_[8168]_ , \new_[8172]_ ,
    \new_[8173]_ , \new_[8176]_ , \new_[8179]_ , \new_[8180]_ ,
    \new_[8181]_ , \new_[8185]_ , \new_[8186]_ , \new_[8189]_ ,
    \new_[8192]_ , \new_[8193]_ , \new_[8194]_ , \new_[8198]_ ,
    \new_[8199]_ , \new_[8202]_ , \new_[8205]_ , \new_[8206]_ ,
    \new_[8207]_ , \new_[8211]_ , \new_[8212]_ , \new_[8215]_ ,
    \new_[8218]_ , \new_[8219]_ , \new_[8220]_ , \new_[8224]_ ,
    \new_[8225]_ , \new_[8228]_ , \new_[8231]_ , \new_[8232]_ ,
    \new_[8233]_ , \new_[8237]_ , \new_[8238]_ , \new_[8241]_ ,
    \new_[8244]_ , \new_[8245]_ , \new_[8246]_ , \new_[8250]_ ,
    \new_[8251]_ , \new_[8254]_ , \new_[8257]_ , \new_[8258]_ ,
    \new_[8259]_ , \new_[8263]_ , \new_[8264]_ , \new_[8267]_ ,
    \new_[8270]_ , \new_[8271]_ , \new_[8272]_ , \new_[8276]_ ,
    \new_[8277]_ , \new_[8280]_ , \new_[8283]_ , \new_[8284]_ ,
    \new_[8285]_ , \new_[8289]_ , \new_[8290]_ , \new_[8293]_ ,
    \new_[8296]_ , \new_[8297]_ , \new_[8298]_ , \new_[8302]_ ,
    \new_[8303]_ , \new_[8306]_ , \new_[8309]_ , \new_[8310]_ ,
    \new_[8311]_ , \new_[8315]_ , \new_[8316]_ , \new_[8319]_ ,
    \new_[8322]_ , \new_[8323]_ , \new_[8324]_ , \new_[8328]_ ,
    \new_[8329]_ , \new_[8332]_ , \new_[8335]_ , \new_[8336]_ ,
    \new_[8337]_ , \new_[8341]_ , \new_[8342]_ , \new_[8345]_ ,
    \new_[8348]_ , \new_[8349]_ , \new_[8350]_ , \new_[8354]_ ,
    \new_[8355]_ , \new_[8358]_ , \new_[8361]_ , \new_[8362]_ ,
    \new_[8363]_ , \new_[8367]_ , \new_[8368]_ , \new_[8371]_ ,
    \new_[8374]_ , \new_[8375]_ , \new_[8376]_ , \new_[8380]_ ,
    \new_[8381]_ , \new_[8384]_ , \new_[8387]_ , \new_[8388]_ ,
    \new_[8389]_ , \new_[8393]_ , \new_[8394]_ , \new_[8397]_ ,
    \new_[8400]_ , \new_[8401]_ , \new_[8402]_ , \new_[8406]_ ,
    \new_[8407]_ , \new_[8410]_ , \new_[8413]_ , \new_[8414]_ ,
    \new_[8415]_ , \new_[8419]_ , \new_[8420]_ , \new_[8423]_ ,
    \new_[8426]_ , \new_[8427]_ , \new_[8428]_ , \new_[8432]_ ,
    \new_[8433]_ , \new_[8436]_ , \new_[8439]_ , \new_[8440]_ ,
    \new_[8441]_ , \new_[8445]_ , \new_[8446]_ , \new_[8449]_ ,
    \new_[8452]_ , \new_[8453]_ , \new_[8454]_ , \new_[8458]_ ,
    \new_[8459]_ , \new_[8462]_ , \new_[8465]_ , \new_[8466]_ ,
    \new_[8467]_ , \new_[8471]_ , \new_[8472]_ , \new_[8475]_ ,
    \new_[8478]_ , \new_[8479]_ , \new_[8480]_ , \new_[8484]_ ,
    \new_[8485]_ , \new_[8488]_ , \new_[8491]_ , \new_[8492]_ ,
    \new_[8493]_ , \new_[8497]_ , \new_[8498]_ , \new_[8501]_ ,
    \new_[8504]_ , \new_[8505]_ , \new_[8506]_ , \new_[8510]_ ,
    \new_[8511]_ , \new_[8514]_ , \new_[8517]_ , \new_[8518]_ ,
    \new_[8519]_ , \new_[8523]_ , \new_[8524]_ , \new_[8527]_ ,
    \new_[8530]_ , \new_[8531]_ , \new_[8532]_ , \new_[8536]_ ,
    \new_[8537]_ , \new_[8540]_ , \new_[8543]_ , \new_[8544]_ ,
    \new_[8545]_ , \new_[8549]_ , \new_[8550]_ , \new_[8553]_ ,
    \new_[8556]_ , \new_[8557]_ , \new_[8558]_ , \new_[8562]_ ,
    \new_[8563]_ , \new_[8566]_ , \new_[8569]_ , \new_[8570]_ ,
    \new_[8571]_ , \new_[8575]_ , \new_[8576]_ , \new_[8579]_ ,
    \new_[8582]_ , \new_[8583]_ , \new_[8584]_ , \new_[8588]_ ,
    \new_[8589]_ , \new_[8592]_ , \new_[8595]_ , \new_[8596]_ ,
    \new_[8597]_ , \new_[8601]_ , \new_[8602]_ , \new_[8605]_ ,
    \new_[8608]_ , \new_[8609]_ , \new_[8610]_ , \new_[8614]_ ,
    \new_[8615]_ , \new_[8618]_ , \new_[8621]_ , \new_[8622]_ ,
    \new_[8623]_ , \new_[8627]_ , \new_[8628]_ , \new_[8631]_ ,
    \new_[8634]_ , \new_[8635]_ , \new_[8636]_ , \new_[8640]_ ,
    \new_[8641]_ , \new_[8644]_ , \new_[8647]_ , \new_[8648]_ ,
    \new_[8649]_ , \new_[8653]_ , \new_[8654]_ , \new_[8657]_ ,
    \new_[8660]_ , \new_[8661]_ , \new_[8662]_ , \new_[8666]_ ,
    \new_[8667]_ , \new_[8670]_ , \new_[8673]_ , \new_[8674]_ ,
    \new_[8675]_ , \new_[8679]_ , \new_[8680]_ , \new_[8683]_ ,
    \new_[8686]_ , \new_[8687]_ , \new_[8688]_ , \new_[8692]_ ,
    \new_[8693]_ , \new_[8696]_ , \new_[8699]_ , \new_[8700]_ ,
    \new_[8701]_ , \new_[8705]_ , \new_[8706]_ , \new_[8709]_ ,
    \new_[8712]_ , \new_[8713]_ , \new_[8714]_ , \new_[8718]_ ,
    \new_[8719]_ , \new_[8722]_ , \new_[8725]_ , \new_[8726]_ ,
    \new_[8727]_ , \new_[8731]_ , \new_[8732]_ , \new_[8735]_ ,
    \new_[8738]_ , \new_[8739]_ , \new_[8740]_ , \new_[8744]_ ,
    \new_[8745]_ , \new_[8748]_ , \new_[8751]_ , \new_[8752]_ ,
    \new_[8753]_ , \new_[8757]_ , \new_[8758]_ , \new_[8761]_ ,
    \new_[8764]_ , \new_[8765]_ , \new_[8766]_ , \new_[8770]_ ,
    \new_[8771]_ , \new_[8774]_ , \new_[8777]_ , \new_[8778]_ ,
    \new_[8779]_ , \new_[8783]_ , \new_[8784]_ , \new_[8787]_ ,
    \new_[8790]_ , \new_[8791]_ , \new_[8792]_ , \new_[8796]_ ,
    \new_[8797]_ , \new_[8800]_ , \new_[8803]_ , \new_[8804]_ ,
    \new_[8805]_ , \new_[8809]_ , \new_[8810]_ , \new_[8813]_ ,
    \new_[8816]_ , \new_[8817]_ , \new_[8818]_ , \new_[8822]_ ,
    \new_[8823]_ , \new_[8826]_ , \new_[8829]_ , \new_[8830]_ ,
    \new_[8831]_ , \new_[8835]_ , \new_[8836]_ , \new_[8839]_ ,
    \new_[8842]_ , \new_[8843]_ , \new_[8844]_ , \new_[8848]_ ,
    \new_[8849]_ , \new_[8852]_ , \new_[8855]_ , \new_[8856]_ ,
    \new_[8857]_ , \new_[8861]_ , \new_[8862]_ , \new_[8865]_ ,
    \new_[8868]_ , \new_[8869]_ , \new_[8870]_ , \new_[8874]_ ,
    \new_[8875]_ , \new_[8878]_ , \new_[8881]_ , \new_[8882]_ ,
    \new_[8883]_ , \new_[8887]_ , \new_[8888]_ , \new_[8891]_ ,
    \new_[8894]_ , \new_[8895]_ , \new_[8896]_ , \new_[8900]_ ,
    \new_[8901]_ , \new_[8904]_ , \new_[8907]_ , \new_[8908]_ ,
    \new_[8909]_ , \new_[8913]_ , \new_[8914]_ , \new_[8917]_ ,
    \new_[8920]_ , \new_[8921]_ , \new_[8922]_ , \new_[8926]_ ,
    \new_[8927]_ , \new_[8930]_ , \new_[8933]_ , \new_[8934]_ ,
    \new_[8935]_ , \new_[8939]_ , \new_[8940]_ , \new_[8943]_ ,
    \new_[8946]_ , \new_[8947]_ , \new_[8948]_ , \new_[8952]_ ,
    \new_[8953]_ , \new_[8956]_ , \new_[8959]_ , \new_[8960]_ ,
    \new_[8961]_ , \new_[8965]_ , \new_[8966]_ , \new_[8969]_ ,
    \new_[8972]_ , \new_[8973]_ , \new_[8974]_ , \new_[8978]_ ,
    \new_[8979]_ , \new_[8982]_ , \new_[8985]_ , \new_[8986]_ ,
    \new_[8987]_ , \new_[8991]_ , \new_[8992]_ , \new_[8995]_ ,
    \new_[8998]_ , \new_[8999]_ , \new_[9000]_ , \new_[9004]_ ,
    \new_[9005]_ , \new_[9008]_ , \new_[9011]_ , \new_[9012]_ ,
    \new_[9013]_ , \new_[9017]_ , \new_[9018]_ , \new_[9021]_ ,
    \new_[9024]_ , \new_[9025]_ , \new_[9026]_ , \new_[9030]_ ,
    \new_[9031]_ , \new_[9034]_ , \new_[9037]_ , \new_[9038]_ ,
    \new_[9039]_ , \new_[9043]_ , \new_[9044]_ , \new_[9047]_ ,
    \new_[9050]_ , \new_[9051]_ , \new_[9052]_ , \new_[9056]_ ,
    \new_[9057]_ , \new_[9060]_ , \new_[9063]_ , \new_[9064]_ ,
    \new_[9065]_ , \new_[9069]_ , \new_[9070]_ , \new_[9073]_ ,
    \new_[9076]_ , \new_[9077]_ , \new_[9078]_ , \new_[9082]_ ,
    \new_[9083]_ , \new_[9086]_ , \new_[9089]_ , \new_[9090]_ ,
    \new_[9091]_ , \new_[9095]_ , \new_[9096]_ , \new_[9099]_ ,
    \new_[9102]_ , \new_[9103]_ , \new_[9104]_ , \new_[9108]_ ,
    \new_[9109]_ , \new_[9112]_ , \new_[9115]_ , \new_[9116]_ ,
    \new_[9117]_ , \new_[9121]_ , \new_[9122]_ , \new_[9125]_ ,
    \new_[9128]_ , \new_[9129]_ , \new_[9130]_ , \new_[9134]_ ,
    \new_[9135]_ , \new_[9138]_ , \new_[9141]_ , \new_[9142]_ ,
    \new_[9143]_ , \new_[9147]_ , \new_[9148]_ , \new_[9151]_ ,
    \new_[9154]_ , \new_[9155]_ , \new_[9156]_ , \new_[9160]_ ,
    \new_[9161]_ , \new_[9164]_ , \new_[9167]_ , \new_[9168]_ ,
    \new_[9169]_ , \new_[9173]_ , \new_[9174]_ , \new_[9177]_ ,
    \new_[9180]_ , \new_[9181]_ , \new_[9182]_ , \new_[9186]_ ,
    \new_[9187]_ , \new_[9190]_ , \new_[9193]_ , \new_[9194]_ ,
    \new_[9195]_ , \new_[9199]_ , \new_[9200]_ , \new_[9203]_ ,
    \new_[9206]_ , \new_[9207]_ , \new_[9208]_ , \new_[9212]_ ,
    \new_[9213]_ , \new_[9216]_ , \new_[9219]_ , \new_[9220]_ ,
    \new_[9221]_ , \new_[9225]_ , \new_[9226]_ , \new_[9229]_ ,
    \new_[9232]_ , \new_[9233]_ , \new_[9234]_ , \new_[9238]_ ,
    \new_[9239]_ , \new_[9242]_ , \new_[9245]_ , \new_[9246]_ ,
    \new_[9247]_ , \new_[9251]_ , \new_[9252]_ , \new_[9255]_ ,
    \new_[9258]_ , \new_[9259]_ , \new_[9260]_ , \new_[9264]_ ,
    \new_[9265]_ , \new_[9268]_ , \new_[9271]_ , \new_[9272]_ ,
    \new_[9273]_ , \new_[9277]_ , \new_[9278]_ , \new_[9281]_ ,
    \new_[9284]_ , \new_[9285]_ , \new_[9286]_ , \new_[9290]_ ,
    \new_[9291]_ , \new_[9294]_ , \new_[9297]_ , \new_[9298]_ ,
    \new_[9299]_ , \new_[9303]_ , \new_[9304]_ , \new_[9307]_ ,
    \new_[9310]_ , \new_[9311]_ , \new_[9312]_ , \new_[9316]_ ,
    \new_[9317]_ , \new_[9320]_ , \new_[9323]_ , \new_[9324]_ ,
    \new_[9325]_ , \new_[9329]_ , \new_[9330]_ , \new_[9333]_ ,
    \new_[9336]_ , \new_[9337]_ , \new_[9338]_ , \new_[9342]_ ,
    \new_[9343]_ , \new_[9346]_ , \new_[9349]_ , \new_[9350]_ ,
    \new_[9351]_ , \new_[9355]_ , \new_[9356]_ , \new_[9359]_ ,
    \new_[9362]_ , \new_[9363]_ , \new_[9364]_ , \new_[9368]_ ,
    \new_[9369]_ , \new_[9372]_ , \new_[9375]_ , \new_[9376]_ ,
    \new_[9377]_ , \new_[9381]_ , \new_[9382]_ , \new_[9385]_ ,
    \new_[9388]_ , \new_[9389]_ , \new_[9390]_ , \new_[9394]_ ,
    \new_[9395]_ , \new_[9398]_ , \new_[9401]_ , \new_[9402]_ ,
    \new_[9403]_ , \new_[9407]_ , \new_[9408]_ , \new_[9411]_ ,
    \new_[9414]_ , \new_[9415]_ , \new_[9416]_ , \new_[9420]_ ,
    \new_[9421]_ , \new_[9424]_ , \new_[9427]_ , \new_[9428]_ ,
    \new_[9429]_ , \new_[9433]_ , \new_[9434]_ , \new_[9437]_ ,
    \new_[9440]_ , \new_[9441]_ , \new_[9442]_ , \new_[9446]_ ,
    \new_[9447]_ , \new_[9450]_ , \new_[9453]_ , \new_[9454]_ ,
    \new_[9455]_ , \new_[9459]_ , \new_[9460]_ , \new_[9463]_ ,
    \new_[9466]_ , \new_[9467]_ , \new_[9468]_ , \new_[9472]_ ,
    \new_[9473]_ , \new_[9476]_ , \new_[9479]_ , \new_[9480]_ ,
    \new_[9481]_ , \new_[9485]_ , \new_[9486]_ , \new_[9489]_ ,
    \new_[9492]_ , \new_[9493]_ , \new_[9494]_ , \new_[9498]_ ,
    \new_[9499]_ , \new_[9502]_ , \new_[9505]_ , \new_[9506]_ ,
    \new_[9507]_ , \new_[9511]_ , \new_[9512]_ , \new_[9515]_ ,
    \new_[9518]_ , \new_[9519]_ , \new_[9520]_ , \new_[9524]_ ,
    \new_[9525]_ , \new_[9528]_ , \new_[9531]_ , \new_[9532]_ ,
    \new_[9533]_ , \new_[9537]_ , \new_[9538]_ , \new_[9541]_ ,
    \new_[9544]_ , \new_[9545]_ , \new_[9546]_ , \new_[9550]_ ,
    \new_[9551]_ , \new_[9554]_ , \new_[9557]_ , \new_[9558]_ ,
    \new_[9559]_ , \new_[9563]_ , \new_[9564]_ , \new_[9567]_ ,
    \new_[9570]_ , \new_[9571]_ , \new_[9572]_ , \new_[9576]_ ,
    \new_[9577]_ , \new_[9580]_ , \new_[9583]_ , \new_[9584]_ ,
    \new_[9585]_ , \new_[9589]_ , \new_[9590]_ , \new_[9593]_ ,
    \new_[9596]_ , \new_[9597]_ , \new_[9598]_ , \new_[9602]_ ,
    \new_[9603]_ , \new_[9606]_ , \new_[9609]_ , \new_[9610]_ ,
    \new_[9611]_ , \new_[9615]_ , \new_[9616]_ , \new_[9619]_ ,
    \new_[9622]_ , \new_[9623]_ , \new_[9624]_ , \new_[9628]_ ,
    \new_[9629]_ , \new_[9632]_ , \new_[9635]_ , \new_[9636]_ ,
    \new_[9637]_ , \new_[9641]_ , \new_[9642]_ , \new_[9645]_ ,
    \new_[9648]_ , \new_[9649]_ , \new_[9650]_ , \new_[9654]_ ,
    \new_[9655]_ , \new_[9658]_ , \new_[9661]_ , \new_[9662]_ ,
    \new_[9663]_ , \new_[9667]_ , \new_[9668]_ , \new_[9671]_ ,
    \new_[9674]_ , \new_[9675]_ , \new_[9676]_ , \new_[9680]_ ,
    \new_[9681]_ , \new_[9684]_ , \new_[9687]_ , \new_[9688]_ ,
    \new_[9689]_ , \new_[9693]_ , \new_[9694]_ , \new_[9697]_ ,
    \new_[9700]_ , \new_[9701]_ , \new_[9702]_ , \new_[9706]_ ,
    \new_[9707]_ , \new_[9710]_ , \new_[9713]_ , \new_[9714]_ ,
    \new_[9715]_ , \new_[9719]_ , \new_[9720]_ , \new_[9723]_ ,
    \new_[9726]_ , \new_[9727]_ , \new_[9728]_ , \new_[9732]_ ,
    \new_[9733]_ , \new_[9736]_ , \new_[9739]_ , \new_[9740]_ ,
    \new_[9741]_ , \new_[9745]_ , \new_[9746]_ , \new_[9749]_ ,
    \new_[9752]_ , \new_[9753]_ , \new_[9754]_ , \new_[9758]_ ,
    \new_[9759]_ , \new_[9762]_ , \new_[9765]_ , \new_[9766]_ ,
    \new_[9767]_ , \new_[9771]_ , \new_[9772]_ , \new_[9775]_ ,
    \new_[9778]_ , \new_[9779]_ , \new_[9780]_ , \new_[9784]_ ,
    \new_[9785]_ , \new_[9788]_ , \new_[9791]_ , \new_[9792]_ ,
    \new_[9793]_ , \new_[9797]_ , \new_[9798]_ , \new_[9801]_ ,
    \new_[9804]_ , \new_[9805]_ , \new_[9806]_ , \new_[9810]_ ,
    \new_[9811]_ , \new_[9814]_ , \new_[9817]_ , \new_[9818]_ ,
    \new_[9819]_ , \new_[9823]_ , \new_[9824]_ , \new_[9827]_ ,
    \new_[9830]_ , \new_[9831]_ , \new_[9832]_ , \new_[9836]_ ,
    \new_[9837]_ , \new_[9840]_ , \new_[9843]_ , \new_[9844]_ ,
    \new_[9845]_ , \new_[9849]_ , \new_[9850]_ , \new_[9853]_ ,
    \new_[9856]_ , \new_[9857]_ , \new_[9858]_ , \new_[9862]_ ,
    \new_[9863]_ , \new_[9866]_ , \new_[9869]_ , \new_[9870]_ ,
    \new_[9871]_ , \new_[9875]_ , \new_[9876]_ , \new_[9879]_ ,
    \new_[9882]_ , \new_[9883]_ , \new_[9884]_ , \new_[9888]_ ,
    \new_[9889]_ , \new_[9892]_ , \new_[9895]_ , \new_[9896]_ ,
    \new_[9897]_ , \new_[9901]_ , \new_[9902]_ , \new_[9905]_ ,
    \new_[9908]_ , \new_[9909]_ , \new_[9910]_ , \new_[9914]_ ,
    \new_[9915]_ , \new_[9918]_ , \new_[9921]_ , \new_[9922]_ ,
    \new_[9923]_ , \new_[9927]_ , \new_[9928]_ , \new_[9931]_ ,
    \new_[9934]_ , \new_[9935]_ , \new_[9936]_ , \new_[9940]_ ,
    \new_[9941]_ , \new_[9944]_ , \new_[9947]_ , \new_[9948]_ ,
    \new_[9949]_ , \new_[9953]_ , \new_[9954]_ , \new_[9957]_ ,
    \new_[9960]_ , \new_[9961]_ , \new_[9962]_ , \new_[9966]_ ,
    \new_[9967]_ , \new_[9970]_ , \new_[9973]_ , \new_[9974]_ ,
    \new_[9975]_ , \new_[9979]_ , \new_[9980]_ , \new_[9983]_ ,
    \new_[9986]_ , \new_[9987]_ , \new_[9988]_ , \new_[9992]_ ,
    \new_[9993]_ , \new_[9996]_ , \new_[9999]_ , \new_[10000]_ ,
    \new_[10001]_ , \new_[10005]_ , \new_[10006]_ , \new_[10009]_ ,
    \new_[10012]_ , \new_[10013]_ , \new_[10014]_ , \new_[10018]_ ,
    \new_[10019]_ , \new_[10022]_ , \new_[10025]_ , \new_[10026]_ ,
    \new_[10027]_ , \new_[10031]_ , \new_[10032]_ , \new_[10035]_ ,
    \new_[10038]_ , \new_[10039]_ , \new_[10040]_ , \new_[10044]_ ,
    \new_[10045]_ , \new_[10048]_ , \new_[10051]_ , \new_[10052]_ ,
    \new_[10053]_ , \new_[10057]_ , \new_[10058]_ , \new_[10061]_ ,
    \new_[10064]_ , \new_[10065]_ , \new_[10066]_ , \new_[10070]_ ,
    \new_[10071]_ , \new_[10074]_ , \new_[10077]_ , \new_[10078]_ ,
    \new_[10079]_ , \new_[10083]_ , \new_[10084]_ , \new_[10087]_ ,
    \new_[10090]_ , \new_[10091]_ , \new_[10092]_ , \new_[10096]_ ,
    \new_[10097]_ , \new_[10100]_ , \new_[10103]_ , \new_[10104]_ ,
    \new_[10105]_ , \new_[10109]_ , \new_[10110]_ , \new_[10113]_ ,
    \new_[10116]_ , \new_[10117]_ , \new_[10118]_ , \new_[10122]_ ,
    \new_[10123]_ , \new_[10126]_ , \new_[10129]_ , \new_[10130]_ ,
    \new_[10131]_ , \new_[10135]_ , \new_[10136]_ , \new_[10139]_ ,
    \new_[10142]_ , \new_[10143]_ , \new_[10144]_ , \new_[10148]_ ,
    \new_[10149]_ , \new_[10152]_ , \new_[10155]_ , \new_[10156]_ ,
    \new_[10157]_ , \new_[10161]_ , \new_[10162]_ , \new_[10165]_ ,
    \new_[10168]_ , \new_[10169]_ , \new_[10170]_ , \new_[10174]_ ,
    \new_[10175]_ , \new_[10178]_ , \new_[10181]_ , \new_[10182]_ ,
    \new_[10183]_ , \new_[10187]_ , \new_[10188]_ , \new_[10191]_ ,
    \new_[10194]_ , \new_[10195]_ , \new_[10196]_ , \new_[10200]_ ,
    \new_[10201]_ , \new_[10204]_ , \new_[10207]_ , \new_[10208]_ ,
    \new_[10209]_ , \new_[10213]_ , \new_[10214]_ , \new_[10217]_ ,
    \new_[10220]_ , \new_[10221]_ , \new_[10222]_ , \new_[10226]_ ,
    \new_[10227]_ , \new_[10230]_ , \new_[10233]_ , \new_[10234]_ ,
    \new_[10235]_ , \new_[10239]_ , \new_[10240]_ , \new_[10243]_ ,
    \new_[10246]_ , \new_[10247]_ , \new_[10248]_ , \new_[10252]_ ,
    \new_[10253]_ , \new_[10256]_ , \new_[10259]_ , \new_[10260]_ ,
    \new_[10261]_ , \new_[10265]_ , \new_[10266]_ , \new_[10269]_ ,
    \new_[10272]_ , \new_[10273]_ , \new_[10274]_ , \new_[10278]_ ,
    \new_[10279]_ , \new_[10282]_ , \new_[10285]_ , \new_[10286]_ ,
    \new_[10287]_ , \new_[10291]_ , \new_[10292]_ , \new_[10295]_ ,
    \new_[10298]_ , \new_[10299]_ , \new_[10300]_ , \new_[10304]_ ,
    \new_[10305]_ , \new_[10308]_ , \new_[10311]_ , \new_[10312]_ ,
    \new_[10313]_ , \new_[10317]_ , \new_[10318]_ , \new_[10321]_ ,
    \new_[10324]_ , \new_[10325]_ , \new_[10326]_ , \new_[10330]_ ,
    \new_[10331]_ , \new_[10334]_ , \new_[10337]_ , \new_[10338]_ ,
    \new_[10339]_ , \new_[10343]_ , \new_[10344]_ , \new_[10347]_ ,
    \new_[10350]_ , \new_[10351]_ , \new_[10352]_ , \new_[10356]_ ,
    \new_[10357]_ , \new_[10360]_ , \new_[10363]_ , \new_[10364]_ ,
    \new_[10365]_ , \new_[10369]_ , \new_[10370]_ , \new_[10373]_ ,
    \new_[10376]_ , \new_[10377]_ , \new_[10378]_ , \new_[10382]_ ,
    \new_[10383]_ , \new_[10386]_ , \new_[10389]_ , \new_[10390]_ ,
    \new_[10391]_ , \new_[10395]_ , \new_[10396]_ , \new_[10399]_ ,
    \new_[10402]_ , \new_[10403]_ , \new_[10404]_ , \new_[10408]_ ,
    \new_[10409]_ , \new_[10412]_ , \new_[10415]_ , \new_[10416]_ ,
    \new_[10417]_ , \new_[10421]_ , \new_[10422]_ , \new_[10425]_ ,
    \new_[10428]_ , \new_[10429]_ , \new_[10430]_ , \new_[10434]_ ,
    \new_[10435]_ , \new_[10438]_ , \new_[10441]_ , \new_[10442]_ ,
    \new_[10443]_ , \new_[10447]_ , \new_[10448]_ , \new_[10451]_ ,
    \new_[10454]_ , \new_[10455]_ , \new_[10456]_ , \new_[10460]_ ,
    \new_[10461]_ , \new_[10464]_ , \new_[10467]_ , \new_[10468]_ ,
    \new_[10469]_ , \new_[10473]_ , \new_[10474]_ , \new_[10477]_ ,
    \new_[10480]_ , \new_[10481]_ , \new_[10482]_ , \new_[10486]_ ,
    \new_[10487]_ , \new_[10490]_ , \new_[10493]_ , \new_[10494]_ ,
    \new_[10495]_ , \new_[10498]_ , \new_[10501]_ , \new_[10502]_ ,
    \new_[10505]_ , \new_[10508]_ , \new_[10509]_ , \new_[10510]_ ,
    \new_[10514]_ , \new_[10515]_ , \new_[10518]_ , \new_[10521]_ ,
    \new_[10522]_ , \new_[10523]_ , \new_[10526]_ , \new_[10529]_ ,
    \new_[10530]_ , \new_[10533]_ , \new_[10536]_ , \new_[10537]_ ,
    \new_[10538]_ , \new_[10542]_ , \new_[10543]_ , \new_[10546]_ ,
    \new_[10549]_ , \new_[10550]_ , \new_[10551]_ , \new_[10554]_ ,
    \new_[10557]_ , \new_[10558]_ , \new_[10561]_ , \new_[10564]_ ,
    \new_[10565]_ , \new_[10566]_ , \new_[10570]_ , \new_[10571]_ ,
    \new_[10574]_ , \new_[10577]_ , \new_[10578]_ , \new_[10579]_ ,
    \new_[10582]_ , \new_[10585]_ , \new_[10586]_ , \new_[10589]_ ,
    \new_[10592]_ , \new_[10593]_ , \new_[10594]_ , \new_[10598]_ ,
    \new_[10599]_ , \new_[10602]_ , \new_[10605]_ , \new_[10606]_ ,
    \new_[10607]_ , \new_[10610]_ , \new_[10613]_ , \new_[10614]_ ,
    \new_[10617]_ , \new_[10620]_ , \new_[10621]_ , \new_[10622]_ ,
    \new_[10626]_ , \new_[10627]_ , \new_[10630]_ , \new_[10633]_ ,
    \new_[10634]_ , \new_[10635]_ , \new_[10638]_ , \new_[10641]_ ,
    \new_[10642]_ , \new_[10645]_ , \new_[10648]_ , \new_[10649]_ ,
    \new_[10650]_ , \new_[10654]_ , \new_[10655]_ , \new_[10658]_ ,
    \new_[10661]_ , \new_[10662]_ , \new_[10663]_ , \new_[10666]_ ,
    \new_[10669]_ , \new_[10670]_ , \new_[10673]_ , \new_[10676]_ ,
    \new_[10677]_ , \new_[10678]_ , \new_[10682]_ , \new_[10683]_ ,
    \new_[10686]_ , \new_[10689]_ , \new_[10690]_ , \new_[10691]_ ,
    \new_[10694]_ , \new_[10697]_ , \new_[10698]_ , \new_[10701]_ ,
    \new_[10704]_ , \new_[10705]_ , \new_[10706]_ , \new_[10710]_ ,
    \new_[10711]_ , \new_[10714]_ , \new_[10717]_ , \new_[10718]_ ,
    \new_[10719]_ , \new_[10722]_ , \new_[10725]_ , \new_[10726]_ ,
    \new_[10729]_ , \new_[10732]_ , \new_[10733]_ , \new_[10734]_ ,
    \new_[10738]_ , \new_[10739]_ , \new_[10742]_ , \new_[10745]_ ,
    \new_[10746]_ , \new_[10747]_ , \new_[10750]_ , \new_[10753]_ ,
    \new_[10754]_ , \new_[10757]_ , \new_[10760]_ , \new_[10761]_ ,
    \new_[10762]_ , \new_[10766]_ , \new_[10767]_ , \new_[10770]_ ,
    \new_[10773]_ , \new_[10774]_ , \new_[10775]_ , \new_[10778]_ ,
    \new_[10781]_ , \new_[10782]_ , \new_[10785]_ , \new_[10788]_ ,
    \new_[10789]_ , \new_[10790]_ , \new_[10794]_ , \new_[10795]_ ,
    \new_[10798]_ , \new_[10801]_ , \new_[10802]_ , \new_[10803]_ ,
    \new_[10806]_ , \new_[10809]_ , \new_[10810]_ , \new_[10813]_ ,
    \new_[10816]_ , \new_[10817]_ , \new_[10818]_ , \new_[10822]_ ,
    \new_[10823]_ , \new_[10826]_ , \new_[10829]_ , \new_[10830]_ ,
    \new_[10831]_ , \new_[10834]_ , \new_[10837]_ , \new_[10838]_ ,
    \new_[10841]_ , \new_[10844]_ , \new_[10845]_ , \new_[10846]_ ,
    \new_[10850]_ , \new_[10851]_ , \new_[10854]_ , \new_[10857]_ ,
    \new_[10858]_ , \new_[10859]_ , \new_[10862]_ , \new_[10865]_ ,
    \new_[10866]_ , \new_[10869]_ , \new_[10872]_ , \new_[10873]_ ,
    \new_[10874]_ , \new_[10878]_ , \new_[10879]_ , \new_[10882]_ ,
    \new_[10885]_ , \new_[10886]_ , \new_[10887]_ , \new_[10890]_ ,
    \new_[10893]_ , \new_[10894]_ , \new_[10897]_ , \new_[10900]_ ,
    \new_[10901]_ , \new_[10902]_ , \new_[10906]_ , \new_[10907]_ ,
    \new_[10910]_ , \new_[10913]_ , \new_[10914]_ , \new_[10915]_ ,
    \new_[10918]_ , \new_[10921]_ , \new_[10922]_ , \new_[10925]_ ,
    \new_[10928]_ , \new_[10929]_ , \new_[10930]_ , \new_[10934]_ ,
    \new_[10935]_ , \new_[10938]_ , \new_[10941]_ , \new_[10942]_ ,
    \new_[10943]_ , \new_[10946]_ , \new_[10949]_ , \new_[10950]_ ,
    \new_[10953]_ , \new_[10956]_ , \new_[10957]_ , \new_[10958]_ ,
    \new_[10962]_ , \new_[10963]_ , \new_[10966]_ , \new_[10969]_ ,
    \new_[10970]_ , \new_[10971]_ , \new_[10974]_ , \new_[10977]_ ,
    \new_[10978]_ , \new_[10981]_ , \new_[10984]_ , \new_[10985]_ ,
    \new_[10986]_ , \new_[10990]_ , \new_[10991]_ , \new_[10994]_ ,
    \new_[10997]_ , \new_[10998]_ , \new_[10999]_ , \new_[11002]_ ,
    \new_[11005]_ , \new_[11006]_ , \new_[11009]_ , \new_[11012]_ ,
    \new_[11013]_ , \new_[11014]_ , \new_[11018]_ , \new_[11019]_ ,
    \new_[11022]_ , \new_[11025]_ , \new_[11026]_ , \new_[11027]_ ,
    \new_[11030]_ , \new_[11033]_ , \new_[11034]_ , \new_[11037]_ ,
    \new_[11040]_ , \new_[11041]_ , \new_[11042]_ , \new_[11046]_ ,
    \new_[11047]_ , \new_[11050]_ , \new_[11053]_ , \new_[11054]_ ,
    \new_[11055]_ , \new_[11058]_ , \new_[11061]_ , \new_[11062]_ ,
    \new_[11065]_ , \new_[11068]_ , \new_[11069]_ , \new_[11070]_ ,
    \new_[11074]_ , \new_[11075]_ , \new_[11078]_ , \new_[11081]_ ,
    \new_[11082]_ , \new_[11083]_ , \new_[11086]_ , \new_[11089]_ ,
    \new_[11090]_ , \new_[11093]_ , \new_[11096]_ , \new_[11097]_ ,
    \new_[11098]_ , \new_[11102]_ , \new_[11103]_ , \new_[11106]_ ,
    \new_[11109]_ , \new_[11110]_ , \new_[11111]_ , \new_[11114]_ ,
    \new_[11117]_ , \new_[11118]_ , \new_[11121]_ , \new_[11124]_ ,
    \new_[11125]_ , \new_[11126]_ , \new_[11130]_ , \new_[11131]_ ,
    \new_[11134]_ , \new_[11137]_ , \new_[11138]_ , \new_[11139]_ ,
    \new_[11142]_ , \new_[11145]_ , \new_[11146]_ , \new_[11149]_ ,
    \new_[11152]_ , \new_[11153]_ , \new_[11154]_ , \new_[11158]_ ,
    \new_[11159]_ , \new_[11162]_ , \new_[11165]_ , \new_[11166]_ ,
    \new_[11167]_ , \new_[11170]_ , \new_[11173]_ , \new_[11174]_ ,
    \new_[11177]_ , \new_[11180]_ , \new_[11181]_ , \new_[11182]_ ,
    \new_[11186]_ , \new_[11187]_ , \new_[11190]_ , \new_[11193]_ ,
    \new_[11194]_ , \new_[11195]_ , \new_[11198]_ , \new_[11201]_ ,
    \new_[11202]_ , \new_[11205]_ , \new_[11208]_ , \new_[11209]_ ,
    \new_[11210]_ , \new_[11214]_ , \new_[11215]_ , \new_[11218]_ ,
    \new_[11221]_ , \new_[11222]_ , \new_[11223]_ , \new_[11226]_ ,
    \new_[11229]_ , \new_[11230]_ , \new_[11233]_ , \new_[11236]_ ,
    \new_[11237]_ , \new_[11238]_ , \new_[11242]_ , \new_[11243]_ ,
    \new_[11246]_ , \new_[11249]_ , \new_[11250]_ , \new_[11251]_ ,
    \new_[11254]_ , \new_[11257]_ , \new_[11258]_ , \new_[11261]_ ,
    \new_[11264]_ , \new_[11265]_ , \new_[11266]_ , \new_[11270]_ ,
    \new_[11271]_ , \new_[11274]_ , \new_[11277]_ , \new_[11278]_ ,
    \new_[11279]_ , \new_[11282]_ , \new_[11285]_ , \new_[11286]_ ,
    \new_[11289]_ , \new_[11292]_ , \new_[11293]_ , \new_[11294]_ ,
    \new_[11298]_ , \new_[11299]_ , \new_[11302]_ , \new_[11305]_ ,
    \new_[11306]_ , \new_[11307]_ , \new_[11310]_ , \new_[11313]_ ,
    \new_[11314]_ , \new_[11317]_ , \new_[11320]_ , \new_[11321]_ ,
    \new_[11322]_ , \new_[11326]_ , \new_[11327]_ , \new_[11330]_ ,
    \new_[11333]_ , \new_[11334]_ , \new_[11335]_ , \new_[11338]_ ,
    \new_[11341]_ , \new_[11342]_ , \new_[11345]_ , \new_[11348]_ ,
    \new_[11349]_ , \new_[11350]_ , \new_[11354]_ , \new_[11355]_ ,
    \new_[11358]_ , \new_[11361]_ , \new_[11362]_ , \new_[11363]_ ,
    \new_[11366]_ , \new_[11369]_ , \new_[11370]_ , \new_[11373]_ ,
    \new_[11376]_ , \new_[11377]_ , \new_[11378]_ ;
  assign A108 = \new_[1366]_  | \new_[911]_ ;
  assign \new_[1]_  = \new_[11378]_  & \new_[11363]_ ;
  assign \new_[2]_  = \new_[11350]_  & \new_[11335]_ ;
  assign \new_[3]_  = \new_[11322]_  & \new_[11307]_ ;
  assign \new_[4]_  = \new_[11294]_  & \new_[11279]_ ;
  assign \new_[5]_  = \new_[11266]_  & \new_[11251]_ ;
  assign \new_[6]_  = \new_[11238]_  & \new_[11223]_ ;
  assign \new_[7]_  = \new_[11210]_  & \new_[11195]_ ;
  assign \new_[8]_  = \new_[11182]_  & \new_[11167]_ ;
  assign \new_[9]_  = \new_[11154]_  & \new_[11139]_ ;
  assign \new_[10]_  = \new_[11126]_  & \new_[11111]_ ;
  assign \new_[11]_  = \new_[11098]_  & \new_[11083]_ ;
  assign \new_[12]_  = \new_[11070]_  & \new_[11055]_ ;
  assign \new_[13]_  = \new_[11042]_  & \new_[11027]_ ;
  assign \new_[14]_  = \new_[11014]_  & \new_[10999]_ ;
  assign \new_[15]_  = \new_[10986]_  & \new_[10971]_ ;
  assign \new_[16]_  = \new_[10958]_  & \new_[10943]_ ;
  assign \new_[17]_  = \new_[10930]_  & \new_[10915]_ ;
  assign \new_[18]_  = \new_[10902]_  & \new_[10887]_ ;
  assign \new_[19]_  = \new_[10874]_  & \new_[10859]_ ;
  assign \new_[20]_  = \new_[10846]_  & \new_[10831]_ ;
  assign \new_[21]_  = \new_[10818]_  & \new_[10803]_ ;
  assign \new_[22]_  = \new_[10790]_  & \new_[10775]_ ;
  assign \new_[23]_  = \new_[10762]_  & \new_[10747]_ ;
  assign \new_[24]_  = \new_[10734]_  & \new_[10719]_ ;
  assign \new_[25]_  = \new_[10706]_  & \new_[10691]_ ;
  assign \new_[26]_  = \new_[10678]_  & \new_[10663]_ ;
  assign \new_[27]_  = \new_[10650]_  & \new_[10635]_ ;
  assign \new_[28]_  = \new_[10622]_  & \new_[10607]_ ;
  assign \new_[29]_  = \new_[10594]_  & \new_[10579]_ ;
  assign \new_[30]_  = \new_[10566]_  & \new_[10551]_ ;
  assign \new_[31]_  = \new_[10538]_  & \new_[10523]_ ;
  assign \new_[32]_  = \new_[10510]_  & \new_[10495]_ ;
  assign \new_[33]_  = \new_[10482]_  & \new_[10469]_ ;
  assign \new_[34]_  = \new_[10456]_  & \new_[10443]_ ;
  assign \new_[35]_  = \new_[10430]_  & \new_[10417]_ ;
  assign \new_[36]_  = \new_[10404]_  & \new_[10391]_ ;
  assign \new_[37]_  = \new_[10378]_  & \new_[10365]_ ;
  assign \new_[38]_  = \new_[10352]_  & \new_[10339]_ ;
  assign \new_[39]_  = \new_[10326]_  & \new_[10313]_ ;
  assign \new_[40]_  = \new_[10300]_  & \new_[10287]_ ;
  assign \new_[41]_  = \new_[10274]_  & \new_[10261]_ ;
  assign \new_[42]_  = \new_[10248]_  & \new_[10235]_ ;
  assign \new_[43]_  = \new_[10222]_  & \new_[10209]_ ;
  assign \new_[44]_  = \new_[10196]_  & \new_[10183]_ ;
  assign \new_[45]_  = \new_[10170]_  & \new_[10157]_ ;
  assign \new_[46]_  = \new_[10144]_  & \new_[10131]_ ;
  assign \new_[47]_  = \new_[10118]_  & \new_[10105]_ ;
  assign \new_[48]_  = \new_[10092]_  & \new_[10079]_ ;
  assign \new_[49]_  = \new_[10066]_  & \new_[10053]_ ;
  assign \new_[50]_  = \new_[10040]_  & \new_[10027]_ ;
  assign \new_[51]_  = \new_[10014]_  & \new_[10001]_ ;
  assign \new_[52]_  = \new_[9988]_  & \new_[9975]_ ;
  assign \new_[53]_  = \new_[9962]_  & \new_[9949]_ ;
  assign \new_[54]_  = \new_[9936]_  & \new_[9923]_ ;
  assign \new_[55]_  = \new_[9910]_  & \new_[9897]_ ;
  assign \new_[56]_  = \new_[9884]_  & \new_[9871]_ ;
  assign \new_[57]_  = \new_[9858]_  & \new_[9845]_ ;
  assign \new_[58]_  = \new_[9832]_  & \new_[9819]_ ;
  assign \new_[59]_  = \new_[9806]_  & \new_[9793]_ ;
  assign \new_[60]_  = \new_[9780]_  & \new_[9767]_ ;
  assign \new_[61]_  = \new_[9754]_  & \new_[9741]_ ;
  assign \new_[62]_  = \new_[9728]_  & \new_[9715]_ ;
  assign \new_[63]_  = \new_[9702]_  & \new_[9689]_ ;
  assign \new_[64]_  = \new_[9676]_  & \new_[9663]_ ;
  assign \new_[65]_  = \new_[9650]_  & \new_[9637]_ ;
  assign \new_[66]_  = \new_[9624]_  & \new_[9611]_ ;
  assign \new_[67]_  = \new_[9598]_  & \new_[9585]_ ;
  assign \new_[68]_  = \new_[9572]_  & \new_[9559]_ ;
  assign \new_[69]_  = \new_[9546]_  & \new_[9533]_ ;
  assign \new_[70]_  = \new_[9520]_  & \new_[9507]_ ;
  assign \new_[71]_  = \new_[9494]_  & \new_[9481]_ ;
  assign \new_[72]_  = \new_[9468]_  & \new_[9455]_ ;
  assign \new_[73]_  = \new_[9442]_  & \new_[9429]_ ;
  assign \new_[74]_  = \new_[9416]_  & \new_[9403]_ ;
  assign \new_[75]_  = \new_[9390]_  & \new_[9377]_ ;
  assign \new_[76]_  = \new_[9364]_  & \new_[9351]_ ;
  assign \new_[77]_  = \new_[9338]_  & \new_[9325]_ ;
  assign \new_[78]_  = \new_[9312]_  & \new_[9299]_ ;
  assign \new_[79]_  = \new_[9286]_  & \new_[9273]_ ;
  assign \new_[80]_  = \new_[9260]_  & \new_[9247]_ ;
  assign \new_[81]_  = \new_[9234]_  & \new_[9221]_ ;
  assign \new_[82]_  = \new_[9208]_  & \new_[9195]_ ;
  assign \new_[83]_  = \new_[9182]_  & \new_[9169]_ ;
  assign \new_[84]_  = \new_[9156]_  & \new_[9143]_ ;
  assign \new_[85]_  = \new_[9130]_  & \new_[9117]_ ;
  assign \new_[86]_  = \new_[9104]_  & \new_[9091]_ ;
  assign \new_[87]_  = \new_[9078]_  & \new_[9065]_ ;
  assign \new_[88]_  = \new_[9052]_  & \new_[9039]_ ;
  assign \new_[89]_  = \new_[9026]_  & \new_[9013]_ ;
  assign \new_[90]_  = \new_[9000]_  & \new_[8987]_ ;
  assign \new_[91]_  = \new_[8974]_  & \new_[8961]_ ;
  assign \new_[92]_  = \new_[8948]_  & \new_[8935]_ ;
  assign \new_[93]_  = \new_[8922]_  & \new_[8909]_ ;
  assign \new_[94]_  = \new_[8896]_  & \new_[8883]_ ;
  assign \new_[95]_  = \new_[8870]_  & \new_[8857]_ ;
  assign \new_[96]_  = \new_[8844]_  & \new_[8831]_ ;
  assign \new_[97]_  = \new_[8818]_  & \new_[8805]_ ;
  assign \new_[98]_  = \new_[8792]_  & \new_[8779]_ ;
  assign \new_[99]_  = \new_[8766]_  & \new_[8753]_ ;
  assign \new_[100]_  = \new_[8740]_  & \new_[8727]_ ;
  assign \new_[101]_  = \new_[8714]_  & \new_[8701]_ ;
  assign \new_[102]_  = \new_[8688]_  & \new_[8675]_ ;
  assign \new_[103]_  = \new_[8662]_  & \new_[8649]_ ;
  assign \new_[104]_  = \new_[8636]_  & \new_[8623]_ ;
  assign \new_[105]_  = \new_[8610]_  & \new_[8597]_ ;
  assign \new_[106]_  = \new_[8584]_  & \new_[8571]_ ;
  assign \new_[107]_  = \new_[8558]_  & \new_[8545]_ ;
  assign \new_[108]_  = \new_[8532]_  & \new_[8519]_ ;
  assign \new_[109]_  = \new_[8506]_  & \new_[8493]_ ;
  assign \new_[110]_  = \new_[8480]_  & \new_[8467]_ ;
  assign \new_[111]_  = \new_[8454]_  & \new_[8441]_ ;
  assign \new_[112]_  = \new_[8428]_  & \new_[8415]_ ;
  assign \new_[113]_  = \new_[8402]_  & \new_[8389]_ ;
  assign \new_[114]_  = \new_[8376]_  & \new_[8363]_ ;
  assign \new_[115]_  = \new_[8350]_  & \new_[8337]_ ;
  assign \new_[116]_  = \new_[8324]_  & \new_[8311]_ ;
  assign \new_[117]_  = \new_[8298]_  & \new_[8285]_ ;
  assign \new_[118]_  = \new_[8272]_  & \new_[8259]_ ;
  assign \new_[119]_  = \new_[8246]_  & \new_[8233]_ ;
  assign \new_[120]_  = \new_[8220]_  & \new_[8207]_ ;
  assign \new_[121]_  = \new_[8194]_  & \new_[8181]_ ;
  assign \new_[122]_  = \new_[8168]_  & \new_[8155]_ ;
  assign \new_[123]_  = \new_[8142]_  & \new_[8129]_ ;
  assign \new_[124]_  = \new_[8116]_  & \new_[8103]_ ;
  assign \new_[125]_  = \new_[8090]_  & \new_[8077]_ ;
  assign \new_[126]_  = \new_[8064]_  & \new_[8051]_ ;
  assign \new_[127]_  = \new_[8038]_  & \new_[8025]_ ;
  assign \new_[128]_  = \new_[8012]_  & \new_[7999]_ ;
  assign \new_[129]_  = \new_[7986]_  & \new_[7973]_ ;
  assign \new_[130]_  = \new_[7962]_  & \new_[7949]_ ;
  assign \new_[131]_  = \new_[7938]_  & \new_[7925]_ ;
  assign \new_[132]_  = \new_[7914]_  & \new_[7901]_ ;
  assign \new_[133]_  = \new_[7890]_  & \new_[7877]_ ;
  assign \new_[134]_  = \new_[7866]_  & \new_[7853]_ ;
  assign \new_[135]_  = \new_[7842]_  & \new_[7829]_ ;
  assign \new_[136]_  = \new_[7818]_  & \new_[7805]_ ;
  assign \new_[137]_  = \new_[7794]_  & \new_[7781]_ ;
  assign \new_[138]_  = \new_[7770]_  & \new_[7757]_ ;
  assign \new_[139]_  = \new_[7746]_  & \new_[7733]_ ;
  assign \new_[140]_  = \new_[7722]_  & \new_[7709]_ ;
  assign \new_[141]_  = \new_[7698]_  & \new_[7685]_ ;
  assign \new_[142]_  = \new_[7674]_  & \new_[7661]_ ;
  assign \new_[143]_  = \new_[7650]_  & \new_[7637]_ ;
  assign \new_[144]_  = \new_[7626]_  & \new_[7613]_ ;
  assign \new_[145]_  = \new_[7602]_  & \new_[7589]_ ;
  assign \new_[146]_  = \new_[7578]_  & \new_[7565]_ ;
  assign \new_[147]_  = \new_[7554]_  & \new_[7541]_ ;
  assign \new_[148]_  = \new_[7530]_  & \new_[7517]_ ;
  assign \new_[149]_  = \new_[7506]_  & \new_[7493]_ ;
  assign \new_[150]_  = \new_[7482]_  & \new_[7469]_ ;
  assign \new_[151]_  = \new_[7458]_  & \new_[7445]_ ;
  assign \new_[152]_  = \new_[7434]_  & \new_[7421]_ ;
  assign \new_[153]_  = \new_[7410]_  & \new_[7397]_ ;
  assign \new_[154]_  = \new_[7386]_  & \new_[7373]_ ;
  assign \new_[155]_  = \new_[7362]_  & \new_[7349]_ ;
  assign \new_[156]_  = \new_[7338]_  & \new_[7325]_ ;
  assign \new_[157]_  = \new_[7314]_  & \new_[7301]_ ;
  assign \new_[158]_  = \new_[7290]_  & \new_[7277]_ ;
  assign \new_[159]_  = \new_[7266]_  & \new_[7253]_ ;
  assign \new_[160]_  = \new_[7242]_  & \new_[7229]_ ;
  assign \new_[161]_  = \new_[7218]_  & \new_[7205]_ ;
  assign \new_[162]_  = \new_[7194]_  & \new_[7181]_ ;
  assign \new_[163]_  = \new_[7170]_  & \new_[7157]_ ;
  assign \new_[164]_  = \new_[7146]_  & \new_[7133]_ ;
  assign \new_[165]_  = \new_[7122]_  & \new_[7109]_ ;
  assign \new_[166]_  = \new_[7098]_  & \new_[7085]_ ;
  assign \new_[167]_  = \new_[7074]_  & \new_[7061]_ ;
  assign \new_[168]_  = \new_[7050]_  & \new_[7037]_ ;
  assign \new_[169]_  = \new_[7026]_  & \new_[7013]_ ;
  assign \new_[170]_  = \new_[7002]_  & \new_[6989]_ ;
  assign \new_[171]_  = \new_[6978]_  & \new_[6965]_ ;
  assign \new_[172]_  = \new_[6954]_  & \new_[6941]_ ;
  assign \new_[173]_  = \new_[6930]_  & \new_[6917]_ ;
  assign \new_[174]_  = \new_[6906]_  & \new_[6893]_ ;
  assign \new_[175]_  = \new_[6882]_  & \new_[6869]_ ;
  assign \new_[176]_  = \new_[6858]_  & \new_[6845]_ ;
  assign \new_[177]_  = \new_[6834]_  & \new_[6823]_ ;
  assign \new_[178]_  = \new_[6812]_  & \new_[6801]_ ;
  assign \new_[179]_  = \new_[6790]_  & \new_[6779]_ ;
  assign \new_[180]_  = \new_[6768]_  & \new_[6757]_ ;
  assign \new_[181]_  = \new_[6746]_  & \new_[6735]_ ;
  assign \new_[182]_  = \new_[6724]_  & \new_[6713]_ ;
  assign \new_[183]_  = \new_[6702]_  & \new_[6691]_ ;
  assign \new_[184]_  = \new_[6680]_  & \new_[6669]_ ;
  assign \new_[185]_  = \new_[6658]_  & \new_[6647]_ ;
  assign \new_[186]_  = \new_[6636]_  & \new_[6625]_ ;
  assign \new_[187]_  = \new_[6614]_  & \new_[6603]_ ;
  assign \new_[188]_  = \new_[6592]_  & \new_[6581]_ ;
  assign \new_[189]_  = \new_[6570]_  & \new_[6559]_ ;
  assign \new_[190]_  = \new_[6548]_  & \new_[6537]_ ;
  assign \new_[191]_  = \new_[6526]_  & \new_[6515]_ ;
  assign \new_[192]_  = \new_[6504]_  & \new_[6493]_ ;
  assign \new_[193]_  = \new_[6482]_  & \new_[6471]_ ;
  assign \new_[194]_  = \new_[6460]_  & \new_[6449]_ ;
  assign \new_[195]_  = \new_[6438]_  & \new_[6427]_ ;
  assign \new_[196]_  = \new_[6416]_  & \new_[6405]_ ;
  assign \new_[197]_  = \new_[6394]_  & \new_[6383]_ ;
  assign \new_[198]_  = \new_[6372]_  & \new_[6361]_ ;
  assign \new_[199]_  = \new_[6350]_  & \new_[6339]_ ;
  assign \new_[200]_  = \new_[6328]_  & \new_[6317]_ ;
  assign \new_[201]_  = \new_[6306]_  & \new_[6295]_ ;
  assign \new_[202]_  = \new_[6284]_  & \new_[6273]_ ;
  assign \new_[203]_  = \new_[6262]_  & \new_[6251]_ ;
  assign \new_[204]_  = \new_[6240]_  & \new_[6229]_ ;
  assign \new_[205]_  = \new_[6218]_  & \new_[6207]_ ;
  assign \new_[206]_  = \new_[6196]_  & \new_[6185]_ ;
  assign \new_[207]_  = \new_[6174]_  & \new_[6163]_ ;
  assign \new_[208]_  = \new_[6152]_  & \new_[6141]_ ;
  assign \new_[209]_  = \new_[6130]_  & \new_[6119]_ ;
  assign \new_[210]_  = \new_[6108]_  & \new_[6097]_ ;
  assign \new_[211]_  = \new_[6086]_  & \new_[6075]_ ;
  assign \new_[212]_  = \new_[6064]_  & \new_[6053]_ ;
  assign \new_[213]_  = \new_[6042]_  & \new_[6031]_ ;
  assign \new_[214]_  = \new_[6020]_  & \new_[6009]_ ;
  assign \new_[215]_  = \new_[5998]_  & \new_[5987]_ ;
  assign \new_[216]_  = \new_[5976]_  & \new_[5965]_ ;
  assign \new_[217]_  = \new_[5954]_  & \new_[5943]_ ;
  assign \new_[218]_  = \new_[5932]_  & \new_[5921]_ ;
  assign \new_[219]_  = \new_[5910]_  & \new_[5899]_ ;
  assign \new_[220]_  = \new_[5888]_  & \new_[5877]_ ;
  assign \new_[221]_  = \new_[5866]_  & \new_[5855]_ ;
  assign \new_[222]_  = \new_[5844]_  & \new_[5833]_ ;
  assign \new_[223]_  = \new_[5822]_  & \new_[5811]_ ;
  assign \new_[224]_  = \new_[5800]_  & \new_[5789]_ ;
  assign \new_[225]_  = \new_[5778]_  & \new_[5767]_ ;
  assign \new_[226]_  = \new_[5756]_  & \new_[5745]_ ;
  assign \new_[227]_  = \new_[5734]_  & \new_[5723]_ ;
  assign \new_[228]_  = \new_[5712]_  & \new_[5701]_ ;
  assign \new_[229]_  = \new_[5690]_  & \new_[5679]_ ;
  assign \new_[230]_  = \new_[5668]_  & \new_[5657]_ ;
  assign \new_[231]_  = \new_[5646]_  & \new_[5635]_ ;
  assign \new_[232]_  = \new_[5624]_  & \new_[5613]_ ;
  assign \new_[233]_  = \new_[5602]_  & \new_[5591]_ ;
  assign \new_[234]_  = \new_[5580]_  & \new_[5569]_ ;
  assign \new_[235]_  = \new_[5558]_  & \new_[5547]_ ;
  assign \new_[236]_  = \new_[5536]_  & \new_[5525]_ ;
  assign \new_[237]_  = \new_[5514]_  & \new_[5503]_ ;
  assign \new_[238]_  = \new_[5492]_  & \new_[5481]_ ;
  assign \new_[239]_  = \new_[5470]_  & \new_[5459]_ ;
  assign \new_[240]_  = \new_[5448]_  & \new_[5437]_ ;
  assign \new_[241]_  = \new_[5426]_  & \new_[5415]_ ;
  assign \new_[242]_  = \new_[5404]_  & \new_[5393]_ ;
  assign \new_[243]_  = \new_[5382]_  & \new_[5371]_ ;
  assign \new_[244]_  = \new_[5360]_  & \new_[5349]_ ;
  assign \new_[245]_  = \new_[5338]_  & \new_[5327]_ ;
  assign \new_[246]_  = \new_[5316]_  & \new_[5305]_ ;
  assign \new_[247]_  = \new_[5294]_  & \new_[5283]_ ;
  assign \new_[248]_  = \new_[5272]_  & \new_[5261]_ ;
  assign \new_[249]_  = \new_[5250]_  & \new_[5239]_ ;
  assign \new_[250]_  = \new_[5228]_  & \new_[5217]_ ;
  assign \new_[251]_  = \new_[5206]_  & \new_[5195]_ ;
  assign \new_[252]_  = \new_[5184]_  & \new_[5173]_ ;
  assign \new_[253]_  = \new_[5162]_  & \new_[5151]_ ;
  assign \new_[254]_  = \new_[5140]_  & \new_[5129]_ ;
  assign \new_[255]_  = \new_[5118]_  & \new_[5107]_ ;
  assign \new_[256]_  = \new_[5096]_  & \new_[5085]_ ;
  assign \new_[257]_  = \new_[5074]_  & \new_[5063]_ ;
  assign \new_[258]_  = \new_[5052]_  & \new_[5041]_ ;
  assign \new_[259]_  = \new_[5030]_  & \new_[5019]_ ;
  assign \new_[260]_  = \new_[5008]_  & \new_[4997]_ ;
  assign \new_[261]_  = \new_[4986]_  & \new_[4975]_ ;
  assign \new_[262]_  = \new_[4964]_  & \new_[4953]_ ;
  assign \new_[263]_  = \new_[4942]_  & \new_[4931]_ ;
  assign \new_[264]_  = \new_[4920]_  & \new_[4909]_ ;
  assign \new_[265]_  = \new_[4898]_  & \new_[4887]_ ;
  assign \new_[266]_  = \new_[4876]_  & \new_[4865]_ ;
  assign \new_[267]_  = \new_[4854]_  & \new_[4843]_ ;
  assign \new_[268]_  = \new_[4832]_  & \new_[4821]_ ;
  assign \new_[269]_  = \new_[4810]_  & \new_[4799]_ ;
  assign \new_[270]_  = \new_[4788]_  & \new_[4777]_ ;
  assign \new_[271]_  = \new_[4766]_  & \new_[4755]_ ;
  assign \new_[272]_  = \new_[4744]_  & \new_[4733]_ ;
  assign \new_[273]_  = \new_[4722]_  & \new_[4711]_ ;
  assign \new_[274]_  = \new_[4700]_  & \new_[4689]_ ;
  assign \new_[275]_  = \new_[4678]_  & \new_[4667]_ ;
  assign \new_[276]_  = \new_[4656]_  & \new_[4645]_ ;
  assign \new_[277]_  = \new_[4634]_  & \new_[4623]_ ;
  assign \new_[278]_  = \new_[4612]_  & \new_[4601]_ ;
  assign \new_[279]_  = \new_[4590]_  & \new_[4579]_ ;
  assign \new_[280]_  = \new_[4568]_  & \new_[4557]_ ;
  assign \new_[281]_  = \new_[4546]_  & \new_[4535]_ ;
  assign \new_[282]_  = \new_[4524]_  & \new_[4513]_ ;
  assign \new_[283]_  = \new_[4502]_  & \new_[4491]_ ;
  assign \new_[284]_  = \new_[4480]_  & \new_[4469]_ ;
  assign \new_[285]_  = \new_[4458]_  & \new_[4447]_ ;
  assign \new_[286]_  = \new_[4436]_  & \new_[4425]_ ;
  assign \new_[287]_  = \new_[4414]_  & \new_[4403]_ ;
  assign \new_[288]_  = \new_[4392]_  & \new_[4381]_ ;
  assign \new_[289]_  = \new_[4370]_  & \new_[4359]_ ;
  assign \new_[290]_  = \new_[4348]_  & \new_[4337]_ ;
  assign \new_[291]_  = \new_[4326]_  & \new_[4315]_ ;
  assign \new_[292]_  = \new_[4304]_  & \new_[4293]_ ;
  assign \new_[293]_  = \new_[4282]_  & \new_[4271]_ ;
  assign \new_[294]_  = \new_[4260]_  & \new_[4249]_ ;
  assign \new_[295]_  = \new_[4238]_  & \new_[4227]_ ;
  assign \new_[296]_  = \new_[4216]_  & \new_[4205]_ ;
  assign \new_[297]_  = \new_[4194]_  & \new_[4183]_ ;
  assign \new_[298]_  = \new_[4172]_  & \new_[4161]_ ;
  assign \new_[299]_  = \new_[4150]_  & \new_[4139]_ ;
  assign \new_[300]_  = \new_[4128]_  & \new_[4117]_ ;
  assign \new_[301]_  = \new_[4106]_  & \new_[4095]_ ;
  assign \new_[302]_  = \new_[4084]_  & \new_[4073]_ ;
  assign \new_[303]_  = \new_[4062]_  & \new_[4051]_ ;
  assign \new_[304]_  = \new_[4040]_  & \new_[4029]_ ;
  assign \new_[305]_  = \new_[4018]_  & \new_[4007]_ ;
  assign \new_[306]_  = \new_[3996]_  & \new_[3985]_ ;
  assign \new_[307]_  = \new_[3974]_  & \new_[3963]_ ;
  assign \new_[308]_  = \new_[3952]_  & \new_[3941]_ ;
  assign \new_[309]_  = \new_[3930]_  & \new_[3919]_ ;
  assign \new_[310]_  = \new_[3908]_  & \new_[3897]_ ;
  assign \new_[311]_  = \new_[3886]_  & \new_[3875]_ ;
  assign \new_[312]_  = \new_[3864]_  & \new_[3853]_ ;
  assign \new_[313]_  = \new_[3842]_  & \new_[3831]_ ;
  assign \new_[314]_  = \new_[3820]_  & \new_[3809]_ ;
  assign \new_[315]_  = \new_[3798]_  & \new_[3787]_ ;
  assign \new_[316]_  = \new_[3776]_  & \new_[3765]_ ;
  assign \new_[317]_  = \new_[3754]_  & \new_[3743]_ ;
  assign \new_[318]_  = \new_[3732]_  & \new_[3721]_ ;
  assign \new_[319]_  = \new_[3710]_  & \new_[3699]_ ;
  assign \new_[320]_  = \new_[3688]_  & \new_[3677]_ ;
  assign \new_[321]_  = \new_[3666]_  & \new_[3655]_ ;
  assign \new_[322]_  = \new_[3646]_  & \new_[3635]_ ;
  assign \new_[323]_  = \new_[3626]_  & \new_[3615]_ ;
  assign \new_[324]_  = \new_[3606]_  & \new_[3595]_ ;
  assign \new_[325]_  = \new_[3586]_  & \new_[3575]_ ;
  assign \new_[326]_  = \new_[3566]_  & \new_[3555]_ ;
  assign \new_[327]_  = \new_[3546]_  & \new_[3535]_ ;
  assign \new_[328]_  = \new_[3526]_  & \new_[3515]_ ;
  assign \new_[329]_  = \new_[3506]_  & \new_[3495]_ ;
  assign \new_[330]_  = \new_[3486]_  & \new_[3475]_ ;
  assign \new_[331]_  = \new_[3466]_  & \new_[3455]_ ;
  assign \new_[332]_  = \new_[3446]_  & \new_[3435]_ ;
  assign \new_[333]_  = \new_[3426]_  & \new_[3415]_ ;
  assign \new_[334]_  = \new_[3406]_  & \new_[3395]_ ;
  assign \new_[335]_  = \new_[3386]_  & \new_[3375]_ ;
  assign \new_[336]_  = \new_[3366]_  & \new_[3355]_ ;
  assign \new_[337]_  = \new_[3346]_  & \new_[3335]_ ;
  assign \new_[338]_  = \new_[3326]_  & \new_[3315]_ ;
  assign \new_[339]_  = \new_[3306]_  & \new_[3295]_ ;
  assign \new_[340]_  = \new_[3286]_  & \new_[3275]_ ;
  assign \new_[341]_  = \new_[3266]_  & \new_[3255]_ ;
  assign \new_[342]_  = \new_[3246]_  & \new_[3235]_ ;
  assign \new_[343]_  = \new_[3226]_  & \new_[3215]_ ;
  assign \new_[344]_  = \new_[3206]_  & \new_[3195]_ ;
  assign \new_[345]_  = \new_[3186]_  & \new_[3177]_ ;
  assign \new_[346]_  = \new_[3168]_  & \new_[3159]_ ;
  assign \new_[347]_  = \new_[3150]_  & \new_[3141]_ ;
  assign \new_[348]_  = \new_[3132]_  & \new_[3123]_ ;
  assign \new_[349]_  = \new_[3114]_  & \new_[3105]_ ;
  assign \new_[350]_  = \new_[3096]_  & \new_[3087]_ ;
  assign \new_[351]_  = \new_[3078]_  & \new_[3069]_ ;
  assign \new_[352]_  = \new_[3060]_  & \new_[3051]_ ;
  assign \new_[353]_  = \new_[3042]_  & \new_[3033]_ ;
  assign \new_[354]_  = \new_[3024]_  & \new_[3015]_ ;
  assign \new_[355]_  = \new_[3006]_  & \new_[2997]_ ;
  assign \new_[356]_  = \new_[2988]_  & \new_[2979]_ ;
  assign \new_[357]_  = \new_[2970]_  & \new_[2961]_ ;
  assign \new_[358]_  = \new_[2952]_  & \new_[2943]_ ;
  assign \new_[359]_  = \new_[2934]_  & \new_[2925]_ ;
  assign \new_[360]_  = \new_[2916]_  & \new_[2907]_ ;
  assign \new_[361]_  = \new_[2898]_  & \new_[2889]_ ;
  assign \new_[362]_  = \new_[2880]_  & \new_[2871]_ ;
  assign \new_[363]_  = \new_[2862]_  & \new_[2853]_ ;
  assign \new_[364]_  = \new_[2844]_  & \new_[2835]_ ;
  assign \new_[365]_  = \new_[2826]_  & \new_[2817]_ ;
  assign \new_[366]_  = \new_[2808]_  & \new_[2799]_ ;
  assign \new_[367]_  = \new_[2790]_  & \new_[2781]_ ;
  assign \new_[368]_  = \new_[2772]_  & \new_[2763]_ ;
  assign \new_[369]_  = \new_[2754]_  & \new_[2745]_ ;
  assign \new_[370]_  = \new_[2736]_  & \new_[2727]_ ;
  assign \new_[371]_  = \new_[2718]_  & \new_[2709]_ ;
  assign \new_[372]_  = \new_[2700]_  & \new_[2691]_ ;
  assign \new_[373]_  = \new_[2682]_  & \new_[2673]_ ;
  assign \new_[374]_  = \new_[2664]_  & \new_[2655]_ ;
  assign \new_[375]_  = \new_[2646]_  & \new_[2637]_ ;
  assign \new_[376]_  = \new_[2628]_  & \new_[2619]_ ;
  assign \new_[377]_  = \new_[2610]_  & \new_[2601]_ ;
  assign \new_[378]_  = \new_[2592]_  & \new_[2583]_ ;
  assign \new_[379]_  = \new_[2574]_  & \new_[2565]_ ;
  assign \new_[380]_  = \new_[2556]_  & \new_[2547]_ ;
  assign \new_[381]_  = \new_[2538]_  & \new_[2529]_ ;
  assign \new_[382]_  = \new_[2520]_  & \new_[2511]_ ;
  assign \new_[383]_  = \new_[2502]_  & \new_[2493]_ ;
  assign \new_[384]_  = \new_[2484]_  & \new_[2475]_ ;
  assign \new_[385]_  = \new_[2466]_  & \new_[2457]_ ;
  assign \new_[386]_  = \new_[2448]_  & \new_[2439]_ ;
  assign \new_[387]_  = \new_[2430]_  & \new_[2421]_ ;
  assign \new_[388]_  = \new_[2412]_  & \new_[2403]_ ;
  assign \new_[389]_  = \new_[2394]_  & \new_[2385]_ ;
  assign \new_[390]_  = \new_[2376]_  & \new_[2367]_ ;
  assign \new_[391]_  = \new_[2358]_  & \new_[2349]_ ;
  assign \new_[392]_  = \new_[2340]_  & \new_[2331]_ ;
  assign \new_[393]_  = \new_[2322]_  & \new_[2313]_ ;
  assign \new_[394]_  = \new_[2304]_  & \new_[2295]_ ;
  assign \new_[395]_  = \new_[2286]_  & \new_[2277]_ ;
  assign \new_[396]_  = \new_[2268]_  & \new_[2259]_ ;
  assign \new_[397]_  = \new_[2250]_  & \new_[2241]_ ;
  assign \new_[398]_  = \new_[2232]_  & \new_[2223]_ ;
  assign \new_[399]_  = \new_[2214]_  & \new_[2205]_ ;
  assign \new_[400]_  = \new_[2196]_  & \new_[2187]_ ;
  assign \new_[401]_  = \new_[2178]_  & \new_[2169]_ ;
  assign \new_[402]_  = \new_[2160]_  & \new_[2151]_ ;
  assign \new_[403]_  = \new_[2142]_  & \new_[2133]_ ;
  assign \new_[404]_  = \new_[2124]_  & \new_[2115]_ ;
  assign \new_[405]_  = \new_[2106]_  & \new_[2097]_ ;
  assign \new_[406]_  = \new_[2088]_  & \new_[2079]_ ;
  assign \new_[407]_  = \new_[2070]_  & \new_[2061]_ ;
  assign \new_[408]_  = \new_[2052]_  & \new_[2043]_ ;
  assign \new_[409]_  = \new_[2034]_  & \new_[2025]_ ;
  assign \new_[410]_  = \new_[2016]_  & \new_[2007]_ ;
  assign \new_[411]_  = \new_[1998]_  & \new_[1989]_ ;
  assign \new_[412]_  = \new_[1980]_  & \new_[1971]_ ;
  assign \new_[413]_  = \new_[1962]_  & \new_[1953]_ ;
  assign \new_[414]_  = \new_[1944]_  & \new_[1935]_ ;
  assign \new_[415]_  = \new_[1926]_  & \new_[1917]_ ;
  assign \new_[416]_  = \new_[1908]_  & \new_[1899]_ ;
  assign \new_[417]_  = \new_[1890]_  & \new_[1881]_ ;
  assign \new_[418]_  = \new_[1874]_  & \new_[1865]_ ;
  assign \new_[419]_  = \new_[1858]_  & \new_[1849]_ ;
  assign \new_[420]_  = \new_[1842]_  & \new_[1833]_ ;
  assign \new_[421]_  = \new_[1826]_  & \new_[1819]_ ;
  assign \new_[422]_  = \new_[1812]_  & \new_[1805]_ ;
  assign \new_[423]_  = \new_[1798]_  & \new_[1791]_ ;
  assign \new_[424]_  = \new_[1784]_  & \new_[1777]_ ;
  assign \new_[425]_  = \new_[1770]_  & \new_[1763]_ ;
  assign \new_[426]_  = \new_[1756]_  & \new_[1749]_ ;
  assign \new_[427]_  = \new_[1742]_  & \new_[1735]_ ;
  assign \new_[428]_  = \new_[1728]_  & \new_[1721]_ ;
  assign \new_[429]_  = \new_[1714]_  & \new_[1707]_ ;
  assign \new_[430]_  = \new_[1700]_  & \new_[1693]_ ;
  assign \new_[431]_  = \new_[1686]_  & \new_[1679]_ ;
  assign \new_[432]_  = \new_[1672]_  & \new_[1665]_ ;
  assign \new_[433]_  = \new_[1658]_  & \new_[1651]_ ;
  assign \new_[434]_  = \new_[1644]_  & \new_[1637]_ ;
  assign \new_[435]_  = \new_[1630]_  & \new_[1623]_ ;
  assign \new_[436]_  = \new_[1616]_  & \new_[1609]_ ;
  assign \new_[437]_  = \new_[1602]_  & \new_[1595]_ ;
  assign \new_[438]_  = \new_[1588]_  & \new_[1581]_ ;
  assign \new_[439]_  = \new_[1574]_  & \new_[1567]_ ;
  assign \new_[440]_  = \new_[1560]_  & \new_[1553]_ ;
  assign \new_[441]_  = \new_[1546]_  & \new_[1539]_ ;
  assign \new_[442]_  = \new_[1532]_  & \new_[1525]_ ;
  assign \new_[443]_  = \new_[1518]_  & \new_[1511]_ ;
  assign \new_[444]_  = \new_[1504]_  & \new_[1497]_ ;
  assign \new_[445]_  = \new_[1490]_  & \new_[1483]_ ;
  assign \new_[446]_  = \new_[1478]_  & \new_[1471]_ ;
  assign \new_[447]_  = \new_[1466]_  & \new_[1459]_ ;
  assign \new_[448]_  = \new_[1454]_  & \new_[1447]_ ;
  assign \new_[449]_  = \new_[1442]_  & \new_[1437]_ ;
  assign \new_[450]_  = \new_[1432]_  & \new_[1427]_ ;
  assign \new_[451]_  = \new_[1422]_  & \new_[1417]_ ;
  assign \new_[452]_  = \new_[1412]_  & \new_[1407]_ ;
  assign \new_[453]_  = \new_[1402]_  & \new_[1397]_ ;
  assign \new_[454]_  = \new_[1392]_  & \new_[1387]_ ;
  assign \new_[455]_  = \new_[1382]_  & \new_[1377]_ ;
  assign \new_[456]_  = \new_[1374]_  & \new_[1369]_ ;
  assign \new_[460]_  = \new_[454]_  | \new_[455]_ ;
  assign \new_[461]_  = \new_[456]_  | \new_[460]_ ;
  assign \new_[464]_  = \new_[452]_  | \new_[453]_ ;
  assign \new_[467]_  = \new_[450]_  | \new_[451]_ ;
  assign \new_[468]_  = \new_[467]_  | \new_[464]_ ;
  assign \new_[469]_  = \new_[468]_  | \new_[461]_ ;
  assign \new_[473]_  = \new_[447]_  | \new_[448]_ ;
  assign \new_[474]_  = \new_[449]_  | \new_[473]_ ;
  assign \new_[477]_  = \new_[445]_  | \new_[446]_ ;
  assign \new_[480]_  = \new_[443]_  | \new_[444]_ ;
  assign \new_[481]_  = \new_[480]_  | \new_[477]_ ;
  assign \new_[482]_  = \new_[481]_  | \new_[474]_ ;
  assign \new_[483]_  = \new_[482]_  | \new_[469]_ ;
  assign \new_[487]_  = \new_[440]_  | \new_[441]_ ;
  assign \new_[488]_  = \new_[442]_  | \new_[487]_ ;
  assign \new_[491]_  = \new_[438]_  | \new_[439]_ ;
  assign \new_[494]_  = \new_[436]_  | \new_[437]_ ;
  assign \new_[495]_  = \new_[494]_  | \new_[491]_ ;
  assign \new_[496]_  = \new_[495]_  | \new_[488]_ ;
  assign \new_[500]_  = \new_[433]_  | \new_[434]_ ;
  assign \new_[501]_  = \new_[435]_  | \new_[500]_ ;
  assign \new_[504]_  = \new_[431]_  | \new_[432]_ ;
  assign \new_[507]_  = \new_[429]_  | \new_[430]_ ;
  assign \new_[508]_  = \new_[507]_  | \new_[504]_ ;
  assign \new_[509]_  = \new_[508]_  | \new_[501]_ ;
  assign \new_[510]_  = \new_[509]_  | \new_[496]_ ;
  assign \new_[511]_  = \new_[510]_  | \new_[483]_ ;
  assign \new_[515]_  = \new_[426]_  | \new_[427]_ ;
  assign \new_[516]_  = \new_[428]_  | \new_[515]_ ;
  assign \new_[519]_  = \new_[424]_  | \new_[425]_ ;
  assign \new_[522]_  = \new_[422]_  | \new_[423]_ ;
  assign \new_[523]_  = \new_[522]_  | \new_[519]_ ;
  assign \new_[524]_  = \new_[523]_  | \new_[516]_ ;
  assign \new_[528]_  = \new_[419]_  | \new_[420]_ ;
  assign \new_[529]_  = \new_[421]_  | \new_[528]_ ;
  assign \new_[532]_  = \new_[417]_  | \new_[418]_ ;
  assign \new_[535]_  = \new_[415]_  | \new_[416]_ ;
  assign \new_[536]_  = \new_[535]_  | \new_[532]_ ;
  assign \new_[537]_  = \new_[536]_  | \new_[529]_ ;
  assign \new_[538]_  = \new_[537]_  | \new_[524]_ ;
  assign \new_[542]_  = \new_[412]_  | \new_[413]_ ;
  assign \new_[543]_  = \new_[414]_  | \new_[542]_ ;
  assign \new_[546]_  = \new_[410]_  | \new_[411]_ ;
  assign \new_[549]_  = \new_[408]_  | \new_[409]_ ;
  assign \new_[550]_  = \new_[549]_  | \new_[546]_ ;
  assign \new_[551]_  = \new_[550]_  | \new_[543]_ ;
  assign \new_[554]_  = \new_[406]_  | \new_[407]_ ;
  assign \new_[557]_  = \new_[404]_  | \new_[405]_ ;
  assign \new_[558]_  = \new_[557]_  | \new_[554]_ ;
  assign \new_[561]_  = \new_[402]_  | \new_[403]_ ;
  assign \new_[564]_  = \new_[400]_  | \new_[401]_ ;
  assign \new_[565]_  = \new_[564]_  | \new_[561]_ ;
  assign \new_[566]_  = \new_[565]_  | \new_[558]_ ;
  assign \new_[567]_  = \new_[566]_  | \new_[551]_ ;
  assign \new_[568]_  = \new_[567]_  | \new_[538]_ ;
  assign \new_[569]_  = \new_[568]_  | \new_[511]_ ;
  assign \new_[573]_  = \new_[397]_  | \new_[398]_ ;
  assign \new_[574]_  = \new_[399]_  | \new_[573]_ ;
  assign \new_[577]_  = \new_[395]_  | \new_[396]_ ;
  assign \new_[580]_  = \new_[393]_  | \new_[394]_ ;
  assign \new_[581]_  = \new_[580]_  | \new_[577]_ ;
  assign \new_[582]_  = \new_[581]_  | \new_[574]_ ;
  assign \new_[586]_  = \new_[390]_  | \new_[391]_ ;
  assign \new_[587]_  = \new_[392]_  | \new_[586]_ ;
  assign \new_[590]_  = \new_[388]_  | \new_[389]_ ;
  assign \new_[593]_  = \new_[386]_  | \new_[387]_ ;
  assign \new_[594]_  = \new_[593]_  | \new_[590]_ ;
  assign \new_[595]_  = \new_[594]_  | \new_[587]_ ;
  assign \new_[596]_  = \new_[595]_  | \new_[582]_ ;
  assign \new_[600]_  = \new_[383]_  | \new_[384]_ ;
  assign \new_[601]_  = \new_[385]_  | \new_[600]_ ;
  assign \new_[604]_  = \new_[381]_  | \new_[382]_ ;
  assign \new_[607]_  = \new_[379]_  | \new_[380]_ ;
  assign \new_[608]_  = \new_[607]_  | \new_[604]_ ;
  assign \new_[609]_  = \new_[608]_  | \new_[601]_ ;
  assign \new_[613]_  = \new_[376]_  | \new_[377]_ ;
  assign \new_[614]_  = \new_[378]_  | \new_[613]_ ;
  assign \new_[617]_  = \new_[374]_  | \new_[375]_ ;
  assign \new_[620]_  = \new_[372]_  | \new_[373]_ ;
  assign \new_[621]_  = \new_[620]_  | \new_[617]_ ;
  assign \new_[622]_  = \new_[621]_  | \new_[614]_ ;
  assign \new_[623]_  = \new_[622]_  | \new_[609]_ ;
  assign \new_[624]_  = \new_[623]_  | \new_[596]_ ;
  assign \new_[628]_  = \new_[369]_  | \new_[370]_ ;
  assign \new_[629]_  = \new_[371]_  | \new_[628]_ ;
  assign \new_[632]_  = \new_[367]_  | \new_[368]_ ;
  assign \new_[635]_  = \new_[365]_  | \new_[366]_ ;
  assign \new_[636]_  = \new_[635]_  | \new_[632]_ ;
  assign \new_[637]_  = \new_[636]_  | \new_[629]_ ;
  assign \new_[641]_  = \new_[362]_  | \new_[363]_ ;
  assign \new_[642]_  = \new_[364]_  | \new_[641]_ ;
  assign \new_[645]_  = \new_[360]_  | \new_[361]_ ;
  assign \new_[648]_  = \new_[358]_  | \new_[359]_ ;
  assign \new_[649]_  = \new_[648]_  | \new_[645]_ ;
  assign \new_[650]_  = \new_[649]_  | \new_[642]_ ;
  assign \new_[651]_  = \new_[650]_  | \new_[637]_ ;
  assign \new_[655]_  = \new_[355]_  | \new_[356]_ ;
  assign \new_[656]_  = \new_[357]_  | \new_[655]_ ;
  assign \new_[659]_  = \new_[353]_  | \new_[354]_ ;
  assign \new_[662]_  = \new_[351]_  | \new_[352]_ ;
  assign \new_[663]_  = \new_[662]_  | \new_[659]_ ;
  assign \new_[664]_  = \new_[663]_  | \new_[656]_ ;
  assign \new_[667]_  = \new_[349]_  | \new_[350]_ ;
  assign \new_[670]_  = \new_[347]_  | \new_[348]_ ;
  assign \new_[671]_  = \new_[670]_  | \new_[667]_ ;
  assign \new_[674]_  = \new_[345]_  | \new_[346]_ ;
  assign \new_[677]_  = \new_[343]_  | \new_[344]_ ;
  assign \new_[678]_  = \new_[677]_  | \new_[674]_ ;
  assign \new_[679]_  = \new_[678]_  | \new_[671]_ ;
  assign \new_[680]_  = \new_[679]_  | \new_[664]_ ;
  assign \new_[681]_  = \new_[680]_  | \new_[651]_ ;
  assign \new_[682]_  = \new_[681]_  | \new_[624]_ ;
  assign \new_[683]_  = \new_[682]_  | \new_[569]_ ;
  assign \new_[687]_  = \new_[340]_  | \new_[341]_ ;
  assign \new_[688]_  = \new_[342]_  | \new_[687]_ ;
  assign \new_[691]_  = \new_[338]_  | \new_[339]_ ;
  assign \new_[694]_  = \new_[336]_  | \new_[337]_ ;
  assign \new_[695]_  = \new_[694]_  | \new_[691]_ ;
  assign \new_[696]_  = \new_[695]_  | \new_[688]_ ;
  assign \new_[700]_  = \new_[333]_  | \new_[334]_ ;
  assign \new_[701]_  = \new_[335]_  | \new_[700]_ ;
  assign \new_[704]_  = \new_[331]_  | \new_[332]_ ;
  assign \new_[707]_  = \new_[329]_  | \new_[330]_ ;
  assign \new_[708]_  = \new_[707]_  | \new_[704]_ ;
  assign \new_[709]_  = \new_[708]_  | \new_[701]_ ;
  assign \new_[710]_  = \new_[709]_  | \new_[696]_ ;
  assign \new_[714]_  = \new_[326]_  | \new_[327]_ ;
  assign \new_[715]_  = \new_[328]_  | \new_[714]_ ;
  assign \new_[718]_  = \new_[324]_  | \new_[325]_ ;
  assign \new_[721]_  = \new_[322]_  | \new_[323]_ ;
  assign \new_[722]_  = \new_[721]_  | \new_[718]_ ;
  assign \new_[723]_  = \new_[722]_  | \new_[715]_ ;
  assign \new_[727]_  = \new_[319]_  | \new_[320]_ ;
  assign \new_[728]_  = \new_[321]_  | \new_[727]_ ;
  assign \new_[731]_  = \new_[317]_  | \new_[318]_ ;
  assign \new_[734]_  = \new_[315]_  | \new_[316]_ ;
  assign \new_[735]_  = \new_[734]_  | \new_[731]_ ;
  assign \new_[736]_  = \new_[735]_  | \new_[728]_ ;
  assign \new_[737]_  = \new_[736]_  | \new_[723]_ ;
  assign \new_[738]_  = \new_[737]_  | \new_[710]_ ;
  assign \new_[742]_  = \new_[312]_  | \new_[313]_ ;
  assign \new_[743]_  = \new_[314]_  | \new_[742]_ ;
  assign \new_[746]_  = \new_[310]_  | \new_[311]_ ;
  assign \new_[749]_  = \new_[308]_  | \new_[309]_ ;
  assign \new_[750]_  = \new_[749]_  | \new_[746]_ ;
  assign \new_[751]_  = \new_[750]_  | \new_[743]_ ;
  assign \new_[755]_  = \new_[305]_  | \new_[306]_ ;
  assign \new_[756]_  = \new_[307]_  | \new_[755]_ ;
  assign \new_[759]_  = \new_[303]_  | \new_[304]_ ;
  assign \new_[762]_  = \new_[301]_  | \new_[302]_ ;
  assign \new_[763]_  = \new_[762]_  | \new_[759]_ ;
  assign \new_[764]_  = \new_[763]_  | \new_[756]_ ;
  assign \new_[765]_  = \new_[764]_  | \new_[751]_ ;
  assign \new_[769]_  = \new_[298]_  | \new_[299]_ ;
  assign \new_[770]_  = \new_[300]_  | \new_[769]_ ;
  assign \new_[773]_  = \new_[296]_  | \new_[297]_ ;
  assign \new_[776]_  = \new_[294]_  | \new_[295]_ ;
  assign \new_[777]_  = \new_[776]_  | \new_[773]_ ;
  assign \new_[778]_  = \new_[777]_  | \new_[770]_ ;
  assign \new_[781]_  = \new_[292]_  | \new_[293]_ ;
  assign \new_[784]_  = \new_[290]_  | \new_[291]_ ;
  assign \new_[785]_  = \new_[784]_  | \new_[781]_ ;
  assign \new_[788]_  = \new_[288]_  | \new_[289]_ ;
  assign \new_[791]_  = \new_[286]_  | \new_[287]_ ;
  assign \new_[792]_  = \new_[791]_  | \new_[788]_ ;
  assign \new_[793]_  = \new_[792]_  | \new_[785]_ ;
  assign \new_[794]_  = \new_[793]_  | \new_[778]_ ;
  assign \new_[795]_  = \new_[794]_  | \new_[765]_ ;
  assign \new_[796]_  = \new_[795]_  | \new_[738]_ ;
  assign \new_[800]_  = \new_[283]_  | \new_[284]_ ;
  assign \new_[801]_  = \new_[285]_  | \new_[800]_ ;
  assign \new_[804]_  = \new_[281]_  | \new_[282]_ ;
  assign \new_[807]_  = \new_[279]_  | \new_[280]_ ;
  assign \new_[808]_  = \new_[807]_  | \new_[804]_ ;
  assign \new_[809]_  = \new_[808]_  | \new_[801]_ ;
  assign \new_[813]_  = \new_[276]_  | \new_[277]_ ;
  assign \new_[814]_  = \new_[278]_  | \new_[813]_ ;
  assign \new_[817]_  = \new_[274]_  | \new_[275]_ ;
  assign \new_[820]_  = \new_[272]_  | \new_[273]_ ;
  assign \new_[821]_  = \new_[820]_  | \new_[817]_ ;
  assign \new_[822]_  = \new_[821]_  | \new_[814]_ ;
  assign \new_[823]_  = \new_[822]_  | \new_[809]_ ;
  assign \new_[827]_  = \new_[269]_  | \new_[270]_ ;
  assign \new_[828]_  = \new_[271]_  | \new_[827]_ ;
  assign \new_[831]_  = \new_[267]_  | \new_[268]_ ;
  assign \new_[834]_  = \new_[265]_  | \new_[266]_ ;
  assign \new_[835]_  = \new_[834]_  | \new_[831]_ ;
  assign \new_[836]_  = \new_[835]_  | \new_[828]_ ;
  assign \new_[840]_  = \new_[262]_  | \new_[263]_ ;
  assign \new_[841]_  = \new_[264]_  | \new_[840]_ ;
  assign \new_[844]_  = \new_[260]_  | \new_[261]_ ;
  assign \new_[847]_  = \new_[258]_  | \new_[259]_ ;
  assign \new_[848]_  = \new_[847]_  | \new_[844]_ ;
  assign \new_[849]_  = \new_[848]_  | \new_[841]_ ;
  assign \new_[850]_  = \new_[849]_  | \new_[836]_ ;
  assign \new_[851]_  = \new_[850]_  | \new_[823]_ ;
  assign \new_[855]_  = \new_[255]_  | \new_[256]_ ;
  assign \new_[856]_  = \new_[257]_  | \new_[855]_ ;
  assign \new_[859]_  = \new_[253]_  | \new_[254]_ ;
  assign \new_[862]_  = \new_[251]_  | \new_[252]_ ;
  assign \new_[863]_  = \new_[862]_  | \new_[859]_ ;
  assign \new_[864]_  = \new_[863]_  | \new_[856]_ ;
  assign \new_[868]_  = \new_[248]_  | \new_[249]_ ;
  assign \new_[869]_  = \new_[250]_  | \new_[868]_ ;
  assign \new_[872]_  = \new_[246]_  | \new_[247]_ ;
  assign \new_[875]_  = \new_[244]_  | \new_[245]_ ;
  assign \new_[876]_  = \new_[875]_  | \new_[872]_ ;
  assign \new_[877]_  = \new_[876]_  | \new_[869]_ ;
  assign \new_[878]_  = \new_[877]_  | \new_[864]_ ;
  assign \new_[882]_  = \new_[241]_  | \new_[242]_ ;
  assign \new_[883]_  = \new_[243]_  | \new_[882]_ ;
  assign \new_[886]_  = \new_[239]_  | \new_[240]_ ;
  assign \new_[889]_  = \new_[237]_  | \new_[238]_ ;
  assign \new_[890]_  = \new_[889]_  | \new_[886]_ ;
  assign \new_[891]_  = \new_[890]_  | \new_[883]_ ;
  assign \new_[894]_  = \new_[235]_  | \new_[236]_ ;
  assign \new_[897]_  = \new_[233]_  | \new_[234]_ ;
  assign \new_[898]_  = \new_[897]_  | \new_[894]_ ;
  assign \new_[901]_  = \new_[231]_  | \new_[232]_ ;
  assign \new_[904]_  = \new_[229]_  | \new_[230]_ ;
  assign \new_[905]_  = \new_[904]_  | \new_[901]_ ;
  assign \new_[906]_  = \new_[905]_  | \new_[898]_ ;
  assign \new_[907]_  = \new_[906]_  | \new_[891]_ ;
  assign \new_[908]_  = \new_[907]_  | \new_[878]_ ;
  assign \new_[909]_  = \new_[908]_  | \new_[851]_ ;
  assign \new_[910]_  = \new_[909]_  | \new_[796]_ ;
  assign \new_[911]_  = \new_[910]_  | \new_[683]_ ;
  assign \new_[915]_  = \new_[226]_  | \new_[227]_ ;
  assign \new_[916]_  = \new_[228]_  | \new_[915]_ ;
  assign \new_[919]_  = \new_[224]_  | \new_[225]_ ;
  assign \new_[922]_  = \new_[222]_  | \new_[223]_ ;
  assign \new_[923]_  = \new_[922]_  | \new_[919]_ ;
  assign \new_[924]_  = \new_[923]_  | \new_[916]_ ;
  assign \new_[928]_  = \new_[219]_  | \new_[220]_ ;
  assign \new_[929]_  = \new_[221]_  | \new_[928]_ ;
  assign \new_[932]_  = \new_[217]_  | \new_[218]_ ;
  assign \new_[935]_  = \new_[215]_  | \new_[216]_ ;
  assign \new_[936]_  = \new_[935]_  | \new_[932]_ ;
  assign \new_[937]_  = \new_[936]_  | \new_[929]_ ;
  assign \new_[938]_  = \new_[937]_  | \new_[924]_ ;
  assign \new_[942]_  = \new_[212]_  | \new_[213]_ ;
  assign \new_[943]_  = \new_[214]_  | \new_[942]_ ;
  assign \new_[946]_  = \new_[210]_  | \new_[211]_ ;
  assign \new_[949]_  = \new_[208]_  | \new_[209]_ ;
  assign \new_[950]_  = \new_[949]_  | \new_[946]_ ;
  assign \new_[951]_  = \new_[950]_  | \new_[943]_ ;
  assign \new_[955]_  = \new_[205]_  | \new_[206]_ ;
  assign \new_[956]_  = \new_[207]_  | \new_[955]_ ;
  assign \new_[959]_  = \new_[203]_  | \new_[204]_ ;
  assign \new_[962]_  = \new_[201]_  | \new_[202]_ ;
  assign \new_[963]_  = \new_[962]_  | \new_[959]_ ;
  assign \new_[964]_  = \new_[963]_  | \new_[956]_ ;
  assign \new_[965]_  = \new_[964]_  | \new_[951]_ ;
  assign \new_[966]_  = \new_[965]_  | \new_[938]_ ;
  assign \new_[970]_  = \new_[198]_  | \new_[199]_ ;
  assign \new_[971]_  = \new_[200]_  | \new_[970]_ ;
  assign \new_[974]_  = \new_[196]_  | \new_[197]_ ;
  assign \new_[977]_  = \new_[194]_  | \new_[195]_ ;
  assign \new_[978]_  = \new_[977]_  | \new_[974]_ ;
  assign \new_[979]_  = \new_[978]_  | \new_[971]_ ;
  assign \new_[983]_  = \new_[191]_  | \new_[192]_ ;
  assign \new_[984]_  = \new_[193]_  | \new_[983]_ ;
  assign \new_[987]_  = \new_[189]_  | \new_[190]_ ;
  assign \new_[990]_  = \new_[187]_  | \new_[188]_ ;
  assign \new_[991]_  = \new_[990]_  | \new_[987]_ ;
  assign \new_[992]_  = \new_[991]_  | \new_[984]_ ;
  assign \new_[993]_  = \new_[992]_  | \new_[979]_ ;
  assign \new_[997]_  = \new_[184]_  | \new_[185]_ ;
  assign \new_[998]_  = \new_[186]_  | \new_[997]_ ;
  assign \new_[1001]_  = \new_[182]_  | \new_[183]_ ;
  assign \new_[1004]_  = \new_[180]_  | \new_[181]_ ;
  assign \new_[1005]_  = \new_[1004]_  | \new_[1001]_ ;
  assign \new_[1006]_  = \new_[1005]_  | \new_[998]_ ;
  assign \new_[1009]_  = \new_[178]_  | \new_[179]_ ;
  assign \new_[1012]_  = \new_[176]_  | \new_[177]_ ;
  assign \new_[1013]_  = \new_[1012]_  | \new_[1009]_ ;
  assign \new_[1016]_  = \new_[174]_  | \new_[175]_ ;
  assign \new_[1019]_  = \new_[172]_  | \new_[173]_ ;
  assign \new_[1020]_  = \new_[1019]_  | \new_[1016]_ ;
  assign \new_[1021]_  = \new_[1020]_  | \new_[1013]_ ;
  assign \new_[1022]_  = \new_[1021]_  | \new_[1006]_ ;
  assign \new_[1023]_  = \new_[1022]_  | \new_[993]_ ;
  assign \new_[1024]_  = \new_[1023]_  | \new_[966]_ ;
  assign \new_[1028]_  = \new_[169]_  | \new_[170]_ ;
  assign \new_[1029]_  = \new_[171]_  | \new_[1028]_ ;
  assign \new_[1032]_  = \new_[167]_  | \new_[168]_ ;
  assign \new_[1035]_  = \new_[165]_  | \new_[166]_ ;
  assign \new_[1036]_  = \new_[1035]_  | \new_[1032]_ ;
  assign \new_[1037]_  = \new_[1036]_  | \new_[1029]_ ;
  assign \new_[1041]_  = \new_[162]_  | \new_[163]_ ;
  assign \new_[1042]_  = \new_[164]_  | \new_[1041]_ ;
  assign \new_[1045]_  = \new_[160]_  | \new_[161]_ ;
  assign \new_[1048]_  = \new_[158]_  | \new_[159]_ ;
  assign \new_[1049]_  = \new_[1048]_  | \new_[1045]_ ;
  assign \new_[1050]_  = \new_[1049]_  | \new_[1042]_ ;
  assign \new_[1051]_  = \new_[1050]_  | \new_[1037]_ ;
  assign \new_[1055]_  = \new_[155]_  | \new_[156]_ ;
  assign \new_[1056]_  = \new_[157]_  | \new_[1055]_ ;
  assign \new_[1059]_  = \new_[153]_  | \new_[154]_ ;
  assign \new_[1062]_  = \new_[151]_  | \new_[152]_ ;
  assign \new_[1063]_  = \new_[1062]_  | \new_[1059]_ ;
  assign \new_[1064]_  = \new_[1063]_  | \new_[1056]_ ;
  assign \new_[1068]_  = \new_[148]_  | \new_[149]_ ;
  assign \new_[1069]_  = \new_[150]_  | \new_[1068]_ ;
  assign \new_[1072]_  = \new_[146]_  | \new_[147]_ ;
  assign \new_[1075]_  = \new_[144]_  | \new_[145]_ ;
  assign \new_[1076]_  = \new_[1075]_  | \new_[1072]_ ;
  assign \new_[1077]_  = \new_[1076]_  | \new_[1069]_ ;
  assign \new_[1078]_  = \new_[1077]_  | \new_[1064]_ ;
  assign \new_[1079]_  = \new_[1078]_  | \new_[1051]_ ;
  assign \new_[1083]_  = \new_[141]_  | \new_[142]_ ;
  assign \new_[1084]_  = \new_[143]_  | \new_[1083]_ ;
  assign \new_[1087]_  = \new_[139]_  | \new_[140]_ ;
  assign \new_[1090]_  = \new_[137]_  | \new_[138]_ ;
  assign \new_[1091]_  = \new_[1090]_  | \new_[1087]_ ;
  assign \new_[1092]_  = \new_[1091]_  | \new_[1084]_ ;
  assign \new_[1096]_  = \new_[134]_  | \new_[135]_ ;
  assign \new_[1097]_  = \new_[136]_  | \new_[1096]_ ;
  assign \new_[1100]_  = \new_[132]_  | \new_[133]_ ;
  assign \new_[1103]_  = \new_[130]_  | \new_[131]_ ;
  assign \new_[1104]_  = \new_[1103]_  | \new_[1100]_ ;
  assign \new_[1105]_  = \new_[1104]_  | \new_[1097]_ ;
  assign \new_[1106]_  = \new_[1105]_  | \new_[1092]_ ;
  assign \new_[1110]_  = \new_[127]_  | \new_[128]_ ;
  assign \new_[1111]_  = \new_[129]_  | \new_[1110]_ ;
  assign \new_[1114]_  = \new_[125]_  | \new_[126]_ ;
  assign \new_[1117]_  = \new_[123]_  | \new_[124]_ ;
  assign \new_[1118]_  = \new_[1117]_  | \new_[1114]_ ;
  assign \new_[1119]_  = \new_[1118]_  | \new_[1111]_ ;
  assign \new_[1122]_  = \new_[121]_  | \new_[122]_ ;
  assign \new_[1125]_  = \new_[119]_  | \new_[120]_ ;
  assign \new_[1126]_  = \new_[1125]_  | \new_[1122]_ ;
  assign \new_[1129]_  = \new_[117]_  | \new_[118]_ ;
  assign \new_[1132]_  = \new_[115]_  | \new_[116]_ ;
  assign \new_[1133]_  = \new_[1132]_  | \new_[1129]_ ;
  assign \new_[1134]_  = \new_[1133]_  | \new_[1126]_ ;
  assign \new_[1135]_  = \new_[1134]_  | \new_[1119]_ ;
  assign \new_[1136]_  = \new_[1135]_  | \new_[1106]_ ;
  assign \new_[1137]_  = \new_[1136]_  | \new_[1079]_ ;
  assign \new_[1138]_  = \new_[1137]_  | \new_[1024]_ ;
  assign \new_[1142]_  = \new_[112]_  | \new_[113]_ ;
  assign \new_[1143]_  = \new_[114]_  | \new_[1142]_ ;
  assign \new_[1146]_  = \new_[110]_  | \new_[111]_ ;
  assign \new_[1149]_  = \new_[108]_  | \new_[109]_ ;
  assign \new_[1150]_  = \new_[1149]_  | \new_[1146]_ ;
  assign \new_[1151]_  = \new_[1150]_  | \new_[1143]_ ;
  assign \new_[1155]_  = \new_[105]_  | \new_[106]_ ;
  assign \new_[1156]_  = \new_[107]_  | \new_[1155]_ ;
  assign \new_[1159]_  = \new_[103]_  | \new_[104]_ ;
  assign \new_[1162]_  = \new_[101]_  | \new_[102]_ ;
  assign \new_[1163]_  = \new_[1162]_  | \new_[1159]_ ;
  assign \new_[1164]_  = \new_[1163]_  | \new_[1156]_ ;
  assign \new_[1165]_  = \new_[1164]_  | \new_[1151]_ ;
  assign \new_[1169]_  = \new_[98]_  | \new_[99]_ ;
  assign \new_[1170]_  = \new_[100]_  | \new_[1169]_ ;
  assign \new_[1173]_  = \new_[96]_  | \new_[97]_ ;
  assign \new_[1176]_  = \new_[94]_  | \new_[95]_ ;
  assign \new_[1177]_  = \new_[1176]_  | \new_[1173]_ ;
  assign \new_[1178]_  = \new_[1177]_  | \new_[1170]_ ;
  assign \new_[1182]_  = \new_[91]_  | \new_[92]_ ;
  assign \new_[1183]_  = \new_[93]_  | \new_[1182]_ ;
  assign \new_[1186]_  = \new_[89]_  | \new_[90]_ ;
  assign \new_[1189]_  = \new_[87]_  | \new_[88]_ ;
  assign \new_[1190]_  = \new_[1189]_  | \new_[1186]_ ;
  assign \new_[1191]_  = \new_[1190]_  | \new_[1183]_ ;
  assign \new_[1192]_  = \new_[1191]_  | \new_[1178]_ ;
  assign \new_[1193]_  = \new_[1192]_  | \new_[1165]_ ;
  assign \new_[1197]_  = \new_[84]_  | \new_[85]_ ;
  assign \new_[1198]_  = \new_[86]_  | \new_[1197]_ ;
  assign \new_[1201]_  = \new_[82]_  | \new_[83]_ ;
  assign \new_[1204]_  = \new_[80]_  | \new_[81]_ ;
  assign \new_[1205]_  = \new_[1204]_  | \new_[1201]_ ;
  assign \new_[1206]_  = \new_[1205]_  | \new_[1198]_ ;
  assign \new_[1210]_  = \new_[77]_  | \new_[78]_ ;
  assign \new_[1211]_  = \new_[79]_  | \new_[1210]_ ;
  assign \new_[1214]_  = \new_[75]_  | \new_[76]_ ;
  assign \new_[1217]_  = \new_[73]_  | \new_[74]_ ;
  assign \new_[1218]_  = \new_[1217]_  | \new_[1214]_ ;
  assign \new_[1219]_  = \new_[1218]_  | \new_[1211]_ ;
  assign \new_[1220]_  = \new_[1219]_  | \new_[1206]_ ;
  assign \new_[1224]_  = \new_[70]_  | \new_[71]_ ;
  assign \new_[1225]_  = \new_[72]_  | \new_[1224]_ ;
  assign \new_[1228]_  = \new_[68]_  | \new_[69]_ ;
  assign \new_[1231]_  = \new_[66]_  | \new_[67]_ ;
  assign \new_[1232]_  = \new_[1231]_  | \new_[1228]_ ;
  assign \new_[1233]_  = \new_[1232]_  | \new_[1225]_ ;
  assign \new_[1236]_  = \new_[64]_  | \new_[65]_ ;
  assign \new_[1239]_  = \new_[62]_  | \new_[63]_ ;
  assign \new_[1240]_  = \new_[1239]_  | \new_[1236]_ ;
  assign \new_[1243]_  = \new_[60]_  | \new_[61]_ ;
  assign \new_[1246]_  = \new_[58]_  | \new_[59]_ ;
  assign \new_[1247]_  = \new_[1246]_  | \new_[1243]_ ;
  assign \new_[1248]_  = \new_[1247]_  | \new_[1240]_ ;
  assign \new_[1249]_  = \new_[1248]_  | \new_[1233]_ ;
  assign \new_[1250]_  = \new_[1249]_  | \new_[1220]_ ;
  assign \new_[1251]_  = \new_[1250]_  | \new_[1193]_ ;
  assign \new_[1255]_  = \new_[55]_  | \new_[56]_ ;
  assign \new_[1256]_  = \new_[57]_  | \new_[1255]_ ;
  assign \new_[1259]_  = \new_[53]_  | \new_[54]_ ;
  assign \new_[1262]_  = \new_[51]_  | \new_[52]_ ;
  assign \new_[1263]_  = \new_[1262]_  | \new_[1259]_ ;
  assign \new_[1264]_  = \new_[1263]_  | \new_[1256]_ ;
  assign \new_[1268]_  = \new_[48]_  | \new_[49]_ ;
  assign \new_[1269]_  = \new_[50]_  | \new_[1268]_ ;
  assign \new_[1272]_  = \new_[46]_  | \new_[47]_ ;
  assign \new_[1275]_  = \new_[44]_  | \new_[45]_ ;
  assign \new_[1276]_  = \new_[1275]_  | \new_[1272]_ ;
  assign \new_[1277]_  = \new_[1276]_  | \new_[1269]_ ;
  assign \new_[1278]_  = \new_[1277]_  | \new_[1264]_ ;
  assign \new_[1282]_  = \new_[41]_  | \new_[42]_ ;
  assign \new_[1283]_  = \new_[43]_  | \new_[1282]_ ;
  assign \new_[1286]_  = \new_[39]_  | \new_[40]_ ;
  assign \new_[1289]_  = \new_[37]_  | \new_[38]_ ;
  assign \new_[1290]_  = \new_[1289]_  | \new_[1286]_ ;
  assign \new_[1291]_  = \new_[1290]_  | \new_[1283]_ ;
  assign \new_[1295]_  = \new_[34]_  | \new_[35]_ ;
  assign \new_[1296]_  = \new_[36]_  | \new_[1295]_ ;
  assign \new_[1299]_  = \new_[32]_  | \new_[33]_ ;
  assign \new_[1302]_  = \new_[30]_  | \new_[31]_ ;
  assign \new_[1303]_  = \new_[1302]_  | \new_[1299]_ ;
  assign \new_[1304]_  = \new_[1303]_  | \new_[1296]_ ;
  assign \new_[1305]_  = \new_[1304]_  | \new_[1291]_ ;
  assign \new_[1306]_  = \new_[1305]_  | \new_[1278]_ ;
  assign \new_[1310]_  = \new_[27]_  | \new_[28]_ ;
  assign \new_[1311]_  = \new_[29]_  | \new_[1310]_ ;
  assign \new_[1314]_  = \new_[25]_  | \new_[26]_ ;
  assign \new_[1317]_  = \new_[23]_  | \new_[24]_ ;
  assign \new_[1318]_  = \new_[1317]_  | \new_[1314]_ ;
  assign \new_[1319]_  = \new_[1318]_  | \new_[1311]_ ;
  assign \new_[1323]_  = \new_[20]_  | \new_[21]_ ;
  assign \new_[1324]_  = \new_[22]_  | \new_[1323]_ ;
  assign \new_[1327]_  = \new_[18]_  | \new_[19]_ ;
  assign \new_[1330]_  = \new_[16]_  | \new_[17]_ ;
  assign \new_[1331]_  = \new_[1330]_  | \new_[1327]_ ;
  assign \new_[1332]_  = \new_[1331]_  | \new_[1324]_ ;
  assign \new_[1333]_  = \new_[1332]_  | \new_[1319]_ ;
  assign \new_[1337]_  = \new_[13]_  | \new_[14]_ ;
  assign \new_[1338]_  = \new_[15]_  | \new_[1337]_ ;
  assign \new_[1341]_  = \new_[11]_  | \new_[12]_ ;
  assign \new_[1344]_  = \new_[9]_  | \new_[10]_ ;
  assign \new_[1345]_  = \new_[1344]_  | \new_[1341]_ ;
  assign \new_[1346]_  = \new_[1345]_  | \new_[1338]_ ;
  assign \new_[1349]_  = \new_[7]_  | \new_[8]_ ;
  assign \new_[1352]_  = \new_[5]_  | \new_[6]_ ;
  assign \new_[1353]_  = \new_[1352]_  | \new_[1349]_ ;
  assign \new_[1356]_  = \new_[3]_  | \new_[4]_ ;
  assign \new_[1359]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[1360]_  = \new_[1359]_  | \new_[1356]_ ;
  assign \new_[1361]_  = \new_[1360]_  | \new_[1353]_ ;
  assign \new_[1362]_  = \new_[1361]_  | \new_[1346]_ ;
  assign \new_[1363]_  = \new_[1362]_  | \new_[1333]_ ;
  assign \new_[1364]_  = \new_[1363]_  | \new_[1306]_ ;
  assign \new_[1365]_  = \new_[1364]_  | \new_[1251]_ ;
  assign \new_[1366]_  = \new_[1365]_  | \new_[1138]_ ;
  assign \new_[1369]_  = ~A167 & A170;
  assign \new_[1373]_  = A200 & ~A199;
  assign \new_[1374]_  = ~A166 & \new_[1373]_ ;
  assign \new_[1377]_  = ~A167 & ~A169;
  assign \new_[1381]_  = A200 & ~A199;
  assign \new_[1382]_  = ~A166 & \new_[1381]_ ;
  assign \new_[1386]_  = A167 & ~A168;
  assign \new_[1387]_  = A170 & \new_[1386]_ ;
  assign \new_[1391]_  = A200 & ~A199;
  assign \new_[1392]_  = A166 & \new_[1391]_ ;
  assign \new_[1396]_  = A167 & ~A168;
  assign \new_[1397]_  = ~A170 & \new_[1396]_ ;
  assign \new_[1401]_  = A200 & ~A199;
  assign \new_[1402]_  = ~A166 & \new_[1401]_ ;
  assign \new_[1406]_  = ~A167 & ~A168;
  assign \new_[1407]_  = ~A170 & \new_[1406]_ ;
  assign \new_[1411]_  = A200 & ~A199;
  assign \new_[1412]_  = A166 & \new_[1411]_ ;
  assign \new_[1416]_  = A167 & ~A168;
  assign \new_[1417]_  = A169 & \new_[1416]_ ;
  assign \new_[1421]_  = A200 & ~A199;
  assign \new_[1422]_  = ~A166 & \new_[1421]_ ;
  assign \new_[1426]_  = ~A167 & ~A168;
  assign \new_[1427]_  = A169 & \new_[1426]_ ;
  assign \new_[1431]_  = A200 & ~A199;
  assign \new_[1432]_  = A166 & \new_[1431]_ ;
  assign \new_[1436]_  = A167 & ~A168;
  assign \new_[1437]_  = ~A169 & \new_[1436]_ ;
  assign \new_[1441]_  = A200 & ~A199;
  assign \new_[1442]_  = A166 & \new_[1441]_ ;
  assign \new_[1446]_  = ~A166 & ~A167;
  assign \new_[1447]_  = A170 & \new_[1446]_ ;
  assign \new_[1450]_  = ~A200 & A199;
  assign \new_[1453]_  = A202 & A201;
  assign \new_[1454]_  = \new_[1453]_  & \new_[1450]_ ;
  assign \new_[1458]_  = ~A166 & ~A167;
  assign \new_[1459]_  = A170 & \new_[1458]_ ;
  assign \new_[1462]_  = ~A200 & A199;
  assign \new_[1465]_  = A203 & A201;
  assign \new_[1466]_  = \new_[1465]_  & \new_[1462]_ ;
  assign \new_[1470]_  = ~A166 & ~A167;
  assign \new_[1471]_  = ~A169 & \new_[1470]_ ;
  assign \new_[1474]_  = ~A200 & A199;
  assign \new_[1477]_  = A202 & A201;
  assign \new_[1478]_  = \new_[1477]_  & \new_[1474]_ ;
  assign \new_[1482]_  = ~A166 & ~A167;
  assign \new_[1483]_  = ~A169 & \new_[1482]_ ;
  assign \new_[1486]_  = ~A200 & A199;
  assign \new_[1489]_  = A203 & A201;
  assign \new_[1490]_  = \new_[1489]_  & \new_[1486]_ ;
  assign \new_[1493]_  = A166 & A168;
  assign \new_[1496]_  = ~A201 & A199;
  assign \new_[1497]_  = \new_[1496]_  & \new_[1493]_ ;
  assign \new_[1500]_  = A233 & ~A232;
  assign \new_[1503]_  = A299 & ~A298;
  assign \new_[1504]_  = \new_[1503]_  & \new_[1500]_ ;
  assign \new_[1507]_  = A166 & A168;
  assign \new_[1510]_  = ~A201 & A199;
  assign \new_[1511]_  = \new_[1510]_  & \new_[1507]_ ;
  assign \new_[1514]_  = A233 & ~A232;
  assign \new_[1517]_  = A266 & ~A265;
  assign \new_[1518]_  = \new_[1517]_  & \new_[1514]_ ;
  assign \new_[1521]_  = A166 & A168;
  assign \new_[1524]_  = A200 & A199;
  assign \new_[1525]_  = \new_[1524]_  & \new_[1521]_ ;
  assign \new_[1528]_  = A233 & ~A232;
  assign \new_[1531]_  = A299 & ~A298;
  assign \new_[1532]_  = \new_[1531]_  & \new_[1528]_ ;
  assign \new_[1535]_  = A166 & A168;
  assign \new_[1538]_  = A200 & A199;
  assign \new_[1539]_  = \new_[1538]_  & \new_[1535]_ ;
  assign \new_[1542]_  = A233 & ~A232;
  assign \new_[1545]_  = A266 & ~A265;
  assign \new_[1546]_  = \new_[1545]_  & \new_[1542]_ ;
  assign \new_[1549]_  = A166 & A168;
  assign \new_[1552]_  = ~A200 & ~A199;
  assign \new_[1553]_  = \new_[1552]_  & \new_[1549]_ ;
  assign \new_[1556]_  = A233 & ~A232;
  assign \new_[1559]_  = A299 & ~A298;
  assign \new_[1560]_  = \new_[1559]_  & \new_[1556]_ ;
  assign \new_[1563]_  = A166 & A168;
  assign \new_[1566]_  = ~A200 & ~A199;
  assign \new_[1567]_  = \new_[1566]_  & \new_[1563]_ ;
  assign \new_[1570]_  = A233 & ~A232;
  assign \new_[1573]_  = A266 & ~A265;
  assign \new_[1574]_  = \new_[1573]_  & \new_[1570]_ ;
  assign \new_[1577]_  = A167 & A168;
  assign \new_[1580]_  = ~A201 & A199;
  assign \new_[1581]_  = \new_[1580]_  & \new_[1577]_ ;
  assign \new_[1584]_  = A233 & ~A232;
  assign \new_[1587]_  = A299 & ~A298;
  assign \new_[1588]_  = \new_[1587]_  & \new_[1584]_ ;
  assign \new_[1591]_  = A167 & A168;
  assign \new_[1594]_  = ~A201 & A199;
  assign \new_[1595]_  = \new_[1594]_  & \new_[1591]_ ;
  assign \new_[1598]_  = A233 & ~A232;
  assign \new_[1601]_  = A266 & ~A265;
  assign \new_[1602]_  = \new_[1601]_  & \new_[1598]_ ;
  assign \new_[1605]_  = A167 & A168;
  assign \new_[1608]_  = A200 & A199;
  assign \new_[1609]_  = \new_[1608]_  & \new_[1605]_ ;
  assign \new_[1612]_  = A233 & ~A232;
  assign \new_[1615]_  = A299 & ~A298;
  assign \new_[1616]_  = \new_[1615]_  & \new_[1612]_ ;
  assign \new_[1619]_  = A167 & A168;
  assign \new_[1622]_  = A200 & A199;
  assign \new_[1623]_  = \new_[1622]_  & \new_[1619]_ ;
  assign \new_[1626]_  = A233 & ~A232;
  assign \new_[1629]_  = A266 & ~A265;
  assign \new_[1630]_  = \new_[1629]_  & \new_[1626]_ ;
  assign \new_[1633]_  = A167 & A168;
  assign \new_[1636]_  = ~A200 & ~A199;
  assign \new_[1637]_  = \new_[1636]_  & \new_[1633]_ ;
  assign \new_[1640]_  = A233 & ~A232;
  assign \new_[1643]_  = A299 & ~A298;
  assign \new_[1644]_  = \new_[1643]_  & \new_[1640]_ ;
  assign \new_[1647]_  = A167 & A168;
  assign \new_[1650]_  = ~A200 & ~A199;
  assign \new_[1651]_  = \new_[1650]_  & \new_[1647]_ ;
  assign \new_[1654]_  = A233 & ~A232;
  assign \new_[1657]_  = A266 & ~A265;
  assign \new_[1658]_  = \new_[1657]_  & \new_[1654]_ ;
  assign \new_[1661]_  = ~A168 & A170;
  assign \new_[1664]_  = A166 & A167;
  assign \new_[1665]_  = \new_[1664]_  & \new_[1661]_ ;
  assign \new_[1668]_  = ~A200 & A199;
  assign \new_[1671]_  = A202 & A201;
  assign \new_[1672]_  = \new_[1671]_  & \new_[1668]_ ;
  assign \new_[1675]_  = ~A168 & A170;
  assign \new_[1678]_  = A166 & A167;
  assign \new_[1679]_  = \new_[1678]_  & \new_[1675]_ ;
  assign \new_[1682]_  = ~A200 & A199;
  assign \new_[1685]_  = A203 & A201;
  assign \new_[1686]_  = \new_[1685]_  & \new_[1682]_ ;
  assign \new_[1689]_  = ~A168 & ~A170;
  assign \new_[1692]_  = ~A166 & A167;
  assign \new_[1693]_  = \new_[1692]_  & \new_[1689]_ ;
  assign \new_[1696]_  = ~A200 & A199;
  assign \new_[1699]_  = A202 & A201;
  assign \new_[1700]_  = \new_[1699]_  & \new_[1696]_ ;
  assign \new_[1703]_  = ~A168 & ~A170;
  assign \new_[1706]_  = ~A166 & A167;
  assign \new_[1707]_  = \new_[1706]_  & \new_[1703]_ ;
  assign \new_[1710]_  = ~A200 & A199;
  assign \new_[1713]_  = A203 & A201;
  assign \new_[1714]_  = \new_[1713]_  & \new_[1710]_ ;
  assign \new_[1717]_  = ~A168 & ~A170;
  assign \new_[1720]_  = A166 & ~A167;
  assign \new_[1721]_  = \new_[1720]_  & \new_[1717]_ ;
  assign \new_[1724]_  = ~A200 & A199;
  assign \new_[1727]_  = A202 & A201;
  assign \new_[1728]_  = \new_[1727]_  & \new_[1724]_ ;
  assign \new_[1731]_  = ~A168 & ~A170;
  assign \new_[1734]_  = A166 & ~A167;
  assign \new_[1735]_  = \new_[1734]_  & \new_[1731]_ ;
  assign \new_[1738]_  = ~A200 & A199;
  assign \new_[1741]_  = A203 & A201;
  assign \new_[1742]_  = \new_[1741]_  & \new_[1738]_ ;
  assign \new_[1745]_  = ~A168 & A169;
  assign \new_[1748]_  = ~A166 & A167;
  assign \new_[1749]_  = \new_[1748]_  & \new_[1745]_ ;
  assign \new_[1752]_  = ~A200 & A199;
  assign \new_[1755]_  = A202 & A201;
  assign \new_[1756]_  = \new_[1755]_  & \new_[1752]_ ;
  assign \new_[1759]_  = ~A168 & A169;
  assign \new_[1762]_  = ~A166 & A167;
  assign \new_[1763]_  = \new_[1762]_  & \new_[1759]_ ;
  assign \new_[1766]_  = ~A200 & A199;
  assign \new_[1769]_  = A203 & A201;
  assign \new_[1770]_  = \new_[1769]_  & \new_[1766]_ ;
  assign \new_[1773]_  = ~A168 & A169;
  assign \new_[1776]_  = A166 & ~A167;
  assign \new_[1777]_  = \new_[1776]_  & \new_[1773]_ ;
  assign \new_[1780]_  = ~A200 & A199;
  assign \new_[1783]_  = A202 & A201;
  assign \new_[1784]_  = \new_[1783]_  & \new_[1780]_ ;
  assign \new_[1787]_  = ~A168 & A169;
  assign \new_[1790]_  = A166 & ~A167;
  assign \new_[1791]_  = \new_[1790]_  & \new_[1787]_ ;
  assign \new_[1794]_  = ~A200 & A199;
  assign \new_[1797]_  = A203 & A201;
  assign \new_[1798]_  = \new_[1797]_  & \new_[1794]_ ;
  assign \new_[1801]_  = ~A168 & ~A169;
  assign \new_[1804]_  = A166 & A167;
  assign \new_[1805]_  = \new_[1804]_  & \new_[1801]_ ;
  assign \new_[1808]_  = ~A200 & A199;
  assign \new_[1811]_  = A202 & A201;
  assign \new_[1812]_  = \new_[1811]_  & \new_[1808]_ ;
  assign \new_[1815]_  = ~A168 & ~A169;
  assign \new_[1818]_  = A166 & A167;
  assign \new_[1819]_  = \new_[1818]_  & \new_[1815]_ ;
  assign \new_[1822]_  = ~A200 & A199;
  assign \new_[1825]_  = A203 & A201;
  assign \new_[1826]_  = \new_[1825]_  & \new_[1822]_ ;
  assign \new_[1829]_  = A166 & A168;
  assign \new_[1832]_  = ~A202 & A199;
  assign \new_[1833]_  = \new_[1832]_  & \new_[1829]_ ;
  assign \new_[1836]_  = ~A232 & ~A203;
  assign \new_[1840]_  = A299 & ~A298;
  assign \new_[1841]_  = A233 & \new_[1840]_ ;
  assign \new_[1842]_  = \new_[1841]_  & \new_[1836]_ ;
  assign \new_[1845]_  = A166 & A168;
  assign \new_[1848]_  = ~A202 & A199;
  assign \new_[1849]_  = \new_[1848]_  & \new_[1845]_ ;
  assign \new_[1852]_  = ~A232 & ~A203;
  assign \new_[1856]_  = A266 & ~A265;
  assign \new_[1857]_  = A233 & \new_[1856]_ ;
  assign \new_[1858]_  = \new_[1857]_  & \new_[1852]_ ;
  assign \new_[1861]_  = A167 & A168;
  assign \new_[1864]_  = ~A202 & A199;
  assign \new_[1865]_  = \new_[1864]_  & \new_[1861]_ ;
  assign \new_[1868]_  = ~A232 & ~A203;
  assign \new_[1872]_  = A299 & ~A298;
  assign \new_[1873]_  = A233 & \new_[1872]_ ;
  assign \new_[1874]_  = \new_[1873]_  & \new_[1868]_ ;
  assign \new_[1877]_  = A167 & A168;
  assign \new_[1880]_  = ~A202 & A199;
  assign \new_[1881]_  = \new_[1880]_  & \new_[1877]_ ;
  assign \new_[1884]_  = ~A232 & ~A203;
  assign \new_[1888]_  = A266 & ~A265;
  assign \new_[1889]_  = A233 & \new_[1888]_ ;
  assign \new_[1890]_  = \new_[1889]_  & \new_[1884]_ ;
  assign \new_[1893]_  = A166 & A168;
  assign \new_[1897]_  = ~A232 & ~A201;
  assign \new_[1898]_  = A199 & \new_[1897]_ ;
  assign \new_[1899]_  = \new_[1898]_  & \new_[1893]_ ;
  assign \new_[1902]_  = A298 & A233;
  assign \new_[1906]_  = A301 & A300;
  assign \new_[1907]_  = ~A299 & \new_[1906]_ ;
  assign \new_[1908]_  = \new_[1907]_  & \new_[1902]_ ;
  assign \new_[1911]_  = A166 & A168;
  assign \new_[1915]_  = ~A232 & ~A201;
  assign \new_[1916]_  = A199 & \new_[1915]_ ;
  assign \new_[1917]_  = \new_[1916]_  & \new_[1911]_ ;
  assign \new_[1920]_  = A298 & A233;
  assign \new_[1924]_  = A302 & A300;
  assign \new_[1925]_  = ~A299 & \new_[1924]_ ;
  assign \new_[1926]_  = \new_[1925]_  & \new_[1920]_ ;
  assign \new_[1929]_  = A166 & A168;
  assign \new_[1933]_  = ~A232 & ~A201;
  assign \new_[1934]_  = A199 & \new_[1933]_ ;
  assign \new_[1935]_  = \new_[1934]_  & \new_[1929]_ ;
  assign \new_[1938]_  = A265 & A233;
  assign \new_[1942]_  = A268 & A267;
  assign \new_[1943]_  = ~A266 & \new_[1942]_ ;
  assign \new_[1944]_  = \new_[1943]_  & \new_[1938]_ ;
  assign \new_[1947]_  = A166 & A168;
  assign \new_[1951]_  = ~A232 & ~A201;
  assign \new_[1952]_  = A199 & \new_[1951]_ ;
  assign \new_[1953]_  = \new_[1952]_  & \new_[1947]_ ;
  assign \new_[1956]_  = A265 & A233;
  assign \new_[1960]_  = A269 & A267;
  assign \new_[1961]_  = ~A266 & \new_[1960]_ ;
  assign \new_[1962]_  = \new_[1961]_  & \new_[1956]_ ;
  assign \new_[1965]_  = A166 & A168;
  assign \new_[1969]_  = A232 & ~A201;
  assign \new_[1970]_  = A199 & \new_[1969]_ ;
  assign \new_[1971]_  = \new_[1970]_  & \new_[1965]_ ;
  assign \new_[1974]_  = A234 & ~A233;
  assign \new_[1978]_  = A299 & ~A298;
  assign \new_[1979]_  = A235 & \new_[1978]_ ;
  assign \new_[1980]_  = \new_[1979]_  & \new_[1974]_ ;
  assign \new_[1983]_  = A166 & A168;
  assign \new_[1987]_  = A232 & ~A201;
  assign \new_[1988]_  = A199 & \new_[1987]_ ;
  assign \new_[1989]_  = \new_[1988]_  & \new_[1983]_ ;
  assign \new_[1992]_  = A234 & ~A233;
  assign \new_[1996]_  = A266 & ~A265;
  assign \new_[1997]_  = A235 & \new_[1996]_ ;
  assign \new_[1998]_  = \new_[1997]_  & \new_[1992]_ ;
  assign \new_[2001]_  = A166 & A168;
  assign \new_[2005]_  = A232 & ~A201;
  assign \new_[2006]_  = A199 & \new_[2005]_ ;
  assign \new_[2007]_  = \new_[2006]_  & \new_[2001]_ ;
  assign \new_[2010]_  = A234 & ~A233;
  assign \new_[2014]_  = A299 & ~A298;
  assign \new_[2015]_  = A236 & \new_[2014]_ ;
  assign \new_[2016]_  = \new_[2015]_  & \new_[2010]_ ;
  assign \new_[2019]_  = A166 & A168;
  assign \new_[2023]_  = A232 & ~A201;
  assign \new_[2024]_  = A199 & \new_[2023]_ ;
  assign \new_[2025]_  = \new_[2024]_  & \new_[2019]_ ;
  assign \new_[2028]_  = A234 & ~A233;
  assign \new_[2032]_  = A266 & ~A265;
  assign \new_[2033]_  = A236 & \new_[2032]_ ;
  assign \new_[2034]_  = \new_[2033]_  & \new_[2028]_ ;
  assign \new_[2037]_  = A166 & A168;
  assign \new_[2041]_  = ~A232 & A200;
  assign \new_[2042]_  = A199 & \new_[2041]_ ;
  assign \new_[2043]_  = \new_[2042]_  & \new_[2037]_ ;
  assign \new_[2046]_  = A298 & A233;
  assign \new_[2050]_  = A301 & A300;
  assign \new_[2051]_  = ~A299 & \new_[2050]_ ;
  assign \new_[2052]_  = \new_[2051]_  & \new_[2046]_ ;
  assign \new_[2055]_  = A166 & A168;
  assign \new_[2059]_  = ~A232 & A200;
  assign \new_[2060]_  = A199 & \new_[2059]_ ;
  assign \new_[2061]_  = \new_[2060]_  & \new_[2055]_ ;
  assign \new_[2064]_  = A298 & A233;
  assign \new_[2068]_  = A302 & A300;
  assign \new_[2069]_  = ~A299 & \new_[2068]_ ;
  assign \new_[2070]_  = \new_[2069]_  & \new_[2064]_ ;
  assign \new_[2073]_  = A166 & A168;
  assign \new_[2077]_  = ~A232 & A200;
  assign \new_[2078]_  = A199 & \new_[2077]_ ;
  assign \new_[2079]_  = \new_[2078]_  & \new_[2073]_ ;
  assign \new_[2082]_  = A265 & A233;
  assign \new_[2086]_  = A268 & A267;
  assign \new_[2087]_  = ~A266 & \new_[2086]_ ;
  assign \new_[2088]_  = \new_[2087]_  & \new_[2082]_ ;
  assign \new_[2091]_  = A166 & A168;
  assign \new_[2095]_  = ~A232 & A200;
  assign \new_[2096]_  = A199 & \new_[2095]_ ;
  assign \new_[2097]_  = \new_[2096]_  & \new_[2091]_ ;
  assign \new_[2100]_  = A265 & A233;
  assign \new_[2104]_  = A269 & A267;
  assign \new_[2105]_  = ~A266 & \new_[2104]_ ;
  assign \new_[2106]_  = \new_[2105]_  & \new_[2100]_ ;
  assign \new_[2109]_  = A166 & A168;
  assign \new_[2113]_  = A232 & A200;
  assign \new_[2114]_  = A199 & \new_[2113]_ ;
  assign \new_[2115]_  = \new_[2114]_  & \new_[2109]_ ;
  assign \new_[2118]_  = A234 & ~A233;
  assign \new_[2122]_  = A299 & ~A298;
  assign \new_[2123]_  = A235 & \new_[2122]_ ;
  assign \new_[2124]_  = \new_[2123]_  & \new_[2118]_ ;
  assign \new_[2127]_  = A166 & A168;
  assign \new_[2131]_  = A232 & A200;
  assign \new_[2132]_  = A199 & \new_[2131]_ ;
  assign \new_[2133]_  = \new_[2132]_  & \new_[2127]_ ;
  assign \new_[2136]_  = A234 & ~A233;
  assign \new_[2140]_  = A266 & ~A265;
  assign \new_[2141]_  = A235 & \new_[2140]_ ;
  assign \new_[2142]_  = \new_[2141]_  & \new_[2136]_ ;
  assign \new_[2145]_  = A166 & A168;
  assign \new_[2149]_  = A232 & A200;
  assign \new_[2150]_  = A199 & \new_[2149]_ ;
  assign \new_[2151]_  = \new_[2150]_  & \new_[2145]_ ;
  assign \new_[2154]_  = A234 & ~A233;
  assign \new_[2158]_  = A299 & ~A298;
  assign \new_[2159]_  = A236 & \new_[2158]_ ;
  assign \new_[2160]_  = \new_[2159]_  & \new_[2154]_ ;
  assign \new_[2163]_  = A166 & A168;
  assign \new_[2167]_  = A232 & A200;
  assign \new_[2168]_  = A199 & \new_[2167]_ ;
  assign \new_[2169]_  = \new_[2168]_  & \new_[2163]_ ;
  assign \new_[2172]_  = A234 & ~A233;
  assign \new_[2176]_  = A266 & ~A265;
  assign \new_[2177]_  = A236 & \new_[2176]_ ;
  assign \new_[2178]_  = \new_[2177]_  & \new_[2172]_ ;
  assign \new_[2181]_  = A166 & A168;
  assign \new_[2185]_  = ~A232 & ~A200;
  assign \new_[2186]_  = ~A199 & \new_[2185]_ ;
  assign \new_[2187]_  = \new_[2186]_  & \new_[2181]_ ;
  assign \new_[2190]_  = A298 & A233;
  assign \new_[2194]_  = A301 & A300;
  assign \new_[2195]_  = ~A299 & \new_[2194]_ ;
  assign \new_[2196]_  = \new_[2195]_  & \new_[2190]_ ;
  assign \new_[2199]_  = A166 & A168;
  assign \new_[2203]_  = ~A232 & ~A200;
  assign \new_[2204]_  = ~A199 & \new_[2203]_ ;
  assign \new_[2205]_  = \new_[2204]_  & \new_[2199]_ ;
  assign \new_[2208]_  = A298 & A233;
  assign \new_[2212]_  = A302 & A300;
  assign \new_[2213]_  = ~A299 & \new_[2212]_ ;
  assign \new_[2214]_  = \new_[2213]_  & \new_[2208]_ ;
  assign \new_[2217]_  = A166 & A168;
  assign \new_[2221]_  = ~A232 & ~A200;
  assign \new_[2222]_  = ~A199 & \new_[2221]_ ;
  assign \new_[2223]_  = \new_[2222]_  & \new_[2217]_ ;
  assign \new_[2226]_  = A265 & A233;
  assign \new_[2230]_  = A268 & A267;
  assign \new_[2231]_  = ~A266 & \new_[2230]_ ;
  assign \new_[2232]_  = \new_[2231]_  & \new_[2226]_ ;
  assign \new_[2235]_  = A166 & A168;
  assign \new_[2239]_  = ~A232 & ~A200;
  assign \new_[2240]_  = ~A199 & \new_[2239]_ ;
  assign \new_[2241]_  = \new_[2240]_  & \new_[2235]_ ;
  assign \new_[2244]_  = A265 & A233;
  assign \new_[2248]_  = A269 & A267;
  assign \new_[2249]_  = ~A266 & \new_[2248]_ ;
  assign \new_[2250]_  = \new_[2249]_  & \new_[2244]_ ;
  assign \new_[2253]_  = A166 & A168;
  assign \new_[2257]_  = A232 & ~A200;
  assign \new_[2258]_  = ~A199 & \new_[2257]_ ;
  assign \new_[2259]_  = \new_[2258]_  & \new_[2253]_ ;
  assign \new_[2262]_  = A234 & ~A233;
  assign \new_[2266]_  = A299 & ~A298;
  assign \new_[2267]_  = A235 & \new_[2266]_ ;
  assign \new_[2268]_  = \new_[2267]_  & \new_[2262]_ ;
  assign \new_[2271]_  = A166 & A168;
  assign \new_[2275]_  = A232 & ~A200;
  assign \new_[2276]_  = ~A199 & \new_[2275]_ ;
  assign \new_[2277]_  = \new_[2276]_  & \new_[2271]_ ;
  assign \new_[2280]_  = A234 & ~A233;
  assign \new_[2284]_  = A266 & ~A265;
  assign \new_[2285]_  = A235 & \new_[2284]_ ;
  assign \new_[2286]_  = \new_[2285]_  & \new_[2280]_ ;
  assign \new_[2289]_  = A166 & A168;
  assign \new_[2293]_  = A232 & ~A200;
  assign \new_[2294]_  = ~A199 & \new_[2293]_ ;
  assign \new_[2295]_  = \new_[2294]_  & \new_[2289]_ ;
  assign \new_[2298]_  = A234 & ~A233;
  assign \new_[2302]_  = A299 & ~A298;
  assign \new_[2303]_  = A236 & \new_[2302]_ ;
  assign \new_[2304]_  = \new_[2303]_  & \new_[2298]_ ;
  assign \new_[2307]_  = A166 & A168;
  assign \new_[2311]_  = A232 & ~A200;
  assign \new_[2312]_  = ~A199 & \new_[2311]_ ;
  assign \new_[2313]_  = \new_[2312]_  & \new_[2307]_ ;
  assign \new_[2316]_  = A234 & ~A233;
  assign \new_[2320]_  = A266 & ~A265;
  assign \new_[2321]_  = A236 & \new_[2320]_ ;
  assign \new_[2322]_  = \new_[2321]_  & \new_[2316]_ ;
  assign \new_[2325]_  = A167 & A168;
  assign \new_[2329]_  = ~A232 & ~A201;
  assign \new_[2330]_  = A199 & \new_[2329]_ ;
  assign \new_[2331]_  = \new_[2330]_  & \new_[2325]_ ;
  assign \new_[2334]_  = A298 & A233;
  assign \new_[2338]_  = A301 & A300;
  assign \new_[2339]_  = ~A299 & \new_[2338]_ ;
  assign \new_[2340]_  = \new_[2339]_  & \new_[2334]_ ;
  assign \new_[2343]_  = A167 & A168;
  assign \new_[2347]_  = ~A232 & ~A201;
  assign \new_[2348]_  = A199 & \new_[2347]_ ;
  assign \new_[2349]_  = \new_[2348]_  & \new_[2343]_ ;
  assign \new_[2352]_  = A298 & A233;
  assign \new_[2356]_  = A302 & A300;
  assign \new_[2357]_  = ~A299 & \new_[2356]_ ;
  assign \new_[2358]_  = \new_[2357]_  & \new_[2352]_ ;
  assign \new_[2361]_  = A167 & A168;
  assign \new_[2365]_  = ~A232 & ~A201;
  assign \new_[2366]_  = A199 & \new_[2365]_ ;
  assign \new_[2367]_  = \new_[2366]_  & \new_[2361]_ ;
  assign \new_[2370]_  = A265 & A233;
  assign \new_[2374]_  = A268 & A267;
  assign \new_[2375]_  = ~A266 & \new_[2374]_ ;
  assign \new_[2376]_  = \new_[2375]_  & \new_[2370]_ ;
  assign \new_[2379]_  = A167 & A168;
  assign \new_[2383]_  = ~A232 & ~A201;
  assign \new_[2384]_  = A199 & \new_[2383]_ ;
  assign \new_[2385]_  = \new_[2384]_  & \new_[2379]_ ;
  assign \new_[2388]_  = A265 & A233;
  assign \new_[2392]_  = A269 & A267;
  assign \new_[2393]_  = ~A266 & \new_[2392]_ ;
  assign \new_[2394]_  = \new_[2393]_  & \new_[2388]_ ;
  assign \new_[2397]_  = A167 & A168;
  assign \new_[2401]_  = A232 & ~A201;
  assign \new_[2402]_  = A199 & \new_[2401]_ ;
  assign \new_[2403]_  = \new_[2402]_  & \new_[2397]_ ;
  assign \new_[2406]_  = A234 & ~A233;
  assign \new_[2410]_  = A299 & ~A298;
  assign \new_[2411]_  = A235 & \new_[2410]_ ;
  assign \new_[2412]_  = \new_[2411]_  & \new_[2406]_ ;
  assign \new_[2415]_  = A167 & A168;
  assign \new_[2419]_  = A232 & ~A201;
  assign \new_[2420]_  = A199 & \new_[2419]_ ;
  assign \new_[2421]_  = \new_[2420]_  & \new_[2415]_ ;
  assign \new_[2424]_  = A234 & ~A233;
  assign \new_[2428]_  = A266 & ~A265;
  assign \new_[2429]_  = A235 & \new_[2428]_ ;
  assign \new_[2430]_  = \new_[2429]_  & \new_[2424]_ ;
  assign \new_[2433]_  = A167 & A168;
  assign \new_[2437]_  = A232 & ~A201;
  assign \new_[2438]_  = A199 & \new_[2437]_ ;
  assign \new_[2439]_  = \new_[2438]_  & \new_[2433]_ ;
  assign \new_[2442]_  = A234 & ~A233;
  assign \new_[2446]_  = A299 & ~A298;
  assign \new_[2447]_  = A236 & \new_[2446]_ ;
  assign \new_[2448]_  = \new_[2447]_  & \new_[2442]_ ;
  assign \new_[2451]_  = A167 & A168;
  assign \new_[2455]_  = A232 & ~A201;
  assign \new_[2456]_  = A199 & \new_[2455]_ ;
  assign \new_[2457]_  = \new_[2456]_  & \new_[2451]_ ;
  assign \new_[2460]_  = A234 & ~A233;
  assign \new_[2464]_  = A266 & ~A265;
  assign \new_[2465]_  = A236 & \new_[2464]_ ;
  assign \new_[2466]_  = \new_[2465]_  & \new_[2460]_ ;
  assign \new_[2469]_  = A167 & A168;
  assign \new_[2473]_  = ~A232 & A200;
  assign \new_[2474]_  = A199 & \new_[2473]_ ;
  assign \new_[2475]_  = \new_[2474]_  & \new_[2469]_ ;
  assign \new_[2478]_  = A298 & A233;
  assign \new_[2482]_  = A301 & A300;
  assign \new_[2483]_  = ~A299 & \new_[2482]_ ;
  assign \new_[2484]_  = \new_[2483]_  & \new_[2478]_ ;
  assign \new_[2487]_  = A167 & A168;
  assign \new_[2491]_  = ~A232 & A200;
  assign \new_[2492]_  = A199 & \new_[2491]_ ;
  assign \new_[2493]_  = \new_[2492]_  & \new_[2487]_ ;
  assign \new_[2496]_  = A298 & A233;
  assign \new_[2500]_  = A302 & A300;
  assign \new_[2501]_  = ~A299 & \new_[2500]_ ;
  assign \new_[2502]_  = \new_[2501]_  & \new_[2496]_ ;
  assign \new_[2505]_  = A167 & A168;
  assign \new_[2509]_  = ~A232 & A200;
  assign \new_[2510]_  = A199 & \new_[2509]_ ;
  assign \new_[2511]_  = \new_[2510]_  & \new_[2505]_ ;
  assign \new_[2514]_  = A265 & A233;
  assign \new_[2518]_  = A268 & A267;
  assign \new_[2519]_  = ~A266 & \new_[2518]_ ;
  assign \new_[2520]_  = \new_[2519]_  & \new_[2514]_ ;
  assign \new_[2523]_  = A167 & A168;
  assign \new_[2527]_  = ~A232 & A200;
  assign \new_[2528]_  = A199 & \new_[2527]_ ;
  assign \new_[2529]_  = \new_[2528]_  & \new_[2523]_ ;
  assign \new_[2532]_  = A265 & A233;
  assign \new_[2536]_  = A269 & A267;
  assign \new_[2537]_  = ~A266 & \new_[2536]_ ;
  assign \new_[2538]_  = \new_[2537]_  & \new_[2532]_ ;
  assign \new_[2541]_  = A167 & A168;
  assign \new_[2545]_  = A232 & A200;
  assign \new_[2546]_  = A199 & \new_[2545]_ ;
  assign \new_[2547]_  = \new_[2546]_  & \new_[2541]_ ;
  assign \new_[2550]_  = A234 & ~A233;
  assign \new_[2554]_  = A299 & ~A298;
  assign \new_[2555]_  = A235 & \new_[2554]_ ;
  assign \new_[2556]_  = \new_[2555]_  & \new_[2550]_ ;
  assign \new_[2559]_  = A167 & A168;
  assign \new_[2563]_  = A232 & A200;
  assign \new_[2564]_  = A199 & \new_[2563]_ ;
  assign \new_[2565]_  = \new_[2564]_  & \new_[2559]_ ;
  assign \new_[2568]_  = A234 & ~A233;
  assign \new_[2572]_  = A266 & ~A265;
  assign \new_[2573]_  = A235 & \new_[2572]_ ;
  assign \new_[2574]_  = \new_[2573]_  & \new_[2568]_ ;
  assign \new_[2577]_  = A167 & A168;
  assign \new_[2581]_  = A232 & A200;
  assign \new_[2582]_  = A199 & \new_[2581]_ ;
  assign \new_[2583]_  = \new_[2582]_  & \new_[2577]_ ;
  assign \new_[2586]_  = A234 & ~A233;
  assign \new_[2590]_  = A299 & ~A298;
  assign \new_[2591]_  = A236 & \new_[2590]_ ;
  assign \new_[2592]_  = \new_[2591]_  & \new_[2586]_ ;
  assign \new_[2595]_  = A167 & A168;
  assign \new_[2599]_  = A232 & A200;
  assign \new_[2600]_  = A199 & \new_[2599]_ ;
  assign \new_[2601]_  = \new_[2600]_  & \new_[2595]_ ;
  assign \new_[2604]_  = A234 & ~A233;
  assign \new_[2608]_  = A266 & ~A265;
  assign \new_[2609]_  = A236 & \new_[2608]_ ;
  assign \new_[2610]_  = \new_[2609]_  & \new_[2604]_ ;
  assign \new_[2613]_  = A167 & A168;
  assign \new_[2617]_  = ~A232 & ~A200;
  assign \new_[2618]_  = ~A199 & \new_[2617]_ ;
  assign \new_[2619]_  = \new_[2618]_  & \new_[2613]_ ;
  assign \new_[2622]_  = A298 & A233;
  assign \new_[2626]_  = A301 & A300;
  assign \new_[2627]_  = ~A299 & \new_[2626]_ ;
  assign \new_[2628]_  = \new_[2627]_  & \new_[2622]_ ;
  assign \new_[2631]_  = A167 & A168;
  assign \new_[2635]_  = ~A232 & ~A200;
  assign \new_[2636]_  = ~A199 & \new_[2635]_ ;
  assign \new_[2637]_  = \new_[2636]_  & \new_[2631]_ ;
  assign \new_[2640]_  = A298 & A233;
  assign \new_[2644]_  = A302 & A300;
  assign \new_[2645]_  = ~A299 & \new_[2644]_ ;
  assign \new_[2646]_  = \new_[2645]_  & \new_[2640]_ ;
  assign \new_[2649]_  = A167 & A168;
  assign \new_[2653]_  = ~A232 & ~A200;
  assign \new_[2654]_  = ~A199 & \new_[2653]_ ;
  assign \new_[2655]_  = \new_[2654]_  & \new_[2649]_ ;
  assign \new_[2658]_  = A265 & A233;
  assign \new_[2662]_  = A268 & A267;
  assign \new_[2663]_  = ~A266 & \new_[2662]_ ;
  assign \new_[2664]_  = \new_[2663]_  & \new_[2658]_ ;
  assign \new_[2667]_  = A167 & A168;
  assign \new_[2671]_  = ~A232 & ~A200;
  assign \new_[2672]_  = ~A199 & \new_[2671]_ ;
  assign \new_[2673]_  = \new_[2672]_  & \new_[2667]_ ;
  assign \new_[2676]_  = A265 & A233;
  assign \new_[2680]_  = A269 & A267;
  assign \new_[2681]_  = ~A266 & \new_[2680]_ ;
  assign \new_[2682]_  = \new_[2681]_  & \new_[2676]_ ;
  assign \new_[2685]_  = A167 & A168;
  assign \new_[2689]_  = A232 & ~A200;
  assign \new_[2690]_  = ~A199 & \new_[2689]_ ;
  assign \new_[2691]_  = \new_[2690]_  & \new_[2685]_ ;
  assign \new_[2694]_  = A234 & ~A233;
  assign \new_[2698]_  = A299 & ~A298;
  assign \new_[2699]_  = A235 & \new_[2698]_ ;
  assign \new_[2700]_  = \new_[2699]_  & \new_[2694]_ ;
  assign \new_[2703]_  = A167 & A168;
  assign \new_[2707]_  = A232 & ~A200;
  assign \new_[2708]_  = ~A199 & \new_[2707]_ ;
  assign \new_[2709]_  = \new_[2708]_  & \new_[2703]_ ;
  assign \new_[2712]_  = A234 & ~A233;
  assign \new_[2716]_  = A266 & ~A265;
  assign \new_[2717]_  = A235 & \new_[2716]_ ;
  assign \new_[2718]_  = \new_[2717]_  & \new_[2712]_ ;
  assign \new_[2721]_  = A167 & A168;
  assign \new_[2725]_  = A232 & ~A200;
  assign \new_[2726]_  = ~A199 & \new_[2725]_ ;
  assign \new_[2727]_  = \new_[2726]_  & \new_[2721]_ ;
  assign \new_[2730]_  = A234 & ~A233;
  assign \new_[2734]_  = A299 & ~A298;
  assign \new_[2735]_  = A236 & \new_[2734]_ ;
  assign \new_[2736]_  = \new_[2735]_  & \new_[2730]_ ;
  assign \new_[2739]_  = A167 & A168;
  assign \new_[2743]_  = A232 & ~A200;
  assign \new_[2744]_  = ~A199 & \new_[2743]_ ;
  assign \new_[2745]_  = \new_[2744]_  & \new_[2739]_ ;
  assign \new_[2748]_  = A234 & ~A233;
  assign \new_[2752]_  = A266 & ~A265;
  assign \new_[2753]_  = A236 & \new_[2752]_ ;
  assign \new_[2754]_  = \new_[2753]_  & \new_[2748]_ ;
  assign \new_[2757]_  = A169 & ~A170;
  assign \new_[2761]_  = A199 & A166;
  assign \new_[2762]_  = A167 & \new_[2761]_ ;
  assign \new_[2763]_  = \new_[2762]_  & \new_[2757]_ ;
  assign \new_[2766]_  = ~A232 & ~A201;
  assign \new_[2770]_  = A299 & ~A298;
  assign \new_[2771]_  = A233 & \new_[2770]_ ;
  assign \new_[2772]_  = \new_[2771]_  & \new_[2766]_ ;
  assign \new_[2775]_  = A169 & ~A170;
  assign \new_[2779]_  = A199 & A166;
  assign \new_[2780]_  = A167 & \new_[2779]_ ;
  assign \new_[2781]_  = \new_[2780]_  & \new_[2775]_ ;
  assign \new_[2784]_  = ~A232 & ~A201;
  assign \new_[2788]_  = A266 & ~A265;
  assign \new_[2789]_  = A233 & \new_[2788]_ ;
  assign \new_[2790]_  = \new_[2789]_  & \new_[2784]_ ;
  assign \new_[2793]_  = A169 & ~A170;
  assign \new_[2797]_  = A199 & A166;
  assign \new_[2798]_  = A167 & \new_[2797]_ ;
  assign \new_[2799]_  = \new_[2798]_  & \new_[2793]_ ;
  assign \new_[2802]_  = ~A232 & A200;
  assign \new_[2806]_  = A299 & ~A298;
  assign \new_[2807]_  = A233 & \new_[2806]_ ;
  assign \new_[2808]_  = \new_[2807]_  & \new_[2802]_ ;
  assign \new_[2811]_  = A169 & ~A170;
  assign \new_[2815]_  = A199 & A166;
  assign \new_[2816]_  = A167 & \new_[2815]_ ;
  assign \new_[2817]_  = \new_[2816]_  & \new_[2811]_ ;
  assign \new_[2820]_  = ~A232 & A200;
  assign \new_[2824]_  = A266 & ~A265;
  assign \new_[2825]_  = A233 & \new_[2824]_ ;
  assign \new_[2826]_  = \new_[2825]_  & \new_[2820]_ ;
  assign \new_[2829]_  = A169 & ~A170;
  assign \new_[2833]_  = ~A199 & A166;
  assign \new_[2834]_  = A167 & \new_[2833]_ ;
  assign \new_[2835]_  = \new_[2834]_  & \new_[2829]_ ;
  assign \new_[2838]_  = ~A232 & ~A200;
  assign \new_[2842]_  = A299 & ~A298;
  assign \new_[2843]_  = A233 & \new_[2842]_ ;
  assign \new_[2844]_  = \new_[2843]_  & \new_[2838]_ ;
  assign \new_[2847]_  = A169 & ~A170;
  assign \new_[2851]_  = ~A199 & A166;
  assign \new_[2852]_  = A167 & \new_[2851]_ ;
  assign \new_[2853]_  = \new_[2852]_  & \new_[2847]_ ;
  assign \new_[2856]_  = ~A232 & ~A200;
  assign \new_[2860]_  = A266 & ~A265;
  assign \new_[2861]_  = A233 & \new_[2860]_ ;
  assign \new_[2862]_  = \new_[2861]_  & \new_[2856]_ ;
  assign \new_[2865]_  = A169 & ~A170;
  assign \new_[2869]_  = A199 & ~A166;
  assign \new_[2870]_  = ~A167 & \new_[2869]_ ;
  assign \new_[2871]_  = \new_[2870]_  & \new_[2865]_ ;
  assign \new_[2874]_  = ~A232 & ~A201;
  assign \new_[2878]_  = A299 & ~A298;
  assign \new_[2879]_  = A233 & \new_[2878]_ ;
  assign \new_[2880]_  = \new_[2879]_  & \new_[2874]_ ;
  assign \new_[2883]_  = A169 & ~A170;
  assign \new_[2887]_  = A199 & ~A166;
  assign \new_[2888]_  = ~A167 & \new_[2887]_ ;
  assign \new_[2889]_  = \new_[2888]_  & \new_[2883]_ ;
  assign \new_[2892]_  = ~A232 & ~A201;
  assign \new_[2896]_  = A266 & ~A265;
  assign \new_[2897]_  = A233 & \new_[2896]_ ;
  assign \new_[2898]_  = \new_[2897]_  & \new_[2892]_ ;
  assign \new_[2901]_  = A169 & ~A170;
  assign \new_[2905]_  = A199 & ~A166;
  assign \new_[2906]_  = ~A167 & \new_[2905]_ ;
  assign \new_[2907]_  = \new_[2906]_  & \new_[2901]_ ;
  assign \new_[2910]_  = ~A232 & A200;
  assign \new_[2914]_  = A299 & ~A298;
  assign \new_[2915]_  = A233 & \new_[2914]_ ;
  assign \new_[2916]_  = \new_[2915]_  & \new_[2910]_ ;
  assign \new_[2919]_  = A169 & ~A170;
  assign \new_[2923]_  = A199 & ~A166;
  assign \new_[2924]_  = ~A167 & \new_[2923]_ ;
  assign \new_[2925]_  = \new_[2924]_  & \new_[2919]_ ;
  assign \new_[2928]_  = ~A232 & A200;
  assign \new_[2932]_  = A266 & ~A265;
  assign \new_[2933]_  = A233 & \new_[2932]_ ;
  assign \new_[2934]_  = \new_[2933]_  & \new_[2928]_ ;
  assign \new_[2937]_  = A169 & ~A170;
  assign \new_[2941]_  = ~A199 & ~A166;
  assign \new_[2942]_  = ~A167 & \new_[2941]_ ;
  assign \new_[2943]_  = \new_[2942]_  & \new_[2937]_ ;
  assign \new_[2946]_  = ~A232 & ~A200;
  assign \new_[2950]_  = A299 & ~A298;
  assign \new_[2951]_  = A233 & \new_[2950]_ ;
  assign \new_[2952]_  = \new_[2951]_  & \new_[2946]_ ;
  assign \new_[2955]_  = A169 & ~A170;
  assign \new_[2959]_  = ~A199 & ~A166;
  assign \new_[2960]_  = ~A167 & \new_[2959]_ ;
  assign \new_[2961]_  = \new_[2960]_  & \new_[2955]_ ;
  assign \new_[2964]_  = ~A232 & ~A200;
  assign \new_[2968]_  = A266 & ~A265;
  assign \new_[2969]_  = A233 & \new_[2968]_ ;
  assign \new_[2970]_  = \new_[2969]_  & \new_[2964]_ ;
  assign \new_[2973]_  = ~A169 & A170;
  assign \new_[2977]_  = A199 & ~A166;
  assign \new_[2978]_  = A167 & \new_[2977]_ ;
  assign \new_[2979]_  = \new_[2978]_  & \new_[2973]_ ;
  assign \new_[2982]_  = ~A232 & ~A201;
  assign \new_[2986]_  = A299 & ~A298;
  assign \new_[2987]_  = A233 & \new_[2986]_ ;
  assign \new_[2988]_  = \new_[2987]_  & \new_[2982]_ ;
  assign \new_[2991]_  = ~A169 & A170;
  assign \new_[2995]_  = A199 & ~A166;
  assign \new_[2996]_  = A167 & \new_[2995]_ ;
  assign \new_[2997]_  = \new_[2996]_  & \new_[2991]_ ;
  assign \new_[3000]_  = ~A232 & ~A201;
  assign \new_[3004]_  = A266 & ~A265;
  assign \new_[3005]_  = A233 & \new_[3004]_ ;
  assign \new_[3006]_  = \new_[3005]_  & \new_[3000]_ ;
  assign \new_[3009]_  = ~A169 & A170;
  assign \new_[3013]_  = A199 & ~A166;
  assign \new_[3014]_  = A167 & \new_[3013]_ ;
  assign \new_[3015]_  = \new_[3014]_  & \new_[3009]_ ;
  assign \new_[3018]_  = ~A232 & A200;
  assign \new_[3022]_  = A299 & ~A298;
  assign \new_[3023]_  = A233 & \new_[3022]_ ;
  assign \new_[3024]_  = \new_[3023]_  & \new_[3018]_ ;
  assign \new_[3027]_  = ~A169 & A170;
  assign \new_[3031]_  = A199 & ~A166;
  assign \new_[3032]_  = A167 & \new_[3031]_ ;
  assign \new_[3033]_  = \new_[3032]_  & \new_[3027]_ ;
  assign \new_[3036]_  = ~A232 & A200;
  assign \new_[3040]_  = A266 & ~A265;
  assign \new_[3041]_  = A233 & \new_[3040]_ ;
  assign \new_[3042]_  = \new_[3041]_  & \new_[3036]_ ;
  assign \new_[3045]_  = ~A169 & A170;
  assign \new_[3049]_  = ~A199 & ~A166;
  assign \new_[3050]_  = A167 & \new_[3049]_ ;
  assign \new_[3051]_  = \new_[3050]_  & \new_[3045]_ ;
  assign \new_[3054]_  = ~A232 & ~A200;
  assign \new_[3058]_  = A299 & ~A298;
  assign \new_[3059]_  = A233 & \new_[3058]_ ;
  assign \new_[3060]_  = \new_[3059]_  & \new_[3054]_ ;
  assign \new_[3063]_  = ~A169 & A170;
  assign \new_[3067]_  = ~A199 & ~A166;
  assign \new_[3068]_  = A167 & \new_[3067]_ ;
  assign \new_[3069]_  = \new_[3068]_  & \new_[3063]_ ;
  assign \new_[3072]_  = ~A232 & ~A200;
  assign \new_[3076]_  = A266 & ~A265;
  assign \new_[3077]_  = A233 & \new_[3076]_ ;
  assign \new_[3078]_  = \new_[3077]_  & \new_[3072]_ ;
  assign \new_[3081]_  = ~A169 & A170;
  assign \new_[3085]_  = A199 & A166;
  assign \new_[3086]_  = ~A167 & \new_[3085]_ ;
  assign \new_[3087]_  = \new_[3086]_  & \new_[3081]_ ;
  assign \new_[3090]_  = ~A232 & ~A201;
  assign \new_[3094]_  = A299 & ~A298;
  assign \new_[3095]_  = A233 & \new_[3094]_ ;
  assign \new_[3096]_  = \new_[3095]_  & \new_[3090]_ ;
  assign \new_[3099]_  = ~A169 & A170;
  assign \new_[3103]_  = A199 & A166;
  assign \new_[3104]_  = ~A167 & \new_[3103]_ ;
  assign \new_[3105]_  = \new_[3104]_  & \new_[3099]_ ;
  assign \new_[3108]_  = ~A232 & ~A201;
  assign \new_[3112]_  = A266 & ~A265;
  assign \new_[3113]_  = A233 & \new_[3112]_ ;
  assign \new_[3114]_  = \new_[3113]_  & \new_[3108]_ ;
  assign \new_[3117]_  = ~A169 & A170;
  assign \new_[3121]_  = A199 & A166;
  assign \new_[3122]_  = ~A167 & \new_[3121]_ ;
  assign \new_[3123]_  = \new_[3122]_  & \new_[3117]_ ;
  assign \new_[3126]_  = ~A232 & A200;
  assign \new_[3130]_  = A299 & ~A298;
  assign \new_[3131]_  = A233 & \new_[3130]_ ;
  assign \new_[3132]_  = \new_[3131]_  & \new_[3126]_ ;
  assign \new_[3135]_  = ~A169 & A170;
  assign \new_[3139]_  = A199 & A166;
  assign \new_[3140]_  = ~A167 & \new_[3139]_ ;
  assign \new_[3141]_  = \new_[3140]_  & \new_[3135]_ ;
  assign \new_[3144]_  = ~A232 & A200;
  assign \new_[3148]_  = A266 & ~A265;
  assign \new_[3149]_  = A233 & \new_[3148]_ ;
  assign \new_[3150]_  = \new_[3149]_  & \new_[3144]_ ;
  assign \new_[3153]_  = ~A169 & A170;
  assign \new_[3157]_  = ~A199 & A166;
  assign \new_[3158]_  = ~A167 & \new_[3157]_ ;
  assign \new_[3159]_  = \new_[3158]_  & \new_[3153]_ ;
  assign \new_[3162]_  = ~A232 & ~A200;
  assign \new_[3166]_  = A299 & ~A298;
  assign \new_[3167]_  = A233 & \new_[3166]_ ;
  assign \new_[3168]_  = \new_[3167]_  & \new_[3162]_ ;
  assign \new_[3171]_  = ~A169 & A170;
  assign \new_[3175]_  = ~A199 & A166;
  assign \new_[3176]_  = ~A167 & \new_[3175]_ ;
  assign \new_[3177]_  = \new_[3176]_  & \new_[3171]_ ;
  assign \new_[3180]_  = ~A232 & ~A200;
  assign \new_[3184]_  = A266 & ~A265;
  assign \new_[3185]_  = A233 & \new_[3184]_ ;
  assign \new_[3186]_  = \new_[3185]_  & \new_[3180]_ ;
  assign \new_[3189]_  = A166 & A168;
  assign \new_[3193]_  = ~A203 & ~A202;
  assign \new_[3194]_  = A199 & \new_[3193]_ ;
  assign \new_[3195]_  = \new_[3194]_  & \new_[3189]_ ;
  assign \new_[3199]_  = A298 & A233;
  assign \new_[3200]_  = ~A232 & \new_[3199]_ ;
  assign \new_[3204]_  = A301 & A300;
  assign \new_[3205]_  = ~A299 & \new_[3204]_ ;
  assign \new_[3206]_  = \new_[3205]_  & \new_[3200]_ ;
  assign \new_[3209]_  = A166 & A168;
  assign \new_[3213]_  = ~A203 & ~A202;
  assign \new_[3214]_  = A199 & \new_[3213]_ ;
  assign \new_[3215]_  = \new_[3214]_  & \new_[3209]_ ;
  assign \new_[3219]_  = A298 & A233;
  assign \new_[3220]_  = ~A232 & \new_[3219]_ ;
  assign \new_[3224]_  = A302 & A300;
  assign \new_[3225]_  = ~A299 & \new_[3224]_ ;
  assign \new_[3226]_  = \new_[3225]_  & \new_[3220]_ ;
  assign \new_[3229]_  = A166 & A168;
  assign \new_[3233]_  = ~A203 & ~A202;
  assign \new_[3234]_  = A199 & \new_[3233]_ ;
  assign \new_[3235]_  = \new_[3234]_  & \new_[3229]_ ;
  assign \new_[3239]_  = A265 & A233;
  assign \new_[3240]_  = ~A232 & \new_[3239]_ ;
  assign \new_[3244]_  = A268 & A267;
  assign \new_[3245]_  = ~A266 & \new_[3244]_ ;
  assign \new_[3246]_  = \new_[3245]_  & \new_[3240]_ ;
  assign \new_[3249]_  = A166 & A168;
  assign \new_[3253]_  = ~A203 & ~A202;
  assign \new_[3254]_  = A199 & \new_[3253]_ ;
  assign \new_[3255]_  = \new_[3254]_  & \new_[3249]_ ;
  assign \new_[3259]_  = A265 & A233;
  assign \new_[3260]_  = ~A232 & \new_[3259]_ ;
  assign \new_[3264]_  = A269 & A267;
  assign \new_[3265]_  = ~A266 & \new_[3264]_ ;
  assign \new_[3266]_  = \new_[3265]_  & \new_[3260]_ ;
  assign \new_[3269]_  = A166 & A168;
  assign \new_[3273]_  = ~A203 & ~A202;
  assign \new_[3274]_  = A199 & \new_[3273]_ ;
  assign \new_[3275]_  = \new_[3274]_  & \new_[3269]_ ;
  assign \new_[3279]_  = A234 & ~A233;
  assign \new_[3280]_  = A232 & \new_[3279]_ ;
  assign \new_[3284]_  = A299 & ~A298;
  assign \new_[3285]_  = A235 & \new_[3284]_ ;
  assign \new_[3286]_  = \new_[3285]_  & \new_[3280]_ ;
  assign \new_[3289]_  = A166 & A168;
  assign \new_[3293]_  = ~A203 & ~A202;
  assign \new_[3294]_  = A199 & \new_[3293]_ ;
  assign \new_[3295]_  = \new_[3294]_  & \new_[3289]_ ;
  assign \new_[3299]_  = A234 & ~A233;
  assign \new_[3300]_  = A232 & \new_[3299]_ ;
  assign \new_[3304]_  = A266 & ~A265;
  assign \new_[3305]_  = A235 & \new_[3304]_ ;
  assign \new_[3306]_  = \new_[3305]_  & \new_[3300]_ ;
  assign \new_[3309]_  = A166 & A168;
  assign \new_[3313]_  = ~A203 & ~A202;
  assign \new_[3314]_  = A199 & \new_[3313]_ ;
  assign \new_[3315]_  = \new_[3314]_  & \new_[3309]_ ;
  assign \new_[3319]_  = A234 & ~A233;
  assign \new_[3320]_  = A232 & \new_[3319]_ ;
  assign \new_[3324]_  = A299 & ~A298;
  assign \new_[3325]_  = A236 & \new_[3324]_ ;
  assign \new_[3326]_  = \new_[3325]_  & \new_[3320]_ ;
  assign \new_[3329]_  = A166 & A168;
  assign \new_[3333]_  = ~A203 & ~A202;
  assign \new_[3334]_  = A199 & \new_[3333]_ ;
  assign \new_[3335]_  = \new_[3334]_  & \new_[3329]_ ;
  assign \new_[3339]_  = A234 & ~A233;
  assign \new_[3340]_  = A232 & \new_[3339]_ ;
  assign \new_[3344]_  = A266 & ~A265;
  assign \new_[3345]_  = A236 & \new_[3344]_ ;
  assign \new_[3346]_  = \new_[3345]_  & \new_[3340]_ ;
  assign \new_[3349]_  = A167 & A168;
  assign \new_[3353]_  = ~A203 & ~A202;
  assign \new_[3354]_  = A199 & \new_[3353]_ ;
  assign \new_[3355]_  = \new_[3354]_  & \new_[3349]_ ;
  assign \new_[3359]_  = A298 & A233;
  assign \new_[3360]_  = ~A232 & \new_[3359]_ ;
  assign \new_[3364]_  = A301 & A300;
  assign \new_[3365]_  = ~A299 & \new_[3364]_ ;
  assign \new_[3366]_  = \new_[3365]_  & \new_[3360]_ ;
  assign \new_[3369]_  = A167 & A168;
  assign \new_[3373]_  = ~A203 & ~A202;
  assign \new_[3374]_  = A199 & \new_[3373]_ ;
  assign \new_[3375]_  = \new_[3374]_  & \new_[3369]_ ;
  assign \new_[3379]_  = A298 & A233;
  assign \new_[3380]_  = ~A232 & \new_[3379]_ ;
  assign \new_[3384]_  = A302 & A300;
  assign \new_[3385]_  = ~A299 & \new_[3384]_ ;
  assign \new_[3386]_  = \new_[3385]_  & \new_[3380]_ ;
  assign \new_[3389]_  = A167 & A168;
  assign \new_[3393]_  = ~A203 & ~A202;
  assign \new_[3394]_  = A199 & \new_[3393]_ ;
  assign \new_[3395]_  = \new_[3394]_  & \new_[3389]_ ;
  assign \new_[3399]_  = A265 & A233;
  assign \new_[3400]_  = ~A232 & \new_[3399]_ ;
  assign \new_[3404]_  = A268 & A267;
  assign \new_[3405]_  = ~A266 & \new_[3404]_ ;
  assign \new_[3406]_  = \new_[3405]_  & \new_[3400]_ ;
  assign \new_[3409]_  = A167 & A168;
  assign \new_[3413]_  = ~A203 & ~A202;
  assign \new_[3414]_  = A199 & \new_[3413]_ ;
  assign \new_[3415]_  = \new_[3414]_  & \new_[3409]_ ;
  assign \new_[3419]_  = A265 & A233;
  assign \new_[3420]_  = ~A232 & \new_[3419]_ ;
  assign \new_[3424]_  = A269 & A267;
  assign \new_[3425]_  = ~A266 & \new_[3424]_ ;
  assign \new_[3426]_  = \new_[3425]_  & \new_[3420]_ ;
  assign \new_[3429]_  = A167 & A168;
  assign \new_[3433]_  = ~A203 & ~A202;
  assign \new_[3434]_  = A199 & \new_[3433]_ ;
  assign \new_[3435]_  = \new_[3434]_  & \new_[3429]_ ;
  assign \new_[3439]_  = A234 & ~A233;
  assign \new_[3440]_  = A232 & \new_[3439]_ ;
  assign \new_[3444]_  = A299 & ~A298;
  assign \new_[3445]_  = A235 & \new_[3444]_ ;
  assign \new_[3446]_  = \new_[3445]_  & \new_[3440]_ ;
  assign \new_[3449]_  = A167 & A168;
  assign \new_[3453]_  = ~A203 & ~A202;
  assign \new_[3454]_  = A199 & \new_[3453]_ ;
  assign \new_[3455]_  = \new_[3454]_  & \new_[3449]_ ;
  assign \new_[3459]_  = A234 & ~A233;
  assign \new_[3460]_  = A232 & \new_[3459]_ ;
  assign \new_[3464]_  = A266 & ~A265;
  assign \new_[3465]_  = A235 & \new_[3464]_ ;
  assign \new_[3466]_  = \new_[3465]_  & \new_[3460]_ ;
  assign \new_[3469]_  = A167 & A168;
  assign \new_[3473]_  = ~A203 & ~A202;
  assign \new_[3474]_  = A199 & \new_[3473]_ ;
  assign \new_[3475]_  = \new_[3474]_  & \new_[3469]_ ;
  assign \new_[3479]_  = A234 & ~A233;
  assign \new_[3480]_  = A232 & \new_[3479]_ ;
  assign \new_[3484]_  = A299 & ~A298;
  assign \new_[3485]_  = A236 & \new_[3484]_ ;
  assign \new_[3486]_  = \new_[3485]_  & \new_[3480]_ ;
  assign \new_[3489]_  = A167 & A168;
  assign \new_[3493]_  = ~A203 & ~A202;
  assign \new_[3494]_  = A199 & \new_[3493]_ ;
  assign \new_[3495]_  = \new_[3494]_  & \new_[3489]_ ;
  assign \new_[3499]_  = A234 & ~A233;
  assign \new_[3500]_  = A232 & \new_[3499]_ ;
  assign \new_[3504]_  = A266 & ~A265;
  assign \new_[3505]_  = A236 & \new_[3504]_ ;
  assign \new_[3506]_  = \new_[3505]_  & \new_[3500]_ ;
  assign \new_[3509]_  = A169 & ~A170;
  assign \new_[3513]_  = A199 & A166;
  assign \new_[3514]_  = A167 & \new_[3513]_ ;
  assign \new_[3515]_  = \new_[3514]_  & \new_[3509]_ ;
  assign \new_[3519]_  = ~A232 & ~A203;
  assign \new_[3520]_  = ~A202 & \new_[3519]_ ;
  assign \new_[3524]_  = A299 & ~A298;
  assign \new_[3525]_  = A233 & \new_[3524]_ ;
  assign \new_[3526]_  = \new_[3525]_  & \new_[3520]_ ;
  assign \new_[3529]_  = A169 & ~A170;
  assign \new_[3533]_  = A199 & A166;
  assign \new_[3534]_  = A167 & \new_[3533]_ ;
  assign \new_[3535]_  = \new_[3534]_  & \new_[3529]_ ;
  assign \new_[3539]_  = ~A232 & ~A203;
  assign \new_[3540]_  = ~A202 & \new_[3539]_ ;
  assign \new_[3544]_  = A266 & ~A265;
  assign \new_[3545]_  = A233 & \new_[3544]_ ;
  assign \new_[3546]_  = \new_[3545]_  & \new_[3540]_ ;
  assign \new_[3549]_  = A169 & ~A170;
  assign \new_[3553]_  = A199 & ~A166;
  assign \new_[3554]_  = ~A167 & \new_[3553]_ ;
  assign \new_[3555]_  = \new_[3554]_  & \new_[3549]_ ;
  assign \new_[3559]_  = ~A232 & ~A203;
  assign \new_[3560]_  = ~A202 & \new_[3559]_ ;
  assign \new_[3564]_  = A299 & ~A298;
  assign \new_[3565]_  = A233 & \new_[3564]_ ;
  assign \new_[3566]_  = \new_[3565]_  & \new_[3560]_ ;
  assign \new_[3569]_  = A169 & ~A170;
  assign \new_[3573]_  = A199 & ~A166;
  assign \new_[3574]_  = ~A167 & \new_[3573]_ ;
  assign \new_[3575]_  = \new_[3574]_  & \new_[3569]_ ;
  assign \new_[3579]_  = ~A232 & ~A203;
  assign \new_[3580]_  = ~A202 & \new_[3579]_ ;
  assign \new_[3584]_  = A266 & ~A265;
  assign \new_[3585]_  = A233 & \new_[3584]_ ;
  assign \new_[3586]_  = \new_[3585]_  & \new_[3580]_ ;
  assign \new_[3589]_  = ~A169 & A170;
  assign \new_[3593]_  = A199 & ~A166;
  assign \new_[3594]_  = A167 & \new_[3593]_ ;
  assign \new_[3595]_  = \new_[3594]_  & \new_[3589]_ ;
  assign \new_[3599]_  = ~A232 & ~A203;
  assign \new_[3600]_  = ~A202 & \new_[3599]_ ;
  assign \new_[3604]_  = A299 & ~A298;
  assign \new_[3605]_  = A233 & \new_[3604]_ ;
  assign \new_[3606]_  = \new_[3605]_  & \new_[3600]_ ;
  assign \new_[3609]_  = ~A169 & A170;
  assign \new_[3613]_  = A199 & ~A166;
  assign \new_[3614]_  = A167 & \new_[3613]_ ;
  assign \new_[3615]_  = \new_[3614]_  & \new_[3609]_ ;
  assign \new_[3619]_  = ~A232 & ~A203;
  assign \new_[3620]_  = ~A202 & \new_[3619]_ ;
  assign \new_[3624]_  = A266 & ~A265;
  assign \new_[3625]_  = A233 & \new_[3624]_ ;
  assign \new_[3626]_  = \new_[3625]_  & \new_[3620]_ ;
  assign \new_[3629]_  = ~A169 & A170;
  assign \new_[3633]_  = A199 & A166;
  assign \new_[3634]_  = ~A167 & \new_[3633]_ ;
  assign \new_[3635]_  = \new_[3634]_  & \new_[3629]_ ;
  assign \new_[3639]_  = ~A232 & ~A203;
  assign \new_[3640]_  = ~A202 & \new_[3639]_ ;
  assign \new_[3644]_  = A299 & ~A298;
  assign \new_[3645]_  = A233 & \new_[3644]_ ;
  assign \new_[3646]_  = \new_[3645]_  & \new_[3640]_ ;
  assign \new_[3649]_  = ~A169 & A170;
  assign \new_[3653]_  = A199 & A166;
  assign \new_[3654]_  = ~A167 & \new_[3653]_ ;
  assign \new_[3655]_  = \new_[3654]_  & \new_[3649]_ ;
  assign \new_[3659]_  = ~A232 & ~A203;
  assign \new_[3660]_  = ~A202 & \new_[3659]_ ;
  assign \new_[3664]_  = A266 & ~A265;
  assign \new_[3665]_  = A233 & \new_[3664]_ ;
  assign \new_[3666]_  = \new_[3665]_  & \new_[3660]_ ;
  assign \new_[3670]_  = A199 & A166;
  assign \new_[3671]_  = A168 & \new_[3670]_ ;
  assign \new_[3675]_  = ~A233 & A232;
  assign \new_[3676]_  = ~A201 & \new_[3675]_ ;
  assign \new_[3677]_  = \new_[3676]_  & \new_[3671]_ ;
  assign \new_[3681]_  = A298 & A235;
  assign \new_[3682]_  = A234 & \new_[3681]_ ;
  assign \new_[3686]_  = A301 & A300;
  assign \new_[3687]_  = ~A299 & \new_[3686]_ ;
  assign \new_[3688]_  = \new_[3687]_  & \new_[3682]_ ;
  assign \new_[3692]_  = A199 & A166;
  assign \new_[3693]_  = A168 & \new_[3692]_ ;
  assign \new_[3697]_  = ~A233 & A232;
  assign \new_[3698]_  = ~A201 & \new_[3697]_ ;
  assign \new_[3699]_  = \new_[3698]_  & \new_[3693]_ ;
  assign \new_[3703]_  = A298 & A235;
  assign \new_[3704]_  = A234 & \new_[3703]_ ;
  assign \new_[3708]_  = A302 & A300;
  assign \new_[3709]_  = ~A299 & \new_[3708]_ ;
  assign \new_[3710]_  = \new_[3709]_  & \new_[3704]_ ;
  assign \new_[3714]_  = A199 & A166;
  assign \new_[3715]_  = A168 & \new_[3714]_ ;
  assign \new_[3719]_  = ~A233 & A232;
  assign \new_[3720]_  = ~A201 & \new_[3719]_ ;
  assign \new_[3721]_  = \new_[3720]_  & \new_[3715]_ ;
  assign \new_[3725]_  = A265 & A235;
  assign \new_[3726]_  = A234 & \new_[3725]_ ;
  assign \new_[3730]_  = A268 & A267;
  assign \new_[3731]_  = ~A266 & \new_[3730]_ ;
  assign \new_[3732]_  = \new_[3731]_  & \new_[3726]_ ;
  assign \new_[3736]_  = A199 & A166;
  assign \new_[3737]_  = A168 & \new_[3736]_ ;
  assign \new_[3741]_  = ~A233 & A232;
  assign \new_[3742]_  = ~A201 & \new_[3741]_ ;
  assign \new_[3743]_  = \new_[3742]_  & \new_[3737]_ ;
  assign \new_[3747]_  = A265 & A235;
  assign \new_[3748]_  = A234 & \new_[3747]_ ;
  assign \new_[3752]_  = A269 & A267;
  assign \new_[3753]_  = ~A266 & \new_[3752]_ ;
  assign \new_[3754]_  = \new_[3753]_  & \new_[3748]_ ;
  assign \new_[3758]_  = A199 & A166;
  assign \new_[3759]_  = A168 & \new_[3758]_ ;
  assign \new_[3763]_  = ~A233 & A232;
  assign \new_[3764]_  = ~A201 & \new_[3763]_ ;
  assign \new_[3765]_  = \new_[3764]_  & \new_[3759]_ ;
  assign \new_[3769]_  = A298 & A236;
  assign \new_[3770]_  = A234 & \new_[3769]_ ;
  assign \new_[3774]_  = A301 & A300;
  assign \new_[3775]_  = ~A299 & \new_[3774]_ ;
  assign \new_[3776]_  = \new_[3775]_  & \new_[3770]_ ;
  assign \new_[3780]_  = A199 & A166;
  assign \new_[3781]_  = A168 & \new_[3780]_ ;
  assign \new_[3785]_  = ~A233 & A232;
  assign \new_[3786]_  = ~A201 & \new_[3785]_ ;
  assign \new_[3787]_  = \new_[3786]_  & \new_[3781]_ ;
  assign \new_[3791]_  = A298 & A236;
  assign \new_[3792]_  = A234 & \new_[3791]_ ;
  assign \new_[3796]_  = A302 & A300;
  assign \new_[3797]_  = ~A299 & \new_[3796]_ ;
  assign \new_[3798]_  = \new_[3797]_  & \new_[3792]_ ;
  assign \new_[3802]_  = A199 & A166;
  assign \new_[3803]_  = A168 & \new_[3802]_ ;
  assign \new_[3807]_  = ~A233 & A232;
  assign \new_[3808]_  = ~A201 & \new_[3807]_ ;
  assign \new_[3809]_  = \new_[3808]_  & \new_[3803]_ ;
  assign \new_[3813]_  = A265 & A236;
  assign \new_[3814]_  = A234 & \new_[3813]_ ;
  assign \new_[3818]_  = A268 & A267;
  assign \new_[3819]_  = ~A266 & \new_[3818]_ ;
  assign \new_[3820]_  = \new_[3819]_  & \new_[3814]_ ;
  assign \new_[3824]_  = A199 & A166;
  assign \new_[3825]_  = A168 & \new_[3824]_ ;
  assign \new_[3829]_  = ~A233 & A232;
  assign \new_[3830]_  = ~A201 & \new_[3829]_ ;
  assign \new_[3831]_  = \new_[3830]_  & \new_[3825]_ ;
  assign \new_[3835]_  = A265 & A236;
  assign \new_[3836]_  = A234 & \new_[3835]_ ;
  assign \new_[3840]_  = A269 & A267;
  assign \new_[3841]_  = ~A266 & \new_[3840]_ ;
  assign \new_[3842]_  = \new_[3841]_  & \new_[3836]_ ;
  assign \new_[3846]_  = A199 & A166;
  assign \new_[3847]_  = A168 & \new_[3846]_ ;
  assign \new_[3851]_  = ~A233 & A232;
  assign \new_[3852]_  = A200 & \new_[3851]_ ;
  assign \new_[3853]_  = \new_[3852]_  & \new_[3847]_ ;
  assign \new_[3857]_  = A298 & A235;
  assign \new_[3858]_  = A234 & \new_[3857]_ ;
  assign \new_[3862]_  = A301 & A300;
  assign \new_[3863]_  = ~A299 & \new_[3862]_ ;
  assign \new_[3864]_  = \new_[3863]_  & \new_[3858]_ ;
  assign \new_[3868]_  = A199 & A166;
  assign \new_[3869]_  = A168 & \new_[3868]_ ;
  assign \new_[3873]_  = ~A233 & A232;
  assign \new_[3874]_  = A200 & \new_[3873]_ ;
  assign \new_[3875]_  = \new_[3874]_  & \new_[3869]_ ;
  assign \new_[3879]_  = A298 & A235;
  assign \new_[3880]_  = A234 & \new_[3879]_ ;
  assign \new_[3884]_  = A302 & A300;
  assign \new_[3885]_  = ~A299 & \new_[3884]_ ;
  assign \new_[3886]_  = \new_[3885]_  & \new_[3880]_ ;
  assign \new_[3890]_  = A199 & A166;
  assign \new_[3891]_  = A168 & \new_[3890]_ ;
  assign \new_[3895]_  = ~A233 & A232;
  assign \new_[3896]_  = A200 & \new_[3895]_ ;
  assign \new_[3897]_  = \new_[3896]_  & \new_[3891]_ ;
  assign \new_[3901]_  = A265 & A235;
  assign \new_[3902]_  = A234 & \new_[3901]_ ;
  assign \new_[3906]_  = A268 & A267;
  assign \new_[3907]_  = ~A266 & \new_[3906]_ ;
  assign \new_[3908]_  = \new_[3907]_  & \new_[3902]_ ;
  assign \new_[3912]_  = A199 & A166;
  assign \new_[3913]_  = A168 & \new_[3912]_ ;
  assign \new_[3917]_  = ~A233 & A232;
  assign \new_[3918]_  = A200 & \new_[3917]_ ;
  assign \new_[3919]_  = \new_[3918]_  & \new_[3913]_ ;
  assign \new_[3923]_  = A265 & A235;
  assign \new_[3924]_  = A234 & \new_[3923]_ ;
  assign \new_[3928]_  = A269 & A267;
  assign \new_[3929]_  = ~A266 & \new_[3928]_ ;
  assign \new_[3930]_  = \new_[3929]_  & \new_[3924]_ ;
  assign \new_[3934]_  = A199 & A166;
  assign \new_[3935]_  = A168 & \new_[3934]_ ;
  assign \new_[3939]_  = ~A233 & A232;
  assign \new_[3940]_  = A200 & \new_[3939]_ ;
  assign \new_[3941]_  = \new_[3940]_  & \new_[3935]_ ;
  assign \new_[3945]_  = A298 & A236;
  assign \new_[3946]_  = A234 & \new_[3945]_ ;
  assign \new_[3950]_  = A301 & A300;
  assign \new_[3951]_  = ~A299 & \new_[3950]_ ;
  assign \new_[3952]_  = \new_[3951]_  & \new_[3946]_ ;
  assign \new_[3956]_  = A199 & A166;
  assign \new_[3957]_  = A168 & \new_[3956]_ ;
  assign \new_[3961]_  = ~A233 & A232;
  assign \new_[3962]_  = A200 & \new_[3961]_ ;
  assign \new_[3963]_  = \new_[3962]_  & \new_[3957]_ ;
  assign \new_[3967]_  = A298 & A236;
  assign \new_[3968]_  = A234 & \new_[3967]_ ;
  assign \new_[3972]_  = A302 & A300;
  assign \new_[3973]_  = ~A299 & \new_[3972]_ ;
  assign \new_[3974]_  = \new_[3973]_  & \new_[3968]_ ;
  assign \new_[3978]_  = A199 & A166;
  assign \new_[3979]_  = A168 & \new_[3978]_ ;
  assign \new_[3983]_  = ~A233 & A232;
  assign \new_[3984]_  = A200 & \new_[3983]_ ;
  assign \new_[3985]_  = \new_[3984]_  & \new_[3979]_ ;
  assign \new_[3989]_  = A265 & A236;
  assign \new_[3990]_  = A234 & \new_[3989]_ ;
  assign \new_[3994]_  = A268 & A267;
  assign \new_[3995]_  = ~A266 & \new_[3994]_ ;
  assign \new_[3996]_  = \new_[3995]_  & \new_[3990]_ ;
  assign \new_[4000]_  = A199 & A166;
  assign \new_[4001]_  = A168 & \new_[4000]_ ;
  assign \new_[4005]_  = ~A233 & A232;
  assign \new_[4006]_  = A200 & \new_[4005]_ ;
  assign \new_[4007]_  = \new_[4006]_  & \new_[4001]_ ;
  assign \new_[4011]_  = A265 & A236;
  assign \new_[4012]_  = A234 & \new_[4011]_ ;
  assign \new_[4016]_  = A269 & A267;
  assign \new_[4017]_  = ~A266 & \new_[4016]_ ;
  assign \new_[4018]_  = \new_[4017]_  & \new_[4012]_ ;
  assign \new_[4022]_  = ~A199 & A166;
  assign \new_[4023]_  = A168 & \new_[4022]_ ;
  assign \new_[4027]_  = ~A233 & A232;
  assign \new_[4028]_  = ~A200 & \new_[4027]_ ;
  assign \new_[4029]_  = \new_[4028]_  & \new_[4023]_ ;
  assign \new_[4033]_  = A298 & A235;
  assign \new_[4034]_  = A234 & \new_[4033]_ ;
  assign \new_[4038]_  = A301 & A300;
  assign \new_[4039]_  = ~A299 & \new_[4038]_ ;
  assign \new_[4040]_  = \new_[4039]_  & \new_[4034]_ ;
  assign \new_[4044]_  = ~A199 & A166;
  assign \new_[4045]_  = A168 & \new_[4044]_ ;
  assign \new_[4049]_  = ~A233 & A232;
  assign \new_[4050]_  = ~A200 & \new_[4049]_ ;
  assign \new_[4051]_  = \new_[4050]_  & \new_[4045]_ ;
  assign \new_[4055]_  = A298 & A235;
  assign \new_[4056]_  = A234 & \new_[4055]_ ;
  assign \new_[4060]_  = A302 & A300;
  assign \new_[4061]_  = ~A299 & \new_[4060]_ ;
  assign \new_[4062]_  = \new_[4061]_  & \new_[4056]_ ;
  assign \new_[4066]_  = ~A199 & A166;
  assign \new_[4067]_  = A168 & \new_[4066]_ ;
  assign \new_[4071]_  = ~A233 & A232;
  assign \new_[4072]_  = ~A200 & \new_[4071]_ ;
  assign \new_[4073]_  = \new_[4072]_  & \new_[4067]_ ;
  assign \new_[4077]_  = A265 & A235;
  assign \new_[4078]_  = A234 & \new_[4077]_ ;
  assign \new_[4082]_  = A268 & A267;
  assign \new_[4083]_  = ~A266 & \new_[4082]_ ;
  assign \new_[4084]_  = \new_[4083]_  & \new_[4078]_ ;
  assign \new_[4088]_  = ~A199 & A166;
  assign \new_[4089]_  = A168 & \new_[4088]_ ;
  assign \new_[4093]_  = ~A233 & A232;
  assign \new_[4094]_  = ~A200 & \new_[4093]_ ;
  assign \new_[4095]_  = \new_[4094]_  & \new_[4089]_ ;
  assign \new_[4099]_  = A265 & A235;
  assign \new_[4100]_  = A234 & \new_[4099]_ ;
  assign \new_[4104]_  = A269 & A267;
  assign \new_[4105]_  = ~A266 & \new_[4104]_ ;
  assign \new_[4106]_  = \new_[4105]_  & \new_[4100]_ ;
  assign \new_[4110]_  = ~A199 & A166;
  assign \new_[4111]_  = A168 & \new_[4110]_ ;
  assign \new_[4115]_  = ~A233 & A232;
  assign \new_[4116]_  = ~A200 & \new_[4115]_ ;
  assign \new_[4117]_  = \new_[4116]_  & \new_[4111]_ ;
  assign \new_[4121]_  = A298 & A236;
  assign \new_[4122]_  = A234 & \new_[4121]_ ;
  assign \new_[4126]_  = A301 & A300;
  assign \new_[4127]_  = ~A299 & \new_[4126]_ ;
  assign \new_[4128]_  = \new_[4127]_  & \new_[4122]_ ;
  assign \new_[4132]_  = ~A199 & A166;
  assign \new_[4133]_  = A168 & \new_[4132]_ ;
  assign \new_[4137]_  = ~A233 & A232;
  assign \new_[4138]_  = ~A200 & \new_[4137]_ ;
  assign \new_[4139]_  = \new_[4138]_  & \new_[4133]_ ;
  assign \new_[4143]_  = A298 & A236;
  assign \new_[4144]_  = A234 & \new_[4143]_ ;
  assign \new_[4148]_  = A302 & A300;
  assign \new_[4149]_  = ~A299 & \new_[4148]_ ;
  assign \new_[4150]_  = \new_[4149]_  & \new_[4144]_ ;
  assign \new_[4154]_  = ~A199 & A166;
  assign \new_[4155]_  = A168 & \new_[4154]_ ;
  assign \new_[4159]_  = ~A233 & A232;
  assign \new_[4160]_  = ~A200 & \new_[4159]_ ;
  assign \new_[4161]_  = \new_[4160]_  & \new_[4155]_ ;
  assign \new_[4165]_  = A265 & A236;
  assign \new_[4166]_  = A234 & \new_[4165]_ ;
  assign \new_[4170]_  = A268 & A267;
  assign \new_[4171]_  = ~A266 & \new_[4170]_ ;
  assign \new_[4172]_  = \new_[4171]_  & \new_[4166]_ ;
  assign \new_[4176]_  = ~A199 & A166;
  assign \new_[4177]_  = A168 & \new_[4176]_ ;
  assign \new_[4181]_  = ~A233 & A232;
  assign \new_[4182]_  = ~A200 & \new_[4181]_ ;
  assign \new_[4183]_  = \new_[4182]_  & \new_[4177]_ ;
  assign \new_[4187]_  = A265 & A236;
  assign \new_[4188]_  = A234 & \new_[4187]_ ;
  assign \new_[4192]_  = A269 & A267;
  assign \new_[4193]_  = ~A266 & \new_[4192]_ ;
  assign \new_[4194]_  = \new_[4193]_  & \new_[4188]_ ;
  assign \new_[4198]_  = A199 & A167;
  assign \new_[4199]_  = A168 & \new_[4198]_ ;
  assign \new_[4203]_  = ~A233 & A232;
  assign \new_[4204]_  = ~A201 & \new_[4203]_ ;
  assign \new_[4205]_  = \new_[4204]_  & \new_[4199]_ ;
  assign \new_[4209]_  = A298 & A235;
  assign \new_[4210]_  = A234 & \new_[4209]_ ;
  assign \new_[4214]_  = A301 & A300;
  assign \new_[4215]_  = ~A299 & \new_[4214]_ ;
  assign \new_[4216]_  = \new_[4215]_  & \new_[4210]_ ;
  assign \new_[4220]_  = A199 & A167;
  assign \new_[4221]_  = A168 & \new_[4220]_ ;
  assign \new_[4225]_  = ~A233 & A232;
  assign \new_[4226]_  = ~A201 & \new_[4225]_ ;
  assign \new_[4227]_  = \new_[4226]_  & \new_[4221]_ ;
  assign \new_[4231]_  = A298 & A235;
  assign \new_[4232]_  = A234 & \new_[4231]_ ;
  assign \new_[4236]_  = A302 & A300;
  assign \new_[4237]_  = ~A299 & \new_[4236]_ ;
  assign \new_[4238]_  = \new_[4237]_  & \new_[4232]_ ;
  assign \new_[4242]_  = A199 & A167;
  assign \new_[4243]_  = A168 & \new_[4242]_ ;
  assign \new_[4247]_  = ~A233 & A232;
  assign \new_[4248]_  = ~A201 & \new_[4247]_ ;
  assign \new_[4249]_  = \new_[4248]_  & \new_[4243]_ ;
  assign \new_[4253]_  = A265 & A235;
  assign \new_[4254]_  = A234 & \new_[4253]_ ;
  assign \new_[4258]_  = A268 & A267;
  assign \new_[4259]_  = ~A266 & \new_[4258]_ ;
  assign \new_[4260]_  = \new_[4259]_  & \new_[4254]_ ;
  assign \new_[4264]_  = A199 & A167;
  assign \new_[4265]_  = A168 & \new_[4264]_ ;
  assign \new_[4269]_  = ~A233 & A232;
  assign \new_[4270]_  = ~A201 & \new_[4269]_ ;
  assign \new_[4271]_  = \new_[4270]_  & \new_[4265]_ ;
  assign \new_[4275]_  = A265 & A235;
  assign \new_[4276]_  = A234 & \new_[4275]_ ;
  assign \new_[4280]_  = A269 & A267;
  assign \new_[4281]_  = ~A266 & \new_[4280]_ ;
  assign \new_[4282]_  = \new_[4281]_  & \new_[4276]_ ;
  assign \new_[4286]_  = A199 & A167;
  assign \new_[4287]_  = A168 & \new_[4286]_ ;
  assign \new_[4291]_  = ~A233 & A232;
  assign \new_[4292]_  = ~A201 & \new_[4291]_ ;
  assign \new_[4293]_  = \new_[4292]_  & \new_[4287]_ ;
  assign \new_[4297]_  = A298 & A236;
  assign \new_[4298]_  = A234 & \new_[4297]_ ;
  assign \new_[4302]_  = A301 & A300;
  assign \new_[4303]_  = ~A299 & \new_[4302]_ ;
  assign \new_[4304]_  = \new_[4303]_  & \new_[4298]_ ;
  assign \new_[4308]_  = A199 & A167;
  assign \new_[4309]_  = A168 & \new_[4308]_ ;
  assign \new_[4313]_  = ~A233 & A232;
  assign \new_[4314]_  = ~A201 & \new_[4313]_ ;
  assign \new_[4315]_  = \new_[4314]_  & \new_[4309]_ ;
  assign \new_[4319]_  = A298 & A236;
  assign \new_[4320]_  = A234 & \new_[4319]_ ;
  assign \new_[4324]_  = A302 & A300;
  assign \new_[4325]_  = ~A299 & \new_[4324]_ ;
  assign \new_[4326]_  = \new_[4325]_  & \new_[4320]_ ;
  assign \new_[4330]_  = A199 & A167;
  assign \new_[4331]_  = A168 & \new_[4330]_ ;
  assign \new_[4335]_  = ~A233 & A232;
  assign \new_[4336]_  = ~A201 & \new_[4335]_ ;
  assign \new_[4337]_  = \new_[4336]_  & \new_[4331]_ ;
  assign \new_[4341]_  = A265 & A236;
  assign \new_[4342]_  = A234 & \new_[4341]_ ;
  assign \new_[4346]_  = A268 & A267;
  assign \new_[4347]_  = ~A266 & \new_[4346]_ ;
  assign \new_[4348]_  = \new_[4347]_  & \new_[4342]_ ;
  assign \new_[4352]_  = A199 & A167;
  assign \new_[4353]_  = A168 & \new_[4352]_ ;
  assign \new_[4357]_  = ~A233 & A232;
  assign \new_[4358]_  = ~A201 & \new_[4357]_ ;
  assign \new_[4359]_  = \new_[4358]_  & \new_[4353]_ ;
  assign \new_[4363]_  = A265 & A236;
  assign \new_[4364]_  = A234 & \new_[4363]_ ;
  assign \new_[4368]_  = A269 & A267;
  assign \new_[4369]_  = ~A266 & \new_[4368]_ ;
  assign \new_[4370]_  = \new_[4369]_  & \new_[4364]_ ;
  assign \new_[4374]_  = A199 & A167;
  assign \new_[4375]_  = A168 & \new_[4374]_ ;
  assign \new_[4379]_  = ~A233 & A232;
  assign \new_[4380]_  = A200 & \new_[4379]_ ;
  assign \new_[4381]_  = \new_[4380]_  & \new_[4375]_ ;
  assign \new_[4385]_  = A298 & A235;
  assign \new_[4386]_  = A234 & \new_[4385]_ ;
  assign \new_[4390]_  = A301 & A300;
  assign \new_[4391]_  = ~A299 & \new_[4390]_ ;
  assign \new_[4392]_  = \new_[4391]_  & \new_[4386]_ ;
  assign \new_[4396]_  = A199 & A167;
  assign \new_[4397]_  = A168 & \new_[4396]_ ;
  assign \new_[4401]_  = ~A233 & A232;
  assign \new_[4402]_  = A200 & \new_[4401]_ ;
  assign \new_[4403]_  = \new_[4402]_  & \new_[4397]_ ;
  assign \new_[4407]_  = A298 & A235;
  assign \new_[4408]_  = A234 & \new_[4407]_ ;
  assign \new_[4412]_  = A302 & A300;
  assign \new_[4413]_  = ~A299 & \new_[4412]_ ;
  assign \new_[4414]_  = \new_[4413]_  & \new_[4408]_ ;
  assign \new_[4418]_  = A199 & A167;
  assign \new_[4419]_  = A168 & \new_[4418]_ ;
  assign \new_[4423]_  = ~A233 & A232;
  assign \new_[4424]_  = A200 & \new_[4423]_ ;
  assign \new_[4425]_  = \new_[4424]_  & \new_[4419]_ ;
  assign \new_[4429]_  = A265 & A235;
  assign \new_[4430]_  = A234 & \new_[4429]_ ;
  assign \new_[4434]_  = A268 & A267;
  assign \new_[4435]_  = ~A266 & \new_[4434]_ ;
  assign \new_[4436]_  = \new_[4435]_  & \new_[4430]_ ;
  assign \new_[4440]_  = A199 & A167;
  assign \new_[4441]_  = A168 & \new_[4440]_ ;
  assign \new_[4445]_  = ~A233 & A232;
  assign \new_[4446]_  = A200 & \new_[4445]_ ;
  assign \new_[4447]_  = \new_[4446]_  & \new_[4441]_ ;
  assign \new_[4451]_  = A265 & A235;
  assign \new_[4452]_  = A234 & \new_[4451]_ ;
  assign \new_[4456]_  = A269 & A267;
  assign \new_[4457]_  = ~A266 & \new_[4456]_ ;
  assign \new_[4458]_  = \new_[4457]_  & \new_[4452]_ ;
  assign \new_[4462]_  = A199 & A167;
  assign \new_[4463]_  = A168 & \new_[4462]_ ;
  assign \new_[4467]_  = ~A233 & A232;
  assign \new_[4468]_  = A200 & \new_[4467]_ ;
  assign \new_[4469]_  = \new_[4468]_  & \new_[4463]_ ;
  assign \new_[4473]_  = A298 & A236;
  assign \new_[4474]_  = A234 & \new_[4473]_ ;
  assign \new_[4478]_  = A301 & A300;
  assign \new_[4479]_  = ~A299 & \new_[4478]_ ;
  assign \new_[4480]_  = \new_[4479]_  & \new_[4474]_ ;
  assign \new_[4484]_  = A199 & A167;
  assign \new_[4485]_  = A168 & \new_[4484]_ ;
  assign \new_[4489]_  = ~A233 & A232;
  assign \new_[4490]_  = A200 & \new_[4489]_ ;
  assign \new_[4491]_  = \new_[4490]_  & \new_[4485]_ ;
  assign \new_[4495]_  = A298 & A236;
  assign \new_[4496]_  = A234 & \new_[4495]_ ;
  assign \new_[4500]_  = A302 & A300;
  assign \new_[4501]_  = ~A299 & \new_[4500]_ ;
  assign \new_[4502]_  = \new_[4501]_  & \new_[4496]_ ;
  assign \new_[4506]_  = A199 & A167;
  assign \new_[4507]_  = A168 & \new_[4506]_ ;
  assign \new_[4511]_  = ~A233 & A232;
  assign \new_[4512]_  = A200 & \new_[4511]_ ;
  assign \new_[4513]_  = \new_[4512]_  & \new_[4507]_ ;
  assign \new_[4517]_  = A265 & A236;
  assign \new_[4518]_  = A234 & \new_[4517]_ ;
  assign \new_[4522]_  = A268 & A267;
  assign \new_[4523]_  = ~A266 & \new_[4522]_ ;
  assign \new_[4524]_  = \new_[4523]_  & \new_[4518]_ ;
  assign \new_[4528]_  = A199 & A167;
  assign \new_[4529]_  = A168 & \new_[4528]_ ;
  assign \new_[4533]_  = ~A233 & A232;
  assign \new_[4534]_  = A200 & \new_[4533]_ ;
  assign \new_[4535]_  = \new_[4534]_  & \new_[4529]_ ;
  assign \new_[4539]_  = A265 & A236;
  assign \new_[4540]_  = A234 & \new_[4539]_ ;
  assign \new_[4544]_  = A269 & A267;
  assign \new_[4545]_  = ~A266 & \new_[4544]_ ;
  assign \new_[4546]_  = \new_[4545]_  & \new_[4540]_ ;
  assign \new_[4550]_  = ~A199 & A167;
  assign \new_[4551]_  = A168 & \new_[4550]_ ;
  assign \new_[4555]_  = ~A233 & A232;
  assign \new_[4556]_  = ~A200 & \new_[4555]_ ;
  assign \new_[4557]_  = \new_[4556]_  & \new_[4551]_ ;
  assign \new_[4561]_  = A298 & A235;
  assign \new_[4562]_  = A234 & \new_[4561]_ ;
  assign \new_[4566]_  = A301 & A300;
  assign \new_[4567]_  = ~A299 & \new_[4566]_ ;
  assign \new_[4568]_  = \new_[4567]_  & \new_[4562]_ ;
  assign \new_[4572]_  = ~A199 & A167;
  assign \new_[4573]_  = A168 & \new_[4572]_ ;
  assign \new_[4577]_  = ~A233 & A232;
  assign \new_[4578]_  = ~A200 & \new_[4577]_ ;
  assign \new_[4579]_  = \new_[4578]_  & \new_[4573]_ ;
  assign \new_[4583]_  = A298 & A235;
  assign \new_[4584]_  = A234 & \new_[4583]_ ;
  assign \new_[4588]_  = A302 & A300;
  assign \new_[4589]_  = ~A299 & \new_[4588]_ ;
  assign \new_[4590]_  = \new_[4589]_  & \new_[4584]_ ;
  assign \new_[4594]_  = ~A199 & A167;
  assign \new_[4595]_  = A168 & \new_[4594]_ ;
  assign \new_[4599]_  = ~A233 & A232;
  assign \new_[4600]_  = ~A200 & \new_[4599]_ ;
  assign \new_[4601]_  = \new_[4600]_  & \new_[4595]_ ;
  assign \new_[4605]_  = A265 & A235;
  assign \new_[4606]_  = A234 & \new_[4605]_ ;
  assign \new_[4610]_  = A268 & A267;
  assign \new_[4611]_  = ~A266 & \new_[4610]_ ;
  assign \new_[4612]_  = \new_[4611]_  & \new_[4606]_ ;
  assign \new_[4616]_  = ~A199 & A167;
  assign \new_[4617]_  = A168 & \new_[4616]_ ;
  assign \new_[4621]_  = ~A233 & A232;
  assign \new_[4622]_  = ~A200 & \new_[4621]_ ;
  assign \new_[4623]_  = \new_[4622]_  & \new_[4617]_ ;
  assign \new_[4627]_  = A265 & A235;
  assign \new_[4628]_  = A234 & \new_[4627]_ ;
  assign \new_[4632]_  = A269 & A267;
  assign \new_[4633]_  = ~A266 & \new_[4632]_ ;
  assign \new_[4634]_  = \new_[4633]_  & \new_[4628]_ ;
  assign \new_[4638]_  = ~A199 & A167;
  assign \new_[4639]_  = A168 & \new_[4638]_ ;
  assign \new_[4643]_  = ~A233 & A232;
  assign \new_[4644]_  = ~A200 & \new_[4643]_ ;
  assign \new_[4645]_  = \new_[4644]_  & \new_[4639]_ ;
  assign \new_[4649]_  = A298 & A236;
  assign \new_[4650]_  = A234 & \new_[4649]_ ;
  assign \new_[4654]_  = A301 & A300;
  assign \new_[4655]_  = ~A299 & \new_[4654]_ ;
  assign \new_[4656]_  = \new_[4655]_  & \new_[4650]_ ;
  assign \new_[4660]_  = ~A199 & A167;
  assign \new_[4661]_  = A168 & \new_[4660]_ ;
  assign \new_[4665]_  = ~A233 & A232;
  assign \new_[4666]_  = ~A200 & \new_[4665]_ ;
  assign \new_[4667]_  = \new_[4666]_  & \new_[4661]_ ;
  assign \new_[4671]_  = A298 & A236;
  assign \new_[4672]_  = A234 & \new_[4671]_ ;
  assign \new_[4676]_  = A302 & A300;
  assign \new_[4677]_  = ~A299 & \new_[4676]_ ;
  assign \new_[4678]_  = \new_[4677]_  & \new_[4672]_ ;
  assign \new_[4682]_  = ~A199 & A167;
  assign \new_[4683]_  = A168 & \new_[4682]_ ;
  assign \new_[4687]_  = ~A233 & A232;
  assign \new_[4688]_  = ~A200 & \new_[4687]_ ;
  assign \new_[4689]_  = \new_[4688]_  & \new_[4683]_ ;
  assign \new_[4693]_  = A265 & A236;
  assign \new_[4694]_  = A234 & \new_[4693]_ ;
  assign \new_[4698]_  = A268 & A267;
  assign \new_[4699]_  = ~A266 & \new_[4698]_ ;
  assign \new_[4700]_  = \new_[4699]_  & \new_[4694]_ ;
  assign \new_[4704]_  = ~A199 & A167;
  assign \new_[4705]_  = A168 & \new_[4704]_ ;
  assign \new_[4709]_  = ~A233 & A232;
  assign \new_[4710]_  = ~A200 & \new_[4709]_ ;
  assign \new_[4711]_  = \new_[4710]_  & \new_[4705]_ ;
  assign \new_[4715]_  = A265 & A236;
  assign \new_[4716]_  = A234 & \new_[4715]_ ;
  assign \new_[4720]_  = A269 & A267;
  assign \new_[4721]_  = ~A266 & \new_[4720]_ ;
  assign \new_[4722]_  = \new_[4721]_  & \new_[4716]_ ;
  assign \new_[4726]_  = A167 & A169;
  assign \new_[4727]_  = ~A170 & \new_[4726]_ ;
  assign \new_[4731]_  = ~A201 & A199;
  assign \new_[4732]_  = A166 & \new_[4731]_ ;
  assign \new_[4733]_  = \new_[4732]_  & \new_[4727]_ ;
  assign \new_[4737]_  = A298 & A233;
  assign \new_[4738]_  = ~A232 & \new_[4737]_ ;
  assign \new_[4742]_  = A301 & A300;
  assign \new_[4743]_  = ~A299 & \new_[4742]_ ;
  assign \new_[4744]_  = \new_[4743]_  & \new_[4738]_ ;
  assign \new_[4748]_  = A167 & A169;
  assign \new_[4749]_  = ~A170 & \new_[4748]_ ;
  assign \new_[4753]_  = ~A201 & A199;
  assign \new_[4754]_  = A166 & \new_[4753]_ ;
  assign \new_[4755]_  = \new_[4754]_  & \new_[4749]_ ;
  assign \new_[4759]_  = A298 & A233;
  assign \new_[4760]_  = ~A232 & \new_[4759]_ ;
  assign \new_[4764]_  = A302 & A300;
  assign \new_[4765]_  = ~A299 & \new_[4764]_ ;
  assign \new_[4766]_  = \new_[4765]_  & \new_[4760]_ ;
  assign \new_[4770]_  = A167 & A169;
  assign \new_[4771]_  = ~A170 & \new_[4770]_ ;
  assign \new_[4775]_  = ~A201 & A199;
  assign \new_[4776]_  = A166 & \new_[4775]_ ;
  assign \new_[4777]_  = \new_[4776]_  & \new_[4771]_ ;
  assign \new_[4781]_  = A265 & A233;
  assign \new_[4782]_  = ~A232 & \new_[4781]_ ;
  assign \new_[4786]_  = A268 & A267;
  assign \new_[4787]_  = ~A266 & \new_[4786]_ ;
  assign \new_[4788]_  = \new_[4787]_  & \new_[4782]_ ;
  assign \new_[4792]_  = A167 & A169;
  assign \new_[4793]_  = ~A170 & \new_[4792]_ ;
  assign \new_[4797]_  = ~A201 & A199;
  assign \new_[4798]_  = A166 & \new_[4797]_ ;
  assign \new_[4799]_  = \new_[4798]_  & \new_[4793]_ ;
  assign \new_[4803]_  = A265 & A233;
  assign \new_[4804]_  = ~A232 & \new_[4803]_ ;
  assign \new_[4808]_  = A269 & A267;
  assign \new_[4809]_  = ~A266 & \new_[4808]_ ;
  assign \new_[4810]_  = \new_[4809]_  & \new_[4804]_ ;
  assign \new_[4814]_  = A167 & A169;
  assign \new_[4815]_  = ~A170 & \new_[4814]_ ;
  assign \new_[4819]_  = ~A201 & A199;
  assign \new_[4820]_  = A166 & \new_[4819]_ ;
  assign \new_[4821]_  = \new_[4820]_  & \new_[4815]_ ;
  assign \new_[4825]_  = A234 & ~A233;
  assign \new_[4826]_  = A232 & \new_[4825]_ ;
  assign \new_[4830]_  = A299 & ~A298;
  assign \new_[4831]_  = A235 & \new_[4830]_ ;
  assign \new_[4832]_  = \new_[4831]_  & \new_[4826]_ ;
  assign \new_[4836]_  = A167 & A169;
  assign \new_[4837]_  = ~A170 & \new_[4836]_ ;
  assign \new_[4841]_  = ~A201 & A199;
  assign \new_[4842]_  = A166 & \new_[4841]_ ;
  assign \new_[4843]_  = \new_[4842]_  & \new_[4837]_ ;
  assign \new_[4847]_  = A234 & ~A233;
  assign \new_[4848]_  = A232 & \new_[4847]_ ;
  assign \new_[4852]_  = A266 & ~A265;
  assign \new_[4853]_  = A235 & \new_[4852]_ ;
  assign \new_[4854]_  = \new_[4853]_  & \new_[4848]_ ;
  assign \new_[4858]_  = A167 & A169;
  assign \new_[4859]_  = ~A170 & \new_[4858]_ ;
  assign \new_[4863]_  = ~A201 & A199;
  assign \new_[4864]_  = A166 & \new_[4863]_ ;
  assign \new_[4865]_  = \new_[4864]_  & \new_[4859]_ ;
  assign \new_[4869]_  = A234 & ~A233;
  assign \new_[4870]_  = A232 & \new_[4869]_ ;
  assign \new_[4874]_  = A299 & ~A298;
  assign \new_[4875]_  = A236 & \new_[4874]_ ;
  assign \new_[4876]_  = \new_[4875]_  & \new_[4870]_ ;
  assign \new_[4880]_  = A167 & A169;
  assign \new_[4881]_  = ~A170 & \new_[4880]_ ;
  assign \new_[4885]_  = ~A201 & A199;
  assign \new_[4886]_  = A166 & \new_[4885]_ ;
  assign \new_[4887]_  = \new_[4886]_  & \new_[4881]_ ;
  assign \new_[4891]_  = A234 & ~A233;
  assign \new_[4892]_  = A232 & \new_[4891]_ ;
  assign \new_[4896]_  = A266 & ~A265;
  assign \new_[4897]_  = A236 & \new_[4896]_ ;
  assign \new_[4898]_  = \new_[4897]_  & \new_[4892]_ ;
  assign \new_[4902]_  = A167 & A169;
  assign \new_[4903]_  = ~A170 & \new_[4902]_ ;
  assign \new_[4907]_  = A200 & A199;
  assign \new_[4908]_  = A166 & \new_[4907]_ ;
  assign \new_[4909]_  = \new_[4908]_  & \new_[4903]_ ;
  assign \new_[4913]_  = A298 & A233;
  assign \new_[4914]_  = ~A232 & \new_[4913]_ ;
  assign \new_[4918]_  = A301 & A300;
  assign \new_[4919]_  = ~A299 & \new_[4918]_ ;
  assign \new_[4920]_  = \new_[4919]_  & \new_[4914]_ ;
  assign \new_[4924]_  = A167 & A169;
  assign \new_[4925]_  = ~A170 & \new_[4924]_ ;
  assign \new_[4929]_  = A200 & A199;
  assign \new_[4930]_  = A166 & \new_[4929]_ ;
  assign \new_[4931]_  = \new_[4930]_  & \new_[4925]_ ;
  assign \new_[4935]_  = A298 & A233;
  assign \new_[4936]_  = ~A232 & \new_[4935]_ ;
  assign \new_[4940]_  = A302 & A300;
  assign \new_[4941]_  = ~A299 & \new_[4940]_ ;
  assign \new_[4942]_  = \new_[4941]_  & \new_[4936]_ ;
  assign \new_[4946]_  = A167 & A169;
  assign \new_[4947]_  = ~A170 & \new_[4946]_ ;
  assign \new_[4951]_  = A200 & A199;
  assign \new_[4952]_  = A166 & \new_[4951]_ ;
  assign \new_[4953]_  = \new_[4952]_  & \new_[4947]_ ;
  assign \new_[4957]_  = A265 & A233;
  assign \new_[4958]_  = ~A232 & \new_[4957]_ ;
  assign \new_[4962]_  = A268 & A267;
  assign \new_[4963]_  = ~A266 & \new_[4962]_ ;
  assign \new_[4964]_  = \new_[4963]_  & \new_[4958]_ ;
  assign \new_[4968]_  = A167 & A169;
  assign \new_[4969]_  = ~A170 & \new_[4968]_ ;
  assign \new_[4973]_  = A200 & A199;
  assign \new_[4974]_  = A166 & \new_[4973]_ ;
  assign \new_[4975]_  = \new_[4974]_  & \new_[4969]_ ;
  assign \new_[4979]_  = A265 & A233;
  assign \new_[4980]_  = ~A232 & \new_[4979]_ ;
  assign \new_[4984]_  = A269 & A267;
  assign \new_[4985]_  = ~A266 & \new_[4984]_ ;
  assign \new_[4986]_  = \new_[4985]_  & \new_[4980]_ ;
  assign \new_[4990]_  = A167 & A169;
  assign \new_[4991]_  = ~A170 & \new_[4990]_ ;
  assign \new_[4995]_  = A200 & A199;
  assign \new_[4996]_  = A166 & \new_[4995]_ ;
  assign \new_[4997]_  = \new_[4996]_  & \new_[4991]_ ;
  assign \new_[5001]_  = A234 & ~A233;
  assign \new_[5002]_  = A232 & \new_[5001]_ ;
  assign \new_[5006]_  = A299 & ~A298;
  assign \new_[5007]_  = A235 & \new_[5006]_ ;
  assign \new_[5008]_  = \new_[5007]_  & \new_[5002]_ ;
  assign \new_[5012]_  = A167 & A169;
  assign \new_[5013]_  = ~A170 & \new_[5012]_ ;
  assign \new_[5017]_  = A200 & A199;
  assign \new_[5018]_  = A166 & \new_[5017]_ ;
  assign \new_[5019]_  = \new_[5018]_  & \new_[5013]_ ;
  assign \new_[5023]_  = A234 & ~A233;
  assign \new_[5024]_  = A232 & \new_[5023]_ ;
  assign \new_[5028]_  = A266 & ~A265;
  assign \new_[5029]_  = A235 & \new_[5028]_ ;
  assign \new_[5030]_  = \new_[5029]_  & \new_[5024]_ ;
  assign \new_[5034]_  = A167 & A169;
  assign \new_[5035]_  = ~A170 & \new_[5034]_ ;
  assign \new_[5039]_  = A200 & A199;
  assign \new_[5040]_  = A166 & \new_[5039]_ ;
  assign \new_[5041]_  = \new_[5040]_  & \new_[5035]_ ;
  assign \new_[5045]_  = A234 & ~A233;
  assign \new_[5046]_  = A232 & \new_[5045]_ ;
  assign \new_[5050]_  = A299 & ~A298;
  assign \new_[5051]_  = A236 & \new_[5050]_ ;
  assign \new_[5052]_  = \new_[5051]_  & \new_[5046]_ ;
  assign \new_[5056]_  = A167 & A169;
  assign \new_[5057]_  = ~A170 & \new_[5056]_ ;
  assign \new_[5061]_  = A200 & A199;
  assign \new_[5062]_  = A166 & \new_[5061]_ ;
  assign \new_[5063]_  = \new_[5062]_  & \new_[5057]_ ;
  assign \new_[5067]_  = A234 & ~A233;
  assign \new_[5068]_  = A232 & \new_[5067]_ ;
  assign \new_[5072]_  = A266 & ~A265;
  assign \new_[5073]_  = A236 & \new_[5072]_ ;
  assign \new_[5074]_  = \new_[5073]_  & \new_[5068]_ ;
  assign \new_[5078]_  = A167 & A169;
  assign \new_[5079]_  = ~A170 & \new_[5078]_ ;
  assign \new_[5083]_  = ~A200 & ~A199;
  assign \new_[5084]_  = A166 & \new_[5083]_ ;
  assign \new_[5085]_  = \new_[5084]_  & \new_[5079]_ ;
  assign \new_[5089]_  = A298 & A233;
  assign \new_[5090]_  = ~A232 & \new_[5089]_ ;
  assign \new_[5094]_  = A301 & A300;
  assign \new_[5095]_  = ~A299 & \new_[5094]_ ;
  assign \new_[5096]_  = \new_[5095]_  & \new_[5090]_ ;
  assign \new_[5100]_  = A167 & A169;
  assign \new_[5101]_  = ~A170 & \new_[5100]_ ;
  assign \new_[5105]_  = ~A200 & ~A199;
  assign \new_[5106]_  = A166 & \new_[5105]_ ;
  assign \new_[5107]_  = \new_[5106]_  & \new_[5101]_ ;
  assign \new_[5111]_  = A298 & A233;
  assign \new_[5112]_  = ~A232 & \new_[5111]_ ;
  assign \new_[5116]_  = A302 & A300;
  assign \new_[5117]_  = ~A299 & \new_[5116]_ ;
  assign \new_[5118]_  = \new_[5117]_  & \new_[5112]_ ;
  assign \new_[5122]_  = A167 & A169;
  assign \new_[5123]_  = ~A170 & \new_[5122]_ ;
  assign \new_[5127]_  = ~A200 & ~A199;
  assign \new_[5128]_  = A166 & \new_[5127]_ ;
  assign \new_[5129]_  = \new_[5128]_  & \new_[5123]_ ;
  assign \new_[5133]_  = A265 & A233;
  assign \new_[5134]_  = ~A232 & \new_[5133]_ ;
  assign \new_[5138]_  = A268 & A267;
  assign \new_[5139]_  = ~A266 & \new_[5138]_ ;
  assign \new_[5140]_  = \new_[5139]_  & \new_[5134]_ ;
  assign \new_[5144]_  = A167 & A169;
  assign \new_[5145]_  = ~A170 & \new_[5144]_ ;
  assign \new_[5149]_  = ~A200 & ~A199;
  assign \new_[5150]_  = A166 & \new_[5149]_ ;
  assign \new_[5151]_  = \new_[5150]_  & \new_[5145]_ ;
  assign \new_[5155]_  = A265 & A233;
  assign \new_[5156]_  = ~A232 & \new_[5155]_ ;
  assign \new_[5160]_  = A269 & A267;
  assign \new_[5161]_  = ~A266 & \new_[5160]_ ;
  assign \new_[5162]_  = \new_[5161]_  & \new_[5156]_ ;
  assign \new_[5166]_  = A167 & A169;
  assign \new_[5167]_  = ~A170 & \new_[5166]_ ;
  assign \new_[5171]_  = ~A200 & ~A199;
  assign \new_[5172]_  = A166 & \new_[5171]_ ;
  assign \new_[5173]_  = \new_[5172]_  & \new_[5167]_ ;
  assign \new_[5177]_  = A234 & ~A233;
  assign \new_[5178]_  = A232 & \new_[5177]_ ;
  assign \new_[5182]_  = A299 & ~A298;
  assign \new_[5183]_  = A235 & \new_[5182]_ ;
  assign \new_[5184]_  = \new_[5183]_  & \new_[5178]_ ;
  assign \new_[5188]_  = A167 & A169;
  assign \new_[5189]_  = ~A170 & \new_[5188]_ ;
  assign \new_[5193]_  = ~A200 & ~A199;
  assign \new_[5194]_  = A166 & \new_[5193]_ ;
  assign \new_[5195]_  = \new_[5194]_  & \new_[5189]_ ;
  assign \new_[5199]_  = A234 & ~A233;
  assign \new_[5200]_  = A232 & \new_[5199]_ ;
  assign \new_[5204]_  = A266 & ~A265;
  assign \new_[5205]_  = A235 & \new_[5204]_ ;
  assign \new_[5206]_  = \new_[5205]_  & \new_[5200]_ ;
  assign \new_[5210]_  = A167 & A169;
  assign \new_[5211]_  = ~A170 & \new_[5210]_ ;
  assign \new_[5215]_  = ~A200 & ~A199;
  assign \new_[5216]_  = A166 & \new_[5215]_ ;
  assign \new_[5217]_  = \new_[5216]_  & \new_[5211]_ ;
  assign \new_[5221]_  = A234 & ~A233;
  assign \new_[5222]_  = A232 & \new_[5221]_ ;
  assign \new_[5226]_  = A299 & ~A298;
  assign \new_[5227]_  = A236 & \new_[5226]_ ;
  assign \new_[5228]_  = \new_[5227]_  & \new_[5222]_ ;
  assign \new_[5232]_  = A167 & A169;
  assign \new_[5233]_  = ~A170 & \new_[5232]_ ;
  assign \new_[5237]_  = ~A200 & ~A199;
  assign \new_[5238]_  = A166 & \new_[5237]_ ;
  assign \new_[5239]_  = \new_[5238]_  & \new_[5233]_ ;
  assign \new_[5243]_  = A234 & ~A233;
  assign \new_[5244]_  = A232 & \new_[5243]_ ;
  assign \new_[5248]_  = A266 & ~A265;
  assign \new_[5249]_  = A236 & \new_[5248]_ ;
  assign \new_[5250]_  = \new_[5249]_  & \new_[5244]_ ;
  assign \new_[5254]_  = ~A167 & A169;
  assign \new_[5255]_  = ~A170 & \new_[5254]_ ;
  assign \new_[5259]_  = ~A201 & A199;
  assign \new_[5260]_  = ~A166 & \new_[5259]_ ;
  assign \new_[5261]_  = \new_[5260]_  & \new_[5255]_ ;
  assign \new_[5265]_  = A298 & A233;
  assign \new_[5266]_  = ~A232 & \new_[5265]_ ;
  assign \new_[5270]_  = A301 & A300;
  assign \new_[5271]_  = ~A299 & \new_[5270]_ ;
  assign \new_[5272]_  = \new_[5271]_  & \new_[5266]_ ;
  assign \new_[5276]_  = ~A167 & A169;
  assign \new_[5277]_  = ~A170 & \new_[5276]_ ;
  assign \new_[5281]_  = ~A201 & A199;
  assign \new_[5282]_  = ~A166 & \new_[5281]_ ;
  assign \new_[5283]_  = \new_[5282]_  & \new_[5277]_ ;
  assign \new_[5287]_  = A298 & A233;
  assign \new_[5288]_  = ~A232 & \new_[5287]_ ;
  assign \new_[5292]_  = A302 & A300;
  assign \new_[5293]_  = ~A299 & \new_[5292]_ ;
  assign \new_[5294]_  = \new_[5293]_  & \new_[5288]_ ;
  assign \new_[5298]_  = ~A167 & A169;
  assign \new_[5299]_  = ~A170 & \new_[5298]_ ;
  assign \new_[5303]_  = ~A201 & A199;
  assign \new_[5304]_  = ~A166 & \new_[5303]_ ;
  assign \new_[5305]_  = \new_[5304]_  & \new_[5299]_ ;
  assign \new_[5309]_  = A265 & A233;
  assign \new_[5310]_  = ~A232 & \new_[5309]_ ;
  assign \new_[5314]_  = A268 & A267;
  assign \new_[5315]_  = ~A266 & \new_[5314]_ ;
  assign \new_[5316]_  = \new_[5315]_  & \new_[5310]_ ;
  assign \new_[5320]_  = ~A167 & A169;
  assign \new_[5321]_  = ~A170 & \new_[5320]_ ;
  assign \new_[5325]_  = ~A201 & A199;
  assign \new_[5326]_  = ~A166 & \new_[5325]_ ;
  assign \new_[5327]_  = \new_[5326]_  & \new_[5321]_ ;
  assign \new_[5331]_  = A265 & A233;
  assign \new_[5332]_  = ~A232 & \new_[5331]_ ;
  assign \new_[5336]_  = A269 & A267;
  assign \new_[5337]_  = ~A266 & \new_[5336]_ ;
  assign \new_[5338]_  = \new_[5337]_  & \new_[5332]_ ;
  assign \new_[5342]_  = ~A167 & A169;
  assign \new_[5343]_  = ~A170 & \new_[5342]_ ;
  assign \new_[5347]_  = ~A201 & A199;
  assign \new_[5348]_  = ~A166 & \new_[5347]_ ;
  assign \new_[5349]_  = \new_[5348]_  & \new_[5343]_ ;
  assign \new_[5353]_  = A234 & ~A233;
  assign \new_[5354]_  = A232 & \new_[5353]_ ;
  assign \new_[5358]_  = A299 & ~A298;
  assign \new_[5359]_  = A235 & \new_[5358]_ ;
  assign \new_[5360]_  = \new_[5359]_  & \new_[5354]_ ;
  assign \new_[5364]_  = ~A167 & A169;
  assign \new_[5365]_  = ~A170 & \new_[5364]_ ;
  assign \new_[5369]_  = ~A201 & A199;
  assign \new_[5370]_  = ~A166 & \new_[5369]_ ;
  assign \new_[5371]_  = \new_[5370]_  & \new_[5365]_ ;
  assign \new_[5375]_  = A234 & ~A233;
  assign \new_[5376]_  = A232 & \new_[5375]_ ;
  assign \new_[5380]_  = A266 & ~A265;
  assign \new_[5381]_  = A235 & \new_[5380]_ ;
  assign \new_[5382]_  = \new_[5381]_  & \new_[5376]_ ;
  assign \new_[5386]_  = ~A167 & A169;
  assign \new_[5387]_  = ~A170 & \new_[5386]_ ;
  assign \new_[5391]_  = ~A201 & A199;
  assign \new_[5392]_  = ~A166 & \new_[5391]_ ;
  assign \new_[5393]_  = \new_[5392]_  & \new_[5387]_ ;
  assign \new_[5397]_  = A234 & ~A233;
  assign \new_[5398]_  = A232 & \new_[5397]_ ;
  assign \new_[5402]_  = A299 & ~A298;
  assign \new_[5403]_  = A236 & \new_[5402]_ ;
  assign \new_[5404]_  = \new_[5403]_  & \new_[5398]_ ;
  assign \new_[5408]_  = ~A167 & A169;
  assign \new_[5409]_  = ~A170 & \new_[5408]_ ;
  assign \new_[5413]_  = ~A201 & A199;
  assign \new_[5414]_  = ~A166 & \new_[5413]_ ;
  assign \new_[5415]_  = \new_[5414]_  & \new_[5409]_ ;
  assign \new_[5419]_  = A234 & ~A233;
  assign \new_[5420]_  = A232 & \new_[5419]_ ;
  assign \new_[5424]_  = A266 & ~A265;
  assign \new_[5425]_  = A236 & \new_[5424]_ ;
  assign \new_[5426]_  = \new_[5425]_  & \new_[5420]_ ;
  assign \new_[5430]_  = ~A167 & A169;
  assign \new_[5431]_  = ~A170 & \new_[5430]_ ;
  assign \new_[5435]_  = A200 & A199;
  assign \new_[5436]_  = ~A166 & \new_[5435]_ ;
  assign \new_[5437]_  = \new_[5436]_  & \new_[5431]_ ;
  assign \new_[5441]_  = A298 & A233;
  assign \new_[5442]_  = ~A232 & \new_[5441]_ ;
  assign \new_[5446]_  = A301 & A300;
  assign \new_[5447]_  = ~A299 & \new_[5446]_ ;
  assign \new_[5448]_  = \new_[5447]_  & \new_[5442]_ ;
  assign \new_[5452]_  = ~A167 & A169;
  assign \new_[5453]_  = ~A170 & \new_[5452]_ ;
  assign \new_[5457]_  = A200 & A199;
  assign \new_[5458]_  = ~A166 & \new_[5457]_ ;
  assign \new_[5459]_  = \new_[5458]_  & \new_[5453]_ ;
  assign \new_[5463]_  = A298 & A233;
  assign \new_[5464]_  = ~A232 & \new_[5463]_ ;
  assign \new_[5468]_  = A302 & A300;
  assign \new_[5469]_  = ~A299 & \new_[5468]_ ;
  assign \new_[5470]_  = \new_[5469]_  & \new_[5464]_ ;
  assign \new_[5474]_  = ~A167 & A169;
  assign \new_[5475]_  = ~A170 & \new_[5474]_ ;
  assign \new_[5479]_  = A200 & A199;
  assign \new_[5480]_  = ~A166 & \new_[5479]_ ;
  assign \new_[5481]_  = \new_[5480]_  & \new_[5475]_ ;
  assign \new_[5485]_  = A265 & A233;
  assign \new_[5486]_  = ~A232 & \new_[5485]_ ;
  assign \new_[5490]_  = A268 & A267;
  assign \new_[5491]_  = ~A266 & \new_[5490]_ ;
  assign \new_[5492]_  = \new_[5491]_  & \new_[5486]_ ;
  assign \new_[5496]_  = ~A167 & A169;
  assign \new_[5497]_  = ~A170 & \new_[5496]_ ;
  assign \new_[5501]_  = A200 & A199;
  assign \new_[5502]_  = ~A166 & \new_[5501]_ ;
  assign \new_[5503]_  = \new_[5502]_  & \new_[5497]_ ;
  assign \new_[5507]_  = A265 & A233;
  assign \new_[5508]_  = ~A232 & \new_[5507]_ ;
  assign \new_[5512]_  = A269 & A267;
  assign \new_[5513]_  = ~A266 & \new_[5512]_ ;
  assign \new_[5514]_  = \new_[5513]_  & \new_[5508]_ ;
  assign \new_[5518]_  = ~A167 & A169;
  assign \new_[5519]_  = ~A170 & \new_[5518]_ ;
  assign \new_[5523]_  = A200 & A199;
  assign \new_[5524]_  = ~A166 & \new_[5523]_ ;
  assign \new_[5525]_  = \new_[5524]_  & \new_[5519]_ ;
  assign \new_[5529]_  = A234 & ~A233;
  assign \new_[5530]_  = A232 & \new_[5529]_ ;
  assign \new_[5534]_  = A299 & ~A298;
  assign \new_[5535]_  = A235 & \new_[5534]_ ;
  assign \new_[5536]_  = \new_[5535]_  & \new_[5530]_ ;
  assign \new_[5540]_  = ~A167 & A169;
  assign \new_[5541]_  = ~A170 & \new_[5540]_ ;
  assign \new_[5545]_  = A200 & A199;
  assign \new_[5546]_  = ~A166 & \new_[5545]_ ;
  assign \new_[5547]_  = \new_[5546]_  & \new_[5541]_ ;
  assign \new_[5551]_  = A234 & ~A233;
  assign \new_[5552]_  = A232 & \new_[5551]_ ;
  assign \new_[5556]_  = A266 & ~A265;
  assign \new_[5557]_  = A235 & \new_[5556]_ ;
  assign \new_[5558]_  = \new_[5557]_  & \new_[5552]_ ;
  assign \new_[5562]_  = ~A167 & A169;
  assign \new_[5563]_  = ~A170 & \new_[5562]_ ;
  assign \new_[5567]_  = A200 & A199;
  assign \new_[5568]_  = ~A166 & \new_[5567]_ ;
  assign \new_[5569]_  = \new_[5568]_  & \new_[5563]_ ;
  assign \new_[5573]_  = A234 & ~A233;
  assign \new_[5574]_  = A232 & \new_[5573]_ ;
  assign \new_[5578]_  = A299 & ~A298;
  assign \new_[5579]_  = A236 & \new_[5578]_ ;
  assign \new_[5580]_  = \new_[5579]_  & \new_[5574]_ ;
  assign \new_[5584]_  = ~A167 & A169;
  assign \new_[5585]_  = ~A170 & \new_[5584]_ ;
  assign \new_[5589]_  = A200 & A199;
  assign \new_[5590]_  = ~A166 & \new_[5589]_ ;
  assign \new_[5591]_  = \new_[5590]_  & \new_[5585]_ ;
  assign \new_[5595]_  = A234 & ~A233;
  assign \new_[5596]_  = A232 & \new_[5595]_ ;
  assign \new_[5600]_  = A266 & ~A265;
  assign \new_[5601]_  = A236 & \new_[5600]_ ;
  assign \new_[5602]_  = \new_[5601]_  & \new_[5596]_ ;
  assign \new_[5606]_  = ~A167 & A169;
  assign \new_[5607]_  = ~A170 & \new_[5606]_ ;
  assign \new_[5611]_  = ~A200 & ~A199;
  assign \new_[5612]_  = ~A166 & \new_[5611]_ ;
  assign \new_[5613]_  = \new_[5612]_  & \new_[5607]_ ;
  assign \new_[5617]_  = A298 & A233;
  assign \new_[5618]_  = ~A232 & \new_[5617]_ ;
  assign \new_[5622]_  = A301 & A300;
  assign \new_[5623]_  = ~A299 & \new_[5622]_ ;
  assign \new_[5624]_  = \new_[5623]_  & \new_[5618]_ ;
  assign \new_[5628]_  = ~A167 & A169;
  assign \new_[5629]_  = ~A170 & \new_[5628]_ ;
  assign \new_[5633]_  = ~A200 & ~A199;
  assign \new_[5634]_  = ~A166 & \new_[5633]_ ;
  assign \new_[5635]_  = \new_[5634]_  & \new_[5629]_ ;
  assign \new_[5639]_  = A298 & A233;
  assign \new_[5640]_  = ~A232 & \new_[5639]_ ;
  assign \new_[5644]_  = A302 & A300;
  assign \new_[5645]_  = ~A299 & \new_[5644]_ ;
  assign \new_[5646]_  = \new_[5645]_  & \new_[5640]_ ;
  assign \new_[5650]_  = ~A167 & A169;
  assign \new_[5651]_  = ~A170 & \new_[5650]_ ;
  assign \new_[5655]_  = ~A200 & ~A199;
  assign \new_[5656]_  = ~A166 & \new_[5655]_ ;
  assign \new_[5657]_  = \new_[5656]_  & \new_[5651]_ ;
  assign \new_[5661]_  = A265 & A233;
  assign \new_[5662]_  = ~A232 & \new_[5661]_ ;
  assign \new_[5666]_  = A268 & A267;
  assign \new_[5667]_  = ~A266 & \new_[5666]_ ;
  assign \new_[5668]_  = \new_[5667]_  & \new_[5662]_ ;
  assign \new_[5672]_  = ~A167 & A169;
  assign \new_[5673]_  = ~A170 & \new_[5672]_ ;
  assign \new_[5677]_  = ~A200 & ~A199;
  assign \new_[5678]_  = ~A166 & \new_[5677]_ ;
  assign \new_[5679]_  = \new_[5678]_  & \new_[5673]_ ;
  assign \new_[5683]_  = A265 & A233;
  assign \new_[5684]_  = ~A232 & \new_[5683]_ ;
  assign \new_[5688]_  = A269 & A267;
  assign \new_[5689]_  = ~A266 & \new_[5688]_ ;
  assign \new_[5690]_  = \new_[5689]_  & \new_[5684]_ ;
  assign \new_[5694]_  = ~A167 & A169;
  assign \new_[5695]_  = ~A170 & \new_[5694]_ ;
  assign \new_[5699]_  = ~A200 & ~A199;
  assign \new_[5700]_  = ~A166 & \new_[5699]_ ;
  assign \new_[5701]_  = \new_[5700]_  & \new_[5695]_ ;
  assign \new_[5705]_  = A234 & ~A233;
  assign \new_[5706]_  = A232 & \new_[5705]_ ;
  assign \new_[5710]_  = A299 & ~A298;
  assign \new_[5711]_  = A235 & \new_[5710]_ ;
  assign \new_[5712]_  = \new_[5711]_  & \new_[5706]_ ;
  assign \new_[5716]_  = ~A167 & A169;
  assign \new_[5717]_  = ~A170 & \new_[5716]_ ;
  assign \new_[5721]_  = ~A200 & ~A199;
  assign \new_[5722]_  = ~A166 & \new_[5721]_ ;
  assign \new_[5723]_  = \new_[5722]_  & \new_[5717]_ ;
  assign \new_[5727]_  = A234 & ~A233;
  assign \new_[5728]_  = A232 & \new_[5727]_ ;
  assign \new_[5732]_  = A266 & ~A265;
  assign \new_[5733]_  = A235 & \new_[5732]_ ;
  assign \new_[5734]_  = \new_[5733]_  & \new_[5728]_ ;
  assign \new_[5738]_  = ~A167 & A169;
  assign \new_[5739]_  = ~A170 & \new_[5738]_ ;
  assign \new_[5743]_  = ~A200 & ~A199;
  assign \new_[5744]_  = ~A166 & \new_[5743]_ ;
  assign \new_[5745]_  = \new_[5744]_  & \new_[5739]_ ;
  assign \new_[5749]_  = A234 & ~A233;
  assign \new_[5750]_  = A232 & \new_[5749]_ ;
  assign \new_[5754]_  = A299 & ~A298;
  assign \new_[5755]_  = A236 & \new_[5754]_ ;
  assign \new_[5756]_  = \new_[5755]_  & \new_[5750]_ ;
  assign \new_[5760]_  = ~A167 & A169;
  assign \new_[5761]_  = ~A170 & \new_[5760]_ ;
  assign \new_[5765]_  = ~A200 & ~A199;
  assign \new_[5766]_  = ~A166 & \new_[5765]_ ;
  assign \new_[5767]_  = \new_[5766]_  & \new_[5761]_ ;
  assign \new_[5771]_  = A234 & ~A233;
  assign \new_[5772]_  = A232 & \new_[5771]_ ;
  assign \new_[5776]_  = A266 & ~A265;
  assign \new_[5777]_  = A236 & \new_[5776]_ ;
  assign \new_[5778]_  = \new_[5777]_  & \new_[5772]_ ;
  assign \new_[5782]_  = A167 & ~A169;
  assign \new_[5783]_  = A170 & \new_[5782]_ ;
  assign \new_[5787]_  = ~A201 & A199;
  assign \new_[5788]_  = ~A166 & \new_[5787]_ ;
  assign \new_[5789]_  = \new_[5788]_  & \new_[5783]_ ;
  assign \new_[5793]_  = A298 & A233;
  assign \new_[5794]_  = ~A232 & \new_[5793]_ ;
  assign \new_[5798]_  = A301 & A300;
  assign \new_[5799]_  = ~A299 & \new_[5798]_ ;
  assign \new_[5800]_  = \new_[5799]_  & \new_[5794]_ ;
  assign \new_[5804]_  = A167 & ~A169;
  assign \new_[5805]_  = A170 & \new_[5804]_ ;
  assign \new_[5809]_  = ~A201 & A199;
  assign \new_[5810]_  = ~A166 & \new_[5809]_ ;
  assign \new_[5811]_  = \new_[5810]_  & \new_[5805]_ ;
  assign \new_[5815]_  = A298 & A233;
  assign \new_[5816]_  = ~A232 & \new_[5815]_ ;
  assign \new_[5820]_  = A302 & A300;
  assign \new_[5821]_  = ~A299 & \new_[5820]_ ;
  assign \new_[5822]_  = \new_[5821]_  & \new_[5816]_ ;
  assign \new_[5826]_  = A167 & ~A169;
  assign \new_[5827]_  = A170 & \new_[5826]_ ;
  assign \new_[5831]_  = ~A201 & A199;
  assign \new_[5832]_  = ~A166 & \new_[5831]_ ;
  assign \new_[5833]_  = \new_[5832]_  & \new_[5827]_ ;
  assign \new_[5837]_  = A265 & A233;
  assign \new_[5838]_  = ~A232 & \new_[5837]_ ;
  assign \new_[5842]_  = A268 & A267;
  assign \new_[5843]_  = ~A266 & \new_[5842]_ ;
  assign \new_[5844]_  = \new_[5843]_  & \new_[5838]_ ;
  assign \new_[5848]_  = A167 & ~A169;
  assign \new_[5849]_  = A170 & \new_[5848]_ ;
  assign \new_[5853]_  = ~A201 & A199;
  assign \new_[5854]_  = ~A166 & \new_[5853]_ ;
  assign \new_[5855]_  = \new_[5854]_  & \new_[5849]_ ;
  assign \new_[5859]_  = A265 & A233;
  assign \new_[5860]_  = ~A232 & \new_[5859]_ ;
  assign \new_[5864]_  = A269 & A267;
  assign \new_[5865]_  = ~A266 & \new_[5864]_ ;
  assign \new_[5866]_  = \new_[5865]_  & \new_[5860]_ ;
  assign \new_[5870]_  = A167 & ~A169;
  assign \new_[5871]_  = A170 & \new_[5870]_ ;
  assign \new_[5875]_  = ~A201 & A199;
  assign \new_[5876]_  = ~A166 & \new_[5875]_ ;
  assign \new_[5877]_  = \new_[5876]_  & \new_[5871]_ ;
  assign \new_[5881]_  = A234 & ~A233;
  assign \new_[5882]_  = A232 & \new_[5881]_ ;
  assign \new_[5886]_  = A299 & ~A298;
  assign \new_[5887]_  = A235 & \new_[5886]_ ;
  assign \new_[5888]_  = \new_[5887]_  & \new_[5882]_ ;
  assign \new_[5892]_  = A167 & ~A169;
  assign \new_[5893]_  = A170 & \new_[5892]_ ;
  assign \new_[5897]_  = ~A201 & A199;
  assign \new_[5898]_  = ~A166 & \new_[5897]_ ;
  assign \new_[5899]_  = \new_[5898]_  & \new_[5893]_ ;
  assign \new_[5903]_  = A234 & ~A233;
  assign \new_[5904]_  = A232 & \new_[5903]_ ;
  assign \new_[5908]_  = A266 & ~A265;
  assign \new_[5909]_  = A235 & \new_[5908]_ ;
  assign \new_[5910]_  = \new_[5909]_  & \new_[5904]_ ;
  assign \new_[5914]_  = A167 & ~A169;
  assign \new_[5915]_  = A170 & \new_[5914]_ ;
  assign \new_[5919]_  = ~A201 & A199;
  assign \new_[5920]_  = ~A166 & \new_[5919]_ ;
  assign \new_[5921]_  = \new_[5920]_  & \new_[5915]_ ;
  assign \new_[5925]_  = A234 & ~A233;
  assign \new_[5926]_  = A232 & \new_[5925]_ ;
  assign \new_[5930]_  = A299 & ~A298;
  assign \new_[5931]_  = A236 & \new_[5930]_ ;
  assign \new_[5932]_  = \new_[5931]_  & \new_[5926]_ ;
  assign \new_[5936]_  = A167 & ~A169;
  assign \new_[5937]_  = A170 & \new_[5936]_ ;
  assign \new_[5941]_  = ~A201 & A199;
  assign \new_[5942]_  = ~A166 & \new_[5941]_ ;
  assign \new_[5943]_  = \new_[5942]_  & \new_[5937]_ ;
  assign \new_[5947]_  = A234 & ~A233;
  assign \new_[5948]_  = A232 & \new_[5947]_ ;
  assign \new_[5952]_  = A266 & ~A265;
  assign \new_[5953]_  = A236 & \new_[5952]_ ;
  assign \new_[5954]_  = \new_[5953]_  & \new_[5948]_ ;
  assign \new_[5958]_  = A167 & ~A169;
  assign \new_[5959]_  = A170 & \new_[5958]_ ;
  assign \new_[5963]_  = A200 & A199;
  assign \new_[5964]_  = ~A166 & \new_[5963]_ ;
  assign \new_[5965]_  = \new_[5964]_  & \new_[5959]_ ;
  assign \new_[5969]_  = A298 & A233;
  assign \new_[5970]_  = ~A232 & \new_[5969]_ ;
  assign \new_[5974]_  = A301 & A300;
  assign \new_[5975]_  = ~A299 & \new_[5974]_ ;
  assign \new_[5976]_  = \new_[5975]_  & \new_[5970]_ ;
  assign \new_[5980]_  = A167 & ~A169;
  assign \new_[5981]_  = A170 & \new_[5980]_ ;
  assign \new_[5985]_  = A200 & A199;
  assign \new_[5986]_  = ~A166 & \new_[5985]_ ;
  assign \new_[5987]_  = \new_[5986]_  & \new_[5981]_ ;
  assign \new_[5991]_  = A298 & A233;
  assign \new_[5992]_  = ~A232 & \new_[5991]_ ;
  assign \new_[5996]_  = A302 & A300;
  assign \new_[5997]_  = ~A299 & \new_[5996]_ ;
  assign \new_[5998]_  = \new_[5997]_  & \new_[5992]_ ;
  assign \new_[6002]_  = A167 & ~A169;
  assign \new_[6003]_  = A170 & \new_[6002]_ ;
  assign \new_[6007]_  = A200 & A199;
  assign \new_[6008]_  = ~A166 & \new_[6007]_ ;
  assign \new_[6009]_  = \new_[6008]_  & \new_[6003]_ ;
  assign \new_[6013]_  = A265 & A233;
  assign \new_[6014]_  = ~A232 & \new_[6013]_ ;
  assign \new_[6018]_  = A268 & A267;
  assign \new_[6019]_  = ~A266 & \new_[6018]_ ;
  assign \new_[6020]_  = \new_[6019]_  & \new_[6014]_ ;
  assign \new_[6024]_  = A167 & ~A169;
  assign \new_[6025]_  = A170 & \new_[6024]_ ;
  assign \new_[6029]_  = A200 & A199;
  assign \new_[6030]_  = ~A166 & \new_[6029]_ ;
  assign \new_[6031]_  = \new_[6030]_  & \new_[6025]_ ;
  assign \new_[6035]_  = A265 & A233;
  assign \new_[6036]_  = ~A232 & \new_[6035]_ ;
  assign \new_[6040]_  = A269 & A267;
  assign \new_[6041]_  = ~A266 & \new_[6040]_ ;
  assign \new_[6042]_  = \new_[6041]_  & \new_[6036]_ ;
  assign \new_[6046]_  = A167 & ~A169;
  assign \new_[6047]_  = A170 & \new_[6046]_ ;
  assign \new_[6051]_  = A200 & A199;
  assign \new_[6052]_  = ~A166 & \new_[6051]_ ;
  assign \new_[6053]_  = \new_[6052]_  & \new_[6047]_ ;
  assign \new_[6057]_  = A234 & ~A233;
  assign \new_[6058]_  = A232 & \new_[6057]_ ;
  assign \new_[6062]_  = A299 & ~A298;
  assign \new_[6063]_  = A235 & \new_[6062]_ ;
  assign \new_[6064]_  = \new_[6063]_  & \new_[6058]_ ;
  assign \new_[6068]_  = A167 & ~A169;
  assign \new_[6069]_  = A170 & \new_[6068]_ ;
  assign \new_[6073]_  = A200 & A199;
  assign \new_[6074]_  = ~A166 & \new_[6073]_ ;
  assign \new_[6075]_  = \new_[6074]_  & \new_[6069]_ ;
  assign \new_[6079]_  = A234 & ~A233;
  assign \new_[6080]_  = A232 & \new_[6079]_ ;
  assign \new_[6084]_  = A266 & ~A265;
  assign \new_[6085]_  = A235 & \new_[6084]_ ;
  assign \new_[6086]_  = \new_[6085]_  & \new_[6080]_ ;
  assign \new_[6090]_  = A167 & ~A169;
  assign \new_[6091]_  = A170 & \new_[6090]_ ;
  assign \new_[6095]_  = A200 & A199;
  assign \new_[6096]_  = ~A166 & \new_[6095]_ ;
  assign \new_[6097]_  = \new_[6096]_  & \new_[6091]_ ;
  assign \new_[6101]_  = A234 & ~A233;
  assign \new_[6102]_  = A232 & \new_[6101]_ ;
  assign \new_[6106]_  = A299 & ~A298;
  assign \new_[6107]_  = A236 & \new_[6106]_ ;
  assign \new_[6108]_  = \new_[6107]_  & \new_[6102]_ ;
  assign \new_[6112]_  = A167 & ~A169;
  assign \new_[6113]_  = A170 & \new_[6112]_ ;
  assign \new_[6117]_  = A200 & A199;
  assign \new_[6118]_  = ~A166 & \new_[6117]_ ;
  assign \new_[6119]_  = \new_[6118]_  & \new_[6113]_ ;
  assign \new_[6123]_  = A234 & ~A233;
  assign \new_[6124]_  = A232 & \new_[6123]_ ;
  assign \new_[6128]_  = A266 & ~A265;
  assign \new_[6129]_  = A236 & \new_[6128]_ ;
  assign \new_[6130]_  = \new_[6129]_  & \new_[6124]_ ;
  assign \new_[6134]_  = A167 & ~A169;
  assign \new_[6135]_  = A170 & \new_[6134]_ ;
  assign \new_[6139]_  = ~A200 & ~A199;
  assign \new_[6140]_  = ~A166 & \new_[6139]_ ;
  assign \new_[6141]_  = \new_[6140]_  & \new_[6135]_ ;
  assign \new_[6145]_  = A298 & A233;
  assign \new_[6146]_  = ~A232 & \new_[6145]_ ;
  assign \new_[6150]_  = A301 & A300;
  assign \new_[6151]_  = ~A299 & \new_[6150]_ ;
  assign \new_[6152]_  = \new_[6151]_  & \new_[6146]_ ;
  assign \new_[6156]_  = A167 & ~A169;
  assign \new_[6157]_  = A170 & \new_[6156]_ ;
  assign \new_[6161]_  = ~A200 & ~A199;
  assign \new_[6162]_  = ~A166 & \new_[6161]_ ;
  assign \new_[6163]_  = \new_[6162]_  & \new_[6157]_ ;
  assign \new_[6167]_  = A298 & A233;
  assign \new_[6168]_  = ~A232 & \new_[6167]_ ;
  assign \new_[6172]_  = A302 & A300;
  assign \new_[6173]_  = ~A299 & \new_[6172]_ ;
  assign \new_[6174]_  = \new_[6173]_  & \new_[6168]_ ;
  assign \new_[6178]_  = A167 & ~A169;
  assign \new_[6179]_  = A170 & \new_[6178]_ ;
  assign \new_[6183]_  = ~A200 & ~A199;
  assign \new_[6184]_  = ~A166 & \new_[6183]_ ;
  assign \new_[6185]_  = \new_[6184]_  & \new_[6179]_ ;
  assign \new_[6189]_  = A265 & A233;
  assign \new_[6190]_  = ~A232 & \new_[6189]_ ;
  assign \new_[6194]_  = A268 & A267;
  assign \new_[6195]_  = ~A266 & \new_[6194]_ ;
  assign \new_[6196]_  = \new_[6195]_  & \new_[6190]_ ;
  assign \new_[6200]_  = A167 & ~A169;
  assign \new_[6201]_  = A170 & \new_[6200]_ ;
  assign \new_[6205]_  = ~A200 & ~A199;
  assign \new_[6206]_  = ~A166 & \new_[6205]_ ;
  assign \new_[6207]_  = \new_[6206]_  & \new_[6201]_ ;
  assign \new_[6211]_  = A265 & A233;
  assign \new_[6212]_  = ~A232 & \new_[6211]_ ;
  assign \new_[6216]_  = A269 & A267;
  assign \new_[6217]_  = ~A266 & \new_[6216]_ ;
  assign \new_[6218]_  = \new_[6217]_  & \new_[6212]_ ;
  assign \new_[6222]_  = A167 & ~A169;
  assign \new_[6223]_  = A170 & \new_[6222]_ ;
  assign \new_[6227]_  = ~A200 & ~A199;
  assign \new_[6228]_  = ~A166 & \new_[6227]_ ;
  assign \new_[6229]_  = \new_[6228]_  & \new_[6223]_ ;
  assign \new_[6233]_  = A234 & ~A233;
  assign \new_[6234]_  = A232 & \new_[6233]_ ;
  assign \new_[6238]_  = A299 & ~A298;
  assign \new_[6239]_  = A235 & \new_[6238]_ ;
  assign \new_[6240]_  = \new_[6239]_  & \new_[6234]_ ;
  assign \new_[6244]_  = A167 & ~A169;
  assign \new_[6245]_  = A170 & \new_[6244]_ ;
  assign \new_[6249]_  = ~A200 & ~A199;
  assign \new_[6250]_  = ~A166 & \new_[6249]_ ;
  assign \new_[6251]_  = \new_[6250]_  & \new_[6245]_ ;
  assign \new_[6255]_  = A234 & ~A233;
  assign \new_[6256]_  = A232 & \new_[6255]_ ;
  assign \new_[6260]_  = A266 & ~A265;
  assign \new_[6261]_  = A235 & \new_[6260]_ ;
  assign \new_[6262]_  = \new_[6261]_  & \new_[6256]_ ;
  assign \new_[6266]_  = A167 & ~A169;
  assign \new_[6267]_  = A170 & \new_[6266]_ ;
  assign \new_[6271]_  = ~A200 & ~A199;
  assign \new_[6272]_  = ~A166 & \new_[6271]_ ;
  assign \new_[6273]_  = \new_[6272]_  & \new_[6267]_ ;
  assign \new_[6277]_  = A234 & ~A233;
  assign \new_[6278]_  = A232 & \new_[6277]_ ;
  assign \new_[6282]_  = A299 & ~A298;
  assign \new_[6283]_  = A236 & \new_[6282]_ ;
  assign \new_[6284]_  = \new_[6283]_  & \new_[6278]_ ;
  assign \new_[6288]_  = A167 & ~A169;
  assign \new_[6289]_  = A170 & \new_[6288]_ ;
  assign \new_[6293]_  = ~A200 & ~A199;
  assign \new_[6294]_  = ~A166 & \new_[6293]_ ;
  assign \new_[6295]_  = \new_[6294]_  & \new_[6289]_ ;
  assign \new_[6299]_  = A234 & ~A233;
  assign \new_[6300]_  = A232 & \new_[6299]_ ;
  assign \new_[6304]_  = A266 & ~A265;
  assign \new_[6305]_  = A236 & \new_[6304]_ ;
  assign \new_[6306]_  = \new_[6305]_  & \new_[6300]_ ;
  assign \new_[6310]_  = ~A167 & ~A169;
  assign \new_[6311]_  = A170 & \new_[6310]_ ;
  assign \new_[6315]_  = ~A201 & A199;
  assign \new_[6316]_  = A166 & \new_[6315]_ ;
  assign \new_[6317]_  = \new_[6316]_  & \new_[6311]_ ;
  assign \new_[6321]_  = A298 & A233;
  assign \new_[6322]_  = ~A232 & \new_[6321]_ ;
  assign \new_[6326]_  = A301 & A300;
  assign \new_[6327]_  = ~A299 & \new_[6326]_ ;
  assign \new_[6328]_  = \new_[6327]_  & \new_[6322]_ ;
  assign \new_[6332]_  = ~A167 & ~A169;
  assign \new_[6333]_  = A170 & \new_[6332]_ ;
  assign \new_[6337]_  = ~A201 & A199;
  assign \new_[6338]_  = A166 & \new_[6337]_ ;
  assign \new_[6339]_  = \new_[6338]_  & \new_[6333]_ ;
  assign \new_[6343]_  = A298 & A233;
  assign \new_[6344]_  = ~A232 & \new_[6343]_ ;
  assign \new_[6348]_  = A302 & A300;
  assign \new_[6349]_  = ~A299 & \new_[6348]_ ;
  assign \new_[6350]_  = \new_[6349]_  & \new_[6344]_ ;
  assign \new_[6354]_  = ~A167 & ~A169;
  assign \new_[6355]_  = A170 & \new_[6354]_ ;
  assign \new_[6359]_  = ~A201 & A199;
  assign \new_[6360]_  = A166 & \new_[6359]_ ;
  assign \new_[6361]_  = \new_[6360]_  & \new_[6355]_ ;
  assign \new_[6365]_  = A265 & A233;
  assign \new_[6366]_  = ~A232 & \new_[6365]_ ;
  assign \new_[6370]_  = A268 & A267;
  assign \new_[6371]_  = ~A266 & \new_[6370]_ ;
  assign \new_[6372]_  = \new_[6371]_  & \new_[6366]_ ;
  assign \new_[6376]_  = ~A167 & ~A169;
  assign \new_[6377]_  = A170 & \new_[6376]_ ;
  assign \new_[6381]_  = ~A201 & A199;
  assign \new_[6382]_  = A166 & \new_[6381]_ ;
  assign \new_[6383]_  = \new_[6382]_  & \new_[6377]_ ;
  assign \new_[6387]_  = A265 & A233;
  assign \new_[6388]_  = ~A232 & \new_[6387]_ ;
  assign \new_[6392]_  = A269 & A267;
  assign \new_[6393]_  = ~A266 & \new_[6392]_ ;
  assign \new_[6394]_  = \new_[6393]_  & \new_[6388]_ ;
  assign \new_[6398]_  = ~A167 & ~A169;
  assign \new_[6399]_  = A170 & \new_[6398]_ ;
  assign \new_[6403]_  = ~A201 & A199;
  assign \new_[6404]_  = A166 & \new_[6403]_ ;
  assign \new_[6405]_  = \new_[6404]_  & \new_[6399]_ ;
  assign \new_[6409]_  = A234 & ~A233;
  assign \new_[6410]_  = A232 & \new_[6409]_ ;
  assign \new_[6414]_  = A299 & ~A298;
  assign \new_[6415]_  = A235 & \new_[6414]_ ;
  assign \new_[6416]_  = \new_[6415]_  & \new_[6410]_ ;
  assign \new_[6420]_  = ~A167 & ~A169;
  assign \new_[6421]_  = A170 & \new_[6420]_ ;
  assign \new_[6425]_  = ~A201 & A199;
  assign \new_[6426]_  = A166 & \new_[6425]_ ;
  assign \new_[6427]_  = \new_[6426]_  & \new_[6421]_ ;
  assign \new_[6431]_  = A234 & ~A233;
  assign \new_[6432]_  = A232 & \new_[6431]_ ;
  assign \new_[6436]_  = A266 & ~A265;
  assign \new_[6437]_  = A235 & \new_[6436]_ ;
  assign \new_[6438]_  = \new_[6437]_  & \new_[6432]_ ;
  assign \new_[6442]_  = ~A167 & ~A169;
  assign \new_[6443]_  = A170 & \new_[6442]_ ;
  assign \new_[6447]_  = ~A201 & A199;
  assign \new_[6448]_  = A166 & \new_[6447]_ ;
  assign \new_[6449]_  = \new_[6448]_  & \new_[6443]_ ;
  assign \new_[6453]_  = A234 & ~A233;
  assign \new_[6454]_  = A232 & \new_[6453]_ ;
  assign \new_[6458]_  = A299 & ~A298;
  assign \new_[6459]_  = A236 & \new_[6458]_ ;
  assign \new_[6460]_  = \new_[6459]_  & \new_[6454]_ ;
  assign \new_[6464]_  = ~A167 & ~A169;
  assign \new_[6465]_  = A170 & \new_[6464]_ ;
  assign \new_[6469]_  = ~A201 & A199;
  assign \new_[6470]_  = A166 & \new_[6469]_ ;
  assign \new_[6471]_  = \new_[6470]_  & \new_[6465]_ ;
  assign \new_[6475]_  = A234 & ~A233;
  assign \new_[6476]_  = A232 & \new_[6475]_ ;
  assign \new_[6480]_  = A266 & ~A265;
  assign \new_[6481]_  = A236 & \new_[6480]_ ;
  assign \new_[6482]_  = \new_[6481]_  & \new_[6476]_ ;
  assign \new_[6486]_  = ~A167 & ~A169;
  assign \new_[6487]_  = A170 & \new_[6486]_ ;
  assign \new_[6491]_  = A200 & A199;
  assign \new_[6492]_  = A166 & \new_[6491]_ ;
  assign \new_[6493]_  = \new_[6492]_  & \new_[6487]_ ;
  assign \new_[6497]_  = A298 & A233;
  assign \new_[6498]_  = ~A232 & \new_[6497]_ ;
  assign \new_[6502]_  = A301 & A300;
  assign \new_[6503]_  = ~A299 & \new_[6502]_ ;
  assign \new_[6504]_  = \new_[6503]_  & \new_[6498]_ ;
  assign \new_[6508]_  = ~A167 & ~A169;
  assign \new_[6509]_  = A170 & \new_[6508]_ ;
  assign \new_[6513]_  = A200 & A199;
  assign \new_[6514]_  = A166 & \new_[6513]_ ;
  assign \new_[6515]_  = \new_[6514]_  & \new_[6509]_ ;
  assign \new_[6519]_  = A298 & A233;
  assign \new_[6520]_  = ~A232 & \new_[6519]_ ;
  assign \new_[6524]_  = A302 & A300;
  assign \new_[6525]_  = ~A299 & \new_[6524]_ ;
  assign \new_[6526]_  = \new_[6525]_  & \new_[6520]_ ;
  assign \new_[6530]_  = ~A167 & ~A169;
  assign \new_[6531]_  = A170 & \new_[6530]_ ;
  assign \new_[6535]_  = A200 & A199;
  assign \new_[6536]_  = A166 & \new_[6535]_ ;
  assign \new_[6537]_  = \new_[6536]_  & \new_[6531]_ ;
  assign \new_[6541]_  = A265 & A233;
  assign \new_[6542]_  = ~A232 & \new_[6541]_ ;
  assign \new_[6546]_  = A268 & A267;
  assign \new_[6547]_  = ~A266 & \new_[6546]_ ;
  assign \new_[6548]_  = \new_[6547]_  & \new_[6542]_ ;
  assign \new_[6552]_  = ~A167 & ~A169;
  assign \new_[6553]_  = A170 & \new_[6552]_ ;
  assign \new_[6557]_  = A200 & A199;
  assign \new_[6558]_  = A166 & \new_[6557]_ ;
  assign \new_[6559]_  = \new_[6558]_  & \new_[6553]_ ;
  assign \new_[6563]_  = A265 & A233;
  assign \new_[6564]_  = ~A232 & \new_[6563]_ ;
  assign \new_[6568]_  = A269 & A267;
  assign \new_[6569]_  = ~A266 & \new_[6568]_ ;
  assign \new_[6570]_  = \new_[6569]_  & \new_[6564]_ ;
  assign \new_[6574]_  = ~A167 & ~A169;
  assign \new_[6575]_  = A170 & \new_[6574]_ ;
  assign \new_[6579]_  = A200 & A199;
  assign \new_[6580]_  = A166 & \new_[6579]_ ;
  assign \new_[6581]_  = \new_[6580]_  & \new_[6575]_ ;
  assign \new_[6585]_  = A234 & ~A233;
  assign \new_[6586]_  = A232 & \new_[6585]_ ;
  assign \new_[6590]_  = A299 & ~A298;
  assign \new_[6591]_  = A235 & \new_[6590]_ ;
  assign \new_[6592]_  = \new_[6591]_  & \new_[6586]_ ;
  assign \new_[6596]_  = ~A167 & ~A169;
  assign \new_[6597]_  = A170 & \new_[6596]_ ;
  assign \new_[6601]_  = A200 & A199;
  assign \new_[6602]_  = A166 & \new_[6601]_ ;
  assign \new_[6603]_  = \new_[6602]_  & \new_[6597]_ ;
  assign \new_[6607]_  = A234 & ~A233;
  assign \new_[6608]_  = A232 & \new_[6607]_ ;
  assign \new_[6612]_  = A266 & ~A265;
  assign \new_[6613]_  = A235 & \new_[6612]_ ;
  assign \new_[6614]_  = \new_[6613]_  & \new_[6608]_ ;
  assign \new_[6618]_  = ~A167 & ~A169;
  assign \new_[6619]_  = A170 & \new_[6618]_ ;
  assign \new_[6623]_  = A200 & A199;
  assign \new_[6624]_  = A166 & \new_[6623]_ ;
  assign \new_[6625]_  = \new_[6624]_  & \new_[6619]_ ;
  assign \new_[6629]_  = A234 & ~A233;
  assign \new_[6630]_  = A232 & \new_[6629]_ ;
  assign \new_[6634]_  = A299 & ~A298;
  assign \new_[6635]_  = A236 & \new_[6634]_ ;
  assign \new_[6636]_  = \new_[6635]_  & \new_[6630]_ ;
  assign \new_[6640]_  = ~A167 & ~A169;
  assign \new_[6641]_  = A170 & \new_[6640]_ ;
  assign \new_[6645]_  = A200 & A199;
  assign \new_[6646]_  = A166 & \new_[6645]_ ;
  assign \new_[6647]_  = \new_[6646]_  & \new_[6641]_ ;
  assign \new_[6651]_  = A234 & ~A233;
  assign \new_[6652]_  = A232 & \new_[6651]_ ;
  assign \new_[6656]_  = A266 & ~A265;
  assign \new_[6657]_  = A236 & \new_[6656]_ ;
  assign \new_[6658]_  = \new_[6657]_  & \new_[6652]_ ;
  assign \new_[6662]_  = ~A167 & ~A169;
  assign \new_[6663]_  = A170 & \new_[6662]_ ;
  assign \new_[6667]_  = ~A200 & ~A199;
  assign \new_[6668]_  = A166 & \new_[6667]_ ;
  assign \new_[6669]_  = \new_[6668]_  & \new_[6663]_ ;
  assign \new_[6673]_  = A298 & A233;
  assign \new_[6674]_  = ~A232 & \new_[6673]_ ;
  assign \new_[6678]_  = A301 & A300;
  assign \new_[6679]_  = ~A299 & \new_[6678]_ ;
  assign \new_[6680]_  = \new_[6679]_  & \new_[6674]_ ;
  assign \new_[6684]_  = ~A167 & ~A169;
  assign \new_[6685]_  = A170 & \new_[6684]_ ;
  assign \new_[6689]_  = ~A200 & ~A199;
  assign \new_[6690]_  = A166 & \new_[6689]_ ;
  assign \new_[6691]_  = \new_[6690]_  & \new_[6685]_ ;
  assign \new_[6695]_  = A298 & A233;
  assign \new_[6696]_  = ~A232 & \new_[6695]_ ;
  assign \new_[6700]_  = A302 & A300;
  assign \new_[6701]_  = ~A299 & \new_[6700]_ ;
  assign \new_[6702]_  = \new_[6701]_  & \new_[6696]_ ;
  assign \new_[6706]_  = ~A167 & ~A169;
  assign \new_[6707]_  = A170 & \new_[6706]_ ;
  assign \new_[6711]_  = ~A200 & ~A199;
  assign \new_[6712]_  = A166 & \new_[6711]_ ;
  assign \new_[6713]_  = \new_[6712]_  & \new_[6707]_ ;
  assign \new_[6717]_  = A265 & A233;
  assign \new_[6718]_  = ~A232 & \new_[6717]_ ;
  assign \new_[6722]_  = A268 & A267;
  assign \new_[6723]_  = ~A266 & \new_[6722]_ ;
  assign \new_[6724]_  = \new_[6723]_  & \new_[6718]_ ;
  assign \new_[6728]_  = ~A167 & ~A169;
  assign \new_[6729]_  = A170 & \new_[6728]_ ;
  assign \new_[6733]_  = ~A200 & ~A199;
  assign \new_[6734]_  = A166 & \new_[6733]_ ;
  assign \new_[6735]_  = \new_[6734]_  & \new_[6729]_ ;
  assign \new_[6739]_  = A265 & A233;
  assign \new_[6740]_  = ~A232 & \new_[6739]_ ;
  assign \new_[6744]_  = A269 & A267;
  assign \new_[6745]_  = ~A266 & \new_[6744]_ ;
  assign \new_[6746]_  = \new_[6745]_  & \new_[6740]_ ;
  assign \new_[6750]_  = ~A167 & ~A169;
  assign \new_[6751]_  = A170 & \new_[6750]_ ;
  assign \new_[6755]_  = ~A200 & ~A199;
  assign \new_[6756]_  = A166 & \new_[6755]_ ;
  assign \new_[6757]_  = \new_[6756]_  & \new_[6751]_ ;
  assign \new_[6761]_  = A234 & ~A233;
  assign \new_[6762]_  = A232 & \new_[6761]_ ;
  assign \new_[6766]_  = A299 & ~A298;
  assign \new_[6767]_  = A235 & \new_[6766]_ ;
  assign \new_[6768]_  = \new_[6767]_  & \new_[6762]_ ;
  assign \new_[6772]_  = ~A167 & ~A169;
  assign \new_[6773]_  = A170 & \new_[6772]_ ;
  assign \new_[6777]_  = ~A200 & ~A199;
  assign \new_[6778]_  = A166 & \new_[6777]_ ;
  assign \new_[6779]_  = \new_[6778]_  & \new_[6773]_ ;
  assign \new_[6783]_  = A234 & ~A233;
  assign \new_[6784]_  = A232 & \new_[6783]_ ;
  assign \new_[6788]_  = A266 & ~A265;
  assign \new_[6789]_  = A235 & \new_[6788]_ ;
  assign \new_[6790]_  = \new_[6789]_  & \new_[6784]_ ;
  assign \new_[6794]_  = ~A167 & ~A169;
  assign \new_[6795]_  = A170 & \new_[6794]_ ;
  assign \new_[6799]_  = ~A200 & ~A199;
  assign \new_[6800]_  = A166 & \new_[6799]_ ;
  assign \new_[6801]_  = \new_[6800]_  & \new_[6795]_ ;
  assign \new_[6805]_  = A234 & ~A233;
  assign \new_[6806]_  = A232 & \new_[6805]_ ;
  assign \new_[6810]_  = A299 & ~A298;
  assign \new_[6811]_  = A236 & \new_[6810]_ ;
  assign \new_[6812]_  = \new_[6811]_  & \new_[6806]_ ;
  assign \new_[6816]_  = ~A167 & ~A169;
  assign \new_[6817]_  = A170 & \new_[6816]_ ;
  assign \new_[6821]_  = ~A200 & ~A199;
  assign \new_[6822]_  = A166 & \new_[6821]_ ;
  assign \new_[6823]_  = \new_[6822]_  & \new_[6817]_ ;
  assign \new_[6827]_  = A234 & ~A233;
  assign \new_[6828]_  = A232 & \new_[6827]_ ;
  assign \new_[6832]_  = A266 & ~A265;
  assign \new_[6833]_  = A236 & \new_[6832]_ ;
  assign \new_[6834]_  = \new_[6833]_  & \new_[6828]_ ;
  assign \new_[6838]_  = A199 & A166;
  assign \new_[6839]_  = A168 & \new_[6838]_ ;
  assign \new_[6843]_  = A232 & ~A203;
  assign \new_[6844]_  = ~A202 & \new_[6843]_ ;
  assign \new_[6845]_  = \new_[6844]_  & \new_[6839]_ ;
  assign \new_[6849]_  = A235 & A234;
  assign \new_[6850]_  = ~A233 & \new_[6849]_ ;
  assign \new_[6853]_  = ~A299 & A298;
  assign \new_[6856]_  = A301 & A300;
  assign \new_[6857]_  = \new_[6856]_  & \new_[6853]_ ;
  assign \new_[6858]_  = \new_[6857]_  & \new_[6850]_ ;
  assign \new_[6862]_  = A199 & A166;
  assign \new_[6863]_  = A168 & \new_[6862]_ ;
  assign \new_[6867]_  = A232 & ~A203;
  assign \new_[6868]_  = ~A202 & \new_[6867]_ ;
  assign \new_[6869]_  = \new_[6868]_  & \new_[6863]_ ;
  assign \new_[6873]_  = A235 & A234;
  assign \new_[6874]_  = ~A233 & \new_[6873]_ ;
  assign \new_[6877]_  = ~A299 & A298;
  assign \new_[6880]_  = A302 & A300;
  assign \new_[6881]_  = \new_[6880]_  & \new_[6877]_ ;
  assign \new_[6882]_  = \new_[6881]_  & \new_[6874]_ ;
  assign \new_[6886]_  = A199 & A166;
  assign \new_[6887]_  = A168 & \new_[6886]_ ;
  assign \new_[6891]_  = A232 & ~A203;
  assign \new_[6892]_  = ~A202 & \new_[6891]_ ;
  assign \new_[6893]_  = \new_[6892]_  & \new_[6887]_ ;
  assign \new_[6897]_  = A235 & A234;
  assign \new_[6898]_  = ~A233 & \new_[6897]_ ;
  assign \new_[6901]_  = ~A266 & A265;
  assign \new_[6904]_  = A268 & A267;
  assign \new_[6905]_  = \new_[6904]_  & \new_[6901]_ ;
  assign \new_[6906]_  = \new_[6905]_  & \new_[6898]_ ;
  assign \new_[6910]_  = A199 & A166;
  assign \new_[6911]_  = A168 & \new_[6910]_ ;
  assign \new_[6915]_  = A232 & ~A203;
  assign \new_[6916]_  = ~A202 & \new_[6915]_ ;
  assign \new_[6917]_  = \new_[6916]_  & \new_[6911]_ ;
  assign \new_[6921]_  = A235 & A234;
  assign \new_[6922]_  = ~A233 & \new_[6921]_ ;
  assign \new_[6925]_  = ~A266 & A265;
  assign \new_[6928]_  = A269 & A267;
  assign \new_[6929]_  = \new_[6928]_  & \new_[6925]_ ;
  assign \new_[6930]_  = \new_[6929]_  & \new_[6922]_ ;
  assign \new_[6934]_  = A199 & A166;
  assign \new_[6935]_  = A168 & \new_[6934]_ ;
  assign \new_[6939]_  = A232 & ~A203;
  assign \new_[6940]_  = ~A202 & \new_[6939]_ ;
  assign \new_[6941]_  = \new_[6940]_  & \new_[6935]_ ;
  assign \new_[6945]_  = A236 & A234;
  assign \new_[6946]_  = ~A233 & \new_[6945]_ ;
  assign \new_[6949]_  = ~A299 & A298;
  assign \new_[6952]_  = A301 & A300;
  assign \new_[6953]_  = \new_[6952]_  & \new_[6949]_ ;
  assign \new_[6954]_  = \new_[6953]_  & \new_[6946]_ ;
  assign \new_[6958]_  = A199 & A166;
  assign \new_[6959]_  = A168 & \new_[6958]_ ;
  assign \new_[6963]_  = A232 & ~A203;
  assign \new_[6964]_  = ~A202 & \new_[6963]_ ;
  assign \new_[6965]_  = \new_[6964]_  & \new_[6959]_ ;
  assign \new_[6969]_  = A236 & A234;
  assign \new_[6970]_  = ~A233 & \new_[6969]_ ;
  assign \new_[6973]_  = ~A299 & A298;
  assign \new_[6976]_  = A302 & A300;
  assign \new_[6977]_  = \new_[6976]_  & \new_[6973]_ ;
  assign \new_[6978]_  = \new_[6977]_  & \new_[6970]_ ;
  assign \new_[6982]_  = A199 & A166;
  assign \new_[6983]_  = A168 & \new_[6982]_ ;
  assign \new_[6987]_  = A232 & ~A203;
  assign \new_[6988]_  = ~A202 & \new_[6987]_ ;
  assign \new_[6989]_  = \new_[6988]_  & \new_[6983]_ ;
  assign \new_[6993]_  = A236 & A234;
  assign \new_[6994]_  = ~A233 & \new_[6993]_ ;
  assign \new_[6997]_  = ~A266 & A265;
  assign \new_[7000]_  = A268 & A267;
  assign \new_[7001]_  = \new_[7000]_  & \new_[6997]_ ;
  assign \new_[7002]_  = \new_[7001]_  & \new_[6994]_ ;
  assign \new_[7006]_  = A199 & A166;
  assign \new_[7007]_  = A168 & \new_[7006]_ ;
  assign \new_[7011]_  = A232 & ~A203;
  assign \new_[7012]_  = ~A202 & \new_[7011]_ ;
  assign \new_[7013]_  = \new_[7012]_  & \new_[7007]_ ;
  assign \new_[7017]_  = A236 & A234;
  assign \new_[7018]_  = ~A233 & \new_[7017]_ ;
  assign \new_[7021]_  = ~A266 & A265;
  assign \new_[7024]_  = A269 & A267;
  assign \new_[7025]_  = \new_[7024]_  & \new_[7021]_ ;
  assign \new_[7026]_  = \new_[7025]_  & \new_[7018]_ ;
  assign \new_[7030]_  = A199 & A167;
  assign \new_[7031]_  = A168 & \new_[7030]_ ;
  assign \new_[7035]_  = A232 & ~A203;
  assign \new_[7036]_  = ~A202 & \new_[7035]_ ;
  assign \new_[7037]_  = \new_[7036]_  & \new_[7031]_ ;
  assign \new_[7041]_  = A235 & A234;
  assign \new_[7042]_  = ~A233 & \new_[7041]_ ;
  assign \new_[7045]_  = ~A299 & A298;
  assign \new_[7048]_  = A301 & A300;
  assign \new_[7049]_  = \new_[7048]_  & \new_[7045]_ ;
  assign \new_[7050]_  = \new_[7049]_  & \new_[7042]_ ;
  assign \new_[7054]_  = A199 & A167;
  assign \new_[7055]_  = A168 & \new_[7054]_ ;
  assign \new_[7059]_  = A232 & ~A203;
  assign \new_[7060]_  = ~A202 & \new_[7059]_ ;
  assign \new_[7061]_  = \new_[7060]_  & \new_[7055]_ ;
  assign \new_[7065]_  = A235 & A234;
  assign \new_[7066]_  = ~A233 & \new_[7065]_ ;
  assign \new_[7069]_  = ~A299 & A298;
  assign \new_[7072]_  = A302 & A300;
  assign \new_[7073]_  = \new_[7072]_  & \new_[7069]_ ;
  assign \new_[7074]_  = \new_[7073]_  & \new_[7066]_ ;
  assign \new_[7078]_  = A199 & A167;
  assign \new_[7079]_  = A168 & \new_[7078]_ ;
  assign \new_[7083]_  = A232 & ~A203;
  assign \new_[7084]_  = ~A202 & \new_[7083]_ ;
  assign \new_[7085]_  = \new_[7084]_  & \new_[7079]_ ;
  assign \new_[7089]_  = A235 & A234;
  assign \new_[7090]_  = ~A233 & \new_[7089]_ ;
  assign \new_[7093]_  = ~A266 & A265;
  assign \new_[7096]_  = A268 & A267;
  assign \new_[7097]_  = \new_[7096]_  & \new_[7093]_ ;
  assign \new_[7098]_  = \new_[7097]_  & \new_[7090]_ ;
  assign \new_[7102]_  = A199 & A167;
  assign \new_[7103]_  = A168 & \new_[7102]_ ;
  assign \new_[7107]_  = A232 & ~A203;
  assign \new_[7108]_  = ~A202 & \new_[7107]_ ;
  assign \new_[7109]_  = \new_[7108]_  & \new_[7103]_ ;
  assign \new_[7113]_  = A235 & A234;
  assign \new_[7114]_  = ~A233 & \new_[7113]_ ;
  assign \new_[7117]_  = ~A266 & A265;
  assign \new_[7120]_  = A269 & A267;
  assign \new_[7121]_  = \new_[7120]_  & \new_[7117]_ ;
  assign \new_[7122]_  = \new_[7121]_  & \new_[7114]_ ;
  assign \new_[7126]_  = A199 & A167;
  assign \new_[7127]_  = A168 & \new_[7126]_ ;
  assign \new_[7131]_  = A232 & ~A203;
  assign \new_[7132]_  = ~A202 & \new_[7131]_ ;
  assign \new_[7133]_  = \new_[7132]_  & \new_[7127]_ ;
  assign \new_[7137]_  = A236 & A234;
  assign \new_[7138]_  = ~A233 & \new_[7137]_ ;
  assign \new_[7141]_  = ~A299 & A298;
  assign \new_[7144]_  = A301 & A300;
  assign \new_[7145]_  = \new_[7144]_  & \new_[7141]_ ;
  assign \new_[7146]_  = \new_[7145]_  & \new_[7138]_ ;
  assign \new_[7150]_  = A199 & A167;
  assign \new_[7151]_  = A168 & \new_[7150]_ ;
  assign \new_[7155]_  = A232 & ~A203;
  assign \new_[7156]_  = ~A202 & \new_[7155]_ ;
  assign \new_[7157]_  = \new_[7156]_  & \new_[7151]_ ;
  assign \new_[7161]_  = A236 & A234;
  assign \new_[7162]_  = ~A233 & \new_[7161]_ ;
  assign \new_[7165]_  = ~A299 & A298;
  assign \new_[7168]_  = A302 & A300;
  assign \new_[7169]_  = \new_[7168]_  & \new_[7165]_ ;
  assign \new_[7170]_  = \new_[7169]_  & \new_[7162]_ ;
  assign \new_[7174]_  = A199 & A167;
  assign \new_[7175]_  = A168 & \new_[7174]_ ;
  assign \new_[7179]_  = A232 & ~A203;
  assign \new_[7180]_  = ~A202 & \new_[7179]_ ;
  assign \new_[7181]_  = \new_[7180]_  & \new_[7175]_ ;
  assign \new_[7185]_  = A236 & A234;
  assign \new_[7186]_  = ~A233 & \new_[7185]_ ;
  assign \new_[7189]_  = ~A266 & A265;
  assign \new_[7192]_  = A268 & A267;
  assign \new_[7193]_  = \new_[7192]_  & \new_[7189]_ ;
  assign \new_[7194]_  = \new_[7193]_  & \new_[7186]_ ;
  assign \new_[7198]_  = A199 & A167;
  assign \new_[7199]_  = A168 & \new_[7198]_ ;
  assign \new_[7203]_  = A232 & ~A203;
  assign \new_[7204]_  = ~A202 & \new_[7203]_ ;
  assign \new_[7205]_  = \new_[7204]_  & \new_[7199]_ ;
  assign \new_[7209]_  = A236 & A234;
  assign \new_[7210]_  = ~A233 & \new_[7209]_ ;
  assign \new_[7213]_  = ~A266 & A265;
  assign \new_[7216]_  = A269 & A267;
  assign \new_[7217]_  = \new_[7216]_  & \new_[7213]_ ;
  assign \new_[7218]_  = \new_[7217]_  & \new_[7210]_ ;
  assign \new_[7222]_  = A167 & A169;
  assign \new_[7223]_  = ~A170 & \new_[7222]_ ;
  assign \new_[7227]_  = ~A202 & A199;
  assign \new_[7228]_  = A166 & \new_[7227]_ ;
  assign \new_[7229]_  = \new_[7228]_  & \new_[7223]_ ;
  assign \new_[7233]_  = A233 & ~A232;
  assign \new_[7234]_  = ~A203 & \new_[7233]_ ;
  assign \new_[7237]_  = ~A299 & A298;
  assign \new_[7240]_  = A301 & A300;
  assign \new_[7241]_  = \new_[7240]_  & \new_[7237]_ ;
  assign \new_[7242]_  = \new_[7241]_  & \new_[7234]_ ;
  assign \new_[7246]_  = A167 & A169;
  assign \new_[7247]_  = ~A170 & \new_[7246]_ ;
  assign \new_[7251]_  = ~A202 & A199;
  assign \new_[7252]_  = A166 & \new_[7251]_ ;
  assign \new_[7253]_  = \new_[7252]_  & \new_[7247]_ ;
  assign \new_[7257]_  = A233 & ~A232;
  assign \new_[7258]_  = ~A203 & \new_[7257]_ ;
  assign \new_[7261]_  = ~A299 & A298;
  assign \new_[7264]_  = A302 & A300;
  assign \new_[7265]_  = \new_[7264]_  & \new_[7261]_ ;
  assign \new_[7266]_  = \new_[7265]_  & \new_[7258]_ ;
  assign \new_[7270]_  = A167 & A169;
  assign \new_[7271]_  = ~A170 & \new_[7270]_ ;
  assign \new_[7275]_  = ~A202 & A199;
  assign \new_[7276]_  = A166 & \new_[7275]_ ;
  assign \new_[7277]_  = \new_[7276]_  & \new_[7271]_ ;
  assign \new_[7281]_  = A233 & ~A232;
  assign \new_[7282]_  = ~A203 & \new_[7281]_ ;
  assign \new_[7285]_  = ~A266 & A265;
  assign \new_[7288]_  = A268 & A267;
  assign \new_[7289]_  = \new_[7288]_  & \new_[7285]_ ;
  assign \new_[7290]_  = \new_[7289]_  & \new_[7282]_ ;
  assign \new_[7294]_  = A167 & A169;
  assign \new_[7295]_  = ~A170 & \new_[7294]_ ;
  assign \new_[7299]_  = ~A202 & A199;
  assign \new_[7300]_  = A166 & \new_[7299]_ ;
  assign \new_[7301]_  = \new_[7300]_  & \new_[7295]_ ;
  assign \new_[7305]_  = A233 & ~A232;
  assign \new_[7306]_  = ~A203 & \new_[7305]_ ;
  assign \new_[7309]_  = ~A266 & A265;
  assign \new_[7312]_  = A269 & A267;
  assign \new_[7313]_  = \new_[7312]_  & \new_[7309]_ ;
  assign \new_[7314]_  = \new_[7313]_  & \new_[7306]_ ;
  assign \new_[7318]_  = A167 & A169;
  assign \new_[7319]_  = ~A170 & \new_[7318]_ ;
  assign \new_[7323]_  = ~A202 & A199;
  assign \new_[7324]_  = A166 & \new_[7323]_ ;
  assign \new_[7325]_  = \new_[7324]_  & \new_[7319]_ ;
  assign \new_[7329]_  = ~A233 & A232;
  assign \new_[7330]_  = ~A203 & \new_[7329]_ ;
  assign \new_[7333]_  = A235 & A234;
  assign \new_[7336]_  = A299 & ~A298;
  assign \new_[7337]_  = \new_[7336]_  & \new_[7333]_ ;
  assign \new_[7338]_  = \new_[7337]_  & \new_[7330]_ ;
  assign \new_[7342]_  = A167 & A169;
  assign \new_[7343]_  = ~A170 & \new_[7342]_ ;
  assign \new_[7347]_  = ~A202 & A199;
  assign \new_[7348]_  = A166 & \new_[7347]_ ;
  assign \new_[7349]_  = \new_[7348]_  & \new_[7343]_ ;
  assign \new_[7353]_  = ~A233 & A232;
  assign \new_[7354]_  = ~A203 & \new_[7353]_ ;
  assign \new_[7357]_  = A235 & A234;
  assign \new_[7360]_  = A266 & ~A265;
  assign \new_[7361]_  = \new_[7360]_  & \new_[7357]_ ;
  assign \new_[7362]_  = \new_[7361]_  & \new_[7354]_ ;
  assign \new_[7366]_  = A167 & A169;
  assign \new_[7367]_  = ~A170 & \new_[7366]_ ;
  assign \new_[7371]_  = ~A202 & A199;
  assign \new_[7372]_  = A166 & \new_[7371]_ ;
  assign \new_[7373]_  = \new_[7372]_  & \new_[7367]_ ;
  assign \new_[7377]_  = ~A233 & A232;
  assign \new_[7378]_  = ~A203 & \new_[7377]_ ;
  assign \new_[7381]_  = A236 & A234;
  assign \new_[7384]_  = A299 & ~A298;
  assign \new_[7385]_  = \new_[7384]_  & \new_[7381]_ ;
  assign \new_[7386]_  = \new_[7385]_  & \new_[7378]_ ;
  assign \new_[7390]_  = A167 & A169;
  assign \new_[7391]_  = ~A170 & \new_[7390]_ ;
  assign \new_[7395]_  = ~A202 & A199;
  assign \new_[7396]_  = A166 & \new_[7395]_ ;
  assign \new_[7397]_  = \new_[7396]_  & \new_[7391]_ ;
  assign \new_[7401]_  = ~A233 & A232;
  assign \new_[7402]_  = ~A203 & \new_[7401]_ ;
  assign \new_[7405]_  = A236 & A234;
  assign \new_[7408]_  = A266 & ~A265;
  assign \new_[7409]_  = \new_[7408]_  & \new_[7405]_ ;
  assign \new_[7410]_  = \new_[7409]_  & \new_[7402]_ ;
  assign \new_[7414]_  = ~A167 & A169;
  assign \new_[7415]_  = ~A170 & \new_[7414]_ ;
  assign \new_[7419]_  = ~A202 & A199;
  assign \new_[7420]_  = ~A166 & \new_[7419]_ ;
  assign \new_[7421]_  = \new_[7420]_  & \new_[7415]_ ;
  assign \new_[7425]_  = A233 & ~A232;
  assign \new_[7426]_  = ~A203 & \new_[7425]_ ;
  assign \new_[7429]_  = ~A299 & A298;
  assign \new_[7432]_  = A301 & A300;
  assign \new_[7433]_  = \new_[7432]_  & \new_[7429]_ ;
  assign \new_[7434]_  = \new_[7433]_  & \new_[7426]_ ;
  assign \new_[7438]_  = ~A167 & A169;
  assign \new_[7439]_  = ~A170 & \new_[7438]_ ;
  assign \new_[7443]_  = ~A202 & A199;
  assign \new_[7444]_  = ~A166 & \new_[7443]_ ;
  assign \new_[7445]_  = \new_[7444]_  & \new_[7439]_ ;
  assign \new_[7449]_  = A233 & ~A232;
  assign \new_[7450]_  = ~A203 & \new_[7449]_ ;
  assign \new_[7453]_  = ~A299 & A298;
  assign \new_[7456]_  = A302 & A300;
  assign \new_[7457]_  = \new_[7456]_  & \new_[7453]_ ;
  assign \new_[7458]_  = \new_[7457]_  & \new_[7450]_ ;
  assign \new_[7462]_  = ~A167 & A169;
  assign \new_[7463]_  = ~A170 & \new_[7462]_ ;
  assign \new_[7467]_  = ~A202 & A199;
  assign \new_[7468]_  = ~A166 & \new_[7467]_ ;
  assign \new_[7469]_  = \new_[7468]_  & \new_[7463]_ ;
  assign \new_[7473]_  = A233 & ~A232;
  assign \new_[7474]_  = ~A203 & \new_[7473]_ ;
  assign \new_[7477]_  = ~A266 & A265;
  assign \new_[7480]_  = A268 & A267;
  assign \new_[7481]_  = \new_[7480]_  & \new_[7477]_ ;
  assign \new_[7482]_  = \new_[7481]_  & \new_[7474]_ ;
  assign \new_[7486]_  = ~A167 & A169;
  assign \new_[7487]_  = ~A170 & \new_[7486]_ ;
  assign \new_[7491]_  = ~A202 & A199;
  assign \new_[7492]_  = ~A166 & \new_[7491]_ ;
  assign \new_[7493]_  = \new_[7492]_  & \new_[7487]_ ;
  assign \new_[7497]_  = A233 & ~A232;
  assign \new_[7498]_  = ~A203 & \new_[7497]_ ;
  assign \new_[7501]_  = ~A266 & A265;
  assign \new_[7504]_  = A269 & A267;
  assign \new_[7505]_  = \new_[7504]_  & \new_[7501]_ ;
  assign \new_[7506]_  = \new_[7505]_  & \new_[7498]_ ;
  assign \new_[7510]_  = ~A167 & A169;
  assign \new_[7511]_  = ~A170 & \new_[7510]_ ;
  assign \new_[7515]_  = ~A202 & A199;
  assign \new_[7516]_  = ~A166 & \new_[7515]_ ;
  assign \new_[7517]_  = \new_[7516]_  & \new_[7511]_ ;
  assign \new_[7521]_  = ~A233 & A232;
  assign \new_[7522]_  = ~A203 & \new_[7521]_ ;
  assign \new_[7525]_  = A235 & A234;
  assign \new_[7528]_  = A299 & ~A298;
  assign \new_[7529]_  = \new_[7528]_  & \new_[7525]_ ;
  assign \new_[7530]_  = \new_[7529]_  & \new_[7522]_ ;
  assign \new_[7534]_  = ~A167 & A169;
  assign \new_[7535]_  = ~A170 & \new_[7534]_ ;
  assign \new_[7539]_  = ~A202 & A199;
  assign \new_[7540]_  = ~A166 & \new_[7539]_ ;
  assign \new_[7541]_  = \new_[7540]_  & \new_[7535]_ ;
  assign \new_[7545]_  = ~A233 & A232;
  assign \new_[7546]_  = ~A203 & \new_[7545]_ ;
  assign \new_[7549]_  = A235 & A234;
  assign \new_[7552]_  = A266 & ~A265;
  assign \new_[7553]_  = \new_[7552]_  & \new_[7549]_ ;
  assign \new_[7554]_  = \new_[7553]_  & \new_[7546]_ ;
  assign \new_[7558]_  = ~A167 & A169;
  assign \new_[7559]_  = ~A170 & \new_[7558]_ ;
  assign \new_[7563]_  = ~A202 & A199;
  assign \new_[7564]_  = ~A166 & \new_[7563]_ ;
  assign \new_[7565]_  = \new_[7564]_  & \new_[7559]_ ;
  assign \new_[7569]_  = ~A233 & A232;
  assign \new_[7570]_  = ~A203 & \new_[7569]_ ;
  assign \new_[7573]_  = A236 & A234;
  assign \new_[7576]_  = A299 & ~A298;
  assign \new_[7577]_  = \new_[7576]_  & \new_[7573]_ ;
  assign \new_[7578]_  = \new_[7577]_  & \new_[7570]_ ;
  assign \new_[7582]_  = ~A167 & A169;
  assign \new_[7583]_  = ~A170 & \new_[7582]_ ;
  assign \new_[7587]_  = ~A202 & A199;
  assign \new_[7588]_  = ~A166 & \new_[7587]_ ;
  assign \new_[7589]_  = \new_[7588]_  & \new_[7583]_ ;
  assign \new_[7593]_  = ~A233 & A232;
  assign \new_[7594]_  = ~A203 & \new_[7593]_ ;
  assign \new_[7597]_  = A236 & A234;
  assign \new_[7600]_  = A266 & ~A265;
  assign \new_[7601]_  = \new_[7600]_  & \new_[7597]_ ;
  assign \new_[7602]_  = \new_[7601]_  & \new_[7594]_ ;
  assign \new_[7606]_  = A167 & ~A169;
  assign \new_[7607]_  = A170 & \new_[7606]_ ;
  assign \new_[7611]_  = ~A202 & A199;
  assign \new_[7612]_  = ~A166 & \new_[7611]_ ;
  assign \new_[7613]_  = \new_[7612]_  & \new_[7607]_ ;
  assign \new_[7617]_  = A233 & ~A232;
  assign \new_[7618]_  = ~A203 & \new_[7617]_ ;
  assign \new_[7621]_  = ~A299 & A298;
  assign \new_[7624]_  = A301 & A300;
  assign \new_[7625]_  = \new_[7624]_  & \new_[7621]_ ;
  assign \new_[7626]_  = \new_[7625]_  & \new_[7618]_ ;
  assign \new_[7630]_  = A167 & ~A169;
  assign \new_[7631]_  = A170 & \new_[7630]_ ;
  assign \new_[7635]_  = ~A202 & A199;
  assign \new_[7636]_  = ~A166 & \new_[7635]_ ;
  assign \new_[7637]_  = \new_[7636]_  & \new_[7631]_ ;
  assign \new_[7641]_  = A233 & ~A232;
  assign \new_[7642]_  = ~A203 & \new_[7641]_ ;
  assign \new_[7645]_  = ~A299 & A298;
  assign \new_[7648]_  = A302 & A300;
  assign \new_[7649]_  = \new_[7648]_  & \new_[7645]_ ;
  assign \new_[7650]_  = \new_[7649]_  & \new_[7642]_ ;
  assign \new_[7654]_  = A167 & ~A169;
  assign \new_[7655]_  = A170 & \new_[7654]_ ;
  assign \new_[7659]_  = ~A202 & A199;
  assign \new_[7660]_  = ~A166 & \new_[7659]_ ;
  assign \new_[7661]_  = \new_[7660]_  & \new_[7655]_ ;
  assign \new_[7665]_  = A233 & ~A232;
  assign \new_[7666]_  = ~A203 & \new_[7665]_ ;
  assign \new_[7669]_  = ~A266 & A265;
  assign \new_[7672]_  = A268 & A267;
  assign \new_[7673]_  = \new_[7672]_  & \new_[7669]_ ;
  assign \new_[7674]_  = \new_[7673]_  & \new_[7666]_ ;
  assign \new_[7678]_  = A167 & ~A169;
  assign \new_[7679]_  = A170 & \new_[7678]_ ;
  assign \new_[7683]_  = ~A202 & A199;
  assign \new_[7684]_  = ~A166 & \new_[7683]_ ;
  assign \new_[7685]_  = \new_[7684]_  & \new_[7679]_ ;
  assign \new_[7689]_  = A233 & ~A232;
  assign \new_[7690]_  = ~A203 & \new_[7689]_ ;
  assign \new_[7693]_  = ~A266 & A265;
  assign \new_[7696]_  = A269 & A267;
  assign \new_[7697]_  = \new_[7696]_  & \new_[7693]_ ;
  assign \new_[7698]_  = \new_[7697]_  & \new_[7690]_ ;
  assign \new_[7702]_  = A167 & ~A169;
  assign \new_[7703]_  = A170 & \new_[7702]_ ;
  assign \new_[7707]_  = ~A202 & A199;
  assign \new_[7708]_  = ~A166 & \new_[7707]_ ;
  assign \new_[7709]_  = \new_[7708]_  & \new_[7703]_ ;
  assign \new_[7713]_  = ~A233 & A232;
  assign \new_[7714]_  = ~A203 & \new_[7713]_ ;
  assign \new_[7717]_  = A235 & A234;
  assign \new_[7720]_  = A299 & ~A298;
  assign \new_[7721]_  = \new_[7720]_  & \new_[7717]_ ;
  assign \new_[7722]_  = \new_[7721]_  & \new_[7714]_ ;
  assign \new_[7726]_  = A167 & ~A169;
  assign \new_[7727]_  = A170 & \new_[7726]_ ;
  assign \new_[7731]_  = ~A202 & A199;
  assign \new_[7732]_  = ~A166 & \new_[7731]_ ;
  assign \new_[7733]_  = \new_[7732]_  & \new_[7727]_ ;
  assign \new_[7737]_  = ~A233 & A232;
  assign \new_[7738]_  = ~A203 & \new_[7737]_ ;
  assign \new_[7741]_  = A235 & A234;
  assign \new_[7744]_  = A266 & ~A265;
  assign \new_[7745]_  = \new_[7744]_  & \new_[7741]_ ;
  assign \new_[7746]_  = \new_[7745]_  & \new_[7738]_ ;
  assign \new_[7750]_  = A167 & ~A169;
  assign \new_[7751]_  = A170 & \new_[7750]_ ;
  assign \new_[7755]_  = ~A202 & A199;
  assign \new_[7756]_  = ~A166 & \new_[7755]_ ;
  assign \new_[7757]_  = \new_[7756]_  & \new_[7751]_ ;
  assign \new_[7761]_  = ~A233 & A232;
  assign \new_[7762]_  = ~A203 & \new_[7761]_ ;
  assign \new_[7765]_  = A236 & A234;
  assign \new_[7768]_  = A299 & ~A298;
  assign \new_[7769]_  = \new_[7768]_  & \new_[7765]_ ;
  assign \new_[7770]_  = \new_[7769]_  & \new_[7762]_ ;
  assign \new_[7774]_  = A167 & ~A169;
  assign \new_[7775]_  = A170 & \new_[7774]_ ;
  assign \new_[7779]_  = ~A202 & A199;
  assign \new_[7780]_  = ~A166 & \new_[7779]_ ;
  assign \new_[7781]_  = \new_[7780]_  & \new_[7775]_ ;
  assign \new_[7785]_  = ~A233 & A232;
  assign \new_[7786]_  = ~A203 & \new_[7785]_ ;
  assign \new_[7789]_  = A236 & A234;
  assign \new_[7792]_  = A266 & ~A265;
  assign \new_[7793]_  = \new_[7792]_  & \new_[7789]_ ;
  assign \new_[7794]_  = \new_[7793]_  & \new_[7786]_ ;
  assign \new_[7798]_  = ~A167 & ~A169;
  assign \new_[7799]_  = A170 & \new_[7798]_ ;
  assign \new_[7803]_  = ~A202 & A199;
  assign \new_[7804]_  = A166 & \new_[7803]_ ;
  assign \new_[7805]_  = \new_[7804]_  & \new_[7799]_ ;
  assign \new_[7809]_  = A233 & ~A232;
  assign \new_[7810]_  = ~A203 & \new_[7809]_ ;
  assign \new_[7813]_  = ~A299 & A298;
  assign \new_[7816]_  = A301 & A300;
  assign \new_[7817]_  = \new_[7816]_  & \new_[7813]_ ;
  assign \new_[7818]_  = \new_[7817]_  & \new_[7810]_ ;
  assign \new_[7822]_  = ~A167 & ~A169;
  assign \new_[7823]_  = A170 & \new_[7822]_ ;
  assign \new_[7827]_  = ~A202 & A199;
  assign \new_[7828]_  = A166 & \new_[7827]_ ;
  assign \new_[7829]_  = \new_[7828]_  & \new_[7823]_ ;
  assign \new_[7833]_  = A233 & ~A232;
  assign \new_[7834]_  = ~A203 & \new_[7833]_ ;
  assign \new_[7837]_  = ~A299 & A298;
  assign \new_[7840]_  = A302 & A300;
  assign \new_[7841]_  = \new_[7840]_  & \new_[7837]_ ;
  assign \new_[7842]_  = \new_[7841]_  & \new_[7834]_ ;
  assign \new_[7846]_  = ~A167 & ~A169;
  assign \new_[7847]_  = A170 & \new_[7846]_ ;
  assign \new_[7851]_  = ~A202 & A199;
  assign \new_[7852]_  = A166 & \new_[7851]_ ;
  assign \new_[7853]_  = \new_[7852]_  & \new_[7847]_ ;
  assign \new_[7857]_  = A233 & ~A232;
  assign \new_[7858]_  = ~A203 & \new_[7857]_ ;
  assign \new_[7861]_  = ~A266 & A265;
  assign \new_[7864]_  = A268 & A267;
  assign \new_[7865]_  = \new_[7864]_  & \new_[7861]_ ;
  assign \new_[7866]_  = \new_[7865]_  & \new_[7858]_ ;
  assign \new_[7870]_  = ~A167 & ~A169;
  assign \new_[7871]_  = A170 & \new_[7870]_ ;
  assign \new_[7875]_  = ~A202 & A199;
  assign \new_[7876]_  = A166 & \new_[7875]_ ;
  assign \new_[7877]_  = \new_[7876]_  & \new_[7871]_ ;
  assign \new_[7881]_  = A233 & ~A232;
  assign \new_[7882]_  = ~A203 & \new_[7881]_ ;
  assign \new_[7885]_  = ~A266 & A265;
  assign \new_[7888]_  = A269 & A267;
  assign \new_[7889]_  = \new_[7888]_  & \new_[7885]_ ;
  assign \new_[7890]_  = \new_[7889]_  & \new_[7882]_ ;
  assign \new_[7894]_  = ~A167 & ~A169;
  assign \new_[7895]_  = A170 & \new_[7894]_ ;
  assign \new_[7899]_  = ~A202 & A199;
  assign \new_[7900]_  = A166 & \new_[7899]_ ;
  assign \new_[7901]_  = \new_[7900]_  & \new_[7895]_ ;
  assign \new_[7905]_  = ~A233 & A232;
  assign \new_[7906]_  = ~A203 & \new_[7905]_ ;
  assign \new_[7909]_  = A235 & A234;
  assign \new_[7912]_  = A299 & ~A298;
  assign \new_[7913]_  = \new_[7912]_  & \new_[7909]_ ;
  assign \new_[7914]_  = \new_[7913]_  & \new_[7906]_ ;
  assign \new_[7918]_  = ~A167 & ~A169;
  assign \new_[7919]_  = A170 & \new_[7918]_ ;
  assign \new_[7923]_  = ~A202 & A199;
  assign \new_[7924]_  = A166 & \new_[7923]_ ;
  assign \new_[7925]_  = \new_[7924]_  & \new_[7919]_ ;
  assign \new_[7929]_  = ~A233 & A232;
  assign \new_[7930]_  = ~A203 & \new_[7929]_ ;
  assign \new_[7933]_  = A235 & A234;
  assign \new_[7936]_  = A266 & ~A265;
  assign \new_[7937]_  = \new_[7936]_  & \new_[7933]_ ;
  assign \new_[7938]_  = \new_[7937]_  & \new_[7930]_ ;
  assign \new_[7942]_  = ~A167 & ~A169;
  assign \new_[7943]_  = A170 & \new_[7942]_ ;
  assign \new_[7947]_  = ~A202 & A199;
  assign \new_[7948]_  = A166 & \new_[7947]_ ;
  assign \new_[7949]_  = \new_[7948]_  & \new_[7943]_ ;
  assign \new_[7953]_  = ~A233 & A232;
  assign \new_[7954]_  = ~A203 & \new_[7953]_ ;
  assign \new_[7957]_  = A236 & A234;
  assign \new_[7960]_  = A299 & ~A298;
  assign \new_[7961]_  = \new_[7960]_  & \new_[7957]_ ;
  assign \new_[7962]_  = \new_[7961]_  & \new_[7954]_ ;
  assign \new_[7966]_  = ~A167 & ~A169;
  assign \new_[7967]_  = A170 & \new_[7966]_ ;
  assign \new_[7971]_  = ~A202 & A199;
  assign \new_[7972]_  = A166 & \new_[7971]_ ;
  assign \new_[7973]_  = \new_[7972]_  & \new_[7967]_ ;
  assign \new_[7977]_  = ~A233 & A232;
  assign \new_[7978]_  = ~A203 & \new_[7977]_ ;
  assign \new_[7981]_  = A236 & A234;
  assign \new_[7984]_  = A266 & ~A265;
  assign \new_[7985]_  = \new_[7984]_  & \new_[7981]_ ;
  assign \new_[7986]_  = \new_[7985]_  & \new_[7978]_ ;
  assign \new_[7990]_  = A167 & A169;
  assign \new_[7991]_  = ~A170 & \new_[7990]_ ;
  assign \new_[7994]_  = A199 & A166;
  assign \new_[7997]_  = A232 & ~A201;
  assign \new_[7998]_  = \new_[7997]_  & \new_[7994]_ ;
  assign \new_[7999]_  = \new_[7998]_  & \new_[7991]_ ;
  assign \new_[8003]_  = A235 & A234;
  assign \new_[8004]_  = ~A233 & \new_[8003]_ ;
  assign \new_[8007]_  = ~A299 & A298;
  assign \new_[8010]_  = A301 & A300;
  assign \new_[8011]_  = \new_[8010]_  & \new_[8007]_ ;
  assign \new_[8012]_  = \new_[8011]_  & \new_[8004]_ ;
  assign \new_[8016]_  = A167 & A169;
  assign \new_[8017]_  = ~A170 & \new_[8016]_ ;
  assign \new_[8020]_  = A199 & A166;
  assign \new_[8023]_  = A232 & ~A201;
  assign \new_[8024]_  = \new_[8023]_  & \new_[8020]_ ;
  assign \new_[8025]_  = \new_[8024]_  & \new_[8017]_ ;
  assign \new_[8029]_  = A235 & A234;
  assign \new_[8030]_  = ~A233 & \new_[8029]_ ;
  assign \new_[8033]_  = ~A299 & A298;
  assign \new_[8036]_  = A302 & A300;
  assign \new_[8037]_  = \new_[8036]_  & \new_[8033]_ ;
  assign \new_[8038]_  = \new_[8037]_  & \new_[8030]_ ;
  assign \new_[8042]_  = A167 & A169;
  assign \new_[8043]_  = ~A170 & \new_[8042]_ ;
  assign \new_[8046]_  = A199 & A166;
  assign \new_[8049]_  = A232 & ~A201;
  assign \new_[8050]_  = \new_[8049]_  & \new_[8046]_ ;
  assign \new_[8051]_  = \new_[8050]_  & \new_[8043]_ ;
  assign \new_[8055]_  = A235 & A234;
  assign \new_[8056]_  = ~A233 & \new_[8055]_ ;
  assign \new_[8059]_  = ~A266 & A265;
  assign \new_[8062]_  = A268 & A267;
  assign \new_[8063]_  = \new_[8062]_  & \new_[8059]_ ;
  assign \new_[8064]_  = \new_[8063]_  & \new_[8056]_ ;
  assign \new_[8068]_  = A167 & A169;
  assign \new_[8069]_  = ~A170 & \new_[8068]_ ;
  assign \new_[8072]_  = A199 & A166;
  assign \new_[8075]_  = A232 & ~A201;
  assign \new_[8076]_  = \new_[8075]_  & \new_[8072]_ ;
  assign \new_[8077]_  = \new_[8076]_  & \new_[8069]_ ;
  assign \new_[8081]_  = A235 & A234;
  assign \new_[8082]_  = ~A233 & \new_[8081]_ ;
  assign \new_[8085]_  = ~A266 & A265;
  assign \new_[8088]_  = A269 & A267;
  assign \new_[8089]_  = \new_[8088]_  & \new_[8085]_ ;
  assign \new_[8090]_  = \new_[8089]_  & \new_[8082]_ ;
  assign \new_[8094]_  = A167 & A169;
  assign \new_[8095]_  = ~A170 & \new_[8094]_ ;
  assign \new_[8098]_  = A199 & A166;
  assign \new_[8101]_  = A232 & ~A201;
  assign \new_[8102]_  = \new_[8101]_  & \new_[8098]_ ;
  assign \new_[8103]_  = \new_[8102]_  & \new_[8095]_ ;
  assign \new_[8107]_  = A236 & A234;
  assign \new_[8108]_  = ~A233 & \new_[8107]_ ;
  assign \new_[8111]_  = ~A299 & A298;
  assign \new_[8114]_  = A301 & A300;
  assign \new_[8115]_  = \new_[8114]_  & \new_[8111]_ ;
  assign \new_[8116]_  = \new_[8115]_  & \new_[8108]_ ;
  assign \new_[8120]_  = A167 & A169;
  assign \new_[8121]_  = ~A170 & \new_[8120]_ ;
  assign \new_[8124]_  = A199 & A166;
  assign \new_[8127]_  = A232 & ~A201;
  assign \new_[8128]_  = \new_[8127]_  & \new_[8124]_ ;
  assign \new_[8129]_  = \new_[8128]_  & \new_[8121]_ ;
  assign \new_[8133]_  = A236 & A234;
  assign \new_[8134]_  = ~A233 & \new_[8133]_ ;
  assign \new_[8137]_  = ~A299 & A298;
  assign \new_[8140]_  = A302 & A300;
  assign \new_[8141]_  = \new_[8140]_  & \new_[8137]_ ;
  assign \new_[8142]_  = \new_[8141]_  & \new_[8134]_ ;
  assign \new_[8146]_  = A167 & A169;
  assign \new_[8147]_  = ~A170 & \new_[8146]_ ;
  assign \new_[8150]_  = A199 & A166;
  assign \new_[8153]_  = A232 & ~A201;
  assign \new_[8154]_  = \new_[8153]_  & \new_[8150]_ ;
  assign \new_[8155]_  = \new_[8154]_  & \new_[8147]_ ;
  assign \new_[8159]_  = A236 & A234;
  assign \new_[8160]_  = ~A233 & \new_[8159]_ ;
  assign \new_[8163]_  = ~A266 & A265;
  assign \new_[8166]_  = A268 & A267;
  assign \new_[8167]_  = \new_[8166]_  & \new_[8163]_ ;
  assign \new_[8168]_  = \new_[8167]_  & \new_[8160]_ ;
  assign \new_[8172]_  = A167 & A169;
  assign \new_[8173]_  = ~A170 & \new_[8172]_ ;
  assign \new_[8176]_  = A199 & A166;
  assign \new_[8179]_  = A232 & ~A201;
  assign \new_[8180]_  = \new_[8179]_  & \new_[8176]_ ;
  assign \new_[8181]_  = \new_[8180]_  & \new_[8173]_ ;
  assign \new_[8185]_  = A236 & A234;
  assign \new_[8186]_  = ~A233 & \new_[8185]_ ;
  assign \new_[8189]_  = ~A266 & A265;
  assign \new_[8192]_  = A269 & A267;
  assign \new_[8193]_  = \new_[8192]_  & \new_[8189]_ ;
  assign \new_[8194]_  = \new_[8193]_  & \new_[8186]_ ;
  assign \new_[8198]_  = A167 & A169;
  assign \new_[8199]_  = ~A170 & \new_[8198]_ ;
  assign \new_[8202]_  = A199 & A166;
  assign \new_[8205]_  = A232 & A200;
  assign \new_[8206]_  = \new_[8205]_  & \new_[8202]_ ;
  assign \new_[8207]_  = \new_[8206]_  & \new_[8199]_ ;
  assign \new_[8211]_  = A235 & A234;
  assign \new_[8212]_  = ~A233 & \new_[8211]_ ;
  assign \new_[8215]_  = ~A299 & A298;
  assign \new_[8218]_  = A301 & A300;
  assign \new_[8219]_  = \new_[8218]_  & \new_[8215]_ ;
  assign \new_[8220]_  = \new_[8219]_  & \new_[8212]_ ;
  assign \new_[8224]_  = A167 & A169;
  assign \new_[8225]_  = ~A170 & \new_[8224]_ ;
  assign \new_[8228]_  = A199 & A166;
  assign \new_[8231]_  = A232 & A200;
  assign \new_[8232]_  = \new_[8231]_  & \new_[8228]_ ;
  assign \new_[8233]_  = \new_[8232]_  & \new_[8225]_ ;
  assign \new_[8237]_  = A235 & A234;
  assign \new_[8238]_  = ~A233 & \new_[8237]_ ;
  assign \new_[8241]_  = ~A299 & A298;
  assign \new_[8244]_  = A302 & A300;
  assign \new_[8245]_  = \new_[8244]_  & \new_[8241]_ ;
  assign \new_[8246]_  = \new_[8245]_  & \new_[8238]_ ;
  assign \new_[8250]_  = A167 & A169;
  assign \new_[8251]_  = ~A170 & \new_[8250]_ ;
  assign \new_[8254]_  = A199 & A166;
  assign \new_[8257]_  = A232 & A200;
  assign \new_[8258]_  = \new_[8257]_  & \new_[8254]_ ;
  assign \new_[8259]_  = \new_[8258]_  & \new_[8251]_ ;
  assign \new_[8263]_  = A235 & A234;
  assign \new_[8264]_  = ~A233 & \new_[8263]_ ;
  assign \new_[8267]_  = ~A266 & A265;
  assign \new_[8270]_  = A268 & A267;
  assign \new_[8271]_  = \new_[8270]_  & \new_[8267]_ ;
  assign \new_[8272]_  = \new_[8271]_  & \new_[8264]_ ;
  assign \new_[8276]_  = A167 & A169;
  assign \new_[8277]_  = ~A170 & \new_[8276]_ ;
  assign \new_[8280]_  = A199 & A166;
  assign \new_[8283]_  = A232 & A200;
  assign \new_[8284]_  = \new_[8283]_  & \new_[8280]_ ;
  assign \new_[8285]_  = \new_[8284]_  & \new_[8277]_ ;
  assign \new_[8289]_  = A235 & A234;
  assign \new_[8290]_  = ~A233 & \new_[8289]_ ;
  assign \new_[8293]_  = ~A266 & A265;
  assign \new_[8296]_  = A269 & A267;
  assign \new_[8297]_  = \new_[8296]_  & \new_[8293]_ ;
  assign \new_[8298]_  = \new_[8297]_  & \new_[8290]_ ;
  assign \new_[8302]_  = A167 & A169;
  assign \new_[8303]_  = ~A170 & \new_[8302]_ ;
  assign \new_[8306]_  = A199 & A166;
  assign \new_[8309]_  = A232 & A200;
  assign \new_[8310]_  = \new_[8309]_  & \new_[8306]_ ;
  assign \new_[8311]_  = \new_[8310]_  & \new_[8303]_ ;
  assign \new_[8315]_  = A236 & A234;
  assign \new_[8316]_  = ~A233 & \new_[8315]_ ;
  assign \new_[8319]_  = ~A299 & A298;
  assign \new_[8322]_  = A301 & A300;
  assign \new_[8323]_  = \new_[8322]_  & \new_[8319]_ ;
  assign \new_[8324]_  = \new_[8323]_  & \new_[8316]_ ;
  assign \new_[8328]_  = A167 & A169;
  assign \new_[8329]_  = ~A170 & \new_[8328]_ ;
  assign \new_[8332]_  = A199 & A166;
  assign \new_[8335]_  = A232 & A200;
  assign \new_[8336]_  = \new_[8335]_  & \new_[8332]_ ;
  assign \new_[8337]_  = \new_[8336]_  & \new_[8329]_ ;
  assign \new_[8341]_  = A236 & A234;
  assign \new_[8342]_  = ~A233 & \new_[8341]_ ;
  assign \new_[8345]_  = ~A299 & A298;
  assign \new_[8348]_  = A302 & A300;
  assign \new_[8349]_  = \new_[8348]_  & \new_[8345]_ ;
  assign \new_[8350]_  = \new_[8349]_  & \new_[8342]_ ;
  assign \new_[8354]_  = A167 & A169;
  assign \new_[8355]_  = ~A170 & \new_[8354]_ ;
  assign \new_[8358]_  = A199 & A166;
  assign \new_[8361]_  = A232 & A200;
  assign \new_[8362]_  = \new_[8361]_  & \new_[8358]_ ;
  assign \new_[8363]_  = \new_[8362]_  & \new_[8355]_ ;
  assign \new_[8367]_  = A236 & A234;
  assign \new_[8368]_  = ~A233 & \new_[8367]_ ;
  assign \new_[8371]_  = ~A266 & A265;
  assign \new_[8374]_  = A268 & A267;
  assign \new_[8375]_  = \new_[8374]_  & \new_[8371]_ ;
  assign \new_[8376]_  = \new_[8375]_  & \new_[8368]_ ;
  assign \new_[8380]_  = A167 & A169;
  assign \new_[8381]_  = ~A170 & \new_[8380]_ ;
  assign \new_[8384]_  = A199 & A166;
  assign \new_[8387]_  = A232 & A200;
  assign \new_[8388]_  = \new_[8387]_  & \new_[8384]_ ;
  assign \new_[8389]_  = \new_[8388]_  & \new_[8381]_ ;
  assign \new_[8393]_  = A236 & A234;
  assign \new_[8394]_  = ~A233 & \new_[8393]_ ;
  assign \new_[8397]_  = ~A266 & A265;
  assign \new_[8400]_  = A269 & A267;
  assign \new_[8401]_  = \new_[8400]_  & \new_[8397]_ ;
  assign \new_[8402]_  = \new_[8401]_  & \new_[8394]_ ;
  assign \new_[8406]_  = A167 & A169;
  assign \new_[8407]_  = ~A170 & \new_[8406]_ ;
  assign \new_[8410]_  = ~A199 & A166;
  assign \new_[8413]_  = A232 & ~A200;
  assign \new_[8414]_  = \new_[8413]_  & \new_[8410]_ ;
  assign \new_[8415]_  = \new_[8414]_  & \new_[8407]_ ;
  assign \new_[8419]_  = A235 & A234;
  assign \new_[8420]_  = ~A233 & \new_[8419]_ ;
  assign \new_[8423]_  = ~A299 & A298;
  assign \new_[8426]_  = A301 & A300;
  assign \new_[8427]_  = \new_[8426]_  & \new_[8423]_ ;
  assign \new_[8428]_  = \new_[8427]_  & \new_[8420]_ ;
  assign \new_[8432]_  = A167 & A169;
  assign \new_[8433]_  = ~A170 & \new_[8432]_ ;
  assign \new_[8436]_  = ~A199 & A166;
  assign \new_[8439]_  = A232 & ~A200;
  assign \new_[8440]_  = \new_[8439]_  & \new_[8436]_ ;
  assign \new_[8441]_  = \new_[8440]_  & \new_[8433]_ ;
  assign \new_[8445]_  = A235 & A234;
  assign \new_[8446]_  = ~A233 & \new_[8445]_ ;
  assign \new_[8449]_  = ~A299 & A298;
  assign \new_[8452]_  = A302 & A300;
  assign \new_[8453]_  = \new_[8452]_  & \new_[8449]_ ;
  assign \new_[8454]_  = \new_[8453]_  & \new_[8446]_ ;
  assign \new_[8458]_  = A167 & A169;
  assign \new_[8459]_  = ~A170 & \new_[8458]_ ;
  assign \new_[8462]_  = ~A199 & A166;
  assign \new_[8465]_  = A232 & ~A200;
  assign \new_[8466]_  = \new_[8465]_  & \new_[8462]_ ;
  assign \new_[8467]_  = \new_[8466]_  & \new_[8459]_ ;
  assign \new_[8471]_  = A235 & A234;
  assign \new_[8472]_  = ~A233 & \new_[8471]_ ;
  assign \new_[8475]_  = ~A266 & A265;
  assign \new_[8478]_  = A268 & A267;
  assign \new_[8479]_  = \new_[8478]_  & \new_[8475]_ ;
  assign \new_[8480]_  = \new_[8479]_  & \new_[8472]_ ;
  assign \new_[8484]_  = A167 & A169;
  assign \new_[8485]_  = ~A170 & \new_[8484]_ ;
  assign \new_[8488]_  = ~A199 & A166;
  assign \new_[8491]_  = A232 & ~A200;
  assign \new_[8492]_  = \new_[8491]_  & \new_[8488]_ ;
  assign \new_[8493]_  = \new_[8492]_  & \new_[8485]_ ;
  assign \new_[8497]_  = A235 & A234;
  assign \new_[8498]_  = ~A233 & \new_[8497]_ ;
  assign \new_[8501]_  = ~A266 & A265;
  assign \new_[8504]_  = A269 & A267;
  assign \new_[8505]_  = \new_[8504]_  & \new_[8501]_ ;
  assign \new_[8506]_  = \new_[8505]_  & \new_[8498]_ ;
  assign \new_[8510]_  = A167 & A169;
  assign \new_[8511]_  = ~A170 & \new_[8510]_ ;
  assign \new_[8514]_  = ~A199 & A166;
  assign \new_[8517]_  = A232 & ~A200;
  assign \new_[8518]_  = \new_[8517]_  & \new_[8514]_ ;
  assign \new_[8519]_  = \new_[8518]_  & \new_[8511]_ ;
  assign \new_[8523]_  = A236 & A234;
  assign \new_[8524]_  = ~A233 & \new_[8523]_ ;
  assign \new_[8527]_  = ~A299 & A298;
  assign \new_[8530]_  = A301 & A300;
  assign \new_[8531]_  = \new_[8530]_  & \new_[8527]_ ;
  assign \new_[8532]_  = \new_[8531]_  & \new_[8524]_ ;
  assign \new_[8536]_  = A167 & A169;
  assign \new_[8537]_  = ~A170 & \new_[8536]_ ;
  assign \new_[8540]_  = ~A199 & A166;
  assign \new_[8543]_  = A232 & ~A200;
  assign \new_[8544]_  = \new_[8543]_  & \new_[8540]_ ;
  assign \new_[8545]_  = \new_[8544]_  & \new_[8537]_ ;
  assign \new_[8549]_  = A236 & A234;
  assign \new_[8550]_  = ~A233 & \new_[8549]_ ;
  assign \new_[8553]_  = ~A299 & A298;
  assign \new_[8556]_  = A302 & A300;
  assign \new_[8557]_  = \new_[8556]_  & \new_[8553]_ ;
  assign \new_[8558]_  = \new_[8557]_  & \new_[8550]_ ;
  assign \new_[8562]_  = A167 & A169;
  assign \new_[8563]_  = ~A170 & \new_[8562]_ ;
  assign \new_[8566]_  = ~A199 & A166;
  assign \new_[8569]_  = A232 & ~A200;
  assign \new_[8570]_  = \new_[8569]_  & \new_[8566]_ ;
  assign \new_[8571]_  = \new_[8570]_  & \new_[8563]_ ;
  assign \new_[8575]_  = A236 & A234;
  assign \new_[8576]_  = ~A233 & \new_[8575]_ ;
  assign \new_[8579]_  = ~A266 & A265;
  assign \new_[8582]_  = A268 & A267;
  assign \new_[8583]_  = \new_[8582]_  & \new_[8579]_ ;
  assign \new_[8584]_  = \new_[8583]_  & \new_[8576]_ ;
  assign \new_[8588]_  = A167 & A169;
  assign \new_[8589]_  = ~A170 & \new_[8588]_ ;
  assign \new_[8592]_  = ~A199 & A166;
  assign \new_[8595]_  = A232 & ~A200;
  assign \new_[8596]_  = \new_[8595]_  & \new_[8592]_ ;
  assign \new_[8597]_  = \new_[8596]_  & \new_[8589]_ ;
  assign \new_[8601]_  = A236 & A234;
  assign \new_[8602]_  = ~A233 & \new_[8601]_ ;
  assign \new_[8605]_  = ~A266 & A265;
  assign \new_[8608]_  = A269 & A267;
  assign \new_[8609]_  = \new_[8608]_  & \new_[8605]_ ;
  assign \new_[8610]_  = \new_[8609]_  & \new_[8602]_ ;
  assign \new_[8614]_  = ~A167 & A169;
  assign \new_[8615]_  = ~A170 & \new_[8614]_ ;
  assign \new_[8618]_  = A199 & ~A166;
  assign \new_[8621]_  = A232 & ~A201;
  assign \new_[8622]_  = \new_[8621]_  & \new_[8618]_ ;
  assign \new_[8623]_  = \new_[8622]_  & \new_[8615]_ ;
  assign \new_[8627]_  = A235 & A234;
  assign \new_[8628]_  = ~A233 & \new_[8627]_ ;
  assign \new_[8631]_  = ~A299 & A298;
  assign \new_[8634]_  = A301 & A300;
  assign \new_[8635]_  = \new_[8634]_  & \new_[8631]_ ;
  assign \new_[8636]_  = \new_[8635]_  & \new_[8628]_ ;
  assign \new_[8640]_  = ~A167 & A169;
  assign \new_[8641]_  = ~A170 & \new_[8640]_ ;
  assign \new_[8644]_  = A199 & ~A166;
  assign \new_[8647]_  = A232 & ~A201;
  assign \new_[8648]_  = \new_[8647]_  & \new_[8644]_ ;
  assign \new_[8649]_  = \new_[8648]_  & \new_[8641]_ ;
  assign \new_[8653]_  = A235 & A234;
  assign \new_[8654]_  = ~A233 & \new_[8653]_ ;
  assign \new_[8657]_  = ~A299 & A298;
  assign \new_[8660]_  = A302 & A300;
  assign \new_[8661]_  = \new_[8660]_  & \new_[8657]_ ;
  assign \new_[8662]_  = \new_[8661]_  & \new_[8654]_ ;
  assign \new_[8666]_  = ~A167 & A169;
  assign \new_[8667]_  = ~A170 & \new_[8666]_ ;
  assign \new_[8670]_  = A199 & ~A166;
  assign \new_[8673]_  = A232 & ~A201;
  assign \new_[8674]_  = \new_[8673]_  & \new_[8670]_ ;
  assign \new_[8675]_  = \new_[8674]_  & \new_[8667]_ ;
  assign \new_[8679]_  = A235 & A234;
  assign \new_[8680]_  = ~A233 & \new_[8679]_ ;
  assign \new_[8683]_  = ~A266 & A265;
  assign \new_[8686]_  = A268 & A267;
  assign \new_[8687]_  = \new_[8686]_  & \new_[8683]_ ;
  assign \new_[8688]_  = \new_[8687]_  & \new_[8680]_ ;
  assign \new_[8692]_  = ~A167 & A169;
  assign \new_[8693]_  = ~A170 & \new_[8692]_ ;
  assign \new_[8696]_  = A199 & ~A166;
  assign \new_[8699]_  = A232 & ~A201;
  assign \new_[8700]_  = \new_[8699]_  & \new_[8696]_ ;
  assign \new_[8701]_  = \new_[8700]_  & \new_[8693]_ ;
  assign \new_[8705]_  = A235 & A234;
  assign \new_[8706]_  = ~A233 & \new_[8705]_ ;
  assign \new_[8709]_  = ~A266 & A265;
  assign \new_[8712]_  = A269 & A267;
  assign \new_[8713]_  = \new_[8712]_  & \new_[8709]_ ;
  assign \new_[8714]_  = \new_[8713]_  & \new_[8706]_ ;
  assign \new_[8718]_  = ~A167 & A169;
  assign \new_[8719]_  = ~A170 & \new_[8718]_ ;
  assign \new_[8722]_  = A199 & ~A166;
  assign \new_[8725]_  = A232 & ~A201;
  assign \new_[8726]_  = \new_[8725]_  & \new_[8722]_ ;
  assign \new_[8727]_  = \new_[8726]_  & \new_[8719]_ ;
  assign \new_[8731]_  = A236 & A234;
  assign \new_[8732]_  = ~A233 & \new_[8731]_ ;
  assign \new_[8735]_  = ~A299 & A298;
  assign \new_[8738]_  = A301 & A300;
  assign \new_[8739]_  = \new_[8738]_  & \new_[8735]_ ;
  assign \new_[8740]_  = \new_[8739]_  & \new_[8732]_ ;
  assign \new_[8744]_  = ~A167 & A169;
  assign \new_[8745]_  = ~A170 & \new_[8744]_ ;
  assign \new_[8748]_  = A199 & ~A166;
  assign \new_[8751]_  = A232 & ~A201;
  assign \new_[8752]_  = \new_[8751]_  & \new_[8748]_ ;
  assign \new_[8753]_  = \new_[8752]_  & \new_[8745]_ ;
  assign \new_[8757]_  = A236 & A234;
  assign \new_[8758]_  = ~A233 & \new_[8757]_ ;
  assign \new_[8761]_  = ~A299 & A298;
  assign \new_[8764]_  = A302 & A300;
  assign \new_[8765]_  = \new_[8764]_  & \new_[8761]_ ;
  assign \new_[8766]_  = \new_[8765]_  & \new_[8758]_ ;
  assign \new_[8770]_  = ~A167 & A169;
  assign \new_[8771]_  = ~A170 & \new_[8770]_ ;
  assign \new_[8774]_  = A199 & ~A166;
  assign \new_[8777]_  = A232 & ~A201;
  assign \new_[8778]_  = \new_[8777]_  & \new_[8774]_ ;
  assign \new_[8779]_  = \new_[8778]_  & \new_[8771]_ ;
  assign \new_[8783]_  = A236 & A234;
  assign \new_[8784]_  = ~A233 & \new_[8783]_ ;
  assign \new_[8787]_  = ~A266 & A265;
  assign \new_[8790]_  = A268 & A267;
  assign \new_[8791]_  = \new_[8790]_  & \new_[8787]_ ;
  assign \new_[8792]_  = \new_[8791]_  & \new_[8784]_ ;
  assign \new_[8796]_  = ~A167 & A169;
  assign \new_[8797]_  = ~A170 & \new_[8796]_ ;
  assign \new_[8800]_  = A199 & ~A166;
  assign \new_[8803]_  = A232 & ~A201;
  assign \new_[8804]_  = \new_[8803]_  & \new_[8800]_ ;
  assign \new_[8805]_  = \new_[8804]_  & \new_[8797]_ ;
  assign \new_[8809]_  = A236 & A234;
  assign \new_[8810]_  = ~A233 & \new_[8809]_ ;
  assign \new_[8813]_  = ~A266 & A265;
  assign \new_[8816]_  = A269 & A267;
  assign \new_[8817]_  = \new_[8816]_  & \new_[8813]_ ;
  assign \new_[8818]_  = \new_[8817]_  & \new_[8810]_ ;
  assign \new_[8822]_  = ~A167 & A169;
  assign \new_[8823]_  = ~A170 & \new_[8822]_ ;
  assign \new_[8826]_  = A199 & ~A166;
  assign \new_[8829]_  = A232 & A200;
  assign \new_[8830]_  = \new_[8829]_  & \new_[8826]_ ;
  assign \new_[8831]_  = \new_[8830]_  & \new_[8823]_ ;
  assign \new_[8835]_  = A235 & A234;
  assign \new_[8836]_  = ~A233 & \new_[8835]_ ;
  assign \new_[8839]_  = ~A299 & A298;
  assign \new_[8842]_  = A301 & A300;
  assign \new_[8843]_  = \new_[8842]_  & \new_[8839]_ ;
  assign \new_[8844]_  = \new_[8843]_  & \new_[8836]_ ;
  assign \new_[8848]_  = ~A167 & A169;
  assign \new_[8849]_  = ~A170 & \new_[8848]_ ;
  assign \new_[8852]_  = A199 & ~A166;
  assign \new_[8855]_  = A232 & A200;
  assign \new_[8856]_  = \new_[8855]_  & \new_[8852]_ ;
  assign \new_[8857]_  = \new_[8856]_  & \new_[8849]_ ;
  assign \new_[8861]_  = A235 & A234;
  assign \new_[8862]_  = ~A233 & \new_[8861]_ ;
  assign \new_[8865]_  = ~A299 & A298;
  assign \new_[8868]_  = A302 & A300;
  assign \new_[8869]_  = \new_[8868]_  & \new_[8865]_ ;
  assign \new_[8870]_  = \new_[8869]_  & \new_[8862]_ ;
  assign \new_[8874]_  = ~A167 & A169;
  assign \new_[8875]_  = ~A170 & \new_[8874]_ ;
  assign \new_[8878]_  = A199 & ~A166;
  assign \new_[8881]_  = A232 & A200;
  assign \new_[8882]_  = \new_[8881]_  & \new_[8878]_ ;
  assign \new_[8883]_  = \new_[8882]_  & \new_[8875]_ ;
  assign \new_[8887]_  = A235 & A234;
  assign \new_[8888]_  = ~A233 & \new_[8887]_ ;
  assign \new_[8891]_  = ~A266 & A265;
  assign \new_[8894]_  = A268 & A267;
  assign \new_[8895]_  = \new_[8894]_  & \new_[8891]_ ;
  assign \new_[8896]_  = \new_[8895]_  & \new_[8888]_ ;
  assign \new_[8900]_  = ~A167 & A169;
  assign \new_[8901]_  = ~A170 & \new_[8900]_ ;
  assign \new_[8904]_  = A199 & ~A166;
  assign \new_[8907]_  = A232 & A200;
  assign \new_[8908]_  = \new_[8907]_  & \new_[8904]_ ;
  assign \new_[8909]_  = \new_[8908]_  & \new_[8901]_ ;
  assign \new_[8913]_  = A235 & A234;
  assign \new_[8914]_  = ~A233 & \new_[8913]_ ;
  assign \new_[8917]_  = ~A266 & A265;
  assign \new_[8920]_  = A269 & A267;
  assign \new_[8921]_  = \new_[8920]_  & \new_[8917]_ ;
  assign \new_[8922]_  = \new_[8921]_  & \new_[8914]_ ;
  assign \new_[8926]_  = ~A167 & A169;
  assign \new_[8927]_  = ~A170 & \new_[8926]_ ;
  assign \new_[8930]_  = A199 & ~A166;
  assign \new_[8933]_  = A232 & A200;
  assign \new_[8934]_  = \new_[8933]_  & \new_[8930]_ ;
  assign \new_[8935]_  = \new_[8934]_  & \new_[8927]_ ;
  assign \new_[8939]_  = A236 & A234;
  assign \new_[8940]_  = ~A233 & \new_[8939]_ ;
  assign \new_[8943]_  = ~A299 & A298;
  assign \new_[8946]_  = A301 & A300;
  assign \new_[8947]_  = \new_[8946]_  & \new_[8943]_ ;
  assign \new_[8948]_  = \new_[8947]_  & \new_[8940]_ ;
  assign \new_[8952]_  = ~A167 & A169;
  assign \new_[8953]_  = ~A170 & \new_[8952]_ ;
  assign \new_[8956]_  = A199 & ~A166;
  assign \new_[8959]_  = A232 & A200;
  assign \new_[8960]_  = \new_[8959]_  & \new_[8956]_ ;
  assign \new_[8961]_  = \new_[8960]_  & \new_[8953]_ ;
  assign \new_[8965]_  = A236 & A234;
  assign \new_[8966]_  = ~A233 & \new_[8965]_ ;
  assign \new_[8969]_  = ~A299 & A298;
  assign \new_[8972]_  = A302 & A300;
  assign \new_[8973]_  = \new_[8972]_  & \new_[8969]_ ;
  assign \new_[8974]_  = \new_[8973]_  & \new_[8966]_ ;
  assign \new_[8978]_  = ~A167 & A169;
  assign \new_[8979]_  = ~A170 & \new_[8978]_ ;
  assign \new_[8982]_  = A199 & ~A166;
  assign \new_[8985]_  = A232 & A200;
  assign \new_[8986]_  = \new_[8985]_  & \new_[8982]_ ;
  assign \new_[8987]_  = \new_[8986]_  & \new_[8979]_ ;
  assign \new_[8991]_  = A236 & A234;
  assign \new_[8992]_  = ~A233 & \new_[8991]_ ;
  assign \new_[8995]_  = ~A266 & A265;
  assign \new_[8998]_  = A268 & A267;
  assign \new_[8999]_  = \new_[8998]_  & \new_[8995]_ ;
  assign \new_[9000]_  = \new_[8999]_  & \new_[8992]_ ;
  assign \new_[9004]_  = ~A167 & A169;
  assign \new_[9005]_  = ~A170 & \new_[9004]_ ;
  assign \new_[9008]_  = A199 & ~A166;
  assign \new_[9011]_  = A232 & A200;
  assign \new_[9012]_  = \new_[9011]_  & \new_[9008]_ ;
  assign \new_[9013]_  = \new_[9012]_  & \new_[9005]_ ;
  assign \new_[9017]_  = A236 & A234;
  assign \new_[9018]_  = ~A233 & \new_[9017]_ ;
  assign \new_[9021]_  = ~A266 & A265;
  assign \new_[9024]_  = A269 & A267;
  assign \new_[9025]_  = \new_[9024]_  & \new_[9021]_ ;
  assign \new_[9026]_  = \new_[9025]_  & \new_[9018]_ ;
  assign \new_[9030]_  = ~A167 & A169;
  assign \new_[9031]_  = ~A170 & \new_[9030]_ ;
  assign \new_[9034]_  = ~A199 & ~A166;
  assign \new_[9037]_  = A232 & ~A200;
  assign \new_[9038]_  = \new_[9037]_  & \new_[9034]_ ;
  assign \new_[9039]_  = \new_[9038]_  & \new_[9031]_ ;
  assign \new_[9043]_  = A235 & A234;
  assign \new_[9044]_  = ~A233 & \new_[9043]_ ;
  assign \new_[9047]_  = ~A299 & A298;
  assign \new_[9050]_  = A301 & A300;
  assign \new_[9051]_  = \new_[9050]_  & \new_[9047]_ ;
  assign \new_[9052]_  = \new_[9051]_  & \new_[9044]_ ;
  assign \new_[9056]_  = ~A167 & A169;
  assign \new_[9057]_  = ~A170 & \new_[9056]_ ;
  assign \new_[9060]_  = ~A199 & ~A166;
  assign \new_[9063]_  = A232 & ~A200;
  assign \new_[9064]_  = \new_[9063]_  & \new_[9060]_ ;
  assign \new_[9065]_  = \new_[9064]_  & \new_[9057]_ ;
  assign \new_[9069]_  = A235 & A234;
  assign \new_[9070]_  = ~A233 & \new_[9069]_ ;
  assign \new_[9073]_  = ~A299 & A298;
  assign \new_[9076]_  = A302 & A300;
  assign \new_[9077]_  = \new_[9076]_  & \new_[9073]_ ;
  assign \new_[9078]_  = \new_[9077]_  & \new_[9070]_ ;
  assign \new_[9082]_  = ~A167 & A169;
  assign \new_[9083]_  = ~A170 & \new_[9082]_ ;
  assign \new_[9086]_  = ~A199 & ~A166;
  assign \new_[9089]_  = A232 & ~A200;
  assign \new_[9090]_  = \new_[9089]_  & \new_[9086]_ ;
  assign \new_[9091]_  = \new_[9090]_  & \new_[9083]_ ;
  assign \new_[9095]_  = A235 & A234;
  assign \new_[9096]_  = ~A233 & \new_[9095]_ ;
  assign \new_[9099]_  = ~A266 & A265;
  assign \new_[9102]_  = A268 & A267;
  assign \new_[9103]_  = \new_[9102]_  & \new_[9099]_ ;
  assign \new_[9104]_  = \new_[9103]_  & \new_[9096]_ ;
  assign \new_[9108]_  = ~A167 & A169;
  assign \new_[9109]_  = ~A170 & \new_[9108]_ ;
  assign \new_[9112]_  = ~A199 & ~A166;
  assign \new_[9115]_  = A232 & ~A200;
  assign \new_[9116]_  = \new_[9115]_  & \new_[9112]_ ;
  assign \new_[9117]_  = \new_[9116]_  & \new_[9109]_ ;
  assign \new_[9121]_  = A235 & A234;
  assign \new_[9122]_  = ~A233 & \new_[9121]_ ;
  assign \new_[9125]_  = ~A266 & A265;
  assign \new_[9128]_  = A269 & A267;
  assign \new_[9129]_  = \new_[9128]_  & \new_[9125]_ ;
  assign \new_[9130]_  = \new_[9129]_  & \new_[9122]_ ;
  assign \new_[9134]_  = ~A167 & A169;
  assign \new_[9135]_  = ~A170 & \new_[9134]_ ;
  assign \new_[9138]_  = ~A199 & ~A166;
  assign \new_[9141]_  = A232 & ~A200;
  assign \new_[9142]_  = \new_[9141]_  & \new_[9138]_ ;
  assign \new_[9143]_  = \new_[9142]_  & \new_[9135]_ ;
  assign \new_[9147]_  = A236 & A234;
  assign \new_[9148]_  = ~A233 & \new_[9147]_ ;
  assign \new_[9151]_  = ~A299 & A298;
  assign \new_[9154]_  = A301 & A300;
  assign \new_[9155]_  = \new_[9154]_  & \new_[9151]_ ;
  assign \new_[9156]_  = \new_[9155]_  & \new_[9148]_ ;
  assign \new_[9160]_  = ~A167 & A169;
  assign \new_[9161]_  = ~A170 & \new_[9160]_ ;
  assign \new_[9164]_  = ~A199 & ~A166;
  assign \new_[9167]_  = A232 & ~A200;
  assign \new_[9168]_  = \new_[9167]_  & \new_[9164]_ ;
  assign \new_[9169]_  = \new_[9168]_  & \new_[9161]_ ;
  assign \new_[9173]_  = A236 & A234;
  assign \new_[9174]_  = ~A233 & \new_[9173]_ ;
  assign \new_[9177]_  = ~A299 & A298;
  assign \new_[9180]_  = A302 & A300;
  assign \new_[9181]_  = \new_[9180]_  & \new_[9177]_ ;
  assign \new_[9182]_  = \new_[9181]_  & \new_[9174]_ ;
  assign \new_[9186]_  = ~A167 & A169;
  assign \new_[9187]_  = ~A170 & \new_[9186]_ ;
  assign \new_[9190]_  = ~A199 & ~A166;
  assign \new_[9193]_  = A232 & ~A200;
  assign \new_[9194]_  = \new_[9193]_  & \new_[9190]_ ;
  assign \new_[9195]_  = \new_[9194]_  & \new_[9187]_ ;
  assign \new_[9199]_  = A236 & A234;
  assign \new_[9200]_  = ~A233 & \new_[9199]_ ;
  assign \new_[9203]_  = ~A266 & A265;
  assign \new_[9206]_  = A268 & A267;
  assign \new_[9207]_  = \new_[9206]_  & \new_[9203]_ ;
  assign \new_[9208]_  = \new_[9207]_  & \new_[9200]_ ;
  assign \new_[9212]_  = ~A167 & A169;
  assign \new_[9213]_  = ~A170 & \new_[9212]_ ;
  assign \new_[9216]_  = ~A199 & ~A166;
  assign \new_[9219]_  = A232 & ~A200;
  assign \new_[9220]_  = \new_[9219]_  & \new_[9216]_ ;
  assign \new_[9221]_  = \new_[9220]_  & \new_[9213]_ ;
  assign \new_[9225]_  = A236 & A234;
  assign \new_[9226]_  = ~A233 & \new_[9225]_ ;
  assign \new_[9229]_  = ~A266 & A265;
  assign \new_[9232]_  = A269 & A267;
  assign \new_[9233]_  = \new_[9232]_  & \new_[9229]_ ;
  assign \new_[9234]_  = \new_[9233]_  & \new_[9226]_ ;
  assign \new_[9238]_  = A167 & ~A169;
  assign \new_[9239]_  = A170 & \new_[9238]_ ;
  assign \new_[9242]_  = A199 & ~A166;
  assign \new_[9245]_  = A232 & ~A201;
  assign \new_[9246]_  = \new_[9245]_  & \new_[9242]_ ;
  assign \new_[9247]_  = \new_[9246]_  & \new_[9239]_ ;
  assign \new_[9251]_  = A235 & A234;
  assign \new_[9252]_  = ~A233 & \new_[9251]_ ;
  assign \new_[9255]_  = ~A299 & A298;
  assign \new_[9258]_  = A301 & A300;
  assign \new_[9259]_  = \new_[9258]_  & \new_[9255]_ ;
  assign \new_[9260]_  = \new_[9259]_  & \new_[9252]_ ;
  assign \new_[9264]_  = A167 & ~A169;
  assign \new_[9265]_  = A170 & \new_[9264]_ ;
  assign \new_[9268]_  = A199 & ~A166;
  assign \new_[9271]_  = A232 & ~A201;
  assign \new_[9272]_  = \new_[9271]_  & \new_[9268]_ ;
  assign \new_[9273]_  = \new_[9272]_  & \new_[9265]_ ;
  assign \new_[9277]_  = A235 & A234;
  assign \new_[9278]_  = ~A233 & \new_[9277]_ ;
  assign \new_[9281]_  = ~A299 & A298;
  assign \new_[9284]_  = A302 & A300;
  assign \new_[9285]_  = \new_[9284]_  & \new_[9281]_ ;
  assign \new_[9286]_  = \new_[9285]_  & \new_[9278]_ ;
  assign \new_[9290]_  = A167 & ~A169;
  assign \new_[9291]_  = A170 & \new_[9290]_ ;
  assign \new_[9294]_  = A199 & ~A166;
  assign \new_[9297]_  = A232 & ~A201;
  assign \new_[9298]_  = \new_[9297]_  & \new_[9294]_ ;
  assign \new_[9299]_  = \new_[9298]_  & \new_[9291]_ ;
  assign \new_[9303]_  = A235 & A234;
  assign \new_[9304]_  = ~A233 & \new_[9303]_ ;
  assign \new_[9307]_  = ~A266 & A265;
  assign \new_[9310]_  = A268 & A267;
  assign \new_[9311]_  = \new_[9310]_  & \new_[9307]_ ;
  assign \new_[9312]_  = \new_[9311]_  & \new_[9304]_ ;
  assign \new_[9316]_  = A167 & ~A169;
  assign \new_[9317]_  = A170 & \new_[9316]_ ;
  assign \new_[9320]_  = A199 & ~A166;
  assign \new_[9323]_  = A232 & ~A201;
  assign \new_[9324]_  = \new_[9323]_  & \new_[9320]_ ;
  assign \new_[9325]_  = \new_[9324]_  & \new_[9317]_ ;
  assign \new_[9329]_  = A235 & A234;
  assign \new_[9330]_  = ~A233 & \new_[9329]_ ;
  assign \new_[9333]_  = ~A266 & A265;
  assign \new_[9336]_  = A269 & A267;
  assign \new_[9337]_  = \new_[9336]_  & \new_[9333]_ ;
  assign \new_[9338]_  = \new_[9337]_  & \new_[9330]_ ;
  assign \new_[9342]_  = A167 & ~A169;
  assign \new_[9343]_  = A170 & \new_[9342]_ ;
  assign \new_[9346]_  = A199 & ~A166;
  assign \new_[9349]_  = A232 & ~A201;
  assign \new_[9350]_  = \new_[9349]_  & \new_[9346]_ ;
  assign \new_[9351]_  = \new_[9350]_  & \new_[9343]_ ;
  assign \new_[9355]_  = A236 & A234;
  assign \new_[9356]_  = ~A233 & \new_[9355]_ ;
  assign \new_[9359]_  = ~A299 & A298;
  assign \new_[9362]_  = A301 & A300;
  assign \new_[9363]_  = \new_[9362]_  & \new_[9359]_ ;
  assign \new_[9364]_  = \new_[9363]_  & \new_[9356]_ ;
  assign \new_[9368]_  = A167 & ~A169;
  assign \new_[9369]_  = A170 & \new_[9368]_ ;
  assign \new_[9372]_  = A199 & ~A166;
  assign \new_[9375]_  = A232 & ~A201;
  assign \new_[9376]_  = \new_[9375]_  & \new_[9372]_ ;
  assign \new_[9377]_  = \new_[9376]_  & \new_[9369]_ ;
  assign \new_[9381]_  = A236 & A234;
  assign \new_[9382]_  = ~A233 & \new_[9381]_ ;
  assign \new_[9385]_  = ~A299 & A298;
  assign \new_[9388]_  = A302 & A300;
  assign \new_[9389]_  = \new_[9388]_  & \new_[9385]_ ;
  assign \new_[9390]_  = \new_[9389]_  & \new_[9382]_ ;
  assign \new_[9394]_  = A167 & ~A169;
  assign \new_[9395]_  = A170 & \new_[9394]_ ;
  assign \new_[9398]_  = A199 & ~A166;
  assign \new_[9401]_  = A232 & ~A201;
  assign \new_[9402]_  = \new_[9401]_  & \new_[9398]_ ;
  assign \new_[9403]_  = \new_[9402]_  & \new_[9395]_ ;
  assign \new_[9407]_  = A236 & A234;
  assign \new_[9408]_  = ~A233 & \new_[9407]_ ;
  assign \new_[9411]_  = ~A266 & A265;
  assign \new_[9414]_  = A268 & A267;
  assign \new_[9415]_  = \new_[9414]_  & \new_[9411]_ ;
  assign \new_[9416]_  = \new_[9415]_  & \new_[9408]_ ;
  assign \new_[9420]_  = A167 & ~A169;
  assign \new_[9421]_  = A170 & \new_[9420]_ ;
  assign \new_[9424]_  = A199 & ~A166;
  assign \new_[9427]_  = A232 & ~A201;
  assign \new_[9428]_  = \new_[9427]_  & \new_[9424]_ ;
  assign \new_[9429]_  = \new_[9428]_  & \new_[9421]_ ;
  assign \new_[9433]_  = A236 & A234;
  assign \new_[9434]_  = ~A233 & \new_[9433]_ ;
  assign \new_[9437]_  = ~A266 & A265;
  assign \new_[9440]_  = A269 & A267;
  assign \new_[9441]_  = \new_[9440]_  & \new_[9437]_ ;
  assign \new_[9442]_  = \new_[9441]_  & \new_[9434]_ ;
  assign \new_[9446]_  = A167 & ~A169;
  assign \new_[9447]_  = A170 & \new_[9446]_ ;
  assign \new_[9450]_  = A199 & ~A166;
  assign \new_[9453]_  = A232 & A200;
  assign \new_[9454]_  = \new_[9453]_  & \new_[9450]_ ;
  assign \new_[9455]_  = \new_[9454]_  & \new_[9447]_ ;
  assign \new_[9459]_  = A235 & A234;
  assign \new_[9460]_  = ~A233 & \new_[9459]_ ;
  assign \new_[9463]_  = ~A299 & A298;
  assign \new_[9466]_  = A301 & A300;
  assign \new_[9467]_  = \new_[9466]_  & \new_[9463]_ ;
  assign \new_[9468]_  = \new_[9467]_  & \new_[9460]_ ;
  assign \new_[9472]_  = A167 & ~A169;
  assign \new_[9473]_  = A170 & \new_[9472]_ ;
  assign \new_[9476]_  = A199 & ~A166;
  assign \new_[9479]_  = A232 & A200;
  assign \new_[9480]_  = \new_[9479]_  & \new_[9476]_ ;
  assign \new_[9481]_  = \new_[9480]_  & \new_[9473]_ ;
  assign \new_[9485]_  = A235 & A234;
  assign \new_[9486]_  = ~A233 & \new_[9485]_ ;
  assign \new_[9489]_  = ~A299 & A298;
  assign \new_[9492]_  = A302 & A300;
  assign \new_[9493]_  = \new_[9492]_  & \new_[9489]_ ;
  assign \new_[9494]_  = \new_[9493]_  & \new_[9486]_ ;
  assign \new_[9498]_  = A167 & ~A169;
  assign \new_[9499]_  = A170 & \new_[9498]_ ;
  assign \new_[9502]_  = A199 & ~A166;
  assign \new_[9505]_  = A232 & A200;
  assign \new_[9506]_  = \new_[9505]_  & \new_[9502]_ ;
  assign \new_[9507]_  = \new_[9506]_  & \new_[9499]_ ;
  assign \new_[9511]_  = A235 & A234;
  assign \new_[9512]_  = ~A233 & \new_[9511]_ ;
  assign \new_[9515]_  = ~A266 & A265;
  assign \new_[9518]_  = A268 & A267;
  assign \new_[9519]_  = \new_[9518]_  & \new_[9515]_ ;
  assign \new_[9520]_  = \new_[9519]_  & \new_[9512]_ ;
  assign \new_[9524]_  = A167 & ~A169;
  assign \new_[9525]_  = A170 & \new_[9524]_ ;
  assign \new_[9528]_  = A199 & ~A166;
  assign \new_[9531]_  = A232 & A200;
  assign \new_[9532]_  = \new_[9531]_  & \new_[9528]_ ;
  assign \new_[9533]_  = \new_[9532]_  & \new_[9525]_ ;
  assign \new_[9537]_  = A235 & A234;
  assign \new_[9538]_  = ~A233 & \new_[9537]_ ;
  assign \new_[9541]_  = ~A266 & A265;
  assign \new_[9544]_  = A269 & A267;
  assign \new_[9545]_  = \new_[9544]_  & \new_[9541]_ ;
  assign \new_[9546]_  = \new_[9545]_  & \new_[9538]_ ;
  assign \new_[9550]_  = A167 & ~A169;
  assign \new_[9551]_  = A170 & \new_[9550]_ ;
  assign \new_[9554]_  = A199 & ~A166;
  assign \new_[9557]_  = A232 & A200;
  assign \new_[9558]_  = \new_[9557]_  & \new_[9554]_ ;
  assign \new_[9559]_  = \new_[9558]_  & \new_[9551]_ ;
  assign \new_[9563]_  = A236 & A234;
  assign \new_[9564]_  = ~A233 & \new_[9563]_ ;
  assign \new_[9567]_  = ~A299 & A298;
  assign \new_[9570]_  = A301 & A300;
  assign \new_[9571]_  = \new_[9570]_  & \new_[9567]_ ;
  assign \new_[9572]_  = \new_[9571]_  & \new_[9564]_ ;
  assign \new_[9576]_  = A167 & ~A169;
  assign \new_[9577]_  = A170 & \new_[9576]_ ;
  assign \new_[9580]_  = A199 & ~A166;
  assign \new_[9583]_  = A232 & A200;
  assign \new_[9584]_  = \new_[9583]_  & \new_[9580]_ ;
  assign \new_[9585]_  = \new_[9584]_  & \new_[9577]_ ;
  assign \new_[9589]_  = A236 & A234;
  assign \new_[9590]_  = ~A233 & \new_[9589]_ ;
  assign \new_[9593]_  = ~A299 & A298;
  assign \new_[9596]_  = A302 & A300;
  assign \new_[9597]_  = \new_[9596]_  & \new_[9593]_ ;
  assign \new_[9598]_  = \new_[9597]_  & \new_[9590]_ ;
  assign \new_[9602]_  = A167 & ~A169;
  assign \new_[9603]_  = A170 & \new_[9602]_ ;
  assign \new_[9606]_  = A199 & ~A166;
  assign \new_[9609]_  = A232 & A200;
  assign \new_[9610]_  = \new_[9609]_  & \new_[9606]_ ;
  assign \new_[9611]_  = \new_[9610]_  & \new_[9603]_ ;
  assign \new_[9615]_  = A236 & A234;
  assign \new_[9616]_  = ~A233 & \new_[9615]_ ;
  assign \new_[9619]_  = ~A266 & A265;
  assign \new_[9622]_  = A268 & A267;
  assign \new_[9623]_  = \new_[9622]_  & \new_[9619]_ ;
  assign \new_[9624]_  = \new_[9623]_  & \new_[9616]_ ;
  assign \new_[9628]_  = A167 & ~A169;
  assign \new_[9629]_  = A170 & \new_[9628]_ ;
  assign \new_[9632]_  = A199 & ~A166;
  assign \new_[9635]_  = A232 & A200;
  assign \new_[9636]_  = \new_[9635]_  & \new_[9632]_ ;
  assign \new_[9637]_  = \new_[9636]_  & \new_[9629]_ ;
  assign \new_[9641]_  = A236 & A234;
  assign \new_[9642]_  = ~A233 & \new_[9641]_ ;
  assign \new_[9645]_  = ~A266 & A265;
  assign \new_[9648]_  = A269 & A267;
  assign \new_[9649]_  = \new_[9648]_  & \new_[9645]_ ;
  assign \new_[9650]_  = \new_[9649]_  & \new_[9642]_ ;
  assign \new_[9654]_  = A167 & ~A169;
  assign \new_[9655]_  = A170 & \new_[9654]_ ;
  assign \new_[9658]_  = ~A199 & ~A166;
  assign \new_[9661]_  = A232 & ~A200;
  assign \new_[9662]_  = \new_[9661]_  & \new_[9658]_ ;
  assign \new_[9663]_  = \new_[9662]_  & \new_[9655]_ ;
  assign \new_[9667]_  = A235 & A234;
  assign \new_[9668]_  = ~A233 & \new_[9667]_ ;
  assign \new_[9671]_  = ~A299 & A298;
  assign \new_[9674]_  = A301 & A300;
  assign \new_[9675]_  = \new_[9674]_  & \new_[9671]_ ;
  assign \new_[9676]_  = \new_[9675]_  & \new_[9668]_ ;
  assign \new_[9680]_  = A167 & ~A169;
  assign \new_[9681]_  = A170 & \new_[9680]_ ;
  assign \new_[9684]_  = ~A199 & ~A166;
  assign \new_[9687]_  = A232 & ~A200;
  assign \new_[9688]_  = \new_[9687]_  & \new_[9684]_ ;
  assign \new_[9689]_  = \new_[9688]_  & \new_[9681]_ ;
  assign \new_[9693]_  = A235 & A234;
  assign \new_[9694]_  = ~A233 & \new_[9693]_ ;
  assign \new_[9697]_  = ~A299 & A298;
  assign \new_[9700]_  = A302 & A300;
  assign \new_[9701]_  = \new_[9700]_  & \new_[9697]_ ;
  assign \new_[9702]_  = \new_[9701]_  & \new_[9694]_ ;
  assign \new_[9706]_  = A167 & ~A169;
  assign \new_[9707]_  = A170 & \new_[9706]_ ;
  assign \new_[9710]_  = ~A199 & ~A166;
  assign \new_[9713]_  = A232 & ~A200;
  assign \new_[9714]_  = \new_[9713]_  & \new_[9710]_ ;
  assign \new_[9715]_  = \new_[9714]_  & \new_[9707]_ ;
  assign \new_[9719]_  = A235 & A234;
  assign \new_[9720]_  = ~A233 & \new_[9719]_ ;
  assign \new_[9723]_  = ~A266 & A265;
  assign \new_[9726]_  = A268 & A267;
  assign \new_[9727]_  = \new_[9726]_  & \new_[9723]_ ;
  assign \new_[9728]_  = \new_[9727]_  & \new_[9720]_ ;
  assign \new_[9732]_  = A167 & ~A169;
  assign \new_[9733]_  = A170 & \new_[9732]_ ;
  assign \new_[9736]_  = ~A199 & ~A166;
  assign \new_[9739]_  = A232 & ~A200;
  assign \new_[9740]_  = \new_[9739]_  & \new_[9736]_ ;
  assign \new_[9741]_  = \new_[9740]_  & \new_[9733]_ ;
  assign \new_[9745]_  = A235 & A234;
  assign \new_[9746]_  = ~A233 & \new_[9745]_ ;
  assign \new_[9749]_  = ~A266 & A265;
  assign \new_[9752]_  = A269 & A267;
  assign \new_[9753]_  = \new_[9752]_  & \new_[9749]_ ;
  assign \new_[9754]_  = \new_[9753]_  & \new_[9746]_ ;
  assign \new_[9758]_  = A167 & ~A169;
  assign \new_[9759]_  = A170 & \new_[9758]_ ;
  assign \new_[9762]_  = ~A199 & ~A166;
  assign \new_[9765]_  = A232 & ~A200;
  assign \new_[9766]_  = \new_[9765]_  & \new_[9762]_ ;
  assign \new_[9767]_  = \new_[9766]_  & \new_[9759]_ ;
  assign \new_[9771]_  = A236 & A234;
  assign \new_[9772]_  = ~A233 & \new_[9771]_ ;
  assign \new_[9775]_  = ~A299 & A298;
  assign \new_[9778]_  = A301 & A300;
  assign \new_[9779]_  = \new_[9778]_  & \new_[9775]_ ;
  assign \new_[9780]_  = \new_[9779]_  & \new_[9772]_ ;
  assign \new_[9784]_  = A167 & ~A169;
  assign \new_[9785]_  = A170 & \new_[9784]_ ;
  assign \new_[9788]_  = ~A199 & ~A166;
  assign \new_[9791]_  = A232 & ~A200;
  assign \new_[9792]_  = \new_[9791]_  & \new_[9788]_ ;
  assign \new_[9793]_  = \new_[9792]_  & \new_[9785]_ ;
  assign \new_[9797]_  = A236 & A234;
  assign \new_[9798]_  = ~A233 & \new_[9797]_ ;
  assign \new_[9801]_  = ~A299 & A298;
  assign \new_[9804]_  = A302 & A300;
  assign \new_[9805]_  = \new_[9804]_  & \new_[9801]_ ;
  assign \new_[9806]_  = \new_[9805]_  & \new_[9798]_ ;
  assign \new_[9810]_  = A167 & ~A169;
  assign \new_[9811]_  = A170 & \new_[9810]_ ;
  assign \new_[9814]_  = ~A199 & ~A166;
  assign \new_[9817]_  = A232 & ~A200;
  assign \new_[9818]_  = \new_[9817]_  & \new_[9814]_ ;
  assign \new_[9819]_  = \new_[9818]_  & \new_[9811]_ ;
  assign \new_[9823]_  = A236 & A234;
  assign \new_[9824]_  = ~A233 & \new_[9823]_ ;
  assign \new_[9827]_  = ~A266 & A265;
  assign \new_[9830]_  = A268 & A267;
  assign \new_[9831]_  = \new_[9830]_  & \new_[9827]_ ;
  assign \new_[9832]_  = \new_[9831]_  & \new_[9824]_ ;
  assign \new_[9836]_  = A167 & ~A169;
  assign \new_[9837]_  = A170 & \new_[9836]_ ;
  assign \new_[9840]_  = ~A199 & ~A166;
  assign \new_[9843]_  = A232 & ~A200;
  assign \new_[9844]_  = \new_[9843]_  & \new_[9840]_ ;
  assign \new_[9845]_  = \new_[9844]_  & \new_[9837]_ ;
  assign \new_[9849]_  = A236 & A234;
  assign \new_[9850]_  = ~A233 & \new_[9849]_ ;
  assign \new_[9853]_  = ~A266 & A265;
  assign \new_[9856]_  = A269 & A267;
  assign \new_[9857]_  = \new_[9856]_  & \new_[9853]_ ;
  assign \new_[9858]_  = \new_[9857]_  & \new_[9850]_ ;
  assign \new_[9862]_  = ~A167 & ~A169;
  assign \new_[9863]_  = A170 & \new_[9862]_ ;
  assign \new_[9866]_  = A199 & A166;
  assign \new_[9869]_  = A232 & ~A201;
  assign \new_[9870]_  = \new_[9869]_  & \new_[9866]_ ;
  assign \new_[9871]_  = \new_[9870]_  & \new_[9863]_ ;
  assign \new_[9875]_  = A235 & A234;
  assign \new_[9876]_  = ~A233 & \new_[9875]_ ;
  assign \new_[9879]_  = ~A299 & A298;
  assign \new_[9882]_  = A301 & A300;
  assign \new_[9883]_  = \new_[9882]_  & \new_[9879]_ ;
  assign \new_[9884]_  = \new_[9883]_  & \new_[9876]_ ;
  assign \new_[9888]_  = ~A167 & ~A169;
  assign \new_[9889]_  = A170 & \new_[9888]_ ;
  assign \new_[9892]_  = A199 & A166;
  assign \new_[9895]_  = A232 & ~A201;
  assign \new_[9896]_  = \new_[9895]_  & \new_[9892]_ ;
  assign \new_[9897]_  = \new_[9896]_  & \new_[9889]_ ;
  assign \new_[9901]_  = A235 & A234;
  assign \new_[9902]_  = ~A233 & \new_[9901]_ ;
  assign \new_[9905]_  = ~A299 & A298;
  assign \new_[9908]_  = A302 & A300;
  assign \new_[9909]_  = \new_[9908]_  & \new_[9905]_ ;
  assign \new_[9910]_  = \new_[9909]_  & \new_[9902]_ ;
  assign \new_[9914]_  = ~A167 & ~A169;
  assign \new_[9915]_  = A170 & \new_[9914]_ ;
  assign \new_[9918]_  = A199 & A166;
  assign \new_[9921]_  = A232 & ~A201;
  assign \new_[9922]_  = \new_[9921]_  & \new_[9918]_ ;
  assign \new_[9923]_  = \new_[9922]_  & \new_[9915]_ ;
  assign \new_[9927]_  = A235 & A234;
  assign \new_[9928]_  = ~A233 & \new_[9927]_ ;
  assign \new_[9931]_  = ~A266 & A265;
  assign \new_[9934]_  = A268 & A267;
  assign \new_[9935]_  = \new_[9934]_  & \new_[9931]_ ;
  assign \new_[9936]_  = \new_[9935]_  & \new_[9928]_ ;
  assign \new_[9940]_  = ~A167 & ~A169;
  assign \new_[9941]_  = A170 & \new_[9940]_ ;
  assign \new_[9944]_  = A199 & A166;
  assign \new_[9947]_  = A232 & ~A201;
  assign \new_[9948]_  = \new_[9947]_  & \new_[9944]_ ;
  assign \new_[9949]_  = \new_[9948]_  & \new_[9941]_ ;
  assign \new_[9953]_  = A235 & A234;
  assign \new_[9954]_  = ~A233 & \new_[9953]_ ;
  assign \new_[9957]_  = ~A266 & A265;
  assign \new_[9960]_  = A269 & A267;
  assign \new_[9961]_  = \new_[9960]_  & \new_[9957]_ ;
  assign \new_[9962]_  = \new_[9961]_  & \new_[9954]_ ;
  assign \new_[9966]_  = ~A167 & ~A169;
  assign \new_[9967]_  = A170 & \new_[9966]_ ;
  assign \new_[9970]_  = A199 & A166;
  assign \new_[9973]_  = A232 & ~A201;
  assign \new_[9974]_  = \new_[9973]_  & \new_[9970]_ ;
  assign \new_[9975]_  = \new_[9974]_  & \new_[9967]_ ;
  assign \new_[9979]_  = A236 & A234;
  assign \new_[9980]_  = ~A233 & \new_[9979]_ ;
  assign \new_[9983]_  = ~A299 & A298;
  assign \new_[9986]_  = A301 & A300;
  assign \new_[9987]_  = \new_[9986]_  & \new_[9983]_ ;
  assign \new_[9988]_  = \new_[9987]_  & \new_[9980]_ ;
  assign \new_[9992]_  = ~A167 & ~A169;
  assign \new_[9993]_  = A170 & \new_[9992]_ ;
  assign \new_[9996]_  = A199 & A166;
  assign \new_[9999]_  = A232 & ~A201;
  assign \new_[10000]_  = \new_[9999]_  & \new_[9996]_ ;
  assign \new_[10001]_  = \new_[10000]_  & \new_[9993]_ ;
  assign \new_[10005]_  = A236 & A234;
  assign \new_[10006]_  = ~A233 & \new_[10005]_ ;
  assign \new_[10009]_  = ~A299 & A298;
  assign \new_[10012]_  = A302 & A300;
  assign \new_[10013]_  = \new_[10012]_  & \new_[10009]_ ;
  assign \new_[10014]_  = \new_[10013]_  & \new_[10006]_ ;
  assign \new_[10018]_  = ~A167 & ~A169;
  assign \new_[10019]_  = A170 & \new_[10018]_ ;
  assign \new_[10022]_  = A199 & A166;
  assign \new_[10025]_  = A232 & ~A201;
  assign \new_[10026]_  = \new_[10025]_  & \new_[10022]_ ;
  assign \new_[10027]_  = \new_[10026]_  & \new_[10019]_ ;
  assign \new_[10031]_  = A236 & A234;
  assign \new_[10032]_  = ~A233 & \new_[10031]_ ;
  assign \new_[10035]_  = ~A266 & A265;
  assign \new_[10038]_  = A268 & A267;
  assign \new_[10039]_  = \new_[10038]_  & \new_[10035]_ ;
  assign \new_[10040]_  = \new_[10039]_  & \new_[10032]_ ;
  assign \new_[10044]_  = ~A167 & ~A169;
  assign \new_[10045]_  = A170 & \new_[10044]_ ;
  assign \new_[10048]_  = A199 & A166;
  assign \new_[10051]_  = A232 & ~A201;
  assign \new_[10052]_  = \new_[10051]_  & \new_[10048]_ ;
  assign \new_[10053]_  = \new_[10052]_  & \new_[10045]_ ;
  assign \new_[10057]_  = A236 & A234;
  assign \new_[10058]_  = ~A233 & \new_[10057]_ ;
  assign \new_[10061]_  = ~A266 & A265;
  assign \new_[10064]_  = A269 & A267;
  assign \new_[10065]_  = \new_[10064]_  & \new_[10061]_ ;
  assign \new_[10066]_  = \new_[10065]_  & \new_[10058]_ ;
  assign \new_[10070]_  = ~A167 & ~A169;
  assign \new_[10071]_  = A170 & \new_[10070]_ ;
  assign \new_[10074]_  = A199 & A166;
  assign \new_[10077]_  = A232 & A200;
  assign \new_[10078]_  = \new_[10077]_  & \new_[10074]_ ;
  assign \new_[10079]_  = \new_[10078]_  & \new_[10071]_ ;
  assign \new_[10083]_  = A235 & A234;
  assign \new_[10084]_  = ~A233 & \new_[10083]_ ;
  assign \new_[10087]_  = ~A299 & A298;
  assign \new_[10090]_  = A301 & A300;
  assign \new_[10091]_  = \new_[10090]_  & \new_[10087]_ ;
  assign \new_[10092]_  = \new_[10091]_  & \new_[10084]_ ;
  assign \new_[10096]_  = ~A167 & ~A169;
  assign \new_[10097]_  = A170 & \new_[10096]_ ;
  assign \new_[10100]_  = A199 & A166;
  assign \new_[10103]_  = A232 & A200;
  assign \new_[10104]_  = \new_[10103]_  & \new_[10100]_ ;
  assign \new_[10105]_  = \new_[10104]_  & \new_[10097]_ ;
  assign \new_[10109]_  = A235 & A234;
  assign \new_[10110]_  = ~A233 & \new_[10109]_ ;
  assign \new_[10113]_  = ~A299 & A298;
  assign \new_[10116]_  = A302 & A300;
  assign \new_[10117]_  = \new_[10116]_  & \new_[10113]_ ;
  assign \new_[10118]_  = \new_[10117]_  & \new_[10110]_ ;
  assign \new_[10122]_  = ~A167 & ~A169;
  assign \new_[10123]_  = A170 & \new_[10122]_ ;
  assign \new_[10126]_  = A199 & A166;
  assign \new_[10129]_  = A232 & A200;
  assign \new_[10130]_  = \new_[10129]_  & \new_[10126]_ ;
  assign \new_[10131]_  = \new_[10130]_  & \new_[10123]_ ;
  assign \new_[10135]_  = A235 & A234;
  assign \new_[10136]_  = ~A233 & \new_[10135]_ ;
  assign \new_[10139]_  = ~A266 & A265;
  assign \new_[10142]_  = A268 & A267;
  assign \new_[10143]_  = \new_[10142]_  & \new_[10139]_ ;
  assign \new_[10144]_  = \new_[10143]_  & \new_[10136]_ ;
  assign \new_[10148]_  = ~A167 & ~A169;
  assign \new_[10149]_  = A170 & \new_[10148]_ ;
  assign \new_[10152]_  = A199 & A166;
  assign \new_[10155]_  = A232 & A200;
  assign \new_[10156]_  = \new_[10155]_  & \new_[10152]_ ;
  assign \new_[10157]_  = \new_[10156]_  & \new_[10149]_ ;
  assign \new_[10161]_  = A235 & A234;
  assign \new_[10162]_  = ~A233 & \new_[10161]_ ;
  assign \new_[10165]_  = ~A266 & A265;
  assign \new_[10168]_  = A269 & A267;
  assign \new_[10169]_  = \new_[10168]_  & \new_[10165]_ ;
  assign \new_[10170]_  = \new_[10169]_  & \new_[10162]_ ;
  assign \new_[10174]_  = ~A167 & ~A169;
  assign \new_[10175]_  = A170 & \new_[10174]_ ;
  assign \new_[10178]_  = A199 & A166;
  assign \new_[10181]_  = A232 & A200;
  assign \new_[10182]_  = \new_[10181]_  & \new_[10178]_ ;
  assign \new_[10183]_  = \new_[10182]_  & \new_[10175]_ ;
  assign \new_[10187]_  = A236 & A234;
  assign \new_[10188]_  = ~A233 & \new_[10187]_ ;
  assign \new_[10191]_  = ~A299 & A298;
  assign \new_[10194]_  = A301 & A300;
  assign \new_[10195]_  = \new_[10194]_  & \new_[10191]_ ;
  assign \new_[10196]_  = \new_[10195]_  & \new_[10188]_ ;
  assign \new_[10200]_  = ~A167 & ~A169;
  assign \new_[10201]_  = A170 & \new_[10200]_ ;
  assign \new_[10204]_  = A199 & A166;
  assign \new_[10207]_  = A232 & A200;
  assign \new_[10208]_  = \new_[10207]_  & \new_[10204]_ ;
  assign \new_[10209]_  = \new_[10208]_  & \new_[10201]_ ;
  assign \new_[10213]_  = A236 & A234;
  assign \new_[10214]_  = ~A233 & \new_[10213]_ ;
  assign \new_[10217]_  = ~A299 & A298;
  assign \new_[10220]_  = A302 & A300;
  assign \new_[10221]_  = \new_[10220]_  & \new_[10217]_ ;
  assign \new_[10222]_  = \new_[10221]_  & \new_[10214]_ ;
  assign \new_[10226]_  = ~A167 & ~A169;
  assign \new_[10227]_  = A170 & \new_[10226]_ ;
  assign \new_[10230]_  = A199 & A166;
  assign \new_[10233]_  = A232 & A200;
  assign \new_[10234]_  = \new_[10233]_  & \new_[10230]_ ;
  assign \new_[10235]_  = \new_[10234]_  & \new_[10227]_ ;
  assign \new_[10239]_  = A236 & A234;
  assign \new_[10240]_  = ~A233 & \new_[10239]_ ;
  assign \new_[10243]_  = ~A266 & A265;
  assign \new_[10246]_  = A268 & A267;
  assign \new_[10247]_  = \new_[10246]_  & \new_[10243]_ ;
  assign \new_[10248]_  = \new_[10247]_  & \new_[10240]_ ;
  assign \new_[10252]_  = ~A167 & ~A169;
  assign \new_[10253]_  = A170 & \new_[10252]_ ;
  assign \new_[10256]_  = A199 & A166;
  assign \new_[10259]_  = A232 & A200;
  assign \new_[10260]_  = \new_[10259]_  & \new_[10256]_ ;
  assign \new_[10261]_  = \new_[10260]_  & \new_[10253]_ ;
  assign \new_[10265]_  = A236 & A234;
  assign \new_[10266]_  = ~A233 & \new_[10265]_ ;
  assign \new_[10269]_  = ~A266 & A265;
  assign \new_[10272]_  = A269 & A267;
  assign \new_[10273]_  = \new_[10272]_  & \new_[10269]_ ;
  assign \new_[10274]_  = \new_[10273]_  & \new_[10266]_ ;
  assign \new_[10278]_  = ~A167 & ~A169;
  assign \new_[10279]_  = A170 & \new_[10278]_ ;
  assign \new_[10282]_  = ~A199 & A166;
  assign \new_[10285]_  = A232 & ~A200;
  assign \new_[10286]_  = \new_[10285]_  & \new_[10282]_ ;
  assign \new_[10287]_  = \new_[10286]_  & \new_[10279]_ ;
  assign \new_[10291]_  = A235 & A234;
  assign \new_[10292]_  = ~A233 & \new_[10291]_ ;
  assign \new_[10295]_  = ~A299 & A298;
  assign \new_[10298]_  = A301 & A300;
  assign \new_[10299]_  = \new_[10298]_  & \new_[10295]_ ;
  assign \new_[10300]_  = \new_[10299]_  & \new_[10292]_ ;
  assign \new_[10304]_  = ~A167 & ~A169;
  assign \new_[10305]_  = A170 & \new_[10304]_ ;
  assign \new_[10308]_  = ~A199 & A166;
  assign \new_[10311]_  = A232 & ~A200;
  assign \new_[10312]_  = \new_[10311]_  & \new_[10308]_ ;
  assign \new_[10313]_  = \new_[10312]_  & \new_[10305]_ ;
  assign \new_[10317]_  = A235 & A234;
  assign \new_[10318]_  = ~A233 & \new_[10317]_ ;
  assign \new_[10321]_  = ~A299 & A298;
  assign \new_[10324]_  = A302 & A300;
  assign \new_[10325]_  = \new_[10324]_  & \new_[10321]_ ;
  assign \new_[10326]_  = \new_[10325]_  & \new_[10318]_ ;
  assign \new_[10330]_  = ~A167 & ~A169;
  assign \new_[10331]_  = A170 & \new_[10330]_ ;
  assign \new_[10334]_  = ~A199 & A166;
  assign \new_[10337]_  = A232 & ~A200;
  assign \new_[10338]_  = \new_[10337]_  & \new_[10334]_ ;
  assign \new_[10339]_  = \new_[10338]_  & \new_[10331]_ ;
  assign \new_[10343]_  = A235 & A234;
  assign \new_[10344]_  = ~A233 & \new_[10343]_ ;
  assign \new_[10347]_  = ~A266 & A265;
  assign \new_[10350]_  = A268 & A267;
  assign \new_[10351]_  = \new_[10350]_  & \new_[10347]_ ;
  assign \new_[10352]_  = \new_[10351]_  & \new_[10344]_ ;
  assign \new_[10356]_  = ~A167 & ~A169;
  assign \new_[10357]_  = A170 & \new_[10356]_ ;
  assign \new_[10360]_  = ~A199 & A166;
  assign \new_[10363]_  = A232 & ~A200;
  assign \new_[10364]_  = \new_[10363]_  & \new_[10360]_ ;
  assign \new_[10365]_  = \new_[10364]_  & \new_[10357]_ ;
  assign \new_[10369]_  = A235 & A234;
  assign \new_[10370]_  = ~A233 & \new_[10369]_ ;
  assign \new_[10373]_  = ~A266 & A265;
  assign \new_[10376]_  = A269 & A267;
  assign \new_[10377]_  = \new_[10376]_  & \new_[10373]_ ;
  assign \new_[10378]_  = \new_[10377]_  & \new_[10370]_ ;
  assign \new_[10382]_  = ~A167 & ~A169;
  assign \new_[10383]_  = A170 & \new_[10382]_ ;
  assign \new_[10386]_  = ~A199 & A166;
  assign \new_[10389]_  = A232 & ~A200;
  assign \new_[10390]_  = \new_[10389]_  & \new_[10386]_ ;
  assign \new_[10391]_  = \new_[10390]_  & \new_[10383]_ ;
  assign \new_[10395]_  = A236 & A234;
  assign \new_[10396]_  = ~A233 & \new_[10395]_ ;
  assign \new_[10399]_  = ~A299 & A298;
  assign \new_[10402]_  = A301 & A300;
  assign \new_[10403]_  = \new_[10402]_  & \new_[10399]_ ;
  assign \new_[10404]_  = \new_[10403]_  & \new_[10396]_ ;
  assign \new_[10408]_  = ~A167 & ~A169;
  assign \new_[10409]_  = A170 & \new_[10408]_ ;
  assign \new_[10412]_  = ~A199 & A166;
  assign \new_[10415]_  = A232 & ~A200;
  assign \new_[10416]_  = \new_[10415]_  & \new_[10412]_ ;
  assign \new_[10417]_  = \new_[10416]_  & \new_[10409]_ ;
  assign \new_[10421]_  = A236 & A234;
  assign \new_[10422]_  = ~A233 & \new_[10421]_ ;
  assign \new_[10425]_  = ~A299 & A298;
  assign \new_[10428]_  = A302 & A300;
  assign \new_[10429]_  = \new_[10428]_  & \new_[10425]_ ;
  assign \new_[10430]_  = \new_[10429]_  & \new_[10422]_ ;
  assign \new_[10434]_  = ~A167 & ~A169;
  assign \new_[10435]_  = A170 & \new_[10434]_ ;
  assign \new_[10438]_  = ~A199 & A166;
  assign \new_[10441]_  = A232 & ~A200;
  assign \new_[10442]_  = \new_[10441]_  & \new_[10438]_ ;
  assign \new_[10443]_  = \new_[10442]_  & \new_[10435]_ ;
  assign \new_[10447]_  = A236 & A234;
  assign \new_[10448]_  = ~A233 & \new_[10447]_ ;
  assign \new_[10451]_  = ~A266 & A265;
  assign \new_[10454]_  = A268 & A267;
  assign \new_[10455]_  = \new_[10454]_  & \new_[10451]_ ;
  assign \new_[10456]_  = \new_[10455]_  & \new_[10448]_ ;
  assign \new_[10460]_  = ~A167 & ~A169;
  assign \new_[10461]_  = A170 & \new_[10460]_ ;
  assign \new_[10464]_  = ~A199 & A166;
  assign \new_[10467]_  = A232 & ~A200;
  assign \new_[10468]_  = \new_[10467]_  & \new_[10464]_ ;
  assign \new_[10469]_  = \new_[10468]_  & \new_[10461]_ ;
  assign \new_[10473]_  = A236 & A234;
  assign \new_[10474]_  = ~A233 & \new_[10473]_ ;
  assign \new_[10477]_  = ~A266 & A265;
  assign \new_[10480]_  = A269 & A267;
  assign \new_[10481]_  = \new_[10480]_  & \new_[10477]_ ;
  assign \new_[10482]_  = \new_[10481]_  & \new_[10474]_ ;
  assign \new_[10486]_  = A167 & A169;
  assign \new_[10487]_  = ~A170 & \new_[10486]_ ;
  assign \new_[10490]_  = A199 & A166;
  assign \new_[10493]_  = ~A203 & ~A202;
  assign \new_[10494]_  = \new_[10493]_  & \new_[10490]_ ;
  assign \new_[10495]_  = \new_[10494]_  & \new_[10487]_ ;
  assign \new_[10498]_  = ~A233 & A232;
  assign \new_[10501]_  = A235 & A234;
  assign \new_[10502]_  = \new_[10501]_  & \new_[10498]_ ;
  assign \new_[10505]_  = ~A299 & A298;
  assign \new_[10508]_  = A301 & A300;
  assign \new_[10509]_  = \new_[10508]_  & \new_[10505]_ ;
  assign \new_[10510]_  = \new_[10509]_  & \new_[10502]_ ;
  assign \new_[10514]_  = A167 & A169;
  assign \new_[10515]_  = ~A170 & \new_[10514]_ ;
  assign \new_[10518]_  = A199 & A166;
  assign \new_[10521]_  = ~A203 & ~A202;
  assign \new_[10522]_  = \new_[10521]_  & \new_[10518]_ ;
  assign \new_[10523]_  = \new_[10522]_  & \new_[10515]_ ;
  assign \new_[10526]_  = ~A233 & A232;
  assign \new_[10529]_  = A235 & A234;
  assign \new_[10530]_  = \new_[10529]_  & \new_[10526]_ ;
  assign \new_[10533]_  = ~A299 & A298;
  assign \new_[10536]_  = A302 & A300;
  assign \new_[10537]_  = \new_[10536]_  & \new_[10533]_ ;
  assign \new_[10538]_  = \new_[10537]_  & \new_[10530]_ ;
  assign \new_[10542]_  = A167 & A169;
  assign \new_[10543]_  = ~A170 & \new_[10542]_ ;
  assign \new_[10546]_  = A199 & A166;
  assign \new_[10549]_  = ~A203 & ~A202;
  assign \new_[10550]_  = \new_[10549]_  & \new_[10546]_ ;
  assign \new_[10551]_  = \new_[10550]_  & \new_[10543]_ ;
  assign \new_[10554]_  = ~A233 & A232;
  assign \new_[10557]_  = A235 & A234;
  assign \new_[10558]_  = \new_[10557]_  & \new_[10554]_ ;
  assign \new_[10561]_  = ~A266 & A265;
  assign \new_[10564]_  = A268 & A267;
  assign \new_[10565]_  = \new_[10564]_  & \new_[10561]_ ;
  assign \new_[10566]_  = \new_[10565]_  & \new_[10558]_ ;
  assign \new_[10570]_  = A167 & A169;
  assign \new_[10571]_  = ~A170 & \new_[10570]_ ;
  assign \new_[10574]_  = A199 & A166;
  assign \new_[10577]_  = ~A203 & ~A202;
  assign \new_[10578]_  = \new_[10577]_  & \new_[10574]_ ;
  assign \new_[10579]_  = \new_[10578]_  & \new_[10571]_ ;
  assign \new_[10582]_  = ~A233 & A232;
  assign \new_[10585]_  = A235 & A234;
  assign \new_[10586]_  = \new_[10585]_  & \new_[10582]_ ;
  assign \new_[10589]_  = ~A266 & A265;
  assign \new_[10592]_  = A269 & A267;
  assign \new_[10593]_  = \new_[10592]_  & \new_[10589]_ ;
  assign \new_[10594]_  = \new_[10593]_  & \new_[10586]_ ;
  assign \new_[10598]_  = A167 & A169;
  assign \new_[10599]_  = ~A170 & \new_[10598]_ ;
  assign \new_[10602]_  = A199 & A166;
  assign \new_[10605]_  = ~A203 & ~A202;
  assign \new_[10606]_  = \new_[10605]_  & \new_[10602]_ ;
  assign \new_[10607]_  = \new_[10606]_  & \new_[10599]_ ;
  assign \new_[10610]_  = ~A233 & A232;
  assign \new_[10613]_  = A236 & A234;
  assign \new_[10614]_  = \new_[10613]_  & \new_[10610]_ ;
  assign \new_[10617]_  = ~A299 & A298;
  assign \new_[10620]_  = A301 & A300;
  assign \new_[10621]_  = \new_[10620]_  & \new_[10617]_ ;
  assign \new_[10622]_  = \new_[10621]_  & \new_[10614]_ ;
  assign \new_[10626]_  = A167 & A169;
  assign \new_[10627]_  = ~A170 & \new_[10626]_ ;
  assign \new_[10630]_  = A199 & A166;
  assign \new_[10633]_  = ~A203 & ~A202;
  assign \new_[10634]_  = \new_[10633]_  & \new_[10630]_ ;
  assign \new_[10635]_  = \new_[10634]_  & \new_[10627]_ ;
  assign \new_[10638]_  = ~A233 & A232;
  assign \new_[10641]_  = A236 & A234;
  assign \new_[10642]_  = \new_[10641]_  & \new_[10638]_ ;
  assign \new_[10645]_  = ~A299 & A298;
  assign \new_[10648]_  = A302 & A300;
  assign \new_[10649]_  = \new_[10648]_  & \new_[10645]_ ;
  assign \new_[10650]_  = \new_[10649]_  & \new_[10642]_ ;
  assign \new_[10654]_  = A167 & A169;
  assign \new_[10655]_  = ~A170 & \new_[10654]_ ;
  assign \new_[10658]_  = A199 & A166;
  assign \new_[10661]_  = ~A203 & ~A202;
  assign \new_[10662]_  = \new_[10661]_  & \new_[10658]_ ;
  assign \new_[10663]_  = \new_[10662]_  & \new_[10655]_ ;
  assign \new_[10666]_  = ~A233 & A232;
  assign \new_[10669]_  = A236 & A234;
  assign \new_[10670]_  = \new_[10669]_  & \new_[10666]_ ;
  assign \new_[10673]_  = ~A266 & A265;
  assign \new_[10676]_  = A268 & A267;
  assign \new_[10677]_  = \new_[10676]_  & \new_[10673]_ ;
  assign \new_[10678]_  = \new_[10677]_  & \new_[10670]_ ;
  assign \new_[10682]_  = A167 & A169;
  assign \new_[10683]_  = ~A170 & \new_[10682]_ ;
  assign \new_[10686]_  = A199 & A166;
  assign \new_[10689]_  = ~A203 & ~A202;
  assign \new_[10690]_  = \new_[10689]_  & \new_[10686]_ ;
  assign \new_[10691]_  = \new_[10690]_  & \new_[10683]_ ;
  assign \new_[10694]_  = ~A233 & A232;
  assign \new_[10697]_  = A236 & A234;
  assign \new_[10698]_  = \new_[10697]_  & \new_[10694]_ ;
  assign \new_[10701]_  = ~A266 & A265;
  assign \new_[10704]_  = A269 & A267;
  assign \new_[10705]_  = \new_[10704]_  & \new_[10701]_ ;
  assign \new_[10706]_  = \new_[10705]_  & \new_[10698]_ ;
  assign \new_[10710]_  = ~A167 & A169;
  assign \new_[10711]_  = ~A170 & \new_[10710]_ ;
  assign \new_[10714]_  = A199 & ~A166;
  assign \new_[10717]_  = ~A203 & ~A202;
  assign \new_[10718]_  = \new_[10717]_  & \new_[10714]_ ;
  assign \new_[10719]_  = \new_[10718]_  & \new_[10711]_ ;
  assign \new_[10722]_  = ~A233 & A232;
  assign \new_[10725]_  = A235 & A234;
  assign \new_[10726]_  = \new_[10725]_  & \new_[10722]_ ;
  assign \new_[10729]_  = ~A299 & A298;
  assign \new_[10732]_  = A301 & A300;
  assign \new_[10733]_  = \new_[10732]_  & \new_[10729]_ ;
  assign \new_[10734]_  = \new_[10733]_  & \new_[10726]_ ;
  assign \new_[10738]_  = ~A167 & A169;
  assign \new_[10739]_  = ~A170 & \new_[10738]_ ;
  assign \new_[10742]_  = A199 & ~A166;
  assign \new_[10745]_  = ~A203 & ~A202;
  assign \new_[10746]_  = \new_[10745]_  & \new_[10742]_ ;
  assign \new_[10747]_  = \new_[10746]_  & \new_[10739]_ ;
  assign \new_[10750]_  = ~A233 & A232;
  assign \new_[10753]_  = A235 & A234;
  assign \new_[10754]_  = \new_[10753]_  & \new_[10750]_ ;
  assign \new_[10757]_  = ~A299 & A298;
  assign \new_[10760]_  = A302 & A300;
  assign \new_[10761]_  = \new_[10760]_  & \new_[10757]_ ;
  assign \new_[10762]_  = \new_[10761]_  & \new_[10754]_ ;
  assign \new_[10766]_  = ~A167 & A169;
  assign \new_[10767]_  = ~A170 & \new_[10766]_ ;
  assign \new_[10770]_  = A199 & ~A166;
  assign \new_[10773]_  = ~A203 & ~A202;
  assign \new_[10774]_  = \new_[10773]_  & \new_[10770]_ ;
  assign \new_[10775]_  = \new_[10774]_  & \new_[10767]_ ;
  assign \new_[10778]_  = ~A233 & A232;
  assign \new_[10781]_  = A235 & A234;
  assign \new_[10782]_  = \new_[10781]_  & \new_[10778]_ ;
  assign \new_[10785]_  = ~A266 & A265;
  assign \new_[10788]_  = A268 & A267;
  assign \new_[10789]_  = \new_[10788]_  & \new_[10785]_ ;
  assign \new_[10790]_  = \new_[10789]_  & \new_[10782]_ ;
  assign \new_[10794]_  = ~A167 & A169;
  assign \new_[10795]_  = ~A170 & \new_[10794]_ ;
  assign \new_[10798]_  = A199 & ~A166;
  assign \new_[10801]_  = ~A203 & ~A202;
  assign \new_[10802]_  = \new_[10801]_  & \new_[10798]_ ;
  assign \new_[10803]_  = \new_[10802]_  & \new_[10795]_ ;
  assign \new_[10806]_  = ~A233 & A232;
  assign \new_[10809]_  = A235 & A234;
  assign \new_[10810]_  = \new_[10809]_  & \new_[10806]_ ;
  assign \new_[10813]_  = ~A266 & A265;
  assign \new_[10816]_  = A269 & A267;
  assign \new_[10817]_  = \new_[10816]_  & \new_[10813]_ ;
  assign \new_[10818]_  = \new_[10817]_  & \new_[10810]_ ;
  assign \new_[10822]_  = ~A167 & A169;
  assign \new_[10823]_  = ~A170 & \new_[10822]_ ;
  assign \new_[10826]_  = A199 & ~A166;
  assign \new_[10829]_  = ~A203 & ~A202;
  assign \new_[10830]_  = \new_[10829]_  & \new_[10826]_ ;
  assign \new_[10831]_  = \new_[10830]_  & \new_[10823]_ ;
  assign \new_[10834]_  = ~A233 & A232;
  assign \new_[10837]_  = A236 & A234;
  assign \new_[10838]_  = \new_[10837]_  & \new_[10834]_ ;
  assign \new_[10841]_  = ~A299 & A298;
  assign \new_[10844]_  = A301 & A300;
  assign \new_[10845]_  = \new_[10844]_  & \new_[10841]_ ;
  assign \new_[10846]_  = \new_[10845]_  & \new_[10838]_ ;
  assign \new_[10850]_  = ~A167 & A169;
  assign \new_[10851]_  = ~A170 & \new_[10850]_ ;
  assign \new_[10854]_  = A199 & ~A166;
  assign \new_[10857]_  = ~A203 & ~A202;
  assign \new_[10858]_  = \new_[10857]_  & \new_[10854]_ ;
  assign \new_[10859]_  = \new_[10858]_  & \new_[10851]_ ;
  assign \new_[10862]_  = ~A233 & A232;
  assign \new_[10865]_  = A236 & A234;
  assign \new_[10866]_  = \new_[10865]_  & \new_[10862]_ ;
  assign \new_[10869]_  = ~A299 & A298;
  assign \new_[10872]_  = A302 & A300;
  assign \new_[10873]_  = \new_[10872]_  & \new_[10869]_ ;
  assign \new_[10874]_  = \new_[10873]_  & \new_[10866]_ ;
  assign \new_[10878]_  = ~A167 & A169;
  assign \new_[10879]_  = ~A170 & \new_[10878]_ ;
  assign \new_[10882]_  = A199 & ~A166;
  assign \new_[10885]_  = ~A203 & ~A202;
  assign \new_[10886]_  = \new_[10885]_  & \new_[10882]_ ;
  assign \new_[10887]_  = \new_[10886]_  & \new_[10879]_ ;
  assign \new_[10890]_  = ~A233 & A232;
  assign \new_[10893]_  = A236 & A234;
  assign \new_[10894]_  = \new_[10893]_  & \new_[10890]_ ;
  assign \new_[10897]_  = ~A266 & A265;
  assign \new_[10900]_  = A268 & A267;
  assign \new_[10901]_  = \new_[10900]_  & \new_[10897]_ ;
  assign \new_[10902]_  = \new_[10901]_  & \new_[10894]_ ;
  assign \new_[10906]_  = ~A167 & A169;
  assign \new_[10907]_  = ~A170 & \new_[10906]_ ;
  assign \new_[10910]_  = A199 & ~A166;
  assign \new_[10913]_  = ~A203 & ~A202;
  assign \new_[10914]_  = \new_[10913]_  & \new_[10910]_ ;
  assign \new_[10915]_  = \new_[10914]_  & \new_[10907]_ ;
  assign \new_[10918]_  = ~A233 & A232;
  assign \new_[10921]_  = A236 & A234;
  assign \new_[10922]_  = \new_[10921]_  & \new_[10918]_ ;
  assign \new_[10925]_  = ~A266 & A265;
  assign \new_[10928]_  = A269 & A267;
  assign \new_[10929]_  = \new_[10928]_  & \new_[10925]_ ;
  assign \new_[10930]_  = \new_[10929]_  & \new_[10922]_ ;
  assign \new_[10934]_  = A167 & ~A169;
  assign \new_[10935]_  = A170 & \new_[10934]_ ;
  assign \new_[10938]_  = A199 & ~A166;
  assign \new_[10941]_  = ~A203 & ~A202;
  assign \new_[10942]_  = \new_[10941]_  & \new_[10938]_ ;
  assign \new_[10943]_  = \new_[10942]_  & \new_[10935]_ ;
  assign \new_[10946]_  = ~A233 & A232;
  assign \new_[10949]_  = A235 & A234;
  assign \new_[10950]_  = \new_[10949]_  & \new_[10946]_ ;
  assign \new_[10953]_  = ~A299 & A298;
  assign \new_[10956]_  = A301 & A300;
  assign \new_[10957]_  = \new_[10956]_  & \new_[10953]_ ;
  assign \new_[10958]_  = \new_[10957]_  & \new_[10950]_ ;
  assign \new_[10962]_  = A167 & ~A169;
  assign \new_[10963]_  = A170 & \new_[10962]_ ;
  assign \new_[10966]_  = A199 & ~A166;
  assign \new_[10969]_  = ~A203 & ~A202;
  assign \new_[10970]_  = \new_[10969]_  & \new_[10966]_ ;
  assign \new_[10971]_  = \new_[10970]_  & \new_[10963]_ ;
  assign \new_[10974]_  = ~A233 & A232;
  assign \new_[10977]_  = A235 & A234;
  assign \new_[10978]_  = \new_[10977]_  & \new_[10974]_ ;
  assign \new_[10981]_  = ~A299 & A298;
  assign \new_[10984]_  = A302 & A300;
  assign \new_[10985]_  = \new_[10984]_  & \new_[10981]_ ;
  assign \new_[10986]_  = \new_[10985]_  & \new_[10978]_ ;
  assign \new_[10990]_  = A167 & ~A169;
  assign \new_[10991]_  = A170 & \new_[10990]_ ;
  assign \new_[10994]_  = A199 & ~A166;
  assign \new_[10997]_  = ~A203 & ~A202;
  assign \new_[10998]_  = \new_[10997]_  & \new_[10994]_ ;
  assign \new_[10999]_  = \new_[10998]_  & \new_[10991]_ ;
  assign \new_[11002]_  = ~A233 & A232;
  assign \new_[11005]_  = A235 & A234;
  assign \new_[11006]_  = \new_[11005]_  & \new_[11002]_ ;
  assign \new_[11009]_  = ~A266 & A265;
  assign \new_[11012]_  = A268 & A267;
  assign \new_[11013]_  = \new_[11012]_  & \new_[11009]_ ;
  assign \new_[11014]_  = \new_[11013]_  & \new_[11006]_ ;
  assign \new_[11018]_  = A167 & ~A169;
  assign \new_[11019]_  = A170 & \new_[11018]_ ;
  assign \new_[11022]_  = A199 & ~A166;
  assign \new_[11025]_  = ~A203 & ~A202;
  assign \new_[11026]_  = \new_[11025]_  & \new_[11022]_ ;
  assign \new_[11027]_  = \new_[11026]_  & \new_[11019]_ ;
  assign \new_[11030]_  = ~A233 & A232;
  assign \new_[11033]_  = A235 & A234;
  assign \new_[11034]_  = \new_[11033]_  & \new_[11030]_ ;
  assign \new_[11037]_  = ~A266 & A265;
  assign \new_[11040]_  = A269 & A267;
  assign \new_[11041]_  = \new_[11040]_  & \new_[11037]_ ;
  assign \new_[11042]_  = \new_[11041]_  & \new_[11034]_ ;
  assign \new_[11046]_  = A167 & ~A169;
  assign \new_[11047]_  = A170 & \new_[11046]_ ;
  assign \new_[11050]_  = A199 & ~A166;
  assign \new_[11053]_  = ~A203 & ~A202;
  assign \new_[11054]_  = \new_[11053]_  & \new_[11050]_ ;
  assign \new_[11055]_  = \new_[11054]_  & \new_[11047]_ ;
  assign \new_[11058]_  = ~A233 & A232;
  assign \new_[11061]_  = A236 & A234;
  assign \new_[11062]_  = \new_[11061]_  & \new_[11058]_ ;
  assign \new_[11065]_  = ~A299 & A298;
  assign \new_[11068]_  = A301 & A300;
  assign \new_[11069]_  = \new_[11068]_  & \new_[11065]_ ;
  assign \new_[11070]_  = \new_[11069]_  & \new_[11062]_ ;
  assign \new_[11074]_  = A167 & ~A169;
  assign \new_[11075]_  = A170 & \new_[11074]_ ;
  assign \new_[11078]_  = A199 & ~A166;
  assign \new_[11081]_  = ~A203 & ~A202;
  assign \new_[11082]_  = \new_[11081]_  & \new_[11078]_ ;
  assign \new_[11083]_  = \new_[11082]_  & \new_[11075]_ ;
  assign \new_[11086]_  = ~A233 & A232;
  assign \new_[11089]_  = A236 & A234;
  assign \new_[11090]_  = \new_[11089]_  & \new_[11086]_ ;
  assign \new_[11093]_  = ~A299 & A298;
  assign \new_[11096]_  = A302 & A300;
  assign \new_[11097]_  = \new_[11096]_  & \new_[11093]_ ;
  assign \new_[11098]_  = \new_[11097]_  & \new_[11090]_ ;
  assign \new_[11102]_  = A167 & ~A169;
  assign \new_[11103]_  = A170 & \new_[11102]_ ;
  assign \new_[11106]_  = A199 & ~A166;
  assign \new_[11109]_  = ~A203 & ~A202;
  assign \new_[11110]_  = \new_[11109]_  & \new_[11106]_ ;
  assign \new_[11111]_  = \new_[11110]_  & \new_[11103]_ ;
  assign \new_[11114]_  = ~A233 & A232;
  assign \new_[11117]_  = A236 & A234;
  assign \new_[11118]_  = \new_[11117]_  & \new_[11114]_ ;
  assign \new_[11121]_  = ~A266 & A265;
  assign \new_[11124]_  = A268 & A267;
  assign \new_[11125]_  = \new_[11124]_  & \new_[11121]_ ;
  assign \new_[11126]_  = \new_[11125]_  & \new_[11118]_ ;
  assign \new_[11130]_  = A167 & ~A169;
  assign \new_[11131]_  = A170 & \new_[11130]_ ;
  assign \new_[11134]_  = A199 & ~A166;
  assign \new_[11137]_  = ~A203 & ~A202;
  assign \new_[11138]_  = \new_[11137]_  & \new_[11134]_ ;
  assign \new_[11139]_  = \new_[11138]_  & \new_[11131]_ ;
  assign \new_[11142]_  = ~A233 & A232;
  assign \new_[11145]_  = A236 & A234;
  assign \new_[11146]_  = \new_[11145]_  & \new_[11142]_ ;
  assign \new_[11149]_  = ~A266 & A265;
  assign \new_[11152]_  = A269 & A267;
  assign \new_[11153]_  = \new_[11152]_  & \new_[11149]_ ;
  assign \new_[11154]_  = \new_[11153]_  & \new_[11146]_ ;
  assign \new_[11158]_  = ~A167 & ~A169;
  assign \new_[11159]_  = A170 & \new_[11158]_ ;
  assign \new_[11162]_  = A199 & A166;
  assign \new_[11165]_  = ~A203 & ~A202;
  assign \new_[11166]_  = \new_[11165]_  & \new_[11162]_ ;
  assign \new_[11167]_  = \new_[11166]_  & \new_[11159]_ ;
  assign \new_[11170]_  = ~A233 & A232;
  assign \new_[11173]_  = A235 & A234;
  assign \new_[11174]_  = \new_[11173]_  & \new_[11170]_ ;
  assign \new_[11177]_  = ~A299 & A298;
  assign \new_[11180]_  = A301 & A300;
  assign \new_[11181]_  = \new_[11180]_  & \new_[11177]_ ;
  assign \new_[11182]_  = \new_[11181]_  & \new_[11174]_ ;
  assign \new_[11186]_  = ~A167 & ~A169;
  assign \new_[11187]_  = A170 & \new_[11186]_ ;
  assign \new_[11190]_  = A199 & A166;
  assign \new_[11193]_  = ~A203 & ~A202;
  assign \new_[11194]_  = \new_[11193]_  & \new_[11190]_ ;
  assign \new_[11195]_  = \new_[11194]_  & \new_[11187]_ ;
  assign \new_[11198]_  = ~A233 & A232;
  assign \new_[11201]_  = A235 & A234;
  assign \new_[11202]_  = \new_[11201]_  & \new_[11198]_ ;
  assign \new_[11205]_  = ~A299 & A298;
  assign \new_[11208]_  = A302 & A300;
  assign \new_[11209]_  = \new_[11208]_  & \new_[11205]_ ;
  assign \new_[11210]_  = \new_[11209]_  & \new_[11202]_ ;
  assign \new_[11214]_  = ~A167 & ~A169;
  assign \new_[11215]_  = A170 & \new_[11214]_ ;
  assign \new_[11218]_  = A199 & A166;
  assign \new_[11221]_  = ~A203 & ~A202;
  assign \new_[11222]_  = \new_[11221]_  & \new_[11218]_ ;
  assign \new_[11223]_  = \new_[11222]_  & \new_[11215]_ ;
  assign \new_[11226]_  = ~A233 & A232;
  assign \new_[11229]_  = A235 & A234;
  assign \new_[11230]_  = \new_[11229]_  & \new_[11226]_ ;
  assign \new_[11233]_  = ~A266 & A265;
  assign \new_[11236]_  = A268 & A267;
  assign \new_[11237]_  = \new_[11236]_  & \new_[11233]_ ;
  assign \new_[11238]_  = \new_[11237]_  & \new_[11230]_ ;
  assign \new_[11242]_  = ~A167 & ~A169;
  assign \new_[11243]_  = A170 & \new_[11242]_ ;
  assign \new_[11246]_  = A199 & A166;
  assign \new_[11249]_  = ~A203 & ~A202;
  assign \new_[11250]_  = \new_[11249]_  & \new_[11246]_ ;
  assign \new_[11251]_  = \new_[11250]_  & \new_[11243]_ ;
  assign \new_[11254]_  = ~A233 & A232;
  assign \new_[11257]_  = A235 & A234;
  assign \new_[11258]_  = \new_[11257]_  & \new_[11254]_ ;
  assign \new_[11261]_  = ~A266 & A265;
  assign \new_[11264]_  = A269 & A267;
  assign \new_[11265]_  = \new_[11264]_  & \new_[11261]_ ;
  assign \new_[11266]_  = \new_[11265]_  & \new_[11258]_ ;
  assign \new_[11270]_  = ~A167 & ~A169;
  assign \new_[11271]_  = A170 & \new_[11270]_ ;
  assign \new_[11274]_  = A199 & A166;
  assign \new_[11277]_  = ~A203 & ~A202;
  assign \new_[11278]_  = \new_[11277]_  & \new_[11274]_ ;
  assign \new_[11279]_  = \new_[11278]_  & \new_[11271]_ ;
  assign \new_[11282]_  = ~A233 & A232;
  assign \new_[11285]_  = A236 & A234;
  assign \new_[11286]_  = \new_[11285]_  & \new_[11282]_ ;
  assign \new_[11289]_  = ~A299 & A298;
  assign \new_[11292]_  = A301 & A300;
  assign \new_[11293]_  = \new_[11292]_  & \new_[11289]_ ;
  assign \new_[11294]_  = \new_[11293]_  & \new_[11286]_ ;
  assign \new_[11298]_  = ~A167 & ~A169;
  assign \new_[11299]_  = A170 & \new_[11298]_ ;
  assign \new_[11302]_  = A199 & A166;
  assign \new_[11305]_  = ~A203 & ~A202;
  assign \new_[11306]_  = \new_[11305]_  & \new_[11302]_ ;
  assign \new_[11307]_  = \new_[11306]_  & \new_[11299]_ ;
  assign \new_[11310]_  = ~A233 & A232;
  assign \new_[11313]_  = A236 & A234;
  assign \new_[11314]_  = \new_[11313]_  & \new_[11310]_ ;
  assign \new_[11317]_  = ~A299 & A298;
  assign \new_[11320]_  = A302 & A300;
  assign \new_[11321]_  = \new_[11320]_  & \new_[11317]_ ;
  assign \new_[11322]_  = \new_[11321]_  & \new_[11314]_ ;
  assign \new_[11326]_  = ~A167 & ~A169;
  assign \new_[11327]_  = A170 & \new_[11326]_ ;
  assign \new_[11330]_  = A199 & A166;
  assign \new_[11333]_  = ~A203 & ~A202;
  assign \new_[11334]_  = \new_[11333]_  & \new_[11330]_ ;
  assign \new_[11335]_  = \new_[11334]_  & \new_[11327]_ ;
  assign \new_[11338]_  = ~A233 & A232;
  assign \new_[11341]_  = A236 & A234;
  assign \new_[11342]_  = \new_[11341]_  & \new_[11338]_ ;
  assign \new_[11345]_  = ~A266 & A265;
  assign \new_[11348]_  = A268 & A267;
  assign \new_[11349]_  = \new_[11348]_  & \new_[11345]_ ;
  assign \new_[11350]_  = \new_[11349]_  & \new_[11342]_ ;
  assign \new_[11354]_  = ~A167 & ~A169;
  assign \new_[11355]_  = A170 & \new_[11354]_ ;
  assign \new_[11358]_  = A199 & A166;
  assign \new_[11361]_  = ~A203 & ~A202;
  assign \new_[11362]_  = \new_[11361]_  & \new_[11358]_ ;
  assign \new_[11363]_  = \new_[11362]_  & \new_[11355]_ ;
  assign \new_[11366]_  = ~A233 & A232;
  assign \new_[11369]_  = A236 & A234;
  assign \new_[11370]_  = \new_[11369]_  & \new_[11366]_ ;
  assign \new_[11373]_  = ~A266 & A265;
  assign \new_[11376]_  = A269 & A267;
  assign \new_[11377]_  = \new_[11376]_  & \new_[11373]_ ;
  assign \new_[11378]_  = \new_[11377]_  & \new_[11370]_ ;
endmodule


