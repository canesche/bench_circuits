module top ( clock, 
    pg7, pg6, pg5, pg4, pg3, pg2, pg1, pg0, pg9, pg8, pclk, pg10, pg12,
    pg11, pg13,
    pg550, pg530, pg539, pg549, pg45, pg542, pg532, pg537, pg548, pg551,
    pg547, pg552, pg535, pg546  );
  input  clock;
  input  pg7, pg6, pg5, pg4, pg3, pg2, pg1, pg0, pg9, pg8, pclk, pg10,
    pg12, pg11, pg13;
  output pg550, pg530, pg539, pg549, pg45, pg542, pg532, pg537, pg548, pg551,
    pg547, pg552, pg535, pg546;
  reg ng38, ng34, ng35, ng36, ng37, ng30, ng31, ng32, ng33, ng29, ng39,
    ng40, ng41, ng42, ng43, ng44, ng45, ng46;
  wire new_n84_, new_n85_1_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_1_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_1_,
    new_n96_, new_n97_, new_n98_, new_n99_, new_n100_1_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_1_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_1_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_1_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_1_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_1_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_1_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_1_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_1_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_1_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n473_, new_n474_, new_n475_,
    new_n477_, new_n478_, new_n480_, new_n482_, new_n484_, new_n485_,
    new_n487_, new_n488_, new_n489_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n496_, new_n497_, new_n498_, new_n500_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n543_,
    new_n544_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, n60, n65, n70, n75, n80,
    n85, n90, n95, n100, n105, n110, n115, n120, n125, n130, n135, n140,
    n145;
  assign new_n84_ = ~pg13 & ~ng33;
  assign new_n85_1_ = pg3 & new_n84_;
  assign new_n86_ = pg5 & pg3;
  assign new_n87_ = pg7 & pg10;
  assign new_n88_ = pg9 & pg11;
  assign new_n89_ = pg8 & new_n88_;
  assign new_n90_1_ = new_n87_ & ~new_n89_;
  assign new_n91_ = pg9 & ~pg10;
  assign new_n92_ = pg7 & new_n91_;
  assign new_n93_ = ~pg7 & pg8;
  assign new_n94_ = ng30 & new_n93_;
  assign new_n95_1_ = ~new_n90_1_ & ~new_n92_;
  assign new_n96_ = ~new_n94_ & new_n95_1_;
  assign new_n97_ = ng32 & ~new_n96_;
  assign new_n98_ = ~pg12 & new_n97_;
  assign new_n99_ = ~pg13 & new_n98_;
  assign new_n100_1_ = pg4 & pg2;
  assign new_n101_ = new_n86_ & new_n99_;
  assign new_n102_ = ~new_n100_1_ & new_n101_;
  assign new_n103_ = ~pg5 & pg4;
  assign new_n104_ = pg4 & ~new_n86_;
  assign new_n105_1_ = pg5 & ~pg1;
  assign new_n106_ = ~new_n104_ & ~new_n105_1_;
  assign new_n107_ = pg2 & ~new_n106_;
  assign new_n108_ = ~pg3 & ~new_n107_;
  assign new_n109_ = ~pg5 & new_n108_;
  assign new_n110_1_ = ~pg4 & ~pg0;
  assign new_n111_ = pg3 & new_n110_1_;
  assign new_n112_ = ~new_n109_ & ~new_n111_;
  assign new_n113_ = ~new_n103_ & ~new_n112_;
  assign new_n114_ = ~pg7 & ~pg11;
  assign new_n115_1_ = pg8 & ~ng31;
  assign new_n116_ = ~pg8 & pg10;
  assign new_n117_ = ~new_n115_1_ & ~new_n116_;
  assign new_n118_ = pg9 & new_n114_;
  assign new_n119_ = ~new_n117_ & new_n118_;
  assign new_n120_1_ = ~pg6 & ~ng30;
  assign new_n121_ = ~pg7 & ~pg8;
  assign new_n122_ = ~pg9 & new_n121_;
  assign new_n123_ = pg7 & ng30;
  assign new_n124_ = ~pg6 & new_n123_;
  assign new_n125_1_ = pg8 & pg10;
  assign new_n126_ = pg9 & ~new_n125_1_;
  assign new_n127_ = new_n115_1_ & ~new_n124_;
  assign new_n128_ = ~new_n126_ & new_n127_;
  assign new_n129_ = ~new_n120_1_ & ~new_n122_;
  assign new_n130_1_ = ~new_n128_ & new_n129_;
  assign new_n131_ = pg11 & ~new_n130_1_;
  assign new_n132_ = pg8 & ng31;
  assign new_n133_ = ~pg10 & ~pg11;
  assign new_n134_ = ~pg9 & new_n133_;
  assign new_n135_1_ = ~new_n124_ & ~new_n132_;
  assign new_n136_ = new_n134_ & new_n135_1_;
  assign new_n137_ = ~new_n113_ & ~new_n119_;
  assign new_n138_ = ~new_n131_ & new_n137_;
  assign new_n139_ = ~new_n136_ & new_n138_;
  assign new_n140_1_ = ng46 & new_n139_;
  assign new_n141_ = pg12 & new_n140_1_;
  assign new_n142_ = ~pg13 & new_n141_;
  assign new_n143_ = pg0 & ~ng29;
  assign new_n144_ = pg4 & pg1;
  assign new_n145_1_ = ~pg0 & new_n144_;
  assign new_n146_ = pg3 & new_n145_1_;
  assign new_n147_ = ~new_n143_ & ~new_n146_;
  assign new_n148_ = new_n142_ & ~new_n147_;
  assign new_n149_ = ~pg6 & pg2;
  assign new_n150_ = new_n144_ & new_n149_;
  assign new_n151_ = pg2 & ~pg1;
  assign new_n152_ = pg6 & ~pg4;
  assign new_n153_ = ~pg5 & ~new_n152_;
  assign new_n154_ = new_n151_ & ~new_n153_;
  assign new_n155_ = ~pg3 & pg2;
  assign new_n156_ = pg3 & ~pg2;
  assign new_n157_ = ~new_n104_ & ~new_n155_;
  assign new_n158_ = ~new_n156_ & new_n157_;
  assign new_n159_ = pg6 & ~new_n158_;
  assign new_n160_ = ~pg6 & ~pg4;
  assign new_n161_ = pg6 & pg4;
  assign new_n162_ = pg3 & ~new_n161_;
  assign new_n163_ = ~new_n160_ & ~new_n162_;
  assign new_n164_ = pg5 & ~new_n163_;
  assign new_n165_ = ~pg3 & new_n103_;
  assign new_n166_ = ~new_n159_ & ~new_n164_;
  assign new_n167_ = ~new_n165_ & new_n166_;
  assign new_n168_ = pg1 & ~new_n167_;
  assign new_n169_ = ~new_n150_ & ~new_n154_;
  assign new_n170_ = ~new_n168_ & new_n169_;
  assign new_n171_ = ~new_n96_ & ~new_n170_;
  assign new_n172_ = new_n144_ & new_n171_;
  assign new_n173_ = ~pg5 & new_n172_;
  assign new_n174_ = ~new_n144_ & new_n171_;
  assign new_n175_ = pg5 & new_n174_;
  assign new_n176_ = ~new_n173_ & ~new_n175_;
  assign new_n177_ = ~pg12 & pg13;
  assign new_n178_ = ~new_n176_ & new_n177_;
  assign new_n179_ = pg2 & new_n178_;
  assign new_n180_ = ~new_n85_1_ & ~new_n102_;
  assign new_n181_ = ~new_n148_ & ~new_n179_;
  assign pg550 = ~new_n180_ | ~new_n181_;
  assign new_n183_ = pg7 & ~pg10;
  assign new_n184_ = ~pg9 & new_n183_;
  assign new_n185_ = pg8 & new_n184_;
  assign new_n186_ = pg9 & new_n116_;
  assign new_n187_ = ~pg7 & new_n186_;
  assign new_n188_ = ~new_n185_ & ~new_n187_;
  assign new_n189_ = pg5 & new_n161_;
  assign new_n190_ = ~new_n188_ & new_n189_;
  assign new_n191_ = pg11 & new_n190_;
  assign new_n192_ = ~pg6 & ng36;
  assign new_n193_ = ~new_n191_ & ~new_n192_;
  assign new_n194_ = ~pg3 & ~new_n193_;
  assign new_n195_ = ~pg13 & ~new_n97_;
  assign new_n196_ = ~pg5 & ~pg4;
  assign new_n197_ = pg11 & new_n196_;
  assign new_n198_ = pg3 & ng35;
  assign new_n199_ = new_n197_ & new_n198_;
  assign new_n200_ = ~pg8 & new_n114_;
  assign new_n201_ = new_n91_ & new_n200_;
  assign new_n202_ = pg5 & new_n201_;
  assign new_n203_ = pg3 & new_n161_;
  assign new_n204_ = new_n202_ & new_n203_;
  assign new_n205_ = new_n87_ & new_n89_;
  assign new_n206_ = new_n161_ & new_n205_;
  assign new_n207_ = new_n86_ & new_n206_;
  assign new_n208_ = ~new_n199_ & ~new_n204_;
  assign new_n209_ = ~new_n207_ & new_n208_;
  assign new_n210_ = pg2 & ~new_n209_;
  assign new_n211_ = ~pg2 & new_n194_;
  assign new_n212_ = new_n91_ & new_n93_;
  assign new_n213_ = new_n188_ & ~new_n212_;
  assign new_n214_ = pg11 & new_n203_;
  assign new_n215_ = ~pg5 & new_n214_;
  assign new_n216_ = ~new_n213_ & new_n215_;
  assign new_n217_ = ~pg2 & new_n216_;
  assign new_n218_ = ~new_n210_ & ~new_n211_;
  assign new_n219_ = ~new_n217_ & new_n218_;
  assign new_n220_ = new_n195_ & ~new_n219_;
  assign new_n221_ = ~pg12 & new_n220_;
  assign new_n222_ = new_n194_ & new_n221_;
  assign new_n223_ = ~pg4 & new_n86_;
  assign new_n224_ = pg3 & pg1;
  assign new_n225_ = ~pg5 & new_n224_;
  assign new_n226_ = new_n106_ & ~new_n223_;
  assign new_n227_ = ~new_n225_ & new_n226_;
  assign new_n228_ = pg0 & ~new_n227_;
  assign new_n229_ = pg1 & ~pg0;
  assign new_n230_ = ~new_n228_ & ~new_n229_;
  assign new_n231_ = new_n142_ & ~new_n230_;
  assign new_n232_ = pg2 & new_n231_;
  assign pg530 = new_n222_ | new_n232_;
  assign new_n234_ = ~pg13 & ~new_n140_1_;
  assign new_n235_ = pg12 & new_n234_;
  assign new_n236_ = pg0 & new_n207_;
  assign new_n237_ = new_n86_ & new_n183_;
  assign new_n238_ = ng37 & new_n237_;
  assign new_n239_ = pg8 & new_n238_;
  assign new_n240_ = pg6 & ~pg9;
  assign new_n241_ = ~pg7 & ~pg5;
  assign new_n242_ = new_n240_ & new_n241_;
  assign new_n243_ = new_n116_ & new_n242_;
  assign new_n244_ = ~pg3 & new_n243_;
  assign new_n245_ = ~new_n239_ & ~new_n244_;
  assign new_n246_ = new_n110_1_ & ~new_n245_;
  assign new_n247_ = pg11 & new_n246_;
  assign new_n248_ = ~new_n236_ & ~new_n247_;
  assign new_n249_ = pg2 & ~new_n248_;
  assign new_n250_ = pg1 & new_n249_;
  assign new_n251_ = new_n235_ & ~new_n250_;
  assign new_n252_ = ~new_n171_ & new_n177_;
  assign new_n253_ = pg2 & new_n161_;
  assign new_n254_ = pg1 & new_n86_;
  assign new_n255_ = ~new_n201_ & ~new_n205_;
  assign new_n256_ = new_n253_ & new_n254_;
  assign new_n257_ = ~new_n255_ & new_n256_;
  assign new_n258_ = pg11 & new_n184_;
  assign new_n259_ = ~pg1 & new_n203_;
  assign new_n260_ = ~pg4 & new_n224_;
  assign new_n261_ = pg6 & new_n260_;
  assign new_n262_ = ~new_n259_ & ~new_n261_;
  assign new_n263_ = pg8 & ~new_n262_;
  assign new_n264_ = pg3 & ~pg1;
  assign new_n265_ = new_n160_ & new_n264_;
  assign new_n266_ = ~pg8 & new_n265_;
  assign new_n267_ = ~new_n263_ & ~new_n266_;
  assign new_n268_ = new_n258_ & ~new_n267_;
  assign new_n269_ = ~pg10 & new_n89_;
  assign new_n270_ = new_n259_ & new_n269_;
  assign new_n271_ = new_n88_ & new_n116_;
  assign new_n272_ = ~new_n262_ & new_n271_;
  assign new_n273_ = ~new_n270_ & ~new_n272_;
  assign new_n274_ = ~pg7 & ~new_n273_;
  assign new_n275_ = ~new_n268_ & ~new_n274_;
  assign new_n276_ = ~pg5 & ~new_n275_;
  assign new_n277_ = pg2 & new_n276_;
  assign new_n278_ = ~new_n257_ & ~new_n277_;
  assign new_n279_ = new_n252_ & new_n278_;
  assign new_n280_ = new_n195_ & new_n219_;
  assign new_n281_ = ~pg12 & new_n280_;
  assign new_n282_ = ~new_n251_ & ~new_n279_;
  assign pg539 = new_n281_ | ~new_n282_;
  assign new_n284_ = pg5 & pg2;
  assign new_n285_ = pg4 & pg3;
  assign new_n286_ = new_n99_ & new_n284_;
  assign new_n287_ = ~new_n285_ & new_n286_;
  assign new_n288_ = pg1 & new_n171_;
  assign new_n289_ = pg2 & new_n103_;
  assign new_n290_ = ~pg5 & ~new_n155_;
  assign new_n291_ = ~pg4 & ~new_n290_;
  assign new_n292_ = ~pg3 & new_n161_;
  assign new_n293_ = ~new_n156_ & ~new_n292_;
  assign new_n294_ = pg5 & ~new_n293_;
  assign new_n295_ = ~new_n289_ & ~new_n291_;
  assign new_n296_ = ~new_n294_ & new_n295_;
  assign new_n297_ = new_n177_ & new_n288_;
  assign new_n298_ = ~new_n296_ & new_n297_;
  assign new_n299_ = pg3 & pg0;
  assign new_n300_ = new_n142_ & new_n144_;
  assign new_n301_ = ~new_n299_ & new_n300_;
  assign new_n302_ = ~new_n85_1_ & ~new_n287_;
  assign new_n303_ = ~new_n298_ & ~new_n301_;
  assign pg549 = ~new_n302_ | ~new_n303_;
  assign new_n305_ = pg6 & new_n142_;
  assign new_n306_ = pg7 & ~pg8;
  assign new_n307_ = ~pg10 & ~new_n306_;
  assign new_n308_ = ~pg9 & ~new_n307_;
  assign new_n309_ = pg7 & pg9;
  assign new_n310_ = new_n125_1_ & ~new_n309_;
  assign new_n311_ = ~new_n271_ & ~new_n308_;
  assign new_n312_ = ~new_n310_ & new_n311_;
  assign new_n313_ = new_n305_ & ~new_n312_;
  assign new_n314_ = pg8 & ng34;
  assign new_n315_ = ~new_n305_ & ~new_n314_;
  assign new_n316_ = new_n92_ & ~new_n315_;
  assign new_n317_ = pg9 & pg8;
  assign new_n318_ = ng34 & new_n87_;
  assign new_n319_ = ~new_n317_ & new_n318_;
  assign new_n320_ = ~new_n313_ & ~new_n316_;
  assign pg542 = new_n319_ | ~new_n320_;
  assign new_n322_ = new_n189_ & new_n258_;
  assign new_n323_ = ~new_n160_ & ~new_n322_;
  assign new_n324_ = new_n220_ & ~new_n323_;
  assign new_n325_ = ~pg3 & new_n324_;
  assign new_n326_ = new_n203_ & new_n220_;
  assign new_n327_ = pg13 & ~new_n278_;
  assign new_n328_ = ~new_n326_ & ~new_n327_;
  assign new_n329_ = new_n271_ & ~new_n328_;
  assign new_n330_ = ~ng43 & new_n171_;
  assign new_n331_ = pg13 & new_n330_;
  assign new_n332_ = ~pg4 & ~new_n188_;
  assign new_n333_ = ~new_n202_ & ~new_n332_;
  assign new_n334_ = ~new_n220_ & ~new_n327_;
  assign new_n335_ = pg6 & ~new_n333_;
  assign new_n336_ = ~new_n334_ & new_n335_;
  assign new_n337_ = ~new_n325_ & ~new_n329_;
  assign new_n338_ = ~new_n331_ & ~new_n336_;
  assign new_n339_ = new_n337_ & new_n338_;
  assign new_n340_ = ~pg12 & ~new_n339_;
  assign new_n341_ = pg2 & ~new_n224_;
  assign new_n342_ = ~pg2 & new_n86_;
  assign new_n343_ = ~pg5 & ~pg3;
  assign new_n344_ = ~new_n341_ & ~new_n342_;
  assign new_n345_ = ~new_n343_ & new_n344_;
  assign new_n346_ = pg4 & ~new_n345_;
  assign new_n347_ = ~pg3 & ~pg2;
  assign new_n348_ = pg1 & new_n347_;
  assign new_n349_ = ~new_n260_ & ~new_n346_;
  assign new_n350_ = ~new_n348_ & new_n349_;
  assign new_n351_ = new_n142_ & ~new_n350_;
  assign new_n352_ = pg0 & new_n351_;
  assign pg532 = new_n340_ | new_n352_;
  assign new_n354_ = ~new_n188_ & new_n203_;
  assign new_n355_ = new_n88_ & new_n189_;
  assign new_n356_ = pg10 & new_n355_;
  assign new_n357_ = ~pg5 & new_n160_;
  assign new_n358_ = new_n133_ & new_n357_;
  assign new_n359_ = ~new_n356_ & ~new_n358_;
  assign new_n360_ = new_n121_ & ~new_n359_;
  assign new_n361_ = ~pg6 & new_n87_;
  assign new_n362_ = new_n103_ & new_n361_;
  assign new_n363_ = new_n89_ & new_n362_;
  assign new_n364_ = ~new_n360_ & ~new_n363_;
  assign new_n365_ = ~new_n354_ & new_n364_;
  assign new_n366_ = new_n221_ & ~new_n365_;
  assign new_n367_ = new_n235_ & new_n250_;
  assign new_n368_ = new_n254_ & new_n367_;
  assign new_n369_ = ng38 & new_n240_;
  assign new_n370_ = ~new_n87_ & ~new_n369_;
  assign new_n371_ = new_n368_ & ~new_n370_;
  assign new_n372_ = new_n327_ & new_n354_;
  assign new_n373_ = pg6 & new_n184_;
  assign new_n374_ = ~new_n86_ & ~new_n373_;
  assign new_n375_ = ~new_n334_ & ~new_n374_;
  assign new_n376_ = pg8 & new_n375_;
  assign new_n377_ = ~new_n372_ & ~new_n376_;
  assign new_n378_ = ~pg12 & ~new_n377_;
  assign new_n379_ = ~new_n371_ & ~new_n378_;
  assign new_n380_ = pg2 & ~new_n379_;
  assign pg537 = new_n366_ | new_n380_;
  assign new_n382_ = ~new_n91_ & new_n93_;
  assign new_n383_ = ~pg9 & new_n87_;
  assign new_n384_ = ~new_n382_ & ~new_n383_;
  assign new_n385_ = pg11 & ~new_n384_;
  assign new_n386_ = pg7 & ~new_n125_1_;
  assign new_n387_ = new_n88_ & new_n386_;
  assign new_n388_ = ~new_n385_ & ~new_n387_;
  assign new_n389_ = ng34 & ~new_n388_;
  assign new_n390_ = ~ng42 & new_n142_;
  assign pg548 = new_n389_ | new_n390_;
  assign new_n392_ = pg2 & pg0;
  assign new_n393_ = pg4 & new_n392_;
  assign new_n394_ = pg1 & ~new_n392_;
  assign new_n395_ = ~new_n393_ & ~new_n394_;
  assign new_n396_ = ~pg3 & ~new_n395_;
  assign new_n397_ = ~new_n144_ & new_n299_;
  assign new_n398_ = ~new_n145_1_ & ~new_n396_;
  assign new_n399_ = ~new_n397_ & new_n398_;
  assign new_n400_ = new_n142_ & ~new_n399_;
  assign new_n401_ = pg5 & new_n400_;
  assign new_n402_ = pg6 & new_n156_;
  assign new_n403_ = ~pg5 & new_n402_;
  assign new_n404_ = ~new_n103_ & ~new_n292_;
  assign new_n405_ = ~new_n403_ & new_n404_;
  assign new_n406_ = new_n288_ & ~new_n405_;
  assign new_n407_ = new_n156_ & new_n172_;
  assign new_n408_ = new_n100_1_ & new_n171_;
  assign new_n409_ = ~pg1 & new_n408_;
  assign new_n410_ = ~new_n407_ & ~new_n409_;
  assign new_n411_ = ~new_n406_ & new_n410_;
  assign new_n412_ = new_n177_ & ~new_n411_;
  assign new_n413_ = ng39 & new_n99_;
  assign new_n414_ = pg4 & new_n413_;
  assign new_n415_ = ~new_n401_ & ~new_n412_;
  assign pg551 = new_n414_ | ~new_n415_;
  assign new_n417_ = ~pg10 & pg11;
  assign new_n418_ = pg9 & pg10;
  assign new_n419_ = ~new_n417_ & ~new_n418_;
  assign new_n420_ = new_n93_ & ~new_n419_;
  assign new_n421_ = new_n91_ & ~new_n93_;
  assign new_n422_ = ~pg8 & new_n88_;
  assign new_n423_ = ~new_n420_ & ~new_n421_;
  assign new_n424_ = ~new_n422_ & new_n423_;
  assign new_n425_ = pg6 & ~new_n424_;
  assign new_n426_ = pg9 & new_n361_;
  assign new_n427_ = ~new_n425_ & ~new_n426_;
  assign new_n428_ = new_n142_ & ~new_n427_;
  assign new_n429_ = ~pg7 & new_n125_1_;
  assign new_n430_ = ~new_n386_ & ~new_n429_;
  assign new_n431_ = ng34 & ~new_n430_;
  assign new_n432_ = pg9 & new_n431_;
  assign pg547 = new_n428_ | new_n432_;
  assign new_n434_ = ~ng40 & new_n142_;
  assign new_n435_ = pg5 & ~pg4;
  assign new_n436_ = ~new_n103_ & ~new_n435_;
  assign new_n437_ = pg6 & ~new_n436_;
  assign new_n438_ = ~new_n292_ & ~new_n437_;
  assign new_n439_ = pg2 & ~new_n438_;
  assign new_n440_ = ~new_n103_ & new_n402_;
  assign new_n441_ = ~new_n439_ & ~new_n440_;
  assign new_n442_ = new_n99_ & ~new_n441_;
  assign new_n443_ = pg2 & ~new_n144_;
  assign new_n444_ = ~new_n86_ & ~new_n443_;
  assign new_n445_ = pg6 & ~new_n444_;
  assign new_n446_ = new_n161_ & ~new_n284_;
  assign new_n447_ = ~new_n445_ & ~new_n446_;
  assign new_n448_ = new_n177_ & ~new_n447_;
  assign new_n449_ = new_n171_ & new_n448_;
  assign new_n450_ = ~new_n434_ & ~new_n442_;
  assign pg552 = new_n449_ | ~new_n450_;
  assign new_n452_ = ~pg3 & ~ng44;
  assign new_n453_ = ~new_n91_ & ~new_n184_;
  assign new_n454_ = new_n215_ & ~new_n453_;
  assign new_n455_ = ~new_n452_ & ~new_n454_;
  assign new_n456_ = new_n221_ & ~new_n455_;
  assign new_n457_ = new_n332_ & ~new_n334_;
  assign new_n458_ = new_n327_ & ~new_n453_;
  assign new_n459_ = new_n103_ & new_n458_;
  assign new_n460_ = ~new_n457_ & ~new_n459_;
  assign new_n461_ = pg6 & ~new_n460_;
  assign new_n462_ = ~pg12 & new_n461_;
  assign new_n463_ = ng38 & new_n368_;
  assign new_n464_ = ng37 & new_n463_;
  assign new_n465_ = ~new_n462_ & ~new_n464_;
  assign pg535 = new_n456_ | ~new_n465_;
  assign n60 = new_n110_1_ & new_n183_;
  assign new_n468_ = ~pg13 & ng32;
  assign new_n469_ = pg13 & ~new_n170_;
  assign new_n470_ = ~new_n468_ & ~new_n469_;
  assign new_n471_ = ~pg12 & ~new_n96_;
  assign n65 = ~new_n470_ & new_n471_;
  assign new_n473_ = pg6 & ~new_n188_;
  assign new_n474_ = ~pg8 & new_n184_;
  assign new_n475_ = ~pg6 & new_n474_;
  assign n70 = new_n473_ | new_n475_;
  assign new_n477_ = ~pg10 & new_n200_;
  assign new_n478_ = ~new_n205_ & ~new_n477_;
  assign n75 = ~pg5 & ~new_n478_;
  assign new_n480_ = ~pg6 & pg9;
  assign n80 = new_n240_ | new_n480_;
  assign new_n482_ = ~pg9 & pg11;
  assign n85 = pg10 | new_n482_;
  assign new_n484_ = ~pg7 & pg11;
  assign new_n485_ = pg10 & ~new_n88_;
  assign n90 = new_n484_ | new_n485_;
  assign new_n487_ = ~new_n153_ & new_n156_;
  assign new_n488_ = ~new_n203_ & new_n284_;
  assign new_n489_ = ~new_n289_ & ~new_n487_;
  assign n95 = new_n488_ | ~new_n489_;
  assign new_n491_ = new_n98_ & new_n289_;
  assign new_n492_ = ~pg4 & pg1;
  assign new_n493_ = new_n141_ & new_n492_;
  assign new_n494_ = pg0 & new_n493_;
  assign n100 = ~new_n491_ & ~new_n494_;
  assign new_n496_ = ~new_n285_ & ~new_n435_;
  assign new_n497_ = new_n151_ & ~new_n496_;
  assign new_n498_ = ~new_n103_ & new_n156_;
  assign n105 = ~new_n497_ & ~new_n498_;
  assign new_n500_ = pg2 & ~new_n86_;
  assign n110 = new_n342_ | new_n500_;
  assign new_n502_ = pg6 & new_n269_;
  assign new_n503_ = pg6 & ng31;
  assign new_n504_ = ~pg6 & ng30;
  assign new_n505_ = pg6 & pg9;
  assign new_n506_ = ~pg11 & new_n505_;
  assign new_n507_ = ~new_n504_ & ~new_n506_;
  assign new_n508_ = pg7 & ~new_n507_;
  assign new_n509_ = ~new_n503_ & ~new_n508_;
  assign new_n510_ = pg8 & ~new_n509_;
  assign n115 = ~new_n502_ & ~new_n510_;
  assign new_n512_ = ng34 & new_n310_;
  assign new_n513_ = new_n87_ & new_n142_;
  assign new_n514_ = ~new_n505_ & new_n513_;
  assign new_n515_ = ~new_n316_ & ~new_n512_;
  assign n120 = ~new_n514_ & new_n515_;
  assign new_n517_ = pg6 & new_n125_1_;
  assign new_n518_ = ~new_n306_ & ~new_n517_;
  assign new_n519_ = ~pg9 & ~new_n518_;
  assign new_n520_ = pg7 & ~new_n91_;
  assign new_n521_ = ~pg6 & new_n520_;
  assign new_n522_ = ~new_n519_ & ~new_n521_;
  assign new_n523_ = pg11 & ~new_n522_;
  assign new_n524_ = ~new_n87_ & new_n88_;
  assign new_n525_ = pg6 & new_n524_;
  assign n125 = ~new_n523_ & ~new_n525_;
  assign new_n527_ = pg6 & new_n103_;
  assign new_n528_ = pg5 & ~new_n161_;
  assign new_n529_ = ~pg6 & new_n100_1_;
  assign new_n530_ = ~new_n527_ & ~new_n528_;
  assign new_n531_ = ~new_n529_ & new_n530_;
  assign new_n532_ = new_n224_ & ~new_n531_;
  assign new_n533_ = pg3 & new_n154_;
  assign new_n534_ = pg1 & new_n402_;
  assign new_n535_ = ~new_n532_ & ~new_n533_;
  assign n130 = ~new_n534_ & new_n535_;
  assign new_n537_ = ~pg6 & new_n134_;
  assign new_n538_ = ~pg5 & new_n537_;
  assign new_n539_ = ~new_n356_ & ~new_n538_;
  assign new_n540_ = new_n121_ & ~new_n539_;
  assign new_n541_ = new_n205_ & new_n357_;
  assign n135 = ~new_n540_ & ~new_n541_;
  assign new_n543_ = new_n252_ & ~new_n278_;
  assign new_n544_ = ~new_n367_ & ~new_n543_;
  assign n140 = new_n221_ | ~new_n544_;
  assign new_n546_ = ~new_n103_ & new_n108_;
  assign new_n547_ = new_n103_ & new_n156_;
  assign new_n548_ = pg0 & ~new_n546_;
  assign new_n549_ = ~new_n547_ & new_n548_;
  assign new_n550_ = ~pg1 & ~new_n549_;
  assign new_n551_ = ~pg7 & ~pg6;
  assign new_n552_ = ~pg10 & new_n120_1_;
  assign new_n553_ = ~pg3 & pg0;
  assign new_n554_ = pg4 & pg0;
  assign new_n555_ = ~new_n264_ & ~new_n553_;
  assign new_n556_ = ~new_n554_ & new_n555_;
  assign new_n557_ = new_n106_ & ~new_n556_;
  assign new_n558_ = pg2 & new_n557_;
  assign new_n559_ = ~new_n550_ & ~new_n551_;
  assign new_n560_ = ~new_n552_ & new_n559_;
  assign n145 = ~new_n558_ & new_n560_;
  assign pg546 = ~ng41;
  assign pg45 = ng45;
  always @ (posedge clock) begin
    ng38 <= n60;
    ng34 <= n65;
    ng35 <= n70;
    ng36 <= n75;
    ng37 <= n80;
    ng30 <= n85;
    ng31 <= n90;
    ng32 <= n95;
    ng33 <= n100;
    ng29 <= n105;
    ng39 <= n110;
    ng40 <= n115;
    ng41 <= n120;
    ng42 <= n125;
    ng43 <= n130;
    ng44 <= n135;
    ng45 <= n140;
    ng46 <= n145;
  end
endmodule

