module top ( clock, 
    pn3083gat, pn3084gat, pn3081gat, pn3082gat, pn3099gat, pn3087gat,
    pn3088gat, pn3070gat, pn3085gat, pn3086gat, pn3094gat, pn3093gat,
    pn3089gat, pn3092gat, pn3091gat, pn3098gat, pn3097gat, pn3095gat,
    pn3079gat, pclk, pn3065gat, pn3090gat, pn3066gat, pn3067gat, pn3068gat,
    pn3069gat, pn3072gat, pn3071gat, pn3074gat, pn3100gat, pn3073gat,
    pn3076gat, pn3075gat, pn3080gat, pn3078gat, pn3077gat,
    pn3113gat, pn3112gat, pn3111gat, pn3110gat, pn3117gat, pn3128gat,
    pn3116gat, pn3129gat, pn3152gat, pn3115gat, pn3151gat, pn3114gat,
    pn3150gat, pn3124gat, pn3125gat, pn3119gat, pn3126gat, pn3118gat,
    pn3127gat, pn3120gat, pn3121gat, pn3122gat, pn3123gat, pn3135gat,
    pn3134gat, pn3108gat, pn3137gat, pn3109gat, pn3136gat, pn3131gat,
    pn3130gat, pn3133gat, pn3148gat, pn3132gat, pn3149gat, pn3146gat,
    pn3147gat, pn3144gat, pn3145gat, pn3106gat, pn3139gat, pn3142gat,
    pn3107gat, pn3138gat, pn3143gat, pn3104gat, pn3140gat, pn3105gat,
    pn3141gat  );
  input  clock;
  input  pn3083gat, pn3084gat, pn3081gat, pn3082gat, pn3099gat,
    pn3087gat, pn3088gat, pn3070gat, pn3085gat, pn3086gat, pn3094gat,
    pn3093gat, pn3089gat, pn3092gat, pn3091gat, pn3098gat, pn3097gat,
    pn3095gat, pn3079gat, pclk, pn3065gat, pn3090gat, pn3066gat, pn3067gat,
    pn3068gat, pn3069gat, pn3072gat, pn3071gat, pn3074gat, pn3100gat,
    pn3073gat, pn3076gat, pn3075gat, pn3080gat, pn3078gat, pn3077gat;
  output pn3113gat, pn3112gat, pn3111gat, pn3110gat, pn3117gat, pn3128gat,
    pn3116gat, pn3129gat, pn3152gat, pn3115gat, pn3151gat, pn3114gat,
    pn3150gat, pn3124gat, pn3125gat, pn3119gat, pn3126gat, pn3118gat,
    pn3127gat, pn3120gat, pn3121gat, pn3122gat, pn3123gat, pn3135gat,
    pn3134gat, pn3108gat, pn3137gat, pn3109gat, pn3136gat, pn3131gat,
    pn3130gat, pn3133gat, pn3148gat, pn3132gat, pn3149gat, pn3146gat,
    pn3147gat, pn3144gat, pn3145gat, pn3106gat, pn3139gat, pn3142gat,
    pn3107gat, pn3138gat, pn3143gat, pn3104gat, pn3140gat, pn3105gat,
    pn3141gat;
  reg nn1332gat, nn1775gat, nn2454gat, nn2117gat, nn470gat, nn1525gat,
    nn1740gat, nn1312gat, nn2040gat, nn2121gat, nn148gat, nn1456gat,
    nn2179gat, nn2592gat, nn2176gat, nn2125gat, nn2190gat, nn1871gat,
    nn2169gat, nn2110gat, nn842gat, nn2021gat, nn1433gat, nn2446gat,
    nn2033gat, nn1394gat, nn2182gat, nn2095gat, nn2266gat, nn1496gat,
    nn1363gat, nn2309gat, nn2099gat, nn2091gat, nn1316gat, nn2450gat,
    nn2025gat, nn2510gat, nn156gat, nn2514gat, nn1588gat, nn271gat,
    nn152gat, nn2458gat, nn160gat, nn331gat, nn1336gat, nn1462gat,
    nn337gat, nn388gat, nn1771gat, nn1596gat, nn398gat, nn2135gat,
    nn1678gat, nn463gat, nn1675gat, nn402gat, nn2262gat, nn1508gat,
    nn327gat, nn1748gat, nn919gat, nn2044gat, nn2644gat, nn384gat,
    nn1340gat, nn846gat, nn2037gat, nn1975gat, nn256gat, nn1807gat,
    nn2630gat, nn931gat, nn322gat, nn2502gat, nn2403gat, nn2543gat,
    nn1226gat, nn318gat, nn2339gat, nn2394gat, nn2102gat, nn1045gat,
    nn561gat, nn2270gat, nn2440gat, nn673gat, nn1880gat, nn1135gat,
    nn366gat, nn2390gat, nn2407gat, nn341gat, nn1241gat, nn680gat,
    nn2343gat, nn2347gat, nn2472gat, nn1294gat, nn816gat, nn2399gat,
    nn1389gat, nn2319gat, nn1080gat, nn614gat, nn2464gat, nn1821gat,
    nn865gat, nn2526gat, nn699gat, nn2029gat, nn2468gat, nn820gat,
    nn2626gat, nn1072gat, nn777gat, nn1829gat, nn1148gat, nn883gat,
    nn2207gat, nn1282gat, nn553gat, nn2476gat, nn707gat, nn580gat,
    nn2562gat, nn2658gat, nn2143gat, nn1068gat, nn834gat, nn824gat,
    nn2203gat, nn2495gat, nn2084gat, nn957gat, nn830gat, nn1763gat,
    nn2518gat, nn2588gat, nn1767gat, nn2061gat, nn861gat, nn838gat,
    nn2155gat, nn1197gat, nn2640gat, nn1834gat, nn2139gat, nn584gat,
    nn2622gat, nn1035gat, nn659gat, nn314gat, nn2506gat, nn1899gat,
    nn684gat, nn2490gat, nn1121gat, nn667gat, nn2599gat, nn2634gat,
    nn1850gat;
  wire new_n576_, new_n577_1_, new_n578_, new_n579_, new_n581_, new_n582_1_,
    new_n583_, new_n584_, new_n586_, new_n587_1_, new_n588_, new_n589_,
    new_n591_, new_n592_1_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_1_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_1_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_1_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_1_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_1_, new_n619_, new_n620_, new_n621_,
    new_n622_1_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_1_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_1_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_1_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_1_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_1_, new_n648_, new_n649_, new_n650_, new_n652_1_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_1_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_1_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_1_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_1_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_1_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_1_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_1_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_1_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_1_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_1_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_1_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_1_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_1_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_1_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_1_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_1_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_1_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_1_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_1_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_1_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_1_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_1_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_1_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_1_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_1_, new_n788_, new_n790_, new_n791_, new_n792_1_, new_n793_,
    new_n795_, new_n796_, new_n797_1_, new_n798_, new_n799_, new_n801_,
    new_n802_1_, new_n804_, new_n805_, new_n806_, new_n807_1_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_1_, new_n813_, new_n815_,
    new_n816_, new_n817_1_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_1_, new_n823_, new_n825_, new_n827_1_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_1_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_1_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_1_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_1_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_1_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_1_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_1_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_1_, new_n868_, new_n869_, new_n871_, new_n872_1_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_1_, new_n878_,
    new_n880_, new_n881_, new_n882_1_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_1_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_1_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_1_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_1_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_1_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_1_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_1_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_1_, new_n924_, new_n925_, new_n926_, new_n927_1_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_1_, new_n938_, new_n939_, new_n940_, new_n942_1_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_1_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_1_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_1_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_1_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_1_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_1_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_1_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_1_, new_n983_, new_n984_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1044_, new_n1045_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1109_, new_n1110_, new_n1111_,
    new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1133_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_,
    new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_,
    new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_,
    new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1335_, new_n1336_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1441_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1546_, new_n1547_, new_n1548_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1557_, new_n1558_, new_n1559_,
    new_n1561_, new_n1563_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1610_, new_n1611_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1624_, new_n1625_,
    new_n1626_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1635_,
    new_n1636_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1644_,
    new_n1647_, new_n1648_, new_n1649_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1681_, new_n1683_,
    new_n1684_, new_n1685_, new_n1689_, new_n1691_, new_n1692_, new_n1693_,
    new_n1696_, new_n1697_, new_n1699_, new_n1701_, new_n1703_, new_n1704_,
    new_n1705_, new_n1707_, new_n1708_, new_n1710_, new_n1711_, new_n1712_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1721_, new_n1722_,
    new_n1724_, new_n1725_, new_n1728_, new_n1729_, new_n1731_, new_n1732_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1745_, new_n1746_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1774_,
    new_n1776_, new_n1777_, new_n1778_, new_n1780_, new_n1781_, new_n1783_,
    new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1791_,
    new_n1793_, new_n1794_, new_n1795_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1806_,
    new_n1807_, new_n1809_, new_n1810_, new_n1812_, new_n1813_, new_n1814_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_,
    new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1835_,
    new_n1836_, new_n1837_, new_n1839_, new_n1840_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_,
    new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_,
    new_n1859_, new_n1860_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1868_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1874_, new_n1875_, new_n1877_, new_n1878_, new_n1881_, new_n1883_,
    new_n1884_, new_n1885_, new_n1887_, new_n1888_, new_n1889_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_,
    new_n1900_, new_n1902_, new_n1903_, new_n1904_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, n172, n177, n182, n187,
    n192, n197, n202, n207, n212, n217, n222, n227, n232, n237, n242, n247,
    n252, n257, n262, n267, n272, n277, n282, n287, n292, n297, n302, n307,
    n312, n317, n322, n327, n332, n337, n342, n347, n352, n357, n362, n367,
    n372, n377, n382, n387, n392, n397, n402, n407, n412, n417, n422, n427,
    n432, n437, n442, n447, n452, n457, n462, n467, n472, n477, n482, n487,
    n492, n497, n502, n507, n512, n517, n522, n527, n532, n537, n542, n547,
    n552, n557, n562, n567, n572, n577, n582, n587, n592, n597, n602, n607,
    n612, n617, n622, n627, n632, n637, n642, n647, n652, n657, n662, n667,
    n672, n677, n682, n687, n692, n697, n702, n707, n712, n717, n722, n727,
    n732, n737, n742, n747, n752, n757, n762, n767, n772, n777, n782, n787,
    n792, n797, n802, n807, n812, n817, n822, n827, n832, n837, n842, n847,
    n852, n857, n862, n867, n872, n877, n882, n887, n892, n897, n902, n907,
    n912, n917, n922, n927, n932, n937, n942, n947, n952, n957, n962, n967,
    n972, n977, n982;
  assign new_n576_ = ~nn2190gat & ~nn2262gat;
  assign new_n577_1_ = ~nn2135gat & ~new_n576_;
  assign new_n578_ = nn2135gat & new_n576_;
  assign new_n579_ = ~new_n577_1_ & ~new_n578_;
  assign pn3113gat = ~nn1135gat | ~new_n579_;
  assign new_n581_ = nn2394gat & ~nn2440gat;
  assign new_n582_1_ = ~nn2394gat & nn2440gat;
  assign new_n583_ = nn2394gat & ~new_n581_;
  assign new_n584_ = ~new_n582_1_ & new_n583_;
  assign pn3111gat = ~nn931gat | ~new_n584_;
  assign new_n586_ = ~nn2394gat & ~nn2440gat;
  assign new_n587_1_ = nn2403gat & new_n586_;
  assign new_n588_ = ~nn2403gat & ~new_n586_;
  assign new_n589_ = ~new_n587_1_ & ~new_n588_;
  assign pn3110gat = ~nn1121gat | ~new_n589_;
  assign new_n591_ = pn3088gat & ~pn3089gat;
  assign new_n592_1_ = ~pn3088gat & pn3089gat;
  assign new_n593_ = ~new_n591_ & ~new_n592_1_;
  assign new_n594_ = pn3087gat & ~pn3086gat;
  assign new_n595_ = ~pn3087gat & pn3086gat;
  assign new_n596_ = ~new_n594_ & ~new_n595_;
  assign new_n597_1_ = pn3084gat & ~pn3085gat;
  assign new_n598_ = ~pn3083gat & new_n597_1_;
  assign new_n599_ = ~pn3084gat & ~pn3085gat;
  assign new_n600_ = pn3083gat & new_n599_;
  assign new_n601_ = ~pn3084gat & pn3085gat;
  assign new_n602_1_ = ~pn3083gat & new_n601_;
  assign new_n603_ = pn3084gat & pn3085gat;
  assign new_n604_ = pn3083gat & new_n603_;
  assign new_n605_ = ~new_n598_ & ~new_n600_;
  assign new_n606_ = ~new_n602_1_ & ~new_n604_;
  assign new_n607_1_ = new_n605_ & new_n606_;
  assign new_n608_ = ~new_n593_ & ~new_n596_;
  assign new_n609_ = new_n607_1_ & new_n608_;
  assign new_n610_ = ~new_n593_ & new_n596_;
  assign new_n611_ = ~new_n607_1_ & new_n610_;
  assign new_n612_1_ = new_n593_ & new_n596_;
  assign new_n613_ = new_n607_1_ & new_n612_1_;
  assign new_n614_ = new_n593_ & ~new_n596_;
  assign new_n615_ = ~new_n607_1_ & new_n614_;
  assign new_n616_ = ~new_n609_ & ~new_n611_;
  assign new_n617_1_ = ~new_n613_ & ~new_n615_;
  assign n357 = ~new_n616_ | ~new_n617_1_;
  assign new_n619_ = pn3086gat & pn3095gat;
  assign new_n620_ = pn3087gat & pn3095gat;
  assign new_n621_ = ~new_n619_ & ~new_n620_;
  assign new_n622_1_ = pn3083gat & pn3095gat;
  assign new_n623_ = pn3084gat & pn3095gat;
  assign new_n624_ = pn3085gat & pn3095gat;
  assign new_n625_ = ~new_n622_1_ & ~new_n623_;
  assign new_n626_ = ~new_n624_ & new_n625_;
  assign new_n627_1_ = ~new_n621_ & new_n626_;
  assign new_n628_ = pn3085gat & pn3093gat;
  assign new_n629_ = ~new_n619_ & ~new_n628_;
  assign new_n630_ = pn3086gat & pn3093gat;
  assign new_n631_ = ~new_n620_ & ~new_n630_;
  assign new_n632_1_ = pn3088gat & pn3095gat;
  assign new_n633_ = pn3087gat & pn3093gat;
  assign new_n634_ = ~new_n632_1_ & ~new_n633_;
  assign new_n635_ = ~new_n629_ & new_n631_;
  assign new_n636_ = ~new_n634_ & new_n635_;
  assign new_n637_1_ = ~nn680gat & new_n636_;
  assign new_n638_ = ~new_n631_ & ~new_n634_;
  assign new_n639_ = new_n629_ & new_n638_;
  assign new_n640_ = ~nn1068gat & new_n639_;
  assign new_n641_ = ~new_n629_ & new_n634_;
  assign new_n642_1_ = ~new_n631_ & new_n641_;
  assign new_n643_ = ~nn659gat & new_n642_1_;
  assign new_n644_ = ~new_n629_ & ~new_n634_;
  assign new_n645_ = ~new_n631_ & new_n644_;
  assign new_n646_ = ~nn271gat & new_n645_;
  assign new_n647_1_ = ~new_n637_1_ & ~new_n640_;
  assign new_n648_ = ~new_n643_ & ~new_n646_;
  assign new_n649_ = new_n647_1_ & new_n648_;
  assign new_n650_ = new_n627_1_ & ~new_n649_;
  assign pn3117gat = ~n357 | new_n650_;
  assign new_n652_1_ = nn1226gat & ~nn1282gat;
  assign new_n653_ = ~nn1226gat & nn1282gat;
  assign new_n654_ = ~new_n652_1_ & ~new_n653_;
  assign new_n655_ = ~nn1045gat & nn1135gat;
  assign new_n656_ = nn931gat & new_n655_;
  assign new_n657_1_ = nn1045gat & nn1135gat;
  assign new_n658_ = ~nn931gat & new_n657_1_;
  assign new_n659_ = nn1045gat & ~nn1135gat;
  assign new_n660_ = nn931gat & new_n659_;
  assign new_n661_ = ~nn1045gat & ~nn1135gat;
  assign new_n662_1_ = ~nn931gat & new_n661_;
  assign new_n663_ = ~new_n656_ & ~new_n658_;
  assign new_n664_ = ~new_n660_ & ~new_n662_1_;
  assign new_n665_ = new_n663_ & new_n664_;
  assign new_n666_ = ~nn1072gat & nn1121gat;
  assign new_n667_1_ = nn1035gat & new_n666_;
  assign new_n668_ = nn1072gat & nn1121gat;
  assign new_n669_ = ~nn1035gat & new_n668_;
  assign new_n670_ = nn1072gat & ~nn1121gat;
  assign new_n671_ = nn1035gat & new_n670_;
  assign new_n672_1_ = ~nn1072gat & ~nn1121gat;
  assign new_n673_ = ~nn1035gat & new_n672_1_;
  assign new_n674_ = ~new_n667_1_ & ~new_n669_;
  assign new_n675_ = ~new_n671_ & ~new_n673_;
  assign new_n676_ = new_n674_ & new_n675_;
  assign new_n677_1_ = ~new_n654_ & ~new_n665_;
  assign new_n678_ = new_n676_ & new_n677_1_;
  assign new_n679_ = ~new_n654_ & new_n665_;
  assign new_n680_ = ~new_n676_ & new_n679_;
  assign new_n681_ = new_n654_ & new_n665_;
  assign new_n682_1_ = new_n676_ & new_n681_;
  assign new_n683_ = new_n654_ & ~new_n665_;
  assign new_n684_ = ~new_n676_ & new_n683_;
  assign new_n685_ = ~new_n678_ & ~new_n680_;
  assign new_n686_ = ~new_n682_1_ & ~new_n684_;
  assign pn3116gat = ~new_n685_ | ~new_n686_;
  assign new_n688_ = ~nn842gat & new_n639_;
  assign new_n689_ = ~nn830gat & new_n636_;
  assign new_n690_ = ~new_n688_ & ~new_n689_;
  assign new_n691_ = new_n642_1_ & pn3116gat;
  assign new_n692_1_ = new_n690_ & ~new_n691_;
  assign new_n693_ = pn3088gat & pn3093gat;
  assign new_n694_ = new_n630_ & new_n693_;
  assign new_n695_ = new_n628_ & new_n694_;
  assign new_n696_ = new_n633_ & new_n695_;
  assign new_n697_1_ = ~new_n628_ & ~new_n630_;
  assign new_n698_ = pn3083gat & pn3093gat;
  assign new_n699_ = pn3084gat & pn3093gat;
  assign new_n700_ = ~new_n698_ & ~new_n699_;
  assign new_n701_ = ~new_n696_ & ~new_n697_1_;
  assign new_n702_1_ = new_n700_ & new_n701_;
  assign new_n703_ = new_n693_ & new_n702_1_;
  assign new_n704_ = ~new_n627_1_ & ~new_n703_;
  assign new_n705_ = ~new_n692_1_ & ~new_n704_;
  assign new_n706_ = new_n620_ & new_n632_1_;
  assign new_n707_1_ = new_n619_ & new_n706_;
  assign new_n708_ = new_n626_ & new_n707_1_;
  assign new_n709_ = ~new_n693_ & new_n702_1_;
  assign new_n710_ = ~new_n708_ & ~new_n709_;
  assign new_n711_ = ~nn561gat & nn366gat;
  assign new_n712_1_ = nn561gat & ~nn366gat;
  assign new_n713_ = ~new_n711_ & ~new_n712_1_;
  assign new_n714_ = nn318gat & ~nn314gat;
  assign new_n715_ = nn322gat & new_n714_;
  assign new_n716_ = nn318gat & nn314gat;
  assign new_n717_1_ = ~nn322gat & new_n716_;
  assign new_n718_ = ~nn318gat & nn314gat;
  assign new_n719_ = nn322gat & new_n718_;
  assign new_n720_ = ~nn318gat & ~nn314gat;
  assign new_n721_ = ~nn322gat & new_n720_;
  assign new_n722_1_ = ~new_n715_ & ~new_n717_1_;
  assign new_n723_ = ~new_n719_ & ~new_n721_;
  assign new_n724_ = new_n722_1_ & new_n723_;
  assign new_n725_ = ~nn777gat & nn553gat;
  assign new_n726_ = nn659gat & new_n725_;
  assign new_n727_1_ = nn777gat & nn553gat;
  assign new_n728_ = ~nn659gat & new_n727_1_;
  assign new_n729_ = nn777gat & ~nn553gat;
  assign new_n730_ = nn659gat & new_n729_;
  assign new_n731_ = ~nn777gat & ~nn553gat;
  assign new_n732_1_ = ~nn659gat & new_n731_;
  assign new_n733_ = ~new_n726_ & ~new_n728_;
  assign new_n734_ = ~new_n730_ & ~new_n732_1_;
  assign new_n735_ = new_n733_ & new_n734_;
  assign new_n736_ = ~new_n713_ & ~new_n724_;
  assign new_n737_1_ = new_n735_ & new_n736_;
  assign new_n738_ = ~new_n713_ & new_n724_;
  assign new_n739_ = ~new_n735_ & new_n738_;
  assign new_n740_ = new_n713_ & new_n724_;
  assign new_n741_ = new_n735_ & new_n740_;
  assign new_n742_1_ = new_n713_ & ~new_n724_;
  assign new_n743_ = ~new_n735_ & new_n742_1_;
  assign new_n744_ = ~new_n737_1_ & ~new_n739_;
  assign new_n745_ = ~new_n741_ & ~new_n743_;
  assign new_n746_ = new_n744_ & new_n745_;
  assign new_n747_1_ = new_n642_1_ & ~new_n746_;
  assign new_n748_ = ~nn1241gat & new_n639_;
  assign new_n749_ = ~nn842gat & new_n645_;
  assign new_n750_ = ~nn820gat & new_n636_;
  assign new_n751_ = ~new_n747_1_ & ~new_n748_;
  assign new_n752_1_ = ~new_n749_ & ~new_n750_;
  assign new_n753_ = new_n751_ & new_n752_1_;
  assign new_n754_ = new_n631_ & new_n634_;
  assign new_n755_ = ~new_n629_ & new_n754_;
  assign new_n756_ = new_n629_ & new_n634_;
  assign new_n757_1_ = ~new_n631_ & new_n756_;
  assign new_n758_ = nn673gat & new_n757_1_;
  assign new_n759_ = ~new_n755_ & ~new_n758_;
  assign new_n760_ = new_n753_ & new_n759_;
  assign new_n761_ = ~new_n710_ & ~new_n760_;
  assign pn3129gat = new_n705_ | new_n761_;
  assign new_n763_ = ~pn3083gat & ~pn3084gat;
  assign new_n764_ = ~pn3085gat & new_n763_;
  assign new_n765_ = nn1871gat & new_n764_;
  assign new_n766_ = pn3095gat & new_n765_;
  assign new_n767_1_ = pn3086gat & new_n766_;
  assign new_n768_ = pn3088gat & new_n766_;
  assign new_n769_ = pn3087gat & new_n766_;
  assign new_n770_ = new_n767_1_ & ~new_n768_;
  assign new_n771_ = ~new_n769_ & new_n770_;
  assign new_n772_1_ = pn3085gat & ~pn3086gat;
  assign new_n773_ = ~pn3087gat & pn3088gat;
  assign new_n774_ = ~pn3084gat & pn3093gat;
  assign new_n775_ = ~pn3083gat & new_n774_;
  assign new_n776_ = nn1871gat & new_n775_;
  assign new_n777_1_ = new_n772_1_ & new_n773_;
  assign new_n778_ = new_n776_ & new_n777_1_;
  assign new_n779_ = ~nn2139gat & nn1899gat;
  assign new_n780_ = nn2139gat & ~nn1899gat;
  assign new_n781_ = ~new_n779_ & ~new_n780_;
  assign new_n782_1_ = nn2139gat & new_n781_;
  assign new_n783_ = ~pn3085gat & pn3086gat;
  assign new_n784_ = new_n773_ & new_n783_;
  assign new_n785_ = new_n776_ & new_n784_;
  assign new_n786_ = ~new_n767_1_ & ~new_n768_;
  assign new_n787_1_ = new_n769_ & new_n786_;
  assign new_n788_ = ~new_n785_ & ~new_n787_1_;
  assign pn3151gat = ~new_n782_1_ | ~new_n788_;
  assign new_n790_ = nn2190gat & ~nn2262gat;
  assign new_n791_ = ~nn2190gat & nn2262gat;
  assign new_n792_1_ = nn2190gat & ~new_n790_;
  assign new_n793_ = ~new_n791_ & new_n792_1_;
  assign pn3114gat = ~nn1282gat | ~new_n793_;
  assign new_n795_ = ~nn2139gat & ~nn1899gat;
  assign new_n796_ = nn2061gat & new_n795_;
  assign new_n797_1_ = ~nn2061gat & ~new_n795_;
  assign new_n798_ = ~new_n796_ & ~new_n797_1_;
  assign new_n799_ = ~nn2454gat & ~nn337gat;
  assign pn3150gat = ~new_n798_ | new_n799_;
  assign new_n801_ = ~nn1197gat & ~pn3116gat;
  assign new_n802_1_ = nn1197gat & pn3116gat;
  assign n862 = new_n801_ | new_n802_1_;
  assign new_n804_ = ~nn673gat & new_n757_1_;
  assign new_n805_ = ~nn366gat & new_n642_1_;
  assign new_n806_ = ~nn883gat & new_n636_;
  assign new_n807_1_ = ~nn919gat & new_n645_;
  assign new_n808_ = ~nn673gat & new_n639_;
  assign new_n809_ = ~new_n805_ & ~new_n806_;
  assign new_n810_ = ~new_n807_1_ & ~new_n808_;
  assign new_n811_ = new_n809_ & new_n810_;
  assign new_n812_1_ = ~new_n804_ & new_n811_;
  assign new_n813_ = new_n627_1_ & ~new_n812_1_;
  assign pn3124gat = ~n862 | new_n813_;
  assign new_n815_ = nn2339gat & ~nn2270gat;
  assign new_n816_ = ~nn2339gat & nn2270gat;
  assign new_n817_1_ = ~new_n815_ & ~new_n816_;
  assign new_n818_ = ~nn2390gat & ~nn2495gat;
  assign new_n819_ = nn2390gat & nn2495gat;
  assign new_n820_ = ~new_n818_ & ~new_n819_;
  assign new_n821_ = new_n817_1_ & new_n820_;
  assign new_n822_1_ = new_n817_1_ & ~new_n821_;
  assign new_n823_ = new_n820_ & ~new_n821_;
  assign n547 = new_n822_1_ | new_n823_;
  assign new_n825_ = new_n627_1_ & ~new_n760_;
  assign pn3125gat = ~n547 | new_n825_;
  assign new_n827_1_ = ~nn673gat & nn1241gat;
  assign new_n828_ = nn1294gat & new_n827_1_;
  assign new_n829_ = nn673gat & nn1241gat;
  assign new_n830_ = ~nn1294gat & new_n829_;
  assign new_n831_ = nn673gat & ~nn1241gat;
  assign new_n832_1_ = nn1294gat & new_n831_;
  assign new_n833_ = ~nn673gat & ~nn1241gat;
  assign new_n834_ = ~nn1294gat & new_n833_;
  assign new_n835_ = ~new_n828_ & ~new_n830_;
  assign new_n836_ = ~new_n832_1_ & ~new_n834_;
  assign new_n837_1_ = new_n835_ & new_n836_;
  assign new_n838_ = nn1080gat & ~nn1148gat;
  assign new_n839_ = nn865gat & new_n838_;
  assign new_n840_ = nn1080gat & nn1148gat;
  assign new_n841_ = ~nn865gat & new_n840_;
  assign new_n842_1_ = ~nn1080gat & nn1148gat;
  assign new_n843_ = nn865gat & new_n842_1_;
  assign new_n844_ = ~nn1080gat & ~nn1148gat;
  assign new_n845_ = ~nn865gat & new_n844_;
  assign new_n846_ = ~new_n839_ & ~new_n841_;
  assign new_n847_1_ = ~new_n843_ & ~new_n845_;
  assign new_n848_ = new_n846_ & new_n847_1_;
  assign new_n849_ = nn957gat & ~nn861gat;
  assign new_n850_ = nn1068gat & new_n849_;
  assign new_n851_ = nn957gat & nn861gat;
  assign new_n852_1_ = ~nn1068gat & new_n851_;
  assign new_n853_ = ~nn957gat & nn861gat;
  assign new_n854_ = nn1068gat & new_n853_;
  assign new_n855_ = ~nn957gat & ~nn861gat;
  assign new_n856_ = ~nn1068gat & new_n855_;
  assign new_n857_1_ = ~new_n850_ & ~new_n852_1_;
  assign new_n858_ = ~new_n854_ & ~new_n856_;
  assign new_n859_ = new_n857_1_ & new_n858_;
  assign new_n860_ = ~new_n837_1_ & ~new_n848_;
  assign new_n861_ = new_n859_ & new_n860_;
  assign new_n862_1_ = ~new_n837_1_ & new_n848_;
  assign new_n863_ = ~new_n859_ & new_n862_1_;
  assign new_n864_ = new_n837_1_ & new_n848_;
  assign new_n865_ = new_n859_ & new_n864_;
  assign new_n866_ = new_n837_1_ & ~new_n848_;
  assign new_n867_1_ = ~new_n859_ & new_n866_;
  assign new_n868_ = ~new_n861_ & ~new_n863_;
  assign new_n869_ = ~new_n865_ & ~new_n867_1_;
  assign n732 = ~new_n868_ | ~new_n869_;
  assign new_n871_ = ~nn160gat & new_n645_;
  assign new_n872_1_ = ~nn553gat & new_n642_1_;
  assign new_n873_ = ~nn816gat & new_n636_;
  assign new_n874_ = ~nn957gat & new_n639_;
  assign new_n875_ = ~new_n871_ & ~new_n872_1_;
  assign new_n876_ = ~new_n873_ & ~new_n874_;
  assign new_n877_1_ = new_n875_ & new_n876_;
  assign new_n878_ = new_n627_1_ & ~new_n877_1_;
  assign pn3119gat = ~n732 | new_n878_;
  assign new_n880_ = nn842gat & ~nn919gat;
  assign new_n881_ = nn846gat & new_n880_;
  assign new_n882_1_ = nn842gat & nn919gat;
  assign new_n883_ = ~nn846gat & new_n882_1_;
  assign new_n884_ = ~nn842gat & nn919gat;
  assign new_n885_ = nn846gat & new_n884_;
  assign new_n886_ = ~nn842gat & ~nn919gat;
  assign new_n887_1_ = ~nn846gat & new_n886_;
  assign new_n888_ = ~new_n881_ & ~new_n883_;
  assign new_n889_ = ~new_n885_ & ~new_n887_1_;
  assign new_n890_ = new_n888_ & new_n889_;
  assign new_n891_ = ~nn398gat & nn402gat;
  assign new_n892_1_ = nn341gat & new_n891_;
  assign new_n893_ = nn398gat & nn402gat;
  assign new_n894_ = ~nn341gat & new_n893_;
  assign new_n895_ = nn398gat & ~nn402gat;
  assign new_n896_ = nn341gat & new_n895_;
  assign new_n897_1_ = ~nn398gat & ~nn402gat;
  assign new_n898_ = ~nn341gat & new_n897_1_;
  assign new_n899_ = ~new_n892_1_ & ~new_n894_;
  assign new_n900_ = ~new_n896_ & ~new_n898_;
  assign new_n901_ = new_n899_ & new_n900_;
  assign new_n902_1_ = nn160gat & ~nn337gat;
  assign new_n903_ = nn271gat & new_n902_1_;
  assign new_n904_ = nn160gat & nn337gat;
  assign new_n905_ = ~nn271gat & new_n904_;
  assign new_n906_ = ~nn160gat & nn337gat;
  assign new_n907_1_ = nn271gat & new_n906_;
  assign new_n908_ = ~nn160gat & ~nn337gat;
  assign new_n909_ = ~nn271gat & new_n908_;
  assign new_n910_ = ~new_n903_ & ~new_n905_;
  assign new_n911_ = ~new_n907_1_ & ~new_n909_;
  assign new_n912_1_ = new_n910_ & new_n911_;
  assign new_n913_ = ~new_n890_ & ~new_n901_;
  assign new_n914_ = new_n912_1_ & new_n913_;
  assign new_n915_ = ~new_n890_ & new_n901_;
  assign new_n916_ = ~new_n912_1_ & new_n915_;
  assign new_n917_1_ = new_n890_ & new_n901_;
  assign new_n918_ = new_n912_1_ & new_n917_1_;
  assign new_n919_ = new_n890_ & ~new_n901_;
  assign new_n920_ = ~new_n912_1_ & new_n919_;
  assign new_n921_ = ~new_n914_ & ~new_n916_;
  assign new_n922_1_ = ~new_n918_ & ~new_n920_;
  assign n787 = ~new_n921_ | ~new_n922_1_;
  assign new_n924_ = ~nn580gat & new_n636_;
  assign new_n925_ = ~nn861gat & new_n639_;
  assign new_n926_ = ~nn777gat & new_n642_1_;
  assign new_n927_1_ = ~nn337gat & new_n645_;
  assign new_n928_ = ~new_n924_ & ~new_n925_;
  assign new_n929_ = ~new_n926_ & ~new_n927_1_;
  assign new_n930_ = new_n928_ & new_n929_;
  assign new_n931_ = new_n627_1_ & ~new_n930_;
  assign pn3118gat = ~n787 | new_n931_;
  assign new_n933_ = ~nn322gat & new_n642_1_;
  assign new_n934_ = ~nn865gat & new_n639_;
  assign new_n935_ = ~nn341gat & new_n645_;
  assign new_n936_ = ~nn584gat & new_n636_;
  assign new_n937_1_ = ~new_n933_ & ~new_n934_;
  assign new_n938_ = ~new_n935_ & ~new_n936_;
  assign new_n939_ = new_n937_1_ & new_n938_;
  assign new_n940_ = new_n627_1_ & ~new_n939_;
  assign pn3120gat = ~n787 | new_n940_;
  assign new_n942_1_ = nn820gat & ~nn883gat;
  assign new_n943_ = nn824gat & new_n942_1_;
  assign new_n944_ = nn820gat & nn883gat;
  assign new_n945_ = ~nn824gat & new_n944_;
  assign new_n946_ = ~nn820gat & nn883gat;
  assign new_n947_1_ = nn824gat & new_n946_;
  assign new_n948_ = ~nn820gat & ~nn883gat;
  assign new_n949_ = ~nn824gat & new_n948_;
  assign new_n950_ = ~new_n943_ & ~new_n945_;
  assign new_n951_ = ~new_n947_1_ & ~new_n949_;
  assign new_n952_1_ = new_n950_ & new_n951_;
  assign new_n953_ = ~nn699gat & nn684gat;
  assign new_n954_ = nn584gat & new_n953_;
  assign new_n955_ = nn699gat & nn684gat;
  assign new_n956_ = ~nn584gat & new_n955_;
  assign new_n957_1_ = nn699gat & ~nn684gat;
  assign new_n958_ = nn584gat & new_n957_1_;
  assign new_n959_ = ~nn699gat & ~nn684gat;
  assign new_n960_ = ~nn584gat & new_n959_;
  assign new_n961_ = ~new_n954_ & ~new_n956_;
  assign new_n962_1_ = ~new_n958_ & ~new_n960_;
  assign new_n963_ = new_n961_ & new_n962_1_;
  assign new_n964_ = nn816gat & ~nn580gat;
  assign new_n965_ = nn680gat & new_n964_;
  assign new_n966_ = nn816gat & nn580gat;
  assign new_n967_1_ = ~nn680gat & new_n966_;
  assign new_n968_ = ~nn816gat & nn580gat;
  assign new_n969_ = nn680gat & new_n968_;
  assign new_n970_ = ~nn816gat & ~nn580gat;
  assign new_n971_ = ~nn680gat & new_n970_;
  assign new_n972_1_ = ~new_n965_ & ~new_n967_1_;
  assign new_n973_ = ~new_n969_ & ~new_n971_;
  assign new_n974_ = new_n972_1_ & new_n973_;
  assign new_n975_ = ~new_n952_1_ & ~new_n963_;
  assign new_n976_ = new_n974_ & new_n975_;
  assign new_n977_1_ = ~new_n952_1_ & new_n963_;
  assign new_n978_ = ~new_n974_ & new_n977_1_;
  assign new_n979_ = new_n952_1_ & new_n963_;
  assign new_n980_ = new_n974_ & new_n979_;
  assign new_n981_ = new_n952_1_ & ~new_n963_;
  assign new_n982_1_ = ~new_n974_ & new_n981_;
  assign new_n983_ = ~new_n976_ & ~new_n978_;
  assign new_n984_ = ~new_n980_ & ~new_n982_1_;
  assign n702 = ~new_n983_ | ~new_n984_;
  assign new_n986_ = ~nn699gat & new_n636_;
  assign new_n987_ = ~nn1148gat & new_n639_;
  assign new_n988_ = ~nn398gat & new_n645_;
  assign new_n989_ = ~nn314gat & new_n642_1_;
  assign new_n990_ = ~new_n986_ & ~new_n987_;
  assign new_n991_ = ~new_n988_ & ~new_n989_;
  assign new_n992_ = new_n990_ & new_n991_;
  assign new_n993_ = new_n627_1_ & ~new_n992_;
  assign pn3121gat = ~n702 | new_n993_;
  assign new_n995_ = ~nn919gat & nn830gat;
  assign new_n996_ = nn846gat & new_n995_;
  assign new_n997_ = nn919gat & nn830gat;
  assign new_n998_ = ~nn846gat & new_n997_;
  assign new_n999_ = nn919gat & ~nn830gat;
  assign new_n1000_ = nn846gat & new_n999_;
  assign new_n1001_ = ~nn919gat & ~nn830gat;
  assign new_n1002_ = ~nn846gat & new_n1001_;
  assign new_n1003_ = ~new_n996_ & ~new_n998_;
  assign new_n1004_ = ~new_n1000_ & ~new_n1002_;
  assign new_n1005_ = new_n1003_ & new_n1004_;
  assign new_n1006_ = nn614gat & new_n891_;
  assign new_n1007_ = ~nn614gat & new_n893_;
  assign new_n1008_ = nn614gat & new_n895_;
  assign new_n1009_ = ~nn614gat & new_n897_1_;
  assign new_n1010_ = ~new_n1006_ & ~new_n1007_;
  assign new_n1011_ = ~new_n1008_ & ~new_n1009_;
  assign new_n1012_ = new_n1010_ & new_n1011_;
  assign new_n1013_ = nn707gat & ~nn838gat;
  assign new_n1014_ = nn834gat & new_n1013_;
  assign new_n1015_ = nn707gat & nn838gat;
  assign new_n1016_ = ~nn834gat & new_n1015_;
  assign new_n1017_ = ~nn707gat & nn838gat;
  assign new_n1018_ = nn834gat & new_n1017_;
  assign new_n1019_ = ~nn707gat & ~nn838gat;
  assign new_n1020_ = ~nn834gat & new_n1019_;
  assign new_n1021_ = ~new_n1014_ & ~new_n1016_;
  assign new_n1022_ = ~new_n1018_ & ~new_n1020_;
  assign new_n1023_ = new_n1021_ & new_n1022_;
  assign new_n1024_ = ~new_n1005_ & ~new_n1012_;
  assign new_n1025_ = new_n1023_ & new_n1024_;
  assign new_n1026_ = ~new_n1005_ & new_n1012_;
  assign new_n1027_ = ~new_n1023_ & new_n1026_;
  assign new_n1028_ = new_n1005_ & new_n1012_;
  assign new_n1029_ = new_n1023_ & new_n1028_;
  assign new_n1030_ = new_n1005_ & ~new_n1012_;
  assign new_n1031_ = ~new_n1023_ & new_n1030_;
  assign new_n1032_ = ~new_n1025_ & ~new_n1027_;
  assign new_n1033_ = ~new_n1029_ & ~new_n1031_;
  assign n717 = ~new_n1032_ | ~new_n1033_;
  assign new_n1035_ = ~nn684gat & new_n636_;
  assign new_n1036_ = ~nn402gat & new_n645_;
  assign new_n1037_ = ~nn1080gat & new_n639_;
  assign new_n1038_ = ~nn318gat & new_n642_1_;
  assign new_n1039_ = ~new_n1035_ & ~new_n1036_;
  assign new_n1040_ = ~new_n1037_ & ~new_n1038_;
  assign new_n1041_ = new_n1039_ & new_n1040_;
  assign new_n1042_ = new_n627_1_ & ~new_n1041_;
  assign pn3122gat = ~n717 | new_n1042_;
  assign new_n1044_ = nn667gat & ~new_n746_;
  assign new_n1045_ = ~nn667gat & new_n746_;
  assign n972 = new_n1044_ | new_n1045_;
  assign new_n1047_ = ~nn561gat & new_n642_1_;
  assign new_n1048_ = ~nn846gat & new_n645_;
  assign new_n1049_ = ~nn824gat & new_n636_;
  assign new_n1050_ = ~nn1294gat & new_n639_;
  assign new_n1051_ = ~new_n1047_ & ~new_n1048_;
  assign new_n1052_ = ~new_n1049_ & ~new_n1050_;
  assign new_n1053_ = new_n1051_ & new_n1052_;
  assign new_n1054_ = new_n627_1_ & ~new_n1053_;
  assign pn3123gat = ~n972 | new_n1054_;
  assign new_n1056_ = ~new_n710_ & ~new_n1041_;
  assign new_n1057_ = ~nn402gat & new_n636_;
  assign new_n1058_ = ~nn402gat & new_n639_;
  assign new_n1059_ = ~new_n1057_ & ~new_n1058_;
  assign new_n1060_ = ~nn1135gat & new_n642_1_;
  assign new_n1061_ = new_n1059_ & ~new_n1060_;
  assign new_n1062_ = ~new_n704_ & ~new_n1061_;
  assign pn3135gat = new_n1056_ | new_n1062_;
  assign new_n1064_ = ~new_n710_ & ~new_n992_;
  assign new_n1065_ = ~nn1045gat & new_n642_1_;
  assign new_n1066_ = ~nn398gat & new_n639_;
  assign new_n1067_ = ~nn398gat & new_n636_;
  assign new_n1068_ = ~new_n1066_ & ~new_n1067_;
  assign new_n1069_ = ~new_n1065_ & new_n1068_;
  assign new_n1070_ = ~new_n704_ & ~new_n1069_;
  assign pn3134gat = new_n1064_ | new_n1070_;
  assign new_n1072_ = ~nn2403gat & new_n586_;
  assign new_n1073_ = ~nn2347gat & new_n1072_;
  assign new_n1074_ = ~nn2407gat & ~new_n1073_;
  assign new_n1075_ = nn2407gat & new_n1073_;
  assign new_n1076_ = ~new_n1074_ & ~new_n1075_;
  assign pn3108gat = ~nn1035gat | ~new_n1076_;
  assign new_n1078_ = ~nn919gat & new_n636_;
  assign new_n1079_ = ~nn919gat & new_n639_;
  assign new_n1080_ = ~new_n1078_ & ~new_n1079_;
  assign new_n1081_ = ~nn1226gat & new_n642_1_;
  assign new_n1082_ = new_n1080_ & ~new_n1081_;
  assign new_n1083_ = ~new_n704_ & ~new_n1082_;
  assign new_n1084_ = ~new_n710_ & ~new_n812_1_;
  assign pn3137gat = new_n1083_ | new_n1084_;
  assign new_n1086_ = nn2403gat & ~nn2347gat;
  assign new_n1087_ = ~nn2347gat & ~new_n586_;
  assign new_n1088_ = nn2347gat & new_n586_;
  assign new_n1089_ = ~nn2403gat & new_n1088_;
  assign new_n1090_ = ~new_n1086_ & ~new_n1087_;
  assign new_n1091_ = ~new_n1089_ & new_n1090_;
  assign pn3109gat = ~nn1072gat | ~new_n1091_;
  assign new_n1093_ = ~nn1282gat & new_n642_1_;
  assign new_n1094_ = ~nn846gat & new_n639_;
  assign new_n1095_ = ~nn846gat & new_n636_;
  assign new_n1096_ = ~new_n1094_ & ~new_n1095_;
  assign new_n1097_ = ~new_n1093_ & new_n1096_;
  assign new_n1098_ = ~new_n704_ & ~new_n1097_;
  assign new_n1099_ = ~new_n710_ & ~new_n1053_;
  assign pn3136gat = new_n1098_ | new_n1099_;
  assign new_n1101_ = ~new_n710_ & ~new_n930_;
  assign new_n1102_ = ~nn1072gat & new_n642_1_;
  assign new_n1103_ = ~nn337gat & new_n639_;
  assign new_n1104_ = ~nn838gat & new_n636_;
  assign new_n1105_ = ~new_n1103_ & ~new_n1104_;
  assign new_n1106_ = ~new_n1102_ & new_n1105_;
  assign new_n1107_ = ~new_n704_ & ~new_n1106_;
  assign pn3131gat = new_n1101_ | new_n1107_;
  assign new_n1109_ = ~nn834gat & new_n636_;
  assign new_n1110_ = ~nn271gat & new_n639_;
  assign new_n1111_ = ~new_n1109_ & ~new_n1110_;
  assign new_n1112_ = ~nn1035gat & new_n642_1_;
  assign new_n1113_ = new_n1111_ & ~new_n1112_;
  assign new_n1114_ = ~new_n704_ & ~new_n1113_;
  assign new_n1115_ = ~new_n649_ & ~new_n710_;
  assign pn3130gat = new_n1114_ | new_n1115_;
  assign new_n1117_ = ~nn931gat & new_n642_1_;
  assign new_n1118_ = ~nn341gat & new_n639_;
  assign new_n1119_ = ~nn614gat & new_n636_;
  assign new_n1120_ = ~new_n1118_ & ~new_n1119_;
  assign new_n1121_ = ~new_n1117_ & new_n1120_;
  assign new_n1122_ = ~new_n704_ & ~new_n1121_;
  assign new_n1123_ = ~new_n710_ & ~new_n939_;
  assign pn3133gat = new_n1122_ | new_n1123_;
  assign new_n1125_ = ~new_n710_ & ~new_n877_1_;
  assign new_n1126_ = ~nn1121gat & new_n642_1_;
  assign new_n1127_ = ~nn160gat & new_n639_;
  assign new_n1128_ = ~nn707gat & new_n636_;
  assign new_n1129_ = ~new_n1127_ & ~new_n1128_;
  assign new_n1130_ = ~new_n1126_ & new_n1129_;
  assign new_n1131_ = ~new_n704_ & ~new_n1130_;
  assign pn3132gat = new_n1125_ | new_n1131_;
  assign new_n1133_ = nn1880gat & nn1767gat;
  assign pn3149gat = ~nn1834gat | ~new_n1133_;
  assign new_n1135_ = nn2176gat & nn2033gat;
  assign new_n1136_ = nn2169gat & new_n1135_;
  assign new_n1137_ = nn2095gat & new_n1136_;
  assign new_n1138_ = nn2110gat & nn2037gat;
  assign new_n1139_ = new_n1137_ & new_n1138_;
  assign new_n1140_ = nn1775gat & nn1771gat;
  assign new_n1141_ = nn2514gat & new_n1140_;
  assign new_n1142_ = nn1871gat & new_n1141_;
  assign pn3146gat = new_n1139_ & ~new_n1142_;
  assign pn3147gat = ~nn2446gat | ~nn2450gat;
  assign new_n1145_ = nn2399gat & ~nn2203gat;
  assign new_n1146_ = nn2207gat & new_n1145_;
  assign new_n1147_ = nn2399gat & nn2203gat;
  assign new_n1148_ = ~nn2207gat & new_n1147_;
  assign new_n1149_ = ~nn2399gat & nn2203gat;
  assign new_n1150_ = nn2207gat & new_n1149_;
  assign new_n1151_ = ~nn2399gat & ~nn2203gat;
  assign new_n1152_ = ~nn2207gat & new_n1151_;
  assign new_n1153_ = ~new_n1146_ & ~new_n1148_;
  assign new_n1154_ = ~new_n1150_ & ~new_n1152_;
  assign new_n1155_ = new_n1153_ & new_n1154_;
  assign new_n1156_ = ~nn2562gat & ~nn2640gat;
  assign new_n1157_ = nn2343gat & new_n1156_;
  assign new_n1158_ = nn2562gat & ~nn2640gat;
  assign new_n1159_ = ~nn2343gat & new_n1158_;
  assign new_n1160_ = nn2562gat & nn2640gat;
  assign new_n1161_ = nn2343gat & new_n1160_;
  assign new_n1162_ = ~nn2562gat & nn2640gat;
  assign new_n1163_ = ~nn2343gat & new_n1162_;
  assign new_n1164_ = ~new_n1157_ & ~new_n1159_;
  assign new_n1165_ = ~new_n1161_ & ~new_n1163_;
  assign new_n1166_ = new_n1164_ & new_n1165_;
  assign new_n1167_ = new_n1155_ & new_n1166_;
  assign new_n1168_ = new_n1155_ & ~new_n1167_;
  assign new_n1169_ = new_n1166_ & ~new_n1167_;
  assign n807 = new_n1168_ | new_n1169_;
  assign new_n1171_ = ~nn699gat & ~pn3149gat;
  assign new_n1172_ = ~nn1148gat & pn3149gat;
  assign new_n1173_ = ~new_n1171_ & ~new_n1172_;
  assign new_n1174_ = nn2207gat & nn2203gat;
  assign new_n1175_ = ~nn2343gat & nn2562gat;
  assign new_n1176_ = ~nn2399gat & new_n1175_;
  assign new_n1177_ = new_n1174_ & new_n1176_;
  assign new_n1178_ = ~new_n1173_ & new_n1177_;
  assign new_n1179_ = ~nn824gat & ~pn3149gat;
  assign new_n1180_ = ~nn1294gat & pn3149gat;
  assign new_n1181_ = ~new_n1179_ & ~new_n1180_;
  assign new_n1182_ = nn2343gat & nn2562gat;
  assign new_n1183_ = nn2399gat & new_n1182_;
  assign new_n1184_ = nn2207gat & ~nn2203gat;
  assign new_n1185_ = new_n1183_ & new_n1184_;
  assign new_n1186_ = ~new_n1181_ & new_n1185_;
  assign new_n1187_ = ~nn684gat & ~pn3149gat;
  assign new_n1188_ = ~nn1080gat & pn3149gat;
  assign new_n1189_ = ~new_n1187_ & ~new_n1188_;
  assign new_n1190_ = ~nn2343gat & ~nn2562gat;
  assign new_n1191_ = ~nn2399gat & new_n1190_;
  assign new_n1192_ = new_n1174_ & new_n1191_;
  assign new_n1193_ = ~new_n1189_ & new_n1192_;
  assign new_n1194_ = nn2343gat & ~nn2562gat;
  assign new_n1195_ = nn2399gat & new_n1194_;
  assign new_n1196_ = new_n1184_ & new_n1195_;
  assign new_n1197_ = ~nn673gat & pn3149gat;
  assign new_n1198_ = ~nn883gat & ~pn3149gat;
  assign new_n1199_ = ~new_n1197_ & ~new_n1198_;
  assign new_n1200_ = new_n1196_ & ~new_n1199_;
  assign new_n1201_ = ~new_n1178_ & ~new_n1186_;
  assign new_n1202_ = ~new_n1193_ & ~new_n1200_;
  assign new_n1203_ = new_n1201_ & new_n1202_;
  assign new_n1204_ = new_n1174_ & new_n1183_;
  assign new_n1205_ = nn919gat & nn846gat;
  assign new_n1206_ = new_n891_ & new_n1205_;
  assign new_n1207_ = ~nn2454gat & new_n1206_;
  assign new_n1208_ = nn2084gat & ~new_n1207_;
  assign new_n1209_ = new_n1204_ & ~new_n1208_;
  assign new_n1210_ = nn919gat & ~nn846gat;
  assign new_n1211_ = new_n893_ & new_n1210_;
  assign new_n1212_ = ~nn2454gat & new_n1211_;
  assign new_n1213_ = ~nn919gat & ~nn846gat;
  assign new_n1214_ = new_n893_ & new_n1213_;
  assign new_n1215_ = ~nn2454gat & new_n1214_;
  assign new_n1216_ = ~new_n1212_ & ~new_n1215_;
  assign new_n1217_ = ~new_n1207_ & new_n1216_;
  assign new_n1218_ = new_n1174_ & new_n1195_;
  assign new_n1219_ = ~new_n1217_ & new_n1218_;
  assign new_n1220_ = ~new_n1209_ & ~new_n1219_;
  assign new_n1221_ = nn2399gat & new_n1190_;
  assign new_n1222_ = new_n1174_ & new_n1221_;
  assign new_n1223_ = ~nn861gat & pn3149gat;
  assign new_n1224_ = ~nn580gat & ~pn3149gat;
  assign new_n1225_ = ~new_n1223_ & ~new_n1224_;
  assign new_n1226_ = new_n1222_ & ~new_n1225_;
  assign new_n1227_ = nn2399gat & new_n1175_;
  assign new_n1228_ = new_n1174_ & new_n1227_;
  assign new_n1229_ = ~nn680gat & ~pn3149gat;
  assign new_n1230_ = ~nn1068gat & pn3149gat;
  assign new_n1231_ = ~new_n1229_ & ~new_n1230_;
  assign new_n1232_ = new_n1228_ & ~new_n1231_;
  assign new_n1233_ = nn2343gat & ~nn2399gat;
  assign new_n1234_ = ~nn2562gat & new_n1233_;
  assign new_n1235_ = new_n1174_ & new_n1234_;
  assign new_n1236_ = ~nn584gat & ~pn3149gat;
  assign new_n1237_ = ~nn865gat & pn3149gat;
  assign new_n1238_ = ~new_n1236_ & ~new_n1237_;
  assign new_n1239_ = new_n1235_ & ~new_n1238_;
  assign new_n1240_ = nn2562gat & new_n1233_;
  assign new_n1241_ = new_n1174_ & new_n1240_;
  assign new_n1242_ = ~nn957gat & pn3149gat;
  assign new_n1243_ = ~nn816gat & ~pn3149gat;
  assign new_n1244_ = ~new_n1242_ & ~new_n1243_;
  assign new_n1245_ = new_n1241_ & ~new_n1244_;
  assign new_n1246_ = ~new_n1226_ & ~new_n1232_;
  assign new_n1247_ = ~new_n1239_ & ~new_n1245_;
  assign new_n1248_ = new_n1246_ & new_n1247_;
  assign new_n1249_ = ~nn271gat & pn3149gat;
  assign new_n1250_ = ~nn834gat & ~pn3149gat;
  assign new_n1251_ = ~new_n1249_ & ~new_n1250_;
  assign new_n1252_ = new_n1184_ & new_n1227_;
  assign new_n1253_ = ~new_n1251_ & new_n1252_;
  assign new_n1254_ = new_n1184_ & new_n1221_;
  assign new_n1255_ = ~nn337gat & pn3149gat;
  assign new_n1256_ = ~nn838gat & ~pn3149gat;
  assign new_n1257_ = ~new_n1255_ & ~new_n1256_;
  assign new_n1258_ = new_n1254_ & ~new_n1257_;
  assign new_n1259_ = ~nn341gat & pn3149gat;
  assign new_n1260_ = ~nn614gat & ~pn3149gat;
  assign new_n1261_ = ~new_n1259_ & ~new_n1260_;
  assign new_n1262_ = new_n1184_ & new_n1234_;
  assign new_n1263_ = ~new_n1261_ & new_n1262_;
  assign new_n1264_ = ~nn160gat & pn3149gat;
  assign new_n1265_ = ~nn707gat & ~pn3149gat;
  assign new_n1266_ = ~new_n1264_ & ~new_n1265_;
  assign new_n1267_ = new_n1184_ & new_n1240_;
  assign new_n1268_ = ~new_n1266_ & new_n1267_;
  assign new_n1269_ = ~new_n1253_ & ~new_n1258_;
  assign new_n1270_ = ~new_n1263_ & ~new_n1268_;
  assign new_n1271_ = new_n1269_ & new_n1270_;
  assign new_n1272_ = new_n1203_ & new_n1220_;
  assign new_n1273_ = new_n1248_ & new_n1272_;
  assign new_n1274_ = new_n1271_ & new_n1273_;
  assign new_n1275_ = nn1389gat & ~new_n1274_;
  assign new_n1276_ = ~nn1880gat & ~nn1763gat;
  assign n892 = ~nn2102gat | new_n1276_;
  assign new_n1278_ = pn3149gat & n892;
  assign new_n1279_ = ~nn1394gat & new_n1278_;
  assign new_n1280_ = ~nn1508gat & new_n1279_;
  assign new_n1281_ = pn3149gat & ~n892;
  assign new_n1282_ = ~nn1678gat & new_n1281_;
  assign new_n1283_ = ~nn1394gat & new_n1282_;
  assign new_n1284_ = ~nn2592gat & ~nn673gat;
  assign new_n1285_ = nn1871gat & new_n1284_;
  assign new_n1286_ = ~new_n1280_ & ~new_n1283_;
  assign new_n1287_ = ~new_n1285_ & new_n1286_;
  assign new_n1288_ = ~nn2207gat & nn2203gat;
  assign new_n1289_ = new_n1176_ & new_n1288_;
  assign new_n1290_ = ~nn561gat & new_n1289_;
  assign new_n1291_ = new_n1240_ & new_n1288_;
  assign new_n1292_ = ~nn314gat & new_n1291_;
  assign new_n1293_ = new_n1234_ & new_n1288_;
  assign new_n1294_ = ~nn318gat & new_n1293_;
  assign new_n1295_ = new_n1191_ & new_n1288_;
  assign new_n1296_ = ~nn366gat & new_n1295_;
  assign new_n1297_ = ~new_n1290_ & ~new_n1292_;
  assign new_n1298_ = ~new_n1294_ & ~new_n1296_;
  assign new_n1299_ = new_n1297_ & new_n1298_;
  assign new_n1300_ = new_n1227_ & new_n1288_;
  assign new_n1301_ = ~nn553gat & new_n1300_;
  assign new_n1302_ = new_n1221_ & new_n1288_;
  assign new_n1303_ = ~nn322gat & new_n1302_;
  assign new_n1304_ = new_n1195_ & new_n1288_;
  assign new_n1305_ = ~nn777gat & new_n1304_;
  assign new_n1306_ = new_n1183_ & new_n1288_;
  assign new_n1307_ = ~nn659gat & new_n1306_;
  assign new_n1308_ = ~new_n1301_ & ~new_n1303_;
  assign new_n1309_ = ~new_n1305_ & ~new_n1307_;
  assign new_n1310_ = new_n1308_ & new_n1309_;
  assign new_n1311_ = ~new_n746_ & ~new_n1215_;
  assign new_n1312_ = new_n746_ & new_n1215_;
  assign new_n1313_ = ~new_n1311_ & ~new_n1312_;
  assign new_n1314_ = ~nn2207gat & ~nn2203gat;
  assign new_n1315_ = new_n1183_ & new_n1314_;
  assign new_n1316_ = ~new_n1313_ & new_n1315_;
  assign new_n1317_ = new_n1299_ & new_n1310_;
  assign new_n1318_ = ~new_n1316_ & new_n1317_;
  assign new_n1319_ = ~new_n1216_ & ~new_n1318_;
  assign new_n1320_ = ~new_n1275_ & new_n1287_;
  assign new_n1321_ = ~new_n1319_ & new_n1320_;
  assign pn3144gat = ~n807 | ~new_n1321_;
  assign new_n1323_ = ~nn919gat & nn846gat;
  assign new_n1324_ = new_n893_ & new_n1323_;
  assign new_n1325_ = ~nn2454gat & new_n1324_;
  assign new_n1326_ = ~new_n1215_ & ~new_n1325_;
  assign new_n1327_ = ~new_n1212_ & new_n1326_;
  assign new_n1328_ = new_n895_ & new_n1323_;
  assign new_n1329_ = ~nn2454gat & new_n1328_;
  assign new_n1330_ = new_n895_ & new_n1205_;
  assign new_n1331_ = ~nn2454gat & new_n1330_;
  assign new_n1332_ = new_n1327_ & ~new_n1329_;
  assign new_n1333_ = ~new_n1207_ & ~new_n1331_;
  assign n212 = ~new_n1332_ | ~new_n1333_;
  assign new_n1335_ = nn1775gat & nn2514gat;
  assign new_n1336_ = nn1771gat & new_n1335_;
  assign pn3145gat = ~n212 & ~new_n1336_;
  assign new_n1338_ = ~nn1588gat & ~n892;
  assign new_n1339_ = nn1596gat & new_n1338_;
  assign new_n1340_ = ~nn1462gat & new_n1278_;
  assign new_n1341_ = nn1394gat & new_n1340_;
  assign new_n1342_ = ~new_n1329_ & new_n1333_;
  assign n337 = new_n1325_ | ~new_n1342_;
  assign new_n1344_ = new_n1216_ & ~n337;
  assign new_n1345_ = ~nn1340gat & ~new_n1344_;
  assign new_n1346_ = n892 & new_n1345_;
  assign new_n1347_ = nn2399gat & ~nn2207gat;
  assign new_n1348_ = ~nn2203gat & new_n1347_;
  assign new_n1349_ = nn2562gat & new_n1348_;
  assign new_n1350_ = ~nn2343gat & new_n1349_;
  assign new_n1351_ = new_n1346_ & ~new_n1350_;
  assign new_n1352_ = ~new_n1341_ & ~new_n1351_;
  assign new_n1353_ = ~nn1508gat & ~new_n1352_;
  assign new_n1354_ = ~nn1394gat & n337;
  assign new_n1355_ = ~n892 & new_n1354_;
  assign new_n1356_ = ~nn1525gat & new_n1355_;
  assign new_n1357_ = ~new_n1216_ & ~n892;
  assign new_n1358_ = ~nn1596gat & new_n1357_;
  assign new_n1359_ = nn1462gat & n892;
  assign new_n1360_ = ~new_n1358_ & ~new_n1359_;
  assign new_n1361_ = ~nn1678gat & ~new_n1360_;
  assign new_n1362_ = nn1821gat & ~nn1829gat;
  assign new_n1363_ = nn2021gat & nn1880gat;
  assign new_n1364_ = ~nn1775gat & new_n1363_;
  assign new_n1365_ = pn3097gat & new_n1364_;
  assign new_n1366_ = nn1821gat & ~new_n1365_;
  assign new_n1367_ = ~pn3098gat & ~new_n1362_;
  assign new_n1368_ = ~new_n1366_ & new_n1367_;
  assign new_n1369_ = nn1871gat & new_n1368_;
  assign new_n1370_ = ~nn1775gat & new_n1369_;
  assign new_n1371_ = ~new_n1353_ & ~new_n1356_;
  assign new_n1372_ = ~new_n1361_ & ~new_n1370_;
  assign new_n1373_ = new_n1371_ & new_n1372_;
  assign new_n1374_ = ~nn1596gat & ~nn1678gat;
  assign new_n1375_ = new_n1216_ & new_n1374_;
  assign new_n1376_ = ~n892 & new_n1375_;
  assign new_n1377_ = nn1394gat & new_n1376_;
  assign new_n1378_ = ~new_n1339_ & new_n1373_;
  assign pn3139gat = new_n1377_ | ~new_n1378_;
  assign new_n1380_ = ~new_n1278_ & ~new_n1346_;
  assign new_n1381_ = ~nn1456gat & ~new_n1380_;
  assign new_n1382_ = ~nn1675gat & new_n1355_;
  assign new_n1383_ = nn1340gat & n892;
  assign new_n1384_ = ~nn1807gat & new_n1383_;
  assign new_n1385_ = ~n892 & n337;
  assign new_n1386_ = nn1336gat & new_n1385_;
  assign new_n1387_ = ~new_n1357_ & ~new_n1386_;
  assign new_n1388_ = ~new_n1281_ & new_n1387_;
  assign new_n1389_ = ~nn1748gat & ~new_n1388_;
  assign new_n1390_ = ~new_n1381_ & ~new_n1382_;
  assign new_n1391_ = ~new_n1384_ & ~new_n1389_;
  assign pn3142gat = ~new_n1390_ | ~new_n1391_;
  assign pn3107gat = nn1871gat & ~new_n1140_;
  assign n232 = new_n1329_ | new_n1331_;
  assign new_n1395_ = nn2343gat & ~nn2203gat;
  assign new_n1396_ = nn2399gat & new_n1395_;
  assign new_n1397_ = ~nn2207gat & new_n1396_;
  assign new_n1398_ = ~nn2562gat & new_n1397_;
  assign new_n1399_ = ~nn2626gat & nn2490gat;
  assign new_n1400_ = nn2622gat & new_n1399_;
  assign new_n1401_ = nn2630gat & nn2543gat;
  assign new_n1402_ = new_n1400_ & new_n1401_;
  assign new_n1403_ = n232 & new_n1398_;
  assign pn3138gat = new_n1402_ & new_n1403_;
  assign new_n1405_ = ~nn2543gat & nn2634gat;
  assign new_n1406_ = nn2630gat & new_n1405_;
  assign new_n1407_ = nn2543gat & nn2634gat;
  assign new_n1408_ = ~nn2630gat & new_n1407_;
  assign new_n1409_ = nn2543gat & ~nn2634gat;
  assign new_n1410_ = nn2630gat & new_n1409_;
  assign new_n1411_ = ~nn2543gat & ~nn2634gat;
  assign new_n1412_ = ~nn2630gat & new_n1411_;
  assign new_n1413_ = ~new_n1406_ & ~new_n1408_;
  assign new_n1414_ = ~new_n1410_ & ~new_n1412_;
  assign new_n1415_ = new_n1413_ & new_n1414_;
  assign new_n1416_ = ~nn2626gat & ~nn2490gat;
  assign new_n1417_ = nn2622gat & new_n1416_;
  assign new_n1418_ = ~nn2622gat & new_n1399_;
  assign new_n1419_ = nn2626gat & nn2490gat;
  assign new_n1420_ = nn2622gat & new_n1419_;
  assign new_n1421_ = nn2626gat & ~nn2490gat;
  assign new_n1422_ = ~nn2622gat & new_n1421_;
  assign new_n1423_ = ~new_n1417_ & ~new_n1418_;
  assign new_n1424_ = ~new_n1420_ & ~new_n1422_;
  assign new_n1425_ = new_n1423_ & new_n1424_;
  assign new_n1426_ = new_n1415_ & new_n1425_;
  assign new_n1427_ = new_n1415_ & ~new_n1426_;
  assign new_n1428_ = new_n1425_ & ~new_n1426_;
  assign n942 = new_n1427_ | new_n1428_;
  assign pn3143gat = ~new_n1321_ | ~n942;
  assign new_n1431_ = pn3094gat & new_n787_1_;
  assign new_n1432_ = ~nn2061gat & new_n795_;
  assign new_n1433_ = ~nn2143gat & new_n1432_;
  assign new_n1434_ = ~nn1850gat & ~new_n1433_;
  assign new_n1435_ = nn1850gat & new_n1433_;
  assign new_n1436_ = ~new_n1434_ & ~new_n1435_;
  assign new_n1437_ = ~pn3092gat & ~pn3091gat;
  assign new_n1438_ = new_n785_ & ~new_n1437_;
  assign new_n1439_ = ~new_n1431_ & new_n1436_;
  assign pn3104gat = new_n1438_ | ~new_n1439_;
  assign new_n1441_ = ~new_n1339_ & ~new_n1377_;
  assign pn3140gat = ~new_n1373_ | ~new_n1441_;
  assign new_n1443_ = pn3094gat & new_n771_;
  assign new_n1444_ = ~nn2143gat & ~new_n795_;
  assign new_n1445_ = ~nn2143gat & nn2061gat;
  assign new_n1446_ = nn2143gat & ~nn2061gat;
  assign new_n1447_ = new_n795_ & new_n1446_;
  assign new_n1448_ = ~new_n1444_ & ~new_n1445_;
  assign new_n1449_ = ~new_n1447_ & new_n1448_;
  assign new_n1450_ = new_n778_ & ~new_n1437_;
  assign new_n1451_ = ~new_n1443_ & new_n1449_;
  assign pn3105gat = new_n1450_ | ~new_n1451_;
  assign new_n1453_ = nn1850gat & new_n795_;
  assign new_n1454_ = nn2061gat & new_n1453_;
  assign new_n1455_ = nn2143gat & new_n1454_;
  assign new_n1456_ = ~nn2403gat & new_n582_1_;
  assign new_n1457_ = nn2407gat & ~nn2347gat;
  assign new_n1458_ = new_n1456_ & new_n1457_;
  assign n172 = new_n1455_ & new_n1458_;
  assign new_n1460_ = ~pn3100gat & pn3147gat;
  assign new_n1461_ = ~new_n1362_ & ~new_n1460_;
  assign new_n1462_ = nn2472gat & new_n1461_;
  assign new_n1463_ = new_n895_ & new_n1210_;
  assign n872 = ~nn2454gat & new_n1463_;
  assign n177 = new_n1462_ & n872;
  assign new_n1466_ = nn2658gat & nn2506gat;
  assign new_n1467_ = nn2502gat & new_n1466_;
  assign new_n1468_ = nn2510gat & new_n1467_;
  assign new_n1469_ = nn2309gat & new_n1468_;
  assign new_n1470_ = nn2588gat & new_n1469_;
  assign new_n1471_ = ~pn3100gat & ~new_n1470_;
  assign new_n1472_ = nn2143gat & new_n795_;
  assign new_n1473_ = nn1850gat & new_n1472_;
  assign new_n1474_ = ~nn2061gat & new_n1473_;
  assign new_n1475_ = ~n892 & new_n1474_;
  assign new_n1476_ = pn3149gat & new_n1475_;
  assign new_n1477_ = nn2061gat & nn2139gat;
  assign new_n1478_ = nn2143gat & new_n1477_;
  assign new_n1479_ = ~nn1850gat & new_n1478_;
  assign new_n1480_ = ~nn1899gat & new_n1479_;
  assign new_n1481_ = new_n1278_ & new_n1480_;
  assign new_n1482_ = ~new_n1476_ & ~new_n1481_;
  assign new_n1483_ = ~nn2403gat & nn2347gat;
  assign new_n1484_ = new_n581_ & new_n1483_;
  assign new_n1485_ = ~nn2407gat & new_n1484_;
  assign new_n1486_ = nn398gat & ~nn846gat;
  assign new_n1487_ = nn398gat & ~nn919gat;
  assign new_n1488_ = new_n895_ & ~new_n1486_;
  assign new_n1489_ = new_n1487_ & new_n1488_;
  assign new_n1490_ = ~new_n1482_ & new_n1485_;
  assign new_n1491_ = new_n1489_ & new_n1490_;
  assign new_n1492_ = new_n895_ & ~new_n1487_;
  assign new_n1493_ = ~new_n1486_ & new_n1492_;
  assign new_n1494_ = nn2394gat & nn2440gat;
  assign new_n1495_ = ~nn2407gat & new_n1483_;
  assign new_n1496_ = new_n1494_ & new_n1495_;
  assign new_n1497_ = ~new_n1482_ & new_n1493_;
  assign new_n1498_ = new_n1496_ & new_n1497_;
  assign new_n1499_ = new_n1486_ & new_n1487_;
  assign new_n1500_ = ~new_n895_ & new_n1499_;
  assign new_n1501_ = nn2403gat & nn2347gat;
  assign new_n1502_ = ~nn2407gat & new_n1501_;
  assign new_n1503_ = new_n586_ & new_n1502_;
  assign new_n1504_ = ~new_n1482_ & new_n1500_;
  assign new_n1505_ = new_n1503_ & new_n1504_;
  assign new_n1506_ = ~new_n1491_ & ~new_n1498_;
  assign new_n1507_ = ~new_n1505_ & new_n1506_;
  assign new_n1508_ = new_n582_1_ & new_n1495_;
  assign new_n1509_ = new_n1486_ & new_n1492_;
  assign new_n1510_ = ~new_n1482_ & new_n1508_;
  assign new_n1511_ = new_n1509_ & new_n1510_;
  assign new_n1512_ = new_n586_ & new_n1483_;
  assign new_n1513_ = ~nn2407gat & new_n1512_;
  assign new_n1514_ = new_n895_ & new_n1499_;
  assign new_n1515_ = ~new_n1482_ & new_n1513_;
  assign new_n1516_ = new_n1514_ & new_n1515_;
  assign new_n1517_ = ~nn2407gat & new_n1494_;
  assign new_n1518_ = new_n1086_ & new_n1517_;
  assign new_n1519_ = ~new_n1482_ & new_n1518_;
  assign new_n1520_ = ~new_n1511_ & ~new_n1516_;
  assign new_n1521_ = ~new_n1519_ & new_n1520_;
  assign new_n1522_ = ~new_n895_ & new_n1486_;
  assign new_n1523_ = ~new_n1487_ & new_n1522_;
  assign new_n1524_ = ~nn2407gat & new_n582_1_;
  assign new_n1525_ = new_n1501_ & new_n1524_;
  assign new_n1526_ = ~new_n1482_ & new_n1523_;
  assign new_n1527_ = new_n1525_ & new_n1526_;
  assign new_n1528_ = nn398gat & ~new_n1487_;
  assign new_n1529_ = ~new_n895_ & new_n1528_;
  assign new_n1530_ = ~new_n1486_ & new_n1529_;
  assign new_n1531_ = new_n1501_ & new_n1517_;
  assign new_n1532_ = ~new_n1482_ & new_n1530_;
  assign new_n1533_ = new_n1531_ & new_n1532_;
  assign new_n1534_ = ~new_n895_ & new_n1487_;
  assign new_n1535_ = ~new_n1486_ & new_n1534_;
  assign new_n1536_ = new_n581_ & new_n1502_;
  assign new_n1537_ = new_n1535_ & new_n1536_;
  assign new_n1538_ = ~new_n1482_ & new_n1537_;
  assign new_n1539_ = ~new_n1527_ & ~new_n1533_;
  assign new_n1540_ = ~new_n1538_ & new_n1539_;
  assign new_n1541_ = new_n1507_ & new_n1521_;
  assign new_n1542_ = new_n1540_ & new_n1541_;
  assign new_n1543_ = nn1312gat & ~nn2169gat;
  assign new_n1544_ = ~new_n1471_ & new_n1543_;
  assign n182 = new_n1542_ & new_n1544_;
  assign new_n1546_ = nn2061gat & nn1899gat;
  assign new_n1547_ = ~nn2139gat & new_n1546_;
  assign new_n1548_ = nn1850gat & new_n1547_;
  assign n197 = nn2143gat & new_n1548_;
  assign new_n1550_ = nn2403gat & nn2440gat;
  assign new_n1551_ = ~nn2394gat & new_n1550_;
  assign new_n1552_ = ~nn2347gat & new_n1551_;
  assign new_n1553_ = ~nn2407gat & new_n1552_;
  assign new_n1554_ = new_n1480_ & ~new_n1553_;
  assign new_n1555_ = new_n1542_ & new_n1554_;
  assign n227 = n892 & new_n1555_;
  assign new_n1557_ = nn1775gat & ~nn1312gat;
  assign new_n1558_ = new_n1542_ & ~new_n1557_;
  assign new_n1559_ = ~new_n1471_ & new_n1558_;
  assign n257 = ~new_n1363_ & new_n1559_;
  assign new_n1561_ = new_n895_ & new_n1213_;
  assign n907 = ~nn2454gat & new_n1561_;
  assign new_n1563_ = ~n872 & ~n907;
  assign n277 = n212 | ~new_n1563_;
  assign new_n1565_ = nn2403gat & nn2394gat;
  assign new_n1566_ = ~nn2440gat & new_n1565_;
  assign new_n1567_ = ~nn2407gat & ~nn2347gat;
  assign new_n1568_ = new_n1566_ & new_n1567_;
  assign new_n1569_ = ~n892 & new_n1568_;
  assign new_n1570_ = n892 & new_n1553_;
  assign new_n1571_ = ~new_n1569_ & ~new_n1570_;
  assign new_n1572_ = ~nn1496gat & ~nn2091gat;
  assign new_n1573_ = ~n892 & new_n1572_;
  assign new_n1574_ = nn2143gat & nn2139gat;
  assign new_n1575_ = nn1850gat & new_n1574_;
  assign new_n1576_ = ~nn1899gat & new_n1575_;
  assign n452 = ~nn2061gat & new_n1576_;
  assign new_n1578_ = new_n1573_ & n452;
  assign new_n1579_ = ~nn2061gat & ~nn2139gat;
  assign new_n1580_ = nn1850gat & new_n1579_;
  assign new_n1581_ = ~nn2143gat & new_n1580_;
  assign n527 = ~nn1899gat & new_n1581_;
  assign new_n1583_ = nn1740gat & n892;
  assign new_n1584_ = n527 & new_n1583_;
  assign new_n1585_ = ~nn1740gat & n892;
  assign new_n1586_ = new_n1480_ & new_n1585_;
  assign new_n1587_ = ~new_n1583_ & ~new_n1585_;
  assign new_n1588_ = ~new_n1573_ & new_n1587_;
  assign new_n1589_ = new_n1474_ & new_n1588_;
  assign new_n1590_ = ~new_n1578_ & ~new_n1584_;
  assign new_n1591_ = ~new_n1586_ & new_n1590_;
  assign new_n1592_ = ~new_n1589_ & new_n1591_;
  assign new_n1593_ = ~nn2182gat & ~new_n1571_;
  assign new_n1594_ = ~new_n1592_ & new_n1593_;
  assign new_n1595_ = ~nn2135gat & ~nn2262gat;
  assign new_n1596_ = ~nn2190gat & new_n1595_;
  assign new_n1597_ = ~nn2179gat & new_n1596_;
  assign new_n1598_ = ~new_n1571_ & new_n1597_;
  assign new_n1599_ = ~new_n1592_ & new_n1598_;
  assign n282 = new_n1594_ | new_n1599_;
  assign n287 = ~nn2588gat | ~new_n1468_;
  assign new_n1602_ = nn2440gat & new_n1565_;
  assign new_n1603_ = ~nn2407gat & new_n1602_;
  assign new_n1604_ = nn2347gat & new_n1603_;
  assign new_n1605_ = nn2143gat & nn2061gat;
  assign new_n1606_ = nn2139gat & new_n1605_;
  assign new_n1607_ = nn1850gat & new_n1606_;
  assign new_n1608_ = ~nn1899gat & new_n1607_;
  assign n297 = new_n1604_ & new_n1608_;
  assign new_n1610_ = ~new_n1212_ & ~new_n1325_;
  assign new_n1611_ = ~new_n1215_ & new_n1610_;
  assign n302 = new_n1207_ | ~new_n1611_;
  assign new_n1613_ = new_n767_1_ & new_n768_;
  assign new_n1614_ = new_n769_ & new_n1613_;
  assign new_n1615_ = pn3094gat & new_n1614_;
  assign new_n1616_ = pn3085gat & pn3086gat;
  assign new_n1617_ = pn3087gat & ~pn3088gat;
  assign new_n1618_ = new_n776_ & new_n1616_;
  assign new_n1619_ = new_n1617_ & new_n1618_;
  assign new_n1620_ = ~new_n1437_ & new_n1619_;
  assign n307 = new_n1615_ | new_n1620_;
  assign n352 = ~new_n1363_ & new_n1542_;
  assign n372 = nn1312gat & new_n1608_;
  assign new_n1624_ = nn2562gat & new_n1288_;
  assign new_n1625_ = nn2343gat & new_n1624_;
  assign new_n1626_ = nn2399gat & new_n1625_;
  assign n402 = new_n1402_ & new_n1626_;
  assign new_n1628_ = ~nn2403gat & ~nn2440gat;
  assign new_n1629_ = nn2394gat & new_n1628_;
  assign new_n1630_ = nn2407gat & new_n1629_;
  assign new_n1631_ = ~nn2347gat & new_n1630_;
  assign n407 = n527 & new_n1631_;
  assign n422 = new_n1462_ & n907;
  assign n427 = new_n1474_ & new_n1631_;
  assign new_n1635_ = nn1899gat & new_n1446_;
  assign new_n1636_ = nn1850gat & new_n1635_;
  assign n442 = nn2139gat & new_n1636_;
  assign new_n1638_ = ~nn1899gat & nn1850gat;
  assign new_n1639_ = nn2139gat & new_n1638_;
  assign new_n1640_ = ~nn2143gat & new_n1639_;
  assign new_n1641_ = nn2061gat & new_n1640_;
  assign n467 = n892 & new_n1641_;
  assign n477 = new_n1474_ & new_n1542_;
  assign new_n1644_ = ~nn1775gat & ~nn1316gat;
  assign n487 = ~nn2040gat & new_n1644_;
  assign n502 = new_n1458_ & n442;
  assign new_n1647_ = nn2099gat & ~new_n1363_;
  assign new_n1648_ = nn2095gat & ~new_n1471_;
  assign new_n1649_ = ~new_n1647_ & new_n1648_;
  assign n627 = nn2037gat & new_n1649_;
  assign n742 = new_n1592_ & n627;
  assign n532 = ~new_n1436_ & n742;
  assign new_n1653_ = new_n773_ & new_n1618_;
  assign new_n1654_ = ~new_n1437_ & new_n1653_;
  assign new_n1655_ = new_n769_ & new_n770_;
  assign new_n1656_ = pn3094gat & new_n1655_;
  assign new_n1657_ = ~new_n1654_ & ~new_n1656_;
  assign new_n1658_ = pn3068gat & ~new_n1657_;
  assign new_n1659_ = ~nn2626gat & ~nn2622gat;
  assign new_n1660_ = nn2490gat & new_n1659_;
  assign new_n1661_ = new_n1401_ & new_n1660_;
  assign new_n1662_ = nn2155gat & new_n1661_;
  assign new_n1663_ = ~nn2622gat & ~nn2490gat;
  assign new_n1664_ = nn2626gat & new_n1663_;
  assign new_n1665_ = nn2630gat & ~nn2543gat;
  assign new_n1666_ = new_n1664_ & new_n1665_;
  assign new_n1667_ = ~nn2155gat & new_n1666_;
  assign new_n1668_ = ~new_n1662_ & ~new_n1667_;
  assign new_n1669_ = ~new_n1350_ & ~new_n1668_;
  assign new_n1670_ = ~new_n1398_ & new_n1669_;
  assign new_n1671_ = ~nn2207gat & new_n1670_;
  assign new_n1672_ = n337 & new_n1671_;
  assign n537 = new_n1658_ | new_n1672_;
  assign new_n1674_ = pn3093gat & ~new_n1672_;
  assign new_n1675_ = pn3068gat & new_n1674_;
  assign new_n1676_ = pn3095gat & ~new_n1672_;
  assign new_n1677_ = pn3077gat & new_n1676_;
  assign new_n1678_ = ~new_n1675_ & ~new_n1677_;
  assign n542 = new_n1672_ | ~new_n1678_;
  assign n557 = ~new_n1449_ & n742;
  assign new_n1681_ = pn3072gat & ~new_n1657_;
  assign n562 = new_n1672_ | new_n1681_;
  assign new_n1683_ = pn3070gat & new_n1674_;
  assign new_n1684_ = pn3079gat & new_n1676_;
  assign new_n1685_ = ~new_n1672_ & ~new_n1683_;
  assign n567 = new_n1684_ | ~new_n1685_;
  assign n572 = ~new_n579_ & n627;
  assign n582 = ~nn2454gat & ~nn271gat;
  assign new_n1689_ = pn3069gat & ~new_n1657_;
  assign n587 = new_n1672_ | new_n1689_;
  assign new_n1691_ = pn3071gat & new_n1674_;
  assign new_n1692_ = pn3080gat & new_n1676_;
  assign new_n1693_ = ~new_n1691_ & ~new_n1692_;
  assign n592 = new_n1672_ | ~new_n1693_;
  assign n597 = ~new_n793_ & n627;
  assign new_n1696_ = pn3081gat & pn3095gat;
  assign new_n1697_ = pn3093gat & pn3072gat;
  assign n607 = new_n1696_ | new_n1697_;
  assign new_n1699_ = nn2117gat & ~new_n1460_;
  assign n612 = ~nn2125gat & new_n1699_;
  assign new_n1701_ = pn3070gat & ~new_n1657_;
  assign n617 = new_n1672_ | new_n1701_;
  assign new_n1703_ = pn3072gat & new_n1674_;
  assign new_n1704_ = pn3081gat & new_n1676_;
  assign new_n1705_ = ~new_n1672_ & ~new_n1703_;
  assign n622 = new_n1704_ | ~new_n1705_;
  assign new_n1707_ = pn3082gat & pn3095gat;
  assign new_n1708_ = pn3093gat & pn3073gat;
  assign n642 = new_n1707_ | new_n1708_;
  assign new_n1710_ = ~new_n769_ & new_n1613_;
  assign new_n1711_ = pn3094gat & new_n1710_;
  assign new_n1712_ = pn3074gat & new_n1711_;
  assign new_n1713_ = new_n772_1_ & new_n776_;
  assign new_n1714_ = new_n1617_ & new_n1713_;
  assign new_n1715_ = ~new_n1437_ & new_n1714_;
  assign new_n1716_ = pn3065gat & new_n1715_;
  assign n647 = new_n1712_ | new_n1716_;
  assign n802 = new_n1571_ & n627;
  assign n652 = ~new_n584_ & n802;
  assign n662 = new_n893_ & new_n1205_;
  assign new_n1721_ = pn3095gat & pn3080gat;
  assign new_n1722_ = pn3093gat & pn3071gat;
  assign n667 = new_n1721_ | new_n1722_;
  assign new_n1724_ = pn3076gat & new_n1711_;
  assign new_n1725_ = pn3067gat & new_n1715_;
  assign n672 = new_n1724_ | new_n1725_;
  assign n677 = ~new_n589_ & n802;
  assign new_n1728_ = n892 & new_n1480_;
  assign new_n1729_ = ~new_n1475_ & ~new_n1728_;
  assign n682 = new_n1458_ & ~new_n1729_;
  assign new_n1731_ = pn3095gat & pn3079gat;
  assign new_n1732_ = pn3070gat & pn3093gat;
  assign n692 = new_n1731_ | new_n1732_;
  assign new_n1734_ = pn3087gat & pn3088gat;
  assign new_n1735_ = new_n1713_ & new_n1734_;
  assign new_n1736_ = ~new_n1437_ & new_n1735_;
  assign new_n1737_ = ~new_n1711_ & ~new_n1736_;
  assign new_n1738_ = pn3068gat & ~new_n1737_;
  assign new_n1739_ = nn156gat & new_n1329_;
  assign new_n1740_ = ~nn156gat & ~new_n1329_;
  assign new_n1741_ = ~new_n1739_ & ~new_n1740_;
  assign new_n1742_ = new_n1737_ & ~new_n1741_;
  assign n697 = new_n1738_ | new_n1742_;
  assign n707 = ~pn3099gat & nn2319gat;
  assign new_n1745_ = pn3095gat & pn3077gat;
  assign new_n1746_ = pn3093gat & pn3068gat;
  assign n712 = new_n1745_ | new_n1746_;
  assign new_n1748_ = ~new_n1711_ & ~new_n1715_;
  assign new_n1749_ = nn327gat & ~nn384gat;
  assign new_n1750_ = ~nn331gat & ~nn388gat;
  assign new_n1751_ = new_n1331_ & new_n1750_;
  assign new_n1752_ = ~nn384gat & ~new_n1751_;
  assign new_n1753_ = ~nn327gat & new_n1751_;
  assign new_n1754_ = nn384gat & new_n1753_;
  assign new_n1755_ = ~new_n1749_ & ~new_n1752_;
  assign new_n1756_ = ~new_n1754_ & new_n1755_;
  assign new_n1757_ = new_n1748_ & ~new_n1756_;
  assign new_n1758_ = pn3069gat & new_n1715_;
  assign new_n1759_ = pn3078gat & new_n1711_;
  assign new_n1760_ = ~new_n1757_ & ~new_n1758_;
  assign n722 = new_n1759_ | ~new_n1760_;
  assign new_n1762_ = nn388gat & new_n1331_;
  assign new_n1763_ = nn327gat & new_n1331_;
  assign new_n1764_ = ~nn331gat & new_n1763_;
  assign new_n1765_ = ~new_n1762_ & ~new_n1764_;
  assign new_n1766_ = nn463gat & ~new_n1765_;
  assign new_n1767_ = ~nn463gat & new_n1765_;
  assign new_n1768_ = ~new_n1766_ & ~new_n1767_;
  assign new_n1769_ = new_n1748_ & ~new_n1768_;
  assign new_n1770_ = pn3073gat & new_n1715_;
  assign new_n1771_ = pn3082gat & new_n1711_;
  assign new_n1772_ = ~new_n1769_ & ~new_n1770_;
  assign n737 = new_n1771_ | ~new_n1772_;
  assign new_n1774_ = pn3066gat & ~new_n1657_;
  assign n747 = new_n1672_ | new_n1774_;
  assign new_n1776_ = pn3066gat & new_n1674_;
  assign new_n1777_ = pn3075gat & new_n1676_;
  assign new_n1778_ = ~new_n1672_ & ~new_n1776_;
  assign n752 = new_n1777_ | ~new_n1778_;
  assign new_n1780_ = pn3095gat & pn3078gat;
  assign new_n1781_ = pn3093gat & pn3069gat;
  assign n762 = new_n1780_ | new_n1781_;
  assign new_n1783_ = ~nn388gat & ~new_n1331_;
  assign new_n1784_ = ~new_n1762_ & ~new_n1783_;
  assign new_n1785_ = new_n1748_ & ~new_n1784_;
  assign new_n1786_ = pn3072gat & new_n1715_;
  assign new_n1787_ = pn3081gat & new_n1711_;
  assign new_n1788_ = ~new_n1785_ & ~new_n1786_;
  assign n767 = new_n1787_ | ~new_n1788_;
  assign n772 = ~new_n1076_ & n802;
  assign new_n1791_ = pn3071gat & ~new_n1657_;
  assign n777 = new_n1672_ | new_n1791_;
  assign new_n1793_ = pn3076gat & new_n1676_;
  assign new_n1794_ = pn3067gat & new_n1674_;
  assign new_n1795_ = ~new_n1672_ & ~new_n1793_;
  assign n782 = new_n1794_ | ~new_n1795_;
  assign new_n1797_ = ~nn152gat & ~new_n1329_;
  assign new_n1798_ = nn156gat & ~nn152gat;
  assign new_n1799_ = nn152gat & new_n1329_;
  assign new_n1800_ = ~nn156gat & new_n1799_;
  assign new_n1801_ = ~new_n1797_ & ~new_n1798_;
  assign new_n1802_ = ~new_n1800_ & new_n1801_;
  assign new_n1803_ = new_n1737_ & ~new_n1802_;
  assign new_n1804_ = pn3067gat & ~new_n1737_;
  assign n792 = new_n1803_ | new_n1804_;
  assign new_n1806_ = pn3066gat & new_n1715_;
  assign new_n1807_ = pn3075gat & new_n1711_;
  assign n797 = new_n1806_ | new_n1807_;
  assign new_n1809_ = pn3095gat & pn3074gat;
  assign new_n1810_ = pn3093gat & pn3065gat;
  assign n817 = new_n1809_ | new_n1810_;
  assign new_n1812_ = pn3065gat & ~new_n1737_;
  assign new_n1813_ = ~nn148gat & nn256gat;
  assign new_n1814_ = ~nn156gat & new_n1329_;
  assign new_n1815_ = ~nn152gat & new_n1814_;
  assign new_n1816_ = ~nn148gat & ~new_n1815_;
  assign new_n1817_ = nn148gat & new_n1815_;
  assign new_n1818_ = ~nn256gat & new_n1817_;
  assign new_n1819_ = ~new_n1813_ & ~new_n1816_;
  assign new_n1820_ = ~new_n1818_ & new_n1819_;
  assign new_n1821_ = new_n1737_ & ~new_n1820_;
  assign n822 = new_n1812_ | new_n1821_;
  assign new_n1823_ = ~nn331gat & nn388gat;
  assign new_n1824_ = ~nn331gat & ~new_n1331_;
  assign new_n1825_ = ~nn388gat & new_n1331_;
  assign new_n1826_ = nn331gat & new_n1825_;
  assign new_n1827_ = ~new_n1823_ & ~new_n1824_;
  assign new_n1828_ = ~new_n1826_ & new_n1827_;
  assign new_n1829_ = new_n1748_ & ~new_n1828_;
  assign new_n1830_ = pn3080gat & new_n1711_;
  assign new_n1831_ = pn3071gat & new_n1715_;
  assign new_n1832_ = ~new_n1829_ & ~new_n1830_;
  assign n827 = new_n1831_ | ~new_n1832_;
  assign n832 = ~new_n1091_ & n802;
  assign new_n1835_ = ~nn2266gat & new_n790_;
  assign new_n1836_ = nn2266gat & ~new_n790_;
  assign new_n1837_ = ~new_n1835_ & ~new_n1836_;
  assign n837 = ~n627 | ~new_n1837_;
  assign new_n1839_ = pn3093gat & pn3067gat;
  assign new_n1840_ = pn3095gat & pn3076gat;
  assign n847 = new_n1839_ | new_n1840_;
  assign new_n1842_ = pn3073gat & ~new_n1737_;
  assign new_n1843_ = ~nn152gat & nn256gat;
  assign new_n1844_ = new_n1329_ & new_n1843_;
  assign new_n1845_ = ~new_n1739_ & ~new_n1844_;
  assign new_n1846_ = ~nn470gat & new_n1845_;
  assign new_n1847_ = nn470gat & ~new_n1845_;
  assign new_n1848_ = ~new_n1846_ & ~new_n1847_;
  assign new_n1849_ = new_n1737_ & ~new_n1848_;
  assign n852 = new_n1842_ | new_n1849_;
  assign n857 = new_n1462_ & n582;
  assign new_n1852_ = nn2476gat & nn2599gat;
  assign new_n1853_ = nn2518gat & new_n1852_;
  assign new_n1854_ = ~pn3090gat & nn2526gat;
  assign new_n1855_ = nn2476gat & new_n1854_;
  assign new_n1856_ = nn2464gat & new_n1855_;
  assign new_n1857_ = nn2468gat & new_n1856_;
  assign n867 = ~new_n1853_ | ~new_n1857_;
  assign new_n1859_ = pn3093gat & pn3066gat;
  assign new_n1860_ = pn3095gat & pn3075gat;
  assign n882 = new_n1859_ | new_n1860_;
  assign new_n1862_ = pn3066gat & ~new_n1737_;
  assign new_n1863_ = ~nn256gat & ~new_n1815_;
  assign new_n1864_ = nn256gat & new_n1815_;
  assign new_n1865_ = ~new_n1863_ & ~new_n1864_;
  assign new_n1866_ = new_n1737_ & ~new_n1865_;
  assign n887 = new_n1862_ | new_n1866_;
  assign new_n1868_ = pn3073gat & ~new_n1657_;
  assign n897 = new_n1672_ | new_n1868_;
  assign new_n1870_ = nn2403gat & ~nn2394gat;
  assign new_n1871_ = ~nn2440gat & ~new_n1870_;
  assign new_n1872_ = ~new_n1073_ & new_n1871_;
  assign new_n1873_ = nn2644gat & ~new_n1872_;
  assign new_n1874_ = ~nn2644gat & new_n1872_;
  assign new_n1875_ = ~new_n1873_ & ~new_n1874_;
  assign n902 = ~n802 | ~new_n1875_;
  assign new_n1877_ = pn3068gat & new_n1715_;
  assign new_n1878_ = pn3077gat & new_n1711_;
  assign n917 = new_n1877_ | new_n1878_;
  assign n922 = ~new_n798_ & n742;
  assign new_n1881_ = pn3065gat & ~new_n1657_;
  assign n927 = new_n1672_ | new_n1881_;
  assign new_n1883_ = pn3074gat & new_n1676_;
  assign new_n1884_ = pn3065gat & new_n1674_;
  assign new_n1885_ = ~new_n1672_ & ~new_n1883_;
  assign n932 = new_n1884_ | ~new_n1885_;
  assign new_n1887_ = pn3069gat & new_n1674_;
  assign new_n1888_ = pn3078gat & new_n1676_;
  assign new_n1889_ = ~new_n1672_ & ~new_n1887_;
  assign n937 = new_n1888_ | ~new_n1889_;
  assign new_n1891_ = ~nn327gat & ~new_n1751_;
  assign new_n1892_ = nn327gat & new_n1751_;
  assign new_n1893_ = ~new_n1891_ & ~new_n1892_;
  assign new_n1894_ = new_n1748_ & ~new_n1893_;
  assign new_n1895_ = pn3070gat & new_n1715_;
  assign new_n1896_ = pn3079gat & new_n1711_;
  assign new_n1897_ = ~new_n1894_ & ~new_n1895_;
  assign n952 = new_n1896_ | ~new_n1897_;
  assign n957 = ~new_n782_1_ & n742;
  assign new_n1900_ = pn3067gat & ~new_n1657_;
  assign n962 = new_n1672_ | new_n1900_;
  assign new_n1902_ = pn3073gat & new_n1674_;
  assign new_n1903_ = pn3082gat & new_n1676_;
  assign new_n1904_ = ~new_n1672_ & ~new_n1902_;
  assign n967 = new_n1903_ | ~new_n1904_;
  assign new_n1906_ = nn2061gat & ~nn2139gat;
  assign new_n1907_ = ~nn1899gat & ~new_n1906_;
  assign new_n1908_ = ~new_n1433_ & new_n1907_;
  assign new_n1909_ = nn1975gat & ~new_n1908_;
  assign new_n1910_ = ~nn1975gat & new_n1908_;
  assign new_n1911_ = ~new_n1909_ & ~new_n1910_;
  assign n977 = ~n742 | ~new_n1911_;
  assign pn3112gat = 1'b1;
  assign pn3152gat = 1'b1;
  assign pn3115gat = 1'b1;
  assign n327 = 1'b1;
  assign pn3128gat = ~nn2390gat;
  assign pn3126gat = ~nn2339gat;
  assign pn3127gat = ~nn2270gat;
  assign pn3148gat = ~nn2450gat;
  assign pn3106gat = ~nn1871gat;
  assign n187 = ~nn2121gat;
  assign n192 = ~nn830gat;
  assign n202 = ~nn1332gat;
  assign n207 = ~nn1363gat;
  assign n217 = ~nn2125gat;
  assign n222 = ~nn834gat;
  assign n237 = ~nn1775gat;
  assign n242 = ~nn2095gat;
  assign n247 = ~nn2110gat;
  assign n262 = ~nn2176gat;
  assign n267 = ~nn2033gat;
  assign n292 = ~nn2037gat;
  assign n312 = ~nn2495gat;
  assign n317 = ~nn1394gat;
  assign n322 = ~nn1316gat;
  assign n332 = ~nn2025gat;
  assign n342 = ~nn1433gat;
  assign n347 = ~nn2309gat;
  assign n362 = ~nn614gat;
  assign n367 = ~nn2458gat;
  assign n382 = ~nn707gat;
  assign n387 = ~nn2592gat;
  assign n397 = ~nn824gat;
  assign n417 = ~nn883gat;
  assign n447 = ~nn820gat;
  assign n472 = ~nn684gat;
  assign n492 = ~nn2640gat;
  assign n497 = ~nn699gat;
  assign n512 = ~nn2044gat;
  assign n517 = ~nn2634gat;
  assign n522 = ~nn838gat;
  assign n552 = ~nn2399gat;
  assign n577 = ~nn2343gat;
  assign n602 = ~nn2562gat;
  assign n632 = ~nn2207gat;
  assign n657 = ~nn2203gat;
  assign n687 = ~nn2472gat;
  assign n727 = ~nn1821gat;
  assign n757 = ~nn2029gat;
  assign n812 = ~nn2543gat;
  assign n877 = ~nn2622gat;
  assign n912 = ~nn2490gat;
  assign n947 = ~nn2626gat;
  assign n982 = ~nn2630gat;
  assign pn3141gat = pn3142gat;
  assign n252 = pn3127gat;
  assign n272 = pn3073gat;
  assign n377 = pn3065gat;
  assign n392 = pn3067gat;
  assign n412 = pn3066gat;
  assign n432 = pn3069gat;
  assign n437 = pn3126gat;
  assign n457 = pn3070gat;
  assign n462 = pn3128gat;
  assign n482 = pn3072gat;
  assign n507 = pn3071gat;
  assign n637 = pn3068gat;
  assign n842 = pn3149gat;
  always @ (posedge clock) begin
    nn1332gat <= n172;
    nn1775gat <= n177;
    nn2454gat <= n182;
    nn2117gat <= n187;
    nn470gat <= n192;
    nn1525gat <= n197;
    nn1740gat <= n202;
    nn1312gat <= n207;
    nn2040gat <= n212;
    nn2121gat <= n217;
    nn148gat <= n222;
    nn1456gat <= n227;
    nn2179gat <= n232;
    nn2592gat <= n237;
    nn2176gat <= n242;
    nn2125gat <= n247;
    nn2190gat <= n252;
    nn1871gat <= n257;
    nn2169gat <= n262;
    nn2110gat <= n267;
    nn842gat <= n272;
    nn2021gat <= n277;
    nn1433gat <= n282;
    nn2446gat <= n287;
    nn2033gat <= n292;
    nn1394gat <= n297;
    nn2182gat <= n302;
    nn2095gat <= n307;
    nn2266gat <= n312;
    nn1496gat <= n317;
    nn1363gat <= n322;
    nn2309gat <= n327;
    nn2099gat <= n332;
    nn2091gat <= n337;
    nn1316gat <= n342;
    nn2450gat <= n347;
    nn2025gat <= n352;
    nn2510gat <= n357;
    nn156gat <= n362;
    nn2514gat <= n367;
    nn1588gat <= n372;
    nn271gat <= n377;
    nn152gat <= n382;
    nn2458gat <= n387;
    nn160gat <= n392;
    nn331gat <= n397;
    nn1336gat <= n402;
    nn1462gat <= n407;
    nn337gat <= n412;
    nn388gat <= n417;
    nn1771gat <= n422;
    nn1596gat <= n427;
    nn398gat <= n432;
    nn2135gat <= n437;
    nn1678gat <= n442;
    nn463gat <= n447;
    nn1675gat <= n452;
    nn402gat <= n457;
    nn2262gat <= n462;
    nn1508gat <= n467;
    nn327gat <= n472;
    nn1748gat <= n477;
    nn919gat <= n482;
    nn2044gat <= n487;
    nn2644gat <= n492;
    nn384gat <= n497;
    nn1340gat <= n502;
    nn846gat <= n507;
    nn2037gat <= n512;
    nn1975gat <= n517;
    nn256gat <= n522;
    nn1807gat <= n527;
    nn2630gat <= n532;
    nn931gat <= n537;
    nn322gat <= n542;
    nn2502gat <= n547;
    nn2403gat <= n552;
    nn2543gat <= n557;
    nn1226gat <= n562;
    nn318gat <= n567;
    nn2339gat <= n572;
    nn2394gat <= n577;
    nn2102gat <= n582;
    nn1045gat <= n587;
    nn561gat <= n592;
    nn2270gat <= n597;
    nn2440gat <= n602;
    nn673gat <= n607;
    nn1880gat <= n612;
    nn1135gat <= n617;
    nn366gat <= n622;
    nn2390gat <= n627;
    nn2407gat <= n632;
    nn341gat <= n637;
    nn1241gat <= n642;
    nn680gat <= n647;
    nn2343gat <= n652;
    nn2347gat <= n657;
    nn2472gat <= n662;
    nn1294gat <= n667;
    nn816gat <= n672;
    nn2399gat <= n677;
    nn1389gat <= n682;
    nn2319gat <= n687;
    nn1080gat <= n692;
    nn614gat <= n697;
    nn2464gat <= n702;
    nn1821gat <= n707;
    nn865gat <= n712;
    nn2526gat <= n717;
    nn699gat <= n722;
    nn2029gat <= n727;
    nn2468gat <= n732;
    nn820gat <= n737;
    nn2626gat <= n742;
    nn1072gat <= n747;
    nn777gat <= n752;
    nn1829gat <= n757;
    nn1148gat <= n762;
    nn883gat <= n767;
    nn2207gat <= n772;
    nn1282gat <= n777;
    nn553gat <= n782;
    nn2476gat <= n787;
    nn707gat <= n792;
    nn580gat <= n797;
    nn2562gat <= n802;
    nn2658gat <= n807;
    nn2143gat <= n812;
    nn1068gat <= n817;
    nn834gat <= n822;
    nn824gat <= n827;
    nn2203gat <= n832;
    nn2495gat <= n837;
    nn2084gat <= n842;
    nn957gat <= n847;
    nn830gat <= n852;
    nn1763gat <= n857;
    nn2518gat <= n862;
    nn2588gat <= n867;
    nn1767gat <= n872;
    nn2061gat <= n877;
    nn861gat <= n882;
    nn838gat <= n887;
    nn2155gat <= n892;
    nn1197gat <= n897;
    nn2640gat <= n902;
    nn1834gat <= n907;
    nn2139gat <= n912;
    nn584gat <= n917;
    nn2622gat <= n922;
    nn1035gat <= n927;
    nn659gat <= n932;
    nn314gat <= n937;
    nn2506gat <= n942;
    nn1899gat <= n947;
    nn684gat <= n952;
    nn2490gat <= n957;
    nn1121gat <= n962;
    nn667gat <= n967;
    nn2599gat <= n972;
    nn2634gat <= n977;
    nn1850gat <= n982;
  end
endmodule

