module top ( 
    _1gat_0_, _85gat_17_, _135gat_32_, _152gat_37_, _210gat_49_,
    _259gat_55_, _36gat_6_, _55gat_9_, _75gat_15_, _159gat_40_,
    _237gat_52_, _138gat_33_, _8gat_1_, _219gat_50_, _26gat_4_, _74gat_14_,
    _153gat_38_, _59gat_10_, _207gat_48_, _261gat_57_, _88gat_20_,
    _183gat_44_, _149gat_36_, _260gat_56_, _13gat_2_, _73gat_13_,
    _116gat_28_, _130gat_31_, _246gat_53_, _89gat_21_, _111gat_27_,
    _189gat_45_, _68gat_11_, _72gat_12_, _268gat_59_, _90gat_22_,
    _143gat_34_, _201gat_47_, _267gat_58_, _101gat_25_, _171gat_42_,
    _29gat_5_, _228gat_51_, _91gat_23_, _146gat_35_, _51gat_8_, _80gat_16_,
    _87gat_19_, _165gat_41_, _255gat_54_, _156gat_39_, _177gat_43_,
    _42gat_7_, _86gat_18_, _17gat_3_, _96gat_24_, _106gat_26_, _121gat_29_,
    _195gat_46_, _126gat_30_,
    _768gat_334_, _388gat_133_, _420gat_158_, _423gat_155_, _419gat_164_,
    _850gat_404_, _389gat_132_, _767gat_349_, _874gat_433_, _418gat_168_,
    _421gat_162_, _422gat_161_, _878gat_442_, _450gat_173_, _447gat_182_,
    _879gat_441_, _449gat_176_, _863gat_424_, _446gat_183_, _866gat_426_,
    _880gat_440_, _391gat_124_, _448gat_179_, _865gat_422_, _390gat_131_,
    _864gat_423_  );
  input  _1gat_0_, _85gat_17_, _135gat_32_, _152gat_37_, _210gat_49_,
    _259gat_55_, _36gat_6_, _55gat_9_, _75gat_15_, _159gat_40_,
    _237gat_52_, _138gat_33_, _8gat_1_, _219gat_50_, _26gat_4_, _74gat_14_,
    _153gat_38_, _59gat_10_, _207gat_48_, _261gat_57_, _88gat_20_,
    _183gat_44_, _149gat_36_, _260gat_56_, _13gat_2_, _73gat_13_,
    _116gat_28_, _130gat_31_, _246gat_53_, _89gat_21_, _111gat_27_,
    _189gat_45_, _68gat_11_, _72gat_12_, _268gat_59_, _90gat_22_,
    _143gat_34_, _201gat_47_, _267gat_58_, _101gat_25_, _171gat_42_,
    _29gat_5_, _228gat_51_, _91gat_23_, _146gat_35_, _51gat_8_, _80gat_16_,
    _87gat_19_, _165gat_41_, _255gat_54_, _156gat_39_, _177gat_43_,
    _42gat_7_, _86gat_18_, _17gat_3_, _96gat_24_, _106gat_26_, _121gat_29_,
    _195gat_46_, _126gat_30_;
  output _768gat_334_, _388gat_133_, _420gat_158_, _423gat_155_, _419gat_164_,
    _850gat_404_, _389gat_132_, _767gat_349_, _874gat_433_, _418gat_168_,
    _421gat_162_, _422gat_161_, _878gat_442_, _450gat_173_, _447gat_182_,
    _879gat_441_, _449gat_176_, _863gat_424_, _446gat_183_, _866gat_426_,
    _880gat_440_, _391gat_124_, _448gat_179_, _865gat_422_, _390gat_131_,
    _864gat_423_;
  wire new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n114_, new_n116_, new_n118_, new_n120_, new_n122_, new_n123_,
    new_n124_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n179_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n265_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n337_, new_n338_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n356_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n375_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_;
  assign new_n87_ = ~_201gat_47_ & ~_195gat_46_;
  assign new_n88_ = _201gat_47_ & _195gat_46_;
  assign new_n89_ = ~new_n87_ & ~new_n88_;
  assign new_n90_ = ~_183gat_44_ & ~_189gat_45_;
  assign new_n91_ = _183gat_44_ & _189gat_45_;
  assign new_n92_ = ~new_n90_ & ~new_n91_;
  assign new_n93_ = new_n89_ & new_n92_;
  assign new_n94_ = ~new_n89_ & ~new_n92_;
  assign new_n95_ = ~new_n93_ & ~new_n94_;
  assign new_n96_ = ~_207gat_48_ & ~new_n95_;
  assign new_n97_ = _207gat_48_ & new_n95_;
  assign new_n98_ = ~new_n96_ & ~new_n97_;
  assign new_n99_ = ~_171gat_42_ & ~_177gat_43_;
  assign new_n100_ = _171gat_42_ & _177gat_43_;
  assign new_n101_ = ~new_n99_ & ~new_n100_;
  assign new_n102_ = ~_159gat_40_ & ~_165gat_41_;
  assign new_n103_ = _159gat_40_ & _165gat_41_;
  assign new_n104_ = ~new_n102_ & ~new_n103_;
  assign new_n105_ = new_n101_ & new_n104_;
  assign new_n106_ = ~new_n101_ & ~new_n104_;
  assign new_n107_ = ~new_n105_ & ~new_n106_;
  assign new_n108_ = ~_130gat_31_ & ~new_n107_;
  assign new_n109_ = _130gat_31_ & new_n107_;
  assign new_n110_ = ~new_n108_ & ~new_n109_;
  assign new_n111_ = new_n98_ & new_n110_;
  assign new_n112_ = ~new_n98_ & ~new_n110_;
  assign _768gat_334_ = ~new_n111_ & ~new_n112_;
  assign new_n114_ = _75gat_15_ & _42gat_7_;
  assign _388gat_133_ = _29gat_5_ & new_n114_;
  assign new_n116_ = _75gat_15_ & _80gat_16_;
  assign _420gat_158_ = ~_59gat_10_ | ~new_n116_;
  assign new_n118_ = ~_88gat_20_ & ~_87gat_19_;
  assign _423gat_155_ = _90gat_22_ & ~new_n118_;
  assign new_n120_ = _36gat_6_ & _42gat_7_;
  assign _390gat_131_ = _29gat_5_ & new_n120_;
  assign new_n122_ = _26gat_4_ & _17gat_3_;
  assign new_n123_ = _13gat_2_ & new_n122_;
  assign new_n124_ = _1gat_0_ & new_n123_;
  assign _419gat_164_ = _390gat_131_ | ~new_n124_;
  assign new_n126_ = _72gat_12_ & _42gat_7_;
  assign new_n127_ = _68gat_11_ & new_n126_;
  assign new_n128_ = _59gat_10_ & new_n127_;
  assign new_n129_ = _55gat_9_ & _8gat_1_;
  assign new_n130_ = _13gat_2_ & new_n129_;
  assign new_n131_ = _1gat_0_ & new_n130_;
  assign new_n132_ = new_n128_ & new_n131_;
  assign new_n133_ = _73gat_13_ & new_n132_;
  assign new_n134_ = _201gat_47_ & new_n133_;
  assign new_n135_ = _59gat_10_ & new_n114_;
  assign new_n136_ = _8gat_1_ & _17gat_3_;
  assign new_n137_ = _51gat_8_ & new_n136_;
  assign new_n138_ = _1gat_0_ & new_n137_;
  assign new_n139_ = ~new_n135_ & new_n138_;
  assign new_n140_ = _26gat_4_ & _51gat_8_;
  assign _447gat_182_ = _1gat_0_ & new_n140_;
  assign new_n142_ = _42gat_7_ & _17gat_3_;
  assign new_n143_ = ~_42gat_7_ & ~_17gat_3_;
  assign new_n144_ = ~new_n142_ & ~new_n143_;
  assign new_n145_ = _59gat_10_ & _447gat_182_;
  assign new_n146_ = _156gat_39_ & new_n145_;
  assign new_n147_ = new_n144_ & new_n146_;
  assign new_n148_ = ~new_n139_ & ~new_n147_;
  assign new_n149_ = _126gat_30_ & ~new_n148_;
  assign new_n150_ = _59gat_10_ & _156gat_39_;
  assign new_n151_ = _17gat_3_ & ~new_n150_;
  assign new_n152_ = _447gat_182_ & new_n151_;
  assign new_n153_ = _1gat_0_ & ~new_n152_;
  assign new_n154_ = _153gat_38_ & ~new_n153_;
  assign new_n155_ = ~new_n149_ & ~new_n154_;
  assign new_n156_ = _29gat_5_ & new_n116_;
  assign new_n157_ = _55gat_9_ & new_n156_;
  assign new_n158_ = _447gat_182_ & new_n157_;
  assign new_n159_ = ~_268gat_59_ & new_n158_;
  assign new_n160_ = new_n155_ & ~new_n159_;
  assign new_n161_ = _201gat_47_ & ~new_n160_;
  assign new_n162_ = _237gat_52_ & new_n161_;
  assign new_n163_ = ~_201gat_47_ & new_n160_;
  assign new_n164_ = ~new_n161_ & ~new_n163_;
  assign new_n165_ = _228gat_51_ & new_n164_;
  assign new_n166_ = ~new_n162_ & ~new_n165_;
  assign new_n167_ = _246gat_53_ & ~new_n160_;
  assign new_n168_ = _267gat_58_ & _255gat_54_;
  assign new_n169_ = ~new_n167_ & ~new_n168_;
  assign new_n170_ = _261gat_57_ & new_n164_;
  assign new_n171_ = ~_261gat_57_ & ~new_n164_;
  assign new_n172_ = ~new_n170_ & ~new_n171_;
  assign new_n173_ = _219gat_50_ & new_n172_;
  assign new_n174_ = _210gat_49_ & _121gat_29_;
  assign new_n175_ = ~new_n173_ & ~new_n174_;
  assign new_n176_ = ~new_n134_ & new_n166_;
  assign new_n177_ = new_n169_ & new_n176_;
  assign _850gat_404_ = ~new_n175_ | ~new_n177_;
  assign new_n179_ = _36gat_6_ & _80gat_16_;
  assign _389gat_132_ = _29gat_5_ & new_n179_;
  assign new_n181_ = ~_121gat_29_ & ~_126gat_30_;
  assign new_n182_ = _121gat_29_ & _126gat_30_;
  assign new_n183_ = ~new_n181_ & ~new_n182_;
  assign new_n184_ = ~_116gat_28_ & ~_111gat_27_;
  assign new_n185_ = _116gat_28_ & _111gat_27_;
  assign new_n186_ = ~new_n184_ & ~new_n185_;
  assign new_n187_ = new_n183_ & new_n186_;
  assign new_n188_ = ~new_n183_ & ~new_n186_;
  assign new_n189_ = ~new_n187_ & ~new_n188_;
  assign new_n190_ = ~_135gat_32_ & ~new_n189_;
  assign new_n191_ = _135gat_32_ & new_n189_;
  assign new_n192_ = ~new_n190_ & ~new_n191_;
  assign new_n193_ = ~_101gat_25_ & ~_106gat_26_;
  assign new_n194_ = _101gat_25_ & _106gat_26_;
  assign new_n195_ = ~new_n193_ & ~new_n194_;
  assign new_n196_ = ~_91gat_23_ & ~_96gat_24_;
  assign new_n197_ = _91gat_23_ & _96gat_24_;
  assign new_n198_ = ~new_n196_ & ~new_n197_;
  assign new_n199_ = new_n195_ & new_n198_;
  assign new_n200_ = ~new_n195_ & ~new_n198_;
  assign new_n201_ = ~new_n199_ & ~new_n200_;
  assign new_n202_ = ~_130gat_31_ & ~new_n201_;
  assign new_n203_ = _130gat_31_ & new_n201_;
  assign new_n204_ = ~new_n202_ & ~new_n203_;
  assign new_n205_ = new_n192_ & new_n204_;
  assign new_n206_ = ~new_n192_ & ~new_n204_;
  assign _767gat_349_ = ~new_n205_ & ~new_n206_;
  assign new_n208_ = _17gat_3_ & new_n156_;
  assign new_n209_ = _447gat_182_ & new_n208_;
  assign new_n210_ = ~_268gat_59_ & new_n209_;
  assign new_n211_ = _55gat_9_ & _447gat_182_;
  assign new_n212_ = ~new_n150_ & new_n211_;
  assign new_n213_ = _153gat_38_ & new_n212_;
  assign new_n214_ = ~new_n210_ & ~new_n213_;
  assign new_n215_ = _106gat_26_ & ~new_n148_;
  assign new_n216_ = _152gat_37_ & _138gat_33_;
  assign new_n217_ = ~new_n215_ & ~new_n216_;
  assign new_n218_ = new_n214_ & new_n217_;
  assign new_n219_ = _177gat_43_ & ~new_n218_;
  assign new_n220_ = _237gat_52_ & new_n219_;
  assign new_n221_ = ~_177gat_43_ & new_n218_;
  assign new_n222_ = ~new_n219_ & ~new_n221_;
  assign new_n223_ = _228gat_51_ & new_n222_;
  assign new_n224_ = ~new_n220_ & ~new_n223_;
  assign new_n225_ = _177gat_43_ & new_n133_;
  assign new_n226_ = _246gat_53_ & ~new_n218_;
  assign new_n227_ = ~new_n225_ & ~new_n226_;
  assign new_n228_ = _111gat_27_ & ~new_n148_;
  assign new_n229_ = _143gat_34_ & ~new_n153_;
  assign new_n230_ = ~new_n228_ & ~new_n229_;
  assign new_n231_ = ~new_n159_ & new_n230_;
  assign new_n232_ = _183gat_44_ & ~new_n231_;
  assign new_n233_ = _121gat_29_ & ~new_n148_;
  assign new_n234_ = _149gat_36_ & ~new_n153_;
  assign new_n235_ = ~new_n233_ & ~new_n234_;
  assign new_n236_ = ~new_n159_ & new_n235_;
  assign new_n237_ = ~_195gat_46_ & new_n236_;
  assign new_n238_ = _116gat_28_ & ~new_n148_;
  assign new_n239_ = _146gat_35_ & ~new_n153_;
  assign new_n240_ = ~new_n238_ & ~new_n239_;
  assign new_n241_ = ~new_n159_ & new_n240_;
  assign new_n242_ = ~_189gat_45_ & new_n241_;
  assign new_n243_ = _261gat_57_ & ~new_n237_;
  assign new_n244_ = ~new_n163_ & new_n243_;
  assign new_n245_ = ~new_n242_ & new_n244_;
  assign new_n246_ = _195gat_46_ & ~new_n236_;
  assign new_n247_ = ~new_n242_ & new_n246_;
  assign new_n248_ = new_n161_ & ~new_n237_;
  assign new_n249_ = ~new_n242_ & new_n248_;
  assign new_n250_ = _189gat_45_ & ~new_n241_;
  assign new_n251_ = ~new_n245_ & ~new_n247_;
  assign new_n252_ = ~new_n249_ & new_n251_;
  assign new_n253_ = ~new_n250_ & new_n252_;
  assign new_n254_ = ~_183gat_44_ & new_n231_;
  assign new_n255_ = ~new_n253_ & ~new_n254_;
  assign new_n256_ = ~new_n232_ & ~new_n255_;
  assign new_n257_ = new_n222_ & ~new_n256_;
  assign new_n258_ = ~new_n222_ & new_n256_;
  assign new_n259_ = ~new_n257_ & ~new_n258_;
  assign new_n260_ = _219gat_50_ & new_n259_;
  assign new_n261_ = _210gat_49_ & _101gat_25_;
  assign new_n262_ = ~new_n260_ & ~new_n261_;
  assign new_n263_ = new_n224_ & new_n227_;
  assign _874gat_433_ = ~new_n262_ | ~new_n263_;
  assign new_n265_ = _13gat_2_ & new_n136_;
  assign _418gat_168_ = _1gat_0_ & new_n265_;
  assign _421gat_162_ = ~_59gat_10_ | ~new_n179_;
  assign _422gat_161_ = ~_59gat_10_ | ~new_n120_;
  assign new_n269_ = _143gat_34_ & new_n212_;
  assign new_n270_ = ~new_n210_ & ~new_n269_;
  assign new_n271_ = _91gat_23_ & ~new_n148_;
  assign new_n272_ = _138gat_33_ & _8gat_1_;
  assign new_n273_ = ~new_n271_ & ~new_n272_;
  assign new_n274_ = new_n270_ & new_n273_;
  assign new_n275_ = _159gat_40_ & ~new_n274_;
  assign new_n276_ = _237gat_52_ & new_n275_;
  assign new_n277_ = ~_159gat_40_ & new_n274_;
  assign new_n278_ = ~new_n275_ & ~new_n277_;
  assign new_n279_ = _228gat_51_ & new_n278_;
  assign new_n280_ = ~new_n276_ & ~new_n279_;
  assign new_n281_ = _159gat_40_ & new_n133_;
  assign new_n282_ = _246gat_53_ & ~new_n274_;
  assign new_n283_ = ~new_n281_ & ~new_n282_;
  assign new_n284_ = _149gat_36_ & new_n212_;
  assign new_n285_ = ~new_n210_ & ~new_n284_;
  assign new_n286_ = _101gat_25_ & ~new_n148_;
  assign new_n287_ = _138gat_33_ & _17gat_3_;
  assign new_n288_ = ~new_n286_ & ~new_n287_;
  assign new_n289_ = new_n285_ & new_n288_;
  assign new_n290_ = ~_171gat_42_ & new_n289_;
  assign new_n291_ = _146gat_35_ & new_n212_;
  assign new_n292_ = ~new_n210_ & ~new_n291_;
  assign new_n293_ = _96gat_24_ & ~new_n148_;
  assign new_n294_ = _138gat_33_ & _51gat_8_;
  assign new_n295_ = ~new_n293_ & ~new_n294_;
  assign new_n296_ = new_n292_ & new_n295_;
  assign new_n297_ = ~_165gat_41_ & new_n296_;
  assign new_n298_ = ~new_n256_ & ~new_n290_;
  assign new_n299_ = ~new_n221_ & new_n298_;
  assign new_n300_ = ~new_n297_ & new_n299_;
  assign new_n301_ = _171gat_42_ & ~new_n289_;
  assign new_n302_ = ~new_n297_ & new_n301_;
  assign new_n303_ = new_n219_ & ~new_n290_;
  assign new_n304_ = ~new_n297_ & new_n303_;
  assign new_n305_ = _165gat_41_ & ~new_n296_;
  assign new_n306_ = ~new_n300_ & ~new_n302_;
  assign new_n307_ = ~new_n304_ & new_n306_;
  assign new_n308_ = ~new_n305_ & new_n307_;
  assign new_n309_ = new_n278_ & ~new_n308_;
  assign new_n310_ = ~new_n278_ & new_n308_;
  assign new_n311_ = ~new_n309_ & ~new_n310_;
  assign new_n312_ = _219gat_50_ & new_n311_;
  assign new_n313_ = _210gat_49_ & _268gat_59_;
  assign new_n314_ = ~new_n312_ & ~new_n313_;
  assign new_n315_ = new_n280_ & new_n283_;
  assign _878gat_442_ = ~new_n314_ | ~new_n315_;
  assign _450gat_173_ = _89gat_21_ & ~new_n118_;
  assign new_n318_ = _237gat_52_ & new_n305_;
  assign new_n319_ = ~new_n297_ & ~new_n305_;
  assign new_n320_ = _228gat_51_ & new_n319_;
  assign new_n321_ = ~new_n318_ & ~new_n320_;
  assign new_n322_ = _165gat_41_ & new_n133_;
  assign new_n323_ = _246gat_53_ & ~new_n296_;
  assign new_n324_ = ~new_n322_ & ~new_n323_;
  assign new_n325_ = ~new_n221_ & ~new_n256_;
  assign new_n326_ = ~new_n290_ & new_n325_;
  assign new_n327_ = ~new_n303_ & ~new_n326_;
  assign new_n328_ = ~new_n301_ & new_n327_;
  assign new_n329_ = new_n319_ & ~new_n328_;
  assign new_n330_ = ~new_n319_ & new_n328_;
  assign new_n331_ = ~new_n329_ & ~new_n330_;
  assign new_n332_ = _219gat_50_ & new_n331_;
  assign new_n333_ = _210gat_49_ & _91gat_23_;
  assign new_n334_ = ~new_n332_ & ~new_n333_;
  assign new_n335_ = new_n321_ & new_n324_;
  assign _879gat_441_ = ~new_n334_ | ~new_n335_;
  assign new_n337_ = _74gat_14_ & _68gat_11_;
  assign new_n338_ = _59gat_10_ & new_n337_;
  assign _449gat_176_ = new_n131_ & new_n338_;
  assign new_n340_ = _237gat_52_ & new_n232_;
  assign new_n341_ = ~new_n232_ & ~new_n254_;
  assign new_n342_ = _228gat_51_ & new_n341_;
  assign new_n343_ = ~new_n340_ & ~new_n342_;
  assign new_n344_ = _183gat_44_ & new_n133_;
  assign new_n345_ = _246gat_53_ & ~new_n231_;
  assign new_n346_ = ~new_n344_ & ~new_n345_;
  assign new_n347_ = ~new_n253_ & new_n341_;
  assign new_n348_ = new_n253_ & ~new_n341_;
  assign new_n349_ = ~new_n347_ & ~new_n348_;
  assign new_n350_ = _219gat_50_ & new_n349_;
  assign new_n351_ = _210gat_49_ & _106gat_26_;
  assign new_n352_ = ~new_n350_ & ~new_n351_;
  assign new_n353_ = new_n343_ & new_n346_;
  assign _863gat_424_ = ~new_n352_ | ~new_n353_;
  assign _446gat_183_ = ~_390gat_131_ | ~new_n124_;
  assign new_n356_ = ~new_n277_ & ~new_n308_;
  assign _866gat_426_ = new_n275_ | new_n356_;
  assign new_n358_ = _237gat_52_ & new_n301_;
  assign new_n359_ = ~new_n290_ & ~new_n301_;
  assign new_n360_ = _228gat_51_ & new_n359_;
  assign new_n361_ = ~new_n358_ & ~new_n360_;
  assign new_n362_ = _171gat_42_ & new_n133_;
  assign new_n363_ = _246gat_53_ & ~new_n289_;
  assign new_n364_ = ~new_n362_ & ~new_n363_;
  assign new_n365_ = ~new_n219_ & ~new_n325_;
  assign new_n366_ = new_n359_ & ~new_n365_;
  assign new_n367_ = ~new_n359_ & new_n365_;
  assign new_n368_ = ~new_n366_ & ~new_n367_;
  assign new_n369_ = _219gat_50_ & new_n368_;
  assign new_n370_ = _210gat_49_ & _96gat_24_;
  assign new_n371_ = ~new_n369_ & ~new_n370_;
  assign new_n372_ = new_n361_ & new_n364_;
  assign _880gat_440_ = ~new_n371_ | ~new_n372_;
  assign _391gat_124_ = _85gat_17_ & _86gat_18_;
  assign new_n375_ = _68gat_11_ & _29gat_5_;
  assign _448gat_179_ = new_n131_ & new_n375_;
  assign new_n377_ = _195gat_46_ & new_n133_;
  assign new_n378_ = _237gat_52_ & new_n246_;
  assign new_n379_ = ~new_n237_ & ~new_n246_;
  assign new_n380_ = _228gat_51_ & new_n379_;
  assign new_n381_ = ~new_n378_ & ~new_n380_;
  assign new_n382_ = _246gat_53_ & ~new_n236_;
  assign new_n383_ = _260gat_56_ & _255gat_54_;
  assign new_n384_ = ~new_n382_ & ~new_n383_;
  assign new_n385_ = _261gat_57_ & ~new_n163_;
  assign new_n386_ = ~new_n161_ & ~new_n385_;
  assign new_n387_ = new_n379_ & ~new_n386_;
  assign new_n388_ = ~new_n379_ & new_n386_;
  assign new_n389_ = ~new_n387_ & ~new_n388_;
  assign new_n390_ = _219gat_50_ & new_n389_;
  assign new_n391_ = _210gat_49_ & _116gat_28_;
  assign new_n392_ = ~new_n390_ & ~new_n391_;
  assign new_n393_ = ~new_n377_ & new_n381_;
  assign new_n394_ = new_n384_ & new_n393_;
  assign _865gat_422_ = ~new_n392_ | ~new_n394_;
  assign new_n396_ = _189gat_45_ & new_n133_;
  assign new_n397_ = _237gat_52_ & new_n250_;
  assign new_n398_ = ~new_n242_ & ~new_n250_;
  assign new_n399_ = _228gat_51_ & new_n398_;
  assign new_n400_ = ~new_n397_ & ~new_n399_;
  assign new_n401_ = _246gat_53_ & ~new_n241_;
  assign new_n402_ = _259gat_55_ & _255gat_54_;
  assign new_n403_ = ~new_n401_ & ~new_n402_;
  assign new_n404_ = ~new_n237_ & new_n385_;
  assign new_n405_ = ~new_n248_ & ~new_n404_;
  assign new_n406_ = ~new_n246_ & new_n405_;
  assign new_n407_ = new_n398_ & ~new_n406_;
  assign new_n408_ = ~new_n398_ & new_n406_;
  assign new_n409_ = ~new_n407_ & ~new_n408_;
  assign new_n410_ = _219gat_50_ & new_n409_;
  assign new_n411_ = _210gat_49_ & _111gat_27_;
  assign new_n412_ = ~new_n410_ & ~new_n411_;
  assign new_n413_ = ~new_n396_ & new_n400_;
  assign new_n414_ = new_n403_ & new_n413_;
  assign _864gat_423_ = ~new_n412_ | ~new_n414_;
endmodule

