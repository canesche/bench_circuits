module top ( 
    pv96_30_, pv96_31_, pv96_10_, pv96_21_, pv138_4_, pv96_11_, pv96_20_,
    pv138_3_, pv138_2_, pv131_18_, pv138_0_, pv131_19_, pv32_7_, pv32_18_,
    pv32_29_, pv64_0_, pv96_9_, pv131_3_, pv131_29_, pv32_6_, pv32_19_,
    pv32_28_, pv64_1_, pv96_8_, pv131_2_, pv131_28_, pv32_5_, pv131_1_,
    pv32_4_, pv131_0_, pv32_3_, pv64_4_, pv96_5_, pv32_2_, pv64_5_,
    pv96_4_, pv32_1_, pv64_2_, pv96_7_, pv32_0_, pv64_3_, pv96_6_,
    pv32_10_, pv32_21_, pv64_8_, pv64_17_, pv64_28_, pv96_1_, pv97_0_,
    pv131_21_, pv32_11_, pv32_20_, pv64_9_, pv64_18_, pv64_27_, pv96_0_,
    pv131_20_, pv32_12_, pv32_23_, pv32_30_, pv64_6_, pv64_15_, pv64_26_,
    pv96_3_, pv99_0_, pv131_9_, pv131_23_, pv134_0_, pv32_13_, pv32_22_,
    pv32_31_, pv64_7_, pv64_16_, pv64_25_, pv96_2_, pv98_0_, pv131_8_,
    pv131_22_, pv32_14_, pv32_25_, pv131_7_, pv131_25_, pv131_30_,
    pv133_1_, pv32_15_, pv32_24_, pv131_6_, pv131_24_, pv131_31_, pv133_0_,
    pv32_9_, pv32_16_, pv32_27_, pv64_19_, pv131_5_, pv131_27_, pv32_8_,
    pv32_17_, pv32_26_, pv64_29_, pv131_4_, pv131_26_, pv64_20_, pv64_31_,
    pv96_16_, pv96_27_, pv131_16_, pv64_10_, pv96_17_, pv96_26_, pv131_17_,
    pv96_18_, pv96_29_, pv131_14_, pv96_19_, pv96_28_, pv131_15_, pv64_13_,
    pv64_24_, pv96_12_, pv96_23_, pv131_12_, pv64_14_, pv64_23_, pv96_13_,
    pv96_22_, pv131_13_, pv64_11_, pv64_22_, pv96_14_, pv96_25_, pv131_10_,
    pv64_12_, pv64_21_, pv64_30_, pv96_15_, pv96_24_, pv131_11_,
    pv198_17_, pv205_3_, pv198_16_, pv205_4_, pv198_19_, pv205_5_,
    pv198_18_, pv205_6_, pv198_8_, pv198_13_, pv198_7_, pv198_12_,
    pv205_0_, pv198_15_, pv205_1_, pv198_9_, pv198_14_, pv205_2_, pv166_7_,
    pv166_10_, pv166_23_, pv198_4_, pv198_22_, pv166_8_, pv166_24_,
    pv198_3_, pv198_23_, pv166_5_, pv166_21_, pv198_6_, pv198_24_,
    pv166_6_, pv166_22_, pv198_5_, pv198_25_, pv166_14_, pv198_0_,
    pv198_26_, pv166_13_, pv166_20_, pv198_27_, pv166_9_, pv166_12_,
    pv198_2_, pv198_28_, pv166_11_, pv198_1_, pv198_29_, pv166_18_,
    pv166_0_, pv166_17_, pv166_16_, pv166_15_, pv166_3_, pv166_27_,
    pv198_31_, pv166_4_, pv198_30_, pv166_1_, pv166_25_, pv198_20_,
    pv166_2_, pv166_19_, pv166_26_, pv198_21_, pv198_11_, pv198_10_  );
  input  pv96_30_, pv96_31_, pv96_10_, pv96_21_, pv138_4_, pv96_11_,
    pv96_20_, pv138_3_, pv138_2_, pv131_18_, pv138_0_, pv131_19_, pv32_7_,
    pv32_18_, pv32_29_, pv64_0_, pv96_9_, pv131_3_, pv131_29_, pv32_6_,
    pv32_19_, pv32_28_, pv64_1_, pv96_8_, pv131_2_, pv131_28_, pv32_5_,
    pv131_1_, pv32_4_, pv131_0_, pv32_3_, pv64_4_, pv96_5_, pv32_2_,
    pv64_5_, pv96_4_, pv32_1_, pv64_2_, pv96_7_, pv32_0_, pv64_3_, pv96_6_,
    pv32_10_, pv32_21_, pv64_8_, pv64_17_, pv64_28_, pv96_1_, pv97_0_,
    pv131_21_, pv32_11_, pv32_20_, pv64_9_, pv64_18_, pv64_27_, pv96_0_,
    pv131_20_, pv32_12_, pv32_23_, pv32_30_, pv64_6_, pv64_15_, pv64_26_,
    pv96_3_, pv99_0_, pv131_9_, pv131_23_, pv134_0_, pv32_13_, pv32_22_,
    pv32_31_, pv64_7_, pv64_16_, pv64_25_, pv96_2_, pv98_0_, pv131_8_,
    pv131_22_, pv32_14_, pv32_25_, pv131_7_, pv131_25_, pv131_30_,
    pv133_1_, pv32_15_, pv32_24_, pv131_6_, pv131_24_, pv131_31_, pv133_0_,
    pv32_9_, pv32_16_, pv32_27_, pv64_19_, pv131_5_, pv131_27_, pv32_8_,
    pv32_17_, pv32_26_, pv64_29_, pv131_4_, pv131_26_, pv64_20_, pv64_31_,
    pv96_16_, pv96_27_, pv131_16_, pv64_10_, pv96_17_, pv96_26_, pv131_17_,
    pv96_18_, pv96_29_, pv131_14_, pv96_19_, pv96_28_, pv131_15_, pv64_13_,
    pv64_24_, pv96_12_, pv96_23_, pv131_12_, pv64_14_, pv64_23_, pv96_13_,
    pv96_22_, pv131_13_, pv64_11_, pv64_22_, pv96_14_, pv96_25_, pv131_10_,
    pv64_12_, pv64_21_, pv64_30_, pv96_15_, pv96_24_, pv131_11_;
  output pv198_17_, pv205_3_, pv198_16_, pv205_4_, pv198_19_, pv205_5_,
    pv198_18_, pv205_6_, pv198_8_, pv198_13_, pv198_7_, pv198_12_,
    pv205_0_, pv198_15_, pv205_1_, pv198_9_, pv198_14_, pv205_2_, pv166_7_,
    pv166_10_, pv166_23_, pv198_4_, pv198_22_, pv166_8_, pv166_24_,
    pv198_3_, pv198_23_, pv166_5_, pv166_21_, pv198_6_, pv198_24_,
    pv166_6_, pv166_22_, pv198_5_, pv198_25_, pv166_14_, pv198_0_,
    pv198_26_, pv166_13_, pv166_20_, pv198_27_, pv166_9_, pv166_12_,
    pv198_2_, pv198_28_, pv166_11_, pv198_1_, pv198_29_, pv166_18_,
    pv166_0_, pv166_17_, pv166_16_, pv166_15_, pv166_3_, pv166_27_,
    pv198_31_, pv166_4_, pv198_30_, pv166_1_, pv166_25_, pv198_20_,
    pv166_2_, pv166_19_, pv166_26_, pv198_21_, pv198_11_, pv198_10_;
  wire new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n459_, new_n460_, new_n461_, new_n462_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n503_, new_n504_, new_n505_, new_n506_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n518_, new_n519_, new_n520_, new_n521_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_;
  assign new_n206_ = pv138_4_ & ~pv138_0_;
  assign new_n207_ = ~pv138_2_ & new_n206_;
  assign new_n208_ = pv96_13_ & new_n207_;
  assign new_n209_ = pv138_4_ & pv138_0_;
  assign new_n210_ = pv138_2_ & new_n209_;
  assign new_n211_ = ~pv131_13_ & new_n210_;
  assign new_n212_ = ~pv138_2_ & new_n209_;
  assign new_n213_ = pv131_13_ & new_n212_;
  assign new_n214_ = ~pv138_4_ & pv138_2_;
  assign new_n215_ = ~new_n208_ & ~new_n211_;
  assign new_n216_ = ~new_n213_ & ~new_n214_;
  assign pv198_17_ = ~new_n215_ | ~new_n216_;
  assign new_n218_ = pv138_3_ & ~pv138_0_;
  assign new_n219_ = ~pv138_2_ & new_n218_;
  assign new_n220_ = pv96_31_ & new_n219_;
  assign new_n221_ = pv138_3_ & pv138_0_;
  assign new_n222_ = pv138_2_ & new_n221_;
  assign new_n223_ = ~pv131_31_ & new_n222_;
  assign new_n224_ = ~pv138_2_ & new_n221_;
  assign new_n225_ = pv131_31_ & new_n224_;
  assign new_n226_ = ~pv138_3_ & pv138_2_;
  assign new_n227_ = ~new_n220_ & ~new_n223_;
  assign new_n228_ = ~new_n225_ & ~new_n226_;
  assign pv205_3_ = ~new_n227_ | ~new_n228_;
  assign new_n230_ = pv96_12_ & new_n207_;
  assign new_n231_ = ~pv131_12_ & new_n210_;
  assign new_n232_ = pv131_12_ & new_n212_;
  assign new_n233_ = ~new_n230_ & ~new_n231_;
  assign new_n234_ = ~new_n214_ & ~new_n232_;
  assign pv198_16_ = ~new_n233_ | ~new_n234_;
  assign new_n236_ = pv97_0_ & new_n219_;
  assign new_n237_ = ~pv133_0_ & new_n222_;
  assign new_n238_ = pv133_0_ & new_n224_;
  assign new_n239_ = ~new_n236_ & ~new_n237_;
  assign new_n240_ = ~new_n226_ & ~new_n238_;
  assign pv205_4_ = ~new_n239_ | ~new_n240_;
  assign new_n242_ = pv96_15_ & new_n207_;
  assign new_n243_ = ~pv131_15_ & new_n210_;
  assign new_n244_ = pv131_15_ & new_n212_;
  assign new_n245_ = ~new_n242_ & ~new_n243_;
  assign new_n246_ = ~new_n214_ & ~new_n244_;
  assign pv198_19_ = ~new_n245_ | ~new_n246_;
  assign new_n248_ = pv98_0_ & new_n219_;
  assign new_n249_ = ~pv133_1_ & new_n222_;
  assign new_n250_ = pv133_1_ & new_n224_;
  assign new_n251_ = ~new_n248_ & ~new_n249_;
  assign new_n252_ = ~new_n226_ & ~new_n250_;
  assign pv205_5_ = ~new_n251_ | ~new_n252_;
  assign new_n254_ = pv96_14_ & new_n207_;
  assign new_n255_ = ~pv131_14_ & new_n210_;
  assign new_n256_ = pv131_14_ & new_n212_;
  assign new_n257_ = ~new_n254_ & ~new_n255_;
  assign new_n258_ = ~new_n214_ & ~new_n256_;
  assign pv198_18_ = ~new_n257_ | ~new_n258_;
  assign new_n260_ = pv134_0_ & new_n224_;
  assign new_n261_ = pv99_0_ & new_n219_;
  assign new_n262_ = pv134_0_ & new_n222_;
  assign new_n263_ = ~new_n260_ & ~new_n261_;
  assign pv205_6_ = new_n262_ | ~new_n263_;
  assign new_n265_ = pv96_4_ & new_n207_;
  assign new_n266_ = ~pv131_4_ & new_n210_;
  assign new_n267_ = pv131_4_ & new_n212_;
  assign new_n268_ = ~new_n265_ & ~new_n266_;
  assign new_n269_ = ~new_n214_ & ~new_n267_;
  assign pv198_8_ = ~new_n268_ | ~new_n269_;
  assign new_n271_ = pv96_9_ & new_n207_;
  assign new_n272_ = ~pv131_9_ & new_n210_;
  assign new_n273_ = pv131_9_ & new_n212_;
  assign new_n274_ = ~new_n271_ & ~new_n272_;
  assign new_n275_ = ~new_n214_ & ~new_n273_;
  assign pv198_13_ = ~new_n274_ | ~new_n275_;
  assign new_n277_ = pv96_3_ & new_n207_;
  assign new_n278_ = ~pv131_3_ & new_n210_;
  assign new_n279_ = pv131_3_ & new_n212_;
  assign new_n280_ = ~new_n277_ & ~new_n278_;
  assign new_n281_ = ~new_n214_ & ~new_n279_;
  assign pv198_7_ = ~new_n280_ | ~new_n281_;
  assign new_n283_ = pv96_8_ & new_n207_;
  assign new_n284_ = ~pv131_8_ & new_n210_;
  assign new_n285_ = pv131_8_ & new_n212_;
  assign new_n286_ = ~new_n283_ & ~new_n284_;
  assign new_n287_ = ~new_n214_ & ~new_n285_;
  assign pv198_12_ = ~new_n286_ | ~new_n287_;
  assign new_n289_ = pv96_28_ & new_n219_;
  assign new_n290_ = ~pv131_28_ & new_n222_;
  assign new_n291_ = pv131_28_ & new_n224_;
  assign new_n292_ = ~new_n289_ & ~new_n290_;
  assign new_n293_ = ~new_n226_ & ~new_n291_;
  assign pv205_0_ = ~new_n292_ | ~new_n293_;
  assign new_n295_ = pv96_11_ & new_n207_;
  assign new_n296_ = ~pv131_11_ & new_n210_;
  assign new_n297_ = pv131_11_ & new_n212_;
  assign new_n298_ = ~new_n295_ & ~new_n296_;
  assign new_n299_ = ~new_n214_ & ~new_n297_;
  assign pv198_15_ = ~new_n298_ | ~new_n299_;
  assign new_n301_ = pv96_29_ & new_n219_;
  assign new_n302_ = ~pv131_29_ & new_n222_;
  assign new_n303_ = pv131_29_ & new_n224_;
  assign new_n304_ = ~new_n301_ & ~new_n302_;
  assign new_n305_ = ~new_n226_ & ~new_n303_;
  assign pv205_1_ = ~new_n304_ | ~new_n305_;
  assign new_n307_ = pv96_5_ & new_n207_;
  assign new_n308_ = ~pv131_5_ & new_n210_;
  assign new_n309_ = pv131_5_ & new_n212_;
  assign new_n310_ = ~new_n307_ & ~new_n308_;
  assign new_n311_ = ~new_n214_ & ~new_n309_;
  assign pv198_9_ = ~new_n310_ | ~new_n311_;
  assign new_n313_ = pv96_10_ & new_n207_;
  assign new_n314_ = ~pv131_10_ & new_n210_;
  assign new_n315_ = pv131_10_ & new_n212_;
  assign new_n316_ = ~new_n313_ & ~new_n314_;
  assign new_n317_ = ~new_n214_ & ~new_n315_;
  assign pv198_14_ = ~new_n316_ | ~new_n317_;
  assign new_n319_ = pv96_30_ & new_n219_;
  assign new_n320_ = ~pv131_30_ & new_n222_;
  assign new_n321_ = pv131_30_ & new_n224_;
  assign new_n322_ = ~new_n319_ & ~new_n320_;
  assign new_n323_ = ~new_n226_ & ~new_n321_;
  assign pv205_2_ = ~new_n322_ | ~new_n323_;
  assign new_n325_ = ~pv138_2_ & pv138_0_;
  assign new_n326_ = pv64_7_ & new_n325_;
  assign new_n327_ = ~pv138_2_ & ~pv138_0_;
  assign new_n328_ = pv32_7_ & new_n327_;
  assign new_n329_ = pv138_2_ & pv138_0_;
  assign new_n330_ = ~pv64_7_ & new_n329_;
  assign new_n331_ = ~new_n326_ & ~new_n328_;
  assign pv166_7_ = new_n330_ | ~new_n331_;
  assign new_n333_ = pv64_10_ & new_n325_;
  assign new_n334_ = pv32_10_ & new_n327_;
  assign new_n335_ = ~pv64_10_ & new_n329_;
  assign new_n336_ = ~new_n333_ & ~new_n334_;
  assign pv166_10_ = new_n335_ | ~new_n336_;
  assign new_n338_ = pv64_23_ & new_n325_;
  assign new_n339_ = pv32_23_ & new_n327_;
  assign new_n340_ = ~pv64_23_ & new_n329_;
  assign new_n341_ = ~new_n338_ & ~new_n339_;
  assign pv166_23_ = new_n340_ | ~new_n341_;
  assign new_n343_ = pv96_0_ & new_n207_;
  assign new_n344_ = ~pv131_0_ & new_n210_;
  assign new_n345_ = pv131_0_ & new_n212_;
  assign new_n346_ = ~new_n343_ & ~new_n344_;
  assign new_n347_ = ~new_n214_ & ~new_n345_;
  assign pv198_4_ = ~new_n346_ | ~new_n347_;
  assign new_n349_ = pv96_18_ & new_n207_;
  assign new_n350_ = ~pv131_18_ & new_n210_;
  assign new_n351_ = pv131_18_ & new_n212_;
  assign new_n352_ = ~new_n349_ & ~new_n350_;
  assign new_n353_ = ~new_n214_ & ~new_n351_;
  assign pv198_22_ = ~new_n352_ | ~new_n353_;
  assign new_n355_ = pv64_8_ & new_n325_;
  assign new_n356_ = pv32_8_ & new_n327_;
  assign new_n357_ = ~pv64_8_ & new_n329_;
  assign new_n358_ = ~new_n355_ & ~new_n356_;
  assign pv166_8_ = new_n357_ | ~new_n358_;
  assign new_n360_ = pv64_24_ & new_n325_;
  assign new_n361_ = pv32_24_ & new_n327_;
  assign new_n362_ = ~pv64_24_ & new_n329_;
  assign new_n363_ = ~new_n360_ & ~new_n361_;
  assign pv166_24_ = new_n362_ | ~new_n363_;
  assign new_n365_ = pv32_31_ & new_n207_;
  assign new_n366_ = ~pv64_31_ & new_n210_;
  assign new_n367_ = pv64_31_ & new_n212_;
  assign new_n368_ = ~new_n365_ & ~new_n366_;
  assign new_n369_ = ~new_n214_ & ~new_n367_;
  assign pv198_3_ = ~new_n368_ | ~new_n369_;
  assign new_n371_ = pv96_19_ & new_n207_;
  assign new_n372_ = ~pv131_19_ & new_n210_;
  assign new_n373_ = pv131_19_ & new_n212_;
  assign new_n374_ = ~new_n371_ & ~new_n372_;
  assign new_n375_ = ~new_n214_ & ~new_n373_;
  assign pv198_23_ = ~new_n374_ | ~new_n375_;
  assign new_n377_ = pv64_5_ & new_n325_;
  assign new_n378_ = pv32_5_ & new_n327_;
  assign new_n379_ = ~pv64_5_ & new_n329_;
  assign new_n380_ = ~new_n377_ & ~new_n378_;
  assign pv166_5_ = new_n379_ | ~new_n380_;
  assign new_n382_ = pv64_21_ & new_n325_;
  assign new_n383_ = pv32_21_ & new_n327_;
  assign new_n384_ = ~pv64_21_ & new_n329_;
  assign new_n385_ = ~new_n382_ & ~new_n383_;
  assign pv166_21_ = new_n384_ | ~new_n385_;
  assign new_n387_ = pv96_2_ & new_n207_;
  assign new_n388_ = ~pv131_2_ & new_n210_;
  assign new_n389_ = pv131_2_ & new_n212_;
  assign new_n390_ = ~new_n387_ & ~new_n388_;
  assign new_n391_ = ~new_n214_ & ~new_n389_;
  assign pv198_6_ = ~new_n390_ | ~new_n391_;
  assign new_n393_ = pv96_20_ & new_n207_;
  assign new_n394_ = ~pv131_20_ & new_n210_;
  assign new_n395_ = pv131_20_ & new_n212_;
  assign new_n396_ = ~new_n393_ & ~new_n394_;
  assign new_n397_ = ~new_n214_ & ~new_n395_;
  assign pv198_24_ = ~new_n396_ | ~new_n397_;
  assign new_n399_ = pv64_6_ & new_n325_;
  assign new_n400_ = pv32_6_ & new_n327_;
  assign new_n401_ = ~pv64_6_ & new_n329_;
  assign new_n402_ = ~new_n399_ & ~new_n400_;
  assign pv166_6_ = new_n401_ | ~new_n402_;
  assign new_n404_ = pv64_22_ & new_n325_;
  assign new_n405_ = pv32_22_ & new_n327_;
  assign new_n406_ = ~pv64_22_ & new_n329_;
  assign new_n407_ = ~new_n404_ & ~new_n405_;
  assign pv166_22_ = new_n406_ | ~new_n407_;
  assign new_n409_ = pv96_1_ & new_n207_;
  assign new_n410_ = ~pv131_1_ & new_n210_;
  assign new_n411_ = pv131_1_ & new_n212_;
  assign new_n412_ = ~new_n409_ & ~new_n410_;
  assign new_n413_ = ~new_n214_ & ~new_n411_;
  assign pv198_5_ = ~new_n412_ | ~new_n413_;
  assign new_n415_ = pv96_21_ & new_n207_;
  assign new_n416_ = ~pv131_21_ & new_n210_;
  assign new_n417_ = pv131_21_ & new_n212_;
  assign new_n418_ = ~new_n415_ & ~new_n416_;
  assign new_n419_ = ~new_n214_ & ~new_n417_;
  assign pv198_25_ = ~new_n418_ | ~new_n419_;
  assign new_n421_ = pv64_14_ & new_n325_;
  assign new_n422_ = pv32_14_ & new_n327_;
  assign new_n423_ = ~pv64_14_ & new_n329_;
  assign new_n424_ = ~new_n421_ & ~new_n422_;
  assign pv166_14_ = new_n423_ | ~new_n424_;
  assign new_n426_ = pv32_28_ & new_n207_;
  assign new_n427_ = ~pv64_28_ & new_n210_;
  assign new_n428_ = pv64_28_ & new_n212_;
  assign new_n429_ = ~new_n426_ & ~new_n427_;
  assign new_n430_ = ~new_n214_ & ~new_n428_;
  assign pv198_0_ = ~new_n429_ | ~new_n430_;
  assign new_n432_ = pv96_22_ & new_n207_;
  assign new_n433_ = ~pv131_22_ & new_n210_;
  assign new_n434_ = pv131_22_ & new_n212_;
  assign new_n435_ = ~new_n432_ & ~new_n433_;
  assign new_n436_ = ~new_n214_ & ~new_n434_;
  assign pv198_26_ = ~new_n435_ | ~new_n436_;
  assign new_n438_ = pv64_13_ & new_n325_;
  assign new_n439_ = pv32_13_ & new_n327_;
  assign new_n440_ = ~pv64_13_ & new_n329_;
  assign new_n441_ = ~new_n438_ & ~new_n439_;
  assign pv166_13_ = new_n440_ | ~new_n441_;
  assign new_n443_ = pv64_20_ & new_n325_;
  assign new_n444_ = pv32_20_ & new_n327_;
  assign new_n445_ = ~pv64_20_ & new_n329_;
  assign new_n446_ = ~new_n443_ & ~new_n444_;
  assign pv166_20_ = new_n445_ | ~new_n446_;
  assign new_n448_ = pv96_23_ & new_n207_;
  assign new_n449_ = ~pv131_23_ & new_n210_;
  assign new_n450_ = pv131_23_ & new_n212_;
  assign new_n451_ = ~new_n448_ & ~new_n449_;
  assign new_n452_ = ~new_n214_ & ~new_n450_;
  assign pv198_27_ = ~new_n451_ | ~new_n452_;
  assign new_n454_ = pv64_9_ & new_n325_;
  assign new_n455_ = pv32_9_ & new_n327_;
  assign new_n456_ = ~pv64_9_ & new_n329_;
  assign new_n457_ = ~new_n454_ & ~new_n455_;
  assign pv166_9_ = new_n456_ | ~new_n457_;
  assign new_n459_ = pv64_12_ & new_n325_;
  assign new_n460_ = pv32_12_ & new_n327_;
  assign new_n461_ = ~pv64_12_ & new_n329_;
  assign new_n462_ = ~new_n459_ & ~new_n460_;
  assign pv166_12_ = new_n461_ | ~new_n462_;
  assign new_n464_ = pv32_30_ & new_n207_;
  assign new_n465_ = ~pv64_30_ & new_n210_;
  assign new_n466_ = pv64_30_ & new_n212_;
  assign new_n467_ = ~new_n464_ & ~new_n465_;
  assign new_n468_ = ~new_n214_ & ~new_n466_;
  assign pv198_2_ = ~new_n467_ | ~new_n468_;
  assign new_n470_ = pv96_24_ & new_n207_;
  assign new_n471_ = ~pv131_24_ & new_n210_;
  assign new_n472_ = pv131_24_ & new_n212_;
  assign new_n473_ = ~new_n470_ & ~new_n471_;
  assign new_n474_ = ~new_n214_ & ~new_n472_;
  assign pv198_28_ = ~new_n473_ | ~new_n474_;
  assign new_n476_ = pv64_11_ & new_n325_;
  assign new_n477_ = pv32_11_ & new_n327_;
  assign new_n478_ = ~pv64_11_ & new_n329_;
  assign new_n479_ = ~new_n476_ & ~new_n477_;
  assign pv166_11_ = new_n478_ | ~new_n479_;
  assign new_n481_ = pv32_29_ & new_n207_;
  assign new_n482_ = ~pv64_29_ & new_n210_;
  assign new_n483_ = pv64_29_ & new_n212_;
  assign new_n484_ = ~new_n481_ & ~new_n482_;
  assign new_n485_ = ~new_n214_ & ~new_n483_;
  assign pv198_1_ = ~new_n484_ | ~new_n485_;
  assign new_n487_ = pv96_25_ & new_n207_;
  assign new_n488_ = ~pv131_25_ & new_n210_;
  assign new_n489_ = pv131_25_ & new_n212_;
  assign new_n490_ = ~new_n487_ & ~new_n488_;
  assign new_n491_ = ~new_n214_ & ~new_n489_;
  assign pv198_29_ = ~new_n490_ | ~new_n491_;
  assign new_n493_ = pv64_18_ & new_n325_;
  assign new_n494_ = pv32_18_ & new_n327_;
  assign new_n495_ = ~pv64_18_ & new_n329_;
  assign new_n496_ = ~new_n493_ & ~new_n494_;
  assign pv166_18_ = new_n495_ | ~new_n496_;
  assign new_n498_ = pv64_0_ & new_n325_;
  assign new_n499_ = pv32_0_ & new_n327_;
  assign new_n500_ = ~pv64_0_ & new_n329_;
  assign new_n501_ = ~new_n498_ & ~new_n499_;
  assign pv166_0_ = new_n500_ | ~new_n501_;
  assign new_n503_ = pv64_17_ & new_n325_;
  assign new_n504_ = pv32_17_ & new_n327_;
  assign new_n505_ = ~pv64_17_ & new_n329_;
  assign new_n506_ = ~new_n503_ & ~new_n504_;
  assign pv166_17_ = new_n505_ | ~new_n506_;
  assign new_n508_ = pv64_16_ & new_n325_;
  assign new_n509_ = pv32_16_ & new_n327_;
  assign new_n510_ = ~pv64_16_ & new_n329_;
  assign new_n511_ = ~new_n508_ & ~new_n509_;
  assign pv166_16_ = new_n510_ | ~new_n511_;
  assign new_n513_ = pv64_15_ & new_n325_;
  assign new_n514_ = pv32_15_ & new_n327_;
  assign new_n515_ = ~pv64_15_ & new_n329_;
  assign new_n516_ = ~new_n513_ & ~new_n514_;
  assign pv166_15_ = new_n515_ | ~new_n516_;
  assign new_n518_ = pv64_3_ & new_n325_;
  assign new_n519_ = pv32_3_ & new_n327_;
  assign new_n520_ = ~pv64_3_ & new_n329_;
  assign new_n521_ = ~new_n518_ & ~new_n519_;
  assign pv166_3_ = new_n520_ | ~new_n521_;
  assign new_n523_ = pv64_27_ & new_n325_;
  assign new_n524_ = pv32_27_ & new_n327_;
  assign new_n525_ = ~pv64_27_ & new_n329_;
  assign new_n526_ = ~new_n523_ & ~new_n524_;
  assign pv166_27_ = new_n525_ | ~new_n526_;
  assign new_n528_ = pv96_27_ & new_n207_;
  assign new_n529_ = ~pv131_27_ & new_n210_;
  assign new_n530_ = pv131_27_ & new_n212_;
  assign new_n531_ = ~new_n528_ & ~new_n529_;
  assign new_n532_ = ~new_n214_ & ~new_n530_;
  assign pv198_31_ = ~new_n531_ | ~new_n532_;
  assign new_n534_ = pv64_4_ & new_n325_;
  assign new_n535_ = pv32_4_ & new_n327_;
  assign new_n536_ = ~pv64_4_ & new_n329_;
  assign new_n537_ = ~new_n534_ & ~new_n535_;
  assign pv166_4_ = new_n536_ | ~new_n537_;
  assign new_n539_ = pv96_26_ & new_n207_;
  assign new_n540_ = ~pv131_26_ & new_n210_;
  assign new_n541_ = pv131_26_ & new_n212_;
  assign new_n542_ = ~new_n539_ & ~new_n540_;
  assign new_n543_ = ~new_n214_ & ~new_n541_;
  assign pv198_30_ = ~new_n542_ | ~new_n543_;
  assign new_n545_ = pv64_1_ & new_n325_;
  assign new_n546_ = pv32_1_ & new_n327_;
  assign new_n547_ = ~pv64_1_ & new_n329_;
  assign new_n548_ = ~new_n545_ & ~new_n546_;
  assign pv166_1_ = new_n547_ | ~new_n548_;
  assign new_n550_ = pv64_25_ & new_n325_;
  assign new_n551_ = pv32_25_ & new_n327_;
  assign new_n552_ = ~pv64_25_ & new_n329_;
  assign new_n553_ = ~new_n550_ & ~new_n551_;
  assign pv166_25_ = new_n552_ | ~new_n553_;
  assign new_n555_ = pv96_16_ & new_n207_;
  assign new_n556_ = ~pv131_16_ & new_n210_;
  assign new_n557_ = pv131_16_ & new_n212_;
  assign new_n558_ = ~new_n555_ & ~new_n556_;
  assign new_n559_ = ~new_n214_ & ~new_n557_;
  assign pv198_20_ = ~new_n558_ | ~new_n559_;
  assign new_n561_ = pv64_2_ & new_n325_;
  assign new_n562_ = pv32_2_ & new_n327_;
  assign new_n563_ = ~pv64_2_ & new_n329_;
  assign new_n564_ = ~new_n561_ & ~new_n562_;
  assign pv166_2_ = new_n563_ | ~new_n564_;
  assign new_n566_ = pv64_19_ & new_n325_;
  assign new_n567_ = pv32_19_ & new_n327_;
  assign new_n568_ = ~pv64_19_ & new_n329_;
  assign new_n569_ = ~new_n566_ & ~new_n567_;
  assign pv166_19_ = new_n568_ | ~new_n569_;
  assign new_n571_ = pv64_26_ & new_n325_;
  assign new_n572_ = pv32_26_ & new_n327_;
  assign new_n573_ = ~pv64_26_ & new_n329_;
  assign new_n574_ = ~new_n571_ & ~new_n572_;
  assign pv166_26_ = new_n573_ | ~new_n574_;
  assign new_n576_ = pv96_17_ & new_n207_;
  assign new_n577_ = ~pv131_17_ & new_n210_;
  assign new_n578_ = pv131_17_ & new_n212_;
  assign new_n579_ = ~new_n576_ & ~new_n577_;
  assign new_n580_ = ~new_n214_ & ~new_n578_;
  assign pv198_21_ = ~new_n579_ | ~new_n580_;
  assign new_n582_ = pv96_7_ & new_n207_;
  assign new_n583_ = ~pv131_7_ & new_n210_;
  assign new_n584_ = pv131_7_ & new_n212_;
  assign new_n585_ = ~new_n582_ & ~new_n583_;
  assign new_n586_ = ~new_n214_ & ~new_n584_;
  assign pv198_11_ = ~new_n585_ | ~new_n586_;
  assign new_n588_ = pv96_6_ & new_n207_;
  assign new_n589_ = ~pv131_6_ & new_n210_;
  assign new_n590_ = pv131_6_ & new_n212_;
  assign new_n591_ = ~new_n588_ & ~new_n589_;
  assign new_n592_ = ~new_n214_ & ~new_n590_;
  assign pv198_10_ = ~new_n591_ | ~new_n592_;
endmodule

