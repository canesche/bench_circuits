module top ( 
    _8, _7, _6, _5, _4, _3, _2, _1,
    _47, _48, _49, _44, _45, _46, _50, _51  );
  input  _8, _7, _6, _5, _4, _3, _2, _1;
  output _47, _48, _49, _44, _45, _46, _50, _51;
  wire new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_,
    new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_,
    new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_,
    new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_,
    new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_,
    new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n66_, new_n67_,
    new_n68_, new_n69_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_,
    new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_;
  assign new_n17_ = ~_7 & ~_5;
  assign new_n18_ = _6 & new_n17_;
  assign new_n19_ = ~_4 & new_n18_;
  assign new_n20_ = _8 & _6;
  assign new_n21_ = _7 & new_n20_;
  assign new_n22_ = _4 & new_n21_;
  assign new_n23_ = _7 & _5;
  assign new_n24_ = _6 & new_n23_;
  assign new_n25_ = _4 & new_n24_;
  assign new_n26_ = ~_6 & new_n23_;
  assign new_n27_ = ~_4 & new_n26_;
  assign new_n28_ = ~_7 & ~_6;
  assign new_n29_ = _4 & new_n28_;
  assign new_n30_ = ~_8 & _6;
  assign new_n31_ = ~_7 & new_n30_;
  assign new_n32_ = ~_4 & new_n31_;
  assign new_n33_ = ~_8 & ~_5;
  assign new_n34_ = _6 & new_n33_;
  assign new_n35_ = ~_4 & new_n34_;
  assign new_n36_ = ~_6 & new_n33_;
  assign new_n37_ = _4 & new_n36_;
  assign new_n38_ = _8 & ~_6;
  assign new_n39_ = _7 & new_n38_;
  assign new_n40_ = ~_4 & new_n39_;
  assign new_n41_ = _8 & _5;
  assign new_n42_ = ~_7 & new_n41_;
  assign new_n43_ = _4 & new_n42_;
  assign new_n44_ = ~new_n27_ & ~new_n29_;
  assign new_n45_ = ~new_n19_ & ~new_n22_;
  assign new_n46_ = ~new_n25_ & new_n45_;
  assign new_n47_ = new_n44_ & new_n46_;
  assign new_n48_ = ~new_n40_ & ~new_n43_;
  assign new_n49_ = ~new_n32_ & ~new_n35_;
  assign new_n50_ = ~new_n37_ & new_n49_;
  assign new_n51_ = new_n48_ & new_n50_;
  assign _47 = ~new_n47_ | ~new_n51_;
  assign new_n53_ = ~_8 & ~_7;
  assign new_n54_ = _5 & new_n53_;
  assign new_n55_ = ~_7 & new_n20_;
  assign new_n56_ = ~_5 & new_n55_;
  assign new_n57_ = _8 & _7;
  assign new_n58_ = _5 & new_n57_;
  assign new_n59_ = ~_8 & _7;
  assign new_n60_ = ~_5 & new_n59_;
  assign new_n61_ = _5 & new_n28_;
  assign new_n62_ = ~new_n60_ & ~new_n61_;
  assign new_n63_ = ~new_n54_ & ~new_n56_;
  assign new_n64_ = ~new_n58_ & new_n63_;
  assign _48 = ~new_n62_ | ~new_n64_;
  assign new_n66_ = _8 & ~_7;
  assign new_n67_ = ~_6 & new_n66_;
  assign new_n68_ = _7 & _6;
  assign new_n69_ = ~new_n30_ & ~new_n67_;
  assign _49 = new_n68_ | ~new_n69_;
  assign new_n71_ = ~_4 & ~_2;
  assign new_n72_ = ~_3 & new_n71_;
  assign new_n73_ = _1 & new_n72_;
  assign new_n74_ = _5 & _2;
  assign new_n75_ = _3 & new_n74_;
  assign new_n76_ = _1 & new_n75_;
  assign new_n77_ = _4 & _2;
  assign new_n78_ = ~_3 & new_n77_;
  assign new_n79_ = ~_1 & new_n78_;
  assign new_n80_ = _3 & new_n71_;
  assign new_n81_ = ~_1 & new_n80_;
  assign new_n82_ = _3 & new_n77_;
  assign new_n83_ = _1 & new_n82_;
  assign new_n84_ = _3 & new_n33_;
  assign new_n85_ = ~_4 & new_n84_;
  assign new_n86_ = ~_1 & new_n85_;
  assign new_n87_ = ~_3 & new_n53_;
  assign new_n88_ = ~_4 & new_n87_;
  assign new_n89_ = _1 & new_n88_;
  assign new_n90_ = _6 & _5;
  assign new_n91_ = _2 & new_n90_;
  assign new_n92_ = ~_3 & new_n91_;
  assign new_n93_ = ~_1 & new_n92_;
  assign new_n94_ = _7 & new_n93_;
  assign new_n95_ = ~_6 & ~_5;
  assign new_n96_ = ~_2 & new_n95_;
  assign new_n97_ = _3 & new_n96_;
  assign new_n98_ = ~_1 & new_n97_;
  assign new_n99_ = ~_7 & new_n98_;
  assign new_n100_ = ~_3 & new_n23_;
  assign new_n101_ = _4 & new_n100_;
  assign new_n102_ = ~_1 & new_n101_;
  assign new_n103_ = ~_8 & new_n98_;
  assign new_n104_ = _3 & new_n17_;
  assign new_n105_ = ~_4 & new_n104_;
  assign new_n106_ = ~_1 & new_n105_;
  assign new_n107_ = ~_2 & new_n28_;
  assign new_n108_ = ~_3 & new_n107_;
  assign new_n109_ = _1 & new_n108_;
  assign new_n110_ = _3 & new_n57_;
  assign new_n111_ = _4 & new_n110_;
  assign new_n112_ = _1 & new_n111_;
  assign new_n113_ = _2 & new_n68_;
  assign new_n114_ = _3 & new_n113_;
  assign new_n115_ = _1 & new_n114_;
  assign new_n116_ = _8 & new_n115_;
  assign new_n117_ = ~_3 & new_n90_;
  assign new_n118_ = _4 & new_n117_;
  assign new_n119_ = ~_1 & new_n118_;
  assign new_n120_ = _8 & new_n93_;
  assign new_n121_ = _3 & new_n95_;
  assign new_n122_ = ~_4 & new_n121_;
  assign new_n123_ = ~_1 & new_n122_;
  assign new_n124_ = ~_6 & ~_3;
  assign new_n125_ = ~_4 & new_n124_;
  assign new_n126_ = _1 & new_n125_;
  assign new_n127_ = ~_5 & ~_3;
  assign new_n128_ = ~_4 & new_n127_;
  assign new_n129_ = _1 & new_n128_;
  assign new_n130_ = _6 & _3;
  assign new_n131_ = _4 & new_n130_;
  assign new_n132_ = _1 & new_n131_;
  assign new_n133_ = _5 & _3;
  assign new_n134_ = _4 & new_n133_;
  assign new_n135_ = _1 & new_n134_;
  assign new_n136_ = ~_5 & ~_2;
  assign new_n137_ = ~_3 & new_n136_;
  assign new_n138_ = _1 & new_n137_;
  assign new_n139_ = ~new_n135_ & ~new_n138_;
  assign new_n140_ = ~new_n126_ & ~new_n129_;
  assign new_n141_ = ~new_n132_ & new_n140_;
  assign new_n142_ = new_n139_ & new_n141_;
  assign new_n143_ = ~new_n119_ & ~new_n120_;
  assign new_n144_ = ~new_n123_ & new_n143_;
  assign new_n145_ = ~new_n109_ & ~new_n112_;
  assign new_n146_ = ~new_n116_ & new_n145_;
  assign new_n147_ = new_n144_ & new_n146_;
  assign new_n148_ = new_n142_ & new_n147_;
  assign new_n149_ = ~new_n102_ & ~new_n103_;
  assign new_n150_ = ~new_n106_ & new_n149_;
  assign new_n151_ = ~new_n89_ & ~new_n94_;
  assign new_n152_ = ~new_n99_ & new_n151_;
  assign new_n153_ = new_n150_ & new_n152_;
  assign new_n154_ = ~new_n73_ & ~new_n76_;
  assign new_n155_ = ~new_n79_ & new_n154_;
  assign new_n156_ = ~new_n81_ & ~new_n83_;
  assign new_n157_ = ~new_n86_ & new_n156_;
  assign new_n158_ = new_n155_ & new_n157_;
  assign new_n159_ = new_n153_ & new_n158_;
  assign _44 = ~new_n148_ | ~new_n159_;
  assign new_n161_ = _2 & new_n128_;
  assign new_n162_ = _2 & new_n131_;
  assign new_n163_ = ~_4 & new_n133_;
  assign new_n164_ = ~_2 & new_n163_;
  assign new_n165_ = _4 & new_n127_;
  assign new_n166_ = ~_2 & new_n165_;
  assign new_n167_ = _2 & new_n134_;
  assign new_n168_ = _3 & new_n68_;
  assign new_n169_ = ~_4 & new_n168_;
  assign new_n170_ = ~_2 & new_n169_;
  assign new_n171_ = _8 & new_n170_;
  assign new_n172_ = _7 & ~_6;
  assign new_n173_ = _3 & new_n172_;
  assign new_n174_ = ~_5 & new_n173_;
  assign new_n175_ = _2 & new_n174_;
  assign new_n176_ = _8 & new_n175_;
  assign new_n177_ = ~_5 & new_n29_;
  assign new_n178_ = ~_2 & new_n177_;
  assign new_n179_ = ~_4 & new_n20_;
  assign new_n180_ = _5 & new_n179_;
  assign new_n181_ = ~_2 & new_n180_;
  assign new_n182_ = ~_8 & ~_6;
  assign new_n183_ = _4 & new_n182_;
  assign new_n184_ = ~_5 & new_n183_;
  assign new_n185_ = ~_2 & new_n184_;
  assign new_n186_ = _2 & new_n88_;
  assign new_n187_ = ~_4 & new_n68_;
  assign new_n188_ = _5 & new_n187_;
  assign new_n189_ = ~_2 & new_n188_;
  assign new_n190_ = ~_3 & new_n28_;
  assign new_n191_ = _4 & new_n190_;
  assign new_n192_ = ~_2 & new_n191_;
  assign new_n193_ = ~_8 & ~_4;
  assign new_n194_ = ~_5 & new_n193_;
  assign new_n195_ = _2 & new_n194_;
  assign new_n196_ = _7 & _4;
  assign new_n197_ = _5 & new_n196_;
  assign new_n198_ = _2 & new_n197_;
  assign new_n199_ = ~_7 & ~_4;
  assign new_n200_ = ~_5 & new_n199_;
  assign new_n201_ = _2 & new_n200_;
  assign new_n202_ = _6 & _4;
  assign new_n203_ = _5 & new_n202_;
  assign new_n204_ = _2 & new_n203_;
  assign new_n205_ = _2 & new_n125_;
  assign new_n206_ = ~new_n204_ & ~new_n205_;
  assign new_n207_ = ~new_n198_ & ~new_n201_;
  assign new_n208_ = new_n206_ & new_n207_;
  assign new_n209_ = ~new_n192_ & ~new_n195_;
  assign new_n210_ = ~new_n185_ & ~new_n186_;
  assign new_n211_ = ~new_n189_ & new_n210_;
  assign new_n212_ = new_n209_ & new_n211_;
  assign new_n213_ = new_n208_ & new_n212_;
  assign new_n214_ = ~new_n166_ & ~new_n167_;
  assign new_n215_ = ~new_n161_ & ~new_n162_;
  assign new_n216_ = ~new_n164_ & new_n215_;
  assign new_n217_ = new_n214_ & new_n216_;
  assign new_n218_ = ~new_n171_ & ~new_n176_;
  assign new_n219_ = ~new_n178_ & ~new_n181_;
  assign new_n220_ = new_n218_ & new_n219_;
  assign new_n221_ = new_n217_ & new_n220_;
  assign _45 = ~new_n213_ | ~new_n221_;
  assign new_n223_ = ~_6 & ~_4;
  assign new_n224_ = ~_5 & new_n223_;
  assign new_n225_ = _3 & new_n224_;
  assign new_n226_ = _3 & new_n197_;
  assign new_n227_ = ~_5 & new_n202_;
  assign new_n228_ = ~_3 & new_n227_;
  assign new_n229_ = _5 & new_n223_;
  assign new_n230_ = ~_3 & new_n229_;
  assign new_n231_ = _3 & new_n203_;
  assign new_n232_ = ~_4 & new_n66_;
  assign new_n233_ = _6 & new_n232_;
  assign new_n234_ = _3 & new_n233_;
  assign new_n235_ = ~_4 & new_n53_;
  assign new_n236_ = _5 & new_n235_;
  assign new_n237_ = ~_3 & new_n236_;
  assign new_n238_ = _4 & new_n57_;
  assign new_n239_ = ~_5 & new_n238_;
  assign new_n240_ = ~_3 & new_n239_;
  assign new_n241_ = ~_5 & new_n57_;
  assign new_n242_ = _6 & new_n241_;
  assign new_n243_ = ~_3 & new_n242_;
  assign new_n244_ = _3 & new_n36_;
  assign new_n245_ = ~_6 & new_n17_;
  assign new_n246_ = _3 & new_n245_;
  assign new_n247_ = _3 & new_n194_;
  assign new_n248_ = _3 & new_n24_;
  assign new_n249_ = ~_7 & _5;
  assign new_n250_ = ~_6 & new_n249_;
  assign new_n251_ = ~_3 & new_n250_;
  assign new_n252_ = ~new_n247_ & ~new_n248_;
  assign new_n253_ = ~new_n251_ & new_n252_;
  assign new_n254_ = ~new_n244_ & ~new_n246_;
  assign new_n255_ = ~new_n240_ & ~new_n243_;
  assign new_n256_ = new_n254_ & new_n255_;
  assign new_n257_ = new_n253_ & new_n256_;
  assign new_n258_ = ~new_n231_ & ~new_n234_;
  assign new_n259_ = ~new_n237_ & new_n258_;
  assign new_n260_ = ~new_n225_ & ~new_n226_;
  assign new_n261_ = ~new_n228_ & ~new_n230_;
  assign new_n262_ = new_n260_ & new_n261_;
  assign new_n263_ = new_n259_ & new_n262_;
  assign _46 = ~new_n257_ | ~new_n263_;
  assign _50 = new_n59_ | new_n66_;
  assign _51 = ~_8;
endmodule

