// Benchmark "testing" written by ABC on Thu Oct  8 22:16:29 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A105  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A105;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ , \new_[350]_ ,
    \new_[351]_ , \new_[352]_ , \new_[353]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[405]_ ,
    \new_[406]_ , \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ ,
    \new_[411]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[436]_ , \new_[437]_ , \new_[438]_ , \new_[439]_ , \new_[440]_ ,
    \new_[441]_ , \new_[442]_ , \new_[443]_ , \new_[444]_ , \new_[445]_ ,
    \new_[446]_ , \new_[447]_ , \new_[448]_ , \new_[449]_ , \new_[450]_ ,
    \new_[451]_ , \new_[452]_ , \new_[453]_ , \new_[454]_ , \new_[455]_ ,
    \new_[456]_ , \new_[457]_ , \new_[458]_ , \new_[459]_ , \new_[460]_ ,
    \new_[461]_ , \new_[462]_ , \new_[463]_ , \new_[464]_ , \new_[465]_ ,
    \new_[466]_ , \new_[467]_ , \new_[468]_ , \new_[469]_ , \new_[470]_ ,
    \new_[471]_ , \new_[472]_ , \new_[473]_ , \new_[474]_ , \new_[475]_ ,
    \new_[476]_ , \new_[477]_ , \new_[478]_ , \new_[479]_ , \new_[480]_ ,
    \new_[481]_ , \new_[482]_ , \new_[483]_ , \new_[484]_ , \new_[485]_ ,
    \new_[486]_ , \new_[487]_ , \new_[488]_ , \new_[489]_ , \new_[490]_ ,
    \new_[491]_ , \new_[492]_ , \new_[493]_ , \new_[494]_ , \new_[495]_ ,
    \new_[496]_ , \new_[497]_ , \new_[498]_ , \new_[499]_ , \new_[500]_ ,
    \new_[501]_ , \new_[502]_ , \new_[503]_ , \new_[504]_ , \new_[505]_ ,
    \new_[506]_ , \new_[507]_ , \new_[508]_ , \new_[509]_ , \new_[510]_ ,
    \new_[511]_ , \new_[512]_ , \new_[513]_ , \new_[514]_ , \new_[515]_ ,
    \new_[516]_ , \new_[517]_ , \new_[518]_ , \new_[519]_ , \new_[520]_ ,
    \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[525]_ ,
    \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ , \new_[530]_ ,
    \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ , \new_[535]_ ,
    \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ , \new_[540]_ ,
    \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ , \new_[545]_ ,
    \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ , \new_[550]_ ,
    \new_[551]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[566]_ , \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ ,
    \new_[571]_ , \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ ,
    \new_[576]_ , \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ ,
    \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[584]_ , \new_[585]_ ,
    \new_[586]_ , \new_[587]_ , \new_[588]_ , \new_[589]_ , \new_[590]_ ,
    \new_[591]_ , \new_[592]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[598]_ , \new_[599]_ , \new_[600]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ ,
    \new_[611]_ , \new_[612]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[616]_ , \new_[617]_ , \new_[618]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[626]_ , \new_[627]_ , \new_[628]_ , \new_[629]_ , \new_[630]_ ,
    \new_[631]_ , \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ ,
    \new_[636]_ , \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ ,
    \new_[641]_ , \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ ,
    \new_[646]_ , \new_[647]_ , \new_[648]_ , \new_[649]_ , \new_[650]_ ,
    \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[655]_ ,
    \new_[656]_ , \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ ,
    \new_[661]_ , \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ ,
    \new_[666]_ , \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ ,
    \new_[671]_ , \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ ,
    \new_[676]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ ,
    \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ ,
    \new_[686]_ , \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ ,
    \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ ,
    \new_[696]_ , \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ ,
    \new_[701]_ , \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ ,
    \new_[706]_ , \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ ,
    \new_[711]_ , \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ ,
    \new_[716]_ , \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ ,
    \new_[726]_ , \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ ,
    \new_[731]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[736]_ , \new_[737]_ , \new_[738]_ , \new_[739]_ , \new_[740]_ ,
    \new_[741]_ , \new_[742]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ ,
    \new_[746]_ , \new_[747]_ , \new_[748]_ , \new_[749]_ , \new_[750]_ ,
    \new_[751]_ , \new_[752]_ , \new_[753]_ , \new_[754]_ , \new_[755]_ ,
    \new_[756]_ , \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ ,
    \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ ,
    \new_[766]_ , \new_[767]_ , \new_[768]_ , \new_[769]_ , \new_[770]_ ,
    \new_[771]_ , \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ ,
    \new_[776]_ , \new_[777]_ , \new_[778]_ , \new_[779]_ , \new_[780]_ ,
    \new_[781]_ , \new_[782]_ , \new_[783]_ , \new_[784]_ , \new_[785]_ ,
    \new_[786]_ , \new_[787]_ , \new_[788]_ , \new_[789]_ , \new_[790]_ ,
    \new_[791]_ , \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ ,
    \new_[796]_ , \new_[797]_ , \new_[798]_ , \new_[799]_ , \new_[800]_ ,
    \new_[801]_ , \new_[802]_ , \new_[803]_ , \new_[804]_ , \new_[805]_ ,
    \new_[806]_ , \new_[807]_ , \new_[808]_ , \new_[809]_ , \new_[810]_ ,
    \new_[811]_ , \new_[812]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ ,
    \new_[816]_ , \new_[817]_ , \new_[818]_ , \new_[819]_ , \new_[820]_ ,
    \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[824]_ , \new_[825]_ ,
    \new_[826]_ , \new_[827]_ , \new_[828]_ , \new_[829]_ , \new_[830]_ ,
    \new_[831]_ , \new_[832]_ , \new_[833]_ , \new_[834]_ , \new_[835]_ ,
    \new_[836]_ , \new_[837]_ , \new_[838]_ , \new_[839]_ , \new_[840]_ ,
    \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[845]_ ,
    \new_[846]_ , \new_[847]_ , \new_[848]_ , \new_[849]_ , \new_[850]_ ,
    \new_[851]_ , \new_[852]_ , \new_[853]_ , \new_[854]_ , \new_[855]_ ,
    \new_[856]_ , \new_[857]_ , \new_[858]_ , \new_[859]_ , \new_[860]_ ,
    \new_[861]_ , \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[865]_ ,
    \new_[866]_ , \new_[867]_ , \new_[868]_ , \new_[869]_ , \new_[870]_ ,
    \new_[871]_ , \new_[872]_ , \new_[873]_ , \new_[874]_ , \new_[875]_ ,
    \new_[876]_ , \new_[877]_ , \new_[878]_ , \new_[879]_ , \new_[880]_ ,
    \new_[881]_ , \new_[882]_ , \new_[883]_ , \new_[884]_ , \new_[885]_ ,
    \new_[886]_ , \new_[887]_ , \new_[888]_ , \new_[889]_ , \new_[890]_ ,
    \new_[891]_ , \new_[892]_ , \new_[893]_ , \new_[894]_ , \new_[895]_ ,
    \new_[896]_ , \new_[897]_ , \new_[898]_ , \new_[899]_ , \new_[900]_ ,
    \new_[901]_ , \new_[902]_ , \new_[903]_ , \new_[904]_ , \new_[905]_ ,
    \new_[906]_ , \new_[907]_ , \new_[908]_ , \new_[909]_ , \new_[910]_ ,
    \new_[911]_ , \new_[912]_ , \new_[913]_ , \new_[914]_ , \new_[915]_ ,
    \new_[916]_ , \new_[917]_ , \new_[918]_ , \new_[919]_ , \new_[920]_ ,
    \new_[921]_ , \new_[922]_ , \new_[923]_ , \new_[924]_ , \new_[925]_ ,
    \new_[926]_ , \new_[927]_ , \new_[928]_ , \new_[929]_ , \new_[930]_ ,
    \new_[931]_ , \new_[932]_ , \new_[933]_ , \new_[934]_ , \new_[935]_ ,
    \new_[936]_ , \new_[937]_ , \new_[938]_ , \new_[939]_ , \new_[940]_ ,
    \new_[941]_ , \new_[942]_ , \new_[943]_ , \new_[944]_ , \new_[945]_ ,
    \new_[946]_ , \new_[947]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ ,
    \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[955]_ ,
    \new_[956]_ , \new_[957]_ , \new_[958]_ , \new_[959]_ , \new_[960]_ ,
    \new_[961]_ , \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ ,
    \new_[966]_ , \new_[967]_ , \new_[968]_ , \new_[969]_ , \new_[970]_ ,
    \new_[971]_ , \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[975]_ ,
    \new_[976]_ , \new_[977]_ , \new_[978]_ , \new_[979]_ , \new_[980]_ ,
    \new_[981]_ , \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ ,
    \new_[986]_ , \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ ,
    \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ ,
    \new_[996]_ , \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ ,
    \new_[1001]_ , \new_[1002]_ , \new_[1003]_ , \new_[1004]_ ,
    \new_[1005]_ , \new_[1006]_ , \new_[1007]_ , \new_[1008]_ ,
    \new_[1009]_ , \new_[1010]_ , \new_[1011]_ , \new_[1012]_ ,
    \new_[1013]_ , \new_[1014]_ , \new_[1015]_ , \new_[1016]_ ,
    \new_[1017]_ , \new_[1018]_ , \new_[1019]_ , \new_[1020]_ ,
    \new_[1021]_ , \new_[1022]_ , \new_[1023]_ , \new_[1024]_ ,
    \new_[1025]_ , \new_[1026]_ , \new_[1027]_ , \new_[1028]_ ,
    \new_[1029]_ , \new_[1030]_ , \new_[1031]_ , \new_[1032]_ ,
    \new_[1033]_ , \new_[1034]_ , \new_[1035]_ , \new_[1036]_ ,
    \new_[1037]_ , \new_[1038]_ , \new_[1039]_ , \new_[1040]_ ,
    \new_[1041]_ , \new_[1042]_ , \new_[1043]_ , \new_[1044]_ ,
    \new_[1045]_ , \new_[1046]_ , \new_[1047]_ , \new_[1048]_ ,
    \new_[1049]_ , \new_[1050]_ , \new_[1051]_ , \new_[1052]_ ,
    \new_[1053]_ , \new_[1054]_ , \new_[1055]_ , \new_[1056]_ ,
    \new_[1057]_ , \new_[1058]_ , \new_[1059]_ , \new_[1060]_ ,
    \new_[1061]_ , \new_[1062]_ , \new_[1063]_ , \new_[1064]_ ,
    \new_[1065]_ , \new_[1066]_ , \new_[1067]_ , \new_[1068]_ ,
    \new_[1069]_ , \new_[1070]_ , \new_[1071]_ , \new_[1072]_ ,
    \new_[1073]_ , \new_[1074]_ , \new_[1075]_ , \new_[1076]_ ,
    \new_[1077]_ , \new_[1078]_ , \new_[1079]_ , \new_[1080]_ ,
    \new_[1081]_ , \new_[1082]_ , \new_[1083]_ , \new_[1084]_ ,
    \new_[1085]_ , \new_[1086]_ , \new_[1087]_ , \new_[1088]_ ,
    \new_[1089]_ , \new_[1090]_ , \new_[1091]_ , \new_[1092]_ ,
    \new_[1093]_ , \new_[1094]_ , \new_[1095]_ , \new_[1096]_ ,
    \new_[1097]_ , \new_[1098]_ , \new_[1099]_ , \new_[1100]_ ,
    \new_[1101]_ , \new_[1102]_ , \new_[1103]_ , \new_[1104]_ ,
    \new_[1105]_ , \new_[1106]_ , \new_[1107]_ , \new_[1108]_ ,
    \new_[1109]_ , \new_[1110]_ , \new_[1111]_ , \new_[1112]_ ,
    \new_[1113]_ , \new_[1114]_ , \new_[1115]_ , \new_[1116]_ ,
    \new_[1117]_ , \new_[1118]_ , \new_[1119]_ , \new_[1120]_ ,
    \new_[1121]_ , \new_[1122]_ , \new_[1123]_ , \new_[1124]_ ,
    \new_[1125]_ , \new_[1126]_ , \new_[1127]_ , \new_[1128]_ ,
    \new_[1129]_ , \new_[1130]_ , \new_[1131]_ , \new_[1132]_ ,
    \new_[1133]_ , \new_[1134]_ , \new_[1135]_ , \new_[1136]_ ,
    \new_[1137]_ , \new_[1138]_ , \new_[1139]_ , \new_[1140]_ ,
    \new_[1141]_ , \new_[1142]_ , \new_[1143]_ , \new_[1144]_ ,
    \new_[1145]_ , \new_[1146]_ , \new_[1147]_ , \new_[1148]_ ,
    \new_[1149]_ , \new_[1150]_ , \new_[1151]_ , \new_[1152]_ ,
    \new_[1153]_ , \new_[1154]_ , \new_[1155]_ , \new_[1156]_ ,
    \new_[1157]_ , \new_[1158]_ , \new_[1159]_ , \new_[1160]_ ,
    \new_[1161]_ , \new_[1162]_ , \new_[1163]_ , \new_[1164]_ ,
    \new_[1165]_ , \new_[1166]_ , \new_[1167]_ , \new_[1168]_ ,
    \new_[1169]_ , \new_[1170]_ , \new_[1171]_ , \new_[1172]_ ,
    \new_[1173]_ , \new_[1174]_ , \new_[1175]_ , \new_[1176]_ ,
    \new_[1177]_ , \new_[1178]_ , \new_[1179]_ , \new_[1180]_ ,
    \new_[1181]_ , \new_[1182]_ , \new_[1183]_ , \new_[1184]_ ,
    \new_[1185]_ , \new_[1186]_ , \new_[1187]_ , \new_[1188]_ ,
    \new_[1189]_ , \new_[1190]_ , \new_[1191]_ , \new_[1192]_ ,
    \new_[1193]_ , \new_[1194]_ , \new_[1195]_ , \new_[1196]_ ,
    \new_[1197]_ , \new_[1198]_ , \new_[1199]_ , \new_[1200]_ ,
    \new_[1201]_ , \new_[1202]_ , \new_[1203]_ , \new_[1204]_ ,
    \new_[1205]_ , \new_[1206]_ , \new_[1207]_ , \new_[1208]_ ,
    \new_[1209]_ , \new_[1210]_ , \new_[1211]_ , \new_[1212]_ ,
    \new_[1213]_ , \new_[1214]_ , \new_[1215]_ , \new_[1216]_ ,
    \new_[1217]_ , \new_[1218]_ , \new_[1219]_ , \new_[1220]_ ,
    \new_[1221]_ , \new_[1222]_ , \new_[1223]_ , \new_[1224]_ ,
    \new_[1225]_ , \new_[1226]_ , \new_[1227]_ , \new_[1228]_ ,
    \new_[1229]_ , \new_[1230]_ , \new_[1231]_ , \new_[1232]_ ,
    \new_[1233]_ , \new_[1234]_ , \new_[1235]_ , \new_[1236]_ ,
    \new_[1237]_ , \new_[1238]_ , \new_[1239]_ , \new_[1240]_ ,
    \new_[1241]_ , \new_[1242]_ , \new_[1243]_ , \new_[1244]_ ,
    \new_[1245]_ , \new_[1246]_ , \new_[1247]_ , \new_[1248]_ ,
    \new_[1249]_ , \new_[1250]_ , \new_[1251]_ , \new_[1252]_ ,
    \new_[1253]_ , \new_[1254]_ , \new_[1255]_ , \new_[1256]_ ,
    \new_[1257]_ , \new_[1258]_ , \new_[1259]_ , \new_[1260]_ ,
    \new_[1261]_ , \new_[1262]_ , \new_[1263]_ , \new_[1264]_ ,
    \new_[1265]_ , \new_[1266]_ , \new_[1267]_ , \new_[1268]_ ,
    \new_[1269]_ , \new_[1270]_ , \new_[1271]_ , \new_[1272]_ ,
    \new_[1273]_ , \new_[1274]_ , \new_[1275]_ , \new_[1276]_ ,
    \new_[1277]_ , \new_[1278]_ , \new_[1279]_ , \new_[1280]_ ,
    \new_[1281]_ , \new_[1282]_ , \new_[1283]_ , \new_[1284]_ ,
    \new_[1285]_ , \new_[1286]_ , \new_[1287]_ , \new_[1288]_ ,
    \new_[1289]_ , \new_[1290]_ , \new_[1291]_ , \new_[1292]_ ,
    \new_[1293]_ , \new_[1294]_ , \new_[1295]_ , \new_[1296]_ ,
    \new_[1297]_ , \new_[1298]_ , \new_[1299]_ , \new_[1300]_ ,
    \new_[1301]_ , \new_[1302]_ , \new_[1303]_ , \new_[1304]_ ,
    \new_[1305]_ , \new_[1306]_ , \new_[1307]_ , \new_[1308]_ ,
    \new_[1309]_ , \new_[1310]_ , \new_[1311]_ , \new_[1312]_ ,
    \new_[1313]_ , \new_[1314]_ , \new_[1315]_ , \new_[1316]_ ,
    \new_[1317]_ , \new_[1318]_ , \new_[1319]_ , \new_[1320]_ ,
    \new_[1321]_ , \new_[1322]_ , \new_[1323]_ , \new_[1324]_ ,
    \new_[1325]_ , \new_[1326]_ , \new_[1327]_ , \new_[1328]_ ,
    \new_[1329]_ , \new_[1330]_ , \new_[1331]_ , \new_[1332]_ ,
    \new_[1333]_ , \new_[1334]_ , \new_[1335]_ , \new_[1336]_ ,
    \new_[1337]_ , \new_[1338]_ , \new_[1339]_ , \new_[1340]_ ,
    \new_[1341]_ , \new_[1342]_ , \new_[1343]_ , \new_[1344]_ ,
    \new_[1345]_ , \new_[1346]_ , \new_[1347]_ , \new_[1348]_ ,
    \new_[1349]_ , \new_[1350]_ , \new_[1351]_ , \new_[1352]_ ,
    \new_[1353]_ , \new_[1354]_ , \new_[1355]_ , \new_[1356]_ ,
    \new_[1357]_ , \new_[1358]_ , \new_[1359]_ , \new_[1360]_ ,
    \new_[1361]_ , \new_[1362]_ , \new_[1363]_ , \new_[1364]_ ,
    \new_[1365]_ , \new_[1366]_ , \new_[1367]_ , \new_[1368]_ ,
    \new_[1369]_ , \new_[1370]_ , \new_[1371]_ , \new_[1372]_ ,
    \new_[1373]_ , \new_[1374]_ , \new_[1375]_ , \new_[1376]_ ,
    \new_[1377]_ , \new_[1378]_ , \new_[1379]_ , \new_[1380]_ ,
    \new_[1381]_ , \new_[1382]_ , \new_[1383]_ , \new_[1384]_ ,
    \new_[1385]_ , \new_[1386]_ , \new_[1387]_ , \new_[1388]_ ,
    \new_[1389]_ , \new_[1390]_ , \new_[1391]_ , \new_[1392]_ ,
    \new_[1393]_ , \new_[1394]_ , \new_[1395]_ , \new_[1396]_ ,
    \new_[1397]_ , \new_[1398]_ , \new_[1399]_ , \new_[1400]_ ,
    \new_[1401]_ , \new_[1402]_ , \new_[1403]_ , \new_[1404]_ ,
    \new_[1405]_ , \new_[1406]_ , \new_[1407]_ , \new_[1408]_ ,
    \new_[1409]_ , \new_[1410]_ , \new_[1411]_ , \new_[1412]_ ,
    \new_[1413]_ , \new_[1414]_ , \new_[1415]_ , \new_[1416]_ ,
    \new_[1417]_ , \new_[1418]_ , \new_[1419]_ , \new_[1420]_ ,
    \new_[1421]_ , \new_[1422]_ , \new_[1423]_ , \new_[1424]_ ,
    \new_[1425]_ , \new_[1426]_ , \new_[1427]_ , \new_[1428]_ ,
    \new_[1429]_ , \new_[1430]_ , \new_[1431]_ , \new_[1432]_ ,
    \new_[1433]_ , \new_[1434]_ , \new_[1435]_ , \new_[1436]_ ,
    \new_[1437]_ , \new_[1438]_ , \new_[1439]_ , \new_[1440]_ ,
    \new_[1441]_ , \new_[1442]_ , \new_[1443]_ , \new_[1444]_ ,
    \new_[1445]_ , \new_[1446]_ , \new_[1447]_ , \new_[1448]_ ,
    \new_[1449]_ , \new_[1450]_ , \new_[1451]_ , \new_[1452]_ ,
    \new_[1453]_ , \new_[1454]_ , \new_[1455]_ , \new_[1456]_ ,
    \new_[1457]_ , \new_[1458]_ , \new_[1459]_ , \new_[1460]_ ,
    \new_[1461]_ , \new_[1462]_ , \new_[1463]_ , \new_[1464]_ ,
    \new_[1465]_ , \new_[1466]_ , \new_[1467]_ , \new_[1468]_ ,
    \new_[1469]_ , \new_[1470]_ , \new_[1471]_ , \new_[1472]_ ,
    \new_[1473]_ , \new_[1474]_ , \new_[1475]_ , \new_[1476]_ ,
    \new_[1477]_ , \new_[1478]_ , \new_[1479]_ , \new_[1480]_ ,
    \new_[1481]_ , \new_[1482]_ , \new_[1483]_ , \new_[1484]_ ,
    \new_[1485]_ , \new_[1486]_ , \new_[1487]_ , \new_[1488]_ ,
    \new_[1489]_ , \new_[1490]_ , \new_[1491]_ , \new_[1492]_ ,
    \new_[1493]_ , \new_[1494]_ , \new_[1495]_ , \new_[1496]_ ,
    \new_[1497]_ , \new_[1498]_ , \new_[1499]_ , \new_[1500]_ ,
    \new_[1501]_ , \new_[1502]_ , \new_[1503]_ , \new_[1504]_ ,
    \new_[1505]_ , \new_[1506]_ , \new_[1507]_ , \new_[1508]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1512]_ ,
    \new_[1513]_ , \new_[1514]_ , \new_[1515]_ , \new_[1516]_ ,
    \new_[1517]_ , \new_[1518]_ , \new_[1519]_ , \new_[1520]_ ,
    \new_[1521]_ , \new_[1522]_ , \new_[1523]_ , \new_[1524]_ ,
    \new_[1525]_ , \new_[1526]_ , \new_[1527]_ , \new_[1528]_ ,
    \new_[1529]_ , \new_[1530]_ , \new_[1531]_ , \new_[1532]_ ,
    \new_[1533]_ , \new_[1534]_ , \new_[1535]_ , \new_[1536]_ ,
    \new_[1537]_ , \new_[1538]_ , \new_[1539]_ , \new_[1540]_ ,
    \new_[1541]_ , \new_[1542]_ , \new_[1543]_ , \new_[1544]_ ,
    \new_[1545]_ , \new_[1546]_ , \new_[1547]_ , \new_[1548]_ ,
    \new_[1549]_ , \new_[1550]_ , \new_[1551]_ , \new_[1552]_ ,
    \new_[1553]_ , \new_[1554]_ , \new_[1555]_ , \new_[1556]_ ,
    \new_[1557]_ , \new_[1558]_ , \new_[1559]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1562]_ , \new_[1563]_ , \new_[1564]_ ,
    \new_[1565]_ , \new_[1566]_ , \new_[1567]_ , \new_[1568]_ ,
    \new_[1569]_ , \new_[1570]_ , \new_[1571]_ , \new_[1572]_ ,
    \new_[1573]_ , \new_[1574]_ , \new_[1575]_ , \new_[1576]_ ,
    \new_[1577]_ , \new_[1578]_ , \new_[1579]_ , \new_[1580]_ ,
    \new_[1581]_ , \new_[1582]_ , \new_[1583]_ , \new_[1584]_ ,
    \new_[1585]_ , \new_[1586]_ , \new_[1587]_ , \new_[1588]_ ,
    \new_[1589]_ , \new_[1590]_ , \new_[1591]_ , \new_[1592]_ ,
    \new_[1593]_ , \new_[1594]_ , \new_[1595]_ , \new_[1596]_ ,
    \new_[1597]_ , \new_[1598]_ , \new_[1599]_ , \new_[1600]_ ,
    \new_[1601]_ , \new_[1602]_ , \new_[1603]_ , \new_[1604]_ ,
    \new_[1605]_ , \new_[1606]_ , \new_[1607]_ , \new_[1608]_ ,
    \new_[1609]_ , \new_[1610]_ , \new_[1611]_ , \new_[1612]_ ,
    \new_[1613]_ , \new_[1614]_ , \new_[1615]_ , \new_[1616]_ ,
    \new_[1617]_ , \new_[1618]_ , \new_[1619]_ , \new_[1620]_ ,
    \new_[1621]_ , \new_[1622]_ , \new_[1623]_ , \new_[1624]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1627]_ , \new_[1628]_ ,
    \new_[1629]_ , \new_[1630]_ , \new_[1631]_ , \new_[1632]_ ,
    \new_[1633]_ , \new_[1634]_ , \new_[1635]_ , \new_[1636]_ ,
    \new_[1637]_ , \new_[1638]_ , \new_[1639]_ , \new_[1640]_ ,
    \new_[1641]_ , \new_[1642]_ , \new_[1643]_ , \new_[1644]_ ,
    \new_[1645]_ , \new_[1646]_ , \new_[1647]_ , \new_[1648]_ ,
    \new_[1649]_ , \new_[1650]_ , \new_[1651]_ , \new_[1652]_ ,
    \new_[1653]_ , \new_[1654]_ , \new_[1655]_ , \new_[1656]_ ,
    \new_[1657]_ , \new_[1658]_ , \new_[1659]_ , \new_[1660]_ ,
    \new_[1661]_ , \new_[1662]_ , \new_[1663]_ , \new_[1664]_ ,
    \new_[1665]_ , \new_[1666]_ , \new_[1667]_ , \new_[1668]_ ,
    \new_[1669]_ , \new_[1670]_ , \new_[1671]_ , \new_[1672]_ ,
    \new_[1673]_ , \new_[1674]_ , \new_[1675]_ , \new_[1676]_ ,
    \new_[1677]_ , \new_[1678]_ , \new_[1679]_ , \new_[1680]_ ,
    \new_[1681]_ , \new_[1682]_ , \new_[1683]_ , \new_[1684]_ ,
    \new_[1685]_ , \new_[1686]_ , \new_[1687]_ , \new_[1688]_ ,
    \new_[1689]_ , \new_[1690]_ , \new_[1691]_ , \new_[1692]_ ,
    \new_[1693]_ , \new_[1694]_ , \new_[1695]_ , \new_[1696]_ ,
    \new_[1697]_ , \new_[1698]_ , \new_[1699]_ , \new_[1700]_ ,
    \new_[1701]_ , \new_[1702]_ , \new_[1703]_ , \new_[1704]_ ,
    \new_[1705]_ , \new_[1706]_ , \new_[1707]_ , \new_[1708]_ ,
    \new_[1709]_ , \new_[1710]_ , \new_[1711]_ , \new_[1712]_ ,
    \new_[1713]_ , \new_[1714]_ , \new_[1715]_ , \new_[1716]_ ,
    \new_[1717]_ , \new_[1718]_ , \new_[1719]_ , \new_[1720]_ ,
    \new_[1721]_ , \new_[1722]_ , \new_[1723]_ , \new_[1724]_ ,
    \new_[1725]_ , \new_[1726]_ , \new_[1727]_ , \new_[1728]_ ,
    \new_[1729]_ , \new_[1730]_ , \new_[1731]_ , \new_[1732]_ ,
    \new_[1733]_ , \new_[1734]_ , \new_[1735]_ , \new_[1736]_ ,
    \new_[1737]_ , \new_[1738]_ , \new_[1739]_ , \new_[1740]_ ,
    \new_[1741]_ , \new_[1742]_ , \new_[1743]_ , \new_[1744]_ ,
    \new_[1745]_ , \new_[1746]_ , \new_[1747]_ , \new_[1748]_ ,
    \new_[1749]_ , \new_[1750]_ , \new_[1751]_ , \new_[1752]_ ,
    \new_[1753]_ , \new_[1754]_ , \new_[1755]_ , \new_[1756]_ ,
    \new_[1757]_ , \new_[1758]_ , \new_[1759]_ , \new_[1760]_ ,
    \new_[1761]_ , \new_[1762]_ , \new_[1763]_ , \new_[1764]_ ,
    \new_[1765]_ , \new_[1766]_ , \new_[1767]_ , \new_[1768]_ ,
    \new_[1769]_ , \new_[1770]_ , \new_[1771]_ , \new_[1772]_ ,
    \new_[1773]_ , \new_[1774]_ , \new_[1775]_ , \new_[1776]_ ,
    \new_[1777]_ , \new_[1778]_ , \new_[1779]_ , \new_[1780]_ ,
    \new_[1781]_ , \new_[1782]_ , \new_[1783]_ , \new_[1784]_ ,
    \new_[1785]_ , \new_[1786]_ , \new_[1787]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1791]_ , \new_[1792]_ ,
    \new_[1793]_ , \new_[1794]_ , \new_[1795]_ , \new_[1796]_ ,
    \new_[1797]_ , \new_[1798]_ , \new_[1799]_ , \new_[1800]_ ,
    \new_[1801]_ , \new_[1802]_ , \new_[1803]_ , \new_[1804]_ ,
    \new_[1805]_ , \new_[1806]_ , \new_[1807]_ , \new_[1808]_ ,
    \new_[1809]_ , \new_[1810]_ , \new_[1811]_ , \new_[1812]_ ,
    \new_[1813]_ , \new_[1814]_ , \new_[1815]_ , \new_[1816]_ ,
    \new_[1817]_ , \new_[1818]_ , \new_[1819]_ , \new_[1820]_ ,
    \new_[1821]_ , \new_[1822]_ , \new_[1823]_ , \new_[1824]_ ,
    \new_[1825]_ , \new_[1826]_ , \new_[1827]_ , \new_[1828]_ ,
    \new_[1829]_ , \new_[1830]_ , \new_[1831]_ , \new_[1832]_ ,
    \new_[1833]_ , \new_[1834]_ , \new_[1835]_ , \new_[1836]_ ,
    \new_[1837]_ , \new_[1838]_ , \new_[1839]_ , \new_[1840]_ ,
    \new_[1841]_ , \new_[1842]_ , \new_[1843]_ , \new_[1844]_ ,
    \new_[1845]_ , \new_[1846]_ , \new_[1847]_ , \new_[1848]_ ,
    \new_[1849]_ , \new_[1850]_ , \new_[1851]_ , \new_[1852]_ ,
    \new_[1853]_ , \new_[1854]_ , \new_[1855]_ , \new_[1856]_ ,
    \new_[1857]_ , \new_[1858]_ , \new_[1859]_ , \new_[1860]_ ,
    \new_[1861]_ , \new_[1862]_ , \new_[1863]_ , \new_[1864]_ ,
    \new_[1865]_ , \new_[1866]_ , \new_[1867]_ , \new_[1868]_ ,
    \new_[1869]_ , \new_[1870]_ , \new_[1871]_ , \new_[1872]_ ,
    \new_[1873]_ , \new_[1874]_ , \new_[1875]_ , \new_[1876]_ ,
    \new_[1877]_ , \new_[1878]_ , \new_[1879]_ , \new_[1880]_ ,
    \new_[1881]_ , \new_[1882]_ , \new_[1883]_ , \new_[1884]_ ,
    \new_[1885]_ , \new_[1886]_ , \new_[1887]_ , \new_[1888]_ ,
    \new_[1889]_ , \new_[1890]_ , \new_[1891]_ , \new_[1892]_ ,
    \new_[1893]_ , \new_[1894]_ , \new_[1895]_ , \new_[1896]_ ,
    \new_[1897]_ , \new_[1898]_ , \new_[1899]_ , \new_[1900]_ ,
    \new_[1901]_ , \new_[1902]_ , \new_[1903]_ , \new_[1904]_ ,
    \new_[1905]_ , \new_[1906]_ , \new_[1907]_ , \new_[1908]_ ,
    \new_[1909]_ , \new_[1910]_ , \new_[1911]_ , \new_[1912]_ ,
    \new_[1913]_ , \new_[1914]_ , \new_[1915]_ , \new_[1916]_ ,
    \new_[1917]_ , \new_[1918]_ , \new_[1919]_ , \new_[1920]_ ,
    \new_[1921]_ , \new_[1922]_ , \new_[1923]_ , \new_[1924]_ ,
    \new_[1925]_ , \new_[1926]_ , \new_[1927]_ , \new_[1928]_ ,
    \new_[1929]_ , \new_[1930]_ , \new_[1931]_ , \new_[1932]_ ,
    \new_[1933]_ , \new_[1934]_ , \new_[1935]_ , \new_[1936]_ ,
    \new_[1937]_ , \new_[1938]_ , \new_[1939]_ , \new_[1940]_ ,
    \new_[1941]_ , \new_[1942]_ , \new_[1943]_ , \new_[1944]_ ,
    \new_[1945]_ , \new_[1946]_ , \new_[1947]_ , \new_[1948]_ ,
    \new_[1949]_ , \new_[1950]_ , \new_[1951]_ , \new_[1952]_ ,
    \new_[1953]_ , \new_[1954]_ , \new_[1955]_ , \new_[1956]_ ,
    \new_[1957]_ , \new_[1958]_ , \new_[1959]_ , \new_[1960]_ ,
    \new_[1961]_ , \new_[1962]_ , \new_[1963]_ , \new_[1964]_ ,
    \new_[1965]_ , \new_[1966]_ , \new_[1967]_ , \new_[1968]_ ,
    \new_[1969]_ , \new_[1970]_ , \new_[1971]_ , \new_[1972]_ ,
    \new_[1973]_ , \new_[1974]_ , \new_[1975]_ , \new_[1976]_ ,
    \new_[1977]_ , \new_[1978]_ , \new_[1979]_ , \new_[1980]_ ,
    \new_[1981]_ , \new_[1982]_ , \new_[1983]_ , \new_[1984]_ ,
    \new_[1985]_ , \new_[1986]_ , \new_[1987]_ , \new_[1988]_ ,
    \new_[1989]_ , \new_[1990]_ , \new_[1991]_ , \new_[1992]_ ,
    \new_[1993]_ , \new_[1994]_ , \new_[1995]_ , \new_[1996]_ ,
    \new_[1997]_ , \new_[1998]_ , \new_[1999]_ , \new_[2000]_ ,
    \new_[2001]_ , \new_[2002]_ , \new_[2003]_ , \new_[2004]_ ,
    \new_[2005]_ , \new_[2006]_ , \new_[2007]_ , \new_[2008]_ ,
    \new_[2009]_ , \new_[2010]_ , \new_[2011]_ , \new_[2012]_ ,
    \new_[2013]_ , \new_[2014]_ , \new_[2015]_ , \new_[2016]_ ,
    \new_[2017]_ , \new_[2018]_ , \new_[2019]_ , \new_[2020]_ ,
    \new_[2021]_ , \new_[2022]_ , \new_[2023]_ , \new_[2024]_ ,
    \new_[2025]_ , \new_[2026]_ , \new_[2027]_ , \new_[2028]_ ,
    \new_[2029]_ , \new_[2030]_ , \new_[2031]_ , \new_[2032]_ ,
    \new_[2033]_ , \new_[2034]_ , \new_[2035]_ , \new_[2036]_ ,
    \new_[2037]_ , \new_[2038]_ , \new_[2039]_ , \new_[2040]_ ,
    \new_[2041]_ , \new_[2042]_ , \new_[2043]_ , \new_[2044]_ ,
    \new_[2045]_ , \new_[2046]_ , \new_[2047]_ , \new_[2048]_ ,
    \new_[2049]_ , \new_[2050]_ , \new_[2051]_ , \new_[2052]_ ,
    \new_[2053]_ , \new_[2054]_ , \new_[2055]_ , \new_[2056]_ ,
    \new_[2057]_ , \new_[2058]_ , \new_[2059]_ , \new_[2060]_ ,
    \new_[2061]_ , \new_[2062]_ , \new_[2063]_ , \new_[2064]_ ,
    \new_[2065]_ , \new_[2066]_ , \new_[2067]_ , \new_[2068]_ ,
    \new_[2069]_ , \new_[2070]_ , \new_[2071]_ , \new_[2072]_ ,
    \new_[2073]_ , \new_[2074]_ , \new_[2075]_ , \new_[2076]_ ,
    \new_[2077]_ , \new_[2078]_ , \new_[2079]_ , \new_[2080]_ ,
    \new_[2081]_ , \new_[2082]_ , \new_[2083]_ , \new_[2084]_ ,
    \new_[2085]_ , \new_[2086]_ , \new_[2087]_ , \new_[2088]_ ,
    \new_[2089]_ , \new_[2090]_ , \new_[2091]_ , \new_[2092]_ ,
    \new_[2093]_ , \new_[2094]_ , \new_[2095]_ , \new_[2096]_ ,
    \new_[2097]_ , \new_[2098]_ , \new_[2099]_ , \new_[2100]_ ,
    \new_[2101]_ , \new_[2102]_ , \new_[2103]_ , \new_[2104]_ ,
    \new_[2105]_ , \new_[2106]_ , \new_[2107]_ , \new_[2108]_ ,
    \new_[2109]_ , \new_[2110]_ , \new_[2111]_ , \new_[2112]_ ,
    \new_[2113]_ , \new_[2114]_ , \new_[2115]_ , \new_[2116]_ ,
    \new_[2117]_ , \new_[2118]_ , \new_[2119]_ , \new_[2120]_ ,
    \new_[2121]_ , \new_[2122]_ , \new_[2123]_ , \new_[2124]_ ,
    \new_[2125]_ , \new_[2126]_ , \new_[2127]_ , \new_[2128]_ ,
    \new_[2129]_ , \new_[2130]_ , \new_[2131]_ , \new_[2132]_ ,
    \new_[2133]_ , \new_[2134]_ , \new_[2135]_ , \new_[2136]_ ,
    \new_[2137]_ , \new_[2138]_ , \new_[2139]_ , \new_[2140]_ ,
    \new_[2141]_ , \new_[2142]_ , \new_[2143]_ , \new_[2144]_ ,
    \new_[2145]_ , \new_[2146]_ , \new_[2147]_ , \new_[2148]_ ,
    \new_[2149]_ , \new_[2150]_ , \new_[2151]_ , \new_[2152]_ ,
    \new_[2153]_ , \new_[2154]_ , \new_[2155]_ , \new_[2156]_ ,
    \new_[2157]_ , \new_[2158]_ , \new_[2159]_ , \new_[2160]_ ,
    \new_[2161]_ , \new_[2162]_ , \new_[2163]_ , \new_[2164]_ ,
    \new_[2165]_ , \new_[2166]_ , \new_[2167]_ , \new_[2168]_ ,
    \new_[2169]_ , \new_[2170]_ , \new_[2171]_ , \new_[2172]_ ,
    \new_[2173]_ , \new_[2174]_ , \new_[2175]_ , \new_[2176]_ ,
    \new_[2177]_ , \new_[2178]_ , \new_[2179]_ , \new_[2180]_ ,
    \new_[2181]_ , \new_[2182]_ , \new_[2183]_ , \new_[2184]_ ,
    \new_[2185]_ , \new_[2186]_ , \new_[2187]_ , \new_[2188]_ ,
    \new_[2189]_ , \new_[2190]_ , \new_[2191]_ , \new_[2192]_ ,
    \new_[2193]_ , \new_[2194]_ , \new_[2195]_ , \new_[2196]_ ,
    \new_[2197]_ , \new_[2198]_ , \new_[2199]_ , \new_[2200]_ ,
    \new_[2201]_ , \new_[2202]_ , \new_[2203]_ , \new_[2204]_ ,
    \new_[2205]_ , \new_[2206]_ , \new_[2207]_ , \new_[2208]_ ,
    \new_[2209]_ , \new_[2210]_ , \new_[2211]_ , \new_[2212]_ ,
    \new_[2213]_ , \new_[2214]_ , \new_[2215]_ , \new_[2216]_ ,
    \new_[2217]_ , \new_[2218]_ , \new_[2219]_ , \new_[2220]_ ,
    \new_[2221]_ , \new_[2222]_ , \new_[2223]_ , \new_[2224]_ ,
    \new_[2225]_ , \new_[2226]_ , \new_[2227]_ , \new_[2228]_ ,
    \new_[2229]_ , \new_[2230]_ , \new_[2231]_ , \new_[2232]_ ,
    \new_[2233]_ , \new_[2234]_ , \new_[2235]_ , \new_[2236]_ ,
    \new_[2237]_ , \new_[2238]_ , \new_[2239]_ , \new_[2240]_ ,
    \new_[2241]_ , \new_[2242]_ , \new_[2243]_ , \new_[2244]_ ,
    \new_[2245]_ , \new_[2246]_ , \new_[2247]_ , \new_[2248]_ ,
    \new_[2249]_ , \new_[2250]_ , \new_[2251]_ , \new_[2252]_ ,
    \new_[2253]_ , \new_[2254]_ , \new_[2255]_ , \new_[2256]_ ,
    \new_[2257]_ , \new_[2258]_ , \new_[2259]_ , \new_[2260]_ ,
    \new_[2261]_ , \new_[2262]_ , \new_[2263]_ , \new_[2264]_ ,
    \new_[2265]_ , \new_[2266]_ , \new_[2267]_ , \new_[2268]_ ,
    \new_[2269]_ , \new_[2270]_ , \new_[2271]_ , \new_[2272]_ ,
    \new_[2273]_ , \new_[2274]_ , \new_[2275]_ , \new_[2276]_ ,
    \new_[2277]_ , \new_[2278]_ , \new_[2279]_ , \new_[2280]_ ,
    \new_[2281]_ , \new_[2282]_ , \new_[2283]_ , \new_[2284]_ ,
    \new_[2285]_ , \new_[2286]_ , \new_[2287]_ , \new_[2288]_ ,
    \new_[2289]_ , \new_[2290]_ , \new_[2291]_ , \new_[2292]_ ,
    \new_[2293]_ , \new_[2294]_ , \new_[2295]_ , \new_[2296]_ ,
    \new_[2297]_ , \new_[2298]_ , \new_[2299]_ , \new_[2300]_ ,
    \new_[2301]_ , \new_[2302]_ , \new_[2303]_ , \new_[2304]_ ,
    \new_[2305]_ , \new_[2306]_ , \new_[2307]_ , \new_[2308]_ ,
    \new_[2309]_ , \new_[2310]_ , \new_[2311]_ , \new_[2312]_ ,
    \new_[2313]_ , \new_[2314]_ , \new_[2315]_ , \new_[2316]_ ,
    \new_[2317]_ , \new_[2318]_ , \new_[2319]_ , \new_[2320]_ ,
    \new_[2321]_ , \new_[2322]_ , \new_[2323]_ , \new_[2324]_ ,
    \new_[2325]_ , \new_[2326]_ , \new_[2327]_ , \new_[2328]_ ,
    \new_[2329]_ , \new_[2330]_ , \new_[2331]_ , \new_[2332]_ ,
    \new_[2333]_ , \new_[2334]_ , \new_[2335]_ , \new_[2336]_ ,
    \new_[2337]_ , \new_[2338]_ , \new_[2339]_ , \new_[2340]_ ,
    \new_[2341]_ , \new_[2342]_ , \new_[2343]_ , \new_[2344]_ ,
    \new_[2345]_ , \new_[2346]_ , \new_[2347]_ , \new_[2348]_ ,
    \new_[2349]_ , \new_[2350]_ , \new_[2351]_ , \new_[2352]_ ,
    \new_[2353]_ , \new_[2354]_ , \new_[2355]_ , \new_[2356]_ ,
    \new_[2357]_ , \new_[2358]_ , \new_[2359]_ , \new_[2360]_ ,
    \new_[2361]_ , \new_[2362]_ , \new_[2363]_ , \new_[2364]_ ,
    \new_[2365]_ , \new_[2366]_ , \new_[2367]_ , \new_[2368]_ ,
    \new_[2369]_ , \new_[2370]_ , \new_[2371]_ , \new_[2372]_ ,
    \new_[2373]_ , \new_[2374]_ , \new_[2375]_ , \new_[2376]_ ,
    \new_[2377]_ , \new_[2378]_ , \new_[2379]_ , \new_[2380]_ ,
    \new_[2381]_ , \new_[2382]_ , \new_[2383]_ , \new_[2384]_ ,
    \new_[2385]_ , \new_[2386]_ , \new_[2387]_ , \new_[2388]_ ,
    \new_[2389]_ , \new_[2390]_ , \new_[2391]_ , \new_[2392]_ ,
    \new_[2393]_ , \new_[2394]_ , \new_[2395]_ , \new_[2396]_ ,
    \new_[2397]_ , \new_[2398]_ , \new_[2399]_ , \new_[2400]_ ,
    \new_[2401]_ , \new_[2402]_ , \new_[2403]_ , \new_[2404]_ ,
    \new_[2405]_ , \new_[2406]_ , \new_[2407]_ , \new_[2408]_ ,
    \new_[2409]_ , \new_[2410]_ , \new_[2411]_ , \new_[2412]_ ,
    \new_[2413]_ , \new_[2414]_ , \new_[2415]_ , \new_[2416]_ ,
    \new_[2417]_ , \new_[2418]_ , \new_[2419]_ , \new_[2420]_ ,
    \new_[2421]_ , \new_[2422]_ , \new_[2423]_ , \new_[2424]_ ,
    \new_[2425]_ , \new_[2426]_ , \new_[2427]_ , \new_[2428]_ ,
    \new_[2429]_ , \new_[2430]_ , \new_[2431]_ , \new_[2432]_ ,
    \new_[2433]_ , \new_[2434]_ , \new_[2435]_ , \new_[2436]_ ,
    \new_[2437]_ , \new_[2438]_ , \new_[2439]_ , \new_[2440]_ ,
    \new_[2441]_ , \new_[2442]_ , \new_[2443]_ , \new_[2444]_ ,
    \new_[2445]_ , \new_[2446]_ , \new_[2447]_ , \new_[2448]_ ,
    \new_[2449]_ , \new_[2450]_ , \new_[2451]_ , \new_[2452]_ ,
    \new_[2453]_ , \new_[2454]_ , \new_[2455]_ , \new_[2456]_ ,
    \new_[2457]_ , \new_[2458]_ , \new_[2459]_ , \new_[2460]_ ,
    \new_[2461]_ , \new_[2462]_ , \new_[2463]_ , \new_[2464]_ ,
    \new_[2465]_ , \new_[2466]_ , \new_[2467]_ , \new_[2468]_ ,
    \new_[2469]_ , \new_[2470]_ , \new_[2471]_ , \new_[2472]_ ,
    \new_[2473]_ , \new_[2474]_ , \new_[2475]_ , \new_[2476]_ ,
    \new_[2477]_ , \new_[2478]_ , \new_[2479]_ , \new_[2480]_ ,
    \new_[2481]_ , \new_[2482]_ , \new_[2483]_ , \new_[2484]_ ,
    \new_[2485]_ , \new_[2486]_ , \new_[2487]_ , \new_[2488]_ ,
    \new_[2489]_ , \new_[2490]_ , \new_[2491]_ , \new_[2492]_ ,
    \new_[2493]_ , \new_[2494]_ , \new_[2495]_ , \new_[2496]_ ,
    \new_[2497]_ , \new_[2498]_ , \new_[2499]_ , \new_[2500]_ ,
    \new_[2501]_ , \new_[2502]_ , \new_[2503]_ , \new_[2504]_ ,
    \new_[2505]_ , \new_[2506]_ , \new_[2507]_ , \new_[2508]_ ,
    \new_[2509]_ , \new_[2510]_ , \new_[2511]_ , \new_[2512]_ ,
    \new_[2513]_ , \new_[2514]_ , \new_[2515]_ , \new_[2516]_ ,
    \new_[2517]_ , \new_[2518]_ , \new_[2519]_ , \new_[2520]_ ,
    \new_[2521]_ , \new_[2522]_ , \new_[2523]_ , \new_[2524]_ ,
    \new_[2525]_ , \new_[2526]_ , \new_[2527]_ , \new_[2528]_ ,
    \new_[2529]_ , \new_[2530]_ , \new_[2531]_ , \new_[2532]_ ,
    \new_[2533]_ , \new_[2534]_ , \new_[2535]_ , \new_[2536]_ ,
    \new_[2537]_ , \new_[2538]_ , \new_[2539]_ , \new_[2540]_ ,
    \new_[2541]_ , \new_[2542]_ , \new_[2543]_ , \new_[2544]_ ,
    \new_[2545]_ , \new_[2546]_ , \new_[2547]_ , \new_[2548]_ ,
    \new_[2549]_ , \new_[2550]_ , \new_[2551]_ , \new_[2552]_ ,
    \new_[2553]_ , \new_[2554]_ , \new_[2555]_ , \new_[2556]_ ,
    \new_[2557]_ , \new_[2558]_ , \new_[2559]_ , \new_[2560]_ ,
    \new_[2561]_ , \new_[2562]_ , \new_[2563]_ , \new_[2564]_ ,
    \new_[2565]_ , \new_[2566]_ , \new_[2567]_ , \new_[2568]_ ,
    \new_[2569]_ , \new_[2570]_ , \new_[2571]_ , \new_[2572]_ ,
    \new_[2573]_ , \new_[2574]_ , \new_[2575]_ , \new_[2576]_ ,
    \new_[2577]_ , \new_[2578]_ , \new_[2579]_ , \new_[2580]_ ,
    \new_[2581]_ , \new_[2582]_ , \new_[2583]_ , \new_[2584]_ ,
    \new_[2585]_ , \new_[2586]_ , \new_[2587]_ , \new_[2588]_ ,
    \new_[2589]_ , \new_[2590]_ , \new_[2591]_ , \new_[2592]_ ,
    \new_[2593]_ , \new_[2594]_ , \new_[2595]_ , \new_[2596]_ ,
    \new_[2597]_ , \new_[2598]_ , \new_[2599]_ , \new_[2600]_ ,
    \new_[2601]_ , \new_[2602]_ , \new_[2603]_ , \new_[2604]_ ,
    \new_[2605]_ , \new_[2606]_ , \new_[2607]_ , \new_[2608]_ ,
    \new_[2609]_ , \new_[2610]_ , \new_[2611]_ , \new_[2612]_ ,
    \new_[2613]_ , \new_[2614]_ , \new_[2615]_ , \new_[2616]_ ,
    \new_[2617]_ , \new_[2618]_ , \new_[2619]_ , \new_[2620]_ ,
    \new_[2621]_ , \new_[2622]_ , \new_[2623]_ , \new_[2624]_ ,
    \new_[2625]_ , \new_[2626]_ , \new_[2627]_ , \new_[2628]_ ,
    \new_[2629]_ , \new_[2630]_ , \new_[2631]_ , \new_[2632]_ ,
    \new_[2633]_ , \new_[2634]_ , \new_[2635]_ , \new_[2636]_ ,
    \new_[2637]_ , \new_[2638]_ , \new_[2639]_ , \new_[2640]_ ,
    \new_[2641]_ , \new_[2642]_ , \new_[2643]_ , \new_[2644]_ ,
    \new_[2645]_ , \new_[2646]_ , \new_[2647]_ , \new_[2648]_ ,
    \new_[2649]_ , \new_[2650]_ , \new_[2651]_ , \new_[2652]_ ,
    \new_[2653]_ , \new_[2654]_ , \new_[2655]_ , \new_[2656]_ ,
    \new_[2657]_ , \new_[2658]_ , \new_[2659]_ , \new_[2660]_ ,
    \new_[2661]_ , \new_[2662]_ , \new_[2663]_ , \new_[2664]_ ,
    \new_[2665]_ , \new_[2666]_ , \new_[2667]_ , \new_[2668]_ ,
    \new_[2669]_ , \new_[2670]_ , \new_[2671]_ , \new_[2672]_ ,
    \new_[2673]_ , \new_[2674]_ , \new_[2675]_ , \new_[2676]_ ,
    \new_[2677]_ , \new_[2678]_ , \new_[2679]_ , \new_[2680]_ ,
    \new_[2681]_ , \new_[2682]_ , \new_[2683]_ , \new_[2684]_ ,
    \new_[2685]_ , \new_[2686]_ , \new_[2687]_ , \new_[2688]_ ,
    \new_[2689]_ , \new_[2690]_ , \new_[2691]_ , \new_[2692]_ ,
    \new_[2693]_ , \new_[2694]_ , \new_[2695]_ , \new_[2696]_ ,
    \new_[2697]_ , \new_[2698]_ , \new_[2699]_ , \new_[2700]_ ,
    \new_[2701]_ , \new_[2702]_ , \new_[2703]_ , \new_[2704]_ ,
    \new_[2705]_ , \new_[2706]_ , \new_[2707]_ , \new_[2708]_ ,
    \new_[2709]_ , \new_[2710]_ , \new_[2711]_ , \new_[2712]_ ,
    \new_[2713]_ , \new_[2714]_ , \new_[2715]_ , \new_[2716]_ ,
    \new_[2717]_ , \new_[2718]_ , \new_[2719]_ , \new_[2720]_ ,
    \new_[2721]_ , \new_[2722]_ , \new_[2723]_ , \new_[2724]_ ,
    \new_[2725]_ , \new_[2726]_ , \new_[2727]_ , \new_[2728]_ ,
    \new_[2729]_ , \new_[2730]_ , \new_[2731]_ , \new_[2732]_ ,
    \new_[2733]_ , \new_[2734]_ , \new_[2735]_ , \new_[2736]_ ,
    \new_[2737]_ , \new_[2738]_ , \new_[2739]_ , \new_[2740]_ ,
    \new_[2741]_ , \new_[2742]_ , \new_[2743]_ , \new_[2744]_ ,
    \new_[2745]_ , \new_[2746]_ , \new_[2747]_ , \new_[2748]_ ,
    \new_[2749]_ , \new_[2750]_ , \new_[2751]_ , \new_[2752]_ ,
    \new_[2753]_ , \new_[2754]_ , \new_[2755]_ , \new_[2756]_ ,
    \new_[2757]_ , \new_[2758]_ , \new_[2759]_ , \new_[2760]_ ,
    \new_[2761]_ , \new_[2762]_ , \new_[2763]_ , \new_[2764]_ ,
    \new_[2765]_ , \new_[2766]_ , \new_[2767]_ , \new_[2768]_ ,
    \new_[2769]_ , \new_[2770]_ , \new_[2771]_ , \new_[2772]_ ,
    \new_[2773]_ , \new_[2774]_ , \new_[2775]_ , \new_[2776]_ ,
    \new_[2777]_ , \new_[2778]_ , \new_[2779]_ , \new_[2780]_ ,
    \new_[2781]_ , \new_[2782]_ , \new_[2783]_ , \new_[2784]_ ,
    \new_[2785]_ , \new_[2786]_ , \new_[2787]_ , \new_[2788]_ ,
    \new_[2789]_ , \new_[2790]_ , \new_[2791]_ , \new_[2792]_ ,
    \new_[2793]_ , \new_[2794]_ , \new_[2795]_ , \new_[2796]_ ,
    \new_[2797]_ , \new_[2798]_ , \new_[2799]_ , \new_[2800]_ ,
    \new_[2801]_ , \new_[2802]_ , \new_[2803]_ , \new_[2804]_ ,
    \new_[2805]_ , \new_[2806]_ , \new_[2807]_ , \new_[2808]_ ,
    \new_[2809]_ , \new_[2810]_ , \new_[2811]_ , \new_[2812]_ ,
    \new_[2813]_ , \new_[2814]_ , \new_[2815]_ , \new_[2816]_ ,
    \new_[2817]_ , \new_[2818]_ , \new_[2819]_ , \new_[2820]_ ,
    \new_[2821]_ , \new_[2822]_ , \new_[2823]_ , \new_[2824]_ ,
    \new_[2825]_ , \new_[2826]_ , \new_[2827]_ , \new_[2828]_ ,
    \new_[2829]_ , \new_[2830]_ , \new_[2831]_ , \new_[2832]_ ,
    \new_[2833]_ , \new_[2834]_ , \new_[2835]_ , \new_[2836]_ ,
    \new_[2837]_ , \new_[2838]_ , \new_[2839]_ , \new_[2840]_ ,
    \new_[2841]_ , \new_[2842]_ , \new_[2843]_ , \new_[2844]_ ,
    \new_[2845]_ , \new_[2846]_ , \new_[2847]_ , \new_[2848]_ ,
    \new_[2849]_ , \new_[2850]_ , \new_[2851]_ , \new_[2852]_ ,
    \new_[2853]_ , \new_[2854]_ , \new_[2855]_ , \new_[2856]_ ,
    \new_[2857]_ , \new_[2858]_ , \new_[2859]_ , \new_[2860]_ ,
    \new_[2861]_ , \new_[2862]_ , \new_[2863]_ , \new_[2864]_ ,
    \new_[2865]_ , \new_[2866]_ , \new_[2867]_ , \new_[2868]_ ,
    \new_[2869]_ , \new_[2870]_ , \new_[2871]_ , \new_[2872]_ ,
    \new_[2873]_ , \new_[2874]_ , \new_[2875]_ , \new_[2876]_ ,
    \new_[2877]_ , \new_[2878]_ , \new_[2879]_ , \new_[2880]_ ,
    \new_[2881]_ , \new_[2882]_ , \new_[2883]_ , \new_[2884]_ ,
    \new_[2885]_ , \new_[2886]_ , \new_[2887]_ , \new_[2888]_ ,
    \new_[2889]_ , \new_[2890]_ , \new_[2891]_ , \new_[2892]_ ,
    \new_[2893]_ , \new_[2894]_ , \new_[2895]_ , \new_[2896]_ ,
    \new_[2897]_ , \new_[2898]_ , \new_[2899]_ , \new_[2900]_ ,
    \new_[2901]_ , \new_[2902]_ , \new_[2903]_ , \new_[2904]_ ,
    \new_[2905]_ , \new_[2906]_ , \new_[2907]_ , \new_[2908]_ ,
    \new_[2909]_ , \new_[2910]_ , \new_[2911]_ , \new_[2912]_ ,
    \new_[2913]_ , \new_[2914]_ , \new_[2915]_ , \new_[2916]_ ,
    \new_[2917]_ , \new_[2918]_ , \new_[2919]_ , \new_[2920]_ ,
    \new_[2921]_ , \new_[2922]_ , \new_[2923]_ , \new_[2924]_ ,
    \new_[2925]_ , \new_[2926]_ , \new_[2927]_ , \new_[2928]_ ,
    \new_[2929]_ , \new_[2930]_ , \new_[2931]_ , \new_[2932]_ ,
    \new_[2933]_ , \new_[2934]_ , \new_[2935]_ , \new_[2936]_ ,
    \new_[2937]_ , \new_[2938]_ , \new_[2939]_ , \new_[2940]_ ,
    \new_[2941]_ , \new_[2942]_ , \new_[2943]_ , \new_[2944]_ ,
    \new_[2945]_ , \new_[2946]_ , \new_[2947]_ , \new_[2948]_ ,
    \new_[2949]_ , \new_[2950]_ , \new_[2951]_ , \new_[2952]_ ,
    \new_[2953]_ , \new_[2954]_ , \new_[2955]_ , \new_[2956]_ ,
    \new_[2957]_ , \new_[2958]_ , \new_[2959]_ , \new_[2960]_ ,
    \new_[2961]_ , \new_[2962]_ , \new_[2963]_ , \new_[2964]_ ,
    \new_[2965]_ , \new_[2966]_ , \new_[2967]_ , \new_[2968]_ ,
    \new_[2969]_ , \new_[2970]_ , \new_[2971]_ , \new_[2972]_ ,
    \new_[2973]_ , \new_[2974]_ , \new_[2975]_ , \new_[2976]_ ,
    \new_[2977]_ , \new_[2978]_ , \new_[2979]_ , \new_[2980]_ ,
    \new_[2981]_ , \new_[2982]_ , \new_[2983]_ , \new_[2984]_ ,
    \new_[2985]_ , \new_[2986]_ , \new_[2987]_ , \new_[2988]_ ,
    \new_[2989]_ , \new_[2990]_ , \new_[2991]_ , \new_[2992]_ ,
    \new_[2993]_ , \new_[2994]_ , \new_[2995]_ , \new_[2996]_ ,
    \new_[2997]_ , \new_[2998]_ , \new_[2999]_ , \new_[3000]_ ,
    \new_[3001]_ , \new_[3002]_ , \new_[3003]_ , \new_[3004]_ ,
    \new_[3005]_ , \new_[3006]_ , \new_[3007]_ , \new_[3008]_ ,
    \new_[3009]_ , \new_[3010]_ , \new_[3011]_ , \new_[3012]_ ,
    \new_[3013]_ , \new_[3014]_ , \new_[3015]_ , \new_[3016]_ ,
    \new_[3017]_ , \new_[3018]_ , \new_[3019]_ , \new_[3020]_ ,
    \new_[3021]_ , \new_[3022]_ , \new_[3023]_ , \new_[3024]_ ,
    \new_[3025]_ , \new_[3026]_ , \new_[3027]_ , \new_[3028]_ ,
    \new_[3029]_ , \new_[3030]_ , \new_[3031]_ , \new_[3032]_ ,
    \new_[3033]_ , \new_[3034]_ , \new_[3035]_ , \new_[3036]_ ,
    \new_[3037]_ , \new_[3038]_ , \new_[3039]_ , \new_[3040]_ ,
    \new_[3041]_ , \new_[3042]_ , \new_[3043]_ , \new_[3044]_ ,
    \new_[3045]_ , \new_[3046]_ , \new_[3047]_ , \new_[3048]_ ,
    \new_[3049]_ , \new_[3050]_ , \new_[3051]_ , \new_[3052]_ ,
    \new_[3053]_ , \new_[3054]_ , \new_[3055]_ , \new_[3056]_ ,
    \new_[3057]_ , \new_[3058]_ , \new_[3059]_ , \new_[3060]_ ,
    \new_[3061]_ , \new_[3062]_ , \new_[3063]_ , \new_[3064]_ ,
    \new_[3065]_ , \new_[3066]_ , \new_[3067]_ , \new_[3068]_ ,
    \new_[3069]_ , \new_[3070]_ , \new_[3071]_ , \new_[3072]_ ,
    \new_[3073]_ , \new_[3074]_ , \new_[3075]_ , \new_[3076]_ ,
    \new_[3077]_ , \new_[3078]_ , \new_[3079]_ , \new_[3080]_ ,
    \new_[3081]_ , \new_[3082]_ , \new_[3083]_ , \new_[3084]_ ,
    \new_[3085]_ , \new_[3086]_ , \new_[3087]_ , \new_[3088]_ ,
    \new_[3089]_ , \new_[3090]_ , \new_[3091]_ , \new_[3092]_ ,
    \new_[3093]_ , \new_[3094]_ , \new_[3095]_ , \new_[3096]_ ,
    \new_[3097]_ , \new_[3098]_ , \new_[3099]_ , \new_[3100]_ ,
    \new_[3101]_ , \new_[3102]_ , \new_[3103]_ , \new_[3104]_ ,
    \new_[3105]_ , \new_[3106]_ , \new_[3107]_ , \new_[3108]_ ,
    \new_[3109]_ , \new_[3110]_ , \new_[3111]_ , \new_[3112]_ ,
    \new_[3113]_ , \new_[3114]_ , \new_[3115]_ , \new_[3116]_ ,
    \new_[3117]_ , \new_[3118]_ , \new_[3119]_ , \new_[3120]_ ,
    \new_[3121]_ , \new_[3122]_ , \new_[3123]_ , \new_[3124]_ ,
    \new_[3125]_ , \new_[3126]_ , \new_[3127]_ , \new_[3128]_ ,
    \new_[3129]_ , \new_[3130]_ , \new_[3131]_ , \new_[3132]_ ,
    \new_[3133]_ , \new_[3134]_ , \new_[3135]_ , \new_[3136]_ ,
    \new_[3137]_ , \new_[3138]_ , \new_[3139]_ , \new_[3140]_ ,
    \new_[3141]_ , \new_[3142]_ , \new_[3143]_ , \new_[3144]_ ,
    \new_[3145]_ , \new_[3146]_ , \new_[3147]_ , \new_[3148]_ ,
    \new_[3149]_ , \new_[3150]_ , \new_[3151]_ , \new_[3152]_ ,
    \new_[3153]_ , \new_[3154]_ , \new_[3155]_ , \new_[3156]_ ,
    \new_[3157]_ , \new_[3158]_ , \new_[3159]_ , \new_[3160]_ ,
    \new_[3161]_ , \new_[3162]_ , \new_[3163]_ , \new_[3164]_ ,
    \new_[3165]_ , \new_[3166]_ , \new_[3167]_ , \new_[3168]_ ,
    \new_[3169]_ , \new_[3170]_ , \new_[3171]_ , \new_[3172]_ ,
    \new_[3173]_ , \new_[3174]_ , \new_[3178]_ , \new_[3179]_ ,
    \new_[3183]_ , \new_[3184]_ , \new_[3185]_ , \new_[3189]_ ,
    \new_[3190]_ , \new_[3194]_ , \new_[3195]_ , \new_[3196]_ ,
    \new_[3197]_ , \new_[3201]_ , \new_[3202]_ , \new_[3206]_ ,
    \new_[3207]_ , \new_[3208]_ , \new_[3212]_ , \new_[3213]_ ,
    \new_[3217]_ , \new_[3218]_ , \new_[3219]_ , \new_[3220]_ ,
    \new_[3221]_ , \new_[3225]_ , \new_[3226]_ , \new_[3230]_ ,
    \new_[3231]_ , \new_[3232]_ , \new_[3236]_ , \new_[3237]_ ,
    \new_[3241]_ , \new_[3242]_ , \new_[3243]_ , \new_[3244]_ ,
    \new_[3248]_ , \new_[3249]_ , \new_[3253]_ , \new_[3254]_ ,
    \new_[3255]_ , \new_[3259]_ , \new_[3260]_ , \new_[3263]_ ,
    \new_[3266]_ , \new_[3267]_ , \new_[3268]_ , \new_[3269]_ ,
    \new_[3270]_ , \new_[3271]_ , \new_[3275]_ , \new_[3276]_ ,
    \new_[3280]_ , \new_[3281]_ , \new_[3282]_ , \new_[3286]_ ,
    \new_[3287]_ , \new_[3291]_ , \new_[3292]_ , \new_[3293]_ ,
    \new_[3294]_ , \new_[3298]_ , \new_[3299]_ , \new_[3303]_ ,
    \new_[3304]_ , \new_[3305]_ , \new_[3309]_ , \new_[3310]_ ,
    \new_[3313]_ , \new_[3316]_ , \new_[3317]_ , \new_[3318]_ ,
    \new_[3319]_ , \new_[3320]_ , \new_[3324]_ , \new_[3325]_ ,
    \new_[3329]_ , \new_[3330]_ , \new_[3331]_ , \new_[3335]_ ,
    \new_[3336]_ , \new_[3340]_ , \new_[3341]_ , \new_[3342]_ ,
    \new_[3343]_ , \new_[3347]_ , \new_[3348]_ , \new_[3352]_ ,
    \new_[3353]_ , \new_[3354]_ , \new_[3358]_ , \new_[3359]_ ,
    \new_[3362]_ , \new_[3365]_ , \new_[3366]_ , \new_[3367]_ ,
    \new_[3368]_ , \new_[3369]_ , \new_[3370]_ , \new_[3371]_ ,
    \new_[3375]_ , \new_[3376]_ , \new_[3380]_ , \new_[3381]_ ,
    \new_[3382]_ , \new_[3386]_ , \new_[3387]_ , \new_[3391]_ ,
    \new_[3392]_ , \new_[3393]_ , \new_[3394]_ , \new_[3398]_ ,
    \new_[3399]_ , \new_[3403]_ , \new_[3404]_ , \new_[3405]_ ,
    \new_[3409]_ , \new_[3410]_ , \new_[3414]_ , \new_[3415]_ ,
    \new_[3416]_ , \new_[3417]_ , \new_[3418]_ , \new_[3422]_ ,
    \new_[3423]_ , \new_[3427]_ , \new_[3428]_ , \new_[3429]_ ,
    \new_[3433]_ , \new_[3434]_ , \new_[3438]_ , \new_[3439]_ ,
    \new_[3440]_ , \new_[3441]_ , \new_[3445]_ , \new_[3446]_ ,
    \new_[3450]_ , \new_[3451]_ , \new_[3452]_ , \new_[3456]_ ,
    \new_[3457]_ , \new_[3460]_ , \new_[3463]_ , \new_[3464]_ ,
    \new_[3465]_ , \new_[3466]_ , \new_[3467]_ , \new_[3468]_ ,
    \new_[3472]_ , \new_[3473]_ , \new_[3477]_ , \new_[3478]_ ,
    \new_[3479]_ , \new_[3483]_ , \new_[3484]_ , \new_[3488]_ ,
    \new_[3489]_ , \new_[3490]_ , \new_[3491]_ , \new_[3495]_ ,
    \new_[3496]_ , \new_[3500]_ , \new_[3501]_ , \new_[3502]_ ,
    \new_[3506]_ , \new_[3507]_ , \new_[3510]_ , \new_[3513]_ ,
    \new_[3514]_ , \new_[3515]_ , \new_[3516]_ , \new_[3517]_ ,
    \new_[3521]_ , \new_[3522]_ , \new_[3526]_ , \new_[3527]_ ,
    \new_[3528]_ , \new_[3532]_ , \new_[3533]_ , \new_[3537]_ ,
    \new_[3538]_ , \new_[3539]_ , \new_[3540]_ , \new_[3544]_ ,
    \new_[3545]_ , \new_[3549]_ , \new_[3550]_ , \new_[3551]_ ,
    \new_[3555]_ , \new_[3556]_ , \new_[3559]_ , \new_[3562]_ ,
    \new_[3563]_ , \new_[3564]_ , \new_[3565]_ , \new_[3566]_ ,
    \new_[3567]_ , \new_[3568]_ , \new_[3569]_ , \new_[3573]_ ,
    \new_[3574]_ , \new_[3578]_ , \new_[3579]_ , \new_[3580]_ ,
    \new_[3584]_ , \new_[3585]_ , \new_[3589]_ , \new_[3590]_ ,
    \new_[3591]_ , \new_[3592]_ , \new_[3596]_ , \new_[3597]_ ,
    \new_[3601]_ , \new_[3602]_ , \new_[3603]_ , \new_[3607]_ ,
    \new_[3608]_ , \new_[3612]_ , \new_[3613]_ , \new_[3614]_ ,
    \new_[3615]_ , \new_[3616]_ , \new_[3620]_ , \new_[3621]_ ,
    \new_[3625]_ , \new_[3626]_ , \new_[3627]_ , \new_[3631]_ ,
    \new_[3632]_ , \new_[3636]_ , \new_[3637]_ , \new_[3638]_ ,
    \new_[3639]_ , \new_[3643]_ , \new_[3644]_ , \new_[3648]_ ,
    \new_[3649]_ , \new_[3650]_ , \new_[3654]_ , \new_[3655]_ ,
    \new_[3658]_ , \new_[3661]_ , \new_[3662]_ , \new_[3663]_ ,
    \new_[3664]_ , \new_[3665]_ , \new_[3666]_ , \new_[3670]_ ,
    \new_[3671]_ , \new_[3675]_ , \new_[3676]_ , \new_[3677]_ ,
    \new_[3681]_ , \new_[3682]_ , \new_[3686]_ , \new_[3687]_ ,
    \new_[3688]_ , \new_[3689]_ , \new_[3693]_ , \new_[3694]_ ,
    \new_[3698]_ , \new_[3699]_ , \new_[3700]_ , \new_[3704]_ ,
    \new_[3705]_ , \new_[3708]_ , \new_[3711]_ , \new_[3712]_ ,
    \new_[3713]_ , \new_[3714]_ , \new_[3715]_ , \new_[3719]_ ,
    \new_[3720]_ , \new_[3724]_ , \new_[3725]_ , \new_[3726]_ ,
    \new_[3730]_ , \new_[3731]_ , \new_[3735]_ , \new_[3736]_ ,
    \new_[3737]_ , \new_[3738]_ , \new_[3742]_ , \new_[3743]_ ,
    \new_[3747]_ , \new_[3748]_ , \new_[3749]_ , \new_[3753]_ ,
    \new_[3754]_ , \new_[3757]_ , \new_[3760]_ , \new_[3761]_ ,
    \new_[3762]_ , \new_[3763]_ , \new_[3764]_ , \new_[3765]_ ,
    \new_[3766]_ , \new_[3770]_ , \new_[3771]_ , \new_[3775]_ ,
    \new_[3776]_ , \new_[3777]_ , \new_[3781]_ , \new_[3782]_ ,
    \new_[3786]_ , \new_[3787]_ , \new_[3788]_ , \new_[3789]_ ,
    \new_[3793]_ , \new_[3794]_ , \new_[3798]_ , \new_[3799]_ ,
    \new_[3800]_ , \new_[3804]_ , \new_[3805]_ , \new_[3809]_ ,
    \new_[3810]_ , \new_[3811]_ , \new_[3812]_ , \new_[3813]_ ,
    \new_[3817]_ , \new_[3818]_ , \new_[3822]_ , \new_[3823]_ ,
    \new_[3824]_ , \new_[3828]_ , \new_[3829]_ , \new_[3833]_ ,
    \new_[3834]_ , \new_[3835]_ , \new_[3836]_ , \new_[3840]_ ,
    \new_[3841]_ , \new_[3845]_ , \new_[3846]_ , \new_[3847]_ ,
    \new_[3851]_ , \new_[3852]_ , \new_[3855]_ , \new_[3858]_ ,
    \new_[3859]_ , \new_[3860]_ , \new_[3861]_ , \new_[3862]_ ,
    \new_[3863]_ , \new_[3867]_ , \new_[3868]_ , \new_[3872]_ ,
    \new_[3873]_ , \new_[3874]_ , \new_[3878]_ , \new_[3879]_ ,
    \new_[3883]_ , \new_[3884]_ , \new_[3885]_ , \new_[3886]_ ,
    \new_[3890]_ , \new_[3891]_ , \new_[3895]_ , \new_[3896]_ ,
    \new_[3897]_ , \new_[3901]_ , \new_[3902]_ , \new_[3905]_ ,
    \new_[3908]_ , \new_[3909]_ , \new_[3910]_ , \new_[3911]_ ,
    \new_[3912]_ , \new_[3916]_ , \new_[3917]_ , \new_[3921]_ ,
    \new_[3922]_ , \new_[3923]_ , \new_[3927]_ , \new_[3928]_ ,
    \new_[3932]_ , \new_[3933]_ , \new_[3934]_ , \new_[3935]_ ,
    \new_[3939]_ , \new_[3940]_ , \new_[3944]_ , \new_[3945]_ ,
    \new_[3946]_ , \new_[3950]_ , \new_[3951]_ , \new_[3954]_ ,
    \new_[3957]_ , \new_[3958]_ , \new_[3959]_ , \new_[3960]_ ,
    \new_[3961]_ , \new_[3962]_ , \new_[3963]_ , \new_[3964]_ ,
    \new_[3965]_ , \new_[3969]_ , \new_[3970]_ , \new_[3974]_ ,
    \new_[3975]_ , \new_[3976]_ , \new_[3980]_ , \new_[3981]_ ,
    \new_[3985]_ , \new_[3986]_ , \new_[3987]_ , \new_[3988]_ ,
    \new_[3992]_ , \new_[3993]_ , \new_[3997]_ , \new_[3998]_ ,
    \new_[3999]_ , \new_[4003]_ , \new_[4004]_ , \new_[4008]_ ,
    \new_[4009]_ , \new_[4010]_ , \new_[4011]_ , \new_[4012]_ ,
    \new_[4016]_ , \new_[4017]_ , \new_[4021]_ , \new_[4022]_ ,
    \new_[4023]_ , \new_[4027]_ , \new_[4028]_ , \new_[4032]_ ,
    \new_[4033]_ , \new_[4034]_ , \new_[4035]_ , \new_[4039]_ ,
    \new_[4040]_ , \new_[4044]_ , \new_[4045]_ , \new_[4046]_ ,
    \new_[4050]_ , \new_[4051]_ , \new_[4054]_ , \new_[4057]_ ,
    \new_[4058]_ , \new_[4059]_ , \new_[4060]_ , \new_[4061]_ ,
    \new_[4062]_ , \new_[4066]_ , \new_[4067]_ , \new_[4071]_ ,
    \new_[4072]_ , \new_[4073]_ , \new_[4077]_ , \new_[4078]_ ,
    \new_[4082]_ , \new_[4083]_ , \new_[4084]_ , \new_[4085]_ ,
    \new_[4089]_ , \new_[4090]_ , \new_[4094]_ , \new_[4095]_ ,
    \new_[4096]_ , \new_[4100]_ , \new_[4101]_ , \new_[4104]_ ,
    \new_[4107]_ , \new_[4108]_ , \new_[4109]_ , \new_[4110]_ ,
    \new_[4111]_ , \new_[4115]_ , \new_[4116]_ , \new_[4120]_ ,
    \new_[4121]_ , \new_[4122]_ , \new_[4126]_ , \new_[4127]_ ,
    \new_[4131]_ , \new_[4132]_ , \new_[4133]_ , \new_[4134]_ ,
    \new_[4138]_ , \new_[4139]_ , \new_[4143]_ , \new_[4144]_ ,
    \new_[4145]_ , \new_[4149]_ , \new_[4150]_ , \new_[4153]_ ,
    \new_[4156]_ , \new_[4157]_ , \new_[4158]_ , \new_[4159]_ ,
    \new_[4160]_ , \new_[4161]_ , \new_[4162]_ , \new_[4166]_ ,
    \new_[4167]_ , \new_[4171]_ , \new_[4172]_ , \new_[4173]_ ,
    \new_[4177]_ , \new_[4178]_ , \new_[4182]_ , \new_[4183]_ ,
    \new_[4184]_ , \new_[4185]_ , \new_[4189]_ , \new_[4190]_ ,
    \new_[4194]_ , \new_[4195]_ , \new_[4196]_ , \new_[4200]_ ,
    \new_[4201]_ , \new_[4205]_ , \new_[4206]_ , \new_[4207]_ ,
    \new_[4208]_ , \new_[4209]_ , \new_[4213]_ , \new_[4214]_ ,
    \new_[4218]_ , \new_[4219]_ , \new_[4220]_ , \new_[4224]_ ,
    \new_[4225]_ , \new_[4229]_ , \new_[4230]_ , \new_[4231]_ ,
    \new_[4232]_ , \new_[4236]_ , \new_[4237]_ , \new_[4241]_ ,
    \new_[4242]_ , \new_[4243]_ , \new_[4247]_ , \new_[4248]_ ,
    \new_[4251]_ , \new_[4254]_ , \new_[4255]_ , \new_[4256]_ ,
    \new_[4257]_ , \new_[4258]_ , \new_[4259]_ , \new_[4263]_ ,
    \new_[4264]_ , \new_[4268]_ , \new_[4269]_ , \new_[4270]_ ,
    \new_[4274]_ , \new_[4275]_ , \new_[4279]_ , \new_[4280]_ ,
    \new_[4281]_ , \new_[4282]_ , \new_[4286]_ , \new_[4287]_ ,
    \new_[4291]_ , \new_[4292]_ , \new_[4293]_ , \new_[4297]_ ,
    \new_[4298]_ , \new_[4301]_ , \new_[4304]_ , \new_[4305]_ ,
    \new_[4306]_ , \new_[4307]_ , \new_[4308]_ , \new_[4312]_ ,
    \new_[4313]_ , \new_[4317]_ , \new_[4318]_ , \new_[4319]_ ,
    \new_[4323]_ , \new_[4324]_ , \new_[4328]_ , \new_[4329]_ ,
    \new_[4330]_ , \new_[4331]_ , \new_[4335]_ , \new_[4336]_ ,
    \new_[4340]_ , \new_[4341]_ , \new_[4342]_ , \new_[4346]_ ,
    \new_[4347]_ , \new_[4350]_ , \new_[4353]_ , \new_[4354]_ ,
    \new_[4355]_ , \new_[4356]_ , \new_[4357]_ , \new_[4358]_ ,
    \new_[4359]_ , \new_[4360]_ , \new_[4364]_ , \new_[4365]_ ,
    \new_[4369]_ , \new_[4370]_ , \new_[4371]_ , \new_[4375]_ ,
    \new_[4376]_ , \new_[4380]_ , \new_[4381]_ , \new_[4382]_ ,
    \new_[4383]_ , \new_[4387]_ , \new_[4388]_ , \new_[4392]_ ,
    \new_[4393]_ , \new_[4394]_ , \new_[4398]_ , \new_[4399]_ ,
    \new_[4403]_ , \new_[4404]_ , \new_[4405]_ , \new_[4406]_ ,
    \new_[4407]_ , \new_[4411]_ , \new_[4412]_ , \new_[4416]_ ,
    \new_[4417]_ , \new_[4418]_ , \new_[4422]_ , \new_[4423]_ ,
    \new_[4427]_ , \new_[4428]_ , \new_[4429]_ , \new_[4430]_ ,
    \new_[4434]_ , \new_[4435]_ , \new_[4439]_ , \new_[4440]_ ,
    \new_[4441]_ , \new_[4445]_ , \new_[4446]_ , \new_[4449]_ ,
    \new_[4452]_ , \new_[4453]_ , \new_[4454]_ , \new_[4455]_ ,
    \new_[4456]_ , \new_[4457]_ , \new_[4461]_ , \new_[4462]_ ,
    \new_[4466]_ , \new_[4467]_ , \new_[4468]_ , \new_[4472]_ ,
    \new_[4473]_ , \new_[4477]_ , \new_[4478]_ , \new_[4479]_ ,
    \new_[4480]_ , \new_[4484]_ , \new_[4485]_ , \new_[4489]_ ,
    \new_[4490]_ , \new_[4491]_ , \new_[4495]_ , \new_[4496]_ ,
    \new_[4499]_ , \new_[4502]_ , \new_[4503]_ , \new_[4504]_ ,
    \new_[4505]_ , \new_[4506]_ , \new_[4510]_ , \new_[4511]_ ,
    \new_[4515]_ , \new_[4516]_ , \new_[4517]_ , \new_[4521]_ ,
    \new_[4522]_ , \new_[4526]_ , \new_[4527]_ , \new_[4528]_ ,
    \new_[4529]_ , \new_[4533]_ , \new_[4534]_ , \new_[4538]_ ,
    \new_[4539]_ , \new_[4540]_ , \new_[4544]_ , \new_[4545]_ ,
    \new_[4548]_ , \new_[4551]_ , \new_[4552]_ , \new_[4553]_ ,
    \new_[4554]_ , \new_[4555]_ , \new_[4556]_ , \new_[4557]_ ,
    \new_[4561]_ , \new_[4562]_ , \new_[4566]_ , \new_[4567]_ ,
    \new_[4568]_ , \new_[4572]_ , \new_[4573]_ , \new_[4577]_ ,
    \new_[4578]_ , \new_[4579]_ , \new_[4580]_ , \new_[4584]_ ,
    \new_[4585]_ , \new_[4589]_ , \new_[4590]_ , \new_[4591]_ ,
    \new_[4595]_ , \new_[4596]_ , \new_[4599]_ , \new_[4602]_ ,
    \new_[4603]_ , \new_[4604]_ , \new_[4605]_ , \new_[4606]_ ,
    \new_[4610]_ , \new_[4611]_ , \new_[4615]_ , \new_[4616]_ ,
    \new_[4617]_ , \new_[4621]_ , \new_[4622]_ , \new_[4626]_ ,
    \new_[4627]_ , \new_[4628]_ , \new_[4629]_ , \new_[4633]_ ,
    \new_[4634]_ , \new_[4638]_ , \new_[4639]_ , \new_[4640]_ ,
    \new_[4644]_ , \new_[4645]_ , \new_[4648]_ , \new_[4651]_ ,
    \new_[4652]_ , \new_[4653]_ , \new_[4654]_ , \new_[4655]_ ,
    \new_[4656]_ , \new_[4660]_ , \new_[4661]_ , \new_[4665]_ ,
    \new_[4666]_ , \new_[4667]_ , \new_[4671]_ , \new_[4672]_ ,
    \new_[4676]_ , \new_[4677]_ , \new_[4678]_ , \new_[4679]_ ,
    \new_[4683]_ , \new_[4684]_ , \new_[4688]_ , \new_[4689]_ ,
    \new_[4690]_ , \new_[4694]_ , \new_[4695]_ , \new_[4698]_ ,
    \new_[4701]_ , \new_[4702]_ , \new_[4703]_ , \new_[4704]_ ,
    \new_[4705]_ , \new_[4709]_ , \new_[4710]_ , \new_[4714]_ ,
    \new_[4715]_ , \new_[4716]_ , \new_[4720]_ , \new_[4721]_ ,
    \new_[4725]_ , \new_[4726]_ , \new_[4727]_ , \new_[4728]_ ,
    \new_[4732]_ , \new_[4733]_ , \new_[4737]_ , \new_[4738]_ ,
    \new_[4739]_ , \new_[4743]_ , \new_[4744]_ , \new_[4747]_ ,
    \new_[4750]_ , \new_[4751]_ , \new_[4752]_ , \new_[4753]_ ,
    \new_[4754]_ , \new_[4755]_ , \new_[4756]_ , \new_[4757]_ ,
    \new_[4758]_ , \new_[4759]_ , \new_[4763]_ , \new_[4764]_ ,
    \new_[4768]_ , \new_[4769]_ , \new_[4770]_ , \new_[4774]_ ,
    \new_[4775]_ , \new_[4779]_ , \new_[4780]_ , \new_[4781]_ ,
    \new_[4782]_ , \new_[4786]_ , \new_[4787]_ , \new_[4791]_ ,
    \new_[4792]_ , \new_[4793]_ , \new_[4797]_ , \new_[4798]_ ,
    \new_[4802]_ , \new_[4803]_ , \new_[4804]_ , \new_[4805]_ ,
    \new_[4806]_ , \new_[4810]_ , \new_[4811]_ , \new_[4815]_ ,
    \new_[4816]_ , \new_[4817]_ , \new_[4821]_ , \new_[4822]_ ,
    \new_[4826]_ , \new_[4827]_ , \new_[4828]_ , \new_[4829]_ ,
    \new_[4833]_ , \new_[4834]_ , \new_[4838]_ , \new_[4839]_ ,
    \new_[4840]_ , \new_[4844]_ , \new_[4845]_ , \new_[4848]_ ,
    \new_[4851]_ , \new_[4852]_ , \new_[4853]_ , \new_[4854]_ ,
    \new_[4855]_ , \new_[4856]_ , \new_[4860]_ , \new_[4861]_ ,
    \new_[4865]_ , \new_[4866]_ , \new_[4867]_ , \new_[4871]_ ,
    \new_[4872]_ , \new_[4876]_ , \new_[4877]_ , \new_[4878]_ ,
    \new_[4879]_ , \new_[4883]_ , \new_[4884]_ , \new_[4888]_ ,
    \new_[4889]_ , \new_[4890]_ , \new_[4894]_ , \new_[4895]_ ,
    \new_[4898]_ , \new_[4901]_ , \new_[4902]_ , \new_[4903]_ ,
    \new_[4904]_ , \new_[4905]_ , \new_[4909]_ , \new_[4910]_ ,
    \new_[4914]_ , \new_[4915]_ , \new_[4916]_ , \new_[4920]_ ,
    \new_[4921]_ , \new_[4925]_ , \new_[4926]_ , \new_[4927]_ ,
    \new_[4928]_ , \new_[4932]_ , \new_[4933]_ , \new_[4937]_ ,
    \new_[4938]_ , \new_[4939]_ , \new_[4943]_ , \new_[4944]_ ,
    \new_[4947]_ , \new_[4950]_ , \new_[4951]_ , \new_[4952]_ ,
    \new_[4953]_ , \new_[4954]_ , \new_[4955]_ , \new_[4956]_ ,
    \new_[4960]_ , \new_[4961]_ , \new_[4965]_ , \new_[4966]_ ,
    \new_[4967]_ , \new_[4971]_ , \new_[4972]_ , \new_[4976]_ ,
    \new_[4977]_ , \new_[4978]_ , \new_[4979]_ , \new_[4983]_ ,
    \new_[4984]_ , \new_[4988]_ , \new_[4989]_ , \new_[4990]_ ,
    \new_[4994]_ , \new_[4995]_ , \new_[4999]_ , \new_[5000]_ ,
    \new_[5001]_ , \new_[5002]_ , \new_[5003]_ , \new_[5007]_ ,
    \new_[5008]_ , \new_[5012]_ , \new_[5013]_ , \new_[5014]_ ,
    \new_[5018]_ , \new_[5019]_ , \new_[5023]_ , \new_[5024]_ ,
    \new_[5025]_ , \new_[5026]_ , \new_[5030]_ , \new_[5031]_ ,
    \new_[5035]_ , \new_[5036]_ , \new_[5037]_ , \new_[5041]_ ,
    \new_[5042]_ , \new_[5045]_ , \new_[5048]_ , \new_[5049]_ ,
    \new_[5050]_ , \new_[5051]_ , \new_[5052]_ , \new_[5053]_ ,
    \new_[5057]_ , \new_[5058]_ , \new_[5062]_ , \new_[5063]_ ,
    \new_[5064]_ , \new_[5068]_ , \new_[5069]_ , \new_[5073]_ ,
    \new_[5074]_ , \new_[5075]_ , \new_[5076]_ , \new_[5080]_ ,
    \new_[5081]_ , \new_[5085]_ , \new_[5086]_ , \new_[5087]_ ,
    \new_[5091]_ , \new_[5092]_ , \new_[5095]_ , \new_[5098]_ ,
    \new_[5099]_ , \new_[5100]_ , \new_[5101]_ , \new_[5102]_ ,
    \new_[5106]_ , \new_[5107]_ , \new_[5111]_ , \new_[5112]_ ,
    \new_[5113]_ , \new_[5117]_ , \new_[5118]_ , \new_[5122]_ ,
    \new_[5123]_ , \new_[5124]_ , \new_[5125]_ , \new_[5129]_ ,
    \new_[5130]_ , \new_[5134]_ , \new_[5135]_ , \new_[5136]_ ,
    \new_[5140]_ , \new_[5141]_ , \new_[5144]_ , \new_[5147]_ ,
    \new_[5148]_ , \new_[5149]_ , \new_[5150]_ , \new_[5151]_ ,
    \new_[5152]_ , \new_[5153]_ , \new_[5154]_ , \new_[5158]_ ,
    \new_[5159]_ , \new_[5163]_ , \new_[5164]_ , \new_[5165]_ ,
    \new_[5169]_ , \new_[5170]_ , \new_[5174]_ , \new_[5175]_ ,
    \new_[5176]_ , \new_[5177]_ , \new_[5181]_ , \new_[5182]_ ,
    \new_[5186]_ , \new_[5187]_ , \new_[5188]_ , \new_[5192]_ ,
    \new_[5193]_ , \new_[5197]_ , \new_[5198]_ , \new_[5199]_ ,
    \new_[5200]_ , \new_[5201]_ , \new_[5205]_ , \new_[5206]_ ,
    \new_[5210]_ , \new_[5211]_ , \new_[5212]_ , \new_[5216]_ ,
    \new_[5217]_ , \new_[5221]_ , \new_[5222]_ , \new_[5223]_ ,
    \new_[5224]_ , \new_[5228]_ , \new_[5229]_ , \new_[5233]_ ,
    \new_[5234]_ , \new_[5235]_ , \new_[5239]_ , \new_[5240]_ ,
    \new_[5243]_ , \new_[5246]_ , \new_[5247]_ , \new_[5248]_ ,
    \new_[5249]_ , \new_[5250]_ , \new_[5251]_ , \new_[5255]_ ,
    \new_[5256]_ , \new_[5260]_ , \new_[5261]_ , \new_[5262]_ ,
    \new_[5266]_ , \new_[5267]_ , \new_[5271]_ , \new_[5272]_ ,
    \new_[5273]_ , \new_[5274]_ , \new_[5278]_ , \new_[5279]_ ,
    \new_[5283]_ , \new_[5284]_ , \new_[5285]_ , \new_[5289]_ ,
    \new_[5290]_ , \new_[5293]_ , \new_[5296]_ , \new_[5297]_ ,
    \new_[5298]_ , \new_[5299]_ , \new_[5300]_ , \new_[5304]_ ,
    \new_[5305]_ , \new_[5309]_ , \new_[5310]_ , \new_[5311]_ ,
    \new_[5315]_ , \new_[5316]_ , \new_[5320]_ , \new_[5321]_ ,
    \new_[5322]_ , \new_[5323]_ , \new_[5327]_ , \new_[5328]_ ,
    \new_[5332]_ , \new_[5333]_ , \new_[5334]_ , \new_[5338]_ ,
    \new_[5339]_ , \new_[5342]_ , \new_[5345]_ , \new_[5346]_ ,
    \new_[5347]_ , \new_[5348]_ , \new_[5349]_ , \new_[5350]_ ,
    \new_[5351]_ , \new_[5355]_ , \new_[5356]_ , \new_[5360]_ ,
    \new_[5361]_ , \new_[5362]_ , \new_[5366]_ , \new_[5367]_ ,
    \new_[5371]_ , \new_[5372]_ , \new_[5373]_ , \new_[5374]_ ,
    \new_[5378]_ , \new_[5379]_ , \new_[5383]_ , \new_[5384]_ ,
    \new_[5385]_ , \new_[5389]_ , \new_[5390]_ , \new_[5393]_ ,
    \new_[5396]_ , \new_[5397]_ , \new_[5398]_ , \new_[5399]_ ,
    \new_[5400]_ , \new_[5404]_ , \new_[5405]_ , \new_[5409]_ ,
    \new_[5410]_ , \new_[5411]_ , \new_[5415]_ , \new_[5416]_ ,
    \new_[5420]_ , \new_[5421]_ , \new_[5422]_ , \new_[5423]_ ,
    \new_[5427]_ , \new_[5428]_ , \new_[5432]_ , \new_[5433]_ ,
    \new_[5434]_ , \new_[5438]_ , \new_[5439]_ , \new_[5442]_ ,
    \new_[5445]_ , \new_[5446]_ , \new_[5447]_ , \new_[5448]_ ,
    \new_[5449]_ , \new_[5450]_ , \new_[5454]_ , \new_[5455]_ ,
    \new_[5459]_ , \new_[5460]_ , \new_[5461]_ , \new_[5465]_ ,
    \new_[5466]_ , \new_[5470]_ , \new_[5471]_ , \new_[5472]_ ,
    \new_[5473]_ , \new_[5477]_ , \new_[5478]_ , \new_[5482]_ ,
    \new_[5483]_ , \new_[5484]_ , \new_[5488]_ , \new_[5489]_ ,
    \new_[5492]_ , \new_[5495]_ , \new_[5496]_ , \new_[5497]_ ,
    \new_[5498]_ , \new_[5499]_ , \new_[5503]_ , \new_[5504]_ ,
    \new_[5508]_ , \new_[5509]_ , \new_[5510]_ , \new_[5514]_ ,
    \new_[5515]_ , \new_[5519]_ , \new_[5520]_ , \new_[5521]_ ,
    \new_[5522]_ , \new_[5526]_ , \new_[5527]_ , \new_[5531]_ ,
    \new_[5532]_ , \new_[5533]_ , \new_[5537]_ , \new_[5538]_ ,
    \new_[5541]_ , \new_[5544]_ , \new_[5545]_ , \new_[5546]_ ,
    \new_[5547]_ , \new_[5548]_ , \new_[5549]_ , \new_[5550]_ ,
    \new_[5551]_ , \new_[5552]_ , \new_[5556]_ , \new_[5557]_ ,
    \new_[5561]_ , \new_[5562]_ , \new_[5563]_ , \new_[5567]_ ,
    \new_[5568]_ , \new_[5572]_ , \new_[5573]_ , \new_[5574]_ ,
    \new_[5575]_ , \new_[5579]_ , \new_[5580]_ , \new_[5584]_ ,
    \new_[5585]_ , \new_[5586]_ , \new_[5590]_ , \new_[5591]_ ,
    \new_[5595]_ , \new_[5596]_ , \new_[5597]_ , \new_[5598]_ ,
    \new_[5599]_ , \new_[5603]_ , \new_[5604]_ , \new_[5608]_ ,
    \new_[5609]_ , \new_[5610]_ , \new_[5614]_ , \new_[5615]_ ,
    \new_[5619]_ , \new_[5620]_ , \new_[5621]_ , \new_[5622]_ ,
    \new_[5626]_ , \new_[5627]_ , \new_[5631]_ , \new_[5632]_ ,
    \new_[5633]_ , \new_[5637]_ , \new_[5638]_ , \new_[5641]_ ,
    \new_[5644]_ , \new_[5645]_ , \new_[5646]_ , \new_[5647]_ ,
    \new_[5648]_ , \new_[5649]_ , \new_[5653]_ , \new_[5654]_ ,
    \new_[5658]_ , \new_[5659]_ , \new_[5660]_ , \new_[5664]_ ,
    \new_[5665]_ , \new_[5669]_ , \new_[5670]_ , \new_[5671]_ ,
    \new_[5672]_ , \new_[5676]_ , \new_[5677]_ , \new_[5681]_ ,
    \new_[5682]_ , \new_[5683]_ , \new_[5687]_ , \new_[5688]_ ,
    \new_[5691]_ , \new_[5694]_ , \new_[5695]_ , \new_[5696]_ ,
    \new_[5697]_ , \new_[5698]_ , \new_[5702]_ , \new_[5703]_ ,
    \new_[5707]_ , \new_[5708]_ , \new_[5709]_ , \new_[5713]_ ,
    \new_[5714]_ , \new_[5718]_ , \new_[5719]_ , \new_[5720]_ ,
    \new_[5721]_ , \new_[5725]_ , \new_[5726]_ , \new_[5730]_ ,
    \new_[5731]_ , \new_[5732]_ , \new_[5736]_ , \new_[5737]_ ,
    \new_[5740]_ , \new_[5743]_ , \new_[5744]_ , \new_[5745]_ ,
    \new_[5746]_ , \new_[5747]_ , \new_[5748]_ , \new_[5749]_ ,
    \new_[5753]_ , \new_[5754]_ , \new_[5758]_ , \new_[5759]_ ,
    \new_[5760]_ , \new_[5764]_ , \new_[5765]_ , \new_[5769]_ ,
    \new_[5770]_ , \new_[5771]_ , \new_[5772]_ , \new_[5776]_ ,
    \new_[5777]_ , \new_[5781]_ , \new_[5782]_ , \new_[5783]_ ,
    \new_[5787]_ , \new_[5788]_ , \new_[5792]_ , \new_[5793]_ ,
    \new_[5794]_ , \new_[5795]_ , \new_[5796]_ , \new_[5800]_ ,
    \new_[5801]_ , \new_[5805]_ , \new_[5806]_ , \new_[5807]_ ,
    \new_[5811]_ , \new_[5812]_ , \new_[5816]_ , \new_[5817]_ ,
    \new_[5818]_ , \new_[5819]_ , \new_[5823]_ , \new_[5824]_ ,
    \new_[5828]_ , \new_[5829]_ , \new_[5830]_ , \new_[5834]_ ,
    \new_[5835]_ , \new_[5838]_ , \new_[5841]_ , \new_[5842]_ ,
    \new_[5843]_ , \new_[5844]_ , \new_[5845]_ , \new_[5846]_ ,
    \new_[5850]_ , \new_[5851]_ , \new_[5855]_ , \new_[5856]_ ,
    \new_[5857]_ , \new_[5861]_ , \new_[5862]_ , \new_[5866]_ ,
    \new_[5867]_ , \new_[5868]_ , \new_[5869]_ , \new_[5873]_ ,
    \new_[5874]_ , \new_[5878]_ , \new_[5879]_ , \new_[5880]_ ,
    \new_[5884]_ , \new_[5885]_ , \new_[5888]_ , \new_[5891]_ ,
    \new_[5892]_ , \new_[5893]_ , \new_[5894]_ , \new_[5895]_ ,
    \new_[5899]_ , \new_[5900]_ , \new_[5904]_ , \new_[5905]_ ,
    \new_[5906]_ , \new_[5910]_ , \new_[5911]_ , \new_[5915]_ ,
    \new_[5916]_ , \new_[5917]_ , \new_[5918]_ , \new_[5922]_ ,
    \new_[5923]_ , \new_[5927]_ , \new_[5928]_ , \new_[5929]_ ,
    \new_[5933]_ , \new_[5934]_ , \new_[5937]_ , \new_[5940]_ ,
    \new_[5941]_ , \new_[5942]_ , \new_[5943]_ , \new_[5944]_ ,
    \new_[5945]_ , \new_[5946]_ , \new_[5947]_ , \new_[5951]_ ,
    \new_[5952]_ , \new_[5956]_ , \new_[5957]_ , \new_[5958]_ ,
    \new_[5962]_ , \new_[5963]_ , \new_[5967]_ , \new_[5968]_ ,
    \new_[5969]_ , \new_[5970]_ , \new_[5974]_ , \new_[5975]_ ,
    \new_[5979]_ , \new_[5980]_ , \new_[5981]_ , \new_[5985]_ ,
    \new_[5986]_ , \new_[5990]_ , \new_[5991]_ , \new_[5992]_ ,
    \new_[5993]_ , \new_[5994]_ , \new_[5998]_ , \new_[5999]_ ,
    \new_[6003]_ , \new_[6004]_ , \new_[6005]_ , \new_[6009]_ ,
    \new_[6010]_ , \new_[6014]_ , \new_[6015]_ , \new_[6016]_ ,
    \new_[6017]_ , \new_[6021]_ , \new_[6022]_ , \new_[6026]_ ,
    \new_[6027]_ , \new_[6028]_ , \new_[6032]_ , \new_[6033]_ ,
    \new_[6036]_ , \new_[6039]_ , \new_[6040]_ , \new_[6041]_ ,
    \new_[6042]_ , \new_[6043]_ , \new_[6044]_ , \new_[6048]_ ,
    \new_[6049]_ , \new_[6053]_ , \new_[6054]_ , \new_[6055]_ ,
    \new_[6059]_ , \new_[6060]_ , \new_[6064]_ , \new_[6065]_ ,
    \new_[6066]_ , \new_[6067]_ , \new_[6071]_ , \new_[6072]_ ,
    \new_[6076]_ , \new_[6077]_ , \new_[6078]_ , \new_[6082]_ ,
    \new_[6083]_ , \new_[6086]_ , \new_[6089]_ , \new_[6090]_ ,
    \new_[6091]_ , \new_[6092]_ , \new_[6093]_ , \new_[6097]_ ,
    \new_[6098]_ , \new_[6102]_ , \new_[6103]_ , \new_[6104]_ ,
    \new_[6108]_ , \new_[6109]_ , \new_[6113]_ , \new_[6114]_ ,
    \new_[6115]_ , \new_[6116]_ , \new_[6120]_ , \new_[6121]_ ,
    \new_[6125]_ , \new_[6126]_ , \new_[6127]_ , \new_[6131]_ ,
    \new_[6132]_ , \new_[6135]_ , \new_[6138]_ , \new_[6139]_ ,
    \new_[6140]_ , \new_[6141]_ , \new_[6142]_ , \new_[6143]_ ,
    \new_[6144]_ , \new_[6148]_ , \new_[6149]_ , \new_[6153]_ ,
    \new_[6154]_ , \new_[6155]_ , \new_[6159]_ , \new_[6160]_ ,
    \new_[6164]_ , \new_[6165]_ , \new_[6166]_ , \new_[6167]_ ,
    \new_[6171]_ , \new_[6172]_ , \new_[6176]_ , \new_[6177]_ ,
    \new_[6178]_ , \new_[6182]_ , \new_[6183]_ , \new_[6186]_ ,
    \new_[6189]_ , \new_[6190]_ , \new_[6191]_ , \new_[6192]_ ,
    \new_[6193]_ , \new_[6197]_ , \new_[6198]_ , \new_[6202]_ ,
    \new_[6203]_ , \new_[6204]_ , \new_[6208]_ , \new_[6209]_ ,
    \new_[6213]_ , \new_[6214]_ , \new_[6215]_ , \new_[6216]_ ,
    \new_[6220]_ , \new_[6221]_ , \new_[6225]_ , \new_[6226]_ ,
    \new_[6227]_ , \new_[6231]_ , \new_[6232]_ , \new_[6235]_ ,
    \new_[6238]_ , \new_[6239]_ , \new_[6240]_ , \new_[6241]_ ,
    \new_[6242]_ , \new_[6243]_ , \new_[6247]_ , \new_[6248]_ ,
    \new_[6252]_ , \new_[6253]_ , \new_[6254]_ , \new_[6258]_ ,
    \new_[6259]_ , \new_[6263]_ , \new_[6264]_ , \new_[6265]_ ,
    \new_[6266]_ , \new_[6270]_ , \new_[6271]_ , \new_[6275]_ ,
    \new_[6276]_ , \new_[6277]_ , \new_[6281]_ , \new_[6282]_ ,
    \new_[6285]_ , \new_[6288]_ , \new_[6289]_ , \new_[6290]_ ,
    \new_[6291]_ , \new_[6292]_ , \new_[6296]_ , \new_[6297]_ ,
    \new_[6301]_ , \new_[6302]_ , \new_[6303]_ , \new_[6307]_ ,
    \new_[6308]_ , \new_[6312]_ , \new_[6313]_ , \new_[6314]_ ,
    \new_[6315]_ , \new_[6319]_ , \new_[6320]_ , \new_[6324]_ ,
    \new_[6325]_ , \new_[6326]_ , \new_[6330]_ , \new_[6331]_ ,
    \new_[6334]_ , \new_[6337]_ , \new_[6338]_ , \new_[6339]_ ,
    \new_[6340]_ , \new_[6341]_ , \new_[6342]_ , \new_[6343]_ ,
    \new_[6344]_ , \new_[6345]_ , \new_[6346]_ , \new_[6347]_ ,
    \new_[6351]_ , \new_[6352]_ , \new_[6356]_ , \new_[6357]_ ,
    \new_[6358]_ , \new_[6362]_ , \new_[6363]_ , \new_[6367]_ ,
    \new_[6368]_ , \new_[6369]_ , \new_[6370]_ , \new_[6374]_ ,
    \new_[6375]_ , \new_[6379]_ , \new_[6380]_ , \new_[6381]_ ,
    \new_[6385]_ , \new_[6386]_ , \new_[6390]_ , \new_[6391]_ ,
    \new_[6392]_ , \new_[6393]_ , \new_[6394]_ , \new_[6398]_ ,
    \new_[6399]_ , \new_[6403]_ , \new_[6404]_ , \new_[6405]_ ,
    \new_[6409]_ , \new_[6410]_ , \new_[6414]_ , \new_[6415]_ ,
    \new_[6416]_ , \new_[6417]_ , \new_[6421]_ , \new_[6422]_ ,
    \new_[6426]_ , \new_[6427]_ , \new_[6428]_ , \new_[6432]_ ,
    \new_[6433]_ , \new_[6436]_ , \new_[6439]_ , \new_[6440]_ ,
    \new_[6441]_ , \new_[6442]_ , \new_[6443]_ , \new_[6444]_ ,
    \new_[6448]_ , \new_[6449]_ , \new_[6453]_ , \new_[6454]_ ,
    \new_[6455]_ , \new_[6459]_ , \new_[6460]_ , \new_[6464]_ ,
    \new_[6465]_ , \new_[6466]_ , \new_[6467]_ , \new_[6471]_ ,
    \new_[6472]_ , \new_[6476]_ , \new_[6477]_ , \new_[6478]_ ,
    \new_[6482]_ , \new_[6483]_ , \new_[6486]_ , \new_[6489]_ ,
    \new_[6490]_ , \new_[6491]_ , \new_[6492]_ , \new_[6493]_ ,
    \new_[6497]_ , \new_[6498]_ , \new_[6502]_ , \new_[6503]_ ,
    \new_[6504]_ , \new_[6508]_ , \new_[6509]_ , \new_[6513]_ ,
    \new_[6514]_ , \new_[6515]_ , \new_[6516]_ , \new_[6520]_ ,
    \new_[6521]_ , \new_[6525]_ , \new_[6526]_ , \new_[6527]_ ,
    \new_[6531]_ , \new_[6532]_ , \new_[6535]_ , \new_[6538]_ ,
    \new_[6539]_ , \new_[6540]_ , \new_[6541]_ , \new_[6542]_ ,
    \new_[6543]_ , \new_[6544]_ , \new_[6548]_ , \new_[6549]_ ,
    \new_[6553]_ , \new_[6554]_ , \new_[6555]_ , \new_[6559]_ ,
    \new_[6560]_ , \new_[6564]_ , \new_[6565]_ , \new_[6566]_ ,
    \new_[6567]_ , \new_[6571]_ , \new_[6572]_ , \new_[6576]_ ,
    \new_[6577]_ , \new_[6578]_ , \new_[6582]_ , \new_[6583]_ ,
    \new_[6587]_ , \new_[6588]_ , \new_[6589]_ , \new_[6590]_ ,
    \new_[6591]_ , \new_[6595]_ , \new_[6596]_ , \new_[6600]_ ,
    \new_[6601]_ , \new_[6602]_ , \new_[6606]_ , \new_[6607]_ ,
    \new_[6611]_ , \new_[6612]_ , \new_[6613]_ , \new_[6614]_ ,
    \new_[6618]_ , \new_[6619]_ , \new_[6623]_ , \new_[6624]_ ,
    \new_[6625]_ , \new_[6629]_ , \new_[6630]_ , \new_[6633]_ ,
    \new_[6636]_ , \new_[6637]_ , \new_[6638]_ , \new_[6639]_ ,
    \new_[6640]_ , \new_[6641]_ , \new_[6645]_ , \new_[6646]_ ,
    \new_[6650]_ , \new_[6651]_ , \new_[6652]_ , \new_[6656]_ ,
    \new_[6657]_ , \new_[6661]_ , \new_[6662]_ , \new_[6663]_ ,
    \new_[6664]_ , \new_[6668]_ , \new_[6669]_ , \new_[6673]_ ,
    \new_[6674]_ , \new_[6675]_ , \new_[6679]_ , \new_[6680]_ ,
    \new_[6683]_ , \new_[6686]_ , \new_[6687]_ , \new_[6688]_ ,
    \new_[6689]_ , \new_[6690]_ , \new_[6694]_ , \new_[6695]_ ,
    \new_[6699]_ , \new_[6700]_ , \new_[6701]_ , \new_[6705]_ ,
    \new_[6706]_ , \new_[6710]_ , \new_[6711]_ , \new_[6712]_ ,
    \new_[6713]_ , \new_[6717]_ , \new_[6718]_ , \new_[6722]_ ,
    \new_[6723]_ , \new_[6724]_ , \new_[6728]_ , \new_[6729]_ ,
    \new_[6732]_ , \new_[6735]_ , \new_[6736]_ , \new_[6737]_ ,
    \new_[6738]_ , \new_[6739]_ , \new_[6740]_ , \new_[6741]_ ,
    \new_[6742]_ , \new_[6746]_ , \new_[6747]_ , \new_[6751]_ ,
    \new_[6752]_ , \new_[6753]_ , \new_[6757]_ , \new_[6758]_ ,
    \new_[6762]_ , \new_[6763]_ , \new_[6764]_ , \new_[6765]_ ,
    \new_[6769]_ , \new_[6770]_ , \new_[6774]_ , \new_[6775]_ ,
    \new_[6776]_ , \new_[6780]_ , \new_[6781]_ , \new_[6785]_ ,
    \new_[6786]_ , \new_[6787]_ , \new_[6788]_ , \new_[6789]_ ,
    \new_[6793]_ , \new_[6794]_ , \new_[6798]_ , \new_[6799]_ ,
    \new_[6800]_ , \new_[6804]_ , \new_[6805]_ , \new_[6809]_ ,
    \new_[6810]_ , \new_[6811]_ , \new_[6812]_ , \new_[6816]_ ,
    \new_[6817]_ , \new_[6821]_ , \new_[6822]_ , \new_[6823]_ ,
    \new_[6827]_ , \new_[6828]_ , \new_[6831]_ , \new_[6834]_ ,
    \new_[6835]_ , \new_[6836]_ , \new_[6837]_ , \new_[6838]_ ,
    \new_[6839]_ , \new_[6843]_ , \new_[6844]_ , \new_[6848]_ ,
    \new_[6849]_ , \new_[6850]_ , \new_[6854]_ , \new_[6855]_ ,
    \new_[6859]_ , \new_[6860]_ , \new_[6861]_ , \new_[6862]_ ,
    \new_[6866]_ , \new_[6867]_ , \new_[6871]_ , \new_[6872]_ ,
    \new_[6873]_ , \new_[6877]_ , \new_[6878]_ , \new_[6881]_ ,
    \new_[6884]_ , \new_[6885]_ , \new_[6886]_ , \new_[6887]_ ,
    \new_[6888]_ , \new_[6892]_ , \new_[6893]_ , \new_[6897]_ ,
    \new_[6898]_ , \new_[6899]_ , \new_[6903]_ , \new_[6904]_ ,
    \new_[6908]_ , \new_[6909]_ , \new_[6910]_ , \new_[6911]_ ,
    \new_[6915]_ , \new_[6916]_ , \new_[6920]_ , \new_[6921]_ ,
    \new_[6922]_ , \new_[6926]_ , \new_[6927]_ , \new_[6930]_ ,
    \new_[6933]_ , \new_[6934]_ , \new_[6935]_ , \new_[6936]_ ,
    \new_[6937]_ , \new_[6938]_ , \new_[6939]_ , \new_[6943]_ ,
    \new_[6944]_ , \new_[6948]_ , \new_[6949]_ , \new_[6950]_ ,
    \new_[6954]_ , \new_[6955]_ , \new_[6959]_ , \new_[6960]_ ,
    \new_[6961]_ , \new_[6962]_ , \new_[6966]_ , \new_[6967]_ ,
    \new_[6971]_ , \new_[6972]_ , \new_[6973]_ , \new_[6977]_ ,
    \new_[6978]_ , \new_[6982]_ , \new_[6983]_ , \new_[6984]_ ,
    \new_[6985]_ , \new_[6986]_ , \new_[6990]_ , \new_[6991]_ ,
    \new_[6995]_ , \new_[6996]_ , \new_[6997]_ , \new_[7001]_ ,
    \new_[7002]_ , \new_[7006]_ , \new_[7007]_ , \new_[7008]_ ,
    \new_[7009]_ , \new_[7013]_ , \new_[7014]_ , \new_[7018]_ ,
    \new_[7019]_ , \new_[7020]_ , \new_[7024]_ , \new_[7025]_ ,
    \new_[7028]_ , \new_[7031]_ , \new_[7032]_ , \new_[7033]_ ,
    \new_[7034]_ , \new_[7035]_ , \new_[7036]_ , \new_[7040]_ ,
    \new_[7041]_ , \new_[7045]_ , \new_[7046]_ , \new_[7047]_ ,
    \new_[7051]_ , \new_[7052]_ , \new_[7056]_ , \new_[7057]_ ,
    \new_[7058]_ , \new_[7059]_ , \new_[7063]_ , \new_[7064]_ ,
    \new_[7068]_ , \new_[7069]_ , \new_[7070]_ , \new_[7074]_ ,
    \new_[7075]_ , \new_[7078]_ , \new_[7081]_ , \new_[7082]_ ,
    \new_[7083]_ , \new_[7084]_ , \new_[7085]_ , \new_[7089]_ ,
    \new_[7090]_ , \new_[7094]_ , \new_[7095]_ , \new_[7096]_ ,
    \new_[7100]_ , \new_[7101]_ , \new_[7105]_ , \new_[7106]_ ,
    \new_[7107]_ , \new_[7108]_ , \new_[7112]_ , \new_[7113]_ ,
    \new_[7117]_ , \new_[7118]_ , \new_[7119]_ , \new_[7123]_ ,
    \new_[7124]_ , \new_[7127]_ , \new_[7130]_ , \new_[7131]_ ,
    \new_[7132]_ , \new_[7133]_ , \new_[7134]_ , \new_[7135]_ ,
    \new_[7136]_ , \new_[7137]_ , \new_[7138]_ , \new_[7142]_ ,
    \new_[7143]_ , \new_[7147]_ , \new_[7148]_ , \new_[7149]_ ,
    \new_[7153]_ , \new_[7154]_ , \new_[7158]_ , \new_[7159]_ ,
    \new_[7160]_ , \new_[7161]_ , \new_[7165]_ , \new_[7166]_ ,
    \new_[7170]_ , \new_[7171]_ , \new_[7172]_ , \new_[7176]_ ,
    \new_[7177]_ , \new_[7181]_ , \new_[7182]_ , \new_[7183]_ ,
    \new_[7184]_ , \new_[7185]_ , \new_[7189]_ , \new_[7190]_ ,
    \new_[7194]_ , \new_[7195]_ , \new_[7196]_ , \new_[7200]_ ,
    \new_[7201]_ , \new_[7205]_ , \new_[7206]_ , \new_[7207]_ ,
    \new_[7208]_ , \new_[7212]_ , \new_[7213]_ , \new_[7217]_ ,
    \new_[7218]_ , \new_[7219]_ , \new_[7223]_ , \new_[7224]_ ,
    \new_[7227]_ , \new_[7230]_ , \new_[7231]_ , \new_[7232]_ ,
    \new_[7233]_ , \new_[7234]_ , \new_[7235]_ , \new_[7239]_ ,
    \new_[7240]_ , \new_[7244]_ , \new_[7245]_ , \new_[7246]_ ,
    \new_[7250]_ , \new_[7251]_ , \new_[7255]_ , \new_[7256]_ ,
    \new_[7257]_ , \new_[7258]_ , \new_[7262]_ , \new_[7263]_ ,
    \new_[7267]_ , \new_[7268]_ , \new_[7269]_ , \new_[7273]_ ,
    \new_[7274]_ , \new_[7277]_ , \new_[7280]_ , \new_[7281]_ ,
    \new_[7282]_ , \new_[7283]_ , \new_[7284]_ , \new_[7288]_ ,
    \new_[7289]_ , \new_[7293]_ , \new_[7294]_ , \new_[7295]_ ,
    \new_[7299]_ , \new_[7300]_ , \new_[7304]_ , \new_[7305]_ ,
    \new_[7306]_ , \new_[7307]_ , \new_[7311]_ , \new_[7312]_ ,
    \new_[7316]_ , \new_[7317]_ , \new_[7318]_ , \new_[7322]_ ,
    \new_[7323]_ , \new_[7326]_ , \new_[7329]_ , \new_[7330]_ ,
    \new_[7331]_ , \new_[7332]_ , \new_[7333]_ , \new_[7334]_ ,
    \new_[7335]_ , \new_[7339]_ , \new_[7340]_ , \new_[7344]_ ,
    \new_[7345]_ , \new_[7346]_ , \new_[7350]_ , \new_[7351]_ ,
    \new_[7355]_ , \new_[7356]_ , \new_[7357]_ , \new_[7358]_ ,
    \new_[7362]_ , \new_[7363]_ , \new_[7367]_ , \new_[7368]_ ,
    \new_[7369]_ , \new_[7373]_ , \new_[7374]_ , \new_[7378]_ ,
    \new_[7379]_ , \new_[7380]_ , \new_[7381]_ , \new_[7382]_ ,
    \new_[7386]_ , \new_[7387]_ , \new_[7391]_ , \new_[7392]_ ,
    \new_[7393]_ , \new_[7397]_ , \new_[7398]_ , \new_[7402]_ ,
    \new_[7403]_ , \new_[7404]_ , \new_[7405]_ , \new_[7409]_ ,
    \new_[7410]_ , \new_[7414]_ , \new_[7415]_ , \new_[7416]_ ,
    \new_[7420]_ , \new_[7421]_ , \new_[7424]_ , \new_[7427]_ ,
    \new_[7428]_ , \new_[7429]_ , \new_[7430]_ , \new_[7431]_ ,
    \new_[7432]_ , \new_[7436]_ , \new_[7437]_ , \new_[7441]_ ,
    \new_[7442]_ , \new_[7443]_ , \new_[7447]_ , \new_[7448]_ ,
    \new_[7452]_ , \new_[7453]_ , \new_[7454]_ , \new_[7455]_ ,
    \new_[7459]_ , \new_[7460]_ , \new_[7464]_ , \new_[7465]_ ,
    \new_[7466]_ , \new_[7470]_ , \new_[7471]_ , \new_[7474]_ ,
    \new_[7477]_ , \new_[7478]_ , \new_[7479]_ , \new_[7480]_ ,
    \new_[7481]_ , \new_[7485]_ , \new_[7486]_ , \new_[7490]_ ,
    \new_[7491]_ , \new_[7492]_ , \new_[7496]_ , \new_[7497]_ ,
    \new_[7501]_ , \new_[7502]_ , \new_[7503]_ , \new_[7504]_ ,
    \new_[7508]_ , \new_[7509]_ , \new_[7513]_ , \new_[7514]_ ,
    \new_[7515]_ , \new_[7519]_ , \new_[7520]_ , \new_[7523]_ ,
    \new_[7526]_ , \new_[7527]_ , \new_[7528]_ , \new_[7529]_ ,
    \new_[7530]_ , \new_[7531]_ , \new_[7532]_ , \new_[7533]_ ,
    \new_[7537]_ , \new_[7538]_ , \new_[7542]_ , \new_[7543]_ ,
    \new_[7544]_ , \new_[7548]_ , \new_[7549]_ , \new_[7553]_ ,
    \new_[7554]_ , \new_[7555]_ , \new_[7556]_ , \new_[7560]_ ,
    \new_[7561]_ , \new_[7565]_ , \new_[7566]_ , \new_[7567]_ ,
    \new_[7571]_ , \new_[7572]_ , \new_[7576]_ , \new_[7577]_ ,
    \new_[7578]_ , \new_[7579]_ , \new_[7580]_ , \new_[7584]_ ,
    \new_[7585]_ , \new_[7589]_ , \new_[7590]_ , \new_[7591]_ ,
    \new_[7595]_ , \new_[7596]_ , \new_[7600]_ , \new_[7601]_ ,
    \new_[7602]_ , \new_[7603]_ , \new_[7607]_ , \new_[7608]_ ,
    \new_[7612]_ , \new_[7613]_ , \new_[7614]_ , \new_[7618]_ ,
    \new_[7619]_ , \new_[7622]_ , \new_[7625]_ , \new_[7626]_ ,
    \new_[7627]_ , \new_[7628]_ , \new_[7629]_ , \new_[7630]_ ,
    \new_[7634]_ , \new_[7635]_ , \new_[7639]_ , \new_[7640]_ ,
    \new_[7641]_ , \new_[7645]_ , \new_[7646]_ , \new_[7650]_ ,
    \new_[7651]_ , \new_[7652]_ , \new_[7653]_ , \new_[7657]_ ,
    \new_[7658]_ , \new_[7662]_ , \new_[7663]_ , \new_[7664]_ ,
    \new_[7668]_ , \new_[7669]_ , \new_[7672]_ , \new_[7675]_ ,
    \new_[7676]_ , \new_[7677]_ , \new_[7678]_ , \new_[7679]_ ,
    \new_[7683]_ , \new_[7684]_ , \new_[7688]_ , \new_[7689]_ ,
    \new_[7690]_ , \new_[7694]_ , \new_[7695]_ , \new_[7699]_ ,
    \new_[7700]_ , \new_[7701]_ , \new_[7702]_ , \new_[7706]_ ,
    \new_[7707]_ , \new_[7711]_ , \new_[7712]_ , \new_[7713]_ ,
    \new_[7717]_ , \new_[7718]_ , \new_[7721]_ , \new_[7724]_ ,
    \new_[7725]_ , \new_[7726]_ , \new_[7727]_ , \new_[7728]_ ,
    \new_[7729]_ , \new_[7730]_ , \new_[7734]_ , \new_[7735]_ ,
    \new_[7739]_ , \new_[7740]_ , \new_[7741]_ , \new_[7745]_ ,
    \new_[7746]_ , \new_[7750]_ , \new_[7751]_ , \new_[7752]_ ,
    \new_[7753]_ , \new_[7757]_ , \new_[7758]_ , \new_[7762]_ ,
    \new_[7763]_ , \new_[7764]_ , \new_[7768]_ , \new_[7769]_ ,
    \new_[7772]_ , \new_[7775]_ , \new_[7776]_ , \new_[7777]_ ,
    \new_[7778]_ , \new_[7779]_ , \new_[7783]_ , \new_[7784]_ ,
    \new_[7788]_ , \new_[7789]_ , \new_[7790]_ , \new_[7794]_ ,
    \new_[7795]_ , \new_[7799]_ , \new_[7800]_ , \new_[7801]_ ,
    \new_[7802]_ , \new_[7806]_ , \new_[7807]_ , \new_[7811]_ ,
    \new_[7812]_ , \new_[7813]_ , \new_[7817]_ , \new_[7818]_ ,
    \new_[7821]_ , \new_[7824]_ , \new_[7825]_ , \new_[7826]_ ,
    \new_[7827]_ , \new_[7828]_ , \new_[7829]_ , \new_[7833]_ ,
    \new_[7834]_ , \new_[7838]_ , \new_[7839]_ , \new_[7840]_ ,
    \new_[7844]_ , \new_[7845]_ , \new_[7849]_ , \new_[7850]_ ,
    \new_[7851]_ , \new_[7852]_ , \new_[7856]_ , \new_[7857]_ ,
    \new_[7861]_ , \new_[7862]_ , \new_[7863]_ , \new_[7867]_ ,
    \new_[7868]_ , \new_[7871]_ , \new_[7874]_ , \new_[7875]_ ,
    \new_[7876]_ , \new_[7877]_ , \new_[7878]_ , \new_[7882]_ ,
    \new_[7883]_ , \new_[7887]_ , \new_[7888]_ , \new_[7889]_ ,
    \new_[7893]_ , \new_[7894]_ , \new_[7898]_ , \new_[7899]_ ,
    \new_[7900]_ , \new_[7901]_ , \new_[7905]_ , \new_[7906]_ ,
    \new_[7910]_ , \new_[7911]_ , \new_[7912]_ , \new_[7916]_ ,
    \new_[7917]_ , \new_[7920]_ , \new_[7923]_ , \new_[7924]_ ,
    \new_[7925]_ , \new_[7926]_ , \new_[7927]_ , \new_[7928]_ ,
    \new_[7929]_ , \new_[7930]_ , \new_[7931]_ , \new_[7932]_ ,
    \new_[7936]_ , \new_[7937]_ , \new_[7941]_ , \new_[7942]_ ,
    \new_[7943]_ , \new_[7947]_ , \new_[7948]_ , \new_[7952]_ ,
    \new_[7953]_ , \new_[7954]_ , \new_[7955]_ , \new_[7959]_ ,
    \new_[7960]_ , \new_[7964]_ , \new_[7965]_ , \new_[7966]_ ,
    \new_[7970]_ , \new_[7971]_ , \new_[7975]_ , \new_[7976]_ ,
    \new_[7977]_ , \new_[7978]_ , \new_[7979]_ , \new_[7983]_ ,
    \new_[7984]_ , \new_[7988]_ , \new_[7989]_ , \new_[7990]_ ,
    \new_[7994]_ , \new_[7995]_ , \new_[7999]_ , \new_[8000]_ ,
    \new_[8001]_ , \new_[8002]_ , \new_[8006]_ , \new_[8007]_ ,
    \new_[8011]_ , \new_[8012]_ , \new_[8013]_ , \new_[8017]_ ,
    \new_[8018]_ , \new_[8021]_ , \new_[8024]_ , \new_[8025]_ ,
    \new_[8026]_ , \new_[8027]_ , \new_[8028]_ , \new_[8029]_ ,
    \new_[8033]_ , \new_[8034]_ , \new_[8038]_ , \new_[8039]_ ,
    \new_[8040]_ , \new_[8044]_ , \new_[8045]_ , \new_[8049]_ ,
    \new_[8050]_ , \new_[8051]_ , \new_[8052]_ , \new_[8056]_ ,
    \new_[8057]_ , \new_[8061]_ , \new_[8062]_ , \new_[8063]_ ,
    \new_[8067]_ , \new_[8068]_ , \new_[8071]_ , \new_[8074]_ ,
    \new_[8075]_ , \new_[8076]_ , \new_[8077]_ , \new_[8078]_ ,
    \new_[8082]_ , \new_[8083]_ , \new_[8087]_ , \new_[8088]_ ,
    \new_[8089]_ , \new_[8093]_ , \new_[8094]_ , \new_[8098]_ ,
    \new_[8099]_ , \new_[8100]_ , \new_[8101]_ , \new_[8105]_ ,
    \new_[8106]_ , \new_[8110]_ , \new_[8111]_ , \new_[8112]_ ,
    \new_[8116]_ , \new_[8117]_ , \new_[8120]_ , \new_[8123]_ ,
    \new_[8124]_ , \new_[8125]_ , \new_[8126]_ , \new_[8127]_ ,
    \new_[8128]_ , \new_[8129]_ , \new_[8133]_ , \new_[8134]_ ,
    \new_[8138]_ , \new_[8139]_ , \new_[8140]_ , \new_[8144]_ ,
    \new_[8145]_ , \new_[8149]_ , \new_[8150]_ , \new_[8151]_ ,
    \new_[8152]_ , \new_[8156]_ , \new_[8157]_ , \new_[8161]_ ,
    \new_[8162]_ , \new_[8163]_ , \new_[8167]_ , \new_[8168]_ ,
    \new_[8172]_ , \new_[8173]_ , \new_[8174]_ , \new_[8175]_ ,
    \new_[8176]_ , \new_[8180]_ , \new_[8181]_ , \new_[8185]_ ,
    \new_[8186]_ , \new_[8187]_ , \new_[8191]_ , \new_[8192]_ ,
    \new_[8196]_ , \new_[8197]_ , \new_[8198]_ , \new_[8199]_ ,
    \new_[8203]_ , \new_[8204]_ , \new_[8208]_ , \new_[8209]_ ,
    \new_[8210]_ , \new_[8214]_ , \new_[8215]_ , \new_[8218]_ ,
    \new_[8221]_ , \new_[8222]_ , \new_[8223]_ , \new_[8224]_ ,
    \new_[8225]_ , \new_[8226]_ , \new_[8230]_ , \new_[8231]_ ,
    \new_[8235]_ , \new_[8236]_ , \new_[8237]_ , \new_[8241]_ ,
    \new_[8242]_ , \new_[8246]_ , \new_[8247]_ , \new_[8248]_ ,
    \new_[8249]_ , \new_[8253]_ , \new_[8254]_ , \new_[8258]_ ,
    \new_[8259]_ , \new_[8260]_ , \new_[8264]_ , \new_[8265]_ ,
    \new_[8268]_ , \new_[8271]_ , \new_[8272]_ , \new_[8273]_ ,
    \new_[8274]_ , \new_[8275]_ , \new_[8279]_ , \new_[8280]_ ,
    \new_[8284]_ , \new_[8285]_ , \new_[8286]_ , \new_[8290]_ ,
    \new_[8291]_ , \new_[8295]_ , \new_[8296]_ , \new_[8297]_ ,
    \new_[8298]_ , \new_[8302]_ , \new_[8303]_ , \new_[8307]_ ,
    \new_[8308]_ , \new_[8309]_ , \new_[8313]_ , \new_[8314]_ ,
    \new_[8317]_ , \new_[8320]_ , \new_[8321]_ , \new_[8322]_ ,
    \new_[8323]_ , \new_[8324]_ , \new_[8325]_ , \new_[8326]_ ,
    \new_[8327]_ , \new_[8331]_ , \new_[8332]_ , \new_[8336]_ ,
    \new_[8337]_ , \new_[8338]_ , \new_[8342]_ , \new_[8343]_ ,
    \new_[8347]_ , \new_[8348]_ , \new_[8349]_ , \new_[8350]_ ,
    \new_[8354]_ , \new_[8355]_ , \new_[8359]_ , \new_[8360]_ ,
    \new_[8361]_ , \new_[8365]_ , \new_[8366]_ , \new_[8370]_ ,
    \new_[8371]_ , \new_[8372]_ , \new_[8373]_ , \new_[8374]_ ,
    \new_[8378]_ , \new_[8379]_ , \new_[8383]_ , \new_[8384]_ ,
    \new_[8385]_ , \new_[8389]_ , \new_[8390]_ , \new_[8394]_ ,
    \new_[8395]_ , \new_[8396]_ , \new_[8397]_ , \new_[8401]_ ,
    \new_[8402]_ , \new_[8406]_ , \new_[8407]_ , \new_[8408]_ ,
    \new_[8412]_ , \new_[8413]_ , \new_[8416]_ , \new_[8419]_ ,
    \new_[8420]_ , \new_[8421]_ , \new_[8422]_ , \new_[8423]_ ,
    \new_[8424]_ , \new_[8428]_ , \new_[8429]_ , \new_[8433]_ ,
    \new_[8434]_ , \new_[8435]_ , \new_[8439]_ , \new_[8440]_ ,
    \new_[8444]_ , \new_[8445]_ , \new_[8446]_ , \new_[8447]_ ,
    \new_[8451]_ , \new_[8452]_ , \new_[8456]_ , \new_[8457]_ ,
    \new_[8458]_ , \new_[8462]_ , \new_[8463]_ , \new_[8466]_ ,
    \new_[8469]_ , \new_[8470]_ , \new_[8471]_ , \new_[8472]_ ,
    \new_[8473]_ , \new_[8477]_ , \new_[8478]_ , \new_[8482]_ ,
    \new_[8483]_ , \new_[8484]_ , \new_[8488]_ , \new_[8489]_ ,
    \new_[8493]_ , \new_[8494]_ , \new_[8495]_ , \new_[8496]_ ,
    \new_[8500]_ , \new_[8501]_ , \new_[8505]_ , \new_[8506]_ ,
    \new_[8507]_ , \new_[8511]_ , \new_[8512]_ , \new_[8515]_ ,
    \new_[8518]_ , \new_[8519]_ , \new_[8520]_ , \new_[8521]_ ,
    \new_[8522]_ , \new_[8523]_ , \new_[8524]_ , \new_[8528]_ ,
    \new_[8529]_ , \new_[8533]_ , \new_[8534]_ , \new_[8535]_ ,
    \new_[8539]_ , \new_[8540]_ , \new_[8544]_ , \new_[8545]_ ,
    \new_[8546]_ , \new_[8547]_ , \new_[8551]_ , \new_[8552]_ ,
    \new_[8556]_ , \new_[8557]_ , \new_[8558]_ , \new_[8562]_ ,
    \new_[8563]_ , \new_[8566]_ , \new_[8569]_ , \new_[8570]_ ,
    \new_[8571]_ , \new_[8572]_ , \new_[8573]_ , \new_[8577]_ ,
    \new_[8578]_ , \new_[8582]_ , \new_[8583]_ , \new_[8584]_ ,
    \new_[8588]_ , \new_[8589]_ , \new_[8593]_ , \new_[8594]_ ,
    \new_[8595]_ , \new_[8596]_ , \new_[8600]_ , \new_[8601]_ ,
    \new_[8605]_ , \new_[8606]_ , \new_[8607]_ , \new_[8611]_ ,
    \new_[8612]_ , \new_[8615]_ , \new_[8618]_ , \new_[8619]_ ,
    \new_[8620]_ , \new_[8621]_ , \new_[8622]_ , \new_[8623]_ ,
    \new_[8627]_ , \new_[8628]_ , \new_[8632]_ , \new_[8633]_ ,
    \new_[8634]_ , \new_[8638]_ , \new_[8639]_ , \new_[8643]_ ,
    \new_[8644]_ , \new_[8645]_ , \new_[8646]_ , \new_[8650]_ ,
    \new_[8651]_ , \new_[8655]_ , \new_[8656]_ , \new_[8657]_ ,
    \new_[8661]_ , \new_[8662]_ , \new_[8665]_ , \new_[8668]_ ,
    \new_[8669]_ , \new_[8670]_ , \new_[8671]_ , \new_[8672]_ ,
    \new_[8676]_ , \new_[8677]_ , \new_[8681]_ , \new_[8682]_ ,
    \new_[8683]_ , \new_[8687]_ , \new_[8688]_ , \new_[8692]_ ,
    \new_[8693]_ , \new_[8694]_ , \new_[8695]_ , \new_[8699]_ ,
    \new_[8700]_ , \new_[8704]_ , \new_[8705]_ , \new_[8706]_ ,
    \new_[8710]_ , \new_[8711]_ , \new_[8714]_ , \new_[8717]_ ,
    \new_[8718]_ , \new_[8719]_ , \new_[8720]_ , \new_[8721]_ ,
    \new_[8722]_ , \new_[8723]_ , \new_[8724]_ , \new_[8725]_ ,
    \new_[8729]_ , \new_[8730]_ , \new_[8734]_ , \new_[8735]_ ,
    \new_[8736]_ , \new_[8740]_ , \new_[8741]_ , \new_[8745]_ ,
    \new_[8746]_ , \new_[8747]_ , \new_[8748]_ , \new_[8752]_ ,
    \new_[8753]_ , \new_[8757]_ , \new_[8758]_ , \new_[8759]_ ,
    \new_[8763]_ , \new_[8764]_ , \new_[8768]_ , \new_[8769]_ ,
    \new_[8770]_ , \new_[8771]_ , \new_[8772]_ , \new_[8776]_ ,
    \new_[8777]_ , \new_[8781]_ , \new_[8782]_ , \new_[8783]_ ,
    \new_[8787]_ , \new_[8788]_ , \new_[8792]_ , \new_[8793]_ ,
    \new_[8794]_ , \new_[8795]_ , \new_[8799]_ , \new_[8800]_ ,
    \new_[8804]_ , \new_[8805]_ , \new_[8806]_ , \new_[8810]_ ,
    \new_[8811]_ , \new_[8814]_ , \new_[8817]_ , \new_[8818]_ ,
    \new_[8819]_ , \new_[8820]_ , \new_[8821]_ , \new_[8822]_ ,
    \new_[8826]_ , \new_[8827]_ , \new_[8831]_ , \new_[8832]_ ,
    \new_[8833]_ , \new_[8837]_ , \new_[8838]_ , \new_[8842]_ ,
    \new_[8843]_ , \new_[8844]_ , \new_[8845]_ , \new_[8849]_ ,
    \new_[8850]_ , \new_[8854]_ , \new_[8855]_ , \new_[8856]_ ,
    \new_[8860]_ , \new_[8861]_ , \new_[8864]_ , \new_[8867]_ ,
    \new_[8868]_ , \new_[8869]_ , \new_[8870]_ , \new_[8871]_ ,
    \new_[8875]_ , \new_[8876]_ , \new_[8880]_ , \new_[8881]_ ,
    \new_[8882]_ , \new_[8886]_ , \new_[8887]_ , \new_[8891]_ ,
    \new_[8892]_ , \new_[8893]_ , \new_[8894]_ , \new_[8898]_ ,
    \new_[8899]_ , \new_[8903]_ , \new_[8904]_ , \new_[8905]_ ,
    \new_[8909]_ , \new_[8910]_ , \new_[8913]_ , \new_[8916]_ ,
    \new_[8917]_ , \new_[8918]_ , \new_[8919]_ , \new_[8920]_ ,
    \new_[8921]_ , \new_[8922]_ , \new_[8926]_ , \new_[8927]_ ,
    \new_[8931]_ , \new_[8932]_ , \new_[8933]_ , \new_[8937]_ ,
    \new_[8938]_ , \new_[8942]_ , \new_[8943]_ , \new_[8944]_ ,
    \new_[8945]_ , \new_[8949]_ , \new_[8950]_ , \new_[8954]_ ,
    \new_[8955]_ , \new_[8956]_ , \new_[8960]_ , \new_[8961]_ ,
    \new_[8965]_ , \new_[8966]_ , \new_[8967]_ , \new_[8968]_ ,
    \new_[8969]_ , \new_[8973]_ , \new_[8974]_ , \new_[8978]_ ,
    \new_[8979]_ , \new_[8980]_ , \new_[8984]_ , \new_[8985]_ ,
    \new_[8989]_ , \new_[8990]_ , \new_[8991]_ , \new_[8992]_ ,
    \new_[8996]_ , \new_[8997]_ , \new_[9001]_ , \new_[9002]_ ,
    \new_[9003]_ , \new_[9007]_ , \new_[9008]_ , \new_[9011]_ ,
    \new_[9014]_ , \new_[9015]_ , \new_[9016]_ , \new_[9017]_ ,
    \new_[9018]_ , \new_[9019]_ , \new_[9023]_ , \new_[9024]_ ,
    \new_[9028]_ , \new_[9029]_ , \new_[9030]_ , \new_[9034]_ ,
    \new_[9035]_ , \new_[9039]_ , \new_[9040]_ , \new_[9041]_ ,
    \new_[9042]_ , \new_[9046]_ , \new_[9047]_ , \new_[9051]_ ,
    \new_[9052]_ , \new_[9053]_ , \new_[9057]_ , \new_[9058]_ ,
    \new_[9061]_ , \new_[9064]_ , \new_[9065]_ , \new_[9066]_ ,
    \new_[9067]_ , \new_[9068]_ , \new_[9072]_ , \new_[9073]_ ,
    \new_[9077]_ , \new_[9078]_ , \new_[9079]_ , \new_[9083]_ ,
    \new_[9084]_ , \new_[9088]_ , \new_[9089]_ , \new_[9090]_ ,
    \new_[9091]_ , \new_[9095]_ , \new_[9096]_ , \new_[9100]_ ,
    \new_[9101]_ , \new_[9102]_ , \new_[9106]_ , \new_[9107]_ ,
    \new_[9110]_ , \new_[9113]_ , \new_[9114]_ , \new_[9115]_ ,
    \new_[9116]_ , \new_[9117]_ , \new_[9118]_ , \new_[9119]_ ,
    \new_[9120]_ , \new_[9124]_ , \new_[9125]_ , \new_[9129]_ ,
    \new_[9130]_ , \new_[9131]_ , \new_[9135]_ , \new_[9136]_ ,
    \new_[9140]_ , \new_[9141]_ , \new_[9142]_ , \new_[9143]_ ,
    \new_[9147]_ , \new_[9148]_ , \new_[9152]_ , \new_[9153]_ ,
    \new_[9154]_ , \new_[9158]_ , \new_[9159]_ , \new_[9163]_ ,
    \new_[9164]_ , \new_[9165]_ , \new_[9166]_ , \new_[9167]_ ,
    \new_[9171]_ , \new_[9172]_ , \new_[9176]_ , \new_[9177]_ ,
    \new_[9178]_ , \new_[9182]_ , \new_[9183]_ , \new_[9187]_ ,
    \new_[9188]_ , \new_[9189]_ , \new_[9190]_ , \new_[9194]_ ,
    \new_[9195]_ , \new_[9199]_ , \new_[9200]_ , \new_[9201]_ ,
    \new_[9205]_ , \new_[9206]_ , \new_[9209]_ , \new_[9212]_ ,
    \new_[9213]_ , \new_[9214]_ , \new_[9215]_ , \new_[9216]_ ,
    \new_[9217]_ , \new_[9221]_ , \new_[9222]_ , \new_[9226]_ ,
    \new_[9227]_ , \new_[9228]_ , \new_[9232]_ , \new_[9233]_ ,
    \new_[9237]_ , \new_[9238]_ , \new_[9239]_ , \new_[9240]_ ,
    \new_[9244]_ , \new_[9245]_ , \new_[9249]_ , \new_[9250]_ ,
    \new_[9251]_ , \new_[9255]_ , \new_[9256]_ , \new_[9259]_ ,
    \new_[9262]_ , \new_[9263]_ , \new_[9264]_ , \new_[9265]_ ,
    \new_[9266]_ , \new_[9270]_ , \new_[9271]_ , \new_[9275]_ ,
    \new_[9276]_ , \new_[9277]_ , \new_[9281]_ , \new_[9282]_ ,
    \new_[9286]_ , \new_[9287]_ , \new_[9288]_ , \new_[9289]_ ,
    \new_[9293]_ , \new_[9294]_ , \new_[9298]_ , \new_[9299]_ ,
    \new_[9300]_ , \new_[9304]_ , \new_[9305]_ , \new_[9308]_ ,
    \new_[9311]_ , \new_[9312]_ , \new_[9313]_ , \new_[9314]_ ,
    \new_[9315]_ , \new_[9316]_ , \new_[9317]_ , \new_[9321]_ ,
    \new_[9322]_ , \new_[9326]_ , \new_[9327]_ , \new_[9328]_ ,
    \new_[9332]_ , \new_[9333]_ , \new_[9337]_ , \new_[9338]_ ,
    \new_[9339]_ , \new_[9340]_ , \new_[9344]_ , \new_[9345]_ ,
    \new_[9349]_ , \new_[9350]_ , \new_[9351]_ , \new_[9355]_ ,
    \new_[9356]_ , \new_[9359]_ , \new_[9362]_ , \new_[9363]_ ,
    \new_[9364]_ , \new_[9365]_ , \new_[9366]_ , \new_[9370]_ ,
    \new_[9371]_ , \new_[9375]_ , \new_[9376]_ , \new_[9377]_ ,
    \new_[9381]_ , \new_[9382]_ , \new_[9386]_ , \new_[9387]_ ,
    \new_[9388]_ , \new_[9389]_ , \new_[9393]_ , \new_[9394]_ ,
    \new_[9398]_ , \new_[9399]_ , \new_[9400]_ , \new_[9404]_ ,
    \new_[9405]_ , \new_[9408]_ , \new_[9411]_ , \new_[9412]_ ,
    \new_[9413]_ , \new_[9414]_ , \new_[9415]_ , \new_[9416]_ ,
    \new_[9420]_ , \new_[9421]_ , \new_[9425]_ , \new_[9426]_ ,
    \new_[9427]_ , \new_[9431]_ , \new_[9432]_ , \new_[9436]_ ,
    \new_[9437]_ , \new_[9438]_ , \new_[9439]_ , \new_[9443]_ ,
    \new_[9444]_ , \new_[9448]_ , \new_[9449]_ , \new_[9450]_ ,
    \new_[9454]_ , \new_[9455]_ , \new_[9458]_ , \new_[9461]_ ,
    \new_[9462]_ , \new_[9463]_ , \new_[9464]_ , \new_[9465]_ ,
    \new_[9469]_ , \new_[9470]_ , \new_[9474]_ , \new_[9475]_ ,
    \new_[9476]_ , \new_[9480]_ , \new_[9481]_ , \new_[9485]_ ,
    \new_[9486]_ , \new_[9487]_ , \new_[9488]_ , \new_[9492]_ ,
    \new_[9493]_ , \new_[9497]_ , \new_[9498]_ , \new_[9499]_ ,
    \new_[9503]_ , \new_[9504]_ , \new_[9507]_ , \new_[9510]_ ,
    \new_[9511]_ , \new_[9512]_ , \new_[9513]_ , \new_[9514]_ ,
    \new_[9515]_ , \new_[9516]_ , \new_[9517]_ , \new_[9518]_ ,
    \new_[9519]_ , \new_[9520]_ , \new_[9523]_ , \new_[9526]_ ,
    \new_[9527]_ , \new_[9530]_ , \new_[9533]_ , \new_[9534]_ ,
    \new_[9537]_ , \new_[9540]_ , \new_[9541]_ , \new_[9544]_ ,
    \new_[9547]_ , \new_[9548]_ , \new_[9551]_ , \new_[9554]_ ,
    \new_[9555]_ , \new_[9558]_ , \new_[9561]_ , \new_[9562]_ ,
    \new_[9565]_ , \new_[9568]_ , \new_[9569]_ , \new_[9572]_ ,
    \new_[9575]_ , \new_[9576]_ , \new_[9579]_ , \new_[9582]_ ,
    \new_[9583]_ , \new_[9586]_ , \new_[9589]_ , \new_[9590]_ ,
    \new_[9593]_ , \new_[9596]_ , \new_[9597]_ , \new_[9600]_ ,
    \new_[9603]_ , \new_[9604]_ , \new_[9607]_ , \new_[9610]_ ,
    \new_[9611]_ , \new_[9614]_ , \new_[9617]_ , \new_[9618]_ ,
    \new_[9621]_ , \new_[9624]_ , \new_[9625]_ , \new_[9628]_ ,
    \new_[9631]_ , \new_[9632]_ , \new_[9635]_ , \new_[9638]_ ,
    \new_[9639]_ , \new_[9642]_ , \new_[9645]_ , \new_[9646]_ ,
    \new_[9649]_ , \new_[9652]_ , \new_[9653]_ , \new_[9656]_ ,
    \new_[9659]_ , \new_[9660]_ , \new_[9663]_ , \new_[9666]_ ,
    \new_[9667]_ , \new_[9670]_ , \new_[9673]_ , \new_[9674]_ ,
    \new_[9677]_ , \new_[9680]_ , \new_[9681]_ , \new_[9684]_ ,
    \new_[9687]_ , \new_[9688]_ , \new_[9691]_ , \new_[9694]_ ,
    \new_[9695]_ , \new_[9698]_ , \new_[9701]_ , \new_[9702]_ ,
    \new_[9705]_ , \new_[9708]_ , \new_[9709]_ , \new_[9712]_ ,
    \new_[9715]_ , \new_[9716]_ , \new_[9719]_ , \new_[9722]_ ,
    \new_[9723]_ , \new_[9726]_ , \new_[9729]_ , \new_[9730]_ ,
    \new_[9733]_ , \new_[9736]_ , \new_[9737]_ , \new_[9740]_ ,
    \new_[9743]_ , \new_[9744]_ , \new_[9747]_ , \new_[9750]_ ,
    \new_[9751]_ , \new_[9754]_ , \new_[9757]_ , \new_[9758]_ ,
    \new_[9761]_ , \new_[9764]_ , \new_[9765]_ , \new_[9768]_ ,
    \new_[9771]_ , \new_[9772]_ , \new_[9775]_ , \new_[9778]_ ,
    \new_[9779]_ , \new_[9782]_ , \new_[9785]_ , \new_[9786]_ ,
    \new_[9789]_ , \new_[9792]_ , \new_[9793]_ , \new_[9796]_ ,
    \new_[9799]_ , \new_[9800]_ , \new_[9803]_ , \new_[9806]_ ,
    \new_[9807]_ , \new_[9810]_ , \new_[9813]_ , \new_[9814]_ ,
    \new_[9817]_ , \new_[9820]_ , \new_[9821]_ , \new_[9824]_ ,
    \new_[9827]_ , \new_[9828]_ , \new_[9831]_ , \new_[9834]_ ,
    \new_[9835]_ , \new_[9838]_ , \new_[9841]_ , \new_[9842]_ ,
    \new_[9845]_ , \new_[9848]_ , \new_[9849]_ , \new_[9852]_ ,
    \new_[9855]_ , \new_[9856]_ , \new_[9859]_ , \new_[9862]_ ,
    \new_[9863]_ , \new_[9866]_ , \new_[9870]_ , \new_[9871]_ ,
    \new_[9872]_ , \new_[9875]_ , \new_[9878]_ , \new_[9879]_ ,
    \new_[9882]_ , \new_[9886]_ , \new_[9887]_ , \new_[9888]_ ,
    \new_[9891]_ , \new_[9894]_ , \new_[9895]_ , \new_[9898]_ ,
    \new_[9902]_ , \new_[9903]_ , \new_[9904]_ , \new_[9907]_ ,
    \new_[9910]_ , \new_[9911]_ , \new_[9914]_ , \new_[9918]_ ,
    \new_[9919]_ , \new_[9920]_ , \new_[9923]_ , \new_[9926]_ ,
    \new_[9927]_ , \new_[9930]_ , \new_[9934]_ , \new_[9935]_ ,
    \new_[9936]_ , \new_[9939]_ , \new_[9942]_ , \new_[9943]_ ,
    \new_[9946]_ , \new_[9950]_ , \new_[9951]_ , \new_[9952]_ ,
    \new_[9955]_ , \new_[9958]_ , \new_[9959]_ , \new_[9962]_ ,
    \new_[9966]_ , \new_[9967]_ , \new_[9968]_ , \new_[9971]_ ,
    \new_[9974]_ , \new_[9975]_ , \new_[9978]_ , \new_[9982]_ ,
    \new_[9983]_ , \new_[9984]_ , \new_[9987]_ , \new_[9990]_ ,
    \new_[9991]_ , \new_[9994]_ , \new_[9998]_ , \new_[9999]_ ,
    \new_[10000]_ , \new_[10003]_ , \new_[10006]_ , \new_[10007]_ ,
    \new_[10010]_ , \new_[10014]_ , \new_[10015]_ , \new_[10016]_ ,
    \new_[10019]_ , \new_[10022]_ , \new_[10023]_ , \new_[10026]_ ,
    \new_[10030]_ , \new_[10031]_ , \new_[10032]_ , \new_[10035]_ ,
    \new_[10038]_ , \new_[10039]_ , \new_[10042]_ , \new_[10046]_ ,
    \new_[10047]_ , \new_[10048]_ , \new_[10051]_ , \new_[10054]_ ,
    \new_[10055]_ , \new_[10058]_ , \new_[10062]_ , \new_[10063]_ ,
    \new_[10064]_ , \new_[10067]_ , \new_[10070]_ , \new_[10071]_ ,
    \new_[10074]_ , \new_[10078]_ , \new_[10079]_ , \new_[10080]_ ,
    \new_[10083]_ , \new_[10086]_ , \new_[10087]_ , \new_[10090]_ ,
    \new_[10094]_ , \new_[10095]_ , \new_[10096]_ , \new_[10099]_ ,
    \new_[10102]_ , \new_[10103]_ , \new_[10106]_ , \new_[10110]_ ,
    \new_[10111]_ , \new_[10112]_ , \new_[10115]_ , \new_[10118]_ ,
    \new_[10119]_ , \new_[10122]_ , \new_[10126]_ , \new_[10127]_ ,
    \new_[10128]_ , \new_[10131]_ , \new_[10134]_ , \new_[10135]_ ,
    \new_[10138]_ , \new_[10142]_ , \new_[10143]_ , \new_[10144]_ ,
    \new_[10147]_ , \new_[10150]_ , \new_[10151]_ , \new_[10154]_ ,
    \new_[10158]_ , \new_[10159]_ , \new_[10160]_ , \new_[10163]_ ,
    \new_[10166]_ , \new_[10167]_ , \new_[10170]_ , \new_[10174]_ ,
    \new_[10175]_ , \new_[10176]_ , \new_[10179]_ , \new_[10182]_ ,
    \new_[10183]_ , \new_[10186]_ , \new_[10190]_ , \new_[10191]_ ,
    \new_[10192]_ , \new_[10195]_ , \new_[10198]_ , \new_[10199]_ ,
    \new_[10202]_ , \new_[10206]_ , \new_[10207]_ , \new_[10208]_ ,
    \new_[10211]_ , \new_[10215]_ , \new_[10216]_ , \new_[10217]_ ,
    \new_[10220]_ , \new_[10224]_ , \new_[10225]_ , \new_[10226]_ ,
    \new_[10229]_ , \new_[10233]_ , \new_[10234]_ , \new_[10235]_ ,
    \new_[10238]_ , \new_[10242]_ , \new_[10243]_ , \new_[10244]_ ,
    \new_[10247]_ , \new_[10251]_ , \new_[10252]_ , \new_[10253]_ ,
    \new_[10256]_ , \new_[10260]_ , \new_[10261]_ , \new_[10262]_ ,
    \new_[10265]_ , \new_[10269]_ , \new_[10270]_ , \new_[10271]_ ,
    \new_[10274]_ , \new_[10278]_ , \new_[10279]_ , \new_[10280]_ ,
    \new_[10283]_ , \new_[10287]_ , \new_[10288]_ , \new_[10289]_ ,
    \new_[10292]_ , \new_[10296]_ , \new_[10297]_ , \new_[10298]_ ,
    \new_[10301]_ , \new_[10305]_ , \new_[10306]_ , \new_[10307]_ ,
    \new_[10310]_ , \new_[10314]_ , \new_[10315]_ , \new_[10316]_ ,
    \new_[10319]_ , \new_[10323]_ , \new_[10324]_ , \new_[10325]_ ,
    \new_[10328]_ , \new_[10332]_ , \new_[10333]_ , \new_[10334]_ ,
    \new_[10337]_ , \new_[10341]_ , \new_[10342]_ , \new_[10343]_ ,
    \new_[10346]_ , \new_[10350]_ , \new_[10351]_ , \new_[10352]_ ,
    \new_[10355]_ , \new_[10359]_ , \new_[10360]_ , \new_[10361]_ ,
    \new_[10364]_ , \new_[10368]_ , \new_[10369]_ , \new_[10370]_ ,
    \new_[10373]_ , \new_[10377]_ , \new_[10378]_ , \new_[10379]_ ,
    \new_[10382]_ , \new_[10386]_ , \new_[10387]_ , \new_[10388]_ ,
    \new_[10391]_ , \new_[10395]_ , \new_[10396]_ , \new_[10397]_ ,
    \new_[10400]_ , \new_[10404]_ , \new_[10405]_ , \new_[10406]_ ,
    \new_[10409]_ , \new_[10413]_ , \new_[10414]_ , \new_[10415]_ ,
    \new_[10418]_ , \new_[10422]_ , \new_[10423]_ , \new_[10424]_ ,
    \new_[10427]_ , \new_[10431]_ , \new_[10432]_ , \new_[10433]_ ,
    \new_[10436]_ , \new_[10440]_ , \new_[10441]_ , \new_[10442]_ ,
    \new_[10445]_ , \new_[10449]_ , \new_[10450]_ , \new_[10451]_ ,
    \new_[10454]_ , \new_[10458]_ , \new_[10459]_ , \new_[10460]_ ,
    \new_[10463]_ , \new_[10467]_ , \new_[10468]_ , \new_[10469]_ ,
    \new_[10472]_ , \new_[10476]_ , \new_[10477]_ , \new_[10478]_ ,
    \new_[10481]_ , \new_[10485]_ , \new_[10486]_ , \new_[10487]_ ,
    \new_[10490]_ , \new_[10494]_ , \new_[10495]_ , \new_[10496]_ ,
    \new_[10499]_ , \new_[10503]_ , \new_[10504]_ , \new_[10505]_ ,
    \new_[10508]_ , \new_[10512]_ , \new_[10513]_ , \new_[10514]_ ,
    \new_[10517]_ , \new_[10521]_ , \new_[10522]_ , \new_[10523]_ ,
    \new_[10526]_ , \new_[10530]_ , \new_[10531]_ , \new_[10532]_ ,
    \new_[10535]_ , \new_[10539]_ , \new_[10540]_ , \new_[10541]_ ,
    \new_[10544]_ , \new_[10548]_ , \new_[10549]_ , \new_[10550]_ ,
    \new_[10553]_ , \new_[10557]_ , \new_[10558]_ , \new_[10559]_ ,
    \new_[10562]_ , \new_[10566]_ , \new_[10567]_ , \new_[10568]_ ,
    \new_[10571]_ , \new_[10575]_ , \new_[10576]_ , \new_[10577]_ ,
    \new_[10580]_ , \new_[10584]_ , \new_[10585]_ , \new_[10586]_ ,
    \new_[10589]_ , \new_[10593]_ , \new_[10594]_ , \new_[10595]_ ,
    \new_[10598]_ , \new_[10602]_ , \new_[10603]_ , \new_[10604]_ ,
    \new_[10607]_ , \new_[10611]_ , \new_[10612]_ , \new_[10613]_ ,
    \new_[10616]_ , \new_[10620]_ , \new_[10621]_ , \new_[10622]_ ,
    \new_[10625]_ , \new_[10629]_ , \new_[10630]_ , \new_[10631]_ ,
    \new_[10634]_ , \new_[10638]_ , \new_[10639]_ , \new_[10640]_ ,
    \new_[10643]_ , \new_[10647]_ , \new_[10648]_ , \new_[10649]_ ,
    \new_[10652]_ , \new_[10656]_ , \new_[10657]_ , \new_[10658]_ ,
    \new_[10661]_ , \new_[10665]_ , \new_[10666]_ , \new_[10667]_ ,
    \new_[10670]_ , \new_[10674]_ , \new_[10675]_ , \new_[10676]_ ,
    \new_[10679]_ , \new_[10683]_ , \new_[10684]_ , \new_[10685]_ ,
    \new_[10688]_ , \new_[10692]_ , \new_[10693]_ , \new_[10694]_ ,
    \new_[10697]_ , \new_[10701]_ , \new_[10702]_ , \new_[10703]_ ,
    \new_[10706]_ , \new_[10710]_ , \new_[10711]_ , \new_[10712]_ ,
    \new_[10715]_ , \new_[10719]_ , \new_[10720]_ , \new_[10721]_ ,
    \new_[10724]_ , \new_[10728]_ , \new_[10729]_ , \new_[10730]_ ,
    \new_[10733]_ , \new_[10737]_ , \new_[10738]_ , \new_[10739]_ ,
    \new_[10742]_ , \new_[10746]_ , \new_[10747]_ , \new_[10748]_ ,
    \new_[10751]_ , \new_[10755]_ , \new_[10756]_ , \new_[10757]_ ,
    \new_[10760]_ , \new_[10764]_ , \new_[10765]_ , \new_[10766]_ ,
    \new_[10769]_ , \new_[10773]_ , \new_[10774]_ , \new_[10775]_ ,
    \new_[10778]_ , \new_[10782]_ , \new_[10783]_ , \new_[10784]_ ,
    \new_[10787]_ , \new_[10791]_ , \new_[10792]_ , \new_[10793]_ ,
    \new_[10796]_ , \new_[10800]_ , \new_[10801]_ , \new_[10802]_ ,
    \new_[10805]_ , \new_[10809]_ , \new_[10810]_ , \new_[10811]_ ,
    \new_[10814]_ , \new_[10818]_ , \new_[10819]_ , \new_[10820]_ ,
    \new_[10823]_ , \new_[10827]_ , \new_[10828]_ , \new_[10829]_ ,
    \new_[10832]_ , \new_[10836]_ , \new_[10837]_ , \new_[10838]_ ,
    \new_[10841]_ , \new_[10845]_ , \new_[10846]_ , \new_[10847]_ ,
    \new_[10850]_ , \new_[10854]_ , \new_[10855]_ , \new_[10856]_ ,
    \new_[10859]_ , \new_[10863]_ , \new_[10864]_ , \new_[10865]_ ,
    \new_[10868]_ , \new_[10872]_ , \new_[10873]_ , \new_[10874]_ ,
    \new_[10877]_ , \new_[10881]_ , \new_[10882]_ , \new_[10883]_ ,
    \new_[10886]_ , \new_[10890]_ , \new_[10891]_ , \new_[10892]_ ,
    \new_[10895]_ , \new_[10899]_ , \new_[10900]_ , \new_[10901]_ ,
    \new_[10904]_ , \new_[10908]_ , \new_[10909]_ , \new_[10910]_ ,
    \new_[10913]_ , \new_[10917]_ , \new_[10918]_ , \new_[10919]_ ,
    \new_[10922]_ , \new_[10926]_ , \new_[10927]_ , \new_[10928]_ ,
    \new_[10931]_ , \new_[10935]_ , \new_[10936]_ , \new_[10937]_ ,
    \new_[10940]_ , \new_[10944]_ , \new_[10945]_ , \new_[10946]_ ,
    \new_[10949]_ , \new_[10953]_ , \new_[10954]_ , \new_[10955]_ ,
    \new_[10958]_ , \new_[10962]_ , \new_[10963]_ , \new_[10964]_ ,
    \new_[10967]_ , \new_[10971]_ , \new_[10972]_ , \new_[10973]_ ,
    \new_[10976]_ , \new_[10980]_ , \new_[10981]_ , \new_[10982]_ ,
    \new_[10985]_ , \new_[10989]_ , \new_[10990]_ , \new_[10991]_ ,
    \new_[10994]_ , \new_[10998]_ , \new_[10999]_ , \new_[11000]_ ,
    \new_[11003]_ , \new_[11007]_ , \new_[11008]_ , \new_[11009]_ ,
    \new_[11012]_ , \new_[11016]_ , \new_[11017]_ , \new_[11018]_ ,
    \new_[11021]_ , \new_[11025]_ , \new_[11026]_ , \new_[11027]_ ,
    \new_[11030]_ , \new_[11034]_ , \new_[11035]_ , \new_[11036]_ ,
    \new_[11039]_ , \new_[11043]_ , \new_[11044]_ , \new_[11045]_ ,
    \new_[11048]_ , \new_[11052]_ , \new_[11053]_ , \new_[11054]_ ,
    \new_[11057]_ , \new_[11061]_ , \new_[11062]_ , \new_[11063]_ ,
    \new_[11066]_ , \new_[11070]_ , \new_[11071]_ , \new_[11072]_ ,
    \new_[11075]_ , \new_[11079]_ , \new_[11080]_ , \new_[11081]_ ,
    \new_[11084]_ , \new_[11088]_ , \new_[11089]_ , \new_[11090]_ ,
    \new_[11093]_ , \new_[11097]_ , \new_[11098]_ , \new_[11099]_ ,
    \new_[11102]_ , \new_[11106]_ , \new_[11107]_ , \new_[11108]_ ,
    \new_[11111]_ , \new_[11115]_ , \new_[11116]_ , \new_[11117]_ ,
    \new_[11120]_ , \new_[11124]_ , \new_[11125]_ , \new_[11126]_ ,
    \new_[11129]_ , \new_[11133]_ , \new_[11134]_ , \new_[11135]_ ,
    \new_[11138]_ , \new_[11142]_ , \new_[11143]_ , \new_[11144]_ ,
    \new_[11147]_ , \new_[11151]_ , \new_[11152]_ , \new_[11153]_ ,
    \new_[11156]_ , \new_[11160]_ , \new_[11161]_ , \new_[11162]_ ,
    \new_[11165]_ , \new_[11169]_ , \new_[11170]_ , \new_[11171]_ ,
    \new_[11174]_ , \new_[11178]_ , \new_[11179]_ , \new_[11180]_ ,
    \new_[11183]_ , \new_[11187]_ , \new_[11188]_ , \new_[11189]_ ,
    \new_[11192]_ , \new_[11196]_ , \new_[11197]_ , \new_[11198]_ ,
    \new_[11201]_ , \new_[11205]_ , \new_[11206]_ , \new_[11207]_ ,
    \new_[11210]_ , \new_[11214]_ , \new_[11215]_ , \new_[11216]_ ,
    \new_[11219]_ , \new_[11223]_ , \new_[11224]_ , \new_[11225]_ ,
    \new_[11228]_ , \new_[11232]_ , \new_[11233]_ , \new_[11234]_ ,
    \new_[11237]_ , \new_[11241]_ , \new_[11242]_ , \new_[11243]_ ,
    \new_[11246]_ , \new_[11250]_ , \new_[11251]_ , \new_[11252]_ ,
    \new_[11255]_ , \new_[11259]_ , \new_[11260]_ , \new_[11261]_ ,
    \new_[11264]_ , \new_[11268]_ , \new_[11269]_ , \new_[11270]_ ,
    \new_[11273]_ , \new_[11277]_ , \new_[11278]_ , \new_[11279]_ ,
    \new_[11282]_ , \new_[11286]_ , \new_[11287]_ , \new_[11288]_ ,
    \new_[11291]_ , \new_[11295]_ , \new_[11296]_ , \new_[11297]_ ,
    \new_[11300]_ , \new_[11304]_ , \new_[11305]_ , \new_[11306]_ ,
    \new_[11309]_ , \new_[11313]_ , \new_[11314]_ , \new_[11315]_ ,
    \new_[11318]_ , \new_[11322]_ , \new_[11323]_ , \new_[11324]_ ,
    \new_[11327]_ , \new_[11331]_ , \new_[11332]_ , \new_[11333]_ ,
    \new_[11336]_ , \new_[11340]_ , \new_[11341]_ , \new_[11342]_ ,
    \new_[11345]_ , \new_[11349]_ , \new_[11350]_ , \new_[11351]_ ,
    \new_[11354]_ , \new_[11358]_ , \new_[11359]_ , \new_[11360]_ ,
    \new_[11363]_ , \new_[11367]_ , \new_[11368]_ , \new_[11369]_ ,
    \new_[11372]_ , \new_[11376]_ , \new_[11377]_ , \new_[11378]_ ,
    \new_[11381]_ , \new_[11385]_ , \new_[11386]_ , \new_[11387]_ ,
    \new_[11390]_ , \new_[11394]_ , \new_[11395]_ , \new_[11396]_ ,
    \new_[11399]_ , \new_[11403]_ , \new_[11404]_ , \new_[11405]_ ,
    \new_[11408]_ , \new_[11412]_ , \new_[11413]_ , \new_[11414]_ ,
    \new_[11417]_ , \new_[11421]_ , \new_[11422]_ , \new_[11423]_ ,
    \new_[11426]_ , \new_[11430]_ , \new_[11431]_ , \new_[11432]_ ,
    \new_[11435]_ , \new_[11439]_ , \new_[11440]_ , \new_[11441]_ ,
    \new_[11444]_ , \new_[11448]_ , \new_[11449]_ , \new_[11450]_ ,
    \new_[11453]_ , \new_[11457]_ , \new_[11458]_ , \new_[11459]_ ,
    \new_[11462]_ , \new_[11466]_ , \new_[11467]_ , \new_[11468]_ ,
    \new_[11471]_ , \new_[11475]_ , \new_[11476]_ , \new_[11477]_ ,
    \new_[11480]_ , \new_[11484]_ , \new_[11485]_ , \new_[11486]_ ,
    \new_[11489]_ , \new_[11493]_ , \new_[11494]_ , \new_[11495]_ ,
    \new_[11498]_ , \new_[11502]_ , \new_[11503]_ , \new_[11504]_ ,
    \new_[11507]_ , \new_[11511]_ , \new_[11512]_ , \new_[11513]_ ,
    \new_[11516]_ , \new_[11520]_ , \new_[11521]_ , \new_[11522]_ ,
    \new_[11525]_ , \new_[11529]_ , \new_[11530]_ , \new_[11531]_ ,
    \new_[11534]_ , \new_[11538]_ , \new_[11539]_ , \new_[11540]_ ,
    \new_[11543]_ , \new_[11547]_ , \new_[11548]_ , \new_[11549]_ ,
    \new_[11552]_ , \new_[11556]_ , \new_[11557]_ , \new_[11558]_ ,
    \new_[11561]_ , \new_[11565]_ , \new_[11566]_ , \new_[11567]_ ,
    \new_[11570]_ , \new_[11574]_ , \new_[11575]_ , \new_[11576]_ ,
    \new_[11579]_ , \new_[11583]_ , \new_[11584]_ , \new_[11585]_ ,
    \new_[11588]_ , \new_[11592]_ , \new_[11593]_ , \new_[11594]_ ,
    \new_[11597]_ , \new_[11601]_ , \new_[11602]_ , \new_[11603]_ ,
    \new_[11606]_ , \new_[11610]_ , \new_[11611]_ , \new_[11612]_ ,
    \new_[11615]_ , \new_[11619]_ , \new_[11620]_ , \new_[11621]_ ,
    \new_[11624]_ , \new_[11628]_ , \new_[11629]_ , \new_[11630]_ ,
    \new_[11633]_ , \new_[11637]_ , \new_[11638]_ , \new_[11639]_ ,
    \new_[11642]_ , \new_[11646]_ , \new_[11647]_ , \new_[11648]_ ,
    \new_[11651]_ , \new_[11655]_ , \new_[11656]_ , \new_[11657]_ ,
    \new_[11660]_ , \new_[11664]_ , \new_[11665]_ , \new_[11666]_ ,
    \new_[11669]_ , \new_[11673]_ , \new_[11674]_ , \new_[11675]_ ,
    \new_[11678]_ , \new_[11682]_ , \new_[11683]_ , \new_[11684]_ ,
    \new_[11687]_ , \new_[11691]_ , \new_[11692]_ , \new_[11693]_ ,
    \new_[11696]_ , \new_[11700]_ , \new_[11701]_ , \new_[11702]_ ,
    \new_[11705]_ , \new_[11709]_ , \new_[11710]_ , \new_[11711]_ ,
    \new_[11714]_ , \new_[11718]_ , \new_[11719]_ , \new_[11720]_ ,
    \new_[11723]_ , \new_[11727]_ , \new_[11728]_ , \new_[11729]_ ,
    \new_[11732]_ , \new_[11736]_ , \new_[11737]_ , \new_[11738]_ ,
    \new_[11741]_ , \new_[11745]_ , \new_[11746]_ , \new_[11747]_ ,
    \new_[11750]_ , \new_[11754]_ , \new_[11755]_ , \new_[11756]_ ,
    \new_[11759]_ , \new_[11763]_ , \new_[11764]_ , \new_[11765]_ ,
    \new_[11768]_ , \new_[11772]_ , \new_[11773]_ , \new_[11774]_ ,
    \new_[11777]_ , \new_[11781]_ , \new_[11782]_ , \new_[11783]_ ,
    \new_[11786]_ , \new_[11790]_ , \new_[11791]_ , \new_[11792]_ ,
    \new_[11795]_ , \new_[11799]_ , \new_[11800]_ , \new_[11801]_ ,
    \new_[11804]_ , \new_[11808]_ , \new_[11809]_ , \new_[11810]_ ,
    \new_[11813]_ , \new_[11817]_ , \new_[11818]_ , \new_[11819]_ ,
    \new_[11822]_ , \new_[11826]_ , \new_[11827]_ , \new_[11828]_ ,
    \new_[11831]_ , \new_[11835]_ , \new_[11836]_ , \new_[11837]_ ,
    \new_[11840]_ , \new_[11844]_ , \new_[11845]_ , \new_[11846]_ ,
    \new_[11849]_ , \new_[11853]_ , \new_[11854]_ , \new_[11855]_ ,
    \new_[11858]_ , \new_[11862]_ , \new_[11863]_ , \new_[11864]_ ,
    \new_[11867]_ , \new_[11871]_ , \new_[11872]_ , \new_[11873]_ ,
    \new_[11876]_ , \new_[11880]_ , \new_[11881]_ , \new_[11882]_ ,
    \new_[11885]_ , \new_[11889]_ , \new_[11890]_ , \new_[11891]_ ,
    \new_[11894]_ , \new_[11898]_ , \new_[11899]_ , \new_[11900]_ ,
    \new_[11903]_ , \new_[11907]_ , \new_[11908]_ , \new_[11909]_ ,
    \new_[11912]_ , \new_[11916]_ , \new_[11917]_ , \new_[11918]_ ,
    \new_[11921]_ , \new_[11925]_ , \new_[11926]_ , \new_[11927]_ ,
    \new_[11930]_ , \new_[11934]_ , \new_[11935]_ , \new_[11936]_ ,
    \new_[11939]_ , \new_[11943]_ , \new_[11944]_ , \new_[11945]_ ,
    \new_[11948]_ , \new_[11952]_ , \new_[11953]_ , \new_[11954]_ ,
    \new_[11957]_ , \new_[11961]_ , \new_[11962]_ , \new_[11963]_ ,
    \new_[11966]_ , \new_[11970]_ , \new_[11971]_ , \new_[11972]_ ,
    \new_[11975]_ , \new_[11979]_ , \new_[11980]_ , \new_[11981]_ ,
    \new_[11984]_ , \new_[11988]_ , \new_[11989]_ , \new_[11990]_ ,
    \new_[11993]_ , \new_[11997]_ , \new_[11998]_ , \new_[11999]_ ,
    \new_[12002]_ , \new_[12006]_ , \new_[12007]_ , \new_[12008]_ ,
    \new_[12011]_ , \new_[12015]_ , \new_[12016]_ , \new_[12017]_ ,
    \new_[12020]_ , \new_[12024]_ , \new_[12025]_ , \new_[12026]_ ,
    \new_[12029]_ , \new_[12033]_ , \new_[12034]_ , \new_[12035]_ ,
    \new_[12038]_ , \new_[12042]_ , \new_[12043]_ , \new_[12044]_ ,
    \new_[12047]_ , \new_[12051]_ , \new_[12052]_ , \new_[12053]_ ,
    \new_[12056]_ , \new_[12060]_ , \new_[12061]_ , \new_[12062]_ ,
    \new_[12065]_ , \new_[12069]_ , \new_[12070]_ , \new_[12071]_ ,
    \new_[12074]_ , \new_[12078]_ , \new_[12079]_ , \new_[12080]_ ,
    \new_[12083]_ , \new_[12087]_ , \new_[12088]_ , \new_[12089]_ ,
    \new_[12092]_ , \new_[12096]_ , \new_[12097]_ , \new_[12098]_ ,
    \new_[12101]_ , \new_[12105]_ , \new_[12106]_ , \new_[12107]_ ,
    \new_[12110]_ , \new_[12114]_ , \new_[12115]_ , \new_[12116]_ ,
    \new_[12119]_ , \new_[12123]_ , \new_[12124]_ , \new_[12125]_ ,
    \new_[12128]_ , \new_[12132]_ , \new_[12133]_ , \new_[12134]_ ,
    \new_[12137]_ , \new_[12141]_ , \new_[12142]_ , \new_[12143]_ ,
    \new_[12146]_ , \new_[12150]_ , \new_[12151]_ , \new_[12152]_ ,
    \new_[12155]_ , \new_[12159]_ , \new_[12160]_ , \new_[12161]_ ,
    \new_[12164]_ , \new_[12168]_ , \new_[12169]_ , \new_[12170]_ ,
    \new_[12173]_ , \new_[12177]_ , \new_[12178]_ , \new_[12179]_ ,
    \new_[12182]_ , \new_[12186]_ , \new_[12187]_ , \new_[12188]_ ,
    \new_[12191]_ , \new_[12195]_ , \new_[12196]_ , \new_[12197]_ ,
    \new_[12200]_ , \new_[12204]_ , \new_[12205]_ , \new_[12206]_ ,
    \new_[12209]_ , \new_[12213]_ , \new_[12214]_ , \new_[12215]_ ,
    \new_[12218]_ , \new_[12222]_ , \new_[12223]_ , \new_[12224]_ ,
    \new_[12227]_ , \new_[12231]_ , \new_[12232]_ , \new_[12233]_ ,
    \new_[12236]_ , \new_[12240]_ , \new_[12241]_ , \new_[12242]_ ,
    \new_[12245]_ , \new_[12249]_ , \new_[12250]_ , \new_[12251]_ ,
    \new_[12254]_ , \new_[12258]_ , \new_[12259]_ , \new_[12260]_ ,
    \new_[12263]_ , \new_[12267]_ , \new_[12268]_ , \new_[12269]_ ,
    \new_[12272]_ , \new_[12276]_ , \new_[12277]_ , \new_[12278]_ ,
    \new_[12281]_ , \new_[12285]_ , \new_[12286]_ , \new_[12287]_ ,
    \new_[12290]_ , \new_[12294]_ , \new_[12295]_ , \new_[12296]_ ,
    \new_[12299]_ , \new_[12303]_ , \new_[12304]_ , \new_[12305]_ ,
    \new_[12308]_ , \new_[12312]_ , \new_[12313]_ , \new_[12314]_ ,
    \new_[12317]_ , \new_[12321]_ , \new_[12322]_ , \new_[12323]_ ,
    \new_[12326]_ , \new_[12330]_ , \new_[12331]_ , \new_[12332]_ ,
    \new_[12335]_ , \new_[12339]_ , \new_[12340]_ , \new_[12341]_ ,
    \new_[12344]_ , \new_[12348]_ , \new_[12349]_ , \new_[12350]_ ,
    \new_[12353]_ , \new_[12357]_ , \new_[12358]_ , \new_[12359]_ ,
    \new_[12362]_ , \new_[12366]_ , \new_[12367]_ , \new_[12368]_ ,
    \new_[12371]_ , \new_[12375]_ , \new_[12376]_ , \new_[12377]_ ,
    \new_[12380]_ , \new_[12384]_ , \new_[12385]_ , \new_[12386]_ ,
    \new_[12389]_ , \new_[12393]_ , \new_[12394]_ , \new_[12395]_ ,
    \new_[12398]_ , \new_[12402]_ , \new_[12403]_ , \new_[12404]_ ,
    \new_[12407]_ , \new_[12411]_ , \new_[12412]_ , \new_[12413]_ ,
    \new_[12416]_ , \new_[12420]_ , \new_[12421]_ , \new_[12422]_ ,
    \new_[12425]_ , \new_[12429]_ , \new_[12430]_ , \new_[12431]_ ,
    \new_[12434]_ , \new_[12438]_ , \new_[12439]_ , \new_[12440]_ ,
    \new_[12443]_ , \new_[12447]_ , \new_[12448]_ , \new_[12449]_ ,
    \new_[12452]_ , \new_[12456]_ , \new_[12457]_ , \new_[12458]_ ,
    \new_[12461]_ , \new_[12465]_ , \new_[12466]_ , \new_[12467]_ ,
    \new_[12470]_ , \new_[12474]_ , \new_[12475]_ , \new_[12476]_ ,
    \new_[12479]_ , \new_[12483]_ , \new_[12484]_ , \new_[12485]_ ,
    \new_[12488]_ , \new_[12492]_ , \new_[12493]_ , \new_[12494]_ ,
    \new_[12497]_ , \new_[12501]_ , \new_[12502]_ , \new_[12503]_ ,
    \new_[12506]_ , \new_[12510]_ , \new_[12511]_ , \new_[12512]_ ,
    \new_[12515]_ , \new_[12519]_ , \new_[12520]_ , \new_[12521]_ ,
    \new_[12524]_ , \new_[12528]_ , \new_[12529]_ , \new_[12530]_ ,
    \new_[12533]_ , \new_[12537]_ , \new_[12538]_ , \new_[12539]_ ,
    \new_[12542]_ , \new_[12546]_ , \new_[12547]_ , \new_[12548]_ ,
    \new_[12551]_ , \new_[12555]_ , \new_[12556]_ , \new_[12557]_ ,
    \new_[12560]_ , \new_[12564]_ , \new_[12565]_ , \new_[12566]_ ,
    \new_[12569]_ , \new_[12573]_ , \new_[12574]_ , \new_[12575]_ ,
    \new_[12578]_ , \new_[12582]_ , \new_[12583]_ , \new_[12584]_ ,
    \new_[12587]_ , \new_[12591]_ , \new_[12592]_ , \new_[12593]_ ,
    \new_[12596]_ , \new_[12600]_ , \new_[12601]_ , \new_[12602]_ ,
    \new_[12605]_ , \new_[12609]_ , \new_[12610]_ , \new_[12611]_ ,
    \new_[12614]_ , \new_[12618]_ , \new_[12619]_ , \new_[12620]_ ,
    \new_[12623]_ , \new_[12627]_ , \new_[12628]_ , \new_[12629]_ ,
    \new_[12632]_ , \new_[12636]_ , \new_[12637]_ , \new_[12638]_ ,
    \new_[12641]_ , \new_[12645]_ , \new_[12646]_ , \new_[12647]_ ,
    \new_[12650]_ , \new_[12654]_ , \new_[12655]_ , \new_[12656]_ ,
    \new_[12659]_ , \new_[12663]_ , \new_[12664]_ , \new_[12665]_ ,
    \new_[12668]_ , \new_[12672]_ , \new_[12673]_ , \new_[12674]_ ,
    \new_[12677]_ , \new_[12681]_ , \new_[12682]_ , \new_[12683]_ ,
    \new_[12686]_ , \new_[12690]_ , \new_[12691]_ , \new_[12692]_ ,
    \new_[12695]_ , \new_[12699]_ , \new_[12700]_ , \new_[12701]_ ,
    \new_[12704]_ , \new_[12708]_ , \new_[12709]_ , \new_[12710]_ ,
    \new_[12713]_ , \new_[12717]_ , \new_[12718]_ , \new_[12719]_ ,
    \new_[12722]_ , \new_[12726]_ , \new_[12727]_ , \new_[12728]_ ,
    \new_[12731]_ , \new_[12735]_ , \new_[12736]_ , \new_[12737]_ ,
    \new_[12740]_ , \new_[12744]_ , \new_[12745]_ , \new_[12746]_ ,
    \new_[12749]_ , \new_[12753]_ , \new_[12754]_ , \new_[12755]_ ,
    \new_[12758]_ , \new_[12762]_ , \new_[12763]_ , \new_[12764]_ ,
    \new_[12767]_ , \new_[12771]_ , \new_[12772]_ , \new_[12773]_ ,
    \new_[12776]_ , \new_[12780]_ , \new_[12781]_ , \new_[12782]_ ,
    \new_[12785]_ , \new_[12789]_ , \new_[12790]_ , \new_[12791]_ ,
    \new_[12794]_ , \new_[12798]_ , \new_[12799]_ , \new_[12800]_ ,
    \new_[12803]_ , \new_[12807]_ , \new_[12808]_ , \new_[12809]_ ,
    \new_[12812]_ , \new_[12816]_ , \new_[12817]_ , \new_[12818]_ ,
    \new_[12821]_ , \new_[12825]_ , \new_[12826]_ , \new_[12827]_ ,
    \new_[12830]_ , \new_[12834]_ , \new_[12835]_ , \new_[12836]_ ,
    \new_[12839]_ , \new_[12843]_ , \new_[12844]_ , \new_[12845]_ ,
    \new_[12848]_ , \new_[12852]_ , \new_[12853]_ , \new_[12854]_ ,
    \new_[12857]_ , \new_[12861]_ , \new_[12862]_ , \new_[12863]_ ,
    \new_[12866]_ , \new_[12870]_ , \new_[12871]_ , \new_[12872]_ ,
    \new_[12875]_ , \new_[12879]_ , \new_[12880]_ , \new_[12881]_ ,
    \new_[12884]_ , \new_[12888]_ , \new_[12889]_ , \new_[12890]_ ,
    \new_[12893]_ , \new_[12897]_ , \new_[12898]_ , \new_[12899]_ ,
    \new_[12902]_ , \new_[12906]_ , \new_[12907]_ , \new_[12908]_ ,
    \new_[12911]_ , \new_[12915]_ , \new_[12916]_ , \new_[12917]_ ,
    \new_[12920]_ , \new_[12924]_ , \new_[12925]_ , \new_[12926]_ ,
    \new_[12929]_ , \new_[12933]_ , \new_[12934]_ , \new_[12935]_ ,
    \new_[12938]_ , \new_[12942]_ , \new_[12943]_ , \new_[12944]_ ,
    \new_[12947]_ , \new_[12951]_ , \new_[12952]_ , \new_[12953]_ ,
    \new_[12956]_ , \new_[12960]_ , \new_[12961]_ , \new_[12962]_ ,
    \new_[12965]_ , \new_[12969]_ , \new_[12970]_ , \new_[12971]_ ,
    \new_[12974]_ , \new_[12978]_ , \new_[12979]_ , \new_[12980]_ ,
    \new_[12983]_ , \new_[12987]_ , \new_[12988]_ , \new_[12989]_ ,
    \new_[12992]_ , \new_[12996]_ , \new_[12997]_ , \new_[12998]_ ,
    \new_[13001]_ , \new_[13005]_ , \new_[13006]_ , \new_[13007]_ ,
    \new_[13010]_ , \new_[13014]_ , \new_[13015]_ , \new_[13016]_ ,
    \new_[13019]_ , \new_[13023]_ , \new_[13024]_ , \new_[13025]_ ,
    \new_[13028]_ , \new_[13032]_ , \new_[13033]_ , \new_[13034]_ ,
    \new_[13037]_ , \new_[13041]_ , \new_[13042]_ , \new_[13043]_ ,
    \new_[13046]_ , \new_[13050]_ , \new_[13051]_ , \new_[13052]_ ,
    \new_[13055]_ , \new_[13059]_ , \new_[13060]_ , \new_[13061]_ ,
    \new_[13064]_ , \new_[13068]_ , \new_[13069]_ , \new_[13070]_ ,
    \new_[13073]_ , \new_[13077]_ , \new_[13078]_ , \new_[13079]_ ,
    \new_[13082]_ , \new_[13086]_ , \new_[13087]_ , \new_[13088]_ ,
    \new_[13091]_ , \new_[13095]_ , \new_[13096]_ , \new_[13097]_ ,
    \new_[13100]_ , \new_[13104]_ , \new_[13105]_ , \new_[13106]_ ,
    \new_[13109]_ , \new_[13113]_ , \new_[13114]_ , \new_[13115]_ ,
    \new_[13118]_ , \new_[13122]_ , \new_[13123]_ , \new_[13124]_ ,
    \new_[13127]_ , \new_[13131]_ , \new_[13132]_ , \new_[13133]_ ,
    \new_[13136]_ , \new_[13140]_ , \new_[13141]_ , \new_[13142]_ ,
    \new_[13145]_ , \new_[13149]_ , \new_[13150]_ , \new_[13151]_ ,
    \new_[13154]_ , \new_[13158]_ , \new_[13159]_ , \new_[13160]_ ,
    \new_[13163]_ , \new_[13167]_ , \new_[13168]_ , \new_[13169]_ ,
    \new_[13172]_ , \new_[13176]_ , \new_[13177]_ , \new_[13178]_ ,
    \new_[13181]_ , \new_[13185]_ , \new_[13186]_ , \new_[13187]_ ,
    \new_[13190]_ , \new_[13194]_ , \new_[13195]_ , \new_[13196]_ ,
    \new_[13199]_ , \new_[13203]_ , \new_[13204]_ , \new_[13205]_ ,
    \new_[13208]_ , \new_[13212]_ , \new_[13213]_ , \new_[13214]_ ,
    \new_[13217]_ , \new_[13221]_ , \new_[13222]_ , \new_[13223]_ ,
    \new_[13226]_ , \new_[13230]_ , \new_[13231]_ , \new_[13232]_ ,
    \new_[13235]_ , \new_[13239]_ , \new_[13240]_ , \new_[13241]_ ,
    \new_[13244]_ , \new_[13248]_ , \new_[13249]_ , \new_[13250]_ ,
    \new_[13253]_ , \new_[13257]_ , \new_[13258]_ , \new_[13259]_ ,
    \new_[13262]_ , \new_[13266]_ , \new_[13267]_ , \new_[13268]_ ,
    \new_[13271]_ , \new_[13275]_ , \new_[13276]_ , \new_[13277]_ ,
    \new_[13280]_ , \new_[13284]_ , \new_[13285]_ , \new_[13286]_ ,
    \new_[13289]_ , \new_[13293]_ , \new_[13294]_ , \new_[13295]_ ,
    \new_[13298]_ , \new_[13302]_ , \new_[13303]_ , \new_[13304]_ ,
    \new_[13307]_ , \new_[13311]_ , \new_[13312]_ , \new_[13313]_ ,
    \new_[13316]_ , \new_[13320]_ , \new_[13321]_ , \new_[13322]_ ,
    \new_[13325]_ , \new_[13329]_ , \new_[13330]_ , \new_[13331]_ ,
    \new_[13334]_ , \new_[13338]_ , \new_[13339]_ , \new_[13340]_ ,
    \new_[13343]_ , \new_[13347]_ , \new_[13348]_ , \new_[13349]_ ,
    \new_[13352]_ , \new_[13356]_ , \new_[13357]_ , \new_[13358]_ ,
    \new_[13361]_ , \new_[13365]_ , \new_[13366]_ , \new_[13367]_ ,
    \new_[13370]_ , \new_[13374]_ , \new_[13375]_ , \new_[13376]_ ,
    \new_[13379]_ , \new_[13383]_ , \new_[13384]_ , \new_[13385]_ ,
    \new_[13388]_ , \new_[13392]_ , \new_[13393]_ , \new_[13394]_ ,
    \new_[13397]_ , \new_[13401]_ , \new_[13402]_ , \new_[13403]_ ,
    \new_[13406]_ , \new_[13410]_ , \new_[13411]_ , \new_[13412]_ ,
    \new_[13415]_ , \new_[13419]_ , \new_[13420]_ , \new_[13421]_ ,
    \new_[13424]_ , \new_[13428]_ , \new_[13429]_ , \new_[13430]_ ,
    \new_[13433]_ , \new_[13437]_ , \new_[13438]_ , \new_[13439]_ ,
    \new_[13442]_ , \new_[13446]_ , \new_[13447]_ , \new_[13448]_ ,
    \new_[13451]_ , \new_[13455]_ , \new_[13456]_ , \new_[13457]_ ,
    \new_[13460]_ , \new_[13464]_ , \new_[13465]_ , \new_[13466]_ ,
    \new_[13469]_ , \new_[13473]_ , \new_[13474]_ , \new_[13475]_ ,
    \new_[13478]_ , \new_[13482]_ , \new_[13483]_ , \new_[13484]_ ,
    \new_[13487]_ , \new_[13491]_ , \new_[13492]_ , \new_[13493]_ ,
    \new_[13496]_ , \new_[13500]_ , \new_[13501]_ , \new_[13502]_ ,
    \new_[13505]_ , \new_[13509]_ , \new_[13510]_ , \new_[13511]_ ,
    \new_[13514]_ , \new_[13518]_ , \new_[13519]_ , \new_[13520]_ ,
    \new_[13523]_ , \new_[13527]_ , \new_[13528]_ , \new_[13529]_ ,
    \new_[13532]_ , \new_[13536]_ , \new_[13537]_ , \new_[13538]_ ,
    \new_[13541]_ , \new_[13545]_ , \new_[13546]_ , \new_[13547]_ ,
    \new_[13550]_ , \new_[13554]_ , \new_[13555]_ , \new_[13556]_ ,
    \new_[13559]_ , \new_[13563]_ , \new_[13564]_ , \new_[13565]_ ,
    \new_[13568]_ , \new_[13572]_ , \new_[13573]_ , \new_[13574]_ ,
    \new_[13577]_ , \new_[13581]_ , \new_[13582]_ , \new_[13583]_ ,
    \new_[13586]_ , \new_[13590]_ , \new_[13591]_ , \new_[13592]_ ,
    \new_[13595]_ , \new_[13599]_ , \new_[13600]_ , \new_[13601]_ ,
    \new_[13604]_ , \new_[13608]_ , \new_[13609]_ , \new_[13610]_ ,
    \new_[13613]_ , \new_[13617]_ , \new_[13618]_ , \new_[13619]_ ,
    \new_[13622]_ , \new_[13626]_ , \new_[13627]_ , \new_[13628]_ ,
    \new_[13631]_ , \new_[13635]_ , \new_[13636]_ , \new_[13637]_ ,
    \new_[13641]_ , \new_[13642]_ , \new_[13646]_ , \new_[13647]_ ,
    \new_[13648]_ , \new_[13651]_ , \new_[13655]_ , \new_[13656]_ ,
    \new_[13657]_ , \new_[13661]_ , \new_[13662]_ , \new_[13666]_ ,
    \new_[13667]_ , \new_[13668]_ , \new_[13671]_ , \new_[13675]_ ,
    \new_[13676]_ , \new_[13677]_ , \new_[13681]_ , \new_[13682]_ ,
    \new_[13686]_ , \new_[13687]_ , \new_[13688]_ , \new_[13691]_ ,
    \new_[13695]_ , \new_[13696]_ , \new_[13697]_ , \new_[13701]_ ,
    \new_[13702]_ , \new_[13706]_ , \new_[13707]_ , \new_[13708]_ ,
    \new_[13711]_ , \new_[13715]_ , \new_[13716]_ , \new_[13717]_ ,
    \new_[13721]_ , \new_[13722]_ , \new_[13726]_ , \new_[13727]_ ,
    \new_[13728]_ , \new_[13731]_ , \new_[13735]_ , \new_[13736]_ ,
    \new_[13737]_ , \new_[13741]_ , \new_[13742]_ , \new_[13746]_ ,
    \new_[13747]_ , \new_[13748]_ , \new_[13751]_ , \new_[13755]_ ,
    \new_[13756]_ , \new_[13757]_ , \new_[13761]_ , \new_[13762]_ ,
    \new_[13766]_ , \new_[13767]_ , \new_[13768]_ , \new_[13771]_ ,
    \new_[13775]_ , \new_[13776]_ , \new_[13777]_ , \new_[13781]_ ,
    \new_[13782]_ , \new_[13786]_ , \new_[13787]_ , \new_[13788]_ ,
    \new_[13791]_ , \new_[13795]_ , \new_[13796]_ , \new_[13797]_ ,
    \new_[13801]_ , \new_[13802]_ , \new_[13806]_ , \new_[13807]_ ,
    \new_[13808]_ , \new_[13811]_ , \new_[13815]_ , \new_[13816]_ ,
    \new_[13817]_ , \new_[13821]_ , \new_[13822]_ , \new_[13826]_ ,
    \new_[13827]_ , \new_[13828]_ , \new_[13831]_ , \new_[13835]_ ,
    \new_[13836]_ , \new_[13837]_ , \new_[13841]_ , \new_[13842]_ ,
    \new_[13846]_ , \new_[13847]_ , \new_[13848]_ , \new_[13851]_ ,
    \new_[13855]_ , \new_[13856]_ , \new_[13857]_ , \new_[13861]_ ,
    \new_[13862]_ , \new_[13866]_ , \new_[13867]_ , \new_[13868]_ ,
    \new_[13871]_ , \new_[13875]_ , \new_[13876]_ , \new_[13877]_ ,
    \new_[13881]_ , \new_[13882]_ , \new_[13886]_ , \new_[13887]_ ,
    \new_[13888]_ , \new_[13891]_ , \new_[13895]_ , \new_[13896]_ ,
    \new_[13897]_ , \new_[13901]_ , \new_[13902]_ , \new_[13906]_ ,
    \new_[13907]_ , \new_[13908]_ , \new_[13911]_ , \new_[13915]_ ,
    \new_[13916]_ , \new_[13917]_ , \new_[13921]_ , \new_[13922]_ ,
    \new_[13926]_ , \new_[13927]_ , \new_[13928]_ , \new_[13931]_ ,
    \new_[13935]_ , \new_[13936]_ , \new_[13937]_ , \new_[13941]_ ,
    \new_[13942]_ , \new_[13946]_ , \new_[13947]_ , \new_[13948]_ ,
    \new_[13951]_ , \new_[13955]_ , \new_[13956]_ , \new_[13957]_ ,
    \new_[13961]_ , \new_[13962]_ , \new_[13966]_ , \new_[13967]_ ,
    \new_[13968]_ , \new_[13971]_ , \new_[13975]_ , \new_[13976]_ ,
    \new_[13977]_ , \new_[13981]_ , \new_[13982]_ , \new_[13986]_ ,
    \new_[13987]_ , \new_[13988]_ , \new_[13991]_ , \new_[13995]_ ,
    \new_[13996]_ , \new_[13997]_ , \new_[14001]_ , \new_[14002]_ ,
    \new_[14006]_ , \new_[14007]_ , \new_[14008]_ , \new_[14011]_ ,
    \new_[14015]_ , \new_[14016]_ , \new_[14017]_ , \new_[14021]_ ,
    \new_[14022]_ , \new_[14026]_ , \new_[14027]_ , \new_[14028]_ ,
    \new_[14031]_ , \new_[14035]_ , \new_[14036]_ , \new_[14037]_ ,
    \new_[14041]_ , \new_[14042]_ , \new_[14046]_ , \new_[14047]_ ,
    \new_[14048]_ , \new_[14051]_ , \new_[14055]_ , \new_[14056]_ ,
    \new_[14057]_ , \new_[14061]_ , \new_[14062]_ , \new_[14066]_ ,
    \new_[14067]_ , \new_[14068]_ , \new_[14071]_ , \new_[14075]_ ,
    \new_[14076]_ , \new_[14077]_ , \new_[14081]_ , \new_[14082]_ ,
    \new_[14086]_ , \new_[14087]_ , \new_[14088]_ , \new_[14091]_ ,
    \new_[14095]_ , \new_[14096]_ , \new_[14097]_ , \new_[14101]_ ,
    \new_[14102]_ , \new_[14106]_ , \new_[14107]_ , \new_[14108]_ ,
    \new_[14111]_ , \new_[14115]_ , \new_[14116]_ , \new_[14117]_ ,
    \new_[14121]_ , \new_[14122]_ , \new_[14126]_ , \new_[14127]_ ,
    \new_[14128]_ , \new_[14131]_ , \new_[14135]_ , \new_[14136]_ ,
    \new_[14137]_ , \new_[14141]_ , \new_[14142]_ , \new_[14146]_ ,
    \new_[14147]_ , \new_[14148]_ , \new_[14151]_ , \new_[14155]_ ,
    \new_[14156]_ , \new_[14157]_ , \new_[14161]_ , \new_[14162]_ ,
    \new_[14166]_ , \new_[14167]_ , \new_[14168]_ , \new_[14171]_ ,
    \new_[14175]_ , \new_[14176]_ , \new_[14177]_ , \new_[14181]_ ,
    \new_[14182]_ , \new_[14186]_ , \new_[14187]_ , \new_[14188]_ ,
    \new_[14191]_ , \new_[14195]_ , \new_[14196]_ , \new_[14197]_ ,
    \new_[14201]_ , \new_[14202]_ , \new_[14206]_ , \new_[14207]_ ,
    \new_[14208]_ , \new_[14211]_ , \new_[14215]_ , \new_[14216]_ ,
    \new_[14217]_ , \new_[14221]_ , \new_[14222]_ , \new_[14226]_ ,
    \new_[14227]_ , \new_[14228]_ , \new_[14231]_ , \new_[14235]_ ,
    \new_[14236]_ , \new_[14237]_ , \new_[14241]_ , \new_[14242]_ ,
    \new_[14246]_ , \new_[14247]_ , \new_[14248]_ , \new_[14251]_ ,
    \new_[14255]_ , \new_[14256]_ , \new_[14257]_ , \new_[14261]_ ,
    \new_[14262]_ , \new_[14266]_ , \new_[14267]_ , \new_[14268]_ ,
    \new_[14271]_ , \new_[14275]_ , \new_[14276]_ , \new_[14277]_ ,
    \new_[14281]_ , \new_[14282]_ , \new_[14286]_ , \new_[14287]_ ,
    \new_[14288]_ , \new_[14291]_ , \new_[14295]_ , \new_[14296]_ ,
    \new_[14297]_ , \new_[14301]_ , \new_[14302]_ , \new_[14306]_ ,
    \new_[14307]_ , \new_[14308]_ , \new_[14311]_ , \new_[14315]_ ,
    \new_[14316]_ , \new_[14317]_ , \new_[14321]_ , \new_[14322]_ ,
    \new_[14326]_ , \new_[14327]_ , \new_[14328]_ , \new_[14331]_ ,
    \new_[14335]_ , \new_[14336]_ , \new_[14337]_ , \new_[14341]_ ,
    \new_[14342]_ , \new_[14346]_ , \new_[14347]_ , \new_[14348]_ ,
    \new_[14351]_ , \new_[14355]_ , \new_[14356]_ , \new_[14357]_ ,
    \new_[14361]_ , \new_[14362]_ , \new_[14366]_ , \new_[14367]_ ,
    \new_[14368]_ , \new_[14371]_ , \new_[14375]_ , \new_[14376]_ ,
    \new_[14377]_ , \new_[14381]_ , \new_[14382]_ , \new_[14386]_ ,
    \new_[14387]_ , \new_[14388]_ , \new_[14391]_ , \new_[14395]_ ,
    \new_[14396]_ , \new_[14397]_ , \new_[14401]_ , \new_[14402]_ ,
    \new_[14406]_ , \new_[14407]_ , \new_[14408]_ , \new_[14411]_ ,
    \new_[14415]_ , \new_[14416]_ , \new_[14417]_ , \new_[14421]_ ,
    \new_[14422]_ , \new_[14426]_ , \new_[14427]_ , \new_[14428]_ ,
    \new_[14431]_ , \new_[14435]_ , \new_[14436]_ , \new_[14437]_ ,
    \new_[14441]_ , \new_[14442]_ , \new_[14446]_ , \new_[14447]_ ,
    \new_[14448]_ , \new_[14451]_ , \new_[14455]_ , \new_[14456]_ ,
    \new_[14457]_ , \new_[14461]_ , \new_[14462]_ , \new_[14466]_ ,
    \new_[14467]_ , \new_[14468]_ , \new_[14471]_ , \new_[14475]_ ,
    \new_[14476]_ , \new_[14477]_ , \new_[14481]_ , \new_[14482]_ ,
    \new_[14486]_ , \new_[14487]_ , \new_[14488]_ , \new_[14491]_ ,
    \new_[14495]_ , \new_[14496]_ , \new_[14497]_ , \new_[14501]_ ,
    \new_[14502]_ , \new_[14506]_ , \new_[14507]_ , \new_[14508]_ ,
    \new_[14511]_ , \new_[14515]_ , \new_[14516]_ , \new_[14517]_ ,
    \new_[14521]_ , \new_[14522]_ , \new_[14526]_ , \new_[14527]_ ,
    \new_[14528]_ , \new_[14531]_ , \new_[14535]_ , \new_[14536]_ ,
    \new_[14537]_ , \new_[14541]_ , \new_[14542]_ , \new_[14546]_ ,
    \new_[14547]_ , \new_[14548]_ , \new_[14551]_ , \new_[14555]_ ,
    \new_[14556]_ , \new_[14557]_ , \new_[14561]_ , \new_[14562]_ ,
    \new_[14566]_ , \new_[14567]_ , \new_[14568]_ , \new_[14571]_ ,
    \new_[14575]_ , \new_[14576]_ , \new_[14577]_ , \new_[14581]_ ,
    \new_[14582]_ , \new_[14586]_ , \new_[14587]_ , \new_[14588]_ ,
    \new_[14591]_ , \new_[14595]_ , \new_[14596]_ , \new_[14597]_ ,
    \new_[14601]_ , \new_[14602]_ , \new_[14606]_ , \new_[14607]_ ,
    \new_[14608]_ , \new_[14611]_ , \new_[14615]_ , \new_[14616]_ ,
    \new_[14617]_ , \new_[14621]_ , \new_[14622]_ , \new_[14626]_ ,
    \new_[14627]_ , \new_[14628]_ , \new_[14631]_ , \new_[14635]_ ,
    \new_[14636]_ , \new_[14637]_ , \new_[14641]_ , \new_[14642]_ ,
    \new_[14646]_ , \new_[14647]_ , \new_[14648]_ , \new_[14651]_ ,
    \new_[14655]_ , \new_[14656]_ , \new_[14657]_ , \new_[14661]_ ,
    \new_[14662]_ , \new_[14666]_ , \new_[14667]_ , \new_[14668]_ ,
    \new_[14671]_ , \new_[14675]_ , \new_[14676]_ , \new_[14677]_ ,
    \new_[14681]_ , \new_[14682]_ , \new_[14686]_ , \new_[14687]_ ,
    \new_[14688]_ , \new_[14691]_ , \new_[14695]_ , \new_[14696]_ ,
    \new_[14697]_ , \new_[14701]_ , \new_[14702]_ , \new_[14706]_ ,
    \new_[14707]_ , \new_[14708]_ , \new_[14711]_ , \new_[14715]_ ,
    \new_[14716]_ , \new_[14717]_ , \new_[14721]_ , \new_[14722]_ ,
    \new_[14726]_ , \new_[14727]_ , \new_[14728]_ , \new_[14731]_ ,
    \new_[14735]_ , \new_[14736]_ , \new_[14737]_ , \new_[14741]_ ,
    \new_[14742]_ , \new_[14746]_ , \new_[14747]_ , \new_[14748]_ ,
    \new_[14751]_ , \new_[14755]_ , \new_[14756]_ , \new_[14757]_ ,
    \new_[14761]_ , \new_[14762]_ , \new_[14766]_ , \new_[14767]_ ,
    \new_[14768]_ , \new_[14771]_ , \new_[14775]_ , \new_[14776]_ ,
    \new_[14777]_ , \new_[14781]_ , \new_[14782]_ , \new_[14786]_ ,
    \new_[14787]_ , \new_[14788]_ , \new_[14791]_ , \new_[14795]_ ,
    \new_[14796]_ , \new_[14797]_ , \new_[14801]_ , \new_[14802]_ ,
    \new_[14806]_ , \new_[14807]_ , \new_[14808]_ , \new_[14811]_ ,
    \new_[14815]_ , \new_[14816]_ , \new_[14817]_ , \new_[14821]_ ,
    \new_[14822]_ , \new_[14826]_ , \new_[14827]_ , \new_[14828]_ ,
    \new_[14831]_ , \new_[14835]_ , \new_[14836]_ , \new_[14837]_ ,
    \new_[14841]_ , \new_[14842]_ , \new_[14846]_ , \new_[14847]_ ,
    \new_[14848]_ , \new_[14851]_ , \new_[14855]_ , \new_[14856]_ ,
    \new_[14857]_ , \new_[14861]_ , \new_[14862]_ , \new_[14866]_ ,
    \new_[14867]_ , \new_[14868]_ , \new_[14871]_ , \new_[14875]_ ,
    \new_[14876]_ , \new_[14877]_ , \new_[14881]_ , \new_[14882]_ ,
    \new_[14886]_ , \new_[14887]_ , \new_[14888]_ , \new_[14891]_ ,
    \new_[14895]_ , \new_[14896]_ , \new_[14897]_ , \new_[14901]_ ,
    \new_[14902]_ , \new_[14906]_ , \new_[14907]_ , \new_[14908]_ ,
    \new_[14911]_ , \new_[14915]_ , \new_[14916]_ , \new_[14917]_ ,
    \new_[14921]_ , \new_[14922]_ , \new_[14926]_ , \new_[14927]_ ,
    \new_[14928]_ , \new_[14931]_ , \new_[14935]_ , \new_[14936]_ ,
    \new_[14937]_ , \new_[14941]_ , \new_[14942]_ , \new_[14946]_ ,
    \new_[14947]_ , \new_[14948]_ , \new_[14951]_ , \new_[14955]_ ,
    \new_[14956]_ , \new_[14957]_ , \new_[14961]_ , \new_[14962]_ ,
    \new_[14966]_ , \new_[14967]_ , \new_[14968]_ , \new_[14971]_ ,
    \new_[14975]_ , \new_[14976]_ , \new_[14977]_ , \new_[14981]_ ,
    \new_[14982]_ , \new_[14986]_ , \new_[14987]_ , \new_[14988]_ ,
    \new_[14991]_ , \new_[14995]_ , \new_[14996]_ , \new_[14997]_ ,
    \new_[15001]_ , \new_[15002]_ , \new_[15006]_ , \new_[15007]_ ,
    \new_[15008]_ , \new_[15011]_ , \new_[15015]_ , \new_[15016]_ ,
    \new_[15017]_ , \new_[15021]_ , \new_[15022]_ , \new_[15026]_ ,
    \new_[15027]_ , \new_[15028]_ , \new_[15031]_ , \new_[15035]_ ,
    \new_[15036]_ , \new_[15037]_ , \new_[15041]_ , \new_[15042]_ ,
    \new_[15046]_ , \new_[15047]_ , \new_[15048]_ , \new_[15051]_ ,
    \new_[15055]_ , \new_[15056]_ , \new_[15057]_ , \new_[15061]_ ,
    \new_[15062]_ , \new_[15066]_ , \new_[15067]_ , \new_[15068]_ ,
    \new_[15071]_ , \new_[15075]_ , \new_[15076]_ , \new_[15077]_ ,
    \new_[15081]_ , \new_[15082]_ , \new_[15086]_ , \new_[15087]_ ,
    \new_[15088]_ , \new_[15091]_ , \new_[15095]_ , \new_[15096]_ ,
    \new_[15097]_ , \new_[15101]_ , \new_[15102]_ , \new_[15106]_ ,
    \new_[15107]_ , \new_[15108]_ , \new_[15111]_ , \new_[15115]_ ,
    \new_[15116]_ , \new_[15117]_ , \new_[15121]_ , \new_[15122]_ ,
    \new_[15126]_ , \new_[15127]_ , \new_[15128]_ , \new_[15131]_ ,
    \new_[15135]_ , \new_[15136]_ , \new_[15137]_ , \new_[15141]_ ,
    \new_[15142]_ , \new_[15146]_ , \new_[15147]_ , \new_[15148]_ ,
    \new_[15151]_ , \new_[15155]_ , \new_[15156]_ , \new_[15157]_ ,
    \new_[15161]_ , \new_[15162]_ , \new_[15166]_ , \new_[15167]_ ,
    \new_[15168]_ , \new_[15171]_ , \new_[15175]_ , \new_[15176]_ ,
    \new_[15177]_ , \new_[15181]_ , \new_[15182]_ , \new_[15186]_ ,
    \new_[15187]_ , \new_[15188]_ , \new_[15191]_ , \new_[15195]_ ,
    \new_[15196]_ , \new_[15197]_ , \new_[15201]_ , \new_[15202]_ ,
    \new_[15206]_ , \new_[15207]_ , \new_[15208]_ , \new_[15211]_ ,
    \new_[15215]_ , \new_[15216]_ , \new_[15217]_ , \new_[15221]_ ,
    \new_[15222]_ , \new_[15226]_ , \new_[15227]_ , \new_[15228]_ ,
    \new_[15231]_ , \new_[15235]_ , \new_[15236]_ , \new_[15237]_ ,
    \new_[15241]_ , \new_[15242]_ , \new_[15246]_ , \new_[15247]_ ,
    \new_[15248]_ , \new_[15251]_ , \new_[15255]_ , \new_[15256]_ ,
    \new_[15257]_ , \new_[15261]_ , \new_[15262]_ , \new_[15266]_ ,
    \new_[15267]_ , \new_[15268]_ , \new_[15271]_ , \new_[15275]_ ,
    \new_[15276]_ , \new_[15277]_ , \new_[15281]_ , \new_[15282]_ ,
    \new_[15286]_ , \new_[15287]_ , \new_[15288]_ , \new_[15291]_ ,
    \new_[15295]_ , \new_[15296]_ , \new_[15297]_ , \new_[15301]_ ,
    \new_[15302]_ , \new_[15306]_ , \new_[15307]_ , \new_[15308]_ ,
    \new_[15311]_ , \new_[15315]_ , \new_[15316]_ , \new_[15317]_ ,
    \new_[15321]_ , \new_[15322]_ , \new_[15326]_ , \new_[15327]_ ,
    \new_[15328]_ , \new_[15331]_ , \new_[15335]_ , \new_[15336]_ ,
    \new_[15337]_ , \new_[15341]_ , \new_[15342]_ , \new_[15346]_ ,
    \new_[15347]_ , \new_[15348]_ , \new_[15351]_ , \new_[15355]_ ,
    \new_[15356]_ , \new_[15357]_ , \new_[15361]_ , \new_[15362]_ ,
    \new_[15366]_ , \new_[15367]_ , \new_[15368]_ , \new_[15371]_ ,
    \new_[15375]_ , \new_[15376]_ , \new_[15377]_ , \new_[15381]_ ,
    \new_[15382]_ , \new_[15386]_ , \new_[15387]_ , \new_[15388]_ ,
    \new_[15391]_ , \new_[15395]_ , \new_[15396]_ , \new_[15397]_ ,
    \new_[15401]_ , \new_[15402]_ , \new_[15406]_ , \new_[15407]_ ,
    \new_[15408]_ , \new_[15411]_ , \new_[15415]_ , \new_[15416]_ ,
    \new_[15417]_ , \new_[15421]_ , \new_[15422]_ , \new_[15426]_ ,
    \new_[15427]_ , \new_[15428]_ , \new_[15431]_ , \new_[15435]_ ,
    \new_[15436]_ , \new_[15437]_ , \new_[15441]_ , \new_[15442]_ ,
    \new_[15446]_ , \new_[15447]_ , \new_[15448]_ , \new_[15451]_ ,
    \new_[15455]_ , \new_[15456]_ , \new_[15457]_ , \new_[15461]_ ,
    \new_[15462]_ , \new_[15466]_ , \new_[15467]_ , \new_[15468]_ ,
    \new_[15471]_ , \new_[15475]_ , \new_[15476]_ , \new_[15477]_ ,
    \new_[15481]_ , \new_[15482]_ , \new_[15486]_ , \new_[15487]_ ,
    \new_[15488]_ , \new_[15491]_ , \new_[15495]_ , \new_[15496]_ ,
    \new_[15497]_ , \new_[15501]_ , \new_[15502]_ , \new_[15506]_ ,
    \new_[15507]_ , \new_[15508]_ , \new_[15511]_ , \new_[15515]_ ,
    \new_[15516]_ , \new_[15517]_ , \new_[15521]_ , \new_[15522]_ ,
    \new_[15526]_ , \new_[15527]_ , \new_[15528]_ , \new_[15531]_ ,
    \new_[15535]_ , \new_[15536]_ , \new_[15537]_ , \new_[15541]_ ,
    \new_[15542]_ , \new_[15546]_ , \new_[15547]_ , \new_[15548]_ ,
    \new_[15551]_ , \new_[15555]_ , \new_[15556]_ , \new_[15557]_ ,
    \new_[15561]_ , \new_[15562]_ , \new_[15566]_ , \new_[15567]_ ,
    \new_[15568]_ , \new_[15571]_ , \new_[15575]_ , \new_[15576]_ ,
    \new_[15577]_ , \new_[15581]_ , \new_[15582]_ , \new_[15586]_ ,
    \new_[15587]_ , \new_[15588]_ , \new_[15591]_ , \new_[15595]_ ,
    \new_[15596]_ , \new_[15597]_ , \new_[15601]_ , \new_[15602]_ ,
    \new_[15606]_ , \new_[15607]_ , \new_[15608]_ , \new_[15611]_ ,
    \new_[15615]_ , \new_[15616]_ , \new_[15617]_ , \new_[15621]_ ,
    \new_[15622]_ , \new_[15626]_ , \new_[15627]_ , \new_[15628]_ ,
    \new_[15631]_ , \new_[15635]_ , \new_[15636]_ , \new_[15637]_ ,
    \new_[15641]_ , \new_[15642]_ , \new_[15646]_ , \new_[15647]_ ,
    \new_[15648]_ , \new_[15651]_ , \new_[15655]_ , \new_[15656]_ ,
    \new_[15657]_ , \new_[15661]_ , \new_[15662]_ , \new_[15666]_ ,
    \new_[15667]_ , \new_[15668]_ , \new_[15671]_ , \new_[15675]_ ,
    \new_[15676]_ , \new_[15677]_ , \new_[15681]_ , \new_[15682]_ ,
    \new_[15686]_ , \new_[15687]_ , \new_[15688]_ , \new_[15691]_ ,
    \new_[15695]_ , \new_[15696]_ , \new_[15697]_ , \new_[15701]_ ,
    \new_[15702]_ , \new_[15706]_ , \new_[15707]_ , \new_[15708]_ ,
    \new_[15711]_ , \new_[15715]_ , \new_[15716]_ , \new_[15717]_ ,
    \new_[15721]_ , \new_[15722]_ , \new_[15726]_ , \new_[15727]_ ,
    \new_[15728]_ , \new_[15731]_ , \new_[15735]_ , \new_[15736]_ ,
    \new_[15737]_ , \new_[15741]_ , \new_[15742]_ , \new_[15746]_ ,
    \new_[15747]_ , \new_[15748]_ , \new_[15751]_ , \new_[15755]_ ,
    \new_[15756]_ , \new_[15757]_ , \new_[15761]_ , \new_[15762]_ ,
    \new_[15766]_ , \new_[15767]_ , \new_[15768]_ , \new_[15771]_ ,
    \new_[15775]_ , \new_[15776]_ , \new_[15777]_ , \new_[15781]_ ,
    \new_[15782]_ , \new_[15786]_ , \new_[15787]_ , \new_[15788]_ ,
    \new_[15791]_ , \new_[15795]_ , \new_[15796]_ , \new_[15797]_ ,
    \new_[15801]_ , \new_[15802]_ , \new_[15806]_ , \new_[15807]_ ,
    \new_[15808]_ , \new_[15811]_ , \new_[15815]_ , \new_[15816]_ ,
    \new_[15817]_ , \new_[15821]_ , \new_[15822]_ , \new_[15826]_ ,
    \new_[15827]_ , \new_[15828]_ , \new_[15831]_ , \new_[15835]_ ,
    \new_[15836]_ , \new_[15837]_ , \new_[15841]_ , \new_[15842]_ ,
    \new_[15846]_ , \new_[15847]_ , \new_[15848]_ , \new_[15851]_ ,
    \new_[15855]_ , \new_[15856]_ , \new_[15857]_ , \new_[15861]_ ,
    \new_[15862]_ , \new_[15866]_ , \new_[15867]_ , \new_[15868]_ ,
    \new_[15871]_ , \new_[15875]_ , \new_[15876]_ , \new_[15877]_ ,
    \new_[15881]_ , \new_[15882]_ , \new_[15886]_ , \new_[15887]_ ,
    \new_[15888]_ , \new_[15891]_ , \new_[15895]_ , \new_[15896]_ ,
    \new_[15897]_ , \new_[15901]_ , \new_[15902]_ , \new_[15906]_ ,
    \new_[15907]_ , \new_[15908]_ , \new_[15911]_ , \new_[15915]_ ,
    \new_[15916]_ , \new_[15917]_ , \new_[15921]_ , \new_[15922]_ ,
    \new_[15926]_ , \new_[15927]_ , \new_[15928]_ , \new_[15931]_ ,
    \new_[15935]_ , \new_[15936]_ , \new_[15937]_ , \new_[15941]_ ,
    \new_[15942]_ , \new_[15946]_ , \new_[15947]_ , \new_[15948]_ ,
    \new_[15951]_ , \new_[15955]_ , \new_[15956]_ , \new_[15957]_ ,
    \new_[15961]_ , \new_[15962]_ , \new_[15966]_ , \new_[15967]_ ,
    \new_[15968]_ , \new_[15971]_ , \new_[15975]_ , \new_[15976]_ ,
    \new_[15977]_ , \new_[15981]_ , \new_[15982]_ , \new_[15986]_ ,
    \new_[15987]_ , \new_[15988]_ , \new_[15991]_ , \new_[15995]_ ,
    \new_[15996]_ , \new_[15997]_ , \new_[16001]_ , \new_[16002]_ ,
    \new_[16006]_ , \new_[16007]_ , \new_[16008]_ , \new_[16011]_ ,
    \new_[16015]_ , \new_[16016]_ , \new_[16017]_ , \new_[16021]_ ,
    \new_[16022]_ , \new_[16026]_ , \new_[16027]_ , \new_[16028]_ ,
    \new_[16031]_ , \new_[16035]_ , \new_[16036]_ , \new_[16037]_ ,
    \new_[16041]_ , \new_[16042]_ , \new_[16046]_ , \new_[16047]_ ,
    \new_[16048]_ , \new_[16051]_ , \new_[16055]_ , \new_[16056]_ ,
    \new_[16057]_ , \new_[16061]_ , \new_[16062]_ , \new_[16066]_ ,
    \new_[16067]_ , \new_[16068]_ , \new_[16071]_ , \new_[16075]_ ,
    \new_[16076]_ , \new_[16077]_ , \new_[16081]_ , \new_[16082]_ ,
    \new_[16086]_ , \new_[16087]_ , \new_[16088]_ , \new_[16091]_ ,
    \new_[16095]_ , \new_[16096]_ , \new_[16097]_ , \new_[16101]_ ,
    \new_[16102]_ , \new_[16106]_ , \new_[16107]_ , \new_[16108]_ ,
    \new_[16111]_ , \new_[16115]_ , \new_[16116]_ , \new_[16117]_ ,
    \new_[16121]_ , \new_[16122]_ , \new_[16126]_ , \new_[16127]_ ,
    \new_[16128]_ , \new_[16131]_ , \new_[16135]_ , \new_[16136]_ ,
    \new_[16137]_ , \new_[16141]_ , \new_[16142]_ , \new_[16146]_ ,
    \new_[16147]_ , \new_[16148]_ , \new_[16151]_ , \new_[16155]_ ,
    \new_[16156]_ , \new_[16157]_ , \new_[16161]_ , \new_[16162]_ ,
    \new_[16166]_ , \new_[16167]_ , \new_[16168]_ , \new_[16171]_ ,
    \new_[16175]_ , \new_[16176]_ , \new_[16177]_ , \new_[16181]_ ,
    \new_[16182]_ , \new_[16186]_ , \new_[16187]_ , \new_[16188]_ ,
    \new_[16191]_ , \new_[16195]_ , \new_[16196]_ , \new_[16197]_ ,
    \new_[16201]_ , \new_[16202]_ , \new_[16206]_ , \new_[16207]_ ,
    \new_[16208]_ , \new_[16211]_ , \new_[16215]_ , \new_[16216]_ ,
    \new_[16217]_ , \new_[16221]_ , \new_[16222]_ , \new_[16226]_ ,
    \new_[16227]_ , \new_[16228]_ , \new_[16231]_ , \new_[16235]_ ,
    \new_[16236]_ , \new_[16237]_ , \new_[16241]_ , \new_[16242]_ ,
    \new_[16246]_ , \new_[16247]_ , \new_[16248]_ , \new_[16251]_ ,
    \new_[16255]_ , \new_[16256]_ , \new_[16257]_ , \new_[16261]_ ,
    \new_[16262]_ , \new_[16266]_ , \new_[16267]_ , \new_[16268]_ ,
    \new_[16271]_ , \new_[16275]_ , \new_[16276]_ , \new_[16277]_ ,
    \new_[16281]_ , \new_[16282]_ , \new_[16286]_ , \new_[16287]_ ,
    \new_[16288]_ , \new_[16291]_ , \new_[16295]_ , \new_[16296]_ ,
    \new_[16297]_ , \new_[16301]_ , \new_[16302]_ , \new_[16306]_ ,
    \new_[16307]_ , \new_[16308]_ , \new_[16311]_ , \new_[16315]_ ,
    \new_[16316]_ , \new_[16317]_ , \new_[16321]_ , \new_[16322]_ ,
    \new_[16326]_ , \new_[16327]_ , \new_[16328]_ , \new_[16331]_ ,
    \new_[16335]_ , \new_[16336]_ , \new_[16337]_ , \new_[16341]_ ,
    \new_[16342]_ , \new_[16346]_ , \new_[16347]_ , \new_[16348]_ ,
    \new_[16351]_ , \new_[16355]_ , \new_[16356]_ , \new_[16357]_ ,
    \new_[16361]_ , \new_[16362]_ , \new_[16366]_ , \new_[16367]_ ,
    \new_[16368]_ , \new_[16371]_ , \new_[16375]_ , \new_[16376]_ ,
    \new_[16377]_ , \new_[16381]_ , \new_[16382]_ , \new_[16386]_ ,
    \new_[16387]_ , \new_[16388]_ , \new_[16391]_ , \new_[16395]_ ,
    \new_[16396]_ , \new_[16397]_ , \new_[16401]_ , \new_[16402]_ ,
    \new_[16406]_ , \new_[16407]_ , \new_[16408]_ , \new_[16411]_ ,
    \new_[16415]_ , \new_[16416]_ , \new_[16417]_ , \new_[16421]_ ,
    \new_[16422]_ , \new_[16426]_ , \new_[16427]_ , \new_[16428]_ ,
    \new_[16431]_ , \new_[16435]_ , \new_[16436]_ , \new_[16437]_ ,
    \new_[16441]_ , \new_[16442]_ , \new_[16446]_ , \new_[16447]_ ,
    \new_[16448]_ , \new_[16451]_ , \new_[16455]_ , \new_[16456]_ ,
    \new_[16457]_ , \new_[16461]_ , \new_[16462]_ , \new_[16466]_ ,
    \new_[16467]_ , \new_[16468]_ , \new_[16471]_ , \new_[16475]_ ,
    \new_[16476]_ , \new_[16477]_ , \new_[16481]_ , \new_[16482]_ ,
    \new_[16486]_ , \new_[16487]_ , \new_[16488]_ , \new_[16491]_ ,
    \new_[16495]_ , \new_[16496]_ , \new_[16497]_ , \new_[16501]_ ,
    \new_[16502]_ , \new_[16506]_ , \new_[16507]_ , \new_[16508]_ ,
    \new_[16511]_ , \new_[16515]_ , \new_[16516]_ , \new_[16517]_ ,
    \new_[16521]_ , \new_[16522]_ , \new_[16526]_ , \new_[16527]_ ,
    \new_[16528]_ , \new_[16531]_ , \new_[16535]_ , \new_[16536]_ ,
    \new_[16537]_ , \new_[16541]_ , \new_[16542]_ , \new_[16546]_ ,
    \new_[16547]_ , \new_[16548]_ , \new_[16551]_ , \new_[16555]_ ,
    \new_[16556]_ , \new_[16557]_ , \new_[16561]_ , \new_[16562]_ ,
    \new_[16566]_ , \new_[16567]_ , \new_[16568]_ , \new_[16571]_ ,
    \new_[16575]_ , \new_[16576]_ , \new_[16577]_ , \new_[16581]_ ,
    \new_[16582]_ , \new_[16586]_ , \new_[16587]_ , \new_[16588]_ ,
    \new_[16591]_ , \new_[16595]_ , \new_[16596]_ , \new_[16597]_ ,
    \new_[16601]_ , \new_[16602]_ , \new_[16606]_ , \new_[16607]_ ,
    \new_[16608]_ , \new_[16611]_ , \new_[16615]_ , \new_[16616]_ ,
    \new_[16617]_ , \new_[16621]_ , \new_[16622]_ , \new_[16626]_ ,
    \new_[16627]_ , \new_[16628]_ , \new_[16631]_ , \new_[16635]_ ,
    \new_[16636]_ , \new_[16637]_ , \new_[16641]_ , \new_[16642]_ ,
    \new_[16646]_ , \new_[16647]_ , \new_[16648]_ , \new_[16651]_ ,
    \new_[16655]_ , \new_[16656]_ , \new_[16657]_ , \new_[16661]_ ,
    \new_[16662]_ , \new_[16666]_ , \new_[16667]_ , \new_[16668]_ ,
    \new_[16671]_ , \new_[16675]_ , \new_[16676]_ , \new_[16677]_ ,
    \new_[16681]_ , \new_[16682]_ , \new_[16686]_ , \new_[16687]_ ,
    \new_[16688]_ , \new_[16691]_ , \new_[16695]_ , \new_[16696]_ ,
    \new_[16697]_ , \new_[16701]_ , \new_[16702]_ , \new_[16706]_ ,
    \new_[16707]_ , \new_[16708]_ , \new_[16711]_ , \new_[16715]_ ,
    \new_[16716]_ , \new_[16717]_ , \new_[16721]_ , \new_[16722]_ ,
    \new_[16726]_ , \new_[16727]_ , \new_[16728]_ , \new_[16731]_ ,
    \new_[16735]_ , \new_[16736]_ , \new_[16737]_ , \new_[16741]_ ,
    \new_[16742]_ , \new_[16746]_ , \new_[16747]_ , \new_[16748]_ ,
    \new_[16751]_ , \new_[16755]_ , \new_[16756]_ , \new_[16757]_ ,
    \new_[16761]_ , \new_[16762]_ , \new_[16766]_ , \new_[16767]_ ,
    \new_[16768]_ , \new_[16771]_ , \new_[16775]_ , \new_[16776]_ ,
    \new_[16777]_ , \new_[16781]_ , \new_[16782]_ , \new_[16786]_ ,
    \new_[16787]_ , \new_[16788]_ , \new_[16791]_ , \new_[16795]_ ,
    \new_[16796]_ , \new_[16797]_ , \new_[16801]_ , \new_[16802]_ ,
    \new_[16806]_ , \new_[16807]_ , \new_[16808]_ , \new_[16811]_ ,
    \new_[16815]_ , \new_[16816]_ , \new_[16817]_ , \new_[16821]_ ,
    \new_[16822]_ , \new_[16826]_ , \new_[16827]_ , \new_[16828]_ ,
    \new_[16831]_ , \new_[16835]_ , \new_[16836]_ , \new_[16837]_ ,
    \new_[16841]_ , \new_[16842]_ , \new_[16846]_ , \new_[16847]_ ,
    \new_[16848]_ , \new_[16851]_ , \new_[16855]_ , \new_[16856]_ ,
    \new_[16857]_ , \new_[16861]_ , \new_[16862]_ , \new_[16866]_ ,
    \new_[16867]_ , \new_[16868]_ , \new_[16871]_ , \new_[16875]_ ,
    \new_[16876]_ , \new_[16877]_ , \new_[16881]_ , \new_[16882]_ ,
    \new_[16886]_ , \new_[16887]_ , \new_[16888]_ , \new_[16891]_ ,
    \new_[16895]_ , \new_[16896]_ , \new_[16897]_ , \new_[16901]_ ,
    \new_[16902]_ , \new_[16906]_ , \new_[16907]_ , \new_[16908]_ ,
    \new_[16911]_ , \new_[16915]_ , \new_[16916]_ , \new_[16917]_ ,
    \new_[16921]_ , \new_[16922]_ , \new_[16926]_ , \new_[16927]_ ,
    \new_[16928]_ , \new_[16931]_ , \new_[16935]_ , \new_[16936]_ ,
    \new_[16937]_ , \new_[16941]_ , \new_[16942]_ , \new_[16946]_ ,
    \new_[16947]_ , \new_[16948]_ , \new_[16951]_ , \new_[16955]_ ,
    \new_[16956]_ , \new_[16957]_ , \new_[16961]_ , \new_[16962]_ ,
    \new_[16966]_ , \new_[16967]_ , \new_[16968]_ , \new_[16971]_ ,
    \new_[16975]_ , \new_[16976]_ , \new_[16977]_ , \new_[16981]_ ,
    \new_[16982]_ , \new_[16986]_ , \new_[16987]_ , \new_[16988]_ ,
    \new_[16991]_ , \new_[16995]_ , \new_[16996]_ , \new_[16997]_ ,
    \new_[17001]_ , \new_[17002]_ , \new_[17006]_ , \new_[17007]_ ,
    \new_[17008]_ , \new_[17011]_ , \new_[17015]_ , \new_[17016]_ ,
    \new_[17017]_ , \new_[17021]_ , \new_[17022]_ , \new_[17026]_ ,
    \new_[17027]_ , \new_[17028]_ , \new_[17031]_ , \new_[17035]_ ,
    \new_[17036]_ , \new_[17037]_ , \new_[17041]_ , \new_[17042]_ ,
    \new_[17046]_ , \new_[17047]_ , \new_[17048]_ , \new_[17051]_ ,
    \new_[17055]_ , \new_[17056]_ , \new_[17057]_ , \new_[17061]_ ,
    \new_[17062]_ , \new_[17066]_ , \new_[17067]_ , \new_[17068]_ ,
    \new_[17071]_ , \new_[17075]_ , \new_[17076]_ , \new_[17077]_ ,
    \new_[17081]_ , \new_[17082]_ , \new_[17086]_ , \new_[17087]_ ,
    \new_[17088]_ , \new_[17091]_ , \new_[17095]_ , \new_[17096]_ ,
    \new_[17097]_ , \new_[17101]_ , \new_[17102]_ , \new_[17106]_ ,
    \new_[17107]_ , \new_[17108]_ , \new_[17111]_ , \new_[17115]_ ,
    \new_[17116]_ , \new_[17117]_ , \new_[17121]_ , \new_[17122]_ ,
    \new_[17126]_ , \new_[17127]_ , \new_[17128]_ , \new_[17131]_ ,
    \new_[17135]_ , \new_[17136]_ , \new_[17137]_ , \new_[17141]_ ,
    \new_[17142]_ , \new_[17146]_ , \new_[17147]_ , \new_[17148]_ ,
    \new_[17151]_ , \new_[17155]_ , \new_[17156]_ , \new_[17157]_ ,
    \new_[17161]_ , \new_[17162]_ , \new_[17166]_ , \new_[17167]_ ,
    \new_[17168]_ , \new_[17171]_ , \new_[17175]_ , \new_[17176]_ ,
    \new_[17177]_ , \new_[17181]_ , \new_[17182]_ , \new_[17186]_ ,
    \new_[17187]_ , \new_[17188]_ , \new_[17191]_ , \new_[17195]_ ,
    \new_[17196]_ , \new_[17197]_ , \new_[17201]_ , \new_[17202]_ ,
    \new_[17206]_ , \new_[17207]_ , \new_[17208]_ , \new_[17211]_ ,
    \new_[17215]_ , \new_[17216]_ , \new_[17217]_ , \new_[17221]_ ,
    \new_[17222]_ , \new_[17226]_ , \new_[17227]_ , \new_[17228]_ ,
    \new_[17231]_ , \new_[17235]_ , \new_[17236]_ , \new_[17237]_ ,
    \new_[17241]_ , \new_[17242]_ , \new_[17246]_ , \new_[17247]_ ,
    \new_[17248]_ , \new_[17251]_ , \new_[17255]_ , \new_[17256]_ ,
    \new_[17257]_ , \new_[17261]_ , \new_[17262]_ , \new_[17266]_ ,
    \new_[17267]_ , \new_[17268]_ , \new_[17271]_ , \new_[17275]_ ,
    \new_[17276]_ , \new_[17277]_ , \new_[17281]_ , \new_[17282]_ ,
    \new_[17286]_ , \new_[17287]_ , \new_[17288]_ , \new_[17291]_ ,
    \new_[17295]_ , \new_[17296]_ , \new_[17297]_ , \new_[17301]_ ,
    \new_[17302]_ , \new_[17306]_ , \new_[17307]_ , \new_[17308]_ ,
    \new_[17311]_ , \new_[17315]_ , \new_[17316]_ , \new_[17317]_ ,
    \new_[17321]_ , \new_[17322]_ , \new_[17326]_ , \new_[17327]_ ,
    \new_[17328]_ , \new_[17331]_ , \new_[17335]_ , \new_[17336]_ ,
    \new_[17337]_ , \new_[17341]_ , \new_[17342]_ , \new_[17346]_ ,
    \new_[17347]_ , \new_[17348]_ , \new_[17351]_ , \new_[17355]_ ,
    \new_[17356]_ , \new_[17357]_ , \new_[17361]_ , \new_[17362]_ ,
    \new_[17366]_ , \new_[17367]_ , \new_[17368]_ , \new_[17371]_ ,
    \new_[17375]_ , \new_[17376]_ , \new_[17377]_ , \new_[17381]_ ,
    \new_[17382]_ , \new_[17386]_ , \new_[17387]_ , \new_[17388]_ ,
    \new_[17391]_ , \new_[17395]_ , \new_[17396]_ , \new_[17397]_ ,
    \new_[17401]_ , \new_[17402]_ , \new_[17406]_ , \new_[17407]_ ,
    \new_[17408]_ , \new_[17411]_ , \new_[17415]_ , \new_[17416]_ ,
    \new_[17417]_ , \new_[17421]_ , \new_[17422]_ , \new_[17426]_ ,
    \new_[17427]_ , \new_[17428]_ , \new_[17432]_ , \new_[17433]_ ,
    \new_[17437]_ , \new_[17438]_ , \new_[17439]_ , \new_[17443]_ ,
    \new_[17444]_ , \new_[17448]_ , \new_[17449]_ , \new_[17450]_ ,
    \new_[17454]_ , \new_[17455]_ , \new_[17459]_ , \new_[17460]_ ,
    \new_[17461]_ , \new_[17465]_ , \new_[17466]_ , \new_[17470]_ ,
    \new_[17471]_ , \new_[17472]_ , \new_[17476]_ , \new_[17477]_ ,
    \new_[17481]_ , \new_[17482]_ , \new_[17483]_ , \new_[17487]_ ,
    \new_[17488]_ , \new_[17492]_ , \new_[17493]_ , \new_[17494]_ ,
    \new_[17498]_ , \new_[17499]_ , \new_[17503]_ , \new_[17504]_ ,
    \new_[17505]_ , \new_[17509]_ , \new_[17510]_ , \new_[17514]_ ,
    \new_[17515]_ , \new_[17516]_ , \new_[17520]_ , \new_[17521]_ ,
    \new_[17525]_ , \new_[17526]_ , \new_[17527]_ , \new_[17531]_ ,
    \new_[17532]_ , \new_[17536]_ , \new_[17537]_ , \new_[17538]_ ,
    \new_[17542]_ , \new_[17543]_ , \new_[17547]_ , \new_[17548]_ ,
    \new_[17549]_ , \new_[17553]_ , \new_[17554]_ , \new_[17558]_ ,
    \new_[17559]_ , \new_[17560]_ , \new_[17564]_ , \new_[17565]_ ,
    \new_[17569]_ , \new_[17570]_ , \new_[17571]_ , \new_[17575]_ ,
    \new_[17576]_ , \new_[17580]_ , \new_[17581]_ , \new_[17582]_ ,
    \new_[17586]_ , \new_[17587]_ , \new_[17591]_ , \new_[17592]_ ,
    \new_[17593]_ , \new_[17597]_ , \new_[17598]_ , \new_[17602]_ ,
    \new_[17603]_ , \new_[17604]_ , \new_[17608]_ , \new_[17609]_ ,
    \new_[17613]_ , \new_[17614]_ , \new_[17615]_ , \new_[17619]_ ,
    \new_[17620]_ , \new_[17624]_ , \new_[17625]_ , \new_[17626]_ ,
    \new_[17630]_ , \new_[17631]_ , \new_[17635]_ , \new_[17636]_ ,
    \new_[17637]_ , \new_[17641]_ , \new_[17642]_ , \new_[17646]_ ,
    \new_[17647]_ , \new_[17648]_ , \new_[17652]_ , \new_[17653]_ ,
    \new_[17657]_ , \new_[17658]_ , \new_[17659]_ , \new_[17663]_ ,
    \new_[17664]_ , \new_[17668]_ , \new_[17669]_ , \new_[17670]_ ,
    \new_[17674]_ , \new_[17675]_ , \new_[17679]_ , \new_[17680]_ ,
    \new_[17681]_ , \new_[17685]_ , \new_[17686]_ , \new_[17690]_ ,
    \new_[17691]_ , \new_[17692]_ , \new_[17696]_ , \new_[17697]_ ,
    \new_[17701]_ , \new_[17702]_ , \new_[17703]_ , \new_[17707]_ ,
    \new_[17708]_ , \new_[17712]_ , \new_[17713]_ , \new_[17714]_ ,
    \new_[17718]_ , \new_[17719]_ , \new_[17723]_ , \new_[17724]_ ,
    \new_[17725]_ , \new_[17729]_ , \new_[17730]_ , \new_[17734]_ ,
    \new_[17735]_ , \new_[17736]_ , \new_[17740]_ , \new_[17741]_ ,
    \new_[17745]_ , \new_[17746]_ , \new_[17747]_ , \new_[17751]_ ,
    \new_[17752]_ , \new_[17756]_ , \new_[17757]_ , \new_[17758]_ ,
    \new_[17762]_ , \new_[17763]_ , \new_[17767]_ , \new_[17768]_ ,
    \new_[17769]_ , \new_[17773]_ , \new_[17774]_ , \new_[17778]_ ,
    \new_[17779]_ , \new_[17780]_ , \new_[17784]_ , \new_[17785]_ ,
    \new_[17789]_ , \new_[17790]_ , \new_[17791]_ , \new_[17795]_ ,
    \new_[17796]_ , \new_[17800]_ , \new_[17801]_ , \new_[17802]_ ,
    \new_[17806]_ , \new_[17807]_ , \new_[17811]_ , \new_[17812]_ ,
    \new_[17813]_ , \new_[17817]_ , \new_[17818]_ , \new_[17822]_ ,
    \new_[17823]_ , \new_[17824]_ , \new_[17828]_ , \new_[17829]_ ,
    \new_[17833]_ , \new_[17834]_ , \new_[17835]_ , \new_[17839]_ ,
    \new_[17840]_ , \new_[17844]_ , \new_[17845]_ , \new_[17846]_ ,
    \new_[17850]_ , \new_[17851]_ , \new_[17855]_ , \new_[17856]_ ,
    \new_[17857]_ , \new_[17861]_ , \new_[17862]_ , \new_[17866]_ ,
    \new_[17867]_ , \new_[17868]_ , \new_[17872]_ , \new_[17873]_ ,
    \new_[17877]_ , \new_[17878]_ , \new_[17879]_ , \new_[17883]_ ,
    \new_[17884]_ , \new_[17888]_ , \new_[17889]_ , \new_[17890]_ ,
    \new_[17894]_ , \new_[17895]_ , \new_[17899]_ , \new_[17900]_ ,
    \new_[17901]_ , \new_[17905]_ , \new_[17906]_ , \new_[17910]_ ,
    \new_[17911]_ , \new_[17912]_ , \new_[17916]_ , \new_[17917]_ ,
    \new_[17921]_ , \new_[17922]_ , \new_[17923]_ , \new_[17927]_ ,
    \new_[17928]_ , \new_[17932]_ , \new_[17933]_ , \new_[17934]_ ,
    \new_[17938]_ , \new_[17939]_ , \new_[17943]_ , \new_[17944]_ ,
    \new_[17945]_ , \new_[17949]_ , \new_[17950]_ , \new_[17954]_ ,
    \new_[17955]_ , \new_[17956]_ , \new_[17960]_ , \new_[17961]_ ,
    \new_[17965]_ , \new_[17966]_ , \new_[17967]_ , \new_[17971]_ ,
    \new_[17972]_ , \new_[17976]_ , \new_[17977]_ , \new_[17978]_ ,
    \new_[17982]_ , \new_[17983]_ , \new_[17987]_ , \new_[17988]_ ,
    \new_[17989]_ , \new_[17993]_ , \new_[17994]_ , \new_[17998]_ ,
    \new_[17999]_ , \new_[18000]_ , \new_[18004]_ , \new_[18005]_ ,
    \new_[18009]_ , \new_[18010]_ , \new_[18011]_ , \new_[18015]_ ,
    \new_[18016]_ , \new_[18020]_ , \new_[18021]_ , \new_[18022]_ ,
    \new_[18026]_ , \new_[18027]_ , \new_[18031]_ , \new_[18032]_ ,
    \new_[18033]_ , \new_[18037]_ , \new_[18038]_ , \new_[18042]_ ,
    \new_[18043]_ , \new_[18044]_ , \new_[18048]_ , \new_[18049]_ ,
    \new_[18053]_ , \new_[18054]_ , \new_[18055]_ , \new_[18059]_ ,
    \new_[18060]_ , \new_[18064]_ , \new_[18065]_ , \new_[18066]_ ,
    \new_[18070]_ , \new_[18071]_ , \new_[18075]_ , \new_[18076]_ ,
    \new_[18077]_ , \new_[18081]_ , \new_[18082]_ , \new_[18086]_ ,
    \new_[18087]_ , \new_[18088]_ , \new_[18092]_ , \new_[18093]_ ,
    \new_[18097]_ , \new_[18098]_ , \new_[18099]_ , \new_[18103]_ ,
    \new_[18104]_ , \new_[18108]_ , \new_[18109]_ , \new_[18110]_ ,
    \new_[18114]_ , \new_[18115]_ , \new_[18119]_ , \new_[18120]_ ,
    \new_[18121]_ , \new_[18125]_ , \new_[18126]_ , \new_[18130]_ ,
    \new_[18131]_ , \new_[18132]_ , \new_[18136]_ , \new_[18137]_ ,
    \new_[18141]_ , \new_[18142]_ , \new_[18143]_ , \new_[18147]_ ,
    \new_[18148]_ , \new_[18152]_ , \new_[18153]_ , \new_[18154]_ ,
    \new_[18158]_ , \new_[18159]_ , \new_[18163]_ , \new_[18164]_ ,
    \new_[18165]_ , \new_[18169]_ , \new_[18170]_ , \new_[18174]_ ,
    \new_[18175]_ , \new_[18176]_ , \new_[18180]_ , \new_[18181]_ ,
    \new_[18185]_ , \new_[18186]_ , \new_[18187]_ , \new_[18191]_ ,
    \new_[18192]_ , \new_[18196]_ , \new_[18197]_ , \new_[18198]_ ,
    \new_[18202]_ , \new_[18203]_ , \new_[18207]_ , \new_[18208]_ ,
    \new_[18209]_ , \new_[18213]_ , \new_[18214]_ , \new_[18218]_ ,
    \new_[18219]_ , \new_[18220]_ , \new_[18224]_ , \new_[18225]_ ,
    \new_[18229]_ , \new_[18230]_ , \new_[18231]_ , \new_[18235]_ ,
    \new_[18236]_ , \new_[18240]_ , \new_[18241]_ , \new_[18242]_ ,
    \new_[18246]_ , \new_[18247]_ , \new_[18251]_ , \new_[18252]_ ,
    \new_[18253]_ , \new_[18257]_ , \new_[18258]_ , \new_[18262]_ ,
    \new_[18263]_ , \new_[18264]_ , \new_[18268]_ , \new_[18269]_ ,
    \new_[18273]_ , \new_[18274]_ , \new_[18275]_ , \new_[18279]_ ,
    \new_[18280]_ , \new_[18284]_ , \new_[18285]_ , \new_[18286]_ ,
    \new_[18290]_ , \new_[18291]_ , \new_[18295]_ , \new_[18296]_ ,
    \new_[18297]_ , \new_[18301]_ , \new_[18302]_ , \new_[18306]_ ,
    \new_[18307]_ , \new_[18308]_ , \new_[18312]_ , \new_[18313]_ ,
    \new_[18317]_ , \new_[18318]_ , \new_[18319]_ , \new_[18323]_ ,
    \new_[18324]_ , \new_[18328]_ , \new_[18329]_ , \new_[18330]_ ,
    \new_[18334]_ , \new_[18335]_ , \new_[18339]_ , \new_[18340]_ ,
    \new_[18341]_ , \new_[18345]_ , \new_[18346]_ , \new_[18350]_ ,
    \new_[18351]_ , \new_[18352]_ , \new_[18356]_ , \new_[18357]_ ,
    \new_[18361]_ , \new_[18362]_ , \new_[18363]_ , \new_[18367]_ ,
    \new_[18368]_ , \new_[18372]_ , \new_[18373]_ , \new_[18374]_ ,
    \new_[18378]_ , \new_[18379]_ , \new_[18383]_ , \new_[18384]_ ,
    \new_[18385]_ , \new_[18389]_ , \new_[18390]_ , \new_[18394]_ ,
    \new_[18395]_ , \new_[18396]_ , \new_[18400]_ , \new_[18401]_ ,
    \new_[18405]_ , \new_[18406]_ , \new_[18407]_ , \new_[18411]_ ,
    \new_[18412]_ , \new_[18416]_ , \new_[18417]_ , \new_[18418]_ ,
    \new_[18422]_ , \new_[18423]_ , \new_[18427]_ , \new_[18428]_ ,
    \new_[18429]_ , \new_[18433]_ , \new_[18434]_ , \new_[18438]_ ,
    \new_[18439]_ , \new_[18440]_ , \new_[18444]_ , \new_[18445]_ ,
    \new_[18449]_ , \new_[18450]_ , \new_[18451]_ , \new_[18455]_ ,
    \new_[18456]_ , \new_[18460]_ , \new_[18461]_ , \new_[18462]_ ,
    \new_[18466]_ , \new_[18467]_ , \new_[18471]_ , \new_[18472]_ ,
    \new_[18473]_ , \new_[18477]_ , \new_[18478]_ , \new_[18482]_ ,
    \new_[18483]_ , \new_[18484]_ , \new_[18488]_ , \new_[18489]_ ,
    \new_[18493]_ , \new_[18494]_ , \new_[18495]_ , \new_[18499]_ ,
    \new_[18500]_ , \new_[18504]_ , \new_[18505]_ , \new_[18506]_ ,
    \new_[18510]_ , \new_[18511]_ , \new_[18515]_ , \new_[18516]_ ,
    \new_[18517]_ , \new_[18521]_ , \new_[18522]_ , \new_[18526]_ ,
    \new_[18527]_ , \new_[18528]_ , \new_[18532]_ , \new_[18533]_ ,
    \new_[18537]_ , \new_[18538]_ , \new_[18539]_ , \new_[18543]_ ,
    \new_[18544]_ , \new_[18548]_ , \new_[18549]_ , \new_[18550]_ ,
    \new_[18554]_ , \new_[18555]_ , \new_[18559]_ , \new_[18560]_ ,
    \new_[18561]_ , \new_[18565]_ , \new_[18566]_ , \new_[18570]_ ,
    \new_[18571]_ , \new_[18572]_ , \new_[18576]_ , \new_[18577]_ ,
    \new_[18581]_ , \new_[18582]_ , \new_[18583]_ , \new_[18587]_ ,
    \new_[18588]_ , \new_[18592]_ , \new_[18593]_ , \new_[18594]_ ,
    \new_[18598]_ , \new_[18599]_ , \new_[18603]_ , \new_[18604]_ ,
    \new_[18605]_ , \new_[18609]_ , \new_[18610]_ , \new_[18614]_ ,
    \new_[18615]_ , \new_[18616]_ , \new_[18620]_ , \new_[18621]_ ,
    \new_[18625]_ , \new_[18626]_ , \new_[18627]_ , \new_[18631]_ ,
    \new_[18632]_ , \new_[18636]_ , \new_[18637]_ , \new_[18638]_ ,
    \new_[18642]_ , \new_[18643]_ , \new_[18647]_ , \new_[18648]_ ,
    \new_[18649]_ , \new_[18653]_ , \new_[18654]_ , \new_[18658]_ ,
    \new_[18659]_ , \new_[18660]_ , \new_[18664]_ , \new_[18665]_ ,
    \new_[18669]_ , \new_[18670]_ , \new_[18671]_ , \new_[18675]_ ,
    \new_[18676]_ , \new_[18680]_ , \new_[18681]_ , \new_[18682]_ ,
    \new_[18686]_ , \new_[18687]_ , \new_[18691]_ , \new_[18692]_ ,
    \new_[18693]_ , \new_[18697]_ , \new_[18698]_ , \new_[18702]_ ,
    \new_[18703]_ , \new_[18704]_ , \new_[18708]_ , \new_[18709]_ ,
    \new_[18713]_ , \new_[18714]_ , \new_[18715]_ , \new_[18719]_ ,
    \new_[18720]_ , \new_[18724]_ , \new_[18725]_ , \new_[18726]_ ,
    \new_[18730]_ , \new_[18731]_ , \new_[18735]_ , \new_[18736]_ ,
    \new_[18737]_ , \new_[18741]_ , \new_[18742]_ , \new_[18746]_ ,
    \new_[18747]_ , \new_[18748]_ , \new_[18752]_ , \new_[18753]_ ,
    \new_[18757]_ , \new_[18758]_ , \new_[18759]_ , \new_[18763]_ ,
    \new_[18764]_ , \new_[18768]_ , \new_[18769]_ , \new_[18770]_ ,
    \new_[18774]_ , \new_[18775]_ , \new_[18779]_ , \new_[18780]_ ,
    \new_[18781]_ , \new_[18785]_ , \new_[18786]_ , \new_[18790]_ ,
    \new_[18791]_ , \new_[18792]_ , \new_[18796]_ , \new_[18797]_ ,
    \new_[18801]_ , \new_[18802]_ , \new_[18803]_ , \new_[18807]_ ,
    \new_[18808]_ , \new_[18812]_ , \new_[18813]_ , \new_[18814]_ ,
    \new_[18818]_ , \new_[18819]_ , \new_[18823]_ , \new_[18824]_ ,
    \new_[18825]_ , \new_[18829]_ , \new_[18830]_ , \new_[18834]_ ,
    \new_[18835]_ , \new_[18836]_ , \new_[18840]_ , \new_[18841]_ ,
    \new_[18845]_ , \new_[18846]_ , \new_[18847]_ , \new_[18851]_ ,
    \new_[18852]_ , \new_[18856]_ , \new_[18857]_ , \new_[18858]_ ,
    \new_[18862]_ , \new_[18863]_ , \new_[18867]_ , \new_[18868]_ ,
    \new_[18869]_ , \new_[18873]_ , \new_[18874]_ , \new_[18878]_ ,
    \new_[18879]_ , \new_[18880]_ , \new_[18884]_ , \new_[18885]_ ,
    \new_[18889]_ , \new_[18890]_ , \new_[18891]_ , \new_[18895]_ ,
    \new_[18896]_ , \new_[18900]_ , \new_[18901]_ , \new_[18902]_ ,
    \new_[18906]_ , \new_[18907]_ , \new_[18911]_ , \new_[18912]_ ,
    \new_[18913]_ , \new_[18917]_ , \new_[18918]_ , \new_[18922]_ ,
    \new_[18923]_ , \new_[18924]_ , \new_[18928]_ , \new_[18929]_ ,
    \new_[18933]_ , \new_[18934]_ , \new_[18935]_ , \new_[18939]_ ,
    \new_[18940]_ , \new_[18944]_ , \new_[18945]_ , \new_[18946]_ ,
    \new_[18950]_ , \new_[18951]_ , \new_[18955]_ , \new_[18956]_ ,
    \new_[18957]_ , \new_[18961]_ , \new_[18962]_ , \new_[18966]_ ,
    \new_[18967]_ , \new_[18968]_ , \new_[18972]_ , \new_[18973]_ ,
    \new_[18977]_ , \new_[18978]_ , \new_[18979]_ , \new_[18983]_ ,
    \new_[18984]_ , \new_[18988]_ , \new_[18989]_ , \new_[18990]_ ,
    \new_[18994]_ , \new_[18995]_ , \new_[18999]_ , \new_[19000]_ ,
    \new_[19001]_ , \new_[19005]_ , \new_[19006]_ , \new_[19010]_ ,
    \new_[19011]_ , \new_[19012]_ , \new_[19016]_ , \new_[19017]_ ,
    \new_[19021]_ , \new_[19022]_ , \new_[19023]_ , \new_[19027]_ ,
    \new_[19028]_ , \new_[19032]_ , \new_[19033]_ , \new_[19034]_ ,
    \new_[19038]_ , \new_[19039]_ , \new_[19043]_ , \new_[19044]_ ,
    \new_[19045]_ , \new_[19049]_ , \new_[19050]_ , \new_[19054]_ ,
    \new_[19055]_ , \new_[19056]_ , \new_[19060]_ , \new_[19061]_ ,
    \new_[19065]_ , \new_[19066]_ , \new_[19067]_ , \new_[19071]_ ,
    \new_[19072]_ , \new_[19076]_ , \new_[19077]_ , \new_[19078]_ ,
    \new_[19082]_ , \new_[19083]_ , \new_[19087]_ , \new_[19088]_ ,
    \new_[19089]_ , \new_[19093]_ , \new_[19094]_ , \new_[19098]_ ,
    \new_[19099]_ , \new_[19100]_ , \new_[19104]_ , \new_[19105]_ ,
    \new_[19109]_ , \new_[19110]_ , \new_[19111]_ , \new_[19115]_ ,
    \new_[19116]_ , \new_[19120]_ , \new_[19121]_ , \new_[19122]_ ,
    \new_[19126]_ , \new_[19127]_ , \new_[19131]_ , \new_[19132]_ ,
    \new_[19133]_ , \new_[19137]_ , \new_[19138]_ , \new_[19142]_ ,
    \new_[19143]_ , \new_[19144]_ , \new_[19148]_ , \new_[19149]_ ,
    \new_[19153]_ , \new_[19154]_ , \new_[19155]_ , \new_[19159]_ ,
    \new_[19160]_ , \new_[19164]_ , \new_[19165]_ , \new_[19166]_ ,
    \new_[19170]_ , \new_[19171]_ , \new_[19175]_ , \new_[19176]_ ,
    \new_[19177]_ , \new_[19181]_ , \new_[19182]_ , \new_[19186]_ ,
    \new_[19187]_ , \new_[19188]_ , \new_[19192]_ , \new_[19193]_ ,
    \new_[19197]_ , \new_[19198]_ , \new_[19199]_ , \new_[19203]_ ,
    \new_[19204]_ , \new_[19208]_ , \new_[19209]_ , \new_[19210]_ ,
    \new_[19214]_ , \new_[19215]_ , \new_[19219]_ , \new_[19220]_ ,
    \new_[19221]_ , \new_[19225]_ , \new_[19226]_ , \new_[19230]_ ,
    \new_[19231]_ , \new_[19232]_ , \new_[19236]_ , \new_[19237]_ ,
    \new_[19241]_ , \new_[19242]_ , \new_[19243]_ , \new_[19247]_ ,
    \new_[19248]_ , \new_[19252]_ , \new_[19253]_ , \new_[19254]_ ,
    \new_[19258]_ , \new_[19259]_ , \new_[19263]_ , \new_[19264]_ ,
    \new_[19265]_ , \new_[19269]_ , \new_[19270]_ , \new_[19274]_ ,
    \new_[19275]_ , \new_[19276]_ , \new_[19280]_ , \new_[19281]_ ,
    \new_[19285]_ , \new_[19286]_ , \new_[19287]_ , \new_[19291]_ ,
    \new_[19292]_ , \new_[19296]_ , \new_[19297]_ , \new_[19298]_ ,
    \new_[19302]_ , \new_[19303]_ , \new_[19307]_ , \new_[19308]_ ,
    \new_[19309]_ , \new_[19313]_ , \new_[19314]_ , \new_[19318]_ ,
    \new_[19319]_ , \new_[19320]_ , \new_[19324]_ , \new_[19325]_ ,
    \new_[19329]_ , \new_[19330]_ , \new_[19331]_ , \new_[19335]_ ,
    \new_[19336]_ , \new_[19340]_ , \new_[19341]_ , \new_[19342]_ ,
    \new_[19346]_ , \new_[19347]_ , \new_[19351]_ , \new_[19352]_ ,
    \new_[19353]_ , \new_[19357]_ , \new_[19358]_ , \new_[19362]_ ,
    \new_[19363]_ , \new_[19364]_ , \new_[19368]_ , \new_[19369]_ ,
    \new_[19373]_ , \new_[19374]_ , \new_[19375]_ , \new_[19379]_ ,
    \new_[19380]_ , \new_[19384]_ , \new_[19385]_ , \new_[19386]_ ,
    \new_[19390]_ , \new_[19391]_ , \new_[19395]_ , \new_[19396]_ ,
    \new_[19397]_ , \new_[19401]_ , \new_[19402]_ , \new_[19406]_ ,
    \new_[19407]_ , \new_[19408]_ , \new_[19412]_ , \new_[19413]_ ,
    \new_[19417]_ , \new_[19418]_ , \new_[19419]_ , \new_[19423]_ ,
    \new_[19424]_ , \new_[19428]_ , \new_[19429]_ , \new_[19430]_ ,
    \new_[19434]_ , \new_[19435]_ , \new_[19439]_ , \new_[19440]_ ,
    \new_[19441]_ , \new_[19445]_ , \new_[19446]_ , \new_[19450]_ ,
    \new_[19451]_ , \new_[19452]_ , \new_[19456]_ , \new_[19457]_ ,
    \new_[19461]_ , \new_[19462]_ , \new_[19463]_ , \new_[19467]_ ,
    \new_[19468]_ , \new_[19472]_ , \new_[19473]_ , \new_[19474]_ ,
    \new_[19478]_ , \new_[19479]_ , \new_[19483]_ , \new_[19484]_ ,
    \new_[19485]_ , \new_[19489]_ , \new_[19490]_ , \new_[19494]_ ,
    \new_[19495]_ , \new_[19496]_ , \new_[19500]_ , \new_[19501]_ ,
    \new_[19505]_ , \new_[19506]_ , \new_[19507]_ , \new_[19511]_ ,
    \new_[19512]_ , \new_[19516]_ , \new_[19517]_ , \new_[19518]_ ,
    \new_[19522]_ , \new_[19523]_ , \new_[19527]_ , \new_[19528]_ ,
    \new_[19529]_ , \new_[19533]_ , \new_[19534]_ , \new_[19538]_ ,
    \new_[19539]_ , \new_[19540]_ , \new_[19544]_ , \new_[19545]_ ,
    \new_[19549]_ , \new_[19550]_ , \new_[19551]_ , \new_[19555]_ ,
    \new_[19556]_ , \new_[19560]_ , \new_[19561]_ , \new_[19562]_ ,
    \new_[19566]_ , \new_[19567]_ , \new_[19571]_ , \new_[19572]_ ,
    \new_[19573]_ , \new_[19577]_ , \new_[19578]_ , \new_[19582]_ ,
    \new_[19583]_ , \new_[19584]_ , \new_[19588]_ , \new_[19589]_ ,
    \new_[19593]_ , \new_[19594]_ , \new_[19595]_ , \new_[19599]_ ,
    \new_[19600]_ , \new_[19604]_ , \new_[19605]_ , \new_[19606]_ ,
    \new_[19610]_ , \new_[19611]_ , \new_[19615]_ , \new_[19616]_ ,
    \new_[19617]_ , \new_[19621]_ , \new_[19622]_ , \new_[19626]_ ,
    \new_[19627]_ , \new_[19628]_ , \new_[19632]_ , \new_[19633]_ ,
    \new_[19637]_ , \new_[19638]_ , \new_[19639]_ , \new_[19643]_ ,
    \new_[19644]_ , \new_[19648]_ , \new_[19649]_ , \new_[19650]_ ,
    \new_[19654]_ , \new_[19655]_ , \new_[19659]_ , \new_[19660]_ ,
    \new_[19661]_ , \new_[19665]_ , \new_[19666]_ , \new_[19670]_ ,
    \new_[19671]_ , \new_[19672]_ , \new_[19676]_ , \new_[19677]_ ,
    \new_[19681]_ , \new_[19682]_ , \new_[19683]_ , \new_[19687]_ ,
    \new_[19688]_ , \new_[19692]_ , \new_[19693]_ , \new_[19694]_ ,
    \new_[19698]_ , \new_[19699]_ , \new_[19703]_ , \new_[19704]_ ,
    \new_[19705]_ , \new_[19709]_ , \new_[19710]_ , \new_[19714]_ ,
    \new_[19715]_ , \new_[19716]_ , \new_[19720]_ , \new_[19721]_ ,
    \new_[19725]_ , \new_[19726]_ , \new_[19727]_ , \new_[19731]_ ,
    \new_[19732]_ , \new_[19736]_ , \new_[19737]_ , \new_[19738]_ ,
    \new_[19742]_ , \new_[19743]_ , \new_[19747]_ , \new_[19748]_ ,
    \new_[19749]_ , \new_[19753]_ , \new_[19754]_ , \new_[19758]_ ,
    \new_[19759]_ , \new_[19760]_ , \new_[19764]_ , \new_[19765]_ ,
    \new_[19769]_ , \new_[19770]_ , \new_[19771]_ , \new_[19775]_ ,
    \new_[19776]_ , \new_[19780]_ , \new_[19781]_ , \new_[19782]_ ,
    \new_[19786]_ , \new_[19787]_ , \new_[19791]_ , \new_[19792]_ ,
    \new_[19793]_ , \new_[19797]_ , \new_[19798]_ , \new_[19802]_ ,
    \new_[19803]_ , \new_[19804]_ , \new_[19808]_ , \new_[19809]_ ,
    \new_[19813]_ , \new_[19814]_ , \new_[19815]_ , \new_[19819]_ ,
    \new_[19820]_ , \new_[19824]_ , \new_[19825]_ , \new_[19826]_ ,
    \new_[19830]_ , \new_[19831]_ , \new_[19835]_ , \new_[19836]_ ,
    \new_[19837]_ , \new_[19841]_ , \new_[19842]_ , \new_[19846]_ ,
    \new_[19847]_ , \new_[19848]_ , \new_[19852]_ , \new_[19853]_ ,
    \new_[19857]_ , \new_[19858]_ , \new_[19859]_ , \new_[19863]_ ,
    \new_[19864]_ , \new_[19868]_ , \new_[19869]_ , \new_[19870]_ ,
    \new_[19874]_ , \new_[19875]_ , \new_[19879]_ , \new_[19880]_ ,
    \new_[19881]_ , \new_[19885]_ , \new_[19886]_ , \new_[19890]_ ,
    \new_[19891]_ , \new_[19892]_ , \new_[19896]_ , \new_[19897]_ ,
    \new_[19901]_ , \new_[19902]_ , \new_[19903]_ , \new_[19907]_ ,
    \new_[19908]_ , \new_[19912]_ , \new_[19913]_ , \new_[19914]_ ,
    \new_[19918]_ , \new_[19919]_ , \new_[19923]_ , \new_[19924]_ ,
    \new_[19925]_ , \new_[19929]_ , \new_[19930]_ , \new_[19934]_ ,
    \new_[19935]_ , \new_[19936]_ , \new_[19940]_ , \new_[19941]_ ,
    \new_[19945]_ , \new_[19946]_ , \new_[19947]_ , \new_[19951]_ ,
    \new_[19952]_ , \new_[19956]_ , \new_[19957]_ , \new_[19958]_ ,
    \new_[19962]_ , \new_[19963]_ , \new_[19967]_ , \new_[19968]_ ,
    \new_[19969]_ , \new_[19973]_ , \new_[19974]_ , \new_[19978]_ ,
    \new_[19979]_ , \new_[19980]_ , \new_[19984]_ , \new_[19985]_ ,
    \new_[19989]_ , \new_[19990]_ , \new_[19991]_ , \new_[19995]_ ,
    \new_[19996]_ , \new_[20000]_ , \new_[20001]_ , \new_[20002]_ ,
    \new_[20006]_ , \new_[20007]_ , \new_[20011]_ , \new_[20012]_ ,
    \new_[20013]_ , \new_[20017]_ , \new_[20018]_ , \new_[20022]_ ,
    \new_[20023]_ , \new_[20024]_ , \new_[20028]_ , \new_[20029]_ ,
    \new_[20033]_ , \new_[20034]_ , \new_[20035]_ , \new_[20039]_ ,
    \new_[20040]_ , \new_[20044]_ , \new_[20045]_ , \new_[20046]_ ,
    \new_[20050]_ , \new_[20051]_ , \new_[20055]_ , \new_[20056]_ ,
    \new_[20057]_ , \new_[20061]_ , \new_[20062]_ , \new_[20066]_ ,
    \new_[20067]_ , \new_[20068]_ , \new_[20072]_ , \new_[20073]_ ,
    \new_[20077]_ , \new_[20078]_ , \new_[20079]_ , \new_[20083]_ ,
    \new_[20084]_ , \new_[20088]_ , \new_[20089]_ , \new_[20090]_ ,
    \new_[20094]_ , \new_[20095]_ , \new_[20099]_ , \new_[20100]_ ,
    \new_[20101]_ , \new_[20105]_ , \new_[20106]_ , \new_[20110]_ ,
    \new_[20111]_ , \new_[20112]_ , \new_[20116]_ , \new_[20117]_ ,
    \new_[20121]_ , \new_[20122]_ , \new_[20123]_ , \new_[20127]_ ,
    \new_[20128]_ , \new_[20132]_ , \new_[20133]_ , \new_[20134]_ ,
    \new_[20138]_ , \new_[20139]_ , \new_[20143]_ , \new_[20144]_ ,
    \new_[20145]_ , \new_[20149]_ , \new_[20150]_ , \new_[20154]_ ,
    \new_[20155]_ , \new_[20156]_ , \new_[20160]_ , \new_[20161]_ ,
    \new_[20165]_ , \new_[20166]_ , \new_[20167]_ , \new_[20171]_ ,
    \new_[20172]_ , \new_[20176]_ , \new_[20177]_ , \new_[20178]_ ,
    \new_[20182]_ , \new_[20183]_ , \new_[20187]_ , \new_[20188]_ ,
    \new_[20189]_ , \new_[20193]_ , \new_[20194]_ , \new_[20198]_ ,
    \new_[20199]_ , \new_[20200]_ , \new_[20204]_ , \new_[20205]_ ,
    \new_[20209]_ , \new_[20210]_ , \new_[20211]_ , \new_[20215]_ ,
    \new_[20216]_ , \new_[20220]_ , \new_[20221]_ , \new_[20222]_ ,
    \new_[20226]_ , \new_[20227]_ , \new_[20231]_ , \new_[20232]_ ,
    \new_[20233]_ , \new_[20237]_ , \new_[20238]_ , \new_[20242]_ ,
    \new_[20243]_ , \new_[20244]_ , \new_[20248]_ , \new_[20249]_ ,
    \new_[20253]_ , \new_[20254]_ , \new_[20255]_ , \new_[20259]_ ,
    \new_[20260]_ , \new_[20264]_ , \new_[20265]_ , \new_[20266]_ ,
    \new_[20270]_ , \new_[20271]_ , \new_[20275]_ , \new_[20276]_ ,
    \new_[20277]_ , \new_[20281]_ , \new_[20282]_ , \new_[20286]_ ,
    \new_[20287]_ , \new_[20288]_ , \new_[20292]_ , \new_[20293]_ ,
    \new_[20297]_ , \new_[20298]_ , \new_[20299]_ , \new_[20303]_ ,
    \new_[20304]_ , \new_[20308]_ , \new_[20309]_ , \new_[20310]_ ,
    \new_[20314]_ , \new_[20315]_ , \new_[20319]_ , \new_[20320]_ ,
    \new_[20321]_ , \new_[20325]_ , \new_[20326]_ , \new_[20330]_ ,
    \new_[20331]_ , \new_[20332]_ , \new_[20336]_ , \new_[20337]_ ,
    \new_[20341]_ , \new_[20342]_ , \new_[20343]_ , \new_[20347]_ ,
    \new_[20348]_ , \new_[20352]_ , \new_[20353]_ , \new_[20354]_ ,
    \new_[20358]_ , \new_[20359]_ , \new_[20363]_ , \new_[20364]_ ,
    \new_[20365]_ , \new_[20369]_ , \new_[20370]_ , \new_[20374]_ ,
    \new_[20375]_ , \new_[20376]_ , \new_[20380]_ , \new_[20381]_ ,
    \new_[20385]_ , \new_[20386]_ , \new_[20387]_ , \new_[20391]_ ,
    \new_[20392]_ , \new_[20396]_ , \new_[20397]_ , \new_[20398]_ ,
    \new_[20402]_ , \new_[20403]_ , \new_[20407]_ , \new_[20408]_ ,
    \new_[20409]_ , \new_[20413]_ , \new_[20414]_ , \new_[20418]_ ,
    \new_[20419]_ , \new_[20420]_ , \new_[20424]_ , \new_[20425]_ ,
    \new_[20429]_ , \new_[20430]_ , \new_[20431]_ , \new_[20435]_ ,
    \new_[20436]_ , \new_[20440]_ , \new_[20441]_ , \new_[20442]_ ,
    \new_[20446]_ , \new_[20447]_ , \new_[20451]_ , \new_[20452]_ ,
    \new_[20453]_ , \new_[20457]_ , \new_[20458]_ , \new_[20462]_ ,
    \new_[20463]_ , \new_[20464]_ , \new_[20468]_ , \new_[20469]_ ,
    \new_[20473]_ , \new_[20474]_ , \new_[20475]_ , \new_[20479]_ ,
    \new_[20480]_ , \new_[20484]_ , \new_[20485]_ , \new_[20486]_ ,
    \new_[20490]_ , \new_[20491]_ , \new_[20495]_ , \new_[20496]_ ,
    \new_[20497]_ , \new_[20501]_ , \new_[20502]_ , \new_[20506]_ ,
    \new_[20507]_ , \new_[20508]_ , \new_[20512]_ , \new_[20513]_ ,
    \new_[20517]_ , \new_[20518]_ , \new_[20519]_ , \new_[20523]_ ,
    \new_[20524]_ , \new_[20528]_ , \new_[20529]_ , \new_[20530]_ ,
    \new_[20534]_ , \new_[20535]_ , \new_[20539]_ , \new_[20540]_ ,
    \new_[20541]_ , \new_[20545]_ , \new_[20546]_ , \new_[20550]_ ,
    \new_[20551]_ , \new_[20552]_ , \new_[20556]_ , \new_[20557]_ ,
    \new_[20561]_ , \new_[20562]_ , \new_[20563]_ , \new_[20567]_ ,
    \new_[20568]_ , \new_[20572]_ , \new_[20573]_ , \new_[20574]_ ,
    \new_[20578]_ , \new_[20579]_ , \new_[20583]_ , \new_[20584]_ ,
    \new_[20585]_ , \new_[20589]_ , \new_[20590]_ , \new_[20594]_ ,
    \new_[20595]_ , \new_[20596]_ , \new_[20600]_ , \new_[20601]_ ,
    \new_[20605]_ , \new_[20606]_ , \new_[20607]_ , \new_[20611]_ ,
    \new_[20612]_ , \new_[20616]_ , \new_[20617]_ , \new_[20618]_ ,
    \new_[20622]_ , \new_[20623]_ , \new_[20627]_ , \new_[20628]_ ,
    \new_[20629]_ , \new_[20633]_ , \new_[20634]_ , \new_[20638]_ ,
    \new_[20639]_ , \new_[20640]_ , \new_[20644]_ , \new_[20645]_ ,
    \new_[20649]_ , \new_[20650]_ , \new_[20651]_ , \new_[20655]_ ,
    \new_[20656]_ , \new_[20660]_ , \new_[20661]_ , \new_[20662]_ ,
    \new_[20666]_ , \new_[20667]_ , \new_[20671]_ , \new_[20672]_ ,
    \new_[20673]_ , \new_[20677]_ , \new_[20678]_ , \new_[20682]_ ,
    \new_[20683]_ , \new_[20684]_ , \new_[20688]_ , \new_[20689]_ ,
    \new_[20693]_ , \new_[20694]_ , \new_[20695]_ , \new_[20699]_ ,
    \new_[20700]_ , \new_[20704]_ , \new_[20705]_ , \new_[20706]_ ,
    \new_[20710]_ , \new_[20711]_ , \new_[20715]_ , \new_[20716]_ ,
    \new_[20717]_ , \new_[20721]_ , \new_[20722]_ , \new_[20726]_ ,
    \new_[20727]_ , \new_[20728]_ , \new_[20732]_ , \new_[20733]_ ,
    \new_[20737]_ , \new_[20738]_ , \new_[20739]_ , \new_[20743]_ ,
    \new_[20744]_ , \new_[20748]_ , \new_[20749]_ , \new_[20750]_ ,
    \new_[20754]_ , \new_[20755]_ , \new_[20759]_ , \new_[20760]_ ,
    \new_[20761]_ , \new_[20765]_ , \new_[20766]_ , \new_[20770]_ ,
    \new_[20771]_ , \new_[20772]_ , \new_[20776]_ , \new_[20777]_ ,
    \new_[20781]_ , \new_[20782]_ , \new_[20783]_ , \new_[20787]_ ,
    \new_[20788]_ , \new_[20792]_ , \new_[20793]_ , \new_[20794]_ ,
    \new_[20798]_ , \new_[20799]_ , \new_[20803]_ , \new_[20804]_ ,
    \new_[20805]_ , \new_[20809]_ , \new_[20810]_ , \new_[20814]_ ,
    \new_[20815]_ , \new_[20816]_ , \new_[20820]_ , \new_[20821]_ ,
    \new_[20825]_ , \new_[20826]_ , \new_[20827]_ , \new_[20831]_ ,
    \new_[20832]_ , \new_[20836]_ , \new_[20837]_ , \new_[20838]_ ,
    \new_[20842]_ , \new_[20843]_ , \new_[20847]_ , \new_[20848]_ ,
    \new_[20849]_ , \new_[20853]_ , \new_[20854]_ , \new_[20858]_ ,
    \new_[20859]_ , \new_[20860]_ , \new_[20864]_ , \new_[20865]_ ,
    \new_[20869]_ , \new_[20870]_ , \new_[20871]_ , \new_[20875]_ ,
    \new_[20876]_ , \new_[20880]_ , \new_[20881]_ , \new_[20882]_ ,
    \new_[20886]_ , \new_[20887]_ , \new_[20891]_ , \new_[20892]_ ,
    \new_[20893]_ , \new_[20897]_ , \new_[20898]_ , \new_[20902]_ ,
    \new_[20903]_ , \new_[20904]_ , \new_[20908]_ , \new_[20909]_ ,
    \new_[20913]_ , \new_[20914]_ , \new_[20915]_ , \new_[20919]_ ,
    \new_[20920]_ , \new_[20924]_ , \new_[20925]_ , \new_[20926]_ ,
    \new_[20930]_ , \new_[20931]_ , \new_[20935]_ , \new_[20936]_ ,
    \new_[20937]_ , \new_[20941]_ , \new_[20942]_ , \new_[20946]_ ,
    \new_[20947]_ , \new_[20948]_ , \new_[20952]_ , \new_[20953]_ ,
    \new_[20957]_ , \new_[20958]_ , \new_[20959]_ , \new_[20963]_ ,
    \new_[20964]_ , \new_[20968]_ , \new_[20969]_ , \new_[20970]_ ,
    \new_[20974]_ , \new_[20975]_ , \new_[20979]_ , \new_[20980]_ ,
    \new_[20981]_ , \new_[20985]_ , \new_[20986]_ , \new_[20990]_ ,
    \new_[20991]_ , \new_[20992]_ , \new_[20996]_ , \new_[20997]_ ,
    \new_[21001]_ , \new_[21002]_ , \new_[21003]_ , \new_[21007]_ ,
    \new_[21008]_ , \new_[21012]_ , \new_[21013]_ , \new_[21014]_ ,
    \new_[21018]_ , \new_[21019]_ , \new_[21023]_ , \new_[21024]_ ,
    \new_[21025]_ , \new_[21029]_ , \new_[21030]_ , \new_[21034]_ ,
    \new_[21035]_ , \new_[21036]_ , \new_[21040]_ , \new_[21041]_ ,
    \new_[21045]_ , \new_[21046]_ , \new_[21047]_ , \new_[21051]_ ,
    \new_[21052]_ , \new_[21056]_ , \new_[21057]_ , \new_[21058]_ ,
    \new_[21062]_ , \new_[21063]_ , \new_[21067]_ , \new_[21068]_ ,
    \new_[21069]_ , \new_[21073]_ , \new_[21074]_ , \new_[21078]_ ,
    \new_[21079]_ , \new_[21080]_ , \new_[21084]_ , \new_[21085]_ ,
    \new_[21089]_ , \new_[21090]_ , \new_[21091]_ , \new_[21095]_ ,
    \new_[21096]_ , \new_[21100]_ , \new_[21101]_ , \new_[21102]_ ,
    \new_[21106]_ , \new_[21107]_ , \new_[21111]_ , \new_[21112]_ ,
    \new_[21113]_ , \new_[21117]_ , \new_[21118]_ , \new_[21122]_ ,
    \new_[21123]_ , \new_[21124]_ , \new_[21128]_ , \new_[21129]_ ,
    \new_[21133]_ , \new_[21134]_ , \new_[21135]_ , \new_[21139]_ ,
    \new_[21140]_ , \new_[21144]_ , \new_[21145]_ , \new_[21146]_ ,
    \new_[21150]_ , \new_[21151]_ , \new_[21155]_ , \new_[21156]_ ,
    \new_[21157]_ , \new_[21161]_ , \new_[21162]_ , \new_[21166]_ ,
    \new_[21167]_ , \new_[21168]_ , \new_[21172]_ , \new_[21173]_ ,
    \new_[21177]_ , \new_[21178]_ , \new_[21179]_ , \new_[21183]_ ,
    \new_[21184]_ , \new_[21188]_ , \new_[21189]_ , \new_[21190]_ ,
    \new_[21194]_ , \new_[21195]_ , \new_[21199]_ , \new_[21200]_ ,
    \new_[21201]_ , \new_[21205]_ , \new_[21206]_ , \new_[21210]_ ,
    \new_[21211]_ , \new_[21212]_ , \new_[21216]_ , \new_[21217]_ ,
    \new_[21221]_ , \new_[21222]_ , \new_[21223]_ , \new_[21227]_ ,
    \new_[21228]_ , \new_[21232]_ , \new_[21233]_ , \new_[21234]_ ,
    \new_[21238]_ , \new_[21239]_ , \new_[21243]_ , \new_[21244]_ ,
    \new_[21245]_ , \new_[21249]_ , \new_[21250]_ , \new_[21254]_ ,
    \new_[21255]_ , \new_[21256]_ , \new_[21260]_ , \new_[21261]_ ,
    \new_[21265]_ , \new_[21266]_ , \new_[21267]_ , \new_[21271]_ ,
    \new_[21272]_ , \new_[21276]_ , \new_[21277]_ , \new_[21278]_ ,
    \new_[21282]_ , \new_[21283]_ , \new_[21287]_ , \new_[21288]_ ,
    \new_[21289]_ , \new_[21293]_ , \new_[21294]_ , \new_[21298]_ ,
    \new_[21299]_ , \new_[21300]_ , \new_[21304]_ , \new_[21305]_ ,
    \new_[21309]_ , \new_[21310]_ , \new_[21311]_ , \new_[21315]_ ,
    \new_[21316]_ , \new_[21320]_ , \new_[21321]_ , \new_[21322]_ ,
    \new_[21326]_ , \new_[21327]_ , \new_[21331]_ , \new_[21332]_ ,
    \new_[21333]_ , \new_[21337]_ , \new_[21338]_ , \new_[21342]_ ,
    \new_[21343]_ , \new_[21344]_ , \new_[21348]_ , \new_[21349]_ ,
    \new_[21353]_ , \new_[21354]_ , \new_[21355]_ , \new_[21359]_ ,
    \new_[21360]_ , \new_[21364]_ , \new_[21365]_ , \new_[21366]_ ,
    \new_[21370]_ , \new_[21371]_ , \new_[21375]_ , \new_[21376]_ ,
    \new_[21377]_ , \new_[21381]_ , \new_[21382]_ , \new_[21386]_ ,
    \new_[21387]_ , \new_[21388]_ , \new_[21392]_ , \new_[21393]_ ,
    \new_[21397]_ , \new_[21398]_ , \new_[21399]_ , \new_[21403]_ ,
    \new_[21404]_ , \new_[21408]_ , \new_[21409]_ , \new_[21410]_ ,
    \new_[21414]_ , \new_[21415]_ , \new_[21419]_ , \new_[21420]_ ,
    \new_[21421]_ , \new_[21425]_ , \new_[21426]_ , \new_[21430]_ ,
    \new_[21431]_ , \new_[21432]_ , \new_[21436]_ , \new_[21437]_ ,
    \new_[21441]_ , \new_[21442]_ , \new_[21443]_ , \new_[21447]_ ,
    \new_[21448]_ , \new_[21452]_ , \new_[21453]_ , \new_[21454]_ ,
    \new_[21458]_ , \new_[21459]_ , \new_[21463]_ , \new_[21464]_ ,
    \new_[21465]_ , \new_[21469]_ , \new_[21470]_ , \new_[21474]_ ,
    \new_[21475]_ , \new_[21476]_ , \new_[21480]_ , \new_[21481]_ ,
    \new_[21485]_ , \new_[21486]_ , \new_[21487]_ , \new_[21491]_ ,
    \new_[21492]_ , \new_[21496]_ , \new_[21497]_ , \new_[21498]_ ,
    \new_[21502]_ , \new_[21503]_ , \new_[21507]_ , \new_[21508]_ ,
    \new_[21509]_ , \new_[21513]_ , \new_[21514]_ , \new_[21518]_ ,
    \new_[21519]_ , \new_[21520]_ , \new_[21524]_ , \new_[21525]_ ,
    \new_[21529]_ , \new_[21530]_ , \new_[21531]_ , \new_[21535]_ ,
    \new_[21536]_ , \new_[21540]_ , \new_[21541]_ , \new_[21542]_ ,
    \new_[21546]_ , \new_[21547]_ , \new_[21551]_ , \new_[21552]_ ,
    \new_[21553]_ , \new_[21557]_ , \new_[21558]_ , \new_[21562]_ ,
    \new_[21563]_ , \new_[21564]_ , \new_[21568]_ , \new_[21569]_ ,
    \new_[21573]_ , \new_[21574]_ , \new_[21575]_ , \new_[21579]_ ,
    \new_[21580]_ , \new_[21584]_ , \new_[21585]_ , \new_[21586]_ ,
    \new_[21590]_ , \new_[21591]_ , \new_[21595]_ , \new_[21596]_ ,
    \new_[21597]_ , \new_[21601]_ , \new_[21602]_ , \new_[21606]_ ,
    \new_[21607]_ , \new_[21608]_ , \new_[21612]_ , \new_[21613]_ ,
    \new_[21617]_ , \new_[21618]_ , \new_[21619]_ , \new_[21623]_ ,
    \new_[21624]_ , \new_[21628]_ , \new_[21629]_ , \new_[21630]_ ,
    \new_[21634]_ , \new_[21635]_ , \new_[21639]_ , \new_[21640]_ ,
    \new_[21641]_ , \new_[21645]_ , \new_[21646]_ , \new_[21650]_ ,
    \new_[21651]_ , \new_[21652]_ , \new_[21656]_ , \new_[21657]_ ,
    \new_[21661]_ , \new_[21662]_ , \new_[21663]_ , \new_[21667]_ ,
    \new_[21668]_ , \new_[21672]_ , \new_[21673]_ , \new_[21674]_ ,
    \new_[21678]_ , \new_[21679]_ , \new_[21683]_ , \new_[21684]_ ,
    \new_[21685]_ , \new_[21689]_ , \new_[21690]_ , \new_[21694]_ ,
    \new_[21695]_ , \new_[21696]_ , \new_[21700]_ , \new_[21701]_ ,
    \new_[21705]_ , \new_[21706]_ , \new_[21707]_ , \new_[21711]_ ,
    \new_[21712]_ , \new_[21716]_ , \new_[21717]_ , \new_[21718]_ ,
    \new_[21722]_ , \new_[21723]_ , \new_[21727]_ , \new_[21728]_ ,
    \new_[21729]_ , \new_[21733]_ , \new_[21734]_ , \new_[21738]_ ,
    \new_[21739]_ , \new_[21740]_ , \new_[21744]_ , \new_[21745]_ ,
    \new_[21749]_ , \new_[21750]_ , \new_[21751]_ , \new_[21755]_ ,
    \new_[21756]_ , \new_[21760]_ , \new_[21761]_ , \new_[21762]_ ,
    \new_[21766]_ , \new_[21767]_ , \new_[21771]_ , \new_[21772]_ ,
    \new_[21773]_ , \new_[21777]_ , \new_[21778]_ , \new_[21782]_ ,
    \new_[21783]_ , \new_[21784]_ , \new_[21788]_ , \new_[21789]_ ,
    \new_[21793]_ , \new_[21794]_ , \new_[21795]_ , \new_[21799]_ ,
    \new_[21800]_ , \new_[21804]_ , \new_[21805]_ , \new_[21806]_ ,
    \new_[21810]_ , \new_[21811]_ , \new_[21815]_ , \new_[21816]_ ,
    \new_[21817]_ , \new_[21821]_ , \new_[21822]_ , \new_[21826]_ ,
    \new_[21827]_ , \new_[21828]_ , \new_[21832]_ , \new_[21833]_ ,
    \new_[21837]_ , \new_[21838]_ , \new_[21839]_ , \new_[21843]_ ,
    \new_[21844]_ , \new_[21848]_ , \new_[21849]_ , \new_[21850]_ ,
    \new_[21854]_ , \new_[21855]_ , \new_[21859]_ , \new_[21860]_ ,
    \new_[21861]_ , \new_[21865]_ , \new_[21866]_ , \new_[21870]_ ,
    \new_[21871]_ , \new_[21872]_ , \new_[21876]_ , \new_[21877]_ ,
    \new_[21881]_ , \new_[21882]_ , \new_[21883]_ , \new_[21887]_ ,
    \new_[21888]_ , \new_[21892]_ , \new_[21893]_ , \new_[21894]_ ,
    \new_[21898]_ , \new_[21899]_ , \new_[21903]_ , \new_[21904]_ ,
    \new_[21905]_ , \new_[21909]_ , \new_[21910]_ , \new_[21914]_ ,
    \new_[21915]_ , \new_[21916]_ , \new_[21920]_ , \new_[21921]_ ,
    \new_[21925]_ , \new_[21926]_ , \new_[21927]_ , \new_[21931]_ ,
    \new_[21932]_ , \new_[21936]_ , \new_[21937]_ , \new_[21938]_ ,
    \new_[21942]_ , \new_[21943]_ , \new_[21947]_ , \new_[21948]_ ,
    \new_[21949]_ , \new_[21953]_ , \new_[21954]_ , \new_[21958]_ ,
    \new_[21959]_ , \new_[21960]_ , \new_[21964]_ , \new_[21965]_ ,
    \new_[21969]_ , \new_[21970]_ , \new_[21971]_ , \new_[21975]_ ,
    \new_[21976]_ , \new_[21980]_ , \new_[21981]_ , \new_[21982]_ ,
    \new_[21986]_ , \new_[21987]_ , \new_[21991]_ , \new_[21992]_ ,
    \new_[21993]_ , \new_[21997]_ , \new_[21998]_ , \new_[22002]_ ,
    \new_[22003]_ , \new_[22004]_ , \new_[22008]_ , \new_[22009]_ ,
    \new_[22013]_ , \new_[22014]_ , \new_[22015]_ , \new_[22019]_ ,
    \new_[22020]_ , \new_[22024]_ , \new_[22025]_ , \new_[22026]_ ,
    \new_[22030]_ , \new_[22031]_ , \new_[22035]_ , \new_[22036]_ ,
    \new_[22037]_ , \new_[22041]_ , \new_[22042]_ , \new_[22046]_ ,
    \new_[22047]_ , \new_[22048]_ , \new_[22052]_ , \new_[22053]_ ,
    \new_[22057]_ , \new_[22058]_ , \new_[22059]_ , \new_[22063]_ ,
    \new_[22064]_ , \new_[22068]_ , \new_[22069]_ , \new_[22070]_ ,
    \new_[22074]_ , \new_[22075]_ , \new_[22079]_ , \new_[22080]_ ,
    \new_[22081]_ , \new_[22085]_ , \new_[22086]_ , \new_[22090]_ ,
    \new_[22091]_ , \new_[22092]_ , \new_[22096]_ , \new_[22097]_ ,
    \new_[22101]_ , \new_[22102]_ , \new_[22103]_ , \new_[22107]_ ,
    \new_[22108]_ , \new_[22112]_ , \new_[22113]_ , \new_[22114]_ ,
    \new_[22118]_ , \new_[22119]_ , \new_[22123]_ , \new_[22124]_ ,
    \new_[22125]_ , \new_[22129]_ , \new_[22130]_ , \new_[22134]_ ,
    \new_[22135]_ , \new_[22136]_ , \new_[22140]_ , \new_[22141]_ ,
    \new_[22145]_ , \new_[22146]_ , \new_[22147]_ , \new_[22151]_ ,
    \new_[22152]_ , \new_[22156]_ , \new_[22157]_ , \new_[22158]_ ,
    \new_[22162]_ , \new_[22163]_ , \new_[22167]_ , \new_[22168]_ ,
    \new_[22169]_ , \new_[22173]_ , \new_[22174]_ , \new_[22178]_ ,
    \new_[22179]_ , \new_[22180]_ , \new_[22184]_ , \new_[22185]_ ,
    \new_[22189]_ , \new_[22190]_ , \new_[22191]_ , \new_[22195]_ ,
    \new_[22196]_ , \new_[22200]_ , \new_[22201]_ , \new_[22202]_ ,
    \new_[22206]_ , \new_[22207]_ , \new_[22211]_ , \new_[22212]_ ,
    \new_[22213]_ , \new_[22217]_ , \new_[22218]_ , \new_[22222]_ ,
    \new_[22223]_ , \new_[22224]_ , \new_[22228]_ , \new_[22229]_ ,
    \new_[22233]_ , \new_[22234]_ , \new_[22235]_ , \new_[22239]_ ,
    \new_[22240]_ , \new_[22244]_ , \new_[22245]_ , \new_[22246]_ ,
    \new_[22250]_ , \new_[22251]_ , \new_[22255]_ , \new_[22256]_ ,
    \new_[22257]_ , \new_[22261]_ , \new_[22262]_ , \new_[22266]_ ,
    \new_[22267]_ , \new_[22268]_ , \new_[22272]_ , \new_[22273]_ ,
    \new_[22277]_ , \new_[22278]_ , \new_[22279]_ , \new_[22283]_ ,
    \new_[22284]_ , \new_[22288]_ , \new_[22289]_ , \new_[22290]_ ,
    \new_[22294]_ , \new_[22295]_ , \new_[22299]_ , \new_[22300]_ ,
    \new_[22301]_ , \new_[22305]_ , \new_[22306]_ , \new_[22310]_ ,
    \new_[22311]_ , \new_[22312]_ , \new_[22316]_ , \new_[22317]_ ,
    \new_[22321]_ , \new_[22322]_ , \new_[22323]_ , \new_[22327]_ ,
    \new_[22328]_ , \new_[22332]_ , \new_[22333]_ , \new_[22334]_ ,
    \new_[22338]_ , \new_[22339]_ , \new_[22343]_ , \new_[22344]_ ,
    \new_[22345]_ , \new_[22349]_ , \new_[22350]_ , \new_[22354]_ ,
    \new_[22355]_ , \new_[22356]_ , \new_[22360]_ , \new_[22361]_ ,
    \new_[22365]_ , \new_[22366]_ , \new_[22367]_ , \new_[22371]_ ,
    \new_[22372]_ , \new_[22376]_ , \new_[22377]_ , \new_[22378]_ ,
    \new_[22382]_ , \new_[22383]_ , \new_[22387]_ , \new_[22388]_ ,
    \new_[22389]_ , \new_[22393]_ , \new_[22394]_ , \new_[22398]_ ,
    \new_[22399]_ , \new_[22400]_ , \new_[22404]_ , \new_[22405]_ ,
    \new_[22409]_ , \new_[22410]_ , \new_[22411]_ , \new_[22415]_ ,
    \new_[22416]_ , \new_[22420]_ , \new_[22421]_ , \new_[22422]_ ,
    \new_[22426]_ , \new_[22427]_ , \new_[22431]_ , \new_[22432]_ ,
    \new_[22433]_ , \new_[22437]_ , \new_[22438]_ , \new_[22442]_ ,
    \new_[22443]_ , \new_[22444]_ , \new_[22448]_ , \new_[22449]_ ,
    \new_[22453]_ , \new_[22454]_ , \new_[22455]_ , \new_[22459]_ ,
    \new_[22460]_ , \new_[22464]_ , \new_[22465]_ , \new_[22466]_ ,
    \new_[22470]_ , \new_[22471]_ , \new_[22475]_ , \new_[22476]_ ,
    \new_[22477]_ , \new_[22481]_ , \new_[22482]_ , \new_[22486]_ ,
    \new_[22487]_ , \new_[22488]_ , \new_[22492]_ , \new_[22493]_ ,
    \new_[22497]_ , \new_[22498]_ , \new_[22499]_ , \new_[22503]_ ,
    \new_[22504]_ , \new_[22508]_ , \new_[22509]_ , \new_[22510]_ ,
    \new_[22514]_ , \new_[22515]_ , \new_[22519]_ , \new_[22520]_ ,
    \new_[22521]_ , \new_[22525]_ , \new_[22526]_ , \new_[22530]_ ,
    \new_[22531]_ , \new_[22532]_ , \new_[22536]_ , \new_[22537]_ ,
    \new_[22541]_ , \new_[22542]_ , \new_[22543]_ , \new_[22547]_ ,
    \new_[22548]_ , \new_[22552]_ , \new_[22553]_ , \new_[22554]_ ,
    \new_[22558]_ , \new_[22559]_ , \new_[22563]_ , \new_[22564]_ ,
    \new_[22565]_ , \new_[22569]_ , \new_[22570]_ , \new_[22574]_ ,
    \new_[22575]_ , \new_[22576]_ , \new_[22580]_ , \new_[22581]_ ,
    \new_[22585]_ , \new_[22586]_ , \new_[22587]_ , \new_[22591]_ ,
    \new_[22592]_ , \new_[22596]_ , \new_[22597]_ , \new_[22598]_ ,
    \new_[22602]_ , \new_[22603]_ , \new_[22607]_ , \new_[22608]_ ,
    \new_[22609]_ , \new_[22613]_ , \new_[22614]_ , \new_[22618]_ ,
    \new_[22619]_ , \new_[22620]_ , \new_[22624]_ , \new_[22625]_ ,
    \new_[22629]_ , \new_[22630]_ , \new_[22631]_ , \new_[22635]_ ,
    \new_[22636]_ , \new_[22640]_ , \new_[22641]_ , \new_[22642]_ ,
    \new_[22646]_ , \new_[22647]_ , \new_[22651]_ , \new_[22652]_ ,
    \new_[22653]_ , \new_[22657]_ , \new_[22658]_ , \new_[22662]_ ,
    \new_[22663]_ , \new_[22664]_ , \new_[22668]_ , \new_[22669]_ ,
    \new_[22673]_ , \new_[22674]_ , \new_[22675]_ , \new_[22679]_ ,
    \new_[22680]_ , \new_[22684]_ , \new_[22685]_ , \new_[22686]_ ,
    \new_[22690]_ , \new_[22691]_ , \new_[22695]_ , \new_[22696]_ ,
    \new_[22697]_ , \new_[22701]_ , \new_[22702]_ , \new_[22706]_ ,
    \new_[22707]_ , \new_[22708]_ , \new_[22712]_ , \new_[22713]_ ,
    \new_[22717]_ , \new_[22718]_ , \new_[22719]_ , \new_[22723]_ ,
    \new_[22724]_ , \new_[22728]_ , \new_[22729]_ , \new_[22730]_ ,
    \new_[22734]_ , \new_[22735]_ , \new_[22739]_ , \new_[22740]_ ,
    \new_[22741]_ , \new_[22745]_ , \new_[22746]_ , \new_[22750]_ ,
    \new_[22751]_ , \new_[22752]_ , \new_[22756]_ , \new_[22757]_ ,
    \new_[22761]_ , \new_[22762]_ , \new_[22763]_ , \new_[22767]_ ,
    \new_[22768]_ , \new_[22772]_ , \new_[22773]_ , \new_[22774]_ ,
    \new_[22778]_ , \new_[22779]_ , \new_[22783]_ , \new_[22784]_ ,
    \new_[22785]_ , \new_[22789]_ , \new_[22790]_ , \new_[22794]_ ,
    \new_[22795]_ , \new_[22796]_ , \new_[22800]_ , \new_[22801]_ ,
    \new_[22805]_ , \new_[22806]_ , \new_[22807]_ , \new_[22811]_ ,
    \new_[22812]_ , \new_[22816]_ , \new_[22817]_ , \new_[22818]_ ,
    \new_[22822]_ , \new_[22823]_ , \new_[22827]_ , \new_[22828]_ ,
    \new_[22829]_ , \new_[22833]_ , \new_[22834]_ , \new_[22838]_ ,
    \new_[22839]_ , \new_[22840]_ , \new_[22844]_ , \new_[22845]_ ,
    \new_[22849]_ , \new_[22850]_ , \new_[22851]_ , \new_[22855]_ ,
    \new_[22856]_ , \new_[22860]_ , \new_[22861]_ , \new_[22862]_ ,
    \new_[22866]_ , \new_[22867]_ , \new_[22871]_ , \new_[22872]_ ,
    \new_[22873]_ , \new_[22877]_ , \new_[22878]_ , \new_[22882]_ ,
    \new_[22883]_ , \new_[22884]_ , \new_[22888]_ , \new_[22889]_ ,
    \new_[22893]_ , \new_[22894]_ , \new_[22895]_ , \new_[22899]_ ,
    \new_[22900]_ , \new_[22904]_ , \new_[22905]_ , \new_[22906]_ ,
    \new_[22910]_ , \new_[22911]_ , \new_[22915]_ , \new_[22916]_ ,
    \new_[22917]_ , \new_[22921]_ , \new_[22922]_ , \new_[22926]_ ,
    \new_[22927]_ , \new_[22928]_ , \new_[22932]_ , \new_[22933]_ ,
    \new_[22937]_ , \new_[22938]_ , \new_[22939]_ , \new_[22943]_ ,
    \new_[22944]_ , \new_[22948]_ , \new_[22949]_ , \new_[22950]_ ,
    \new_[22954]_ , \new_[22955]_ , \new_[22959]_ , \new_[22960]_ ,
    \new_[22961]_ , \new_[22965]_ , \new_[22966]_ , \new_[22970]_ ,
    \new_[22971]_ , \new_[22972]_ , \new_[22976]_ , \new_[22977]_ ,
    \new_[22981]_ , \new_[22982]_ , \new_[22983]_ , \new_[22987]_ ,
    \new_[22988]_ , \new_[22992]_ , \new_[22993]_ , \new_[22994]_ ,
    \new_[22998]_ , \new_[22999]_ , \new_[23003]_ , \new_[23004]_ ,
    \new_[23005]_ , \new_[23009]_ , \new_[23010]_ , \new_[23014]_ ,
    \new_[23015]_ , \new_[23016]_ , \new_[23020]_ , \new_[23021]_ ,
    \new_[23025]_ , \new_[23026]_ , \new_[23027]_ , \new_[23031]_ ,
    \new_[23032]_ , \new_[23036]_ , \new_[23037]_ , \new_[23038]_ ,
    \new_[23042]_ , \new_[23043]_ , \new_[23047]_ , \new_[23048]_ ,
    \new_[23049]_ , \new_[23053]_ , \new_[23054]_ , \new_[23058]_ ,
    \new_[23059]_ , \new_[23060]_ , \new_[23064]_ , \new_[23065]_ ,
    \new_[23069]_ , \new_[23070]_ , \new_[23071]_ , \new_[23075]_ ,
    \new_[23076]_ , \new_[23080]_ , \new_[23081]_ , \new_[23082]_ ,
    \new_[23086]_ , \new_[23087]_ , \new_[23091]_ , \new_[23092]_ ,
    \new_[23093]_ , \new_[23097]_ , \new_[23098]_ , \new_[23102]_ ,
    \new_[23103]_ , \new_[23104]_ , \new_[23108]_ , \new_[23109]_ ,
    \new_[23113]_ , \new_[23114]_ , \new_[23115]_ , \new_[23119]_ ,
    \new_[23120]_ , \new_[23124]_ , \new_[23125]_ , \new_[23126]_ ,
    \new_[23130]_ , \new_[23131]_ , \new_[23135]_ , \new_[23136]_ ,
    \new_[23137]_ , \new_[23141]_ , \new_[23142]_ , \new_[23146]_ ,
    \new_[23147]_ , \new_[23148]_ , \new_[23152]_ , \new_[23153]_ ,
    \new_[23157]_ , \new_[23158]_ , \new_[23159]_ , \new_[23163]_ ,
    \new_[23164]_ , \new_[23168]_ , \new_[23169]_ , \new_[23170]_ ,
    \new_[23174]_ , \new_[23175]_ , \new_[23179]_ , \new_[23180]_ ,
    \new_[23181]_ , \new_[23185]_ , \new_[23186]_ , \new_[23190]_ ,
    \new_[23191]_ , \new_[23192]_ , \new_[23196]_ , \new_[23197]_ ,
    \new_[23201]_ , \new_[23202]_ , \new_[23203]_ , \new_[23207]_ ,
    \new_[23208]_ , \new_[23212]_ , \new_[23213]_ , \new_[23214]_ ,
    \new_[23218]_ , \new_[23219]_ , \new_[23223]_ , \new_[23224]_ ,
    \new_[23225]_ , \new_[23229]_ , \new_[23230]_ , \new_[23234]_ ,
    \new_[23235]_ , \new_[23236]_ , \new_[23240]_ , \new_[23241]_ ,
    \new_[23245]_ , \new_[23246]_ , \new_[23247]_ , \new_[23251]_ ,
    \new_[23252]_ , \new_[23256]_ , \new_[23257]_ , \new_[23258]_ ,
    \new_[23262]_ , \new_[23263]_ , \new_[23267]_ , \new_[23268]_ ,
    \new_[23269]_ , \new_[23273]_ , \new_[23274]_ , \new_[23278]_ ,
    \new_[23279]_ , \new_[23280]_ , \new_[23284]_ , \new_[23285]_ ,
    \new_[23289]_ , \new_[23290]_ , \new_[23291]_ , \new_[23295]_ ,
    \new_[23296]_ , \new_[23300]_ , \new_[23301]_ , \new_[23302]_ ,
    \new_[23306]_ , \new_[23307]_ , \new_[23311]_ , \new_[23312]_ ,
    \new_[23313]_ , \new_[23317]_ , \new_[23318]_ , \new_[23322]_ ,
    \new_[23323]_ , \new_[23324]_ , \new_[23328]_ , \new_[23329]_ ,
    \new_[23333]_ , \new_[23334]_ , \new_[23335]_ , \new_[23339]_ ,
    \new_[23340]_ , \new_[23344]_ , \new_[23345]_ , \new_[23346]_ ,
    \new_[23350]_ , \new_[23351]_ , \new_[23355]_ , \new_[23356]_ ,
    \new_[23357]_ , \new_[23361]_ , \new_[23362]_ , \new_[23366]_ ,
    \new_[23367]_ , \new_[23368]_ , \new_[23372]_ , \new_[23373]_ ,
    \new_[23377]_ , \new_[23378]_ , \new_[23379]_ , \new_[23383]_ ,
    \new_[23384]_ , \new_[23388]_ , \new_[23389]_ , \new_[23390]_ ,
    \new_[23394]_ , \new_[23395]_ , \new_[23399]_ , \new_[23400]_ ,
    \new_[23401]_ , \new_[23405]_ , \new_[23406]_ , \new_[23410]_ ,
    \new_[23411]_ , \new_[23412]_ , \new_[23416]_ , \new_[23417]_ ,
    \new_[23421]_ , \new_[23422]_ , \new_[23423]_ , \new_[23427]_ ,
    \new_[23428]_ , \new_[23432]_ , \new_[23433]_ , \new_[23434]_ ,
    \new_[23438]_ , \new_[23439]_ , \new_[23443]_ , \new_[23444]_ ,
    \new_[23445]_ , \new_[23449]_ , \new_[23450]_ , \new_[23454]_ ,
    \new_[23455]_ , \new_[23456]_ , \new_[23460]_ , \new_[23461]_ ,
    \new_[23465]_ , \new_[23466]_ , \new_[23467]_ , \new_[23471]_ ,
    \new_[23472]_ , \new_[23476]_ , \new_[23477]_ , \new_[23478]_ ,
    \new_[23482]_ , \new_[23483]_ , \new_[23487]_ , \new_[23488]_ ,
    \new_[23489]_ , \new_[23493]_ , \new_[23494]_ , \new_[23498]_ ,
    \new_[23499]_ , \new_[23500]_ , \new_[23504]_ , \new_[23505]_ ,
    \new_[23509]_ , \new_[23510]_ , \new_[23511]_ , \new_[23515]_ ,
    \new_[23516]_ , \new_[23520]_ , \new_[23521]_ , \new_[23522]_ ,
    \new_[23526]_ , \new_[23527]_ , \new_[23531]_ , \new_[23532]_ ,
    \new_[23533]_ , \new_[23537]_ , \new_[23538]_ , \new_[23542]_ ,
    \new_[23543]_ , \new_[23544]_ , \new_[23548]_ , \new_[23549]_ ,
    \new_[23553]_ , \new_[23554]_ , \new_[23555]_ , \new_[23559]_ ,
    \new_[23560]_ , \new_[23564]_ , \new_[23565]_ , \new_[23566]_ ,
    \new_[23570]_ , \new_[23571]_ , \new_[23575]_ , \new_[23576]_ ,
    \new_[23577]_ , \new_[23581]_ , \new_[23582]_ , \new_[23586]_ ,
    \new_[23587]_ , \new_[23588]_ , \new_[23592]_ , \new_[23593]_ ,
    \new_[23597]_ , \new_[23598]_ , \new_[23599]_ , \new_[23603]_ ,
    \new_[23604]_ , \new_[23608]_ , \new_[23609]_ , \new_[23610]_ ,
    \new_[23614]_ , \new_[23615]_ , \new_[23619]_ , \new_[23620]_ ,
    \new_[23621]_ , \new_[23625]_ , \new_[23626]_ , \new_[23630]_ ,
    \new_[23631]_ , \new_[23632]_ , \new_[23636]_ , \new_[23637]_ ,
    \new_[23641]_ , \new_[23642]_ , \new_[23643]_ , \new_[23647]_ ,
    \new_[23648]_ , \new_[23652]_ , \new_[23653]_ , \new_[23654]_ ,
    \new_[23658]_ , \new_[23659]_ , \new_[23663]_ , \new_[23664]_ ,
    \new_[23665]_ , \new_[23669]_ , \new_[23670]_ , \new_[23674]_ ,
    \new_[23675]_ , \new_[23676]_ , \new_[23680]_ , \new_[23681]_ ,
    \new_[23685]_ , \new_[23686]_ , \new_[23687]_ , \new_[23691]_ ,
    \new_[23692]_ , \new_[23696]_ , \new_[23697]_ , \new_[23698]_ ,
    \new_[23702]_ , \new_[23703]_ , \new_[23707]_ , \new_[23708]_ ,
    \new_[23709]_ , \new_[23713]_ , \new_[23714]_ , \new_[23718]_ ,
    \new_[23719]_ , \new_[23720]_ , \new_[23724]_ , \new_[23725]_ ,
    \new_[23729]_ , \new_[23730]_ , \new_[23731]_ , \new_[23735]_ ,
    \new_[23736]_ , \new_[23740]_ , \new_[23741]_ , \new_[23742]_ ,
    \new_[23746]_ , \new_[23747]_ , \new_[23751]_ , \new_[23752]_ ,
    \new_[23753]_ , \new_[23757]_ , \new_[23758]_ , \new_[23762]_ ,
    \new_[23763]_ , \new_[23764]_ , \new_[23768]_ , \new_[23769]_ ,
    \new_[23773]_ , \new_[23774]_ , \new_[23775]_ , \new_[23779]_ ,
    \new_[23780]_ , \new_[23784]_ , \new_[23785]_ , \new_[23786]_ ,
    \new_[23790]_ , \new_[23791]_ , \new_[23795]_ , \new_[23796]_ ,
    \new_[23797]_ , \new_[23801]_ , \new_[23802]_ , \new_[23806]_ ,
    \new_[23807]_ , \new_[23808]_ , \new_[23812]_ , \new_[23813]_ ,
    \new_[23817]_ , \new_[23818]_ , \new_[23819]_ , \new_[23823]_ ,
    \new_[23824]_ , \new_[23828]_ , \new_[23829]_ , \new_[23830]_ ,
    \new_[23834]_ , \new_[23835]_ , \new_[23839]_ , \new_[23840]_ ,
    \new_[23841]_ , \new_[23845]_ , \new_[23846]_ , \new_[23850]_ ,
    \new_[23851]_ , \new_[23852]_ , \new_[23856]_ , \new_[23857]_ ,
    \new_[23861]_ , \new_[23862]_ , \new_[23863]_ , \new_[23867]_ ,
    \new_[23868]_ , \new_[23872]_ , \new_[23873]_ , \new_[23874]_ ,
    \new_[23878]_ , \new_[23879]_ , \new_[23883]_ , \new_[23884]_ ,
    \new_[23885]_ , \new_[23889]_ , \new_[23890]_ , \new_[23894]_ ,
    \new_[23895]_ , \new_[23896]_ , \new_[23900]_ , \new_[23901]_ ,
    \new_[23905]_ , \new_[23906]_ , \new_[23907]_ , \new_[23911]_ ,
    \new_[23912]_ , \new_[23916]_ , \new_[23917]_ , \new_[23918]_ ,
    \new_[23922]_ , \new_[23923]_ , \new_[23927]_ , \new_[23928]_ ,
    \new_[23929]_ , \new_[23933]_ , \new_[23934]_ , \new_[23938]_ ,
    \new_[23939]_ , \new_[23940]_ , \new_[23944]_ , \new_[23945]_ ,
    \new_[23949]_ , \new_[23950]_ , \new_[23951]_ , \new_[23955]_ ,
    \new_[23956]_ , \new_[23960]_ , \new_[23961]_ , \new_[23962]_ ,
    \new_[23966]_ , \new_[23967]_ , \new_[23971]_ , \new_[23972]_ ,
    \new_[23973]_ , \new_[23977]_ , \new_[23978]_ , \new_[23982]_ ,
    \new_[23983]_ , \new_[23984]_ , \new_[23988]_ , \new_[23989]_ ,
    \new_[23993]_ , \new_[23994]_ , \new_[23995]_ , \new_[23999]_ ,
    \new_[24000]_ , \new_[24004]_ , \new_[24005]_ , \new_[24006]_ ,
    \new_[24010]_ , \new_[24011]_ , \new_[24015]_ , \new_[24016]_ ,
    \new_[24017]_ , \new_[24021]_ , \new_[24022]_ , \new_[24026]_ ,
    \new_[24027]_ , \new_[24028]_ , \new_[24032]_ , \new_[24033]_ ,
    \new_[24037]_ , \new_[24038]_ , \new_[24039]_ , \new_[24043]_ ,
    \new_[24044]_ , \new_[24048]_ , \new_[24049]_ , \new_[24050]_ ,
    \new_[24054]_ , \new_[24055]_ , \new_[24059]_ , \new_[24060]_ ,
    \new_[24061]_ , \new_[24065]_ , \new_[24066]_ , \new_[24070]_ ,
    \new_[24071]_ , \new_[24072]_ , \new_[24076]_ , \new_[24077]_ ,
    \new_[24081]_ , \new_[24082]_ , \new_[24083]_ , \new_[24087]_ ,
    \new_[24088]_ , \new_[24092]_ , \new_[24093]_ , \new_[24094]_ ,
    \new_[24098]_ , \new_[24099]_ , \new_[24103]_ , \new_[24104]_ ,
    \new_[24105]_ , \new_[24109]_ , \new_[24110]_ , \new_[24114]_ ,
    \new_[24115]_ , \new_[24116]_ , \new_[24120]_ , \new_[24121]_ ,
    \new_[24125]_ , \new_[24126]_ , \new_[24127]_ , \new_[24131]_ ,
    \new_[24132]_ , \new_[24136]_ , \new_[24137]_ , \new_[24138]_ ,
    \new_[24142]_ , \new_[24143]_ , \new_[24147]_ , \new_[24148]_ ,
    \new_[24149]_ , \new_[24153]_ , \new_[24154]_ , \new_[24158]_ ,
    \new_[24159]_ , \new_[24160]_ , \new_[24164]_ , \new_[24165]_ ,
    \new_[24169]_ , \new_[24170]_ , \new_[24171]_ , \new_[24175]_ ,
    \new_[24176]_ , \new_[24180]_ , \new_[24181]_ , \new_[24182]_ ,
    \new_[24186]_ , \new_[24187]_ , \new_[24191]_ , \new_[24192]_ ,
    \new_[24193]_ , \new_[24197]_ , \new_[24198]_ , \new_[24202]_ ,
    \new_[24203]_ , \new_[24204]_ , \new_[24208]_ , \new_[24209]_ ,
    \new_[24213]_ , \new_[24214]_ , \new_[24215]_ , \new_[24219]_ ,
    \new_[24220]_ , \new_[24224]_ , \new_[24225]_ , \new_[24226]_ ,
    \new_[24230]_ , \new_[24231]_ , \new_[24235]_ , \new_[24236]_ ,
    \new_[24237]_ , \new_[24241]_ , \new_[24242]_ , \new_[24246]_ ,
    \new_[24247]_ , \new_[24248]_ , \new_[24252]_ , \new_[24253]_ ,
    \new_[24257]_ , \new_[24258]_ , \new_[24259]_ , \new_[24263]_ ,
    \new_[24264]_ , \new_[24268]_ , \new_[24269]_ , \new_[24270]_ ,
    \new_[24274]_ , \new_[24275]_ , \new_[24279]_ , \new_[24280]_ ,
    \new_[24281]_ , \new_[24285]_ , \new_[24286]_ , \new_[24290]_ ,
    \new_[24291]_ , \new_[24292]_ , \new_[24296]_ , \new_[24297]_ ,
    \new_[24301]_ , \new_[24302]_ , \new_[24303]_ , \new_[24307]_ ,
    \new_[24308]_ , \new_[24312]_ , \new_[24313]_ , \new_[24314]_ ,
    \new_[24318]_ , \new_[24319]_ , \new_[24323]_ , \new_[24324]_ ,
    \new_[24325]_ , \new_[24329]_ , \new_[24330]_ , \new_[24334]_ ,
    \new_[24335]_ , \new_[24336]_ , \new_[24340]_ , \new_[24341]_ ,
    \new_[24345]_ , \new_[24346]_ , \new_[24347]_ , \new_[24351]_ ,
    \new_[24352]_ , \new_[24356]_ , \new_[24357]_ , \new_[24358]_ ,
    \new_[24362]_ , \new_[24363]_ , \new_[24367]_ , \new_[24368]_ ,
    \new_[24369]_ , \new_[24373]_ , \new_[24374]_ , \new_[24378]_ ,
    \new_[24379]_ , \new_[24380]_ , \new_[24384]_ , \new_[24385]_ ,
    \new_[24389]_ , \new_[24390]_ , \new_[24391]_ , \new_[24395]_ ,
    \new_[24396]_ , \new_[24400]_ , \new_[24401]_ , \new_[24402]_ ,
    \new_[24406]_ , \new_[24407]_ , \new_[24411]_ , \new_[24412]_ ,
    \new_[24413]_ , \new_[24417]_ , \new_[24418]_ , \new_[24422]_ ,
    \new_[24423]_ , \new_[24424]_ , \new_[24428]_ , \new_[24429]_ ,
    \new_[24433]_ , \new_[24434]_ , \new_[24435]_ , \new_[24439]_ ,
    \new_[24440]_ , \new_[24444]_ , \new_[24445]_ , \new_[24446]_ ,
    \new_[24450]_ , \new_[24451]_ , \new_[24455]_ , \new_[24456]_ ,
    \new_[24457]_ , \new_[24461]_ , \new_[24462]_ , \new_[24466]_ ,
    \new_[24467]_ , \new_[24468]_ , \new_[24472]_ , \new_[24473]_ ,
    \new_[24477]_ , \new_[24478]_ , \new_[24479]_ , \new_[24483]_ ,
    \new_[24484]_ , \new_[24488]_ , \new_[24489]_ , \new_[24490]_ ,
    \new_[24494]_ , \new_[24495]_ , \new_[24499]_ , \new_[24500]_ ,
    \new_[24501]_ , \new_[24505]_ , \new_[24506]_ , \new_[24510]_ ,
    \new_[24511]_ , \new_[24512]_ , \new_[24516]_ , \new_[24517]_ ,
    \new_[24521]_ , \new_[24522]_ , \new_[24523]_ , \new_[24527]_ ,
    \new_[24528]_ , \new_[24532]_ , \new_[24533]_ , \new_[24534]_ ,
    \new_[24538]_ , \new_[24539]_ , \new_[24543]_ , \new_[24544]_ ,
    \new_[24545]_ , \new_[24549]_ , \new_[24550]_ , \new_[24554]_ ,
    \new_[24555]_ , \new_[24556]_ , \new_[24560]_ , \new_[24561]_ ,
    \new_[24565]_ , \new_[24566]_ , \new_[24567]_ , \new_[24571]_ ,
    \new_[24572]_ , \new_[24576]_ , \new_[24577]_ , \new_[24578]_ ,
    \new_[24582]_ , \new_[24583]_ , \new_[24587]_ , \new_[24588]_ ,
    \new_[24589]_ , \new_[24593]_ , \new_[24594]_ , \new_[24598]_ ,
    \new_[24599]_ , \new_[24600]_ , \new_[24604]_ , \new_[24605]_ ,
    \new_[24609]_ , \new_[24610]_ , \new_[24611]_ , \new_[24615]_ ,
    \new_[24616]_ , \new_[24620]_ , \new_[24621]_ , \new_[24622]_ ,
    \new_[24626]_ , \new_[24627]_ , \new_[24631]_ , \new_[24632]_ ,
    \new_[24633]_ , \new_[24637]_ , \new_[24638]_ , \new_[24642]_ ,
    \new_[24643]_ , \new_[24644]_ , \new_[24648]_ , \new_[24649]_ ,
    \new_[24653]_ , \new_[24654]_ , \new_[24655]_ , \new_[24659]_ ,
    \new_[24660]_ , \new_[24664]_ , \new_[24665]_ , \new_[24666]_ ,
    \new_[24670]_ , \new_[24671]_ , \new_[24675]_ , \new_[24676]_ ,
    \new_[24677]_ , \new_[24681]_ , \new_[24682]_ , \new_[24686]_ ,
    \new_[24687]_ , \new_[24688]_ , \new_[24692]_ , \new_[24693]_ ,
    \new_[24697]_ , \new_[24698]_ , \new_[24699]_ , \new_[24703]_ ,
    \new_[24704]_ , \new_[24708]_ , \new_[24709]_ , \new_[24710]_ ,
    \new_[24714]_ , \new_[24715]_ , \new_[24719]_ , \new_[24720]_ ,
    \new_[24721]_ , \new_[24725]_ , \new_[24726]_ , \new_[24730]_ ,
    \new_[24731]_ , \new_[24732]_ , \new_[24736]_ , \new_[24737]_ ,
    \new_[24741]_ , \new_[24742]_ , \new_[24743]_ , \new_[24747]_ ,
    \new_[24748]_ , \new_[24752]_ , \new_[24753]_ , \new_[24754]_ ,
    \new_[24758]_ , \new_[24759]_ , \new_[24763]_ , \new_[24764]_ ,
    \new_[24765]_ , \new_[24769]_ , \new_[24770]_ , \new_[24774]_ ,
    \new_[24775]_ , \new_[24776]_ , \new_[24780]_ , \new_[24781]_ ,
    \new_[24785]_ , \new_[24786]_ , \new_[24787]_ , \new_[24791]_ ,
    \new_[24792]_ , \new_[24796]_ , \new_[24797]_ , \new_[24798]_ ,
    \new_[24802]_ , \new_[24803]_ , \new_[24807]_ , \new_[24808]_ ,
    \new_[24809]_ , \new_[24813]_ , \new_[24814]_ , \new_[24818]_ ,
    \new_[24819]_ , \new_[24820]_ , \new_[24824]_ , \new_[24825]_ ,
    \new_[24829]_ , \new_[24830]_ , \new_[24831]_ , \new_[24835]_ ,
    \new_[24836]_ , \new_[24840]_ , \new_[24841]_ , \new_[24842]_ ,
    \new_[24846]_ , \new_[24847]_ , \new_[24851]_ , \new_[24852]_ ,
    \new_[24853]_ , \new_[24857]_ , \new_[24858]_ , \new_[24862]_ ,
    \new_[24863]_ , \new_[24864]_ , \new_[24868]_ , \new_[24869]_ ,
    \new_[24873]_ , \new_[24874]_ , \new_[24875]_ , \new_[24879]_ ,
    \new_[24880]_ , \new_[24884]_ , \new_[24885]_ , \new_[24886]_ ,
    \new_[24890]_ , \new_[24891]_ , \new_[24895]_ , \new_[24896]_ ,
    \new_[24897]_ , \new_[24901]_ , \new_[24902]_ , \new_[24906]_ ,
    \new_[24907]_ , \new_[24908]_ , \new_[24912]_ , \new_[24913]_ ,
    \new_[24917]_ , \new_[24918]_ , \new_[24919]_ , \new_[24923]_ ,
    \new_[24924]_ , \new_[24928]_ , \new_[24929]_ , \new_[24930]_ ,
    \new_[24934]_ , \new_[24935]_ , \new_[24939]_ , \new_[24940]_ ,
    \new_[24941]_ , \new_[24945]_ , \new_[24946]_ , \new_[24950]_ ,
    \new_[24951]_ , \new_[24952]_ , \new_[24956]_ , \new_[24957]_ ,
    \new_[24961]_ , \new_[24962]_ , \new_[24963]_ , \new_[24967]_ ,
    \new_[24968]_ , \new_[24972]_ , \new_[24973]_ , \new_[24974]_ ,
    \new_[24978]_ , \new_[24979]_ , \new_[24983]_ , \new_[24984]_ ,
    \new_[24985]_ , \new_[24989]_ , \new_[24990]_ , \new_[24994]_ ,
    \new_[24995]_ , \new_[24996]_ , \new_[25000]_ , \new_[25001]_ ,
    \new_[25005]_ , \new_[25006]_ , \new_[25007]_ , \new_[25011]_ ,
    \new_[25012]_ , \new_[25016]_ , \new_[25017]_ , \new_[25018]_ ,
    \new_[25022]_ , \new_[25023]_ , \new_[25027]_ , \new_[25028]_ ,
    \new_[25029]_ , \new_[25033]_ , \new_[25034]_ , \new_[25038]_ ,
    \new_[25039]_ , \new_[25040]_ , \new_[25044]_ , \new_[25045]_ ,
    \new_[25049]_ , \new_[25050]_ , \new_[25051]_ , \new_[25055]_ ,
    \new_[25056]_ , \new_[25060]_ , \new_[25061]_ , \new_[25062]_ ,
    \new_[25066]_ , \new_[25067]_ , \new_[25071]_ , \new_[25072]_ ,
    \new_[25073]_ , \new_[25077]_ , \new_[25078]_ , \new_[25082]_ ,
    \new_[25083]_ , \new_[25084]_ , \new_[25088]_ , \new_[25089]_ ,
    \new_[25093]_ , \new_[25094]_ , \new_[25095]_ , \new_[25099]_ ,
    \new_[25100]_ , \new_[25104]_ , \new_[25105]_ , \new_[25106]_ ,
    \new_[25110]_ , \new_[25111]_ , \new_[25115]_ , \new_[25116]_ ,
    \new_[25117]_ , \new_[25121]_ , \new_[25122]_ , \new_[25126]_ ,
    \new_[25127]_ , \new_[25128]_ , \new_[25132]_ , \new_[25133]_ ,
    \new_[25137]_ , \new_[25138]_ , \new_[25139]_ , \new_[25143]_ ,
    \new_[25144]_ , \new_[25148]_ , \new_[25149]_ , \new_[25150]_ ,
    \new_[25154]_ , \new_[25155]_ , \new_[25159]_ , \new_[25160]_ ,
    \new_[25161]_ , \new_[25165]_ , \new_[25166]_ , \new_[25170]_ ,
    \new_[25171]_ , \new_[25172]_ , \new_[25176]_ , \new_[25177]_ ,
    \new_[25181]_ , \new_[25182]_ , \new_[25183]_ , \new_[25187]_ ,
    \new_[25188]_ , \new_[25192]_ , \new_[25193]_ , \new_[25194]_ ,
    \new_[25198]_ , \new_[25199]_ , \new_[25203]_ , \new_[25204]_ ,
    \new_[25205]_ , \new_[25209]_ , \new_[25210]_ , \new_[25214]_ ,
    \new_[25215]_ , \new_[25216]_ , \new_[25220]_ , \new_[25221]_ ,
    \new_[25225]_ , \new_[25226]_ , \new_[25227]_ , \new_[25231]_ ,
    \new_[25232]_ , \new_[25236]_ , \new_[25237]_ , \new_[25238]_ ,
    \new_[25242]_ , \new_[25243]_ , \new_[25247]_ , \new_[25248]_ ,
    \new_[25249]_ , \new_[25253]_ , \new_[25254]_ , \new_[25258]_ ,
    \new_[25259]_ , \new_[25260]_ , \new_[25264]_ , \new_[25265]_ ,
    \new_[25269]_ , \new_[25270]_ , \new_[25271]_ , \new_[25275]_ ,
    \new_[25276]_ , \new_[25280]_ , \new_[25281]_ , \new_[25282]_ ,
    \new_[25286]_ , \new_[25287]_ , \new_[25291]_ , \new_[25292]_ ,
    \new_[25293]_ , \new_[25297]_ , \new_[25298]_ , \new_[25302]_ ,
    \new_[25303]_ , \new_[25304]_ , \new_[25308]_ , \new_[25309]_ ,
    \new_[25313]_ , \new_[25314]_ , \new_[25315]_ , \new_[25319]_ ,
    \new_[25320]_ , \new_[25324]_ , \new_[25325]_ , \new_[25326]_ ,
    \new_[25330]_ , \new_[25331]_ , \new_[25335]_ , \new_[25336]_ ,
    \new_[25337]_ , \new_[25341]_ , \new_[25342]_ , \new_[25346]_ ,
    \new_[25347]_ , \new_[25348]_ , \new_[25352]_ , \new_[25353]_ ,
    \new_[25357]_ , \new_[25358]_ , \new_[25359]_ , \new_[25363]_ ,
    \new_[25364]_ , \new_[25368]_ , \new_[25369]_ , \new_[25370]_ ,
    \new_[25374]_ , \new_[25375]_ , \new_[25379]_ , \new_[25380]_ ,
    \new_[25381]_ , \new_[25385]_ , \new_[25386]_ , \new_[25390]_ ,
    \new_[25391]_ , \new_[25392]_ , \new_[25396]_ , \new_[25397]_ ,
    \new_[25401]_ , \new_[25402]_ , \new_[25403]_ , \new_[25407]_ ,
    \new_[25408]_ , \new_[25412]_ , \new_[25413]_ , \new_[25414]_ ,
    \new_[25418]_ , \new_[25419]_ , \new_[25423]_ , \new_[25424]_ ,
    \new_[25425]_ , \new_[25429]_ , \new_[25430]_ , \new_[25434]_ ,
    \new_[25435]_ , \new_[25436]_ , \new_[25440]_ , \new_[25441]_ ,
    \new_[25445]_ , \new_[25446]_ , \new_[25447]_ , \new_[25451]_ ,
    \new_[25452]_ , \new_[25456]_ , \new_[25457]_ , \new_[25458]_ ,
    \new_[25462]_ , \new_[25463]_ , \new_[25467]_ , \new_[25468]_ ,
    \new_[25469]_ , \new_[25473]_ , \new_[25474]_ , \new_[25478]_ ,
    \new_[25479]_ , \new_[25480]_ , \new_[25484]_ , \new_[25485]_ ,
    \new_[25489]_ , \new_[25490]_ , \new_[25491]_ , \new_[25495]_ ,
    \new_[25496]_ , \new_[25500]_ , \new_[25501]_ , \new_[25502]_ ,
    \new_[25506]_ , \new_[25507]_ , \new_[25511]_ , \new_[25512]_ ,
    \new_[25513]_ , \new_[25517]_ , \new_[25518]_ , \new_[25522]_ ,
    \new_[25523]_ , \new_[25524]_ , \new_[25528]_ , \new_[25529]_ ,
    \new_[25533]_ , \new_[25534]_ , \new_[25535]_ , \new_[25539]_ ,
    \new_[25540]_ , \new_[25544]_ , \new_[25545]_ , \new_[25546]_ ,
    \new_[25550]_ , \new_[25551]_ , \new_[25555]_ , \new_[25556]_ ,
    \new_[25557]_ , \new_[25561]_ , \new_[25562]_ , \new_[25566]_ ,
    \new_[25567]_ , \new_[25568]_ , \new_[25572]_ , \new_[25573]_ ,
    \new_[25577]_ , \new_[25578]_ , \new_[25579]_ , \new_[25583]_ ,
    \new_[25584]_ , \new_[25588]_ , \new_[25589]_ , \new_[25590]_ ,
    \new_[25594]_ , \new_[25595]_ , \new_[25599]_ , \new_[25600]_ ,
    \new_[25601]_ , \new_[25605]_ , \new_[25606]_ , \new_[25610]_ ,
    \new_[25611]_ , \new_[25612]_ , \new_[25616]_ , \new_[25617]_ ,
    \new_[25621]_ , \new_[25622]_ , \new_[25623]_ , \new_[25627]_ ,
    \new_[25628]_ , \new_[25632]_ , \new_[25633]_ , \new_[25634]_ ,
    \new_[25638]_ , \new_[25639]_ , \new_[25643]_ , \new_[25644]_ ,
    \new_[25645]_ , \new_[25649]_ , \new_[25650]_ , \new_[25654]_ ,
    \new_[25655]_ , \new_[25656]_ , \new_[25660]_ , \new_[25661]_ ,
    \new_[25665]_ , \new_[25666]_ , \new_[25667]_ , \new_[25671]_ ,
    \new_[25672]_ , \new_[25676]_ , \new_[25677]_ , \new_[25678]_ ,
    \new_[25682]_ , \new_[25683]_ , \new_[25687]_ , \new_[25688]_ ,
    \new_[25689]_ , \new_[25693]_ , \new_[25694]_ , \new_[25698]_ ,
    \new_[25699]_ , \new_[25700]_ , \new_[25704]_ , \new_[25705]_ ,
    \new_[25709]_ , \new_[25710]_ , \new_[25711]_ , \new_[25715]_ ,
    \new_[25716]_ , \new_[25720]_ , \new_[25721]_ , \new_[25722]_ ,
    \new_[25726]_ , \new_[25727]_ , \new_[25731]_ , \new_[25732]_ ,
    \new_[25733]_ , \new_[25737]_ , \new_[25738]_ , \new_[25742]_ ,
    \new_[25743]_ , \new_[25744]_ , \new_[25748]_ , \new_[25749]_ ,
    \new_[25753]_ , \new_[25754]_ , \new_[25755]_ , \new_[25759]_ ,
    \new_[25760]_ , \new_[25764]_ , \new_[25765]_ , \new_[25766]_ ,
    \new_[25770]_ , \new_[25771]_ , \new_[25775]_ , \new_[25776]_ ,
    \new_[25777]_ , \new_[25781]_ , \new_[25782]_ , \new_[25786]_ ,
    \new_[25787]_ , \new_[25788]_ , \new_[25792]_ , \new_[25793]_ ,
    \new_[25797]_ , \new_[25798]_ , \new_[25799]_ , \new_[25803]_ ,
    \new_[25804]_ , \new_[25808]_ , \new_[25809]_ , \new_[25810]_ ,
    \new_[25814]_ , \new_[25815]_ , \new_[25819]_ , \new_[25820]_ ,
    \new_[25821]_ , \new_[25825]_ , \new_[25826]_ , \new_[25830]_ ,
    \new_[25831]_ , \new_[25832]_ , \new_[25836]_ , \new_[25837]_ ,
    \new_[25841]_ , \new_[25842]_ , \new_[25843]_ , \new_[25847]_ ,
    \new_[25848]_ , \new_[25852]_ , \new_[25853]_ , \new_[25854]_ ,
    \new_[25858]_ , \new_[25859]_ , \new_[25863]_ , \new_[25864]_ ,
    \new_[25865]_ , \new_[25869]_ , \new_[25870]_ , \new_[25874]_ ,
    \new_[25875]_ , \new_[25876]_ , \new_[25880]_ , \new_[25881]_ ,
    \new_[25885]_ , \new_[25886]_ , \new_[25887]_ , \new_[25891]_ ,
    \new_[25892]_ , \new_[25896]_ , \new_[25897]_ , \new_[25898]_ ,
    \new_[25902]_ , \new_[25903]_ , \new_[25907]_ , \new_[25908]_ ,
    \new_[25909]_ , \new_[25913]_ , \new_[25914]_ , \new_[25918]_ ,
    \new_[25919]_ , \new_[25920]_ , \new_[25924]_ , \new_[25925]_ ,
    \new_[25929]_ , \new_[25930]_ , \new_[25931]_ , \new_[25935]_ ,
    \new_[25936]_ , \new_[25940]_ , \new_[25941]_ , \new_[25942]_ ,
    \new_[25946]_ , \new_[25947]_ , \new_[25951]_ , \new_[25952]_ ,
    \new_[25953]_ , \new_[25957]_ , \new_[25958]_ , \new_[25962]_ ,
    \new_[25963]_ , \new_[25964]_ , \new_[25968]_ , \new_[25969]_ ,
    \new_[25973]_ , \new_[25974]_ , \new_[25975]_ , \new_[25979]_ ,
    \new_[25980]_ , \new_[25984]_ , \new_[25985]_ , \new_[25986]_ ,
    \new_[25990]_ , \new_[25991]_ , \new_[25995]_ , \new_[25996]_ ,
    \new_[25997]_ , \new_[26001]_ , \new_[26002]_ , \new_[26006]_ ,
    \new_[26007]_ , \new_[26008]_ , \new_[26012]_ , \new_[26013]_ ,
    \new_[26017]_ , \new_[26018]_ , \new_[26019]_ , \new_[26023]_ ,
    \new_[26024]_ , \new_[26028]_ , \new_[26029]_ , \new_[26030]_ ,
    \new_[26034]_ , \new_[26035]_ , \new_[26039]_ , \new_[26040]_ ,
    \new_[26041]_ , \new_[26045]_ , \new_[26046]_ , \new_[26050]_ ,
    \new_[26051]_ , \new_[26052]_ , \new_[26056]_ , \new_[26057]_ ,
    \new_[26061]_ , \new_[26062]_ , \new_[26063]_ , \new_[26067]_ ,
    \new_[26068]_ , \new_[26072]_ , \new_[26073]_ , \new_[26074]_ ,
    \new_[26078]_ , \new_[26079]_ , \new_[26083]_ , \new_[26084]_ ,
    \new_[26085]_ , \new_[26089]_ , \new_[26090]_ , \new_[26094]_ ,
    \new_[26095]_ , \new_[26096]_ , \new_[26100]_ , \new_[26101]_ ,
    \new_[26105]_ , \new_[26106]_ , \new_[26107]_ , \new_[26111]_ ,
    \new_[26112]_ , \new_[26116]_ , \new_[26117]_ , \new_[26118]_ ,
    \new_[26122]_ , \new_[26123]_ , \new_[26127]_ , \new_[26128]_ ,
    \new_[26129]_ , \new_[26133]_ , \new_[26134]_ , \new_[26138]_ ,
    \new_[26139]_ , \new_[26140]_ , \new_[26144]_ , \new_[26145]_ ,
    \new_[26149]_ , \new_[26150]_ , \new_[26151]_ , \new_[26155]_ ,
    \new_[26156]_ , \new_[26160]_ , \new_[26161]_ , \new_[26162]_ ,
    \new_[26166]_ , \new_[26167]_ , \new_[26171]_ , \new_[26172]_ ,
    \new_[26173]_ , \new_[26177]_ , \new_[26178]_ , \new_[26182]_ ,
    \new_[26183]_ , \new_[26184]_ , \new_[26188]_ , \new_[26189]_ ,
    \new_[26193]_ , \new_[26194]_ , \new_[26195]_ , \new_[26199]_ ,
    \new_[26200]_ , \new_[26204]_ , \new_[26205]_ , \new_[26206]_ ,
    \new_[26210]_ , \new_[26211]_ , \new_[26215]_ , \new_[26216]_ ,
    \new_[26217]_ , \new_[26221]_ , \new_[26222]_ , \new_[26226]_ ,
    \new_[26227]_ , \new_[26228]_ , \new_[26232]_ , \new_[26233]_ ,
    \new_[26237]_ , \new_[26238]_ , \new_[26239]_ , \new_[26243]_ ,
    \new_[26244]_ , \new_[26248]_ , \new_[26249]_ , \new_[26250]_ ,
    \new_[26254]_ , \new_[26255]_ , \new_[26259]_ , \new_[26260]_ ,
    \new_[26261]_ , \new_[26265]_ , \new_[26266]_ , \new_[26270]_ ,
    \new_[26271]_ , \new_[26272]_ , \new_[26276]_ , \new_[26277]_ ,
    \new_[26281]_ , \new_[26282]_ , \new_[26283]_ , \new_[26287]_ ,
    \new_[26288]_ , \new_[26292]_ , \new_[26293]_ , \new_[26294]_ ,
    \new_[26298]_ , \new_[26299]_ , \new_[26303]_ , \new_[26304]_ ,
    \new_[26305]_ , \new_[26309]_ , \new_[26310]_ , \new_[26314]_ ,
    \new_[26315]_ , \new_[26316]_ , \new_[26320]_ , \new_[26321]_ ,
    \new_[26325]_ , \new_[26326]_ , \new_[26327]_ , \new_[26331]_ ,
    \new_[26332]_ , \new_[26336]_ , \new_[26337]_ , \new_[26338]_ ,
    \new_[26342]_ , \new_[26343]_ , \new_[26347]_ , \new_[26348]_ ,
    \new_[26349]_ , \new_[26353]_ , \new_[26354]_ , \new_[26358]_ ,
    \new_[26359]_ , \new_[26360]_ , \new_[26364]_ , \new_[26365]_ ,
    \new_[26369]_ , \new_[26370]_ , \new_[26371]_ , \new_[26375]_ ,
    \new_[26376]_ , \new_[26380]_ , \new_[26381]_ , \new_[26382]_ ,
    \new_[26386]_ , \new_[26387]_ , \new_[26391]_ , \new_[26392]_ ,
    \new_[26393]_ , \new_[26397]_ , \new_[26398]_ , \new_[26402]_ ,
    \new_[26403]_ , \new_[26404]_ , \new_[26408]_ , \new_[26409]_ ,
    \new_[26413]_ , \new_[26414]_ , \new_[26415]_ , \new_[26419]_ ,
    \new_[26420]_ , \new_[26424]_ , \new_[26425]_ , \new_[26426]_ ,
    \new_[26430]_ , \new_[26431]_ , \new_[26435]_ , \new_[26436]_ ,
    \new_[26437]_ , \new_[26441]_ , \new_[26442]_ , \new_[26446]_ ,
    \new_[26447]_ , \new_[26448]_ , \new_[26452]_ , \new_[26453]_ ,
    \new_[26457]_ , \new_[26458]_ , \new_[26459]_ , \new_[26463]_ ,
    \new_[26464]_ , \new_[26468]_ , \new_[26469]_ , \new_[26470]_ ,
    \new_[26474]_ , \new_[26475]_ , \new_[26479]_ , \new_[26480]_ ,
    \new_[26481]_ , \new_[26485]_ , \new_[26486]_ , \new_[26490]_ ,
    \new_[26491]_ , \new_[26492]_ , \new_[26496]_ , \new_[26497]_ ,
    \new_[26501]_ , \new_[26502]_ , \new_[26503]_ , \new_[26507]_ ,
    \new_[26508]_ , \new_[26512]_ , \new_[26513]_ , \new_[26514]_ ,
    \new_[26518]_ , \new_[26519]_ , \new_[26523]_ , \new_[26524]_ ,
    \new_[26525]_ , \new_[26529]_ , \new_[26530]_ , \new_[26534]_ ,
    \new_[26535]_ , \new_[26536]_ , \new_[26540]_ , \new_[26541]_ ,
    \new_[26545]_ , \new_[26546]_ , \new_[26547]_ , \new_[26551]_ ,
    \new_[26552]_ , \new_[26556]_ , \new_[26557]_ , \new_[26558]_ ,
    \new_[26562]_ , \new_[26563]_ , \new_[26567]_ , \new_[26568]_ ,
    \new_[26569]_ , \new_[26573]_ , \new_[26574]_ , \new_[26578]_ ,
    \new_[26579]_ , \new_[26580]_ , \new_[26584]_ , \new_[26585]_ ,
    \new_[26589]_ , \new_[26590]_ , \new_[26591]_ , \new_[26595]_ ,
    \new_[26596]_ , \new_[26600]_ , \new_[26601]_ , \new_[26602]_ ,
    \new_[26606]_ , \new_[26607]_ , \new_[26611]_ , \new_[26612]_ ,
    \new_[26613]_ , \new_[26617]_ , \new_[26618]_ , \new_[26622]_ ,
    \new_[26623]_ , \new_[26624]_ , \new_[26628]_ , \new_[26629]_ ,
    \new_[26633]_ , \new_[26634]_ , \new_[26635]_ , \new_[26639]_ ,
    \new_[26640]_ , \new_[26644]_ , \new_[26645]_ , \new_[26646]_ ,
    \new_[26650]_ , \new_[26651]_ , \new_[26655]_ , \new_[26656]_ ,
    \new_[26657]_ , \new_[26661]_ , \new_[26662]_ , \new_[26666]_ ,
    \new_[26667]_ , \new_[26668]_ , \new_[26672]_ , \new_[26673]_ ,
    \new_[26677]_ , \new_[26678]_ , \new_[26679]_ , \new_[26683]_ ,
    \new_[26684]_ , \new_[26688]_ , \new_[26689]_ , \new_[26690]_ ,
    \new_[26694]_ , \new_[26695]_ , \new_[26699]_ , \new_[26700]_ ,
    \new_[26701]_ , \new_[26705]_ , \new_[26706]_ , \new_[26710]_ ,
    \new_[26711]_ , \new_[26712]_ , \new_[26716]_ , \new_[26717]_ ,
    \new_[26721]_ , \new_[26722]_ , \new_[26723]_ , \new_[26727]_ ,
    \new_[26728]_ , \new_[26732]_ , \new_[26733]_ , \new_[26734]_ ,
    \new_[26738]_ , \new_[26739]_ , \new_[26743]_ , \new_[26744]_ ,
    \new_[26745]_ , \new_[26749]_ , \new_[26750]_ , \new_[26754]_ ,
    \new_[26755]_ , \new_[26756]_ , \new_[26760]_ , \new_[26761]_ ,
    \new_[26765]_ , \new_[26766]_ , \new_[26767]_ , \new_[26771]_ ,
    \new_[26772]_ , \new_[26776]_ , \new_[26777]_ , \new_[26778]_ ,
    \new_[26782]_ , \new_[26783]_ , \new_[26787]_ , \new_[26788]_ ,
    \new_[26789]_ , \new_[26793]_ , \new_[26794]_ , \new_[26798]_ ,
    \new_[26799]_ , \new_[26800]_ , \new_[26804]_ , \new_[26805]_ ,
    \new_[26809]_ , \new_[26810]_ , \new_[26811]_ , \new_[26815]_ ,
    \new_[26816]_ , \new_[26820]_ , \new_[26821]_ , \new_[26822]_ ,
    \new_[26826]_ , \new_[26827]_ , \new_[26831]_ , \new_[26832]_ ,
    \new_[26833]_ , \new_[26837]_ , \new_[26838]_ , \new_[26842]_ ,
    \new_[26843]_ , \new_[26844]_ , \new_[26848]_ , \new_[26849]_ ,
    \new_[26853]_ , \new_[26854]_ , \new_[26855]_ , \new_[26859]_ ,
    \new_[26860]_ , \new_[26864]_ , \new_[26865]_ , \new_[26866]_ ,
    \new_[26870]_ , \new_[26871]_ , \new_[26875]_ , \new_[26876]_ ,
    \new_[26877]_ , \new_[26881]_ , \new_[26882]_ , \new_[26886]_ ,
    \new_[26887]_ , \new_[26888]_ , \new_[26892]_ , \new_[26893]_ ,
    \new_[26897]_ , \new_[26898]_ , \new_[26899]_ , \new_[26903]_ ,
    \new_[26904]_ , \new_[26908]_ , \new_[26909]_ , \new_[26910]_ ,
    \new_[26914]_ , \new_[26915]_ , \new_[26919]_ , \new_[26920]_ ,
    \new_[26921]_ , \new_[26925]_ , \new_[26926]_ , \new_[26930]_ ,
    \new_[26931]_ , \new_[26932]_ , \new_[26936]_ , \new_[26937]_ ,
    \new_[26941]_ , \new_[26942]_ , \new_[26943]_ , \new_[26947]_ ,
    \new_[26948]_ , \new_[26952]_ , \new_[26953]_ , \new_[26954]_ ,
    \new_[26958]_ , \new_[26959]_ , \new_[26963]_ , \new_[26964]_ ,
    \new_[26965]_ , \new_[26969]_ , \new_[26970]_ , \new_[26974]_ ,
    \new_[26975]_ , \new_[26976]_ , \new_[26980]_ , \new_[26981]_ ,
    \new_[26985]_ , \new_[26986]_ , \new_[26987]_ , \new_[26991]_ ,
    \new_[26992]_ , \new_[26996]_ , \new_[26997]_ , \new_[26998]_ ,
    \new_[27002]_ , \new_[27003]_ , \new_[27007]_ , \new_[27008]_ ,
    \new_[27009]_ , \new_[27013]_ , \new_[27014]_ , \new_[27018]_ ,
    \new_[27019]_ , \new_[27020]_ , \new_[27024]_ , \new_[27025]_ ,
    \new_[27029]_ , \new_[27030]_ , \new_[27031]_ , \new_[27035]_ ,
    \new_[27036]_ , \new_[27040]_ , \new_[27041]_ , \new_[27042]_ ,
    \new_[27046]_ , \new_[27047]_ , \new_[27051]_ , \new_[27052]_ ,
    \new_[27053]_ , \new_[27057]_ , \new_[27058]_ , \new_[27062]_ ,
    \new_[27063]_ , \new_[27064]_ , \new_[27068]_ , \new_[27069]_ ,
    \new_[27073]_ , \new_[27074]_ , \new_[27075]_ , \new_[27079]_ ,
    \new_[27080]_ , \new_[27084]_ , \new_[27085]_ , \new_[27086]_ ,
    \new_[27090]_ , \new_[27091]_ , \new_[27095]_ , \new_[27096]_ ,
    \new_[27097]_ , \new_[27101]_ , \new_[27102]_ , \new_[27106]_ ,
    \new_[27107]_ , \new_[27108]_ , \new_[27112]_ , \new_[27113]_ ,
    \new_[27117]_ , \new_[27118]_ , \new_[27119]_ , \new_[27123]_ ,
    \new_[27124]_ , \new_[27128]_ , \new_[27129]_ , \new_[27130]_ ,
    \new_[27134]_ , \new_[27135]_ , \new_[27139]_ , \new_[27140]_ ,
    \new_[27141]_ , \new_[27145]_ , \new_[27146]_ , \new_[27150]_ ,
    \new_[27151]_ , \new_[27152]_ , \new_[27156]_ , \new_[27157]_ ,
    \new_[27161]_ , \new_[27162]_ , \new_[27163]_ , \new_[27167]_ ,
    \new_[27168]_ , \new_[27172]_ , \new_[27173]_ , \new_[27174]_ ,
    \new_[27178]_ , \new_[27179]_ , \new_[27183]_ , \new_[27184]_ ,
    \new_[27185]_ , \new_[27189]_ , \new_[27190]_ , \new_[27194]_ ,
    \new_[27195]_ , \new_[27196]_ , \new_[27200]_ , \new_[27201]_ ,
    \new_[27205]_ , \new_[27206]_ , \new_[27207]_ , \new_[27211]_ ,
    \new_[27212]_ , \new_[27216]_ , \new_[27217]_ , \new_[27218]_ ,
    \new_[27222]_ , \new_[27223]_ , \new_[27227]_ , \new_[27228]_ ,
    \new_[27229]_ , \new_[27233]_ , \new_[27234]_ , \new_[27238]_ ,
    \new_[27239]_ , \new_[27240]_ , \new_[27244]_ , \new_[27245]_ ,
    \new_[27249]_ , \new_[27250]_ , \new_[27251]_ , \new_[27255]_ ,
    \new_[27256]_ , \new_[27260]_ , \new_[27261]_ , \new_[27262]_ ,
    \new_[27266]_ , \new_[27267]_ , \new_[27271]_ , \new_[27272]_ ,
    \new_[27273]_ , \new_[27277]_ , \new_[27278]_ , \new_[27282]_ ,
    \new_[27283]_ , \new_[27284]_ , \new_[27288]_ , \new_[27289]_ ,
    \new_[27293]_ , \new_[27294]_ , \new_[27295]_ , \new_[27299]_ ,
    \new_[27300]_ , \new_[27304]_ , \new_[27305]_ , \new_[27306]_ ,
    \new_[27310]_ , \new_[27311]_ , \new_[27315]_ , \new_[27316]_ ,
    \new_[27317]_ , \new_[27321]_ , \new_[27322]_ , \new_[27326]_ ,
    \new_[27327]_ , \new_[27328]_ , \new_[27332]_ , \new_[27333]_ ,
    \new_[27337]_ , \new_[27338]_ , \new_[27339]_ , \new_[27343]_ ,
    \new_[27344]_ , \new_[27348]_ , \new_[27349]_ , \new_[27350]_ ,
    \new_[27354]_ , \new_[27355]_ , \new_[27359]_ , \new_[27360]_ ,
    \new_[27361]_ , \new_[27365]_ , \new_[27366]_ , \new_[27370]_ ,
    \new_[27371]_ , \new_[27372]_ , \new_[27376]_ , \new_[27377]_ ,
    \new_[27381]_ , \new_[27382]_ , \new_[27383]_ , \new_[27387]_ ,
    \new_[27388]_ , \new_[27392]_ , \new_[27393]_ , \new_[27394]_ ,
    \new_[27398]_ , \new_[27399]_ , \new_[27403]_ , \new_[27404]_ ,
    \new_[27405]_ , \new_[27409]_ , \new_[27410]_ , \new_[27414]_ ,
    \new_[27415]_ , \new_[27416]_ , \new_[27420]_ , \new_[27421]_ ,
    \new_[27425]_ , \new_[27426]_ , \new_[27427]_ , \new_[27431]_ ,
    \new_[27432]_ , \new_[27436]_ , \new_[27437]_ , \new_[27438]_ ,
    \new_[27442]_ , \new_[27443]_ , \new_[27447]_ , \new_[27448]_ ,
    \new_[27449]_ , \new_[27453]_ , \new_[27454]_ , \new_[27458]_ ,
    \new_[27459]_ , \new_[27460]_ , \new_[27464]_ , \new_[27465]_ ,
    \new_[27469]_ , \new_[27470]_ , \new_[27471]_ , \new_[27475]_ ,
    \new_[27476]_ , \new_[27480]_ , \new_[27481]_ , \new_[27482]_ ,
    \new_[27486]_ , \new_[27487]_ , \new_[27491]_ , \new_[27492]_ ,
    \new_[27493]_ , \new_[27497]_ , \new_[27498]_ , \new_[27502]_ ,
    \new_[27503]_ , \new_[27504]_ , \new_[27508]_ , \new_[27509]_ ,
    \new_[27513]_ , \new_[27514]_ , \new_[27515]_ , \new_[27519]_ ,
    \new_[27520]_ , \new_[27524]_ , \new_[27525]_ , \new_[27526]_ ,
    \new_[27530]_ , \new_[27531]_ , \new_[27535]_ , \new_[27536]_ ,
    \new_[27537]_ , \new_[27541]_ , \new_[27542]_ , \new_[27546]_ ,
    \new_[27547]_ , \new_[27548]_ , \new_[27552]_ , \new_[27553]_ ,
    \new_[27557]_ , \new_[27558]_ , \new_[27559]_ , \new_[27563]_ ,
    \new_[27564]_ , \new_[27568]_ , \new_[27569]_ , \new_[27570]_ ,
    \new_[27574]_ , \new_[27575]_ , \new_[27579]_ , \new_[27580]_ ,
    \new_[27581]_ , \new_[27585]_ , \new_[27586]_ , \new_[27590]_ ,
    \new_[27591]_ , \new_[27592]_ , \new_[27596]_ , \new_[27597]_ ,
    \new_[27601]_ , \new_[27602]_ , \new_[27603]_ , \new_[27607]_ ,
    \new_[27608]_ , \new_[27612]_ , \new_[27613]_ , \new_[27614]_ ,
    \new_[27618]_ , \new_[27619]_ , \new_[27623]_ , \new_[27624]_ ,
    \new_[27625]_ , \new_[27629]_ , \new_[27630]_ , \new_[27634]_ ,
    \new_[27635]_ , \new_[27636]_ , \new_[27640]_ , \new_[27641]_ ,
    \new_[27645]_ , \new_[27646]_ , \new_[27647]_ , \new_[27651]_ ,
    \new_[27652]_ , \new_[27656]_ , \new_[27657]_ , \new_[27658]_ ,
    \new_[27662]_ , \new_[27663]_ , \new_[27667]_ , \new_[27668]_ ,
    \new_[27669]_ , \new_[27673]_ , \new_[27674]_ , \new_[27678]_ ,
    \new_[27679]_ , \new_[27680]_ , \new_[27684]_ , \new_[27685]_ ,
    \new_[27689]_ , \new_[27690]_ , \new_[27691]_ , \new_[27695]_ ,
    \new_[27696]_ , \new_[27700]_ , \new_[27701]_ , \new_[27702]_ ,
    \new_[27706]_ , \new_[27707]_ , \new_[27711]_ , \new_[27712]_ ,
    \new_[27713]_ , \new_[27717]_ , \new_[27718]_ , \new_[27722]_ ,
    \new_[27723]_ , \new_[27724]_ , \new_[27728]_ , \new_[27729]_ ,
    \new_[27733]_ , \new_[27734]_ , \new_[27735]_ , \new_[27739]_ ,
    \new_[27740]_ , \new_[27744]_ , \new_[27745]_ , \new_[27746]_ ,
    \new_[27750]_ , \new_[27751]_ , \new_[27755]_ , \new_[27756]_ ,
    \new_[27757]_ , \new_[27761]_ , \new_[27762]_ , \new_[27766]_ ,
    \new_[27767]_ , \new_[27768]_ , \new_[27772]_ , \new_[27773]_ ,
    \new_[27777]_ , \new_[27778]_ , \new_[27779]_ , \new_[27783]_ ,
    \new_[27784]_ , \new_[27788]_ , \new_[27789]_ , \new_[27790]_ ,
    \new_[27794]_ , \new_[27795]_ , \new_[27799]_ , \new_[27800]_ ,
    \new_[27801]_ , \new_[27805]_ , \new_[27806]_ , \new_[27810]_ ,
    \new_[27811]_ , \new_[27812]_ , \new_[27816]_ , \new_[27817]_ ,
    \new_[27821]_ , \new_[27822]_ , \new_[27823]_ , \new_[27827]_ ,
    \new_[27828]_ , \new_[27832]_ , \new_[27833]_ , \new_[27834]_ ,
    \new_[27838]_ , \new_[27839]_ , \new_[27843]_ , \new_[27844]_ ,
    \new_[27845]_ , \new_[27849]_ , \new_[27850]_ , \new_[27854]_ ,
    \new_[27855]_ , \new_[27856]_ , \new_[27860]_ , \new_[27861]_ ,
    \new_[27865]_ , \new_[27866]_ , \new_[27867]_ , \new_[27871]_ ,
    \new_[27872]_ , \new_[27876]_ , \new_[27877]_ , \new_[27878]_ ,
    \new_[27882]_ , \new_[27883]_ , \new_[27887]_ , \new_[27888]_ ,
    \new_[27889]_ , \new_[27893]_ , \new_[27894]_ , \new_[27898]_ ,
    \new_[27899]_ , \new_[27900]_ , \new_[27904]_ , \new_[27905]_ ,
    \new_[27909]_ , \new_[27910]_ , \new_[27911]_ , \new_[27915]_ ,
    \new_[27916]_ , \new_[27920]_ , \new_[27921]_ , \new_[27922]_ ,
    \new_[27926]_ , \new_[27927]_ , \new_[27931]_ , \new_[27932]_ ,
    \new_[27933]_ , \new_[27937]_ , \new_[27938]_ , \new_[27942]_ ,
    \new_[27943]_ , \new_[27944]_ , \new_[27948]_ , \new_[27949]_ ,
    \new_[27953]_ , \new_[27954]_ , \new_[27955]_ , \new_[27959]_ ,
    \new_[27960]_ , \new_[27964]_ , \new_[27965]_ , \new_[27966]_ ,
    \new_[27970]_ , \new_[27971]_ , \new_[27975]_ , \new_[27976]_ ,
    \new_[27977]_ , \new_[27981]_ , \new_[27982]_ , \new_[27986]_ ,
    \new_[27987]_ , \new_[27988]_ , \new_[27992]_ , \new_[27993]_ ,
    \new_[27997]_ , \new_[27998]_ , \new_[27999]_ , \new_[28003]_ ,
    \new_[28004]_ , \new_[28008]_ , \new_[28009]_ , \new_[28010]_ ,
    \new_[28014]_ , \new_[28015]_ , \new_[28019]_ , \new_[28020]_ ,
    \new_[28021]_ , \new_[28025]_ , \new_[28026]_ , \new_[28030]_ ,
    \new_[28031]_ , \new_[28032]_ , \new_[28036]_ , \new_[28037]_ ,
    \new_[28041]_ , \new_[28042]_ , \new_[28043]_ , \new_[28047]_ ,
    \new_[28048]_ , \new_[28052]_ , \new_[28053]_ , \new_[28054]_ ,
    \new_[28058]_ , \new_[28059]_ , \new_[28063]_ , \new_[28064]_ ,
    \new_[28065]_ , \new_[28069]_ , \new_[28070]_ , \new_[28074]_ ,
    \new_[28075]_ , \new_[28076]_ , \new_[28080]_ , \new_[28081]_ ,
    \new_[28085]_ , \new_[28086]_ , \new_[28087]_ , \new_[28091]_ ,
    \new_[28092]_ , \new_[28096]_ , \new_[28097]_ , \new_[28098]_ ,
    \new_[28102]_ , \new_[28103]_ , \new_[28107]_ , \new_[28108]_ ,
    \new_[28109]_ , \new_[28113]_ , \new_[28114]_ , \new_[28118]_ ,
    \new_[28119]_ , \new_[28120]_ , \new_[28124]_ , \new_[28125]_ ,
    \new_[28129]_ , \new_[28130]_ , \new_[28131]_ , \new_[28135]_ ,
    \new_[28136]_ , \new_[28140]_ , \new_[28141]_ , \new_[28142]_ ,
    \new_[28146]_ , \new_[28147]_ , \new_[28151]_ , \new_[28152]_ ,
    \new_[28153]_ , \new_[28157]_ , \new_[28158]_ , \new_[28162]_ ,
    \new_[28163]_ , \new_[28164]_ , \new_[28168]_ , \new_[28169]_ ,
    \new_[28173]_ , \new_[28174]_ , \new_[28175]_ , \new_[28179]_ ,
    \new_[28180]_ , \new_[28184]_ , \new_[28185]_ , \new_[28186]_ ,
    \new_[28190]_ , \new_[28191]_ , \new_[28195]_ , \new_[28196]_ ,
    \new_[28197]_ , \new_[28201]_ , \new_[28202]_ , \new_[28206]_ ,
    \new_[28207]_ , \new_[28208]_ , \new_[28212]_ , \new_[28213]_ ,
    \new_[28217]_ , \new_[28218]_ , \new_[28219]_ , \new_[28223]_ ,
    \new_[28224]_ , \new_[28228]_ , \new_[28229]_ , \new_[28230]_ ,
    \new_[28234]_ , \new_[28235]_ , \new_[28239]_ , \new_[28240]_ ,
    \new_[28241]_ , \new_[28245]_ , \new_[28246]_ , \new_[28250]_ ,
    \new_[28251]_ , \new_[28252]_ , \new_[28256]_ , \new_[28257]_ ,
    \new_[28261]_ , \new_[28262]_ , \new_[28263]_ , \new_[28267]_ ,
    \new_[28268]_ , \new_[28272]_ , \new_[28273]_ , \new_[28274]_ ,
    \new_[28278]_ , \new_[28279]_ , \new_[28283]_ , \new_[28284]_ ,
    \new_[28285]_ , \new_[28289]_ , \new_[28290]_ , \new_[28294]_ ,
    \new_[28295]_ , \new_[28296]_ , \new_[28300]_ , \new_[28301]_ ,
    \new_[28305]_ , \new_[28306]_ , \new_[28307]_ , \new_[28311]_ ,
    \new_[28312]_ , \new_[28316]_ , \new_[28317]_ , \new_[28318]_ ,
    \new_[28322]_ , \new_[28323]_ , \new_[28327]_ , \new_[28328]_ ,
    \new_[28329]_ , \new_[28333]_ , \new_[28334]_ , \new_[28338]_ ,
    \new_[28339]_ , \new_[28340]_ , \new_[28344]_ , \new_[28345]_ ,
    \new_[28349]_ , \new_[28350]_ , \new_[28351]_ , \new_[28355]_ ,
    \new_[28356]_ , \new_[28360]_ , \new_[28361]_ , \new_[28362]_ ,
    \new_[28366]_ , \new_[28367]_ , \new_[28371]_ , \new_[28372]_ ,
    \new_[28373]_ , \new_[28377]_ , \new_[28378]_ , \new_[28382]_ ,
    \new_[28383]_ , \new_[28384]_ , \new_[28388]_ , \new_[28389]_ ,
    \new_[28393]_ , \new_[28394]_ , \new_[28395]_ , \new_[28399]_ ,
    \new_[28400]_ , \new_[28404]_ , \new_[28405]_ , \new_[28406]_ ,
    \new_[28410]_ , \new_[28411]_ , \new_[28415]_ , \new_[28416]_ ,
    \new_[28417]_ , \new_[28421]_ , \new_[28422]_ , \new_[28426]_ ,
    \new_[28427]_ , \new_[28428]_ , \new_[28432]_ , \new_[28433]_ ,
    \new_[28437]_ , \new_[28438]_ , \new_[28439]_ , \new_[28443]_ ,
    \new_[28444]_ , \new_[28448]_ , \new_[28449]_ , \new_[28450]_ ,
    \new_[28454]_ , \new_[28455]_ , \new_[28459]_ , \new_[28460]_ ,
    \new_[28461]_ , \new_[28465]_ , \new_[28466]_ , \new_[28470]_ ,
    \new_[28471]_ , \new_[28472]_ , \new_[28476]_ , \new_[28477]_ ,
    \new_[28481]_ , \new_[28482]_ , \new_[28483]_ , \new_[28487]_ ,
    \new_[28488]_ , \new_[28492]_ , \new_[28493]_ , \new_[28494]_ ,
    \new_[28498]_ , \new_[28499]_ , \new_[28503]_ , \new_[28504]_ ,
    \new_[28505]_ , \new_[28509]_ , \new_[28510]_ , \new_[28514]_ ,
    \new_[28515]_ , \new_[28516]_ , \new_[28520]_ , \new_[28521]_ ,
    \new_[28525]_ , \new_[28526]_ , \new_[28527]_ , \new_[28531]_ ,
    \new_[28532]_ , \new_[28536]_ , \new_[28537]_ , \new_[28538]_ ,
    \new_[28542]_ , \new_[28543]_ , \new_[28547]_ , \new_[28548]_ ,
    \new_[28549]_ , \new_[28553]_ , \new_[28554]_ , \new_[28558]_ ,
    \new_[28559]_ , \new_[28560]_ , \new_[28564]_ , \new_[28565]_ ,
    \new_[28569]_ , \new_[28570]_ , \new_[28571]_ , \new_[28575]_ ,
    \new_[28576]_ , \new_[28580]_ , \new_[28581]_ , \new_[28582]_ ,
    \new_[28586]_ , \new_[28587]_ , \new_[28591]_ , \new_[28592]_ ,
    \new_[28593]_ , \new_[28597]_ , \new_[28598]_ , \new_[28602]_ ,
    \new_[28603]_ , \new_[28604]_ , \new_[28608]_ , \new_[28609]_ ,
    \new_[28613]_ , \new_[28614]_ , \new_[28615]_ , \new_[28619]_ ,
    \new_[28620]_ , \new_[28624]_ , \new_[28625]_ , \new_[28626]_ ,
    \new_[28630]_ , \new_[28631]_ , \new_[28635]_ , \new_[28636]_ ,
    \new_[28637]_ , \new_[28641]_ , \new_[28642]_ , \new_[28646]_ ,
    \new_[28647]_ , \new_[28648]_ , \new_[28652]_ , \new_[28653]_ ,
    \new_[28657]_ , \new_[28658]_ , \new_[28659]_ , \new_[28663]_ ,
    \new_[28664]_ , \new_[28668]_ , \new_[28669]_ , \new_[28670]_ ,
    \new_[28674]_ , \new_[28675]_ , \new_[28679]_ , \new_[28680]_ ,
    \new_[28681]_ , \new_[28685]_ , \new_[28686]_ , \new_[28690]_ ,
    \new_[28691]_ , \new_[28692]_ , \new_[28696]_ , \new_[28697]_ ,
    \new_[28701]_ , \new_[28702]_ , \new_[28703]_ , \new_[28707]_ ,
    \new_[28708]_ , \new_[28712]_ , \new_[28713]_ , \new_[28714]_ ,
    \new_[28718]_ , \new_[28719]_ , \new_[28723]_ , \new_[28724]_ ,
    \new_[28725]_ , \new_[28729]_ , \new_[28730]_ , \new_[28734]_ ,
    \new_[28735]_ , \new_[28736]_ , \new_[28740]_ , \new_[28741]_ ,
    \new_[28745]_ , \new_[28746]_ , \new_[28747]_ , \new_[28751]_ ,
    \new_[28752]_ , \new_[28756]_ , \new_[28757]_ , \new_[28758]_ ,
    \new_[28762]_ , \new_[28763]_ , \new_[28767]_ , \new_[28768]_ ,
    \new_[28769]_ , \new_[28773]_ , \new_[28774]_ , \new_[28778]_ ,
    \new_[28779]_ , \new_[28780]_ , \new_[28784]_ , \new_[28785]_ ,
    \new_[28789]_ , \new_[28790]_ , \new_[28791]_ , \new_[28795]_ ,
    \new_[28796]_ , \new_[28800]_ , \new_[28801]_ , \new_[28802]_ ,
    \new_[28806]_ , \new_[28807]_ , \new_[28811]_ , \new_[28812]_ ,
    \new_[28813]_ , \new_[28817]_ , \new_[28818]_ , \new_[28822]_ ,
    \new_[28823]_ , \new_[28824]_ , \new_[28828]_ , \new_[28829]_ ,
    \new_[28833]_ , \new_[28834]_ , \new_[28835]_ , \new_[28839]_ ,
    \new_[28840]_ , \new_[28844]_ , \new_[28845]_ , \new_[28846]_ ,
    \new_[28850]_ , \new_[28851]_ , \new_[28855]_ , \new_[28856]_ ,
    \new_[28857]_ , \new_[28861]_ , \new_[28862]_ , \new_[28866]_ ,
    \new_[28867]_ , \new_[28868]_ , \new_[28872]_ , \new_[28873]_ ,
    \new_[28877]_ , \new_[28878]_ , \new_[28879]_ , \new_[28883]_ ,
    \new_[28884]_ , \new_[28888]_ , \new_[28889]_ , \new_[28890]_ ,
    \new_[28894]_ , \new_[28895]_ , \new_[28899]_ , \new_[28900]_ ,
    \new_[28901]_ , \new_[28905]_ , \new_[28906]_ , \new_[28910]_ ,
    \new_[28911]_ , \new_[28912]_ , \new_[28916]_ , \new_[28917]_ ,
    \new_[28921]_ , \new_[28922]_ , \new_[28923]_ , \new_[28927]_ ,
    \new_[28928]_ , \new_[28932]_ , \new_[28933]_ , \new_[28934]_ ,
    \new_[28938]_ , \new_[28939]_ , \new_[28943]_ , \new_[28944]_ ,
    \new_[28945]_ , \new_[28949]_ , \new_[28950]_ , \new_[28954]_ ,
    \new_[28955]_ , \new_[28956]_ , \new_[28960]_ , \new_[28961]_ ,
    \new_[28965]_ , \new_[28966]_ , \new_[28967]_ , \new_[28971]_ ,
    \new_[28972]_ , \new_[28976]_ , \new_[28977]_ , \new_[28978]_ ,
    \new_[28982]_ , \new_[28983]_ , \new_[28987]_ , \new_[28988]_ ,
    \new_[28989]_ , \new_[28993]_ , \new_[28994]_ , \new_[28998]_ ,
    \new_[28999]_ , \new_[29000]_ , \new_[29004]_ , \new_[29005]_ ,
    \new_[29009]_ , \new_[29010]_ , \new_[29011]_ , \new_[29015]_ ,
    \new_[29016]_ , \new_[29020]_ , \new_[29021]_ , \new_[29022]_ ,
    \new_[29026]_ , \new_[29027]_ , \new_[29031]_ , \new_[29032]_ ,
    \new_[29033]_ , \new_[29037]_ , \new_[29038]_ , \new_[29042]_ ,
    \new_[29043]_ , \new_[29044]_ , \new_[29048]_ , \new_[29049]_ ,
    \new_[29053]_ , \new_[29054]_ , \new_[29055]_ , \new_[29059]_ ,
    \new_[29060]_ , \new_[29064]_ , \new_[29065]_ , \new_[29066]_ ,
    \new_[29070]_ , \new_[29071]_ , \new_[29075]_ , \new_[29076]_ ,
    \new_[29077]_ , \new_[29081]_ , \new_[29082]_ , \new_[29086]_ ,
    \new_[29087]_ , \new_[29088]_ , \new_[29092]_ , \new_[29093]_ ,
    \new_[29097]_ , \new_[29098]_ , \new_[29099]_ , \new_[29103]_ ,
    \new_[29104]_ , \new_[29108]_ , \new_[29109]_ , \new_[29110]_ ,
    \new_[29114]_ , \new_[29115]_ , \new_[29119]_ , \new_[29120]_ ,
    \new_[29121]_ , \new_[29125]_ , \new_[29126]_ , \new_[29130]_ ,
    \new_[29131]_ , \new_[29132]_ , \new_[29136]_ , \new_[29137]_ ,
    \new_[29141]_ , \new_[29142]_ , \new_[29143]_ , \new_[29147]_ ,
    \new_[29148]_ , \new_[29152]_ , \new_[29153]_ , \new_[29154]_ ,
    \new_[29158]_ , \new_[29159]_ , \new_[29163]_ , \new_[29164]_ ,
    \new_[29165]_ , \new_[29169]_ , \new_[29170]_ , \new_[29174]_ ,
    \new_[29175]_ , \new_[29176]_ , \new_[29180]_ , \new_[29181]_ ,
    \new_[29185]_ , \new_[29186]_ , \new_[29187]_ , \new_[29191]_ ,
    \new_[29192]_ , \new_[29196]_ , \new_[29197]_ , \new_[29198]_ ,
    \new_[29202]_ , \new_[29203]_ , \new_[29207]_ , \new_[29208]_ ,
    \new_[29209]_ , \new_[29213]_ , \new_[29214]_ , \new_[29218]_ ,
    \new_[29219]_ , \new_[29220]_ , \new_[29224]_ , \new_[29225]_ ,
    \new_[29229]_ , \new_[29230]_ , \new_[29231]_ , \new_[29235]_ ,
    \new_[29236]_ , \new_[29240]_ , \new_[29241]_ , \new_[29242]_ ,
    \new_[29246]_ , \new_[29247]_ , \new_[29251]_ , \new_[29252]_ ,
    \new_[29253]_ , \new_[29257]_ , \new_[29258]_ , \new_[29262]_ ,
    \new_[29263]_ , \new_[29264]_ , \new_[29268]_ , \new_[29269]_ ,
    \new_[29273]_ , \new_[29274]_ , \new_[29275]_ , \new_[29279]_ ,
    \new_[29280]_ , \new_[29284]_ , \new_[29285]_ , \new_[29286]_ ,
    \new_[29290]_ , \new_[29291]_ , \new_[29295]_ , \new_[29296]_ ,
    \new_[29297]_ , \new_[29301]_ , \new_[29302]_ , \new_[29306]_ ,
    \new_[29307]_ , \new_[29308]_ , \new_[29312]_ , \new_[29313]_ ,
    \new_[29317]_ , \new_[29318]_ , \new_[29319]_ , \new_[29323]_ ,
    \new_[29324]_ , \new_[29328]_ , \new_[29329]_ , \new_[29330]_ ,
    \new_[29334]_ , \new_[29335]_ , \new_[29339]_ , \new_[29340]_ ,
    \new_[29341]_ , \new_[29345]_ , \new_[29346]_ , \new_[29350]_ ,
    \new_[29351]_ , \new_[29352]_ , \new_[29356]_ , \new_[29357]_ ,
    \new_[29361]_ , \new_[29362]_ , \new_[29363]_ , \new_[29367]_ ,
    \new_[29368]_ , \new_[29372]_ , \new_[29373]_ , \new_[29374]_ ,
    \new_[29378]_ , \new_[29379]_ , \new_[29383]_ , \new_[29384]_ ,
    \new_[29385]_ , \new_[29389]_ , \new_[29390]_ , \new_[29394]_ ,
    \new_[29395]_ , \new_[29396]_ , \new_[29400]_ , \new_[29401]_ ,
    \new_[29405]_ , \new_[29406]_ , \new_[29407]_ , \new_[29411]_ ,
    \new_[29412]_ , \new_[29416]_ , \new_[29417]_ , \new_[29418]_ ,
    \new_[29422]_ , \new_[29423]_ , \new_[29427]_ , \new_[29428]_ ,
    \new_[29429]_ , \new_[29433]_ , \new_[29434]_ , \new_[29438]_ ,
    \new_[29439]_ , \new_[29440]_ , \new_[29444]_ , \new_[29445]_ ,
    \new_[29449]_ , \new_[29450]_ , \new_[29451]_ , \new_[29455]_ ,
    \new_[29456]_ , \new_[29460]_ , \new_[29461]_ , \new_[29462]_ ,
    \new_[29466]_ , \new_[29467]_ , \new_[29471]_ , \new_[29472]_ ,
    \new_[29473]_ , \new_[29477]_ , \new_[29478]_ , \new_[29482]_ ,
    \new_[29483]_ , \new_[29484]_ , \new_[29488]_ , \new_[29489]_ ,
    \new_[29493]_ , \new_[29494]_ , \new_[29495]_ , \new_[29499]_ ,
    \new_[29500]_ , \new_[29503]_ , \new_[29506]_ , \new_[29507]_ ,
    \new_[29508]_ , \new_[29512]_ , \new_[29513]_ , \new_[29517]_ ,
    \new_[29518]_ , \new_[29519]_ , \new_[29523]_ , \new_[29524]_ ,
    \new_[29527]_ , \new_[29530]_ , \new_[29531]_ , \new_[29532]_ ,
    \new_[29536]_ , \new_[29537]_ , \new_[29541]_ , \new_[29542]_ ,
    \new_[29543]_ , \new_[29547]_ , \new_[29548]_ , \new_[29551]_ ,
    \new_[29554]_ , \new_[29555]_ , \new_[29556]_ , \new_[29560]_ ,
    \new_[29561]_ , \new_[29565]_ , \new_[29566]_ , \new_[29567]_ ,
    \new_[29571]_ , \new_[29572]_ , \new_[29575]_ , \new_[29578]_ ,
    \new_[29579]_ , \new_[29580]_ , \new_[29584]_ , \new_[29585]_ ,
    \new_[29589]_ , \new_[29590]_ , \new_[29591]_ , \new_[29595]_ ,
    \new_[29596]_ , \new_[29599]_ , \new_[29602]_ , \new_[29603]_ ,
    \new_[29604]_ , \new_[29608]_ , \new_[29609]_ , \new_[29613]_ ,
    \new_[29614]_ , \new_[29615]_ , \new_[29619]_ , \new_[29620]_ ,
    \new_[29623]_ , \new_[29626]_ , \new_[29627]_ , \new_[29628]_ ,
    \new_[29632]_ , \new_[29633]_ , \new_[29637]_ , \new_[29638]_ ,
    \new_[29639]_ , \new_[29643]_ , \new_[29644]_ , \new_[29647]_ ,
    \new_[29650]_ , \new_[29651]_ , \new_[29652]_ , \new_[29656]_ ,
    \new_[29657]_ , \new_[29661]_ , \new_[29662]_ , \new_[29663]_ ,
    \new_[29667]_ , \new_[29668]_ , \new_[29671]_ , \new_[29674]_ ,
    \new_[29675]_ , \new_[29676]_ , \new_[29680]_ , \new_[29681]_ ,
    \new_[29685]_ , \new_[29686]_ , \new_[29687]_ , \new_[29691]_ ,
    \new_[29692]_ , \new_[29695]_ , \new_[29698]_ , \new_[29699]_ ,
    \new_[29700]_ , \new_[29704]_ , \new_[29705]_ , \new_[29709]_ ,
    \new_[29710]_ , \new_[29711]_ , \new_[29715]_ , \new_[29716]_ ,
    \new_[29719]_ , \new_[29722]_ , \new_[29723]_ , \new_[29724]_ ,
    \new_[29728]_ , \new_[29729]_ , \new_[29733]_ , \new_[29734]_ ,
    \new_[29735]_ , \new_[29739]_ , \new_[29740]_ , \new_[29743]_ ,
    \new_[29746]_ , \new_[29747]_ , \new_[29748]_ , \new_[29752]_ ,
    \new_[29753]_ , \new_[29757]_ , \new_[29758]_ , \new_[29759]_ ,
    \new_[29763]_ , \new_[29764]_ , \new_[29767]_ , \new_[29770]_ ,
    \new_[29771]_ , \new_[29772]_ , \new_[29776]_ , \new_[29777]_ ,
    \new_[29781]_ , \new_[29782]_ , \new_[29783]_ , \new_[29787]_ ,
    \new_[29788]_ , \new_[29791]_ , \new_[29794]_ , \new_[29795]_ ,
    \new_[29796]_ , \new_[29800]_ , \new_[29801]_ , \new_[29805]_ ,
    \new_[29806]_ , \new_[29807]_ , \new_[29811]_ , \new_[29812]_ ,
    \new_[29815]_ , \new_[29818]_ , \new_[29819]_ , \new_[29820]_ ,
    \new_[29824]_ , \new_[29825]_ , \new_[29829]_ , \new_[29830]_ ,
    \new_[29831]_ , \new_[29835]_ , \new_[29836]_ , \new_[29839]_ ,
    \new_[29842]_ , \new_[29843]_ , \new_[29844]_ , \new_[29848]_ ,
    \new_[29849]_ , \new_[29853]_ , \new_[29854]_ , \new_[29855]_ ,
    \new_[29859]_ , \new_[29860]_ , \new_[29863]_ , \new_[29866]_ ,
    \new_[29867]_ , \new_[29868]_ , \new_[29872]_ , \new_[29873]_ ,
    \new_[29877]_ , \new_[29878]_ , \new_[29879]_ , \new_[29883]_ ,
    \new_[29884]_ , \new_[29887]_ , \new_[29890]_ , \new_[29891]_ ,
    \new_[29892]_ , \new_[29896]_ , \new_[29897]_ , \new_[29901]_ ,
    \new_[29902]_ , \new_[29903]_ , \new_[29907]_ , \new_[29908]_ ,
    \new_[29911]_ , \new_[29914]_ , \new_[29915]_ , \new_[29916]_ ,
    \new_[29920]_ , \new_[29921]_ , \new_[29925]_ , \new_[29926]_ ,
    \new_[29927]_ , \new_[29931]_ , \new_[29932]_ , \new_[29935]_ ,
    \new_[29938]_ , \new_[29939]_ , \new_[29940]_ , \new_[29944]_ ,
    \new_[29945]_ , \new_[29949]_ , \new_[29950]_ , \new_[29951]_ ,
    \new_[29955]_ , \new_[29956]_ , \new_[29959]_ , \new_[29962]_ ,
    \new_[29963]_ , \new_[29964]_ , \new_[29968]_ , \new_[29969]_ ,
    \new_[29973]_ , \new_[29974]_ , \new_[29975]_ , \new_[29979]_ ,
    \new_[29980]_ , \new_[29983]_ , \new_[29986]_ , \new_[29987]_ ,
    \new_[29988]_ , \new_[29992]_ , \new_[29993]_ , \new_[29997]_ ,
    \new_[29998]_ , \new_[29999]_ , \new_[30003]_ , \new_[30004]_ ,
    \new_[30007]_ , \new_[30010]_ , \new_[30011]_ , \new_[30012]_ ,
    \new_[30016]_ , \new_[30017]_ , \new_[30021]_ , \new_[30022]_ ,
    \new_[30023]_ , \new_[30027]_ , \new_[30028]_ , \new_[30031]_ ,
    \new_[30034]_ , \new_[30035]_ , \new_[30036]_ , \new_[30040]_ ,
    \new_[30041]_ , \new_[30045]_ , \new_[30046]_ , \new_[30047]_ ,
    \new_[30051]_ , \new_[30052]_ , \new_[30055]_ , \new_[30058]_ ,
    \new_[30059]_ , \new_[30060]_ , \new_[30064]_ , \new_[30065]_ ,
    \new_[30069]_ , \new_[30070]_ , \new_[30071]_ , \new_[30075]_ ,
    \new_[30076]_ , \new_[30079]_ , \new_[30082]_ , \new_[30083]_ ,
    \new_[30084]_ , \new_[30088]_ , \new_[30089]_ , \new_[30093]_ ,
    \new_[30094]_ , \new_[30095]_ , \new_[30099]_ , \new_[30100]_ ,
    \new_[30103]_ , \new_[30106]_ , \new_[30107]_ , \new_[30108]_ ,
    \new_[30112]_ , \new_[30113]_ , \new_[30117]_ , \new_[30118]_ ,
    \new_[30119]_ , \new_[30123]_ , \new_[30124]_ , \new_[30127]_ ,
    \new_[30130]_ , \new_[30131]_ , \new_[30132]_ , \new_[30136]_ ,
    \new_[30137]_ , \new_[30141]_ , \new_[30142]_ , \new_[30143]_ ,
    \new_[30147]_ , \new_[30148]_ , \new_[30151]_ , \new_[30154]_ ,
    \new_[30155]_ , \new_[30156]_ , \new_[30160]_ , \new_[30161]_ ,
    \new_[30165]_ , \new_[30166]_ , \new_[30167]_ , \new_[30171]_ ,
    \new_[30172]_ , \new_[30175]_ , \new_[30178]_ , \new_[30179]_ ,
    \new_[30180]_ , \new_[30184]_ , \new_[30185]_ , \new_[30189]_ ,
    \new_[30190]_ , \new_[30191]_ , \new_[30195]_ , \new_[30196]_ ,
    \new_[30199]_ , \new_[30202]_ , \new_[30203]_ , \new_[30204]_ ,
    \new_[30208]_ , \new_[30209]_ , \new_[30213]_ , \new_[30214]_ ,
    \new_[30215]_ , \new_[30219]_ , \new_[30220]_ , \new_[30223]_ ,
    \new_[30226]_ , \new_[30227]_ , \new_[30228]_ , \new_[30232]_ ,
    \new_[30233]_ , \new_[30237]_ , \new_[30238]_ , \new_[30239]_ ,
    \new_[30243]_ , \new_[30244]_ , \new_[30247]_ , \new_[30250]_ ,
    \new_[30251]_ , \new_[30252]_ , \new_[30256]_ , \new_[30257]_ ,
    \new_[30261]_ , \new_[30262]_ , \new_[30263]_ , \new_[30267]_ ,
    \new_[30268]_ , \new_[30271]_ , \new_[30274]_ , \new_[30275]_ ,
    \new_[30276]_ , \new_[30280]_ , \new_[30281]_ , \new_[30285]_ ,
    \new_[30286]_ , \new_[30287]_ , \new_[30291]_ , \new_[30292]_ ,
    \new_[30295]_ , \new_[30298]_ , \new_[30299]_ , \new_[30300]_ ,
    \new_[30304]_ , \new_[30305]_ , \new_[30309]_ , \new_[30310]_ ,
    \new_[30311]_ , \new_[30315]_ , \new_[30316]_ , \new_[30319]_ ,
    \new_[30322]_ , \new_[30323]_ , \new_[30324]_ , \new_[30328]_ ,
    \new_[30329]_ , \new_[30333]_ , \new_[30334]_ , \new_[30335]_ ,
    \new_[30339]_ , \new_[30340]_ , \new_[30343]_ , \new_[30346]_ ,
    \new_[30347]_ , \new_[30348]_ , \new_[30352]_ , \new_[30353]_ ,
    \new_[30357]_ , \new_[30358]_ , \new_[30359]_ , \new_[30363]_ ,
    \new_[30364]_ , \new_[30367]_ , \new_[30370]_ , \new_[30371]_ ,
    \new_[30372]_ , \new_[30376]_ , \new_[30377]_ , \new_[30381]_ ,
    \new_[30382]_ , \new_[30383]_ , \new_[30387]_ , \new_[30388]_ ,
    \new_[30391]_ , \new_[30394]_ , \new_[30395]_ , \new_[30396]_ ,
    \new_[30400]_ , \new_[30401]_ , \new_[30405]_ , \new_[30406]_ ,
    \new_[30407]_ , \new_[30411]_ , \new_[30412]_ , \new_[30415]_ ,
    \new_[30418]_ , \new_[30419]_ , \new_[30420]_ , \new_[30424]_ ,
    \new_[30425]_ , \new_[30429]_ , \new_[30430]_ , \new_[30431]_ ,
    \new_[30435]_ , \new_[30436]_ , \new_[30439]_ , \new_[30442]_ ,
    \new_[30443]_ , \new_[30444]_ , \new_[30448]_ , \new_[30449]_ ,
    \new_[30453]_ , \new_[30454]_ , \new_[30455]_ , \new_[30459]_ ,
    \new_[30460]_ , \new_[30463]_ , \new_[30466]_ , \new_[30467]_ ,
    \new_[30468]_ , \new_[30472]_ , \new_[30473]_ , \new_[30477]_ ,
    \new_[30478]_ , \new_[30479]_ , \new_[30483]_ , \new_[30484]_ ,
    \new_[30487]_ , \new_[30490]_ , \new_[30491]_ , \new_[30492]_ ,
    \new_[30496]_ , \new_[30497]_ , \new_[30501]_ , \new_[30502]_ ,
    \new_[30503]_ , \new_[30507]_ , \new_[30508]_ , \new_[30511]_ ,
    \new_[30514]_ , \new_[30515]_ , \new_[30516]_ , \new_[30520]_ ,
    \new_[30521]_ , \new_[30525]_ , \new_[30526]_ , \new_[30527]_ ,
    \new_[30531]_ , \new_[30532]_ , \new_[30535]_ , \new_[30538]_ ,
    \new_[30539]_ , \new_[30540]_ , \new_[30544]_ , \new_[30545]_ ,
    \new_[30549]_ , \new_[30550]_ , \new_[30551]_ , \new_[30555]_ ,
    \new_[30556]_ , \new_[30559]_ , \new_[30562]_ , \new_[30563]_ ,
    \new_[30564]_ , \new_[30568]_ , \new_[30569]_ , \new_[30573]_ ,
    \new_[30574]_ , \new_[30575]_ , \new_[30579]_ , \new_[30580]_ ,
    \new_[30583]_ , \new_[30586]_ , \new_[30587]_ , \new_[30588]_ ,
    \new_[30592]_ , \new_[30593]_ , \new_[30597]_ , \new_[30598]_ ,
    \new_[30599]_ , \new_[30603]_ , \new_[30604]_ , \new_[30607]_ ,
    \new_[30610]_ , \new_[30611]_ , \new_[30612]_ , \new_[30616]_ ,
    \new_[30617]_ , \new_[30621]_ , \new_[30622]_ , \new_[30623]_ ,
    \new_[30627]_ , \new_[30628]_ , \new_[30631]_ , \new_[30634]_ ,
    \new_[30635]_ , \new_[30636]_ , \new_[30640]_ , \new_[30641]_ ,
    \new_[30645]_ , \new_[30646]_ , \new_[30647]_ , \new_[30651]_ ,
    \new_[30652]_ , \new_[30655]_ , \new_[30658]_ , \new_[30659]_ ,
    \new_[30660]_ , \new_[30664]_ , \new_[30665]_ , \new_[30669]_ ,
    \new_[30670]_ , \new_[30671]_ , \new_[30675]_ , \new_[30676]_ ,
    \new_[30679]_ , \new_[30682]_ , \new_[30683]_ , \new_[30684]_ ,
    \new_[30688]_ , \new_[30689]_ , \new_[30693]_ , \new_[30694]_ ,
    \new_[30695]_ , \new_[30699]_ , \new_[30700]_ , \new_[30703]_ ,
    \new_[30706]_ , \new_[30707]_ , \new_[30708]_ , \new_[30712]_ ,
    \new_[30713]_ , \new_[30717]_ , \new_[30718]_ , \new_[30719]_ ,
    \new_[30723]_ , \new_[30724]_ , \new_[30727]_ , \new_[30730]_ ,
    \new_[30731]_ , \new_[30732]_ , \new_[30736]_ , \new_[30737]_ ,
    \new_[30741]_ , \new_[30742]_ , \new_[30743]_ , \new_[30747]_ ,
    \new_[30748]_ , \new_[30751]_ , \new_[30754]_ , \new_[30755]_ ,
    \new_[30756]_ , \new_[30760]_ , \new_[30761]_ , \new_[30765]_ ,
    \new_[30766]_ , \new_[30767]_ , \new_[30771]_ , \new_[30772]_ ,
    \new_[30775]_ , \new_[30778]_ , \new_[30779]_ , \new_[30780]_ ,
    \new_[30784]_ , \new_[30785]_ , \new_[30789]_ , \new_[30790]_ ,
    \new_[30791]_ , \new_[30795]_ , \new_[30796]_ , \new_[30799]_ ,
    \new_[30802]_ , \new_[30803]_ , \new_[30804]_ , \new_[30808]_ ,
    \new_[30809]_ , \new_[30813]_ , \new_[30814]_ , \new_[30815]_ ,
    \new_[30819]_ , \new_[30820]_ , \new_[30823]_ , \new_[30826]_ ,
    \new_[30827]_ , \new_[30828]_ , \new_[30832]_ , \new_[30833]_ ,
    \new_[30837]_ , \new_[30838]_ , \new_[30839]_ , \new_[30843]_ ,
    \new_[30844]_ , \new_[30847]_ , \new_[30850]_ , \new_[30851]_ ,
    \new_[30852]_ , \new_[30856]_ , \new_[30857]_ , \new_[30861]_ ,
    \new_[30862]_ , \new_[30863]_ , \new_[30867]_ , \new_[30868]_ ,
    \new_[30871]_ , \new_[30874]_ , \new_[30875]_ , \new_[30876]_ ,
    \new_[30880]_ , \new_[30881]_ , \new_[30885]_ , \new_[30886]_ ,
    \new_[30887]_ , \new_[30891]_ , \new_[30892]_ , \new_[30895]_ ,
    \new_[30898]_ , \new_[30899]_ , \new_[30900]_ , \new_[30904]_ ,
    \new_[30905]_ , \new_[30909]_ , \new_[30910]_ , \new_[30911]_ ,
    \new_[30915]_ , \new_[30916]_ , \new_[30919]_ , \new_[30922]_ ,
    \new_[30923]_ , \new_[30924]_ , \new_[30928]_ , \new_[30929]_ ,
    \new_[30933]_ , \new_[30934]_ , \new_[30935]_ , \new_[30939]_ ,
    \new_[30940]_ , \new_[30943]_ , \new_[30946]_ , \new_[30947]_ ,
    \new_[30948]_ , \new_[30952]_ , \new_[30953]_ , \new_[30957]_ ,
    \new_[30958]_ , \new_[30959]_ , \new_[30963]_ , \new_[30964]_ ,
    \new_[30967]_ , \new_[30970]_ , \new_[30971]_ , \new_[30972]_ ,
    \new_[30976]_ , \new_[30977]_ , \new_[30981]_ , \new_[30982]_ ,
    \new_[30983]_ , \new_[30987]_ , \new_[30988]_ , \new_[30991]_ ,
    \new_[30994]_ , \new_[30995]_ , \new_[30996]_ , \new_[31000]_ ,
    \new_[31001]_ , \new_[31005]_ , \new_[31006]_ , \new_[31007]_ ,
    \new_[31011]_ , \new_[31012]_ , \new_[31015]_ , \new_[31018]_ ,
    \new_[31019]_ , \new_[31020]_ , \new_[31024]_ , \new_[31025]_ ,
    \new_[31029]_ , \new_[31030]_ , \new_[31031]_ , \new_[31035]_ ,
    \new_[31036]_ , \new_[31039]_ , \new_[31042]_ , \new_[31043]_ ,
    \new_[31044]_ , \new_[31048]_ , \new_[31049]_ , \new_[31053]_ ,
    \new_[31054]_ , \new_[31055]_ , \new_[31059]_ , \new_[31060]_ ,
    \new_[31063]_ , \new_[31066]_ , \new_[31067]_ , \new_[31068]_ ,
    \new_[31072]_ , \new_[31073]_ , \new_[31077]_ , \new_[31078]_ ,
    \new_[31079]_ , \new_[31083]_ , \new_[31084]_ , \new_[31087]_ ,
    \new_[31090]_ , \new_[31091]_ , \new_[31092]_ , \new_[31096]_ ,
    \new_[31097]_ , \new_[31101]_ , \new_[31102]_ , \new_[31103]_ ,
    \new_[31107]_ , \new_[31108]_ , \new_[31111]_ , \new_[31114]_ ,
    \new_[31115]_ , \new_[31116]_ , \new_[31120]_ , \new_[31121]_ ,
    \new_[31125]_ , \new_[31126]_ , \new_[31127]_ , \new_[31131]_ ,
    \new_[31132]_ , \new_[31135]_ , \new_[31138]_ , \new_[31139]_ ,
    \new_[31140]_ , \new_[31144]_ , \new_[31145]_ , \new_[31149]_ ,
    \new_[31150]_ , \new_[31151]_ , \new_[31155]_ , \new_[31156]_ ,
    \new_[31159]_ , \new_[31162]_ , \new_[31163]_ , \new_[31164]_ ,
    \new_[31168]_ , \new_[31169]_ , \new_[31173]_ , \new_[31174]_ ,
    \new_[31175]_ , \new_[31179]_ , \new_[31180]_ , \new_[31183]_ ,
    \new_[31186]_ , \new_[31187]_ , \new_[31188]_ , \new_[31192]_ ,
    \new_[31193]_ , \new_[31197]_ , \new_[31198]_ , \new_[31199]_ ,
    \new_[31203]_ , \new_[31204]_ , \new_[31207]_ , \new_[31210]_ ,
    \new_[31211]_ , \new_[31212]_ , \new_[31216]_ , \new_[31217]_ ,
    \new_[31221]_ , \new_[31222]_ , \new_[31223]_ , \new_[31227]_ ,
    \new_[31228]_ , \new_[31231]_ , \new_[31234]_ , \new_[31235]_ ,
    \new_[31236]_ , \new_[31240]_ , \new_[31241]_ , \new_[31245]_ ,
    \new_[31246]_ , \new_[31247]_ , \new_[31251]_ , \new_[31252]_ ,
    \new_[31255]_ , \new_[31258]_ , \new_[31259]_ , \new_[31260]_ ,
    \new_[31264]_ , \new_[31265]_ , \new_[31269]_ , \new_[31270]_ ,
    \new_[31271]_ , \new_[31275]_ , \new_[31276]_ , \new_[31279]_ ,
    \new_[31282]_ , \new_[31283]_ , \new_[31284]_ , \new_[31288]_ ,
    \new_[31289]_ , \new_[31293]_ , \new_[31294]_ , \new_[31295]_ ,
    \new_[31299]_ , \new_[31300]_ , \new_[31303]_ , \new_[31306]_ ,
    \new_[31307]_ , \new_[31308]_ , \new_[31312]_ , \new_[31313]_ ,
    \new_[31317]_ , \new_[31318]_ , \new_[31319]_ , \new_[31323]_ ,
    \new_[31324]_ , \new_[31327]_ , \new_[31330]_ , \new_[31331]_ ,
    \new_[31332]_ , \new_[31336]_ , \new_[31337]_ , \new_[31341]_ ,
    \new_[31342]_ , \new_[31343]_ , \new_[31347]_ , \new_[31348]_ ,
    \new_[31351]_ , \new_[31354]_ , \new_[31355]_ , \new_[31356]_ ,
    \new_[31360]_ , \new_[31361]_ , \new_[31365]_ , \new_[31366]_ ,
    \new_[31367]_ , \new_[31371]_ , \new_[31372]_ , \new_[31375]_ ,
    \new_[31378]_ , \new_[31379]_ , \new_[31380]_ , \new_[31384]_ ,
    \new_[31385]_ , \new_[31389]_ , \new_[31390]_ , \new_[31391]_ ,
    \new_[31395]_ , \new_[31396]_ , \new_[31399]_ , \new_[31402]_ ,
    \new_[31403]_ , \new_[31404]_ , \new_[31408]_ , \new_[31409]_ ,
    \new_[31413]_ , \new_[31414]_ , \new_[31415]_ , \new_[31419]_ ,
    \new_[31420]_ , \new_[31423]_ , \new_[31426]_ , \new_[31427]_ ,
    \new_[31428]_ , \new_[31432]_ , \new_[31433]_ , \new_[31437]_ ,
    \new_[31438]_ , \new_[31439]_ , \new_[31443]_ , \new_[31444]_ ,
    \new_[31447]_ , \new_[31450]_ , \new_[31451]_ , \new_[31452]_ ,
    \new_[31456]_ , \new_[31457]_ , \new_[31461]_ , \new_[31462]_ ,
    \new_[31463]_ , \new_[31467]_ , \new_[31468]_ , \new_[31471]_ ,
    \new_[31474]_ , \new_[31475]_ , \new_[31476]_ , \new_[31480]_ ,
    \new_[31481]_ , \new_[31485]_ , \new_[31486]_ , \new_[31487]_ ,
    \new_[31491]_ , \new_[31492]_ , \new_[31495]_ , \new_[31498]_ ,
    \new_[31499]_ , \new_[31500]_ , \new_[31504]_ , \new_[31505]_ ,
    \new_[31509]_ , \new_[31510]_ , \new_[31511]_ , \new_[31515]_ ,
    \new_[31516]_ , \new_[31519]_ , \new_[31522]_ , \new_[31523]_ ,
    \new_[31524]_ , \new_[31528]_ , \new_[31529]_ , \new_[31533]_ ,
    \new_[31534]_ , \new_[31535]_ , \new_[31539]_ , \new_[31540]_ ,
    \new_[31543]_ , \new_[31546]_ , \new_[31547]_ , \new_[31548]_ ,
    \new_[31552]_ , \new_[31553]_ , \new_[31557]_ , \new_[31558]_ ,
    \new_[31559]_ , \new_[31563]_ , \new_[31564]_ , \new_[31567]_ ,
    \new_[31570]_ , \new_[31571]_ , \new_[31572]_ , \new_[31576]_ ,
    \new_[31577]_ , \new_[31581]_ , \new_[31582]_ , \new_[31583]_ ,
    \new_[31587]_ , \new_[31588]_ , \new_[31591]_ , \new_[31594]_ ,
    \new_[31595]_ , \new_[31596]_ , \new_[31600]_ , \new_[31601]_ ,
    \new_[31605]_ , \new_[31606]_ , \new_[31607]_ , \new_[31611]_ ,
    \new_[31612]_ , \new_[31615]_ , \new_[31618]_ , \new_[31619]_ ,
    \new_[31620]_ , \new_[31624]_ , \new_[31625]_ , \new_[31629]_ ,
    \new_[31630]_ , \new_[31631]_ , \new_[31635]_ , \new_[31636]_ ,
    \new_[31639]_ , \new_[31642]_ , \new_[31643]_ , \new_[31644]_ ,
    \new_[31648]_ , \new_[31649]_ , \new_[31653]_ , \new_[31654]_ ,
    \new_[31655]_ , \new_[31659]_ , \new_[31660]_ , \new_[31663]_ ,
    \new_[31666]_ , \new_[31667]_ , \new_[31668]_ , \new_[31672]_ ,
    \new_[31673]_ , \new_[31677]_ , \new_[31678]_ , \new_[31679]_ ,
    \new_[31683]_ , \new_[31684]_ , \new_[31687]_ , \new_[31690]_ ,
    \new_[31691]_ , \new_[31692]_ , \new_[31696]_ , \new_[31697]_ ,
    \new_[31701]_ , \new_[31702]_ , \new_[31703]_ , \new_[31707]_ ,
    \new_[31708]_ , \new_[31711]_ , \new_[31714]_ , \new_[31715]_ ,
    \new_[31716]_ , \new_[31720]_ , \new_[31721]_ , \new_[31725]_ ,
    \new_[31726]_ , \new_[31727]_ , \new_[31731]_ , \new_[31732]_ ,
    \new_[31735]_ , \new_[31738]_ , \new_[31739]_ , \new_[31740]_ ,
    \new_[31744]_ , \new_[31745]_ , \new_[31749]_ , \new_[31750]_ ,
    \new_[31751]_ , \new_[31755]_ , \new_[31756]_ , \new_[31759]_ ,
    \new_[31762]_ , \new_[31763]_ , \new_[31764]_ , \new_[31768]_ ,
    \new_[31769]_ , \new_[31773]_ , \new_[31774]_ , \new_[31775]_ ,
    \new_[31779]_ , \new_[31780]_ , \new_[31783]_ , \new_[31786]_ ,
    \new_[31787]_ , \new_[31788]_ , \new_[31792]_ , \new_[31793]_ ,
    \new_[31797]_ , \new_[31798]_ , \new_[31799]_ , \new_[31803]_ ,
    \new_[31804]_ , \new_[31807]_ , \new_[31810]_ , \new_[31811]_ ,
    \new_[31812]_ , \new_[31816]_ , \new_[31817]_ , \new_[31821]_ ,
    \new_[31822]_ , \new_[31823]_ , \new_[31827]_ , \new_[31828]_ ,
    \new_[31831]_ , \new_[31834]_ , \new_[31835]_ , \new_[31836]_ ,
    \new_[31840]_ , \new_[31841]_ , \new_[31845]_ , \new_[31846]_ ,
    \new_[31847]_ , \new_[31851]_ , \new_[31852]_ , \new_[31855]_ ,
    \new_[31858]_ , \new_[31859]_ , \new_[31860]_ , \new_[31864]_ ,
    \new_[31865]_ , \new_[31869]_ , \new_[31870]_ , \new_[31871]_ ,
    \new_[31875]_ , \new_[31876]_ , \new_[31879]_ , \new_[31882]_ ,
    \new_[31883]_ , \new_[31884]_ , \new_[31888]_ , \new_[31889]_ ,
    \new_[31893]_ , \new_[31894]_ , \new_[31895]_ , \new_[31899]_ ,
    \new_[31900]_ , \new_[31903]_ , \new_[31906]_ , \new_[31907]_ ,
    \new_[31908]_ , \new_[31912]_ , \new_[31913]_ , \new_[31917]_ ,
    \new_[31918]_ , \new_[31919]_ , \new_[31923]_ , \new_[31924]_ ,
    \new_[31927]_ , \new_[31930]_ , \new_[31931]_ , \new_[31932]_ ,
    \new_[31936]_ , \new_[31937]_ , \new_[31941]_ , \new_[31942]_ ,
    \new_[31943]_ , \new_[31947]_ , \new_[31948]_ , \new_[31951]_ ,
    \new_[31954]_ , \new_[31955]_ , \new_[31956]_ , \new_[31960]_ ,
    \new_[31961]_ , \new_[31965]_ , \new_[31966]_ , \new_[31967]_ ,
    \new_[31971]_ , \new_[31972]_ , \new_[31975]_ , \new_[31978]_ ,
    \new_[31979]_ , \new_[31980]_ , \new_[31984]_ , \new_[31985]_ ,
    \new_[31989]_ , \new_[31990]_ , \new_[31991]_ , \new_[31995]_ ,
    \new_[31996]_ , \new_[31999]_ , \new_[32002]_ , \new_[32003]_ ,
    \new_[32004]_ , \new_[32008]_ , \new_[32009]_ , \new_[32013]_ ,
    \new_[32014]_ , \new_[32015]_ , \new_[32019]_ , \new_[32020]_ ,
    \new_[32023]_ , \new_[32026]_ , \new_[32027]_ , \new_[32028]_ ,
    \new_[32032]_ , \new_[32033]_ , \new_[32037]_ , \new_[32038]_ ,
    \new_[32039]_ , \new_[32043]_ , \new_[32044]_ , \new_[32047]_ ,
    \new_[32050]_ , \new_[32051]_ , \new_[32052]_ , \new_[32056]_ ,
    \new_[32057]_ , \new_[32061]_ , \new_[32062]_ , \new_[32063]_ ,
    \new_[32067]_ , \new_[32068]_ , \new_[32071]_ , \new_[32074]_ ,
    \new_[32075]_ , \new_[32076]_ , \new_[32080]_ , \new_[32081]_ ,
    \new_[32085]_ , \new_[32086]_ , \new_[32087]_ , \new_[32091]_ ,
    \new_[32092]_ , \new_[32095]_ , \new_[32098]_ , \new_[32099]_ ,
    \new_[32100]_ , \new_[32104]_ , \new_[32105]_ , \new_[32109]_ ,
    \new_[32110]_ , \new_[32111]_ , \new_[32115]_ , \new_[32116]_ ,
    \new_[32119]_ , \new_[32122]_ , \new_[32123]_ , \new_[32124]_ ,
    \new_[32128]_ , \new_[32129]_ , \new_[32133]_ , \new_[32134]_ ,
    \new_[32135]_ , \new_[32139]_ , \new_[32140]_ , \new_[32143]_ ,
    \new_[32146]_ , \new_[32147]_ , \new_[32148]_ , \new_[32152]_ ,
    \new_[32153]_ , \new_[32157]_ , \new_[32158]_ , \new_[32159]_ ,
    \new_[32163]_ , \new_[32164]_ , \new_[32167]_ , \new_[32170]_ ,
    \new_[32171]_ , \new_[32172]_ , \new_[32176]_ , \new_[32177]_ ,
    \new_[32181]_ , \new_[32182]_ , \new_[32183]_ , \new_[32187]_ ,
    \new_[32188]_ , \new_[32191]_ , \new_[32194]_ , \new_[32195]_ ,
    \new_[32196]_ , \new_[32200]_ , \new_[32201]_ , \new_[32205]_ ,
    \new_[32206]_ , \new_[32207]_ , \new_[32211]_ , \new_[32212]_ ,
    \new_[32215]_ , \new_[32218]_ , \new_[32219]_ , \new_[32220]_ ,
    \new_[32224]_ , \new_[32225]_ , \new_[32229]_ , \new_[32230]_ ,
    \new_[32231]_ , \new_[32235]_ , \new_[32236]_ , \new_[32239]_ ,
    \new_[32242]_ , \new_[32243]_ , \new_[32244]_ , \new_[32248]_ ,
    \new_[32249]_ , \new_[32253]_ , \new_[32254]_ , \new_[32255]_ ,
    \new_[32259]_ , \new_[32260]_ , \new_[32263]_ , \new_[32266]_ ,
    \new_[32267]_ , \new_[32268]_ , \new_[32272]_ , \new_[32273]_ ,
    \new_[32277]_ , \new_[32278]_ , \new_[32279]_ , \new_[32283]_ ,
    \new_[32284]_ , \new_[32287]_ , \new_[32290]_ , \new_[32291]_ ,
    \new_[32292]_ , \new_[32296]_ , \new_[32297]_ , \new_[32301]_ ,
    \new_[32302]_ , \new_[32303]_ , \new_[32307]_ , \new_[32308]_ ,
    \new_[32311]_ , \new_[32314]_ , \new_[32315]_ , \new_[32316]_ ,
    \new_[32320]_ , \new_[32321]_ , \new_[32325]_ , \new_[32326]_ ,
    \new_[32327]_ , \new_[32331]_ , \new_[32332]_ , \new_[32335]_ ,
    \new_[32338]_ , \new_[32339]_ , \new_[32340]_ , \new_[32344]_ ,
    \new_[32345]_ , \new_[32349]_ , \new_[32350]_ , \new_[32351]_ ,
    \new_[32355]_ , \new_[32356]_ , \new_[32359]_ , \new_[32362]_ ,
    \new_[32363]_ , \new_[32364]_ , \new_[32368]_ , \new_[32369]_ ,
    \new_[32373]_ , \new_[32374]_ , \new_[32375]_ , \new_[32379]_ ,
    \new_[32380]_ , \new_[32383]_ , \new_[32386]_ , \new_[32387]_ ,
    \new_[32388]_ , \new_[32392]_ , \new_[32393]_ , \new_[32397]_ ,
    \new_[32398]_ , \new_[32399]_ , \new_[32403]_ , \new_[32404]_ ,
    \new_[32407]_ , \new_[32410]_ , \new_[32411]_ , \new_[32412]_ ,
    \new_[32416]_ , \new_[32417]_ , \new_[32421]_ , \new_[32422]_ ,
    \new_[32423]_ , \new_[32427]_ , \new_[32428]_ , \new_[32431]_ ,
    \new_[32434]_ , \new_[32435]_ , \new_[32436]_ , \new_[32440]_ ,
    \new_[32441]_ , \new_[32445]_ , \new_[32446]_ , \new_[32447]_ ,
    \new_[32451]_ , \new_[32452]_ , \new_[32455]_ , \new_[32458]_ ,
    \new_[32459]_ , \new_[32460]_ , \new_[32464]_ , \new_[32465]_ ,
    \new_[32469]_ , \new_[32470]_ , \new_[32471]_ , \new_[32475]_ ,
    \new_[32476]_ , \new_[32479]_ , \new_[32482]_ , \new_[32483]_ ,
    \new_[32484]_ , \new_[32488]_ , \new_[32489]_ , \new_[32493]_ ,
    \new_[32494]_ , \new_[32495]_ , \new_[32499]_ , \new_[32500]_ ,
    \new_[32503]_ , \new_[32506]_ , \new_[32507]_ , \new_[32508]_ ,
    \new_[32512]_ , \new_[32513]_ , \new_[32517]_ , \new_[32518]_ ,
    \new_[32519]_ , \new_[32523]_ , \new_[32524]_ , \new_[32527]_ ,
    \new_[32530]_ , \new_[32531]_ , \new_[32532]_ , \new_[32536]_ ,
    \new_[32537]_ , \new_[32541]_ , \new_[32542]_ , \new_[32543]_ ,
    \new_[32547]_ , \new_[32548]_ , \new_[32551]_ , \new_[32554]_ ,
    \new_[32555]_ , \new_[32556]_ , \new_[32560]_ , \new_[32561]_ ,
    \new_[32565]_ , \new_[32566]_ , \new_[32567]_ , \new_[32571]_ ,
    \new_[32572]_ , \new_[32575]_ , \new_[32578]_ , \new_[32579]_ ,
    \new_[32580]_ , \new_[32584]_ , \new_[32585]_ , \new_[32589]_ ,
    \new_[32590]_ , \new_[32591]_ , \new_[32595]_ , \new_[32596]_ ,
    \new_[32599]_ , \new_[32602]_ , \new_[32603]_ , \new_[32604]_ ,
    \new_[32608]_ , \new_[32609]_ , \new_[32613]_ , \new_[32614]_ ,
    \new_[32615]_ , \new_[32619]_ , \new_[32620]_ , \new_[32623]_ ,
    \new_[32626]_ , \new_[32627]_ , \new_[32628]_ , \new_[32632]_ ,
    \new_[32633]_ , \new_[32637]_ , \new_[32638]_ , \new_[32639]_ ,
    \new_[32643]_ , \new_[32644]_ , \new_[32647]_ , \new_[32650]_ ,
    \new_[32651]_ , \new_[32652]_ , \new_[32656]_ , \new_[32657]_ ,
    \new_[32661]_ , \new_[32662]_ , \new_[32663]_ , \new_[32667]_ ,
    \new_[32668]_ , \new_[32671]_ , \new_[32674]_ , \new_[32675]_ ,
    \new_[32676]_ , \new_[32680]_ , \new_[32681]_ , \new_[32685]_ ,
    \new_[32686]_ , \new_[32687]_ , \new_[32691]_ , \new_[32692]_ ,
    \new_[32695]_ , \new_[32698]_ , \new_[32699]_ , \new_[32700]_ ,
    \new_[32704]_ , \new_[32705]_ , \new_[32709]_ , \new_[32710]_ ,
    \new_[32711]_ , \new_[32715]_ , \new_[32716]_ , \new_[32719]_ ,
    \new_[32722]_ , \new_[32723]_ , \new_[32724]_ , \new_[32728]_ ,
    \new_[32729]_ , \new_[32733]_ , \new_[32734]_ , \new_[32735]_ ,
    \new_[32739]_ , \new_[32740]_ , \new_[32743]_ , \new_[32746]_ ,
    \new_[32747]_ , \new_[32748]_ , \new_[32752]_ , \new_[32753]_ ,
    \new_[32757]_ , \new_[32758]_ , \new_[32759]_ , \new_[32763]_ ,
    \new_[32764]_ , \new_[32767]_ , \new_[32770]_ , \new_[32771]_ ,
    \new_[32772]_ , \new_[32776]_ , \new_[32777]_ , \new_[32781]_ ,
    \new_[32782]_ , \new_[32783]_ , \new_[32787]_ , \new_[32788]_ ,
    \new_[32791]_ , \new_[32794]_ , \new_[32795]_ , \new_[32796]_ ,
    \new_[32800]_ , \new_[32801]_ , \new_[32805]_ , \new_[32806]_ ,
    \new_[32807]_ , \new_[32811]_ , \new_[32812]_ , \new_[32815]_ ,
    \new_[32818]_ , \new_[32819]_ , \new_[32820]_ , \new_[32824]_ ,
    \new_[32825]_ , \new_[32829]_ , \new_[32830]_ , \new_[32831]_ ,
    \new_[32835]_ , \new_[32836]_ , \new_[32839]_ , \new_[32842]_ ,
    \new_[32843]_ , \new_[32844]_ , \new_[32848]_ , \new_[32849]_ ,
    \new_[32853]_ , \new_[32854]_ , \new_[32855]_ , \new_[32859]_ ,
    \new_[32860]_ , \new_[32863]_ , \new_[32866]_ , \new_[32867]_ ,
    \new_[32868]_ , \new_[32872]_ , \new_[32873]_ , \new_[32877]_ ,
    \new_[32878]_ , \new_[32879]_ , \new_[32883]_ , \new_[32884]_ ,
    \new_[32887]_ , \new_[32890]_ , \new_[32891]_ , \new_[32892]_ ,
    \new_[32896]_ , \new_[32897]_ , \new_[32901]_ , \new_[32902]_ ,
    \new_[32903]_ , \new_[32907]_ , \new_[32908]_ , \new_[32911]_ ,
    \new_[32914]_ , \new_[32915]_ , \new_[32916]_ , \new_[32920]_ ,
    \new_[32921]_ , \new_[32925]_ , \new_[32926]_ , \new_[32927]_ ,
    \new_[32931]_ , \new_[32932]_ , \new_[32935]_ , \new_[32938]_ ,
    \new_[32939]_ , \new_[32940]_ , \new_[32944]_ , \new_[32945]_ ,
    \new_[32949]_ , \new_[32950]_ , \new_[32951]_ , \new_[32955]_ ,
    \new_[32956]_ , \new_[32959]_ , \new_[32962]_ , \new_[32963]_ ,
    \new_[32964]_ , \new_[32968]_ , \new_[32969]_ , \new_[32973]_ ,
    \new_[32974]_ , \new_[32975]_ , \new_[32979]_ , \new_[32980]_ ,
    \new_[32983]_ , \new_[32986]_ , \new_[32987]_ , \new_[32988]_ ,
    \new_[32992]_ , \new_[32993]_ , \new_[32997]_ , \new_[32998]_ ,
    \new_[32999]_ , \new_[33003]_ , \new_[33004]_ , \new_[33007]_ ,
    \new_[33010]_ , \new_[33011]_ , \new_[33012]_ , \new_[33016]_ ,
    \new_[33017]_ , \new_[33021]_ , \new_[33022]_ , \new_[33023]_ ,
    \new_[33027]_ , \new_[33028]_ , \new_[33031]_ , \new_[33034]_ ,
    \new_[33035]_ , \new_[33036]_ , \new_[33040]_ , \new_[33041]_ ,
    \new_[33045]_ , \new_[33046]_ , \new_[33047]_ , \new_[33051]_ ,
    \new_[33052]_ , \new_[33055]_ , \new_[33058]_ , \new_[33059]_ ,
    \new_[33060]_ , \new_[33064]_ , \new_[33065]_ , \new_[33069]_ ,
    \new_[33070]_ , \new_[33071]_ , \new_[33075]_ , \new_[33076]_ ,
    \new_[33079]_ , \new_[33082]_ , \new_[33083]_ , \new_[33084]_ ,
    \new_[33088]_ , \new_[33089]_ , \new_[33093]_ , \new_[33094]_ ,
    \new_[33095]_ , \new_[33099]_ , \new_[33100]_ , \new_[33103]_ ,
    \new_[33106]_ , \new_[33107]_ , \new_[33108]_ , \new_[33112]_ ,
    \new_[33113]_ , \new_[33117]_ , \new_[33118]_ , \new_[33119]_ ,
    \new_[33123]_ , \new_[33124]_ , \new_[33127]_ , \new_[33130]_ ,
    \new_[33131]_ , \new_[33132]_ , \new_[33136]_ , \new_[33137]_ ,
    \new_[33141]_ , \new_[33142]_ , \new_[33143]_ , \new_[33147]_ ,
    \new_[33148]_ , \new_[33151]_ , \new_[33154]_ , \new_[33155]_ ,
    \new_[33156]_ , \new_[33160]_ , \new_[33161]_ , \new_[33165]_ ,
    \new_[33166]_ , \new_[33167]_ , \new_[33171]_ , \new_[33172]_ ,
    \new_[33175]_ , \new_[33178]_ , \new_[33179]_ , \new_[33180]_ ,
    \new_[33184]_ , \new_[33185]_ , \new_[33189]_ , \new_[33190]_ ,
    \new_[33191]_ , \new_[33195]_ , \new_[33196]_ , \new_[33199]_ ,
    \new_[33202]_ , \new_[33203]_ , \new_[33204]_ , \new_[33208]_ ,
    \new_[33209]_ , \new_[33213]_ , \new_[33214]_ , \new_[33215]_ ,
    \new_[33219]_ , \new_[33220]_ , \new_[33223]_ , \new_[33226]_ ,
    \new_[33227]_ , \new_[33228]_ , \new_[33232]_ , \new_[33233]_ ,
    \new_[33237]_ , \new_[33238]_ , \new_[33239]_ , \new_[33243]_ ,
    \new_[33244]_ , \new_[33247]_ , \new_[33250]_ , \new_[33251]_ ,
    \new_[33252]_ , \new_[33256]_ , \new_[33257]_ , \new_[33261]_ ,
    \new_[33262]_ , \new_[33263]_ , \new_[33267]_ , \new_[33268]_ ,
    \new_[33271]_ , \new_[33274]_ , \new_[33275]_ , \new_[33276]_ ,
    \new_[33280]_ , \new_[33281]_ , \new_[33285]_ , \new_[33286]_ ,
    \new_[33287]_ , \new_[33291]_ , \new_[33292]_ , \new_[33295]_ ,
    \new_[33298]_ , \new_[33299]_ , \new_[33300]_ , \new_[33304]_ ,
    \new_[33305]_ , \new_[33309]_ , \new_[33310]_ , \new_[33311]_ ,
    \new_[33315]_ , \new_[33316]_ , \new_[33319]_ , \new_[33322]_ ,
    \new_[33323]_ , \new_[33324]_ , \new_[33328]_ , \new_[33329]_ ,
    \new_[33333]_ , \new_[33334]_ , \new_[33335]_ , \new_[33339]_ ,
    \new_[33340]_ , \new_[33343]_ , \new_[33346]_ , \new_[33347]_ ,
    \new_[33348]_ , \new_[33352]_ , \new_[33353]_ , \new_[33357]_ ,
    \new_[33358]_ , \new_[33359]_ , \new_[33363]_ , \new_[33364]_ ,
    \new_[33367]_ , \new_[33370]_ , \new_[33371]_ , \new_[33372]_ ,
    \new_[33376]_ , \new_[33377]_ , \new_[33381]_ , \new_[33382]_ ,
    \new_[33383]_ , \new_[33387]_ , \new_[33388]_ , \new_[33391]_ ,
    \new_[33394]_ , \new_[33395]_ , \new_[33396]_ , \new_[33400]_ ,
    \new_[33401]_ , \new_[33405]_ , \new_[33406]_ , \new_[33407]_ ,
    \new_[33411]_ , \new_[33412]_ , \new_[33415]_ , \new_[33418]_ ,
    \new_[33419]_ , \new_[33420]_ , \new_[33424]_ , \new_[33425]_ ,
    \new_[33429]_ , \new_[33430]_ , \new_[33431]_ , \new_[33435]_ ,
    \new_[33436]_ , \new_[33439]_ , \new_[33442]_ , \new_[33443]_ ,
    \new_[33444]_ , \new_[33448]_ , \new_[33449]_ , \new_[33453]_ ,
    \new_[33454]_ , \new_[33455]_ , \new_[33459]_ , \new_[33460]_ ,
    \new_[33463]_ , \new_[33466]_ , \new_[33467]_ , \new_[33468]_ ,
    \new_[33472]_ , \new_[33473]_ , \new_[33477]_ , \new_[33478]_ ,
    \new_[33479]_ , \new_[33483]_ , \new_[33484]_ , \new_[33487]_ ,
    \new_[33490]_ , \new_[33491]_ , \new_[33492]_ , \new_[33496]_ ,
    \new_[33497]_ , \new_[33501]_ , \new_[33502]_ , \new_[33503]_ ,
    \new_[33507]_ , \new_[33508]_ , \new_[33511]_ , \new_[33514]_ ,
    \new_[33515]_ , \new_[33516]_ , \new_[33520]_ , \new_[33521]_ ,
    \new_[33525]_ , \new_[33526]_ , \new_[33527]_ , \new_[33531]_ ,
    \new_[33532]_ , \new_[33535]_ , \new_[33538]_ , \new_[33539]_ ,
    \new_[33540]_ , \new_[33544]_ , \new_[33545]_ , \new_[33549]_ ,
    \new_[33550]_ , \new_[33551]_ , \new_[33555]_ , \new_[33556]_ ,
    \new_[33559]_ , \new_[33562]_ , \new_[33563]_ , \new_[33564]_ ,
    \new_[33568]_ , \new_[33569]_ , \new_[33573]_ , \new_[33574]_ ,
    \new_[33575]_ , \new_[33579]_ , \new_[33580]_ , \new_[33583]_ ,
    \new_[33586]_ , \new_[33587]_ , \new_[33588]_ , \new_[33592]_ ,
    \new_[33593]_ , \new_[33597]_ , \new_[33598]_ , \new_[33599]_ ,
    \new_[33603]_ , \new_[33604]_ , \new_[33607]_ , \new_[33610]_ ,
    \new_[33611]_ , \new_[33612]_ , \new_[33616]_ , \new_[33617]_ ,
    \new_[33621]_ , \new_[33622]_ , \new_[33623]_ , \new_[33627]_ ,
    \new_[33628]_ , \new_[33631]_ , \new_[33634]_ , \new_[33635]_ ,
    \new_[33636]_ , \new_[33640]_ , \new_[33641]_ , \new_[33645]_ ,
    \new_[33646]_ , \new_[33647]_ , \new_[33651]_ , \new_[33652]_ ,
    \new_[33655]_ , \new_[33658]_ , \new_[33659]_ , \new_[33660]_ ,
    \new_[33664]_ , \new_[33665]_ , \new_[33669]_ , \new_[33670]_ ,
    \new_[33671]_ , \new_[33675]_ , \new_[33676]_ , \new_[33679]_ ,
    \new_[33682]_ , \new_[33683]_ , \new_[33684]_ , \new_[33688]_ ,
    \new_[33689]_ , \new_[33693]_ , \new_[33694]_ , \new_[33695]_ ,
    \new_[33699]_ , \new_[33700]_ , \new_[33703]_ , \new_[33706]_ ,
    \new_[33707]_ , \new_[33708]_ , \new_[33712]_ , \new_[33713]_ ,
    \new_[33717]_ , \new_[33718]_ , \new_[33719]_ , \new_[33723]_ ,
    \new_[33724]_ , \new_[33727]_ , \new_[33730]_ , \new_[33731]_ ,
    \new_[33732]_ , \new_[33736]_ , \new_[33737]_ , \new_[33741]_ ,
    \new_[33742]_ , \new_[33743]_ , \new_[33747]_ , \new_[33748]_ ,
    \new_[33751]_ , \new_[33754]_ , \new_[33755]_ , \new_[33756]_ ,
    \new_[33760]_ , \new_[33761]_ , \new_[33765]_ , \new_[33766]_ ,
    \new_[33767]_ , \new_[33771]_ , \new_[33772]_ , \new_[33775]_ ,
    \new_[33778]_ , \new_[33779]_ , \new_[33780]_ , \new_[33784]_ ,
    \new_[33785]_ , \new_[33789]_ , \new_[33790]_ , \new_[33791]_ ,
    \new_[33795]_ , \new_[33796]_ , \new_[33799]_ , \new_[33802]_ ,
    \new_[33803]_ , \new_[33804]_ , \new_[33808]_ , \new_[33809]_ ,
    \new_[33813]_ , \new_[33814]_ , \new_[33815]_ , \new_[33819]_ ,
    \new_[33820]_ , \new_[33823]_ , \new_[33826]_ , \new_[33827]_ ,
    \new_[33828]_ , \new_[33832]_ , \new_[33833]_ , \new_[33837]_ ,
    \new_[33838]_ , \new_[33839]_ , \new_[33843]_ , \new_[33844]_ ,
    \new_[33847]_ , \new_[33850]_ , \new_[33851]_ , \new_[33852]_ ,
    \new_[33856]_ , \new_[33857]_ , \new_[33861]_ , \new_[33862]_ ,
    \new_[33863]_ , \new_[33867]_ , \new_[33868]_ , \new_[33871]_ ,
    \new_[33874]_ , \new_[33875]_ , \new_[33876]_ , \new_[33880]_ ,
    \new_[33881]_ , \new_[33885]_ , \new_[33886]_ , \new_[33887]_ ,
    \new_[33891]_ , \new_[33892]_ , \new_[33895]_ , \new_[33898]_ ,
    \new_[33899]_ , \new_[33900]_ , \new_[33904]_ , \new_[33905]_ ,
    \new_[33909]_ , \new_[33910]_ , \new_[33911]_ , \new_[33915]_ ,
    \new_[33916]_ , \new_[33919]_ , \new_[33922]_ , \new_[33923]_ ,
    \new_[33924]_ , \new_[33928]_ , \new_[33929]_ , \new_[33933]_ ,
    \new_[33934]_ , \new_[33935]_ , \new_[33939]_ , \new_[33940]_ ,
    \new_[33943]_ , \new_[33946]_ , \new_[33947]_ , \new_[33948]_ ,
    \new_[33952]_ , \new_[33953]_ , \new_[33957]_ , \new_[33958]_ ,
    \new_[33959]_ , \new_[33963]_ , \new_[33964]_ , \new_[33967]_ ,
    \new_[33970]_ , \new_[33971]_ , \new_[33972]_ , \new_[33976]_ ,
    \new_[33977]_ , \new_[33981]_ , \new_[33982]_ , \new_[33983]_ ,
    \new_[33987]_ , \new_[33988]_ , \new_[33991]_ , \new_[33994]_ ,
    \new_[33995]_ , \new_[33996]_ , \new_[34000]_ , \new_[34001]_ ,
    \new_[34005]_ , \new_[34006]_ , \new_[34007]_ , \new_[34011]_ ,
    \new_[34012]_ , \new_[34015]_ , \new_[34018]_ , \new_[34019]_ ,
    \new_[34020]_ , \new_[34024]_ , \new_[34025]_ , \new_[34029]_ ,
    \new_[34030]_ , \new_[34031]_ , \new_[34035]_ , \new_[34036]_ ,
    \new_[34039]_ , \new_[34042]_ , \new_[34043]_ , \new_[34044]_ ,
    \new_[34048]_ , \new_[34049]_ , \new_[34053]_ , \new_[34054]_ ,
    \new_[34055]_ , \new_[34059]_ , \new_[34060]_ , \new_[34063]_ ,
    \new_[34066]_ , \new_[34067]_ , \new_[34068]_ , \new_[34072]_ ,
    \new_[34073]_ , \new_[34077]_ , \new_[34078]_ , \new_[34079]_ ,
    \new_[34083]_ , \new_[34084]_ , \new_[34087]_ , \new_[34090]_ ,
    \new_[34091]_ , \new_[34092]_ , \new_[34096]_ , \new_[34097]_ ,
    \new_[34101]_ , \new_[34102]_ , \new_[34103]_ , \new_[34107]_ ,
    \new_[34108]_ , \new_[34111]_ , \new_[34114]_ , \new_[34115]_ ,
    \new_[34116]_ , \new_[34120]_ , \new_[34121]_ , \new_[34125]_ ,
    \new_[34126]_ , \new_[34127]_ , \new_[34131]_ , \new_[34132]_ ,
    \new_[34135]_ , \new_[34138]_ , \new_[34139]_ , \new_[34140]_ ,
    \new_[34144]_ , \new_[34145]_ , \new_[34149]_ , \new_[34150]_ ,
    \new_[34151]_ , \new_[34155]_ , \new_[34156]_ , \new_[34159]_ ,
    \new_[34162]_ , \new_[34163]_ , \new_[34164]_ , \new_[34168]_ ,
    \new_[34169]_ , \new_[34173]_ , \new_[34174]_ , \new_[34175]_ ,
    \new_[34179]_ , \new_[34180]_ , \new_[34183]_ , \new_[34186]_ ,
    \new_[34187]_ , \new_[34188]_ , \new_[34192]_ , \new_[34193]_ ,
    \new_[34197]_ , \new_[34198]_ , \new_[34199]_ , \new_[34203]_ ,
    \new_[34204]_ , \new_[34207]_ , \new_[34210]_ , \new_[34211]_ ,
    \new_[34212]_ , \new_[34216]_ , \new_[34217]_ , \new_[34221]_ ,
    \new_[34222]_ , \new_[34223]_ , \new_[34227]_ , \new_[34228]_ ,
    \new_[34231]_ , \new_[34234]_ , \new_[34235]_ , \new_[34236]_ ,
    \new_[34240]_ , \new_[34241]_ , \new_[34245]_ , \new_[34246]_ ,
    \new_[34247]_ , \new_[34251]_ , \new_[34252]_ , \new_[34255]_ ,
    \new_[34258]_ , \new_[34259]_ , \new_[34260]_ , \new_[34264]_ ,
    \new_[34265]_ , \new_[34269]_ , \new_[34270]_ , \new_[34271]_ ,
    \new_[34275]_ , \new_[34276]_ , \new_[34279]_ , \new_[34282]_ ,
    \new_[34283]_ , \new_[34284]_ , \new_[34288]_ , \new_[34289]_ ,
    \new_[34293]_ , \new_[34294]_ , \new_[34295]_ , \new_[34299]_ ,
    \new_[34300]_ , \new_[34303]_ , \new_[34306]_ , \new_[34307]_ ,
    \new_[34308]_ , \new_[34312]_ , \new_[34313]_ , \new_[34317]_ ,
    \new_[34318]_ , \new_[34319]_ , \new_[34323]_ , \new_[34324]_ ,
    \new_[34327]_ , \new_[34330]_ , \new_[34331]_ , \new_[34332]_ ,
    \new_[34336]_ , \new_[34337]_ , \new_[34341]_ , \new_[34342]_ ,
    \new_[34343]_ , \new_[34347]_ , \new_[34348]_ , \new_[34351]_ ,
    \new_[34354]_ , \new_[34355]_ , \new_[34356]_ , \new_[34360]_ ,
    \new_[34361]_ , \new_[34365]_ , \new_[34366]_ , \new_[34367]_ ,
    \new_[34371]_ , \new_[34372]_ , \new_[34375]_ , \new_[34378]_ ,
    \new_[34379]_ , \new_[34380]_ , \new_[34384]_ , \new_[34385]_ ,
    \new_[34389]_ , \new_[34390]_ , \new_[34391]_ , \new_[34395]_ ,
    \new_[34396]_ , \new_[34399]_ , \new_[34402]_ , \new_[34403]_ ,
    \new_[34404]_ , \new_[34408]_ , \new_[34409]_ , \new_[34413]_ ,
    \new_[34414]_ , \new_[34415]_ , \new_[34419]_ , \new_[34420]_ ,
    \new_[34423]_ , \new_[34426]_ , \new_[34427]_ , \new_[34428]_ ,
    \new_[34432]_ , \new_[34433]_ , \new_[34437]_ , \new_[34438]_ ,
    \new_[34439]_ , \new_[34443]_ , \new_[34444]_ , \new_[34447]_ ,
    \new_[34450]_ , \new_[34451]_ , \new_[34452]_ , \new_[34456]_ ,
    \new_[34457]_ , \new_[34461]_ , \new_[34462]_ , \new_[34463]_ ,
    \new_[34467]_ , \new_[34468]_ , \new_[34471]_ , \new_[34474]_ ,
    \new_[34475]_ , \new_[34476]_ , \new_[34480]_ , \new_[34481]_ ,
    \new_[34485]_ , \new_[34486]_ , \new_[34487]_ , \new_[34491]_ ,
    \new_[34492]_ , \new_[34495]_ , \new_[34498]_ , \new_[34499]_ ,
    \new_[34500]_ , \new_[34504]_ , \new_[34505]_ , \new_[34509]_ ,
    \new_[34510]_ , \new_[34511]_ , \new_[34515]_ , \new_[34516]_ ,
    \new_[34519]_ , \new_[34522]_ , \new_[34523]_ , \new_[34524]_ ,
    \new_[34528]_ , \new_[34529]_ , \new_[34533]_ , \new_[34534]_ ,
    \new_[34535]_ , \new_[34539]_ , \new_[34540]_ , \new_[34543]_ ,
    \new_[34546]_ , \new_[34547]_ , \new_[34548]_ , \new_[34552]_ ,
    \new_[34553]_ , \new_[34557]_ , \new_[34558]_ , \new_[34559]_ ,
    \new_[34563]_ , \new_[34564]_ , \new_[34567]_ , \new_[34570]_ ,
    \new_[34571]_ , \new_[34572]_ , \new_[34576]_ , \new_[34577]_ ,
    \new_[34581]_ , \new_[34582]_ , \new_[34583]_ , \new_[34587]_ ,
    \new_[34588]_ , \new_[34591]_ , \new_[34594]_ , \new_[34595]_ ,
    \new_[34596]_ , \new_[34600]_ , \new_[34601]_ , \new_[34605]_ ,
    \new_[34606]_ , \new_[34607]_ , \new_[34611]_ , \new_[34612]_ ,
    \new_[34615]_ , \new_[34618]_ , \new_[34619]_ , \new_[34620]_ ,
    \new_[34624]_ , \new_[34625]_ , \new_[34629]_ , \new_[34630]_ ,
    \new_[34631]_ , \new_[34635]_ , \new_[34636]_ , \new_[34639]_ ,
    \new_[34642]_ , \new_[34643]_ , \new_[34644]_ , \new_[34648]_ ,
    \new_[34649]_ , \new_[34653]_ , \new_[34654]_ , \new_[34655]_ ,
    \new_[34659]_ , \new_[34660]_ , \new_[34663]_ , \new_[34666]_ ,
    \new_[34667]_ , \new_[34668]_ , \new_[34672]_ , \new_[34673]_ ,
    \new_[34677]_ , \new_[34678]_ , \new_[34679]_ , \new_[34683]_ ,
    \new_[34684]_ , \new_[34687]_ , \new_[34690]_ , \new_[34691]_ ,
    \new_[34692]_ , \new_[34696]_ , \new_[34697]_ , \new_[34701]_ ,
    \new_[34702]_ , \new_[34703]_ , \new_[34707]_ , \new_[34708]_ ,
    \new_[34711]_ , \new_[34714]_ , \new_[34715]_ , \new_[34716]_ ,
    \new_[34720]_ , \new_[34721]_ , \new_[34725]_ , \new_[34726]_ ,
    \new_[34727]_ , \new_[34731]_ , \new_[34732]_ , \new_[34735]_ ,
    \new_[34738]_ , \new_[34739]_ , \new_[34740]_ , \new_[34744]_ ,
    \new_[34745]_ , \new_[34749]_ , \new_[34750]_ , \new_[34751]_ ,
    \new_[34755]_ , \new_[34756]_ , \new_[34759]_ , \new_[34762]_ ,
    \new_[34763]_ , \new_[34764]_ , \new_[34768]_ , \new_[34769]_ ,
    \new_[34773]_ , \new_[34774]_ , \new_[34775]_ , \new_[34779]_ ,
    \new_[34780]_ , \new_[34783]_ , \new_[34786]_ , \new_[34787]_ ,
    \new_[34788]_ , \new_[34792]_ , \new_[34793]_ , \new_[34797]_ ,
    \new_[34798]_ , \new_[34799]_ , \new_[34803]_ , \new_[34804]_ ,
    \new_[34807]_ , \new_[34810]_ , \new_[34811]_ , \new_[34812]_ ,
    \new_[34816]_ , \new_[34817]_ , \new_[34821]_ , \new_[34822]_ ,
    \new_[34823]_ , \new_[34827]_ , \new_[34828]_ , \new_[34831]_ ,
    \new_[34834]_ , \new_[34835]_ , \new_[34836]_ , \new_[34840]_ ,
    \new_[34841]_ , \new_[34845]_ , \new_[34846]_ , \new_[34847]_ ,
    \new_[34851]_ , \new_[34852]_ , \new_[34855]_ , \new_[34858]_ ,
    \new_[34859]_ , \new_[34860]_ , \new_[34864]_ , \new_[34865]_ ,
    \new_[34869]_ , \new_[34870]_ , \new_[34871]_ , \new_[34875]_ ,
    \new_[34876]_ , \new_[34879]_ , \new_[34882]_ , \new_[34883]_ ,
    \new_[34884]_ , \new_[34888]_ , \new_[34889]_ , \new_[34893]_ ,
    \new_[34894]_ , \new_[34895]_ , \new_[34899]_ , \new_[34900]_ ,
    \new_[34903]_ , \new_[34906]_ , \new_[34907]_ , \new_[34908]_ ,
    \new_[34912]_ , \new_[34913]_ , \new_[34917]_ , \new_[34918]_ ,
    \new_[34919]_ , \new_[34923]_ , \new_[34924]_ , \new_[34927]_ ,
    \new_[34930]_ , \new_[34931]_ , \new_[34932]_ , \new_[34936]_ ,
    \new_[34937]_ , \new_[34941]_ , \new_[34942]_ , \new_[34943]_ ,
    \new_[34947]_ , \new_[34948]_ , \new_[34951]_ , \new_[34954]_ ,
    \new_[34955]_ , \new_[34956]_ , \new_[34960]_ , \new_[34961]_ ,
    \new_[34965]_ , \new_[34966]_ , \new_[34967]_ , \new_[34971]_ ,
    \new_[34972]_ , \new_[34975]_ , \new_[34978]_ , \new_[34979]_ ,
    \new_[34980]_ , \new_[34984]_ , \new_[34985]_ , \new_[34989]_ ,
    \new_[34990]_ , \new_[34991]_ , \new_[34995]_ , \new_[34996]_ ,
    \new_[34999]_ , \new_[35002]_ , \new_[35003]_ , \new_[35004]_ ,
    \new_[35008]_ , \new_[35009]_ , \new_[35013]_ , \new_[35014]_ ,
    \new_[35015]_ , \new_[35019]_ , \new_[35020]_ , \new_[35023]_ ,
    \new_[35026]_ , \new_[35027]_ , \new_[35028]_ , \new_[35032]_ ,
    \new_[35033]_ , \new_[35037]_ , \new_[35038]_ , \new_[35039]_ ,
    \new_[35043]_ , \new_[35044]_ , \new_[35047]_ , \new_[35050]_ ,
    \new_[35051]_ , \new_[35052]_ , \new_[35056]_ , \new_[35057]_ ,
    \new_[35061]_ , \new_[35062]_ , \new_[35063]_ , \new_[35067]_ ,
    \new_[35068]_ , \new_[35071]_ , \new_[35074]_ , \new_[35075]_ ,
    \new_[35076]_ , \new_[35080]_ , \new_[35081]_ , \new_[35085]_ ,
    \new_[35086]_ , \new_[35087]_ , \new_[35091]_ , \new_[35092]_ ,
    \new_[35095]_ , \new_[35098]_ , \new_[35099]_ , \new_[35100]_ ,
    \new_[35104]_ , \new_[35105]_ , \new_[35109]_ , \new_[35110]_ ,
    \new_[35111]_ , \new_[35115]_ , \new_[35116]_ , \new_[35119]_ ,
    \new_[35122]_ , \new_[35123]_ , \new_[35124]_ , \new_[35128]_ ,
    \new_[35129]_ , \new_[35133]_ , \new_[35134]_ , \new_[35135]_ ,
    \new_[35139]_ , \new_[35140]_ , \new_[35143]_ , \new_[35146]_ ,
    \new_[35147]_ , \new_[35148]_ , \new_[35152]_ , \new_[35153]_ ,
    \new_[35157]_ , \new_[35158]_ , \new_[35159]_ , \new_[35163]_ ,
    \new_[35164]_ , \new_[35167]_ , \new_[35170]_ , \new_[35171]_ ,
    \new_[35172]_ , \new_[35176]_ , \new_[35177]_ , \new_[35181]_ ,
    \new_[35182]_ , \new_[35183]_ , \new_[35187]_ , \new_[35188]_ ,
    \new_[35191]_ , \new_[35194]_ , \new_[35195]_ , \new_[35196]_ ,
    \new_[35200]_ , \new_[35201]_ , \new_[35205]_ , \new_[35206]_ ,
    \new_[35207]_ , \new_[35211]_ , \new_[35212]_ , \new_[35215]_ ,
    \new_[35218]_ , \new_[35219]_ , \new_[35220]_ , \new_[35224]_ ,
    \new_[35225]_ , \new_[35229]_ , \new_[35230]_ , \new_[35231]_ ,
    \new_[35235]_ , \new_[35236]_ , \new_[35239]_ , \new_[35242]_ ,
    \new_[35243]_ , \new_[35244]_ , \new_[35248]_ , \new_[35249]_ ,
    \new_[35253]_ , \new_[35254]_ , \new_[35255]_ , \new_[35259]_ ,
    \new_[35260]_ , \new_[35263]_ , \new_[35266]_ , \new_[35267]_ ,
    \new_[35268]_ , \new_[35272]_ , \new_[35273]_ , \new_[35277]_ ,
    \new_[35278]_ , \new_[35279]_ , \new_[35283]_ , \new_[35284]_ ,
    \new_[35287]_ , \new_[35290]_ , \new_[35291]_ , \new_[35292]_ ,
    \new_[35296]_ , \new_[35297]_ , \new_[35301]_ , \new_[35302]_ ,
    \new_[35303]_ , \new_[35307]_ , \new_[35308]_ , \new_[35311]_ ,
    \new_[35314]_ , \new_[35315]_ , \new_[35316]_ , \new_[35320]_ ,
    \new_[35321]_ , \new_[35325]_ , \new_[35326]_ , \new_[35327]_ ,
    \new_[35331]_ , \new_[35332]_ , \new_[35335]_ , \new_[35338]_ ,
    \new_[35339]_ , \new_[35340]_ , \new_[35344]_ , \new_[35345]_ ,
    \new_[35349]_ , \new_[35350]_ , \new_[35351]_ , \new_[35355]_ ,
    \new_[35356]_ , \new_[35359]_ , \new_[35362]_ , \new_[35363]_ ,
    \new_[35364]_ , \new_[35368]_ , \new_[35369]_ , \new_[35373]_ ,
    \new_[35374]_ , \new_[35375]_ , \new_[35379]_ , \new_[35380]_ ,
    \new_[35383]_ , \new_[35386]_ , \new_[35387]_ , \new_[35388]_ ,
    \new_[35392]_ , \new_[35393]_ , \new_[35397]_ , \new_[35398]_ ,
    \new_[35399]_ , \new_[35403]_ , \new_[35404]_ , \new_[35407]_ ,
    \new_[35410]_ , \new_[35411]_ , \new_[35412]_ , \new_[35416]_ ,
    \new_[35417]_ , \new_[35421]_ , \new_[35422]_ , \new_[35423]_ ,
    \new_[35427]_ , \new_[35428]_ , \new_[35431]_ , \new_[35434]_ ,
    \new_[35435]_ , \new_[35436]_ , \new_[35440]_ , \new_[35441]_ ,
    \new_[35445]_ , \new_[35446]_ , \new_[35447]_ , \new_[35451]_ ,
    \new_[35452]_ , \new_[35455]_ , \new_[35458]_ , \new_[35459]_ ,
    \new_[35460]_ , \new_[35464]_ , \new_[35465]_ , \new_[35469]_ ,
    \new_[35470]_ , \new_[35471]_ , \new_[35475]_ , \new_[35476]_ ,
    \new_[35479]_ , \new_[35482]_ , \new_[35483]_ , \new_[35484]_ ,
    \new_[35488]_ , \new_[35489]_ , \new_[35493]_ , \new_[35494]_ ,
    \new_[35495]_ , \new_[35499]_ , \new_[35500]_ , \new_[35503]_ ,
    \new_[35506]_ , \new_[35507]_ , \new_[35508]_ , \new_[35512]_ ,
    \new_[35513]_ , \new_[35517]_ , \new_[35518]_ , \new_[35519]_ ,
    \new_[35523]_ , \new_[35524]_ , \new_[35527]_ , \new_[35530]_ ,
    \new_[35531]_ , \new_[35532]_ , \new_[35536]_ , \new_[35537]_ ,
    \new_[35541]_ , \new_[35542]_ , \new_[35543]_ , \new_[35547]_ ,
    \new_[35548]_ , \new_[35551]_ , \new_[35554]_ , \new_[35555]_ ,
    \new_[35556]_ , \new_[35560]_ , \new_[35561]_ , \new_[35565]_ ,
    \new_[35566]_ , \new_[35567]_ , \new_[35571]_ , \new_[35572]_ ,
    \new_[35575]_ , \new_[35578]_ , \new_[35579]_ , \new_[35580]_ ,
    \new_[35584]_ , \new_[35585]_ , \new_[35589]_ , \new_[35590]_ ,
    \new_[35591]_ , \new_[35595]_ , \new_[35596]_ , \new_[35599]_ ,
    \new_[35602]_ , \new_[35603]_ , \new_[35604]_ , \new_[35608]_ ,
    \new_[35609]_ , \new_[35613]_ , \new_[35614]_ , \new_[35615]_ ,
    \new_[35619]_ , \new_[35620]_ , \new_[35623]_ , \new_[35626]_ ,
    \new_[35627]_ , \new_[35628]_ , \new_[35632]_ , \new_[35633]_ ,
    \new_[35637]_ , \new_[35638]_ , \new_[35639]_ , \new_[35643]_ ,
    \new_[35644]_ , \new_[35647]_ , \new_[35650]_ , \new_[35651]_ ,
    \new_[35652]_ , \new_[35656]_ , \new_[35657]_ , \new_[35661]_ ,
    \new_[35662]_ , \new_[35663]_ , \new_[35667]_ , \new_[35668]_ ,
    \new_[35671]_ , \new_[35674]_ , \new_[35675]_ , \new_[35676]_ ,
    \new_[35680]_ , \new_[35681]_ , \new_[35685]_ , \new_[35686]_ ,
    \new_[35687]_ , \new_[35691]_ , \new_[35692]_ , \new_[35695]_ ,
    \new_[35698]_ , \new_[35699]_ , \new_[35700]_ , \new_[35704]_ ,
    \new_[35705]_ , \new_[35709]_ , \new_[35710]_ , \new_[35711]_ ,
    \new_[35715]_ , \new_[35716]_ , \new_[35719]_ , \new_[35722]_ ,
    \new_[35723]_ , \new_[35724]_ , \new_[35728]_ , \new_[35729]_ ,
    \new_[35733]_ , \new_[35734]_ , \new_[35735]_ , \new_[35739]_ ,
    \new_[35740]_ , \new_[35743]_ , \new_[35746]_ , \new_[35747]_ ,
    \new_[35748]_ , \new_[35752]_ , \new_[35753]_ , \new_[35757]_ ,
    \new_[35758]_ , \new_[35759]_ , \new_[35763]_ , \new_[35764]_ ,
    \new_[35767]_ , \new_[35770]_ , \new_[35771]_ , \new_[35772]_ ,
    \new_[35776]_ , \new_[35777]_ , \new_[35781]_ , \new_[35782]_ ,
    \new_[35783]_ , \new_[35787]_ , \new_[35788]_ , \new_[35791]_ ,
    \new_[35794]_ , \new_[35795]_ , \new_[35796]_ , \new_[35800]_ ,
    \new_[35801]_ , \new_[35805]_ , \new_[35806]_ , \new_[35807]_ ,
    \new_[35811]_ , \new_[35812]_ , \new_[35815]_ , \new_[35818]_ ,
    \new_[35819]_ , \new_[35820]_ , \new_[35824]_ , \new_[35825]_ ,
    \new_[35829]_ , \new_[35830]_ , \new_[35831]_ , \new_[35835]_ ,
    \new_[35836]_ , \new_[35839]_ , \new_[35842]_ , \new_[35843]_ ,
    \new_[35844]_ , \new_[35848]_ , \new_[35849]_ , \new_[35853]_ ,
    \new_[35854]_ , \new_[35855]_ , \new_[35859]_ , \new_[35860]_ ,
    \new_[35863]_ , \new_[35866]_ , \new_[35867]_ , \new_[35868]_ ,
    \new_[35872]_ , \new_[35873]_ , \new_[35877]_ , \new_[35878]_ ,
    \new_[35879]_ , \new_[35883]_ , \new_[35884]_ , \new_[35887]_ ,
    \new_[35890]_ , \new_[35891]_ , \new_[35892]_ , \new_[35896]_ ,
    \new_[35897]_ , \new_[35901]_ , \new_[35902]_ , \new_[35903]_ ,
    \new_[35907]_ , \new_[35908]_ , \new_[35911]_ , \new_[35914]_ ,
    \new_[35915]_ , \new_[35916]_ , \new_[35920]_ , \new_[35921]_ ,
    \new_[35925]_ , \new_[35926]_ , \new_[35927]_ , \new_[35931]_ ,
    \new_[35932]_ , \new_[35935]_ , \new_[35938]_ , \new_[35939]_ ,
    \new_[35940]_ , \new_[35944]_ , \new_[35945]_ , \new_[35949]_ ,
    \new_[35950]_ , \new_[35951]_ , \new_[35955]_ , \new_[35956]_ ,
    \new_[35959]_ , \new_[35962]_ , \new_[35963]_ , \new_[35964]_ ,
    \new_[35968]_ , \new_[35969]_ , \new_[35973]_ , \new_[35974]_ ,
    \new_[35975]_ , \new_[35979]_ , \new_[35980]_ , \new_[35983]_ ,
    \new_[35986]_ , \new_[35987]_ , \new_[35988]_ , \new_[35992]_ ,
    \new_[35993]_ , \new_[35997]_ , \new_[35998]_ , \new_[35999]_ ,
    \new_[36003]_ , \new_[36004]_ , \new_[36007]_ , \new_[36010]_ ,
    \new_[36011]_ , \new_[36012]_ , \new_[36016]_ , \new_[36017]_ ,
    \new_[36021]_ , \new_[36022]_ , \new_[36023]_ , \new_[36027]_ ,
    \new_[36028]_ , \new_[36031]_ , \new_[36034]_ , \new_[36035]_ ,
    \new_[36036]_ , \new_[36040]_ , \new_[36041]_ , \new_[36045]_ ,
    \new_[36046]_ , \new_[36047]_ , \new_[36051]_ , \new_[36052]_ ,
    \new_[36055]_ , \new_[36058]_ , \new_[36059]_ , \new_[36060]_ ,
    \new_[36064]_ , \new_[36065]_ , \new_[36069]_ , \new_[36070]_ ,
    \new_[36071]_ , \new_[36075]_ , \new_[36076]_ , \new_[36079]_ ,
    \new_[36082]_ , \new_[36083]_ , \new_[36084]_ , \new_[36088]_ ,
    \new_[36089]_ , \new_[36093]_ , \new_[36094]_ , \new_[36095]_ ,
    \new_[36099]_ , \new_[36100]_ , \new_[36103]_ , \new_[36106]_ ,
    \new_[36107]_ , \new_[36108]_ , \new_[36112]_ , \new_[36113]_ ,
    \new_[36117]_ , \new_[36118]_ , \new_[36119]_ , \new_[36123]_ ,
    \new_[36124]_ , \new_[36127]_ , \new_[36130]_ , \new_[36131]_ ,
    \new_[36132]_ , \new_[36136]_ , \new_[36137]_ , \new_[36141]_ ,
    \new_[36142]_ , \new_[36143]_ , \new_[36147]_ , \new_[36148]_ ,
    \new_[36151]_ , \new_[36154]_ , \new_[36155]_ , \new_[36156]_ ,
    \new_[36160]_ , \new_[36161]_ , \new_[36165]_ , \new_[36166]_ ,
    \new_[36167]_ , \new_[36171]_ , \new_[36172]_ , \new_[36175]_ ,
    \new_[36178]_ , \new_[36179]_ , \new_[36180]_ , \new_[36184]_ ,
    \new_[36185]_ , \new_[36189]_ , \new_[36190]_ , \new_[36191]_ ,
    \new_[36195]_ , \new_[36196]_ , \new_[36199]_ , \new_[36202]_ ,
    \new_[36203]_ , \new_[36204]_ , \new_[36208]_ , \new_[36209]_ ,
    \new_[36213]_ , \new_[36214]_ , \new_[36215]_ , \new_[36219]_ ,
    \new_[36220]_ , \new_[36223]_ , \new_[36226]_ , \new_[36227]_ ,
    \new_[36228]_ , \new_[36232]_ , \new_[36233]_ , \new_[36237]_ ,
    \new_[36238]_ , \new_[36239]_ , \new_[36243]_ , \new_[36244]_ ,
    \new_[36247]_ , \new_[36250]_ , \new_[36251]_ , \new_[36252]_ ,
    \new_[36256]_ , \new_[36257]_ , \new_[36261]_ , \new_[36262]_ ,
    \new_[36263]_ , \new_[36267]_ , \new_[36268]_ , \new_[36271]_ ,
    \new_[36274]_ , \new_[36275]_ , \new_[36276]_ , \new_[36280]_ ,
    \new_[36281]_ , \new_[36285]_ , \new_[36286]_ , \new_[36287]_ ,
    \new_[36291]_ , \new_[36292]_ , \new_[36295]_ , \new_[36298]_ ,
    \new_[36299]_ , \new_[36300]_ , \new_[36304]_ , \new_[36305]_ ,
    \new_[36309]_ , \new_[36310]_ , \new_[36311]_ , \new_[36315]_ ,
    \new_[36316]_ , \new_[36319]_ , \new_[36322]_ , \new_[36323]_ ,
    \new_[36324]_ , \new_[36328]_ , \new_[36329]_ , \new_[36333]_ ,
    \new_[36334]_ , \new_[36335]_ , \new_[36339]_ , \new_[36340]_ ,
    \new_[36343]_ , \new_[36346]_ , \new_[36347]_ , \new_[36348]_ ,
    \new_[36352]_ , \new_[36353]_ , \new_[36357]_ , \new_[36358]_ ,
    \new_[36359]_ , \new_[36363]_ , \new_[36364]_ , \new_[36367]_ ,
    \new_[36370]_ , \new_[36371]_ , \new_[36372]_ , \new_[36376]_ ,
    \new_[36377]_ , \new_[36381]_ , \new_[36382]_ , \new_[36383]_ ,
    \new_[36387]_ , \new_[36388]_ , \new_[36391]_ , \new_[36394]_ ,
    \new_[36395]_ , \new_[36396]_ , \new_[36400]_ , \new_[36401]_ ,
    \new_[36405]_ , \new_[36406]_ , \new_[36407]_ , \new_[36411]_ ,
    \new_[36412]_ , \new_[36415]_ , \new_[36418]_ , \new_[36419]_ ,
    \new_[36420]_ , \new_[36424]_ , \new_[36425]_ , \new_[36429]_ ,
    \new_[36430]_ , \new_[36431]_ , \new_[36435]_ , \new_[36436]_ ,
    \new_[36439]_ , \new_[36442]_ , \new_[36443]_ , \new_[36444]_ ,
    \new_[36448]_ , \new_[36449]_ , \new_[36453]_ , \new_[36454]_ ,
    \new_[36455]_ , \new_[36459]_ , \new_[36460]_ , \new_[36463]_ ,
    \new_[36466]_ , \new_[36467]_ , \new_[36468]_ , \new_[36472]_ ,
    \new_[36473]_ , \new_[36477]_ , \new_[36478]_ , \new_[36479]_ ,
    \new_[36483]_ , \new_[36484]_ , \new_[36487]_ , \new_[36490]_ ,
    \new_[36491]_ , \new_[36492]_ , \new_[36496]_ , \new_[36497]_ ,
    \new_[36501]_ , \new_[36502]_ , \new_[36503]_ , \new_[36507]_ ,
    \new_[36508]_ , \new_[36511]_ , \new_[36514]_ , \new_[36515]_ ,
    \new_[36516]_ , \new_[36520]_ , \new_[36521]_ , \new_[36525]_ ,
    \new_[36526]_ , \new_[36527]_ , \new_[36531]_ , \new_[36532]_ ,
    \new_[36535]_ , \new_[36538]_ , \new_[36539]_ , \new_[36540]_ ,
    \new_[36544]_ , \new_[36545]_ , \new_[36549]_ , \new_[36550]_ ,
    \new_[36551]_ , \new_[36555]_ , \new_[36556]_ , \new_[36559]_ ,
    \new_[36562]_ , \new_[36563]_ , \new_[36564]_ , \new_[36568]_ ,
    \new_[36569]_ , \new_[36573]_ , \new_[36574]_ , \new_[36575]_ ,
    \new_[36579]_ , \new_[36580]_ , \new_[36583]_ , \new_[36586]_ ,
    \new_[36587]_ , \new_[36588]_ , \new_[36592]_ , \new_[36593]_ ,
    \new_[36597]_ , \new_[36598]_ , \new_[36599]_ , \new_[36603]_ ,
    \new_[36604]_ , \new_[36607]_ , \new_[36610]_ , \new_[36611]_ ,
    \new_[36612]_ , \new_[36616]_ , \new_[36617]_ , \new_[36621]_ ,
    \new_[36622]_ , \new_[36623]_ , \new_[36627]_ , \new_[36628]_ ,
    \new_[36631]_ , \new_[36634]_ , \new_[36635]_ , \new_[36636]_ ,
    \new_[36640]_ , \new_[36641]_ , \new_[36645]_ , \new_[36646]_ ,
    \new_[36647]_ , \new_[36651]_ , \new_[36652]_ , \new_[36655]_ ,
    \new_[36658]_ , \new_[36659]_ , \new_[36660]_ , \new_[36664]_ ,
    \new_[36665]_ , \new_[36669]_ , \new_[36670]_ , \new_[36671]_ ,
    \new_[36675]_ , \new_[36676]_ , \new_[36679]_ , \new_[36682]_ ,
    \new_[36683]_ , \new_[36684]_ , \new_[36688]_ , \new_[36689]_ ,
    \new_[36693]_ , \new_[36694]_ , \new_[36695]_ , \new_[36699]_ ,
    \new_[36700]_ , \new_[36703]_ , \new_[36706]_ , \new_[36707]_ ,
    \new_[36708]_ , \new_[36712]_ , \new_[36713]_ , \new_[36717]_ ,
    \new_[36718]_ , \new_[36719]_ , \new_[36723]_ , \new_[36724]_ ,
    \new_[36727]_ , \new_[36730]_ , \new_[36731]_ , \new_[36732]_ ,
    \new_[36736]_ , \new_[36737]_ , \new_[36741]_ , \new_[36742]_ ,
    \new_[36743]_ , \new_[36747]_ , \new_[36748]_ , \new_[36751]_ ,
    \new_[36754]_ , \new_[36755]_ , \new_[36756]_ , \new_[36760]_ ,
    \new_[36761]_ , \new_[36765]_ , \new_[36766]_ , \new_[36767]_ ,
    \new_[36771]_ , \new_[36772]_ , \new_[36775]_ , \new_[36778]_ ,
    \new_[36779]_ , \new_[36780]_ , \new_[36784]_ , \new_[36785]_ ,
    \new_[36789]_ , \new_[36790]_ , \new_[36791]_ , \new_[36795]_ ,
    \new_[36796]_ , \new_[36799]_ , \new_[36802]_ , \new_[36803]_ ,
    \new_[36804]_ , \new_[36808]_ , \new_[36809]_ , \new_[36813]_ ,
    \new_[36814]_ , \new_[36815]_ , \new_[36819]_ , \new_[36820]_ ,
    \new_[36823]_ , \new_[36826]_ , \new_[36827]_ , \new_[36828]_ ,
    \new_[36832]_ , \new_[36833]_ , \new_[36837]_ , \new_[36838]_ ,
    \new_[36839]_ , \new_[36843]_ , \new_[36844]_ , \new_[36847]_ ,
    \new_[36850]_ , \new_[36851]_ , \new_[36852]_ , \new_[36856]_ ,
    \new_[36857]_ , \new_[36861]_ , \new_[36862]_ , \new_[36863]_ ,
    \new_[36867]_ , \new_[36868]_ , \new_[36871]_ , \new_[36874]_ ,
    \new_[36875]_ , \new_[36876]_ , \new_[36880]_ , \new_[36881]_ ,
    \new_[36885]_ , \new_[36886]_ , \new_[36887]_ , \new_[36891]_ ,
    \new_[36892]_ , \new_[36895]_ , \new_[36898]_ , \new_[36899]_ ,
    \new_[36900]_ , \new_[36904]_ , \new_[36905]_ , \new_[36909]_ ,
    \new_[36910]_ , \new_[36911]_ , \new_[36915]_ , \new_[36916]_ ,
    \new_[36919]_ , \new_[36922]_ , \new_[36923]_ , \new_[36924]_ ,
    \new_[36928]_ , \new_[36929]_ , \new_[36933]_ , \new_[36934]_ ,
    \new_[36935]_ , \new_[36939]_ , \new_[36940]_ , \new_[36943]_ ,
    \new_[36946]_ , \new_[36947]_ , \new_[36948]_ , \new_[36952]_ ,
    \new_[36953]_ , \new_[36957]_ , \new_[36958]_ , \new_[36959]_ ,
    \new_[36963]_ , \new_[36964]_ , \new_[36967]_ , \new_[36970]_ ,
    \new_[36971]_ , \new_[36972]_ , \new_[36976]_ , \new_[36977]_ ,
    \new_[36981]_ , \new_[36982]_ , \new_[36983]_ , \new_[36987]_ ,
    \new_[36988]_ , \new_[36991]_ , \new_[36994]_ , \new_[36995]_ ,
    \new_[36996]_ , \new_[37000]_ , \new_[37001]_ , \new_[37005]_ ,
    \new_[37006]_ , \new_[37007]_ , \new_[37011]_ , \new_[37012]_ ,
    \new_[37015]_ , \new_[37018]_ , \new_[37019]_ , \new_[37020]_ ,
    \new_[37024]_ , \new_[37025]_ , \new_[37029]_ , \new_[37030]_ ,
    \new_[37031]_ , \new_[37035]_ , \new_[37036]_ , \new_[37039]_ ,
    \new_[37042]_ , \new_[37043]_ , \new_[37044]_ , \new_[37048]_ ,
    \new_[37049]_ , \new_[37053]_ , \new_[37054]_ , \new_[37055]_ ,
    \new_[37059]_ , \new_[37060]_ , \new_[37063]_ , \new_[37066]_ ,
    \new_[37067]_ , \new_[37068]_ , \new_[37072]_ , \new_[37073]_ ,
    \new_[37077]_ , \new_[37078]_ , \new_[37079]_ , \new_[37083]_ ,
    \new_[37084]_ , \new_[37087]_ , \new_[37090]_ , \new_[37091]_ ,
    \new_[37092]_ , \new_[37096]_ , \new_[37097]_ , \new_[37101]_ ,
    \new_[37102]_ , \new_[37103]_ , \new_[37107]_ , \new_[37108]_ ,
    \new_[37111]_ , \new_[37114]_ , \new_[37115]_ , \new_[37116]_ ,
    \new_[37120]_ , \new_[37121]_ , \new_[37125]_ , \new_[37126]_ ,
    \new_[37127]_ , \new_[37131]_ , \new_[37132]_ , \new_[37135]_ ,
    \new_[37138]_ , \new_[37139]_ , \new_[37140]_ , \new_[37144]_ ,
    \new_[37145]_ , \new_[37149]_ , \new_[37150]_ , \new_[37151]_ ,
    \new_[37155]_ , \new_[37156]_ , \new_[37159]_ , \new_[37162]_ ,
    \new_[37163]_ , \new_[37164]_ , \new_[37168]_ , \new_[37169]_ ,
    \new_[37173]_ , \new_[37174]_ , \new_[37175]_ , \new_[37179]_ ,
    \new_[37180]_ , \new_[37183]_ , \new_[37186]_ , \new_[37187]_ ,
    \new_[37188]_ , \new_[37192]_ , \new_[37193]_ , \new_[37197]_ ,
    \new_[37198]_ , \new_[37199]_ , \new_[37203]_ , \new_[37204]_ ,
    \new_[37207]_ , \new_[37210]_ , \new_[37211]_ , \new_[37212]_ ,
    \new_[37216]_ , \new_[37217]_ , \new_[37221]_ , \new_[37222]_ ,
    \new_[37223]_ , \new_[37227]_ , \new_[37228]_ , \new_[37231]_ ,
    \new_[37234]_ , \new_[37235]_ , \new_[37236]_ , \new_[37240]_ ,
    \new_[37241]_ , \new_[37245]_ , \new_[37246]_ , \new_[37247]_ ,
    \new_[37251]_ , \new_[37252]_ , \new_[37255]_ , \new_[37258]_ ,
    \new_[37259]_ , \new_[37260]_ , \new_[37264]_ , \new_[37265]_ ,
    \new_[37269]_ , \new_[37270]_ , \new_[37271]_ , \new_[37275]_ ,
    \new_[37276]_ , \new_[37279]_ , \new_[37282]_ , \new_[37283]_ ,
    \new_[37284]_ , \new_[37288]_ , \new_[37289]_ , \new_[37293]_ ,
    \new_[37294]_ , \new_[37295]_ , \new_[37299]_ , \new_[37300]_ ,
    \new_[37303]_ , \new_[37306]_ , \new_[37307]_ , \new_[37308]_ ,
    \new_[37312]_ , \new_[37313]_ , \new_[37317]_ , \new_[37318]_ ,
    \new_[37319]_ , \new_[37323]_ , \new_[37324]_ , \new_[37327]_ ,
    \new_[37330]_ , \new_[37331]_ , \new_[37332]_ , \new_[37336]_ ,
    \new_[37337]_ , \new_[37341]_ , \new_[37342]_ , \new_[37343]_ ,
    \new_[37347]_ , \new_[37348]_ , \new_[37351]_ , \new_[37354]_ ,
    \new_[37355]_ , \new_[37356]_ , \new_[37360]_ , \new_[37361]_ ,
    \new_[37365]_ , \new_[37366]_ , \new_[37367]_ , \new_[37371]_ ,
    \new_[37372]_ , \new_[37375]_ , \new_[37378]_ , \new_[37379]_ ,
    \new_[37380]_ , \new_[37384]_ , \new_[37385]_ , \new_[37389]_ ,
    \new_[37390]_ , \new_[37391]_ , \new_[37395]_ , \new_[37396]_ ,
    \new_[37399]_ , \new_[37402]_ , \new_[37403]_ , \new_[37404]_ ,
    \new_[37408]_ , \new_[37409]_ , \new_[37413]_ , \new_[37414]_ ,
    \new_[37415]_ , \new_[37419]_ , \new_[37420]_ , \new_[37423]_ ,
    \new_[37426]_ , \new_[37427]_ , \new_[37428]_ , \new_[37432]_ ,
    \new_[37433]_ , \new_[37437]_ , \new_[37438]_ , \new_[37439]_ ,
    \new_[37443]_ , \new_[37444]_ , \new_[37447]_ , \new_[37450]_ ,
    \new_[37451]_ , \new_[37452]_ , \new_[37456]_ , \new_[37457]_ ,
    \new_[37461]_ , \new_[37462]_ , \new_[37463]_ , \new_[37467]_ ,
    \new_[37468]_ , \new_[37471]_ , \new_[37474]_ , \new_[37475]_ ,
    \new_[37476]_ , \new_[37480]_ , \new_[37481]_ , \new_[37485]_ ,
    \new_[37486]_ , \new_[37487]_ , \new_[37491]_ , \new_[37492]_ ,
    \new_[37495]_ , \new_[37498]_ , \new_[37499]_ , \new_[37500]_ ,
    \new_[37504]_ , \new_[37505]_ , \new_[37509]_ , \new_[37510]_ ,
    \new_[37511]_ , \new_[37515]_ , \new_[37516]_ , \new_[37519]_ ,
    \new_[37522]_ , \new_[37523]_ , \new_[37524]_ , \new_[37528]_ ,
    \new_[37529]_ , \new_[37533]_ , \new_[37534]_ , \new_[37535]_ ,
    \new_[37539]_ , \new_[37540]_ , \new_[37543]_ , \new_[37546]_ ,
    \new_[37547]_ , \new_[37548]_ , \new_[37552]_ , \new_[37553]_ ,
    \new_[37557]_ , \new_[37558]_ , \new_[37559]_ , \new_[37563]_ ,
    \new_[37564]_ , \new_[37567]_ , \new_[37570]_ , \new_[37571]_ ,
    \new_[37572]_ , \new_[37576]_ , \new_[37577]_ , \new_[37581]_ ,
    \new_[37582]_ , \new_[37583]_ , \new_[37587]_ , \new_[37588]_ ,
    \new_[37591]_ , \new_[37594]_ , \new_[37595]_ , \new_[37596]_ ,
    \new_[37600]_ , \new_[37601]_ , \new_[37605]_ , \new_[37606]_ ,
    \new_[37607]_ , \new_[37611]_ , \new_[37612]_ , \new_[37615]_ ,
    \new_[37618]_ , \new_[37619]_ , \new_[37620]_ , \new_[37624]_ ,
    \new_[37625]_ , \new_[37629]_ , \new_[37630]_ , \new_[37631]_ ,
    \new_[37635]_ , \new_[37636]_ , \new_[37639]_ , \new_[37642]_ ,
    \new_[37643]_ , \new_[37644]_ , \new_[37648]_ , \new_[37649]_ ,
    \new_[37653]_ , \new_[37654]_ , \new_[37655]_ , \new_[37659]_ ,
    \new_[37660]_ , \new_[37663]_ , \new_[37666]_ , \new_[37667]_ ,
    \new_[37668]_ , \new_[37672]_ , \new_[37673]_ , \new_[37677]_ ,
    \new_[37678]_ , \new_[37679]_ , \new_[37683]_ , \new_[37684]_ ,
    \new_[37687]_ , \new_[37690]_ , \new_[37691]_ , \new_[37692]_ ,
    \new_[37696]_ , \new_[37697]_ , \new_[37701]_ , \new_[37702]_ ,
    \new_[37703]_ , \new_[37707]_ , \new_[37708]_ , \new_[37711]_ ,
    \new_[37714]_ , \new_[37715]_ , \new_[37716]_ , \new_[37720]_ ,
    \new_[37721]_ , \new_[37725]_ , \new_[37726]_ , \new_[37727]_ ,
    \new_[37731]_ , \new_[37732]_ , \new_[37735]_ , \new_[37738]_ ,
    \new_[37739]_ , \new_[37740]_ , \new_[37744]_ , \new_[37745]_ ,
    \new_[37749]_ , \new_[37750]_ , \new_[37751]_ , \new_[37755]_ ,
    \new_[37756]_ , \new_[37759]_ , \new_[37762]_ , \new_[37763]_ ,
    \new_[37764]_ , \new_[37768]_ , \new_[37769]_ , \new_[37773]_ ,
    \new_[37774]_ , \new_[37775]_ , \new_[37779]_ , \new_[37780]_ ,
    \new_[37783]_ , \new_[37786]_ , \new_[37787]_ , \new_[37788]_ ,
    \new_[37792]_ , \new_[37793]_ , \new_[37797]_ , \new_[37798]_ ,
    \new_[37799]_ , \new_[37803]_ , \new_[37804]_ , \new_[37807]_ ,
    \new_[37810]_ , \new_[37811]_ , \new_[37812]_ , \new_[37816]_ ,
    \new_[37817]_ , \new_[37821]_ , \new_[37822]_ , \new_[37823]_ ,
    \new_[37827]_ , \new_[37828]_ , \new_[37831]_ , \new_[37834]_ ,
    \new_[37835]_ , \new_[37836]_ , \new_[37840]_ , \new_[37841]_ ,
    \new_[37845]_ , \new_[37846]_ , \new_[37847]_ , \new_[37851]_ ,
    \new_[37852]_ , \new_[37855]_ , \new_[37858]_ , \new_[37859]_ ,
    \new_[37860]_ , \new_[37864]_ , \new_[37865]_ , \new_[37869]_ ,
    \new_[37870]_ , \new_[37871]_ , \new_[37875]_ , \new_[37876]_ ,
    \new_[37879]_ , \new_[37882]_ , \new_[37883]_ , \new_[37884]_ ,
    \new_[37888]_ , \new_[37889]_ , \new_[37893]_ , \new_[37894]_ ,
    \new_[37895]_ , \new_[37899]_ , \new_[37900]_ , \new_[37903]_ ,
    \new_[37906]_ , \new_[37907]_ , \new_[37908]_ , \new_[37912]_ ,
    \new_[37913]_ , \new_[37917]_ , \new_[37918]_ , \new_[37919]_ ,
    \new_[37923]_ , \new_[37924]_ , \new_[37927]_ , \new_[37930]_ ,
    \new_[37931]_ , \new_[37932]_ , \new_[37936]_ , \new_[37937]_ ,
    \new_[37941]_ , \new_[37942]_ , \new_[37943]_ , \new_[37947]_ ,
    \new_[37948]_ , \new_[37951]_ , \new_[37954]_ , \new_[37955]_ ,
    \new_[37956]_ , \new_[37960]_ , \new_[37961]_ , \new_[37965]_ ,
    \new_[37966]_ , \new_[37967]_ , \new_[37971]_ , \new_[37972]_ ,
    \new_[37975]_ , \new_[37978]_ , \new_[37979]_ , \new_[37980]_ ,
    \new_[37984]_ , \new_[37985]_ , \new_[37989]_ , \new_[37990]_ ,
    \new_[37991]_ , \new_[37995]_ , \new_[37996]_ , \new_[37999]_ ,
    \new_[38002]_ , \new_[38003]_ , \new_[38004]_ , \new_[38008]_ ,
    \new_[38009]_ , \new_[38013]_ , \new_[38014]_ , \new_[38015]_ ,
    \new_[38019]_ , \new_[38020]_ , \new_[38023]_ , \new_[38026]_ ,
    \new_[38027]_ , \new_[38028]_ , \new_[38032]_ , \new_[38033]_ ,
    \new_[38037]_ , \new_[38038]_ , \new_[38039]_ , \new_[38043]_ ,
    \new_[38044]_ , \new_[38047]_ , \new_[38050]_ , \new_[38051]_ ,
    \new_[38052]_ , \new_[38056]_ , \new_[38057]_ , \new_[38061]_ ,
    \new_[38062]_ , \new_[38063]_ , \new_[38067]_ , \new_[38068]_ ,
    \new_[38071]_ , \new_[38074]_ , \new_[38075]_ , \new_[38076]_ ,
    \new_[38080]_ , \new_[38081]_ , \new_[38085]_ , \new_[38086]_ ,
    \new_[38087]_ , \new_[38091]_ , \new_[38092]_ , \new_[38095]_ ,
    \new_[38098]_ , \new_[38099]_ , \new_[38100]_ , \new_[38104]_ ,
    \new_[38105]_ , \new_[38109]_ , \new_[38110]_ , \new_[38111]_ ,
    \new_[38115]_ , \new_[38116]_ , \new_[38119]_ , \new_[38122]_ ,
    \new_[38123]_ , \new_[38124]_ , \new_[38128]_ , \new_[38129]_ ,
    \new_[38133]_ , \new_[38134]_ , \new_[38135]_ , \new_[38139]_ ,
    \new_[38140]_ , \new_[38143]_ , \new_[38146]_ , \new_[38147]_ ,
    \new_[38148]_ , \new_[38152]_ , \new_[38153]_ , \new_[38157]_ ,
    \new_[38158]_ , \new_[38159]_ , \new_[38163]_ , \new_[38164]_ ,
    \new_[38167]_ , \new_[38170]_ , \new_[38171]_ , \new_[38172]_ ,
    \new_[38176]_ , \new_[38177]_ , \new_[38181]_ , \new_[38182]_ ,
    \new_[38183]_ , \new_[38187]_ , \new_[38188]_ , \new_[38191]_ ,
    \new_[38194]_ , \new_[38195]_ , \new_[38196]_ , \new_[38200]_ ,
    \new_[38201]_ , \new_[38205]_ , \new_[38206]_ , \new_[38207]_ ,
    \new_[38211]_ , \new_[38212]_ , \new_[38215]_ , \new_[38218]_ ,
    \new_[38219]_ , \new_[38220]_ , \new_[38224]_ , \new_[38225]_ ,
    \new_[38229]_ , \new_[38230]_ , \new_[38231]_ , \new_[38235]_ ,
    \new_[38236]_ , \new_[38239]_ , \new_[38242]_ , \new_[38243]_ ,
    \new_[38244]_ , \new_[38248]_ , \new_[38249]_ , \new_[38253]_ ,
    \new_[38254]_ , \new_[38255]_ , \new_[38259]_ , \new_[38260]_ ,
    \new_[38263]_ , \new_[38266]_ , \new_[38267]_ , \new_[38268]_ ,
    \new_[38272]_ , \new_[38273]_ , \new_[38277]_ , \new_[38278]_ ,
    \new_[38279]_ , \new_[38283]_ , \new_[38284]_ , \new_[38287]_ ,
    \new_[38290]_ , \new_[38291]_ , \new_[38292]_ , \new_[38296]_ ,
    \new_[38297]_ , \new_[38301]_ , \new_[38302]_ , \new_[38303]_ ,
    \new_[38307]_ , \new_[38308]_ , \new_[38311]_ , \new_[38314]_ ,
    \new_[38315]_ , \new_[38316]_ , \new_[38320]_ , \new_[38321]_ ,
    \new_[38325]_ , \new_[38326]_ , \new_[38327]_ , \new_[38331]_ ,
    \new_[38332]_ , \new_[38335]_ , \new_[38338]_ , \new_[38339]_ ,
    \new_[38340]_ , \new_[38344]_ , \new_[38345]_ , \new_[38349]_ ,
    \new_[38350]_ , \new_[38351]_ , \new_[38355]_ , \new_[38356]_ ,
    \new_[38359]_ , \new_[38362]_ , \new_[38363]_ , \new_[38364]_ ,
    \new_[38368]_ , \new_[38369]_ , \new_[38373]_ , \new_[38374]_ ,
    \new_[38375]_ , \new_[38379]_ , \new_[38380]_ , \new_[38383]_ ,
    \new_[38386]_ , \new_[38387]_ , \new_[38388]_ , \new_[38392]_ ,
    \new_[38393]_ , \new_[38397]_ , \new_[38398]_ , \new_[38399]_ ,
    \new_[38403]_ , \new_[38404]_ , \new_[38407]_ , \new_[38410]_ ,
    \new_[38411]_ , \new_[38412]_ , \new_[38416]_ , \new_[38417]_ ,
    \new_[38421]_ , \new_[38422]_ , \new_[38423]_ , \new_[38427]_ ,
    \new_[38428]_ , \new_[38431]_ , \new_[38434]_ , \new_[38435]_ ,
    \new_[38436]_ , \new_[38440]_ , \new_[38441]_ , \new_[38445]_ ,
    \new_[38446]_ , \new_[38447]_ , \new_[38451]_ , \new_[38452]_ ,
    \new_[38455]_ , \new_[38458]_ , \new_[38459]_ , \new_[38460]_ ,
    \new_[38464]_ , \new_[38465]_ , \new_[38469]_ , \new_[38470]_ ,
    \new_[38471]_ , \new_[38475]_ , \new_[38476]_ , \new_[38479]_ ,
    \new_[38482]_ , \new_[38483]_ , \new_[38484]_ , \new_[38488]_ ,
    \new_[38489]_ , \new_[38493]_ , \new_[38494]_ , \new_[38495]_ ,
    \new_[38499]_ , \new_[38500]_ , \new_[38503]_ , \new_[38506]_ ,
    \new_[38507]_ , \new_[38508]_ , \new_[38512]_ , \new_[38513]_ ,
    \new_[38517]_ , \new_[38518]_ , \new_[38519]_ , \new_[38523]_ ,
    \new_[38524]_ , \new_[38527]_ , \new_[38530]_ , \new_[38531]_ ,
    \new_[38532]_ , \new_[38536]_ , \new_[38537]_ , \new_[38541]_ ,
    \new_[38542]_ , \new_[38543]_ , \new_[38547]_ , \new_[38548]_ ,
    \new_[38551]_ , \new_[38554]_ , \new_[38555]_ , \new_[38556]_ ,
    \new_[38560]_ , \new_[38561]_ , \new_[38565]_ , \new_[38566]_ ,
    \new_[38567]_ , \new_[38571]_ , \new_[38572]_ , \new_[38575]_ ,
    \new_[38578]_ , \new_[38579]_ , \new_[38580]_ , \new_[38584]_ ,
    \new_[38585]_ , \new_[38589]_ , \new_[38590]_ , \new_[38591]_ ,
    \new_[38595]_ , \new_[38596]_ , \new_[38599]_ , \new_[38602]_ ,
    \new_[38603]_ , \new_[38604]_ , \new_[38608]_ , \new_[38609]_ ,
    \new_[38613]_ , \new_[38614]_ , \new_[38615]_ , \new_[38619]_ ,
    \new_[38620]_ , \new_[38623]_ , \new_[38626]_ , \new_[38627]_ ,
    \new_[38628]_ , \new_[38632]_ , \new_[38633]_ , \new_[38637]_ ,
    \new_[38638]_ , \new_[38639]_ , \new_[38643]_ , \new_[38644]_ ,
    \new_[38647]_ , \new_[38650]_ , \new_[38651]_ , \new_[38652]_ ,
    \new_[38656]_ , \new_[38657]_ , \new_[38661]_ , \new_[38662]_ ,
    \new_[38663]_ , \new_[38667]_ , \new_[38668]_ , \new_[38671]_ ,
    \new_[38674]_ , \new_[38675]_ , \new_[38676]_ , \new_[38680]_ ,
    \new_[38681]_ , \new_[38685]_ , \new_[38686]_ , \new_[38687]_ ,
    \new_[38691]_ , \new_[38692]_ , \new_[38695]_ , \new_[38698]_ ,
    \new_[38699]_ , \new_[38700]_ , \new_[38704]_ , \new_[38705]_ ,
    \new_[38709]_ , \new_[38710]_ , \new_[38711]_ , \new_[38715]_ ,
    \new_[38716]_ , \new_[38719]_ , \new_[38722]_ , \new_[38723]_ ,
    \new_[38724]_ , \new_[38728]_ , \new_[38729]_ , \new_[38733]_ ,
    \new_[38734]_ , \new_[38735]_ , \new_[38739]_ , \new_[38740]_ ,
    \new_[38743]_ , \new_[38746]_ , \new_[38747]_ , \new_[38748]_ ,
    \new_[38752]_ , \new_[38753]_ , \new_[38757]_ , \new_[38758]_ ,
    \new_[38759]_ , \new_[38763]_ , \new_[38764]_ , \new_[38767]_ ,
    \new_[38770]_ , \new_[38771]_ , \new_[38772]_ , \new_[38776]_ ,
    \new_[38777]_ , \new_[38781]_ , \new_[38782]_ , \new_[38783]_ ,
    \new_[38787]_ , \new_[38788]_ , \new_[38791]_ , \new_[38794]_ ,
    \new_[38795]_ , \new_[38796]_ , \new_[38800]_ , \new_[38801]_ ,
    \new_[38805]_ , \new_[38806]_ , \new_[38807]_ , \new_[38811]_ ,
    \new_[38812]_ , \new_[38815]_ , \new_[38818]_ , \new_[38819]_ ,
    \new_[38820]_ , \new_[38824]_ , \new_[38825]_ , \new_[38829]_ ,
    \new_[38830]_ , \new_[38831]_ , \new_[38835]_ , \new_[38836]_ ,
    \new_[38839]_ , \new_[38842]_ , \new_[38843]_ , \new_[38844]_ ,
    \new_[38848]_ , \new_[38849]_ , \new_[38853]_ , \new_[38854]_ ,
    \new_[38855]_ , \new_[38859]_ , \new_[38860]_ , \new_[38863]_ ,
    \new_[38866]_ , \new_[38867]_ , \new_[38868]_ , \new_[38872]_ ,
    \new_[38873]_ , \new_[38877]_ , \new_[38878]_ , \new_[38879]_ ,
    \new_[38883]_ , \new_[38884]_ , \new_[38887]_ , \new_[38890]_ ,
    \new_[38891]_ , \new_[38892]_ , \new_[38896]_ , \new_[38897]_ ,
    \new_[38901]_ , \new_[38902]_ , \new_[38903]_ , \new_[38907]_ ,
    \new_[38908]_ , \new_[38911]_ , \new_[38914]_ , \new_[38915]_ ,
    \new_[38916]_ , \new_[38920]_ , \new_[38921]_ , \new_[38925]_ ,
    \new_[38926]_ , \new_[38927]_ , \new_[38931]_ , \new_[38932]_ ,
    \new_[38935]_ , \new_[38938]_ , \new_[38939]_ , \new_[38940]_ ,
    \new_[38944]_ , \new_[38945]_ , \new_[38949]_ , \new_[38950]_ ,
    \new_[38951]_ , \new_[38955]_ , \new_[38956]_ , \new_[38959]_ ,
    \new_[38962]_ , \new_[38963]_ , \new_[38964]_ , \new_[38968]_ ,
    \new_[38969]_ , \new_[38973]_ , \new_[38974]_ , \new_[38975]_ ,
    \new_[38979]_ , \new_[38980]_ , \new_[38983]_ , \new_[38986]_ ,
    \new_[38987]_ , \new_[38988]_ , \new_[38992]_ , \new_[38993]_ ,
    \new_[38997]_ , \new_[38998]_ , \new_[38999]_ , \new_[39003]_ ,
    \new_[39004]_ , \new_[39007]_ , \new_[39010]_ , \new_[39011]_ ,
    \new_[39012]_ , \new_[39016]_ , \new_[39017]_ , \new_[39021]_ ,
    \new_[39022]_ , \new_[39023]_ , \new_[39027]_ , \new_[39028]_ ,
    \new_[39031]_ , \new_[39034]_ , \new_[39035]_ , \new_[39036]_ ,
    \new_[39040]_ , \new_[39041]_ , \new_[39045]_ , \new_[39046]_ ,
    \new_[39047]_ , \new_[39051]_ , \new_[39052]_ , \new_[39055]_ ,
    \new_[39058]_ , \new_[39059]_ , \new_[39060]_ , \new_[39064]_ ,
    \new_[39065]_ , \new_[39069]_ , \new_[39070]_ , \new_[39071]_ ,
    \new_[39075]_ , \new_[39076]_ , \new_[39079]_ , \new_[39082]_ ,
    \new_[39083]_ , \new_[39084]_ , \new_[39088]_ , \new_[39089]_ ,
    \new_[39093]_ , \new_[39094]_ , \new_[39095]_ , \new_[39099]_ ,
    \new_[39100]_ , \new_[39103]_ , \new_[39106]_ , \new_[39107]_ ,
    \new_[39108]_ , \new_[39112]_ , \new_[39113]_ , \new_[39117]_ ,
    \new_[39118]_ , \new_[39119]_ , \new_[39123]_ , \new_[39124]_ ,
    \new_[39127]_ , \new_[39130]_ , \new_[39131]_ , \new_[39132]_ ,
    \new_[39136]_ , \new_[39137]_ , \new_[39141]_ , \new_[39142]_ ,
    \new_[39143]_ , \new_[39147]_ , \new_[39148]_ , \new_[39151]_ ,
    \new_[39154]_ , \new_[39155]_ , \new_[39156]_ , \new_[39160]_ ,
    \new_[39161]_ , \new_[39165]_ , \new_[39166]_ , \new_[39167]_ ,
    \new_[39171]_ , \new_[39172]_ , \new_[39175]_ , \new_[39178]_ ,
    \new_[39179]_ , \new_[39180]_ , \new_[39184]_ , \new_[39185]_ ,
    \new_[39189]_ , \new_[39190]_ , \new_[39191]_ , \new_[39195]_ ,
    \new_[39196]_ , \new_[39199]_ , \new_[39202]_ , \new_[39203]_ ,
    \new_[39204]_ , \new_[39208]_ , \new_[39209]_ , \new_[39213]_ ,
    \new_[39214]_ , \new_[39215]_ , \new_[39219]_ , \new_[39220]_ ,
    \new_[39223]_ , \new_[39226]_ , \new_[39227]_ , \new_[39228]_ ,
    \new_[39232]_ , \new_[39233]_ , \new_[39237]_ , \new_[39238]_ ,
    \new_[39239]_ , \new_[39243]_ , \new_[39244]_ , \new_[39247]_ ,
    \new_[39250]_ , \new_[39251]_ , \new_[39252]_ , \new_[39256]_ ,
    \new_[39257]_ , \new_[39261]_ , \new_[39262]_ , \new_[39263]_ ,
    \new_[39267]_ , \new_[39268]_ , \new_[39271]_ , \new_[39274]_ ,
    \new_[39275]_ , \new_[39276]_ , \new_[39280]_ , \new_[39281]_ ,
    \new_[39285]_ , \new_[39286]_ , \new_[39287]_ , \new_[39291]_ ,
    \new_[39292]_ , \new_[39295]_ , \new_[39298]_ , \new_[39299]_ ,
    \new_[39300]_ , \new_[39304]_ , \new_[39305]_ , \new_[39309]_ ,
    \new_[39310]_ , \new_[39311]_ , \new_[39315]_ , \new_[39316]_ ,
    \new_[39319]_ , \new_[39322]_ , \new_[39323]_ , \new_[39324]_ ,
    \new_[39328]_ , \new_[39329]_ , \new_[39333]_ , \new_[39334]_ ,
    \new_[39335]_ , \new_[39339]_ , \new_[39340]_ , \new_[39343]_ ,
    \new_[39346]_ , \new_[39347]_ , \new_[39348]_ , \new_[39352]_ ,
    \new_[39353]_ , \new_[39357]_ , \new_[39358]_ , \new_[39359]_ ,
    \new_[39363]_ , \new_[39364]_ , \new_[39367]_ , \new_[39370]_ ,
    \new_[39371]_ , \new_[39372]_ , \new_[39376]_ , \new_[39377]_ ,
    \new_[39381]_ , \new_[39382]_ , \new_[39383]_ , \new_[39387]_ ,
    \new_[39388]_ , \new_[39391]_ , \new_[39394]_ , \new_[39395]_ ,
    \new_[39396]_ , \new_[39400]_ , \new_[39401]_ , \new_[39405]_ ,
    \new_[39406]_ , \new_[39407]_ , \new_[39411]_ , \new_[39412]_ ,
    \new_[39415]_ , \new_[39418]_ , \new_[39419]_ , \new_[39420]_ ,
    \new_[39424]_ , \new_[39425]_ , \new_[39429]_ , \new_[39430]_ ,
    \new_[39431]_ , \new_[39435]_ , \new_[39436]_ , \new_[39439]_ ,
    \new_[39442]_ , \new_[39443]_ , \new_[39444]_ , \new_[39448]_ ,
    \new_[39449]_ , \new_[39453]_ , \new_[39454]_ , \new_[39455]_ ,
    \new_[39459]_ , \new_[39460]_ , \new_[39463]_ , \new_[39466]_ ,
    \new_[39467]_ , \new_[39468]_ , \new_[39472]_ , \new_[39473]_ ,
    \new_[39477]_ , \new_[39478]_ , \new_[39479]_ , \new_[39483]_ ,
    \new_[39484]_ , \new_[39487]_ , \new_[39490]_ , \new_[39491]_ ,
    \new_[39492]_ , \new_[39496]_ , \new_[39497]_ , \new_[39501]_ ,
    \new_[39502]_ , \new_[39503]_ , \new_[39507]_ , \new_[39508]_ ,
    \new_[39511]_ , \new_[39514]_ , \new_[39515]_ , \new_[39516]_ ,
    \new_[39520]_ , \new_[39521]_ , \new_[39525]_ , \new_[39526]_ ,
    \new_[39527]_ , \new_[39531]_ , \new_[39532]_ , \new_[39535]_ ,
    \new_[39538]_ , \new_[39539]_ , \new_[39540]_ , \new_[39544]_ ,
    \new_[39545]_ , \new_[39549]_ , \new_[39550]_ , \new_[39551]_ ,
    \new_[39555]_ , \new_[39556]_ , \new_[39559]_ , \new_[39562]_ ,
    \new_[39563]_ , \new_[39564]_ , \new_[39568]_ , \new_[39569]_ ,
    \new_[39573]_ , \new_[39574]_ , \new_[39575]_ , \new_[39579]_ ,
    \new_[39580]_ , \new_[39583]_ , \new_[39586]_ , \new_[39587]_ ,
    \new_[39588]_ , \new_[39592]_ , \new_[39593]_ , \new_[39597]_ ,
    \new_[39598]_ , \new_[39599]_ , \new_[39603]_ , \new_[39604]_ ,
    \new_[39607]_ , \new_[39610]_ , \new_[39611]_ , \new_[39612]_ ,
    \new_[39616]_ , \new_[39617]_ , \new_[39621]_ , \new_[39622]_ ,
    \new_[39623]_ , \new_[39627]_ , \new_[39628]_ , \new_[39631]_ ,
    \new_[39634]_ , \new_[39635]_ , \new_[39636]_ , \new_[39640]_ ,
    \new_[39641]_ , \new_[39645]_ , \new_[39646]_ , \new_[39647]_ ,
    \new_[39651]_ , \new_[39652]_ , \new_[39655]_ , \new_[39658]_ ,
    \new_[39659]_ , \new_[39660]_ , \new_[39664]_ , \new_[39665]_ ,
    \new_[39669]_ , \new_[39670]_ , \new_[39671]_ , \new_[39675]_ ,
    \new_[39676]_ , \new_[39679]_ , \new_[39682]_ , \new_[39683]_ ,
    \new_[39684]_ , \new_[39688]_ , \new_[39689]_ , \new_[39693]_ ,
    \new_[39694]_ , \new_[39695]_ , \new_[39699]_ , \new_[39700]_ ,
    \new_[39703]_ , \new_[39706]_ , \new_[39707]_ , \new_[39708]_ ,
    \new_[39712]_ , \new_[39713]_ , \new_[39717]_ , \new_[39718]_ ,
    \new_[39719]_ , \new_[39723]_ , \new_[39724]_ , \new_[39727]_ ,
    \new_[39730]_ , \new_[39731]_ , \new_[39732]_ , \new_[39736]_ ,
    \new_[39737]_ , \new_[39741]_ , \new_[39742]_ , \new_[39743]_ ,
    \new_[39747]_ , \new_[39748]_ , \new_[39751]_ , \new_[39754]_ ,
    \new_[39755]_ , \new_[39756]_ , \new_[39760]_ , \new_[39761]_ ,
    \new_[39765]_ , \new_[39766]_ , \new_[39767]_ , \new_[39771]_ ,
    \new_[39772]_ , \new_[39775]_ , \new_[39778]_ , \new_[39779]_ ,
    \new_[39780]_ , \new_[39784]_ , \new_[39785]_ , \new_[39789]_ ,
    \new_[39790]_ , \new_[39791]_ , \new_[39795]_ , \new_[39796]_ ,
    \new_[39799]_ , \new_[39802]_ , \new_[39803]_ , \new_[39804]_ ,
    \new_[39808]_ , \new_[39809]_ , \new_[39813]_ , \new_[39814]_ ,
    \new_[39815]_ , \new_[39819]_ , \new_[39820]_ , \new_[39823]_ ,
    \new_[39826]_ , \new_[39827]_ , \new_[39828]_ , \new_[39832]_ ,
    \new_[39833]_ , \new_[39837]_ , \new_[39838]_ , \new_[39839]_ ,
    \new_[39843]_ , \new_[39844]_ , \new_[39847]_ , \new_[39850]_ ,
    \new_[39851]_ , \new_[39852]_ , \new_[39856]_ , \new_[39857]_ ,
    \new_[39861]_ , \new_[39862]_ , \new_[39863]_ , \new_[39867]_ ,
    \new_[39868]_ , \new_[39871]_ , \new_[39874]_ , \new_[39875]_ ,
    \new_[39876]_ , \new_[39880]_ , \new_[39881]_ , \new_[39885]_ ,
    \new_[39886]_ , \new_[39887]_ , \new_[39891]_ , \new_[39892]_ ,
    \new_[39895]_ , \new_[39898]_ , \new_[39899]_ , \new_[39900]_ ,
    \new_[39904]_ , \new_[39905]_ , \new_[39909]_ , \new_[39910]_ ,
    \new_[39911]_ , \new_[39915]_ , \new_[39916]_ , \new_[39919]_ ,
    \new_[39922]_ , \new_[39923]_ , \new_[39924]_ , \new_[39928]_ ,
    \new_[39929]_ , \new_[39933]_ , \new_[39934]_ , \new_[39935]_ ,
    \new_[39939]_ , \new_[39940]_ , \new_[39943]_ , \new_[39946]_ ,
    \new_[39947]_ , \new_[39948]_ , \new_[39952]_ , \new_[39953]_ ,
    \new_[39957]_ , \new_[39958]_ , \new_[39959]_ , \new_[39963]_ ,
    \new_[39964]_ , \new_[39967]_ , \new_[39970]_ , \new_[39971]_ ,
    \new_[39972]_ , \new_[39976]_ , \new_[39977]_ , \new_[39981]_ ,
    \new_[39982]_ , \new_[39983]_ , \new_[39987]_ , \new_[39988]_ ,
    \new_[39991]_ , \new_[39994]_ , \new_[39995]_ , \new_[39996]_ ,
    \new_[40000]_ , \new_[40001]_ , \new_[40005]_ , \new_[40006]_ ,
    \new_[40007]_ , \new_[40011]_ , \new_[40012]_ , \new_[40015]_ ,
    \new_[40018]_ , \new_[40019]_ , \new_[40020]_ , \new_[40024]_ ,
    \new_[40025]_ , \new_[40029]_ , \new_[40030]_ , \new_[40031]_ ,
    \new_[40035]_ , \new_[40036]_ , \new_[40039]_ , \new_[40042]_ ,
    \new_[40043]_ , \new_[40044]_ , \new_[40048]_ , \new_[40049]_ ,
    \new_[40053]_ , \new_[40054]_ , \new_[40055]_ , \new_[40059]_ ,
    \new_[40060]_ , \new_[40063]_ , \new_[40066]_ , \new_[40067]_ ,
    \new_[40068]_ , \new_[40072]_ , \new_[40073]_ , \new_[40077]_ ,
    \new_[40078]_ , \new_[40079]_ , \new_[40083]_ , \new_[40084]_ ,
    \new_[40087]_ , \new_[40090]_ , \new_[40091]_ , \new_[40092]_ ,
    \new_[40096]_ , \new_[40097]_ , \new_[40101]_ , \new_[40102]_ ,
    \new_[40103]_ , \new_[40107]_ , \new_[40108]_ , \new_[40111]_ ,
    \new_[40114]_ , \new_[40115]_ , \new_[40116]_ , \new_[40120]_ ,
    \new_[40121]_ , \new_[40125]_ , \new_[40126]_ , \new_[40127]_ ,
    \new_[40131]_ , \new_[40132]_ , \new_[40135]_ , \new_[40138]_ ,
    \new_[40139]_ , \new_[40140]_ , \new_[40144]_ , \new_[40145]_ ,
    \new_[40149]_ , \new_[40150]_ , \new_[40151]_ , \new_[40155]_ ,
    \new_[40156]_ , \new_[40159]_ , \new_[40162]_ , \new_[40163]_ ,
    \new_[40164]_ , \new_[40168]_ , \new_[40169]_ , \new_[40173]_ ,
    \new_[40174]_ , \new_[40175]_ , \new_[40179]_ , \new_[40180]_ ,
    \new_[40183]_ , \new_[40186]_ , \new_[40187]_ , \new_[40188]_ ,
    \new_[40192]_ , \new_[40193]_ , \new_[40197]_ , \new_[40198]_ ,
    \new_[40199]_ , \new_[40203]_ , \new_[40204]_ , \new_[40207]_ ,
    \new_[40210]_ , \new_[40211]_ , \new_[40212]_ , \new_[40216]_ ,
    \new_[40217]_ , \new_[40221]_ , \new_[40222]_ , \new_[40223]_ ,
    \new_[40227]_ , \new_[40228]_ , \new_[40231]_ , \new_[40234]_ ,
    \new_[40235]_ , \new_[40236]_ , \new_[40240]_ , \new_[40241]_ ,
    \new_[40245]_ , \new_[40246]_ , \new_[40247]_ , \new_[40251]_ ,
    \new_[40252]_ , \new_[40255]_ , \new_[40258]_ , \new_[40259]_ ,
    \new_[40260]_ , \new_[40264]_ , \new_[40265]_ , \new_[40269]_ ,
    \new_[40270]_ , \new_[40271]_ , \new_[40275]_ , \new_[40276]_ ,
    \new_[40279]_ , \new_[40282]_ , \new_[40283]_ , \new_[40284]_ ,
    \new_[40288]_ , \new_[40289]_ , \new_[40293]_ , \new_[40294]_ ,
    \new_[40295]_ , \new_[40299]_ , \new_[40300]_ , \new_[40303]_ ,
    \new_[40306]_ , \new_[40307]_ , \new_[40308]_ , \new_[40312]_ ,
    \new_[40313]_ , \new_[40317]_ , \new_[40318]_ , \new_[40319]_ ,
    \new_[40323]_ , \new_[40324]_ , \new_[40327]_ , \new_[40330]_ ,
    \new_[40331]_ , \new_[40332]_ , \new_[40336]_ , \new_[40337]_ ,
    \new_[40341]_ , \new_[40342]_ , \new_[40343]_ , \new_[40347]_ ,
    \new_[40348]_ , \new_[40351]_ , \new_[40354]_ , \new_[40355]_ ,
    \new_[40356]_ , \new_[40360]_ , \new_[40361]_ , \new_[40365]_ ,
    \new_[40366]_ , \new_[40367]_ , \new_[40371]_ , \new_[40372]_ ,
    \new_[40375]_ , \new_[40378]_ , \new_[40379]_ , \new_[40380]_ ,
    \new_[40384]_ , \new_[40385]_ , \new_[40389]_ , \new_[40390]_ ,
    \new_[40391]_ , \new_[40395]_ , \new_[40396]_ , \new_[40399]_ ,
    \new_[40402]_ , \new_[40403]_ , \new_[40404]_ , \new_[40408]_ ,
    \new_[40409]_ , \new_[40413]_ , \new_[40414]_ , \new_[40415]_ ,
    \new_[40419]_ , \new_[40420]_ , \new_[40423]_ , \new_[40426]_ ,
    \new_[40427]_ , \new_[40428]_ , \new_[40432]_ , \new_[40433]_ ,
    \new_[40437]_ , \new_[40438]_ , \new_[40439]_ , \new_[40443]_ ,
    \new_[40444]_ , \new_[40447]_ , \new_[40450]_ , \new_[40451]_ ,
    \new_[40452]_ , \new_[40456]_ , \new_[40457]_ , \new_[40461]_ ,
    \new_[40462]_ , \new_[40463]_ , \new_[40467]_ , \new_[40468]_ ,
    \new_[40471]_ , \new_[40474]_ , \new_[40475]_ , \new_[40476]_ ,
    \new_[40480]_ , \new_[40481]_ , \new_[40485]_ , \new_[40486]_ ,
    \new_[40487]_ , \new_[40491]_ , \new_[40492]_ , \new_[40495]_ ,
    \new_[40498]_ , \new_[40499]_ , \new_[40500]_ , \new_[40504]_ ,
    \new_[40505]_ , \new_[40509]_ , \new_[40510]_ , \new_[40511]_ ,
    \new_[40515]_ , \new_[40516]_ , \new_[40519]_ , \new_[40522]_ ,
    \new_[40523]_ , \new_[40524]_ , \new_[40528]_ , \new_[40529]_ ,
    \new_[40533]_ , \new_[40534]_ , \new_[40535]_ , \new_[40539]_ ,
    \new_[40540]_ , \new_[40543]_ , \new_[40546]_ , \new_[40547]_ ,
    \new_[40548]_ , \new_[40552]_ , \new_[40553]_ , \new_[40557]_ ,
    \new_[40558]_ , \new_[40559]_ , \new_[40563]_ , \new_[40564]_ ,
    \new_[40567]_ , \new_[40570]_ , \new_[40571]_ , \new_[40572]_ ,
    \new_[40576]_ , \new_[40577]_ , \new_[40581]_ , \new_[40582]_ ,
    \new_[40583]_ , \new_[40587]_ , \new_[40588]_ , \new_[40591]_ ,
    \new_[40594]_ , \new_[40595]_ , \new_[40596]_ , \new_[40600]_ ,
    \new_[40601]_ , \new_[40605]_ , \new_[40606]_ , \new_[40607]_ ,
    \new_[40611]_ , \new_[40612]_ , \new_[40615]_ , \new_[40618]_ ,
    \new_[40619]_ , \new_[40620]_ , \new_[40624]_ , \new_[40625]_ ,
    \new_[40629]_ , \new_[40630]_ , \new_[40631]_ , \new_[40635]_ ,
    \new_[40636]_ , \new_[40639]_ , \new_[40642]_ , \new_[40643]_ ,
    \new_[40644]_ , \new_[40648]_ , \new_[40649]_ , \new_[40653]_ ,
    \new_[40654]_ , \new_[40655]_ , \new_[40659]_ , \new_[40660]_ ,
    \new_[40663]_ , \new_[40666]_ , \new_[40667]_ , \new_[40668]_ ,
    \new_[40672]_ , \new_[40673]_ , \new_[40677]_ , \new_[40678]_ ,
    \new_[40679]_ , \new_[40683]_ , \new_[40684]_ , \new_[40687]_ ,
    \new_[40690]_ , \new_[40691]_ , \new_[40692]_ , \new_[40696]_ ,
    \new_[40697]_ , \new_[40701]_ , \new_[40702]_ , \new_[40703]_ ,
    \new_[40707]_ , \new_[40708]_ , \new_[40711]_ , \new_[40714]_ ,
    \new_[40715]_ , \new_[40716]_ , \new_[40720]_ , \new_[40721]_ ,
    \new_[40725]_ , \new_[40726]_ , \new_[40727]_ , \new_[40731]_ ,
    \new_[40732]_ , \new_[40735]_ , \new_[40738]_ , \new_[40739]_ ,
    \new_[40740]_ , \new_[40744]_ , \new_[40745]_ , \new_[40749]_ ,
    \new_[40750]_ , \new_[40751]_ , \new_[40755]_ , \new_[40756]_ ,
    \new_[40759]_ , \new_[40762]_ , \new_[40763]_ , \new_[40764]_ ,
    \new_[40768]_ , \new_[40769]_ , \new_[40773]_ , \new_[40774]_ ,
    \new_[40775]_ , \new_[40779]_ , \new_[40780]_ , \new_[40783]_ ,
    \new_[40786]_ , \new_[40787]_ , \new_[40788]_ , \new_[40792]_ ,
    \new_[40793]_ , \new_[40797]_ , \new_[40798]_ , \new_[40799]_ ,
    \new_[40803]_ , \new_[40804]_ , \new_[40807]_ , \new_[40810]_ ,
    \new_[40811]_ , \new_[40812]_ , \new_[40816]_ , \new_[40817]_ ,
    \new_[40821]_ , \new_[40822]_ , \new_[40823]_ , \new_[40827]_ ,
    \new_[40828]_ , \new_[40831]_ , \new_[40834]_ , \new_[40835]_ ,
    \new_[40836]_ , \new_[40840]_ , \new_[40841]_ , \new_[40845]_ ,
    \new_[40846]_ , \new_[40847]_ , \new_[40851]_ , \new_[40852]_ ,
    \new_[40855]_ , \new_[40858]_ , \new_[40859]_ , \new_[40860]_ ,
    \new_[40864]_ , \new_[40865]_ , \new_[40869]_ , \new_[40870]_ ,
    \new_[40871]_ , \new_[40875]_ , \new_[40876]_ , \new_[40879]_ ,
    \new_[40882]_ , \new_[40883]_ , \new_[40884]_ , \new_[40888]_ ,
    \new_[40889]_ , \new_[40893]_ , \new_[40894]_ , \new_[40895]_ ,
    \new_[40899]_ , \new_[40900]_ , \new_[40903]_ , \new_[40906]_ ,
    \new_[40907]_ , \new_[40908]_ , \new_[40912]_ , \new_[40913]_ ,
    \new_[40917]_ , \new_[40918]_ , \new_[40919]_ , \new_[40923]_ ,
    \new_[40924]_ , \new_[40927]_ , \new_[40930]_ , \new_[40931]_ ,
    \new_[40932]_ , \new_[40936]_ , \new_[40937]_ , \new_[40941]_ ,
    \new_[40942]_ , \new_[40943]_ , \new_[40947]_ , \new_[40948]_ ,
    \new_[40951]_ , \new_[40954]_ , \new_[40955]_ , \new_[40956]_ ,
    \new_[40960]_ , \new_[40961]_ , \new_[40965]_ , \new_[40966]_ ,
    \new_[40967]_ , \new_[40971]_ , \new_[40972]_ , \new_[40975]_ ,
    \new_[40978]_ , \new_[40979]_ , \new_[40980]_ , \new_[40984]_ ,
    \new_[40985]_ , \new_[40989]_ , \new_[40990]_ , \new_[40991]_ ,
    \new_[40995]_ , \new_[40996]_ , \new_[40999]_ , \new_[41002]_ ,
    \new_[41003]_ , \new_[41004]_ , \new_[41008]_ , \new_[41009]_ ,
    \new_[41013]_ , \new_[41014]_ , \new_[41015]_ , \new_[41019]_ ,
    \new_[41020]_ , \new_[41023]_ , \new_[41026]_ , \new_[41027]_ ,
    \new_[41028]_ , \new_[41032]_ , \new_[41033]_ , \new_[41037]_ ,
    \new_[41038]_ , \new_[41039]_ , \new_[41043]_ , \new_[41044]_ ,
    \new_[41047]_ , \new_[41050]_ , \new_[41051]_ , \new_[41052]_ ,
    \new_[41056]_ , \new_[41057]_ , \new_[41061]_ , \new_[41062]_ ,
    \new_[41063]_ , \new_[41067]_ , \new_[41068]_ , \new_[41071]_ ,
    \new_[41074]_ , \new_[41075]_ , \new_[41076]_ , \new_[41080]_ ,
    \new_[41081]_ , \new_[41085]_ , \new_[41086]_ , \new_[41087]_ ,
    \new_[41091]_ , \new_[41092]_ , \new_[41095]_ , \new_[41098]_ ,
    \new_[41099]_ , \new_[41100]_ , \new_[41104]_ , \new_[41105]_ ,
    \new_[41109]_ , \new_[41110]_ , \new_[41111]_ , \new_[41115]_ ,
    \new_[41116]_ , \new_[41119]_ , \new_[41122]_ , \new_[41123]_ ,
    \new_[41124]_ , \new_[41128]_ , \new_[41129]_ , \new_[41133]_ ,
    \new_[41134]_ , \new_[41135]_ , \new_[41139]_ , \new_[41140]_ ,
    \new_[41143]_ , \new_[41146]_ , \new_[41147]_ , \new_[41148]_ ,
    \new_[41152]_ , \new_[41153]_ , \new_[41157]_ , \new_[41158]_ ,
    \new_[41159]_ , \new_[41163]_ , \new_[41164]_ , \new_[41167]_ ,
    \new_[41170]_ , \new_[41171]_ , \new_[41172]_ , \new_[41176]_ ,
    \new_[41177]_ , \new_[41181]_ , \new_[41182]_ , \new_[41183]_ ,
    \new_[41187]_ , \new_[41188]_ , \new_[41191]_ , \new_[41194]_ ,
    \new_[41195]_ , \new_[41196]_ , \new_[41200]_ , \new_[41201]_ ,
    \new_[41205]_ , \new_[41206]_ , \new_[41207]_ , \new_[41211]_ ,
    \new_[41212]_ , \new_[41215]_ , \new_[41218]_ , \new_[41219]_ ,
    \new_[41220]_ , \new_[41224]_ , \new_[41225]_ , \new_[41229]_ ,
    \new_[41230]_ , \new_[41231]_ , \new_[41235]_ , \new_[41236]_ ,
    \new_[41239]_ , \new_[41242]_ , \new_[41243]_ , \new_[41244]_ ,
    \new_[41248]_ , \new_[41249]_ , \new_[41253]_ , \new_[41254]_ ,
    \new_[41255]_ , \new_[41259]_ , \new_[41260]_ , \new_[41263]_ ,
    \new_[41266]_ , \new_[41267]_ , \new_[41268]_ , \new_[41272]_ ,
    \new_[41273]_ , \new_[41277]_ , \new_[41278]_ , \new_[41279]_ ,
    \new_[41283]_ , \new_[41284]_ , \new_[41287]_ , \new_[41290]_ ,
    \new_[41291]_ , \new_[41292]_ , \new_[41296]_ , \new_[41297]_ ,
    \new_[41301]_ , \new_[41302]_ , \new_[41303]_ , \new_[41307]_ ,
    \new_[41308]_ , \new_[41311]_ , \new_[41314]_ , \new_[41315]_ ,
    \new_[41316]_ , \new_[41320]_ , \new_[41321]_ , \new_[41325]_ ,
    \new_[41326]_ , \new_[41327]_ , \new_[41331]_ , \new_[41332]_ ,
    \new_[41335]_ , \new_[41338]_ , \new_[41339]_ , \new_[41340]_ ,
    \new_[41344]_ , \new_[41345]_ , \new_[41349]_ , \new_[41350]_ ,
    \new_[41351]_ , \new_[41355]_ , \new_[41356]_ , \new_[41359]_ ,
    \new_[41362]_ , \new_[41363]_ , \new_[41364]_ , \new_[41368]_ ,
    \new_[41369]_ , \new_[41373]_ , \new_[41374]_ , \new_[41375]_ ,
    \new_[41379]_ , \new_[41380]_ , \new_[41383]_ , \new_[41386]_ ,
    \new_[41387]_ , \new_[41388]_ , \new_[41392]_ , \new_[41393]_ ,
    \new_[41397]_ , \new_[41398]_ , \new_[41399]_ , \new_[41403]_ ,
    \new_[41404]_ , \new_[41407]_ , \new_[41410]_ , \new_[41411]_ ,
    \new_[41412]_ , \new_[41416]_ , \new_[41417]_ , \new_[41421]_ ,
    \new_[41422]_ , \new_[41423]_ , \new_[41427]_ , \new_[41428]_ ,
    \new_[41431]_ , \new_[41434]_ , \new_[41435]_ , \new_[41436]_ ,
    \new_[41440]_ , \new_[41441]_ , \new_[41445]_ , \new_[41446]_ ,
    \new_[41447]_ , \new_[41451]_ , \new_[41452]_ , \new_[41455]_ ,
    \new_[41458]_ , \new_[41459]_ , \new_[41460]_ , \new_[41464]_ ,
    \new_[41465]_ , \new_[41469]_ , \new_[41470]_ , \new_[41471]_ ,
    \new_[41475]_ , \new_[41476]_ , \new_[41479]_ , \new_[41482]_ ,
    \new_[41483]_ , \new_[41484]_ , \new_[41488]_ , \new_[41489]_ ,
    \new_[41493]_ , \new_[41494]_ , \new_[41495]_ , \new_[41499]_ ,
    \new_[41500]_ , \new_[41503]_ , \new_[41506]_ , \new_[41507]_ ,
    \new_[41508]_ , \new_[41512]_ , \new_[41513]_ , \new_[41517]_ ,
    \new_[41518]_ , \new_[41519]_ , \new_[41523]_ , \new_[41524]_ ,
    \new_[41527]_ , \new_[41530]_ , \new_[41531]_ , \new_[41532]_ ,
    \new_[41536]_ , \new_[41537]_ , \new_[41541]_ , \new_[41542]_ ,
    \new_[41543]_ , \new_[41547]_ , \new_[41548]_ , \new_[41551]_ ,
    \new_[41554]_ , \new_[41555]_ , \new_[41556]_ , \new_[41560]_ ,
    \new_[41561]_ , \new_[41565]_ , \new_[41566]_ , \new_[41567]_ ,
    \new_[41571]_ , \new_[41572]_ , \new_[41575]_ , \new_[41578]_ ,
    \new_[41579]_ , \new_[41580]_ , \new_[41584]_ , \new_[41585]_ ,
    \new_[41589]_ , \new_[41590]_ , \new_[41591]_ , \new_[41595]_ ,
    \new_[41596]_ , \new_[41599]_ , \new_[41602]_ , \new_[41603]_ ,
    \new_[41604]_ , \new_[41608]_ , \new_[41609]_ , \new_[41613]_ ,
    \new_[41614]_ , \new_[41615]_ , \new_[41619]_ , \new_[41620]_ ,
    \new_[41623]_ , \new_[41626]_ , \new_[41627]_ , \new_[41628]_ ,
    \new_[41632]_ , \new_[41633]_ , \new_[41637]_ , \new_[41638]_ ,
    \new_[41639]_ , \new_[41643]_ , \new_[41644]_ , \new_[41647]_ ,
    \new_[41650]_ , \new_[41651]_ , \new_[41652]_ , \new_[41656]_ ,
    \new_[41657]_ , \new_[41661]_ , \new_[41662]_ , \new_[41663]_ ,
    \new_[41667]_ , \new_[41668]_ , \new_[41671]_ , \new_[41674]_ ,
    \new_[41675]_ , \new_[41676]_ , \new_[41680]_ , \new_[41681]_ ,
    \new_[41685]_ , \new_[41686]_ , \new_[41687]_ , \new_[41691]_ ,
    \new_[41692]_ , \new_[41695]_ , \new_[41698]_ , \new_[41699]_ ,
    \new_[41700]_ , \new_[41704]_ , \new_[41705]_ , \new_[41709]_ ,
    \new_[41710]_ , \new_[41711]_ , \new_[41715]_ , \new_[41716]_ ,
    \new_[41719]_ , \new_[41722]_ , \new_[41723]_ , \new_[41724]_ ,
    \new_[41728]_ , \new_[41729]_ , \new_[41733]_ , \new_[41734]_ ,
    \new_[41735]_ , \new_[41739]_ , \new_[41740]_ , \new_[41743]_ ,
    \new_[41746]_ , \new_[41747]_ , \new_[41748]_ , \new_[41752]_ ,
    \new_[41753]_ , \new_[41757]_ , \new_[41758]_ , \new_[41759]_ ,
    \new_[41763]_ , \new_[41764]_ , \new_[41767]_ , \new_[41770]_ ,
    \new_[41771]_ , \new_[41772]_ , \new_[41776]_ , \new_[41777]_ ,
    \new_[41781]_ , \new_[41782]_ , \new_[41783]_ , \new_[41787]_ ,
    \new_[41788]_ , \new_[41791]_ , \new_[41794]_ , \new_[41795]_ ,
    \new_[41796]_ , \new_[41800]_ , \new_[41801]_ , \new_[41805]_ ,
    \new_[41806]_ , \new_[41807]_ , \new_[41811]_ , \new_[41812]_ ,
    \new_[41815]_ , \new_[41818]_ , \new_[41819]_ , \new_[41820]_ ,
    \new_[41824]_ , \new_[41825]_ , \new_[41829]_ , \new_[41830]_ ,
    \new_[41831]_ , \new_[41835]_ , \new_[41836]_ , \new_[41839]_ ,
    \new_[41842]_ , \new_[41843]_ , \new_[41844]_ , \new_[41848]_ ,
    \new_[41849]_ , \new_[41853]_ , \new_[41854]_ , \new_[41855]_ ,
    \new_[41859]_ , \new_[41860]_ , \new_[41863]_ , \new_[41866]_ ,
    \new_[41867]_ , \new_[41868]_ , \new_[41872]_ , \new_[41873]_ ,
    \new_[41877]_ , \new_[41878]_ , \new_[41879]_ , \new_[41883]_ ,
    \new_[41884]_ , \new_[41887]_ , \new_[41890]_ , \new_[41891]_ ,
    \new_[41892]_ , \new_[41896]_ , \new_[41897]_ , \new_[41901]_ ,
    \new_[41902]_ , \new_[41903]_ , \new_[41907]_ , \new_[41908]_ ,
    \new_[41911]_ , \new_[41914]_ , \new_[41915]_ , \new_[41916]_ ,
    \new_[41920]_ , \new_[41921]_ , \new_[41925]_ , \new_[41926]_ ,
    \new_[41927]_ , \new_[41931]_ , \new_[41932]_ , \new_[41935]_ ,
    \new_[41938]_ , \new_[41939]_ , \new_[41940]_ , \new_[41944]_ ,
    \new_[41945]_ , \new_[41949]_ , \new_[41950]_ , \new_[41951]_ ,
    \new_[41955]_ , \new_[41956]_ , \new_[41959]_ , \new_[41962]_ ,
    \new_[41963]_ , \new_[41964]_ , \new_[41968]_ , \new_[41969]_ ,
    \new_[41973]_ , \new_[41974]_ , \new_[41975]_ , \new_[41979]_ ,
    \new_[41980]_ , \new_[41983]_ , \new_[41986]_ , \new_[41987]_ ,
    \new_[41988]_ , \new_[41992]_ , \new_[41993]_ , \new_[41997]_ ,
    \new_[41998]_ , \new_[41999]_ , \new_[42003]_ , \new_[42004]_ ,
    \new_[42007]_ , \new_[42010]_ , \new_[42011]_ , \new_[42012]_ ,
    \new_[42016]_ , \new_[42017]_ , \new_[42021]_ , \new_[42022]_ ,
    \new_[42023]_ , \new_[42027]_ , \new_[42028]_ , \new_[42031]_ ,
    \new_[42034]_ , \new_[42035]_ , \new_[42036]_ , \new_[42040]_ ,
    \new_[42041]_ , \new_[42045]_ , \new_[42046]_ , \new_[42047]_ ,
    \new_[42051]_ , \new_[42052]_ , \new_[42055]_ , \new_[42058]_ ,
    \new_[42059]_ , \new_[42060]_ , \new_[42064]_ , \new_[42065]_ ,
    \new_[42069]_ , \new_[42070]_ , \new_[42071]_ , \new_[42075]_ ,
    \new_[42076]_ , \new_[42079]_ , \new_[42082]_ , \new_[42083]_ ,
    \new_[42084]_ , \new_[42088]_ , \new_[42089]_ , \new_[42093]_ ,
    \new_[42094]_ , \new_[42095]_ , \new_[42099]_ , \new_[42100]_ ,
    \new_[42103]_ , \new_[42106]_ , \new_[42107]_ , \new_[42108]_ ,
    \new_[42112]_ , \new_[42113]_ , \new_[42117]_ , \new_[42118]_ ,
    \new_[42119]_ , \new_[42123]_ , \new_[42124]_ , \new_[42127]_ ,
    \new_[42130]_ , \new_[42131]_ , \new_[42132]_ , \new_[42136]_ ,
    \new_[42137]_ , \new_[42141]_ , \new_[42142]_ , \new_[42143]_ ,
    \new_[42147]_ , \new_[42148]_ , \new_[42151]_ , \new_[42154]_ ,
    \new_[42155]_ , \new_[42156]_ , \new_[42160]_ , \new_[42161]_ ,
    \new_[42165]_ , \new_[42166]_ , \new_[42167]_ , \new_[42171]_ ,
    \new_[42172]_ , \new_[42175]_ , \new_[42178]_ , \new_[42179]_ ,
    \new_[42180]_ , \new_[42184]_ , \new_[42185]_ , \new_[42189]_ ,
    \new_[42190]_ , \new_[42191]_ , \new_[42195]_ , \new_[42196]_ ,
    \new_[42199]_ , \new_[42202]_ , \new_[42203]_ , \new_[42204]_ ,
    \new_[42208]_ , \new_[42209]_ , \new_[42213]_ , \new_[42214]_ ,
    \new_[42215]_ , \new_[42219]_ , \new_[42220]_ , \new_[42223]_ ,
    \new_[42226]_ , \new_[42227]_ , \new_[42228]_ , \new_[42232]_ ,
    \new_[42233]_ , \new_[42237]_ , \new_[42238]_ , \new_[42239]_ ,
    \new_[42243]_ , \new_[42244]_ , \new_[42247]_ , \new_[42250]_ ,
    \new_[42251]_ , \new_[42252]_ , \new_[42256]_ , \new_[42257]_ ,
    \new_[42261]_ , \new_[42262]_ , \new_[42263]_ , \new_[42267]_ ,
    \new_[42268]_ , \new_[42271]_ , \new_[42274]_ , \new_[42275]_ ,
    \new_[42276]_ , \new_[42280]_ , \new_[42281]_ , \new_[42285]_ ,
    \new_[42286]_ , \new_[42287]_ , \new_[42291]_ , \new_[42292]_ ,
    \new_[42295]_ , \new_[42298]_ , \new_[42299]_ , \new_[42300]_ ,
    \new_[42304]_ , \new_[42305]_ , \new_[42309]_ , \new_[42310]_ ,
    \new_[42311]_ , \new_[42315]_ , \new_[42316]_ , \new_[42319]_ ,
    \new_[42322]_ , \new_[42323]_ , \new_[42324]_ , \new_[42328]_ ,
    \new_[42329]_ , \new_[42333]_ , \new_[42334]_ , \new_[42335]_ ,
    \new_[42339]_ , \new_[42340]_ , \new_[42343]_ , \new_[42346]_ ,
    \new_[42347]_ , \new_[42348]_ , \new_[42352]_ , \new_[42353]_ ,
    \new_[42357]_ , \new_[42358]_ , \new_[42359]_ , \new_[42363]_ ,
    \new_[42364]_ , \new_[42367]_ , \new_[42370]_ , \new_[42371]_ ,
    \new_[42372]_ , \new_[42376]_ , \new_[42377]_ , \new_[42381]_ ,
    \new_[42382]_ , \new_[42383]_ , \new_[42387]_ , \new_[42388]_ ,
    \new_[42391]_ , \new_[42394]_ , \new_[42395]_ , \new_[42396]_ ,
    \new_[42400]_ , \new_[42401]_ , \new_[42405]_ , \new_[42406]_ ,
    \new_[42407]_ , \new_[42411]_ , \new_[42412]_ , \new_[42415]_ ,
    \new_[42418]_ , \new_[42419]_ , \new_[42420]_ , \new_[42424]_ ,
    \new_[42425]_ , \new_[42429]_ , \new_[42430]_ , \new_[42431]_ ,
    \new_[42435]_ , \new_[42436]_ , \new_[42439]_ , \new_[42442]_ ,
    \new_[42443]_ , \new_[42444]_ , \new_[42448]_ , \new_[42449]_ ,
    \new_[42453]_ , \new_[42454]_ , \new_[42455]_ , \new_[42459]_ ,
    \new_[42460]_ , \new_[42463]_ , \new_[42466]_ , \new_[42467]_ ,
    \new_[42468]_ , \new_[42472]_ , \new_[42473]_ , \new_[42477]_ ,
    \new_[42478]_ , \new_[42479]_ , \new_[42483]_ , \new_[42484]_ ,
    \new_[42487]_ , \new_[42490]_ , \new_[42491]_ , \new_[42492]_ ,
    \new_[42496]_ , \new_[42497]_ , \new_[42500]_ , \new_[42503]_ ,
    \new_[42504]_ , \new_[42505]_ , \new_[42509]_ , \new_[42510]_ ,
    \new_[42513]_ , \new_[42516]_ , \new_[42517]_ , \new_[42518]_ ,
    \new_[42522]_ , \new_[42523]_ , \new_[42526]_ , \new_[42529]_ ,
    \new_[42530]_ , \new_[42531]_ , \new_[42535]_ , \new_[42536]_ ,
    \new_[42539]_ , \new_[42542]_ , \new_[42543]_ , \new_[42544]_ ,
    \new_[42548]_ , \new_[42549]_ , \new_[42552]_ , \new_[42555]_ ,
    \new_[42556]_ , \new_[42557]_ , \new_[42561]_ , \new_[42562]_ ,
    \new_[42565]_ , \new_[42568]_ , \new_[42569]_ , \new_[42570]_ ,
    \new_[42574]_ , \new_[42575]_ , \new_[42578]_ , \new_[42581]_ ,
    \new_[42582]_ , \new_[42583]_ , \new_[42587]_ , \new_[42588]_ ,
    \new_[42591]_ , \new_[42594]_ , \new_[42595]_ , \new_[42596]_ ,
    \new_[42600]_ , \new_[42601]_ , \new_[42604]_ , \new_[42607]_ ,
    \new_[42608]_ , \new_[42609]_ , \new_[42613]_ , \new_[42614]_ ,
    \new_[42617]_ , \new_[42620]_ , \new_[42621]_ , \new_[42622]_ ,
    \new_[42626]_ , \new_[42627]_ , \new_[42630]_ , \new_[42633]_ ,
    \new_[42634]_ , \new_[42635]_ , \new_[42639]_ , \new_[42640]_ ,
    \new_[42643]_ , \new_[42646]_ , \new_[42647]_ , \new_[42648]_ ,
    \new_[42652]_ , \new_[42653]_ , \new_[42656]_ , \new_[42659]_ ,
    \new_[42660]_ , \new_[42661]_ , \new_[42665]_ , \new_[42666]_ ,
    \new_[42669]_ , \new_[42672]_ , \new_[42673]_ , \new_[42674]_ ,
    \new_[42678]_ , \new_[42679]_ , \new_[42682]_ , \new_[42685]_ ,
    \new_[42686]_ , \new_[42687]_ , \new_[42691]_ , \new_[42692]_ ,
    \new_[42695]_ , \new_[42698]_ , \new_[42699]_ , \new_[42700]_ ,
    \new_[42704]_ , \new_[42705]_ , \new_[42708]_ , \new_[42711]_ ,
    \new_[42712]_ , \new_[42713]_ , \new_[42717]_ , \new_[42718]_ ,
    \new_[42721]_ , \new_[42724]_ , \new_[42725]_ , \new_[42726]_ ,
    \new_[42730]_ , \new_[42731]_ , \new_[42734]_ , \new_[42737]_ ,
    \new_[42738]_ , \new_[42739]_ , \new_[42743]_ , \new_[42744]_ ,
    \new_[42747]_ , \new_[42750]_ , \new_[42751]_ , \new_[42752]_ ,
    \new_[42756]_ , \new_[42757]_ , \new_[42760]_ , \new_[42763]_ ,
    \new_[42764]_ , \new_[42765]_ , \new_[42769]_ , \new_[42770]_ ,
    \new_[42773]_ , \new_[42776]_ , \new_[42777]_ , \new_[42778]_ ,
    \new_[42782]_ , \new_[42783]_ , \new_[42786]_ , \new_[42789]_ ,
    \new_[42790]_ , \new_[42791]_ , \new_[42795]_ , \new_[42796]_ ,
    \new_[42799]_ , \new_[42802]_ , \new_[42803]_ , \new_[42804]_ ,
    \new_[42808]_ , \new_[42809]_ , \new_[42812]_ , \new_[42815]_ ,
    \new_[42816]_ , \new_[42817]_ , \new_[42821]_ , \new_[42822]_ ,
    \new_[42825]_ , \new_[42828]_ , \new_[42829]_ , \new_[42830]_ ,
    \new_[42834]_ , \new_[42835]_ , \new_[42838]_ , \new_[42841]_ ,
    \new_[42842]_ , \new_[42843]_ , \new_[42847]_ , \new_[42848]_ ,
    \new_[42851]_ , \new_[42854]_ , \new_[42855]_ , \new_[42856]_ ,
    \new_[42860]_ , \new_[42861]_ , \new_[42864]_ , \new_[42867]_ ,
    \new_[42868]_ , \new_[42869]_ , \new_[42873]_ , \new_[42874]_ ,
    \new_[42877]_ , \new_[42880]_ , \new_[42881]_ , \new_[42882]_ ,
    \new_[42886]_ , \new_[42887]_ , \new_[42890]_ , \new_[42893]_ ,
    \new_[42894]_ , \new_[42895]_ , \new_[42899]_ , \new_[42900]_ ,
    \new_[42903]_ , \new_[42906]_ , \new_[42907]_ , \new_[42908]_ ,
    \new_[42912]_ , \new_[42913]_ , \new_[42916]_ , \new_[42919]_ ,
    \new_[42920]_ , \new_[42921]_ , \new_[42925]_ , \new_[42926]_ ,
    \new_[42929]_ , \new_[42932]_ , \new_[42933]_ , \new_[42934]_ ,
    \new_[42938]_ , \new_[42939]_ , \new_[42942]_ , \new_[42945]_ ,
    \new_[42946]_ , \new_[42947]_ , \new_[42951]_ , \new_[42952]_ ,
    \new_[42955]_ , \new_[42958]_ , \new_[42959]_ , \new_[42960]_ ,
    \new_[42964]_ , \new_[42965]_ , \new_[42968]_ , \new_[42971]_ ,
    \new_[42972]_ , \new_[42973]_ , \new_[42977]_ , \new_[42978]_ ,
    \new_[42981]_ , \new_[42984]_ , \new_[42985]_ , \new_[42986]_ ,
    \new_[42990]_ , \new_[42991]_ , \new_[42994]_ , \new_[42997]_ ,
    \new_[42998]_ , \new_[42999]_ , \new_[43003]_ , \new_[43004]_ ,
    \new_[43007]_ , \new_[43010]_ , \new_[43011]_ , \new_[43012]_ ,
    \new_[43016]_ , \new_[43017]_ , \new_[43020]_ , \new_[43023]_ ,
    \new_[43024]_ , \new_[43025]_ , \new_[43029]_ , \new_[43030]_ ,
    \new_[43033]_ , \new_[43036]_ , \new_[43037]_ , \new_[43038]_ ,
    \new_[43042]_ , \new_[43043]_ , \new_[43046]_ , \new_[43049]_ ,
    \new_[43050]_ , \new_[43051]_ , \new_[43055]_ , \new_[43056]_ ,
    \new_[43059]_ , \new_[43062]_ , \new_[43063]_ , \new_[43064]_ ,
    \new_[43068]_ , \new_[43069]_ , \new_[43072]_ , \new_[43075]_ ,
    \new_[43076]_ , \new_[43077]_ , \new_[43081]_ , \new_[43082]_ ,
    \new_[43085]_ , \new_[43088]_ , \new_[43089]_ , \new_[43090]_ ,
    \new_[43094]_ , \new_[43095]_ , \new_[43098]_ , \new_[43101]_ ,
    \new_[43102]_ , \new_[43103]_ , \new_[43107]_ , \new_[43108]_ ,
    \new_[43111]_ , \new_[43114]_ , \new_[43115]_ , \new_[43116]_ ,
    \new_[43120]_ , \new_[43121]_ , \new_[43124]_ , \new_[43127]_ ,
    \new_[43128]_ , \new_[43129]_ , \new_[43133]_ , \new_[43134]_ ,
    \new_[43137]_ , \new_[43140]_ , \new_[43141]_ , \new_[43142]_ ,
    \new_[43146]_ , \new_[43147]_ , \new_[43150]_ , \new_[43153]_ ,
    \new_[43154]_ , \new_[43155]_ , \new_[43159]_ , \new_[43160]_ ,
    \new_[43163]_ , \new_[43166]_ , \new_[43167]_ , \new_[43168]_ ,
    \new_[43172]_ , \new_[43173]_ , \new_[43176]_ , \new_[43179]_ ,
    \new_[43180]_ , \new_[43181]_ , \new_[43185]_ , \new_[43186]_ ,
    \new_[43189]_ , \new_[43192]_ , \new_[43193]_ , \new_[43194]_ ,
    \new_[43198]_ , \new_[43199]_ , \new_[43202]_ , \new_[43205]_ ,
    \new_[43206]_ , \new_[43207]_ , \new_[43211]_ , \new_[43212]_ ,
    \new_[43215]_ , \new_[43218]_ , \new_[43219]_ , \new_[43220]_ ,
    \new_[43224]_ , \new_[43225]_ , \new_[43228]_ , \new_[43231]_ ,
    \new_[43232]_ , \new_[43233]_ , \new_[43237]_ , \new_[43238]_ ,
    \new_[43241]_ , \new_[43244]_ , \new_[43245]_ , \new_[43246]_ ,
    \new_[43250]_ , \new_[43251]_ , \new_[43254]_ , \new_[43257]_ ,
    \new_[43258]_ , \new_[43259]_ , \new_[43263]_ , \new_[43264]_ ,
    \new_[43267]_ , \new_[43270]_ , \new_[43271]_ , \new_[43272]_ ,
    \new_[43276]_ , \new_[43277]_ , \new_[43280]_ , \new_[43283]_ ,
    \new_[43284]_ , \new_[43285]_ , \new_[43289]_ , \new_[43290]_ ,
    \new_[43293]_ , \new_[43296]_ , \new_[43297]_ , \new_[43298]_ ,
    \new_[43302]_ , \new_[43303]_ , \new_[43306]_ , \new_[43309]_ ,
    \new_[43310]_ , \new_[43311]_ , \new_[43315]_ , \new_[43316]_ ,
    \new_[43319]_ , \new_[43322]_ , \new_[43323]_ , \new_[43324]_ ,
    \new_[43328]_ , \new_[43329]_ , \new_[43332]_ , \new_[43335]_ ,
    \new_[43336]_ , \new_[43337]_ , \new_[43341]_ , \new_[43342]_ ,
    \new_[43345]_ , \new_[43348]_ , \new_[43349]_ , \new_[43350]_ ,
    \new_[43354]_ , \new_[43355]_ , \new_[43358]_ , \new_[43361]_ ,
    \new_[43362]_ , \new_[43363]_ , \new_[43367]_ , \new_[43368]_ ,
    \new_[43371]_ , \new_[43374]_ , \new_[43375]_ , \new_[43376]_ ,
    \new_[43380]_ , \new_[43381]_ , \new_[43384]_ , \new_[43387]_ ,
    \new_[43388]_ , \new_[43389]_ , \new_[43393]_ , \new_[43394]_ ,
    \new_[43397]_ , \new_[43400]_ , \new_[43401]_ , \new_[43402]_ ,
    \new_[43406]_ , \new_[43407]_ , \new_[43410]_ , \new_[43413]_ ,
    \new_[43414]_ , \new_[43415]_ , \new_[43419]_ , \new_[43420]_ ,
    \new_[43423]_ , \new_[43426]_ , \new_[43427]_ , \new_[43428]_ ,
    \new_[43432]_ , \new_[43433]_ , \new_[43436]_ , \new_[43439]_ ,
    \new_[43440]_ , \new_[43441]_ , \new_[43445]_ , \new_[43446]_ ,
    \new_[43449]_ , \new_[43452]_ , \new_[43453]_ , \new_[43454]_ ,
    \new_[43458]_ , \new_[43459]_ , \new_[43462]_ , \new_[43465]_ ,
    \new_[43466]_ , \new_[43467]_ , \new_[43471]_ , \new_[43472]_ ,
    \new_[43475]_ , \new_[43478]_ , \new_[43479]_ , \new_[43480]_ ,
    \new_[43484]_ , \new_[43485]_ , \new_[43488]_ , \new_[43491]_ ,
    \new_[43492]_ , \new_[43493]_ , \new_[43497]_ , \new_[43498]_ ,
    \new_[43501]_ , \new_[43504]_ , \new_[43505]_ , \new_[43506]_ ,
    \new_[43510]_ , \new_[43511]_ , \new_[43514]_ , \new_[43517]_ ,
    \new_[43518]_ , \new_[43519]_ , \new_[43523]_ , \new_[43524]_ ,
    \new_[43527]_ , \new_[43530]_ , \new_[43531]_ , \new_[43532]_ ,
    \new_[43536]_ , \new_[43537]_ , \new_[43540]_ , \new_[43543]_ ,
    \new_[43544]_ , \new_[43545]_ , \new_[43549]_ , \new_[43550]_ ,
    \new_[43553]_ , \new_[43556]_ , \new_[43557]_ , \new_[43558]_ ,
    \new_[43562]_ , \new_[43563]_ , \new_[43566]_ , \new_[43569]_ ,
    \new_[43570]_ , \new_[43571]_ , \new_[43575]_ , \new_[43576]_ ,
    \new_[43579]_ , \new_[43582]_ , \new_[43583]_ , \new_[43584]_ ,
    \new_[43588]_ , \new_[43589]_ , \new_[43592]_ , \new_[43595]_ ,
    \new_[43596]_ , \new_[43597]_ , \new_[43601]_ , \new_[43602]_ ,
    \new_[43605]_ , \new_[43608]_ , \new_[43609]_ , \new_[43610]_ ,
    \new_[43614]_ , \new_[43615]_ , \new_[43618]_ , \new_[43621]_ ,
    \new_[43622]_ , \new_[43623]_ , \new_[43627]_ , \new_[43628]_ ,
    \new_[43631]_ , \new_[43634]_ , \new_[43635]_ , \new_[43636]_ ,
    \new_[43640]_ , \new_[43641]_ , \new_[43644]_ , \new_[43647]_ ,
    \new_[43648]_ , \new_[43649]_ , \new_[43653]_ , \new_[43654]_ ,
    \new_[43657]_ , \new_[43660]_ , \new_[43661]_ , \new_[43662]_ ,
    \new_[43666]_ , \new_[43667]_ , \new_[43670]_ , \new_[43673]_ ,
    \new_[43674]_ , \new_[43675]_ , \new_[43679]_ , \new_[43680]_ ,
    \new_[43683]_ , \new_[43686]_ , \new_[43687]_ , \new_[43688]_ ,
    \new_[43692]_ , \new_[43693]_ , \new_[43696]_ , \new_[43699]_ ,
    \new_[43700]_ , \new_[43701]_ , \new_[43705]_ , \new_[43706]_ ,
    \new_[43709]_ , \new_[43712]_ , \new_[43713]_ , \new_[43714]_ ,
    \new_[43718]_ , \new_[43719]_ , \new_[43722]_ , \new_[43725]_ ,
    \new_[43726]_ , \new_[43727]_ , \new_[43731]_ , \new_[43732]_ ,
    \new_[43735]_ , \new_[43738]_ , \new_[43739]_ , \new_[43740]_ ,
    \new_[43744]_ , \new_[43745]_ , \new_[43748]_ , \new_[43751]_ ,
    \new_[43752]_ , \new_[43753]_ , \new_[43757]_ , \new_[43758]_ ,
    \new_[43761]_ , \new_[43764]_ , \new_[43765]_ , \new_[43766]_ ,
    \new_[43770]_ , \new_[43771]_ , \new_[43774]_ , \new_[43777]_ ,
    \new_[43778]_ , \new_[43779]_ , \new_[43783]_ , \new_[43784]_ ,
    \new_[43787]_ , \new_[43790]_ , \new_[43791]_ , \new_[43792]_ ,
    \new_[43796]_ , \new_[43797]_ , \new_[43800]_ , \new_[43803]_ ,
    \new_[43804]_ , \new_[43805]_ , \new_[43809]_ , \new_[43810]_ ,
    \new_[43813]_ , \new_[43816]_ , \new_[43817]_ , \new_[43818]_ ,
    \new_[43822]_ , \new_[43823]_ , \new_[43826]_ , \new_[43829]_ ,
    \new_[43830]_ , \new_[43831]_ , \new_[43835]_ , \new_[43836]_ ,
    \new_[43839]_ , \new_[43842]_ , \new_[43843]_ , \new_[43844]_ ,
    \new_[43848]_ , \new_[43849]_ , \new_[43852]_ , \new_[43855]_ ,
    \new_[43856]_ , \new_[43857]_ , \new_[43861]_ , \new_[43862]_ ,
    \new_[43865]_ , \new_[43868]_ , \new_[43869]_ , \new_[43870]_ ,
    \new_[43874]_ , \new_[43875]_ , \new_[43878]_ , \new_[43881]_ ,
    \new_[43882]_ , \new_[43883]_ , \new_[43887]_ , \new_[43888]_ ,
    \new_[43891]_ , \new_[43894]_ , \new_[43895]_ , \new_[43896]_ ,
    \new_[43900]_ , \new_[43901]_ , \new_[43904]_ , \new_[43907]_ ,
    \new_[43908]_ , \new_[43909]_ , \new_[43913]_ , \new_[43914]_ ,
    \new_[43917]_ , \new_[43920]_ , \new_[43921]_ , \new_[43922]_ ,
    \new_[43926]_ , \new_[43927]_ , \new_[43930]_ , \new_[43933]_ ,
    \new_[43934]_ , \new_[43935]_ , \new_[43939]_ , \new_[43940]_ ,
    \new_[43943]_ , \new_[43946]_ , \new_[43947]_ , \new_[43948]_ ,
    \new_[43952]_ , \new_[43953]_ , \new_[43956]_ , \new_[43959]_ ,
    \new_[43960]_ , \new_[43961]_ , \new_[43965]_ , \new_[43966]_ ,
    \new_[43969]_ , \new_[43972]_ , \new_[43973]_ , \new_[43974]_ ,
    \new_[43978]_ , \new_[43979]_ , \new_[43982]_ , \new_[43985]_ ,
    \new_[43986]_ , \new_[43987]_ , \new_[43991]_ , \new_[43992]_ ,
    \new_[43995]_ , \new_[43998]_ , \new_[43999]_ , \new_[44000]_ ,
    \new_[44004]_ , \new_[44005]_ , \new_[44008]_ , \new_[44011]_ ,
    \new_[44012]_ , \new_[44013]_ , \new_[44017]_ , \new_[44018]_ ,
    \new_[44021]_ , \new_[44024]_ , \new_[44025]_ , \new_[44026]_ ,
    \new_[44030]_ , \new_[44031]_ , \new_[44034]_ , \new_[44037]_ ,
    \new_[44038]_ , \new_[44039]_ , \new_[44043]_ , \new_[44044]_ ,
    \new_[44047]_ , \new_[44050]_ , \new_[44051]_ , \new_[44052]_ ,
    \new_[44056]_ , \new_[44057]_ , \new_[44060]_ , \new_[44063]_ ,
    \new_[44064]_ , \new_[44065]_ , \new_[44069]_ , \new_[44070]_ ,
    \new_[44073]_ , \new_[44076]_ , \new_[44077]_ , \new_[44078]_ ,
    \new_[44082]_ , \new_[44083]_ , \new_[44086]_ , \new_[44089]_ ,
    \new_[44090]_ , \new_[44091]_ , \new_[44095]_ , \new_[44096]_ ,
    \new_[44099]_ , \new_[44102]_ , \new_[44103]_ , \new_[44104]_ ,
    \new_[44108]_ , \new_[44109]_ , \new_[44112]_ , \new_[44115]_ ,
    \new_[44116]_ , \new_[44117]_ , \new_[44121]_ , \new_[44122]_ ,
    \new_[44125]_ , \new_[44128]_ , \new_[44129]_ , \new_[44130]_ ,
    \new_[44134]_ , \new_[44135]_ , \new_[44138]_ , \new_[44141]_ ,
    \new_[44142]_ , \new_[44143]_ , \new_[44147]_ , \new_[44148]_ ,
    \new_[44151]_ , \new_[44154]_ , \new_[44155]_ , \new_[44156]_ ,
    \new_[44160]_ , \new_[44161]_ , \new_[44164]_ , \new_[44167]_ ,
    \new_[44168]_ , \new_[44169]_ , \new_[44173]_ , \new_[44174]_ ,
    \new_[44177]_ , \new_[44180]_ , \new_[44181]_ , \new_[44182]_ ,
    \new_[44186]_ , \new_[44187]_ , \new_[44190]_ , \new_[44193]_ ,
    \new_[44194]_ , \new_[44195]_ , \new_[44199]_ , \new_[44200]_ ,
    \new_[44203]_ , \new_[44206]_ , \new_[44207]_ , \new_[44208]_ ,
    \new_[44212]_ , \new_[44213]_ , \new_[44216]_ , \new_[44219]_ ,
    \new_[44220]_ , \new_[44221]_ , \new_[44225]_ , \new_[44226]_ ,
    \new_[44229]_ , \new_[44232]_ , \new_[44233]_ , \new_[44234]_ ,
    \new_[44238]_ , \new_[44239]_ , \new_[44242]_ , \new_[44245]_ ,
    \new_[44246]_ , \new_[44247]_ , \new_[44251]_ , \new_[44252]_ ,
    \new_[44255]_ , \new_[44258]_ , \new_[44259]_ , \new_[44260]_ ,
    \new_[44264]_ , \new_[44265]_ , \new_[44268]_ , \new_[44271]_ ,
    \new_[44272]_ , \new_[44273]_ , \new_[44277]_ , \new_[44278]_ ,
    \new_[44281]_ , \new_[44284]_ , \new_[44285]_ , \new_[44286]_ ,
    \new_[44290]_ , \new_[44291]_ , \new_[44294]_ , \new_[44297]_ ,
    \new_[44298]_ , \new_[44299]_ , \new_[44303]_ , \new_[44304]_ ,
    \new_[44307]_ , \new_[44310]_ , \new_[44311]_ , \new_[44312]_ ,
    \new_[44316]_ , \new_[44317]_ , \new_[44320]_ , \new_[44323]_ ,
    \new_[44324]_ , \new_[44325]_ , \new_[44329]_ , \new_[44330]_ ,
    \new_[44333]_ , \new_[44336]_ , \new_[44337]_ , \new_[44338]_ ,
    \new_[44342]_ , \new_[44343]_ , \new_[44346]_ , \new_[44349]_ ,
    \new_[44350]_ , \new_[44351]_ , \new_[44355]_ , \new_[44356]_ ,
    \new_[44359]_ , \new_[44362]_ , \new_[44363]_ , \new_[44364]_ ,
    \new_[44368]_ , \new_[44369]_ , \new_[44372]_ , \new_[44375]_ ,
    \new_[44376]_ , \new_[44377]_ , \new_[44381]_ , \new_[44382]_ ,
    \new_[44385]_ , \new_[44388]_ , \new_[44389]_ , \new_[44390]_ ,
    \new_[44394]_ , \new_[44395]_ , \new_[44398]_ , \new_[44401]_ ,
    \new_[44402]_ , \new_[44403]_ , \new_[44407]_ , \new_[44408]_ ,
    \new_[44411]_ , \new_[44414]_ , \new_[44415]_ , \new_[44416]_ ,
    \new_[44420]_ , \new_[44421]_ , \new_[44424]_ , \new_[44427]_ ,
    \new_[44428]_ , \new_[44429]_ , \new_[44433]_ , \new_[44434]_ ,
    \new_[44437]_ , \new_[44440]_ , \new_[44441]_ , \new_[44442]_ ,
    \new_[44446]_ , \new_[44447]_ , \new_[44450]_ , \new_[44453]_ ,
    \new_[44454]_ , \new_[44455]_ , \new_[44459]_ , \new_[44460]_ ,
    \new_[44463]_ , \new_[44466]_ , \new_[44467]_ , \new_[44468]_ ,
    \new_[44472]_ , \new_[44473]_ , \new_[44476]_ , \new_[44479]_ ,
    \new_[44480]_ , \new_[44481]_ , \new_[44485]_ , \new_[44486]_ ,
    \new_[44489]_ , \new_[44492]_ , \new_[44493]_ , \new_[44494]_ ,
    \new_[44498]_ , \new_[44499]_ , \new_[44502]_ , \new_[44505]_ ,
    \new_[44506]_ , \new_[44507]_ , \new_[44511]_ , \new_[44512]_ ,
    \new_[44515]_ , \new_[44518]_ , \new_[44519]_ , \new_[44520]_ ,
    \new_[44524]_ , \new_[44525]_ , \new_[44528]_ , \new_[44531]_ ,
    \new_[44532]_ , \new_[44533]_ , \new_[44537]_ , \new_[44538]_ ,
    \new_[44541]_ , \new_[44544]_ , \new_[44545]_ , \new_[44546]_ ,
    \new_[44550]_ , \new_[44551]_ , \new_[44554]_ , \new_[44557]_ ,
    \new_[44558]_ , \new_[44559]_ , \new_[44563]_ , \new_[44564]_ ,
    \new_[44567]_ , \new_[44570]_ , \new_[44571]_ , \new_[44572]_ ,
    \new_[44576]_ , \new_[44577]_ , \new_[44580]_ , \new_[44583]_ ,
    \new_[44584]_ , \new_[44585]_ , \new_[44589]_ , \new_[44590]_ ,
    \new_[44593]_ , \new_[44596]_ , \new_[44597]_ , \new_[44598]_ ,
    \new_[44602]_ , \new_[44603]_ , \new_[44606]_ , \new_[44609]_ ,
    \new_[44610]_ , \new_[44611]_ , \new_[44615]_ , \new_[44616]_ ,
    \new_[44619]_ , \new_[44622]_ , \new_[44623]_ , \new_[44624]_ ,
    \new_[44628]_ , \new_[44629]_ , \new_[44632]_ , \new_[44635]_ ,
    \new_[44636]_ , \new_[44637]_ , \new_[44641]_ , \new_[44642]_ ,
    \new_[44645]_ , \new_[44648]_ , \new_[44649]_ , \new_[44650]_ ,
    \new_[44654]_ , \new_[44655]_ , \new_[44658]_ , \new_[44661]_ ,
    \new_[44662]_ , \new_[44663]_ , \new_[44667]_ , \new_[44668]_ ,
    \new_[44671]_ , \new_[44674]_ , \new_[44675]_ , \new_[44676]_ ,
    \new_[44680]_ , \new_[44681]_ , \new_[44684]_ , \new_[44687]_ ,
    \new_[44688]_ , \new_[44689]_ , \new_[44693]_ , \new_[44694]_ ,
    \new_[44697]_ , \new_[44700]_ , \new_[44701]_ , \new_[44702]_ ,
    \new_[44706]_ , \new_[44707]_ , \new_[44710]_ , \new_[44713]_ ,
    \new_[44714]_ , \new_[44715]_ , \new_[44719]_ , \new_[44720]_ ,
    \new_[44723]_ , \new_[44726]_ , \new_[44727]_ , \new_[44728]_ ,
    \new_[44732]_ , \new_[44733]_ , \new_[44736]_ , \new_[44739]_ ,
    \new_[44740]_ , \new_[44741]_ , \new_[44745]_ , \new_[44746]_ ,
    \new_[44749]_ , \new_[44752]_ , \new_[44753]_ , \new_[44754]_ ,
    \new_[44758]_ , \new_[44759]_ , \new_[44762]_ , \new_[44765]_ ,
    \new_[44766]_ , \new_[44767]_ , \new_[44771]_ , \new_[44772]_ ,
    \new_[44775]_ , \new_[44778]_ , \new_[44779]_ , \new_[44780]_ ,
    \new_[44784]_ , \new_[44785]_ , \new_[44788]_ , \new_[44791]_ ,
    \new_[44792]_ , \new_[44793]_ , \new_[44797]_ , \new_[44798]_ ,
    \new_[44801]_ , \new_[44804]_ , \new_[44805]_ , \new_[44806]_ ,
    \new_[44810]_ , \new_[44811]_ , \new_[44814]_ , \new_[44817]_ ,
    \new_[44818]_ , \new_[44819]_ , \new_[44823]_ , \new_[44824]_ ,
    \new_[44827]_ , \new_[44830]_ , \new_[44831]_ , \new_[44832]_ ,
    \new_[44836]_ , \new_[44837]_ , \new_[44840]_ , \new_[44843]_ ,
    \new_[44844]_ , \new_[44845]_ , \new_[44849]_ , \new_[44850]_ ,
    \new_[44853]_ , \new_[44856]_ , \new_[44857]_ , \new_[44858]_ ,
    \new_[44862]_ , \new_[44863]_ , \new_[44866]_ , \new_[44869]_ ,
    \new_[44870]_ , \new_[44871]_ , \new_[44875]_ , \new_[44876]_ ,
    \new_[44879]_ , \new_[44882]_ , \new_[44883]_ , \new_[44884]_ ,
    \new_[44888]_ , \new_[44889]_ , \new_[44892]_ , \new_[44895]_ ,
    \new_[44896]_ , \new_[44897]_ , \new_[44901]_ , \new_[44902]_ ,
    \new_[44905]_ , \new_[44908]_ , \new_[44909]_ , \new_[44910]_ ,
    \new_[44914]_ , \new_[44915]_ , \new_[44918]_ , \new_[44921]_ ,
    \new_[44922]_ , \new_[44923]_ , \new_[44927]_ , \new_[44928]_ ,
    \new_[44931]_ , \new_[44934]_ , \new_[44935]_ , \new_[44936]_ ,
    \new_[44940]_ , \new_[44941]_ , \new_[44944]_ , \new_[44947]_ ,
    \new_[44948]_ , \new_[44949]_ , \new_[44953]_ , \new_[44954]_ ,
    \new_[44957]_ , \new_[44960]_ , \new_[44961]_ , \new_[44962]_ ,
    \new_[44966]_ , \new_[44967]_ , \new_[44970]_ , \new_[44973]_ ,
    \new_[44974]_ , \new_[44975]_ , \new_[44979]_ , \new_[44980]_ ,
    \new_[44983]_ , \new_[44986]_ , \new_[44987]_ , \new_[44988]_ ,
    \new_[44992]_ , \new_[44993]_ , \new_[44996]_ , \new_[44999]_ ,
    \new_[45000]_ , \new_[45001]_ , \new_[45005]_ , \new_[45006]_ ,
    \new_[45009]_ , \new_[45012]_ , \new_[45013]_ , \new_[45014]_ ,
    \new_[45018]_ , \new_[45019]_ , \new_[45022]_ , \new_[45025]_ ,
    \new_[45026]_ , \new_[45027]_ , \new_[45031]_ , \new_[45032]_ ,
    \new_[45035]_ , \new_[45038]_ , \new_[45039]_ , \new_[45040]_ ,
    \new_[45044]_ , \new_[45045]_ , \new_[45048]_ , \new_[45051]_ ,
    \new_[45052]_ , \new_[45053]_ , \new_[45057]_ , \new_[45058]_ ,
    \new_[45061]_ , \new_[45064]_ , \new_[45065]_ , \new_[45066]_ ,
    \new_[45070]_ , \new_[45071]_ , \new_[45074]_ , \new_[45077]_ ,
    \new_[45078]_ , \new_[45079]_ , \new_[45083]_ , \new_[45084]_ ,
    \new_[45087]_ , \new_[45090]_ , \new_[45091]_ , \new_[45092]_ ,
    \new_[45096]_ , \new_[45097]_ , \new_[45100]_ , \new_[45103]_ ,
    \new_[45104]_ , \new_[45105]_ , \new_[45109]_ , \new_[45110]_ ,
    \new_[45113]_ , \new_[45116]_ , \new_[45117]_ , \new_[45118]_ ,
    \new_[45122]_ , \new_[45123]_ , \new_[45126]_ , \new_[45129]_ ,
    \new_[45130]_ , \new_[45131]_ , \new_[45135]_ , \new_[45136]_ ,
    \new_[45139]_ , \new_[45142]_ , \new_[45143]_ , \new_[45144]_ ,
    \new_[45148]_ , \new_[45149]_ , \new_[45152]_ , \new_[45155]_ ,
    \new_[45156]_ , \new_[45157]_ , \new_[45161]_ , \new_[45162]_ ,
    \new_[45165]_ , \new_[45168]_ , \new_[45169]_ , \new_[45170]_ ,
    \new_[45174]_ , \new_[45175]_ , \new_[45178]_ , \new_[45181]_ ,
    \new_[45182]_ , \new_[45183]_ , \new_[45187]_ , \new_[45188]_ ,
    \new_[45191]_ , \new_[45194]_ , \new_[45195]_ , \new_[45196]_ ,
    \new_[45200]_ , \new_[45201]_ , \new_[45204]_ , \new_[45207]_ ,
    \new_[45208]_ , \new_[45209]_ , \new_[45213]_ , \new_[45214]_ ,
    \new_[45217]_ , \new_[45220]_ , \new_[45221]_ , \new_[45222]_ ,
    \new_[45226]_ , \new_[45227]_ , \new_[45230]_ , \new_[45233]_ ,
    \new_[45234]_ , \new_[45235]_ , \new_[45239]_ , \new_[45240]_ ,
    \new_[45243]_ , \new_[45246]_ , \new_[45247]_ , \new_[45248]_ ,
    \new_[45252]_ , \new_[45253]_ , \new_[45256]_ , \new_[45259]_ ,
    \new_[45260]_ , \new_[45261]_ , \new_[45265]_ , \new_[45266]_ ,
    \new_[45269]_ , \new_[45272]_ , \new_[45273]_ , \new_[45274]_ ,
    \new_[45278]_ , \new_[45279]_ , \new_[45282]_ , \new_[45285]_ ,
    \new_[45286]_ , \new_[45287]_ , \new_[45291]_ , \new_[45292]_ ,
    \new_[45295]_ , \new_[45298]_ , \new_[45299]_ , \new_[45300]_ ,
    \new_[45304]_ , \new_[45305]_ , \new_[45308]_ , \new_[45311]_ ,
    \new_[45312]_ , \new_[45313]_ , \new_[45317]_ , \new_[45318]_ ,
    \new_[45321]_ , \new_[45324]_ , \new_[45325]_ , \new_[45326]_ ,
    \new_[45330]_ , \new_[45331]_ , \new_[45334]_ , \new_[45337]_ ,
    \new_[45338]_ , \new_[45339]_ , \new_[45343]_ , \new_[45344]_ ,
    \new_[45347]_ , \new_[45350]_ , \new_[45351]_ , \new_[45352]_ ,
    \new_[45356]_ , \new_[45357]_ , \new_[45360]_ , \new_[45363]_ ,
    \new_[45364]_ , \new_[45365]_ , \new_[45369]_ , \new_[45370]_ ,
    \new_[45373]_ , \new_[45376]_ , \new_[45377]_ , \new_[45378]_ ,
    \new_[45382]_ , \new_[45383]_ , \new_[45386]_ , \new_[45389]_ ,
    \new_[45390]_ , \new_[45391]_ , \new_[45395]_ , \new_[45396]_ ,
    \new_[45399]_ , \new_[45402]_ , \new_[45403]_ , \new_[45404]_ ,
    \new_[45408]_ , \new_[45409]_ , \new_[45412]_ , \new_[45415]_ ,
    \new_[45416]_ , \new_[45417]_ , \new_[45421]_ , \new_[45422]_ ,
    \new_[45425]_ , \new_[45428]_ , \new_[45429]_ , \new_[45430]_ ,
    \new_[45434]_ , \new_[45435]_ , \new_[45438]_ , \new_[45441]_ ,
    \new_[45442]_ , \new_[45443]_ , \new_[45447]_ , \new_[45448]_ ,
    \new_[45451]_ , \new_[45454]_ , \new_[45455]_ , \new_[45456]_ ,
    \new_[45460]_ , \new_[45461]_ , \new_[45464]_ , \new_[45467]_ ,
    \new_[45468]_ , \new_[45469]_ , \new_[45473]_ , \new_[45474]_ ,
    \new_[45477]_ , \new_[45480]_ , \new_[45481]_ , \new_[45482]_ ,
    \new_[45486]_ , \new_[45487]_ , \new_[45490]_ , \new_[45493]_ ,
    \new_[45494]_ , \new_[45495]_ , \new_[45499]_ , \new_[45500]_ ,
    \new_[45503]_ , \new_[45506]_ , \new_[45507]_ , \new_[45508]_ ,
    \new_[45512]_ , \new_[45513]_ , \new_[45516]_ , \new_[45519]_ ,
    \new_[45520]_ , \new_[45521]_ , \new_[45525]_ , \new_[45526]_ ,
    \new_[45529]_ , \new_[45532]_ , \new_[45533]_ , \new_[45534]_ ,
    \new_[45538]_ , \new_[45539]_ , \new_[45542]_ , \new_[45545]_ ,
    \new_[45546]_ , \new_[45547]_ , \new_[45551]_ , \new_[45552]_ ,
    \new_[45555]_ , \new_[45558]_ , \new_[45559]_ , \new_[45560]_ ,
    \new_[45564]_ , \new_[45565]_ , \new_[45568]_ , \new_[45571]_ ,
    \new_[45572]_ , \new_[45573]_ , \new_[45577]_ , \new_[45578]_ ,
    \new_[45581]_ , \new_[45584]_ , \new_[45585]_ , \new_[45586]_ ,
    \new_[45590]_ , \new_[45591]_ , \new_[45594]_ , \new_[45597]_ ,
    \new_[45598]_ , \new_[45599]_ , \new_[45603]_ , \new_[45604]_ ,
    \new_[45607]_ , \new_[45610]_ , \new_[45611]_ , \new_[45612]_ ,
    \new_[45616]_ , \new_[45617]_ , \new_[45620]_ , \new_[45623]_ ,
    \new_[45624]_ , \new_[45625]_ , \new_[45629]_ , \new_[45630]_ ,
    \new_[45633]_ , \new_[45636]_ , \new_[45637]_ , \new_[45638]_ ,
    \new_[45642]_ , \new_[45643]_ , \new_[45646]_ , \new_[45649]_ ,
    \new_[45650]_ , \new_[45651]_ , \new_[45655]_ , \new_[45656]_ ,
    \new_[45659]_ , \new_[45662]_ , \new_[45663]_ , \new_[45664]_ ,
    \new_[45668]_ , \new_[45669]_ , \new_[45672]_ , \new_[45675]_ ,
    \new_[45676]_ , \new_[45677]_ , \new_[45681]_ , \new_[45682]_ ,
    \new_[45685]_ , \new_[45688]_ , \new_[45689]_ , \new_[45690]_ ,
    \new_[45694]_ , \new_[45695]_ , \new_[45698]_ , \new_[45701]_ ,
    \new_[45702]_ , \new_[45703]_ , \new_[45707]_ , \new_[45708]_ ,
    \new_[45711]_ , \new_[45714]_ , \new_[45715]_ , \new_[45716]_ ,
    \new_[45720]_ , \new_[45721]_ , \new_[45724]_ , \new_[45727]_ ,
    \new_[45728]_ , \new_[45729]_ , \new_[45733]_ , \new_[45734]_ ,
    \new_[45737]_ , \new_[45740]_ , \new_[45741]_ , \new_[45742]_ ,
    \new_[45746]_ , \new_[45747]_ , \new_[45750]_ , \new_[45753]_ ,
    \new_[45754]_ , \new_[45755]_ , \new_[45759]_ , \new_[45760]_ ,
    \new_[45763]_ , \new_[45766]_ , \new_[45767]_ , \new_[45768]_ ,
    \new_[45772]_ , \new_[45773]_ , \new_[45776]_ , \new_[45779]_ ,
    \new_[45780]_ , \new_[45781]_ , \new_[45785]_ , \new_[45786]_ ,
    \new_[45789]_ , \new_[45792]_ , \new_[45793]_ , \new_[45794]_ ,
    \new_[45798]_ , \new_[45799]_ , \new_[45802]_ , \new_[45805]_ ,
    \new_[45806]_ , \new_[45807]_ , \new_[45811]_ , \new_[45812]_ ,
    \new_[45815]_ , \new_[45818]_ , \new_[45819]_ , \new_[45820]_ ,
    \new_[45824]_ , \new_[45825]_ , \new_[45828]_ , \new_[45831]_ ,
    \new_[45832]_ , \new_[45833]_ , \new_[45837]_ , \new_[45838]_ ,
    \new_[45841]_ , \new_[45844]_ , \new_[45845]_ , \new_[45846]_ ,
    \new_[45850]_ , \new_[45851]_ , \new_[45854]_ , \new_[45857]_ ,
    \new_[45858]_ , \new_[45859]_ , \new_[45863]_ , \new_[45864]_ ,
    \new_[45867]_ , \new_[45870]_ , \new_[45871]_ , \new_[45872]_ ,
    \new_[45876]_ , \new_[45877]_ , \new_[45880]_ , \new_[45883]_ ,
    \new_[45884]_ , \new_[45885]_ , \new_[45889]_ , \new_[45890]_ ,
    \new_[45893]_ , \new_[45896]_ , \new_[45897]_ , \new_[45898]_ ,
    \new_[45902]_ , \new_[45903]_ , \new_[45906]_ , \new_[45909]_ ,
    \new_[45910]_ , \new_[45911]_ , \new_[45915]_ , \new_[45916]_ ,
    \new_[45919]_ , \new_[45922]_ , \new_[45923]_ , \new_[45924]_ ,
    \new_[45928]_ , \new_[45929]_ , \new_[45932]_ , \new_[45935]_ ,
    \new_[45936]_ , \new_[45937]_ , \new_[45941]_ , \new_[45942]_ ,
    \new_[45945]_ , \new_[45948]_ , \new_[45949]_ , \new_[45950]_ ,
    \new_[45954]_ , \new_[45955]_ , \new_[45958]_ , \new_[45961]_ ,
    \new_[45962]_ , \new_[45963]_ , \new_[45967]_ , \new_[45968]_ ,
    \new_[45971]_ , \new_[45974]_ , \new_[45975]_ , \new_[45976]_ ,
    \new_[45980]_ , \new_[45981]_ , \new_[45984]_ , \new_[45987]_ ,
    \new_[45988]_ , \new_[45989]_ , \new_[45993]_ , \new_[45994]_ ,
    \new_[45997]_ , \new_[46000]_ , \new_[46001]_ , \new_[46002]_ ,
    \new_[46006]_ , \new_[46007]_ , \new_[46010]_ , \new_[46013]_ ,
    \new_[46014]_ , \new_[46015]_ , \new_[46019]_ , \new_[46020]_ ,
    \new_[46023]_ , \new_[46026]_ , \new_[46027]_ , \new_[46028]_ ,
    \new_[46032]_ , \new_[46033]_ , \new_[46036]_ , \new_[46039]_ ,
    \new_[46040]_ , \new_[46041]_ , \new_[46045]_ , \new_[46046]_ ,
    \new_[46049]_ , \new_[46052]_ , \new_[46053]_ , \new_[46054]_ ,
    \new_[46058]_ , \new_[46059]_ , \new_[46062]_ , \new_[46065]_ ,
    \new_[46066]_ , \new_[46067]_ , \new_[46071]_ , \new_[46072]_ ,
    \new_[46075]_ , \new_[46078]_ , \new_[46079]_ , \new_[46080]_ ,
    \new_[46084]_ , \new_[46085]_ , \new_[46088]_ , \new_[46091]_ ,
    \new_[46092]_ , \new_[46093]_ , \new_[46097]_ , \new_[46098]_ ,
    \new_[46101]_ , \new_[46104]_ , \new_[46105]_ , \new_[46106]_ ,
    \new_[46110]_ , \new_[46111]_ , \new_[46114]_ , \new_[46117]_ ,
    \new_[46118]_ , \new_[46119]_ , \new_[46123]_ , \new_[46124]_ ,
    \new_[46127]_ , \new_[46130]_ , \new_[46131]_ , \new_[46132]_ ,
    \new_[46136]_ , \new_[46137]_ , \new_[46140]_ , \new_[46143]_ ,
    \new_[46144]_ , \new_[46145]_ , \new_[46149]_ , \new_[46150]_ ,
    \new_[46153]_ , \new_[46156]_ , \new_[46157]_ , \new_[46158]_ ,
    \new_[46162]_ , \new_[46163]_ , \new_[46166]_ , \new_[46169]_ ,
    \new_[46170]_ , \new_[46171]_ , \new_[46175]_ , \new_[46176]_ ,
    \new_[46179]_ , \new_[46182]_ , \new_[46183]_ , \new_[46184]_ ,
    \new_[46188]_ , \new_[46189]_ , \new_[46192]_ , \new_[46195]_ ,
    \new_[46196]_ , \new_[46197]_ , \new_[46201]_ , \new_[46202]_ ,
    \new_[46205]_ , \new_[46208]_ , \new_[46209]_ , \new_[46210]_ ,
    \new_[46214]_ , \new_[46215]_ , \new_[46218]_ , \new_[46221]_ ,
    \new_[46222]_ , \new_[46223]_ , \new_[46227]_ , \new_[46228]_ ,
    \new_[46231]_ , \new_[46234]_ , \new_[46235]_ , \new_[46236]_ ,
    \new_[46240]_ , \new_[46241]_ , \new_[46244]_ , \new_[46247]_ ,
    \new_[46248]_ , \new_[46249]_ , \new_[46253]_ , \new_[46254]_ ,
    \new_[46257]_ , \new_[46260]_ , \new_[46261]_ , \new_[46262]_ ,
    \new_[46266]_ , \new_[46267]_ , \new_[46270]_ , \new_[46273]_ ,
    \new_[46274]_ , \new_[46275]_ , \new_[46279]_ , \new_[46280]_ ,
    \new_[46283]_ , \new_[46286]_ , \new_[46287]_ , \new_[46288]_ ,
    \new_[46292]_ , \new_[46293]_ , \new_[46296]_ , \new_[46299]_ ,
    \new_[46300]_ , \new_[46301]_ , \new_[46305]_ , \new_[46306]_ ,
    \new_[46309]_ , \new_[46312]_ , \new_[46313]_ , \new_[46314]_ ,
    \new_[46318]_ , \new_[46319]_ , \new_[46322]_ , \new_[46325]_ ,
    \new_[46326]_ , \new_[46327]_ , \new_[46331]_ , \new_[46332]_ ,
    \new_[46335]_ , \new_[46338]_ , \new_[46339]_ , \new_[46340]_ ,
    \new_[46344]_ , \new_[46345]_ , \new_[46348]_ , \new_[46351]_ ,
    \new_[46352]_ , \new_[46353]_ , \new_[46357]_ , \new_[46358]_ ,
    \new_[46361]_ , \new_[46364]_ , \new_[46365]_ , \new_[46366]_ ,
    \new_[46370]_ , \new_[46371]_ , \new_[46374]_ , \new_[46377]_ ,
    \new_[46378]_ , \new_[46379]_ , \new_[46383]_ , \new_[46384]_ ,
    \new_[46387]_ , \new_[46390]_ , \new_[46391]_ , \new_[46392]_ ,
    \new_[46396]_ , \new_[46397]_ , \new_[46400]_ , \new_[46403]_ ,
    \new_[46404]_ , \new_[46405]_ , \new_[46409]_ , \new_[46410]_ ,
    \new_[46413]_ , \new_[46416]_ , \new_[46417]_ , \new_[46418]_ ,
    \new_[46422]_ , \new_[46423]_ , \new_[46426]_ , \new_[46429]_ ,
    \new_[46430]_ , \new_[46431]_ , \new_[46435]_ , \new_[46436]_ ,
    \new_[46439]_ , \new_[46442]_ , \new_[46443]_ , \new_[46444]_ ,
    \new_[46448]_ , \new_[46449]_ , \new_[46452]_ , \new_[46455]_ ,
    \new_[46456]_ , \new_[46457]_ , \new_[46461]_ , \new_[46462]_ ,
    \new_[46465]_ , \new_[46468]_ , \new_[46469]_ , \new_[46470]_ ,
    \new_[46474]_ , \new_[46475]_ , \new_[46478]_ , \new_[46481]_ ,
    \new_[46482]_ , \new_[46483]_ , \new_[46487]_ , \new_[46488]_ ,
    \new_[46491]_ , \new_[46494]_ , \new_[46495]_ , \new_[46496]_ ,
    \new_[46500]_ , \new_[46501]_ , \new_[46504]_ , \new_[46507]_ ,
    \new_[46508]_ , \new_[46509]_ , \new_[46513]_ , \new_[46514]_ ,
    \new_[46517]_ , \new_[46520]_ , \new_[46521]_ , \new_[46522]_ ,
    \new_[46526]_ , \new_[46527]_ , \new_[46530]_ , \new_[46533]_ ,
    \new_[46534]_ , \new_[46535]_ , \new_[46539]_ , \new_[46540]_ ,
    \new_[46543]_ , \new_[46546]_ , \new_[46547]_ , \new_[46548]_ ,
    \new_[46552]_ , \new_[46553]_ , \new_[46556]_ , \new_[46559]_ ,
    \new_[46560]_ , \new_[46561]_ , \new_[46565]_ , \new_[46566]_ ,
    \new_[46569]_ , \new_[46572]_ , \new_[46573]_ , \new_[46574]_ ,
    \new_[46578]_ , \new_[46579]_ , \new_[46582]_ , \new_[46585]_ ,
    \new_[46586]_ , \new_[46587]_ , \new_[46591]_ , \new_[46592]_ ,
    \new_[46595]_ , \new_[46598]_ , \new_[46599]_ , \new_[46600]_ ,
    \new_[46604]_ , \new_[46605]_ , \new_[46608]_ , \new_[46611]_ ,
    \new_[46612]_ , \new_[46613]_ , \new_[46617]_ , \new_[46618]_ ,
    \new_[46621]_ , \new_[46624]_ , \new_[46625]_ , \new_[46626]_ ,
    \new_[46630]_ , \new_[46631]_ , \new_[46634]_ , \new_[46637]_ ,
    \new_[46638]_ , \new_[46639]_ , \new_[46643]_ , \new_[46644]_ ,
    \new_[46647]_ , \new_[46650]_ , \new_[46651]_ , \new_[46652]_ ,
    \new_[46656]_ , \new_[46657]_ , \new_[46660]_ , \new_[46663]_ ,
    \new_[46664]_ , \new_[46665]_ , \new_[46669]_ , \new_[46670]_ ,
    \new_[46673]_ , \new_[46676]_ , \new_[46677]_ , \new_[46678]_ ,
    \new_[46682]_ , \new_[46683]_ , \new_[46686]_ , \new_[46689]_ ,
    \new_[46690]_ , \new_[46691]_ , \new_[46695]_ , \new_[46696]_ ,
    \new_[46699]_ , \new_[46702]_ , \new_[46703]_ , \new_[46704]_ ,
    \new_[46708]_ , \new_[46709]_ , \new_[46712]_ , \new_[46715]_ ,
    \new_[46716]_ , \new_[46717]_ , \new_[46721]_ , \new_[46722]_ ,
    \new_[46725]_ , \new_[46728]_ , \new_[46729]_ , \new_[46730]_ ,
    \new_[46734]_ , \new_[46735]_ , \new_[46738]_ , \new_[46741]_ ,
    \new_[46742]_ , \new_[46743]_ , \new_[46747]_ , \new_[46748]_ ,
    \new_[46751]_ , \new_[46754]_ , \new_[46755]_ , \new_[46756]_ ,
    \new_[46760]_ , \new_[46761]_ , \new_[46764]_ , \new_[46767]_ ,
    \new_[46768]_ , \new_[46769]_ , \new_[46773]_ , \new_[46774]_ ,
    \new_[46777]_ , \new_[46780]_ , \new_[46781]_ , \new_[46782]_ ,
    \new_[46786]_ , \new_[46787]_ , \new_[46790]_ , \new_[46793]_ ,
    \new_[46794]_ , \new_[46795]_ , \new_[46799]_ , \new_[46800]_ ,
    \new_[46803]_ , \new_[46806]_ , \new_[46807]_ , \new_[46808]_ ,
    \new_[46812]_ , \new_[46813]_ , \new_[46816]_ , \new_[46819]_ ,
    \new_[46820]_ , \new_[46821]_ , \new_[46825]_ , \new_[46826]_ ,
    \new_[46829]_ , \new_[46832]_ , \new_[46833]_ , \new_[46834]_ ,
    \new_[46838]_ , \new_[46839]_ , \new_[46842]_ , \new_[46845]_ ,
    \new_[46846]_ , \new_[46847]_ , \new_[46851]_ , \new_[46852]_ ,
    \new_[46855]_ , \new_[46858]_ , \new_[46859]_ , \new_[46860]_ ,
    \new_[46864]_ , \new_[46865]_ , \new_[46868]_ , \new_[46871]_ ,
    \new_[46872]_ , \new_[46873]_ , \new_[46877]_ , \new_[46878]_ ,
    \new_[46881]_ , \new_[46884]_ , \new_[46885]_ , \new_[46886]_ ,
    \new_[46890]_ , \new_[46891]_ , \new_[46894]_ , \new_[46897]_ ,
    \new_[46898]_ , \new_[46899]_ , \new_[46903]_ , \new_[46904]_ ,
    \new_[46907]_ , \new_[46910]_ , \new_[46911]_ , \new_[46912]_ ,
    \new_[46916]_ , \new_[46917]_ , \new_[46920]_ , \new_[46923]_ ,
    \new_[46924]_ , \new_[46925]_ , \new_[46929]_ , \new_[46930]_ ,
    \new_[46933]_ , \new_[46936]_ , \new_[46937]_ , \new_[46938]_ ,
    \new_[46942]_ , \new_[46943]_ , \new_[46946]_ , \new_[46949]_ ,
    \new_[46950]_ , \new_[46951]_ , \new_[46955]_ , \new_[46956]_ ,
    \new_[46959]_ , \new_[46962]_ , \new_[46963]_ , \new_[46964]_ ,
    \new_[46968]_ , \new_[46969]_ , \new_[46972]_ , \new_[46975]_ ,
    \new_[46976]_ , \new_[46977]_ , \new_[46981]_ , \new_[46982]_ ,
    \new_[46985]_ , \new_[46988]_ , \new_[46989]_ , \new_[46990]_ ,
    \new_[46994]_ , \new_[46995]_ , \new_[46998]_ , \new_[47001]_ ,
    \new_[47002]_ , \new_[47003]_ , \new_[47007]_ , \new_[47008]_ ,
    \new_[47011]_ , \new_[47014]_ , \new_[47015]_ , \new_[47016]_ ,
    \new_[47020]_ , \new_[47021]_ , \new_[47024]_ , \new_[47027]_ ,
    \new_[47028]_ , \new_[47029]_ , \new_[47033]_ , \new_[47034]_ ,
    \new_[47037]_ , \new_[47040]_ , \new_[47041]_ , \new_[47042]_ ,
    \new_[47046]_ , \new_[47047]_ , \new_[47050]_ , \new_[47053]_ ,
    \new_[47054]_ , \new_[47055]_ , \new_[47059]_ , \new_[47060]_ ,
    \new_[47063]_ , \new_[47066]_ , \new_[47067]_ , \new_[47068]_ ,
    \new_[47072]_ , \new_[47073]_ , \new_[47076]_ , \new_[47079]_ ,
    \new_[47080]_ , \new_[47081]_ , \new_[47085]_ , \new_[47086]_ ,
    \new_[47089]_ , \new_[47092]_ , \new_[47093]_ , \new_[47094]_ ,
    \new_[47098]_ , \new_[47099]_ , \new_[47102]_ , \new_[47105]_ ,
    \new_[47106]_ , \new_[47107]_ , \new_[47111]_ , \new_[47112]_ ,
    \new_[47115]_ , \new_[47118]_ , \new_[47119]_ , \new_[47120]_ ,
    \new_[47124]_ , \new_[47125]_ , \new_[47128]_ , \new_[47131]_ ,
    \new_[47132]_ , \new_[47133]_ , \new_[47137]_ , \new_[47138]_ ,
    \new_[47141]_ , \new_[47144]_ , \new_[47145]_ , \new_[47146]_ ,
    \new_[47150]_ , \new_[47151]_ , \new_[47154]_ , \new_[47157]_ ,
    \new_[47158]_ , \new_[47159]_ , \new_[47163]_ , \new_[47164]_ ,
    \new_[47167]_ , \new_[47170]_ , \new_[47171]_ , \new_[47172]_ ,
    \new_[47176]_ , \new_[47177]_ , \new_[47180]_ , \new_[47183]_ ,
    \new_[47184]_ , \new_[47185]_ , \new_[47189]_ , \new_[47190]_ ,
    \new_[47193]_ , \new_[47196]_ , \new_[47197]_ , \new_[47198]_ ,
    \new_[47202]_ , \new_[47203]_ , \new_[47206]_ , \new_[47209]_ ,
    \new_[47210]_ , \new_[47211]_ , \new_[47215]_ , \new_[47216]_ ,
    \new_[47219]_ , \new_[47222]_ , \new_[47223]_ , \new_[47224]_ ,
    \new_[47228]_ , \new_[47229]_ , \new_[47232]_ , \new_[47235]_ ,
    \new_[47236]_ , \new_[47237]_ , \new_[47241]_ , \new_[47242]_ ,
    \new_[47245]_ , \new_[47248]_ , \new_[47249]_ , \new_[47250]_ ,
    \new_[47254]_ , \new_[47255]_ , \new_[47258]_ , \new_[47261]_ ,
    \new_[47262]_ , \new_[47263]_ , \new_[47267]_ , \new_[47268]_ ,
    \new_[47271]_ , \new_[47274]_ , \new_[47275]_ , \new_[47276]_ ,
    \new_[47280]_ , \new_[47281]_ , \new_[47284]_ , \new_[47287]_ ,
    \new_[47288]_ , \new_[47289]_ , \new_[47293]_ , \new_[47294]_ ,
    \new_[47297]_ , \new_[47300]_ , \new_[47301]_ , \new_[47302]_ ,
    \new_[47306]_ , \new_[47307]_ , \new_[47310]_ , \new_[47313]_ ,
    \new_[47314]_ , \new_[47315]_ , \new_[47319]_ , \new_[47320]_ ,
    \new_[47323]_ , \new_[47326]_ , \new_[47327]_ , \new_[47328]_ ,
    \new_[47332]_ , \new_[47333]_ , \new_[47336]_ , \new_[47339]_ ,
    \new_[47340]_ , \new_[47341]_ , \new_[47345]_ , \new_[47346]_ ,
    \new_[47349]_ , \new_[47352]_ , \new_[47353]_ , \new_[47354]_ ,
    \new_[47358]_ , \new_[47359]_ , \new_[47362]_ , \new_[47365]_ ,
    \new_[47366]_ , \new_[47367]_ , \new_[47371]_ , \new_[47372]_ ,
    \new_[47375]_ , \new_[47378]_ , \new_[47379]_ , \new_[47380]_ ,
    \new_[47384]_ , \new_[47385]_ , \new_[47388]_ , \new_[47391]_ ,
    \new_[47392]_ , \new_[47393]_ , \new_[47397]_ , \new_[47398]_ ,
    \new_[47401]_ , \new_[47404]_ , \new_[47405]_ , \new_[47406]_ ,
    \new_[47410]_ , \new_[47411]_ , \new_[47414]_ , \new_[47417]_ ,
    \new_[47418]_ , \new_[47419]_ , \new_[47423]_ , \new_[47424]_ ,
    \new_[47427]_ , \new_[47430]_ , \new_[47431]_ , \new_[47432]_ ,
    \new_[47436]_ , \new_[47437]_ , \new_[47440]_ , \new_[47443]_ ,
    \new_[47444]_ , \new_[47445]_ , \new_[47449]_ , \new_[47450]_ ,
    \new_[47453]_ , \new_[47456]_ , \new_[47457]_ , \new_[47458]_ ,
    \new_[47462]_ , \new_[47463]_ , \new_[47466]_ , \new_[47469]_ ,
    \new_[47470]_ , \new_[47471]_ , \new_[47475]_ , \new_[47476]_ ,
    \new_[47479]_ , \new_[47482]_ , \new_[47483]_ , \new_[47484]_ ,
    \new_[47488]_ , \new_[47489]_ , \new_[47492]_ , \new_[47495]_ ,
    \new_[47496]_ , \new_[47497]_ , \new_[47501]_ , \new_[47502]_ ,
    \new_[47505]_ , \new_[47508]_ , \new_[47509]_ , \new_[47510]_ ,
    \new_[47514]_ , \new_[47515]_ , \new_[47518]_ , \new_[47521]_ ,
    \new_[47522]_ , \new_[47523]_ , \new_[47527]_ , \new_[47528]_ ,
    \new_[47531]_ , \new_[47534]_ , \new_[47535]_ , \new_[47536]_ ,
    \new_[47540]_ , \new_[47541]_ , \new_[47544]_ , \new_[47547]_ ,
    \new_[47548]_ , \new_[47549]_ , \new_[47553]_ , \new_[47554]_ ,
    \new_[47557]_ , \new_[47560]_ , \new_[47561]_ , \new_[47562]_ ,
    \new_[47566]_ , \new_[47567]_ , \new_[47570]_ , \new_[47573]_ ,
    \new_[47574]_ , \new_[47575]_ , \new_[47579]_ , \new_[47580]_ ,
    \new_[47583]_ , \new_[47586]_ , \new_[47587]_ , \new_[47588]_ ,
    \new_[47592]_ , \new_[47593]_ , \new_[47596]_ , \new_[47599]_ ,
    \new_[47600]_ , \new_[47601]_ , \new_[47605]_ , \new_[47606]_ ,
    \new_[47609]_ , \new_[47612]_ , \new_[47613]_ , \new_[47614]_ ,
    \new_[47618]_ , \new_[47619]_ , \new_[47622]_ , \new_[47625]_ ,
    \new_[47626]_ , \new_[47627]_ , \new_[47631]_ , \new_[47632]_ ,
    \new_[47635]_ , \new_[47638]_ , \new_[47639]_ , \new_[47640]_ ,
    \new_[47644]_ , \new_[47645]_ , \new_[47648]_ , \new_[47651]_ ,
    \new_[47652]_ , \new_[47653]_ , \new_[47657]_ , \new_[47658]_ ,
    \new_[47661]_ , \new_[47664]_ , \new_[47665]_ , \new_[47666]_ ,
    \new_[47670]_ , \new_[47671]_ , \new_[47674]_ , \new_[47677]_ ,
    \new_[47678]_ , \new_[47679]_ , \new_[47683]_ , \new_[47684]_ ,
    \new_[47687]_ , \new_[47690]_ , \new_[47691]_ , \new_[47692]_ ,
    \new_[47696]_ , \new_[47697]_ , \new_[47700]_ , \new_[47703]_ ,
    \new_[47704]_ , \new_[47705]_ , \new_[47709]_ , \new_[47710]_ ,
    \new_[47713]_ , \new_[47716]_ , \new_[47717]_ , \new_[47718]_ ,
    \new_[47722]_ , \new_[47723]_ , \new_[47726]_ , \new_[47729]_ ,
    \new_[47730]_ , \new_[47731]_ , \new_[47735]_ , \new_[47736]_ ,
    \new_[47739]_ , \new_[47742]_ , \new_[47743]_ , \new_[47744]_ ,
    \new_[47748]_ , \new_[47749]_ , \new_[47752]_ , \new_[47755]_ ,
    \new_[47756]_ , \new_[47757]_ , \new_[47761]_ , \new_[47762]_ ,
    \new_[47765]_ , \new_[47768]_ , \new_[47769]_ , \new_[47770]_ ,
    \new_[47774]_ , \new_[47775]_ , \new_[47778]_ , \new_[47781]_ ,
    \new_[47782]_ , \new_[47783]_ , \new_[47787]_ , \new_[47788]_ ,
    \new_[47791]_ , \new_[47794]_ , \new_[47795]_ , \new_[47796]_ ,
    \new_[47800]_ , \new_[47801]_ , \new_[47804]_ , \new_[47807]_ ,
    \new_[47808]_ , \new_[47809]_ , \new_[47813]_ , \new_[47814]_ ,
    \new_[47817]_ , \new_[47820]_ , \new_[47821]_ , \new_[47822]_ ,
    \new_[47826]_ , \new_[47827]_ , \new_[47830]_ , \new_[47833]_ ,
    \new_[47834]_ , \new_[47835]_ , \new_[47839]_ , \new_[47840]_ ,
    \new_[47843]_ , \new_[47846]_ , \new_[47847]_ , \new_[47848]_ ,
    \new_[47852]_ , \new_[47853]_ , \new_[47856]_ , \new_[47859]_ ,
    \new_[47860]_ , \new_[47861]_ , \new_[47865]_ , \new_[47866]_ ,
    \new_[47869]_ , \new_[47872]_ , \new_[47873]_ , \new_[47874]_ ,
    \new_[47878]_ , \new_[47879]_ , \new_[47882]_ , \new_[47885]_ ,
    \new_[47886]_ , \new_[47887]_ , \new_[47891]_ , \new_[47892]_ ,
    \new_[47895]_ , \new_[47898]_ , \new_[47899]_ , \new_[47900]_ ,
    \new_[47904]_ , \new_[47905]_ , \new_[47908]_ , \new_[47911]_ ,
    \new_[47912]_ , \new_[47913]_ , \new_[47917]_ , \new_[47918]_ ,
    \new_[47921]_ , \new_[47924]_ , \new_[47925]_ , \new_[47926]_ ,
    \new_[47930]_ , \new_[47931]_ , \new_[47934]_ , \new_[47937]_ ,
    \new_[47938]_ , \new_[47939]_ , \new_[47943]_ , \new_[47944]_ ,
    \new_[47947]_ , \new_[47950]_ , \new_[47951]_ , \new_[47952]_ ,
    \new_[47956]_ , \new_[47957]_ , \new_[47960]_ , \new_[47963]_ ,
    \new_[47964]_ , \new_[47965]_ , \new_[47969]_ , \new_[47970]_ ,
    \new_[47973]_ , \new_[47976]_ , \new_[47977]_ , \new_[47978]_ ,
    \new_[47982]_ , \new_[47983]_ , \new_[47986]_ , \new_[47989]_ ,
    \new_[47990]_ , \new_[47991]_ , \new_[47995]_ , \new_[47996]_ ,
    \new_[47999]_ , \new_[48002]_ , \new_[48003]_ , \new_[48004]_ ,
    \new_[48008]_ , \new_[48009]_ , \new_[48012]_ , \new_[48015]_ ,
    \new_[48016]_ , \new_[48017]_ , \new_[48021]_ , \new_[48022]_ ,
    \new_[48025]_ , \new_[48028]_ , \new_[48029]_ , \new_[48030]_ ,
    \new_[48034]_ , \new_[48035]_ , \new_[48038]_ , \new_[48041]_ ,
    \new_[48042]_ , \new_[48043]_ , \new_[48047]_ , \new_[48048]_ ,
    \new_[48051]_ , \new_[48054]_ , \new_[48055]_ , \new_[48056]_ ,
    \new_[48060]_ , \new_[48061]_ , \new_[48064]_ , \new_[48067]_ ,
    \new_[48068]_ , \new_[48069]_ , \new_[48073]_ , \new_[48074]_ ,
    \new_[48077]_ , \new_[48080]_ , \new_[48081]_ , \new_[48082]_ ,
    \new_[48086]_ , \new_[48087]_ , \new_[48090]_ , \new_[48093]_ ,
    \new_[48094]_ , \new_[48095]_ , \new_[48099]_ , \new_[48100]_ ,
    \new_[48103]_ , \new_[48106]_ , \new_[48107]_ , \new_[48108]_ ,
    \new_[48112]_ , \new_[48113]_ , \new_[48116]_ , \new_[48119]_ ,
    \new_[48120]_ , \new_[48121]_ , \new_[48125]_ , \new_[48126]_ ,
    \new_[48129]_ , \new_[48132]_ , \new_[48133]_ , \new_[48134]_ ,
    \new_[48138]_ , \new_[48139]_ , \new_[48142]_ , \new_[48145]_ ,
    \new_[48146]_ , \new_[48147]_ , \new_[48151]_ , \new_[48152]_ ,
    \new_[48155]_ , \new_[48158]_ , \new_[48159]_ , \new_[48160]_ ,
    \new_[48164]_ , \new_[48165]_ , \new_[48168]_ , \new_[48171]_ ,
    \new_[48172]_ , \new_[48173]_ , \new_[48177]_ , \new_[48178]_ ,
    \new_[48181]_ , \new_[48184]_ , \new_[48185]_ , \new_[48186]_ ,
    \new_[48190]_ , \new_[48191]_ , \new_[48194]_ , \new_[48197]_ ,
    \new_[48198]_ , \new_[48199]_ , \new_[48203]_ , \new_[48204]_ ,
    \new_[48207]_ , \new_[48210]_ , \new_[48211]_ , \new_[48212]_ ,
    \new_[48216]_ , \new_[48217]_ , \new_[48220]_ , \new_[48223]_ ,
    \new_[48224]_ , \new_[48225]_ , \new_[48229]_ , \new_[48230]_ ,
    \new_[48233]_ , \new_[48236]_ , \new_[48237]_ , \new_[48238]_ ,
    \new_[48242]_ , \new_[48243]_ , \new_[48246]_ , \new_[48249]_ ,
    \new_[48250]_ , \new_[48251]_ , \new_[48255]_ , \new_[48256]_ ,
    \new_[48259]_ , \new_[48262]_ , \new_[48263]_ , \new_[48264]_ ,
    \new_[48268]_ , \new_[48269]_ , \new_[48272]_ , \new_[48275]_ ,
    \new_[48276]_ , \new_[48277]_ , \new_[48281]_ , \new_[48282]_ ,
    \new_[48285]_ , \new_[48288]_ , \new_[48289]_ , \new_[48290]_ ,
    \new_[48294]_ , \new_[48295]_ , \new_[48298]_ , \new_[48301]_ ,
    \new_[48302]_ , \new_[48303]_ , \new_[48307]_ , \new_[48308]_ ,
    \new_[48311]_ , \new_[48314]_ , \new_[48315]_ , \new_[48316]_ ,
    \new_[48320]_ , \new_[48321]_ , \new_[48324]_ , \new_[48327]_ ,
    \new_[48328]_ , \new_[48329]_ , \new_[48333]_ , \new_[48334]_ ,
    \new_[48337]_ , \new_[48340]_ , \new_[48341]_ , \new_[48342]_ ,
    \new_[48346]_ , \new_[48347]_ , \new_[48350]_ , \new_[48353]_ ,
    \new_[48354]_ , \new_[48355]_ , \new_[48359]_ , \new_[48360]_ ,
    \new_[48363]_ , \new_[48366]_ , \new_[48367]_ , \new_[48368]_ ,
    \new_[48372]_ , \new_[48373]_ , \new_[48376]_ , \new_[48379]_ ,
    \new_[48380]_ , \new_[48381]_ , \new_[48385]_ , \new_[48386]_ ,
    \new_[48389]_ , \new_[48392]_ , \new_[48393]_ , \new_[48394]_ ,
    \new_[48398]_ , \new_[48399]_ , \new_[48402]_ , \new_[48405]_ ,
    \new_[48406]_ , \new_[48407]_ , \new_[48411]_ , \new_[48412]_ ,
    \new_[48415]_ , \new_[48418]_ , \new_[48419]_ , \new_[48420]_ ,
    \new_[48424]_ , \new_[48425]_ , \new_[48428]_ , \new_[48431]_ ,
    \new_[48432]_ , \new_[48433]_ , \new_[48437]_ , \new_[48438]_ ,
    \new_[48441]_ , \new_[48444]_ , \new_[48445]_ , \new_[48446]_ ,
    \new_[48450]_ , \new_[48451]_ , \new_[48454]_ , \new_[48457]_ ,
    \new_[48458]_ , \new_[48459]_ , \new_[48463]_ , \new_[48464]_ ,
    \new_[48467]_ , \new_[48470]_ , \new_[48471]_ , \new_[48472]_ ,
    \new_[48476]_ , \new_[48477]_ , \new_[48480]_ , \new_[48483]_ ,
    \new_[48484]_ , \new_[48485]_ , \new_[48489]_ , \new_[48490]_ ,
    \new_[48493]_ , \new_[48496]_ , \new_[48497]_ , \new_[48498]_ ,
    \new_[48502]_ , \new_[48503]_ , \new_[48506]_ , \new_[48509]_ ,
    \new_[48510]_ , \new_[48511]_ , \new_[48515]_ , \new_[48516]_ ,
    \new_[48519]_ , \new_[48522]_ , \new_[48523]_ , \new_[48524]_ ,
    \new_[48528]_ , \new_[48529]_ , \new_[48532]_ , \new_[48535]_ ,
    \new_[48536]_ , \new_[48537]_ , \new_[48541]_ , \new_[48542]_ ,
    \new_[48545]_ , \new_[48548]_ , \new_[48549]_ , \new_[48550]_ ,
    \new_[48554]_ , \new_[48555]_ , \new_[48558]_ , \new_[48561]_ ,
    \new_[48562]_ , \new_[48563]_ , \new_[48567]_ , \new_[48568]_ ,
    \new_[48571]_ , \new_[48574]_ , \new_[48575]_ , \new_[48576]_ ,
    \new_[48580]_ , \new_[48581]_ , \new_[48584]_ , \new_[48587]_ ,
    \new_[48588]_ , \new_[48589]_ , \new_[48593]_ , \new_[48594]_ ,
    \new_[48597]_ , \new_[48600]_ , \new_[48601]_ , \new_[48602]_ ,
    \new_[48606]_ , \new_[48607]_ , \new_[48610]_ , \new_[48613]_ ,
    \new_[48614]_ , \new_[48615]_ , \new_[48619]_ , \new_[48620]_ ,
    \new_[48623]_ , \new_[48626]_ , \new_[48627]_ , \new_[48628]_ ,
    \new_[48632]_ , \new_[48633]_ , \new_[48636]_ , \new_[48639]_ ,
    \new_[48640]_ , \new_[48641]_ , \new_[48645]_ , \new_[48646]_ ,
    \new_[48649]_ , \new_[48652]_ , \new_[48653]_ , \new_[48654]_ ,
    \new_[48658]_ , \new_[48659]_ , \new_[48662]_ , \new_[48665]_ ,
    \new_[48666]_ , \new_[48667]_ , \new_[48671]_ , \new_[48672]_ ,
    \new_[48675]_ , \new_[48678]_ , \new_[48679]_ , \new_[48680]_ ,
    \new_[48684]_ , \new_[48685]_ , \new_[48688]_ , \new_[48691]_ ,
    \new_[48692]_ , \new_[48693]_ , \new_[48697]_ , \new_[48698]_ ,
    \new_[48701]_ , \new_[48704]_ , \new_[48705]_ , \new_[48706]_ ,
    \new_[48710]_ , \new_[48711]_ , \new_[48714]_ , \new_[48717]_ ,
    \new_[48718]_ , \new_[48719]_ , \new_[48723]_ , \new_[48724]_ ,
    \new_[48727]_ , \new_[48730]_ , \new_[48731]_ , \new_[48732]_ ,
    \new_[48736]_ , \new_[48737]_ , \new_[48740]_ , \new_[48743]_ ,
    \new_[48744]_ , \new_[48745]_ , \new_[48749]_ , \new_[48750]_ ,
    \new_[48753]_ , \new_[48756]_ , \new_[48757]_ , \new_[48758]_ ,
    \new_[48762]_ , \new_[48763]_ , \new_[48766]_ , \new_[48769]_ ,
    \new_[48770]_ , \new_[48771]_ , \new_[48775]_ , \new_[48776]_ ,
    \new_[48779]_ , \new_[48782]_ , \new_[48783]_ , \new_[48784]_ ,
    \new_[48788]_ , \new_[48789]_ , \new_[48792]_ , \new_[48795]_ ,
    \new_[48796]_ , \new_[48797]_ , \new_[48801]_ , \new_[48802]_ ,
    \new_[48805]_ , \new_[48808]_ , \new_[48809]_ , \new_[48810]_ ,
    \new_[48814]_ , \new_[48815]_ , \new_[48818]_ , \new_[48821]_ ,
    \new_[48822]_ , \new_[48823]_ , \new_[48827]_ , \new_[48828]_ ,
    \new_[48831]_ , \new_[48834]_ , \new_[48835]_ , \new_[48836]_ ,
    \new_[48840]_ , \new_[48841]_ , \new_[48844]_ , \new_[48847]_ ,
    \new_[48848]_ , \new_[48849]_ , \new_[48853]_ , \new_[48854]_ ,
    \new_[48857]_ , \new_[48860]_ , \new_[48861]_ , \new_[48862]_ ,
    \new_[48866]_ , \new_[48867]_ , \new_[48870]_ , \new_[48873]_ ,
    \new_[48874]_ , \new_[48875]_ , \new_[48879]_ , \new_[48880]_ ,
    \new_[48883]_ , \new_[48886]_ , \new_[48887]_ , \new_[48888]_ ,
    \new_[48892]_ , \new_[48893]_ , \new_[48896]_ , \new_[48899]_ ,
    \new_[48900]_ , \new_[48901]_ , \new_[48905]_ , \new_[48906]_ ,
    \new_[48909]_ , \new_[48912]_ , \new_[48913]_ , \new_[48914]_ ,
    \new_[48918]_ , \new_[48919]_ , \new_[48922]_ , \new_[48925]_ ,
    \new_[48926]_ , \new_[48927]_ , \new_[48931]_ , \new_[48932]_ ,
    \new_[48935]_ , \new_[48938]_ , \new_[48939]_ , \new_[48940]_ ,
    \new_[48944]_ , \new_[48945]_ , \new_[48948]_ , \new_[48951]_ ,
    \new_[48952]_ , \new_[48953]_ , \new_[48957]_ , \new_[48958]_ ,
    \new_[48961]_ , \new_[48964]_ , \new_[48965]_ , \new_[48966]_ ,
    \new_[48970]_ , \new_[48971]_ , \new_[48974]_ , \new_[48977]_ ,
    \new_[48978]_ , \new_[48979]_ , \new_[48983]_ , \new_[48984]_ ,
    \new_[48987]_ , \new_[48990]_ , \new_[48991]_ , \new_[48992]_ ,
    \new_[48996]_ , \new_[48997]_ , \new_[49000]_ , \new_[49003]_ ,
    \new_[49004]_ , \new_[49005]_ , \new_[49009]_ , \new_[49010]_ ,
    \new_[49013]_ , \new_[49016]_ , \new_[49017]_ , \new_[49018]_ ,
    \new_[49022]_ , \new_[49023]_ , \new_[49026]_ , \new_[49029]_ ,
    \new_[49030]_ , \new_[49031]_ , \new_[49035]_ , \new_[49036]_ ,
    \new_[49039]_ , \new_[49042]_ , \new_[49043]_ , \new_[49044]_ ,
    \new_[49048]_ , \new_[49049]_ , \new_[49052]_ , \new_[49055]_ ,
    \new_[49056]_ , \new_[49057]_ , \new_[49061]_ , \new_[49062]_ ,
    \new_[49065]_ , \new_[49068]_ , \new_[49069]_ , \new_[49070]_ ,
    \new_[49074]_ , \new_[49075]_ , \new_[49078]_ , \new_[49081]_ ,
    \new_[49082]_ , \new_[49083]_ , \new_[49087]_ , \new_[49088]_ ,
    \new_[49091]_ , \new_[49094]_ , \new_[49095]_ , \new_[49096]_ ,
    \new_[49100]_ , \new_[49101]_ , \new_[49104]_ , \new_[49107]_ ,
    \new_[49108]_ , \new_[49109]_ , \new_[49113]_ , \new_[49114]_ ,
    \new_[49117]_ , \new_[49120]_ , \new_[49121]_ , \new_[49122]_ ,
    \new_[49126]_ , \new_[49127]_ , \new_[49130]_ , \new_[49133]_ ,
    \new_[49134]_ , \new_[49135]_ , \new_[49139]_ , \new_[49140]_ ,
    \new_[49143]_ , \new_[49146]_ , \new_[49147]_ , \new_[49148]_ ,
    \new_[49152]_ , \new_[49153]_ , \new_[49156]_ , \new_[49159]_ ,
    \new_[49160]_ , \new_[49161]_ , \new_[49165]_ , \new_[49166]_ ,
    \new_[49169]_ , \new_[49172]_ , \new_[49173]_ , \new_[49174]_ ,
    \new_[49178]_ , \new_[49179]_ , \new_[49182]_ , \new_[49185]_ ,
    \new_[49186]_ , \new_[49187]_ , \new_[49191]_ , \new_[49192]_ ,
    \new_[49195]_ , \new_[49198]_ , \new_[49199]_ , \new_[49200]_ ,
    \new_[49204]_ , \new_[49205]_ , \new_[49208]_ , \new_[49211]_ ,
    \new_[49212]_ , \new_[49213]_ , \new_[49217]_ , \new_[49218]_ ,
    \new_[49221]_ , \new_[49224]_ , \new_[49225]_ , \new_[49226]_ ,
    \new_[49230]_ , \new_[49231]_ , \new_[49234]_ , \new_[49237]_ ,
    \new_[49238]_ , \new_[49239]_ , \new_[49243]_ , \new_[49244]_ ,
    \new_[49247]_ , \new_[49250]_ , \new_[49251]_ , \new_[49252]_ ,
    \new_[49256]_ , \new_[49257]_ , \new_[49260]_ , \new_[49263]_ ,
    \new_[49264]_ , \new_[49265]_ , \new_[49269]_ , \new_[49270]_ ,
    \new_[49273]_ , \new_[49276]_ , \new_[49277]_ , \new_[49278]_ ,
    \new_[49282]_ , \new_[49283]_ , \new_[49286]_ , \new_[49289]_ ,
    \new_[49290]_ , \new_[49291]_ , \new_[49295]_ , \new_[49296]_ ,
    \new_[49299]_ , \new_[49302]_ , \new_[49303]_ , \new_[49304]_ ,
    \new_[49308]_ , \new_[49309]_ , \new_[49312]_ , \new_[49315]_ ,
    \new_[49316]_ , \new_[49317]_ , \new_[49321]_ , \new_[49322]_ ,
    \new_[49325]_ , \new_[49328]_ , \new_[49329]_ , \new_[49330]_ ,
    \new_[49334]_ , \new_[49335]_ , \new_[49338]_ , \new_[49341]_ ,
    \new_[49342]_ , \new_[49343]_ , \new_[49347]_ , \new_[49348]_ ,
    \new_[49351]_ , \new_[49354]_ , \new_[49355]_ , \new_[49356]_ ,
    \new_[49360]_ , \new_[49361]_ , \new_[49364]_ , \new_[49367]_ ,
    \new_[49368]_ , \new_[49369]_ , \new_[49373]_ , \new_[49374]_ ,
    \new_[49377]_ , \new_[49380]_ , \new_[49381]_ , \new_[49382]_ ,
    \new_[49386]_ , \new_[49387]_ , \new_[49390]_ , \new_[49393]_ ,
    \new_[49394]_ , \new_[49395]_ , \new_[49399]_ , \new_[49400]_ ,
    \new_[49403]_ , \new_[49406]_ , \new_[49407]_ , \new_[49408]_ ,
    \new_[49412]_ , \new_[49413]_ , \new_[49416]_ , \new_[49419]_ ,
    \new_[49420]_ , \new_[49421]_ , \new_[49425]_ , \new_[49426]_ ,
    \new_[49429]_ , \new_[49432]_ , \new_[49433]_ , \new_[49434]_ ,
    \new_[49438]_ , \new_[49439]_ , \new_[49442]_ , \new_[49445]_ ,
    \new_[49446]_ , \new_[49447]_ , \new_[49451]_ , \new_[49452]_ ,
    \new_[49455]_ , \new_[49458]_ , \new_[49459]_ , \new_[49460]_ ,
    \new_[49464]_ , \new_[49465]_ , \new_[49468]_ , \new_[49471]_ ,
    \new_[49472]_ , \new_[49473]_ , \new_[49477]_ , \new_[49478]_ ,
    \new_[49481]_ , \new_[49484]_ , \new_[49485]_ , \new_[49486]_ ,
    \new_[49490]_ , \new_[49491]_ , \new_[49494]_ , \new_[49497]_ ,
    \new_[49498]_ , \new_[49499]_ , \new_[49503]_ , \new_[49504]_ ,
    \new_[49507]_ , \new_[49510]_ , \new_[49511]_ , \new_[49512]_ ,
    \new_[49516]_ , \new_[49517]_ , \new_[49520]_ , \new_[49523]_ ,
    \new_[49524]_ , \new_[49525]_ , \new_[49529]_ , \new_[49530]_ ,
    \new_[49533]_ , \new_[49536]_ , \new_[49537]_ , \new_[49538]_ ,
    \new_[49542]_ , \new_[49543]_ , \new_[49546]_ , \new_[49549]_ ,
    \new_[49550]_ , \new_[49551]_ , \new_[49555]_ , \new_[49556]_ ,
    \new_[49559]_ , \new_[49562]_ , \new_[49563]_ , \new_[49564]_ ,
    \new_[49568]_ , \new_[49569]_ , \new_[49572]_ , \new_[49575]_ ,
    \new_[49576]_ , \new_[49577]_ , \new_[49581]_ , \new_[49582]_ ,
    \new_[49585]_ , \new_[49588]_ , \new_[49589]_ , \new_[49590]_ ,
    \new_[49594]_ , \new_[49595]_ , \new_[49598]_ , \new_[49601]_ ,
    \new_[49602]_ , \new_[49603]_ , \new_[49607]_ , \new_[49608]_ ,
    \new_[49611]_ , \new_[49614]_ , \new_[49615]_ , \new_[49616]_ ,
    \new_[49620]_ , \new_[49621]_ , \new_[49624]_ , \new_[49627]_ ,
    \new_[49628]_ , \new_[49629]_ , \new_[49633]_ , \new_[49634]_ ,
    \new_[49637]_ , \new_[49640]_ , \new_[49641]_ , \new_[49642]_ ,
    \new_[49646]_ , \new_[49647]_ , \new_[49650]_ , \new_[49653]_ ,
    \new_[49654]_ , \new_[49655]_ , \new_[49659]_ , \new_[49660]_ ,
    \new_[49663]_ , \new_[49666]_ , \new_[49667]_ , \new_[49668]_ ,
    \new_[49672]_ , \new_[49673]_ , \new_[49676]_ , \new_[49679]_ ,
    \new_[49680]_ , \new_[49681]_ , \new_[49685]_ , \new_[49686]_ ,
    \new_[49689]_ , \new_[49692]_ , \new_[49693]_ , \new_[49694]_ ,
    \new_[49698]_ , \new_[49699]_ , \new_[49702]_ , \new_[49705]_ ,
    \new_[49706]_ , \new_[49707]_ , \new_[49711]_ , \new_[49712]_ ,
    \new_[49715]_ , \new_[49718]_ , \new_[49719]_ , \new_[49720]_ ,
    \new_[49724]_ , \new_[49725]_ , \new_[49728]_ , \new_[49731]_ ,
    \new_[49732]_ , \new_[49733]_ , \new_[49737]_ , \new_[49738]_ ,
    \new_[49741]_ , \new_[49744]_ , \new_[49745]_ , \new_[49746]_ ,
    \new_[49750]_ , \new_[49751]_ , \new_[49754]_ , \new_[49757]_ ,
    \new_[49758]_ , \new_[49759]_ , \new_[49763]_ , \new_[49764]_ ,
    \new_[49767]_ , \new_[49770]_ , \new_[49771]_ , \new_[49772]_ ,
    \new_[49776]_ , \new_[49777]_ , \new_[49780]_ , \new_[49783]_ ,
    \new_[49784]_ , \new_[49785]_ , \new_[49789]_ , \new_[49790]_ ,
    \new_[49793]_ , \new_[49796]_ , \new_[49797]_ , \new_[49798]_ ,
    \new_[49802]_ , \new_[49803]_ , \new_[49806]_ , \new_[49809]_ ,
    \new_[49810]_ , \new_[49811]_ , \new_[49815]_ , \new_[49816]_ ,
    \new_[49819]_ , \new_[49822]_ , \new_[49823]_ , \new_[49824]_ ,
    \new_[49828]_ , \new_[49829]_ , \new_[49832]_ , \new_[49835]_ ,
    \new_[49836]_ , \new_[49837]_ , \new_[49841]_ , \new_[49842]_ ,
    \new_[49845]_ , \new_[49848]_ , \new_[49849]_ , \new_[49850]_ ,
    \new_[49854]_ , \new_[49855]_ , \new_[49858]_ , \new_[49861]_ ,
    \new_[49862]_ , \new_[49863]_ , \new_[49867]_ , \new_[49868]_ ,
    \new_[49871]_ , \new_[49874]_ , \new_[49875]_ , \new_[49876]_ ,
    \new_[49880]_ , \new_[49881]_ , \new_[49884]_ , \new_[49887]_ ,
    \new_[49888]_ , \new_[49889]_ , \new_[49893]_ , \new_[49894]_ ,
    \new_[49897]_ , \new_[49900]_ , \new_[49901]_ , \new_[49902]_ ,
    \new_[49906]_ , \new_[49907]_ , \new_[49910]_ , \new_[49913]_ ,
    \new_[49914]_ , \new_[49915]_ , \new_[49919]_ , \new_[49920]_ ,
    \new_[49923]_ , \new_[49926]_ , \new_[49927]_ , \new_[49928]_ ,
    \new_[49932]_ , \new_[49933]_ , \new_[49936]_ , \new_[49939]_ ,
    \new_[49940]_ , \new_[49941]_ , \new_[49945]_ , \new_[49946]_ ,
    \new_[49949]_ , \new_[49952]_ , \new_[49953]_ , \new_[49954]_ ,
    \new_[49958]_ , \new_[49959]_ , \new_[49962]_ , \new_[49965]_ ,
    \new_[49966]_ , \new_[49967]_ , \new_[49971]_ , \new_[49972]_ ,
    \new_[49975]_ , \new_[49978]_ , \new_[49979]_ , \new_[49980]_ ,
    \new_[49984]_ , \new_[49985]_ , \new_[49988]_ , \new_[49991]_ ,
    \new_[49992]_ , \new_[49993]_ , \new_[49997]_ , \new_[49998]_ ,
    \new_[50001]_ , \new_[50004]_ , \new_[50005]_ , \new_[50006]_ ,
    \new_[50010]_ , \new_[50011]_ , \new_[50014]_ , \new_[50017]_ ,
    \new_[50018]_ , \new_[50019]_ , \new_[50023]_ , \new_[50024]_ ,
    \new_[50027]_ , \new_[50030]_ , \new_[50031]_ , \new_[50032]_ ,
    \new_[50036]_ , \new_[50037]_ , \new_[50040]_ , \new_[50043]_ ,
    \new_[50044]_ , \new_[50045]_ , \new_[50049]_ , \new_[50050]_ ,
    \new_[50053]_ , \new_[50056]_ , \new_[50057]_ , \new_[50058]_ ,
    \new_[50062]_ , \new_[50063]_ , \new_[50066]_ , \new_[50069]_ ,
    \new_[50070]_ , \new_[50071]_ , \new_[50075]_ , \new_[50076]_ ,
    \new_[50079]_ , \new_[50082]_ , \new_[50083]_ , \new_[50084]_ ,
    \new_[50088]_ , \new_[50089]_ , \new_[50092]_ , \new_[50095]_ ,
    \new_[50096]_ , \new_[50097]_ , \new_[50101]_ , \new_[50102]_ ,
    \new_[50105]_ , \new_[50108]_ , \new_[50109]_ , \new_[50110]_ ,
    \new_[50114]_ , \new_[50115]_ , \new_[50118]_ , \new_[50121]_ ,
    \new_[50122]_ , \new_[50123]_ , \new_[50127]_ , \new_[50128]_ ,
    \new_[50131]_ , \new_[50134]_ , \new_[50135]_ , \new_[50136]_ ,
    \new_[50140]_ , \new_[50141]_ , \new_[50144]_ , \new_[50147]_ ,
    \new_[50148]_ , \new_[50149]_ , \new_[50153]_ , \new_[50154]_ ,
    \new_[50157]_ , \new_[50160]_ , \new_[50161]_ , \new_[50162]_ ,
    \new_[50166]_ , \new_[50167]_ , \new_[50170]_ , \new_[50173]_ ,
    \new_[50174]_ , \new_[50175]_ , \new_[50179]_ , \new_[50180]_ ,
    \new_[50183]_ , \new_[50186]_ , \new_[50187]_ , \new_[50188]_ ,
    \new_[50192]_ , \new_[50193]_ , \new_[50196]_ , \new_[50199]_ ,
    \new_[50200]_ , \new_[50201]_ , \new_[50205]_ , \new_[50206]_ ,
    \new_[50209]_ , \new_[50212]_ , \new_[50213]_ , \new_[50214]_ ,
    \new_[50218]_ , \new_[50219]_ , \new_[50222]_ , \new_[50225]_ ,
    \new_[50226]_ , \new_[50227]_ , \new_[50231]_ , \new_[50232]_ ,
    \new_[50235]_ , \new_[50238]_ , \new_[50239]_ , \new_[50240]_ ,
    \new_[50244]_ , \new_[50245]_ , \new_[50248]_ , \new_[50251]_ ,
    \new_[50252]_ , \new_[50253]_ , \new_[50257]_ , \new_[50258]_ ,
    \new_[50261]_ , \new_[50264]_ , \new_[50265]_ , \new_[50266]_ ,
    \new_[50270]_ , \new_[50271]_ , \new_[50274]_ , \new_[50277]_ ,
    \new_[50278]_ , \new_[50279]_ , \new_[50283]_ , \new_[50284]_ ,
    \new_[50287]_ , \new_[50290]_ , \new_[50291]_ , \new_[50292]_ ,
    \new_[50296]_ , \new_[50297]_ , \new_[50300]_ , \new_[50303]_ ,
    \new_[50304]_ , \new_[50305]_ , \new_[50309]_ , \new_[50310]_ ,
    \new_[50313]_ , \new_[50316]_ , \new_[50317]_ , \new_[50318]_ ,
    \new_[50322]_ , \new_[50323]_ , \new_[50326]_ , \new_[50329]_ ,
    \new_[50330]_ , \new_[50331]_ , \new_[50335]_ , \new_[50336]_ ,
    \new_[50339]_ , \new_[50342]_ , \new_[50343]_ , \new_[50344]_ ,
    \new_[50348]_ , \new_[50349]_ , \new_[50352]_ , \new_[50355]_ ,
    \new_[50356]_ , \new_[50357]_ , \new_[50361]_ , \new_[50362]_ ,
    \new_[50365]_ , \new_[50368]_ , \new_[50369]_ , \new_[50370]_ ,
    \new_[50374]_ , \new_[50375]_ , \new_[50378]_ , \new_[50381]_ ,
    \new_[50382]_ , \new_[50383]_ , \new_[50387]_ , \new_[50388]_ ,
    \new_[50391]_ , \new_[50394]_ , \new_[50395]_ , \new_[50396]_ ,
    \new_[50400]_ , \new_[50401]_ , \new_[50404]_ , \new_[50407]_ ,
    \new_[50408]_ , \new_[50409]_ , \new_[50413]_ , \new_[50414]_ ,
    \new_[50417]_ , \new_[50420]_ , \new_[50421]_ , \new_[50422]_ ,
    \new_[50426]_ , \new_[50427]_ , \new_[50430]_ , \new_[50433]_ ,
    \new_[50434]_ , \new_[50435]_ , \new_[50439]_ , \new_[50440]_ ,
    \new_[50443]_ , \new_[50446]_ , \new_[50447]_ , \new_[50448]_ ,
    \new_[50452]_ , \new_[50453]_ , \new_[50456]_ , \new_[50459]_ ,
    \new_[50460]_ , \new_[50461]_ , \new_[50465]_ , \new_[50466]_ ,
    \new_[50469]_ , \new_[50472]_ , \new_[50473]_ , \new_[50474]_ ,
    \new_[50478]_ , \new_[50479]_ , \new_[50482]_ , \new_[50485]_ ,
    \new_[50486]_ , \new_[50487]_ , \new_[50491]_ , \new_[50492]_ ,
    \new_[50495]_ , \new_[50498]_ , \new_[50499]_ , \new_[50500]_ ,
    \new_[50504]_ , \new_[50505]_ , \new_[50508]_ , \new_[50511]_ ,
    \new_[50512]_ , \new_[50513]_ , \new_[50517]_ , \new_[50518]_ ,
    \new_[50521]_ , \new_[50524]_ , \new_[50525]_ , \new_[50526]_ ,
    \new_[50530]_ , \new_[50531]_ , \new_[50534]_ , \new_[50537]_ ,
    \new_[50538]_ , \new_[50539]_ , \new_[50543]_ , \new_[50544]_ ,
    \new_[50547]_ , \new_[50550]_ , \new_[50551]_ , \new_[50552]_ ,
    \new_[50556]_ , \new_[50557]_ , \new_[50560]_ , \new_[50563]_ ,
    \new_[50564]_ , \new_[50565]_ , \new_[50569]_ , \new_[50570]_ ,
    \new_[50573]_ , \new_[50576]_ , \new_[50577]_ , \new_[50578]_ ,
    \new_[50582]_ , \new_[50583]_ , \new_[50586]_ , \new_[50589]_ ,
    \new_[50590]_ , \new_[50591]_ , \new_[50595]_ , \new_[50596]_ ,
    \new_[50599]_ , \new_[50602]_ , \new_[50603]_ , \new_[50604]_ ,
    \new_[50608]_ , \new_[50609]_ , \new_[50612]_ , \new_[50615]_ ,
    \new_[50616]_ , \new_[50617]_ , \new_[50621]_ , \new_[50622]_ ,
    \new_[50625]_ , \new_[50628]_ , \new_[50629]_ , \new_[50630]_ ,
    \new_[50634]_ , \new_[50635]_ , \new_[50638]_ , \new_[50641]_ ,
    \new_[50642]_ , \new_[50643]_ , \new_[50647]_ , \new_[50648]_ ,
    \new_[50651]_ , \new_[50654]_ , \new_[50655]_ , \new_[50656]_ ,
    \new_[50660]_ , \new_[50661]_ , \new_[50664]_ , \new_[50667]_ ,
    \new_[50668]_ , \new_[50669]_ , \new_[50673]_ , \new_[50674]_ ,
    \new_[50677]_ , \new_[50680]_ , \new_[50681]_ , \new_[50682]_ ,
    \new_[50686]_ , \new_[50687]_ , \new_[50690]_ , \new_[50693]_ ,
    \new_[50694]_ , \new_[50695]_ , \new_[50699]_ , \new_[50700]_ ,
    \new_[50703]_ , \new_[50706]_ , \new_[50707]_ , \new_[50708]_ ,
    \new_[50712]_ , \new_[50713]_ , \new_[50716]_ , \new_[50719]_ ,
    \new_[50720]_ , \new_[50721]_ , \new_[50725]_ , \new_[50726]_ ,
    \new_[50729]_ , \new_[50732]_ , \new_[50733]_ , \new_[50734]_ ,
    \new_[50738]_ , \new_[50739]_ , \new_[50742]_ , \new_[50745]_ ,
    \new_[50746]_ , \new_[50747]_ , \new_[50751]_ , \new_[50752]_ ,
    \new_[50755]_ , \new_[50758]_ , \new_[50759]_ , \new_[50760]_ ,
    \new_[50764]_ , \new_[50765]_ , \new_[50768]_ , \new_[50771]_ ,
    \new_[50772]_ , \new_[50773]_ , \new_[50777]_ , \new_[50778]_ ,
    \new_[50781]_ , \new_[50784]_ , \new_[50785]_ , \new_[50786]_ ,
    \new_[50790]_ , \new_[50791]_ , \new_[50794]_ , \new_[50797]_ ,
    \new_[50798]_ , \new_[50799]_ , \new_[50803]_ , \new_[50804]_ ,
    \new_[50807]_ , \new_[50810]_ , \new_[50811]_ , \new_[50812]_ ,
    \new_[50816]_ , \new_[50817]_ , \new_[50820]_ , \new_[50823]_ ,
    \new_[50824]_ , \new_[50825]_ , \new_[50829]_ , \new_[50830]_ ,
    \new_[50833]_ , \new_[50836]_ , \new_[50837]_ , \new_[50838]_ ,
    \new_[50842]_ , \new_[50843]_ , \new_[50846]_ , \new_[50849]_ ,
    \new_[50850]_ , \new_[50851]_ , \new_[50855]_ , \new_[50856]_ ,
    \new_[50859]_ , \new_[50862]_ , \new_[50863]_ , \new_[50864]_ ,
    \new_[50868]_ , \new_[50869]_ , \new_[50872]_ , \new_[50875]_ ,
    \new_[50876]_ , \new_[50877]_ , \new_[50881]_ , \new_[50882]_ ,
    \new_[50885]_ , \new_[50888]_ , \new_[50889]_ , \new_[50890]_ ,
    \new_[50894]_ , \new_[50895]_ , \new_[50898]_ , \new_[50901]_ ,
    \new_[50902]_ , \new_[50903]_ , \new_[50907]_ , \new_[50908]_ ,
    \new_[50911]_ , \new_[50914]_ , \new_[50915]_ , \new_[50916]_ ,
    \new_[50920]_ , \new_[50921]_ , \new_[50924]_ , \new_[50927]_ ,
    \new_[50928]_ , \new_[50929]_ , \new_[50933]_ , \new_[50934]_ ,
    \new_[50937]_ , \new_[50940]_ , \new_[50941]_ , \new_[50942]_ ,
    \new_[50946]_ , \new_[50947]_ , \new_[50950]_ , \new_[50953]_ ,
    \new_[50954]_ , \new_[50955]_ , \new_[50959]_ , \new_[50960]_ ,
    \new_[50963]_ , \new_[50966]_ , \new_[50967]_ , \new_[50968]_ ,
    \new_[50972]_ , \new_[50973]_ , \new_[50976]_ , \new_[50979]_ ,
    \new_[50980]_ , \new_[50981]_ , \new_[50985]_ , \new_[50986]_ ,
    \new_[50989]_ , \new_[50992]_ , \new_[50993]_ , \new_[50994]_ ,
    \new_[50998]_ , \new_[50999]_ , \new_[51002]_ , \new_[51005]_ ,
    \new_[51006]_ , \new_[51007]_ , \new_[51011]_ , \new_[51012]_ ,
    \new_[51015]_ , \new_[51018]_ , \new_[51019]_ , \new_[51020]_ ,
    \new_[51024]_ , \new_[51025]_ , \new_[51028]_ , \new_[51031]_ ,
    \new_[51032]_ , \new_[51033]_ , \new_[51037]_ , \new_[51038]_ ,
    \new_[51041]_ , \new_[51044]_ , \new_[51045]_ , \new_[51046]_ ,
    \new_[51050]_ , \new_[51051]_ , \new_[51054]_ , \new_[51057]_ ,
    \new_[51058]_ , \new_[51059]_ , \new_[51063]_ , \new_[51064]_ ,
    \new_[51067]_ , \new_[51070]_ , \new_[51071]_ , \new_[51072]_ ,
    \new_[51076]_ , \new_[51077]_ , \new_[51080]_ , \new_[51083]_ ,
    \new_[51084]_ , \new_[51085]_ , \new_[51089]_ , \new_[51090]_ ,
    \new_[51093]_ , \new_[51096]_ , \new_[51097]_ , \new_[51098]_ ,
    \new_[51102]_ , \new_[51103]_ , \new_[51106]_ , \new_[51109]_ ,
    \new_[51110]_ , \new_[51111]_ , \new_[51115]_ , \new_[51116]_ ,
    \new_[51119]_ , \new_[51122]_ , \new_[51123]_ , \new_[51124]_ ,
    \new_[51128]_ , \new_[51129]_ , \new_[51132]_ , \new_[51135]_ ,
    \new_[51136]_ , \new_[51137]_ , \new_[51141]_ , \new_[51142]_ ,
    \new_[51145]_ , \new_[51148]_ , \new_[51149]_ , \new_[51150]_ ,
    \new_[51154]_ , \new_[51155]_ , \new_[51158]_ , \new_[51161]_ ,
    \new_[51162]_ , \new_[51163]_ , \new_[51167]_ , \new_[51168]_ ,
    \new_[51171]_ , \new_[51174]_ , \new_[51175]_ , \new_[51176]_ ,
    \new_[51180]_ , \new_[51181]_ , \new_[51184]_ , \new_[51187]_ ,
    \new_[51188]_ , \new_[51189]_ , \new_[51193]_ , \new_[51194]_ ,
    \new_[51197]_ , \new_[51200]_ , \new_[51201]_ , \new_[51202]_ ,
    \new_[51206]_ , \new_[51207]_ , \new_[51210]_ , \new_[51213]_ ,
    \new_[51214]_ , \new_[51215]_ , \new_[51219]_ , \new_[51220]_ ,
    \new_[51223]_ , \new_[51226]_ , \new_[51227]_ , \new_[51228]_ ,
    \new_[51232]_ , \new_[51233]_ , \new_[51236]_ , \new_[51239]_ ,
    \new_[51240]_ , \new_[51241]_ , \new_[51245]_ , \new_[51246]_ ,
    \new_[51249]_ , \new_[51252]_ , \new_[51253]_ , \new_[51254]_ ,
    \new_[51258]_ , \new_[51259]_ , \new_[51262]_ , \new_[51265]_ ,
    \new_[51266]_ , \new_[51267]_ , \new_[51271]_ , \new_[51272]_ ,
    \new_[51275]_ , \new_[51278]_ , \new_[51279]_ , \new_[51280]_ ,
    \new_[51284]_ , \new_[51285]_ , \new_[51288]_ , \new_[51291]_ ,
    \new_[51292]_ , \new_[51293]_ , \new_[51297]_ , \new_[51298]_ ,
    \new_[51301]_ , \new_[51304]_ , \new_[51305]_ , \new_[51306]_ ,
    \new_[51310]_ , \new_[51311]_ , \new_[51314]_ , \new_[51317]_ ,
    \new_[51318]_ , \new_[51319]_ , \new_[51323]_ , \new_[51324]_ ,
    \new_[51327]_ , \new_[51330]_ , \new_[51331]_ , \new_[51332]_ ,
    \new_[51336]_ , \new_[51337]_ , \new_[51340]_ , \new_[51343]_ ,
    \new_[51344]_ , \new_[51345]_ , \new_[51349]_ , \new_[51350]_ ,
    \new_[51353]_ , \new_[51356]_ , \new_[51357]_ , \new_[51358]_ ,
    \new_[51362]_ , \new_[51363]_ , \new_[51366]_ , \new_[51369]_ ,
    \new_[51370]_ , \new_[51371]_ , \new_[51375]_ , \new_[51376]_ ,
    \new_[51379]_ , \new_[51382]_ , \new_[51383]_ , \new_[51384]_ ,
    \new_[51388]_ , \new_[51389]_ , \new_[51392]_ , \new_[51395]_ ,
    \new_[51396]_ , \new_[51397]_ , \new_[51401]_ , \new_[51402]_ ,
    \new_[51405]_ , \new_[51408]_ , \new_[51409]_ , \new_[51410]_ ,
    \new_[51414]_ , \new_[51415]_ , \new_[51418]_ , \new_[51421]_ ,
    \new_[51422]_ , \new_[51423]_ , \new_[51427]_ , \new_[51428]_ ,
    \new_[51431]_ , \new_[51434]_ , \new_[51435]_ , \new_[51436]_ ,
    \new_[51440]_ , \new_[51441]_ , \new_[51444]_ , \new_[51447]_ ,
    \new_[51448]_ , \new_[51449]_ , \new_[51453]_ , \new_[51454]_ ,
    \new_[51457]_ , \new_[51460]_ , \new_[51461]_ , \new_[51462]_ ,
    \new_[51466]_ , \new_[51467]_ , \new_[51470]_ , \new_[51473]_ ,
    \new_[51474]_ , \new_[51475]_ , \new_[51479]_ , \new_[51480]_ ,
    \new_[51483]_ , \new_[51486]_ , \new_[51487]_ , \new_[51488]_ ,
    \new_[51492]_ , \new_[51493]_ , \new_[51496]_ , \new_[51499]_ ,
    \new_[51500]_ , \new_[51501]_ , \new_[51505]_ , \new_[51506]_ ,
    \new_[51509]_ , \new_[51512]_ , \new_[51513]_ , \new_[51514]_ ,
    \new_[51518]_ , \new_[51519]_ , \new_[51522]_ , \new_[51525]_ ,
    \new_[51526]_ , \new_[51527]_ , \new_[51531]_ , \new_[51532]_ ,
    \new_[51535]_ , \new_[51538]_ , \new_[51539]_ , \new_[51540]_ ,
    \new_[51544]_ , \new_[51545]_ , \new_[51548]_ , \new_[51551]_ ,
    \new_[51552]_ , \new_[51553]_ , \new_[51557]_ , \new_[51558]_ ,
    \new_[51561]_ , \new_[51564]_ , \new_[51565]_ , \new_[51566]_ ,
    \new_[51570]_ , \new_[51571]_ , \new_[51574]_ , \new_[51577]_ ,
    \new_[51578]_ , \new_[51579]_ , \new_[51583]_ , \new_[51584]_ ,
    \new_[51587]_ , \new_[51590]_ , \new_[51591]_ , \new_[51592]_ ,
    \new_[51596]_ , \new_[51597]_ , \new_[51600]_ , \new_[51603]_ ,
    \new_[51604]_ , \new_[51605]_ , \new_[51609]_ , \new_[51610]_ ,
    \new_[51613]_ , \new_[51616]_ , \new_[51617]_ , \new_[51618]_ ,
    \new_[51622]_ , \new_[51623]_ , \new_[51626]_ , \new_[51629]_ ,
    \new_[51630]_ , \new_[51631]_ , \new_[51635]_ , \new_[51636]_ ,
    \new_[51639]_ , \new_[51642]_ , \new_[51643]_ , \new_[51644]_ ,
    \new_[51648]_ , \new_[51649]_ , \new_[51652]_ , \new_[51655]_ ,
    \new_[51656]_ , \new_[51657]_ , \new_[51661]_ , \new_[51662]_ ,
    \new_[51665]_ , \new_[51668]_ , \new_[51669]_ , \new_[51670]_ ,
    \new_[51674]_ , \new_[51675]_ , \new_[51678]_ , \new_[51681]_ ,
    \new_[51682]_ , \new_[51683]_ , \new_[51687]_ , \new_[51688]_ ,
    \new_[51691]_ , \new_[51694]_ , \new_[51695]_ , \new_[51696]_ ,
    \new_[51700]_ , \new_[51701]_ , \new_[51704]_ , \new_[51707]_ ,
    \new_[51708]_ , \new_[51709]_ , \new_[51713]_ , \new_[51714]_ ,
    \new_[51717]_ , \new_[51720]_ , \new_[51721]_ , \new_[51722]_ ,
    \new_[51726]_ , \new_[51727]_ , \new_[51730]_ , \new_[51733]_ ,
    \new_[51734]_ , \new_[51735]_ , \new_[51739]_ , \new_[51740]_ ,
    \new_[51743]_ , \new_[51746]_ , \new_[51747]_ , \new_[51748]_ ,
    \new_[51752]_ , \new_[51753]_ , \new_[51756]_ , \new_[51759]_ ,
    \new_[51760]_ , \new_[51761]_ , \new_[51765]_ , \new_[51766]_ ,
    \new_[51769]_ , \new_[51772]_ , \new_[51773]_ , \new_[51774]_ ,
    \new_[51778]_ , \new_[51779]_ , \new_[51782]_ , \new_[51785]_ ,
    \new_[51786]_ , \new_[51787]_ , \new_[51791]_ , \new_[51792]_ ,
    \new_[51795]_ , \new_[51798]_ , \new_[51799]_ , \new_[51800]_ ,
    \new_[51804]_ , \new_[51805]_ , \new_[51808]_ , \new_[51811]_ ,
    \new_[51812]_ , \new_[51813]_ , \new_[51817]_ , \new_[51818]_ ,
    \new_[51821]_ , \new_[51824]_ , \new_[51825]_ , \new_[51826]_ ,
    \new_[51830]_ , \new_[51831]_ , \new_[51834]_ , \new_[51837]_ ,
    \new_[51838]_ , \new_[51839]_ , \new_[51843]_ , \new_[51844]_ ,
    \new_[51847]_ , \new_[51850]_ , \new_[51851]_ , \new_[51852]_ ,
    \new_[51856]_ , \new_[51857]_ , \new_[51860]_ , \new_[51863]_ ,
    \new_[51864]_ , \new_[51865]_ , \new_[51869]_ , \new_[51870]_ ,
    \new_[51873]_ , \new_[51876]_ , \new_[51877]_ , \new_[51878]_ ,
    \new_[51882]_ , \new_[51883]_ , \new_[51886]_ , \new_[51889]_ ,
    \new_[51890]_ , \new_[51891]_ , \new_[51895]_ , \new_[51896]_ ,
    \new_[51899]_ , \new_[51902]_ , \new_[51903]_ , \new_[51904]_ ,
    \new_[51908]_ , \new_[51909]_ , \new_[51912]_ , \new_[51915]_ ,
    \new_[51916]_ , \new_[51917]_ , \new_[51921]_ , \new_[51922]_ ,
    \new_[51925]_ , \new_[51928]_ , \new_[51929]_ , \new_[51930]_ ,
    \new_[51934]_ , \new_[51935]_ , \new_[51938]_ , \new_[51941]_ ,
    \new_[51942]_ , \new_[51943]_ , \new_[51947]_ , \new_[51948]_ ,
    \new_[51951]_ , \new_[51954]_ , \new_[51955]_ , \new_[51956]_ ,
    \new_[51960]_ , \new_[51961]_ , \new_[51964]_ , \new_[51967]_ ,
    \new_[51968]_ , \new_[51969]_ , \new_[51973]_ , \new_[51974]_ ,
    \new_[51977]_ , \new_[51980]_ , \new_[51981]_ , \new_[51982]_ ,
    \new_[51986]_ , \new_[51987]_ , \new_[51990]_ , \new_[51993]_ ,
    \new_[51994]_ , \new_[51995]_ , \new_[51999]_ , \new_[52000]_ ,
    \new_[52003]_ , \new_[52006]_ , \new_[52007]_ , \new_[52008]_ ,
    \new_[52012]_ , \new_[52013]_ , \new_[52016]_ , \new_[52019]_ ,
    \new_[52020]_ , \new_[52021]_ , \new_[52025]_ , \new_[52026]_ ,
    \new_[52029]_ , \new_[52032]_ , \new_[52033]_ , \new_[52034]_ ,
    \new_[52038]_ , \new_[52039]_ , \new_[52042]_ , \new_[52045]_ ,
    \new_[52046]_ , \new_[52047]_ , \new_[52051]_ , \new_[52052]_ ,
    \new_[52055]_ , \new_[52058]_ , \new_[52059]_ , \new_[52060]_ ,
    \new_[52064]_ , \new_[52065]_ , \new_[52068]_ , \new_[52071]_ ,
    \new_[52072]_ , \new_[52073]_ , \new_[52077]_ , \new_[52078]_ ,
    \new_[52081]_ , \new_[52084]_ , \new_[52085]_ , \new_[52086]_ ,
    \new_[52090]_ , \new_[52091]_ , \new_[52094]_ , \new_[52097]_ ,
    \new_[52098]_ , \new_[52099]_ , \new_[52103]_ , \new_[52104]_ ,
    \new_[52107]_ , \new_[52110]_ , \new_[52111]_ , \new_[52112]_ ,
    \new_[52116]_ , \new_[52117]_ , \new_[52120]_ , \new_[52123]_ ,
    \new_[52124]_ , \new_[52125]_ , \new_[52129]_ , \new_[52130]_ ,
    \new_[52133]_ , \new_[52136]_ , \new_[52137]_ , \new_[52138]_ ,
    \new_[52142]_ , \new_[52143]_ , \new_[52146]_ , \new_[52149]_ ,
    \new_[52150]_ , \new_[52151]_ , \new_[52155]_ , \new_[52156]_ ,
    \new_[52159]_ , \new_[52162]_ , \new_[52163]_ , \new_[52164]_ ,
    \new_[52168]_ , \new_[52169]_ , \new_[52172]_ , \new_[52175]_ ,
    \new_[52176]_ , \new_[52177]_ , \new_[52181]_ , \new_[52182]_ ,
    \new_[52185]_ , \new_[52188]_ , \new_[52189]_ , \new_[52190]_ ,
    \new_[52194]_ , \new_[52195]_ , \new_[52198]_ , \new_[52201]_ ,
    \new_[52202]_ , \new_[52203]_ , \new_[52207]_ , \new_[52208]_ ,
    \new_[52211]_ , \new_[52214]_ , \new_[52215]_ , \new_[52216]_ ,
    \new_[52220]_ , \new_[52221]_ , \new_[52224]_ , \new_[52227]_ ,
    \new_[52228]_ , \new_[52229]_ , \new_[52233]_ , \new_[52234]_ ,
    \new_[52237]_ , \new_[52240]_ , \new_[52241]_ , \new_[52242]_ ,
    \new_[52246]_ , \new_[52247]_ , \new_[52250]_ , \new_[52253]_ ,
    \new_[52254]_ , \new_[52255]_ , \new_[52259]_ , \new_[52260]_ ,
    \new_[52263]_ , \new_[52266]_ , \new_[52267]_ , \new_[52268]_ ,
    \new_[52272]_ , \new_[52273]_ , \new_[52276]_ , \new_[52279]_ ,
    \new_[52280]_ , \new_[52281]_ , \new_[52285]_ , \new_[52286]_ ,
    \new_[52289]_ , \new_[52292]_ , \new_[52293]_ , \new_[52294]_ ,
    \new_[52298]_ , \new_[52299]_ , \new_[52302]_ , \new_[52305]_ ,
    \new_[52306]_ , \new_[52307]_ , \new_[52311]_ , \new_[52312]_ ,
    \new_[52315]_ , \new_[52318]_ , \new_[52319]_ , \new_[52320]_ ,
    \new_[52324]_ , \new_[52325]_ , \new_[52328]_ , \new_[52331]_ ,
    \new_[52332]_ , \new_[52333]_ , \new_[52337]_ , \new_[52338]_ ,
    \new_[52341]_ , \new_[52344]_ , \new_[52345]_ , \new_[52346]_ ,
    \new_[52350]_ , \new_[52351]_ , \new_[52354]_ , \new_[52357]_ ,
    \new_[52358]_ , \new_[52359]_ , \new_[52363]_ , \new_[52364]_ ,
    \new_[52367]_ , \new_[52370]_ , \new_[52371]_ , \new_[52372]_ ,
    \new_[52376]_ , \new_[52377]_ , \new_[52380]_ , \new_[52383]_ ,
    \new_[52384]_ , \new_[52385]_ , \new_[52389]_ , \new_[52390]_ ,
    \new_[52393]_ , \new_[52396]_ , \new_[52397]_ , \new_[52398]_ ,
    \new_[52402]_ , \new_[52403]_ , \new_[52406]_ , \new_[52409]_ ,
    \new_[52410]_ , \new_[52411]_ , \new_[52415]_ , \new_[52416]_ ,
    \new_[52419]_ , \new_[52422]_ , \new_[52423]_ , \new_[52424]_ ,
    \new_[52428]_ , \new_[52429]_ , \new_[52432]_ , \new_[52435]_ ,
    \new_[52436]_ , \new_[52437]_ , \new_[52441]_ , \new_[52442]_ ,
    \new_[52445]_ , \new_[52448]_ , \new_[52449]_ , \new_[52450]_ ,
    \new_[52454]_ , \new_[52455]_ , \new_[52458]_ , \new_[52461]_ ,
    \new_[52462]_ , \new_[52463]_ , \new_[52467]_ , \new_[52468]_ ,
    \new_[52471]_ , \new_[52474]_ , \new_[52475]_ , \new_[52476]_ ,
    \new_[52480]_ , \new_[52481]_ , \new_[52484]_ , \new_[52487]_ ,
    \new_[52488]_ , \new_[52489]_ , \new_[52493]_ , \new_[52494]_ ,
    \new_[52497]_ , \new_[52500]_ , \new_[52501]_ , \new_[52502]_ ,
    \new_[52506]_ , \new_[52507]_ , \new_[52510]_ , \new_[52513]_ ,
    \new_[52514]_ , \new_[52515]_ , \new_[52519]_ , \new_[52520]_ ,
    \new_[52523]_ , \new_[52526]_ , \new_[52527]_ , \new_[52528]_ ,
    \new_[52532]_ , \new_[52533]_ , \new_[52536]_ , \new_[52539]_ ,
    \new_[52540]_ , \new_[52541]_ , \new_[52545]_ , \new_[52546]_ ,
    \new_[52549]_ , \new_[52552]_ , \new_[52553]_ , \new_[52554]_ ,
    \new_[52558]_ , \new_[52559]_ , \new_[52562]_ , \new_[52565]_ ,
    \new_[52566]_ , \new_[52567]_ , \new_[52571]_ , \new_[52572]_ ,
    \new_[52575]_ , \new_[52578]_ , \new_[52579]_ , \new_[52580]_ ,
    \new_[52584]_ , \new_[52585]_ , \new_[52588]_ , \new_[52591]_ ,
    \new_[52592]_ , \new_[52593]_ , \new_[52597]_ , \new_[52598]_ ,
    \new_[52601]_ , \new_[52604]_ , \new_[52605]_ , \new_[52606]_ ,
    \new_[52610]_ , \new_[52611]_ , \new_[52614]_ , \new_[52617]_ ,
    \new_[52618]_ , \new_[52619]_ , \new_[52623]_ , \new_[52624]_ ,
    \new_[52627]_ , \new_[52630]_ , \new_[52631]_ , \new_[52632]_ ,
    \new_[52636]_ , \new_[52637]_ , \new_[52640]_ , \new_[52643]_ ,
    \new_[52644]_ , \new_[52645]_ , \new_[52649]_ , \new_[52650]_ ,
    \new_[52653]_ , \new_[52656]_ , \new_[52657]_ , \new_[52658]_ ,
    \new_[52662]_ , \new_[52663]_ , \new_[52666]_ , \new_[52669]_ ,
    \new_[52670]_ , \new_[52671]_ , \new_[52675]_ , \new_[52676]_ ,
    \new_[52679]_ , \new_[52682]_ , \new_[52683]_ , \new_[52684]_ ,
    \new_[52688]_ , \new_[52689]_ , \new_[52692]_ , \new_[52695]_ ,
    \new_[52696]_ , \new_[52697]_ , \new_[52701]_ , \new_[52702]_ ,
    \new_[52705]_ , \new_[52708]_ , \new_[52709]_ , \new_[52710]_ ,
    \new_[52714]_ , \new_[52715]_ , \new_[52718]_ , \new_[52721]_ ,
    \new_[52722]_ , \new_[52723]_ , \new_[52727]_ , \new_[52728]_ ,
    \new_[52731]_ , \new_[52734]_ , \new_[52735]_ , \new_[52736]_ ,
    \new_[52740]_ , \new_[52741]_ , \new_[52744]_ , \new_[52747]_ ,
    \new_[52748]_ , \new_[52749]_ , \new_[52753]_ , \new_[52754]_ ,
    \new_[52757]_ , \new_[52760]_ , \new_[52761]_ , \new_[52762]_ ,
    \new_[52766]_ , \new_[52767]_ , \new_[52770]_ , \new_[52773]_ ,
    \new_[52774]_ , \new_[52775]_ , \new_[52779]_ , \new_[52780]_ ,
    \new_[52783]_ , \new_[52786]_ , \new_[52787]_ , \new_[52788]_ ,
    \new_[52792]_ , \new_[52793]_ , \new_[52796]_ , \new_[52799]_ ,
    \new_[52800]_ , \new_[52801]_ , \new_[52805]_ , \new_[52806]_ ,
    \new_[52809]_ , \new_[52812]_ , \new_[52813]_ , \new_[52814]_ ,
    \new_[52818]_ , \new_[52819]_ , \new_[52822]_ , \new_[52825]_ ,
    \new_[52826]_ , \new_[52827]_ , \new_[52831]_ , \new_[52832]_ ,
    \new_[52835]_ , \new_[52838]_ , \new_[52839]_ , \new_[52840]_ ,
    \new_[52844]_ , \new_[52845]_ , \new_[52848]_ , \new_[52851]_ ,
    \new_[52852]_ , \new_[52853]_ , \new_[52857]_ , \new_[52858]_ ,
    \new_[52861]_ , \new_[52864]_ , \new_[52865]_ , \new_[52866]_ ,
    \new_[52870]_ , \new_[52871]_ , \new_[52874]_ , \new_[52877]_ ,
    \new_[52878]_ , \new_[52879]_ , \new_[52883]_ , \new_[52884]_ ,
    \new_[52887]_ , \new_[52890]_ , \new_[52891]_ , \new_[52892]_ ,
    \new_[52896]_ , \new_[52897]_ , \new_[52900]_ , \new_[52903]_ ,
    \new_[52904]_ , \new_[52905]_ , \new_[52909]_ , \new_[52910]_ ,
    \new_[52913]_ , \new_[52916]_ , \new_[52917]_ , \new_[52918]_ ,
    \new_[52922]_ , \new_[52923]_ , \new_[52926]_ , \new_[52929]_ ,
    \new_[52930]_ , \new_[52931]_ , \new_[52935]_ , \new_[52936]_ ,
    \new_[52939]_ , \new_[52942]_ , \new_[52943]_ , \new_[52944]_ ,
    \new_[52948]_ , \new_[52949]_ , \new_[52952]_ , \new_[52955]_ ,
    \new_[52956]_ , \new_[52957]_ , \new_[52961]_ , \new_[52962]_ ,
    \new_[52965]_ , \new_[52968]_ , \new_[52969]_ , \new_[52970]_ ,
    \new_[52974]_ , \new_[52975]_ , \new_[52978]_ , \new_[52981]_ ,
    \new_[52982]_ , \new_[52983]_ , \new_[52987]_ , \new_[52988]_ ,
    \new_[52991]_ , \new_[52994]_ , \new_[52995]_ , \new_[52996]_ ,
    \new_[53000]_ , \new_[53001]_ , \new_[53004]_ , \new_[53007]_ ,
    \new_[53008]_ , \new_[53009]_ , \new_[53013]_ , \new_[53014]_ ,
    \new_[53017]_ , \new_[53020]_ , \new_[53021]_ , \new_[53022]_ ,
    \new_[53026]_ , \new_[53027]_ , \new_[53030]_ , \new_[53033]_ ,
    \new_[53034]_ , \new_[53035]_ , \new_[53039]_ , \new_[53040]_ ,
    \new_[53043]_ , \new_[53046]_ , \new_[53047]_ , \new_[53048]_ ,
    \new_[53052]_ , \new_[53053]_ , \new_[53056]_ , \new_[53059]_ ,
    \new_[53060]_ , \new_[53061]_ , \new_[53065]_ , \new_[53066]_ ,
    \new_[53069]_ , \new_[53072]_ , \new_[53073]_ , \new_[53074]_ ,
    \new_[53078]_ , \new_[53079]_ , \new_[53082]_ , \new_[53085]_ ,
    \new_[53086]_ , \new_[53087]_ , \new_[53091]_ , \new_[53092]_ ,
    \new_[53095]_ , \new_[53098]_ , \new_[53099]_ , \new_[53100]_ ,
    \new_[53104]_ , \new_[53105]_ , \new_[53108]_ , \new_[53111]_ ,
    \new_[53112]_ , \new_[53113]_ , \new_[53117]_ , \new_[53118]_ ,
    \new_[53121]_ , \new_[53124]_ , \new_[53125]_ , \new_[53126]_ ,
    \new_[53130]_ , \new_[53131]_ , \new_[53134]_ , \new_[53137]_ ,
    \new_[53138]_ , \new_[53139]_ , \new_[53143]_ , \new_[53144]_ ,
    \new_[53147]_ , \new_[53150]_ , \new_[53151]_ , \new_[53152]_ ,
    \new_[53156]_ , \new_[53157]_ , \new_[53160]_ , \new_[53163]_ ,
    \new_[53164]_ , \new_[53165]_ , \new_[53169]_ , \new_[53170]_ ,
    \new_[53173]_ , \new_[53176]_ , \new_[53177]_ , \new_[53178]_ ,
    \new_[53182]_ , \new_[53183]_ , \new_[53186]_ , \new_[53189]_ ,
    \new_[53190]_ , \new_[53191]_ , \new_[53195]_ , \new_[53196]_ ,
    \new_[53199]_ , \new_[53202]_ , \new_[53203]_ , \new_[53204]_ ,
    \new_[53208]_ , \new_[53209]_ , \new_[53212]_ , \new_[53215]_ ,
    \new_[53216]_ , \new_[53217]_ , \new_[53221]_ , \new_[53222]_ ,
    \new_[53225]_ , \new_[53228]_ , \new_[53229]_ , \new_[53230]_ ,
    \new_[53234]_ , \new_[53235]_ , \new_[53238]_ , \new_[53241]_ ,
    \new_[53242]_ , \new_[53243]_ , \new_[53247]_ , \new_[53248]_ ,
    \new_[53251]_ , \new_[53254]_ , \new_[53255]_ , \new_[53256]_ ,
    \new_[53260]_ , \new_[53261]_ , \new_[53264]_ , \new_[53267]_ ,
    \new_[53268]_ , \new_[53269]_ , \new_[53273]_ , \new_[53274]_ ,
    \new_[53277]_ , \new_[53280]_ , \new_[53281]_ , \new_[53282]_ ,
    \new_[53286]_ , \new_[53287]_ , \new_[53290]_ , \new_[53293]_ ,
    \new_[53294]_ , \new_[53295]_ , \new_[53299]_ , \new_[53300]_ ,
    \new_[53303]_ , \new_[53306]_ , \new_[53307]_ , \new_[53308]_ ,
    \new_[53312]_ , \new_[53313]_ , \new_[53316]_ , \new_[53319]_ ,
    \new_[53320]_ , \new_[53321]_ , \new_[53325]_ , \new_[53326]_ ,
    \new_[53329]_ , \new_[53332]_ , \new_[53333]_ , \new_[53334]_ ,
    \new_[53338]_ , \new_[53339]_ , \new_[53342]_ , \new_[53345]_ ,
    \new_[53346]_ , \new_[53347]_ , \new_[53351]_ , \new_[53352]_ ,
    \new_[53355]_ , \new_[53358]_ , \new_[53359]_ , \new_[53360]_ ,
    \new_[53364]_ , \new_[53365]_ , \new_[53368]_ , \new_[53371]_ ,
    \new_[53372]_ , \new_[53373]_ , \new_[53377]_ , \new_[53378]_ ,
    \new_[53381]_ , \new_[53384]_ , \new_[53385]_ , \new_[53386]_ ,
    \new_[53390]_ , \new_[53391]_ , \new_[53394]_ , \new_[53397]_ ,
    \new_[53398]_ , \new_[53399]_ , \new_[53403]_ , \new_[53404]_ ,
    \new_[53407]_ , \new_[53410]_ , \new_[53411]_ , \new_[53412]_ ,
    \new_[53416]_ , \new_[53417]_ , \new_[53420]_ , \new_[53423]_ ,
    \new_[53424]_ , \new_[53425]_ , \new_[53429]_ , \new_[53430]_ ,
    \new_[53433]_ , \new_[53436]_ , \new_[53437]_ , \new_[53438]_ ,
    \new_[53442]_ , \new_[53443]_ , \new_[53446]_ , \new_[53449]_ ,
    \new_[53450]_ , \new_[53451]_ , \new_[53455]_ , \new_[53456]_ ,
    \new_[53459]_ , \new_[53462]_ , \new_[53463]_ , \new_[53464]_ ,
    \new_[53468]_ , \new_[53469]_ , \new_[53472]_ , \new_[53475]_ ,
    \new_[53476]_ , \new_[53477]_ , \new_[53481]_ , \new_[53482]_ ,
    \new_[53485]_ , \new_[53488]_ , \new_[53489]_ , \new_[53490]_ ,
    \new_[53494]_ , \new_[53495]_ , \new_[53498]_ , \new_[53501]_ ,
    \new_[53502]_ , \new_[53503]_ , \new_[53507]_ , \new_[53508]_ ,
    \new_[53511]_ , \new_[53514]_ , \new_[53515]_ , \new_[53516]_ ,
    \new_[53520]_ , \new_[53521]_ , \new_[53524]_ , \new_[53527]_ ,
    \new_[53528]_ , \new_[53529]_ , \new_[53533]_ , \new_[53534]_ ,
    \new_[53537]_ , \new_[53540]_ , \new_[53541]_ , \new_[53542]_ ,
    \new_[53546]_ , \new_[53547]_ , \new_[53550]_ , \new_[53553]_ ,
    \new_[53554]_ , \new_[53555]_ , \new_[53559]_ , \new_[53560]_ ,
    \new_[53563]_ , \new_[53566]_ , \new_[53567]_ , \new_[53568]_ ,
    \new_[53572]_ , \new_[53573]_ , \new_[53576]_ , \new_[53579]_ ,
    \new_[53580]_ , \new_[53581]_ , \new_[53585]_ , \new_[53586]_ ,
    \new_[53589]_ , \new_[53592]_ , \new_[53593]_ , \new_[53594]_ ,
    \new_[53598]_ , \new_[53599]_ , \new_[53602]_ , \new_[53605]_ ,
    \new_[53606]_ , \new_[53607]_ , \new_[53611]_ , \new_[53612]_ ,
    \new_[53615]_ , \new_[53618]_ , \new_[53619]_ , \new_[53620]_ ,
    \new_[53624]_ , \new_[53625]_ , \new_[53628]_ , \new_[53631]_ ,
    \new_[53632]_ , \new_[53633]_ , \new_[53637]_ , \new_[53638]_ ,
    \new_[53641]_ , \new_[53644]_ , \new_[53645]_ , \new_[53646]_ ,
    \new_[53650]_ , \new_[53651]_ , \new_[53654]_ , \new_[53657]_ ,
    \new_[53658]_ , \new_[53659]_ , \new_[53663]_ , \new_[53664]_ ,
    \new_[53667]_ , \new_[53670]_ , \new_[53671]_ , \new_[53672]_ ,
    \new_[53676]_ , \new_[53677]_ , \new_[53680]_ , \new_[53683]_ ,
    \new_[53684]_ , \new_[53685]_ , \new_[53689]_ , \new_[53690]_ ,
    \new_[53693]_ , \new_[53696]_ , \new_[53697]_ , \new_[53698]_ ,
    \new_[53702]_ , \new_[53703]_ , \new_[53706]_ , \new_[53709]_ ,
    \new_[53710]_ , \new_[53711]_ , \new_[53715]_ , \new_[53716]_ ,
    \new_[53719]_ , \new_[53722]_ , \new_[53723]_ , \new_[53724]_ ,
    \new_[53728]_ , \new_[53729]_ , \new_[53732]_ , \new_[53735]_ ,
    \new_[53736]_ , \new_[53737]_ , \new_[53741]_ , \new_[53742]_ ,
    \new_[53745]_ , \new_[53748]_ , \new_[53749]_ , \new_[53750]_ ,
    \new_[53754]_ , \new_[53755]_ , \new_[53758]_ , \new_[53761]_ ,
    \new_[53762]_ , \new_[53763]_ , \new_[53767]_ , \new_[53768]_ ,
    \new_[53771]_ , \new_[53774]_ , \new_[53775]_ , \new_[53776]_ ,
    \new_[53780]_ , \new_[53781]_ , \new_[53784]_ , \new_[53787]_ ,
    \new_[53788]_ , \new_[53789]_ , \new_[53793]_ , \new_[53794]_ ,
    \new_[53797]_ , \new_[53800]_ , \new_[53801]_ , \new_[53802]_ ,
    \new_[53806]_ , \new_[53807]_ , \new_[53810]_ , \new_[53813]_ ,
    \new_[53814]_ , \new_[53815]_ , \new_[53819]_ , \new_[53820]_ ,
    \new_[53823]_ , \new_[53826]_ , \new_[53827]_ , \new_[53828]_ ,
    \new_[53832]_ , \new_[53833]_ , \new_[53836]_ , \new_[53839]_ ,
    \new_[53840]_ , \new_[53841]_ , \new_[53845]_ , \new_[53846]_ ,
    \new_[53849]_ , \new_[53852]_ , \new_[53853]_ , \new_[53854]_ ,
    \new_[53858]_ , \new_[53859]_ , \new_[53862]_ , \new_[53865]_ ,
    \new_[53866]_ , \new_[53867]_ , \new_[53871]_ , \new_[53872]_ ,
    \new_[53875]_ , \new_[53878]_ , \new_[53879]_ , \new_[53880]_ ,
    \new_[53884]_ , \new_[53885]_ , \new_[53888]_ , \new_[53891]_ ,
    \new_[53892]_ , \new_[53893]_ , \new_[53897]_ , \new_[53898]_ ,
    \new_[53901]_ , \new_[53904]_ , \new_[53905]_ , \new_[53906]_ ,
    \new_[53910]_ , \new_[53911]_ , \new_[53914]_ , \new_[53917]_ ,
    \new_[53918]_ , \new_[53919]_ , \new_[53923]_ , \new_[53924]_ ,
    \new_[53927]_ , \new_[53930]_ , \new_[53931]_ , \new_[53932]_ ,
    \new_[53936]_ , \new_[53937]_ , \new_[53940]_ , \new_[53943]_ ,
    \new_[53944]_ , \new_[53945]_ , \new_[53949]_ , \new_[53950]_ ,
    \new_[53953]_ , \new_[53956]_ , \new_[53957]_ , \new_[53958]_ ,
    \new_[53962]_ , \new_[53963]_ , \new_[53966]_ , \new_[53969]_ ,
    \new_[53970]_ , \new_[53971]_ , \new_[53975]_ , \new_[53976]_ ,
    \new_[53979]_ , \new_[53982]_ , \new_[53983]_ , \new_[53984]_ ,
    \new_[53988]_ , \new_[53989]_ , \new_[53992]_ , \new_[53995]_ ,
    \new_[53996]_ , \new_[53997]_ , \new_[54001]_ , \new_[54002]_ ,
    \new_[54005]_ , \new_[54008]_ , \new_[54009]_ , \new_[54010]_ ,
    \new_[54014]_ , \new_[54015]_ , \new_[54018]_ , \new_[54021]_ ,
    \new_[54022]_ , \new_[54023]_ , \new_[54027]_ , \new_[54028]_ ,
    \new_[54031]_ , \new_[54034]_ , \new_[54035]_ , \new_[54036]_ ,
    \new_[54040]_ , \new_[54041]_ , \new_[54044]_ , \new_[54047]_ ,
    \new_[54048]_ , \new_[54049]_ , \new_[54053]_ , \new_[54054]_ ,
    \new_[54057]_ , \new_[54060]_ , \new_[54061]_ , \new_[54062]_ ,
    \new_[54066]_ , \new_[54067]_ , \new_[54070]_ , \new_[54073]_ ,
    \new_[54074]_ , \new_[54075]_ , \new_[54079]_ , \new_[54080]_ ,
    \new_[54083]_ , \new_[54086]_ , \new_[54087]_ , \new_[54088]_ ,
    \new_[54092]_ , \new_[54093]_ , \new_[54096]_ , \new_[54099]_ ,
    \new_[54100]_ , \new_[54101]_ , \new_[54105]_ , \new_[54106]_ ,
    \new_[54109]_ , \new_[54112]_ , \new_[54113]_ , \new_[54114]_ ,
    \new_[54118]_ , \new_[54119]_ , \new_[54122]_ , \new_[54125]_ ,
    \new_[54126]_ , \new_[54127]_ , \new_[54131]_ , \new_[54132]_ ,
    \new_[54135]_ , \new_[54138]_ , \new_[54139]_ , \new_[54140]_ ,
    \new_[54144]_ , \new_[54145]_ , \new_[54148]_ , \new_[54151]_ ,
    \new_[54152]_ , \new_[54153]_ , \new_[54157]_ , \new_[54158]_ ,
    \new_[54161]_ , \new_[54164]_ , \new_[54165]_ , \new_[54166]_ ,
    \new_[54170]_ , \new_[54171]_ , \new_[54174]_ , \new_[54177]_ ,
    \new_[54178]_ , \new_[54179]_ , \new_[54183]_ , \new_[54184]_ ,
    \new_[54187]_ , \new_[54190]_ , \new_[54191]_ , \new_[54192]_ ,
    \new_[54196]_ , \new_[54197]_ , \new_[54200]_ , \new_[54203]_ ,
    \new_[54204]_ , \new_[54205]_ , \new_[54209]_ , \new_[54210]_ ,
    \new_[54213]_ , \new_[54216]_ , \new_[54217]_ , \new_[54218]_ ,
    \new_[54222]_ , \new_[54223]_ , \new_[54226]_ , \new_[54229]_ ,
    \new_[54230]_ , \new_[54231]_ , \new_[54235]_ , \new_[54236]_ ,
    \new_[54239]_ , \new_[54242]_ , \new_[54243]_ , \new_[54244]_ ,
    \new_[54248]_ , \new_[54249]_ , \new_[54252]_ , \new_[54255]_ ,
    \new_[54256]_ , \new_[54257]_ , \new_[54261]_ , \new_[54262]_ ,
    \new_[54265]_ , \new_[54268]_ , \new_[54269]_ , \new_[54270]_ ,
    \new_[54274]_ , \new_[54275]_ , \new_[54278]_ , \new_[54281]_ ,
    \new_[54282]_ , \new_[54283]_ , \new_[54287]_ , \new_[54288]_ ,
    \new_[54291]_ , \new_[54294]_ , \new_[54295]_ , \new_[54296]_ ,
    \new_[54300]_ , \new_[54301]_ , \new_[54304]_ , \new_[54307]_ ,
    \new_[54308]_ , \new_[54309]_ , \new_[54313]_ , \new_[54314]_ ,
    \new_[54317]_ , \new_[54320]_ , \new_[54321]_ , \new_[54322]_ ,
    \new_[54326]_ , \new_[54327]_ , \new_[54330]_ , \new_[54333]_ ,
    \new_[54334]_ , \new_[54335]_ , \new_[54339]_ , \new_[54340]_ ,
    \new_[54343]_ , \new_[54346]_ , \new_[54347]_ , \new_[54348]_ ,
    \new_[54352]_ , \new_[54353]_ , \new_[54356]_ , \new_[54359]_ ,
    \new_[54360]_ , \new_[54361]_ , \new_[54365]_ , \new_[54366]_ ,
    \new_[54369]_ , \new_[54372]_ , \new_[54373]_ , \new_[54374]_ ,
    \new_[54378]_ , \new_[54379]_ , \new_[54382]_ , \new_[54385]_ ,
    \new_[54386]_ , \new_[54387]_ , \new_[54391]_ , \new_[54392]_ ,
    \new_[54395]_ , \new_[54398]_ , \new_[54399]_ , \new_[54400]_ ,
    \new_[54404]_ , \new_[54405]_ , \new_[54408]_ , \new_[54411]_ ,
    \new_[54412]_ , \new_[54413]_ , \new_[54417]_ , \new_[54418]_ ,
    \new_[54421]_ , \new_[54424]_ , \new_[54425]_ , \new_[54426]_ ,
    \new_[54430]_ , \new_[54431]_ , \new_[54434]_ , \new_[54437]_ ,
    \new_[54438]_ , \new_[54439]_ , \new_[54443]_ , \new_[54444]_ ,
    \new_[54447]_ , \new_[54450]_ , \new_[54451]_ , \new_[54452]_ ,
    \new_[54456]_ , \new_[54457]_ , \new_[54460]_ , \new_[54463]_ ,
    \new_[54464]_ , \new_[54465]_ , \new_[54469]_ , \new_[54470]_ ,
    \new_[54473]_ , \new_[54476]_ , \new_[54477]_ , \new_[54478]_ ,
    \new_[54482]_ , \new_[54483]_ , \new_[54486]_ , \new_[54489]_ ,
    \new_[54490]_ , \new_[54491]_ , \new_[54495]_ , \new_[54496]_ ,
    \new_[54499]_ , \new_[54502]_ , \new_[54503]_ , \new_[54504]_ ,
    \new_[54508]_ , \new_[54509]_ , \new_[54512]_ , \new_[54515]_ ,
    \new_[54516]_ , \new_[54517]_ , \new_[54521]_ , \new_[54522]_ ,
    \new_[54525]_ , \new_[54528]_ , \new_[54529]_ , \new_[54530]_ ,
    \new_[54534]_ , \new_[54535]_ , \new_[54538]_ , \new_[54541]_ ,
    \new_[54542]_ , \new_[54543]_ , \new_[54547]_ , \new_[54548]_ ,
    \new_[54551]_ , \new_[54554]_ , \new_[54555]_ , \new_[54556]_ ,
    \new_[54560]_ , \new_[54561]_ , \new_[54564]_ , \new_[54567]_ ,
    \new_[54568]_ , \new_[54569]_ , \new_[54573]_ , \new_[54574]_ ,
    \new_[54577]_ , \new_[54580]_ , \new_[54581]_ , \new_[54582]_ ,
    \new_[54586]_ , \new_[54587]_ , \new_[54590]_ , \new_[54593]_ ,
    \new_[54594]_ , \new_[54595]_ , \new_[54599]_ , \new_[54600]_ ,
    \new_[54603]_ , \new_[54606]_ , \new_[54607]_ , \new_[54608]_ ,
    \new_[54612]_ , \new_[54613]_ , \new_[54616]_ , \new_[54619]_ ,
    \new_[54620]_ , \new_[54621]_ , \new_[54625]_ , \new_[54626]_ ,
    \new_[54629]_ , \new_[54632]_ , \new_[54633]_ , \new_[54634]_ ,
    \new_[54638]_ , \new_[54639]_ , \new_[54642]_ , \new_[54645]_ ,
    \new_[54646]_ , \new_[54647]_ , \new_[54651]_ , \new_[54652]_ ,
    \new_[54655]_ , \new_[54658]_ , \new_[54659]_ , \new_[54660]_ ,
    \new_[54664]_ , \new_[54665]_ , \new_[54668]_ , \new_[54671]_ ,
    \new_[54672]_ , \new_[54673]_ , \new_[54677]_ , \new_[54678]_ ,
    \new_[54681]_ , \new_[54684]_ , \new_[54685]_ , \new_[54686]_ ,
    \new_[54690]_ , \new_[54691]_ , \new_[54694]_ , \new_[54697]_ ,
    \new_[54698]_ , \new_[54699]_ , \new_[54703]_ , \new_[54704]_ ,
    \new_[54707]_ , \new_[54710]_ , \new_[54711]_ , \new_[54712]_ ,
    \new_[54716]_ , \new_[54717]_ , \new_[54720]_ , \new_[54723]_ ,
    \new_[54724]_ , \new_[54725]_ , \new_[54729]_ , \new_[54730]_ ,
    \new_[54733]_ , \new_[54736]_ , \new_[54737]_ , \new_[54738]_ ,
    \new_[54742]_ , \new_[54743]_ , \new_[54746]_ , \new_[54749]_ ,
    \new_[54750]_ , \new_[54751]_ , \new_[54755]_ , \new_[54756]_ ,
    \new_[54759]_ , \new_[54762]_ , \new_[54763]_ , \new_[54764]_ ,
    \new_[54768]_ , \new_[54769]_ , \new_[54772]_ , \new_[54775]_ ,
    \new_[54776]_ , \new_[54777]_ , \new_[54781]_ , \new_[54782]_ ,
    \new_[54785]_ , \new_[54788]_ , \new_[54789]_ , \new_[54790]_ ,
    \new_[54794]_ , \new_[54795]_ , \new_[54798]_ , \new_[54801]_ ,
    \new_[54802]_ , \new_[54803]_ , \new_[54807]_ , \new_[54808]_ ,
    \new_[54811]_ , \new_[54814]_ , \new_[54815]_ , \new_[54816]_ ,
    \new_[54820]_ , \new_[54821]_ , \new_[54824]_ , \new_[54827]_ ,
    \new_[54828]_ , \new_[54829]_ , \new_[54833]_ , \new_[54834]_ ,
    \new_[54837]_ , \new_[54840]_ , \new_[54841]_ , \new_[54842]_ ,
    \new_[54846]_ , \new_[54847]_ , \new_[54850]_ , \new_[54853]_ ,
    \new_[54854]_ , \new_[54855]_ , \new_[54859]_ , \new_[54860]_ ,
    \new_[54863]_ , \new_[54866]_ , \new_[54867]_ , \new_[54868]_ ,
    \new_[54872]_ , \new_[54873]_ , \new_[54876]_ , \new_[54879]_ ,
    \new_[54880]_ , \new_[54881]_ , \new_[54885]_ , \new_[54886]_ ,
    \new_[54889]_ , \new_[54892]_ , \new_[54893]_ , \new_[54894]_ ,
    \new_[54898]_ , \new_[54899]_ , \new_[54902]_ , \new_[54905]_ ,
    \new_[54906]_ , \new_[54907]_ , \new_[54911]_ , \new_[54912]_ ,
    \new_[54915]_ , \new_[54918]_ , \new_[54919]_ , \new_[54920]_ ,
    \new_[54924]_ , \new_[54925]_ , \new_[54928]_ , \new_[54931]_ ,
    \new_[54932]_ , \new_[54933]_ , \new_[54937]_ , \new_[54938]_ ,
    \new_[54941]_ , \new_[54944]_ , \new_[54945]_ , \new_[54946]_ ,
    \new_[54950]_ , \new_[54951]_ , \new_[54954]_ , \new_[54957]_ ,
    \new_[54958]_ , \new_[54959]_ , \new_[54963]_ , \new_[54964]_ ,
    \new_[54967]_ , \new_[54970]_ , \new_[54971]_ , \new_[54972]_ ,
    \new_[54976]_ , \new_[54977]_ , \new_[54980]_ , \new_[54983]_ ,
    \new_[54984]_ , \new_[54985]_ , \new_[54989]_ , \new_[54990]_ ,
    \new_[54993]_ , \new_[54996]_ , \new_[54997]_ , \new_[54998]_ ,
    \new_[55002]_ , \new_[55003]_ , \new_[55006]_ , \new_[55009]_ ,
    \new_[55010]_ , \new_[55011]_ , \new_[55015]_ , \new_[55016]_ ,
    \new_[55019]_ , \new_[55022]_ , \new_[55023]_ , \new_[55024]_ ,
    \new_[55028]_ , \new_[55029]_ , \new_[55032]_ , \new_[55035]_ ,
    \new_[55036]_ , \new_[55037]_ , \new_[55041]_ , \new_[55042]_ ,
    \new_[55045]_ , \new_[55048]_ , \new_[55049]_ , \new_[55050]_ ,
    \new_[55054]_ , \new_[55055]_ , \new_[55058]_ , \new_[55061]_ ,
    \new_[55062]_ , \new_[55063]_ , \new_[55067]_ , \new_[55068]_ ,
    \new_[55071]_ , \new_[55074]_ , \new_[55075]_ , \new_[55076]_ ,
    \new_[55080]_ , \new_[55081]_ , \new_[55084]_ , \new_[55087]_ ,
    \new_[55088]_ , \new_[55089]_ , \new_[55093]_ , \new_[55094]_ ,
    \new_[55097]_ , \new_[55100]_ , \new_[55101]_ , \new_[55102]_ ,
    \new_[55106]_ , \new_[55107]_ , \new_[55110]_ , \new_[55113]_ ,
    \new_[55114]_ , \new_[55115]_ , \new_[55119]_ , \new_[55120]_ ,
    \new_[55123]_ , \new_[55126]_ , \new_[55127]_ , \new_[55128]_ ,
    \new_[55132]_ , \new_[55133]_ , \new_[55136]_ , \new_[55139]_ ,
    \new_[55140]_ , \new_[55141]_ , \new_[55145]_ , \new_[55146]_ ,
    \new_[55149]_ , \new_[55152]_ , \new_[55153]_ , \new_[55154]_ ,
    \new_[55158]_ , \new_[55159]_ , \new_[55162]_ , \new_[55165]_ ,
    \new_[55166]_ , \new_[55167]_ , \new_[55171]_ , \new_[55172]_ ,
    \new_[55175]_ , \new_[55178]_ , \new_[55179]_ , \new_[55180]_ ,
    \new_[55184]_ , \new_[55185]_ , \new_[55188]_ , \new_[55191]_ ,
    \new_[55192]_ , \new_[55193]_ , \new_[55197]_ , \new_[55198]_ ,
    \new_[55201]_ , \new_[55204]_ , \new_[55205]_ , \new_[55206]_ ,
    \new_[55210]_ , \new_[55211]_ , \new_[55214]_ , \new_[55217]_ ,
    \new_[55218]_ , \new_[55219]_ , \new_[55223]_ , \new_[55224]_ ,
    \new_[55227]_ , \new_[55230]_ , \new_[55231]_ , \new_[55232]_ ,
    \new_[55236]_ , \new_[55237]_ , \new_[55240]_ , \new_[55243]_ ,
    \new_[55244]_ , \new_[55245]_ , \new_[55249]_ , \new_[55250]_ ,
    \new_[55253]_ , \new_[55256]_ , \new_[55257]_ , \new_[55258]_ ,
    \new_[55262]_ , \new_[55263]_ , \new_[55266]_ , \new_[55269]_ ,
    \new_[55270]_ , \new_[55271]_ , \new_[55275]_ , \new_[55276]_ ,
    \new_[55279]_ , \new_[55282]_ , \new_[55283]_ , \new_[55284]_ ,
    \new_[55288]_ , \new_[55289]_ , \new_[55292]_ , \new_[55295]_ ,
    \new_[55296]_ , \new_[55297]_ , \new_[55301]_ , \new_[55302]_ ,
    \new_[55305]_ , \new_[55308]_ , \new_[55309]_ , \new_[55310]_ ,
    \new_[55314]_ , \new_[55315]_ , \new_[55318]_ , \new_[55321]_ ,
    \new_[55322]_ , \new_[55323]_ , \new_[55327]_ , \new_[55328]_ ,
    \new_[55331]_ , \new_[55334]_ , \new_[55335]_ , \new_[55336]_ ,
    \new_[55340]_ , \new_[55341]_ , \new_[55344]_ , \new_[55347]_ ,
    \new_[55348]_ , \new_[55349]_ , \new_[55353]_ , \new_[55354]_ ,
    \new_[55357]_ , \new_[55360]_ , \new_[55361]_ , \new_[55362]_ ,
    \new_[55366]_ , \new_[55367]_ , \new_[55370]_ , \new_[55373]_ ,
    \new_[55374]_ , \new_[55375]_ , \new_[55379]_ , \new_[55380]_ ,
    \new_[55383]_ , \new_[55386]_ , \new_[55387]_ , \new_[55388]_ ,
    \new_[55392]_ , \new_[55393]_ , \new_[55396]_ , \new_[55399]_ ,
    \new_[55400]_ , \new_[55401]_ , \new_[55405]_ , \new_[55406]_ ,
    \new_[55409]_ , \new_[55412]_ , \new_[55413]_ , \new_[55414]_ ,
    \new_[55418]_ , \new_[55419]_ , \new_[55422]_ , \new_[55425]_ ,
    \new_[55426]_ , \new_[55427]_ , \new_[55431]_ , \new_[55432]_ ,
    \new_[55435]_ , \new_[55438]_ , \new_[55439]_ , \new_[55440]_ ,
    \new_[55444]_ , \new_[55445]_ , \new_[55448]_ , \new_[55451]_ ,
    \new_[55452]_ , \new_[55453]_ , \new_[55457]_ , \new_[55458]_ ,
    \new_[55461]_ , \new_[55464]_ , \new_[55465]_ , \new_[55466]_ ,
    \new_[55470]_ , \new_[55471]_ , \new_[55474]_ , \new_[55477]_ ,
    \new_[55478]_ , \new_[55479]_ , \new_[55483]_ , \new_[55484]_ ,
    \new_[55487]_ , \new_[55490]_ , \new_[55491]_ , \new_[55492]_ ,
    \new_[55496]_ , \new_[55497]_ , \new_[55500]_ , \new_[55503]_ ,
    \new_[55504]_ , \new_[55505]_ , \new_[55509]_ , \new_[55510]_ ,
    \new_[55513]_ , \new_[55516]_ , \new_[55517]_ , \new_[55518]_ ,
    \new_[55522]_ , \new_[55523]_ , \new_[55526]_ , \new_[55529]_ ,
    \new_[55530]_ , \new_[55531]_ , \new_[55535]_ , \new_[55536]_ ,
    \new_[55539]_ , \new_[55542]_ , \new_[55543]_ , \new_[55544]_ ,
    \new_[55548]_ , \new_[55549]_ , \new_[55552]_ , \new_[55555]_ ,
    \new_[55556]_ , \new_[55557]_ , \new_[55561]_ , \new_[55562]_ ,
    \new_[55565]_ , \new_[55568]_ , \new_[55569]_ , \new_[55570]_ ,
    \new_[55574]_ , \new_[55575]_ , \new_[55578]_ , \new_[55581]_ ,
    \new_[55582]_ , \new_[55583]_ , \new_[55587]_ , \new_[55588]_ ,
    \new_[55591]_ , \new_[55594]_ , \new_[55595]_ , \new_[55596]_ ,
    \new_[55600]_ , \new_[55601]_ , \new_[55604]_ , \new_[55607]_ ,
    \new_[55608]_ , \new_[55609]_ , \new_[55613]_ , \new_[55614]_ ,
    \new_[55617]_ , \new_[55620]_ , \new_[55621]_ , \new_[55622]_ ,
    \new_[55626]_ , \new_[55627]_ , \new_[55630]_ , \new_[55633]_ ,
    \new_[55634]_ , \new_[55635]_ , \new_[55639]_ , \new_[55640]_ ,
    \new_[55643]_ , \new_[55646]_ , \new_[55647]_ , \new_[55648]_ ,
    \new_[55652]_ , \new_[55653]_ , \new_[55656]_ , \new_[55659]_ ,
    \new_[55660]_ , \new_[55661]_ , \new_[55665]_ , \new_[55666]_ ,
    \new_[55669]_ , \new_[55672]_ , \new_[55673]_ , \new_[55674]_ ,
    \new_[55678]_ , \new_[55679]_ , \new_[55682]_ , \new_[55685]_ ,
    \new_[55686]_ , \new_[55687]_ , \new_[55691]_ , \new_[55692]_ ,
    \new_[55695]_ , \new_[55698]_ , \new_[55699]_ , \new_[55700]_ ,
    \new_[55704]_ , \new_[55705]_ , \new_[55708]_ , \new_[55711]_ ,
    \new_[55712]_ , \new_[55713]_ , \new_[55717]_ , \new_[55718]_ ,
    \new_[55721]_ , \new_[55724]_ , \new_[55725]_ , \new_[55726]_ ,
    \new_[55730]_ , \new_[55731]_ , \new_[55734]_ , \new_[55737]_ ,
    \new_[55738]_ , \new_[55739]_ , \new_[55743]_ , \new_[55744]_ ,
    \new_[55747]_ , \new_[55750]_ , \new_[55751]_ , \new_[55752]_ ,
    \new_[55756]_ , \new_[55757]_ , \new_[55760]_ , \new_[55763]_ ,
    \new_[55764]_ , \new_[55765]_ , \new_[55769]_ , \new_[55770]_ ,
    \new_[55773]_ , \new_[55776]_ , \new_[55777]_ , \new_[55778]_ ,
    \new_[55782]_ , \new_[55783]_ , \new_[55786]_ , \new_[55789]_ ,
    \new_[55790]_ , \new_[55791]_ , \new_[55795]_ , \new_[55796]_ ,
    \new_[55799]_ , \new_[55802]_ , \new_[55803]_ , \new_[55804]_ ,
    \new_[55808]_ , \new_[55809]_ , \new_[55812]_ , \new_[55815]_ ,
    \new_[55816]_ , \new_[55817]_ , \new_[55821]_ , \new_[55822]_ ,
    \new_[55825]_ , \new_[55828]_ , \new_[55829]_ , \new_[55830]_ ,
    \new_[55834]_ , \new_[55835]_ , \new_[55838]_ , \new_[55841]_ ,
    \new_[55842]_ , \new_[55843]_ , \new_[55847]_ , \new_[55848]_ ,
    \new_[55851]_ , \new_[55854]_ , \new_[55855]_ , \new_[55856]_ ,
    \new_[55860]_ , \new_[55861]_ , \new_[55864]_ , \new_[55867]_ ,
    \new_[55868]_ , \new_[55869]_ , \new_[55873]_ , \new_[55874]_ ,
    \new_[55877]_ , \new_[55880]_ , \new_[55881]_ , \new_[55882]_ ,
    \new_[55886]_ , \new_[55887]_ , \new_[55890]_ , \new_[55893]_ ,
    \new_[55894]_ , \new_[55895]_ , \new_[55899]_ , \new_[55900]_ ,
    \new_[55903]_ , \new_[55906]_ , \new_[55907]_ , \new_[55908]_ ,
    \new_[55912]_ , \new_[55913]_ , \new_[55916]_ , \new_[55919]_ ,
    \new_[55920]_ , \new_[55921]_ , \new_[55925]_ , \new_[55926]_ ,
    \new_[55929]_ , \new_[55932]_ , \new_[55933]_ , \new_[55934]_ ,
    \new_[55938]_ , \new_[55939]_ , \new_[55942]_ , \new_[55945]_ ,
    \new_[55946]_ , \new_[55947]_ , \new_[55951]_ , \new_[55952]_ ,
    \new_[55955]_ , \new_[55958]_ , \new_[55959]_ , \new_[55960]_ ,
    \new_[55964]_ , \new_[55965]_ , \new_[55968]_ , \new_[55971]_ ,
    \new_[55972]_ , \new_[55973]_ , \new_[55977]_ , \new_[55978]_ ,
    \new_[55981]_ , \new_[55984]_ , \new_[55985]_ , \new_[55986]_ ,
    \new_[55990]_ , \new_[55991]_ , \new_[55994]_ , \new_[55997]_ ,
    \new_[55998]_ , \new_[55999]_ , \new_[56003]_ , \new_[56004]_ ,
    \new_[56007]_ , \new_[56010]_ , \new_[56011]_ , \new_[56012]_ ,
    \new_[56016]_ , \new_[56017]_ , \new_[56020]_ , \new_[56023]_ ,
    \new_[56024]_ , \new_[56025]_ , \new_[56029]_ , \new_[56030]_ ,
    \new_[56033]_ , \new_[56036]_ , \new_[56037]_ , \new_[56038]_ ,
    \new_[56042]_ , \new_[56043]_ , \new_[56046]_ , \new_[56049]_ ,
    \new_[56050]_ , \new_[56051]_ , \new_[56055]_ , \new_[56056]_ ,
    \new_[56059]_ , \new_[56062]_ , \new_[56063]_ , \new_[56064]_ ,
    \new_[56068]_ , \new_[56069]_ , \new_[56072]_ , \new_[56075]_ ,
    \new_[56076]_ , \new_[56077]_ , \new_[56081]_ , \new_[56082]_ ,
    \new_[56085]_ , \new_[56088]_ , \new_[56089]_ , \new_[56090]_ ,
    \new_[56094]_ , \new_[56095]_ , \new_[56098]_ , \new_[56101]_ ,
    \new_[56102]_ , \new_[56103]_ , \new_[56107]_ , \new_[56108]_ ,
    \new_[56111]_ , \new_[56114]_ , \new_[56115]_ , \new_[56116]_ ,
    \new_[56120]_ , \new_[56121]_ , \new_[56124]_ , \new_[56127]_ ,
    \new_[56128]_ , \new_[56129]_ , \new_[56133]_ , \new_[56134]_ ,
    \new_[56137]_ , \new_[56140]_ , \new_[56141]_ , \new_[56142]_ ,
    \new_[56146]_ , \new_[56147]_ , \new_[56150]_ , \new_[56153]_ ,
    \new_[56154]_ , \new_[56155]_ , \new_[56159]_ , \new_[56160]_ ,
    \new_[56163]_ , \new_[56166]_ , \new_[56167]_ , \new_[56168]_ ,
    \new_[56172]_ , \new_[56173]_ , \new_[56176]_ , \new_[56179]_ ,
    \new_[56180]_ , \new_[56181]_ , \new_[56185]_ , \new_[56186]_ ,
    \new_[56189]_ , \new_[56192]_ , \new_[56193]_ , \new_[56194]_ ,
    \new_[56198]_ , \new_[56199]_ , \new_[56202]_ , \new_[56205]_ ,
    \new_[56206]_ , \new_[56207]_ , \new_[56211]_ , \new_[56212]_ ,
    \new_[56215]_ , \new_[56218]_ , \new_[56219]_ , \new_[56220]_ ,
    \new_[56224]_ , \new_[56225]_ , \new_[56228]_ , \new_[56231]_ ,
    \new_[56232]_ , \new_[56233]_ , \new_[56237]_ , \new_[56238]_ ,
    \new_[56241]_ , \new_[56244]_ , \new_[56245]_ , \new_[56246]_ ,
    \new_[56250]_ , \new_[56251]_ , \new_[56254]_ , \new_[56257]_ ,
    \new_[56258]_ , \new_[56259]_ , \new_[56263]_ , \new_[56264]_ ,
    \new_[56267]_ , \new_[56270]_ , \new_[56271]_ , \new_[56272]_ ,
    \new_[56276]_ , \new_[56277]_ , \new_[56280]_ , \new_[56283]_ ,
    \new_[56284]_ , \new_[56285]_ , \new_[56289]_ , \new_[56290]_ ,
    \new_[56293]_ , \new_[56296]_ , \new_[56297]_ , \new_[56298]_ ,
    \new_[56302]_ , \new_[56303]_ , \new_[56306]_ , \new_[56309]_ ,
    \new_[56310]_ , \new_[56311]_ , \new_[56315]_ , \new_[56316]_ ,
    \new_[56319]_ , \new_[56322]_ , \new_[56323]_ , \new_[56324]_ ,
    \new_[56328]_ , \new_[56329]_ , \new_[56332]_ , \new_[56335]_ ,
    \new_[56336]_ , \new_[56337]_ , \new_[56341]_ , \new_[56342]_ ,
    \new_[56345]_ , \new_[56348]_ , \new_[56349]_ , \new_[56350]_ ,
    \new_[56354]_ , \new_[56355]_ , \new_[56358]_ , \new_[56361]_ ,
    \new_[56362]_ , \new_[56363]_ , \new_[56367]_ , \new_[56368]_ ,
    \new_[56371]_ , \new_[56374]_ , \new_[56375]_ , \new_[56376]_ ,
    \new_[56380]_ , \new_[56381]_ , \new_[56384]_ , \new_[56387]_ ,
    \new_[56388]_ , \new_[56389]_ , \new_[56393]_ , \new_[56394]_ ,
    \new_[56397]_ , \new_[56400]_ , \new_[56401]_ , \new_[56402]_ ,
    \new_[56406]_ , \new_[56407]_ , \new_[56410]_ , \new_[56413]_ ,
    \new_[56414]_ , \new_[56415]_ , \new_[56419]_ , \new_[56420]_ ,
    \new_[56423]_ , \new_[56426]_ , \new_[56427]_ , \new_[56428]_ ,
    \new_[56432]_ , \new_[56433]_ , \new_[56436]_ , \new_[56439]_ ,
    \new_[56440]_ , \new_[56441]_ , \new_[56445]_ , \new_[56446]_ ,
    \new_[56449]_ , \new_[56452]_ , \new_[56453]_ , \new_[56454]_ ,
    \new_[56458]_ , \new_[56459]_ , \new_[56462]_ , \new_[56465]_ ,
    \new_[56466]_ , \new_[56467]_ , \new_[56471]_ , \new_[56472]_ ,
    \new_[56475]_ , \new_[56478]_ , \new_[56479]_ , \new_[56480]_ ,
    \new_[56484]_ , \new_[56485]_ , \new_[56488]_ , \new_[56491]_ ,
    \new_[56492]_ , \new_[56493]_ , \new_[56497]_ , \new_[56498]_ ,
    \new_[56501]_ , \new_[56504]_ , \new_[56505]_ , \new_[56506]_ ,
    \new_[56510]_ , \new_[56511]_ , \new_[56514]_ , \new_[56517]_ ,
    \new_[56518]_ , \new_[56519]_ , \new_[56523]_ , \new_[56524]_ ,
    \new_[56527]_ , \new_[56530]_ , \new_[56531]_ , \new_[56532]_ ,
    \new_[56536]_ , \new_[56537]_ , \new_[56540]_ , \new_[56543]_ ,
    \new_[56544]_ , \new_[56545]_ , \new_[56549]_ , \new_[56550]_ ,
    \new_[56553]_ , \new_[56556]_ , \new_[56557]_ , \new_[56558]_ ,
    \new_[56562]_ , \new_[56563]_ , \new_[56566]_ , \new_[56569]_ ,
    \new_[56570]_ , \new_[56571]_ , \new_[56575]_ , \new_[56576]_ ,
    \new_[56579]_ , \new_[56582]_ , \new_[56583]_ , \new_[56584]_ ,
    \new_[56588]_ , \new_[56589]_ , \new_[56592]_ , \new_[56595]_ ,
    \new_[56596]_ , \new_[56597]_ , \new_[56601]_ , \new_[56602]_ ,
    \new_[56605]_ , \new_[56608]_ , \new_[56609]_ , \new_[56610]_ ,
    \new_[56614]_ , \new_[56615]_ , \new_[56618]_ , \new_[56621]_ ,
    \new_[56622]_ , \new_[56623]_ , \new_[56627]_ , \new_[56628]_ ,
    \new_[56631]_ , \new_[56634]_ , \new_[56635]_ , \new_[56636]_ ,
    \new_[56640]_ , \new_[56641]_ , \new_[56644]_ , \new_[56647]_ ,
    \new_[56648]_ , \new_[56649]_ , \new_[56653]_ , \new_[56654]_ ,
    \new_[56657]_ , \new_[56660]_ , \new_[56661]_ , \new_[56662]_ ,
    \new_[56666]_ , \new_[56667]_ , \new_[56670]_ , \new_[56673]_ ,
    \new_[56674]_ , \new_[56675]_ , \new_[56679]_ , \new_[56680]_ ,
    \new_[56683]_ , \new_[56686]_ , \new_[56687]_ , \new_[56688]_ ,
    \new_[56692]_ , \new_[56693]_ , \new_[56696]_ , \new_[56699]_ ,
    \new_[56700]_ , \new_[56701]_ , \new_[56705]_ , \new_[56706]_ ,
    \new_[56709]_ , \new_[56712]_ , \new_[56713]_ , \new_[56714]_ ,
    \new_[56718]_ , \new_[56719]_ , \new_[56722]_ , \new_[56725]_ ,
    \new_[56726]_ , \new_[56727]_ , \new_[56731]_ , \new_[56732]_ ,
    \new_[56735]_ , \new_[56738]_ , \new_[56739]_ , \new_[56740]_ ,
    \new_[56744]_ , \new_[56745]_ , \new_[56748]_ , \new_[56751]_ ,
    \new_[56752]_ , \new_[56753]_ , \new_[56757]_ , \new_[56758]_ ,
    \new_[56761]_ , \new_[56764]_ , \new_[56765]_ , \new_[56766]_ ,
    \new_[56770]_ , \new_[56771]_ , \new_[56774]_ , \new_[56777]_ ,
    \new_[56778]_ , \new_[56779]_ , \new_[56783]_ , \new_[56784]_ ,
    \new_[56787]_ , \new_[56790]_ , \new_[56791]_ , \new_[56792]_ ,
    \new_[56796]_ , \new_[56797]_ , \new_[56800]_ , \new_[56803]_ ,
    \new_[56804]_ , \new_[56805]_ , \new_[56809]_ , \new_[56810]_ ,
    \new_[56813]_ , \new_[56816]_ , \new_[56817]_ , \new_[56818]_ ,
    \new_[56822]_ , \new_[56823]_ , \new_[56826]_ , \new_[56829]_ ,
    \new_[56830]_ , \new_[56831]_ , \new_[56835]_ , \new_[56836]_ ,
    \new_[56839]_ , \new_[56842]_ , \new_[56843]_ , \new_[56844]_ ,
    \new_[56848]_ , \new_[56849]_ , \new_[56852]_ , \new_[56855]_ ,
    \new_[56856]_ , \new_[56857]_ , \new_[56861]_ , \new_[56862]_ ,
    \new_[56865]_ , \new_[56868]_ , \new_[56869]_ , \new_[56870]_ ,
    \new_[56874]_ , \new_[56875]_ , \new_[56878]_ , \new_[56881]_ ,
    \new_[56882]_ , \new_[56883]_ , \new_[56887]_ , \new_[56888]_ ,
    \new_[56891]_ , \new_[56894]_ , \new_[56895]_ , \new_[56896]_ ,
    \new_[56900]_ , \new_[56901]_ , \new_[56904]_ , \new_[56907]_ ,
    \new_[56908]_ , \new_[56909]_ , \new_[56913]_ , \new_[56914]_ ,
    \new_[56917]_ , \new_[56920]_ , \new_[56921]_ , \new_[56922]_ ,
    \new_[56926]_ , \new_[56927]_ , \new_[56930]_ , \new_[56933]_ ,
    \new_[56934]_ , \new_[56935]_ , \new_[56939]_ , \new_[56940]_ ,
    \new_[56943]_ , \new_[56946]_ , \new_[56947]_ , \new_[56948]_ ,
    \new_[56952]_ , \new_[56953]_ , \new_[56956]_ , \new_[56959]_ ,
    \new_[56960]_ , \new_[56961]_ , \new_[56965]_ , \new_[56966]_ ,
    \new_[56969]_ , \new_[56972]_ , \new_[56973]_ , \new_[56974]_ ,
    \new_[56978]_ , \new_[56979]_ , \new_[56982]_ , \new_[56985]_ ,
    \new_[56986]_ , \new_[56987]_ , \new_[56991]_ , \new_[56992]_ ,
    \new_[56995]_ , \new_[56998]_ , \new_[56999]_ , \new_[57000]_ ,
    \new_[57004]_ , \new_[57005]_ , \new_[57008]_ , \new_[57011]_ ,
    \new_[57012]_ , \new_[57013]_ , \new_[57017]_ , \new_[57018]_ ,
    \new_[57021]_ , \new_[57024]_ , \new_[57025]_ , \new_[57026]_ ,
    \new_[57030]_ , \new_[57031]_ , \new_[57034]_ , \new_[57037]_ ,
    \new_[57038]_ , \new_[57039]_ , \new_[57043]_ , \new_[57044]_ ,
    \new_[57047]_ , \new_[57050]_ , \new_[57051]_ , \new_[57052]_ ,
    \new_[57056]_ , \new_[57057]_ , \new_[57060]_ , \new_[57063]_ ,
    \new_[57064]_ , \new_[57065]_ , \new_[57069]_ , \new_[57070]_ ,
    \new_[57073]_ , \new_[57076]_ , \new_[57077]_ , \new_[57078]_ ,
    \new_[57082]_ , \new_[57083]_ , \new_[57086]_ , \new_[57089]_ ,
    \new_[57090]_ , \new_[57091]_ , \new_[57095]_ , \new_[57096]_ ,
    \new_[57099]_ , \new_[57102]_ , \new_[57103]_ , \new_[57104]_ ,
    \new_[57108]_ , \new_[57109]_ , \new_[57112]_ , \new_[57115]_ ,
    \new_[57116]_ , \new_[57117]_ , \new_[57121]_ , \new_[57122]_ ,
    \new_[57125]_ , \new_[57128]_ , \new_[57129]_ , \new_[57130]_ ,
    \new_[57134]_ , \new_[57135]_ , \new_[57138]_ , \new_[57141]_ ,
    \new_[57142]_ , \new_[57143]_ , \new_[57147]_ , \new_[57148]_ ,
    \new_[57151]_ , \new_[57154]_ , \new_[57155]_ , \new_[57156]_ ,
    \new_[57160]_ , \new_[57161]_ , \new_[57164]_ , \new_[57167]_ ,
    \new_[57168]_ , \new_[57169]_ , \new_[57173]_ , \new_[57174]_ ,
    \new_[57177]_ , \new_[57180]_ , \new_[57181]_ , \new_[57182]_ ,
    \new_[57186]_ , \new_[57187]_ , \new_[57190]_ , \new_[57193]_ ,
    \new_[57194]_ , \new_[57195]_ , \new_[57199]_ , \new_[57200]_ ,
    \new_[57203]_ , \new_[57206]_ , \new_[57207]_ , \new_[57208]_ ,
    \new_[57212]_ , \new_[57213]_ , \new_[57216]_ , \new_[57219]_ ,
    \new_[57220]_ , \new_[57221]_ , \new_[57225]_ , \new_[57226]_ ,
    \new_[57229]_ , \new_[57232]_ , \new_[57233]_ , \new_[57234]_ ,
    \new_[57238]_ , \new_[57239]_ , \new_[57242]_ , \new_[57245]_ ,
    \new_[57246]_ , \new_[57247]_ , \new_[57251]_ , \new_[57252]_ ,
    \new_[57255]_ , \new_[57258]_ , \new_[57259]_ , \new_[57260]_ ,
    \new_[57264]_ , \new_[57265]_ , \new_[57268]_ , \new_[57271]_ ,
    \new_[57272]_ , \new_[57273]_ , \new_[57277]_ , \new_[57278]_ ,
    \new_[57281]_ , \new_[57284]_ , \new_[57285]_ , \new_[57286]_ ,
    \new_[57290]_ , \new_[57291]_ , \new_[57294]_ , \new_[57297]_ ,
    \new_[57298]_ , \new_[57299]_ , \new_[57303]_ , \new_[57304]_ ,
    \new_[57307]_ , \new_[57310]_ , \new_[57311]_ , \new_[57312]_ ,
    \new_[57316]_ , \new_[57317]_ , \new_[57320]_ , \new_[57323]_ ,
    \new_[57324]_ , \new_[57325]_ , \new_[57329]_ , \new_[57330]_ ,
    \new_[57333]_ , \new_[57336]_ , \new_[57337]_ , \new_[57338]_ ,
    \new_[57342]_ , \new_[57343]_ , \new_[57346]_ , \new_[57349]_ ,
    \new_[57350]_ , \new_[57351]_ , \new_[57355]_ , \new_[57356]_ ,
    \new_[57359]_ , \new_[57362]_ , \new_[57363]_ , \new_[57364]_ ,
    \new_[57368]_ , \new_[57369]_ , \new_[57372]_ , \new_[57375]_ ,
    \new_[57376]_ , \new_[57377]_ , \new_[57381]_ , \new_[57382]_ ,
    \new_[57385]_ , \new_[57388]_ , \new_[57389]_ , \new_[57390]_ ,
    \new_[57394]_ , \new_[57395]_ , \new_[57398]_ , \new_[57401]_ ,
    \new_[57402]_ , \new_[57403]_ , \new_[57407]_ , \new_[57408]_ ,
    \new_[57411]_ , \new_[57414]_ , \new_[57415]_ , \new_[57416]_ ,
    \new_[57420]_ , \new_[57421]_ , \new_[57424]_ , \new_[57427]_ ,
    \new_[57428]_ , \new_[57429]_ , \new_[57433]_ , \new_[57434]_ ,
    \new_[57437]_ , \new_[57440]_ , \new_[57441]_ , \new_[57442]_ ,
    \new_[57446]_ , \new_[57447]_ , \new_[57450]_ , \new_[57453]_ ,
    \new_[57454]_ , \new_[57455]_ , \new_[57459]_ , \new_[57460]_ ,
    \new_[57463]_ , \new_[57466]_ , \new_[57467]_ , \new_[57468]_ ,
    \new_[57472]_ , \new_[57473]_ , \new_[57476]_ , \new_[57479]_ ,
    \new_[57480]_ , \new_[57481]_ , \new_[57485]_ , \new_[57486]_ ,
    \new_[57489]_ , \new_[57492]_ , \new_[57493]_ , \new_[57494]_ ,
    \new_[57498]_ , \new_[57499]_ , \new_[57502]_ , \new_[57505]_ ,
    \new_[57506]_ , \new_[57507]_ , \new_[57511]_ , \new_[57512]_ ,
    \new_[57515]_ , \new_[57518]_ , \new_[57519]_ , \new_[57520]_ ,
    \new_[57524]_ , \new_[57525]_ , \new_[57528]_ , \new_[57531]_ ,
    \new_[57532]_ , \new_[57533]_ , \new_[57537]_ , \new_[57538]_ ,
    \new_[57541]_ , \new_[57544]_ , \new_[57545]_ , \new_[57546]_ ,
    \new_[57550]_ , \new_[57551]_ , \new_[57554]_ , \new_[57557]_ ,
    \new_[57558]_ , \new_[57559]_ , \new_[57563]_ , \new_[57564]_ ,
    \new_[57567]_ , \new_[57570]_ , \new_[57571]_ , \new_[57572]_ ,
    \new_[57576]_ , \new_[57577]_ , \new_[57580]_ , \new_[57583]_ ,
    \new_[57584]_ , \new_[57585]_ , \new_[57589]_ , \new_[57590]_ ,
    \new_[57593]_ , \new_[57596]_ , \new_[57597]_ , \new_[57598]_ ,
    \new_[57602]_ , \new_[57603]_ , \new_[57606]_ , \new_[57609]_ ,
    \new_[57610]_ , \new_[57611]_ , \new_[57615]_ , \new_[57616]_ ,
    \new_[57619]_ , \new_[57622]_ , \new_[57623]_ , \new_[57624]_ ,
    \new_[57628]_ , \new_[57629]_ , \new_[57632]_ , \new_[57635]_ ,
    \new_[57636]_ , \new_[57637]_ , \new_[57641]_ , \new_[57642]_ ,
    \new_[57645]_ , \new_[57648]_ , \new_[57649]_ , \new_[57650]_ ,
    \new_[57654]_ , \new_[57655]_ , \new_[57658]_ , \new_[57661]_ ,
    \new_[57662]_ , \new_[57663]_ , \new_[57667]_ , \new_[57668]_ ,
    \new_[57671]_ , \new_[57674]_ , \new_[57675]_ , \new_[57676]_ ,
    \new_[57680]_ , \new_[57681]_ , \new_[57684]_ , \new_[57687]_ ,
    \new_[57688]_ , \new_[57689]_ , \new_[57693]_ , \new_[57694]_ ,
    \new_[57697]_ , \new_[57700]_ , \new_[57701]_ , \new_[57702]_ ,
    \new_[57706]_ , \new_[57707]_ , \new_[57710]_ , \new_[57713]_ ,
    \new_[57714]_ , \new_[57715]_ , \new_[57719]_ , \new_[57720]_ ,
    \new_[57723]_ , \new_[57726]_ , \new_[57727]_ , \new_[57728]_ ,
    \new_[57732]_ , \new_[57733]_ , \new_[57736]_ , \new_[57739]_ ,
    \new_[57740]_ , \new_[57741]_ , \new_[57745]_ , \new_[57746]_ ,
    \new_[57749]_ , \new_[57752]_ , \new_[57753]_ , \new_[57754]_ ,
    \new_[57758]_ , \new_[57759]_ , \new_[57762]_ , \new_[57765]_ ,
    \new_[57766]_ , \new_[57767]_ , \new_[57771]_ , \new_[57772]_ ,
    \new_[57775]_ , \new_[57778]_ , \new_[57779]_ , \new_[57780]_ ,
    \new_[57784]_ , \new_[57785]_ , \new_[57788]_ , \new_[57791]_ ,
    \new_[57792]_ , \new_[57793]_ , \new_[57797]_ , \new_[57798]_ ,
    \new_[57801]_ , \new_[57804]_ , \new_[57805]_ , \new_[57806]_ ,
    \new_[57810]_ , \new_[57811]_ , \new_[57814]_ , \new_[57817]_ ,
    \new_[57818]_ , \new_[57819]_ , \new_[57823]_ , \new_[57824]_ ,
    \new_[57827]_ , \new_[57830]_ , \new_[57831]_ , \new_[57832]_ ,
    \new_[57836]_ , \new_[57837]_ , \new_[57840]_ , \new_[57843]_ ,
    \new_[57844]_ , \new_[57845]_ , \new_[57849]_ , \new_[57850]_ ,
    \new_[57853]_ , \new_[57856]_ , \new_[57857]_ , \new_[57858]_ ,
    \new_[57862]_ , \new_[57863]_ , \new_[57866]_ , \new_[57869]_ ,
    \new_[57870]_ , \new_[57871]_ , \new_[57875]_ , \new_[57876]_ ,
    \new_[57879]_ , \new_[57882]_ , \new_[57883]_ , \new_[57884]_ ,
    \new_[57888]_ , \new_[57889]_ , \new_[57892]_ , \new_[57895]_ ,
    \new_[57896]_ , \new_[57897]_ , \new_[57901]_ , \new_[57902]_ ,
    \new_[57905]_ , \new_[57908]_ , \new_[57909]_ , \new_[57910]_ ,
    \new_[57914]_ , \new_[57915]_ , \new_[57918]_ , \new_[57921]_ ,
    \new_[57922]_ , \new_[57923]_ , \new_[57927]_ , \new_[57928]_ ,
    \new_[57931]_ , \new_[57934]_ , \new_[57935]_ , \new_[57936]_ ,
    \new_[57940]_ , \new_[57941]_ , \new_[57944]_ , \new_[57947]_ ,
    \new_[57948]_ , \new_[57949]_ , \new_[57953]_ , \new_[57954]_ ,
    \new_[57957]_ , \new_[57960]_ , \new_[57961]_ , \new_[57962]_ ,
    \new_[57966]_ , \new_[57967]_ , \new_[57970]_ , \new_[57973]_ ,
    \new_[57974]_ , \new_[57975]_ , \new_[57979]_ , \new_[57980]_ ,
    \new_[57983]_ , \new_[57986]_ , \new_[57987]_ , \new_[57988]_ ,
    \new_[57992]_ , \new_[57993]_ , \new_[57996]_ , \new_[57999]_ ,
    \new_[58000]_ , \new_[58001]_ , \new_[58005]_ , \new_[58006]_ ,
    \new_[58009]_ , \new_[58012]_ , \new_[58013]_ , \new_[58014]_ ,
    \new_[58018]_ , \new_[58019]_ , \new_[58022]_ , \new_[58025]_ ,
    \new_[58026]_ , \new_[58027]_ , \new_[58031]_ , \new_[58032]_ ,
    \new_[58035]_ , \new_[58038]_ , \new_[58039]_ , \new_[58040]_ ,
    \new_[58044]_ , \new_[58045]_ , \new_[58048]_ , \new_[58051]_ ,
    \new_[58052]_ , \new_[58053]_ , \new_[58057]_ , \new_[58058]_ ,
    \new_[58061]_ , \new_[58064]_ , \new_[58065]_ , \new_[58066]_ ,
    \new_[58070]_ , \new_[58071]_ , \new_[58074]_ , \new_[58077]_ ,
    \new_[58078]_ , \new_[58079]_ , \new_[58083]_ , \new_[58084]_ ,
    \new_[58087]_ , \new_[58090]_ , \new_[58091]_ , \new_[58092]_ ,
    \new_[58096]_ , \new_[58097]_ , \new_[58100]_ , \new_[58103]_ ,
    \new_[58104]_ , \new_[58105]_ , \new_[58109]_ , \new_[58110]_ ,
    \new_[58113]_ , \new_[58116]_ , \new_[58117]_ , \new_[58118]_ ,
    \new_[58122]_ , \new_[58123]_ , \new_[58126]_ , \new_[58129]_ ,
    \new_[58130]_ , \new_[58131]_ , \new_[58135]_ , \new_[58136]_ ,
    \new_[58139]_ , \new_[58142]_ , \new_[58143]_ , \new_[58144]_ ,
    \new_[58148]_ , \new_[58149]_ , \new_[58152]_ , \new_[58155]_ ,
    \new_[58156]_ , \new_[58157]_ , \new_[58161]_ , \new_[58162]_ ,
    \new_[58165]_ , \new_[58168]_ , \new_[58169]_ , \new_[58170]_ ,
    \new_[58174]_ , \new_[58175]_ , \new_[58178]_ , \new_[58181]_ ,
    \new_[58182]_ , \new_[58183]_ , \new_[58187]_ , \new_[58188]_ ,
    \new_[58191]_ , \new_[58194]_ , \new_[58195]_ , \new_[58196]_ ,
    \new_[58200]_ , \new_[58201]_ , \new_[58204]_ , \new_[58207]_ ,
    \new_[58208]_ , \new_[58209]_ , \new_[58213]_ , \new_[58214]_ ,
    \new_[58217]_ , \new_[58220]_ , \new_[58221]_ , \new_[58222]_ ,
    \new_[58226]_ , \new_[58227]_ , \new_[58230]_ , \new_[58233]_ ,
    \new_[58234]_ , \new_[58235]_ , \new_[58239]_ , \new_[58240]_ ,
    \new_[58243]_ , \new_[58246]_ , \new_[58247]_ , \new_[58248]_ ,
    \new_[58252]_ , \new_[58253]_ , \new_[58256]_ , \new_[58259]_ ,
    \new_[58260]_ , \new_[58261]_ , \new_[58265]_ , \new_[58266]_ ,
    \new_[58269]_ , \new_[58272]_ , \new_[58273]_ , \new_[58274]_ ,
    \new_[58278]_ , \new_[58279]_ , \new_[58282]_ , \new_[58285]_ ,
    \new_[58286]_ , \new_[58287]_ , \new_[58291]_ , \new_[58292]_ ,
    \new_[58295]_ , \new_[58298]_ , \new_[58299]_ , \new_[58300]_ ,
    \new_[58304]_ , \new_[58305]_ , \new_[58308]_ , \new_[58311]_ ,
    \new_[58312]_ , \new_[58313]_ , \new_[58317]_ , \new_[58318]_ ,
    \new_[58321]_ , \new_[58324]_ , \new_[58325]_ , \new_[58326]_ ,
    \new_[58330]_ , \new_[58331]_ , \new_[58334]_ , \new_[58337]_ ,
    \new_[58338]_ , \new_[58339]_ , \new_[58343]_ , \new_[58344]_ ,
    \new_[58347]_ , \new_[58350]_ , \new_[58351]_ , \new_[58352]_ ,
    \new_[58356]_ , \new_[58357]_ , \new_[58360]_ , \new_[58363]_ ,
    \new_[58364]_ , \new_[58365]_ , \new_[58369]_ , \new_[58370]_ ,
    \new_[58373]_ , \new_[58376]_ , \new_[58377]_ , \new_[58378]_ ,
    \new_[58382]_ , \new_[58383]_ , \new_[58386]_ , \new_[58389]_ ,
    \new_[58390]_ , \new_[58391]_ , \new_[58395]_ , \new_[58396]_ ,
    \new_[58399]_ , \new_[58402]_ , \new_[58403]_ , \new_[58404]_ ,
    \new_[58408]_ , \new_[58409]_ , \new_[58412]_ , \new_[58415]_ ,
    \new_[58416]_ , \new_[58417]_ , \new_[58421]_ , \new_[58422]_ ,
    \new_[58425]_ , \new_[58428]_ , \new_[58429]_ , \new_[58430]_ ,
    \new_[58434]_ , \new_[58435]_ , \new_[58438]_ , \new_[58441]_ ,
    \new_[58442]_ , \new_[58443]_ , \new_[58447]_ , \new_[58448]_ ,
    \new_[58451]_ , \new_[58454]_ , \new_[58455]_ , \new_[58456]_ ,
    \new_[58460]_ , \new_[58461]_ , \new_[58464]_ , \new_[58467]_ ,
    \new_[58468]_ , \new_[58469]_ , \new_[58473]_ , \new_[58474]_ ,
    \new_[58477]_ , \new_[58480]_ , \new_[58481]_ , \new_[58482]_ ,
    \new_[58486]_ , \new_[58487]_ , \new_[58490]_ , \new_[58493]_ ,
    \new_[58494]_ , \new_[58495]_ , \new_[58499]_ , \new_[58500]_ ,
    \new_[58503]_ , \new_[58506]_ , \new_[58507]_ , \new_[58508]_ ,
    \new_[58512]_ , \new_[58513]_ , \new_[58516]_ , \new_[58519]_ ,
    \new_[58520]_ , \new_[58521]_ , \new_[58525]_ , \new_[58526]_ ,
    \new_[58529]_ , \new_[58532]_ , \new_[58533]_ , \new_[58534]_ ,
    \new_[58538]_ , \new_[58539]_ , \new_[58542]_ , \new_[58545]_ ,
    \new_[58546]_ , \new_[58547]_ , \new_[58551]_ , \new_[58552]_ ,
    \new_[58555]_ , \new_[58558]_ , \new_[58559]_ , \new_[58560]_ ,
    \new_[58564]_ , \new_[58565]_ , \new_[58568]_ , \new_[58571]_ ,
    \new_[58572]_ , \new_[58573]_ , \new_[58577]_ , \new_[58578]_ ,
    \new_[58581]_ , \new_[58584]_ , \new_[58585]_ , \new_[58586]_ ,
    \new_[58590]_ , \new_[58591]_ , \new_[58594]_ , \new_[58597]_ ,
    \new_[58598]_ , \new_[58599]_ , \new_[58603]_ , \new_[58604]_ ,
    \new_[58607]_ , \new_[58610]_ , \new_[58611]_ , \new_[58612]_ ,
    \new_[58616]_ , \new_[58617]_ , \new_[58620]_ , \new_[58623]_ ,
    \new_[58624]_ , \new_[58625]_ , \new_[58629]_ , \new_[58630]_ ,
    \new_[58633]_ , \new_[58636]_ , \new_[58637]_ , \new_[58638]_ ,
    \new_[58642]_ , \new_[58643]_ , \new_[58646]_ , \new_[58649]_ ,
    \new_[58650]_ , \new_[58651]_ , \new_[58655]_ , \new_[58656]_ ,
    \new_[58659]_ , \new_[58662]_ , \new_[58663]_ , \new_[58664]_ ,
    \new_[58668]_ , \new_[58669]_ , \new_[58672]_ , \new_[58675]_ ,
    \new_[58676]_ , \new_[58677]_ , \new_[58681]_ , \new_[58682]_ ,
    \new_[58685]_ , \new_[58688]_ , \new_[58689]_ , \new_[58690]_ ,
    \new_[58694]_ , \new_[58695]_ , \new_[58698]_ , \new_[58701]_ ,
    \new_[58702]_ , \new_[58703]_ , \new_[58707]_ , \new_[58708]_ ,
    \new_[58711]_ , \new_[58714]_ , \new_[58715]_ , \new_[58716]_ ,
    \new_[58720]_ , \new_[58721]_ , \new_[58724]_ , \new_[58727]_ ,
    \new_[58728]_ , \new_[58729]_ , \new_[58733]_ , \new_[58734]_ ,
    \new_[58737]_ , \new_[58740]_ , \new_[58741]_ , \new_[58742]_ ,
    \new_[58746]_ , \new_[58747]_ , \new_[58750]_ , \new_[58753]_ ,
    \new_[58754]_ , \new_[58755]_ , \new_[58759]_ , \new_[58760]_ ,
    \new_[58763]_ , \new_[58766]_ , \new_[58767]_ , \new_[58768]_ ,
    \new_[58772]_ , \new_[58773]_ , \new_[58776]_ , \new_[58779]_ ,
    \new_[58780]_ , \new_[58781]_ , \new_[58785]_ , \new_[58786]_ ,
    \new_[58789]_ , \new_[58792]_ , \new_[58793]_ , \new_[58794]_ ,
    \new_[58798]_ , \new_[58799]_ , \new_[58802]_ , \new_[58805]_ ,
    \new_[58806]_ , \new_[58807]_ , \new_[58811]_ , \new_[58812]_ ,
    \new_[58815]_ , \new_[58818]_ , \new_[58819]_ , \new_[58820]_ ,
    \new_[58824]_ , \new_[58825]_ , \new_[58828]_ , \new_[58831]_ ,
    \new_[58832]_ , \new_[58833]_ , \new_[58837]_ , \new_[58838]_ ,
    \new_[58841]_ , \new_[58844]_ , \new_[58845]_ , \new_[58846]_ ,
    \new_[58850]_ , \new_[58851]_ , \new_[58854]_ , \new_[58857]_ ,
    \new_[58858]_ , \new_[58859]_ , \new_[58863]_ , \new_[58864]_ ,
    \new_[58867]_ , \new_[58870]_ , \new_[58871]_ , \new_[58872]_ ,
    \new_[58876]_ , \new_[58877]_ , \new_[58880]_ , \new_[58883]_ ,
    \new_[58884]_ , \new_[58885]_ , \new_[58889]_ , \new_[58890]_ ,
    \new_[58893]_ , \new_[58896]_ , \new_[58897]_ , \new_[58898]_ ,
    \new_[58902]_ , \new_[58903]_ , \new_[58906]_ , \new_[58909]_ ,
    \new_[58910]_ , \new_[58911]_ , \new_[58915]_ , \new_[58916]_ ,
    \new_[58919]_ , \new_[58922]_ , \new_[58923]_ , \new_[58924]_ ,
    \new_[58928]_ , \new_[58929]_ , \new_[58932]_ , \new_[58935]_ ,
    \new_[58936]_ , \new_[58937]_ , \new_[58941]_ , \new_[58942]_ ,
    \new_[58945]_ , \new_[58948]_ , \new_[58949]_ , \new_[58950]_ ,
    \new_[58954]_ , \new_[58955]_ , \new_[58958]_ , \new_[58961]_ ,
    \new_[58962]_ , \new_[58963]_ , \new_[58967]_ , \new_[58968]_ ,
    \new_[58971]_ , \new_[58974]_ , \new_[58975]_ , \new_[58976]_ ,
    \new_[58980]_ , \new_[58981]_ , \new_[58984]_ , \new_[58987]_ ,
    \new_[58988]_ , \new_[58989]_ , \new_[58993]_ , \new_[58994]_ ,
    \new_[58997]_ , \new_[59000]_ , \new_[59001]_ , \new_[59002]_ ,
    \new_[59006]_ , \new_[59007]_ , \new_[59010]_ , \new_[59013]_ ,
    \new_[59014]_ , \new_[59015]_ , \new_[59019]_ , \new_[59020]_ ,
    \new_[59023]_ , \new_[59026]_ , \new_[59027]_ , \new_[59028]_ ,
    \new_[59032]_ , \new_[59033]_ , \new_[59036]_ , \new_[59039]_ ,
    \new_[59040]_ , \new_[59041]_ , \new_[59045]_ , \new_[59046]_ ,
    \new_[59049]_ , \new_[59052]_ , \new_[59053]_ , \new_[59054]_ ,
    \new_[59058]_ , \new_[59059]_ , \new_[59062]_ , \new_[59065]_ ,
    \new_[59066]_ , \new_[59067]_ , \new_[59071]_ , \new_[59072]_ ,
    \new_[59075]_ , \new_[59078]_ , \new_[59079]_ , \new_[59080]_ ,
    \new_[59084]_ , \new_[59085]_ , \new_[59088]_ , \new_[59091]_ ,
    \new_[59092]_ , \new_[59093]_ , \new_[59097]_ , \new_[59098]_ ,
    \new_[59101]_ , \new_[59104]_ , \new_[59105]_ , \new_[59106]_ ,
    \new_[59110]_ , \new_[59111]_ , \new_[59114]_ , \new_[59117]_ ,
    \new_[59118]_ , \new_[59119]_ , \new_[59123]_ , \new_[59124]_ ,
    \new_[59127]_ , \new_[59130]_ , \new_[59131]_ , \new_[59132]_ ,
    \new_[59136]_ , \new_[59137]_ , \new_[59140]_ , \new_[59143]_ ,
    \new_[59144]_ , \new_[59145]_ , \new_[59149]_ , \new_[59150]_ ,
    \new_[59153]_ , \new_[59156]_ , \new_[59157]_ , \new_[59158]_ ,
    \new_[59162]_ , \new_[59163]_ , \new_[59166]_ , \new_[59169]_ ,
    \new_[59170]_ , \new_[59171]_ , \new_[59175]_ , \new_[59176]_ ,
    \new_[59179]_ , \new_[59182]_ , \new_[59183]_ , \new_[59184]_ ,
    \new_[59188]_ , \new_[59189]_ , \new_[59192]_ , \new_[59195]_ ,
    \new_[59196]_ , \new_[59197]_ , \new_[59201]_ , \new_[59202]_ ,
    \new_[59205]_ , \new_[59208]_ , \new_[59209]_ , \new_[59210]_ ,
    \new_[59214]_ , \new_[59215]_ , \new_[59218]_ , \new_[59221]_ ,
    \new_[59222]_ , \new_[59223]_ , \new_[59227]_ , \new_[59228]_ ,
    \new_[59231]_ , \new_[59234]_ , \new_[59235]_ , \new_[59236]_ ,
    \new_[59240]_ , \new_[59241]_ , \new_[59244]_ , \new_[59247]_ ,
    \new_[59248]_ , \new_[59249]_ , \new_[59253]_ , \new_[59254]_ ,
    \new_[59257]_ , \new_[59260]_ , \new_[59261]_ , \new_[59262]_ ,
    \new_[59266]_ , \new_[59267]_ , \new_[59270]_ , \new_[59273]_ ,
    \new_[59274]_ , \new_[59275]_ , \new_[59279]_ , \new_[59280]_ ,
    \new_[59283]_ , \new_[59286]_ , \new_[59287]_ , \new_[59288]_ ,
    \new_[59292]_ , \new_[59293]_ , \new_[59296]_ , \new_[59299]_ ,
    \new_[59300]_ , \new_[59301]_ , \new_[59305]_ , \new_[59306]_ ,
    \new_[59309]_ , \new_[59312]_ , \new_[59313]_ , \new_[59314]_ ,
    \new_[59318]_ , \new_[59319]_ , \new_[59322]_ , \new_[59325]_ ,
    \new_[59326]_ , \new_[59327]_ , \new_[59331]_ , \new_[59332]_ ,
    \new_[59335]_ , \new_[59338]_ , \new_[59339]_ , \new_[59340]_ ,
    \new_[59344]_ , \new_[59345]_ , \new_[59348]_ , \new_[59351]_ ,
    \new_[59352]_ , \new_[59353]_ , \new_[59357]_ , \new_[59358]_ ,
    \new_[59361]_ , \new_[59364]_ , \new_[59365]_ , \new_[59366]_ ,
    \new_[59370]_ , \new_[59371]_ , \new_[59374]_ , \new_[59377]_ ,
    \new_[59378]_ , \new_[59379]_ , \new_[59383]_ , \new_[59384]_ ,
    \new_[59387]_ , \new_[59390]_ , \new_[59391]_ , \new_[59392]_ ,
    \new_[59396]_ , \new_[59397]_ , \new_[59400]_ , \new_[59403]_ ,
    \new_[59404]_ , \new_[59405]_ , \new_[59409]_ , \new_[59410]_ ,
    \new_[59413]_ , \new_[59416]_ , \new_[59417]_ , \new_[59418]_ ,
    \new_[59422]_ , \new_[59423]_ , \new_[59426]_ , \new_[59429]_ ,
    \new_[59430]_ , \new_[59431]_ , \new_[59435]_ , \new_[59436]_ ,
    \new_[59439]_ , \new_[59442]_ , \new_[59443]_ , \new_[59444]_ ,
    \new_[59448]_ , \new_[59449]_ , \new_[59452]_ , \new_[59455]_ ,
    \new_[59456]_ , \new_[59457]_ , \new_[59461]_ , \new_[59462]_ ,
    \new_[59465]_ , \new_[59468]_ , \new_[59469]_ , \new_[59470]_ ,
    \new_[59474]_ , \new_[59475]_ , \new_[59478]_ , \new_[59481]_ ,
    \new_[59482]_ , \new_[59483]_ , \new_[59487]_ , \new_[59488]_ ,
    \new_[59491]_ , \new_[59494]_ , \new_[59495]_ , \new_[59496]_ ,
    \new_[59500]_ , \new_[59501]_ , \new_[59504]_ , \new_[59507]_ ,
    \new_[59508]_ , \new_[59509]_ , \new_[59513]_ , \new_[59514]_ ,
    \new_[59517]_ , \new_[59520]_ , \new_[59521]_ , \new_[59522]_ ,
    \new_[59526]_ , \new_[59527]_ , \new_[59530]_ , \new_[59533]_ ,
    \new_[59534]_ , \new_[59535]_ , \new_[59539]_ , \new_[59540]_ ,
    \new_[59543]_ , \new_[59546]_ , \new_[59547]_ , \new_[59548]_ ,
    \new_[59552]_ , \new_[59553]_ , \new_[59556]_ , \new_[59559]_ ,
    \new_[59560]_ , \new_[59561]_ , \new_[59565]_ , \new_[59566]_ ,
    \new_[59569]_ , \new_[59572]_ , \new_[59573]_ , \new_[59574]_ ,
    \new_[59578]_ , \new_[59579]_ , \new_[59582]_ , \new_[59585]_ ,
    \new_[59586]_ , \new_[59587]_ , \new_[59591]_ , \new_[59592]_ ,
    \new_[59595]_ , \new_[59598]_ , \new_[59599]_ , \new_[59600]_ ,
    \new_[59604]_ , \new_[59605]_ , \new_[59608]_ , \new_[59611]_ ,
    \new_[59612]_ , \new_[59613]_ , \new_[59617]_ , \new_[59618]_ ,
    \new_[59621]_ , \new_[59624]_ , \new_[59625]_ , \new_[59626]_ ,
    \new_[59630]_ , \new_[59631]_ , \new_[59634]_ , \new_[59637]_ ,
    \new_[59638]_ , \new_[59639]_ , \new_[59643]_ , \new_[59644]_ ,
    \new_[59647]_ , \new_[59650]_ , \new_[59651]_ , \new_[59652]_ ,
    \new_[59656]_ , \new_[59657]_ , \new_[59660]_ , \new_[59663]_ ,
    \new_[59664]_ , \new_[59665]_ , \new_[59669]_ , \new_[59670]_ ,
    \new_[59673]_ , \new_[59676]_ , \new_[59677]_ , \new_[59678]_ ,
    \new_[59682]_ , \new_[59683]_ , \new_[59686]_ , \new_[59689]_ ,
    \new_[59690]_ , \new_[59691]_ , \new_[59695]_ , \new_[59696]_ ,
    \new_[59699]_ , \new_[59702]_ , \new_[59703]_ , \new_[59704]_ ,
    \new_[59708]_ , \new_[59709]_ , \new_[59712]_ , \new_[59715]_ ,
    \new_[59716]_ , \new_[59717]_ , \new_[59721]_ , \new_[59722]_ ,
    \new_[59725]_ , \new_[59728]_ , \new_[59729]_ , \new_[59730]_ ,
    \new_[59734]_ , \new_[59735]_ , \new_[59738]_ , \new_[59741]_ ,
    \new_[59742]_ , \new_[59743]_ , \new_[59747]_ , \new_[59748]_ ,
    \new_[59751]_ , \new_[59754]_ , \new_[59755]_ , \new_[59756]_ ,
    \new_[59760]_ , \new_[59761]_ , \new_[59764]_ , \new_[59767]_ ,
    \new_[59768]_ , \new_[59769]_ , \new_[59773]_ , \new_[59774]_ ,
    \new_[59777]_ , \new_[59780]_ , \new_[59781]_ , \new_[59782]_ ,
    \new_[59786]_ , \new_[59787]_ , \new_[59790]_ , \new_[59793]_ ,
    \new_[59794]_ , \new_[59795]_ , \new_[59799]_ , \new_[59800]_ ,
    \new_[59803]_ , \new_[59806]_ , \new_[59807]_ , \new_[59808]_ ,
    \new_[59812]_ , \new_[59813]_ , \new_[59816]_ , \new_[59819]_ ,
    \new_[59820]_ , \new_[59821]_ , \new_[59825]_ , \new_[59826]_ ,
    \new_[59829]_ , \new_[59832]_ , \new_[59833]_ , \new_[59834]_ ,
    \new_[59838]_ , \new_[59839]_ , \new_[59842]_ , \new_[59845]_ ,
    \new_[59846]_ , \new_[59847]_ , \new_[59851]_ , \new_[59852]_ ,
    \new_[59855]_ , \new_[59858]_ , \new_[59859]_ , \new_[59860]_ ,
    \new_[59864]_ , \new_[59865]_ , \new_[59868]_ , \new_[59871]_ ,
    \new_[59872]_ , \new_[59873]_ , \new_[59877]_ , \new_[59878]_ ,
    \new_[59881]_ , \new_[59884]_ , \new_[59885]_ , \new_[59886]_ ,
    \new_[59890]_ , \new_[59891]_ , \new_[59894]_ , \new_[59897]_ ,
    \new_[59898]_ , \new_[59899]_ , \new_[59903]_ , \new_[59904]_ ,
    \new_[59907]_ , \new_[59910]_ , \new_[59911]_ , \new_[59912]_ ,
    \new_[59916]_ , \new_[59917]_ , \new_[59920]_ , \new_[59923]_ ,
    \new_[59924]_ , \new_[59925]_ , \new_[59929]_ , \new_[59930]_ ,
    \new_[59933]_ , \new_[59936]_ , \new_[59937]_ , \new_[59938]_ ,
    \new_[59942]_ , \new_[59943]_ , \new_[59946]_ , \new_[59949]_ ,
    \new_[59950]_ , \new_[59951]_ , \new_[59955]_ , \new_[59956]_ ,
    \new_[59959]_ , \new_[59962]_ , \new_[59963]_ , \new_[59964]_ ,
    \new_[59968]_ , \new_[59969]_ , \new_[59972]_ , \new_[59975]_ ,
    \new_[59976]_ , \new_[59977]_ , \new_[59981]_ , \new_[59982]_ ,
    \new_[59985]_ , \new_[59988]_ , \new_[59989]_ , \new_[59990]_ ,
    \new_[59994]_ , \new_[59995]_ , \new_[59998]_ , \new_[60001]_ ,
    \new_[60002]_ , \new_[60003]_ , \new_[60007]_ , \new_[60008]_ ,
    \new_[60011]_ , \new_[60014]_ , \new_[60015]_ , \new_[60016]_ ,
    \new_[60020]_ , \new_[60021]_ , \new_[60024]_ , \new_[60027]_ ,
    \new_[60028]_ , \new_[60029]_ , \new_[60033]_ , \new_[60034]_ ,
    \new_[60037]_ , \new_[60040]_ , \new_[60041]_ , \new_[60042]_ ,
    \new_[60046]_ , \new_[60047]_ , \new_[60050]_ , \new_[60053]_ ,
    \new_[60054]_ , \new_[60055]_ , \new_[60059]_ , \new_[60060]_ ,
    \new_[60063]_ , \new_[60066]_ , \new_[60067]_ , \new_[60068]_ ,
    \new_[60072]_ , \new_[60073]_ , \new_[60076]_ , \new_[60079]_ ,
    \new_[60080]_ , \new_[60081]_ , \new_[60085]_ , \new_[60086]_ ,
    \new_[60089]_ , \new_[60092]_ , \new_[60093]_ , \new_[60094]_ ,
    \new_[60098]_ , \new_[60099]_ , \new_[60102]_ , \new_[60105]_ ,
    \new_[60106]_ , \new_[60107]_ , \new_[60111]_ , \new_[60112]_ ,
    \new_[60115]_ , \new_[60118]_ , \new_[60119]_ , \new_[60120]_ ,
    \new_[60124]_ , \new_[60125]_ , \new_[60128]_ , \new_[60131]_ ,
    \new_[60132]_ , \new_[60133]_ , \new_[60137]_ , \new_[60138]_ ,
    \new_[60141]_ , \new_[60144]_ , \new_[60145]_ , \new_[60146]_ ,
    \new_[60150]_ , \new_[60151]_ , \new_[60154]_ , \new_[60157]_ ,
    \new_[60158]_ , \new_[60159]_ , \new_[60163]_ , \new_[60164]_ ,
    \new_[60167]_ , \new_[60170]_ , \new_[60171]_ , \new_[60172]_ ,
    \new_[60176]_ , \new_[60177]_ , \new_[60180]_ , \new_[60183]_ ,
    \new_[60184]_ , \new_[60185]_ , \new_[60189]_ , \new_[60190]_ ,
    \new_[60193]_ , \new_[60196]_ , \new_[60197]_ , \new_[60198]_ ,
    \new_[60202]_ , \new_[60203]_ , \new_[60206]_ , \new_[60209]_ ,
    \new_[60210]_ , \new_[60211]_ , \new_[60215]_ , \new_[60216]_ ,
    \new_[60219]_ , \new_[60222]_ , \new_[60223]_ , \new_[60224]_ ,
    \new_[60228]_ , \new_[60229]_ , \new_[60232]_ , \new_[60235]_ ,
    \new_[60236]_ , \new_[60237]_ , \new_[60241]_ , \new_[60242]_ ,
    \new_[60245]_ , \new_[60248]_ , \new_[60249]_ , \new_[60250]_ ,
    \new_[60254]_ , \new_[60255]_ , \new_[60258]_ , \new_[60261]_ ,
    \new_[60262]_ , \new_[60263]_ , \new_[60267]_ , \new_[60268]_ ,
    \new_[60271]_ , \new_[60274]_ , \new_[60275]_ , \new_[60276]_ ,
    \new_[60280]_ , \new_[60281]_ , \new_[60284]_ , \new_[60287]_ ,
    \new_[60288]_ , \new_[60289]_ , \new_[60292]_ , \new_[60295]_ ,
    \new_[60296]_ , \new_[60299]_ , \new_[60302]_ , \new_[60303]_ ,
    \new_[60304]_ , \new_[60308]_ , \new_[60309]_ , \new_[60312]_ ,
    \new_[60315]_ , \new_[60316]_ , \new_[60317]_ , \new_[60320]_ ,
    \new_[60323]_ , \new_[60324]_ , \new_[60327]_ , \new_[60330]_ ,
    \new_[60331]_ , \new_[60332]_ , \new_[60336]_ , \new_[60337]_ ,
    \new_[60340]_ , \new_[60343]_ , \new_[60344]_ , \new_[60345]_ ,
    \new_[60348]_ , \new_[60351]_ , \new_[60352]_ , \new_[60355]_ ,
    \new_[60358]_ , \new_[60359]_ , \new_[60360]_ , \new_[60364]_ ,
    \new_[60365]_ , \new_[60368]_ , \new_[60371]_ , \new_[60372]_ ,
    \new_[60373]_ , \new_[60376]_ , \new_[60379]_ , \new_[60380]_ ,
    \new_[60383]_ , \new_[60386]_ , \new_[60387]_ , \new_[60388]_ ,
    \new_[60392]_ , \new_[60393]_ , \new_[60396]_ , \new_[60399]_ ,
    \new_[60400]_ , \new_[60401]_ , \new_[60404]_ , \new_[60407]_ ,
    \new_[60408]_ , \new_[60411]_ , \new_[60414]_ , \new_[60415]_ ,
    \new_[60416]_ , \new_[60420]_ , \new_[60421]_ , \new_[60424]_ ,
    \new_[60427]_ , \new_[60428]_ , \new_[60429]_ , \new_[60432]_ ,
    \new_[60435]_ , \new_[60436]_ , \new_[60439]_ , \new_[60442]_ ,
    \new_[60443]_ , \new_[60444]_ , \new_[60448]_ , \new_[60449]_ ,
    \new_[60452]_ , \new_[60455]_ , \new_[60456]_ , \new_[60457]_ ,
    \new_[60460]_ , \new_[60463]_ , \new_[60464]_ , \new_[60467]_ ,
    \new_[60470]_ , \new_[60471]_ , \new_[60472]_ , \new_[60476]_ ,
    \new_[60477]_ , \new_[60480]_ , \new_[60483]_ , \new_[60484]_ ,
    \new_[60485]_ , \new_[60488]_ , \new_[60491]_ , \new_[60492]_ ,
    \new_[60495]_ , \new_[60498]_ , \new_[60499]_ , \new_[60500]_ ,
    \new_[60504]_ , \new_[60505]_ , \new_[60508]_ , \new_[60511]_ ,
    \new_[60512]_ , \new_[60513]_ , \new_[60516]_ , \new_[60519]_ ,
    \new_[60520]_ , \new_[60523]_ , \new_[60526]_ , \new_[60527]_ ,
    \new_[60528]_ , \new_[60532]_ , \new_[60533]_ , \new_[60536]_ ,
    \new_[60539]_ , \new_[60540]_ , \new_[60541]_ , \new_[60544]_ ,
    \new_[60547]_ , \new_[60548]_ , \new_[60551]_ , \new_[60554]_ ,
    \new_[60555]_ , \new_[60556]_ , \new_[60560]_ , \new_[60561]_ ,
    \new_[60564]_ , \new_[60567]_ , \new_[60568]_ , \new_[60569]_ ,
    \new_[60572]_ , \new_[60575]_ , \new_[60576]_ , \new_[60579]_ ,
    \new_[60582]_ , \new_[60583]_ , \new_[60584]_ , \new_[60588]_ ,
    \new_[60589]_ , \new_[60592]_ , \new_[60595]_ , \new_[60596]_ ,
    \new_[60597]_ , \new_[60600]_ , \new_[60603]_ , \new_[60604]_ ,
    \new_[60607]_ , \new_[60610]_ , \new_[60611]_ , \new_[60612]_ ,
    \new_[60616]_ , \new_[60617]_ , \new_[60620]_ , \new_[60623]_ ,
    \new_[60624]_ , \new_[60625]_ , \new_[60628]_ , \new_[60631]_ ,
    \new_[60632]_ , \new_[60635]_ , \new_[60638]_ , \new_[60639]_ ,
    \new_[60640]_ , \new_[60644]_ , \new_[60645]_ , \new_[60648]_ ,
    \new_[60651]_ , \new_[60652]_ , \new_[60653]_ , \new_[60656]_ ,
    \new_[60659]_ , \new_[60660]_ , \new_[60663]_ , \new_[60666]_ ,
    \new_[60667]_ , \new_[60668]_ , \new_[60672]_ , \new_[60673]_ ,
    \new_[60676]_ , \new_[60679]_ , \new_[60680]_ , \new_[60681]_ ,
    \new_[60684]_ , \new_[60687]_ , \new_[60688]_ , \new_[60691]_ ,
    \new_[60694]_ , \new_[60695]_ , \new_[60696]_ , \new_[60700]_ ,
    \new_[60701]_ , \new_[60704]_ , \new_[60707]_ , \new_[60708]_ ,
    \new_[60709]_ , \new_[60712]_ , \new_[60715]_ , \new_[60716]_ ,
    \new_[60719]_ , \new_[60722]_ , \new_[60723]_ , \new_[60724]_ ,
    \new_[60728]_ , \new_[60729]_ , \new_[60732]_ , \new_[60735]_ ,
    \new_[60736]_ , \new_[60737]_ , \new_[60740]_ , \new_[60743]_ ,
    \new_[60744]_ , \new_[60747]_ , \new_[60750]_ , \new_[60751]_ ,
    \new_[60752]_ , \new_[60756]_ , \new_[60757]_ , \new_[60760]_ ,
    \new_[60763]_ , \new_[60764]_ , \new_[60765]_ , \new_[60768]_ ,
    \new_[60771]_ , \new_[60772]_ , \new_[60775]_ , \new_[60778]_ ,
    \new_[60779]_ , \new_[60780]_ , \new_[60784]_ , \new_[60785]_ ,
    \new_[60788]_ , \new_[60791]_ , \new_[60792]_ , \new_[60793]_ ,
    \new_[60796]_ , \new_[60799]_ , \new_[60800]_ , \new_[60803]_ ,
    \new_[60806]_ , \new_[60807]_ , \new_[60808]_ , \new_[60812]_ ,
    \new_[60813]_ , \new_[60816]_ , \new_[60819]_ , \new_[60820]_ ,
    \new_[60821]_ , \new_[60824]_ , \new_[60827]_ , \new_[60828]_ ,
    \new_[60831]_ , \new_[60834]_ , \new_[60835]_ , \new_[60836]_ ,
    \new_[60840]_ , \new_[60841]_ , \new_[60844]_ , \new_[60847]_ ,
    \new_[60848]_ , \new_[60849]_ , \new_[60852]_ , \new_[60855]_ ,
    \new_[60856]_ , \new_[60859]_ , \new_[60862]_ , \new_[60863]_ ,
    \new_[60864]_ , \new_[60868]_ , \new_[60869]_ , \new_[60872]_ ,
    \new_[60875]_ , \new_[60876]_ , \new_[60877]_ , \new_[60880]_ ,
    \new_[60883]_ , \new_[60884]_ , \new_[60887]_ , \new_[60890]_ ,
    \new_[60891]_ , \new_[60892]_ , \new_[60896]_ , \new_[60897]_ ,
    \new_[60900]_ , \new_[60903]_ , \new_[60904]_ , \new_[60905]_ ,
    \new_[60908]_ , \new_[60911]_ , \new_[60912]_ , \new_[60915]_ ,
    \new_[60918]_ , \new_[60919]_ , \new_[60920]_ , \new_[60924]_ ,
    \new_[60925]_ , \new_[60928]_ , \new_[60931]_ , \new_[60932]_ ,
    \new_[60933]_ , \new_[60936]_ , \new_[60939]_ , \new_[60940]_ ,
    \new_[60943]_ , \new_[60946]_ , \new_[60947]_ , \new_[60948]_ ,
    \new_[60952]_ , \new_[60953]_ , \new_[60956]_ , \new_[60959]_ ,
    \new_[60960]_ , \new_[60961]_ , \new_[60964]_ , \new_[60967]_ ,
    \new_[60968]_ , \new_[60971]_ , \new_[60974]_ , \new_[60975]_ ,
    \new_[60976]_ , \new_[60980]_ , \new_[60981]_ , \new_[60984]_ ,
    \new_[60987]_ , \new_[60988]_ , \new_[60989]_ , \new_[60992]_ ,
    \new_[60995]_ , \new_[60996]_ , \new_[60999]_ , \new_[61002]_ ,
    \new_[61003]_ , \new_[61004]_ , \new_[61008]_ , \new_[61009]_ ,
    \new_[61012]_ , \new_[61015]_ , \new_[61016]_ , \new_[61017]_ ,
    \new_[61020]_ , \new_[61023]_ , \new_[61024]_ , \new_[61027]_ ,
    \new_[61030]_ , \new_[61031]_ , \new_[61032]_ , \new_[61036]_ ,
    \new_[61037]_ , \new_[61040]_ , \new_[61043]_ , \new_[61044]_ ,
    \new_[61045]_ , \new_[61048]_ , \new_[61051]_ , \new_[61052]_ ,
    \new_[61055]_ , \new_[61058]_ , \new_[61059]_ , \new_[61060]_ ,
    \new_[61064]_ , \new_[61065]_ , \new_[61068]_ , \new_[61071]_ ,
    \new_[61072]_ , \new_[61073]_ , \new_[61076]_ , \new_[61079]_ ,
    \new_[61080]_ , \new_[61083]_ , \new_[61086]_ , \new_[61087]_ ,
    \new_[61088]_ , \new_[61092]_ , \new_[61093]_ , \new_[61096]_ ,
    \new_[61099]_ , \new_[61100]_ , \new_[61101]_ , \new_[61104]_ ,
    \new_[61107]_ , \new_[61108]_ , \new_[61111]_ , \new_[61114]_ ,
    \new_[61115]_ , \new_[61116]_ , \new_[61120]_ , \new_[61121]_ ,
    \new_[61124]_ , \new_[61127]_ , \new_[61128]_ , \new_[61129]_ ,
    \new_[61132]_ , \new_[61135]_ , \new_[61136]_ , \new_[61139]_ ,
    \new_[61142]_ , \new_[61143]_ , \new_[61144]_ , \new_[61148]_ ,
    \new_[61149]_ , \new_[61152]_ , \new_[61155]_ , \new_[61156]_ ,
    \new_[61157]_ , \new_[61160]_ , \new_[61163]_ , \new_[61164]_ ,
    \new_[61167]_ , \new_[61170]_ , \new_[61171]_ , \new_[61172]_ ,
    \new_[61176]_ , \new_[61177]_ , \new_[61180]_ , \new_[61183]_ ,
    \new_[61184]_ , \new_[61185]_ , \new_[61188]_ , \new_[61191]_ ,
    \new_[61192]_ , \new_[61195]_ , \new_[61198]_ , \new_[61199]_ ,
    \new_[61200]_ , \new_[61204]_ , \new_[61205]_ , \new_[61208]_ ,
    \new_[61211]_ , \new_[61212]_ , \new_[61213]_ , \new_[61216]_ ,
    \new_[61219]_ , \new_[61220]_ , \new_[61223]_ , \new_[61226]_ ,
    \new_[61227]_ , \new_[61228]_ , \new_[61232]_ , \new_[61233]_ ,
    \new_[61236]_ , \new_[61239]_ , \new_[61240]_ , \new_[61241]_ ,
    \new_[61244]_ , \new_[61247]_ , \new_[61248]_ , \new_[61251]_ ,
    \new_[61254]_ , \new_[61255]_ , \new_[61256]_ , \new_[61260]_ ,
    \new_[61261]_ , \new_[61264]_ , \new_[61267]_ , \new_[61268]_ ,
    \new_[61269]_ , \new_[61272]_ , \new_[61275]_ , \new_[61276]_ ,
    \new_[61279]_ , \new_[61282]_ , \new_[61283]_ , \new_[61284]_ ,
    \new_[61288]_ , \new_[61289]_ , \new_[61292]_ , \new_[61295]_ ,
    \new_[61296]_ , \new_[61297]_ , \new_[61300]_ , \new_[61303]_ ,
    \new_[61304]_ , \new_[61307]_ , \new_[61310]_ , \new_[61311]_ ,
    \new_[61312]_ , \new_[61316]_ , \new_[61317]_ , \new_[61320]_ ,
    \new_[61323]_ , \new_[61324]_ , \new_[61325]_ , \new_[61328]_ ,
    \new_[61331]_ , \new_[61332]_ , \new_[61335]_ , \new_[61338]_ ,
    \new_[61339]_ , \new_[61340]_ , \new_[61344]_ , \new_[61345]_ ,
    \new_[61348]_ , \new_[61351]_ , \new_[61352]_ , \new_[61353]_ ,
    \new_[61356]_ , \new_[61359]_ , \new_[61360]_ , \new_[61363]_ ,
    \new_[61366]_ , \new_[61367]_ , \new_[61368]_ , \new_[61372]_ ,
    \new_[61373]_ , \new_[61376]_ , \new_[61379]_ , \new_[61380]_ ,
    \new_[61381]_ , \new_[61384]_ , \new_[61387]_ , \new_[61388]_ ,
    \new_[61391]_ , \new_[61394]_ , \new_[61395]_ , \new_[61396]_ ,
    \new_[61400]_ , \new_[61401]_ , \new_[61404]_ , \new_[61407]_ ,
    \new_[61408]_ , \new_[61409]_ , \new_[61412]_ , \new_[61415]_ ,
    \new_[61416]_ , \new_[61419]_ , \new_[61422]_ , \new_[61423]_ ,
    \new_[61424]_ , \new_[61428]_ , \new_[61429]_ , \new_[61432]_ ,
    \new_[61435]_ , \new_[61436]_ , \new_[61437]_ , \new_[61440]_ ,
    \new_[61443]_ , \new_[61444]_ , \new_[61447]_ , \new_[61450]_ ,
    \new_[61451]_ , \new_[61452]_ , \new_[61456]_ , \new_[61457]_ ,
    \new_[61460]_ , \new_[61463]_ , \new_[61464]_ , \new_[61465]_ ,
    \new_[61468]_ , \new_[61471]_ , \new_[61472]_ , \new_[61475]_ ,
    \new_[61478]_ , \new_[61479]_ , \new_[61480]_ , \new_[61484]_ ,
    \new_[61485]_ , \new_[61488]_ , \new_[61491]_ , \new_[61492]_ ,
    \new_[61493]_ , \new_[61496]_ , \new_[61499]_ , \new_[61500]_ ,
    \new_[61503]_ , \new_[61506]_ , \new_[61507]_ , \new_[61508]_ ,
    \new_[61512]_ , \new_[61513]_ , \new_[61516]_ , \new_[61519]_ ,
    \new_[61520]_ , \new_[61521]_ , \new_[61524]_ , \new_[61527]_ ,
    \new_[61528]_ , \new_[61531]_ , \new_[61534]_ , \new_[61535]_ ,
    \new_[61536]_ , \new_[61540]_ , \new_[61541]_ , \new_[61544]_ ,
    \new_[61547]_ , \new_[61548]_ , \new_[61549]_ , \new_[61552]_ ,
    \new_[61555]_ , \new_[61556]_ , \new_[61559]_ , \new_[61562]_ ,
    \new_[61563]_ , \new_[61564]_ , \new_[61568]_ , \new_[61569]_ ,
    \new_[61572]_ , \new_[61575]_ , \new_[61576]_ , \new_[61577]_ ,
    \new_[61580]_ , \new_[61583]_ , \new_[61584]_ , \new_[61587]_ ,
    \new_[61590]_ , \new_[61591]_ , \new_[61592]_ , \new_[61596]_ ,
    \new_[61597]_ , \new_[61600]_ , \new_[61603]_ , \new_[61604]_ ,
    \new_[61605]_ , \new_[61608]_ , \new_[61611]_ , \new_[61612]_ ,
    \new_[61615]_ , \new_[61618]_ , \new_[61619]_ , \new_[61620]_ ,
    \new_[61624]_ , \new_[61625]_ , \new_[61628]_ , \new_[61631]_ ,
    \new_[61632]_ , \new_[61633]_ , \new_[61636]_ , \new_[61639]_ ,
    \new_[61640]_ , \new_[61643]_ , \new_[61646]_ , \new_[61647]_ ,
    \new_[61648]_ , \new_[61652]_ , \new_[61653]_ , \new_[61656]_ ,
    \new_[61659]_ , \new_[61660]_ , \new_[61661]_ , \new_[61664]_ ,
    \new_[61667]_ , \new_[61668]_ , \new_[61671]_ , \new_[61674]_ ,
    \new_[61675]_ , \new_[61676]_ , \new_[61680]_ , \new_[61681]_ ,
    \new_[61684]_ , \new_[61687]_ , \new_[61688]_ , \new_[61689]_ ,
    \new_[61692]_ , \new_[61695]_ , \new_[61696]_ , \new_[61699]_ ,
    \new_[61702]_ , \new_[61703]_ , \new_[61704]_ , \new_[61708]_ ,
    \new_[61709]_ , \new_[61712]_ , \new_[61715]_ , \new_[61716]_ ,
    \new_[61717]_ , \new_[61720]_ , \new_[61723]_ , \new_[61724]_ ,
    \new_[61727]_ , \new_[61730]_ , \new_[61731]_ , \new_[61732]_ ,
    \new_[61736]_ , \new_[61737]_ , \new_[61740]_ , \new_[61743]_ ,
    \new_[61744]_ , \new_[61745]_ , \new_[61748]_ , \new_[61751]_ ,
    \new_[61752]_ , \new_[61755]_ , \new_[61758]_ , \new_[61759]_ ,
    \new_[61760]_ , \new_[61764]_ , \new_[61765]_ , \new_[61768]_ ,
    \new_[61771]_ , \new_[61772]_ , \new_[61773]_ , \new_[61776]_ ,
    \new_[61779]_ , \new_[61780]_ , \new_[61783]_ , \new_[61786]_ ,
    \new_[61787]_ , \new_[61788]_ , \new_[61792]_ , \new_[61793]_ ,
    \new_[61796]_ , \new_[61799]_ , \new_[61800]_ , \new_[61801]_ ,
    \new_[61804]_ , \new_[61807]_ , \new_[61808]_ , \new_[61811]_ ,
    \new_[61814]_ , \new_[61815]_ , \new_[61816]_ , \new_[61820]_ ,
    \new_[61821]_ , \new_[61824]_ , \new_[61827]_ , \new_[61828]_ ,
    \new_[61829]_ , \new_[61832]_ , \new_[61835]_ , \new_[61836]_ ,
    \new_[61839]_ , \new_[61842]_ , \new_[61843]_ , \new_[61844]_ ,
    \new_[61848]_ , \new_[61849]_ , \new_[61852]_ , \new_[61855]_ ,
    \new_[61856]_ , \new_[61857]_ , \new_[61860]_ , \new_[61863]_ ,
    \new_[61864]_ , \new_[61867]_ , \new_[61870]_ , \new_[61871]_ ,
    \new_[61872]_ , \new_[61876]_ , \new_[61877]_ , \new_[61880]_ ,
    \new_[61883]_ , \new_[61884]_ , \new_[61885]_ , \new_[61888]_ ,
    \new_[61891]_ , \new_[61892]_ , \new_[61895]_ , \new_[61898]_ ,
    \new_[61899]_ , \new_[61900]_ , \new_[61904]_ , \new_[61905]_ ,
    \new_[61908]_ , \new_[61911]_ , \new_[61912]_ , \new_[61913]_ ,
    \new_[61916]_ , \new_[61919]_ , \new_[61920]_ , \new_[61923]_ ,
    \new_[61926]_ , \new_[61927]_ , \new_[61928]_ , \new_[61932]_ ,
    \new_[61933]_ , \new_[61936]_ , \new_[61939]_ , \new_[61940]_ ,
    \new_[61941]_ , \new_[61944]_ , \new_[61947]_ , \new_[61948]_ ,
    \new_[61951]_ , \new_[61954]_ , \new_[61955]_ , \new_[61956]_ ,
    \new_[61960]_ , \new_[61961]_ , \new_[61964]_ , \new_[61967]_ ,
    \new_[61968]_ , \new_[61969]_ , \new_[61972]_ , \new_[61975]_ ,
    \new_[61976]_ , \new_[61979]_ , \new_[61982]_ , \new_[61983]_ ,
    \new_[61984]_ , \new_[61988]_ , \new_[61989]_ , \new_[61992]_ ,
    \new_[61995]_ , \new_[61996]_ , \new_[61997]_ , \new_[62000]_ ,
    \new_[62003]_ , \new_[62004]_ , \new_[62007]_ , \new_[62010]_ ,
    \new_[62011]_ , \new_[62012]_ , \new_[62016]_ , \new_[62017]_ ,
    \new_[62020]_ , \new_[62023]_ , \new_[62024]_ , \new_[62025]_ ,
    \new_[62028]_ , \new_[62031]_ , \new_[62032]_ , \new_[62035]_ ,
    \new_[62038]_ , \new_[62039]_ , \new_[62040]_ , \new_[62044]_ ,
    \new_[62045]_ , \new_[62048]_ , \new_[62051]_ , \new_[62052]_ ,
    \new_[62053]_ , \new_[62056]_ , \new_[62059]_ , \new_[62060]_ ,
    \new_[62063]_ , \new_[62066]_ , \new_[62067]_ , \new_[62068]_ ,
    \new_[62072]_ , \new_[62073]_ , \new_[62076]_ , \new_[62079]_ ,
    \new_[62080]_ , \new_[62081]_ , \new_[62084]_ , \new_[62087]_ ,
    \new_[62088]_ , \new_[62091]_ , \new_[62094]_ , \new_[62095]_ ,
    \new_[62096]_ , \new_[62100]_ , \new_[62101]_ , \new_[62104]_ ,
    \new_[62107]_ , \new_[62108]_ , \new_[62109]_ , \new_[62112]_ ,
    \new_[62115]_ , \new_[62116]_ , \new_[62119]_ , \new_[62122]_ ,
    \new_[62123]_ , \new_[62124]_ , \new_[62128]_ , \new_[62129]_ ,
    \new_[62132]_ , \new_[62135]_ , \new_[62136]_ , \new_[62137]_ ,
    \new_[62140]_ , \new_[62143]_ , \new_[62144]_ , \new_[62147]_ ,
    \new_[62150]_ , \new_[62151]_ , \new_[62152]_ , \new_[62156]_ ,
    \new_[62157]_ , \new_[62160]_ , \new_[62163]_ , \new_[62164]_ ,
    \new_[62165]_ , \new_[62168]_ , \new_[62171]_ , \new_[62172]_ ,
    \new_[62175]_ , \new_[62178]_ , \new_[62179]_ , \new_[62180]_ ,
    \new_[62184]_ , \new_[62185]_ , \new_[62188]_ , \new_[62191]_ ,
    \new_[62192]_ , \new_[62193]_ , \new_[62196]_ , \new_[62199]_ ,
    \new_[62200]_ , \new_[62203]_ , \new_[62206]_ , \new_[62207]_ ,
    \new_[62208]_ , \new_[62212]_ , \new_[62213]_ , \new_[62216]_ ,
    \new_[62219]_ , \new_[62220]_ , \new_[62221]_ , \new_[62224]_ ,
    \new_[62227]_ , \new_[62228]_ , \new_[62231]_ , \new_[62234]_ ,
    \new_[62235]_ , \new_[62236]_ , \new_[62240]_ , \new_[62241]_ ,
    \new_[62244]_ , \new_[62247]_ , \new_[62248]_ , \new_[62249]_ ,
    \new_[62252]_ , \new_[62255]_ , \new_[62256]_ , \new_[62259]_ ,
    \new_[62262]_ , \new_[62263]_ , \new_[62264]_ , \new_[62268]_ ,
    \new_[62269]_ , \new_[62272]_ , \new_[62275]_ , \new_[62276]_ ,
    \new_[62277]_ , \new_[62280]_ , \new_[62283]_ , \new_[62284]_ ,
    \new_[62287]_ , \new_[62290]_ , \new_[62291]_ , \new_[62292]_ ,
    \new_[62296]_ , \new_[62297]_ , \new_[62300]_ , \new_[62303]_ ,
    \new_[62304]_ , \new_[62305]_ , \new_[62308]_ , \new_[62311]_ ,
    \new_[62312]_ , \new_[62315]_ , \new_[62318]_ , \new_[62319]_ ,
    \new_[62320]_ , \new_[62324]_ , \new_[62325]_ , \new_[62328]_ ,
    \new_[62331]_ , \new_[62332]_ , \new_[62333]_ , \new_[62336]_ ,
    \new_[62339]_ , \new_[62340]_ , \new_[62343]_ , \new_[62346]_ ,
    \new_[62347]_ , \new_[62348]_ , \new_[62352]_ , \new_[62353]_ ,
    \new_[62356]_ , \new_[62359]_ , \new_[62360]_ , \new_[62361]_ ,
    \new_[62364]_ , \new_[62367]_ , \new_[62368]_ , \new_[62371]_ ,
    \new_[62374]_ , \new_[62375]_ , \new_[62376]_ , \new_[62380]_ ,
    \new_[62381]_ , \new_[62384]_ , \new_[62387]_ , \new_[62388]_ ,
    \new_[62389]_ , \new_[62392]_ , \new_[62395]_ , \new_[62396]_ ,
    \new_[62399]_ , \new_[62402]_ , \new_[62403]_ , \new_[62404]_ ,
    \new_[62408]_ , \new_[62409]_ , \new_[62412]_ , \new_[62415]_ ,
    \new_[62416]_ , \new_[62417]_ , \new_[62420]_ , \new_[62423]_ ,
    \new_[62424]_ , \new_[62427]_ , \new_[62430]_ , \new_[62431]_ ,
    \new_[62432]_ , \new_[62436]_ , \new_[62437]_ , \new_[62440]_ ,
    \new_[62443]_ , \new_[62444]_ , \new_[62445]_ , \new_[62448]_ ,
    \new_[62451]_ , \new_[62452]_ , \new_[62455]_ , \new_[62458]_ ,
    \new_[62459]_ , \new_[62460]_ , \new_[62464]_ , \new_[62465]_ ,
    \new_[62468]_ , \new_[62471]_ , \new_[62472]_ , \new_[62473]_ ,
    \new_[62476]_ , \new_[62479]_ , \new_[62480]_ , \new_[62483]_ ,
    \new_[62486]_ , \new_[62487]_ , \new_[62488]_ , \new_[62492]_ ,
    \new_[62493]_ , \new_[62496]_ , \new_[62499]_ , \new_[62500]_ ,
    \new_[62501]_ , \new_[62504]_ , \new_[62507]_ , \new_[62508]_ ,
    \new_[62511]_ , \new_[62514]_ , \new_[62515]_ , \new_[62516]_ ,
    \new_[62520]_ , \new_[62521]_ , \new_[62524]_ , \new_[62527]_ ,
    \new_[62528]_ , \new_[62529]_ , \new_[62532]_ , \new_[62535]_ ,
    \new_[62536]_ , \new_[62539]_ , \new_[62542]_ , \new_[62543]_ ,
    \new_[62544]_ , \new_[62548]_ , \new_[62549]_ , \new_[62552]_ ,
    \new_[62555]_ , \new_[62556]_ , \new_[62557]_ , \new_[62560]_ ,
    \new_[62563]_ , \new_[62564]_ , \new_[62567]_ , \new_[62570]_ ,
    \new_[62571]_ , \new_[62572]_ , \new_[62576]_ , \new_[62577]_ ,
    \new_[62580]_ , \new_[62583]_ , \new_[62584]_ , \new_[62585]_ ,
    \new_[62588]_ , \new_[62591]_ , \new_[62592]_ , \new_[62595]_ ,
    \new_[62598]_ , \new_[62599]_ , \new_[62600]_ , \new_[62604]_ ,
    \new_[62605]_ , \new_[62608]_ , \new_[62611]_ , \new_[62612]_ ,
    \new_[62613]_ , \new_[62616]_ , \new_[62619]_ , \new_[62620]_ ,
    \new_[62623]_ , \new_[62626]_ , \new_[62627]_ , \new_[62628]_ ,
    \new_[62632]_ , \new_[62633]_ , \new_[62636]_ , \new_[62639]_ ,
    \new_[62640]_ , \new_[62641]_ , \new_[62644]_ , \new_[62647]_ ,
    \new_[62648]_ , \new_[62651]_ , \new_[62654]_ , \new_[62655]_ ,
    \new_[62656]_ , \new_[62660]_ , \new_[62661]_ , \new_[62664]_ ,
    \new_[62667]_ , \new_[62668]_ , \new_[62669]_ , \new_[62672]_ ,
    \new_[62675]_ , \new_[62676]_ , \new_[62679]_ , \new_[62682]_ ,
    \new_[62683]_ , \new_[62684]_ , \new_[62688]_ , \new_[62689]_ ,
    \new_[62692]_ , \new_[62695]_ , \new_[62696]_ , \new_[62697]_ ,
    \new_[62700]_ , \new_[62703]_ , \new_[62704]_ , \new_[62707]_ ,
    \new_[62710]_ , \new_[62711]_ , \new_[62712]_ , \new_[62716]_ ,
    \new_[62717]_ , \new_[62720]_ , \new_[62723]_ , \new_[62724]_ ,
    \new_[62725]_ , \new_[62728]_ , \new_[62731]_ , \new_[62732]_ ,
    \new_[62735]_ , \new_[62738]_ , \new_[62739]_ , \new_[62740]_ ,
    \new_[62744]_ , \new_[62745]_ , \new_[62748]_ , \new_[62751]_ ,
    \new_[62752]_ , \new_[62753]_ , \new_[62756]_ , \new_[62759]_ ,
    \new_[62760]_ , \new_[62763]_ , \new_[62766]_ , \new_[62767]_ ,
    \new_[62768]_ , \new_[62772]_ , \new_[62773]_ , \new_[62776]_ ,
    \new_[62779]_ , \new_[62780]_ , \new_[62781]_ , \new_[62784]_ ,
    \new_[62787]_ , \new_[62788]_ , \new_[62791]_ , \new_[62794]_ ,
    \new_[62795]_ , \new_[62796]_ , \new_[62800]_ , \new_[62801]_ ,
    \new_[62804]_ , \new_[62807]_ , \new_[62808]_ , \new_[62809]_ ,
    \new_[62812]_ , \new_[62815]_ , \new_[62816]_ , \new_[62819]_ ,
    \new_[62822]_ , \new_[62823]_ , \new_[62824]_ , \new_[62828]_ ,
    \new_[62829]_ , \new_[62832]_ , \new_[62835]_ , \new_[62836]_ ,
    \new_[62837]_ , \new_[62840]_ , \new_[62843]_ , \new_[62844]_ ,
    \new_[62847]_ , \new_[62850]_ , \new_[62851]_ , \new_[62852]_ ,
    \new_[62856]_ , \new_[62857]_ , \new_[62860]_ , \new_[62863]_ ,
    \new_[62864]_ , \new_[62865]_ , \new_[62868]_ , \new_[62871]_ ,
    \new_[62872]_ , \new_[62875]_ , \new_[62878]_ , \new_[62879]_ ,
    \new_[62880]_ , \new_[62884]_ , \new_[62885]_ , \new_[62888]_ ,
    \new_[62891]_ , \new_[62892]_ , \new_[62893]_ , \new_[62896]_ ,
    \new_[62899]_ , \new_[62900]_ , \new_[62903]_ , \new_[62906]_ ,
    \new_[62907]_ , \new_[62908]_ , \new_[62912]_ , \new_[62913]_ ,
    \new_[62916]_ , \new_[62919]_ , \new_[62920]_ , \new_[62921]_ ,
    \new_[62924]_ , \new_[62927]_ , \new_[62928]_ , \new_[62931]_ ,
    \new_[62934]_ , \new_[62935]_ , \new_[62936]_ , \new_[62940]_ ,
    \new_[62941]_ , \new_[62944]_ , \new_[62947]_ , \new_[62948]_ ,
    \new_[62949]_ , \new_[62952]_ , \new_[62955]_ , \new_[62956]_ ,
    \new_[62959]_ , \new_[62962]_ , \new_[62963]_ , \new_[62964]_ ,
    \new_[62968]_ , \new_[62969]_ , \new_[62972]_ , \new_[62975]_ ,
    \new_[62976]_ , \new_[62977]_ , \new_[62980]_ , \new_[62983]_ ,
    \new_[62984]_ , \new_[62987]_ , \new_[62990]_ , \new_[62991]_ ,
    \new_[62992]_ , \new_[62996]_ , \new_[62997]_ , \new_[63000]_ ,
    \new_[63003]_ , \new_[63004]_ , \new_[63005]_ , \new_[63008]_ ,
    \new_[63011]_ , \new_[63012]_ , \new_[63015]_ , \new_[63018]_ ,
    \new_[63019]_ , \new_[63020]_ , \new_[63024]_ , \new_[63025]_ ,
    \new_[63028]_ , \new_[63031]_ , \new_[63032]_ , \new_[63033]_ ,
    \new_[63036]_ , \new_[63039]_ , \new_[63040]_ , \new_[63043]_ ,
    \new_[63046]_ , \new_[63047]_ , \new_[63048]_ , \new_[63052]_ ,
    \new_[63053]_ , \new_[63056]_ , \new_[63059]_ , \new_[63060]_ ,
    \new_[63061]_ , \new_[63064]_ , \new_[63067]_ , \new_[63068]_ ,
    \new_[63071]_ , \new_[63074]_ , \new_[63075]_ , \new_[63076]_ ,
    \new_[63080]_ , \new_[63081]_ , \new_[63084]_ , \new_[63087]_ ,
    \new_[63088]_ , \new_[63089]_ , \new_[63092]_ , \new_[63095]_ ,
    \new_[63096]_ , \new_[63099]_ , \new_[63102]_ , \new_[63103]_ ,
    \new_[63104]_ , \new_[63108]_ , \new_[63109]_ , \new_[63112]_ ,
    \new_[63115]_ , \new_[63116]_ , \new_[63117]_ , \new_[63120]_ ,
    \new_[63123]_ , \new_[63124]_ , \new_[63127]_ , \new_[63130]_ ,
    \new_[63131]_ , \new_[63132]_ , \new_[63136]_ , \new_[63137]_ ,
    \new_[63140]_ , \new_[63143]_ , \new_[63144]_ , \new_[63145]_ ,
    \new_[63148]_ , \new_[63151]_ , \new_[63152]_ , \new_[63155]_ ,
    \new_[63158]_ , \new_[63159]_ , \new_[63160]_ , \new_[63164]_ ,
    \new_[63165]_ , \new_[63168]_ , \new_[63171]_ , \new_[63172]_ ,
    \new_[63173]_ , \new_[63176]_ , \new_[63179]_ , \new_[63180]_ ,
    \new_[63183]_ , \new_[63186]_ , \new_[63187]_ , \new_[63188]_ ,
    \new_[63192]_ , \new_[63193]_ , \new_[63196]_ , \new_[63199]_ ,
    \new_[63200]_ , \new_[63201]_ , \new_[63204]_ , \new_[63207]_ ,
    \new_[63208]_ , \new_[63211]_ , \new_[63214]_ , \new_[63215]_ ,
    \new_[63216]_ , \new_[63220]_ , \new_[63221]_ , \new_[63224]_ ,
    \new_[63227]_ , \new_[63228]_ , \new_[63229]_ , \new_[63232]_ ,
    \new_[63235]_ , \new_[63236]_ , \new_[63239]_ , \new_[63242]_ ,
    \new_[63243]_ , \new_[63244]_ , \new_[63248]_ , \new_[63249]_ ,
    \new_[63252]_ , \new_[63255]_ , \new_[63256]_ , \new_[63257]_ ,
    \new_[63260]_ , \new_[63263]_ , \new_[63264]_ , \new_[63267]_ ,
    \new_[63270]_ , \new_[63271]_ , \new_[63272]_ , \new_[63276]_ ,
    \new_[63277]_ , \new_[63280]_ , \new_[63283]_ , \new_[63284]_ ,
    \new_[63285]_ , \new_[63288]_ , \new_[63291]_ , \new_[63292]_ ,
    \new_[63295]_ , \new_[63298]_ , \new_[63299]_ , \new_[63300]_ ,
    \new_[63304]_ , \new_[63305]_ , \new_[63308]_ , \new_[63311]_ ,
    \new_[63312]_ , \new_[63313]_ , \new_[63316]_ , \new_[63319]_ ,
    \new_[63320]_ , \new_[63323]_ , \new_[63326]_ , \new_[63327]_ ,
    \new_[63328]_ , \new_[63332]_ , \new_[63333]_ , \new_[63336]_ ,
    \new_[63339]_ , \new_[63340]_ , \new_[63341]_ , \new_[63344]_ ,
    \new_[63347]_ , \new_[63348]_ , \new_[63351]_ , \new_[63354]_ ,
    \new_[63355]_ , \new_[63356]_ , \new_[63360]_ , \new_[63361]_ ,
    \new_[63364]_ , \new_[63367]_ , \new_[63368]_ , \new_[63369]_ ,
    \new_[63372]_ , \new_[63375]_ , \new_[63376]_ , \new_[63379]_ ,
    \new_[63382]_ , \new_[63383]_ , \new_[63384]_ , \new_[63388]_ ,
    \new_[63389]_ , \new_[63392]_ , \new_[63395]_ , \new_[63396]_ ,
    \new_[63397]_ , \new_[63400]_ , \new_[63403]_ , \new_[63404]_ ,
    \new_[63407]_ , \new_[63410]_ , \new_[63411]_ , \new_[63412]_ ,
    \new_[63416]_ , \new_[63417]_ , \new_[63420]_ , \new_[63423]_ ,
    \new_[63424]_ , \new_[63425]_ , \new_[63428]_ , \new_[63431]_ ,
    \new_[63432]_ , \new_[63435]_ , \new_[63438]_ , \new_[63439]_ ,
    \new_[63440]_ , \new_[63444]_ , \new_[63445]_ , \new_[63448]_ ,
    \new_[63451]_ , \new_[63452]_ , \new_[63453]_ , \new_[63456]_ ,
    \new_[63459]_ , \new_[63460]_ , \new_[63463]_ , \new_[63466]_ ,
    \new_[63467]_ , \new_[63468]_ , \new_[63472]_ , \new_[63473]_ ,
    \new_[63476]_ , \new_[63479]_ , \new_[63480]_ , \new_[63481]_ ,
    \new_[63484]_ , \new_[63487]_ , \new_[63488]_ , \new_[63491]_ ,
    \new_[63494]_ , \new_[63495]_ , \new_[63496]_ , \new_[63500]_ ,
    \new_[63501]_ , \new_[63504]_ , \new_[63507]_ , \new_[63508]_ ,
    \new_[63509]_ , \new_[63512]_ , \new_[63515]_ , \new_[63516]_ ,
    \new_[63519]_ , \new_[63522]_ , \new_[63523]_ , \new_[63524]_ ,
    \new_[63528]_ , \new_[63529]_ , \new_[63532]_ , \new_[63535]_ ,
    \new_[63536]_ , \new_[63537]_ , \new_[63540]_ , \new_[63543]_ ,
    \new_[63544]_ , \new_[63547]_ , \new_[63550]_ , \new_[63551]_ ,
    \new_[63552]_ , \new_[63556]_ , \new_[63557]_ , \new_[63560]_ ,
    \new_[63563]_ , \new_[63564]_ , \new_[63565]_ , \new_[63568]_ ,
    \new_[63571]_ , \new_[63572]_ , \new_[63575]_ , \new_[63578]_ ,
    \new_[63579]_ , \new_[63580]_ , \new_[63584]_ , \new_[63585]_ ,
    \new_[63588]_ , \new_[63591]_ , \new_[63592]_ , \new_[63593]_ ,
    \new_[63596]_ , \new_[63599]_ , \new_[63600]_ , \new_[63603]_ ,
    \new_[63606]_ , \new_[63607]_ , \new_[63608]_ , \new_[63612]_ ,
    \new_[63613]_ , \new_[63616]_ , \new_[63619]_ , \new_[63620]_ ,
    \new_[63621]_ , \new_[63624]_ , \new_[63627]_ , \new_[63628]_ ,
    \new_[63631]_ , \new_[63634]_ , \new_[63635]_ , \new_[63636]_ ,
    \new_[63640]_ , \new_[63641]_ , \new_[63644]_ , \new_[63647]_ ,
    \new_[63648]_ , \new_[63649]_ , \new_[63652]_ , \new_[63655]_ ,
    \new_[63656]_ , \new_[63659]_ , \new_[63662]_ , \new_[63663]_ ,
    \new_[63664]_ , \new_[63668]_ , \new_[63669]_ , \new_[63672]_ ,
    \new_[63675]_ , \new_[63676]_ , \new_[63677]_ , \new_[63680]_ ,
    \new_[63683]_ , \new_[63684]_ , \new_[63687]_ , \new_[63690]_ ,
    \new_[63691]_ , \new_[63692]_ , \new_[63696]_ , \new_[63697]_ ,
    \new_[63700]_ , \new_[63703]_ , \new_[63704]_ , \new_[63705]_ ,
    \new_[63708]_ , \new_[63711]_ , \new_[63712]_ , \new_[63715]_ ,
    \new_[63718]_ , \new_[63719]_ , \new_[63720]_ , \new_[63724]_ ,
    \new_[63725]_ , \new_[63728]_ , \new_[63731]_ , \new_[63732]_ ,
    \new_[63733]_ , \new_[63736]_ , \new_[63739]_ , \new_[63740]_ ,
    \new_[63743]_ , \new_[63746]_ , \new_[63747]_ , \new_[63748]_ ,
    \new_[63752]_ , \new_[63753]_ , \new_[63756]_ , \new_[63759]_ ,
    \new_[63760]_ , \new_[63761]_ , \new_[63764]_ , \new_[63767]_ ,
    \new_[63768]_ , \new_[63771]_ , \new_[63774]_ , \new_[63775]_ ,
    \new_[63776]_ , \new_[63780]_ , \new_[63781]_ , \new_[63784]_ ,
    \new_[63787]_ , \new_[63788]_ , \new_[63789]_ , \new_[63792]_ ,
    \new_[63795]_ , \new_[63796]_ , \new_[63799]_ , \new_[63802]_ ,
    \new_[63803]_ , \new_[63804]_ , \new_[63808]_ , \new_[63809]_ ,
    \new_[63812]_ , \new_[63815]_ , \new_[63816]_ , \new_[63817]_ ,
    \new_[63820]_ , \new_[63823]_ , \new_[63824]_ , \new_[63827]_ ,
    \new_[63830]_ , \new_[63831]_ , \new_[63832]_ , \new_[63836]_ ,
    \new_[63837]_ , \new_[63840]_ , \new_[63843]_ , \new_[63844]_ ,
    \new_[63845]_ , \new_[63848]_ , \new_[63851]_ , \new_[63852]_ ,
    \new_[63855]_ , \new_[63858]_ , \new_[63859]_ , \new_[63860]_ ,
    \new_[63864]_ , \new_[63865]_ , \new_[63868]_ , \new_[63871]_ ,
    \new_[63872]_ , \new_[63873]_ , \new_[63876]_ , \new_[63879]_ ,
    \new_[63880]_ , \new_[63883]_ , \new_[63886]_ , \new_[63887]_ ,
    \new_[63888]_ , \new_[63892]_ , \new_[63893]_ , \new_[63896]_ ,
    \new_[63899]_ , \new_[63900]_ , \new_[63901]_ , \new_[63904]_ ,
    \new_[63907]_ , \new_[63908]_ , \new_[63911]_ , \new_[63914]_ ,
    \new_[63915]_ , \new_[63916]_ , \new_[63920]_ , \new_[63921]_ ,
    \new_[63924]_ , \new_[63927]_ , \new_[63928]_ , \new_[63929]_ ,
    \new_[63932]_ , \new_[63935]_ , \new_[63936]_ , \new_[63939]_ ,
    \new_[63942]_ , \new_[63943]_ , \new_[63944]_ , \new_[63948]_ ,
    \new_[63949]_ , \new_[63952]_ , \new_[63955]_ , \new_[63956]_ ,
    \new_[63957]_ , \new_[63960]_ , \new_[63963]_ , \new_[63964]_ ,
    \new_[63967]_ , \new_[63970]_ , \new_[63971]_ , \new_[63972]_ ,
    \new_[63976]_ , \new_[63977]_ , \new_[63980]_ , \new_[63983]_ ,
    \new_[63984]_ , \new_[63985]_ , \new_[63988]_ , \new_[63991]_ ,
    \new_[63992]_ , \new_[63995]_ , \new_[63998]_ , \new_[63999]_ ,
    \new_[64000]_ , \new_[64004]_ , \new_[64005]_ , \new_[64008]_ ,
    \new_[64011]_ , \new_[64012]_ , \new_[64013]_ , \new_[64016]_ ,
    \new_[64019]_ , \new_[64020]_ , \new_[64023]_ , \new_[64026]_ ,
    \new_[64027]_ , \new_[64028]_ , \new_[64032]_ , \new_[64033]_ ,
    \new_[64036]_ , \new_[64039]_ , \new_[64040]_ , \new_[64041]_ ,
    \new_[64044]_ , \new_[64047]_ , \new_[64048]_ , \new_[64051]_ ,
    \new_[64054]_ , \new_[64055]_ , \new_[64056]_ , \new_[64060]_ ,
    \new_[64061]_ , \new_[64064]_ , \new_[64067]_ , \new_[64068]_ ,
    \new_[64069]_ , \new_[64072]_ , \new_[64075]_ , \new_[64076]_ ,
    \new_[64079]_ , \new_[64082]_ , \new_[64083]_ , \new_[64084]_ ,
    \new_[64088]_ , \new_[64089]_ , \new_[64092]_ , \new_[64095]_ ,
    \new_[64096]_ , \new_[64097]_ , \new_[64100]_ , \new_[64103]_ ,
    \new_[64104]_ , \new_[64107]_ , \new_[64110]_ , \new_[64111]_ ,
    \new_[64112]_ , \new_[64116]_ , \new_[64117]_ , \new_[64120]_ ,
    \new_[64123]_ , \new_[64124]_ , \new_[64125]_ , \new_[64128]_ ,
    \new_[64131]_ , \new_[64132]_ , \new_[64135]_ , \new_[64138]_ ,
    \new_[64139]_ , \new_[64140]_ , \new_[64144]_ , \new_[64145]_ ,
    \new_[64148]_ , \new_[64151]_ , \new_[64152]_ , \new_[64153]_ ,
    \new_[64156]_ , \new_[64159]_ , \new_[64160]_ , \new_[64163]_ ,
    \new_[64166]_ , \new_[64167]_ , \new_[64168]_ , \new_[64172]_ ,
    \new_[64173]_ , \new_[64176]_ , \new_[64179]_ , \new_[64180]_ ,
    \new_[64181]_ , \new_[64184]_ , \new_[64187]_ , \new_[64188]_ ,
    \new_[64191]_ , \new_[64194]_ , \new_[64195]_ , \new_[64196]_ ,
    \new_[64200]_ , \new_[64201]_ , \new_[64204]_ , \new_[64207]_ ,
    \new_[64208]_ , \new_[64209]_ , \new_[64212]_ , \new_[64215]_ ,
    \new_[64216]_ , \new_[64219]_ , \new_[64222]_ , \new_[64223]_ ,
    \new_[64224]_ , \new_[64228]_ , \new_[64229]_ , \new_[64232]_ ,
    \new_[64235]_ , \new_[64236]_ , \new_[64237]_ , \new_[64240]_ ,
    \new_[64243]_ , \new_[64244]_ , \new_[64247]_ , \new_[64250]_ ,
    \new_[64251]_ , \new_[64252]_ , \new_[64256]_ , \new_[64257]_ ,
    \new_[64260]_ , \new_[64263]_ , \new_[64264]_ , \new_[64265]_ ,
    \new_[64268]_ , \new_[64271]_ , \new_[64272]_ , \new_[64275]_ ,
    \new_[64278]_ , \new_[64279]_ , \new_[64280]_ , \new_[64284]_ ,
    \new_[64285]_ , \new_[64288]_ , \new_[64291]_ , \new_[64292]_ ,
    \new_[64293]_ , \new_[64296]_ , \new_[64299]_ , \new_[64300]_ ,
    \new_[64303]_ , \new_[64306]_ , \new_[64307]_ , \new_[64308]_ ,
    \new_[64312]_ , \new_[64313]_ , \new_[64316]_ , \new_[64319]_ ,
    \new_[64320]_ , \new_[64321]_ , \new_[64324]_ , \new_[64327]_ ,
    \new_[64328]_ , \new_[64331]_ , \new_[64334]_ , \new_[64335]_ ,
    \new_[64336]_ , \new_[64340]_ , \new_[64341]_ , \new_[64344]_ ,
    \new_[64347]_ , \new_[64348]_ , \new_[64349]_ , \new_[64352]_ ,
    \new_[64355]_ , \new_[64356]_ , \new_[64359]_ , \new_[64362]_ ,
    \new_[64363]_ , \new_[64364]_ , \new_[64368]_ , \new_[64369]_ ,
    \new_[64372]_ , \new_[64375]_ , \new_[64376]_ , \new_[64377]_ ,
    \new_[64380]_ , \new_[64383]_ , \new_[64384]_ , \new_[64387]_ ,
    \new_[64390]_ , \new_[64391]_ , \new_[64392]_ , \new_[64396]_ ,
    \new_[64397]_ , \new_[64400]_ , \new_[64403]_ , \new_[64404]_ ,
    \new_[64405]_ , \new_[64408]_ , \new_[64411]_ , \new_[64412]_ ,
    \new_[64415]_ , \new_[64418]_ , \new_[64419]_ , \new_[64420]_ ,
    \new_[64424]_ , \new_[64425]_ , \new_[64428]_ , \new_[64431]_ ,
    \new_[64432]_ , \new_[64433]_ , \new_[64436]_ , \new_[64439]_ ,
    \new_[64440]_ , \new_[64443]_ , \new_[64446]_ , \new_[64447]_ ,
    \new_[64448]_ , \new_[64452]_ , \new_[64453]_ , \new_[64456]_ ,
    \new_[64459]_ , \new_[64460]_ , \new_[64461]_ , \new_[64464]_ ,
    \new_[64467]_ , \new_[64468]_ , \new_[64471]_ , \new_[64474]_ ,
    \new_[64475]_ , \new_[64476]_ , \new_[64480]_ , \new_[64481]_ ,
    \new_[64484]_ , \new_[64487]_ , \new_[64488]_ , \new_[64489]_ ,
    \new_[64492]_ , \new_[64495]_ , \new_[64496]_ , \new_[64499]_ ,
    \new_[64502]_ , \new_[64503]_ , \new_[64504]_ , \new_[64508]_ ,
    \new_[64509]_ , \new_[64512]_ , \new_[64515]_ , \new_[64516]_ ,
    \new_[64517]_ , \new_[64520]_ , \new_[64523]_ , \new_[64524]_ ,
    \new_[64527]_ , \new_[64530]_ , \new_[64531]_ , \new_[64532]_ ,
    \new_[64536]_ , \new_[64537]_ , \new_[64540]_ , \new_[64543]_ ,
    \new_[64544]_ , \new_[64545]_ , \new_[64548]_ , \new_[64551]_ ,
    \new_[64552]_ , \new_[64555]_ , \new_[64558]_ , \new_[64559]_ ,
    \new_[64560]_ , \new_[64564]_ , \new_[64565]_ , \new_[64568]_ ,
    \new_[64571]_ , \new_[64572]_ , \new_[64573]_ , \new_[64576]_ ,
    \new_[64579]_ , \new_[64580]_ , \new_[64583]_ , \new_[64586]_ ,
    \new_[64587]_ , \new_[64588]_ , \new_[64592]_ , \new_[64593]_ ,
    \new_[64596]_ , \new_[64599]_ , \new_[64600]_ , \new_[64601]_ ,
    \new_[64604]_ , \new_[64607]_ , \new_[64608]_ , \new_[64611]_ ,
    \new_[64614]_ , \new_[64615]_ , \new_[64616]_ , \new_[64620]_ ,
    \new_[64621]_ , \new_[64624]_ , \new_[64627]_ , \new_[64628]_ ,
    \new_[64629]_ , \new_[64632]_ , \new_[64635]_ , \new_[64636]_ ,
    \new_[64639]_ , \new_[64642]_ , \new_[64643]_ , \new_[64644]_ ,
    \new_[64648]_ , \new_[64649]_ , \new_[64652]_ , \new_[64655]_ ,
    \new_[64656]_ , \new_[64657]_ , \new_[64660]_ , \new_[64663]_ ,
    \new_[64664]_ , \new_[64667]_ , \new_[64670]_ , \new_[64671]_ ,
    \new_[64672]_ , \new_[64676]_ , \new_[64677]_ , \new_[64680]_ ,
    \new_[64683]_ , \new_[64684]_ , \new_[64685]_ , \new_[64688]_ ,
    \new_[64691]_ , \new_[64692]_ , \new_[64695]_ , \new_[64698]_ ,
    \new_[64699]_ , \new_[64700]_ , \new_[64704]_ , \new_[64705]_ ,
    \new_[64708]_ , \new_[64711]_ , \new_[64712]_ , \new_[64713]_ ,
    \new_[64716]_ , \new_[64719]_ , \new_[64720]_ , \new_[64723]_ ,
    \new_[64726]_ , \new_[64727]_ , \new_[64728]_ , \new_[64732]_ ,
    \new_[64733]_ , \new_[64736]_ , \new_[64739]_ , \new_[64740]_ ,
    \new_[64741]_ , \new_[64744]_ , \new_[64747]_ , \new_[64748]_ ,
    \new_[64751]_ , \new_[64754]_ , \new_[64755]_ , \new_[64756]_ ,
    \new_[64760]_ , \new_[64761]_ , \new_[64764]_ , \new_[64767]_ ,
    \new_[64768]_ , \new_[64769]_ , \new_[64772]_ , \new_[64775]_ ,
    \new_[64776]_ , \new_[64779]_ , \new_[64782]_ , \new_[64783]_ ,
    \new_[64784]_ , \new_[64788]_ , \new_[64789]_ , \new_[64792]_ ,
    \new_[64795]_ , \new_[64796]_ , \new_[64797]_ , \new_[64800]_ ,
    \new_[64803]_ , \new_[64804]_ , \new_[64807]_ , \new_[64810]_ ,
    \new_[64811]_ , \new_[64812]_ , \new_[64816]_ , \new_[64817]_ ,
    \new_[64820]_ , \new_[64823]_ , \new_[64824]_ , \new_[64825]_ ,
    \new_[64828]_ , \new_[64831]_ , \new_[64832]_ , \new_[64835]_ ,
    \new_[64838]_ , \new_[64839]_ , \new_[64840]_ , \new_[64844]_ ,
    \new_[64845]_ , \new_[64848]_ , \new_[64851]_ , \new_[64852]_ ,
    \new_[64853]_ , \new_[64856]_ , \new_[64859]_ , \new_[64860]_ ,
    \new_[64863]_ , \new_[64866]_ , \new_[64867]_ , \new_[64868]_ ,
    \new_[64872]_ , \new_[64873]_ , \new_[64876]_ , \new_[64879]_ ,
    \new_[64880]_ , \new_[64881]_ , \new_[64884]_ , \new_[64887]_ ,
    \new_[64888]_ , \new_[64891]_ , \new_[64894]_ , \new_[64895]_ ,
    \new_[64896]_ , \new_[64900]_ , \new_[64901]_ , \new_[64904]_ ,
    \new_[64907]_ , \new_[64908]_ , \new_[64909]_ , \new_[64912]_ ,
    \new_[64915]_ , \new_[64916]_ , \new_[64919]_ , \new_[64922]_ ,
    \new_[64923]_ , \new_[64924]_ , \new_[64928]_ , \new_[64929]_ ,
    \new_[64932]_ , \new_[64935]_ , \new_[64936]_ , \new_[64937]_ ,
    \new_[64940]_ , \new_[64943]_ , \new_[64944]_ , \new_[64947]_ ,
    \new_[64950]_ , \new_[64951]_ , \new_[64952]_ , \new_[64956]_ ,
    \new_[64957]_ , \new_[64960]_ , \new_[64963]_ , \new_[64964]_ ,
    \new_[64965]_ , \new_[64968]_ , \new_[64971]_ , \new_[64972]_ ,
    \new_[64975]_ , \new_[64978]_ , \new_[64979]_ , \new_[64980]_ ,
    \new_[64984]_ , \new_[64985]_ , \new_[64988]_ , \new_[64991]_ ,
    \new_[64992]_ , \new_[64993]_ , \new_[64996]_ , \new_[64999]_ ,
    \new_[65000]_ , \new_[65003]_ , \new_[65006]_ , \new_[65007]_ ,
    \new_[65008]_ , \new_[65012]_ , \new_[65013]_ , \new_[65016]_ ,
    \new_[65019]_ , \new_[65020]_ , \new_[65021]_ , \new_[65024]_ ,
    \new_[65027]_ , \new_[65028]_ , \new_[65031]_ , \new_[65034]_ ,
    \new_[65035]_ , \new_[65036]_ , \new_[65040]_ , \new_[65041]_ ,
    \new_[65044]_ , \new_[65047]_ , \new_[65048]_ , \new_[65049]_ ,
    \new_[65052]_ , \new_[65055]_ , \new_[65056]_ , \new_[65059]_ ,
    \new_[65062]_ , \new_[65063]_ , \new_[65064]_ , \new_[65068]_ ,
    \new_[65069]_ , \new_[65072]_ , \new_[65075]_ , \new_[65076]_ ,
    \new_[65077]_ , \new_[65080]_ , \new_[65083]_ , \new_[65084]_ ,
    \new_[65087]_ , \new_[65090]_ , \new_[65091]_ , \new_[65092]_ ,
    \new_[65096]_ , \new_[65097]_ , \new_[65100]_ , \new_[65103]_ ,
    \new_[65104]_ , \new_[65105]_ , \new_[65108]_ , \new_[65111]_ ,
    \new_[65112]_ , \new_[65115]_ , \new_[65118]_ , \new_[65119]_ ,
    \new_[65120]_ , \new_[65124]_ , \new_[65125]_ , \new_[65128]_ ,
    \new_[65131]_ , \new_[65132]_ , \new_[65133]_ , \new_[65136]_ ,
    \new_[65139]_ , \new_[65140]_ , \new_[65143]_ , \new_[65146]_ ,
    \new_[65147]_ , \new_[65148]_ , \new_[65152]_ , \new_[65153]_ ,
    \new_[65156]_ , \new_[65159]_ , \new_[65160]_ , \new_[65161]_ ,
    \new_[65164]_ , \new_[65167]_ , \new_[65168]_ , \new_[65171]_ ,
    \new_[65174]_ , \new_[65175]_ , \new_[65176]_ , \new_[65180]_ ,
    \new_[65181]_ , \new_[65184]_ , \new_[65187]_ , \new_[65188]_ ,
    \new_[65189]_ , \new_[65192]_ , \new_[65195]_ , \new_[65196]_ ,
    \new_[65199]_ , \new_[65202]_ , \new_[65203]_ , \new_[65204]_ ,
    \new_[65208]_ , \new_[65209]_ , \new_[65212]_ , \new_[65215]_ ,
    \new_[65216]_ , \new_[65217]_ , \new_[65220]_ , \new_[65223]_ ,
    \new_[65224]_ , \new_[65227]_ , \new_[65230]_ , \new_[65231]_ ,
    \new_[65232]_ , \new_[65236]_ , \new_[65237]_ , \new_[65240]_ ,
    \new_[65243]_ , \new_[65244]_ , \new_[65245]_ , \new_[65248]_ ,
    \new_[65251]_ , \new_[65252]_ , \new_[65255]_ , \new_[65258]_ ,
    \new_[65259]_ , \new_[65260]_ , \new_[65264]_ , \new_[65265]_ ,
    \new_[65268]_ , \new_[65271]_ , \new_[65272]_ , \new_[65273]_ ,
    \new_[65276]_ , \new_[65279]_ , \new_[65280]_ , \new_[65283]_ ,
    \new_[65286]_ , \new_[65287]_ , \new_[65288]_ , \new_[65292]_ ,
    \new_[65293]_ , \new_[65296]_ , \new_[65299]_ , \new_[65300]_ ,
    \new_[65301]_ , \new_[65304]_ , \new_[65307]_ , \new_[65308]_ ,
    \new_[65311]_ , \new_[65314]_ , \new_[65315]_ , \new_[65316]_ ,
    \new_[65320]_ , \new_[65321]_ , \new_[65324]_ , \new_[65327]_ ,
    \new_[65328]_ , \new_[65329]_ , \new_[65332]_ , \new_[65335]_ ,
    \new_[65336]_ , \new_[65339]_ , \new_[65342]_ , \new_[65343]_ ,
    \new_[65344]_ , \new_[65348]_ , \new_[65349]_ , \new_[65352]_ ,
    \new_[65355]_ , \new_[65356]_ , \new_[65357]_ , \new_[65360]_ ,
    \new_[65363]_ , \new_[65364]_ , \new_[65367]_ , \new_[65370]_ ,
    \new_[65371]_ , \new_[65372]_ , \new_[65376]_ , \new_[65377]_ ,
    \new_[65380]_ , \new_[65383]_ , \new_[65384]_ , \new_[65385]_ ,
    \new_[65388]_ , \new_[65391]_ , \new_[65392]_ , \new_[65395]_ ,
    \new_[65398]_ , \new_[65399]_ , \new_[65400]_ , \new_[65404]_ ,
    \new_[65405]_ , \new_[65408]_ , \new_[65411]_ , \new_[65412]_ ,
    \new_[65413]_ , \new_[65416]_ , \new_[65419]_ , \new_[65420]_ ,
    \new_[65423]_ , \new_[65426]_ , \new_[65427]_ , \new_[65428]_ ,
    \new_[65432]_ , \new_[65433]_ , \new_[65436]_ , \new_[65439]_ ,
    \new_[65440]_ , \new_[65441]_ , \new_[65444]_ , \new_[65447]_ ,
    \new_[65448]_ , \new_[65451]_ , \new_[65454]_ , \new_[65455]_ ,
    \new_[65456]_ , \new_[65460]_ , \new_[65461]_ , \new_[65464]_ ,
    \new_[65467]_ , \new_[65468]_ , \new_[65469]_ , \new_[65472]_ ,
    \new_[65475]_ , \new_[65476]_ , \new_[65479]_ , \new_[65482]_ ,
    \new_[65483]_ , \new_[65484]_ , \new_[65488]_ , \new_[65489]_ ,
    \new_[65492]_ , \new_[65495]_ , \new_[65496]_ , \new_[65497]_ ,
    \new_[65500]_ , \new_[65503]_ , \new_[65504]_ , \new_[65507]_ ,
    \new_[65510]_ , \new_[65511]_ , \new_[65512]_ , \new_[65516]_ ,
    \new_[65517]_ , \new_[65520]_ , \new_[65523]_ , \new_[65524]_ ,
    \new_[65525]_ , \new_[65528]_ , \new_[65531]_ , \new_[65532]_ ,
    \new_[65535]_ , \new_[65538]_ , \new_[65539]_ , \new_[65540]_ ,
    \new_[65544]_ , \new_[65545]_ , \new_[65548]_ , \new_[65551]_ ,
    \new_[65552]_ , \new_[65553]_ , \new_[65556]_ , \new_[65559]_ ,
    \new_[65560]_ , \new_[65563]_ , \new_[65566]_ , \new_[65567]_ ,
    \new_[65568]_ , \new_[65572]_ , \new_[65573]_ , \new_[65576]_ ,
    \new_[65579]_ , \new_[65580]_ , \new_[65581]_ , \new_[65584]_ ,
    \new_[65587]_ , \new_[65588]_ , \new_[65591]_ , \new_[65594]_ ,
    \new_[65595]_ , \new_[65596]_ , \new_[65600]_ , \new_[65601]_ ,
    \new_[65604]_ , \new_[65607]_ , \new_[65608]_ , \new_[65609]_ ,
    \new_[65612]_ , \new_[65615]_ , \new_[65616]_ , \new_[65619]_ ,
    \new_[65622]_ , \new_[65623]_ , \new_[65624]_ , \new_[65628]_ ,
    \new_[65629]_ , \new_[65632]_ , \new_[65635]_ , \new_[65636]_ ,
    \new_[65637]_ , \new_[65640]_ , \new_[65643]_ , \new_[65644]_ ,
    \new_[65647]_ , \new_[65650]_ , \new_[65651]_ , \new_[65652]_ ,
    \new_[65656]_ , \new_[65657]_ , \new_[65660]_ , \new_[65663]_ ,
    \new_[65664]_ , \new_[65665]_ , \new_[65668]_ , \new_[65671]_ ,
    \new_[65672]_ , \new_[65675]_ , \new_[65678]_ , \new_[65679]_ ,
    \new_[65680]_ , \new_[65684]_ , \new_[65685]_ , \new_[65688]_ ,
    \new_[65691]_ , \new_[65692]_ , \new_[65693]_ , \new_[65696]_ ,
    \new_[65699]_ , \new_[65700]_ , \new_[65703]_ , \new_[65706]_ ,
    \new_[65707]_ , \new_[65708]_ , \new_[65712]_ , \new_[65713]_ ,
    \new_[65716]_ , \new_[65719]_ , \new_[65720]_ , \new_[65721]_ ,
    \new_[65724]_ , \new_[65727]_ , \new_[65728]_ , \new_[65731]_ ,
    \new_[65734]_ , \new_[65735]_ , \new_[65736]_ , \new_[65740]_ ,
    \new_[65741]_ , \new_[65744]_ , \new_[65747]_ , \new_[65748]_ ,
    \new_[65749]_ , \new_[65752]_ , \new_[65755]_ , \new_[65756]_ ,
    \new_[65759]_ , \new_[65762]_ , \new_[65763]_ , \new_[65764]_ ,
    \new_[65768]_ , \new_[65769]_ , \new_[65772]_ , \new_[65775]_ ,
    \new_[65776]_ , \new_[65777]_ , \new_[65780]_ , \new_[65783]_ ,
    \new_[65784]_ , \new_[65787]_ , \new_[65790]_ , \new_[65791]_ ,
    \new_[65792]_ , \new_[65796]_ , \new_[65797]_ , \new_[65800]_ ,
    \new_[65803]_ , \new_[65804]_ , \new_[65805]_ , \new_[65808]_ ,
    \new_[65811]_ , \new_[65812]_ , \new_[65815]_ , \new_[65818]_ ,
    \new_[65819]_ , \new_[65820]_ , \new_[65824]_ , \new_[65825]_ ,
    \new_[65828]_ , \new_[65831]_ , \new_[65832]_ , \new_[65833]_ ,
    \new_[65836]_ , \new_[65839]_ , \new_[65840]_ , \new_[65843]_ ,
    \new_[65846]_ , \new_[65847]_ , \new_[65848]_ , \new_[65852]_ ,
    \new_[65853]_ , \new_[65856]_ , \new_[65859]_ , \new_[65860]_ ,
    \new_[65861]_ , \new_[65864]_ , \new_[65867]_ , \new_[65868]_ ,
    \new_[65871]_ , \new_[65874]_ , \new_[65875]_ , \new_[65876]_ ,
    \new_[65880]_ , \new_[65881]_ , \new_[65884]_ , \new_[65887]_ ,
    \new_[65888]_ , \new_[65889]_ , \new_[65892]_ , \new_[65895]_ ,
    \new_[65896]_ , \new_[65899]_ , \new_[65902]_ , \new_[65903]_ ,
    \new_[65904]_ , \new_[65908]_ , \new_[65909]_ , \new_[65912]_ ,
    \new_[65915]_ , \new_[65916]_ , \new_[65917]_ , \new_[65920]_ ,
    \new_[65923]_ , \new_[65924]_ , \new_[65927]_ , \new_[65930]_ ,
    \new_[65931]_ , \new_[65932]_ , \new_[65936]_ , \new_[65937]_ ,
    \new_[65940]_ , \new_[65943]_ , \new_[65944]_ , \new_[65945]_ ,
    \new_[65948]_ , \new_[65951]_ , \new_[65952]_ , \new_[65955]_ ,
    \new_[65958]_ , \new_[65959]_ , \new_[65960]_ , \new_[65964]_ ,
    \new_[65965]_ , \new_[65968]_ , \new_[65971]_ , \new_[65972]_ ,
    \new_[65973]_ , \new_[65976]_ , \new_[65979]_ , \new_[65980]_ ,
    \new_[65983]_ , \new_[65986]_ , \new_[65987]_ , \new_[65988]_ ,
    \new_[65992]_ , \new_[65993]_ , \new_[65996]_ , \new_[65999]_ ,
    \new_[66000]_ , \new_[66001]_ , \new_[66004]_ , \new_[66007]_ ,
    \new_[66008]_ , \new_[66011]_ , \new_[66014]_ , \new_[66015]_ ,
    \new_[66016]_ , \new_[66020]_ , \new_[66021]_ , \new_[66024]_ ,
    \new_[66027]_ , \new_[66028]_ , \new_[66029]_ , \new_[66032]_ ,
    \new_[66035]_ , \new_[66036]_ , \new_[66039]_ , \new_[66042]_ ,
    \new_[66043]_ , \new_[66044]_ , \new_[66048]_ , \new_[66049]_ ,
    \new_[66052]_ , \new_[66055]_ , \new_[66056]_ , \new_[66057]_ ,
    \new_[66060]_ , \new_[66063]_ , \new_[66064]_ , \new_[66067]_ ,
    \new_[66070]_ , \new_[66071]_ , \new_[66072]_ , \new_[66076]_ ,
    \new_[66077]_ , \new_[66080]_ , \new_[66083]_ , \new_[66084]_ ,
    \new_[66085]_ , \new_[66088]_ , \new_[66091]_ , \new_[66092]_ ,
    \new_[66095]_ , \new_[66098]_ , \new_[66099]_ , \new_[66100]_ ,
    \new_[66104]_ , \new_[66105]_ , \new_[66108]_ , \new_[66111]_ ,
    \new_[66112]_ , \new_[66113]_ , \new_[66116]_ , \new_[66119]_ ,
    \new_[66120]_ , \new_[66123]_ , \new_[66126]_ , \new_[66127]_ ,
    \new_[66128]_ , \new_[66132]_ , \new_[66133]_ , \new_[66136]_ ,
    \new_[66139]_ , \new_[66140]_ , \new_[66141]_ , \new_[66144]_ ,
    \new_[66147]_ , \new_[66148]_ , \new_[66151]_ , \new_[66154]_ ,
    \new_[66155]_ , \new_[66156]_ , \new_[66160]_ , \new_[66161]_ ,
    \new_[66164]_ , \new_[66167]_ , \new_[66168]_ , \new_[66169]_ ,
    \new_[66172]_ , \new_[66175]_ , \new_[66176]_ , \new_[66179]_ ,
    \new_[66182]_ , \new_[66183]_ , \new_[66184]_ , \new_[66188]_ ,
    \new_[66189]_ , \new_[66192]_ , \new_[66195]_ , \new_[66196]_ ,
    \new_[66197]_ , \new_[66200]_ , \new_[66203]_ , \new_[66204]_ ,
    \new_[66207]_ , \new_[66210]_ , \new_[66211]_ , \new_[66212]_ ,
    \new_[66216]_ , \new_[66217]_ , \new_[66220]_ , \new_[66223]_ ,
    \new_[66224]_ , \new_[66225]_ , \new_[66228]_ , \new_[66231]_ ,
    \new_[66232]_ , \new_[66235]_ , \new_[66238]_ , \new_[66239]_ ,
    \new_[66240]_ , \new_[66244]_ , \new_[66245]_ , \new_[66248]_ ,
    \new_[66251]_ , \new_[66252]_ , \new_[66253]_ , \new_[66256]_ ,
    \new_[66259]_ , \new_[66260]_ , \new_[66263]_ , \new_[66266]_ ,
    \new_[66267]_ , \new_[66268]_ , \new_[66272]_ , \new_[66273]_ ,
    \new_[66276]_ , \new_[66279]_ , \new_[66280]_ , \new_[66281]_ ,
    \new_[66284]_ , \new_[66287]_ , \new_[66288]_ , \new_[66291]_ ,
    \new_[66294]_ , \new_[66295]_ , \new_[66296]_ , \new_[66300]_ ,
    \new_[66301]_ , \new_[66304]_ , \new_[66307]_ , \new_[66308]_ ,
    \new_[66309]_ , \new_[66312]_ , \new_[66315]_ , \new_[66316]_ ,
    \new_[66319]_ , \new_[66322]_ , \new_[66323]_ , \new_[66324]_ ,
    \new_[66328]_ , \new_[66329]_ , \new_[66332]_ , \new_[66335]_ ,
    \new_[66336]_ , \new_[66337]_ , \new_[66340]_ , \new_[66343]_ ,
    \new_[66344]_ , \new_[66347]_ , \new_[66350]_ , \new_[66351]_ ,
    \new_[66352]_ , \new_[66356]_ , \new_[66357]_ , \new_[66360]_ ,
    \new_[66363]_ , \new_[66364]_ , \new_[66365]_ , \new_[66368]_ ,
    \new_[66371]_ , \new_[66372]_ , \new_[66375]_ , \new_[66378]_ ,
    \new_[66379]_ , \new_[66380]_ , \new_[66384]_ , \new_[66385]_ ,
    \new_[66388]_ , \new_[66391]_ , \new_[66392]_ , \new_[66393]_ ,
    \new_[66396]_ , \new_[66399]_ , \new_[66400]_ , \new_[66403]_ ,
    \new_[66406]_ , \new_[66407]_ , \new_[66408]_ , \new_[66412]_ ,
    \new_[66413]_ , \new_[66416]_ , \new_[66419]_ , \new_[66420]_ ,
    \new_[66421]_ , \new_[66424]_ , \new_[66427]_ , \new_[66428]_ ,
    \new_[66431]_ , \new_[66434]_ , \new_[66435]_ , \new_[66436]_ ,
    \new_[66440]_ , \new_[66441]_ , \new_[66444]_ , \new_[66447]_ ,
    \new_[66448]_ , \new_[66449]_ , \new_[66452]_ , \new_[66455]_ ,
    \new_[66456]_ , \new_[66459]_ , \new_[66462]_ , \new_[66463]_ ,
    \new_[66464]_ , \new_[66468]_ , \new_[66469]_ , \new_[66472]_ ,
    \new_[66475]_ , \new_[66476]_ , \new_[66477]_ , \new_[66480]_ ,
    \new_[66483]_ , \new_[66484]_ , \new_[66487]_ , \new_[66490]_ ,
    \new_[66491]_ , \new_[66492]_ , \new_[66496]_ , \new_[66497]_ ,
    \new_[66500]_ , \new_[66503]_ , \new_[66504]_ , \new_[66505]_ ,
    \new_[66508]_ , \new_[66511]_ , \new_[66512]_ , \new_[66515]_ ,
    \new_[66518]_ , \new_[66519]_ , \new_[66520]_ , \new_[66524]_ ,
    \new_[66525]_ , \new_[66528]_ , \new_[66531]_ , \new_[66532]_ ,
    \new_[66533]_ , \new_[66536]_ , \new_[66539]_ , \new_[66540]_ ,
    \new_[66543]_ , \new_[66546]_ , \new_[66547]_ , \new_[66548]_ ,
    \new_[66552]_ , \new_[66553]_ , \new_[66556]_ , \new_[66559]_ ,
    \new_[66560]_ , \new_[66561]_ , \new_[66564]_ , \new_[66567]_ ,
    \new_[66568]_ , \new_[66571]_ , \new_[66574]_ , \new_[66575]_ ,
    \new_[66576]_ , \new_[66580]_ , \new_[66581]_ , \new_[66584]_ ,
    \new_[66587]_ , \new_[66588]_ , \new_[66589]_ , \new_[66592]_ ,
    \new_[66595]_ , \new_[66596]_ , \new_[66599]_ , \new_[66602]_ ,
    \new_[66603]_ , \new_[66604]_ , \new_[66608]_ , \new_[66609]_ ,
    \new_[66612]_ , \new_[66615]_ , \new_[66616]_ , \new_[66617]_ ,
    \new_[66620]_ , \new_[66623]_ , \new_[66624]_ , \new_[66627]_ ,
    \new_[66630]_ , \new_[66631]_ , \new_[66632]_ , \new_[66636]_ ,
    \new_[66637]_ , \new_[66640]_ , \new_[66643]_ , \new_[66644]_ ,
    \new_[66645]_ , \new_[66648]_ , \new_[66651]_ , \new_[66652]_ ,
    \new_[66655]_ , \new_[66658]_ , \new_[66659]_ , \new_[66660]_ ,
    \new_[66664]_ , \new_[66665]_ , \new_[66668]_ , \new_[66671]_ ,
    \new_[66672]_ , \new_[66673]_ , \new_[66676]_ , \new_[66679]_ ,
    \new_[66680]_ , \new_[66683]_ , \new_[66686]_ , \new_[66687]_ ,
    \new_[66688]_ , \new_[66692]_ , \new_[66693]_ , \new_[66696]_ ,
    \new_[66699]_ , \new_[66700]_ , \new_[66701]_ , \new_[66704]_ ,
    \new_[66707]_ , \new_[66708]_ , \new_[66711]_ , \new_[66714]_ ,
    \new_[66715]_ , \new_[66716]_ , \new_[66720]_ , \new_[66721]_ ,
    \new_[66724]_ , \new_[66727]_ , \new_[66728]_ , \new_[66729]_ ,
    \new_[66732]_ , \new_[66735]_ , \new_[66736]_ , \new_[66739]_ ,
    \new_[66742]_ , \new_[66743]_ , \new_[66744]_ , \new_[66748]_ ,
    \new_[66749]_ , \new_[66752]_ , \new_[66755]_ , \new_[66756]_ ,
    \new_[66757]_ , \new_[66760]_ , \new_[66763]_ , \new_[66764]_ ,
    \new_[66767]_ , \new_[66770]_ , \new_[66771]_ , \new_[66772]_ ,
    \new_[66776]_ , \new_[66777]_ , \new_[66780]_ , \new_[66783]_ ,
    \new_[66784]_ , \new_[66785]_ , \new_[66788]_ , \new_[66791]_ ,
    \new_[66792]_ , \new_[66795]_ , \new_[66798]_ , \new_[66799]_ ,
    \new_[66800]_ , \new_[66804]_ , \new_[66805]_ , \new_[66808]_ ,
    \new_[66811]_ , \new_[66812]_ , \new_[66813]_ , \new_[66816]_ ,
    \new_[66819]_ , \new_[66820]_ , \new_[66823]_ , \new_[66826]_ ,
    \new_[66827]_ , \new_[66828]_ , \new_[66832]_ , \new_[66833]_ ,
    \new_[66836]_ , \new_[66839]_ , \new_[66840]_ , \new_[66841]_ ,
    \new_[66844]_ , \new_[66847]_ , \new_[66848]_ , \new_[66851]_ ,
    \new_[66854]_ , \new_[66855]_ , \new_[66856]_ , \new_[66860]_ ,
    \new_[66861]_ , \new_[66864]_ , \new_[66867]_ , \new_[66868]_ ,
    \new_[66869]_ , \new_[66872]_ , \new_[66875]_ , \new_[66876]_ ,
    \new_[66879]_ , \new_[66882]_ , \new_[66883]_ , \new_[66884]_ ,
    \new_[66888]_ , \new_[66889]_ , \new_[66892]_ , \new_[66895]_ ,
    \new_[66896]_ , \new_[66897]_ , \new_[66900]_ , \new_[66903]_ ,
    \new_[66904]_ , \new_[66907]_ , \new_[66910]_ , \new_[66911]_ ,
    \new_[66912]_ , \new_[66916]_ , \new_[66917]_ , \new_[66920]_ ,
    \new_[66923]_ , \new_[66924]_ , \new_[66925]_ , \new_[66928]_ ,
    \new_[66931]_ , \new_[66932]_ , \new_[66935]_ , \new_[66938]_ ,
    \new_[66939]_ , \new_[66940]_ , \new_[66944]_ , \new_[66945]_ ,
    \new_[66948]_ , \new_[66951]_ , \new_[66952]_ , \new_[66953]_ ,
    \new_[66956]_ , \new_[66959]_ , \new_[66960]_ , \new_[66963]_ ,
    \new_[66966]_ , \new_[66967]_ , \new_[66968]_ , \new_[66972]_ ,
    \new_[66973]_ , \new_[66976]_ , \new_[66979]_ , \new_[66980]_ ,
    \new_[66981]_ , \new_[66984]_ , \new_[66987]_ , \new_[66988]_ ,
    \new_[66991]_ , \new_[66994]_ , \new_[66995]_ , \new_[66996]_ ,
    \new_[67000]_ , \new_[67001]_ , \new_[67004]_ , \new_[67007]_ ,
    \new_[67008]_ , \new_[67009]_ , \new_[67012]_ , \new_[67015]_ ,
    \new_[67016]_ , \new_[67019]_ , \new_[67022]_ , \new_[67023]_ ,
    \new_[67024]_ , \new_[67028]_ , \new_[67029]_ , \new_[67032]_ ,
    \new_[67035]_ , \new_[67036]_ , \new_[67037]_ , \new_[67040]_ ,
    \new_[67043]_ , \new_[67044]_ , \new_[67047]_ , \new_[67050]_ ,
    \new_[67051]_ , \new_[67052]_ , \new_[67056]_ , \new_[67057]_ ,
    \new_[67060]_ , \new_[67063]_ , \new_[67064]_ , \new_[67065]_ ,
    \new_[67068]_ , \new_[67071]_ , \new_[67072]_ , \new_[67075]_ ,
    \new_[67078]_ , \new_[67079]_ , \new_[67080]_ , \new_[67084]_ ,
    \new_[67085]_ , \new_[67088]_ , \new_[67091]_ , \new_[67092]_ ,
    \new_[67093]_ , \new_[67096]_ , \new_[67099]_ , \new_[67100]_ ,
    \new_[67103]_ , \new_[67106]_ , \new_[67107]_ , \new_[67108]_ ,
    \new_[67112]_ , \new_[67113]_ , \new_[67116]_ , \new_[67119]_ ,
    \new_[67120]_ , \new_[67121]_ , \new_[67124]_ , \new_[67127]_ ,
    \new_[67128]_ , \new_[67131]_ , \new_[67134]_ , \new_[67135]_ ,
    \new_[67136]_ , \new_[67140]_ , \new_[67141]_ , \new_[67144]_ ,
    \new_[67147]_ , \new_[67148]_ , \new_[67149]_ , \new_[67152]_ ,
    \new_[67155]_ , \new_[67156]_ , \new_[67159]_ , \new_[67162]_ ,
    \new_[67163]_ , \new_[67164]_ , \new_[67168]_ , \new_[67169]_ ,
    \new_[67172]_ , \new_[67175]_ , \new_[67176]_ , \new_[67177]_ ,
    \new_[67180]_ , \new_[67183]_ , \new_[67184]_ , \new_[67187]_ ,
    \new_[67190]_ , \new_[67191]_ , \new_[67192]_ , \new_[67196]_ ,
    \new_[67197]_ , \new_[67200]_ , \new_[67203]_ , \new_[67204]_ ,
    \new_[67205]_ , \new_[67208]_ , \new_[67211]_ , \new_[67212]_ ,
    \new_[67215]_ , \new_[67218]_ , \new_[67219]_ , \new_[67220]_ ,
    \new_[67224]_ , \new_[67225]_ , \new_[67228]_ , \new_[67231]_ ,
    \new_[67232]_ , \new_[67233]_ , \new_[67236]_ , \new_[67239]_ ,
    \new_[67240]_ , \new_[67243]_ , \new_[67246]_ , \new_[67247]_ ,
    \new_[67248]_ , \new_[67252]_ , \new_[67253]_ , \new_[67256]_ ,
    \new_[67259]_ , \new_[67260]_ , \new_[67261]_ , \new_[67264]_ ,
    \new_[67267]_ , \new_[67268]_ , \new_[67271]_ , \new_[67274]_ ,
    \new_[67275]_ , \new_[67276]_ , \new_[67280]_ , \new_[67281]_ ,
    \new_[67284]_ , \new_[67287]_ , \new_[67288]_ , \new_[67289]_ ,
    \new_[67292]_ , \new_[67295]_ , \new_[67296]_ , \new_[67299]_ ,
    \new_[67302]_ , \new_[67303]_ , \new_[67304]_ , \new_[67308]_ ,
    \new_[67309]_ , \new_[67312]_ , \new_[67315]_ , \new_[67316]_ ,
    \new_[67317]_ , \new_[67320]_ , \new_[67323]_ , \new_[67324]_ ,
    \new_[67327]_ , \new_[67330]_ , \new_[67331]_ , \new_[67332]_ ,
    \new_[67336]_ , \new_[67337]_ , \new_[67340]_ , \new_[67343]_ ,
    \new_[67344]_ , \new_[67345]_ , \new_[67348]_ , \new_[67351]_ ,
    \new_[67352]_ , \new_[67355]_ , \new_[67358]_ , \new_[67359]_ ,
    \new_[67360]_ , \new_[67364]_ , \new_[67365]_ , \new_[67368]_ ,
    \new_[67371]_ , \new_[67372]_ , \new_[67373]_ , \new_[67376]_ ,
    \new_[67379]_ , \new_[67380]_ , \new_[67383]_ , \new_[67386]_ ,
    \new_[67387]_ , \new_[67388]_ , \new_[67392]_ , \new_[67393]_ ,
    \new_[67396]_ , \new_[67399]_ , \new_[67400]_ , \new_[67401]_ ,
    \new_[67404]_ , \new_[67407]_ , \new_[67408]_ , \new_[67411]_ ,
    \new_[67414]_ , \new_[67415]_ , \new_[67416]_ , \new_[67420]_ ,
    \new_[67421]_ , \new_[67424]_ , \new_[67427]_ , \new_[67428]_ ,
    \new_[67429]_ , \new_[67432]_ , \new_[67435]_ , \new_[67436]_ ,
    \new_[67439]_ , \new_[67442]_ , \new_[67443]_ , \new_[67444]_ ,
    \new_[67448]_ , \new_[67449]_ , \new_[67452]_ , \new_[67455]_ ,
    \new_[67456]_ , \new_[67457]_ , \new_[67460]_ , \new_[67463]_ ,
    \new_[67464]_ , \new_[67467]_ , \new_[67470]_ , \new_[67471]_ ,
    \new_[67472]_ , \new_[67476]_ , \new_[67477]_ , \new_[67480]_ ,
    \new_[67483]_ , \new_[67484]_ , \new_[67485]_ , \new_[67488]_ ,
    \new_[67491]_ , \new_[67492]_ , \new_[67495]_ , \new_[67498]_ ,
    \new_[67499]_ , \new_[67500]_ , \new_[67504]_ , \new_[67505]_ ,
    \new_[67508]_ , \new_[67511]_ , \new_[67512]_ , \new_[67513]_ ,
    \new_[67516]_ , \new_[67519]_ , \new_[67520]_ , \new_[67523]_ ,
    \new_[67526]_ , \new_[67527]_ , \new_[67528]_ , \new_[67532]_ ,
    \new_[67533]_ , \new_[67536]_ , \new_[67539]_ , \new_[67540]_ ,
    \new_[67541]_ , \new_[67544]_ , \new_[67547]_ , \new_[67548]_ ,
    \new_[67551]_ , \new_[67554]_ , \new_[67555]_ , \new_[67556]_ ,
    \new_[67560]_ , \new_[67561]_ , \new_[67564]_ , \new_[67567]_ ,
    \new_[67568]_ , \new_[67569]_ , \new_[67572]_ , \new_[67575]_ ,
    \new_[67576]_ , \new_[67579]_ , \new_[67582]_ , \new_[67583]_ ,
    \new_[67584]_ , \new_[67588]_ , \new_[67589]_ , \new_[67592]_ ,
    \new_[67595]_ , \new_[67596]_ , \new_[67597]_ , \new_[67600]_ ,
    \new_[67603]_ , \new_[67604]_ , \new_[67607]_ , \new_[67610]_ ,
    \new_[67611]_ , \new_[67612]_ , \new_[67616]_ , \new_[67617]_ ,
    \new_[67620]_ , \new_[67623]_ , \new_[67624]_ , \new_[67625]_ ,
    \new_[67628]_ , \new_[67631]_ , \new_[67632]_ , \new_[67635]_ ,
    \new_[67638]_ , \new_[67639]_ , \new_[67640]_ , \new_[67644]_ ,
    \new_[67645]_ , \new_[67648]_ , \new_[67651]_ , \new_[67652]_ ,
    \new_[67653]_ , \new_[67656]_ , \new_[67659]_ , \new_[67660]_ ,
    \new_[67663]_ , \new_[67666]_ , \new_[67667]_ , \new_[67668]_ ,
    \new_[67672]_ , \new_[67673]_ , \new_[67676]_ , \new_[67679]_ ,
    \new_[67680]_ , \new_[67681]_ , \new_[67684]_ , \new_[67687]_ ,
    \new_[67688]_ , \new_[67691]_ , \new_[67694]_ , \new_[67695]_ ,
    \new_[67696]_ , \new_[67700]_ , \new_[67701]_ , \new_[67704]_ ,
    \new_[67707]_ , \new_[67708]_ , \new_[67709]_ , \new_[67712]_ ,
    \new_[67715]_ , \new_[67716]_ , \new_[67719]_ , \new_[67722]_ ,
    \new_[67723]_ , \new_[67724]_ , \new_[67728]_ , \new_[67729]_ ,
    \new_[67732]_ , \new_[67735]_ , \new_[67736]_ , \new_[67737]_ ,
    \new_[67740]_ , \new_[67743]_ , \new_[67744]_ , \new_[67747]_ ,
    \new_[67750]_ , \new_[67751]_ , \new_[67752]_ , \new_[67756]_ ,
    \new_[67757]_ , \new_[67760]_ , \new_[67763]_ , \new_[67764]_ ,
    \new_[67765]_ , \new_[67768]_ , \new_[67771]_ , \new_[67772]_ ,
    \new_[67775]_ , \new_[67778]_ , \new_[67779]_ , \new_[67780]_ ,
    \new_[67784]_ , \new_[67785]_ , \new_[67788]_ , \new_[67791]_ ,
    \new_[67792]_ , \new_[67793]_ , \new_[67796]_ , \new_[67799]_ ,
    \new_[67800]_ , \new_[67803]_ , \new_[67806]_ , \new_[67807]_ ,
    \new_[67808]_ , \new_[67812]_ , \new_[67813]_ , \new_[67816]_ ,
    \new_[67819]_ , \new_[67820]_ , \new_[67821]_ , \new_[67824]_ ,
    \new_[67827]_ , \new_[67828]_ , \new_[67831]_ , \new_[67834]_ ,
    \new_[67835]_ , \new_[67836]_ , \new_[67840]_ , \new_[67841]_ ,
    \new_[67844]_ , \new_[67847]_ , \new_[67848]_ , \new_[67849]_ ,
    \new_[67852]_ , \new_[67855]_ , \new_[67856]_ , \new_[67859]_ ,
    \new_[67862]_ , \new_[67863]_ , \new_[67864]_ , \new_[67868]_ ,
    \new_[67869]_ , \new_[67872]_ , \new_[67875]_ , \new_[67876]_ ,
    \new_[67877]_ , \new_[67880]_ , \new_[67883]_ , \new_[67884]_ ,
    \new_[67887]_ , \new_[67890]_ , \new_[67891]_ , \new_[67892]_ ,
    \new_[67896]_ , \new_[67897]_ , \new_[67900]_ , \new_[67903]_ ,
    \new_[67904]_ , \new_[67905]_ , \new_[67908]_ , \new_[67911]_ ,
    \new_[67912]_ , \new_[67915]_ , \new_[67918]_ , \new_[67919]_ ,
    \new_[67920]_ , \new_[67924]_ , \new_[67925]_ , \new_[67928]_ ,
    \new_[67931]_ , \new_[67932]_ , \new_[67933]_ , \new_[67936]_ ,
    \new_[67939]_ , \new_[67940]_ , \new_[67943]_ , \new_[67946]_ ,
    \new_[67947]_ , \new_[67948]_ , \new_[67952]_ , \new_[67953]_ ,
    \new_[67956]_ , \new_[67959]_ , \new_[67960]_ , \new_[67961]_ ,
    \new_[67964]_ , \new_[67967]_ , \new_[67968]_ , \new_[67971]_ ,
    \new_[67974]_ , \new_[67975]_ , \new_[67976]_ , \new_[67980]_ ,
    \new_[67981]_ , \new_[67984]_ , \new_[67987]_ , \new_[67988]_ ,
    \new_[67989]_ , \new_[67992]_ , \new_[67995]_ , \new_[67996]_ ,
    \new_[67999]_ , \new_[68002]_ , \new_[68003]_ , \new_[68004]_ ,
    \new_[68008]_ , \new_[68009]_ , \new_[68012]_ , \new_[68015]_ ,
    \new_[68016]_ , \new_[68017]_ , \new_[68020]_ , \new_[68023]_ ,
    \new_[68024]_ , \new_[68027]_ , \new_[68030]_ , \new_[68031]_ ,
    \new_[68032]_ , \new_[68036]_ , \new_[68037]_ , \new_[68040]_ ,
    \new_[68043]_ , \new_[68044]_ , \new_[68045]_ , \new_[68048]_ ,
    \new_[68051]_ , \new_[68052]_ , \new_[68055]_ , \new_[68058]_ ,
    \new_[68059]_ , \new_[68060]_ , \new_[68064]_ , \new_[68065]_ ,
    \new_[68068]_ , \new_[68071]_ , \new_[68072]_ , \new_[68073]_ ,
    \new_[68076]_ , \new_[68079]_ , \new_[68080]_ , \new_[68083]_ ,
    \new_[68086]_ , \new_[68087]_ , \new_[68088]_ , \new_[68092]_ ,
    \new_[68093]_ , \new_[68096]_ , \new_[68099]_ , \new_[68100]_ ,
    \new_[68101]_ , \new_[68104]_ , \new_[68107]_ , \new_[68108]_ ,
    \new_[68111]_ , \new_[68114]_ , \new_[68115]_ , \new_[68116]_ ,
    \new_[68120]_ , \new_[68121]_ , \new_[68124]_ , \new_[68127]_ ,
    \new_[68128]_ , \new_[68129]_ , \new_[68132]_ , \new_[68135]_ ,
    \new_[68136]_ , \new_[68139]_ , \new_[68142]_ , \new_[68143]_ ,
    \new_[68144]_ , \new_[68148]_ , \new_[68149]_ , \new_[68152]_ ,
    \new_[68155]_ , \new_[68156]_ , \new_[68157]_ , \new_[68160]_ ,
    \new_[68163]_ , \new_[68164]_ , \new_[68167]_ , \new_[68170]_ ,
    \new_[68171]_ , \new_[68172]_ , \new_[68176]_ , \new_[68177]_ ,
    \new_[68180]_ , \new_[68183]_ , \new_[68184]_ , \new_[68185]_ ,
    \new_[68188]_ , \new_[68191]_ , \new_[68192]_ , \new_[68195]_ ,
    \new_[68198]_ , \new_[68199]_ , \new_[68200]_ , \new_[68204]_ ,
    \new_[68205]_ , \new_[68208]_ , \new_[68211]_ , \new_[68212]_ ,
    \new_[68213]_ , \new_[68216]_ , \new_[68219]_ , \new_[68220]_ ,
    \new_[68223]_ , \new_[68226]_ , \new_[68227]_ , \new_[68228]_ ,
    \new_[68232]_ , \new_[68233]_ , \new_[68236]_ , \new_[68239]_ ,
    \new_[68240]_ , \new_[68241]_ , \new_[68244]_ , \new_[68247]_ ,
    \new_[68248]_ , \new_[68251]_ , \new_[68254]_ , \new_[68255]_ ,
    \new_[68256]_ , \new_[68260]_ , \new_[68261]_ , \new_[68264]_ ,
    \new_[68267]_ , \new_[68268]_ , \new_[68269]_ , \new_[68272]_ ,
    \new_[68275]_ , \new_[68276]_ , \new_[68279]_ , \new_[68282]_ ,
    \new_[68283]_ , \new_[68284]_ , \new_[68288]_ , \new_[68289]_ ,
    \new_[68292]_ , \new_[68295]_ , \new_[68296]_ , \new_[68297]_ ,
    \new_[68300]_ , \new_[68303]_ , \new_[68304]_ , \new_[68307]_ ,
    \new_[68310]_ , \new_[68311]_ , \new_[68312]_ , \new_[68316]_ ,
    \new_[68317]_ , \new_[68320]_ , \new_[68323]_ , \new_[68324]_ ,
    \new_[68325]_ , \new_[68328]_ , \new_[68331]_ , \new_[68332]_ ,
    \new_[68335]_ , \new_[68338]_ , \new_[68339]_ , \new_[68340]_ ,
    \new_[68344]_ , \new_[68345]_ , \new_[68348]_ , \new_[68351]_ ,
    \new_[68352]_ , \new_[68353]_ , \new_[68356]_ , \new_[68359]_ ,
    \new_[68360]_ , \new_[68363]_ , \new_[68366]_ , \new_[68367]_ ,
    \new_[68368]_ , \new_[68372]_ , \new_[68373]_ , \new_[68376]_ ,
    \new_[68379]_ , \new_[68380]_ , \new_[68381]_ , \new_[68384]_ ,
    \new_[68387]_ , \new_[68388]_ , \new_[68391]_ , \new_[68394]_ ,
    \new_[68395]_ , \new_[68396]_ , \new_[68400]_ , \new_[68401]_ ,
    \new_[68404]_ , \new_[68407]_ , \new_[68408]_ , \new_[68409]_ ,
    \new_[68412]_ , \new_[68415]_ , \new_[68416]_ , \new_[68419]_ ,
    \new_[68422]_ , \new_[68423]_ , \new_[68424]_ , \new_[68428]_ ,
    \new_[68429]_ , \new_[68432]_ , \new_[68435]_ , \new_[68436]_ ,
    \new_[68437]_ , \new_[68440]_ , \new_[68443]_ , \new_[68444]_ ,
    \new_[68447]_ , \new_[68450]_ , \new_[68451]_ , \new_[68452]_ ,
    \new_[68456]_ , \new_[68457]_ , \new_[68460]_ , \new_[68463]_ ,
    \new_[68464]_ , \new_[68465]_ , \new_[68468]_ , \new_[68471]_ ,
    \new_[68472]_ , \new_[68475]_ , \new_[68478]_ , \new_[68479]_ ,
    \new_[68480]_ , \new_[68484]_ , \new_[68485]_ , \new_[68488]_ ,
    \new_[68491]_ , \new_[68492]_ , \new_[68493]_ , \new_[68496]_ ,
    \new_[68499]_ , \new_[68500]_ , \new_[68503]_ , \new_[68506]_ ,
    \new_[68507]_ , \new_[68508]_ , \new_[68512]_ , \new_[68513]_ ,
    \new_[68516]_ , \new_[68519]_ , \new_[68520]_ , \new_[68521]_ ,
    \new_[68524]_ , \new_[68527]_ , \new_[68528]_ , \new_[68531]_ ,
    \new_[68534]_ , \new_[68535]_ , \new_[68536]_ , \new_[68540]_ ,
    \new_[68541]_ , \new_[68544]_ , \new_[68547]_ , \new_[68548]_ ,
    \new_[68549]_ , \new_[68552]_ , \new_[68555]_ , \new_[68556]_ ,
    \new_[68559]_ , \new_[68562]_ , \new_[68563]_ , \new_[68564]_ ,
    \new_[68568]_ , \new_[68569]_ , \new_[68572]_ , \new_[68575]_ ,
    \new_[68576]_ , \new_[68577]_ , \new_[68580]_ , \new_[68583]_ ,
    \new_[68584]_ , \new_[68587]_ , \new_[68590]_ , \new_[68591]_ ,
    \new_[68592]_ , \new_[68596]_ , \new_[68597]_ , \new_[68600]_ ,
    \new_[68603]_ , \new_[68604]_ , \new_[68605]_ , \new_[68608]_ ,
    \new_[68611]_ , \new_[68612]_ , \new_[68615]_ , \new_[68618]_ ,
    \new_[68619]_ , \new_[68620]_ , \new_[68624]_ , \new_[68625]_ ,
    \new_[68628]_ , \new_[68631]_ , \new_[68632]_ , \new_[68633]_ ,
    \new_[68636]_ , \new_[68639]_ , \new_[68640]_ , \new_[68643]_ ,
    \new_[68646]_ , \new_[68647]_ , \new_[68648]_ , \new_[68652]_ ,
    \new_[68653]_ , \new_[68656]_ , \new_[68659]_ , \new_[68660]_ ,
    \new_[68661]_ , \new_[68664]_ , \new_[68667]_ , \new_[68668]_ ,
    \new_[68671]_ , \new_[68674]_ , \new_[68675]_ , \new_[68676]_ ,
    \new_[68680]_ , \new_[68681]_ , \new_[68684]_ , \new_[68687]_ ,
    \new_[68688]_ , \new_[68689]_ , \new_[68692]_ , \new_[68695]_ ,
    \new_[68696]_ , \new_[68699]_ , \new_[68702]_ , \new_[68703]_ ,
    \new_[68704]_ , \new_[68708]_ , \new_[68709]_ , \new_[68712]_ ,
    \new_[68715]_ , \new_[68716]_ , \new_[68717]_ , \new_[68720]_ ,
    \new_[68723]_ , \new_[68724]_ , \new_[68727]_ , \new_[68730]_ ,
    \new_[68731]_ , \new_[68732]_ , \new_[68736]_ , \new_[68737]_ ,
    \new_[68740]_ , \new_[68743]_ , \new_[68744]_ , \new_[68745]_ ,
    \new_[68748]_ , \new_[68751]_ , \new_[68752]_ , \new_[68755]_ ,
    \new_[68758]_ , \new_[68759]_ , \new_[68760]_ , \new_[68764]_ ,
    \new_[68765]_ , \new_[68768]_ , \new_[68771]_ , \new_[68772]_ ,
    \new_[68773]_ , \new_[68776]_ , \new_[68779]_ , \new_[68780]_ ,
    \new_[68783]_ , \new_[68786]_ , \new_[68787]_ , \new_[68788]_ ,
    \new_[68792]_ , \new_[68793]_ , \new_[68796]_ , \new_[68799]_ ,
    \new_[68800]_ , \new_[68801]_ , \new_[68804]_ , \new_[68807]_ ,
    \new_[68808]_ , \new_[68811]_ , \new_[68814]_ , \new_[68815]_ ,
    \new_[68816]_ , \new_[68820]_ , \new_[68821]_ , \new_[68824]_ ,
    \new_[68827]_ , \new_[68828]_ , \new_[68829]_ , \new_[68832]_ ,
    \new_[68835]_ , \new_[68836]_ , \new_[68839]_ , \new_[68842]_ ,
    \new_[68843]_ , \new_[68844]_ , \new_[68848]_ , \new_[68849]_ ,
    \new_[68852]_ , \new_[68855]_ , \new_[68856]_ , \new_[68857]_ ,
    \new_[68860]_ , \new_[68863]_ , \new_[68864]_ , \new_[68867]_ ,
    \new_[68870]_ , \new_[68871]_ , \new_[68872]_ , \new_[68876]_ ,
    \new_[68877]_ , \new_[68880]_ , \new_[68883]_ , \new_[68884]_ ,
    \new_[68885]_ , \new_[68888]_ , \new_[68891]_ , \new_[68892]_ ,
    \new_[68895]_ , \new_[68898]_ , \new_[68899]_ , \new_[68900]_ ,
    \new_[68904]_ , \new_[68905]_ , \new_[68908]_ , \new_[68911]_ ,
    \new_[68912]_ , \new_[68913]_ , \new_[68916]_ , \new_[68919]_ ,
    \new_[68920]_ , \new_[68923]_ , \new_[68926]_ , \new_[68927]_ ,
    \new_[68928]_ , \new_[68932]_ , \new_[68933]_ , \new_[68936]_ ,
    \new_[68939]_ , \new_[68940]_ , \new_[68941]_ , \new_[68944]_ ,
    \new_[68947]_ , \new_[68948]_ , \new_[68951]_ , \new_[68954]_ ,
    \new_[68955]_ , \new_[68956]_ , \new_[68960]_ , \new_[68961]_ ,
    \new_[68964]_ , \new_[68967]_ , \new_[68968]_ , \new_[68969]_ ,
    \new_[68972]_ , \new_[68975]_ , \new_[68976]_ , \new_[68979]_ ,
    \new_[68982]_ , \new_[68983]_ , \new_[68984]_ , \new_[68988]_ ,
    \new_[68989]_ , \new_[68992]_ , \new_[68995]_ , \new_[68996]_ ,
    \new_[68997]_ , \new_[69000]_ , \new_[69003]_ , \new_[69004]_ ,
    \new_[69007]_ , \new_[69010]_ , \new_[69011]_ , \new_[69012]_ ,
    \new_[69016]_ , \new_[69017]_ , \new_[69020]_ , \new_[69023]_ ,
    \new_[69024]_ , \new_[69025]_ , \new_[69028]_ , \new_[69031]_ ,
    \new_[69032]_ , \new_[69035]_ , \new_[69038]_ , \new_[69039]_ ,
    \new_[69040]_ , \new_[69044]_ , \new_[69045]_ , \new_[69048]_ ,
    \new_[69051]_ , \new_[69052]_ , \new_[69053]_ , \new_[69056]_ ,
    \new_[69059]_ , \new_[69060]_ , \new_[69063]_ , \new_[69066]_ ,
    \new_[69067]_ , \new_[69068]_ , \new_[69072]_ , \new_[69073]_ ,
    \new_[69076]_ , \new_[69079]_ , \new_[69080]_ , \new_[69081]_ ,
    \new_[69084]_ , \new_[69087]_ , \new_[69088]_ , \new_[69091]_ ,
    \new_[69094]_ , \new_[69095]_ , \new_[69096]_ , \new_[69100]_ ,
    \new_[69101]_ , \new_[69104]_ , \new_[69107]_ , \new_[69108]_ ,
    \new_[69109]_ , \new_[69112]_ , \new_[69115]_ , \new_[69116]_ ,
    \new_[69119]_ , \new_[69122]_ , \new_[69123]_ , \new_[69124]_ ,
    \new_[69128]_ , \new_[69129]_ , \new_[69132]_ , \new_[69135]_ ,
    \new_[69136]_ , \new_[69137]_ , \new_[69140]_ , \new_[69143]_ ,
    \new_[69144]_ , \new_[69147]_ , \new_[69150]_ , \new_[69151]_ ,
    \new_[69152]_ , \new_[69156]_ , \new_[69157]_ , \new_[69160]_ ,
    \new_[69163]_ , \new_[69164]_ , \new_[69165]_ , \new_[69168]_ ,
    \new_[69171]_ , \new_[69172]_ , \new_[69175]_ , \new_[69178]_ ,
    \new_[69179]_ , \new_[69180]_ , \new_[69184]_ , \new_[69185]_ ,
    \new_[69188]_ , \new_[69191]_ , \new_[69192]_ , \new_[69193]_ ,
    \new_[69196]_ , \new_[69199]_ , \new_[69200]_ , \new_[69203]_ ,
    \new_[69206]_ , \new_[69207]_ , \new_[69208]_ , \new_[69212]_ ,
    \new_[69213]_ , \new_[69216]_ , \new_[69219]_ , \new_[69220]_ ,
    \new_[69221]_ , \new_[69224]_ , \new_[69227]_ , \new_[69228]_ ,
    \new_[69231]_ , \new_[69234]_ , \new_[69235]_ , \new_[69236]_ ,
    \new_[69240]_ , \new_[69241]_ , \new_[69244]_ , \new_[69247]_ ,
    \new_[69248]_ , \new_[69249]_ , \new_[69252]_ , \new_[69255]_ ,
    \new_[69256]_ , \new_[69259]_ , \new_[69262]_ , \new_[69263]_ ,
    \new_[69264]_ , \new_[69268]_ , \new_[69269]_ , \new_[69272]_ ,
    \new_[69275]_ , \new_[69276]_ , \new_[69277]_ , \new_[69280]_ ,
    \new_[69283]_ , \new_[69284]_ , \new_[69287]_ , \new_[69290]_ ,
    \new_[69291]_ , \new_[69292]_ , \new_[69296]_ , \new_[69297]_ ,
    \new_[69300]_ , \new_[69303]_ , \new_[69304]_ , \new_[69305]_ ,
    \new_[69308]_ , \new_[69311]_ , \new_[69312]_ , \new_[69315]_ ,
    \new_[69318]_ , \new_[69319]_ , \new_[69320]_ , \new_[69324]_ ,
    \new_[69325]_ , \new_[69328]_ , \new_[69331]_ , \new_[69332]_ ,
    \new_[69333]_ , \new_[69336]_ , \new_[69339]_ , \new_[69340]_ ,
    \new_[69343]_ , \new_[69346]_ , \new_[69347]_ , \new_[69348]_ ,
    \new_[69352]_ , \new_[69353]_ , \new_[69356]_ , \new_[69359]_ ,
    \new_[69360]_ , \new_[69361]_ , \new_[69364]_ , \new_[69367]_ ,
    \new_[69368]_ , \new_[69371]_ , \new_[69374]_ , \new_[69375]_ ,
    \new_[69376]_ , \new_[69380]_ , \new_[69381]_ , \new_[69384]_ ,
    \new_[69387]_ , \new_[69388]_ , \new_[69389]_ , \new_[69392]_ ,
    \new_[69395]_ , \new_[69396]_ , \new_[69399]_ , \new_[69402]_ ,
    \new_[69403]_ , \new_[69404]_ , \new_[69408]_ , \new_[69409]_ ,
    \new_[69412]_ , \new_[69415]_ , \new_[69416]_ , \new_[69417]_ ,
    \new_[69420]_ , \new_[69423]_ , \new_[69424]_ , \new_[69427]_ ,
    \new_[69430]_ , \new_[69431]_ , \new_[69432]_ , \new_[69436]_ ,
    \new_[69437]_ , \new_[69440]_ , \new_[69443]_ , \new_[69444]_ ,
    \new_[69445]_ , \new_[69448]_ , \new_[69451]_ , \new_[69452]_ ,
    \new_[69455]_ , \new_[69458]_ , \new_[69459]_ , \new_[69460]_ ,
    \new_[69464]_ , \new_[69465]_ , \new_[69468]_ , \new_[69471]_ ,
    \new_[69472]_ , \new_[69473]_ , \new_[69476]_ , \new_[69479]_ ,
    \new_[69480]_ , \new_[69483]_ , \new_[69486]_ , \new_[69487]_ ,
    \new_[69488]_ , \new_[69492]_ , \new_[69493]_ , \new_[69496]_ ,
    \new_[69499]_ , \new_[69500]_ , \new_[69501]_ , \new_[69504]_ ,
    \new_[69507]_ , \new_[69508]_ , \new_[69511]_ , \new_[69514]_ ,
    \new_[69515]_ , \new_[69516]_ , \new_[69520]_ , \new_[69521]_ ,
    \new_[69524]_ , \new_[69527]_ , \new_[69528]_ , \new_[69529]_ ,
    \new_[69532]_ , \new_[69535]_ , \new_[69536]_ , \new_[69539]_ ,
    \new_[69542]_ , \new_[69543]_ , \new_[69544]_ , \new_[69548]_ ,
    \new_[69549]_ , \new_[69552]_ , \new_[69555]_ , \new_[69556]_ ,
    \new_[69557]_ , \new_[69560]_ , \new_[69563]_ , \new_[69564]_ ,
    \new_[69567]_ , \new_[69570]_ , \new_[69571]_ , \new_[69572]_ ,
    \new_[69576]_ , \new_[69577]_ , \new_[69580]_ , \new_[69583]_ ,
    \new_[69584]_ , \new_[69585]_ , \new_[69588]_ , \new_[69591]_ ,
    \new_[69592]_ , \new_[69595]_ , \new_[69598]_ , \new_[69599]_ ,
    \new_[69600]_ , \new_[69604]_ , \new_[69605]_ , \new_[69608]_ ,
    \new_[69611]_ , \new_[69612]_ , \new_[69613]_ , \new_[69616]_ ,
    \new_[69619]_ , \new_[69620]_ , \new_[69623]_ , \new_[69626]_ ,
    \new_[69627]_ , \new_[69628]_ , \new_[69632]_ , \new_[69633]_ ,
    \new_[69636]_ , \new_[69639]_ , \new_[69640]_ , \new_[69641]_ ,
    \new_[69644]_ , \new_[69647]_ , \new_[69648]_ , \new_[69651]_ ,
    \new_[69654]_ , \new_[69655]_ , \new_[69656]_ , \new_[69660]_ ,
    \new_[69661]_ , \new_[69664]_ , \new_[69667]_ , \new_[69668]_ ,
    \new_[69669]_ , \new_[69672]_ , \new_[69675]_ , \new_[69676]_ ,
    \new_[69679]_ , \new_[69682]_ , \new_[69683]_ , \new_[69684]_ ,
    \new_[69688]_ , \new_[69689]_ , \new_[69692]_ , \new_[69695]_ ,
    \new_[69696]_ , \new_[69697]_ , \new_[69700]_ , \new_[69703]_ ,
    \new_[69704]_ , \new_[69707]_ , \new_[69710]_ , \new_[69711]_ ,
    \new_[69712]_ , \new_[69716]_ , \new_[69717]_ , \new_[69720]_ ,
    \new_[69723]_ , \new_[69724]_ , \new_[69725]_ , \new_[69728]_ ,
    \new_[69731]_ , \new_[69732]_ , \new_[69735]_ , \new_[69738]_ ,
    \new_[69739]_ , \new_[69740]_ , \new_[69744]_ , \new_[69745]_ ,
    \new_[69748]_ , \new_[69751]_ , \new_[69752]_ , \new_[69753]_ ,
    \new_[69756]_ , \new_[69759]_ , \new_[69760]_ , \new_[69763]_ ,
    \new_[69766]_ , \new_[69767]_ , \new_[69768]_ , \new_[69772]_ ,
    \new_[69773]_ , \new_[69776]_ , \new_[69779]_ , \new_[69780]_ ,
    \new_[69781]_ , \new_[69784]_ , \new_[69787]_ , \new_[69788]_ ,
    \new_[69791]_ , \new_[69794]_ , \new_[69795]_ , \new_[69796]_ ,
    \new_[69800]_ , \new_[69801]_ , \new_[69804]_ , \new_[69807]_ ,
    \new_[69808]_ , \new_[69809]_ , \new_[69812]_ , \new_[69815]_ ,
    \new_[69816]_ , \new_[69819]_ , \new_[69822]_ , \new_[69823]_ ,
    \new_[69824]_ , \new_[69828]_ , \new_[69829]_ , \new_[69832]_ ,
    \new_[69835]_ , \new_[69836]_ , \new_[69837]_ , \new_[69840]_ ,
    \new_[69843]_ , \new_[69844]_ , \new_[69847]_ , \new_[69850]_ ,
    \new_[69851]_ , \new_[69852]_ , \new_[69856]_ , \new_[69857]_ ,
    \new_[69860]_ , \new_[69863]_ , \new_[69864]_ , \new_[69865]_ ,
    \new_[69868]_ , \new_[69871]_ , \new_[69872]_ , \new_[69875]_ ,
    \new_[69878]_ , \new_[69879]_ , \new_[69880]_ , \new_[69884]_ ,
    \new_[69885]_ , \new_[69888]_ , \new_[69891]_ , \new_[69892]_ ,
    \new_[69893]_ , \new_[69896]_ , \new_[69899]_ , \new_[69900]_ ,
    \new_[69903]_ , \new_[69906]_ , \new_[69907]_ , \new_[69908]_ ,
    \new_[69912]_ , \new_[69913]_ , \new_[69916]_ , \new_[69919]_ ,
    \new_[69920]_ , \new_[69921]_ , \new_[69924]_ , \new_[69927]_ ,
    \new_[69928]_ , \new_[69931]_ , \new_[69934]_ , \new_[69935]_ ,
    \new_[69936]_ , \new_[69940]_ , \new_[69941]_ , \new_[69944]_ ,
    \new_[69947]_ , \new_[69948]_ , \new_[69949]_ , \new_[69952]_ ,
    \new_[69955]_ , \new_[69956]_ , \new_[69959]_ , \new_[69962]_ ,
    \new_[69963]_ , \new_[69964]_ , \new_[69968]_ , \new_[69969]_ ,
    \new_[69972]_ , \new_[69975]_ , \new_[69976]_ , \new_[69977]_ ,
    \new_[69980]_ , \new_[69983]_ , \new_[69984]_ , \new_[69987]_ ,
    \new_[69990]_ , \new_[69991]_ , \new_[69992]_ , \new_[69996]_ ,
    \new_[69997]_ , \new_[70000]_ , \new_[70003]_ , \new_[70004]_ ,
    \new_[70005]_ , \new_[70008]_ , \new_[70011]_ , \new_[70012]_ ,
    \new_[70015]_ , \new_[70018]_ , \new_[70019]_ , \new_[70020]_ ,
    \new_[70024]_ , \new_[70025]_ , \new_[70028]_ , \new_[70031]_ ,
    \new_[70032]_ , \new_[70033]_ , \new_[70036]_ , \new_[70039]_ ,
    \new_[70040]_ , \new_[70043]_ , \new_[70046]_ , \new_[70047]_ ,
    \new_[70048]_ , \new_[70052]_ , \new_[70053]_ , \new_[70056]_ ,
    \new_[70059]_ , \new_[70060]_ , \new_[70061]_ , \new_[70064]_ ,
    \new_[70067]_ , \new_[70068]_ , \new_[70071]_ , \new_[70074]_ ,
    \new_[70075]_ , \new_[70076]_ , \new_[70080]_ , \new_[70081]_ ,
    \new_[70084]_ , \new_[70087]_ , \new_[70088]_ , \new_[70089]_ ,
    \new_[70092]_ , \new_[70095]_ , \new_[70096]_ , \new_[70099]_ ,
    \new_[70102]_ , \new_[70103]_ , \new_[70104]_ , \new_[70108]_ ,
    \new_[70109]_ , \new_[70112]_ , \new_[70115]_ , \new_[70116]_ ,
    \new_[70117]_ , \new_[70120]_ , \new_[70123]_ , \new_[70124]_ ,
    \new_[70127]_ , \new_[70130]_ , \new_[70131]_ , \new_[70132]_ ,
    \new_[70136]_ , \new_[70137]_ , \new_[70140]_ , \new_[70143]_ ,
    \new_[70144]_ , \new_[70145]_ , \new_[70148]_ , \new_[70151]_ ,
    \new_[70152]_ , \new_[70155]_ , \new_[70158]_ , \new_[70159]_ ,
    \new_[70160]_ , \new_[70164]_ , \new_[70165]_ , \new_[70168]_ ,
    \new_[70171]_ , \new_[70172]_ , \new_[70173]_ , \new_[70176]_ ,
    \new_[70179]_ , \new_[70180]_ , \new_[70183]_ , \new_[70186]_ ,
    \new_[70187]_ , \new_[70188]_ , \new_[70192]_ , \new_[70193]_ ,
    \new_[70196]_ , \new_[70199]_ , \new_[70200]_ , \new_[70201]_ ,
    \new_[70204]_ , \new_[70207]_ , \new_[70208]_ , \new_[70211]_ ,
    \new_[70214]_ , \new_[70215]_ , \new_[70216]_ , \new_[70220]_ ,
    \new_[70221]_ , \new_[70224]_ , \new_[70227]_ , \new_[70228]_ ,
    \new_[70229]_ , \new_[70232]_ , \new_[70235]_ , \new_[70236]_ ,
    \new_[70239]_ , \new_[70242]_ , \new_[70243]_ , \new_[70244]_ ,
    \new_[70248]_ , \new_[70249]_ , \new_[70252]_ , \new_[70255]_ ,
    \new_[70256]_ , \new_[70257]_ , \new_[70260]_ , \new_[70263]_ ,
    \new_[70264]_ , \new_[70267]_ , \new_[70270]_ , \new_[70271]_ ,
    \new_[70272]_ , \new_[70276]_ , \new_[70277]_ , \new_[70280]_ ,
    \new_[70283]_ , \new_[70284]_ , \new_[70285]_ , \new_[70288]_ ,
    \new_[70291]_ , \new_[70292]_ , \new_[70295]_ , \new_[70298]_ ,
    \new_[70299]_ , \new_[70300]_ , \new_[70304]_ , \new_[70305]_ ,
    \new_[70308]_ , \new_[70311]_ , \new_[70312]_ , \new_[70313]_ ,
    \new_[70316]_ , \new_[70319]_ , \new_[70320]_ , \new_[70323]_ ,
    \new_[70326]_ , \new_[70327]_ , \new_[70328]_ , \new_[70332]_ ,
    \new_[70333]_ , \new_[70336]_ , \new_[70339]_ , \new_[70340]_ ,
    \new_[70341]_ , \new_[70344]_ , \new_[70347]_ , \new_[70348]_ ,
    \new_[70351]_ , \new_[70354]_ , \new_[70355]_ , \new_[70356]_ ,
    \new_[70360]_ , \new_[70361]_ , \new_[70364]_ , \new_[70367]_ ,
    \new_[70368]_ , \new_[70369]_ , \new_[70372]_ , \new_[70375]_ ,
    \new_[70376]_ , \new_[70379]_ , \new_[70382]_ , \new_[70383]_ ,
    \new_[70384]_ , \new_[70388]_ , \new_[70389]_ , \new_[70392]_ ,
    \new_[70395]_ , \new_[70396]_ , \new_[70397]_ , \new_[70400]_ ,
    \new_[70403]_ , \new_[70404]_ , \new_[70407]_ , \new_[70410]_ ,
    \new_[70411]_ , \new_[70412]_ , \new_[70416]_ , \new_[70417]_ ,
    \new_[70420]_ , \new_[70423]_ , \new_[70424]_ , \new_[70425]_ ,
    \new_[70428]_ , \new_[70431]_ , \new_[70432]_ , \new_[70435]_ ,
    \new_[70438]_ , \new_[70439]_ , \new_[70440]_ , \new_[70444]_ ,
    \new_[70445]_ , \new_[70448]_ , \new_[70451]_ , \new_[70452]_ ,
    \new_[70453]_ , \new_[70456]_ , \new_[70459]_ , \new_[70460]_ ,
    \new_[70463]_ , \new_[70466]_ , \new_[70467]_ , \new_[70468]_ ,
    \new_[70472]_ , \new_[70473]_ , \new_[70476]_ , \new_[70479]_ ,
    \new_[70480]_ , \new_[70481]_ , \new_[70484]_ , \new_[70487]_ ,
    \new_[70488]_ , \new_[70491]_ , \new_[70494]_ , \new_[70495]_ ,
    \new_[70496]_ , \new_[70500]_ , \new_[70501]_ , \new_[70504]_ ,
    \new_[70507]_ , \new_[70508]_ , \new_[70509]_ , \new_[70512]_ ,
    \new_[70515]_ , \new_[70516]_ , \new_[70519]_ , \new_[70522]_ ,
    \new_[70523]_ , \new_[70524]_ , \new_[70528]_ , \new_[70529]_ ,
    \new_[70532]_ , \new_[70535]_ , \new_[70536]_ , \new_[70537]_ ,
    \new_[70540]_ , \new_[70543]_ , \new_[70544]_ , \new_[70547]_ ,
    \new_[70550]_ , \new_[70551]_ , \new_[70552]_ , \new_[70556]_ ,
    \new_[70557]_ , \new_[70560]_ , \new_[70563]_ , \new_[70564]_ ,
    \new_[70565]_ , \new_[70568]_ , \new_[70571]_ , \new_[70572]_ ,
    \new_[70575]_ , \new_[70578]_ , \new_[70579]_ , \new_[70580]_ ,
    \new_[70584]_ , \new_[70585]_ , \new_[70588]_ , \new_[70591]_ ,
    \new_[70592]_ , \new_[70593]_ , \new_[70596]_ , \new_[70599]_ ,
    \new_[70600]_ , \new_[70603]_ , \new_[70606]_ , \new_[70607]_ ,
    \new_[70608]_ , \new_[70612]_ , \new_[70613]_ , \new_[70616]_ ,
    \new_[70619]_ , \new_[70620]_ , \new_[70621]_ , \new_[70624]_ ,
    \new_[70627]_ , \new_[70628]_ , \new_[70631]_ , \new_[70634]_ ,
    \new_[70635]_ , \new_[70636]_ , \new_[70640]_ , \new_[70641]_ ,
    \new_[70644]_ , \new_[70647]_ , \new_[70648]_ , \new_[70649]_ ,
    \new_[70652]_ , \new_[70655]_ , \new_[70656]_ , \new_[70659]_ ,
    \new_[70662]_ , \new_[70663]_ , \new_[70664]_ , \new_[70668]_ ,
    \new_[70669]_ , \new_[70672]_ , \new_[70675]_ , \new_[70676]_ ,
    \new_[70677]_ , \new_[70680]_ , \new_[70683]_ , \new_[70684]_ ,
    \new_[70687]_ , \new_[70690]_ , \new_[70691]_ , \new_[70692]_ ,
    \new_[70696]_ , \new_[70697]_ , \new_[70700]_ , \new_[70703]_ ,
    \new_[70704]_ , \new_[70705]_ , \new_[70708]_ , \new_[70711]_ ,
    \new_[70712]_ , \new_[70715]_ , \new_[70718]_ , \new_[70719]_ ,
    \new_[70720]_ , \new_[70724]_ , \new_[70725]_ , \new_[70728]_ ,
    \new_[70731]_ , \new_[70732]_ , \new_[70733]_ , \new_[70736]_ ,
    \new_[70739]_ , \new_[70740]_ , \new_[70743]_ , \new_[70746]_ ,
    \new_[70747]_ , \new_[70748]_ , \new_[70752]_ , \new_[70753]_ ,
    \new_[70756]_ , \new_[70759]_ , \new_[70760]_ , \new_[70761]_ ,
    \new_[70764]_ , \new_[70767]_ , \new_[70768]_ , \new_[70771]_ ,
    \new_[70774]_ , \new_[70775]_ , \new_[70776]_ , \new_[70780]_ ,
    \new_[70781]_ , \new_[70784]_ , \new_[70787]_ , \new_[70788]_ ,
    \new_[70789]_ , \new_[70792]_ , \new_[70795]_ , \new_[70796]_ ,
    \new_[70799]_ , \new_[70802]_ , \new_[70803]_ , \new_[70804]_ ,
    \new_[70808]_ , \new_[70809]_ , \new_[70812]_ , \new_[70815]_ ,
    \new_[70816]_ , \new_[70817]_ , \new_[70820]_ , \new_[70823]_ ,
    \new_[70824]_ , \new_[70827]_ , \new_[70830]_ , \new_[70831]_ ,
    \new_[70832]_ , \new_[70836]_ , \new_[70837]_ , \new_[70840]_ ,
    \new_[70843]_ , \new_[70844]_ , \new_[70845]_ , \new_[70848]_ ,
    \new_[70851]_ , \new_[70852]_ , \new_[70855]_ , \new_[70858]_ ,
    \new_[70859]_ , \new_[70860]_ , \new_[70864]_ , \new_[70865]_ ,
    \new_[70868]_ , \new_[70871]_ , \new_[70872]_ , \new_[70873]_ ,
    \new_[70876]_ , \new_[70879]_ , \new_[70880]_ , \new_[70883]_ ,
    \new_[70886]_ , \new_[70887]_ , \new_[70888]_ , \new_[70892]_ ,
    \new_[70893]_ , \new_[70896]_ , \new_[70899]_ , \new_[70900]_ ,
    \new_[70901]_ , \new_[70904]_ , \new_[70907]_ , \new_[70908]_ ,
    \new_[70911]_ , \new_[70914]_ , \new_[70915]_ , \new_[70916]_ ,
    \new_[70920]_ , \new_[70921]_ , \new_[70924]_ , \new_[70927]_ ,
    \new_[70928]_ , \new_[70929]_ , \new_[70932]_ , \new_[70935]_ ,
    \new_[70936]_ , \new_[70939]_ , \new_[70942]_ , \new_[70943]_ ,
    \new_[70944]_ , \new_[70948]_ , \new_[70949]_ , \new_[70952]_ ,
    \new_[70955]_ , \new_[70956]_ , \new_[70957]_ , \new_[70960]_ ,
    \new_[70963]_ , \new_[70964]_ , \new_[70967]_ , \new_[70970]_ ,
    \new_[70971]_ , \new_[70972]_ , \new_[70976]_ , \new_[70977]_ ,
    \new_[70980]_ , \new_[70983]_ , \new_[70984]_ , \new_[70985]_ ,
    \new_[70988]_ , \new_[70991]_ , \new_[70992]_ , \new_[70995]_ ,
    \new_[70998]_ , \new_[70999]_ , \new_[71000]_ , \new_[71004]_ ,
    \new_[71005]_ , \new_[71008]_ , \new_[71011]_ , \new_[71012]_ ,
    \new_[71013]_ , \new_[71016]_ , \new_[71019]_ , \new_[71020]_ ,
    \new_[71023]_ , \new_[71026]_ , \new_[71027]_ , \new_[71028]_ ,
    \new_[71032]_ , \new_[71033]_ , \new_[71036]_ , \new_[71039]_ ,
    \new_[71040]_ , \new_[71041]_ , \new_[71044]_ , \new_[71047]_ ,
    \new_[71048]_ , \new_[71051]_ , \new_[71054]_ , \new_[71055]_ ,
    \new_[71056]_ , \new_[71060]_ , \new_[71061]_ , \new_[71064]_ ,
    \new_[71067]_ , \new_[71068]_ , \new_[71069]_ , \new_[71072]_ ,
    \new_[71075]_ , \new_[71076]_ , \new_[71079]_ , \new_[71082]_ ,
    \new_[71083]_ , \new_[71084]_ , \new_[71088]_ , \new_[71089]_ ,
    \new_[71092]_ , \new_[71095]_ , \new_[71096]_ , \new_[71097]_ ,
    \new_[71100]_ , \new_[71103]_ , \new_[71104]_ , \new_[71107]_ ,
    \new_[71110]_ , \new_[71111]_ , \new_[71112]_ , \new_[71116]_ ,
    \new_[71117]_ , \new_[71120]_ , \new_[71123]_ , \new_[71124]_ ,
    \new_[71125]_ , \new_[71128]_ , \new_[71131]_ , \new_[71132]_ ,
    \new_[71135]_ , \new_[71138]_ , \new_[71139]_ , \new_[71140]_ ,
    \new_[71144]_ , \new_[71145]_ , \new_[71148]_ , \new_[71151]_ ,
    \new_[71152]_ , \new_[71153]_ , \new_[71156]_ , \new_[71159]_ ,
    \new_[71160]_ , \new_[71163]_ , \new_[71166]_ , \new_[71167]_ ,
    \new_[71168]_ , \new_[71172]_ , \new_[71173]_ , \new_[71176]_ ,
    \new_[71179]_ , \new_[71180]_ , \new_[71181]_ , \new_[71184]_ ,
    \new_[71187]_ , \new_[71188]_ , \new_[71191]_ , \new_[71194]_ ,
    \new_[71195]_ , \new_[71196]_ , \new_[71200]_ , \new_[71201]_ ,
    \new_[71204]_ , \new_[71207]_ , \new_[71208]_ , \new_[71209]_ ,
    \new_[71212]_ , \new_[71215]_ , \new_[71216]_ , \new_[71219]_ ,
    \new_[71222]_ , \new_[71223]_ , \new_[71224]_ , \new_[71228]_ ,
    \new_[71229]_ , \new_[71232]_ , \new_[71235]_ , \new_[71236]_ ,
    \new_[71237]_ , \new_[71240]_ , \new_[71243]_ , \new_[71244]_ ,
    \new_[71247]_ , \new_[71250]_ , \new_[71251]_ , \new_[71252]_ ,
    \new_[71256]_ , \new_[71257]_ , \new_[71260]_ , \new_[71263]_ ,
    \new_[71264]_ , \new_[71265]_ , \new_[71268]_ , \new_[71271]_ ,
    \new_[71272]_ , \new_[71275]_ , \new_[71278]_ , \new_[71279]_ ,
    \new_[71280]_ , \new_[71284]_ , \new_[71285]_ , \new_[71288]_ ,
    \new_[71291]_ , \new_[71292]_ , \new_[71293]_ , \new_[71296]_ ,
    \new_[71299]_ , \new_[71300]_ , \new_[71303]_ , \new_[71306]_ ,
    \new_[71307]_ , \new_[71308]_ , \new_[71312]_ , \new_[71313]_ ,
    \new_[71316]_ , \new_[71319]_ , \new_[71320]_ , \new_[71321]_ ,
    \new_[71324]_ , \new_[71327]_ , \new_[71328]_ , \new_[71331]_ ,
    \new_[71334]_ , \new_[71335]_ , \new_[71336]_ , \new_[71340]_ ,
    \new_[71341]_ , \new_[71344]_ , \new_[71347]_ , \new_[71348]_ ,
    \new_[71349]_ , \new_[71352]_ , \new_[71355]_ , \new_[71356]_ ,
    \new_[71359]_ , \new_[71362]_ , \new_[71363]_ , \new_[71364]_ ,
    \new_[71368]_ , \new_[71369]_ , \new_[71372]_ , \new_[71375]_ ,
    \new_[71376]_ , \new_[71377]_ , \new_[71380]_ , \new_[71383]_ ,
    \new_[71384]_ , \new_[71387]_ , \new_[71390]_ , \new_[71391]_ ,
    \new_[71392]_ , \new_[71396]_ , \new_[71397]_ , \new_[71400]_ ,
    \new_[71403]_ , \new_[71404]_ , \new_[71405]_ , \new_[71408]_ ,
    \new_[71411]_ , \new_[71412]_ , \new_[71415]_ , \new_[71418]_ ,
    \new_[71419]_ , \new_[71420]_ , \new_[71424]_ , \new_[71425]_ ,
    \new_[71428]_ , \new_[71431]_ , \new_[71432]_ , \new_[71433]_ ,
    \new_[71436]_ , \new_[71439]_ , \new_[71440]_ , \new_[71443]_ ,
    \new_[71446]_ , \new_[71447]_ , \new_[71448]_ , \new_[71452]_ ,
    \new_[71453]_ , \new_[71456]_ , \new_[71459]_ , \new_[71460]_ ,
    \new_[71461]_ , \new_[71464]_ , \new_[71467]_ , \new_[71468]_ ,
    \new_[71471]_ , \new_[71474]_ , \new_[71475]_ , \new_[71476]_ ,
    \new_[71480]_ , \new_[71481]_ , \new_[71484]_ , \new_[71487]_ ,
    \new_[71488]_ , \new_[71489]_ , \new_[71492]_ , \new_[71495]_ ,
    \new_[71496]_ , \new_[71499]_ , \new_[71502]_ , \new_[71503]_ ,
    \new_[71504]_ , \new_[71508]_ , \new_[71509]_ , \new_[71512]_ ,
    \new_[71515]_ , \new_[71516]_ , \new_[71517]_ , \new_[71520]_ ,
    \new_[71523]_ , \new_[71524]_ , \new_[71527]_ , \new_[71530]_ ,
    \new_[71531]_ , \new_[71532]_ , \new_[71536]_ , \new_[71537]_ ,
    \new_[71540]_ , \new_[71543]_ , \new_[71544]_ , \new_[71545]_ ,
    \new_[71548]_ , \new_[71551]_ , \new_[71552]_ , \new_[71555]_ ,
    \new_[71558]_ , \new_[71559]_ , \new_[71560]_ , \new_[71564]_ ,
    \new_[71565]_ , \new_[71568]_ , \new_[71571]_ , \new_[71572]_ ,
    \new_[71573]_ , \new_[71576]_ , \new_[71579]_ , \new_[71580]_ ,
    \new_[71583]_ , \new_[71586]_ , \new_[71587]_ , \new_[71588]_ ,
    \new_[71592]_ , \new_[71593]_ , \new_[71596]_ , \new_[71599]_ ,
    \new_[71600]_ , \new_[71601]_ , \new_[71604]_ , \new_[71607]_ ,
    \new_[71608]_ , \new_[71611]_ , \new_[71614]_ , \new_[71615]_ ,
    \new_[71616]_ , \new_[71620]_ , \new_[71621]_ , \new_[71624]_ ,
    \new_[71627]_ , \new_[71628]_ , \new_[71629]_ , \new_[71632]_ ,
    \new_[71635]_ , \new_[71636]_ , \new_[71639]_ , \new_[71642]_ ,
    \new_[71643]_ , \new_[71644]_ , \new_[71648]_ , \new_[71649]_ ,
    \new_[71652]_ , \new_[71655]_ , \new_[71656]_ , \new_[71657]_ ,
    \new_[71660]_ , \new_[71663]_ , \new_[71664]_ , \new_[71667]_ ,
    \new_[71670]_ , \new_[71671]_ , \new_[71672]_ , \new_[71676]_ ,
    \new_[71677]_ , \new_[71680]_ , \new_[71683]_ , \new_[71684]_ ,
    \new_[71685]_ , \new_[71688]_ , \new_[71691]_ , \new_[71692]_ ,
    \new_[71695]_ , \new_[71698]_ , \new_[71699]_ , \new_[71700]_ ,
    \new_[71704]_ , \new_[71705]_ , \new_[71708]_ , \new_[71711]_ ,
    \new_[71712]_ , \new_[71713]_ , \new_[71716]_ , \new_[71719]_ ,
    \new_[71720]_ , \new_[71723]_ , \new_[71726]_ , \new_[71727]_ ,
    \new_[71728]_ , \new_[71732]_ , \new_[71733]_ , \new_[71736]_ ,
    \new_[71739]_ , \new_[71740]_ , \new_[71741]_ , \new_[71744]_ ,
    \new_[71747]_ , \new_[71748]_ , \new_[71751]_ , \new_[71754]_ ,
    \new_[71755]_ , \new_[71756]_ , \new_[71760]_ , \new_[71761]_ ,
    \new_[71764]_ , \new_[71767]_ , \new_[71768]_ , \new_[71769]_ ,
    \new_[71772]_ , \new_[71775]_ , \new_[71776]_ , \new_[71779]_ ,
    \new_[71782]_ , \new_[71783]_ , \new_[71784]_ , \new_[71788]_ ,
    \new_[71789]_ , \new_[71792]_ , \new_[71795]_ , \new_[71796]_ ,
    \new_[71797]_ , \new_[71800]_ , \new_[71803]_ , \new_[71804]_ ,
    \new_[71807]_ , \new_[71810]_ , \new_[71811]_ , \new_[71812]_ ,
    \new_[71816]_ , \new_[71817]_ , \new_[71820]_ , \new_[71823]_ ,
    \new_[71824]_ , \new_[71825]_ , \new_[71828]_ , \new_[71831]_ ,
    \new_[71832]_ , \new_[71835]_ , \new_[71838]_ , \new_[71839]_ ,
    \new_[71840]_ , \new_[71844]_ , \new_[71845]_ , \new_[71848]_ ,
    \new_[71851]_ , \new_[71852]_ , \new_[71853]_ , \new_[71856]_ ,
    \new_[71859]_ , \new_[71860]_ , \new_[71863]_ , \new_[71866]_ ,
    \new_[71867]_ , \new_[71868]_ , \new_[71872]_ , \new_[71873]_ ,
    \new_[71876]_ , \new_[71879]_ , \new_[71880]_ , \new_[71881]_ ,
    \new_[71884]_ , \new_[71887]_ , \new_[71888]_ , \new_[71891]_ ,
    \new_[71894]_ , \new_[71895]_ , \new_[71896]_ , \new_[71900]_ ,
    \new_[71901]_ , \new_[71904]_ , \new_[71907]_ , \new_[71908]_ ,
    \new_[71909]_ , \new_[71912]_ , \new_[71915]_ , \new_[71916]_ ,
    \new_[71919]_ , \new_[71922]_ , \new_[71923]_ , \new_[71924]_ ,
    \new_[71928]_ , \new_[71929]_ , \new_[71932]_ , \new_[71935]_ ,
    \new_[71936]_ , \new_[71937]_ , \new_[71940]_ , \new_[71943]_ ,
    \new_[71944]_ , \new_[71947]_ , \new_[71950]_ , \new_[71951]_ ,
    \new_[71952]_ , \new_[71956]_ , \new_[71957]_ , \new_[71960]_ ,
    \new_[71963]_ , \new_[71964]_ , \new_[71965]_ , \new_[71968]_ ,
    \new_[71971]_ , \new_[71972]_ , \new_[71975]_ , \new_[71978]_ ,
    \new_[71979]_ , \new_[71980]_ , \new_[71984]_ , \new_[71985]_ ,
    \new_[71988]_ , \new_[71991]_ , \new_[71992]_ , \new_[71993]_ ,
    \new_[71996]_ , \new_[71999]_ , \new_[72000]_ , \new_[72003]_ ,
    \new_[72006]_ , \new_[72007]_ , \new_[72008]_ , \new_[72012]_ ,
    \new_[72013]_ , \new_[72016]_ , \new_[72019]_ , \new_[72020]_ ,
    \new_[72021]_ , \new_[72024]_ , \new_[72027]_ , \new_[72028]_ ,
    \new_[72031]_ , \new_[72034]_ , \new_[72035]_ , \new_[72036]_ ,
    \new_[72040]_ , \new_[72041]_ , \new_[72044]_ , \new_[72047]_ ,
    \new_[72048]_ , \new_[72049]_ , \new_[72052]_ , \new_[72055]_ ,
    \new_[72056]_ , \new_[72059]_ , \new_[72062]_ , \new_[72063]_ ,
    \new_[72064]_ , \new_[72068]_ , \new_[72069]_ , \new_[72072]_ ,
    \new_[72075]_ , \new_[72076]_ , \new_[72077]_ , \new_[72080]_ ,
    \new_[72083]_ , \new_[72084]_ , \new_[72087]_ , \new_[72090]_ ,
    \new_[72091]_ , \new_[72092]_ , \new_[72096]_ , \new_[72097]_ ,
    \new_[72100]_ , \new_[72103]_ , \new_[72104]_ , \new_[72105]_ ,
    \new_[72108]_ , \new_[72111]_ , \new_[72112]_ , \new_[72115]_ ,
    \new_[72118]_ , \new_[72119]_ , \new_[72120]_ , \new_[72124]_ ,
    \new_[72125]_ , \new_[72128]_ , \new_[72131]_ , \new_[72132]_ ,
    \new_[72133]_ , \new_[72136]_ , \new_[72139]_ , \new_[72140]_ ,
    \new_[72143]_ , \new_[72146]_ , \new_[72147]_ , \new_[72148]_ ,
    \new_[72152]_ , \new_[72153]_ , \new_[72156]_ , \new_[72159]_ ,
    \new_[72160]_ , \new_[72161]_ , \new_[72164]_ , \new_[72167]_ ,
    \new_[72168]_ , \new_[72171]_ , \new_[72174]_ , \new_[72175]_ ,
    \new_[72176]_ , \new_[72180]_ , \new_[72181]_ , \new_[72184]_ ,
    \new_[72187]_ , \new_[72188]_ , \new_[72189]_ , \new_[72192]_ ,
    \new_[72195]_ , \new_[72196]_ , \new_[72199]_ , \new_[72202]_ ,
    \new_[72203]_ , \new_[72204]_ , \new_[72208]_ , \new_[72209]_ ,
    \new_[72212]_ , \new_[72215]_ , \new_[72216]_ , \new_[72217]_ ,
    \new_[72220]_ , \new_[72223]_ , \new_[72224]_ , \new_[72227]_ ,
    \new_[72230]_ , \new_[72231]_ , \new_[72232]_ , \new_[72236]_ ,
    \new_[72237]_ , \new_[72240]_ , \new_[72243]_ , \new_[72244]_ ,
    \new_[72245]_ , \new_[72248]_ , \new_[72251]_ , \new_[72252]_ ,
    \new_[72255]_ , \new_[72258]_ , \new_[72259]_ , \new_[72260]_ ,
    \new_[72264]_ , \new_[72265]_ , \new_[72268]_ , \new_[72271]_ ,
    \new_[72272]_ , \new_[72273]_ , \new_[72276]_ , \new_[72279]_ ,
    \new_[72280]_ , \new_[72283]_ , \new_[72286]_ , \new_[72287]_ ,
    \new_[72288]_ , \new_[72292]_ , \new_[72293]_ , \new_[72296]_ ,
    \new_[72299]_ , \new_[72300]_ , \new_[72301]_ , \new_[72304]_ ,
    \new_[72307]_ , \new_[72308]_ , \new_[72311]_ , \new_[72314]_ ,
    \new_[72315]_ , \new_[72316]_ , \new_[72320]_ , \new_[72321]_ ,
    \new_[72324]_ , \new_[72327]_ , \new_[72328]_ , \new_[72329]_ ,
    \new_[72332]_ , \new_[72335]_ , \new_[72336]_ , \new_[72339]_ ,
    \new_[72342]_ , \new_[72343]_ , \new_[72344]_ , \new_[72348]_ ,
    \new_[72349]_ , \new_[72352]_ , \new_[72355]_ , \new_[72356]_ ,
    \new_[72357]_ , \new_[72360]_ , \new_[72363]_ , \new_[72364]_ ,
    \new_[72367]_ , \new_[72370]_ , \new_[72371]_ , \new_[72372]_ ,
    \new_[72376]_ , \new_[72377]_ , \new_[72380]_ , \new_[72383]_ ,
    \new_[72384]_ , \new_[72385]_ , \new_[72388]_ , \new_[72391]_ ,
    \new_[72392]_ , \new_[72395]_ , \new_[72398]_ , \new_[72399]_ ,
    \new_[72400]_ , \new_[72404]_ , \new_[72405]_ , \new_[72408]_ ,
    \new_[72411]_ , \new_[72412]_ , \new_[72413]_ , \new_[72416]_ ,
    \new_[72419]_ , \new_[72420]_ , \new_[72423]_ , \new_[72426]_ ,
    \new_[72427]_ , \new_[72428]_ , \new_[72432]_ , \new_[72433]_ ,
    \new_[72436]_ , \new_[72439]_ , \new_[72440]_ , \new_[72441]_ ,
    \new_[72444]_ , \new_[72447]_ , \new_[72448]_ , \new_[72451]_ ,
    \new_[72454]_ , \new_[72455]_ , \new_[72456]_ , \new_[72460]_ ,
    \new_[72461]_ , \new_[72464]_ , \new_[72467]_ , \new_[72468]_ ,
    \new_[72469]_ , \new_[72472]_ , \new_[72475]_ , \new_[72476]_ ,
    \new_[72479]_ , \new_[72482]_ , \new_[72483]_ , \new_[72484]_ ,
    \new_[72488]_ , \new_[72489]_ , \new_[72492]_ , \new_[72495]_ ,
    \new_[72496]_ , \new_[72497]_ , \new_[72500]_ , \new_[72503]_ ,
    \new_[72504]_ , \new_[72507]_ , \new_[72510]_ , \new_[72511]_ ,
    \new_[72512]_ , \new_[72516]_ , \new_[72517]_ , \new_[72520]_ ,
    \new_[72523]_ , \new_[72524]_ , \new_[72525]_ , \new_[72528]_ ,
    \new_[72531]_ , \new_[72532]_ , \new_[72535]_ , \new_[72538]_ ,
    \new_[72539]_ , \new_[72540]_ , \new_[72544]_ , \new_[72545]_ ,
    \new_[72548]_ , \new_[72551]_ , \new_[72552]_ , \new_[72553]_ ,
    \new_[72556]_ , \new_[72559]_ , \new_[72560]_ , \new_[72563]_ ,
    \new_[72566]_ , \new_[72567]_ , \new_[72568]_ , \new_[72572]_ ,
    \new_[72573]_ , \new_[72576]_ , \new_[72579]_ , \new_[72580]_ ,
    \new_[72581]_ , \new_[72584]_ , \new_[72587]_ , \new_[72588]_ ,
    \new_[72591]_ , \new_[72594]_ , \new_[72595]_ , \new_[72596]_ ,
    \new_[72600]_ , \new_[72601]_ , \new_[72604]_ , \new_[72607]_ ,
    \new_[72608]_ , \new_[72609]_ , \new_[72612]_ , \new_[72615]_ ,
    \new_[72616]_ , \new_[72619]_ , \new_[72622]_ , \new_[72623]_ ,
    \new_[72624]_ , \new_[72628]_ , \new_[72629]_ , \new_[72632]_ ,
    \new_[72635]_ , \new_[72636]_ , \new_[72637]_ , \new_[72640]_ ,
    \new_[72643]_ , \new_[72644]_ , \new_[72647]_ , \new_[72650]_ ,
    \new_[72651]_ , \new_[72652]_ , \new_[72656]_ , \new_[72657]_ ,
    \new_[72660]_ , \new_[72663]_ , \new_[72664]_ , \new_[72665]_ ,
    \new_[72668]_ , \new_[72671]_ , \new_[72672]_ , \new_[72675]_ ,
    \new_[72678]_ , \new_[72679]_ , \new_[72680]_ , \new_[72684]_ ,
    \new_[72685]_ , \new_[72688]_ , \new_[72691]_ , \new_[72692]_ ,
    \new_[72693]_ , \new_[72696]_ , \new_[72699]_ , \new_[72700]_ ,
    \new_[72703]_ , \new_[72706]_ , \new_[72707]_ , \new_[72708]_ ,
    \new_[72712]_ , \new_[72713]_ , \new_[72716]_ , \new_[72719]_ ,
    \new_[72720]_ , \new_[72721]_ , \new_[72724]_ , \new_[72727]_ ,
    \new_[72728]_ , \new_[72731]_ , \new_[72734]_ , \new_[72735]_ ,
    \new_[72736]_ , \new_[72740]_ , \new_[72741]_ , \new_[72744]_ ,
    \new_[72747]_ , \new_[72748]_ , \new_[72749]_ , \new_[72752]_ ,
    \new_[72755]_ , \new_[72756]_ , \new_[72759]_ , \new_[72762]_ ,
    \new_[72763]_ , \new_[72764]_ , \new_[72768]_ , \new_[72769]_ ,
    \new_[72772]_ , \new_[72775]_ , \new_[72776]_ , \new_[72777]_ ,
    \new_[72780]_ , \new_[72783]_ , \new_[72784]_ , \new_[72787]_ ,
    \new_[72790]_ , \new_[72791]_ , \new_[72792]_ , \new_[72796]_ ,
    \new_[72797]_ , \new_[72800]_ , \new_[72803]_ , \new_[72804]_ ,
    \new_[72805]_ , \new_[72808]_ , \new_[72811]_ , \new_[72812]_ ,
    \new_[72815]_ , \new_[72818]_ , \new_[72819]_ , \new_[72820]_ ,
    \new_[72824]_ , \new_[72825]_ , \new_[72828]_ , \new_[72831]_ ,
    \new_[72832]_ , \new_[72833]_ , \new_[72836]_ , \new_[72839]_ ,
    \new_[72840]_ , \new_[72843]_ , \new_[72846]_ , \new_[72847]_ ,
    \new_[72848]_ , \new_[72852]_ , \new_[72853]_ , \new_[72856]_ ,
    \new_[72859]_ , \new_[72860]_ , \new_[72861]_ , \new_[72864]_ ,
    \new_[72867]_ , \new_[72868]_ , \new_[72871]_ , \new_[72874]_ ,
    \new_[72875]_ , \new_[72876]_ , \new_[72880]_ , \new_[72881]_ ,
    \new_[72884]_ , \new_[72887]_ , \new_[72888]_ , \new_[72889]_ ,
    \new_[72892]_ , \new_[72895]_ , \new_[72896]_ , \new_[72899]_ ,
    \new_[72902]_ , \new_[72903]_ , \new_[72904]_ , \new_[72908]_ ,
    \new_[72909]_ , \new_[72912]_ , \new_[72915]_ , \new_[72916]_ ,
    \new_[72917]_ , \new_[72920]_ , \new_[72923]_ , \new_[72924]_ ,
    \new_[72927]_ , \new_[72930]_ , \new_[72931]_ , \new_[72932]_ ,
    \new_[72936]_ , \new_[72937]_ , \new_[72940]_ , \new_[72943]_ ,
    \new_[72944]_ , \new_[72945]_ , \new_[72948]_ , \new_[72951]_ ,
    \new_[72952]_ , \new_[72955]_ , \new_[72958]_ , \new_[72959]_ ,
    \new_[72960]_ , \new_[72964]_ , \new_[72965]_ , \new_[72968]_ ,
    \new_[72971]_ , \new_[72972]_ , \new_[72973]_ , \new_[72976]_ ,
    \new_[72979]_ , \new_[72980]_ , \new_[72983]_ , \new_[72986]_ ,
    \new_[72987]_ , \new_[72988]_ , \new_[72992]_ , \new_[72993]_ ,
    \new_[72996]_ , \new_[72999]_ , \new_[73000]_ , \new_[73001]_ ,
    \new_[73004]_ , \new_[73007]_ , \new_[73008]_ , \new_[73011]_ ,
    \new_[73014]_ , \new_[73015]_ , \new_[73016]_ , \new_[73020]_ ,
    \new_[73021]_ , \new_[73024]_ , \new_[73027]_ , \new_[73028]_ ,
    \new_[73029]_ , \new_[73032]_ , \new_[73035]_ , \new_[73036]_ ,
    \new_[73039]_ , \new_[73042]_ , \new_[73043]_ , \new_[73044]_ ,
    \new_[73048]_ , \new_[73049]_ , \new_[73052]_ , \new_[73055]_ ,
    \new_[73056]_ , \new_[73057]_ , \new_[73060]_ , \new_[73063]_ ,
    \new_[73064]_ , \new_[73067]_ , \new_[73070]_ , \new_[73071]_ ,
    \new_[73072]_ , \new_[73076]_ , \new_[73077]_ , \new_[73080]_ ,
    \new_[73083]_ , \new_[73084]_ , \new_[73085]_ , \new_[73088]_ ,
    \new_[73091]_ , \new_[73092]_ , \new_[73095]_ , \new_[73098]_ ,
    \new_[73099]_ , \new_[73100]_ , \new_[73104]_ , \new_[73105]_ ,
    \new_[73108]_ , \new_[73111]_ , \new_[73112]_ , \new_[73113]_ ,
    \new_[73116]_ , \new_[73119]_ , \new_[73120]_ , \new_[73123]_ ,
    \new_[73126]_ , \new_[73127]_ , \new_[73128]_ , \new_[73132]_ ,
    \new_[73133]_ , \new_[73136]_ , \new_[73139]_ , \new_[73140]_ ,
    \new_[73141]_ , \new_[73144]_ , \new_[73147]_ , \new_[73148]_ ,
    \new_[73151]_ , \new_[73154]_ , \new_[73155]_ , \new_[73156]_ ,
    \new_[73160]_ , \new_[73161]_ , \new_[73164]_ , \new_[73167]_ ,
    \new_[73168]_ , \new_[73169]_ , \new_[73172]_ , \new_[73175]_ ,
    \new_[73176]_ , \new_[73179]_ , \new_[73182]_ , \new_[73183]_ ,
    \new_[73184]_ , \new_[73188]_ , \new_[73189]_ , \new_[73192]_ ,
    \new_[73195]_ , \new_[73196]_ , \new_[73197]_ , \new_[73200]_ ,
    \new_[73203]_ , \new_[73204]_ , \new_[73207]_ , \new_[73210]_ ,
    \new_[73211]_ , \new_[73212]_ , \new_[73216]_ , \new_[73217]_ ,
    \new_[73220]_ , \new_[73223]_ , \new_[73224]_ , \new_[73225]_ ,
    \new_[73228]_ , \new_[73231]_ , \new_[73232]_ , \new_[73235]_ ,
    \new_[73238]_ , \new_[73239]_ , \new_[73240]_ , \new_[73244]_ ,
    \new_[73245]_ , \new_[73248]_ , \new_[73251]_ , \new_[73252]_ ,
    \new_[73253]_ , \new_[73256]_ , \new_[73259]_ , \new_[73260]_ ,
    \new_[73263]_ , \new_[73266]_ , \new_[73267]_ , \new_[73268]_ ,
    \new_[73272]_ , \new_[73273]_ , \new_[73276]_ , \new_[73279]_ ,
    \new_[73280]_ , \new_[73281]_ , \new_[73284]_ , \new_[73287]_ ,
    \new_[73288]_ , \new_[73291]_ , \new_[73294]_ , \new_[73295]_ ,
    \new_[73296]_ , \new_[73300]_ , \new_[73301]_ , \new_[73304]_ ,
    \new_[73307]_ , \new_[73308]_ , \new_[73309]_ , \new_[73312]_ ,
    \new_[73315]_ , \new_[73316]_ , \new_[73319]_ , \new_[73322]_ ,
    \new_[73323]_ , \new_[73324]_ , \new_[73328]_ , \new_[73329]_ ,
    \new_[73332]_ , \new_[73335]_ , \new_[73336]_ , \new_[73337]_ ,
    \new_[73340]_ , \new_[73343]_ , \new_[73344]_ , \new_[73347]_ ,
    \new_[73350]_ , \new_[73351]_ , \new_[73352]_ , \new_[73356]_ ,
    \new_[73357]_ , \new_[73360]_ , \new_[73363]_ , \new_[73364]_ ,
    \new_[73365]_ , \new_[73368]_ , \new_[73371]_ , \new_[73372]_ ,
    \new_[73375]_ , \new_[73378]_ , \new_[73379]_ , \new_[73380]_ ,
    \new_[73384]_ , \new_[73385]_ , \new_[73388]_ , \new_[73391]_ ,
    \new_[73392]_ , \new_[73393]_ , \new_[73396]_ , \new_[73399]_ ,
    \new_[73400]_ , \new_[73403]_ , \new_[73406]_ , \new_[73407]_ ,
    \new_[73408]_ , \new_[73412]_ , \new_[73413]_ , \new_[73416]_ ,
    \new_[73419]_ , \new_[73420]_ , \new_[73421]_ , \new_[73424]_ ,
    \new_[73427]_ , \new_[73428]_ , \new_[73431]_ , \new_[73434]_ ,
    \new_[73435]_ , \new_[73436]_ , \new_[73440]_ , \new_[73441]_ ,
    \new_[73444]_ , \new_[73447]_ , \new_[73448]_ , \new_[73449]_ ,
    \new_[73452]_ , \new_[73455]_ , \new_[73456]_ , \new_[73459]_ ,
    \new_[73462]_ , \new_[73463]_ , \new_[73464]_ , \new_[73468]_ ,
    \new_[73469]_ , \new_[73472]_ , \new_[73475]_ , \new_[73476]_ ,
    \new_[73477]_ , \new_[73480]_ , \new_[73483]_ , \new_[73484]_ ,
    \new_[73487]_ , \new_[73490]_ , \new_[73491]_ , \new_[73492]_ ,
    \new_[73496]_ , \new_[73497]_ , \new_[73500]_ , \new_[73503]_ ,
    \new_[73504]_ , \new_[73505]_ , \new_[73508]_ , \new_[73511]_ ,
    \new_[73512]_ , \new_[73515]_ , \new_[73518]_ , \new_[73519]_ ,
    \new_[73520]_ , \new_[73524]_ , \new_[73525]_ , \new_[73528]_ ,
    \new_[73531]_ , \new_[73532]_ , \new_[73533]_ , \new_[73536]_ ,
    \new_[73539]_ , \new_[73540]_ , \new_[73543]_ , \new_[73546]_ ,
    \new_[73547]_ , \new_[73548]_ , \new_[73552]_ , \new_[73553]_ ,
    \new_[73556]_ , \new_[73559]_ , \new_[73560]_ , \new_[73561]_ ,
    \new_[73564]_ , \new_[73567]_ , \new_[73568]_ , \new_[73571]_ ,
    \new_[73574]_ , \new_[73575]_ , \new_[73576]_ , \new_[73580]_ ,
    \new_[73581]_ , \new_[73584]_ , \new_[73587]_ , \new_[73588]_ ,
    \new_[73589]_ , \new_[73592]_ , \new_[73595]_ , \new_[73596]_ ,
    \new_[73599]_ , \new_[73602]_ , \new_[73603]_ , \new_[73604]_ ,
    \new_[73608]_ , \new_[73609]_ , \new_[73612]_ , \new_[73615]_ ,
    \new_[73616]_ , \new_[73617]_ , \new_[73620]_ , \new_[73623]_ ,
    \new_[73624]_ , \new_[73627]_ , \new_[73630]_ , \new_[73631]_ ,
    \new_[73632]_ , \new_[73636]_ , \new_[73637]_ , \new_[73640]_ ,
    \new_[73643]_ , \new_[73644]_ , \new_[73645]_ , \new_[73648]_ ,
    \new_[73651]_ , \new_[73652]_ , \new_[73655]_ , \new_[73658]_ ,
    \new_[73659]_ , \new_[73660]_ , \new_[73664]_ , \new_[73665]_ ,
    \new_[73668]_ , \new_[73671]_ , \new_[73672]_ , \new_[73673]_ ,
    \new_[73676]_ , \new_[73679]_ , \new_[73680]_ , \new_[73683]_ ,
    \new_[73686]_ , \new_[73687]_ , \new_[73688]_ , \new_[73692]_ ,
    \new_[73693]_ , \new_[73696]_ , \new_[73699]_ , \new_[73700]_ ,
    \new_[73701]_ , \new_[73704]_ , \new_[73707]_ , \new_[73708]_ ,
    \new_[73711]_ , \new_[73714]_ , \new_[73715]_ , \new_[73716]_ ,
    \new_[73720]_ , \new_[73721]_ , \new_[73724]_ , \new_[73727]_ ,
    \new_[73728]_ , \new_[73729]_ , \new_[73732]_ , \new_[73735]_ ,
    \new_[73736]_ , \new_[73739]_ , \new_[73742]_ , \new_[73743]_ ,
    \new_[73744]_ , \new_[73748]_ , \new_[73749]_ , \new_[73752]_ ,
    \new_[73755]_ , \new_[73756]_ , \new_[73757]_ , \new_[73760]_ ,
    \new_[73763]_ , \new_[73764]_ , \new_[73767]_ , \new_[73770]_ ,
    \new_[73771]_ , \new_[73772]_ , \new_[73776]_ , \new_[73777]_ ,
    \new_[73780]_ , \new_[73783]_ , \new_[73784]_ , \new_[73785]_ ,
    \new_[73788]_ , \new_[73791]_ , \new_[73792]_ , \new_[73795]_ ,
    \new_[73798]_ , \new_[73799]_ , \new_[73800]_ , \new_[73804]_ ,
    \new_[73805]_ , \new_[73808]_ , \new_[73811]_ , \new_[73812]_ ,
    \new_[73813]_ , \new_[73816]_ , \new_[73819]_ , \new_[73820]_ ,
    \new_[73823]_ , \new_[73826]_ , \new_[73827]_ , \new_[73828]_ ,
    \new_[73832]_ , \new_[73833]_ , \new_[73836]_ , \new_[73839]_ ,
    \new_[73840]_ , \new_[73841]_ , \new_[73844]_ , \new_[73847]_ ,
    \new_[73848]_ , \new_[73851]_ , \new_[73854]_ , \new_[73855]_ ,
    \new_[73856]_ , \new_[73860]_ , \new_[73861]_ , \new_[73864]_ ,
    \new_[73867]_ , \new_[73868]_ , \new_[73869]_ , \new_[73872]_ ,
    \new_[73875]_ , \new_[73876]_ , \new_[73879]_ , \new_[73882]_ ,
    \new_[73883]_ , \new_[73884]_ , \new_[73888]_ , \new_[73889]_ ,
    \new_[73892]_ , \new_[73895]_ , \new_[73896]_ , \new_[73897]_ ,
    \new_[73900]_ , \new_[73903]_ , \new_[73904]_ , \new_[73907]_ ,
    \new_[73910]_ , \new_[73911]_ , \new_[73912]_ , \new_[73916]_ ,
    \new_[73917]_ , \new_[73920]_ , \new_[73923]_ , \new_[73924]_ ,
    \new_[73925]_ , \new_[73928]_ , \new_[73931]_ , \new_[73932]_ ,
    \new_[73935]_ , \new_[73938]_ , \new_[73939]_ , \new_[73940]_ ,
    \new_[73944]_ , \new_[73945]_ , \new_[73948]_ , \new_[73951]_ ,
    \new_[73952]_ , \new_[73953]_ , \new_[73956]_ , \new_[73959]_ ,
    \new_[73960]_ , \new_[73963]_ , \new_[73966]_ , \new_[73967]_ ,
    \new_[73968]_ , \new_[73972]_ , \new_[73973]_ , \new_[73976]_ ,
    \new_[73979]_ , \new_[73980]_ , \new_[73981]_ , \new_[73984]_ ,
    \new_[73987]_ , \new_[73988]_ , \new_[73991]_ , \new_[73994]_ ,
    \new_[73995]_ , \new_[73996]_ , \new_[74000]_ , \new_[74001]_ ,
    \new_[74004]_ , \new_[74007]_ , \new_[74008]_ , \new_[74009]_ ,
    \new_[74012]_ , \new_[74015]_ , \new_[74016]_ , \new_[74019]_ ,
    \new_[74022]_ , \new_[74023]_ , \new_[74024]_ , \new_[74028]_ ,
    \new_[74029]_ , \new_[74032]_ , \new_[74035]_ , \new_[74036]_ ,
    \new_[74037]_ , \new_[74040]_ , \new_[74043]_ , \new_[74044]_ ,
    \new_[74047]_ , \new_[74050]_ , \new_[74051]_ , \new_[74052]_ ,
    \new_[74056]_ , \new_[74057]_ , \new_[74060]_ , \new_[74063]_ ,
    \new_[74064]_ , \new_[74065]_ , \new_[74068]_ , \new_[74071]_ ,
    \new_[74072]_ , \new_[74075]_ , \new_[74078]_ , \new_[74079]_ ,
    \new_[74080]_ , \new_[74084]_ , \new_[74085]_ , \new_[74088]_ ,
    \new_[74091]_ , \new_[74092]_ , \new_[74093]_ , \new_[74096]_ ,
    \new_[74099]_ , \new_[74100]_ , \new_[74103]_ , \new_[74106]_ ,
    \new_[74107]_ , \new_[74108]_ , \new_[74112]_ , \new_[74113]_ ,
    \new_[74116]_ , \new_[74119]_ , \new_[74120]_ , \new_[74121]_ ,
    \new_[74124]_ , \new_[74127]_ , \new_[74128]_ , \new_[74131]_ ,
    \new_[74134]_ , \new_[74135]_ , \new_[74136]_ , \new_[74140]_ ,
    \new_[74141]_ , \new_[74144]_ , \new_[74147]_ , \new_[74148]_ ,
    \new_[74149]_ , \new_[74152]_ , \new_[74155]_ , \new_[74156]_ ,
    \new_[74159]_ , \new_[74162]_ , \new_[74163]_ , \new_[74164]_ ,
    \new_[74168]_ , \new_[74169]_ , \new_[74172]_ , \new_[74175]_ ,
    \new_[74176]_ , \new_[74177]_ , \new_[74180]_ , \new_[74183]_ ,
    \new_[74184]_ , \new_[74187]_ , \new_[74190]_ , \new_[74191]_ ,
    \new_[74192]_ , \new_[74196]_ , \new_[74197]_ , \new_[74200]_ ,
    \new_[74203]_ , \new_[74204]_ , \new_[74205]_ , \new_[74208]_ ,
    \new_[74211]_ , \new_[74212]_ , \new_[74215]_ , \new_[74218]_ ,
    \new_[74219]_ , \new_[74220]_ , \new_[74224]_ , \new_[74225]_ ,
    \new_[74228]_ , \new_[74231]_ , \new_[74232]_ , \new_[74233]_ ,
    \new_[74236]_ , \new_[74239]_ , \new_[74240]_ , \new_[74243]_ ,
    \new_[74246]_ , \new_[74247]_ , \new_[74248]_ , \new_[74252]_ ,
    \new_[74253]_ , \new_[74256]_ , \new_[74259]_ , \new_[74260]_ ,
    \new_[74261]_ , \new_[74264]_ , \new_[74267]_ , \new_[74268]_ ,
    \new_[74271]_ , \new_[74274]_ , \new_[74275]_ , \new_[74276]_ ,
    \new_[74280]_ , \new_[74281]_ , \new_[74284]_ , \new_[74287]_ ,
    \new_[74288]_ , \new_[74289]_ , \new_[74292]_ , \new_[74295]_ ,
    \new_[74296]_ , \new_[74299]_ , \new_[74302]_ , \new_[74303]_ ,
    \new_[74304]_ , \new_[74308]_ , \new_[74309]_ , \new_[74312]_ ,
    \new_[74315]_ , \new_[74316]_ , \new_[74317]_ , \new_[74320]_ ,
    \new_[74323]_ , \new_[74324]_ , \new_[74327]_ , \new_[74330]_ ,
    \new_[74331]_ , \new_[74332]_ , \new_[74336]_ , \new_[74337]_ ,
    \new_[74340]_ , \new_[74343]_ , \new_[74344]_ , \new_[74345]_ ,
    \new_[74348]_ , \new_[74351]_ , \new_[74352]_ , \new_[74355]_ ,
    \new_[74358]_ , \new_[74359]_ , \new_[74360]_ , \new_[74364]_ ,
    \new_[74365]_ , \new_[74368]_ , \new_[74371]_ , \new_[74372]_ ,
    \new_[74373]_ , \new_[74376]_ , \new_[74379]_ , \new_[74380]_ ,
    \new_[74383]_ , \new_[74386]_ , \new_[74387]_ , \new_[74388]_ ,
    \new_[74392]_ , \new_[74393]_ , \new_[74396]_ , \new_[74399]_ ,
    \new_[74400]_ , \new_[74401]_ , \new_[74404]_ , \new_[74407]_ ,
    \new_[74408]_ , \new_[74411]_ , \new_[74414]_ , \new_[74415]_ ,
    \new_[74416]_ , \new_[74420]_ , \new_[74421]_ , \new_[74424]_ ,
    \new_[74427]_ , \new_[74428]_ , \new_[74429]_ , \new_[74432]_ ,
    \new_[74435]_ , \new_[74436]_ , \new_[74439]_ , \new_[74442]_ ,
    \new_[74443]_ , \new_[74444]_ , \new_[74448]_ , \new_[74449]_ ,
    \new_[74452]_ , \new_[74455]_ , \new_[74456]_ , \new_[74457]_ ,
    \new_[74460]_ , \new_[74463]_ , \new_[74464]_ , \new_[74467]_ ,
    \new_[74470]_ , \new_[74471]_ , \new_[74472]_ , \new_[74476]_ ,
    \new_[74477]_ , \new_[74480]_ , \new_[74483]_ , \new_[74484]_ ,
    \new_[74485]_ , \new_[74488]_ , \new_[74491]_ , \new_[74492]_ ,
    \new_[74495]_ , \new_[74498]_ , \new_[74499]_ , \new_[74500]_ ,
    \new_[74504]_ , \new_[74505]_ , \new_[74508]_ , \new_[74511]_ ,
    \new_[74512]_ , \new_[74513]_ , \new_[74516]_ , \new_[74519]_ ,
    \new_[74520]_ , \new_[74523]_ , \new_[74526]_ , \new_[74527]_ ,
    \new_[74528]_ , \new_[74532]_ , \new_[74533]_ , \new_[74536]_ ,
    \new_[74539]_ , \new_[74540]_ , \new_[74541]_ , \new_[74544]_ ,
    \new_[74547]_ , \new_[74548]_ , \new_[74551]_ , \new_[74554]_ ,
    \new_[74555]_ , \new_[74556]_ , \new_[74560]_ , \new_[74561]_ ,
    \new_[74564]_ , \new_[74567]_ , \new_[74568]_ , \new_[74569]_ ,
    \new_[74572]_ , \new_[74575]_ , \new_[74576]_ , \new_[74579]_ ,
    \new_[74582]_ , \new_[74583]_ , \new_[74584]_ , \new_[74588]_ ,
    \new_[74589]_ , \new_[74592]_ , \new_[74595]_ , \new_[74596]_ ,
    \new_[74597]_ , \new_[74600]_ , \new_[74603]_ , \new_[74604]_ ,
    \new_[74607]_ , \new_[74610]_ , \new_[74611]_ , \new_[74612]_ ,
    \new_[74616]_ , \new_[74617]_ , \new_[74620]_ , \new_[74623]_ ,
    \new_[74624]_ , \new_[74625]_ , \new_[74628]_ , \new_[74631]_ ,
    \new_[74632]_ , \new_[74635]_ , \new_[74638]_ , \new_[74639]_ ,
    \new_[74640]_ , \new_[74644]_ , \new_[74645]_ , \new_[74648]_ ,
    \new_[74651]_ , \new_[74652]_ , \new_[74653]_ , \new_[74656]_ ,
    \new_[74659]_ , \new_[74660]_ , \new_[74663]_ , \new_[74666]_ ,
    \new_[74667]_ , \new_[74668]_ , \new_[74672]_ , \new_[74673]_ ,
    \new_[74676]_ , \new_[74679]_ , \new_[74680]_ , \new_[74681]_ ,
    \new_[74684]_ , \new_[74687]_ , \new_[74688]_ , \new_[74691]_ ,
    \new_[74694]_ , \new_[74695]_ , \new_[74696]_ , \new_[74700]_ ,
    \new_[74701]_ , \new_[74704]_ , \new_[74707]_ , \new_[74708]_ ,
    \new_[74709]_ , \new_[74712]_ , \new_[74715]_ , \new_[74716]_ ,
    \new_[74719]_ , \new_[74722]_ , \new_[74723]_ , \new_[74724]_ ,
    \new_[74728]_ , \new_[74729]_ , \new_[74732]_ , \new_[74735]_ ,
    \new_[74736]_ , \new_[74737]_ , \new_[74740]_ , \new_[74743]_ ,
    \new_[74744]_ , \new_[74747]_ , \new_[74750]_ , \new_[74751]_ ,
    \new_[74752]_ , \new_[74756]_ , \new_[74757]_ , \new_[74760]_ ,
    \new_[74763]_ , \new_[74764]_ , \new_[74765]_ , \new_[74768]_ ,
    \new_[74771]_ , \new_[74772]_ , \new_[74775]_ , \new_[74778]_ ,
    \new_[74779]_ , \new_[74780]_ , \new_[74784]_ , \new_[74785]_ ,
    \new_[74788]_ , \new_[74791]_ , \new_[74792]_ , \new_[74793]_ ,
    \new_[74796]_ , \new_[74799]_ , \new_[74800]_ , \new_[74803]_ ,
    \new_[74806]_ , \new_[74807]_ , \new_[74808]_ , \new_[74812]_ ,
    \new_[74813]_ , \new_[74816]_ , \new_[74819]_ , \new_[74820]_ ,
    \new_[74821]_ , \new_[74824]_ , \new_[74827]_ , \new_[74828]_ ,
    \new_[74831]_ , \new_[74834]_ , \new_[74835]_ , \new_[74836]_ ,
    \new_[74840]_ , \new_[74841]_ , \new_[74844]_ , \new_[74847]_ ,
    \new_[74848]_ , \new_[74849]_ , \new_[74852]_ , \new_[74855]_ ,
    \new_[74856]_ , \new_[74859]_ , \new_[74862]_ , \new_[74863]_ ,
    \new_[74864]_ , \new_[74868]_ , \new_[74869]_ , \new_[74872]_ ,
    \new_[74875]_ , \new_[74876]_ , \new_[74877]_ , \new_[74880]_ ,
    \new_[74883]_ , \new_[74884]_ , \new_[74887]_ , \new_[74890]_ ,
    \new_[74891]_ , \new_[74892]_ , \new_[74896]_ , \new_[74897]_ ,
    \new_[74900]_ , \new_[74903]_ , \new_[74904]_ , \new_[74905]_ ,
    \new_[74908]_ , \new_[74911]_ , \new_[74912]_ , \new_[74915]_ ,
    \new_[74918]_ , \new_[74919]_ , \new_[74920]_ , \new_[74924]_ ,
    \new_[74925]_ , \new_[74928]_ , \new_[74931]_ , \new_[74932]_ ,
    \new_[74933]_ , \new_[74936]_ , \new_[74939]_ , \new_[74940]_ ,
    \new_[74943]_ , \new_[74946]_ , \new_[74947]_ , \new_[74948]_ ,
    \new_[74952]_ , \new_[74953]_ , \new_[74956]_ , \new_[74959]_ ,
    \new_[74960]_ , \new_[74961]_ , \new_[74964]_ , \new_[74967]_ ,
    \new_[74968]_ , \new_[74971]_ , \new_[74974]_ , \new_[74975]_ ,
    \new_[74976]_ , \new_[74980]_ , \new_[74981]_ , \new_[74984]_ ,
    \new_[74987]_ , \new_[74988]_ , \new_[74989]_ , \new_[74992]_ ,
    \new_[74995]_ , \new_[74996]_ , \new_[74999]_ , \new_[75002]_ ,
    \new_[75003]_ , \new_[75004]_ , \new_[75008]_ , \new_[75009]_ ,
    \new_[75012]_ , \new_[75015]_ , \new_[75016]_ , \new_[75017]_ ,
    \new_[75020]_ , \new_[75023]_ , \new_[75024]_ , \new_[75027]_ ,
    \new_[75030]_ , \new_[75031]_ , \new_[75032]_ , \new_[75036]_ ,
    \new_[75037]_ , \new_[75040]_ , \new_[75043]_ , \new_[75044]_ ,
    \new_[75045]_ , \new_[75048]_ , \new_[75051]_ , \new_[75052]_ ,
    \new_[75055]_ , \new_[75058]_ , \new_[75059]_ , \new_[75060]_ ,
    \new_[75064]_ , \new_[75065]_ , \new_[75068]_ , \new_[75071]_ ,
    \new_[75072]_ , \new_[75073]_ , \new_[75076]_ , \new_[75079]_ ,
    \new_[75080]_ , \new_[75083]_ , \new_[75086]_ , \new_[75087]_ ,
    \new_[75088]_ , \new_[75092]_ , \new_[75093]_ , \new_[75096]_ ,
    \new_[75099]_ , \new_[75100]_ , \new_[75101]_ , \new_[75104]_ ,
    \new_[75107]_ , \new_[75108]_ , \new_[75111]_ , \new_[75114]_ ,
    \new_[75115]_ , \new_[75116]_ , \new_[75120]_ , \new_[75121]_ ,
    \new_[75124]_ , \new_[75127]_ , \new_[75128]_ , \new_[75129]_ ,
    \new_[75132]_ , \new_[75135]_ , \new_[75136]_ , \new_[75139]_ ,
    \new_[75142]_ , \new_[75143]_ , \new_[75144]_ , \new_[75148]_ ,
    \new_[75149]_ , \new_[75152]_ , \new_[75155]_ , \new_[75156]_ ,
    \new_[75157]_ , \new_[75160]_ , \new_[75163]_ , \new_[75164]_ ,
    \new_[75167]_ , \new_[75170]_ , \new_[75171]_ , \new_[75172]_ ,
    \new_[75175]_ , \new_[75178]_ , \new_[75179]_ , \new_[75182]_ ,
    \new_[75185]_ , \new_[75186]_ , \new_[75187]_ , \new_[75190]_ ,
    \new_[75193]_ , \new_[75194]_ , \new_[75197]_ , \new_[75200]_ ,
    \new_[75201]_ , \new_[75202]_ , \new_[75205]_ , \new_[75208]_ ,
    \new_[75209]_ , \new_[75212]_ , \new_[75215]_ , \new_[75216]_ ,
    \new_[75217]_ , \new_[75220]_ , \new_[75223]_ , \new_[75224]_ ,
    \new_[75227]_ , \new_[75230]_ , \new_[75231]_ , \new_[75232]_ ,
    \new_[75235]_ , \new_[75238]_ , \new_[75239]_ , \new_[75242]_ ,
    \new_[75245]_ , \new_[75246]_ , \new_[75247]_ , \new_[75250]_ ,
    \new_[75253]_ , \new_[75254]_ , \new_[75257]_ , \new_[75260]_ ,
    \new_[75261]_ , \new_[75262]_ , \new_[75265]_ , \new_[75268]_ ,
    \new_[75269]_ , \new_[75272]_ , \new_[75275]_ , \new_[75276]_ ,
    \new_[75277]_ , \new_[75280]_ , \new_[75283]_ , \new_[75284]_ ,
    \new_[75287]_ , \new_[75290]_ , \new_[75291]_ , \new_[75292]_ ,
    \new_[75295]_ , \new_[75298]_ , \new_[75299]_ , \new_[75302]_ ,
    \new_[75305]_ , \new_[75306]_ , \new_[75307]_ , \new_[75310]_ ,
    \new_[75313]_ , \new_[75314]_ , \new_[75317]_ , \new_[75320]_ ,
    \new_[75321]_ , \new_[75322]_ , \new_[75325]_ , \new_[75328]_ ,
    \new_[75329]_ , \new_[75332]_ , \new_[75335]_ , \new_[75336]_ ,
    \new_[75337]_ , \new_[75340]_ , \new_[75343]_ , \new_[75344]_ ,
    \new_[75347]_ , \new_[75350]_ , \new_[75351]_ , \new_[75352]_ ,
    \new_[75355]_ , \new_[75358]_ , \new_[75359]_ , \new_[75362]_ ,
    \new_[75365]_ , \new_[75366]_ , \new_[75367]_ , \new_[75370]_ ,
    \new_[75373]_ , \new_[75374]_ , \new_[75377]_ , \new_[75380]_ ,
    \new_[75381]_ , \new_[75382]_ , \new_[75385]_ , \new_[75388]_ ,
    \new_[75389]_ , \new_[75392]_ , \new_[75395]_ , \new_[75396]_ ,
    \new_[75397]_ , \new_[75400]_ , \new_[75403]_ , \new_[75404]_ ,
    \new_[75407]_ , \new_[75410]_ , \new_[75411]_ , \new_[75412]_ ,
    \new_[75415]_ , \new_[75418]_ , \new_[75419]_ , \new_[75422]_ ,
    \new_[75425]_ , \new_[75426]_ , \new_[75427]_ , \new_[75430]_ ,
    \new_[75433]_ , \new_[75434]_ , \new_[75437]_ , \new_[75440]_ ,
    \new_[75441]_ , \new_[75442]_ , \new_[75445]_ , \new_[75448]_ ,
    \new_[75449]_ , \new_[75452]_ , \new_[75455]_ , \new_[75456]_ ,
    \new_[75457]_ , \new_[75460]_ , \new_[75463]_ , \new_[75464]_ ,
    \new_[75467]_ , \new_[75470]_ , \new_[75471]_ , \new_[75472]_ ,
    \new_[75475]_ , \new_[75478]_ , \new_[75479]_ , \new_[75482]_ ,
    \new_[75485]_ , \new_[75486]_ , \new_[75487]_ , \new_[75490]_ ,
    \new_[75493]_ , \new_[75494]_ , \new_[75497]_ , \new_[75500]_ ,
    \new_[75501]_ , \new_[75502]_ , \new_[75505]_ , \new_[75508]_ ,
    \new_[75509]_ , \new_[75512]_ , \new_[75515]_ , \new_[75516]_ ,
    \new_[75517]_ , \new_[75520]_ , \new_[75523]_ , \new_[75524]_ ,
    \new_[75527]_ , \new_[75530]_ , \new_[75531]_ , \new_[75532]_ ,
    \new_[75535]_ , \new_[75538]_ , \new_[75539]_ , \new_[75542]_ ,
    \new_[75545]_ , \new_[75546]_ , \new_[75547]_ , \new_[75550]_ ,
    \new_[75553]_ , \new_[75554]_ , \new_[75557]_ , \new_[75560]_ ,
    \new_[75561]_ , \new_[75562]_ , \new_[75565]_ , \new_[75568]_ ,
    \new_[75569]_ , \new_[75572]_ , \new_[75575]_ , \new_[75576]_ ,
    \new_[75577]_ , \new_[75580]_ , \new_[75583]_ , \new_[75584]_ ,
    \new_[75587]_ , \new_[75590]_ , \new_[75591]_ , \new_[75592]_ ,
    \new_[75595]_ , \new_[75598]_ , \new_[75599]_ , \new_[75602]_ ,
    \new_[75605]_ , \new_[75606]_ , \new_[75607]_ , \new_[75610]_ ,
    \new_[75613]_ , \new_[75614]_ , \new_[75617]_ , \new_[75620]_ ,
    \new_[75621]_ , \new_[75622]_ , \new_[75625]_ , \new_[75628]_ ,
    \new_[75629]_ , \new_[75632]_ , \new_[75635]_ , \new_[75636]_ ,
    \new_[75637]_ , \new_[75640]_ , \new_[75643]_ , \new_[75644]_ ,
    \new_[75647]_ , \new_[75650]_ , \new_[75651]_ , \new_[75652]_ ,
    \new_[75655]_ , \new_[75658]_ , \new_[75659]_ , \new_[75662]_ ,
    \new_[75665]_ , \new_[75666]_ , \new_[75667]_ , \new_[75670]_ ,
    \new_[75673]_ , \new_[75674]_ , \new_[75677]_ , \new_[75680]_ ,
    \new_[75681]_ , \new_[75682]_ , \new_[75685]_ , \new_[75688]_ ,
    \new_[75689]_ , \new_[75692]_ , \new_[75695]_ , \new_[75696]_ ,
    \new_[75697]_ , \new_[75700]_ , \new_[75703]_ , \new_[75704]_ ,
    \new_[75707]_ , \new_[75710]_ , \new_[75711]_ , \new_[75712]_ ,
    \new_[75715]_ , \new_[75718]_ , \new_[75719]_ , \new_[75722]_ ,
    \new_[75725]_ , \new_[75726]_ , \new_[75727]_ , \new_[75730]_ ,
    \new_[75733]_ , \new_[75734]_ , \new_[75737]_ , \new_[75740]_ ,
    \new_[75741]_ , \new_[75742]_ , \new_[75745]_ , \new_[75748]_ ,
    \new_[75749]_ , \new_[75752]_ , \new_[75755]_ , \new_[75756]_ ,
    \new_[75757]_ , \new_[75760]_ , \new_[75763]_ , \new_[75764]_ ,
    \new_[75767]_ , \new_[75770]_ , \new_[75771]_ , \new_[75772]_ ,
    \new_[75775]_ , \new_[75778]_ , \new_[75779]_ , \new_[75782]_ ,
    \new_[75785]_ , \new_[75786]_ , \new_[75787]_ , \new_[75790]_ ,
    \new_[75793]_ , \new_[75794]_ , \new_[75797]_ , \new_[75800]_ ,
    \new_[75801]_ , \new_[75802]_ , \new_[75805]_ , \new_[75808]_ ,
    \new_[75809]_ , \new_[75812]_ , \new_[75815]_ , \new_[75816]_ ,
    \new_[75817]_ , \new_[75820]_ , \new_[75823]_ , \new_[75824]_ ,
    \new_[75827]_ , \new_[75830]_ , \new_[75831]_ , \new_[75832]_ ,
    \new_[75835]_ , \new_[75838]_ , \new_[75839]_ , \new_[75842]_ ,
    \new_[75845]_ , \new_[75846]_ , \new_[75847]_ , \new_[75850]_ ,
    \new_[75853]_ , \new_[75854]_ , \new_[75857]_ , \new_[75860]_ ,
    \new_[75861]_ , \new_[75862]_ , \new_[75865]_ , \new_[75868]_ ,
    \new_[75869]_ , \new_[75872]_ , \new_[75875]_ , \new_[75876]_ ,
    \new_[75877]_ , \new_[75880]_ , \new_[75883]_ , \new_[75884]_ ,
    \new_[75887]_ , \new_[75890]_ , \new_[75891]_ , \new_[75892]_ ,
    \new_[75895]_ , \new_[75898]_ , \new_[75899]_ , \new_[75902]_ ,
    \new_[75905]_ , \new_[75906]_ , \new_[75907]_ , \new_[75910]_ ,
    \new_[75913]_ , \new_[75914]_ , \new_[75917]_ , \new_[75920]_ ,
    \new_[75921]_ , \new_[75922]_ , \new_[75925]_ , \new_[75928]_ ,
    \new_[75929]_ , \new_[75932]_ , \new_[75935]_ , \new_[75936]_ ,
    \new_[75937]_ , \new_[75940]_ , \new_[75943]_ , \new_[75944]_ ,
    \new_[75947]_ , \new_[75950]_ , \new_[75951]_ , \new_[75952]_ ,
    \new_[75955]_ , \new_[75958]_ , \new_[75959]_ , \new_[75962]_ ,
    \new_[75965]_ , \new_[75966]_ , \new_[75967]_ , \new_[75970]_ ,
    \new_[75973]_ , \new_[75974]_ , \new_[75977]_ , \new_[75980]_ ,
    \new_[75981]_ , \new_[75982]_ , \new_[75985]_ , \new_[75988]_ ,
    \new_[75989]_ , \new_[75992]_ , \new_[75995]_ , \new_[75996]_ ,
    \new_[75997]_ , \new_[76000]_ , \new_[76003]_ , \new_[76004]_ ,
    \new_[76007]_ , \new_[76010]_ , \new_[76011]_ , \new_[76012]_ ,
    \new_[76015]_ , \new_[76018]_ , \new_[76019]_ , \new_[76022]_ ,
    \new_[76025]_ , \new_[76026]_ , \new_[76027]_ , \new_[76030]_ ,
    \new_[76033]_ , \new_[76034]_ , \new_[76037]_ , \new_[76040]_ ,
    \new_[76041]_ , \new_[76042]_ , \new_[76045]_ , \new_[76048]_ ,
    \new_[76049]_ , \new_[76052]_ , \new_[76055]_ , \new_[76056]_ ,
    \new_[76057]_ , \new_[76060]_ , \new_[76063]_ , \new_[76064]_ ,
    \new_[76067]_ , \new_[76070]_ , \new_[76071]_ , \new_[76072]_ ,
    \new_[76075]_ , \new_[76078]_ , \new_[76079]_ , \new_[76082]_ ,
    \new_[76085]_ , \new_[76086]_ , \new_[76087]_ , \new_[76090]_ ,
    \new_[76093]_ , \new_[76094]_ , \new_[76097]_ , \new_[76100]_ ,
    \new_[76101]_ , \new_[76102]_ , \new_[76105]_ , \new_[76108]_ ,
    \new_[76109]_ , \new_[76112]_ , \new_[76115]_ , \new_[76116]_ ,
    \new_[76117]_ , \new_[76120]_ , \new_[76123]_ , \new_[76124]_ ,
    \new_[76127]_ , \new_[76130]_ , \new_[76131]_ , \new_[76132]_ ,
    \new_[76135]_ , \new_[76138]_ , \new_[76139]_ , \new_[76142]_ ,
    \new_[76145]_ , \new_[76146]_ , \new_[76147]_ , \new_[76150]_ ,
    \new_[76153]_ , \new_[76154]_ , \new_[76157]_ , \new_[76160]_ ,
    \new_[76161]_ , \new_[76162]_ , \new_[76165]_ , \new_[76168]_ ,
    \new_[76169]_ , \new_[76172]_ , \new_[76175]_ , \new_[76176]_ ,
    \new_[76177]_ , \new_[76180]_ , \new_[76183]_ , \new_[76184]_ ,
    \new_[76187]_ , \new_[76190]_ , \new_[76191]_ , \new_[76192]_ ,
    \new_[76195]_ , \new_[76198]_ , \new_[76199]_ , \new_[76202]_ ,
    \new_[76205]_ , \new_[76206]_ , \new_[76207]_ , \new_[76210]_ ,
    \new_[76213]_ , \new_[76214]_ , \new_[76217]_ , \new_[76220]_ ,
    \new_[76221]_ , \new_[76222]_ , \new_[76225]_ , \new_[76228]_ ,
    \new_[76229]_ , \new_[76232]_ , \new_[76235]_ , \new_[76236]_ ,
    \new_[76237]_ , \new_[76240]_ , \new_[76243]_ , \new_[76244]_ ,
    \new_[76247]_ , \new_[76250]_ , \new_[76251]_ , \new_[76252]_ ,
    \new_[76255]_ , \new_[76258]_ , \new_[76259]_ , \new_[76262]_ ,
    \new_[76265]_ , \new_[76266]_ , \new_[76267]_ , \new_[76270]_ ,
    \new_[76273]_ , \new_[76274]_ , \new_[76277]_ , \new_[76280]_ ,
    \new_[76281]_ , \new_[76282]_ , \new_[76285]_ , \new_[76288]_ ,
    \new_[76289]_ , \new_[76292]_ , \new_[76295]_ , \new_[76296]_ ,
    \new_[76297]_ , \new_[76300]_ , \new_[76303]_ , \new_[76304]_ ,
    \new_[76307]_ , \new_[76310]_ , \new_[76311]_ , \new_[76312]_ ,
    \new_[76315]_ , \new_[76318]_ , \new_[76319]_ , \new_[76322]_ ,
    \new_[76325]_ , \new_[76326]_ , \new_[76327]_ , \new_[76330]_ ,
    \new_[76333]_ , \new_[76334]_ , \new_[76337]_ , \new_[76340]_ ,
    \new_[76341]_ , \new_[76342]_ , \new_[76345]_ , \new_[76348]_ ,
    \new_[76349]_ , \new_[76352]_ , \new_[76355]_ , \new_[76356]_ ,
    \new_[76357]_ , \new_[76360]_ , \new_[76363]_ , \new_[76364]_ ,
    \new_[76367]_ , \new_[76370]_ , \new_[76371]_ , \new_[76372]_ ,
    \new_[76375]_ , \new_[76378]_ , \new_[76379]_ , \new_[76382]_ ,
    \new_[76385]_ , \new_[76386]_ , \new_[76387]_ , \new_[76390]_ ,
    \new_[76393]_ , \new_[76394]_ , \new_[76397]_ , \new_[76400]_ ,
    \new_[76401]_ , \new_[76402]_ , \new_[76405]_ , \new_[76408]_ ,
    \new_[76409]_ , \new_[76412]_ , \new_[76415]_ , \new_[76416]_ ,
    \new_[76417]_ , \new_[76420]_ , \new_[76423]_ , \new_[76424]_ ,
    \new_[76427]_ , \new_[76430]_ , \new_[76431]_ , \new_[76432]_ ,
    \new_[76435]_ , \new_[76438]_ , \new_[76439]_ , \new_[76442]_ ,
    \new_[76445]_ , \new_[76446]_ , \new_[76447]_ , \new_[76450]_ ,
    \new_[76453]_ , \new_[76454]_ , \new_[76457]_ , \new_[76460]_ ,
    \new_[76461]_ , \new_[76462]_ , \new_[76465]_ , \new_[76468]_ ,
    \new_[76469]_ , \new_[76472]_ , \new_[76475]_ , \new_[76476]_ ,
    \new_[76477]_ , \new_[76480]_ , \new_[76483]_ , \new_[76484]_ ,
    \new_[76487]_ , \new_[76490]_ , \new_[76491]_ , \new_[76492]_ ,
    \new_[76495]_ , \new_[76498]_ , \new_[76499]_ , \new_[76502]_ ,
    \new_[76505]_ , \new_[76506]_ , \new_[76507]_ , \new_[76510]_ ,
    \new_[76513]_ , \new_[76514]_ , \new_[76517]_ , \new_[76520]_ ,
    \new_[76521]_ , \new_[76522]_ , \new_[76525]_ , \new_[76528]_ ,
    \new_[76529]_ , \new_[76532]_ , \new_[76535]_ , \new_[76536]_ ,
    \new_[76537]_ , \new_[76540]_ , \new_[76543]_ , \new_[76544]_ ,
    \new_[76547]_ , \new_[76550]_ , \new_[76551]_ , \new_[76552]_ ,
    \new_[76555]_ , \new_[76558]_ , \new_[76559]_ , \new_[76562]_ ,
    \new_[76565]_ , \new_[76566]_ , \new_[76567]_ , \new_[76570]_ ,
    \new_[76573]_ , \new_[76574]_ , \new_[76577]_ , \new_[76580]_ ,
    \new_[76581]_ , \new_[76582]_ , \new_[76585]_ , \new_[76588]_ ,
    \new_[76589]_ , \new_[76592]_ , \new_[76595]_ , \new_[76596]_ ,
    \new_[76597]_ , \new_[76600]_ , \new_[76603]_ , \new_[76604]_ ,
    \new_[76607]_ , \new_[76610]_ , \new_[76611]_ , \new_[76612]_ ,
    \new_[76615]_ , \new_[76618]_ , \new_[76619]_ , \new_[76622]_ ,
    \new_[76625]_ , \new_[76626]_ , \new_[76627]_ , \new_[76630]_ ,
    \new_[76633]_ , \new_[76634]_ , \new_[76637]_ , \new_[76640]_ ,
    \new_[76641]_ , \new_[76642]_ , \new_[76645]_ , \new_[76648]_ ,
    \new_[76649]_ , \new_[76652]_ , \new_[76655]_ , \new_[76656]_ ,
    \new_[76657]_ , \new_[76660]_ , \new_[76663]_ , \new_[76664]_ ,
    \new_[76667]_ , \new_[76670]_ , \new_[76671]_ , \new_[76672]_ ,
    \new_[76675]_ , \new_[76678]_ , \new_[76679]_ , \new_[76682]_ ,
    \new_[76685]_ , \new_[76686]_ , \new_[76687]_ , \new_[76690]_ ,
    \new_[76693]_ , \new_[76694]_ , \new_[76697]_ , \new_[76700]_ ,
    \new_[76701]_ , \new_[76702]_ , \new_[76705]_ , \new_[76708]_ ,
    \new_[76709]_ , \new_[76712]_ , \new_[76715]_ , \new_[76716]_ ,
    \new_[76717]_ , \new_[76720]_ , \new_[76723]_ , \new_[76724]_ ,
    \new_[76727]_ , \new_[76730]_ , \new_[76731]_ , \new_[76732]_ ,
    \new_[76735]_ , \new_[76738]_ , \new_[76739]_ , \new_[76742]_ ,
    \new_[76745]_ , \new_[76746]_ , \new_[76747]_ , \new_[76750]_ ,
    \new_[76753]_ , \new_[76754]_ , \new_[76757]_ , \new_[76760]_ ,
    \new_[76761]_ , \new_[76762]_ , \new_[76765]_ , \new_[76768]_ ,
    \new_[76769]_ , \new_[76772]_ , \new_[76775]_ , \new_[76776]_ ,
    \new_[76777]_ , \new_[76780]_ , \new_[76783]_ , \new_[76784]_ ,
    \new_[76787]_ , \new_[76790]_ , \new_[76791]_ , \new_[76792]_ ,
    \new_[76795]_ , \new_[76798]_ , \new_[76799]_ , \new_[76802]_ ,
    \new_[76805]_ , \new_[76806]_ , \new_[76807]_ , \new_[76810]_ ,
    \new_[76813]_ , \new_[76814]_ , \new_[76817]_ , \new_[76820]_ ,
    \new_[76821]_ , \new_[76822]_ , \new_[76825]_ , \new_[76828]_ ,
    \new_[76829]_ , \new_[76832]_ , \new_[76835]_ , \new_[76836]_ ,
    \new_[76837]_ , \new_[76840]_ , \new_[76843]_ , \new_[76844]_ ,
    \new_[76847]_ , \new_[76850]_ , \new_[76851]_ , \new_[76852]_ ,
    \new_[76855]_ , \new_[76858]_ , \new_[76859]_ , \new_[76862]_ ,
    \new_[76865]_ , \new_[76866]_ , \new_[76867]_ , \new_[76870]_ ,
    \new_[76873]_ , \new_[76874]_ , \new_[76877]_ , \new_[76880]_ ,
    \new_[76881]_ , \new_[76882]_ , \new_[76885]_ , \new_[76888]_ ,
    \new_[76889]_ , \new_[76892]_ , \new_[76895]_ , \new_[76896]_ ,
    \new_[76897]_ , \new_[76900]_ , \new_[76903]_ , \new_[76904]_ ,
    \new_[76907]_ , \new_[76910]_ , \new_[76911]_ , \new_[76912]_ ,
    \new_[76915]_ , \new_[76918]_ , \new_[76919]_ , \new_[76922]_ ,
    \new_[76925]_ , \new_[76926]_ , \new_[76927]_ , \new_[76930]_ ,
    \new_[76933]_ , \new_[76934]_ , \new_[76937]_ , \new_[76940]_ ,
    \new_[76941]_ , \new_[76942]_ , \new_[76945]_ , \new_[76948]_ ,
    \new_[76949]_ , \new_[76952]_ , \new_[76955]_ , \new_[76956]_ ,
    \new_[76957]_ , \new_[76960]_ , \new_[76963]_ , \new_[76964]_ ,
    \new_[76967]_ , \new_[76970]_ , \new_[76971]_ , \new_[76972]_ ,
    \new_[76975]_ , \new_[76978]_ , \new_[76979]_ , \new_[76982]_ ,
    \new_[76985]_ , \new_[76986]_ , \new_[76987]_ , \new_[76990]_ ,
    \new_[76993]_ , \new_[76994]_ , \new_[76997]_ , \new_[77000]_ ,
    \new_[77001]_ , \new_[77002]_ , \new_[77005]_ , \new_[77008]_ ,
    \new_[77009]_ , \new_[77012]_ , \new_[77015]_ , \new_[77016]_ ,
    \new_[77017]_ , \new_[77020]_ , \new_[77023]_ , \new_[77024]_ ,
    \new_[77027]_ , \new_[77030]_ , \new_[77031]_ , \new_[77032]_ ,
    \new_[77035]_ , \new_[77038]_ , \new_[77039]_ , \new_[77042]_ ,
    \new_[77045]_ , \new_[77046]_ , \new_[77047]_ , \new_[77050]_ ,
    \new_[77053]_ , \new_[77054]_ , \new_[77057]_ , \new_[77060]_ ,
    \new_[77061]_ , \new_[77062]_ , \new_[77065]_ , \new_[77068]_ ,
    \new_[77069]_ , \new_[77072]_ , \new_[77075]_ , \new_[77076]_ ,
    \new_[77077]_ , \new_[77080]_ , \new_[77083]_ , \new_[77084]_ ,
    \new_[77087]_ , \new_[77090]_ , \new_[77091]_ , \new_[77092]_ ,
    \new_[77095]_ , \new_[77098]_ , \new_[77099]_ , \new_[77102]_ ,
    \new_[77105]_ , \new_[77106]_ , \new_[77107]_ , \new_[77110]_ ,
    \new_[77113]_ , \new_[77114]_ , \new_[77117]_ , \new_[77120]_ ,
    \new_[77121]_ , \new_[77122]_ , \new_[77125]_ , \new_[77128]_ ,
    \new_[77129]_ , \new_[77132]_ , \new_[77135]_ , \new_[77136]_ ,
    \new_[77137]_ , \new_[77140]_ , \new_[77143]_ , \new_[77144]_ ,
    \new_[77147]_ , \new_[77150]_ , \new_[77151]_ , \new_[77152]_ ,
    \new_[77155]_ , \new_[77158]_ , \new_[77159]_ , \new_[77162]_ ,
    \new_[77165]_ , \new_[77166]_ , \new_[77167]_ , \new_[77170]_ ,
    \new_[77173]_ , \new_[77174]_ , \new_[77177]_ , \new_[77180]_ ,
    \new_[77181]_ , \new_[77182]_ , \new_[77185]_ , \new_[77188]_ ,
    \new_[77189]_ , \new_[77192]_ , \new_[77195]_ , \new_[77196]_ ,
    \new_[77197]_ , \new_[77200]_ , \new_[77203]_ , \new_[77204]_ ,
    \new_[77207]_ , \new_[77210]_ , \new_[77211]_ , \new_[77212]_ ,
    \new_[77215]_ , \new_[77218]_ , \new_[77219]_ , \new_[77222]_ ,
    \new_[77225]_ , \new_[77226]_ , \new_[77227]_ , \new_[77230]_ ,
    \new_[77233]_ , \new_[77234]_ , \new_[77237]_ , \new_[77240]_ ,
    \new_[77241]_ , \new_[77242]_ , \new_[77245]_ , \new_[77248]_ ,
    \new_[77249]_ , \new_[77252]_ , \new_[77255]_ , \new_[77256]_ ,
    \new_[77257]_ , \new_[77260]_ , \new_[77263]_ , \new_[77264]_ ,
    \new_[77267]_ , \new_[77270]_ , \new_[77271]_ , \new_[77272]_ ,
    \new_[77275]_ , \new_[77278]_ , \new_[77279]_ , \new_[77282]_ ,
    \new_[77285]_ , \new_[77286]_ , \new_[77287]_ , \new_[77290]_ ,
    \new_[77293]_ , \new_[77294]_ , \new_[77297]_ , \new_[77300]_ ,
    \new_[77301]_ , \new_[77302]_ , \new_[77305]_ , \new_[77308]_ ,
    \new_[77309]_ , \new_[77312]_ , \new_[77315]_ , \new_[77316]_ ,
    \new_[77317]_ , \new_[77320]_ , \new_[77323]_ , \new_[77324]_ ,
    \new_[77327]_ , \new_[77330]_ , \new_[77331]_ , \new_[77332]_ ,
    \new_[77335]_ , \new_[77338]_ , \new_[77339]_ , \new_[77342]_ ,
    \new_[77345]_ , \new_[77346]_ , \new_[77347]_ , \new_[77350]_ ,
    \new_[77353]_ , \new_[77354]_ , \new_[77357]_ , \new_[77360]_ ,
    \new_[77361]_ , \new_[77362]_ , \new_[77365]_ , \new_[77368]_ ,
    \new_[77369]_ , \new_[77372]_ , \new_[77375]_ , \new_[77376]_ ,
    \new_[77377]_ , \new_[77380]_ , \new_[77383]_ , \new_[77384]_ ,
    \new_[77387]_ , \new_[77390]_ , \new_[77391]_ , \new_[77392]_ ,
    \new_[77395]_ , \new_[77398]_ , \new_[77399]_ , \new_[77402]_ ,
    \new_[77405]_ , \new_[77406]_ , \new_[77407]_ , \new_[77410]_ ,
    \new_[77413]_ , \new_[77414]_ , \new_[77417]_ , \new_[77420]_ ,
    \new_[77421]_ , \new_[77422]_ , \new_[77425]_ , \new_[77428]_ ,
    \new_[77429]_ , \new_[77432]_ , \new_[77435]_ , \new_[77436]_ ,
    \new_[77437]_ , \new_[77440]_ , \new_[77443]_ , \new_[77444]_ ,
    \new_[77447]_ , \new_[77450]_ , \new_[77451]_ , \new_[77452]_ ,
    \new_[77455]_ , \new_[77458]_ , \new_[77459]_ , \new_[77462]_ ,
    \new_[77465]_ , \new_[77466]_ , \new_[77467]_ , \new_[77470]_ ,
    \new_[77473]_ , \new_[77474]_ , \new_[77477]_ , \new_[77480]_ ,
    \new_[77481]_ , \new_[77482]_ , \new_[77485]_ , \new_[77488]_ ,
    \new_[77489]_ , \new_[77492]_ , \new_[77495]_ , \new_[77496]_ ,
    \new_[77497]_ , \new_[77500]_ , \new_[77503]_ , \new_[77504]_ ,
    \new_[77507]_ , \new_[77510]_ , \new_[77511]_ , \new_[77512]_ ,
    \new_[77515]_ , \new_[77518]_ , \new_[77519]_ , \new_[77522]_ ,
    \new_[77525]_ , \new_[77526]_ , \new_[77527]_ , \new_[77530]_ ,
    \new_[77533]_ , \new_[77534]_ , \new_[77537]_ , \new_[77540]_ ,
    \new_[77541]_ , \new_[77542]_ , \new_[77545]_ , \new_[77548]_ ,
    \new_[77549]_ , \new_[77552]_ , \new_[77555]_ , \new_[77556]_ ,
    \new_[77557]_ , \new_[77560]_ , \new_[77563]_ , \new_[77564]_ ,
    \new_[77567]_ , \new_[77570]_ , \new_[77571]_ , \new_[77572]_ ,
    \new_[77575]_ , \new_[77578]_ , \new_[77579]_ , \new_[77582]_ ,
    \new_[77585]_ , \new_[77586]_ , \new_[77587]_ , \new_[77590]_ ,
    \new_[77593]_ , \new_[77594]_ , \new_[77597]_ , \new_[77600]_ ,
    \new_[77601]_ , \new_[77602]_ , \new_[77605]_ , \new_[77608]_ ,
    \new_[77609]_ , \new_[77612]_ , \new_[77615]_ , \new_[77616]_ ,
    \new_[77617]_ , \new_[77620]_ , \new_[77623]_ , \new_[77624]_ ,
    \new_[77627]_ , \new_[77630]_ , \new_[77631]_ , \new_[77632]_ ,
    \new_[77635]_ , \new_[77638]_ , \new_[77639]_ , \new_[77642]_ ,
    \new_[77645]_ , \new_[77646]_ , \new_[77647]_ , \new_[77650]_ ,
    \new_[77653]_ , \new_[77654]_ , \new_[77657]_ , \new_[77660]_ ,
    \new_[77661]_ , \new_[77662]_ , \new_[77665]_ , \new_[77668]_ ,
    \new_[77669]_ , \new_[77672]_ , \new_[77675]_ , \new_[77676]_ ,
    \new_[77677]_ , \new_[77680]_ , \new_[77683]_ , \new_[77684]_ ,
    \new_[77687]_ , \new_[77690]_ , \new_[77691]_ , \new_[77692]_ ,
    \new_[77695]_ , \new_[77698]_ , \new_[77699]_ , \new_[77702]_ ,
    \new_[77705]_ , \new_[77706]_ , \new_[77707]_ , \new_[77710]_ ,
    \new_[77713]_ , \new_[77714]_ , \new_[77717]_ , \new_[77720]_ ,
    \new_[77721]_ , \new_[77722]_ , \new_[77725]_ , \new_[77728]_ ,
    \new_[77729]_ , \new_[77732]_ , \new_[77735]_ , \new_[77736]_ ,
    \new_[77737]_ , \new_[77740]_ , \new_[77743]_ , \new_[77744]_ ,
    \new_[77747]_ , \new_[77750]_ , \new_[77751]_ , \new_[77752]_ ,
    \new_[77755]_ , \new_[77758]_ , \new_[77759]_ , \new_[77762]_ ,
    \new_[77765]_ , \new_[77766]_ , \new_[77767]_ , \new_[77770]_ ,
    \new_[77773]_ , \new_[77774]_ , \new_[77777]_ , \new_[77780]_ ,
    \new_[77781]_ , \new_[77782]_ , \new_[77785]_ , \new_[77788]_ ,
    \new_[77789]_ , \new_[77792]_ , \new_[77795]_ , \new_[77796]_ ,
    \new_[77797]_ , \new_[77800]_ , \new_[77803]_ , \new_[77804]_ ,
    \new_[77807]_ , \new_[77810]_ , \new_[77811]_ , \new_[77812]_ ,
    \new_[77815]_ , \new_[77818]_ , \new_[77819]_ , \new_[77822]_ ,
    \new_[77825]_ , \new_[77826]_ , \new_[77827]_ , \new_[77830]_ ,
    \new_[77833]_ , \new_[77834]_ , \new_[77837]_ , \new_[77840]_ ,
    \new_[77841]_ , \new_[77842]_ , \new_[77845]_ , \new_[77848]_ ,
    \new_[77849]_ , \new_[77852]_ , \new_[77855]_ , \new_[77856]_ ,
    \new_[77857]_ , \new_[77860]_ , \new_[77863]_ , \new_[77864]_ ,
    \new_[77867]_ , \new_[77870]_ , \new_[77871]_ , \new_[77872]_ ,
    \new_[77875]_ , \new_[77878]_ , \new_[77879]_ , \new_[77882]_ ,
    \new_[77885]_ , \new_[77886]_ , \new_[77887]_ , \new_[77890]_ ,
    \new_[77893]_ , \new_[77894]_ , \new_[77897]_ , \new_[77900]_ ,
    \new_[77901]_ , \new_[77902]_ , \new_[77905]_ , \new_[77908]_ ,
    \new_[77909]_ , \new_[77912]_ , \new_[77915]_ , \new_[77916]_ ,
    \new_[77917]_ , \new_[77920]_ , \new_[77923]_ , \new_[77924]_ ,
    \new_[77927]_ , \new_[77930]_ , \new_[77931]_ , \new_[77932]_ ,
    \new_[77935]_ , \new_[77938]_ , \new_[77939]_ , \new_[77942]_ ,
    \new_[77945]_ , \new_[77946]_ , \new_[77947]_ , \new_[77950]_ ,
    \new_[77953]_ , \new_[77954]_ , \new_[77957]_ , \new_[77960]_ ,
    \new_[77961]_ , \new_[77962]_ , \new_[77965]_ , \new_[77968]_ ,
    \new_[77969]_ , \new_[77972]_ , \new_[77975]_ , \new_[77976]_ ,
    \new_[77977]_ , \new_[77980]_ , \new_[77983]_ , \new_[77984]_ ,
    \new_[77987]_ , \new_[77990]_ , \new_[77991]_ , \new_[77992]_ ,
    \new_[77995]_ , \new_[77998]_ , \new_[77999]_ , \new_[78002]_ ,
    \new_[78005]_ , \new_[78006]_ , \new_[78007]_ , \new_[78010]_ ,
    \new_[78013]_ , \new_[78014]_ , \new_[78017]_ , \new_[78020]_ ,
    \new_[78021]_ , \new_[78022]_ , \new_[78025]_ , \new_[78028]_ ,
    \new_[78029]_ , \new_[78032]_ , \new_[78035]_ , \new_[78036]_ ,
    \new_[78037]_ , \new_[78040]_ , \new_[78043]_ , \new_[78044]_ ,
    \new_[78047]_ , \new_[78050]_ , \new_[78051]_ , \new_[78052]_ ,
    \new_[78055]_ , \new_[78058]_ , \new_[78059]_ , \new_[78062]_ ,
    \new_[78065]_ , \new_[78066]_ , \new_[78067]_ , \new_[78070]_ ,
    \new_[78073]_ , \new_[78074]_ , \new_[78077]_ , \new_[78080]_ ,
    \new_[78081]_ , \new_[78082]_ , \new_[78085]_ , \new_[78088]_ ,
    \new_[78089]_ , \new_[78092]_ , \new_[78095]_ , \new_[78096]_ ,
    \new_[78097]_ , \new_[78100]_ , \new_[78103]_ , \new_[78104]_ ,
    \new_[78107]_ , \new_[78110]_ , \new_[78111]_ , \new_[78112]_ ,
    \new_[78115]_ , \new_[78118]_ , \new_[78119]_ , \new_[78122]_ ,
    \new_[78125]_ , \new_[78126]_ , \new_[78127]_ , \new_[78130]_ ,
    \new_[78133]_ , \new_[78134]_ , \new_[78137]_ , \new_[78140]_ ,
    \new_[78141]_ , \new_[78142]_ , \new_[78145]_ , \new_[78148]_ ,
    \new_[78149]_ , \new_[78152]_ , \new_[78155]_ , \new_[78156]_ ,
    \new_[78157]_ , \new_[78160]_ , \new_[78163]_ , \new_[78164]_ ,
    \new_[78167]_ , \new_[78170]_ , \new_[78171]_ , \new_[78172]_ ,
    \new_[78175]_ , \new_[78178]_ , \new_[78179]_ , \new_[78182]_ ,
    \new_[78185]_ , \new_[78186]_ , \new_[78187]_ , \new_[78190]_ ,
    \new_[78193]_ , \new_[78194]_ , \new_[78197]_ , \new_[78200]_ ,
    \new_[78201]_ , \new_[78202]_ , \new_[78205]_ , \new_[78208]_ ,
    \new_[78209]_ , \new_[78212]_ , \new_[78215]_ , \new_[78216]_ ,
    \new_[78217]_ , \new_[78220]_ , \new_[78223]_ , \new_[78224]_ ,
    \new_[78227]_ , \new_[78230]_ , \new_[78231]_ , \new_[78232]_ ,
    \new_[78235]_ , \new_[78238]_ , \new_[78239]_ , \new_[78242]_ ,
    \new_[78245]_ , \new_[78246]_ , \new_[78247]_ , \new_[78250]_ ,
    \new_[78253]_ , \new_[78254]_ , \new_[78257]_ , \new_[78260]_ ,
    \new_[78261]_ , \new_[78262]_ , \new_[78265]_ , \new_[78268]_ ,
    \new_[78269]_ , \new_[78272]_ , \new_[78275]_ , \new_[78276]_ ,
    \new_[78277]_ , \new_[78280]_ , \new_[78283]_ , \new_[78284]_ ,
    \new_[78287]_ , \new_[78290]_ , \new_[78291]_ , \new_[78292]_ ,
    \new_[78295]_ , \new_[78298]_ , \new_[78299]_ , \new_[78302]_ ,
    \new_[78305]_ , \new_[78306]_ , \new_[78307]_ , \new_[78310]_ ,
    \new_[78313]_ , \new_[78314]_ , \new_[78317]_ , \new_[78320]_ ,
    \new_[78321]_ , \new_[78322]_ , \new_[78325]_ , \new_[78328]_ ,
    \new_[78329]_ , \new_[78332]_ , \new_[78335]_ , \new_[78336]_ ,
    \new_[78337]_ , \new_[78340]_ , \new_[78343]_ , \new_[78344]_ ,
    \new_[78347]_ , \new_[78350]_ , \new_[78351]_ , \new_[78352]_ ,
    \new_[78355]_ , \new_[78358]_ , \new_[78359]_ , \new_[78362]_ ,
    \new_[78365]_ , \new_[78366]_ , \new_[78367]_ , \new_[78370]_ ,
    \new_[78373]_ , \new_[78374]_ , \new_[78377]_ , \new_[78380]_ ,
    \new_[78381]_ , \new_[78382]_ , \new_[78385]_ , \new_[78388]_ ,
    \new_[78389]_ , \new_[78392]_ , \new_[78395]_ , \new_[78396]_ ,
    \new_[78397]_ , \new_[78400]_ , \new_[78403]_ , \new_[78404]_ ,
    \new_[78407]_ , \new_[78410]_ , \new_[78411]_ , \new_[78412]_ ,
    \new_[78415]_ , \new_[78418]_ , \new_[78419]_ , \new_[78422]_ ,
    \new_[78425]_ , \new_[78426]_ , \new_[78427]_ , \new_[78430]_ ,
    \new_[78433]_ , \new_[78434]_ , \new_[78437]_ , \new_[78440]_ ,
    \new_[78441]_ , \new_[78442]_ , \new_[78445]_ , \new_[78448]_ ,
    \new_[78449]_ , \new_[78452]_ , \new_[78455]_ , \new_[78456]_ ,
    \new_[78457]_ , \new_[78460]_ , \new_[78463]_ , \new_[78464]_ ,
    \new_[78467]_ , \new_[78470]_ , \new_[78471]_ , \new_[78472]_ ,
    \new_[78475]_ , \new_[78478]_ , \new_[78479]_ , \new_[78482]_ ,
    \new_[78485]_ , \new_[78486]_ , \new_[78487]_ , \new_[78490]_ ,
    \new_[78493]_ , \new_[78494]_ , \new_[78497]_ , \new_[78500]_ ,
    \new_[78501]_ , \new_[78502]_ , \new_[78505]_ , \new_[78508]_ ,
    \new_[78509]_ , \new_[78512]_ , \new_[78515]_ , \new_[78516]_ ,
    \new_[78517]_ , \new_[78520]_ , \new_[78523]_ , \new_[78524]_ ,
    \new_[78527]_ , \new_[78530]_ , \new_[78531]_ , \new_[78532]_ ,
    \new_[78535]_ , \new_[78538]_ , \new_[78539]_ , \new_[78542]_ ,
    \new_[78545]_ , \new_[78546]_ , \new_[78547]_ , \new_[78550]_ ,
    \new_[78553]_ , \new_[78554]_ , \new_[78557]_ , \new_[78560]_ ,
    \new_[78561]_ , \new_[78562]_ , \new_[78565]_ , \new_[78568]_ ,
    \new_[78569]_ , \new_[78572]_ , \new_[78575]_ , \new_[78576]_ ,
    \new_[78577]_ , \new_[78580]_ , \new_[78583]_ , \new_[78584]_ ,
    \new_[78587]_ , \new_[78590]_ , \new_[78591]_ , \new_[78592]_ ,
    \new_[78595]_ , \new_[78598]_ , \new_[78599]_ , \new_[78602]_ ,
    \new_[78605]_ , \new_[78606]_ , \new_[78607]_ , \new_[78610]_ ,
    \new_[78613]_ , \new_[78614]_ , \new_[78617]_ , \new_[78620]_ ,
    \new_[78621]_ , \new_[78622]_ , \new_[78625]_ , \new_[78628]_ ,
    \new_[78629]_ , \new_[78632]_ , \new_[78635]_ , \new_[78636]_ ,
    \new_[78637]_ , \new_[78640]_ , \new_[78643]_ , \new_[78644]_ ,
    \new_[78647]_ , \new_[78650]_ , \new_[78651]_ , \new_[78652]_ ,
    \new_[78655]_ , \new_[78658]_ , \new_[78659]_ , \new_[78662]_ ,
    \new_[78665]_ , \new_[78666]_ , \new_[78667]_ , \new_[78670]_ ,
    \new_[78673]_ , \new_[78674]_ , \new_[78677]_ , \new_[78680]_ ,
    \new_[78681]_ , \new_[78682]_ , \new_[78685]_ , \new_[78688]_ ,
    \new_[78689]_ , \new_[78692]_ , \new_[78695]_ , \new_[78696]_ ,
    \new_[78697]_ , \new_[78700]_ , \new_[78703]_ , \new_[78704]_ ,
    \new_[78707]_ , \new_[78710]_ , \new_[78711]_ , \new_[78712]_ ,
    \new_[78715]_ , \new_[78718]_ , \new_[78719]_ , \new_[78722]_ ,
    \new_[78725]_ , \new_[78726]_ , \new_[78727]_ , \new_[78730]_ ,
    \new_[78733]_ , \new_[78734]_ , \new_[78737]_ , \new_[78740]_ ,
    \new_[78741]_ , \new_[78742]_ , \new_[78745]_ , \new_[78748]_ ,
    \new_[78749]_ , \new_[78752]_ , \new_[78755]_ , \new_[78756]_ ,
    \new_[78757]_ , \new_[78760]_ , \new_[78763]_ , \new_[78764]_ ,
    \new_[78767]_ , \new_[78770]_ , \new_[78771]_ , \new_[78772]_ ,
    \new_[78775]_ , \new_[78778]_ , \new_[78779]_ , \new_[78782]_ ,
    \new_[78785]_ , \new_[78786]_ , \new_[78787]_ , \new_[78790]_ ,
    \new_[78793]_ , \new_[78794]_ , \new_[78797]_ , \new_[78800]_ ,
    \new_[78801]_ , \new_[78802]_ , \new_[78805]_ , \new_[78808]_ ,
    \new_[78809]_ , \new_[78812]_ , \new_[78815]_ , \new_[78816]_ ,
    \new_[78817]_ , \new_[78820]_ , \new_[78823]_ , \new_[78824]_ ,
    \new_[78827]_ , \new_[78830]_ , \new_[78831]_ , \new_[78832]_ ,
    \new_[78835]_ , \new_[78838]_ , \new_[78839]_ , \new_[78842]_ ,
    \new_[78845]_ , \new_[78846]_ , \new_[78847]_ , \new_[78850]_ ,
    \new_[78853]_ , \new_[78854]_ , \new_[78857]_ , \new_[78860]_ ,
    \new_[78861]_ , \new_[78862]_ , \new_[78865]_ , \new_[78868]_ ,
    \new_[78869]_ , \new_[78872]_ , \new_[78875]_ , \new_[78876]_ ,
    \new_[78877]_ , \new_[78880]_ , \new_[78883]_ , \new_[78884]_ ,
    \new_[78887]_ , \new_[78890]_ , \new_[78891]_ , \new_[78892]_ ,
    \new_[78895]_ , \new_[78898]_ , \new_[78899]_ , \new_[78902]_ ,
    \new_[78905]_ , \new_[78906]_ , \new_[78907]_ , \new_[78910]_ ,
    \new_[78913]_ , \new_[78914]_ , \new_[78917]_ , \new_[78920]_ ,
    \new_[78921]_ , \new_[78922]_ , \new_[78925]_ , \new_[78928]_ ,
    \new_[78929]_ , \new_[78932]_ , \new_[78935]_ , \new_[78936]_ ,
    \new_[78937]_ , \new_[78940]_ , \new_[78943]_ , \new_[78944]_ ,
    \new_[78947]_ , \new_[78950]_ , \new_[78951]_ , \new_[78952]_ ,
    \new_[78955]_ , \new_[78958]_ , \new_[78959]_ , \new_[78962]_ ,
    \new_[78965]_ , \new_[78966]_ , \new_[78967]_ , \new_[78970]_ ,
    \new_[78973]_ , \new_[78974]_ , \new_[78977]_ , \new_[78980]_ ,
    \new_[78981]_ , \new_[78982]_ , \new_[78985]_ , \new_[78988]_ ,
    \new_[78989]_ , \new_[78992]_ , \new_[78995]_ , \new_[78996]_ ,
    \new_[78997]_ , \new_[79000]_ , \new_[79003]_ , \new_[79004]_ ,
    \new_[79007]_ , \new_[79010]_ , \new_[79011]_ , \new_[79012]_ ,
    \new_[79015]_ , \new_[79018]_ , \new_[79019]_ , \new_[79022]_ ,
    \new_[79025]_ , \new_[79026]_ , \new_[79027]_ , \new_[79030]_ ,
    \new_[79033]_ , \new_[79034]_ , \new_[79037]_ , \new_[79040]_ ,
    \new_[79041]_ , \new_[79042]_ , \new_[79045]_ , \new_[79048]_ ,
    \new_[79049]_ , \new_[79052]_ , \new_[79055]_ , \new_[79056]_ ,
    \new_[79057]_ , \new_[79060]_ , \new_[79063]_ , \new_[79064]_ ,
    \new_[79067]_ , \new_[79070]_ , \new_[79071]_ , \new_[79072]_ ,
    \new_[79075]_ , \new_[79078]_ , \new_[79079]_ , \new_[79082]_ ,
    \new_[79085]_ , \new_[79086]_ , \new_[79087]_ , \new_[79090]_ ,
    \new_[79093]_ , \new_[79094]_ , \new_[79097]_ , \new_[79100]_ ,
    \new_[79101]_ , \new_[79102]_ , \new_[79105]_ , \new_[79108]_ ,
    \new_[79109]_ , \new_[79112]_ , \new_[79115]_ , \new_[79116]_ ,
    \new_[79117]_ , \new_[79120]_ , \new_[79123]_ , \new_[79124]_ ,
    \new_[79127]_ , \new_[79130]_ , \new_[79131]_ , \new_[79132]_ ,
    \new_[79135]_ , \new_[79138]_ , \new_[79139]_ , \new_[79142]_ ,
    \new_[79145]_ , \new_[79146]_ , \new_[79147]_ , \new_[79150]_ ,
    \new_[79153]_ , \new_[79154]_ , \new_[79157]_ , \new_[79160]_ ,
    \new_[79161]_ , \new_[79162]_ , \new_[79165]_ , \new_[79168]_ ,
    \new_[79169]_ , \new_[79172]_ , \new_[79175]_ , \new_[79176]_ ,
    \new_[79177]_ , \new_[79180]_ , \new_[79183]_ , \new_[79184]_ ,
    \new_[79187]_ , \new_[79190]_ , \new_[79191]_ , \new_[79192]_ ,
    \new_[79195]_ , \new_[79198]_ , \new_[79199]_ , \new_[79202]_ ,
    \new_[79205]_ , \new_[79206]_ , \new_[79207]_ , \new_[79210]_ ,
    \new_[79213]_ , \new_[79214]_ , \new_[79217]_ , \new_[79220]_ ,
    \new_[79221]_ , \new_[79222]_ , \new_[79225]_ , \new_[79228]_ ,
    \new_[79229]_ , \new_[79232]_ , \new_[79235]_ , \new_[79236]_ ,
    \new_[79237]_ , \new_[79240]_ , \new_[79243]_ , \new_[79244]_ ,
    \new_[79247]_ , \new_[79250]_ , \new_[79251]_ , \new_[79252]_ ,
    \new_[79255]_ , \new_[79258]_ , \new_[79259]_ , \new_[79262]_ ,
    \new_[79265]_ , \new_[79266]_ , \new_[79267]_ , \new_[79270]_ ,
    \new_[79273]_ , \new_[79274]_ , \new_[79277]_ , \new_[79280]_ ,
    \new_[79281]_ , \new_[79282]_ , \new_[79285]_ , \new_[79288]_ ,
    \new_[79289]_ , \new_[79292]_ , \new_[79295]_ , \new_[79296]_ ,
    \new_[79297]_ , \new_[79300]_ , \new_[79303]_ , \new_[79304]_ ,
    \new_[79307]_ , \new_[79310]_ , \new_[79311]_ , \new_[79312]_ ,
    \new_[79315]_ , \new_[79318]_ , \new_[79319]_ , \new_[79322]_ ,
    \new_[79325]_ , \new_[79326]_ , \new_[79327]_ , \new_[79330]_ ,
    \new_[79333]_ , \new_[79334]_ , \new_[79337]_ , \new_[79340]_ ,
    \new_[79341]_ , \new_[79342]_ , \new_[79345]_ , \new_[79348]_ ,
    \new_[79349]_ , \new_[79352]_ , \new_[79355]_ , \new_[79356]_ ,
    \new_[79357]_ , \new_[79360]_ , \new_[79363]_ , \new_[79364]_ ,
    \new_[79367]_ , \new_[79370]_ , \new_[79371]_ , \new_[79372]_ ,
    \new_[79375]_ , \new_[79378]_ , \new_[79379]_ , \new_[79382]_ ,
    \new_[79385]_ , \new_[79386]_ , \new_[79387]_ , \new_[79390]_ ,
    \new_[79393]_ , \new_[79394]_ , \new_[79397]_ , \new_[79400]_ ,
    \new_[79401]_ , \new_[79402]_ , \new_[79405]_ , \new_[79408]_ ,
    \new_[79409]_ , \new_[79412]_ , \new_[79415]_ , \new_[79416]_ ,
    \new_[79417]_ , \new_[79420]_ , \new_[79423]_ , \new_[79424]_ ,
    \new_[79427]_ , \new_[79430]_ , \new_[79431]_ , \new_[79432]_ ,
    \new_[79435]_ , \new_[79438]_ , \new_[79439]_ , \new_[79442]_ ,
    \new_[79445]_ , \new_[79446]_ , \new_[79447]_ , \new_[79450]_ ,
    \new_[79453]_ , \new_[79454]_ , \new_[79457]_ , \new_[79460]_ ,
    \new_[79461]_ , \new_[79462]_ , \new_[79465]_ , \new_[79468]_ ,
    \new_[79469]_ , \new_[79472]_ , \new_[79475]_ , \new_[79476]_ ,
    \new_[79477]_ , \new_[79480]_ , \new_[79483]_ , \new_[79484]_ ,
    \new_[79487]_ , \new_[79490]_ , \new_[79491]_ , \new_[79492]_ ,
    \new_[79495]_ , \new_[79498]_ , \new_[79499]_ , \new_[79502]_ ,
    \new_[79505]_ , \new_[79506]_ , \new_[79507]_ , \new_[79510]_ ,
    \new_[79513]_ , \new_[79514]_ , \new_[79517]_ , \new_[79520]_ ,
    \new_[79521]_ , \new_[79522]_ , \new_[79525]_ , \new_[79528]_ ,
    \new_[79529]_ , \new_[79532]_ , \new_[79535]_ , \new_[79536]_ ,
    \new_[79537]_ , \new_[79540]_ , \new_[79543]_ , \new_[79544]_ ,
    \new_[79547]_ , \new_[79550]_ , \new_[79551]_ , \new_[79552]_ ,
    \new_[79555]_ , \new_[79558]_ , \new_[79559]_ , \new_[79562]_ ,
    \new_[79565]_ , \new_[79566]_ , \new_[79567]_ , \new_[79570]_ ,
    \new_[79573]_ , \new_[79574]_ , \new_[79577]_ , \new_[79580]_ ,
    \new_[79581]_ , \new_[79582]_ , \new_[79585]_ , \new_[79588]_ ,
    \new_[79589]_ , \new_[79592]_ , \new_[79595]_ , \new_[79596]_ ,
    \new_[79597]_ , \new_[79600]_ , \new_[79603]_ , \new_[79604]_ ,
    \new_[79607]_ , \new_[79610]_ , \new_[79611]_ , \new_[79612]_ ,
    \new_[79615]_ , \new_[79618]_ , \new_[79619]_ , \new_[79622]_ ,
    \new_[79625]_ , \new_[79626]_ , \new_[79627]_ , \new_[79630]_ ,
    \new_[79633]_ , \new_[79634]_ , \new_[79637]_ , \new_[79640]_ ,
    \new_[79641]_ , \new_[79642]_ , \new_[79645]_ , \new_[79648]_ ,
    \new_[79649]_ , \new_[79652]_ , \new_[79655]_ , \new_[79656]_ ,
    \new_[79657]_ , \new_[79660]_ , \new_[79663]_ , \new_[79664]_ ,
    \new_[79667]_ , \new_[79670]_ , \new_[79671]_ , \new_[79672]_ ,
    \new_[79675]_ , \new_[79678]_ , \new_[79679]_ , \new_[79682]_ ,
    \new_[79685]_ , \new_[79686]_ , \new_[79687]_ , \new_[79690]_ ,
    \new_[79693]_ , \new_[79694]_ , \new_[79697]_ , \new_[79700]_ ,
    \new_[79701]_ , \new_[79702]_ , \new_[79705]_ , \new_[79708]_ ,
    \new_[79709]_ , \new_[79712]_ , \new_[79715]_ , \new_[79716]_ ,
    \new_[79717]_ , \new_[79720]_ , \new_[79723]_ , \new_[79724]_ ,
    \new_[79727]_ , \new_[79730]_ , \new_[79731]_ , \new_[79732]_ ,
    \new_[79735]_ , \new_[79738]_ , \new_[79739]_ , \new_[79742]_ ,
    \new_[79745]_ , \new_[79746]_ , \new_[79747]_ , \new_[79750]_ ,
    \new_[79753]_ , \new_[79754]_ , \new_[79757]_ , \new_[79760]_ ,
    \new_[79761]_ , \new_[79762]_ , \new_[79765]_ , \new_[79768]_ ,
    \new_[79769]_ , \new_[79772]_ , \new_[79775]_ , \new_[79776]_ ,
    \new_[79777]_ , \new_[79780]_ , \new_[79783]_ , \new_[79784]_ ,
    \new_[79787]_ , \new_[79790]_ , \new_[79791]_ , \new_[79792]_ ,
    \new_[79795]_ , \new_[79798]_ , \new_[79799]_ , \new_[79802]_ ,
    \new_[79805]_ , \new_[79806]_ , \new_[79807]_ , \new_[79810]_ ,
    \new_[79813]_ , \new_[79814]_ , \new_[79817]_ , \new_[79820]_ ,
    \new_[79821]_ , \new_[79822]_ , \new_[79825]_ , \new_[79828]_ ,
    \new_[79829]_ , \new_[79832]_ , \new_[79835]_ , \new_[79836]_ ,
    \new_[79837]_ , \new_[79840]_ , \new_[79843]_ , \new_[79844]_ ,
    \new_[79847]_ , \new_[79850]_ , \new_[79851]_ , \new_[79852]_ ,
    \new_[79855]_ , \new_[79858]_ , \new_[79859]_ , \new_[79862]_ ,
    \new_[79865]_ , \new_[79866]_ , \new_[79867]_ , \new_[79870]_ ,
    \new_[79873]_ , \new_[79874]_ , \new_[79877]_ , \new_[79880]_ ,
    \new_[79881]_ , \new_[79882]_ , \new_[79885]_ , \new_[79888]_ ,
    \new_[79889]_ , \new_[79892]_ , \new_[79895]_ , \new_[79896]_ ,
    \new_[79897]_ , \new_[79900]_ , \new_[79903]_ , \new_[79904]_ ,
    \new_[79907]_ , \new_[79910]_ , \new_[79911]_ , \new_[79912]_ ,
    \new_[79915]_ , \new_[79918]_ , \new_[79919]_ , \new_[79922]_ ,
    \new_[79925]_ , \new_[79926]_ , \new_[79927]_ , \new_[79930]_ ,
    \new_[79933]_ , \new_[79934]_ , \new_[79937]_ , \new_[79940]_ ,
    \new_[79941]_ , \new_[79942]_ , \new_[79945]_ , \new_[79948]_ ,
    \new_[79949]_ , \new_[79952]_ , \new_[79955]_ , \new_[79956]_ ,
    \new_[79957]_ , \new_[79960]_ , \new_[79963]_ , \new_[79964]_ ,
    \new_[79967]_ , \new_[79970]_ , \new_[79971]_ , \new_[79972]_ ,
    \new_[79975]_ , \new_[79978]_ , \new_[79979]_ , \new_[79982]_ ,
    \new_[79985]_ , \new_[79986]_ , \new_[79987]_ , \new_[79990]_ ,
    \new_[79993]_ , \new_[79994]_ , \new_[79997]_ , \new_[80000]_ ,
    \new_[80001]_ , \new_[80002]_ , \new_[80005]_ , \new_[80008]_ ,
    \new_[80009]_ , \new_[80012]_ , \new_[80015]_ , \new_[80016]_ ,
    \new_[80017]_ , \new_[80020]_ , \new_[80023]_ , \new_[80024]_ ,
    \new_[80027]_ , \new_[80030]_ , \new_[80031]_ , \new_[80032]_ ,
    \new_[80035]_ , \new_[80038]_ , \new_[80039]_ , \new_[80042]_ ,
    \new_[80045]_ , \new_[80046]_ , \new_[80047]_ , \new_[80050]_ ,
    \new_[80053]_ , \new_[80054]_ , \new_[80057]_ , \new_[80060]_ ,
    \new_[80061]_ , \new_[80062]_ , \new_[80065]_ , \new_[80068]_ ,
    \new_[80069]_ , \new_[80072]_ , \new_[80075]_ , \new_[80076]_ ,
    \new_[80077]_ , \new_[80080]_ , \new_[80083]_ , \new_[80084]_ ,
    \new_[80087]_ , \new_[80090]_ , \new_[80091]_ , \new_[80092]_ ,
    \new_[80095]_ , \new_[80098]_ , \new_[80099]_ , \new_[80102]_ ,
    \new_[80105]_ , \new_[80106]_ , \new_[80107]_ , \new_[80110]_ ,
    \new_[80113]_ , \new_[80114]_ , \new_[80117]_ , \new_[80120]_ ,
    \new_[80121]_ , \new_[80122]_ , \new_[80125]_ , \new_[80128]_ ,
    \new_[80129]_ , \new_[80132]_ , \new_[80135]_ , \new_[80136]_ ,
    \new_[80137]_ , \new_[80140]_ , \new_[80143]_ , \new_[80144]_ ,
    \new_[80147]_ , \new_[80150]_ , \new_[80151]_ , \new_[80152]_ ,
    \new_[80155]_ , \new_[80158]_ , \new_[80159]_ , \new_[80162]_ ,
    \new_[80165]_ , \new_[80166]_ , \new_[80167]_ , \new_[80170]_ ,
    \new_[80173]_ , \new_[80174]_ , \new_[80177]_ , \new_[80180]_ ,
    \new_[80181]_ , \new_[80182]_ , \new_[80185]_ , \new_[80188]_ ,
    \new_[80189]_ , \new_[80192]_ , \new_[80195]_ , \new_[80196]_ ,
    \new_[80197]_ , \new_[80200]_ , \new_[80203]_ , \new_[80204]_ ,
    \new_[80207]_ , \new_[80210]_ , \new_[80211]_ , \new_[80212]_ ,
    \new_[80215]_ , \new_[80218]_ , \new_[80219]_ , \new_[80222]_ ,
    \new_[80225]_ , \new_[80226]_ , \new_[80227]_ , \new_[80230]_ ,
    \new_[80233]_ , \new_[80234]_ , \new_[80237]_ , \new_[80240]_ ,
    \new_[80241]_ , \new_[80242]_ , \new_[80245]_ , \new_[80248]_ ,
    \new_[80249]_ , \new_[80252]_ , \new_[80255]_ , \new_[80256]_ ,
    \new_[80257]_ , \new_[80260]_ , \new_[80263]_ , \new_[80264]_ ,
    \new_[80267]_ , \new_[80270]_ , \new_[80271]_ , \new_[80272]_ ,
    \new_[80275]_ , \new_[80278]_ , \new_[80279]_ , \new_[80282]_ ,
    \new_[80285]_ , \new_[80286]_ , \new_[80287]_ , \new_[80290]_ ,
    \new_[80293]_ , \new_[80294]_ , \new_[80297]_ , \new_[80300]_ ,
    \new_[80301]_ , \new_[80302]_ , \new_[80305]_ , \new_[80308]_ ,
    \new_[80309]_ , \new_[80312]_ , \new_[80315]_ , \new_[80316]_ ,
    \new_[80317]_ , \new_[80320]_ , \new_[80323]_ , \new_[80324]_ ,
    \new_[80327]_ , \new_[80330]_ , \new_[80331]_ , \new_[80332]_ ,
    \new_[80335]_ , \new_[80338]_ , \new_[80339]_ , \new_[80342]_ ,
    \new_[80345]_ , \new_[80346]_ , \new_[80347]_ , \new_[80350]_ ,
    \new_[80353]_ , \new_[80354]_ , \new_[80357]_ , \new_[80360]_ ,
    \new_[80361]_ , \new_[80362]_ , \new_[80365]_ , \new_[80368]_ ,
    \new_[80369]_ , \new_[80372]_ , \new_[80375]_ , \new_[80376]_ ,
    \new_[80377]_ , \new_[80380]_ , \new_[80383]_ , \new_[80384]_ ,
    \new_[80387]_ , \new_[80390]_ , \new_[80391]_ , \new_[80392]_ ,
    \new_[80395]_ , \new_[80398]_ , \new_[80399]_ , \new_[80402]_ ,
    \new_[80405]_ , \new_[80406]_ , \new_[80407]_ , \new_[80410]_ ,
    \new_[80413]_ , \new_[80414]_ , \new_[80417]_ , \new_[80420]_ ,
    \new_[80421]_ , \new_[80422]_ , \new_[80425]_ , \new_[80428]_ ,
    \new_[80429]_ , \new_[80432]_ , \new_[80435]_ , \new_[80436]_ ,
    \new_[80437]_ , \new_[80440]_ , \new_[80443]_ , \new_[80444]_ ,
    \new_[80447]_ , \new_[80450]_ , \new_[80451]_ , \new_[80452]_ ,
    \new_[80455]_ , \new_[80458]_ , \new_[80459]_ , \new_[80462]_ ,
    \new_[80465]_ , \new_[80466]_ , \new_[80467]_ , \new_[80470]_ ,
    \new_[80473]_ , \new_[80474]_ , \new_[80477]_ , \new_[80480]_ ,
    \new_[80481]_ , \new_[80482]_ , \new_[80485]_ , \new_[80488]_ ,
    \new_[80489]_ , \new_[80492]_ , \new_[80495]_ , \new_[80496]_ ,
    \new_[80497]_ , \new_[80500]_ , \new_[80503]_ , \new_[80504]_ ,
    \new_[80507]_ , \new_[80510]_ , \new_[80511]_ , \new_[80512]_ ,
    \new_[80515]_ , \new_[80518]_ , \new_[80519]_ , \new_[80522]_ ,
    \new_[80525]_ , \new_[80526]_ , \new_[80527]_ , \new_[80530]_ ,
    \new_[80533]_ , \new_[80534]_ , \new_[80537]_ , \new_[80540]_ ,
    \new_[80541]_ , \new_[80542]_ , \new_[80545]_ , \new_[80548]_ ,
    \new_[80549]_ , \new_[80552]_ , \new_[80555]_ , \new_[80556]_ ,
    \new_[80557]_ , \new_[80560]_ , \new_[80563]_ , \new_[80564]_ ,
    \new_[80567]_ , \new_[80570]_ , \new_[80571]_ , \new_[80572]_ ,
    \new_[80575]_ , \new_[80578]_ , \new_[80579]_ , \new_[80582]_ ,
    \new_[80585]_ , \new_[80586]_ , \new_[80587]_ , \new_[80590]_ ,
    \new_[80593]_ , \new_[80594]_ , \new_[80597]_ , \new_[80600]_ ,
    \new_[80601]_ , \new_[80602]_ , \new_[80605]_ , \new_[80608]_ ,
    \new_[80609]_ , \new_[80612]_ , \new_[80615]_ , \new_[80616]_ ,
    \new_[80617]_ , \new_[80620]_ , \new_[80623]_ , \new_[80624]_ ,
    \new_[80627]_ , \new_[80630]_ , \new_[80631]_ , \new_[80632]_ ,
    \new_[80635]_ , \new_[80638]_ , \new_[80639]_ , \new_[80642]_ ,
    \new_[80645]_ , \new_[80646]_ , \new_[80647]_ , \new_[80650]_ ,
    \new_[80653]_ , \new_[80654]_ , \new_[80657]_ , \new_[80660]_ ,
    \new_[80661]_ , \new_[80662]_ , \new_[80665]_ , \new_[80668]_ ,
    \new_[80669]_ , \new_[80672]_ , \new_[80675]_ , \new_[80676]_ ,
    \new_[80677]_ , \new_[80680]_ , \new_[80683]_ , \new_[80684]_ ,
    \new_[80687]_ , \new_[80690]_ , \new_[80691]_ , \new_[80692]_ ,
    \new_[80695]_ , \new_[80698]_ , \new_[80699]_ , \new_[80702]_ ,
    \new_[80705]_ , \new_[80706]_ , \new_[80707]_ , \new_[80710]_ ,
    \new_[80713]_ , \new_[80714]_ , \new_[80717]_ , \new_[80720]_ ,
    \new_[80721]_ , \new_[80722]_ , \new_[80725]_ , \new_[80728]_ ,
    \new_[80729]_ , \new_[80732]_ , \new_[80735]_ , \new_[80736]_ ,
    \new_[80737]_ , \new_[80740]_ , \new_[80743]_ , \new_[80744]_ ,
    \new_[80747]_ , \new_[80750]_ , \new_[80751]_ , \new_[80752]_ ,
    \new_[80755]_ , \new_[80758]_ , \new_[80759]_ , \new_[80762]_ ,
    \new_[80765]_ , \new_[80766]_ , \new_[80767]_ , \new_[80770]_ ,
    \new_[80773]_ , \new_[80774]_ , \new_[80777]_ , \new_[80780]_ ,
    \new_[80781]_ , \new_[80782]_ , \new_[80785]_ , \new_[80788]_ ,
    \new_[80789]_ , \new_[80792]_ , \new_[80795]_ , \new_[80796]_ ,
    \new_[80797]_ , \new_[80800]_ , \new_[80803]_ , \new_[80804]_ ,
    \new_[80807]_ , \new_[80810]_ , \new_[80811]_ , \new_[80812]_ ,
    \new_[80815]_ , \new_[80818]_ , \new_[80819]_ , \new_[80822]_ ,
    \new_[80825]_ , \new_[80826]_ , \new_[80827]_ , \new_[80830]_ ,
    \new_[80833]_ , \new_[80834]_ , \new_[80837]_ , \new_[80840]_ ,
    \new_[80841]_ , \new_[80842]_ , \new_[80845]_ , \new_[80848]_ ,
    \new_[80849]_ , \new_[80852]_ , \new_[80855]_ , \new_[80856]_ ,
    \new_[80857]_ , \new_[80860]_ , \new_[80863]_ , \new_[80864]_ ,
    \new_[80867]_ , \new_[80870]_ , \new_[80871]_ , \new_[80872]_ ,
    \new_[80875]_ , \new_[80878]_ , \new_[80879]_ , \new_[80882]_ ,
    \new_[80885]_ , \new_[80886]_ , \new_[80887]_ , \new_[80890]_ ,
    \new_[80893]_ , \new_[80894]_ , \new_[80897]_ , \new_[80900]_ ,
    \new_[80901]_ , \new_[80902]_ , \new_[80905]_ , \new_[80908]_ ,
    \new_[80909]_ , \new_[80912]_ , \new_[80915]_ , \new_[80916]_ ,
    \new_[80917]_ , \new_[80920]_ , \new_[80923]_ , \new_[80924]_ ,
    \new_[80927]_ , \new_[80930]_ , \new_[80931]_ , \new_[80932]_ ,
    \new_[80935]_ , \new_[80938]_ , \new_[80939]_ , \new_[80942]_ ,
    \new_[80945]_ , \new_[80946]_ , \new_[80947]_ , \new_[80950]_ ,
    \new_[80953]_ , \new_[80954]_ , \new_[80957]_ , \new_[80960]_ ,
    \new_[80961]_ , \new_[80962]_ , \new_[80965]_ , \new_[80968]_ ,
    \new_[80969]_ , \new_[80972]_ , \new_[80975]_ , \new_[80976]_ ,
    \new_[80977]_ , \new_[80980]_ , \new_[80983]_ , \new_[80984]_ ,
    \new_[80987]_ , \new_[80990]_ , \new_[80991]_ , \new_[80992]_ ,
    \new_[80995]_ , \new_[80998]_ , \new_[80999]_ , \new_[81002]_ ,
    \new_[81005]_ , \new_[81006]_ , \new_[81007]_ , \new_[81010]_ ,
    \new_[81013]_ , \new_[81014]_ , \new_[81017]_ , \new_[81020]_ ,
    \new_[81021]_ , \new_[81022]_ , \new_[81025]_ , \new_[81028]_ ,
    \new_[81029]_ , \new_[81032]_ , \new_[81035]_ , \new_[81036]_ ,
    \new_[81037]_ , \new_[81040]_ , \new_[81043]_ , \new_[81044]_ ,
    \new_[81047]_ , \new_[81050]_ , \new_[81051]_ , \new_[81052]_ ,
    \new_[81055]_ , \new_[81058]_ , \new_[81059]_ , \new_[81062]_ ,
    \new_[81065]_ , \new_[81066]_ , \new_[81067]_ , \new_[81070]_ ,
    \new_[81073]_ , \new_[81074]_ , \new_[81077]_ , \new_[81080]_ ,
    \new_[81081]_ , \new_[81082]_ , \new_[81085]_ , \new_[81088]_ ,
    \new_[81089]_ , \new_[81092]_ , \new_[81095]_ , \new_[81096]_ ,
    \new_[81097]_ , \new_[81100]_ , \new_[81103]_ , \new_[81104]_ ,
    \new_[81107]_ , \new_[81110]_ , \new_[81111]_ , \new_[81112]_ ,
    \new_[81115]_ , \new_[81118]_ , \new_[81119]_ , \new_[81122]_ ,
    \new_[81125]_ , \new_[81126]_ , \new_[81127]_ , \new_[81130]_ ,
    \new_[81133]_ , \new_[81134]_ , \new_[81137]_ , \new_[81140]_ ,
    \new_[81141]_ , \new_[81142]_ , \new_[81145]_ , \new_[81148]_ ,
    \new_[81149]_ , \new_[81152]_ , \new_[81155]_ , \new_[81156]_ ,
    \new_[81157]_ , \new_[81160]_ , \new_[81163]_ , \new_[81164]_ ,
    \new_[81167]_ , \new_[81170]_ , \new_[81171]_ , \new_[81172]_ ,
    \new_[81175]_ , \new_[81178]_ , \new_[81179]_ , \new_[81182]_ ,
    \new_[81185]_ , \new_[81186]_ , \new_[81187]_ , \new_[81190]_ ,
    \new_[81193]_ , \new_[81194]_ , \new_[81197]_ , \new_[81200]_ ,
    \new_[81201]_ , \new_[81202]_ , \new_[81205]_ , \new_[81208]_ ,
    \new_[81209]_ , \new_[81212]_ , \new_[81215]_ , \new_[81216]_ ,
    \new_[81217]_ , \new_[81220]_ , \new_[81223]_ , \new_[81224]_ ,
    \new_[81227]_ , \new_[81230]_ , \new_[81231]_ , \new_[81232]_ ,
    \new_[81235]_ , \new_[81238]_ , \new_[81239]_ , \new_[81242]_ ,
    \new_[81245]_ , \new_[81246]_ , \new_[81247]_ , \new_[81250]_ ,
    \new_[81253]_ , \new_[81254]_ , \new_[81257]_ , \new_[81260]_ ,
    \new_[81261]_ , \new_[81262]_ , \new_[81265]_ , \new_[81268]_ ,
    \new_[81269]_ , \new_[81272]_ , \new_[81275]_ , \new_[81276]_ ,
    \new_[81277]_ , \new_[81280]_ , \new_[81283]_ , \new_[81284]_ ,
    \new_[81287]_ , \new_[81290]_ , \new_[81291]_ , \new_[81292]_ ,
    \new_[81295]_ , \new_[81298]_ , \new_[81299]_ , \new_[81302]_ ,
    \new_[81305]_ , \new_[81306]_ , \new_[81307]_ , \new_[81310]_ ,
    \new_[81313]_ , \new_[81314]_ , \new_[81317]_ , \new_[81320]_ ,
    \new_[81321]_ , \new_[81322]_ , \new_[81325]_ , \new_[81328]_ ,
    \new_[81329]_ , \new_[81332]_ , \new_[81335]_ , \new_[81336]_ ,
    \new_[81337]_ , \new_[81340]_ , \new_[81343]_ , \new_[81344]_ ,
    \new_[81347]_ , \new_[81350]_ , \new_[81351]_ , \new_[81352]_ ,
    \new_[81355]_ , \new_[81358]_ , \new_[81359]_ , \new_[81362]_ ,
    \new_[81365]_ , \new_[81366]_ , \new_[81367]_ , \new_[81370]_ ,
    \new_[81373]_ , \new_[81374]_ , \new_[81377]_ , \new_[81380]_ ,
    \new_[81381]_ , \new_[81382]_ , \new_[81385]_ , \new_[81388]_ ,
    \new_[81389]_ , \new_[81392]_ , \new_[81395]_ , \new_[81396]_ ,
    \new_[81397]_ , \new_[81400]_ , \new_[81403]_ , \new_[81404]_ ,
    \new_[81407]_ , \new_[81410]_ , \new_[81411]_ , \new_[81412]_ ,
    \new_[81415]_ , \new_[81418]_ , \new_[81419]_ , \new_[81422]_ ,
    \new_[81425]_ , \new_[81426]_ , \new_[81427]_ , \new_[81430]_ ,
    \new_[81433]_ , \new_[81434]_ , \new_[81437]_ , \new_[81440]_ ,
    \new_[81441]_ , \new_[81442]_ , \new_[81445]_ , \new_[81448]_ ,
    \new_[81449]_ , \new_[81452]_ , \new_[81455]_ , \new_[81456]_ ,
    \new_[81457]_ , \new_[81460]_ , \new_[81463]_ , \new_[81464]_ ,
    \new_[81467]_ , \new_[81470]_ , \new_[81471]_ , \new_[81472]_ ,
    \new_[81475]_ , \new_[81478]_ , \new_[81479]_ , \new_[81482]_ ,
    \new_[81485]_ , \new_[81486]_ , \new_[81487]_ , \new_[81490]_ ,
    \new_[81493]_ , \new_[81494]_ , \new_[81497]_ , \new_[81500]_ ,
    \new_[81501]_ , \new_[81502]_ , \new_[81505]_ , \new_[81508]_ ,
    \new_[81509]_ , \new_[81512]_ , \new_[81515]_ , \new_[81516]_ ,
    \new_[81517]_ , \new_[81520]_ , \new_[81523]_ , \new_[81524]_ ,
    \new_[81527]_ , \new_[81530]_ , \new_[81531]_ , \new_[81532]_ ,
    \new_[81535]_ , \new_[81538]_ , \new_[81539]_ , \new_[81542]_ ,
    \new_[81545]_ , \new_[81546]_ , \new_[81547]_ , \new_[81550]_ ,
    \new_[81553]_ , \new_[81554]_ , \new_[81557]_ , \new_[81560]_ ,
    \new_[81561]_ , \new_[81562]_ , \new_[81565]_ , \new_[81568]_ ,
    \new_[81569]_ , \new_[81572]_ , \new_[81575]_ , \new_[81576]_ ,
    \new_[81577]_ , \new_[81580]_ , \new_[81583]_ , \new_[81584]_ ,
    \new_[81587]_ , \new_[81590]_ , \new_[81591]_ , \new_[81592]_ ,
    \new_[81595]_ , \new_[81598]_ , \new_[81599]_ , \new_[81602]_ ,
    \new_[81605]_ , \new_[81606]_ , \new_[81607]_ , \new_[81610]_ ,
    \new_[81613]_ , \new_[81614]_ , \new_[81617]_ , \new_[81620]_ ,
    \new_[81621]_ , \new_[81622]_ , \new_[81625]_ , \new_[81628]_ ,
    \new_[81629]_ , \new_[81632]_ , \new_[81635]_ , \new_[81636]_ ,
    \new_[81637]_ , \new_[81640]_ , \new_[81643]_ , \new_[81644]_ ,
    \new_[81647]_ , \new_[81650]_ , \new_[81651]_ , \new_[81652]_ ,
    \new_[81655]_ , \new_[81658]_ , \new_[81659]_ , \new_[81662]_ ,
    \new_[81665]_ , \new_[81666]_ , \new_[81667]_ , \new_[81670]_ ,
    \new_[81673]_ , \new_[81674]_ , \new_[81677]_ , \new_[81680]_ ,
    \new_[81681]_ , \new_[81682]_ , \new_[81685]_ , \new_[81688]_ ,
    \new_[81689]_ , \new_[81692]_ , \new_[81695]_ , \new_[81696]_ ,
    \new_[81697]_ , \new_[81700]_ , \new_[81703]_ , \new_[81704]_ ,
    \new_[81707]_ , \new_[81710]_ , \new_[81711]_ , \new_[81712]_ ,
    \new_[81715]_ , \new_[81718]_ , \new_[81719]_ , \new_[81722]_ ,
    \new_[81725]_ , \new_[81726]_ , \new_[81727]_ , \new_[81730]_ ,
    \new_[81733]_ , \new_[81734]_ , \new_[81737]_ , \new_[81740]_ ,
    \new_[81741]_ , \new_[81742]_ , \new_[81745]_ , \new_[81748]_ ,
    \new_[81749]_ , \new_[81752]_ , \new_[81755]_ , \new_[81756]_ ,
    \new_[81757]_ , \new_[81760]_ , \new_[81763]_ , \new_[81764]_ ,
    \new_[81767]_ , \new_[81770]_ , \new_[81771]_ , \new_[81772]_ ,
    \new_[81775]_ , \new_[81778]_ , \new_[81779]_ , \new_[81782]_ ,
    \new_[81785]_ , \new_[81786]_ , \new_[81787]_ , \new_[81790]_ ,
    \new_[81793]_ , \new_[81794]_ , \new_[81797]_ , \new_[81800]_ ,
    \new_[81801]_ , \new_[81802]_ , \new_[81805]_ , \new_[81808]_ ,
    \new_[81809]_ , \new_[81812]_ , \new_[81815]_ , \new_[81816]_ ,
    \new_[81817]_ , \new_[81820]_ , \new_[81823]_ , \new_[81824]_ ,
    \new_[81827]_ , \new_[81830]_ , \new_[81831]_ , \new_[81832]_ ,
    \new_[81835]_ , \new_[81838]_ , \new_[81839]_ , \new_[81842]_ ,
    \new_[81845]_ , \new_[81846]_ , \new_[81847]_ , \new_[81850]_ ,
    \new_[81853]_ , \new_[81854]_ , \new_[81857]_ , \new_[81860]_ ,
    \new_[81861]_ , \new_[81862]_ , \new_[81865]_ , \new_[81868]_ ,
    \new_[81869]_ , \new_[81872]_ , \new_[81875]_ , \new_[81876]_ ,
    \new_[81877]_ , \new_[81880]_ , \new_[81883]_ , \new_[81884]_ ,
    \new_[81887]_ , \new_[81890]_ , \new_[81891]_ , \new_[81892]_ ,
    \new_[81895]_ , \new_[81898]_ , \new_[81899]_ , \new_[81902]_ ,
    \new_[81905]_ , \new_[81906]_ , \new_[81907]_ , \new_[81910]_ ,
    \new_[81913]_ , \new_[81914]_ , \new_[81917]_ , \new_[81920]_ ,
    \new_[81921]_ , \new_[81922]_ , \new_[81925]_ , \new_[81928]_ ,
    \new_[81929]_ , \new_[81932]_ , \new_[81935]_ , \new_[81936]_ ,
    \new_[81937]_ , \new_[81940]_ , \new_[81943]_ , \new_[81944]_ ,
    \new_[81947]_ , \new_[81950]_ , \new_[81951]_ , \new_[81952]_ ,
    \new_[81955]_ , \new_[81958]_ , \new_[81959]_ , \new_[81962]_ ,
    \new_[81965]_ , \new_[81966]_ , \new_[81967]_ , \new_[81970]_ ,
    \new_[81973]_ , \new_[81974]_ , \new_[81977]_ , \new_[81980]_ ,
    \new_[81981]_ , \new_[81982]_ , \new_[81985]_ , \new_[81988]_ ,
    \new_[81989]_ , \new_[81992]_ , \new_[81995]_ , \new_[81996]_ ,
    \new_[81997]_ , \new_[82000]_ , \new_[82003]_ , \new_[82004]_ ,
    \new_[82007]_ , \new_[82010]_ , \new_[82011]_ , \new_[82012]_ ,
    \new_[82015]_ , \new_[82018]_ , \new_[82019]_ , \new_[82022]_ ,
    \new_[82025]_ , \new_[82026]_ , \new_[82027]_ , \new_[82030]_ ,
    \new_[82033]_ , \new_[82034]_ , \new_[82037]_ , \new_[82040]_ ,
    \new_[82041]_ , \new_[82042]_ , \new_[82045]_ , \new_[82048]_ ,
    \new_[82049]_ , \new_[82052]_ , \new_[82055]_ , \new_[82056]_ ,
    \new_[82057]_ , \new_[82060]_ , \new_[82063]_ , \new_[82064]_ ,
    \new_[82067]_ , \new_[82070]_ , \new_[82071]_ , \new_[82072]_ ,
    \new_[82075]_ , \new_[82078]_ , \new_[82079]_ , \new_[82082]_ ,
    \new_[82085]_ , \new_[82086]_ , \new_[82087]_ , \new_[82090]_ ,
    \new_[82093]_ , \new_[82094]_ , \new_[82097]_ , \new_[82100]_ ,
    \new_[82101]_ , \new_[82102]_ , \new_[82105]_ , \new_[82108]_ ,
    \new_[82109]_ , \new_[82112]_ , \new_[82115]_ , \new_[82116]_ ,
    \new_[82117]_ , \new_[82120]_ , \new_[82123]_ , \new_[82124]_ ,
    \new_[82127]_ , \new_[82130]_ , \new_[82131]_ , \new_[82132]_ ,
    \new_[82135]_ , \new_[82138]_ , \new_[82139]_ , \new_[82142]_ ,
    \new_[82145]_ , \new_[82146]_ , \new_[82147]_ , \new_[82150]_ ,
    \new_[82153]_ , \new_[82154]_ , \new_[82157]_ , \new_[82160]_ ,
    \new_[82161]_ , \new_[82162]_ , \new_[82165]_ , \new_[82168]_ ,
    \new_[82169]_ , \new_[82172]_ , \new_[82175]_ , \new_[82176]_ ,
    \new_[82177]_ , \new_[82180]_ , \new_[82183]_ , \new_[82184]_ ,
    \new_[82187]_ , \new_[82190]_ , \new_[82191]_ , \new_[82192]_ ,
    \new_[82195]_ , \new_[82198]_ , \new_[82199]_ , \new_[82202]_ ,
    \new_[82205]_ , \new_[82206]_ , \new_[82207]_ , \new_[82210]_ ,
    \new_[82213]_ , \new_[82214]_ , \new_[82217]_ , \new_[82220]_ ,
    \new_[82221]_ , \new_[82222]_ , \new_[82225]_ , \new_[82228]_ ,
    \new_[82229]_ , \new_[82232]_ , \new_[82235]_ , \new_[82236]_ ,
    \new_[82237]_ , \new_[82240]_ , \new_[82243]_ , \new_[82244]_ ,
    \new_[82247]_ , \new_[82250]_ , \new_[82251]_ , \new_[82252]_ ,
    \new_[82255]_ , \new_[82258]_ , \new_[82259]_ , \new_[82262]_ ,
    \new_[82265]_ , \new_[82266]_ , \new_[82267]_ , \new_[82270]_ ,
    \new_[82273]_ , \new_[82274]_ , \new_[82277]_ , \new_[82280]_ ,
    \new_[82281]_ , \new_[82282]_ , \new_[82285]_ , \new_[82288]_ ,
    \new_[82289]_ , \new_[82292]_ , \new_[82295]_ , \new_[82296]_ ,
    \new_[82297]_ , \new_[82300]_ , \new_[82303]_ , \new_[82304]_ ,
    \new_[82307]_ , \new_[82310]_ , \new_[82311]_ , \new_[82312]_ ,
    \new_[82315]_ , \new_[82318]_ , \new_[82319]_ , \new_[82322]_ ,
    \new_[82325]_ , \new_[82326]_ , \new_[82327]_ , \new_[82330]_ ,
    \new_[82333]_ , \new_[82334]_ , \new_[82337]_ , \new_[82340]_ ,
    \new_[82341]_ , \new_[82342]_ , \new_[82345]_ , \new_[82348]_ ,
    \new_[82349]_ , \new_[82352]_ , \new_[82355]_ , \new_[82356]_ ,
    \new_[82357]_ , \new_[82360]_ , \new_[82363]_ , \new_[82364]_ ,
    \new_[82367]_ , \new_[82370]_ , \new_[82371]_ , \new_[82372]_ ,
    \new_[82375]_ , \new_[82378]_ , \new_[82379]_ , \new_[82382]_ ,
    \new_[82385]_ , \new_[82386]_ , \new_[82387]_ , \new_[82390]_ ,
    \new_[82393]_ , \new_[82394]_ , \new_[82397]_ , \new_[82400]_ ,
    \new_[82401]_ , \new_[82402]_ , \new_[82405]_ , \new_[82408]_ ,
    \new_[82409]_ , \new_[82412]_ , \new_[82415]_ , \new_[82416]_ ,
    \new_[82417]_ , \new_[82420]_ , \new_[82423]_ , \new_[82424]_ ,
    \new_[82427]_ , \new_[82430]_ , \new_[82431]_ , \new_[82432]_ ,
    \new_[82435]_ , \new_[82438]_ , \new_[82439]_ , \new_[82442]_ ,
    \new_[82445]_ , \new_[82446]_ , \new_[82447]_ , \new_[82450]_ ,
    \new_[82453]_ , \new_[82454]_ , \new_[82457]_ , \new_[82460]_ ,
    \new_[82461]_ , \new_[82462]_ , \new_[82465]_ , \new_[82468]_ ,
    \new_[82469]_ , \new_[82472]_ , \new_[82475]_ , \new_[82476]_ ,
    \new_[82477]_ , \new_[82480]_ , \new_[82483]_ , \new_[82484]_ ,
    \new_[82487]_ , \new_[82490]_ , \new_[82491]_ , \new_[82492]_ ,
    \new_[82495]_ , \new_[82498]_ , \new_[82499]_ , \new_[82502]_ ,
    \new_[82505]_ , \new_[82506]_ , \new_[82507]_ , \new_[82510]_ ,
    \new_[82513]_ , \new_[82514]_ , \new_[82517]_ , \new_[82520]_ ,
    \new_[82521]_ , \new_[82522]_ , \new_[82525]_ , \new_[82528]_ ,
    \new_[82529]_ , \new_[82532]_ , \new_[82535]_ , \new_[82536]_ ,
    \new_[82537]_ , \new_[82540]_ , \new_[82543]_ , \new_[82544]_ ,
    \new_[82547]_ , \new_[82550]_ , \new_[82551]_ , \new_[82552]_ ,
    \new_[82555]_ , \new_[82558]_ , \new_[82559]_ , \new_[82562]_ ,
    \new_[82565]_ , \new_[82566]_ , \new_[82567]_ , \new_[82570]_ ,
    \new_[82573]_ , \new_[82574]_ , \new_[82577]_ , \new_[82580]_ ,
    \new_[82581]_ , \new_[82582]_ , \new_[82585]_ , \new_[82588]_ ,
    \new_[82589]_ , \new_[82592]_ , \new_[82595]_ , \new_[82596]_ ,
    \new_[82597]_ , \new_[82600]_ , \new_[82603]_ , \new_[82604]_ ,
    \new_[82607]_ , \new_[82610]_ , \new_[82611]_ , \new_[82612]_ ,
    \new_[82615]_ , \new_[82618]_ , \new_[82619]_ , \new_[82622]_ ,
    \new_[82625]_ , \new_[82626]_ , \new_[82627]_ , \new_[82630]_ ,
    \new_[82633]_ , \new_[82634]_ , \new_[82637]_ , \new_[82640]_ ,
    \new_[82641]_ , \new_[82642]_ , \new_[82645]_ , \new_[82648]_ ,
    \new_[82649]_ , \new_[82652]_ , \new_[82655]_ , \new_[82656]_ ,
    \new_[82657]_ , \new_[82660]_ , \new_[82663]_ , \new_[82664]_ ,
    \new_[82667]_ , \new_[82670]_ , \new_[82671]_ , \new_[82672]_ ,
    \new_[82675]_ , \new_[82678]_ , \new_[82679]_ , \new_[82682]_ ,
    \new_[82685]_ , \new_[82686]_ , \new_[82687]_ , \new_[82690]_ ,
    \new_[82693]_ , \new_[82694]_ , \new_[82697]_ , \new_[82700]_ ,
    \new_[82701]_ , \new_[82702]_ , \new_[82705]_ , \new_[82708]_ ,
    \new_[82709]_ , \new_[82712]_ , \new_[82715]_ , \new_[82716]_ ,
    \new_[82717]_ , \new_[82720]_ , \new_[82723]_ , \new_[82724]_ ,
    \new_[82727]_ , \new_[82730]_ , \new_[82731]_ , \new_[82732]_ ,
    \new_[82735]_ , \new_[82738]_ , \new_[82739]_ , \new_[82742]_ ,
    \new_[82745]_ , \new_[82746]_ , \new_[82747]_ , \new_[82750]_ ,
    \new_[82753]_ , \new_[82754]_ , \new_[82757]_ , \new_[82760]_ ,
    \new_[82761]_ , \new_[82762]_ , \new_[82765]_ , \new_[82768]_ ,
    \new_[82769]_ , \new_[82772]_ , \new_[82775]_ , \new_[82776]_ ,
    \new_[82777]_ , \new_[82780]_ , \new_[82783]_ , \new_[82784]_ ,
    \new_[82787]_ , \new_[82790]_ , \new_[82791]_ , \new_[82792]_ ,
    \new_[82795]_ , \new_[82798]_ , \new_[82799]_ , \new_[82802]_ ,
    \new_[82805]_ , \new_[82806]_ , \new_[82807]_ , \new_[82810]_ ,
    \new_[82813]_ , \new_[82814]_ , \new_[82817]_ , \new_[82820]_ ,
    \new_[82821]_ , \new_[82822]_ , \new_[82825]_ , \new_[82828]_ ,
    \new_[82829]_ , \new_[82832]_ , \new_[82835]_ , \new_[82836]_ ,
    \new_[82837]_ , \new_[82840]_ , \new_[82843]_ , \new_[82844]_ ,
    \new_[82847]_ , \new_[82850]_ , \new_[82851]_ , \new_[82852]_ ,
    \new_[82855]_ , \new_[82858]_ , \new_[82859]_ , \new_[82862]_ ,
    \new_[82865]_ , \new_[82866]_ , \new_[82867]_ , \new_[82870]_ ,
    \new_[82873]_ , \new_[82874]_ , \new_[82877]_ , \new_[82880]_ ,
    \new_[82881]_ , \new_[82882]_ , \new_[82885]_ , \new_[82888]_ ,
    \new_[82889]_ , \new_[82892]_ , \new_[82895]_ , \new_[82896]_ ,
    \new_[82897]_ , \new_[82900]_ , \new_[82903]_ , \new_[82904]_ ,
    \new_[82907]_ , \new_[82910]_ , \new_[82911]_ , \new_[82912]_ ,
    \new_[82915]_ , \new_[82918]_ , \new_[82919]_ , \new_[82922]_ ,
    \new_[82925]_ , \new_[82926]_ , \new_[82927]_ , \new_[82930]_ ,
    \new_[82933]_ , \new_[82934]_ , \new_[82937]_ , \new_[82940]_ ,
    \new_[82941]_ , \new_[82942]_ , \new_[82945]_ , \new_[82948]_ ,
    \new_[82949]_ , \new_[82952]_ , \new_[82955]_ , \new_[82956]_ ,
    \new_[82957]_ , \new_[82960]_ , \new_[82963]_ , \new_[82964]_ ,
    \new_[82967]_ , \new_[82970]_ , \new_[82971]_ , \new_[82972]_ ,
    \new_[82975]_ , \new_[82978]_ , \new_[82979]_ , \new_[82982]_ ,
    \new_[82985]_ , \new_[82986]_ , \new_[82987]_ , \new_[82990]_ ,
    \new_[82993]_ , \new_[82994]_ , \new_[82997]_ , \new_[83000]_ ,
    \new_[83001]_ , \new_[83002]_ , \new_[83005]_ , \new_[83008]_ ,
    \new_[83009]_ , \new_[83012]_ , \new_[83015]_ , \new_[83016]_ ,
    \new_[83017]_ , \new_[83020]_ , \new_[83023]_ , \new_[83024]_ ,
    \new_[83027]_ , \new_[83030]_ , \new_[83031]_ , \new_[83032]_ ,
    \new_[83035]_ , \new_[83038]_ , \new_[83039]_ , \new_[83042]_ ,
    \new_[83045]_ , \new_[83046]_ , \new_[83047]_ , \new_[83050]_ ,
    \new_[83053]_ , \new_[83054]_ , \new_[83057]_ , \new_[83060]_ ,
    \new_[83061]_ , \new_[83062]_ , \new_[83065]_ , \new_[83068]_ ,
    \new_[83069]_ , \new_[83072]_ , \new_[83075]_ , \new_[83076]_ ,
    \new_[83077]_ , \new_[83080]_ , \new_[83083]_ , \new_[83084]_ ,
    \new_[83087]_ , \new_[83090]_ , \new_[83091]_ , \new_[83092]_ ,
    \new_[83095]_ , \new_[83098]_ , \new_[83099]_ , \new_[83102]_ ,
    \new_[83105]_ , \new_[83106]_ , \new_[83107]_ , \new_[83110]_ ,
    \new_[83113]_ , \new_[83114]_ , \new_[83117]_ , \new_[83120]_ ,
    \new_[83121]_ , \new_[83122]_ , \new_[83125]_ , \new_[83128]_ ,
    \new_[83129]_ , \new_[83132]_ , \new_[83135]_ , \new_[83136]_ ,
    \new_[83137]_ , \new_[83140]_ , \new_[83143]_ , \new_[83144]_ ,
    \new_[83147]_ , \new_[83150]_ , \new_[83151]_ , \new_[83152]_ ,
    \new_[83155]_ , \new_[83158]_ , \new_[83159]_ , \new_[83162]_ ,
    \new_[83165]_ , \new_[83166]_ , \new_[83167]_ , \new_[83170]_ ,
    \new_[83173]_ , \new_[83174]_ , \new_[83177]_ , \new_[83180]_ ,
    \new_[83181]_ , \new_[83182]_ , \new_[83185]_ , \new_[83188]_ ,
    \new_[83189]_ , \new_[83192]_ , \new_[83195]_ , \new_[83196]_ ,
    \new_[83197]_ , \new_[83200]_ , \new_[83203]_ , \new_[83204]_ ,
    \new_[83207]_ , \new_[83210]_ , \new_[83211]_ , \new_[83212]_ ,
    \new_[83215]_ , \new_[83218]_ , \new_[83219]_ , \new_[83222]_ ,
    \new_[83225]_ , \new_[83226]_ , \new_[83227]_ , \new_[83230]_ ,
    \new_[83233]_ , \new_[83234]_ , \new_[83237]_ , \new_[83240]_ ,
    \new_[83241]_ , \new_[83242]_ , \new_[83245]_ , \new_[83248]_ ,
    \new_[83249]_ , \new_[83252]_ , \new_[83255]_ , \new_[83256]_ ,
    \new_[83257]_ , \new_[83260]_ , \new_[83263]_ , \new_[83264]_ ,
    \new_[83267]_ , \new_[83270]_ , \new_[83271]_ , \new_[83272]_ ,
    \new_[83275]_ , \new_[83278]_ , \new_[83279]_ , \new_[83282]_ ,
    \new_[83285]_ , \new_[83286]_ , \new_[83287]_ , \new_[83290]_ ,
    \new_[83293]_ , \new_[83294]_ , \new_[83297]_ , \new_[83300]_ ,
    \new_[83301]_ , \new_[83302]_ , \new_[83305]_ , \new_[83308]_ ,
    \new_[83309]_ , \new_[83312]_ , \new_[83315]_ , \new_[83316]_ ,
    \new_[83317]_ , \new_[83320]_ , \new_[83323]_ , \new_[83324]_ ,
    \new_[83327]_ , \new_[83330]_ , \new_[83331]_ , \new_[83332]_ ,
    \new_[83335]_ , \new_[83338]_ , \new_[83339]_ , \new_[83342]_ ,
    \new_[83345]_ , \new_[83346]_ , \new_[83347]_ , \new_[83350]_ ,
    \new_[83353]_ , \new_[83354]_ , \new_[83357]_ , \new_[83360]_ ,
    \new_[83361]_ , \new_[83362]_ , \new_[83365]_ , \new_[83368]_ ,
    \new_[83369]_ , \new_[83372]_ , \new_[83375]_ , \new_[83376]_ ,
    \new_[83377]_ , \new_[83380]_ , \new_[83383]_ , \new_[83384]_ ,
    \new_[83387]_ , \new_[83390]_ , \new_[83391]_ , \new_[83392]_ ,
    \new_[83395]_ , \new_[83398]_ , \new_[83399]_ , \new_[83402]_ ,
    \new_[83405]_ , \new_[83406]_ , \new_[83407]_ , \new_[83410]_ ,
    \new_[83413]_ , \new_[83414]_ , \new_[83417]_ , \new_[83420]_ ,
    \new_[83421]_ , \new_[83422]_ , \new_[83425]_ , \new_[83428]_ ,
    \new_[83429]_ , \new_[83432]_ , \new_[83435]_ , \new_[83436]_ ,
    \new_[83437]_ , \new_[83440]_ , \new_[83443]_ , \new_[83444]_ ,
    \new_[83447]_ , \new_[83450]_ , \new_[83451]_ , \new_[83452]_ ,
    \new_[83455]_ , \new_[83458]_ , \new_[83459]_ , \new_[83462]_ ,
    \new_[83465]_ , \new_[83466]_ , \new_[83467]_ , \new_[83470]_ ,
    \new_[83473]_ , \new_[83474]_ , \new_[83477]_ , \new_[83480]_ ,
    \new_[83481]_ , \new_[83482]_ , \new_[83485]_ , \new_[83488]_ ,
    \new_[83489]_ , \new_[83492]_ , \new_[83495]_ , \new_[83496]_ ,
    \new_[83497]_ , \new_[83500]_ , \new_[83503]_ , \new_[83504]_ ,
    \new_[83507]_ , \new_[83510]_ , \new_[83511]_ , \new_[83512]_ ,
    \new_[83515]_ , \new_[83518]_ , \new_[83519]_ , \new_[83522]_ ,
    \new_[83525]_ , \new_[83526]_ , \new_[83527]_ , \new_[83530]_ ,
    \new_[83533]_ , \new_[83534]_ , \new_[83537]_ , \new_[83540]_ ,
    \new_[83541]_ , \new_[83542]_ , \new_[83545]_ , \new_[83548]_ ,
    \new_[83549]_ , \new_[83552]_ , \new_[83555]_ , \new_[83556]_ ,
    \new_[83557]_ , \new_[83560]_ , \new_[83563]_ , \new_[83564]_ ,
    \new_[83567]_ , \new_[83570]_ , \new_[83571]_ , \new_[83572]_ ,
    \new_[83575]_ , \new_[83578]_ , \new_[83579]_ , \new_[83582]_ ,
    \new_[83585]_ , \new_[83586]_ , \new_[83587]_ , \new_[83590]_ ,
    \new_[83593]_ , \new_[83594]_ , \new_[83597]_ , \new_[83600]_ ,
    \new_[83601]_ , \new_[83602]_ , \new_[83605]_ , \new_[83608]_ ,
    \new_[83609]_ , \new_[83612]_ , \new_[83615]_ , \new_[83616]_ ,
    \new_[83617]_ , \new_[83620]_ , \new_[83623]_ , \new_[83624]_ ,
    \new_[83627]_ , \new_[83630]_ , \new_[83631]_ , \new_[83632]_ ,
    \new_[83635]_ , \new_[83638]_ , \new_[83639]_ , \new_[83642]_ ,
    \new_[83645]_ , \new_[83646]_ , \new_[83647]_ , \new_[83650]_ ,
    \new_[83653]_ , \new_[83654]_ , \new_[83657]_ , \new_[83660]_ ,
    \new_[83661]_ , \new_[83662]_ , \new_[83665]_ , \new_[83668]_ ,
    \new_[83669]_ , \new_[83672]_ , \new_[83675]_ , \new_[83676]_ ,
    \new_[83677]_ , \new_[83680]_ , \new_[83683]_ , \new_[83684]_ ,
    \new_[83687]_ , \new_[83690]_ , \new_[83691]_ , \new_[83692]_ ,
    \new_[83695]_ , \new_[83698]_ , \new_[83699]_ , \new_[83702]_ ,
    \new_[83705]_ , \new_[83706]_ , \new_[83707]_ , \new_[83710]_ ,
    \new_[83713]_ , \new_[83714]_ , \new_[83717]_ , \new_[83720]_ ,
    \new_[83721]_ , \new_[83722]_ , \new_[83725]_ , \new_[83728]_ ,
    \new_[83729]_ , \new_[83732]_ , \new_[83735]_ , \new_[83736]_ ,
    \new_[83737]_ , \new_[83740]_ , \new_[83743]_ , \new_[83744]_ ,
    \new_[83747]_ , \new_[83750]_ , \new_[83751]_ , \new_[83752]_ ,
    \new_[83755]_ , \new_[83758]_ , \new_[83759]_ , \new_[83762]_ ,
    \new_[83765]_ , \new_[83766]_ , \new_[83767]_ , \new_[83770]_ ,
    \new_[83773]_ , \new_[83774]_ , \new_[83777]_ , \new_[83780]_ ,
    \new_[83781]_ , \new_[83782]_ , \new_[83785]_ , \new_[83788]_ ,
    \new_[83789]_ , \new_[83792]_ , \new_[83795]_ , \new_[83796]_ ,
    \new_[83797]_ , \new_[83800]_ , \new_[83803]_ , \new_[83804]_ ,
    \new_[83807]_ , \new_[83810]_ , \new_[83811]_ , \new_[83812]_ ,
    \new_[83815]_ , \new_[83818]_ , \new_[83819]_ , \new_[83822]_ ,
    \new_[83825]_ , \new_[83826]_ , \new_[83827]_ , \new_[83830]_ ,
    \new_[83833]_ , \new_[83834]_ , \new_[83837]_ , \new_[83840]_ ,
    \new_[83841]_ , \new_[83842]_ , \new_[83845]_ , \new_[83848]_ ,
    \new_[83849]_ , \new_[83852]_ , \new_[83855]_ , \new_[83856]_ ,
    \new_[83857]_ , \new_[83860]_ , \new_[83863]_ , \new_[83864]_ ,
    \new_[83867]_ , \new_[83870]_ , \new_[83871]_ , \new_[83872]_ ,
    \new_[83875]_ , \new_[83878]_ , \new_[83879]_ , \new_[83882]_ ,
    \new_[83885]_ , \new_[83886]_ , \new_[83887]_ , \new_[83890]_ ,
    \new_[83893]_ , \new_[83894]_ , \new_[83897]_ , \new_[83900]_ ,
    \new_[83901]_ , \new_[83902]_ , \new_[83905]_ , \new_[83908]_ ,
    \new_[83909]_ , \new_[83912]_ , \new_[83915]_ , \new_[83916]_ ,
    \new_[83917]_ , \new_[83920]_ , \new_[83923]_ , \new_[83924]_ ,
    \new_[83927]_ , \new_[83930]_ , \new_[83931]_ , \new_[83932]_ ,
    \new_[83935]_ , \new_[83938]_ , \new_[83939]_ , \new_[83942]_ ,
    \new_[83945]_ , \new_[83946]_ , \new_[83947]_ , \new_[83950]_ ,
    \new_[83953]_ , \new_[83954]_ , \new_[83957]_ , \new_[83960]_ ,
    \new_[83961]_ , \new_[83962]_ , \new_[83965]_ , \new_[83968]_ ,
    \new_[83969]_ , \new_[83972]_ , \new_[83975]_ , \new_[83976]_ ,
    \new_[83977]_ , \new_[83980]_ , \new_[83983]_ , \new_[83984]_ ,
    \new_[83987]_ , \new_[83990]_ , \new_[83991]_ , \new_[83992]_ ,
    \new_[83995]_ , \new_[83998]_ , \new_[83999]_ , \new_[84002]_ ,
    \new_[84005]_ , \new_[84006]_ , \new_[84007]_ , \new_[84010]_ ,
    \new_[84013]_ , \new_[84014]_ , \new_[84017]_ , \new_[84020]_ ,
    \new_[84021]_ , \new_[84022]_ , \new_[84025]_ , \new_[84028]_ ,
    \new_[84029]_ , \new_[84032]_ , \new_[84035]_ , \new_[84036]_ ,
    \new_[84037]_ , \new_[84040]_ , \new_[84043]_ , \new_[84044]_ ,
    \new_[84047]_ , \new_[84050]_ , \new_[84051]_ , \new_[84052]_ ,
    \new_[84055]_ , \new_[84058]_ , \new_[84059]_ , \new_[84062]_ ,
    \new_[84065]_ , \new_[84066]_ , \new_[84067]_ , \new_[84070]_ ,
    \new_[84073]_ , \new_[84074]_ , \new_[84077]_ , \new_[84080]_ ,
    \new_[84081]_ , \new_[84082]_ , \new_[84085]_ , \new_[84088]_ ,
    \new_[84089]_ , \new_[84092]_ , \new_[84095]_ , \new_[84096]_ ,
    \new_[84097]_ , \new_[84100]_ , \new_[84103]_ , \new_[84104]_ ,
    \new_[84107]_ , \new_[84110]_ , \new_[84111]_ , \new_[84112]_ ,
    \new_[84115]_ , \new_[84118]_ , \new_[84119]_ , \new_[84122]_ ,
    \new_[84125]_ , \new_[84126]_ , \new_[84127]_ , \new_[84130]_ ,
    \new_[84133]_ , \new_[84134]_ , \new_[84137]_ , \new_[84140]_ ,
    \new_[84141]_ , \new_[84142]_ , \new_[84145]_ , \new_[84148]_ ,
    \new_[84149]_ , \new_[84152]_ , \new_[84155]_ , \new_[84156]_ ,
    \new_[84157]_ , \new_[84160]_ , \new_[84163]_ , \new_[84164]_ ,
    \new_[84167]_ , \new_[84170]_ , \new_[84171]_ , \new_[84172]_ ,
    \new_[84175]_ , \new_[84178]_ , \new_[84179]_ , \new_[84182]_ ,
    \new_[84185]_ , \new_[84186]_ , \new_[84187]_ , \new_[84190]_ ,
    \new_[84193]_ , \new_[84194]_ , \new_[84197]_ , \new_[84200]_ ,
    \new_[84201]_ , \new_[84202]_ , \new_[84205]_ , \new_[84208]_ ,
    \new_[84209]_ , \new_[84212]_ , \new_[84215]_ , \new_[84216]_ ,
    \new_[84217]_ , \new_[84220]_ , \new_[84223]_ , \new_[84224]_ ,
    \new_[84227]_ , \new_[84230]_ , \new_[84231]_ , \new_[84232]_ ,
    \new_[84235]_ , \new_[84238]_ , \new_[84239]_ , \new_[84242]_ ,
    \new_[84245]_ , \new_[84246]_ , \new_[84247]_ , \new_[84250]_ ,
    \new_[84253]_ , \new_[84254]_ , \new_[84257]_ , \new_[84260]_ ,
    \new_[84261]_ , \new_[84262]_ , \new_[84265]_ , \new_[84268]_ ,
    \new_[84269]_ , \new_[84272]_ , \new_[84275]_ , \new_[84276]_ ,
    \new_[84277]_ , \new_[84280]_ , \new_[84283]_ , \new_[84284]_ ,
    \new_[84287]_ , \new_[84290]_ , \new_[84291]_ , \new_[84292]_ ,
    \new_[84295]_ , \new_[84298]_ , \new_[84299]_ , \new_[84302]_ ,
    \new_[84305]_ , \new_[84306]_ , \new_[84307]_ , \new_[84310]_ ,
    \new_[84313]_ , \new_[84314]_ , \new_[84317]_ , \new_[84320]_ ,
    \new_[84321]_ , \new_[84322]_ , \new_[84325]_ , \new_[84328]_ ,
    \new_[84329]_ , \new_[84332]_ , \new_[84335]_ , \new_[84336]_ ,
    \new_[84337]_ , \new_[84340]_ , \new_[84343]_ , \new_[84344]_ ,
    \new_[84347]_ , \new_[84350]_ , \new_[84351]_ , \new_[84352]_ ,
    \new_[84355]_ , \new_[84358]_ , \new_[84359]_ , \new_[84362]_ ,
    \new_[84365]_ , \new_[84366]_ , \new_[84367]_ , \new_[84370]_ ,
    \new_[84373]_ , \new_[84374]_ , \new_[84377]_ , \new_[84380]_ ,
    \new_[84381]_ , \new_[84382]_ , \new_[84385]_ , \new_[84388]_ ,
    \new_[84389]_ , \new_[84392]_ , \new_[84395]_ , \new_[84396]_ ,
    \new_[84397]_ , \new_[84400]_ , \new_[84403]_ , \new_[84404]_ ,
    \new_[84407]_ , \new_[84410]_ , \new_[84411]_ , \new_[84412]_ ,
    \new_[84415]_ , \new_[84418]_ , \new_[84419]_ , \new_[84422]_ ,
    \new_[84425]_ , \new_[84426]_ , \new_[84427]_ , \new_[84430]_ ,
    \new_[84433]_ , \new_[84434]_ , \new_[84437]_ , \new_[84440]_ ,
    \new_[84441]_ , \new_[84442]_ , \new_[84445]_ , \new_[84448]_ ,
    \new_[84449]_ , \new_[84452]_ , \new_[84455]_ , \new_[84456]_ ,
    \new_[84457]_ , \new_[84460]_ , \new_[84463]_ , \new_[84464]_ ,
    \new_[84467]_ , \new_[84470]_ , \new_[84471]_ , \new_[84472]_ ,
    \new_[84475]_ , \new_[84478]_ , \new_[84479]_ , \new_[84482]_ ,
    \new_[84485]_ , \new_[84486]_ , \new_[84487]_ , \new_[84490]_ ,
    \new_[84493]_ , \new_[84494]_ , \new_[84497]_ , \new_[84500]_ ,
    \new_[84501]_ , \new_[84502]_ , \new_[84505]_ , \new_[84508]_ ,
    \new_[84509]_ , \new_[84512]_ , \new_[84515]_ , \new_[84516]_ ,
    \new_[84517]_ , \new_[84520]_ , \new_[84523]_ , \new_[84524]_ ,
    \new_[84527]_ , \new_[84530]_ , \new_[84531]_ , \new_[84532]_ ,
    \new_[84535]_ , \new_[84538]_ , \new_[84539]_ , \new_[84542]_ ,
    \new_[84545]_ , \new_[84546]_ , \new_[84547]_ , \new_[84550]_ ,
    \new_[84553]_ , \new_[84554]_ , \new_[84557]_ , \new_[84560]_ ,
    \new_[84561]_ , \new_[84562]_ , \new_[84565]_ , \new_[84568]_ ,
    \new_[84569]_ , \new_[84572]_ , \new_[84575]_ , \new_[84576]_ ,
    \new_[84577]_ , \new_[84580]_ , \new_[84583]_ , \new_[84584]_ ,
    \new_[84587]_ , \new_[84590]_ , \new_[84591]_ , \new_[84592]_ ,
    \new_[84595]_ , \new_[84598]_ , \new_[84599]_ , \new_[84602]_ ,
    \new_[84605]_ , \new_[84606]_ , \new_[84607]_ , \new_[84610]_ ,
    \new_[84613]_ , \new_[84614]_ , \new_[84617]_ , \new_[84620]_ ,
    \new_[84621]_ , \new_[84622]_ , \new_[84625]_ , \new_[84628]_ ,
    \new_[84629]_ , \new_[84632]_ , \new_[84635]_ , \new_[84636]_ ,
    \new_[84637]_ , \new_[84640]_ , \new_[84643]_ , \new_[84644]_ ,
    \new_[84647]_ , \new_[84650]_ , \new_[84651]_ , \new_[84652]_ ,
    \new_[84655]_ , \new_[84658]_ , \new_[84659]_ , \new_[84662]_ ,
    \new_[84665]_ , \new_[84666]_ , \new_[84667]_ , \new_[84670]_ ,
    \new_[84673]_ , \new_[84674]_ , \new_[84677]_ , \new_[84680]_ ,
    \new_[84681]_ , \new_[84682]_ , \new_[84685]_ , \new_[84688]_ ,
    \new_[84689]_ , \new_[84692]_ , \new_[84695]_ , \new_[84696]_ ,
    \new_[84697]_ , \new_[84700]_ , \new_[84703]_ , \new_[84704]_ ,
    \new_[84707]_ , \new_[84710]_ , \new_[84711]_ , \new_[84712]_ ,
    \new_[84715]_ , \new_[84718]_ , \new_[84719]_ , \new_[84722]_ ,
    \new_[84725]_ , \new_[84726]_ , \new_[84727]_ , \new_[84730]_ ,
    \new_[84733]_ , \new_[84734]_ , \new_[84737]_ , \new_[84740]_ ,
    \new_[84741]_ , \new_[84742]_ , \new_[84745]_ , \new_[84748]_ ,
    \new_[84749]_ , \new_[84752]_ , \new_[84755]_ , \new_[84756]_ ,
    \new_[84757]_ , \new_[84760]_ , \new_[84763]_ , \new_[84764]_ ,
    \new_[84767]_ , \new_[84770]_ , \new_[84771]_ , \new_[84772]_ ,
    \new_[84775]_ , \new_[84778]_ , \new_[84779]_ , \new_[84782]_ ,
    \new_[84785]_ , \new_[84786]_ , \new_[84787]_ , \new_[84790]_ ,
    \new_[84793]_ , \new_[84794]_ , \new_[84797]_ , \new_[84800]_ ,
    \new_[84801]_ , \new_[84802]_ , \new_[84805]_ , \new_[84808]_ ,
    \new_[84809]_ , \new_[84812]_ , \new_[84815]_ , \new_[84816]_ ,
    \new_[84817]_ , \new_[84820]_ , \new_[84823]_ , \new_[84824]_ ,
    \new_[84827]_ , \new_[84830]_ , \new_[84831]_ , \new_[84832]_ ,
    \new_[84835]_ , \new_[84838]_ , \new_[84839]_ , \new_[84842]_ ,
    \new_[84845]_ , \new_[84846]_ , \new_[84847]_ , \new_[84850]_ ,
    \new_[84853]_ , \new_[84854]_ , \new_[84857]_ , \new_[84860]_ ,
    \new_[84861]_ , \new_[84862]_ , \new_[84865]_ , \new_[84868]_ ,
    \new_[84869]_ , \new_[84872]_ , \new_[84875]_ , \new_[84876]_ ,
    \new_[84877]_ , \new_[84880]_ , \new_[84883]_ , \new_[84884]_ ,
    \new_[84887]_ , \new_[84890]_ , \new_[84891]_ , \new_[84892]_ ,
    \new_[84895]_ , \new_[84898]_ , \new_[84899]_ , \new_[84902]_ ,
    \new_[84905]_ , \new_[84906]_ , \new_[84907]_ , \new_[84910]_ ,
    \new_[84913]_ , \new_[84914]_ , \new_[84917]_ , \new_[84920]_ ,
    \new_[84921]_ , \new_[84922]_ , \new_[84925]_ , \new_[84928]_ ,
    \new_[84929]_ , \new_[84932]_ , \new_[84935]_ , \new_[84936]_ ,
    \new_[84937]_ , \new_[84940]_ , \new_[84943]_ , \new_[84944]_ ,
    \new_[84947]_ , \new_[84950]_ , \new_[84951]_ , \new_[84952]_ ,
    \new_[84955]_ , \new_[84958]_ , \new_[84959]_ , \new_[84962]_ ,
    \new_[84965]_ , \new_[84966]_ , \new_[84967]_ , \new_[84970]_ ,
    \new_[84973]_ , \new_[84974]_ , \new_[84977]_ , \new_[84981]_ ,
    \new_[84982]_ , \new_[84983]_ , \new_[84984]_ , \new_[84987]_ ,
    \new_[84990]_ , \new_[84991]_ , \new_[84994]_ , \new_[84997]_ ,
    \new_[84998]_ , \new_[84999]_ , \new_[85002]_ , \new_[85005]_ ,
    \new_[85006]_ , \new_[85009]_ , \new_[85013]_ , \new_[85014]_ ,
    \new_[85015]_ , \new_[85016]_ , \new_[85019]_ , \new_[85022]_ ,
    \new_[85023]_ , \new_[85026]_ , \new_[85029]_ , \new_[85030]_ ,
    \new_[85031]_ , \new_[85034]_ , \new_[85037]_ , \new_[85038]_ ,
    \new_[85041]_ , \new_[85045]_ , \new_[85046]_ , \new_[85047]_ ,
    \new_[85048]_ , \new_[85051]_ , \new_[85054]_ , \new_[85055]_ ,
    \new_[85058]_ , \new_[85061]_ , \new_[85062]_ , \new_[85063]_ ,
    \new_[85066]_ , \new_[85069]_ , \new_[85070]_ , \new_[85073]_ ,
    \new_[85077]_ , \new_[85078]_ , \new_[85079]_ , \new_[85080]_ ,
    \new_[85083]_ , \new_[85086]_ , \new_[85087]_ , \new_[85090]_ ,
    \new_[85093]_ , \new_[85094]_ , \new_[85095]_ , \new_[85098]_ ,
    \new_[85101]_ , \new_[85102]_ , \new_[85105]_ , \new_[85109]_ ,
    \new_[85110]_ , \new_[85111]_ , \new_[85112]_ , \new_[85115]_ ,
    \new_[85118]_ , \new_[85119]_ , \new_[85122]_ , \new_[85125]_ ,
    \new_[85126]_ , \new_[85127]_ , \new_[85130]_ , \new_[85133]_ ,
    \new_[85134]_ , \new_[85137]_ , \new_[85141]_ , \new_[85142]_ ,
    \new_[85143]_ , \new_[85144]_ , \new_[85147]_ , \new_[85150]_ ,
    \new_[85151]_ , \new_[85154]_ , \new_[85157]_ , \new_[85158]_ ,
    \new_[85159]_ , \new_[85162]_ , \new_[85165]_ , \new_[85166]_ ,
    \new_[85169]_ , \new_[85173]_ , \new_[85174]_ , \new_[85175]_ ,
    \new_[85176]_ , \new_[85179]_ , \new_[85182]_ , \new_[85183]_ ,
    \new_[85186]_ , \new_[85189]_ , \new_[85190]_ , \new_[85191]_ ,
    \new_[85194]_ , \new_[85197]_ , \new_[85198]_ , \new_[85201]_ ,
    \new_[85205]_ , \new_[85206]_ , \new_[85207]_ , \new_[85208]_ ,
    \new_[85211]_ , \new_[85214]_ , \new_[85215]_ , \new_[85218]_ ,
    \new_[85221]_ , \new_[85222]_ , \new_[85223]_ , \new_[85226]_ ,
    \new_[85229]_ , \new_[85230]_ , \new_[85233]_ , \new_[85237]_ ,
    \new_[85238]_ , \new_[85239]_ , \new_[85240]_ , \new_[85243]_ ,
    \new_[85246]_ , \new_[85247]_ , \new_[85250]_ , \new_[85253]_ ,
    \new_[85254]_ , \new_[85255]_ , \new_[85258]_ , \new_[85261]_ ,
    \new_[85262]_ , \new_[85265]_ , \new_[85269]_ , \new_[85270]_ ,
    \new_[85271]_ , \new_[85272]_ , \new_[85275]_ , \new_[85278]_ ,
    \new_[85279]_ , \new_[85282]_ , \new_[85285]_ , \new_[85286]_ ,
    \new_[85287]_ , \new_[85290]_ , \new_[85293]_ , \new_[85294]_ ,
    \new_[85297]_ , \new_[85301]_ , \new_[85302]_ , \new_[85303]_ ,
    \new_[85304]_ , \new_[85307]_ , \new_[85310]_ , \new_[85311]_ ,
    \new_[85314]_ , \new_[85317]_ , \new_[85318]_ , \new_[85319]_ ,
    \new_[85322]_ , \new_[85325]_ , \new_[85326]_ , \new_[85329]_ ,
    \new_[85333]_ , \new_[85334]_ , \new_[85335]_ , \new_[85336]_ ,
    \new_[85339]_ , \new_[85342]_ , \new_[85343]_ , \new_[85346]_ ,
    \new_[85349]_ , \new_[85350]_ , \new_[85351]_ , \new_[85354]_ ,
    \new_[85357]_ , \new_[85358]_ , \new_[85361]_ , \new_[85365]_ ,
    \new_[85366]_ , \new_[85367]_ , \new_[85368]_ , \new_[85371]_ ,
    \new_[85374]_ , \new_[85375]_ , \new_[85378]_ , \new_[85381]_ ,
    \new_[85382]_ , \new_[85383]_ , \new_[85386]_ , \new_[85389]_ ,
    \new_[85390]_ , \new_[85393]_ , \new_[85397]_ , \new_[85398]_ ,
    \new_[85399]_ , \new_[85400]_ , \new_[85403]_ , \new_[85406]_ ,
    \new_[85407]_ , \new_[85410]_ , \new_[85413]_ , \new_[85414]_ ,
    \new_[85415]_ , \new_[85418]_ , \new_[85421]_ , \new_[85422]_ ,
    \new_[85425]_ , \new_[85429]_ , \new_[85430]_ , \new_[85431]_ ,
    \new_[85432]_ , \new_[85435]_ , \new_[85438]_ , \new_[85439]_ ,
    \new_[85442]_ , \new_[85445]_ , \new_[85446]_ , \new_[85447]_ ,
    \new_[85450]_ , \new_[85453]_ , \new_[85454]_ , \new_[85457]_ ,
    \new_[85461]_ , \new_[85462]_ , \new_[85463]_ , \new_[85464]_ ,
    \new_[85467]_ , \new_[85470]_ , \new_[85471]_ , \new_[85474]_ ,
    \new_[85477]_ , \new_[85478]_ , \new_[85479]_ , \new_[85482]_ ,
    \new_[85485]_ , \new_[85486]_ , \new_[85489]_ , \new_[85493]_ ,
    \new_[85494]_ , \new_[85495]_ , \new_[85496]_ , \new_[85499]_ ,
    \new_[85502]_ , \new_[85503]_ , \new_[85506]_ , \new_[85509]_ ,
    \new_[85510]_ , \new_[85511]_ , \new_[85514]_ , \new_[85517]_ ,
    \new_[85518]_ , \new_[85521]_ , \new_[85525]_ , \new_[85526]_ ,
    \new_[85527]_ , \new_[85528]_ , \new_[85531]_ , \new_[85534]_ ,
    \new_[85535]_ , \new_[85538]_ , \new_[85541]_ , \new_[85542]_ ,
    \new_[85543]_ , \new_[85546]_ , \new_[85549]_ , \new_[85550]_ ,
    \new_[85553]_ , \new_[85557]_ , \new_[85558]_ , \new_[85559]_ ,
    \new_[85560]_ , \new_[85563]_ , \new_[85566]_ , \new_[85567]_ ,
    \new_[85570]_ , \new_[85573]_ , \new_[85574]_ , \new_[85575]_ ,
    \new_[85578]_ , \new_[85581]_ , \new_[85582]_ , \new_[85585]_ ,
    \new_[85589]_ , \new_[85590]_ , \new_[85591]_ , \new_[85592]_ ,
    \new_[85595]_ , \new_[85598]_ , \new_[85599]_ , \new_[85602]_ ,
    \new_[85605]_ , \new_[85606]_ , \new_[85607]_ , \new_[85610]_ ,
    \new_[85613]_ , \new_[85614]_ , \new_[85617]_ , \new_[85621]_ ,
    \new_[85622]_ , \new_[85623]_ , \new_[85624]_ , \new_[85627]_ ,
    \new_[85630]_ , \new_[85631]_ , \new_[85634]_ , \new_[85637]_ ,
    \new_[85638]_ , \new_[85639]_ , \new_[85642]_ , \new_[85645]_ ,
    \new_[85646]_ , \new_[85649]_ , \new_[85653]_ , \new_[85654]_ ,
    \new_[85655]_ , \new_[85656]_ , \new_[85659]_ , \new_[85662]_ ,
    \new_[85663]_ , \new_[85666]_ , \new_[85669]_ , \new_[85670]_ ,
    \new_[85671]_ , \new_[85674]_ , \new_[85677]_ , \new_[85678]_ ,
    \new_[85681]_ , \new_[85685]_ , \new_[85686]_ , \new_[85687]_ ,
    \new_[85688]_ , \new_[85691]_ , \new_[85694]_ , \new_[85695]_ ,
    \new_[85698]_ , \new_[85701]_ , \new_[85702]_ , \new_[85703]_ ,
    \new_[85706]_ , \new_[85709]_ , \new_[85710]_ , \new_[85713]_ ,
    \new_[85717]_ , \new_[85718]_ , \new_[85719]_ , \new_[85720]_ ,
    \new_[85723]_ , \new_[85726]_ , \new_[85727]_ , \new_[85730]_ ,
    \new_[85733]_ , \new_[85734]_ , \new_[85735]_ , \new_[85738]_ ,
    \new_[85741]_ , \new_[85742]_ , \new_[85745]_ , \new_[85749]_ ,
    \new_[85750]_ , \new_[85751]_ , \new_[85752]_ , \new_[85755]_ ,
    \new_[85758]_ , \new_[85759]_ , \new_[85762]_ , \new_[85765]_ ,
    \new_[85766]_ , \new_[85767]_ , \new_[85770]_ , \new_[85773]_ ,
    \new_[85774]_ , \new_[85777]_ , \new_[85781]_ , \new_[85782]_ ,
    \new_[85783]_ , \new_[85784]_ , \new_[85787]_ , \new_[85790]_ ,
    \new_[85791]_ , \new_[85794]_ , \new_[85797]_ , \new_[85798]_ ,
    \new_[85799]_ , \new_[85802]_ , \new_[85805]_ , \new_[85806]_ ,
    \new_[85809]_ , \new_[85813]_ , \new_[85814]_ , \new_[85815]_ ,
    \new_[85816]_ , \new_[85819]_ , \new_[85822]_ , \new_[85823]_ ,
    \new_[85826]_ , \new_[85829]_ , \new_[85830]_ , \new_[85831]_ ,
    \new_[85834]_ , \new_[85837]_ , \new_[85838]_ , \new_[85841]_ ,
    \new_[85845]_ , \new_[85846]_ , \new_[85847]_ , \new_[85848]_ ,
    \new_[85851]_ , \new_[85854]_ , \new_[85855]_ , \new_[85858]_ ,
    \new_[85861]_ , \new_[85862]_ , \new_[85863]_ , \new_[85866]_ ,
    \new_[85869]_ , \new_[85870]_ , \new_[85873]_ , \new_[85877]_ ,
    \new_[85878]_ , \new_[85879]_ , \new_[85880]_ , \new_[85883]_ ,
    \new_[85886]_ , \new_[85887]_ , \new_[85890]_ , \new_[85893]_ ,
    \new_[85894]_ , \new_[85895]_ , \new_[85898]_ , \new_[85901]_ ,
    \new_[85902]_ , \new_[85905]_ , \new_[85909]_ , \new_[85910]_ ,
    \new_[85911]_ , \new_[85912]_ , \new_[85915]_ , \new_[85918]_ ,
    \new_[85919]_ , \new_[85922]_ , \new_[85925]_ , \new_[85926]_ ,
    \new_[85927]_ , \new_[85930]_ , \new_[85933]_ , \new_[85934]_ ,
    \new_[85937]_ , \new_[85941]_ , \new_[85942]_ , \new_[85943]_ ,
    \new_[85944]_ , \new_[85947]_ , \new_[85950]_ , \new_[85951]_ ,
    \new_[85954]_ , \new_[85957]_ , \new_[85958]_ , \new_[85959]_ ,
    \new_[85962]_ , \new_[85965]_ , \new_[85966]_ , \new_[85969]_ ,
    \new_[85973]_ , \new_[85974]_ , \new_[85975]_ , \new_[85976]_ ,
    \new_[85979]_ , \new_[85982]_ , \new_[85983]_ , \new_[85986]_ ,
    \new_[85989]_ , \new_[85990]_ , \new_[85991]_ , \new_[85994]_ ,
    \new_[85997]_ , \new_[85998]_ , \new_[86001]_ , \new_[86005]_ ,
    \new_[86006]_ , \new_[86007]_ , \new_[86008]_ , \new_[86011]_ ,
    \new_[86014]_ , \new_[86015]_ , \new_[86018]_ , \new_[86021]_ ,
    \new_[86022]_ , \new_[86023]_ , \new_[86026]_ , \new_[86029]_ ,
    \new_[86030]_ , \new_[86033]_ , \new_[86037]_ , \new_[86038]_ ,
    \new_[86039]_ , \new_[86040]_ , \new_[86043]_ , \new_[86046]_ ,
    \new_[86047]_ , \new_[86050]_ , \new_[86053]_ , \new_[86054]_ ,
    \new_[86055]_ , \new_[86058]_ , \new_[86061]_ , \new_[86062]_ ,
    \new_[86065]_ , \new_[86069]_ , \new_[86070]_ , \new_[86071]_ ,
    \new_[86072]_ , \new_[86075]_ , \new_[86078]_ , \new_[86079]_ ,
    \new_[86082]_ , \new_[86085]_ , \new_[86086]_ , \new_[86087]_ ,
    \new_[86090]_ , \new_[86093]_ , \new_[86094]_ , \new_[86097]_ ,
    \new_[86101]_ , \new_[86102]_ , \new_[86103]_ , \new_[86104]_ ,
    \new_[86107]_ , \new_[86110]_ , \new_[86111]_ , \new_[86114]_ ,
    \new_[86117]_ , \new_[86118]_ , \new_[86119]_ , \new_[86122]_ ,
    \new_[86125]_ , \new_[86126]_ , \new_[86129]_ , \new_[86133]_ ,
    \new_[86134]_ , \new_[86135]_ , \new_[86136]_ , \new_[86139]_ ,
    \new_[86142]_ , \new_[86143]_ , \new_[86146]_ , \new_[86149]_ ,
    \new_[86150]_ , \new_[86151]_ , \new_[86154]_ , \new_[86157]_ ,
    \new_[86158]_ , \new_[86161]_ , \new_[86165]_ , \new_[86166]_ ,
    \new_[86167]_ , \new_[86168]_ , \new_[86171]_ , \new_[86174]_ ,
    \new_[86175]_ , \new_[86178]_ , \new_[86181]_ , \new_[86182]_ ,
    \new_[86183]_ , \new_[86186]_ , \new_[86189]_ , \new_[86190]_ ,
    \new_[86193]_ , \new_[86197]_ , \new_[86198]_ , \new_[86199]_ ,
    \new_[86200]_ , \new_[86203]_ , \new_[86206]_ , \new_[86207]_ ,
    \new_[86210]_ , \new_[86213]_ , \new_[86214]_ , \new_[86215]_ ,
    \new_[86218]_ , \new_[86221]_ , \new_[86222]_ , \new_[86225]_ ,
    \new_[86229]_ , \new_[86230]_ , \new_[86231]_ , \new_[86232]_ ,
    \new_[86235]_ , \new_[86238]_ , \new_[86239]_ , \new_[86242]_ ,
    \new_[86245]_ , \new_[86246]_ , \new_[86247]_ , \new_[86250]_ ,
    \new_[86253]_ , \new_[86254]_ , \new_[86257]_ , \new_[86261]_ ,
    \new_[86262]_ , \new_[86263]_ , \new_[86264]_ , \new_[86267]_ ,
    \new_[86270]_ , \new_[86271]_ , \new_[86274]_ , \new_[86277]_ ,
    \new_[86278]_ , \new_[86279]_ , \new_[86282]_ , \new_[86285]_ ,
    \new_[86286]_ , \new_[86289]_ , \new_[86293]_ , \new_[86294]_ ,
    \new_[86295]_ , \new_[86296]_ , \new_[86299]_ , \new_[86302]_ ,
    \new_[86303]_ , \new_[86306]_ , \new_[86309]_ , \new_[86310]_ ,
    \new_[86311]_ , \new_[86314]_ , \new_[86317]_ , \new_[86318]_ ,
    \new_[86321]_ , \new_[86325]_ , \new_[86326]_ , \new_[86327]_ ,
    \new_[86328]_ , \new_[86331]_ , \new_[86334]_ , \new_[86335]_ ,
    \new_[86338]_ , \new_[86341]_ , \new_[86342]_ , \new_[86343]_ ,
    \new_[86346]_ , \new_[86349]_ , \new_[86350]_ , \new_[86353]_ ,
    \new_[86357]_ , \new_[86358]_ , \new_[86359]_ , \new_[86360]_ ,
    \new_[86363]_ , \new_[86366]_ , \new_[86367]_ , \new_[86370]_ ,
    \new_[86373]_ , \new_[86374]_ , \new_[86375]_ , \new_[86378]_ ,
    \new_[86381]_ , \new_[86382]_ , \new_[86385]_ , \new_[86389]_ ,
    \new_[86390]_ , \new_[86391]_ , \new_[86392]_ , \new_[86395]_ ,
    \new_[86398]_ , \new_[86399]_ , \new_[86402]_ , \new_[86405]_ ,
    \new_[86406]_ , \new_[86407]_ , \new_[86410]_ , \new_[86413]_ ,
    \new_[86414]_ , \new_[86417]_ , \new_[86421]_ , \new_[86422]_ ,
    \new_[86423]_ , \new_[86424]_ , \new_[86427]_ , \new_[86430]_ ,
    \new_[86431]_ , \new_[86434]_ , \new_[86437]_ , \new_[86438]_ ,
    \new_[86439]_ , \new_[86442]_ , \new_[86445]_ , \new_[86446]_ ,
    \new_[86449]_ , \new_[86453]_ , \new_[86454]_ , \new_[86455]_ ,
    \new_[86456]_ , \new_[86459]_ , \new_[86462]_ , \new_[86463]_ ,
    \new_[86466]_ , \new_[86469]_ , \new_[86470]_ , \new_[86471]_ ,
    \new_[86474]_ , \new_[86477]_ , \new_[86478]_ , \new_[86481]_ ,
    \new_[86485]_ , \new_[86486]_ , \new_[86487]_ , \new_[86488]_ ,
    \new_[86491]_ , \new_[86494]_ , \new_[86495]_ , \new_[86498]_ ,
    \new_[86501]_ , \new_[86502]_ , \new_[86503]_ , \new_[86506]_ ,
    \new_[86509]_ , \new_[86510]_ , \new_[86513]_ , \new_[86517]_ ,
    \new_[86518]_ , \new_[86519]_ , \new_[86520]_ , \new_[86523]_ ,
    \new_[86526]_ , \new_[86527]_ , \new_[86530]_ , \new_[86533]_ ,
    \new_[86534]_ , \new_[86535]_ , \new_[86538]_ , \new_[86541]_ ,
    \new_[86542]_ , \new_[86545]_ , \new_[86549]_ , \new_[86550]_ ,
    \new_[86551]_ , \new_[86552]_ , \new_[86555]_ , \new_[86558]_ ,
    \new_[86559]_ , \new_[86562]_ , \new_[86565]_ , \new_[86566]_ ,
    \new_[86567]_ , \new_[86570]_ , \new_[86573]_ , \new_[86574]_ ,
    \new_[86577]_ , \new_[86581]_ , \new_[86582]_ , \new_[86583]_ ,
    \new_[86584]_ , \new_[86587]_ , \new_[86590]_ , \new_[86591]_ ,
    \new_[86594]_ , \new_[86597]_ , \new_[86598]_ , \new_[86599]_ ,
    \new_[86602]_ , \new_[86605]_ , \new_[86606]_ , \new_[86609]_ ,
    \new_[86613]_ , \new_[86614]_ , \new_[86615]_ , \new_[86616]_ ,
    \new_[86619]_ , \new_[86622]_ , \new_[86623]_ , \new_[86626]_ ,
    \new_[86629]_ , \new_[86630]_ , \new_[86631]_ , \new_[86634]_ ,
    \new_[86637]_ , \new_[86638]_ , \new_[86641]_ , \new_[86645]_ ,
    \new_[86646]_ , \new_[86647]_ , \new_[86648]_ , \new_[86651]_ ,
    \new_[86654]_ , \new_[86655]_ , \new_[86658]_ , \new_[86661]_ ,
    \new_[86662]_ , \new_[86663]_ , \new_[86666]_ , \new_[86669]_ ,
    \new_[86670]_ , \new_[86673]_ , \new_[86677]_ , \new_[86678]_ ,
    \new_[86679]_ , \new_[86680]_ , \new_[86683]_ , \new_[86686]_ ,
    \new_[86687]_ , \new_[86690]_ , \new_[86693]_ , \new_[86694]_ ,
    \new_[86695]_ , \new_[86698]_ , \new_[86701]_ , \new_[86702]_ ,
    \new_[86705]_ , \new_[86709]_ , \new_[86710]_ , \new_[86711]_ ,
    \new_[86712]_ , \new_[86715]_ , \new_[86718]_ , \new_[86719]_ ,
    \new_[86722]_ , \new_[86725]_ , \new_[86726]_ , \new_[86727]_ ,
    \new_[86730]_ , \new_[86733]_ , \new_[86734]_ , \new_[86737]_ ,
    \new_[86741]_ , \new_[86742]_ , \new_[86743]_ , \new_[86744]_ ,
    \new_[86747]_ , \new_[86750]_ , \new_[86751]_ , \new_[86754]_ ,
    \new_[86757]_ , \new_[86758]_ , \new_[86759]_ , \new_[86762]_ ,
    \new_[86765]_ , \new_[86766]_ , \new_[86769]_ , \new_[86773]_ ,
    \new_[86774]_ , \new_[86775]_ , \new_[86776]_ , \new_[86779]_ ,
    \new_[86782]_ , \new_[86783]_ , \new_[86786]_ , \new_[86789]_ ,
    \new_[86790]_ , \new_[86791]_ , \new_[86794]_ , \new_[86797]_ ,
    \new_[86798]_ , \new_[86801]_ , \new_[86805]_ , \new_[86806]_ ,
    \new_[86807]_ , \new_[86808]_ , \new_[86811]_ , \new_[86814]_ ,
    \new_[86815]_ , \new_[86818]_ , \new_[86821]_ , \new_[86822]_ ,
    \new_[86823]_ , \new_[86826]_ , \new_[86829]_ , \new_[86830]_ ,
    \new_[86833]_ , \new_[86837]_ , \new_[86838]_ , \new_[86839]_ ,
    \new_[86840]_ , \new_[86843]_ , \new_[86846]_ , \new_[86847]_ ,
    \new_[86850]_ , \new_[86853]_ , \new_[86854]_ , \new_[86855]_ ,
    \new_[86858]_ , \new_[86861]_ , \new_[86862]_ , \new_[86865]_ ,
    \new_[86869]_ , \new_[86870]_ , \new_[86871]_ , \new_[86872]_ ,
    \new_[86875]_ , \new_[86878]_ , \new_[86879]_ , \new_[86882]_ ,
    \new_[86885]_ , \new_[86886]_ , \new_[86887]_ , \new_[86890]_ ,
    \new_[86893]_ , \new_[86894]_ , \new_[86897]_ , \new_[86901]_ ,
    \new_[86902]_ , \new_[86903]_ , \new_[86904]_ , \new_[86907]_ ,
    \new_[86910]_ , \new_[86911]_ , \new_[86914]_ , \new_[86917]_ ,
    \new_[86918]_ , \new_[86919]_ , \new_[86922]_ , \new_[86925]_ ,
    \new_[86926]_ , \new_[86929]_ , \new_[86933]_ , \new_[86934]_ ,
    \new_[86935]_ , \new_[86936]_ , \new_[86939]_ , \new_[86942]_ ,
    \new_[86943]_ , \new_[86946]_ , \new_[86949]_ , \new_[86950]_ ,
    \new_[86951]_ , \new_[86954]_ , \new_[86957]_ , \new_[86958]_ ,
    \new_[86961]_ , \new_[86965]_ , \new_[86966]_ , \new_[86967]_ ,
    \new_[86968]_ , \new_[86971]_ , \new_[86974]_ , \new_[86975]_ ,
    \new_[86978]_ , \new_[86981]_ , \new_[86982]_ , \new_[86983]_ ,
    \new_[86986]_ , \new_[86989]_ , \new_[86990]_ , \new_[86993]_ ,
    \new_[86997]_ , \new_[86998]_ , \new_[86999]_ , \new_[87000]_ ,
    \new_[87003]_ , \new_[87006]_ , \new_[87007]_ , \new_[87010]_ ,
    \new_[87013]_ , \new_[87014]_ , \new_[87015]_ , \new_[87018]_ ,
    \new_[87021]_ , \new_[87022]_ , \new_[87025]_ , \new_[87029]_ ,
    \new_[87030]_ , \new_[87031]_ , \new_[87032]_ , \new_[87035]_ ,
    \new_[87038]_ , \new_[87039]_ , \new_[87042]_ , \new_[87045]_ ,
    \new_[87046]_ , \new_[87047]_ , \new_[87050]_ , \new_[87053]_ ,
    \new_[87054]_ , \new_[87057]_ , \new_[87061]_ , \new_[87062]_ ,
    \new_[87063]_ , \new_[87064]_ , \new_[87067]_ , \new_[87070]_ ,
    \new_[87071]_ , \new_[87074]_ , \new_[87077]_ , \new_[87078]_ ,
    \new_[87079]_ , \new_[87082]_ , \new_[87085]_ , \new_[87086]_ ,
    \new_[87089]_ , \new_[87093]_ , \new_[87094]_ , \new_[87095]_ ,
    \new_[87096]_ , \new_[87099]_ , \new_[87102]_ , \new_[87103]_ ,
    \new_[87106]_ , \new_[87109]_ , \new_[87110]_ , \new_[87111]_ ,
    \new_[87114]_ , \new_[87117]_ , \new_[87118]_ , \new_[87121]_ ,
    \new_[87125]_ , \new_[87126]_ , \new_[87127]_ , \new_[87128]_ ,
    \new_[87131]_ , \new_[87134]_ , \new_[87135]_ , \new_[87138]_ ,
    \new_[87141]_ , \new_[87142]_ , \new_[87143]_ , \new_[87146]_ ,
    \new_[87149]_ , \new_[87150]_ , \new_[87153]_ , \new_[87157]_ ,
    \new_[87158]_ , \new_[87159]_ , \new_[87160]_ , \new_[87163]_ ,
    \new_[87166]_ , \new_[87167]_ , \new_[87170]_ , \new_[87173]_ ,
    \new_[87174]_ , \new_[87175]_ , \new_[87178]_ , \new_[87181]_ ,
    \new_[87182]_ , \new_[87185]_ , \new_[87189]_ , \new_[87190]_ ,
    \new_[87191]_ , \new_[87192]_ , \new_[87195]_ , \new_[87198]_ ,
    \new_[87199]_ , \new_[87202]_ , \new_[87205]_ , \new_[87206]_ ,
    \new_[87207]_ , \new_[87210]_ , \new_[87213]_ , \new_[87214]_ ,
    \new_[87217]_ , \new_[87221]_ , \new_[87222]_ , \new_[87223]_ ,
    \new_[87224]_ , \new_[87227]_ , \new_[87230]_ , \new_[87231]_ ,
    \new_[87234]_ , \new_[87237]_ , \new_[87238]_ , \new_[87239]_ ,
    \new_[87242]_ , \new_[87245]_ , \new_[87246]_ , \new_[87249]_ ,
    \new_[87253]_ , \new_[87254]_ , \new_[87255]_ , \new_[87256]_ ,
    \new_[87259]_ , \new_[87262]_ , \new_[87263]_ , \new_[87266]_ ,
    \new_[87269]_ , \new_[87270]_ , \new_[87271]_ , \new_[87274]_ ,
    \new_[87277]_ , \new_[87278]_ , \new_[87281]_ , \new_[87285]_ ,
    \new_[87286]_ , \new_[87287]_ , \new_[87288]_ , \new_[87291]_ ,
    \new_[87294]_ , \new_[87295]_ , \new_[87298]_ , \new_[87301]_ ,
    \new_[87302]_ , \new_[87303]_ , \new_[87306]_ , \new_[87309]_ ,
    \new_[87310]_ , \new_[87313]_ , \new_[87317]_ , \new_[87318]_ ,
    \new_[87319]_ , \new_[87320]_ , \new_[87323]_ , \new_[87326]_ ,
    \new_[87327]_ , \new_[87330]_ , \new_[87333]_ , \new_[87334]_ ,
    \new_[87335]_ , \new_[87338]_ , \new_[87341]_ , \new_[87342]_ ,
    \new_[87345]_ , \new_[87349]_ , \new_[87350]_ , \new_[87351]_ ,
    \new_[87352]_ , \new_[87355]_ , \new_[87358]_ , \new_[87359]_ ,
    \new_[87362]_ , \new_[87365]_ , \new_[87366]_ , \new_[87367]_ ,
    \new_[87370]_ , \new_[87373]_ , \new_[87374]_ , \new_[87377]_ ,
    \new_[87381]_ , \new_[87382]_ , \new_[87383]_ , \new_[87384]_ ,
    \new_[87387]_ , \new_[87390]_ , \new_[87391]_ , \new_[87394]_ ,
    \new_[87397]_ , \new_[87398]_ , \new_[87399]_ , \new_[87402]_ ,
    \new_[87405]_ , \new_[87406]_ , \new_[87409]_ , \new_[87413]_ ,
    \new_[87414]_ , \new_[87415]_ , \new_[87416]_ , \new_[87419]_ ,
    \new_[87422]_ , \new_[87423]_ , \new_[87426]_ , \new_[87429]_ ,
    \new_[87430]_ , \new_[87431]_ , \new_[87434]_ , \new_[87437]_ ,
    \new_[87438]_ , \new_[87441]_ , \new_[87445]_ , \new_[87446]_ ,
    \new_[87447]_ , \new_[87448]_ , \new_[87451]_ , \new_[87454]_ ,
    \new_[87455]_ , \new_[87458]_ , \new_[87461]_ , \new_[87462]_ ,
    \new_[87463]_ , \new_[87466]_ , \new_[87469]_ , \new_[87470]_ ,
    \new_[87473]_ , \new_[87477]_ , \new_[87478]_ , \new_[87479]_ ,
    \new_[87480]_ , \new_[87483]_ , \new_[87486]_ , \new_[87487]_ ,
    \new_[87490]_ , \new_[87493]_ , \new_[87494]_ , \new_[87495]_ ,
    \new_[87498]_ , \new_[87501]_ , \new_[87502]_ , \new_[87505]_ ,
    \new_[87509]_ , \new_[87510]_ , \new_[87511]_ , \new_[87512]_ ,
    \new_[87515]_ , \new_[87518]_ , \new_[87519]_ , \new_[87522]_ ,
    \new_[87525]_ , \new_[87526]_ , \new_[87527]_ , \new_[87530]_ ,
    \new_[87533]_ , \new_[87534]_ , \new_[87537]_ , \new_[87541]_ ,
    \new_[87542]_ , \new_[87543]_ , \new_[87544]_ , \new_[87547]_ ,
    \new_[87550]_ , \new_[87551]_ , \new_[87554]_ , \new_[87557]_ ,
    \new_[87558]_ , \new_[87559]_ , \new_[87562]_ , \new_[87565]_ ,
    \new_[87566]_ , \new_[87569]_ , \new_[87573]_ , \new_[87574]_ ,
    \new_[87575]_ , \new_[87576]_ , \new_[87579]_ , \new_[87582]_ ,
    \new_[87583]_ , \new_[87586]_ , \new_[87589]_ , \new_[87590]_ ,
    \new_[87591]_ , \new_[87594]_ , \new_[87597]_ , \new_[87598]_ ,
    \new_[87601]_ , \new_[87605]_ , \new_[87606]_ , \new_[87607]_ ,
    \new_[87608]_ , \new_[87611]_ , \new_[87614]_ , \new_[87615]_ ,
    \new_[87618]_ , \new_[87621]_ , \new_[87622]_ , \new_[87623]_ ,
    \new_[87626]_ , \new_[87629]_ , \new_[87630]_ , \new_[87633]_ ,
    \new_[87637]_ , \new_[87638]_ , \new_[87639]_ , \new_[87640]_ ,
    \new_[87643]_ , \new_[87646]_ , \new_[87647]_ , \new_[87650]_ ,
    \new_[87653]_ , \new_[87654]_ , \new_[87655]_ , \new_[87658]_ ,
    \new_[87661]_ , \new_[87662]_ , \new_[87665]_ , \new_[87669]_ ,
    \new_[87670]_ , \new_[87671]_ , \new_[87672]_ , \new_[87675]_ ,
    \new_[87678]_ , \new_[87679]_ , \new_[87682]_ , \new_[87685]_ ,
    \new_[87686]_ , \new_[87687]_ , \new_[87690]_ , \new_[87693]_ ,
    \new_[87694]_ , \new_[87697]_ , \new_[87701]_ , \new_[87702]_ ,
    \new_[87703]_ , \new_[87704]_ , \new_[87707]_ , \new_[87710]_ ,
    \new_[87711]_ , \new_[87714]_ , \new_[87717]_ , \new_[87718]_ ,
    \new_[87719]_ , \new_[87722]_ , \new_[87725]_ , \new_[87726]_ ,
    \new_[87729]_ , \new_[87733]_ , \new_[87734]_ , \new_[87735]_ ,
    \new_[87736]_ , \new_[87739]_ , \new_[87742]_ , \new_[87743]_ ,
    \new_[87746]_ , \new_[87749]_ , \new_[87750]_ , \new_[87751]_ ,
    \new_[87754]_ , \new_[87757]_ , \new_[87758]_ , \new_[87761]_ ,
    \new_[87765]_ , \new_[87766]_ , \new_[87767]_ , \new_[87768]_ ,
    \new_[87771]_ , \new_[87774]_ , \new_[87775]_ , \new_[87778]_ ,
    \new_[87781]_ , \new_[87782]_ , \new_[87783]_ , \new_[87786]_ ,
    \new_[87789]_ , \new_[87790]_ , \new_[87793]_ , \new_[87797]_ ,
    \new_[87798]_ , \new_[87799]_ , \new_[87800]_ , \new_[87803]_ ,
    \new_[87806]_ , \new_[87807]_ , \new_[87810]_ , \new_[87813]_ ,
    \new_[87814]_ , \new_[87815]_ , \new_[87818]_ , \new_[87821]_ ,
    \new_[87822]_ , \new_[87825]_ , \new_[87829]_ , \new_[87830]_ ,
    \new_[87831]_ , \new_[87832]_ , \new_[87835]_ , \new_[87838]_ ,
    \new_[87839]_ , \new_[87842]_ , \new_[87845]_ , \new_[87846]_ ,
    \new_[87847]_ , \new_[87850]_ , \new_[87853]_ , \new_[87854]_ ,
    \new_[87857]_ , \new_[87861]_ , \new_[87862]_ , \new_[87863]_ ,
    \new_[87864]_ , \new_[87867]_ , \new_[87870]_ , \new_[87871]_ ,
    \new_[87874]_ , \new_[87877]_ , \new_[87878]_ , \new_[87879]_ ,
    \new_[87882]_ , \new_[87885]_ , \new_[87886]_ , \new_[87889]_ ,
    \new_[87893]_ , \new_[87894]_ , \new_[87895]_ , \new_[87896]_ ,
    \new_[87899]_ , \new_[87902]_ , \new_[87903]_ , \new_[87906]_ ,
    \new_[87909]_ , \new_[87910]_ , \new_[87911]_ , \new_[87914]_ ,
    \new_[87917]_ , \new_[87918]_ , \new_[87921]_ , \new_[87925]_ ,
    \new_[87926]_ , \new_[87927]_ , \new_[87928]_ , \new_[87931]_ ,
    \new_[87934]_ , \new_[87935]_ , \new_[87938]_ , \new_[87941]_ ,
    \new_[87942]_ , \new_[87943]_ , \new_[87946]_ , \new_[87949]_ ,
    \new_[87950]_ , \new_[87953]_ , \new_[87957]_ , \new_[87958]_ ,
    \new_[87959]_ , \new_[87960]_ , \new_[87963]_ , \new_[87966]_ ,
    \new_[87967]_ , \new_[87970]_ , \new_[87973]_ , \new_[87974]_ ,
    \new_[87975]_ , \new_[87978]_ , \new_[87981]_ , \new_[87982]_ ,
    \new_[87985]_ , \new_[87989]_ , \new_[87990]_ , \new_[87991]_ ,
    \new_[87992]_ , \new_[87995]_ , \new_[87998]_ , \new_[87999]_ ,
    \new_[88002]_ , \new_[88005]_ , \new_[88006]_ , \new_[88007]_ ,
    \new_[88010]_ , \new_[88013]_ , \new_[88014]_ , \new_[88017]_ ,
    \new_[88021]_ , \new_[88022]_ , \new_[88023]_ , \new_[88024]_ ,
    \new_[88027]_ , \new_[88030]_ , \new_[88031]_ , \new_[88034]_ ,
    \new_[88037]_ , \new_[88038]_ , \new_[88039]_ , \new_[88042]_ ,
    \new_[88045]_ , \new_[88046]_ , \new_[88049]_ , \new_[88053]_ ,
    \new_[88054]_ , \new_[88055]_ , \new_[88056]_ , \new_[88059]_ ,
    \new_[88062]_ , \new_[88063]_ , \new_[88066]_ , \new_[88069]_ ,
    \new_[88070]_ , \new_[88071]_ , \new_[88074]_ , \new_[88077]_ ,
    \new_[88078]_ , \new_[88081]_ , \new_[88085]_ , \new_[88086]_ ,
    \new_[88087]_ , \new_[88088]_ , \new_[88091]_ , \new_[88094]_ ,
    \new_[88095]_ , \new_[88098]_ , \new_[88101]_ , \new_[88102]_ ,
    \new_[88103]_ , \new_[88106]_ , \new_[88109]_ , \new_[88110]_ ,
    \new_[88113]_ , \new_[88117]_ , \new_[88118]_ , \new_[88119]_ ,
    \new_[88120]_ , \new_[88123]_ , \new_[88126]_ , \new_[88127]_ ,
    \new_[88130]_ , \new_[88133]_ , \new_[88134]_ , \new_[88135]_ ,
    \new_[88138]_ , \new_[88141]_ , \new_[88142]_ , \new_[88145]_ ,
    \new_[88149]_ , \new_[88150]_ , \new_[88151]_ , \new_[88152]_ ,
    \new_[88155]_ , \new_[88158]_ , \new_[88159]_ , \new_[88162]_ ,
    \new_[88165]_ , \new_[88166]_ , \new_[88167]_ , \new_[88170]_ ,
    \new_[88173]_ , \new_[88174]_ , \new_[88177]_ , \new_[88181]_ ,
    \new_[88182]_ , \new_[88183]_ , \new_[88184]_ , \new_[88187]_ ,
    \new_[88190]_ , \new_[88191]_ , \new_[88194]_ , \new_[88197]_ ,
    \new_[88198]_ , \new_[88199]_ , \new_[88202]_ , \new_[88205]_ ,
    \new_[88206]_ , \new_[88209]_ , \new_[88213]_ , \new_[88214]_ ,
    \new_[88215]_ , \new_[88216]_ , \new_[88219]_ , \new_[88222]_ ,
    \new_[88223]_ , \new_[88226]_ , \new_[88229]_ , \new_[88230]_ ,
    \new_[88231]_ , \new_[88234]_ , \new_[88237]_ , \new_[88238]_ ,
    \new_[88241]_ , \new_[88245]_ , \new_[88246]_ , \new_[88247]_ ,
    \new_[88248]_ , \new_[88251]_ , \new_[88254]_ , \new_[88255]_ ,
    \new_[88258]_ , \new_[88261]_ , \new_[88262]_ , \new_[88263]_ ,
    \new_[88266]_ , \new_[88269]_ , \new_[88270]_ , \new_[88273]_ ,
    \new_[88277]_ , \new_[88278]_ , \new_[88279]_ , \new_[88280]_ ,
    \new_[88283]_ , \new_[88286]_ , \new_[88287]_ , \new_[88290]_ ,
    \new_[88294]_ , \new_[88295]_ , \new_[88296]_ , \new_[88297]_ ,
    \new_[88300]_ , \new_[88303]_ , \new_[88304]_ , \new_[88307]_ ,
    \new_[88311]_ , \new_[88312]_ , \new_[88313]_ , \new_[88314]_ ,
    \new_[88317]_ , \new_[88320]_ , \new_[88321]_ , \new_[88324]_ ,
    \new_[88328]_ , \new_[88329]_ , \new_[88330]_ , \new_[88331]_ ,
    \new_[88334]_ , \new_[88337]_ , \new_[88338]_ , \new_[88341]_ ,
    \new_[88345]_ , \new_[88346]_ , \new_[88347]_ , \new_[88348]_ ,
    \new_[88351]_ , \new_[88354]_ , \new_[88355]_ , \new_[88358]_ ,
    \new_[88362]_ , \new_[88363]_ , \new_[88364]_ , \new_[88365]_ ,
    \new_[88368]_ , \new_[88371]_ , \new_[88372]_ , \new_[88375]_ ,
    \new_[88379]_ , \new_[88380]_ , \new_[88381]_ , \new_[88382]_ ,
    \new_[88385]_ , \new_[88388]_ , \new_[88389]_ , \new_[88392]_ ,
    \new_[88396]_ , \new_[88397]_ , \new_[88398]_ , \new_[88399]_ ,
    \new_[88402]_ , \new_[88405]_ , \new_[88406]_ , \new_[88409]_ ,
    \new_[88413]_ , \new_[88414]_ , \new_[88415]_ , \new_[88416]_ ,
    \new_[88419]_ , \new_[88422]_ , \new_[88423]_ , \new_[88426]_ ,
    \new_[88430]_ , \new_[88431]_ , \new_[88432]_ , \new_[88433]_ ,
    \new_[88436]_ , \new_[88439]_ , \new_[88440]_ , \new_[88443]_ ,
    \new_[88447]_ , \new_[88448]_ , \new_[88449]_ , \new_[88450]_ ,
    \new_[88453]_ , \new_[88456]_ , \new_[88457]_ , \new_[88460]_ ,
    \new_[88464]_ , \new_[88465]_ , \new_[88466]_ , \new_[88467]_ ,
    \new_[88470]_ , \new_[88473]_ , \new_[88474]_ , \new_[88477]_ ,
    \new_[88481]_ , \new_[88482]_ , \new_[88483]_ , \new_[88484]_ ,
    \new_[88487]_ , \new_[88490]_ , \new_[88491]_ , \new_[88494]_ ,
    \new_[88498]_ , \new_[88499]_ , \new_[88500]_ , \new_[88501]_ ,
    \new_[88504]_ , \new_[88507]_ , \new_[88508]_ , \new_[88511]_ ,
    \new_[88515]_ , \new_[88516]_ , \new_[88517]_ , \new_[88518]_ ,
    \new_[88521]_ , \new_[88524]_ , \new_[88525]_ , \new_[88528]_ ,
    \new_[88532]_ , \new_[88533]_ , \new_[88534]_ , \new_[88535]_ ,
    \new_[88538]_ , \new_[88541]_ , \new_[88542]_ , \new_[88545]_ ,
    \new_[88549]_ , \new_[88550]_ , \new_[88551]_ , \new_[88552]_ ,
    \new_[88555]_ , \new_[88558]_ , \new_[88559]_ , \new_[88562]_ ,
    \new_[88566]_ , \new_[88567]_ , \new_[88568]_ , \new_[88569]_ ,
    \new_[88572]_ , \new_[88575]_ , \new_[88576]_ , \new_[88579]_ ,
    \new_[88583]_ , \new_[88584]_ , \new_[88585]_ , \new_[88586]_ ,
    \new_[88589]_ , \new_[88592]_ , \new_[88593]_ , \new_[88596]_ ,
    \new_[88600]_ , \new_[88601]_ , \new_[88602]_ , \new_[88603]_ ,
    \new_[88606]_ , \new_[88609]_ , \new_[88610]_ , \new_[88613]_ ,
    \new_[88617]_ , \new_[88618]_ , \new_[88619]_ , \new_[88620]_ ,
    \new_[88623]_ , \new_[88626]_ , \new_[88627]_ , \new_[88630]_ ,
    \new_[88634]_ , \new_[88635]_ , \new_[88636]_ , \new_[88637]_ ,
    \new_[88640]_ , \new_[88643]_ , \new_[88644]_ , \new_[88647]_ ,
    \new_[88651]_ , \new_[88652]_ , \new_[88653]_ , \new_[88654]_ ,
    \new_[88657]_ , \new_[88660]_ , \new_[88661]_ , \new_[88664]_ ,
    \new_[88668]_ , \new_[88669]_ , \new_[88670]_ , \new_[88671]_ ,
    \new_[88674]_ , \new_[88677]_ , \new_[88678]_ , \new_[88681]_ ,
    \new_[88685]_ , \new_[88686]_ , \new_[88687]_ , \new_[88688]_ ;
  assign A105 = \new_[9520]_  | \new_[6347]_ ;
  assign \new_[1]_  = \new_[88688]_  & \new_[88671]_ ;
  assign \new_[2]_  = \new_[88654]_  & \new_[88637]_ ;
  assign \new_[3]_  = \new_[88620]_  & \new_[88603]_ ;
  assign \new_[4]_  = \new_[88586]_  & \new_[88569]_ ;
  assign \new_[5]_  = \new_[88552]_  & \new_[88535]_ ;
  assign \new_[6]_  = \new_[88518]_  & \new_[88501]_ ;
  assign \new_[7]_  = \new_[88484]_  & \new_[88467]_ ;
  assign \new_[8]_  = \new_[88450]_  & \new_[88433]_ ;
  assign \new_[9]_  = \new_[88416]_  & \new_[88399]_ ;
  assign \new_[10]_  = \new_[88382]_  & \new_[88365]_ ;
  assign \new_[11]_  = \new_[88348]_  & \new_[88331]_ ;
  assign \new_[12]_  = \new_[88314]_  & \new_[88297]_ ;
  assign \new_[13]_  = \new_[88280]_  & \new_[88263]_ ;
  assign \new_[14]_  = \new_[88248]_  & \new_[88231]_ ;
  assign \new_[15]_  = \new_[88216]_  & \new_[88199]_ ;
  assign \new_[16]_  = \new_[88184]_  & \new_[88167]_ ;
  assign \new_[17]_  = \new_[88152]_  & \new_[88135]_ ;
  assign \new_[18]_  = \new_[88120]_  & \new_[88103]_ ;
  assign \new_[19]_  = \new_[88088]_  & \new_[88071]_ ;
  assign \new_[20]_  = \new_[88056]_  & \new_[88039]_ ;
  assign \new_[21]_  = \new_[88024]_  & \new_[88007]_ ;
  assign \new_[22]_  = \new_[87992]_  & \new_[87975]_ ;
  assign \new_[23]_  = \new_[87960]_  & \new_[87943]_ ;
  assign \new_[24]_  = \new_[87928]_  & \new_[87911]_ ;
  assign \new_[25]_  = \new_[87896]_  & \new_[87879]_ ;
  assign \new_[26]_  = \new_[87864]_  & \new_[87847]_ ;
  assign \new_[27]_  = \new_[87832]_  & \new_[87815]_ ;
  assign \new_[28]_  = \new_[87800]_  & \new_[87783]_ ;
  assign \new_[29]_  = \new_[87768]_  & \new_[87751]_ ;
  assign \new_[30]_  = \new_[87736]_  & \new_[87719]_ ;
  assign \new_[31]_  = \new_[87704]_  & \new_[87687]_ ;
  assign \new_[32]_  = \new_[87672]_  & \new_[87655]_ ;
  assign \new_[33]_  = \new_[87640]_  & \new_[87623]_ ;
  assign \new_[34]_  = \new_[87608]_  & \new_[87591]_ ;
  assign \new_[35]_  = \new_[87576]_  & \new_[87559]_ ;
  assign \new_[36]_  = \new_[87544]_  & \new_[87527]_ ;
  assign \new_[37]_  = \new_[87512]_  & \new_[87495]_ ;
  assign \new_[38]_  = \new_[87480]_  & \new_[87463]_ ;
  assign \new_[39]_  = \new_[87448]_  & \new_[87431]_ ;
  assign \new_[40]_  = \new_[87416]_  & \new_[87399]_ ;
  assign \new_[41]_  = \new_[87384]_  & \new_[87367]_ ;
  assign \new_[42]_  = \new_[87352]_  & \new_[87335]_ ;
  assign \new_[43]_  = \new_[87320]_  & \new_[87303]_ ;
  assign \new_[44]_  = \new_[87288]_  & \new_[87271]_ ;
  assign \new_[45]_  = \new_[87256]_  & \new_[87239]_ ;
  assign \new_[46]_  = \new_[87224]_  & \new_[87207]_ ;
  assign \new_[47]_  = \new_[87192]_  & \new_[87175]_ ;
  assign \new_[48]_  = \new_[87160]_  & \new_[87143]_ ;
  assign \new_[49]_  = \new_[87128]_  & \new_[87111]_ ;
  assign \new_[50]_  = \new_[87096]_  & \new_[87079]_ ;
  assign \new_[51]_  = \new_[87064]_  & \new_[87047]_ ;
  assign \new_[52]_  = \new_[87032]_  & \new_[87015]_ ;
  assign \new_[53]_  = \new_[87000]_  & \new_[86983]_ ;
  assign \new_[54]_  = \new_[86968]_  & \new_[86951]_ ;
  assign \new_[55]_  = \new_[86936]_  & \new_[86919]_ ;
  assign \new_[56]_  = \new_[86904]_  & \new_[86887]_ ;
  assign \new_[57]_  = \new_[86872]_  & \new_[86855]_ ;
  assign \new_[58]_  = \new_[86840]_  & \new_[86823]_ ;
  assign \new_[59]_  = \new_[86808]_  & \new_[86791]_ ;
  assign \new_[60]_  = \new_[86776]_  & \new_[86759]_ ;
  assign \new_[61]_  = \new_[86744]_  & \new_[86727]_ ;
  assign \new_[62]_  = \new_[86712]_  & \new_[86695]_ ;
  assign \new_[63]_  = \new_[86680]_  & \new_[86663]_ ;
  assign \new_[64]_  = \new_[86648]_  & \new_[86631]_ ;
  assign \new_[65]_  = \new_[86616]_  & \new_[86599]_ ;
  assign \new_[66]_  = \new_[86584]_  & \new_[86567]_ ;
  assign \new_[67]_  = \new_[86552]_  & \new_[86535]_ ;
  assign \new_[68]_  = \new_[86520]_  & \new_[86503]_ ;
  assign \new_[69]_  = \new_[86488]_  & \new_[86471]_ ;
  assign \new_[70]_  = \new_[86456]_  & \new_[86439]_ ;
  assign \new_[71]_  = \new_[86424]_  & \new_[86407]_ ;
  assign \new_[72]_  = \new_[86392]_  & \new_[86375]_ ;
  assign \new_[73]_  = \new_[86360]_  & \new_[86343]_ ;
  assign \new_[74]_  = \new_[86328]_  & \new_[86311]_ ;
  assign \new_[75]_  = \new_[86296]_  & \new_[86279]_ ;
  assign \new_[76]_  = \new_[86264]_  & \new_[86247]_ ;
  assign \new_[77]_  = \new_[86232]_  & \new_[86215]_ ;
  assign \new_[78]_  = \new_[86200]_  & \new_[86183]_ ;
  assign \new_[79]_  = \new_[86168]_  & \new_[86151]_ ;
  assign \new_[80]_  = \new_[86136]_  & \new_[86119]_ ;
  assign \new_[81]_  = \new_[86104]_  & \new_[86087]_ ;
  assign \new_[82]_  = \new_[86072]_  & \new_[86055]_ ;
  assign \new_[83]_  = \new_[86040]_  & \new_[86023]_ ;
  assign \new_[84]_  = \new_[86008]_  & \new_[85991]_ ;
  assign \new_[85]_  = \new_[85976]_  & \new_[85959]_ ;
  assign \new_[86]_  = \new_[85944]_  & \new_[85927]_ ;
  assign \new_[87]_  = \new_[85912]_  & \new_[85895]_ ;
  assign \new_[88]_  = \new_[85880]_  & \new_[85863]_ ;
  assign \new_[89]_  = \new_[85848]_  & \new_[85831]_ ;
  assign \new_[90]_  = \new_[85816]_  & \new_[85799]_ ;
  assign \new_[91]_  = \new_[85784]_  & \new_[85767]_ ;
  assign \new_[92]_  = \new_[85752]_  & \new_[85735]_ ;
  assign \new_[93]_  = \new_[85720]_  & \new_[85703]_ ;
  assign \new_[94]_  = \new_[85688]_  & \new_[85671]_ ;
  assign \new_[95]_  = \new_[85656]_  & \new_[85639]_ ;
  assign \new_[96]_  = \new_[85624]_  & \new_[85607]_ ;
  assign \new_[97]_  = \new_[85592]_  & \new_[85575]_ ;
  assign \new_[98]_  = \new_[85560]_  & \new_[85543]_ ;
  assign \new_[99]_  = \new_[85528]_  & \new_[85511]_ ;
  assign \new_[100]_  = \new_[85496]_  & \new_[85479]_ ;
  assign \new_[101]_  = \new_[85464]_  & \new_[85447]_ ;
  assign \new_[102]_  = \new_[85432]_  & \new_[85415]_ ;
  assign \new_[103]_  = \new_[85400]_  & \new_[85383]_ ;
  assign \new_[104]_  = \new_[85368]_  & \new_[85351]_ ;
  assign \new_[105]_  = \new_[85336]_  & \new_[85319]_ ;
  assign \new_[106]_  = \new_[85304]_  & \new_[85287]_ ;
  assign \new_[107]_  = \new_[85272]_  & \new_[85255]_ ;
  assign \new_[108]_  = \new_[85240]_  & \new_[85223]_ ;
  assign \new_[109]_  = \new_[85208]_  & \new_[85191]_ ;
  assign \new_[110]_  = \new_[85176]_  & \new_[85159]_ ;
  assign \new_[111]_  = \new_[85144]_  & \new_[85127]_ ;
  assign \new_[112]_  = \new_[85112]_  & \new_[85095]_ ;
  assign \new_[113]_  = \new_[85080]_  & \new_[85063]_ ;
  assign \new_[114]_  = \new_[85048]_  & \new_[85031]_ ;
  assign \new_[115]_  = \new_[85016]_  & \new_[84999]_ ;
  assign \new_[116]_  = \new_[84984]_  & \new_[84967]_ ;
  assign \new_[117]_  = \new_[84952]_  & \new_[84937]_ ;
  assign \new_[118]_  = \new_[84922]_  & \new_[84907]_ ;
  assign \new_[119]_  = \new_[84892]_  & \new_[84877]_ ;
  assign \new_[120]_  = \new_[84862]_  & \new_[84847]_ ;
  assign \new_[121]_  = \new_[84832]_  & \new_[84817]_ ;
  assign \new_[122]_  = \new_[84802]_  & \new_[84787]_ ;
  assign \new_[123]_  = \new_[84772]_  & \new_[84757]_ ;
  assign \new_[124]_  = \new_[84742]_  & \new_[84727]_ ;
  assign \new_[125]_  = \new_[84712]_  & \new_[84697]_ ;
  assign \new_[126]_  = \new_[84682]_  & \new_[84667]_ ;
  assign \new_[127]_  = \new_[84652]_  & \new_[84637]_ ;
  assign \new_[128]_  = \new_[84622]_  & \new_[84607]_ ;
  assign \new_[129]_  = \new_[84592]_  & \new_[84577]_ ;
  assign \new_[130]_  = \new_[84562]_  & \new_[84547]_ ;
  assign \new_[131]_  = \new_[84532]_  & \new_[84517]_ ;
  assign \new_[132]_  = \new_[84502]_  & \new_[84487]_ ;
  assign \new_[133]_  = \new_[84472]_  & \new_[84457]_ ;
  assign \new_[134]_  = \new_[84442]_  & \new_[84427]_ ;
  assign \new_[135]_  = \new_[84412]_  & \new_[84397]_ ;
  assign \new_[136]_  = \new_[84382]_  & \new_[84367]_ ;
  assign \new_[137]_  = \new_[84352]_  & \new_[84337]_ ;
  assign \new_[138]_  = \new_[84322]_  & \new_[84307]_ ;
  assign \new_[139]_  = \new_[84292]_  & \new_[84277]_ ;
  assign \new_[140]_  = \new_[84262]_  & \new_[84247]_ ;
  assign \new_[141]_  = \new_[84232]_  & \new_[84217]_ ;
  assign \new_[142]_  = \new_[84202]_  & \new_[84187]_ ;
  assign \new_[143]_  = \new_[84172]_  & \new_[84157]_ ;
  assign \new_[144]_  = \new_[84142]_  & \new_[84127]_ ;
  assign \new_[145]_  = \new_[84112]_  & \new_[84097]_ ;
  assign \new_[146]_  = \new_[84082]_  & \new_[84067]_ ;
  assign \new_[147]_  = \new_[84052]_  & \new_[84037]_ ;
  assign \new_[148]_  = \new_[84022]_  & \new_[84007]_ ;
  assign \new_[149]_  = \new_[83992]_  & \new_[83977]_ ;
  assign \new_[150]_  = \new_[83962]_  & \new_[83947]_ ;
  assign \new_[151]_  = \new_[83932]_  & \new_[83917]_ ;
  assign \new_[152]_  = \new_[83902]_  & \new_[83887]_ ;
  assign \new_[153]_  = \new_[83872]_  & \new_[83857]_ ;
  assign \new_[154]_  = \new_[83842]_  & \new_[83827]_ ;
  assign \new_[155]_  = \new_[83812]_  & \new_[83797]_ ;
  assign \new_[156]_  = \new_[83782]_  & \new_[83767]_ ;
  assign \new_[157]_  = \new_[83752]_  & \new_[83737]_ ;
  assign \new_[158]_  = \new_[83722]_  & \new_[83707]_ ;
  assign \new_[159]_  = \new_[83692]_  & \new_[83677]_ ;
  assign \new_[160]_  = \new_[83662]_  & \new_[83647]_ ;
  assign \new_[161]_  = \new_[83632]_  & \new_[83617]_ ;
  assign \new_[162]_  = \new_[83602]_  & \new_[83587]_ ;
  assign \new_[163]_  = \new_[83572]_  & \new_[83557]_ ;
  assign \new_[164]_  = \new_[83542]_  & \new_[83527]_ ;
  assign \new_[165]_  = \new_[83512]_  & \new_[83497]_ ;
  assign \new_[166]_  = \new_[83482]_  & \new_[83467]_ ;
  assign \new_[167]_  = \new_[83452]_  & \new_[83437]_ ;
  assign \new_[168]_  = \new_[83422]_  & \new_[83407]_ ;
  assign \new_[169]_  = \new_[83392]_  & \new_[83377]_ ;
  assign \new_[170]_  = \new_[83362]_  & \new_[83347]_ ;
  assign \new_[171]_  = \new_[83332]_  & \new_[83317]_ ;
  assign \new_[172]_  = \new_[83302]_  & \new_[83287]_ ;
  assign \new_[173]_  = \new_[83272]_  & \new_[83257]_ ;
  assign \new_[174]_  = \new_[83242]_  & \new_[83227]_ ;
  assign \new_[175]_  = \new_[83212]_  & \new_[83197]_ ;
  assign \new_[176]_  = \new_[83182]_  & \new_[83167]_ ;
  assign \new_[177]_  = \new_[83152]_  & \new_[83137]_ ;
  assign \new_[178]_  = \new_[83122]_  & \new_[83107]_ ;
  assign \new_[179]_  = \new_[83092]_  & \new_[83077]_ ;
  assign \new_[180]_  = \new_[83062]_  & \new_[83047]_ ;
  assign \new_[181]_  = \new_[83032]_  & \new_[83017]_ ;
  assign \new_[182]_  = \new_[83002]_  & \new_[82987]_ ;
  assign \new_[183]_  = \new_[82972]_  & \new_[82957]_ ;
  assign \new_[184]_  = \new_[82942]_  & \new_[82927]_ ;
  assign \new_[185]_  = \new_[82912]_  & \new_[82897]_ ;
  assign \new_[186]_  = \new_[82882]_  & \new_[82867]_ ;
  assign \new_[187]_  = \new_[82852]_  & \new_[82837]_ ;
  assign \new_[188]_  = \new_[82822]_  & \new_[82807]_ ;
  assign \new_[189]_  = \new_[82792]_  & \new_[82777]_ ;
  assign \new_[190]_  = \new_[82762]_  & \new_[82747]_ ;
  assign \new_[191]_  = \new_[82732]_  & \new_[82717]_ ;
  assign \new_[192]_  = \new_[82702]_  & \new_[82687]_ ;
  assign \new_[193]_  = \new_[82672]_  & \new_[82657]_ ;
  assign \new_[194]_  = \new_[82642]_  & \new_[82627]_ ;
  assign \new_[195]_  = \new_[82612]_  & \new_[82597]_ ;
  assign \new_[196]_  = \new_[82582]_  & \new_[82567]_ ;
  assign \new_[197]_  = \new_[82552]_  & \new_[82537]_ ;
  assign \new_[198]_  = \new_[82522]_  & \new_[82507]_ ;
  assign \new_[199]_  = \new_[82492]_  & \new_[82477]_ ;
  assign \new_[200]_  = \new_[82462]_  & \new_[82447]_ ;
  assign \new_[201]_  = \new_[82432]_  & \new_[82417]_ ;
  assign \new_[202]_  = \new_[82402]_  & \new_[82387]_ ;
  assign \new_[203]_  = \new_[82372]_  & \new_[82357]_ ;
  assign \new_[204]_  = \new_[82342]_  & \new_[82327]_ ;
  assign \new_[205]_  = \new_[82312]_  & \new_[82297]_ ;
  assign \new_[206]_  = \new_[82282]_  & \new_[82267]_ ;
  assign \new_[207]_  = \new_[82252]_  & \new_[82237]_ ;
  assign \new_[208]_  = \new_[82222]_  & \new_[82207]_ ;
  assign \new_[209]_  = \new_[82192]_  & \new_[82177]_ ;
  assign \new_[210]_  = \new_[82162]_  & \new_[82147]_ ;
  assign \new_[211]_  = \new_[82132]_  & \new_[82117]_ ;
  assign \new_[212]_  = \new_[82102]_  & \new_[82087]_ ;
  assign \new_[213]_  = \new_[82072]_  & \new_[82057]_ ;
  assign \new_[214]_  = \new_[82042]_  & \new_[82027]_ ;
  assign \new_[215]_  = \new_[82012]_  & \new_[81997]_ ;
  assign \new_[216]_  = \new_[81982]_  & \new_[81967]_ ;
  assign \new_[217]_  = \new_[81952]_  & \new_[81937]_ ;
  assign \new_[218]_  = \new_[81922]_  & \new_[81907]_ ;
  assign \new_[219]_  = \new_[81892]_  & \new_[81877]_ ;
  assign \new_[220]_  = \new_[81862]_  & \new_[81847]_ ;
  assign \new_[221]_  = \new_[81832]_  & \new_[81817]_ ;
  assign \new_[222]_  = \new_[81802]_  & \new_[81787]_ ;
  assign \new_[223]_  = \new_[81772]_  & \new_[81757]_ ;
  assign \new_[224]_  = \new_[81742]_  & \new_[81727]_ ;
  assign \new_[225]_  = \new_[81712]_  & \new_[81697]_ ;
  assign \new_[226]_  = \new_[81682]_  & \new_[81667]_ ;
  assign \new_[227]_  = \new_[81652]_  & \new_[81637]_ ;
  assign \new_[228]_  = \new_[81622]_  & \new_[81607]_ ;
  assign \new_[229]_  = \new_[81592]_  & \new_[81577]_ ;
  assign \new_[230]_  = \new_[81562]_  & \new_[81547]_ ;
  assign \new_[231]_  = \new_[81532]_  & \new_[81517]_ ;
  assign \new_[232]_  = \new_[81502]_  & \new_[81487]_ ;
  assign \new_[233]_  = \new_[81472]_  & \new_[81457]_ ;
  assign \new_[234]_  = \new_[81442]_  & \new_[81427]_ ;
  assign \new_[235]_  = \new_[81412]_  & \new_[81397]_ ;
  assign \new_[236]_  = \new_[81382]_  & \new_[81367]_ ;
  assign \new_[237]_  = \new_[81352]_  & \new_[81337]_ ;
  assign \new_[238]_  = \new_[81322]_  & \new_[81307]_ ;
  assign \new_[239]_  = \new_[81292]_  & \new_[81277]_ ;
  assign \new_[240]_  = \new_[81262]_  & \new_[81247]_ ;
  assign \new_[241]_  = \new_[81232]_  & \new_[81217]_ ;
  assign \new_[242]_  = \new_[81202]_  & \new_[81187]_ ;
  assign \new_[243]_  = \new_[81172]_  & \new_[81157]_ ;
  assign \new_[244]_  = \new_[81142]_  & \new_[81127]_ ;
  assign \new_[245]_  = \new_[81112]_  & \new_[81097]_ ;
  assign \new_[246]_  = \new_[81082]_  & \new_[81067]_ ;
  assign \new_[247]_  = \new_[81052]_  & \new_[81037]_ ;
  assign \new_[248]_  = \new_[81022]_  & \new_[81007]_ ;
  assign \new_[249]_  = \new_[80992]_  & \new_[80977]_ ;
  assign \new_[250]_  = \new_[80962]_  & \new_[80947]_ ;
  assign \new_[251]_  = \new_[80932]_  & \new_[80917]_ ;
  assign \new_[252]_  = \new_[80902]_  & \new_[80887]_ ;
  assign \new_[253]_  = \new_[80872]_  & \new_[80857]_ ;
  assign \new_[254]_  = \new_[80842]_  & \new_[80827]_ ;
  assign \new_[255]_  = \new_[80812]_  & \new_[80797]_ ;
  assign \new_[256]_  = \new_[80782]_  & \new_[80767]_ ;
  assign \new_[257]_  = \new_[80752]_  & \new_[80737]_ ;
  assign \new_[258]_  = \new_[80722]_  & \new_[80707]_ ;
  assign \new_[259]_  = \new_[80692]_  & \new_[80677]_ ;
  assign \new_[260]_  = \new_[80662]_  & \new_[80647]_ ;
  assign \new_[261]_  = \new_[80632]_  & \new_[80617]_ ;
  assign \new_[262]_  = \new_[80602]_  & \new_[80587]_ ;
  assign \new_[263]_  = \new_[80572]_  & \new_[80557]_ ;
  assign \new_[264]_  = \new_[80542]_  & \new_[80527]_ ;
  assign \new_[265]_  = \new_[80512]_  & \new_[80497]_ ;
  assign \new_[266]_  = \new_[80482]_  & \new_[80467]_ ;
  assign \new_[267]_  = \new_[80452]_  & \new_[80437]_ ;
  assign \new_[268]_  = \new_[80422]_  & \new_[80407]_ ;
  assign \new_[269]_  = \new_[80392]_  & \new_[80377]_ ;
  assign \new_[270]_  = \new_[80362]_  & \new_[80347]_ ;
  assign \new_[271]_  = \new_[80332]_  & \new_[80317]_ ;
  assign \new_[272]_  = \new_[80302]_  & \new_[80287]_ ;
  assign \new_[273]_  = \new_[80272]_  & \new_[80257]_ ;
  assign \new_[274]_  = \new_[80242]_  & \new_[80227]_ ;
  assign \new_[275]_  = \new_[80212]_  & \new_[80197]_ ;
  assign \new_[276]_  = \new_[80182]_  & \new_[80167]_ ;
  assign \new_[277]_  = \new_[80152]_  & \new_[80137]_ ;
  assign \new_[278]_  = \new_[80122]_  & \new_[80107]_ ;
  assign \new_[279]_  = \new_[80092]_  & \new_[80077]_ ;
  assign \new_[280]_  = \new_[80062]_  & \new_[80047]_ ;
  assign \new_[281]_  = \new_[80032]_  & \new_[80017]_ ;
  assign \new_[282]_  = \new_[80002]_  & \new_[79987]_ ;
  assign \new_[283]_  = \new_[79972]_  & \new_[79957]_ ;
  assign \new_[284]_  = \new_[79942]_  & \new_[79927]_ ;
  assign \new_[285]_  = \new_[79912]_  & \new_[79897]_ ;
  assign \new_[286]_  = \new_[79882]_  & \new_[79867]_ ;
  assign \new_[287]_  = \new_[79852]_  & \new_[79837]_ ;
  assign \new_[288]_  = \new_[79822]_  & \new_[79807]_ ;
  assign \new_[289]_  = \new_[79792]_  & \new_[79777]_ ;
  assign \new_[290]_  = \new_[79762]_  & \new_[79747]_ ;
  assign \new_[291]_  = \new_[79732]_  & \new_[79717]_ ;
  assign \new_[292]_  = \new_[79702]_  & \new_[79687]_ ;
  assign \new_[293]_  = \new_[79672]_  & \new_[79657]_ ;
  assign \new_[294]_  = \new_[79642]_  & \new_[79627]_ ;
  assign \new_[295]_  = \new_[79612]_  & \new_[79597]_ ;
  assign \new_[296]_  = \new_[79582]_  & \new_[79567]_ ;
  assign \new_[297]_  = \new_[79552]_  & \new_[79537]_ ;
  assign \new_[298]_  = \new_[79522]_  & \new_[79507]_ ;
  assign \new_[299]_  = \new_[79492]_  & \new_[79477]_ ;
  assign \new_[300]_  = \new_[79462]_  & \new_[79447]_ ;
  assign \new_[301]_  = \new_[79432]_  & \new_[79417]_ ;
  assign \new_[302]_  = \new_[79402]_  & \new_[79387]_ ;
  assign \new_[303]_  = \new_[79372]_  & \new_[79357]_ ;
  assign \new_[304]_  = \new_[79342]_  & \new_[79327]_ ;
  assign \new_[305]_  = \new_[79312]_  & \new_[79297]_ ;
  assign \new_[306]_  = \new_[79282]_  & \new_[79267]_ ;
  assign \new_[307]_  = \new_[79252]_  & \new_[79237]_ ;
  assign \new_[308]_  = \new_[79222]_  & \new_[79207]_ ;
  assign \new_[309]_  = \new_[79192]_  & \new_[79177]_ ;
  assign \new_[310]_  = \new_[79162]_  & \new_[79147]_ ;
  assign \new_[311]_  = \new_[79132]_  & \new_[79117]_ ;
  assign \new_[312]_  = \new_[79102]_  & \new_[79087]_ ;
  assign \new_[313]_  = \new_[79072]_  & \new_[79057]_ ;
  assign \new_[314]_  = \new_[79042]_  & \new_[79027]_ ;
  assign \new_[315]_  = \new_[79012]_  & \new_[78997]_ ;
  assign \new_[316]_  = \new_[78982]_  & \new_[78967]_ ;
  assign \new_[317]_  = \new_[78952]_  & \new_[78937]_ ;
  assign \new_[318]_  = \new_[78922]_  & \new_[78907]_ ;
  assign \new_[319]_  = \new_[78892]_  & \new_[78877]_ ;
  assign \new_[320]_  = \new_[78862]_  & \new_[78847]_ ;
  assign \new_[321]_  = \new_[78832]_  & \new_[78817]_ ;
  assign \new_[322]_  = \new_[78802]_  & \new_[78787]_ ;
  assign \new_[323]_  = \new_[78772]_  & \new_[78757]_ ;
  assign \new_[324]_  = \new_[78742]_  & \new_[78727]_ ;
  assign \new_[325]_  = \new_[78712]_  & \new_[78697]_ ;
  assign \new_[326]_  = \new_[78682]_  & \new_[78667]_ ;
  assign \new_[327]_  = \new_[78652]_  & \new_[78637]_ ;
  assign \new_[328]_  = \new_[78622]_  & \new_[78607]_ ;
  assign \new_[329]_  = \new_[78592]_  & \new_[78577]_ ;
  assign \new_[330]_  = \new_[78562]_  & \new_[78547]_ ;
  assign \new_[331]_  = \new_[78532]_  & \new_[78517]_ ;
  assign \new_[332]_  = \new_[78502]_  & \new_[78487]_ ;
  assign \new_[333]_  = \new_[78472]_  & \new_[78457]_ ;
  assign \new_[334]_  = \new_[78442]_  & \new_[78427]_ ;
  assign \new_[335]_  = \new_[78412]_  & \new_[78397]_ ;
  assign \new_[336]_  = \new_[78382]_  & \new_[78367]_ ;
  assign \new_[337]_  = \new_[78352]_  & \new_[78337]_ ;
  assign \new_[338]_  = \new_[78322]_  & \new_[78307]_ ;
  assign \new_[339]_  = \new_[78292]_  & \new_[78277]_ ;
  assign \new_[340]_  = \new_[78262]_  & \new_[78247]_ ;
  assign \new_[341]_  = \new_[78232]_  & \new_[78217]_ ;
  assign \new_[342]_  = \new_[78202]_  & \new_[78187]_ ;
  assign \new_[343]_  = \new_[78172]_  & \new_[78157]_ ;
  assign \new_[344]_  = \new_[78142]_  & \new_[78127]_ ;
  assign \new_[345]_  = \new_[78112]_  & \new_[78097]_ ;
  assign \new_[346]_  = \new_[78082]_  & \new_[78067]_ ;
  assign \new_[347]_  = \new_[78052]_  & \new_[78037]_ ;
  assign \new_[348]_  = \new_[78022]_  & \new_[78007]_ ;
  assign \new_[349]_  = \new_[77992]_  & \new_[77977]_ ;
  assign \new_[350]_  = \new_[77962]_  & \new_[77947]_ ;
  assign \new_[351]_  = \new_[77932]_  & \new_[77917]_ ;
  assign \new_[352]_  = \new_[77902]_  & \new_[77887]_ ;
  assign \new_[353]_  = \new_[77872]_  & \new_[77857]_ ;
  assign \new_[354]_  = \new_[77842]_  & \new_[77827]_ ;
  assign \new_[355]_  = \new_[77812]_  & \new_[77797]_ ;
  assign \new_[356]_  = \new_[77782]_  & \new_[77767]_ ;
  assign \new_[357]_  = \new_[77752]_  & \new_[77737]_ ;
  assign \new_[358]_  = \new_[77722]_  & \new_[77707]_ ;
  assign \new_[359]_  = \new_[77692]_  & \new_[77677]_ ;
  assign \new_[360]_  = \new_[77662]_  & \new_[77647]_ ;
  assign \new_[361]_  = \new_[77632]_  & \new_[77617]_ ;
  assign \new_[362]_  = \new_[77602]_  & \new_[77587]_ ;
  assign \new_[363]_  = \new_[77572]_  & \new_[77557]_ ;
  assign \new_[364]_  = \new_[77542]_  & \new_[77527]_ ;
  assign \new_[365]_  = \new_[77512]_  & \new_[77497]_ ;
  assign \new_[366]_  = \new_[77482]_  & \new_[77467]_ ;
  assign \new_[367]_  = \new_[77452]_  & \new_[77437]_ ;
  assign \new_[368]_  = \new_[77422]_  & \new_[77407]_ ;
  assign \new_[369]_  = \new_[77392]_  & \new_[77377]_ ;
  assign \new_[370]_  = \new_[77362]_  & \new_[77347]_ ;
  assign \new_[371]_  = \new_[77332]_  & \new_[77317]_ ;
  assign \new_[372]_  = \new_[77302]_  & \new_[77287]_ ;
  assign \new_[373]_  = \new_[77272]_  & \new_[77257]_ ;
  assign \new_[374]_  = \new_[77242]_  & \new_[77227]_ ;
  assign \new_[375]_  = \new_[77212]_  & \new_[77197]_ ;
  assign \new_[376]_  = \new_[77182]_  & \new_[77167]_ ;
  assign \new_[377]_  = \new_[77152]_  & \new_[77137]_ ;
  assign \new_[378]_  = \new_[77122]_  & \new_[77107]_ ;
  assign \new_[379]_  = \new_[77092]_  & \new_[77077]_ ;
  assign \new_[380]_  = \new_[77062]_  & \new_[77047]_ ;
  assign \new_[381]_  = \new_[77032]_  & \new_[77017]_ ;
  assign \new_[382]_  = \new_[77002]_  & \new_[76987]_ ;
  assign \new_[383]_  = \new_[76972]_  & \new_[76957]_ ;
  assign \new_[384]_  = \new_[76942]_  & \new_[76927]_ ;
  assign \new_[385]_  = \new_[76912]_  & \new_[76897]_ ;
  assign \new_[386]_  = \new_[76882]_  & \new_[76867]_ ;
  assign \new_[387]_  = \new_[76852]_  & \new_[76837]_ ;
  assign \new_[388]_  = \new_[76822]_  & \new_[76807]_ ;
  assign \new_[389]_  = \new_[76792]_  & \new_[76777]_ ;
  assign \new_[390]_  = \new_[76762]_  & \new_[76747]_ ;
  assign \new_[391]_  = \new_[76732]_  & \new_[76717]_ ;
  assign \new_[392]_  = \new_[76702]_  & \new_[76687]_ ;
  assign \new_[393]_  = \new_[76672]_  & \new_[76657]_ ;
  assign \new_[394]_  = \new_[76642]_  & \new_[76627]_ ;
  assign \new_[395]_  = \new_[76612]_  & \new_[76597]_ ;
  assign \new_[396]_  = \new_[76582]_  & \new_[76567]_ ;
  assign \new_[397]_  = \new_[76552]_  & \new_[76537]_ ;
  assign \new_[398]_  = \new_[76522]_  & \new_[76507]_ ;
  assign \new_[399]_  = \new_[76492]_  & \new_[76477]_ ;
  assign \new_[400]_  = \new_[76462]_  & \new_[76447]_ ;
  assign \new_[401]_  = \new_[76432]_  & \new_[76417]_ ;
  assign \new_[402]_  = \new_[76402]_  & \new_[76387]_ ;
  assign \new_[403]_  = \new_[76372]_  & \new_[76357]_ ;
  assign \new_[404]_  = \new_[76342]_  & \new_[76327]_ ;
  assign \new_[405]_  = \new_[76312]_  & \new_[76297]_ ;
  assign \new_[406]_  = \new_[76282]_  & \new_[76267]_ ;
  assign \new_[407]_  = \new_[76252]_  & \new_[76237]_ ;
  assign \new_[408]_  = \new_[76222]_  & \new_[76207]_ ;
  assign \new_[409]_  = \new_[76192]_  & \new_[76177]_ ;
  assign \new_[410]_  = \new_[76162]_  & \new_[76147]_ ;
  assign \new_[411]_  = \new_[76132]_  & \new_[76117]_ ;
  assign \new_[412]_  = \new_[76102]_  & \new_[76087]_ ;
  assign \new_[413]_  = \new_[76072]_  & \new_[76057]_ ;
  assign \new_[414]_  = \new_[76042]_  & \new_[76027]_ ;
  assign \new_[415]_  = \new_[76012]_  & \new_[75997]_ ;
  assign \new_[416]_  = \new_[75982]_  & \new_[75967]_ ;
  assign \new_[417]_  = \new_[75952]_  & \new_[75937]_ ;
  assign \new_[418]_  = \new_[75922]_  & \new_[75907]_ ;
  assign \new_[419]_  = \new_[75892]_  & \new_[75877]_ ;
  assign \new_[420]_  = \new_[75862]_  & \new_[75847]_ ;
  assign \new_[421]_  = \new_[75832]_  & \new_[75817]_ ;
  assign \new_[422]_  = \new_[75802]_  & \new_[75787]_ ;
  assign \new_[423]_  = \new_[75772]_  & \new_[75757]_ ;
  assign \new_[424]_  = \new_[75742]_  & \new_[75727]_ ;
  assign \new_[425]_  = \new_[75712]_  & \new_[75697]_ ;
  assign \new_[426]_  = \new_[75682]_  & \new_[75667]_ ;
  assign \new_[427]_  = \new_[75652]_  & \new_[75637]_ ;
  assign \new_[428]_  = \new_[75622]_  & \new_[75607]_ ;
  assign \new_[429]_  = \new_[75592]_  & \new_[75577]_ ;
  assign \new_[430]_  = \new_[75562]_  & \new_[75547]_ ;
  assign \new_[431]_  = \new_[75532]_  & \new_[75517]_ ;
  assign \new_[432]_  = \new_[75502]_  & \new_[75487]_ ;
  assign \new_[433]_  = \new_[75472]_  & \new_[75457]_ ;
  assign \new_[434]_  = \new_[75442]_  & \new_[75427]_ ;
  assign \new_[435]_  = \new_[75412]_  & \new_[75397]_ ;
  assign \new_[436]_  = \new_[75382]_  & \new_[75367]_ ;
  assign \new_[437]_  = \new_[75352]_  & \new_[75337]_ ;
  assign \new_[438]_  = \new_[75322]_  & \new_[75307]_ ;
  assign \new_[439]_  = \new_[75292]_  & \new_[75277]_ ;
  assign \new_[440]_  = \new_[75262]_  & \new_[75247]_ ;
  assign \new_[441]_  = \new_[75232]_  & \new_[75217]_ ;
  assign \new_[442]_  = \new_[75202]_  & \new_[75187]_ ;
  assign \new_[443]_  = \new_[75172]_  & \new_[75157]_ ;
  assign \new_[444]_  = \new_[75144]_  & \new_[75129]_ ;
  assign \new_[445]_  = \new_[75116]_  & \new_[75101]_ ;
  assign \new_[446]_  = \new_[75088]_  & \new_[75073]_ ;
  assign \new_[447]_  = \new_[75060]_  & \new_[75045]_ ;
  assign \new_[448]_  = \new_[75032]_  & \new_[75017]_ ;
  assign \new_[449]_  = \new_[75004]_  & \new_[74989]_ ;
  assign \new_[450]_  = \new_[74976]_  & \new_[74961]_ ;
  assign \new_[451]_  = \new_[74948]_  & \new_[74933]_ ;
  assign \new_[452]_  = \new_[74920]_  & \new_[74905]_ ;
  assign \new_[453]_  = \new_[74892]_  & \new_[74877]_ ;
  assign \new_[454]_  = \new_[74864]_  & \new_[74849]_ ;
  assign \new_[455]_  = \new_[74836]_  & \new_[74821]_ ;
  assign \new_[456]_  = \new_[74808]_  & \new_[74793]_ ;
  assign \new_[457]_  = \new_[74780]_  & \new_[74765]_ ;
  assign \new_[458]_  = \new_[74752]_  & \new_[74737]_ ;
  assign \new_[459]_  = \new_[74724]_  & \new_[74709]_ ;
  assign \new_[460]_  = \new_[74696]_  & \new_[74681]_ ;
  assign \new_[461]_  = \new_[74668]_  & \new_[74653]_ ;
  assign \new_[462]_  = \new_[74640]_  & \new_[74625]_ ;
  assign \new_[463]_  = \new_[74612]_  & \new_[74597]_ ;
  assign \new_[464]_  = \new_[74584]_  & \new_[74569]_ ;
  assign \new_[465]_  = \new_[74556]_  & \new_[74541]_ ;
  assign \new_[466]_  = \new_[74528]_  & \new_[74513]_ ;
  assign \new_[467]_  = \new_[74500]_  & \new_[74485]_ ;
  assign \new_[468]_  = \new_[74472]_  & \new_[74457]_ ;
  assign \new_[469]_  = \new_[74444]_  & \new_[74429]_ ;
  assign \new_[470]_  = \new_[74416]_  & \new_[74401]_ ;
  assign \new_[471]_  = \new_[74388]_  & \new_[74373]_ ;
  assign \new_[472]_  = \new_[74360]_  & \new_[74345]_ ;
  assign \new_[473]_  = \new_[74332]_  & \new_[74317]_ ;
  assign \new_[474]_  = \new_[74304]_  & \new_[74289]_ ;
  assign \new_[475]_  = \new_[74276]_  & \new_[74261]_ ;
  assign \new_[476]_  = \new_[74248]_  & \new_[74233]_ ;
  assign \new_[477]_  = \new_[74220]_  & \new_[74205]_ ;
  assign \new_[478]_  = \new_[74192]_  & \new_[74177]_ ;
  assign \new_[479]_  = \new_[74164]_  & \new_[74149]_ ;
  assign \new_[480]_  = \new_[74136]_  & \new_[74121]_ ;
  assign \new_[481]_  = \new_[74108]_  & \new_[74093]_ ;
  assign \new_[482]_  = \new_[74080]_  & \new_[74065]_ ;
  assign \new_[483]_  = \new_[74052]_  & \new_[74037]_ ;
  assign \new_[484]_  = \new_[74024]_  & \new_[74009]_ ;
  assign \new_[485]_  = \new_[73996]_  & \new_[73981]_ ;
  assign \new_[486]_  = \new_[73968]_  & \new_[73953]_ ;
  assign \new_[487]_  = \new_[73940]_  & \new_[73925]_ ;
  assign \new_[488]_  = \new_[73912]_  & \new_[73897]_ ;
  assign \new_[489]_  = \new_[73884]_  & \new_[73869]_ ;
  assign \new_[490]_  = \new_[73856]_  & \new_[73841]_ ;
  assign \new_[491]_  = \new_[73828]_  & \new_[73813]_ ;
  assign \new_[492]_  = \new_[73800]_  & \new_[73785]_ ;
  assign \new_[493]_  = \new_[73772]_  & \new_[73757]_ ;
  assign \new_[494]_  = \new_[73744]_  & \new_[73729]_ ;
  assign \new_[495]_  = \new_[73716]_  & \new_[73701]_ ;
  assign \new_[496]_  = \new_[73688]_  & \new_[73673]_ ;
  assign \new_[497]_  = \new_[73660]_  & \new_[73645]_ ;
  assign \new_[498]_  = \new_[73632]_  & \new_[73617]_ ;
  assign \new_[499]_  = \new_[73604]_  & \new_[73589]_ ;
  assign \new_[500]_  = \new_[73576]_  & \new_[73561]_ ;
  assign \new_[501]_  = \new_[73548]_  & \new_[73533]_ ;
  assign \new_[502]_  = \new_[73520]_  & \new_[73505]_ ;
  assign \new_[503]_  = \new_[73492]_  & \new_[73477]_ ;
  assign \new_[504]_  = \new_[73464]_  & \new_[73449]_ ;
  assign \new_[505]_  = \new_[73436]_  & \new_[73421]_ ;
  assign \new_[506]_  = \new_[73408]_  & \new_[73393]_ ;
  assign \new_[507]_  = \new_[73380]_  & \new_[73365]_ ;
  assign \new_[508]_  = \new_[73352]_  & \new_[73337]_ ;
  assign \new_[509]_  = \new_[73324]_  & \new_[73309]_ ;
  assign \new_[510]_  = \new_[73296]_  & \new_[73281]_ ;
  assign \new_[511]_  = \new_[73268]_  & \new_[73253]_ ;
  assign \new_[512]_  = \new_[73240]_  & \new_[73225]_ ;
  assign \new_[513]_  = \new_[73212]_  & \new_[73197]_ ;
  assign \new_[514]_  = \new_[73184]_  & \new_[73169]_ ;
  assign \new_[515]_  = \new_[73156]_  & \new_[73141]_ ;
  assign \new_[516]_  = \new_[73128]_  & \new_[73113]_ ;
  assign \new_[517]_  = \new_[73100]_  & \new_[73085]_ ;
  assign \new_[518]_  = \new_[73072]_  & \new_[73057]_ ;
  assign \new_[519]_  = \new_[73044]_  & \new_[73029]_ ;
  assign \new_[520]_  = \new_[73016]_  & \new_[73001]_ ;
  assign \new_[521]_  = \new_[72988]_  & \new_[72973]_ ;
  assign \new_[522]_  = \new_[72960]_  & \new_[72945]_ ;
  assign \new_[523]_  = \new_[72932]_  & \new_[72917]_ ;
  assign \new_[524]_  = \new_[72904]_  & \new_[72889]_ ;
  assign \new_[525]_  = \new_[72876]_  & \new_[72861]_ ;
  assign \new_[526]_  = \new_[72848]_  & \new_[72833]_ ;
  assign \new_[527]_  = \new_[72820]_  & \new_[72805]_ ;
  assign \new_[528]_  = \new_[72792]_  & \new_[72777]_ ;
  assign \new_[529]_  = \new_[72764]_  & \new_[72749]_ ;
  assign \new_[530]_  = \new_[72736]_  & \new_[72721]_ ;
  assign \new_[531]_  = \new_[72708]_  & \new_[72693]_ ;
  assign \new_[532]_  = \new_[72680]_  & \new_[72665]_ ;
  assign \new_[533]_  = \new_[72652]_  & \new_[72637]_ ;
  assign \new_[534]_  = \new_[72624]_  & \new_[72609]_ ;
  assign \new_[535]_  = \new_[72596]_  & \new_[72581]_ ;
  assign \new_[536]_  = \new_[72568]_  & \new_[72553]_ ;
  assign \new_[537]_  = \new_[72540]_  & \new_[72525]_ ;
  assign \new_[538]_  = \new_[72512]_  & \new_[72497]_ ;
  assign \new_[539]_  = \new_[72484]_  & \new_[72469]_ ;
  assign \new_[540]_  = \new_[72456]_  & \new_[72441]_ ;
  assign \new_[541]_  = \new_[72428]_  & \new_[72413]_ ;
  assign \new_[542]_  = \new_[72400]_  & \new_[72385]_ ;
  assign \new_[543]_  = \new_[72372]_  & \new_[72357]_ ;
  assign \new_[544]_  = \new_[72344]_  & \new_[72329]_ ;
  assign \new_[545]_  = \new_[72316]_  & \new_[72301]_ ;
  assign \new_[546]_  = \new_[72288]_  & \new_[72273]_ ;
  assign \new_[547]_  = \new_[72260]_  & \new_[72245]_ ;
  assign \new_[548]_  = \new_[72232]_  & \new_[72217]_ ;
  assign \new_[549]_  = \new_[72204]_  & \new_[72189]_ ;
  assign \new_[550]_  = \new_[72176]_  & \new_[72161]_ ;
  assign \new_[551]_  = \new_[72148]_  & \new_[72133]_ ;
  assign \new_[552]_  = \new_[72120]_  & \new_[72105]_ ;
  assign \new_[553]_  = \new_[72092]_  & \new_[72077]_ ;
  assign \new_[554]_  = \new_[72064]_  & \new_[72049]_ ;
  assign \new_[555]_  = \new_[72036]_  & \new_[72021]_ ;
  assign \new_[556]_  = \new_[72008]_  & \new_[71993]_ ;
  assign \new_[557]_  = \new_[71980]_  & \new_[71965]_ ;
  assign \new_[558]_  = \new_[71952]_  & \new_[71937]_ ;
  assign \new_[559]_  = \new_[71924]_  & \new_[71909]_ ;
  assign \new_[560]_  = \new_[71896]_  & \new_[71881]_ ;
  assign \new_[561]_  = \new_[71868]_  & \new_[71853]_ ;
  assign \new_[562]_  = \new_[71840]_  & \new_[71825]_ ;
  assign \new_[563]_  = \new_[71812]_  & \new_[71797]_ ;
  assign \new_[564]_  = \new_[71784]_  & \new_[71769]_ ;
  assign \new_[565]_  = \new_[71756]_  & \new_[71741]_ ;
  assign \new_[566]_  = \new_[71728]_  & \new_[71713]_ ;
  assign \new_[567]_  = \new_[71700]_  & \new_[71685]_ ;
  assign \new_[568]_  = \new_[71672]_  & \new_[71657]_ ;
  assign \new_[569]_  = \new_[71644]_  & \new_[71629]_ ;
  assign \new_[570]_  = \new_[71616]_  & \new_[71601]_ ;
  assign \new_[571]_  = \new_[71588]_  & \new_[71573]_ ;
  assign \new_[572]_  = \new_[71560]_  & \new_[71545]_ ;
  assign \new_[573]_  = \new_[71532]_  & \new_[71517]_ ;
  assign \new_[574]_  = \new_[71504]_  & \new_[71489]_ ;
  assign \new_[575]_  = \new_[71476]_  & \new_[71461]_ ;
  assign \new_[576]_  = \new_[71448]_  & \new_[71433]_ ;
  assign \new_[577]_  = \new_[71420]_  & \new_[71405]_ ;
  assign \new_[578]_  = \new_[71392]_  & \new_[71377]_ ;
  assign \new_[579]_  = \new_[71364]_  & \new_[71349]_ ;
  assign \new_[580]_  = \new_[71336]_  & \new_[71321]_ ;
  assign \new_[581]_  = \new_[71308]_  & \new_[71293]_ ;
  assign \new_[582]_  = \new_[71280]_  & \new_[71265]_ ;
  assign \new_[583]_  = \new_[71252]_  & \new_[71237]_ ;
  assign \new_[584]_  = \new_[71224]_  & \new_[71209]_ ;
  assign \new_[585]_  = \new_[71196]_  & \new_[71181]_ ;
  assign \new_[586]_  = \new_[71168]_  & \new_[71153]_ ;
  assign \new_[587]_  = \new_[71140]_  & \new_[71125]_ ;
  assign \new_[588]_  = \new_[71112]_  & \new_[71097]_ ;
  assign \new_[589]_  = \new_[71084]_  & \new_[71069]_ ;
  assign \new_[590]_  = \new_[71056]_  & \new_[71041]_ ;
  assign \new_[591]_  = \new_[71028]_  & \new_[71013]_ ;
  assign \new_[592]_  = \new_[71000]_  & \new_[70985]_ ;
  assign \new_[593]_  = \new_[70972]_  & \new_[70957]_ ;
  assign \new_[594]_  = \new_[70944]_  & \new_[70929]_ ;
  assign \new_[595]_  = \new_[70916]_  & \new_[70901]_ ;
  assign \new_[596]_  = \new_[70888]_  & \new_[70873]_ ;
  assign \new_[597]_  = \new_[70860]_  & \new_[70845]_ ;
  assign \new_[598]_  = \new_[70832]_  & \new_[70817]_ ;
  assign \new_[599]_  = \new_[70804]_  & \new_[70789]_ ;
  assign \new_[600]_  = \new_[70776]_  & \new_[70761]_ ;
  assign \new_[601]_  = \new_[70748]_  & \new_[70733]_ ;
  assign \new_[602]_  = \new_[70720]_  & \new_[70705]_ ;
  assign \new_[603]_  = \new_[70692]_  & \new_[70677]_ ;
  assign \new_[604]_  = \new_[70664]_  & \new_[70649]_ ;
  assign \new_[605]_  = \new_[70636]_  & \new_[70621]_ ;
  assign \new_[606]_  = \new_[70608]_  & \new_[70593]_ ;
  assign \new_[607]_  = \new_[70580]_  & \new_[70565]_ ;
  assign \new_[608]_  = \new_[70552]_  & \new_[70537]_ ;
  assign \new_[609]_  = \new_[70524]_  & \new_[70509]_ ;
  assign \new_[610]_  = \new_[70496]_  & \new_[70481]_ ;
  assign \new_[611]_  = \new_[70468]_  & \new_[70453]_ ;
  assign \new_[612]_  = \new_[70440]_  & \new_[70425]_ ;
  assign \new_[613]_  = \new_[70412]_  & \new_[70397]_ ;
  assign \new_[614]_  = \new_[70384]_  & \new_[70369]_ ;
  assign \new_[615]_  = \new_[70356]_  & \new_[70341]_ ;
  assign \new_[616]_  = \new_[70328]_  & \new_[70313]_ ;
  assign \new_[617]_  = \new_[70300]_  & \new_[70285]_ ;
  assign \new_[618]_  = \new_[70272]_  & \new_[70257]_ ;
  assign \new_[619]_  = \new_[70244]_  & \new_[70229]_ ;
  assign \new_[620]_  = \new_[70216]_  & \new_[70201]_ ;
  assign \new_[621]_  = \new_[70188]_  & \new_[70173]_ ;
  assign \new_[622]_  = \new_[70160]_  & \new_[70145]_ ;
  assign \new_[623]_  = \new_[70132]_  & \new_[70117]_ ;
  assign \new_[624]_  = \new_[70104]_  & \new_[70089]_ ;
  assign \new_[625]_  = \new_[70076]_  & \new_[70061]_ ;
  assign \new_[626]_  = \new_[70048]_  & \new_[70033]_ ;
  assign \new_[627]_  = \new_[70020]_  & \new_[70005]_ ;
  assign \new_[628]_  = \new_[69992]_  & \new_[69977]_ ;
  assign \new_[629]_  = \new_[69964]_  & \new_[69949]_ ;
  assign \new_[630]_  = \new_[69936]_  & \new_[69921]_ ;
  assign \new_[631]_  = \new_[69908]_  & \new_[69893]_ ;
  assign \new_[632]_  = \new_[69880]_  & \new_[69865]_ ;
  assign \new_[633]_  = \new_[69852]_  & \new_[69837]_ ;
  assign \new_[634]_  = \new_[69824]_  & \new_[69809]_ ;
  assign \new_[635]_  = \new_[69796]_  & \new_[69781]_ ;
  assign \new_[636]_  = \new_[69768]_  & \new_[69753]_ ;
  assign \new_[637]_  = \new_[69740]_  & \new_[69725]_ ;
  assign \new_[638]_  = \new_[69712]_  & \new_[69697]_ ;
  assign \new_[639]_  = \new_[69684]_  & \new_[69669]_ ;
  assign \new_[640]_  = \new_[69656]_  & \new_[69641]_ ;
  assign \new_[641]_  = \new_[69628]_  & \new_[69613]_ ;
  assign \new_[642]_  = \new_[69600]_  & \new_[69585]_ ;
  assign \new_[643]_  = \new_[69572]_  & \new_[69557]_ ;
  assign \new_[644]_  = \new_[69544]_  & \new_[69529]_ ;
  assign \new_[645]_  = \new_[69516]_  & \new_[69501]_ ;
  assign \new_[646]_  = \new_[69488]_  & \new_[69473]_ ;
  assign \new_[647]_  = \new_[69460]_  & \new_[69445]_ ;
  assign \new_[648]_  = \new_[69432]_  & \new_[69417]_ ;
  assign \new_[649]_  = \new_[69404]_  & \new_[69389]_ ;
  assign \new_[650]_  = \new_[69376]_  & \new_[69361]_ ;
  assign \new_[651]_  = \new_[69348]_  & \new_[69333]_ ;
  assign \new_[652]_  = \new_[69320]_  & \new_[69305]_ ;
  assign \new_[653]_  = \new_[69292]_  & \new_[69277]_ ;
  assign \new_[654]_  = \new_[69264]_  & \new_[69249]_ ;
  assign \new_[655]_  = \new_[69236]_  & \new_[69221]_ ;
  assign \new_[656]_  = \new_[69208]_  & \new_[69193]_ ;
  assign \new_[657]_  = \new_[69180]_  & \new_[69165]_ ;
  assign \new_[658]_  = \new_[69152]_  & \new_[69137]_ ;
  assign \new_[659]_  = \new_[69124]_  & \new_[69109]_ ;
  assign \new_[660]_  = \new_[69096]_  & \new_[69081]_ ;
  assign \new_[661]_  = \new_[69068]_  & \new_[69053]_ ;
  assign \new_[662]_  = \new_[69040]_  & \new_[69025]_ ;
  assign \new_[663]_  = \new_[69012]_  & \new_[68997]_ ;
  assign \new_[664]_  = \new_[68984]_  & \new_[68969]_ ;
  assign \new_[665]_  = \new_[68956]_  & \new_[68941]_ ;
  assign \new_[666]_  = \new_[68928]_  & \new_[68913]_ ;
  assign \new_[667]_  = \new_[68900]_  & \new_[68885]_ ;
  assign \new_[668]_  = \new_[68872]_  & \new_[68857]_ ;
  assign \new_[669]_  = \new_[68844]_  & \new_[68829]_ ;
  assign \new_[670]_  = \new_[68816]_  & \new_[68801]_ ;
  assign \new_[671]_  = \new_[68788]_  & \new_[68773]_ ;
  assign \new_[672]_  = \new_[68760]_  & \new_[68745]_ ;
  assign \new_[673]_  = \new_[68732]_  & \new_[68717]_ ;
  assign \new_[674]_  = \new_[68704]_  & \new_[68689]_ ;
  assign \new_[675]_  = \new_[68676]_  & \new_[68661]_ ;
  assign \new_[676]_  = \new_[68648]_  & \new_[68633]_ ;
  assign \new_[677]_  = \new_[68620]_  & \new_[68605]_ ;
  assign \new_[678]_  = \new_[68592]_  & \new_[68577]_ ;
  assign \new_[679]_  = \new_[68564]_  & \new_[68549]_ ;
  assign \new_[680]_  = \new_[68536]_  & \new_[68521]_ ;
  assign \new_[681]_  = \new_[68508]_  & \new_[68493]_ ;
  assign \new_[682]_  = \new_[68480]_  & \new_[68465]_ ;
  assign \new_[683]_  = \new_[68452]_  & \new_[68437]_ ;
  assign \new_[684]_  = \new_[68424]_  & \new_[68409]_ ;
  assign \new_[685]_  = \new_[68396]_  & \new_[68381]_ ;
  assign \new_[686]_  = \new_[68368]_  & \new_[68353]_ ;
  assign \new_[687]_  = \new_[68340]_  & \new_[68325]_ ;
  assign \new_[688]_  = \new_[68312]_  & \new_[68297]_ ;
  assign \new_[689]_  = \new_[68284]_  & \new_[68269]_ ;
  assign \new_[690]_  = \new_[68256]_  & \new_[68241]_ ;
  assign \new_[691]_  = \new_[68228]_  & \new_[68213]_ ;
  assign \new_[692]_  = \new_[68200]_  & \new_[68185]_ ;
  assign \new_[693]_  = \new_[68172]_  & \new_[68157]_ ;
  assign \new_[694]_  = \new_[68144]_  & \new_[68129]_ ;
  assign \new_[695]_  = \new_[68116]_  & \new_[68101]_ ;
  assign \new_[696]_  = \new_[68088]_  & \new_[68073]_ ;
  assign \new_[697]_  = \new_[68060]_  & \new_[68045]_ ;
  assign \new_[698]_  = \new_[68032]_  & \new_[68017]_ ;
  assign \new_[699]_  = \new_[68004]_  & \new_[67989]_ ;
  assign \new_[700]_  = \new_[67976]_  & \new_[67961]_ ;
  assign \new_[701]_  = \new_[67948]_  & \new_[67933]_ ;
  assign \new_[702]_  = \new_[67920]_  & \new_[67905]_ ;
  assign \new_[703]_  = \new_[67892]_  & \new_[67877]_ ;
  assign \new_[704]_  = \new_[67864]_  & \new_[67849]_ ;
  assign \new_[705]_  = \new_[67836]_  & \new_[67821]_ ;
  assign \new_[706]_  = \new_[67808]_  & \new_[67793]_ ;
  assign \new_[707]_  = \new_[67780]_  & \new_[67765]_ ;
  assign \new_[708]_  = \new_[67752]_  & \new_[67737]_ ;
  assign \new_[709]_  = \new_[67724]_  & \new_[67709]_ ;
  assign \new_[710]_  = \new_[67696]_  & \new_[67681]_ ;
  assign \new_[711]_  = \new_[67668]_  & \new_[67653]_ ;
  assign \new_[712]_  = \new_[67640]_  & \new_[67625]_ ;
  assign \new_[713]_  = \new_[67612]_  & \new_[67597]_ ;
  assign \new_[714]_  = \new_[67584]_  & \new_[67569]_ ;
  assign \new_[715]_  = \new_[67556]_  & \new_[67541]_ ;
  assign \new_[716]_  = \new_[67528]_  & \new_[67513]_ ;
  assign \new_[717]_  = \new_[67500]_  & \new_[67485]_ ;
  assign \new_[718]_  = \new_[67472]_  & \new_[67457]_ ;
  assign \new_[719]_  = \new_[67444]_  & \new_[67429]_ ;
  assign \new_[720]_  = \new_[67416]_  & \new_[67401]_ ;
  assign \new_[721]_  = \new_[67388]_  & \new_[67373]_ ;
  assign \new_[722]_  = \new_[67360]_  & \new_[67345]_ ;
  assign \new_[723]_  = \new_[67332]_  & \new_[67317]_ ;
  assign \new_[724]_  = \new_[67304]_  & \new_[67289]_ ;
  assign \new_[725]_  = \new_[67276]_  & \new_[67261]_ ;
  assign \new_[726]_  = \new_[67248]_  & \new_[67233]_ ;
  assign \new_[727]_  = \new_[67220]_  & \new_[67205]_ ;
  assign \new_[728]_  = \new_[67192]_  & \new_[67177]_ ;
  assign \new_[729]_  = \new_[67164]_  & \new_[67149]_ ;
  assign \new_[730]_  = \new_[67136]_  & \new_[67121]_ ;
  assign \new_[731]_  = \new_[67108]_  & \new_[67093]_ ;
  assign \new_[732]_  = \new_[67080]_  & \new_[67065]_ ;
  assign \new_[733]_  = \new_[67052]_  & \new_[67037]_ ;
  assign \new_[734]_  = \new_[67024]_  & \new_[67009]_ ;
  assign \new_[735]_  = \new_[66996]_  & \new_[66981]_ ;
  assign \new_[736]_  = \new_[66968]_  & \new_[66953]_ ;
  assign \new_[737]_  = \new_[66940]_  & \new_[66925]_ ;
  assign \new_[738]_  = \new_[66912]_  & \new_[66897]_ ;
  assign \new_[739]_  = \new_[66884]_  & \new_[66869]_ ;
  assign \new_[740]_  = \new_[66856]_  & \new_[66841]_ ;
  assign \new_[741]_  = \new_[66828]_  & \new_[66813]_ ;
  assign \new_[742]_  = \new_[66800]_  & \new_[66785]_ ;
  assign \new_[743]_  = \new_[66772]_  & \new_[66757]_ ;
  assign \new_[744]_  = \new_[66744]_  & \new_[66729]_ ;
  assign \new_[745]_  = \new_[66716]_  & \new_[66701]_ ;
  assign \new_[746]_  = \new_[66688]_  & \new_[66673]_ ;
  assign \new_[747]_  = \new_[66660]_  & \new_[66645]_ ;
  assign \new_[748]_  = \new_[66632]_  & \new_[66617]_ ;
  assign \new_[749]_  = \new_[66604]_  & \new_[66589]_ ;
  assign \new_[750]_  = \new_[66576]_  & \new_[66561]_ ;
  assign \new_[751]_  = \new_[66548]_  & \new_[66533]_ ;
  assign \new_[752]_  = \new_[66520]_  & \new_[66505]_ ;
  assign \new_[753]_  = \new_[66492]_  & \new_[66477]_ ;
  assign \new_[754]_  = \new_[66464]_  & \new_[66449]_ ;
  assign \new_[755]_  = \new_[66436]_  & \new_[66421]_ ;
  assign \new_[756]_  = \new_[66408]_  & \new_[66393]_ ;
  assign \new_[757]_  = \new_[66380]_  & \new_[66365]_ ;
  assign \new_[758]_  = \new_[66352]_  & \new_[66337]_ ;
  assign \new_[759]_  = \new_[66324]_  & \new_[66309]_ ;
  assign \new_[760]_  = \new_[66296]_  & \new_[66281]_ ;
  assign \new_[761]_  = \new_[66268]_  & \new_[66253]_ ;
  assign \new_[762]_  = \new_[66240]_  & \new_[66225]_ ;
  assign \new_[763]_  = \new_[66212]_  & \new_[66197]_ ;
  assign \new_[764]_  = \new_[66184]_  & \new_[66169]_ ;
  assign \new_[765]_  = \new_[66156]_  & \new_[66141]_ ;
  assign \new_[766]_  = \new_[66128]_  & \new_[66113]_ ;
  assign \new_[767]_  = \new_[66100]_  & \new_[66085]_ ;
  assign \new_[768]_  = \new_[66072]_  & \new_[66057]_ ;
  assign \new_[769]_  = \new_[66044]_  & \new_[66029]_ ;
  assign \new_[770]_  = \new_[66016]_  & \new_[66001]_ ;
  assign \new_[771]_  = \new_[65988]_  & \new_[65973]_ ;
  assign \new_[772]_  = \new_[65960]_  & \new_[65945]_ ;
  assign \new_[773]_  = \new_[65932]_  & \new_[65917]_ ;
  assign \new_[774]_  = \new_[65904]_  & \new_[65889]_ ;
  assign \new_[775]_  = \new_[65876]_  & \new_[65861]_ ;
  assign \new_[776]_  = \new_[65848]_  & \new_[65833]_ ;
  assign \new_[777]_  = \new_[65820]_  & \new_[65805]_ ;
  assign \new_[778]_  = \new_[65792]_  & \new_[65777]_ ;
  assign \new_[779]_  = \new_[65764]_  & \new_[65749]_ ;
  assign \new_[780]_  = \new_[65736]_  & \new_[65721]_ ;
  assign \new_[781]_  = \new_[65708]_  & \new_[65693]_ ;
  assign \new_[782]_  = \new_[65680]_  & \new_[65665]_ ;
  assign \new_[783]_  = \new_[65652]_  & \new_[65637]_ ;
  assign \new_[784]_  = \new_[65624]_  & \new_[65609]_ ;
  assign \new_[785]_  = \new_[65596]_  & \new_[65581]_ ;
  assign \new_[786]_  = \new_[65568]_  & \new_[65553]_ ;
  assign \new_[787]_  = \new_[65540]_  & \new_[65525]_ ;
  assign \new_[788]_  = \new_[65512]_  & \new_[65497]_ ;
  assign \new_[789]_  = \new_[65484]_  & \new_[65469]_ ;
  assign \new_[790]_  = \new_[65456]_  & \new_[65441]_ ;
  assign \new_[791]_  = \new_[65428]_  & \new_[65413]_ ;
  assign \new_[792]_  = \new_[65400]_  & \new_[65385]_ ;
  assign \new_[793]_  = \new_[65372]_  & \new_[65357]_ ;
  assign \new_[794]_  = \new_[65344]_  & \new_[65329]_ ;
  assign \new_[795]_  = \new_[65316]_  & \new_[65301]_ ;
  assign \new_[796]_  = \new_[65288]_  & \new_[65273]_ ;
  assign \new_[797]_  = \new_[65260]_  & \new_[65245]_ ;
  assign \new_[798]_  = \new_[65232]_  & \new_[65217]_ ;
  assign \new_[799]_  = \new_[65204]_  & \new_[65189]_ ;
  assign \new_[800]_  = \new_[65176]_  & \new_[65161]_ ;
  assign \new_[801]_  = \new_[65148]_  & \new_[65133]_ ;
  assign \new_[802]_  = \new_[65120]_  & \new_[65105]_ ;
  assign \new_[803]_  = \new_[65092]_  & \new_[65077]_ ;
  assign \new_[804]_  = \new_[65064]_  & \new_[65049]_ ;
  assign \new_[805]_  = \new_[65036]_  & \new_[65021]_ ;
  assign \new_[806]_  = \new_[65008]_  & \new_[64993]_ ;
  assign \new_[807]_  = \new_[64980]_  & \new_[64965]_ ;
  assign \new_[808]_  = \new_[64952]_  & \new_[64937]_ ;
  assign \new_[809]_  = \new_[64924]_  & \new_[64909]_ ;
  assign \new_[810]_  = \new_[64896]_  & \new_[64881]_ ;
  assign \new_[811]_  = \new_[64868]_  & \new_[64853]_ ;
  assign \new_[812]_  = \new_[64840]_  & \new_[64825]_ ;
  assign \new_[813]_  = \new_[64812]_  & \new_[64797]_ ;
  assign \new_[814]_  = \new_[64784]_  & \new_[64769]_ ;
  assign \new_[815]_  = \new_[64756]_  & \new_[64741]_ ;
  assign \new_[816]_  = \new_[64728]_  & \new_[64713]_ ;
  assign \new_[817]_  = \new_[64700]_  & \new_[64685]_ ;
  assign \new_[818]_  = \new_[64672]_  & \new_[64657]_ ;
  assign \new_[819]_  = \new_[64644]_  & \new_[64629]_ ;
  assign \new_[820]_  = \new_[64616]_  & \new_[64601]_ ;
  assign \new_[821]_  = \new_[64588]_  & \new_[64573]_ ;
  assign \new_[822]_  = \new_[64560]_  & \new_[64545]_ ;
  assign \new_[823]_  = \new_[64532]_  & \new_[64517]_ ;
  assign \new_[824]_  = \new_[64504]_  & \new_[64489]_ ;
  assign \new_[825]_  = \new_[64476]_  & \new_[64461]_ ;
  assign \new_[826]_  = \new_[64448]_  & \new_[64433]_ ;
  assign \new_[827]_  = \new_[64420]_  & \new_[64405]_ ;
  assign \new_[828]_  = \new_[64392]_  & \new_[64377]_ ;
  assign \new_[829]_  = \new_[64364]_  & \new_[64349]_ ;
  assign \new_[830]_  = \new_[64336]_  & \new_[64321]_ ;
  assign \new_[831]_  = \new_[64308]_  & \new_[64293]_ ;
  assign \new_[832]_  = \new_[64280]_  & \new_[64265]_ ;
  assign \new_[833]_  = \new_[64252]_  & \new_[64237]_ ;
  assign \new_[834]_  = \new_[64224]_  & \new_[64209]_ ;
  assign \new_[835]_  = \new_[64196]_  & \new_[64181]_ ;
  assign \new_[836]_  = \new_[64168]_  & \new_[64153]_ ;
  assign \new_[837]_  = \new_[64140]_  & \new_[64125]_ ;
  assign \new_[838]_  = \new_[64112]_  & \new_[64097]_ ;
  assign \new_[839]_  = \new_[64084]_  & \new_[64069]_ ;
  assign \new_[840]_  = \new_[64056]_  & \new_[64041]_ ;
  assign \new_[841]_  = \new_[64028]_  & \new_[64013]_ ;
  assign \new_[842]_  = \new_[64000]_  & \new_[63985]_ ;
  assign \new_[843]_  = \new_[63972]_  & \new_[63957]_ ;
  assign \new_[844]_  = \new_[63944]_  & \new_[63929]_ ;
  assign \new_[845]_  = \new_[63916]_  & \new_[63901]_ ;
  assign \new_[846]_  = \new_[63888]_  & \new_[63873]_ ;
  assign \new_[847]_  = \new_[63860]_  & \new_[63845]_ ;
  assign \new_[848]_  = \new_[63832]_  & \new_[63817]_ ;
  assign \new_[849]_  = \new_[63804]_  & \new_[63789]_ ;
  assign \new_[850]_  = \new_[63776]_  & \new_[63761]_ ;
  assign \new_[851]_  = \new_[63748]_  & \new_[63733]_ ;
  assign \new_[852]_  = \new_[63720]_  & \new_[63705]_ ;
  assign \new_[853]_  = \new_[63692]_  & \new_[63677]_ ;
  assign \new_[854]_  = \new_[63664]_  & \new_[63649]_ ;
  assign \new_[855]_  = \new_[63636]_  & \new_[63621]_ ;
  assign \new_[856]_  = \new_[63608]_  & \new_[63593]_ ;
  assign \new_[857]_  = \new_[63580]_  & \new_[63565]_ ;
  assign \new_[858]_  = \new_[63552]_  & \new_[63537]_ ;
  assign \new_[859]_  = \new_[63524]_  & \new_[63509]_ ;
  assign \new_[860]_  = \new_[63496]_  & \new_[63481]_ ;
  assign \new_[861]_  = \new_[63468]_  & \new_[63453]_ ;
  assign \new_[862]_  = \new_[63440]_  & \new_[63425]_ ;
  assign \new_[863]_  = \new_[63412]_  & \new_[63397]_ ;
  assign \new_[864]_  = \new_[63384]_  & \new_[63369]_ ;
  assign \new_[865]_  = \new_[63356]_  & \new_[63341]_ ;
  assign \new_[866]_  = \new_[63328]_  & \new_[63313]_ ;
  assign \new_[867]_  = \new_[63300]_  & \new_[63285]_ ;
  assign \new_[868]_  = \new_[63272]_  & \new_[63257]_ ;
  assign \new_[869]_  = \new_[63244]_  & \new_[63229]_ ;
  assign \new_[870]_  = \new_[63216]_  & \new_[63201]_ ;
  assign \new_[871]_  = \new_[63188]_  & \new_[63173]_ ;
  assign \new_[872]_  = \new_[63160]_  & \new_[63145]_ ;
  assign \new_[873]_  = \new_[63132]_  & \new_[63117]_ ;
  assign \new_[874]_  = \new_[63104]_  & \new_[63089]_ ;
  assign \new_[875]_  = \new_[63076]_  & \new_[63061]_ ;
  assign \new_[876]_  = \new_[63048]_  & \new_[63033]_ ;
  assign \new_[877]_  = \new_[63020]_  & \new_[63005]_ ;
  assign \new_[878]_  = \new_[62992]_  & \new_[62977]_ ;
  assign \new_[879]_  = \new_[62964]_  & \new_[62949]_ ;
  assign \new_[880]_  = \new_[62936]_  & \new_[62921]_ ;
  assign \new_[881]_  = \new_[62908]_  & \new_[62893]_ ;
  assign \new_[882]_  = \new_[62880]_  & \new_[62865]_ ;
  assign \new_[883]_  = \new_[62852]_  & \new_[62837]_ ;
  assign \new_[884]_  = \new_[62824]_  & \new_[62809]_ ;
  assign \new_[885]_  = \new_[62796]_  & \new_[62781]_ ;
  assign \new_[886]_  = \new_[62768]_  & \new_[62753]_ ;
  assign \new_[887]_  = \new_[62740]_  & \new_[62725]_ ;
  assign \new_[888]_  = \new_[62712]_  & \new_[62697]_ ;
  assign \new_[889]_  = \new_[62684]_  & \new_[62669]_ ;
  assign \new_[890]_  = \new_[62656]_  & \new_[62641]_ ;
  assign \new_[891]_  = \new_[62628]_  & \new_[62613]_ ;
  assign \new_[892]_  = \new_[62600]_  & \new_[62585]_ ;
  assign \new_[893]_  = \new_[62572]_  & \new_[62557]_ ;
  assign \new_[894]_  = \new_[62544]_  & \new_[62529]_ ;
  assign \new_[895]_  = \new_[62516]_  & \new_[62501]_ ;
  assign \new_[896]_  = \new_[62488]_  & \new_[62473]_ ;
  assign \new_[897]_  = \new_[62460]_  & \new_[62445]_ ;
  assign \new_[898]_  = \new_[62432]_  & \new_[62417]_ ;
  assign \new_[899]_  = \new_[62404]_  & \new_[62389]_ ;
  assign \new_[900]_  = \new_[62376]_  & \new_[62361]_ ;
  assign \new_[901]_  = \new_[62348]_  & \new_[62333]_ ;
  assign \new_[902]_  = \new_[62320]_  & \new_[62305]_ ;
  assign \new_[903]_  = \new_[62292]_  & \new_[62277]_ ;
  assign \new_[904]_  = \new_[62264]_  & \new_[62249]_ ;
  assign \new_[905]_  = \new_[62236]_  & \new_[62221]_ ;
  assign \new_[906]_  = \new_[62208]_  & \new_[62193]_ ;
  assign \new_[907]_  = \new_[62180]_  & \new_[62165]_ ;
  assign \new_[908]_  = \new_[62152]_  & \new_[62137]_ ;
  assign \new_[909]_  = \new_[62124]_  & \new_[62109]_ ;
  assign \new_[910]_  = \new_[62096]_  & \new_[62081]_ ;
  assign \new_[911]_  = \new_[62068]_  & \new_[62053]_ ;
  assign \new_[912]_  = \new_[62040]_  & \new_[62025]_ ;
  assign \new_[913]_  = \new_[62012]_  & \new_[61997]_ ;
  assign \new_[914]_  = \new_[61984]_  & \new_[61969]_ ;
  assign \new_[915]_  = \new_[61956]_  & \new_[61941]_ ;
  assign \new_[916]_  = \new_[61928]_  & \new_[61913]_ ;
  assign \new_[917]_  = \new_[61900]_  & \new_[61885]_ ;
  assign \new_[918]_  = \new_[61872]_  & \new_[61857]_ ;
  assign \new_[919]_  = \new_[61844]_  & \new_[61829]_ ;
  assign \new_[920]_  = \new_[61816]_  & \new_[61801]_ ;
  assign \new_[921]_  = \new_[61788]_  & \new_[61773]_ ;
  assign \new_[922]_  = \new_[61760]_  & \new_[61745]_ ;
  assign \new_[923]_  = \new_[61732]_  & \new_[61717]_ ;
  assign \new_[924]_  = \new_[61704]_  & \new_[61689]_ ;
  assign \new_[925]_  = \new_[61676]_  & \new_[61661]_ ;
  assign \new_[926]_  = \new_[61648]_  & \new_[61633]_ ;
  assign \new_[927]_  = \new_[61620]_  & \new_[61605]_ ;
  assign \new_[928]_  = \new_[61592]_  & \new_[61577]_ ;
  assign \new_[929]_  = \new_[61564]_  & \new_[61549]_ ;
  assign \new_[930]_  = \new_[61536]_  & \new_[61521]_ ;
  assign \new_[931]_  = \new_[61508]_  & \new_[61493]_ ;
  assign \new_[932]_  = \new_[61480]_  & \new_[61465]_ ;
  assign \new_[933]_  = \new_[61452]_  & \new_[61437]_ ;
  assign \new_[934]_  = \new_[61424]_  & \new_[61409]_ ;
  assign \new_[935]_  = \new_[61396]_  & \new_[61381]_ ;
  assign \new_[936]_  = \new_[61368]_  & \new_[61353]_ ;
  assign \new_[937]_  = \new_[61340]_  & \new_[61325]_ ;
  assign \new_[938]_  = \new_[61312]_  & \new_[61297]_ ;
  assign \new_[939]_  = \new_[61284]_  & \new_[61269]_ ;
  assign \new_[940]_  = \new_[61256]_  & \new_[61241]_ ;
  assign \new_[941]_  = \new_[61228]_  & \new_[61213]_ ;
  assign \new_[942]_  = \new_[61200]_  & \new_[61185]_ ;
  assign \new_[943]_  = \new_[61172]_  & \new_[61157]_ ;
  assign \new_[944]_  = \new_[61144]_  & \new_[61129]_ ;
  assign \new_[945]_  = \new_[61116]_  & \new_[61101]_ ;
  assign \new_[946]_  = \new_[61088]_  & \new_[61073]_ ;
  assign \new_[947]_  = \new_[61060]_  & \new_[61045]_ ;
  assign \new_[948]_  = \new_[61032]_  & \new_[61017]_ ;
  assign \new_[949]_  = \new_[61004]_  & \new_[60989]_ ;
  assign \new_[950]_  = \new_[60976]_  & \new_[60961]_ ;
  assign \new_[951]_  = \new_[60948]_  & \new_[60933]_ ;
  assign \new_[952]_  = \new_[60920]_  & \new_[60905]_ ;
  assign \new_[953]_  = \new_[60892]_  & \new_[60877]_ ;
  assign \new_[954]_  = \new_[60864]_  & \new_[60849]_ ;
  assign \new_[955]_  = \new_[60836]_  & \new_[60821]_ ;
  assign \new_[956]_  = \new_[60808]_  & \new_[60793]_ ;
  assign \new_[957]_  = \new_[60780]_  & \new_[60765]_ ;
  assign \new_[958]_  = \new_[60752]_  & \new_[60737]_ ;
  assign \new_[959]_  = \new_[60724]_  & \new_[60709]_ ;
  assign \new_[960]_  = \new_[60696]_  & \new_[60681]_ ;
  assign \new_[961]_  = \new_[60668]_  & \new_[60653]_ ;
  assign \new_[962]_  = \new_[60640]_  & \new_[60625]_ ;
  assign \new_[963]_  = \new_[60612]_  & \new_[60597]_ ;
  assign \new_[964]_  = \new_[60584]_  & \new_[60569]_ ;
  assign \new_[965]_  = \new_[60556]_  & \new_[60541]_ ;
  assign \new_[966]_  = \new_[60528]_  & \new_[60513]_ ;
  assign \new_[967]_  = \new_[60500]_  & \new_[60485]_ ;
  assign \new_[968]_  = \new_[60472]_  & \new_[60457]_ ;
  assign \new_[969]_  = \new_[60444]_  & \new_[60429]_ ;
  assign \new_[970]_  = \new_[60416]_  & \new_[60401]_ ;
  assign \new_[971]_  = \new_[60388]_  & \new_[60373]_ ;
  assign \new_[972]_  = \new_[60360]_  & \new_[60345]_ ;
  assign \new_[973]_  = \new_[60332]_  & \new_[60317]_ ;
  assign \new_[974]_  = \new_[60304]_  & \new_[60289]_ ;
  assign \new_[975]_  = \new_[60276]_  & \new_[60263]_ ;
  assign \new_[976]_  = \new_[60250]_  & \new_[60237]_ ;
  assign \new_[977]_  = \new_[60224]_  & \new_[60211]_ ;
  assign \new_[978]_  = \new_[60198]_  & \new_[60185]_ ;
  assign \new_[979]_  = \new_[60172]_  & \new_[60159]_ ;
  assign \new_[980]_  = \new_[60146]_  & \new_[60133]_ ;
  assign \new_[981]_  = \new_[60120]_  & \new_[60107]_ ;
  assign \new_[982]_  = \new_[60094]_  & \new_[60081]_ ;
  assign \new_[983]_  = \new_[60068]_  & \new_[60055]_ ;
  assign \new_[984]_  = \new_[60042]_  & \new_[60029]_ ;
  assign \new_[985]_  = \new_[60016]_  & \new_[60003]_ ;
  assign \new_[986]_  = \new_[59990]_  & \new_[59977]_ ;
  assign \new_[987]_  = \new_[59964]_  & \new_[59951]_ ;
  assign \new_[988]_  = \new_[59938]_  & \new_[59925]_ ;
  assign \new_[989]_  = \new_[59912]_  & \new_[59899]_ ;
  assign \new_[990]_  = \new_[59886]_  & \new_[59873]_ ;
  assign \new_[991]_  = \new_[59860]_  & \new_[59847]_ ;
  assign \new_[992]_  = \new_[59834]_  & \new_[59821]_ ;
  assign \new_[993]_  = \new_[59808]_  & \new_[59795]_ ;
  assign \new_[994]_  = \new_[59782]_  & \new_[59769]_ ;
  assign \new_[995]_  = \new_[59756]_  & \new_[59743]_ ;
  assign \new_[996]_  = \new_[59730]_  & \new_[59717]_ ;
  assign \new_[997]_  = \new_[59704]_  & \new_[59691]_ ;
  assign \new_[998]_  = \new_[59678]_  & \new_[59665]_ ;
  assign \new_[999]_  = \new_[59652]_  & \new_[59639]_ ;
  assign \new_[1000]_  = \new_[59626]_  & \new_[59613]_ ;
  assign \new_[1001]_  = \new_[59600]_  & \new_[59587]_ ;
  assign \new_[1002]_  = \new_[59574]_  & \new_[59561]_ ;
  assign \new_[1003]_  = \new_[59548]_  & \new_[59535]_ ;
  assign \new_[1004]_  = \new_[59522]_  & \new_[59509]_ ;
  assign \new_[1005]_  = \new_[59496]_  & \new_[59483]_ ;
  assign \new_[1006]_  = \new_[59470]_  & \new_[59457]_ ;
  assign \new_[1007]_  = \new_[59444]_  & \new_[59431]_ ;
  assign \new_[1008]_  = \new_[59418]_  & \new_[59405]_ ;
  assign \new_[1009]_  = \new_[59392]_  & \new_[59379]_ ;
  assign \new_[1010]_  = \new_[59366]_  & \new_[59353]_ ;
  assign \new_[1011]_  = \new_[59340]_  & \new_[59327]_ ;
  assign \new_[1012]_  = \new_[59314]_  & \new_[59301]_ ;
  assign \new_[1013]_  = \new_[59288]_  & \new_[59275]_ ;
  assign \new_[1014]_  = \new_[59262]_  & \new_[59249]_ ;
  assign \new_[1015]_  = \new_[59236]_  & \new_[59223]_ ;
  assign \new_[1016]_  = \new_[59210]_  & \new_[59197]_ ;
  assign \new_[1017]_  = \new_[59184]_  & \new_[59171]_ ;
  assign \new_[1018]_  = \new_[59158]_  & \new_[59145]_ ;
  assign \new_[1019]_  = \new_[59132]_  & \new_[59119]_ ;
  assign \new_[1020]_  = \new_[59106]_  & \new_[59093]_ ;
  assign \new_[1021]_  = \new_[59080]_  & \new_[59067]_ ;
  assign \new_[1022]_  = \new_[59054]_  & \new_[59041]_ ;
  assign \new_[1023]_  = \new_[59028]_  & \new_[59015]_ ;
  assign \new_[1024]_  = \new_[59002]_  & \new_[58989]_ ;
  assign \new_[1025]_  = \new_[58976]_  & \new_[58963]_ ;
  assign \new_[1026]_  = \new_[58950]_  & \new_[58937]_ ;
  assign \new_[1027]_  = \new_[58924]_  & \new_[58911]_ ;
  assign \new_[1028]_  = \new_[58898]_  & \new_[58885]_ ;
  assign \new_[1029]_  = \new_[58872]_  & \new_[58859]_ ;
  assign \new_[1030]_  = \new_[58846]_  & \new_[58833]_ ;
  assign \new_[1031]_  = \new_[58820]_  & \new_[58807]_ ;
  assign \new_[1032]_  = \new_[58794]_  & \new_[58781]_ ;
  assign \new_[1033]_  = \new_[58768]_  & \new_[58755]_ ;
  assign \new_[1034]_  = \new_[58742]_  & \new_[58729]_ ;
  assign \new_[1035]_  = \new_[58716]_  & \new_[58703]_ ;
  assign \new_[1036]_  = \new_[58690]_  & \new_[58677]_ ;
  assign \new_[1037]_  = \new_[58664]_  & \new_[58651]_ ;
  assign \new_[1038]_  = \new_[58638]_  & \new_[58625]_ ;
  assign \new_[1039]_  = \new_[58612]_  & \new_[58599]_ ;
  assign \new_[1040]_  = \new_[58586]_  & \new_[58573]_ ;
  assign \new_[1041]_  = \new_[58560]_  & \new_[58547]_ ;
  assign \new_[1042]_  = \new_[58534]_  & \new_[58521]_ ;
  assign \new_[1043]_  = \new_[58508]_  & \new_[58495]_ ;
  assign \new_[1044]_  = \new_[58482]_  & \new_[58469]_ ;
  assign \new_[1045]_  = \new_[58456]_  & \new_[58443]_ ;
  assign \new_[1046]_  = \new_[58430]_  & \new_[58417]_ ;
  assign \new_[1047]_  = \new_[58404]_  & \new_[58391]_ ;
  assign \new_[1048]_  = \new_[58378]_  & \new_[58365]_ ;
  assign \new_[1049]_  = \new_[58352]_  & \new_[58339]_ ;
  assign \new_[1050]_  = \new_[58326]_  & \new_[58313]_ ;
  assign \new_[1051]_  = \new_[58300]_  & \new_[58287]_ ;
  assign \new_[1052]_  = \new_[58274]_  & \new_[58261]_ ;
  assign \new_[1053]_  = \new_[58248]_  & \new_[58235]_ ;
  assign \new_[1054]_  = \new_[58222]_  & \new_[58209]_ ;
  assign \new_[1055]_  = \new_[58196]_  & \new_[58183]_ ;
  assign \new_[1056]_  = \new_[58170]_  & \new_[58157]_ ;
  assign \new_[1057]_  = \new_[58144]_  & \new_[58131]_ ;
  assign \new_[1058]_  = \new_[58118]_  & \new_[58105]_ ;
  assign \new_[1059]_  = \new_[58092]_  & \new_[58079]_ ;
  assign \new_[1060]_  = \new_[58066]_  & \new_[58053]_ ;
  assign \new_[1061]_  = \new_[58040]_  & \new_[58027]_ ;
  assign \new_[1062]_  = \new_[58014]_  & \new_[58001]_ ;
  assign \new_[1063]_  = \new_[57988]_  & \new_[57975]_ ;
  assign \new_[1064]_  = \new_[57962]_  & \new_[57949]_ ;
  assign \new_[1065]_  = \new_[57936]_  & \new_[57923]_ ;
  assign \new_[1066]_  = \new_[57910]_  & \new_[57897]_ ;
  assign \new_[1067]_  = \new_[57884]_  & \new_[57871]_ ;
  assign \new_[1068]_  = \new_[57858]_  & \new_[57845]_ ;
  assign \new_[1069]_  = \new_[57832]_  & \new_[57819]_ ;
  assign \new_[1070]_  = \new_[57806]_  & \new_[57793]_ ;
  assign \new_[1071]_  = \new_[57780]_  & \new_[57767]_ ;
  assign \new_[1072]_  = \new_[57754]_  & \new_[57741]_ ;
  assign \new_[1073]_  = \new_[57728]_  & \new_[57715]_ ;
  assign \new_[1074]_  = \new_[57702]_  & \new_[57689]_ ;
  assign \new_[1075]_  = \new_[57676]_  & \new_[57663]_ ;
  assign \new_[1076]_  = \new_[57650]_  & \new_[57637]_ ;
  assign \new_[1077]_  = \new_[57624]_  & \new_[57611]_ ;
  assign \new_[1078]_  = \new_[57598]_  & \new_[57585]_ ;
  assign \new_[1079]_  = \new_[57572]_  & \new_[57559]_ ;
  assign \new_[1080]_  = \new_[57546]_  & \new_[57533]_ ;
  assign \new_[1081]_  = \new_[57520]_  & \new_[57507]_ ;
  assign \new_[1082]_  = \new_[57494]_  & \new_[57481]_ ;
  assign \new_[1083]_  = \new_[57468]_  & \new_[57455]_ ;
  assign \new_[1084]_  = \new_[57442]_  & \new_[57429]_ ;
  assign \new_[1085]_  = \new_[57416]_  & \new_[57403]_ ;
  assign \new_[1086]_  = \new_[57390]_  & \new_[57377]_ ;
  assign \new_[1087]_  = \new_[57364]_  & \new_[57351]_ ;
  assign \new_[1088]_  = \new_[57338]_  & \new_[57325]_ ;
  assign \new_[1089]_  = \new_[57312]_  & \new_[57299]_ ;
  assign \new_[1090]_  = \new_[57286]_  & \new_[57273]_ ;
  assign \new_[1091]_  = \new_[57260]_  & \new_[57247]_ ;
  assign \new_[1092]_  = \new_[57234]_  & \new_[57221]_ ;
  assign \new_[1093]_  = \new_[57208]_  & \new_[57195]_ ;
  assign \new_[1094]_  = \new_[57182]_  & \new_[57169]_ ;
  assign \new_[1095]_  = \new_[57156]_  & \new_[57143]_ ;
  assign \new_[1096]_  = \new_[57130]_  & \new_[57117]_ ;
  assign \new_[1097]_  = \new_[57104]_  & \new_[57091]_ ;
  assign \new_[1098]_  = \new_[57078]_  & \new_[57065]_ ;
  assign \new_[1099]_  = \new_[57052]_  & \new_[57039]_ ;
  assign \new_[1100]_  = \new_[57026]_  & \new_[57013]_ ;
  assign \new_[1101]_  = \new_[57000]_  & \new_[56987]_ ;
  assign \new_[1102]_  = \new_[56974]_  & \new_[56961]_ ;
  assign \new_[1103]_  = \new_[56948]_  & \new_[56935]_ ;
  assign \new_[1104]_  = \new_[56922]_  & \new_[56909]_ ;
  assign \new_[1105]_  = \new_[56896]_  & \new_[56883]_ ;
  assign \new_[1106]_  = \new_[56870]_  & \new_[56857]_ ;
  assign \new_[1107]_  = \new_[56844]_  & \new_[56831]_ ;
  assign \new_[1108]_  = \new_[56818]_  & \new_[56805]_ ;
  assign \new_[1109]_  = \new_[56792]_  & \new_[56779]_ ;
  assign \new_[1110]_  = \new_[56766]_  & \new_[56753]_ ;
  assign \new_[1111]_  = \new_[56740]_  & \new_[56727]_ ;
  assign \new_[1112]_  = \new_[56714]_  & \new_[56701]_ ;
  assign \new_[1113]_  = \new_[56688]_  & \new_[56675]_ ;
  assign \new_[1114]_  = \new_[56662]_  & \new_[56649]_ ;
  assign \new_[1115]_  = \new_[56636]_  & \new_[56623]_ ;
  assign \new_[1116]_  = \new_[56610]_  & \new_[56597]_ ;
  assign \new_[1117]_  = \new_[56584]_  & \new_[56571]_ ;
  assign \new_[1118]_  = \new_[56558]_  & \new_[56545]_ ;
  assign \new_[1119]_  = \new_[56532]_  & \new_[56519]_ ;
  assign \new_[1120]_  = \new_[56506]_  & \new_[56493]_ ;
  assign \new_[1121]_  = \new_[56480]_  & \new_[56467]_ ;
  assign \new_[1122]_  = \new_[56454]_  & \new_[56441]_ ;
  assign \new_[1123]_  = \new_[56428]_  & \new_[56415]_ ;
  assign \new_[1124]_  = \new_[56402]_  & \new_[56389]_ ;
  assign \new_[1125]_  = \new_[56376]_  & \new_[56363]_ ;
  assign \new_[1126]_  = \new_[56350]_  & \new_[56337]_ ;
  assign \new_[1127]_  = \new_[56324]_  & \new_[56311]_ ;
  assign \new_[1128]_  = \new_[56298]_  & \new_[56285]_ ;
  assign \new_[1129]_  = \new_[56272]_  & \new_[56259]_ ;
  assign \new_[1130]_  = \new_[56246]_  & \new_[56233]_ ;
  assign \new_[1131]_  = \new_[56220]_  & \new_[56207]_ ;
  assign \new_[1132]_  = \new_[56194]_  & \new_[56181]_ ;
  assign \new_[1133]_  = \new_[56168]_  & \new_[56155]_ ;
  assign \new_[1134]_  = \new_[56142]_  & \new_[56129]_ ;
  assign \new_[1135]_  = \new_[56116]_  & \new_[56103]_ ;
  assign \new_[1136]_  = \new_[56090]_  & \new_[56077]_ ;
  assign \new_[1137]_  = \new_[56064]_  & \new_[56051]_ ;
  assign \new_[1138]_  = \new_[56038]_  & \new_[56025]_ ;
  assign \new_[1139]_  = \new_[56012]_  & \new_[55999]_ ;
  assign \new_[1140]_  = \new_[55986]_  & \new_[55973]_ ;
  assign \new_[1141]_  = \new_[55960]_  & \new_[55947]_ ;
  assign \new_[1142]_  = \new_[55934]_  & \new_[55921]_ ;
  assign \new_[1143]_  = \new_[55908]_  & \new_[55895]_ ;
  assign \new_[1144]_  = \new_[55882]_  & \new_[55869]_ ;
  assign \new_[1145]_  = \new_[55856]_  & \new_[55843]_ ;
  assign \new_[1146]_  = \new_[55830]_  & \new_[55817]_ ;
  assign \new_[1147]_  = \new_[55804]_  & \new_[55791]_ ;
  assign \new_[1148]_  = \new_[55778]_  & \new_[55765]_ ;
  assign \new_[1149]_  = \new_[55752]_  & \new_[55739]_ ;
  assign \new_[1150]_  = \new_[55726]_  & \new_[55713]_ ;
  assign \new_[1151]_  = \new_[55700]_  & \new_[55687]_ ;
  assign \new_[1152]_  = \new_[55674]_  & \new_[55661]_ ;
  assign \new_[1153]_  = \new_[55648]_  & \new_[55635]_ ;
  assign \new_[1154]_  = \new_[55622]_  & \new_[55609]_ ;
  assign \new_[1155]_  = \new_[55596]_  & \new_[55583]_ ;
  assign \new_[1156]_  = \new_[55570]_  & \new_[55557]_ ;
  assign \new_[1157]_  = \new_[55544]_  & \new_[55531]_ ;
  assign \new_[1158]_  = \new_[55518]_  & \new_[55505]_ ;
  assign \new_[1159]_  = \new_[55492]_  & \new_[55479]_ ;
  assign \new_[1160]_  = \new_[55466]_  & \new_[55453]_ ;
  assign \new_[1161]_  = \new_[55440]_  & \new_[55427]_ ;
  assign \new_[1162]_  = \new_[55414]_  & \new_[55401]_ ;
  assign \new_[1163]_  = \new_[55388]_  & \new_[55375]_ ;
  assign \new_[1164]_  = \new_[55362]_  & \new_[55349]_ ;
  assign \new_[1165]_  = \new_[55336]_  & \new_[55323]_ ;
  assign \new_[1166]_  = \new_[55310]_  & \new_[55297]_ ;
  assign \new_[1167]_  = \new_[55284]_  & \new_[55271]_ ;
  assign \new_[1168]_  = \new_[55258]_  & \new_[55245]_ ;
  assign \new_[1169]_  = \new_[55232]_  & \new_[55219]_ ;
  assign \new_[1170]_  = \new_[55206]_  & \new_[55193]_ ;
  assign \new_[1171]_  = \new_[55180]_  & \new_[55167]_ ;
  assign \new_[1172]_  = \new_[55154]_  & \new_[55141]_ ;
  assign \new_[1173]_  = \new_[55128]_  & \new_[55115]_ ;
  assign \new_[1174]_  = \new_[55102]_  & \new_[55089]_ ;
  assign \new_[1175]_  = \new_[55076]_  & \new_[55063]_ ;
  assign \new_[1176]_  = \new_[55050]_  & \new_[55037]_ ;
  assign \new_[1177]_  = \new_[55024]_  & \new_[55011]_ ;
  assign \new_[1178]_  = \new_[54998]_  & \new_[54985]_ ;
  assign \new_[1179]_  = \new_[54972]_  & \new_[54959]_ ;
  assign \new_[1180]_  = \new_[54946]_  & \new_[54933]_ ;
  assign \new_[1181]_  = \new_[54920]_  & \new_[54907]_ ;
  assign \new_[1182]_  = \new_[54894]_  & \new_[54881]_ ;
  assign \new_[1183]_  = \new_[54868]_  & \new_[54855]_ ;
  assign \new_[1184]_  = \new_[54842]_  & \new_[54829]_ ;
  assign \new_[1185]_  = \new_[54816]_  & \new_[54803]_ ;
  assign \new_[1186]_  = \new_[54790]_  & \new_[54777]_ ;
  assign \new_[1187]_  = \new_[54764]_  & \new_[54751]_ ;
  assign \new_[1188]_  = \new_[54738]_  & \new_[54725]_ ;
  assign \new_[1189]_  = \new_[54712]_  & \new_[54699]_ ;
  assign \new_[1190]_  = \new_[54686]_  & \new_[54673]_ ;
  assign \new_[1191]_  = \new_[54660]_  & \new_[54647]_ ;
  assign \new_[1192]_  = \new_[54634]_  & \new_[54621]_ ;
  assign \new_[1193]_  = \new_[54608]_  & \new_[54595]_ ;
  assign \new_[1194]_  = \new_[54582]_  & \new_[54569]_ ;
  assign \new_[1195]_  = \new_[54556]_  & \new_[54543]_ ;
  assign \new_[1196]_  = \new_[54530]_  & \new_[54517]_ ;
  assign \new_[1197]_  = \new_[54504]_  & \new_[54491]_ ;
  assign \new_[1198]_  = \new_[54478]_  & \new_[54465]_ ;
  assign \new_[1199]_  = \new_[54452]_  & \new_[54439]_ ;
  assign \new_[1200]_  = \new_[54426]_  & \new_[54413]_ ;
  assign \new_[1201]_  = \new_[54400]_  & \new_[54387]_ ;
  assign \new_[1202]_  = \new_[54374]_  & \new_[54361]_ ;
  assign \new_[1203]_  = \new_[54348]_  & \new_[54335]_ ;
  assign \new_[1204]_  = \new_[54322]_  & \new_[54309]_ ;
  assign \new_[1205]_  = \new_[54296]_  & \new_[54283]_ ;
  assign \new_[1206]_  = \new_[54270]_  & \new_[54257]_ ;
  assign \new_[1207]_  = \new_[54244]_  & \new_[54231]_ ;
  assign \new_[1208]_  = \new_[54218]_  & \new_[54205]_ ;
  assign \new_[1209]_  = \new_[54192]_  & \new_[54179]_ ;
  assign \new_[1210]_  = \new_[54166]_  & \new_[54153]_ ;
  assign \new_[1211]_  = \new_[54140]_  & \new_[54127]_ ;
  assign \new_[1212]_  = \new_[54114]_  & \new_[54101]_ ;
  assign \new_[1213]_  = \new_[54088]_  & \new_[54075]_ ;
  assign \new_[1214]_  = \new_[54062]_  & \new_[54049]_ ;
  assign \new_[1215]_  = \new_[54036]_  & \new_[54023]_ ;
  assign \new_[1216]_  = \new_[54010]_  & \new_[53997]_ ;
  assign \new_[1217]_  = \new_[53984]_  & \new_[53971]_ ;
  assign \new_[1218]_  = \new_[53958]_  & \new_[53945]_ ;
  assign \new_[1219]_  = \new_[53932]_  & \new_[53919]_ ;
  assign \new_[1220]_  = \new_[53906]_  & \new_[53893]_ ;
  assign \new_[1221]_  = \new_[53880]_  & \new_[53867]_ ;
  assign \new_[1222]_  = \new_[53854]_  & \new_[53841]_ ;
  assign \new_[1223]_  = \new_[53828]_  & \new_[53815]_ ;
  assign \new_[1224]_  = \new_[53802]_  & \new_[53789]_ ;
  assign \new_[1225]_  = \new_[53776]_  & \new_[53763]_ ;
  assign \new_[1226]_  = \new_[53750]_  & \new_[53737]_ ;
  assign \new_[1227]_  = \new_[53724]_  & \new_[53711]_ ;
  assign \new_[1228]_  = \new_[53698]_  & \new_[53685]_ ;
  assign \new_[1229]_  = \new_[53672]_  & \new_[53659]_ ;
  assign \new_[1230]_  = \new_[53646]_  & \new_[53633]_ ;
  assign \new_[1231]_  = \new_[53620]_  & \new_[53607]_ ;
  assign \new_[1232]_  = \new_[53594]_  & \new_[53581]_ ;
  assign \new_[1233]_  = \new_[53568]_  & \new_[53555]_ ;
  assign \new_[1234]_  = \new_[53542]_  & \new_[53529]_ ;
  assign \new_[1235]_  = \new_[53516]_  & \new_[53503]_ ;
  assign \new_[1236]_  = \new_[53490]_  & \new_[53477]_ ;
  assign \new_[1237]_  = \new_[53464]_  & \new_[53451]_ ;
  assign \new_[1238]_  = \new_[53438]_  & \new_[53425]_ ;
  assign \new_[1239]_  = \new_[53412]_  & \new_[53399]_ ;
  assign \new_[1240]_  = \new_[53386]_  & \new_[53373]_ ;
  assign \new_[1241]_  = \new_[53360]_  & \new_[53347]_ ;
  assign \new_[1242]_  = \new_[53334]_  & \new_[53321]_ ;
  assign \new_[1243]_  = \new_[53308]_  & \new_[53295]_ ;
  assign \new_[1244]_  = \new_[53282]_  & \new_[53269]_ ;
  assign \new_[1245]_  = \new_[53256]_  & \new_[53243]_ ;
  assign \new_[1246]_  = \new_[53230]_  & \new_[53217]_ ;
  assign \new_[1247]_  = \new_[53204]_  & \new_[53191]_ ;
  assign \new_[1248]_  = \new_[53178]_  & \new_[53165]_ ;
  assign \new_[1249]_  = \new_[53152]_  & \new_[53139]_ ;
  assign \new_[1250]_  = \new_[53126]_  & \new_[53113]_ ;
  assign \new_[1251]_  = \new_[53100]_  & \new_[53087]_ ;
  assign \new_[1252]_  = \new_[53074]_  & \new_[53061]_ ;
  assign \new_[1253]_  = \new_[53048]_  & \new_[53035]_ ;
  assign \new_[1254]_  = \new_[53022]_  & \new_[53009]_ ;
  assign \new_[1255]_  = \new_[52996]_  & \new_[52983]_ ;
  assign \new_[1256]_  = \new_[52970]_  & \new_[52957]_ ;
  assign \new_[1257]_  = \new_[52944]_  & \new_[52931]_ ;
  assign \new_[1258]_  = \new_[52918]_  & \new_[52905]_ ;
  assign \new_[1259]_  = \new_[52892]_  & \new_[52879]_ ;
  assign \new_[1260]_  = \new_[52866]_  & \new_[52853]_ ;
  assign \new_[1261]_  = \new_[52840]_  & \new_[52827]_ ;
  assign \new_[1262]_  = \new_[52814]_  & \new_[52801]_ ;
  assign \new_[1263]_  = \new_[52788]_  & \new_[52775]_ ;
  assign \new_[1264]_  = \new_[52762]_  & \new_[52749]_ ;
  assign \new_[1265]_  = \new_[52736]_  & \new_[52723]_ ;
  assign \new_[1266]_  = \new_[52710]_  & \new_[52697]_ ;
  assign \new_[1267]_  = \new_[52684]_  & \new_[52671]_ ;
  assign \new_[1268]_  = \new_[52658]_  & \new_[52645]_ ;
  assign \new_[1269]_  = \new_[52632]_  & \new_[52619]_ ;
  assign \new_[1270]_  = \new_[52606]_  & \new_[52593]_ ;
  assign \new_[1271]_  = \new_[52580]_  & \new_[52567]_ ;
  assign \new_[1272]_  = \new_[52554]_  & \new_[52541]_ ;
  assign \new_[1273]_  = \new_[52528]_  & \new_[52515]_ ;
  assign \new_[1274]_  = \new_[52502]_  & \new_[52489]_ ;
  assign \new_[1275]_  = \new_[52476]_  & \new_[52463]_ ;
  assign \new_[1276]_  = \new_[52450]_  & \new_[52437]_ ;
  assign \new_[1277]_  = \new_[52424]_  & \new_[52411]_ ;
  assign \new_[1278]_  = \new_[52398]_  & \new_[52385]_ ;
  assign \new_[1279]_  = \new_[52372]_  & \new_[52359]_ ;
  assign \new_[1280]_  = \new_[52346]_  & \new_[52333]_ ;
  assign \new_[1281]_  = \new_[52320]_  & \new_[52307]_ ;
  assign \new_[1282]_  = \new_[52294]_  & \new_[52281]_ ;
  assign \new_[1283]_  = \new_[52268]_  & \new_[52255]_ ;
  assign \new_[1284]_  = \new_[52242]_  & \new_[52229]_ ;
  assign \new_[1285]_  = \new_[52216]_  & \new_[52203]_ ;
  assign \new_[1286]_  = \new_[52190]_  & \new_[52177]_ ;
  assign \new_[1287]_  = \new_[52164]_  & \new_[52151]_ ;
  assign \new_[1288]_  = \new_[52138]_  & \new_[52125]_ ;
  assign \new_[1289]_  = \new_[52112]_  & \new_[52099]_ ;
  assign \new_[1290]_  = \new_[52086]_  & \new_[52073]_ ;
  assign \new_[1291]_  = \new_[52060]_  & \new_[52047]_ ;
  assign \new_[1292]_  = \new_[52034]_  & \new_[52021]_ ;
  assign \new_[1293]_  = \new_[52008]_  & \new_[51995]_ ;
  assign \new_[1294]_  = \new_[51982]_  & \new_[51969]_ ;
  assign \new_[1295]_  = \new_[51956]_  & \new_[51943]_ ;
  assign \new_[1296]_  = \new_[51930]_  & \new_[51917]_ ;
  assign \new_[1297]_  = \new_[51904]_  & \new_[51891]_ ;
  assign \new_[1298]_  = \new_[51878]_  & \new_[51865]_ ;
  assign \new_[1299]_  = \new_[51852]_  & \new_[51839]_ ;
  assign \new_[1300]_  = \new_[51826]_  & \new_[51813]_ ;
  assign \new_[1301]_  = \new_[51800]_  & \new_[51787]_ ;
  assign \new_[1302]_  = \new_[51774]_  & \new_[51761]_ ;
  assign \new_[1303]_  = \new_[51748]_  & \new_[51735]_ ;
  assign \new_[1304]_  = \new_[51722]_  & \new_[51709]_ ;
  assign \new_[1305]_  = \new_[51696]_  & \new_[51683]_ ;
  assign \new_[1306]_  = \new_[51670]_  & \new_[51657]_ ;
  assign \new_[1307]_  = \new_[51644]_  & \new_[51631]_ ;
  assign \new_[1308]_  = \new_[51618]_  & \new_[51605]_ ;
  assign \new_[1309]_  = \new_[51592]_  & \new_[51579]_ ;
  assign \new_[1310]_  = \new_[51566]_  & \new_[51553]_ ;
  assign \new_[1311]_  = \new_[51540]_  & \new_[51527]_ ;
  assign \new_[1312]_  = \new_[51514]_  & \new_[51501]_ ;
  assign \new_[1313]_  = \new_[51488]_  & \new_[51475]_ ;
  assign \new_[1314]_  = \new_[51462]_  & \new_[51449]_ ;
  assign \new_[1315]_  = \new_[51436]_  & \new_[51423]_ ;
  assign \new_[1316]_  = \new_[51410]_  & \new_[51397]_ ;
  assign \new_[1317]_  = \new_[51384]_  & \new_[51371]_ ;
  assign \new_[1318]_  = \new_[51358]_  & \new_[51345]_ ;
  assign \new_[1319]_  = \new_[51332]_  & \new_[51319]_ ;
  assign \new_[1320]_  = \new_[51306]_  & \new_[51293]_ ;
  assign \new_[1321]_  = \new_[51280]_  & \new_[51267]_ ;
  assign \new_[1322]_  = \new_[51254]_  & \new_[51241]_ ;
  assign \new_[1323]_  = \new_[51228]_  & \new_[51215]_ ;
  assign \new_[1324]_  = \new_[51202]_  & \new_[51189]_ ;
  assign \new_[1325]_  = \new_[51176]_  & \new_[51163]_ ;
  assign \new_[1326]_  = \new_[51150]_  & \new_[51137]_ ;
  assign \new_[1327]_  = \new_[51124]_  & \new_[51111]_ ;
  assign \new_[1328]_  = \new_[51098]_  & \new_[51085]_ ;
  assign \new_[1329]_  = \new_[51072]_  & \new_[51059]_ ;
  assign \new_[1330]_  = \new_[51046]_  & \new_[51033]_ ;
  assign \new_[1331]_  = \new_[51020]_  & \new_[51007]_ ;
  assign \new_[1332]_  = \new_[50994]_  & \new_[50981]_ ;
  assign \new_[1333]_  = \new_[50968]_  & \new_[50955]_ ;
  assign \new_[1334]_  = \new_[50942]_  & \new_[50929]_ ;
  assign \new_[1335]_  = \new_[50916]_  & \new_[50903]_ ;
  assign \new_[1336]_  = \new_[50890]_  & \new_[50877]_ ;
  assign \new_[1337]_  = \new_[50864]_  & \new_[50851]_ ;
  assign \new_[1338]_  = \new_[50838]_  & \new_[50825]_ ;
  assign \new_[1339]_  = \new_[50812]_  & \new_[50799]_ ;
  assign \new_[1340]_  = \new_[50786]_  & \new_[50773]_ ;
  assign \new_[1341]_  = \new_[50760]_  & \new_[50747]_ ;
  assign \new_[1342]_  = \new_[50734]_  & \new_[50721]_ ;
  assign \new_[1343]_  = \new_[50708]_  & \new_[50695]_ ;
  assign \new_[1344]_  = \new_[50682]_  & \new_[50669]_ ;
  assign \new_[1345]_  = \new_[50656]_  & \new_[50643]_ ;
  assign \new_[1346]_  = \new_[50630]_  & \new_[50617]_ ;
  assign \new_[1347]_  = \new_[50604]_  & \new_[50591]_ ;
  assign \new_[1348]_  = \new_[50578]_  & \new_[50565]_ ;
  assign \new_[1349]_  = \new_[50552]_  & \new_[50539]_ ;
  assign \new_[1350]_  = \new_[50526]_  & \new_[50513]_ ;
  assign \new_[1351]_  = \new_[50500]_  & \new_[50487]_ ;
  assign \new_[1352]_  = \new_[50474]_  & \new_[50461]_ ;
  assign \new_[1353]_  = \new_[50448]_  & \new_[50435]_ ;
  assign \new_[1354]_  = \new_[50422]_  & \new_[50409]_ ;
  assign \new_[1355]_  = \new_[50396]_  & \new_[50383]_ ;
  assign \new_[1356]_  = \new_[50370]_  & \new_[50357]_ ;
  assign \new_[1357]_  = \new_[50344]_  & \new_[50331]_ ;
  assign \new_[1358]_  = \new_[50318]_  & \new_[50305]_ ;
  assign \new_[1359]_  = \new_[50292]_  & \new_[50279]_ ;
  assign \new_[1360]_  = \new_[50266]_  & \new_[50253]_ ;
  assign \new_[1361]_  = \new_[50240]_  & \new_[50227]_ ;
  assign \new_[1362]_  = \new_[50214]_  & \new_[50201]_ ;
  assign \new_[1363]_  = \new_[50188]_  & \new_[50175]_ ;
  assign \new_[1364]_  = \new_[50162]_  & \new_[50149]_ ;
  assign \new_[1365]_  = \new_[50136]_  & \new_[50123]_ ;
  assign \new_[1366]_  = \new_[50110]_  & \new_[50097]_ ;
  assign \new_[1367]_  = \new_[50084]_  & \new_[50071]_ ;
  assign \new_[1368]_  = \new_[50058]_  & \new_[50045]_ ;
  assign \new_[1369]_  = \new_[50032]_  & \new_[50019]_ ;
  assign \new_[1370]_  = \new_[50006]_  & \new_[49993]_ ;
  assign \new_[1371]_  = \new_[49980]_  & \new_[49967]_ ;
  assign \new_[1372]_  = \new_[49954]_  & \new_[49941]_ ;
  assign \new_[1373]_  = \new_[49928]_  & \new_[49915]_ ;
  assign \new_[1374]_  = \new_[49902]_  & \new_[49889]_ ;
  assign \new_[1375]_  = \new_[49876]_  & \new_[49863]_ ;
  assign \new_[1376]_  = \new_[49850]_  & \new_[49837]_ ;
  assign \new_[1377]_  = \new_[49824]_  & \new_[49811]_ ;
  assign \new_[1378]_  = \new_[49798]_  & \new_[49785]_ ;
  assign \new_[1379]_  = \new_[49772]_  & \new_[49759]_ ;
  assign \new_[1380]_  = \new_[49746]_  & \new_[49733]_ ;
  assign \new_[1381]_  = \new_[49720]_  & \new_[49707]_ ;
  assign \new_[1382]_  = \new_[49694]_  & \new_[49681]_ ;
  assign \new_[1383]_  = \new_[49668]_  & \new_[49655]_ ;
  assign \new_[1384]_  = \new_[49642]_  & \new_[49629]_ ;
  assign \new_[1385]_  = \new_[49616]_  & \new_[49603]_ ;
  assign \new_[1386]_  = \new_[49590]_  & \new_[49577]_ ;
  assign \new_[1387]_  = \new_[49564]_  & \new_[49551]_ ;
  assign \new_[1388]_  = \new_[49538]_  & \new_[49525]_ ;
  assign \new_[1389]_  = \new_[49512]_  & \new_[49499]_ ;
  assign \new_[1390]_  = \new_[49486]_  & \new_[49473]_ ;
  assign \new_[1391]_  = \new_[49460]_  & \new_[49447]_ ;
  assign \new_[1392]_  = \new_[49434]_  & \new_[49421]_ ;
  assign \new_[1393]_  = \new_[49408]_  & \new_[49395]_ ;
  assign \new_[1394]_  = \new_[49382]_  & \new_[49369]_ ;
  assign \new_[1395]_  = \new_[49356]_  & \new_[49343]_ ;
  assign \new_[1396]_  = \new_[49330]_  & \new_[49317]_ ;
  assign \new_[1397]_  = \new_[49304]_  & \new_[49291]_ ;
  assign \new_[1398]_  = \new_[49278]_  & \new_[49265]_ ;
  assign \new_[1399]_  = \new_[49252]_  & \new_[49239]_ ;
  assign \new_[1400]_  = \new_[49226]_  & \new_[49213]_ ;
  assign \new_[1401]_  = \new_[49200]_  & \new_[49187]_ ;
  assign \new_[1402]_  = \new_[49174]_  & \new_[49161]_ ;
  assign \new_[1403]_  = \new_[49148]_  & \new_[49135]_ ;
  assign \new_[1404]_  = \new_[49122]_  & \new_[49109]_ ;
  assign \new_[1405]_  = \new_[49096]_  & \new_[49083]_ ;
  assign \new_[1406]_  = \new_[49070]_  & \new_[49057]_ ;
  assign \new_[1407]_  = \new_[49044]_  & \new_[49031]_ ;
  assign \new_[1408]_  = \new_[49018]_  & \new_[49005]_ ;
  assign \new_[1409]_  = \new_[48992]_  & \new_[48979]_ ;
  assign \new_[1410]_  = \new_[48966]_  & \new_[48953]_ ;
  assign \new_[1411]_  = \new_[48940]_  & \new_[48927]_ ;
  assign \new_[1412]_  = \new_[48914]_  & \new_[48901]_ ;
  assign \new_[1413]_  = \new_[48888]_  & \new_[48875]_ ;
  assign \new_[1414]_  = \new_[48862]_  & \new_[48849]_ ;
  assign \new_[1415]_  = \new_[48836]_  & \new_[48823]_ ;
  assign \new_[1416]_  = \new_[48810]_  & \new_[48797]_ ;
  assign \new_[1417]_  = \new_[48784]_  & \new_[48771]_ ;
  assign \new_[1418]_  = \new_[48758]_  & \new_[48745]_ ;
  assign \new_[1419]_  = \new_[48732]_  & \new_[48719]_ ;
  assign \new_[1420]_  = \new_[48706]_  & \new_[48693]_ ;
  assign \new_[1421]_  = \new_[48680]_  & \new_[48667]_ ;
  assign \new_[1422]_  = \new_[48654]_  & \new_[48641]_ ;
  assign \new_[1423]_  = \new_[48628]_  & \new_[48615]_ ;
  assign \new_[1424]_  = \new_[48602]_  & \new_[48589]_ ;
  assign \new_[1425]_  = \new_[48576]_  & \new_[48563]_ ;
  assign \new_[1426]_  = \new_[48550]_  & \new_[48537]_ ;
  assign \new_[1427]_  = \new_[48524]_  & \new_[48511]_ ;
  assign \new_[1428]_  = \new_[48498]_  & \new_[48485]_ ;
  assign \new_[1429]_  = \new_[48472]_  & \new_[48459]_ ;
  assign \new_[1430]_  = \new_[48446]_  & \new_[48433]_ ;
  assign \new_[1431]_  = \new_[48420]_  & \new_[48407]_ ;
  assign \new_[1432]_  = \new_[48394]_  & \new_[48381]_ ;
  assign \new_[1433]_  = \new_[48368]_  & \new_[48355]_ ;
  assign \new_[1434]_  = \new_[48342]_  & \new_[48329]_ ;
  assign \new_[1435]_  = \new_[48316]_  & \new_[48303]_ ;
  assign \new_[1436]_  = \new_[48290]_  & \new_[48277]_ ;
  assign \new_[1437]_  = \new_[48264]_  & \new_[48251]_ ;
  assign \new_[1438]_  = \new_[48238]_  & \new_[48225]_ ;
  assign \new_[1439]_  = \new_[48212]_  & \new_[48199]_ ;
  assign \new_[1440]_  = \new_[48186]_  & \new_[48173]_ ;
  assign \new_[1441]_  = \new_[48160]_  & \new_[48147]_ ;
  assign \new_[1442]_  = \new_[48134]_  & \new_[48121]_ ;
  assign \new_[1443]_  = \new_[48108]_  & \new_[48095]_ ;
  assign \new_[1444]_  = \new_[48082]_  & \new_[48069]_ ;
  assign \new_[1445]_  = \new_[48056]_  & \new_[48043]_ ;
  assign \new_[1446]_  = \new_[48030]_  & \new_[48017]_ ;
  assign \new_[1447]_  = \new_[48004]_  & \new_[47991]_ ;
  assign \new_[1448]_  = \new_[47978]_  & \new_[47965]_ ;
  assign \new_[1449]_  = \new_[47952]_  & \new_[47939]_ ;
  assign \new_[1450]_  = \new_[47926]_  & \new_[47913]_ ;
  assign \new_[1451]_  = \new_[47900]_  & \new_[47887]_ ;
  assign \new_[1452]_  = \new_[47874]_  & \new_[47861]_ ;
  assign \new_[1453]_  = \new_[47848]_  & \new_[47835]_ ;
  assign \new_[1454]_  = \new_[47822]_  & \new_[47809]_ ;
  assign \new_[1455]_  = \new_[47796]_  & \new_[47783]_ ;
  assign \new_[1456]_  = \new_[47770]_  & \new_[47757]_ ;
  assign \new_[1457]_  = \new_[47744]_  & \new_[47731]_ ;
  assign \new_[1458]_  = \new_[47718]_  & \new_[47705]_ ;
  assign \new_[1459]_  = \new_[47692]_  & \new_[47679]_ ;
  assign \new_[1460]_  = \new_[47666]_  & \new_[47653]_ ;
  assign \new_[1461]_  = \new_[47640]_  & \new_[47627]_ ;
  assign \new_[1462]_  = \new_[47614]_  & \new_[47601]_ ;
  assign \new_[1463]_  = \new_[47588]_  & \new_[47575]_ ;
  assign \new_[1464]_  = \new_[47562]_  & \new_[47549]_ ;
  assign \new_[1465]_  = \new_[47536]_  & \new_[47523]_ ;
  assign \new_[1466]_  = \new_[47510]_  & \new_[47497]_ ;
  assign \new_[1467]_  = \new_[47484]_  & \new_[47471]_ ;
  assign \new_[1468]_  = \new_[47458]_  & \new_[47445]_ ;
  assign \new_[1469]_  = \new_[47432]_  & \new_[47419]_ ;
  assign \new_[1470]_  = \new_[47406]_  & \new_[47393]_ ;
  assign \new_[1471]_  = \new_[47380]_  & \new_[47367]_ ;
  assign \new_[1472]_  = \new_[47354]_  & \new_[47341]_ ;
  assign \new_[1473]_  = \new_[47328]_  & \new_[47315]_ ;
  assign \new_[1474]_  = \new_[47302]_  & \new_[47289]_ ;
  assign \new_[1475]_  = \new_[47276]_  & \new_[47263]_ ;
  assign \new_[1476]_  = \new_[47250]_  & \new_[47237]_ ;
  assign \new_[1477]_  = \new_[47224]_  & \new_[47211]_ ;
  assign \new_[1478]_  = \new_[47198]_  & \new_[47185]_ ;
  assign \new_[1479]_  = \new_[47172]_  & \new_[47159]_ ;
  assign \new_[1480]_  = \new_[47146]_  & \new_[47133]_ ;
  assign \new_[1481]_  = \new_[47120]_  & \new_[47107]_ ;
  assign \new_[1482]_  = \new_[47094]_  & \new_[47081]_ ;
  assign \new_[1483]_  = \new_[47068]_  & \new_[47055]_ ;
  assign \new_[1484]_  = \new_[47042]_  & \new_[47029]_ ;
  assign \new_[1485]_  = \new_[47016]_  & \new_[47003]_ ;
  assign \new_[1486]_  = \new_[46990]_  & \new_[46977]_ ;
  assign \new_[1487]_  = \new_[46964]_  & \new_[46951]_ ;
  assign \new_[1488]_  = \new_[46938]_  & \new_[46925]_ ;
  assign \new_[1489]_  = \new_[46912]_  & \new_[46899]_ ;
  assign \new_[1490]_  = \new_[46886]_  & \new_[46873]_ ;
  assign \new_[1491]_  = \new_[46860]_  & \new_[46847]_ ;
  assign \new_[1492]_  = \new_[46834]_  & \new_[46821]_ ;
  assign \new_[1493]_  = \new_[46808]_  & \new_[46795]_ ;
  assign \new_[1494]_  = \new_[46782]_  & \new_[46769]_ ;
  assign \new_[1495]_  = \new_[46756]_  & \new_[46743]_ ;
  assign \new_[1496]_  = \new_[46730]_  & \new_[46717]_ ;
  assign \new_[1497]_  = \new_[46704]_  & \new_[46691]_ ;
  assign \new_[1498]_  = \new_[46678]_  & \new_[46665]_ ;
  assign \new_[1499]_  = \new_[46652]_  & \new_[46639]_ ;
  assign \new_[1500]_  = \new_[46626]_  & \new_[46613]_ ;
  assign \new_[1501]_  = \new_[46600]_  & \new_[46587]_ ;
  assign \new_[1502]_  = \new_[46574]_  & \new_[46561]_ ;
  assign \new_[1503]_  = \new_[46548]_  & \new_[46535]_ ;
  assign \new_[1504]_  = \new_[46522]_  & \new_[46509]_ ;
  assign \new_[1505]_  = \new_[46496]_  & \new_[46483]_ ;
  assign \new_[1506]_  = \new_[46470]_  & \new_[46457]_ ;
  assign \new_[1507]_  = \new_[46444]_  & \new_[46431]_ ;
  assign \new_[1508]_  = \new_[46418]_  & \new_[46405]_ ;
  assign \new_[1509]_  = \new_[46392]_  & \new_[46379]_ ;
  assign \new_[1510]_  = \new_[46366]_  & \new_[46353]_ ;
  assign \new_[1511]_  = \new_[46340]_  & \new_[46327]_ ;
  assign \new_[1512]_  = \new_[46314]_  & \new_[46301]_ ;
  assign \new_[1513]_  = \new_[46288]_  & \new_[46275]_ ;
  assign \new_[1514]_  = \new_[46262]_  & \new_[46249]_ ;
  assign \new_[1515]_  = \new_[46236]_  & \new_[46223]_ ;
  assign \new_[1516]_  = \new_[46210]_  & \new_[46197]_ ;
  assign \new_[1517]_  = \new_[46184]_  & \new_[46171]_ ;
  assign \new_[1518]_  = \new_[46158]_  & \new_[46145]_ ;
  assign \new_[1519]_  = \new_[46132]_  & \new_[46119]_ ;
  assign \new_[1520]_  = \new_[46106]_  & \new_[46093]_ ;
  assign \new_[1521]_  = \new_[46080]_  & \new_[46067]_ ;
  assign \new_[1522]_  = \new_[46054]_  & \new_[46041]_ ;
  assign \new_[1523]_  = \new_[46028]_  & \new_[46015]_ ;
  assign \new_[1524]_  = \new_[46002]_  & \new_[45989]_ ;
  assign \new_[1525]_  = \new_[45976]_  & \new_[45963]_ ;
  assign \new_[1526]_  = \new_[45950]_  & \new_[45937]_ ;
  assign \new_[1527]_  = \new_[45924]_  & \new_[45911]_ ;
  assign \new_[1528]_  = \new_[45898]_  & \new_[45885]_ ;
  assign \new_[1529]_  = \new_[45872]_  & \new_[45859]_ ;
  assign \new_[1530]_  = \new_[45846]_  & \new_[45833]_ ;
  assign \new_[1531]_  = \new_[45820]_  & \new_[45807]_ ;
  assign \new_[1532]_  = \new_[45794]_  & \new_[45781]_ ;
  assign \new_[1533]_  = \new_[45768]_  & \new_[45755]_ ;
  assign \new_[1534]_  = \new_[45742]_  & \new_[45729]_ ;
  assign \new_[1535]_  = \new_[45716]_  & \new_[45703]_ ;
  assign \new_[1536]_  = \new_[45690]_  & \new_[45677]_ ;
  assign \new_[1537]_  = \new_[45664]_  & \new_[45651]_ ;
  assign \new_[1538]_  = \new_[45638]_  & \new_[45625]_ ;
  assign \new_[1539]_  = \new_[45612]_  & \new_[45599]_ ;
  assign \new_[1540]_  = \new_[45586]_  & \new_[45573]_ ;
  assign \new_[1541]_  = \new_[45560]_  & \new_[45547]_ ;
  assign \new_[1542]_  = \new_[45534]_  & \new_[45521]_ ;
  assign \new_[1543]_  = \new_[45508]_  & \new_[45495]_ ;
  assign \new_[1544]_  = \new_[45482]_  & \new_[45469]_ ;
  assign \new_[1545]_  = \new_[45456]_  & \new_[45443]_ ;
  assign \new_[1546]_  = \new_[45430]_  & \new_[45417]_ ;
  assign \new_[1547]_  = \new_[45404]_  & \new_[45391]_ ;
  assign \new_[1548]_  = \new_[45378]_  & \new_[45365]_ ;
  assign \new_[1549]_  = \new_[45352]_  & \new_[45339]_ ;
  assign \new_[1550]_  = \new_[45326]_  & \new_[45313]_ ;
  assign \new_[1551]_  = \new_[45300]_  & \new_[45287]_ ;
  assign \new_[1552]_  = \new_[45274]_  & \new_[45261]_ ;
  assign \new_[1553]_  = \new_[45248]_  & \new_[45235]_ ;
  assign \new_[1554]_  = \new_[45222]_  & \new_[45209]_ ;
  assign \new_[1555]_  = \new_[45196]_  & \new_[45183]_ ;
  assign \new_[1556]_  = \new_[45170]_  & \new_[45157]_ ;
  assign \new_[1557]_  = \new_[45144]_  & \new_[45131]_ ;
  assign \new_[1558]_  = \new_[45118]_  & \new_[45105]_ ;
  assign \new_[1559]_  = \new_[45092]_  & \new_[45079]_ ;
  assign \new_[1560]_  = \new_[45066]_  & \new_[45053]_ ;
  assign \new_[1561]_  = \new_[45040]_  & \new_[45027]_ ;
  assign \new_[1562]_  = \new_[45014]_  & \new_[45001]_ ;
  assign \new_[1563]_  = \new_[44988]_  & \new_[44975]_ ;
  assign \new_[1564]_  = \new_[44962]_  & \new_[44949]_ ;
  assign \new_[1565]_  = \new_[44936]_  & \new_[44923]_ ;
  assign \new_[1566]_  = \new_[44910]_  & \new_[44897]_ ;
  assign \new_[1567]_  = \new_[44884]_  & \new_[44871]_ ;
  assign \new_[1568]_  = \new_[44858]_  & \new_[44845]_ ;
  assign \new_[1569]_  = \new_[44832]_  & \new_[44819]_ ;
  assign \new_[1570]_  = \new_[44806]_  & \new_[44793]_ ;
  assign \new_[1571]_  = \new_[44780]_  & \new_[44767]_ ;
  assign \new_[1572]_  = \new_[44754]_  & \new_[44741]_ ;
  assign \new_[1573]_  = \new_[44728]_  & \new_[44715]_ ;
  assign \new_[1574]_  = \new_[44702]_  & \new_[44689]_ ;
  assign \new_[1575]_  = \new_[44676]_  & \new_[44663]_ ;
  assign \new_[1576]_  = \new_[44650]_  & \new_[44637]_ ;
  assign \new_[1577]_  = \new_[44624]_  & \new_[44611]_ ;
  assign \new_[1578]_  = \new_[44598]_  & \new_[44585]_ ;
  assign \new_[1579]_  = \new_[44572]_  & \new_[44559]_ ;
  assign \new_[1580]_  = \new_[44546]_  & \new_[44533]_ ;
  assign \new_[1581]_  = \new_[44520]_  & \new_[44507]_ ;
  assign \new_[1582]_  = \new_[44494]_  & \new_[44481]_ ;
  assign \new_[1583]_  = \new_[44468]_  & \new_[44455]_ ;
  assign \new_[1584]_  = \new_[44442]_  & \new_[44429]_ ;
  assign \new_[1585]_  = \new_[44416]_  & \new_[44403]_ ;
  assign \new_[1586]_  = \new_[44390]_  & \new_[44377]_ ;
  assign \new_[1587]_  = \new_[44364]_  & \new_[44351]_ ;
  assign \new_[1588]_  = \new_[44338]_  & \new_[44325]_ ;
  assign \new_[1589]_  = \new_[44312]_  & \new_[44299]_ ;
  assign \new_[1590]_  = \new_[44286]_  & \new_[44273]_ ;
  assign \new_[1591]_  = \new_[44260]_  & \new_[44247]_ ;
  assign \new_[1592]_  = \new_[44234]_  & \new_[44221]_ ;
  assign \new_[1593]_  = \new_[44208]_  & \new_[44195]_ ;
  assign \new_[1594]_  = \new_[44182]_  & \new_[44169]_ ;
  assign \new_[1595]_  = \new_[44156]_  & \new_[44143]_ ;
  assign \new_[1596]_  = \new_[44130]_  & \new_[44117]_ ;
  assign \new_[1597]_  = \new_[44104]_  & \new_[44091]_ ;
  assign \new_[1598]_  = \new_[44078]_  & \new_[44065]_ ;
  assign \new_[1599]_  = \new_[44052]_  & \new_[44039]_ ;
  assign \new_[1600]_  = \new_[44026]_  & \new_[44013]_ ;
  assign \new_[1601]_  = \new_[44000]_  & \new_[43987]_ ;
  assign \new_[1602]_  = \new_[43974]_  & \new_[43961]_ ;
  assign \new_[1603]_  = \new_[43948]_  & \new_[43935]_ ;
  assign \new_[1604]_  = \new_[43922]_  & \new_[43909]_ ;
  assign \new_[1605]_  = \new_[43896]_  & \new_[43883]_ ;
  assign \new_[1606]_  = \new_[43870]_  & \new_[43857]_ ;
  assign \new_[1607]_  = \new_[43844]_  & \new_[43831]_ ;
  assign \new_[1608]_  = \new_[43818]_  & \new_[43805]_ ;
  assign \new_[1609]_  = \new_[43792]_  & \new_[43779]_ ;
  assign \new_[1610]_  = \new_[43766]_  & \new_[43753]_ ;
  assign \new_[1611]_  = \new_[43740]_  & \new_[43727]_ ;
  assign \new_[1612]_  = \new_[43714]_  & \new_[43701]_ ;
  assign \new_[1613]_  = \new_[43688]_  & \new_[43675]_ ;
  assign \new_[1614]_  = \new_[43662]_  & \new_[43649]_ ;
  assign \new_[1615]_  = \new_[43636]_  & \new_[43623]_ ;
  assign \new_[1616]_  = \new_[43610]_  & \new_[43597]_ ;
  assign \new_[1617]_  = \new_[43584]_  & \new_[43571]_ ;
  assign \new_[1618]_  = \new_[43558]_  & \new_[43545]_ ;
  assign \new_[1619]_  = \new_[43532]_  & \new_[43519]_ ;
  assign \new_[1620]_  = \new_[43506]_  & \new_[43493]_ ;
  assign \new_[1621]_  = \new_[43480]_  & \new_[43467]_ ;
  assign \new_[1622]_  = \new_[43454]_  & \new_[43441]_ ;
  assign \new_[1623]_  = \new_[43428]_  & \new_[43415]_ ;
  assign \new_[1624]_  = \new_[43402]_  & \new_[43389]_ ;
  assign \new_[1625]_  = \new_[43376]_  & \new_[43363]_ ;
  assign \new_[1626]_  = \new_[43350]_  & \new_[43337]_ ;
  assign \new_[1627]_  = \new_[43324]_  & \new_[43311]_ ;
  assign \new_[1628]_  = \new_[43298]_  & \new_[43285]_ ;
  assign \new_[1629]_  = \new_[43272]_  & \new_[43259]_ ;
  assign \new_[1630]_  = \new_[43246]_  & \new_[43233]_ ;
  assign \new_[1631]_  = \new_[43220]_  & \new_[43207]_ ;
  assign \new_[1632]_  = \new_[43194]_  & \new_[43181]_ ;
  assign \new_[1633]_  = \new_[43168]_  & \new_[43155]_ ;
  assign \new_[1634]_  = \new_[43142]_  & \new_[43129]_ ;
  assign \new_[1635]_  = \new_[43116]_  & \new_[43103]_ ;
  assign \new_[1636]_  = \new_[43090]_  & \new_[43077]_ ;
  assign \new_[1637]_  = \new_[43064]_  & \new_[43051]_ ;
  assign \new_[1638]_  = \new_[43038]_  & \new_[43025]_ ;
  assign \new_[1639]_  = \new_[43012]_  & \new_[42999]_ ;
  assign \new_[1640]_  = \new_[42986]_  & \new_[42973]_ ;
  assign \new_[1641]_  = \new_[42960]_  & \new_[42947]_ ;
  assign \new_[1642]_  = \new_[42934]_  & \new_[42921]_ ;
  assign \new_[1643]_  = \new_[42908]_  & \new_[42895]_ ;
  assign \new_[1644]_  = \new_[42882]_  & \new_[42869]_ ;
  assign \new_[1645]_  = \new_[42856]_  & \new_[42843]_ ;
  assign \new_[1646]_  = \new_[42830]_  & \new_[42817]_ ;
  assign \new_[1647]_  = \new_[42804]_  & \new_[42791]_ ;
  assign \new_[1648]_  = \new_[42778]_  & \new_[42765]_ ;
  assign \new_[1649]_  = \new_[42752]_  & \new_[42739]_ ;
  assign \new_[1650]_  = \new_[42726]_  & \new_[42713]_ ;
  assign \new_[1651]_  = \new_[42700]_  & \new_[42687]_ ;
  assign \new_[1652]_  = \new_[42674]_  & \new_[42661]_ ;
  assign \new_[1653]_  = \new_[42648]_  & \new_[42635]_ ;
  assign \new_[1654]_  = \new_[42622]_  & \new_[42609]_ ;
  assign \new_[1655]_  = \new_[42596]_  & \new_[42583]_ ;
  assign \new_[1656]_  = \new_[42570]_  & \new_[42557]_ ;
  assign \new_[1657]_  = \new_[42544]_  & \new_[42531]_ ;
  assign \new_[1658]_  = \new_[42518]_  & \new_[42505]_ ;
  assign \new_[1659]_  = \new_[42492]_  & \new_[42479]_ ;
  assign \new_[1660]_  = \new_[42468]_  & \new_[42455]_ ;
  assign \new_[1661]_  = \new_[42444]_  & \new_[42431]_ ;
  assign \new_[1662]_  = \new_[42420]_  & \new_[42407]_ ;
  assign \new_[1663]_  = \new_[42396]_  & \new_[42383]_ ;
  assign \new_[1664]_  = \new_[42372]_  & \new_[42359]_ ;
  assign \new_[1665]_  = \new_[42348]_  & \new_[42335]_ ;
  assign \new_[1666]_  = \new_[42324]_  & \new_[42311]_ ;
  assign \new_[1667]_  = \new_[42300]_  & \new_[42287]_ ;
  assign \new_[1668]_  = \new_[42276]_  & \new_[42263]_ ;
  assign \new_[1669]_  = \new_[42252]_  & \new_[42239]_ ;
  assign \new_[1670]_  = \new_[42228]_  & \new_[42215]_ ;
  assign \new_[1671]_  = \new_[42204]_  & \new_[42191]_ ;
  assign \new_[1672]_  = \new_[42180]_  & \new_[42167]_ ;
  assign \new_[1673]_  = \new_[42156]_  & \new_[42143]_ ;
  assign \new_[1674]_  = \new_[42132]_  & \new_[42119]_ ;
  assign \new_[1675]_  = \new_[42108]_  & \new_[42095]_ ;
  assign \new_[1676]_  = \new_[42084]_  & \new_[42071]_ ;
  assign \new_[1677]_  = \new_[42060]_  & \new_[42047]_ ;
  assign \new_[1678]_  = \new_[42036]_  & \new_[42023]_ ;
  assign \new_[1679]_  = \new_[42012]_  & \new_[41999]_ ;
  assign \new_[1680]_  = \new_[41988]_  & \new_[41975]_ ;
  assign \new_[1681]_  = \new_[41964]_  & \new_[41951]_ ;
  assign \new_[1682]_  = \new_[41940]_  & \new_[41927]_ ;
  assign \new_[1683]_  = \new_[41916]_  & \new_[41903]_ ;
  assign \new_[1684]_  = \new_[41892]_  & \new_[41879]_ ;
  assign \new_[1685]_  = \new_[41868]_  & \new_[41855]_ ;
  assign \new_[1686]_  = \new_[41844]_  & \new_[41831]_ ;
  assign \new_[1687]_  = \new_[41820]_  & \new_[41807]_ ;
  assign \new_[1688]_  = \new_[41796]_  & \new_[41783]_ ;
  assign \new_[1689]_  = \new_[41772]_  & \new_[41759]_ ;
  assign \new_[1690]_  = \new_[41748]_  & \new_[41735]_ ;
  assign \new_[1691]_  = \new_[41724]_  & \new_[41711]_ ;
  assign \new_[1692]_  = \new_[41700]_  & \new_[41687]_ ;
  assign \new_[1693]_  = \new_[41676]_  & \new_[41663]_ ;
  assign \new_[1694]_  = \new_[41652]_  & \new_[41639]_ ;
  assign \new_[1695]_  = \new_[41628]_  & \new_[41615]_ ;
  assign \new_[1696]_  = \new_[41604]_  & \new_[41591]_ ;
  assign \new_[1697]_  = \new_[41580]_  & \new_[41567]_ ;
  assign \new_[1698]_  = \new_[41556]_  & \new_[41543]_ ;
  assign \new_[1699]_  = \new_[41532]_  & \new_[41519]_ ;
  assign \new_[1700]_  = \new_[41508]_  & \new_[41495]_ ;
  assign \new_[1701]_  = \new_[41484]_  & \new_[41471]_ ;
  assign \new_[1702]_  = \new_[41460]_  & \new_[41447]_ ;
  assign \new_[1703]_  = \new_[41436]_  & \new_[41423]_ ;
  assign \new_[1704]_  = \new_[41412]_  & \new_[41399]_ ;
  assign \new_[1705]_  = \new_[41388]_  & \new_[41375]_ ;
  assign \new_[1706]_  = \new_[41364]_  & \new_[41351]_ ;
  assign \new_[1707]_  = \new_[41340]_  & \new_[41327]_ ;
  assign \new_[1708]_  = \new_[41316]_  & \new_[41303]_ ;
  assign \new_[1709]_  = \new_[41292]_  & \new_[41279]_ ;
  assign \new_[1710]_  = \new_[41268]_  & \new_[41255]_ ;
  assign \new_[1711]_  = \new_[41244]_  & \new_[41231]_ ;
  assign \new_[1712]_  = \new_[41220]_  & \new_[41207]_ ;
  assign \new_[1713]_  = \new_[41196]_  & \new_[41183]_ ;
  assign \new_[1714]_  = \new_[41172]_  & \new_[41159]_ ;
  assign \new_[1715]_  = \new_[41148]_  & \new_[41135]_ ;
  assign \new_[1716]_  = \new_[41124]_  & \new_[41111]_ ;
  assign \new_[1717]_  = \new_[41100]_  & \new_[41087]_ ;
  assign \new_[1718]_  = \new_[41076]_  & \new_[41063]_ ;
  assign \new_[1719]_  = \new_[41052]_  & \new_[41039]_ ;
  assign \new_[1720]_  = \new_[41028]_  & \new_[41015]_ ;
  assign \new_[1721]_  = \new_[41004]_  & \new_[40991]_ ;
  assign \new_[1722]_  = \new_[40980]_  & \new_[40967]_ ;
  assign \new_[1723]_  = \new_[40956]_  & \new_[40943]_ ;
  assign \new_[1724]_  = \new_[40932]_  & \new_[40919]_ ;
  assign \new_[1725]_  = \new_[40908]_  & \new_[40895]_ ;
  assign \new_[1726]_  = \new_[40884]_  & \new_[40871]_ ;
  assign \new_[1727]_  = \new_[40860]_  & \new_[40847]_ ;
  assign \new_[1728]_  = \new_[40836]_  & \new_[40823]_ ;
  assign \new_[1729]_  = \new_[40812]_  & \new_[40799]_ ;
  assign \new_[1730]_  = \new_[40788]_  & \new_[40775]_ ;
  assign \new_[1731]_  = \new_[40764]_  & \new_[40751]_ ;
  assign \new_[1732]_  = \new_[40740]_  & \new_[40727]_ ;
  assign \new_[1733]_  = \new_[40716]_  & \new_[40703]_ ;
  assign \new_[1734]_  = \new_[40692]_  & \new_[40679]_ ;
  assign \new_[1735]_  = \new_[40668]_  & \new_[40655]_ ;
  assign \new_[1736]_  = \new_[40644]_  & \new_[40631]_ ;
  assign \new_[1737]_  = \new_[40620]_  & \new_[40607]_ ;
  assign \new_[1738]_  = \new_[40596]_  & \new_[40583]_ ;
  assign \new_[1739]_  = \new_[40572]_  & \new_[40559]_ ;
  assign \new_[1740]_  = \new_[40548]_  & \new_[40535]_ ;
  assign \new_[1741]_  = \new_[40524]_  & \new_[40511]_ ;
  assign \new_[1742]_  = \new_[40500]_  & \new_[40487]_ ;
  assign \new_[1743]_  = \new_[40476]_  & \new_[40463]_ ;
  assign \new_[1744]_  = \new_[40452]_  & \new_[40439]_ ;
  assign \new_[1745]_  = \new_[40428]_  & \new_[40415]_ ;
  assign \new_[1746]_  = \new_[40404]_  & \new_[40391]_ ;
  assign \new_[1747]_  = \new_[40380]_  & \new_[40367]_ ;
  assign \new_[1748]_  = \new_[40356]_  & \new_[40343]_ ;
  assign \new_[1749]_  = \new_[40332]_  & \new_[40319]_ ;
  assign \new_[1750]_  = \new_[40308]_  & \new_[40295]_ ;
  assign \new_[1751]_  = \new_[40284]_  & \new_[40271]_ ;
  assign \new_[1752]_  = \new_[40260]_  & \new_[40247]_ ;
  assign \new_[1753]_  = \new_[40236]_  & \new_[40223]_ ;
  assign \new_[1754]_  = \new_[40212]_  & \new_[40199]_ ;
  assign \new_[1755]_  = \new_[40188]_  & \new_[40175]_ ;
  assign \new_[1756]_  = \new_[40164]_  & \new_[40151]_ ;
  assign \new_[1757]_  = \new_[40140]_  & \new_[40127]_ ;
  assign \new_[1758]_  = \new_[40116]_  & \new_[40103]_ ;
  assign \new_[1759]_  = \new_[40092]_  & \new_[40079]_ ;
  assign \new_[1760]_  = \new_[40068]_  & \new_[40055]_ ;
  assign \new_[1761]_  = \new_[40044]_  & \new_[40031]_ ;
  assign \new_[1762]_  = \new_[40020]_  & \new_[40007]_ ;
  assign \new_[1763]_  = \new_[39996]_  & \new_[39983]_ ;
  assign \new_[1764]_  = \new_[39972]_  & \new_[39959]_ ;
  assign \new_[1765]_  = \new_[39948]_  & \new_[39935]_ ;
  assign \new_[1766]_  = \new_[39924]_  & \new_[39911]_ ;
  assign \new_[1767]_  = \new_[39900]_  & \new_[39887]_ ;
  assign \new_[1768]_  = \new_[39876]_  & \new_[39863]_ ;
  assign \new_[1769]_  = \new_[39852]_  & \new_[39839]_ ;
  assign \new_[1770]_  = \new_[39828]_  & \new_[39815]_ ;
  assign \new_[1771]_  = \new_[39804]_  & \new_[39791]_ ;
  assign \new_[1772]_  = \new_[39780]_  & \new_[39767]_ ;
  assign \new_[1773]_  = \new_[39756]_  & \new_[39743]_ ;
  assign \new_[1774]_  = \new_[39732]_  & \new_[39719]_ ;
  assign \new_[1775]_  = \new_[39708]_  & \new_[39695]_ ;
  assign \new_[1776]_  = \new_[39684]_  & \new_[39671]_ ;
  assign \new_[1777]_  = \new_[39660]_  & \new_[39647]_ ;
  assign \new_[1778]_  = \new_[39636]_  & \new_[39623]_ ;
  assign \new_[1779]_  = \new_[39612]_  & \new_[39599]_ ;
  assign \new_[1780]_  = \new_[39588]_  & \new_[39575]_ ;
  assign \new_[1781]_  = \new_[39564]_  & \new_[39551]_ ;
  assign \new_[1782]_  = \new_[39540]_  & \new_[39527]_ ;
  assign \new_[1783]_  = \new_[39516]_  & \new_[39503]_ ;
  assign \new_[1784]_  = \new_[39492]_  & \new_[39479]_ ;
  assign \new_[1785]_  = \new_[39468]_  & \new_[39455]_ ;
  assign \new_[1786]_  = \new_[39444]_  & \new_[39431]_ ;
  assign \new_[1787]_  = \new_[39420]_  & \new_[39407]_ ;
  assign \new_[1788]_  = \new_[39396]_  & \new_[39383]_ ;
  assign \new_[1789]_  = \new_[39372]_  & \new_[39359]_ ;
  assign \new_[1790]_  = \new_[39348]_  & \new_[39335]_ ;
  assign \new_[1791]_  = \new_[39324]_  & \new_[39311]_ ;
  assign \new_[1792]_  = \new_[39300]_  & \new_[39287]_ ;
  assign \new_[1793]_  = \new_[39276]_  & \new_[39263]_ ;
  assign \new_[1794]_  = \new_[39252]_  & \new_[39239]_ ;
  assign \new_[1795]_  = \new_[39228]_  & \new_[39215]_ ;
  assign \new_[1796]_  = \new_[39204]_  & \new_[39191]_ ;
  assign \new_[1797]_  = \new_[39180]_  & \new_[39167]_ ;
  assign \new_[1798]_  = \new_[39156]_  & \new_[39143]_ ;
  assign \new_[1799]_  = \new_[39132]_  & \new_[39119]_ ;
  assign \new_[1800]_  = \new_[39108]_  & \new_[39095]_ ;
  assign \new_[1801]_  = \new_[39084]_  & \new_[39071]_ ;
  assign \new_[1802]_  = \new_[39060]_  & \new_[39047]_ ;
  assign \new_[1803]_  = \new_[39036]_  & \new_[39023]_ ;
  assign \new_[1804]_  = \new_[39012]_  & \new_[38999]_ ;
  assign \new_[1805]_  = \new_[38988]_  & \new_[38975]_ ;
  assign \new_[1806]_  = \new_[38964]_  & \new_[38951]_ ;
  assign \new_[1807]_  = \new_[38940]_  & \new_[38927]_ ;
  assign \new_[1808]_  = \new_[38916]_  & \new_[38903]_ ;
  assign \new_[1809]_  = \new_[38892]_  & \new_[38879]_ ;
  assign \new_[1810]_  = \new_[38868]_  & \new_[38855]_ ;
  assign \new_[1811]_  = \new_[38844]_  & \new_[38831]_ ;
  assign \new_[1812]_  = \new_[38820]_  & \new_[38807]_ ;
  assign \new_[1813]_  = \new_[38796]_  & \new_[38783]_ ;
  assign \new_[1814]_  = \new_[38772]_  & \new_[38759]_ ;
  assign \new_[1815]_  = \new_[38748]_  & \new_[38735]_ ;
  assign \new_[1816]_  = \new_[38724]_  & \new_[38711]_ ;
  assign \new_[1817]_  = \new_[38700]_  & \new_[38687]_ ;
  assign \new_[1818]_  = \new_[38676]_  & \new_[38663]_ ;
  assign \new_[1819]_  = \new_[38652]_  & \new_[38639]_ ;
  assign \new_[1820]_  = \new_[38628]_  & \new_[38615]_ ;
  assign \new_[1821]_  = \new_[38604]_  & \new_[38591]_ ;
  assign \new_[1822]_  = \new_[38580]_  & \new_[38567]_ ;
  assign \new_[1823]_  = \new_[38556]_  & \new_[38543]_ ;
  assign \new_[1824]_  = \new_[38532]_  & \new_[38519]_ ;
  assign \new_[1825]_  = \new_[38508]_  & \new_[38495]_ ;
  assign \new_[1826]_  = \new_[38484]_  & \new_[38471]_ ;
  assign \new_[1827]_  = \new_[38460]_  & \new_[38447]_ ;
  assign \new_[1828]_  = \new_[38436]_  & \new_[38423]_ ;
  assign \new_[1829]_  = \new_[38412]_  & \new_[38399]_ ;
  assign \new_[1830]_  = \new_[38388]_  & \new_[38375]_ ;
  assign \new_[1831]_  = \new_[38364]_  & \new_[38351]_ ;
  assign \new_[1832]_  = \new_[38340]_  & \new_[38327]_ ;
  assign \new_[1833]_  = \new_[38316]_  & \new_[38303]_ ;
  assign \new_[1834]_  = \new_[38292]_  & \new_[38279]_ ;
  assign \new_[1835]_  = \new_[38268]_  & \new_[38255]_ ;
  assign \new_[1836]_  = \new_[38244]_  & \new_[38231]_ ;
  assign \new_[1837]_  = \new_[38220]_  & \new_[38207]_ ;
  assign \new_[1838]_  = \new_[38196]_  & \new_[38183]_ ;
  assign \new_[1839]_  = \new_[38172]_  & \new_[38159]_ ;
  assign \new_[1840]_  = \new_[38148]_  & \new_[38135]_ ;
  assign \new_[1841]_  = \new_[38124]_  & \new_[38111]_ ;
  assign \new_[1842]_  = \new_[38100]_  & \new_[38087]_ ;
  assign \new_[1843]_  = \new_[38076]_  & \new_[38063]_ ;
  assign \new_[1844]_  = \new_[38052]_  & \new_[38039]_ ;
  assign \new_[1845]_  = \new_[38028]_  & \new_[38015]_ ;
  assign \new_[1846]_  = \new_[38004]_  & \new_[37991]_ ;
  assign \new_[1847]_  = \new_[37980]_  & \new_[37967]_ ;
  assign \new_[1848]_  = \new_[37956]_  & \new_[37943]_ ;
  assign \new_[1849]_  = \new_[37932]_  & \new_[37919]_ ;
  assign \new_[1850]_  = \new_[37908]_  & \new_[37895]_ ;
  assign \new_[1851]_  = \new_[37884]_  & \new_[37871]_ ;
  assign \new_[1852]_  = \new_[37860]_  & \new_[37847]_ ;
  assign \new_[1853]_  = \new_[37836]_  & \new_[37823]_ ;
  assign \new_[1854]_  = \new_[37812]_  & \new_[37799]_ ;
  assign \new_[1855]_  = \new_[37788]_  & \new_[37775]_ ;
  assign \new_[1856]_  = \new_[37764]_  & \new_[37751]_ ;
  assign \new_[1857]_  = \new_[37740]_  & \new_[37727]_ ;
  assign \new_[1858]_  = \new_[37716]_  & \new_[37703]_ ;
  assign \new_[1859]_  = \new_[37692]_  & \new_[37679]_ ;
  assign \new_[1860]_  = \new_[37668]_  & \new_[37655]_ ;
  assign \new_[1861]_  = \new_[37644]_  & \new_[37631]_ ;
  assign \new_[1862]_  = \new_[37620]_  & \new_[37607]_ ;
  assign \new_[1863]_  = \new_[37596]_  & \new_[37583]_ ;
  assign \new_[1864]_  = \new_[37572]_  & \new_[37559]_ ;
  assign \new_[1865]_  = \new_[37548]_  & \new_[37535]_ ;
  assign \new_[1866]_  = \new_[37524]_  & \new_[37511]_ ;
  assign \new_[1867]_  = \new_[37500]_  & \new_[37487]_ ;
  assign \new_[1868]_  = \new_[37476]_  & \new_[37463]_ ;
  assign \new_[1869]_  = \new_[37452]_  & \new_[37439]_ ;
  assign \new_[1870]_  = \new_[37428]_  & \new_[37415]_ ;
  assign \new_[1871]_  = \new_[37404]_  & \new_[37391]_ ;
  assign \new_[1872]_  = \new_[37380]_  & \new_[37367]_ ;
  assign \new_[1873]_  = \new_[37356]_  & \new_[37343]_ ;
  assign \new_[1874]_  = \new_[37332]_  & \new_[37319]_ ;
  assign \new_[1875]_  = \new_[37308]_  & \new_[37295]_ ;
  assign \new_[1876]_  = \new_[37284]_  & \new_[37271]_ ;
  assign \new_[1877]_  = \new_[37260]_  & \new_[37247]_ ;
  assign \new_[1878]_  = \new_[37236]_  & \new_[37223]_ ;
  assign \new_[1879]_  = \new_[37212]_  & \new_[37199]_ ;
  assign \new_[1880]_  = \new_[37188]_  & \new_[37175]_ ;
  assign \new_[1881]_  = \new_[37164]_  & \new_[37151]_ ;
  assign \new_[1882]_  = \new_[37140]_  & \new_[37127]_ ;
  assign \new_[1883]_  = \new_[37116]_  & \new_[37103]_ ;
  assign \new_[1884]_  = \new_[37092]_  & \new_[37079]_ ;
  assign \new_[1885]_  = \new_[37068]_  & \new_[37055]_ ;
  assign \new_[1886]_  = \new_[37044]_  & \new_[37031]_ ;
  assign \new_[1887]_  = \new_[37020]_  & \new_[37007]_ ;
  assign \new_[1888]_  = \new_[36996]_  & \new_[36983]_ ;
  assign \new_[1889]_  = \new_[36972]_  & \new_[36959]_ ;
  assign \new_[1890]_  = \new_[36948]_  & \new_[36935]_ ;
  assign \new_[1891]_  = \new_[36924]_  & \new_[36911]_ ;
  assign \new_[1892]_  = \new_[36900]_  & \new_[36887]_ ;
  assign \new_[1893]_  = \new_[36876]_  & \new_[36863]_ ;
  assign \new_[1894]_  = \new_[36852]_  & \new_[36839]_ ;
  assign \new_[1895]_  = \new_[36828]_  & \new_[36815]_ ;
  assign \new_[1896]_  = \new_[36804]_  & \new_[36791]_ ;
  assign \new_[1897]_  = \new_[36780]_  & \new_[36767]_ ;
  assign \new_[1898]_  = \new_[36756]_  & \new_[36743]_ ;
  assign \new_[1899]_  = \new_[36732]_  & \new_[36719]_ ;
  assign \new_[1900]_  = \new_[36708]_  & \new_[36695]_ ;
  assign \new_[1901]_  = \new_[36684]_  & \new_[36671]_ ;
  assign \new_[1902]_  = \new_[36660]_  & \new_[36647]_ ;
  assign \new_[1903]_  = \new_[36636]_  & \new_[36623]_ ;
  assign \new_[1904]_  = \new_[36612]_  & \new_[36599]_ ;
  assign \new_[1905]_  = \new_[36588]_  & \new_[36575]_ ;
  assign \new_[1906]_  = \new_[36564]_  & \new_[36551]_ ;
  assign \new_[1907]_  = \new_[36540]_  & \new_[36527]_ ;
  assign \new_[1908]_  = \new_[36516]_  & \new_[36503]_ ;
  assign \new_[1909]_  = \new_[36492]_  & \new_[36479]_ ;
  assign \new_[1910]_  = \new_[36468]_  & \new_[36455]_ ;
  assign \new_[1911]_  = \new_[36444]_  & \new_[36431]_ ;
  assign \new_[1912]_  = \new_[36420]_  & \new_[36407]_ ;
  assign \new_[1913]_  = \new_[36396]_  & \new_[36383]_ ;
  assign \new_[1914]_  = \new_[36372]_  & \new_[36359]_ ;
  assign \new_[1915]_  = \new_[36348]_  & \new_[36335]_ ;
  assign \new_[1916]_  = \new_[36324]_  & \new_[36311]_ ;
  assign \new_[1917]_  = \new_[36300]_  & \new_[36287]_ ;
  assign \new_[1918]_  = \new_[36276]_  & \new_[36263]_ ;
  assign \new_[1919]_  = \new_[36252]_  & \new_[36239]_ ;
  assign \new_[1920]_  = \new_[36228]_  & \new_[36215]_ ;
  assign \new_[1921]_  = \new_[36204]_  & \new_[36191]_ ;
  assign \new_[1922]_  = \new_[36180]_  & \new_[36167]_ ;
  assign \new_[1923]_  = \new_[36156]_  & \new_[36143]_ ;
  assign \new_[1924]_  = \new_[36132]_  & \new_[36119]_ ;
  assign \new_[1925]_  = \new_[36108]_  & \new_[36095]_ ;
  assign \new_[1926]_  = \new_[36084]_  & \new_[36071]_ ;
  assign \new_[1927]_  = \new_[36060]_  & \new_[36047]_ ;
  assign \new_[1928]_  = \new_[36036]_  & \new_[36023]_ ;
  assign \new_[1929]_  = \new_[36012]_  & \new_[35999]_ ;
  assign \new_[1930]_  = \new_[35988]_  & \new_[35975]_ ;
  assign \new_[1931]_  = \new_[35964]_  & \new_[35951]_ ;
  assign \new_[1932]_  = \new_[35940]_  & \new_[35927]_ ;
  assign \new_[1933]_  = \new_[35916]_  & \new_[35903]_ ;
  assign \new_[1934]_  = \new_[35892]_  & \new_[35879]_ ;
  assign \new_[1935]_  = \new_[35868]_  & \new_[35855]_ ;
  assign \new_[1936]_  = \new_[35844]_  & \new_[35831]_ ;
  assign \new_[1937]_  = \new_[35820]_  & \new_[35807]_ ;
  assign \new_[1938]_  = \new_[35796]_  & \new_[35783]_ ;
  assign \new_[1939]_  = \new_[35772]_  & \new_[35759]_ ;
  assign \new_[1940]_  = \new_[35748]_  & \new_[35735]_ ;
  assign \new_[1941]_  = \new_[35724]_  & \new_[35711]_ ;
  assign \new_[1942]_  = \new_[35700]_  & \new_[35687]_ ;
  assign \new_[1943]_  = \new_[35676]_  & \new_[35663]_ ;
  assign \new_[1944]_  = \new_[35652]_  & \new_[35639]_ ;
  assign \new_[1945]_  = \new_[35628]_  & \new_[35615]_ ;
  assign \new_[1946]_  = \new_[35604]_  & \new_[35591]_ ;
  assign \new_[1947]_  = \new_[35580]_  & \new_[35567]_ ;
  assign \new_[1948]_  = \new_[35556]_  & \new_[35543]_ ;
  assign \new_[1949]_  = \new_[35532]_  & \new_[35519]_ ;
  assign \new_[1950]_  = \new_[35508]_  & \new_[35495]_ ;
  assign \new_[1951]_  = \new_[35484]_  & \new_[35471]_ ;
  assign \new_[1952]_  = \new_[35460]_  & \new_[35447]_ ;
  assign \new_[1953]_  = \new_[35436]_  & \new_[35423]_ ;
  assign \new_[1954]_  = \new_[35412]_  & \new_[35399]_ ;
  assign \new_[1955]_  = \new_[35388]_  & \new_[35375]_ ;
  assign \new_[1956]_  = \new_[35364]_  & \new_[35351]_ ;
  assign \new_[1957]_  = \new_[35340]_  & \new_[35327]_ ;
  assign \new_[1958]_  = \new_[35316]_  & \new_[35303]_ ;
  assign \new_[1959]_  = \new_[35292]_  & \new_[35279]_ ;
  assign \new_[1960]_  = \new_[35268]_  & \new_[35255]_ ;
  assign \new_[1961]_  = \new_[35244]_  & \new_[35231]_ ;
  assign \new_[1962]_  = \new_[35220]_  & \new_[35207]_ ;
  assign \new_[1963]_  = \new_[35196]_  & \new_[35183]_ ;
  assign \new_[1964]_  = \new_[35172]_  & \new_[35159]_ ;
  assign \new_[1965]_  = \new_[35148]_  & \new_[35135]_ ;
  assign \new_[1966]_  = \new_[35124]_  & \new_[35111]_ ;
  assign \new_[1967]_  = \new_[35100]_  & \new_[35087]_ ;
  assign \new_[1968]_  = \new_[35076]_  & \new_[35063]_ ;
  assign \new_[1969]_  = \new_[35052]_  & \new_[35039]_ ;
  assign \new_[1970]_  = \new_[35028]_  & \new_[35015]_ ;
  assign \new_[1971]_  = \new_[35004]_  & \new_[34991]_ ;
  assign \new_[1972]_  = \new_[34980]_  & \new_[34967]_ ;
  assign \new_[1973]_  = \new_[34956]_  & \new_[34943]_ ;
  assign \new_[1974]_  = \new_[34932]_  & \new_[34919]_ ;
  assign \new_[1975]_  = \new_[34908]_  & \new_[34895]_ ;
  assign \new_[1976]_  = \new_[34884]_  & \new_[34871]_ ;
  assign \new_[1977]_  = \new_[34860]_  & \new_[34847]_ ;
  assign \new_[1978]_  = \new_[34836]_  & \new_[34823]_ ;
  assign \new_[1979]_  = \new_[34812]_  & \new_[34799]_ ;
  assign \new_[1980]_  = \new_[34788]_  & \new_[34775]_ ;
  assign \new_[1981]_  = \new_[34764]_  & \new_[34751]_ ;
  assign \new_[1982]_  = \new_[34740]_  & \new_[34727]_ ;
  assign \new_[1983]_  = \new_[34716]_  & \new_[34703]_ ;
  assign \new_[1984]_  = \new_[34692]_  & \new_[34679]_ ;
  assign \new_[1985]_  = \new_[34668]_  & \new_[34655]_ ;
  assign \new_[1986]_  = \new_[34644]_  & \new_[34631]_ ;
  assign \new_[1987]_  = \new_[34620]_  & \new_[34607]_ ;
  assign \new_[1988]_  = \new_[34596]_  & \new_[34583]_ ;
  assign \new_[1989]_  = \new_[34572]_  & \new_[34559]_ ;
  assign \new_[1990]_  = \new_[34548]_  & \new_[34535]_ ;
  assign \new_[1991]_  = \new_[34524]_  & \new_[34511]_ ;
  assign \new_[1992]_  = \new_[34500]_  & \new_[34487]_ ;
  assign \new_[1993]_  = \new_[34476]_  & \new_[34463]_ ;
  assign \new_[1994]_  = \new_[34452]_  & \new_[34439]_ ;
  assign \new_[1995]_  = \new_[34428]_  & \new_[34415]_ ;
  assign \new_[1996]_  = \new_[34404]_  & \new_[34391]_ ;
  assign \new_[1997]_  = \new_[34380]_  & \new_[34367]_ ;
  assign \new_[1998]_  = \new_[34356]_  & \new_[34343]_ ;
  assign \new_[1999]_  = \new_[34332]_  & \new_[34319]_ ;
  assign \new_[2000]_  = \new_[34308]_  & \new_[34295]_ ;
  assign \new_[2001]_  = \new_[34284]_  & \new_[34271]_ ;
  assign \new_[2002]_  = \new_[34260]_  & \new_[34247]_ ;
  assign \new_[2003]_  = \new_[34236]_  & \new_[34223]_ ;
  assign \new_[2004]_  = \new_[34212]_  & \new_[34199]_ ;
  assign \new_[2005]_  = \new_[34188]_  & \new_[34175]_ ;
  assign \new_[2006]_  = \new_[34164]_  & \new_[34151]_ ;
  assign \new_[2007]_  = \new_[34140]_  & \new_[34127]_ ;
  assign \new_[2008]_  = \new_[34116]_  & \new_[34103]_ ;
  assign \new_[2009]_  = \new_[34092]_  & \new_[34079]_ ;
  assign \new_[2010]_  = \new_[34068]_  & \new_[34055]_ ;
  assign \new_[2011]_  = \new_[34044]_  & \new_[34031]_ ;
  assign \new_[2012]_  = \new_[34020]_  & \new_[34007]_ ;
  assign \new_[2013]_  = \new_[33996]_  & \new_[33983]_ ;
  assign \new_[2014]_  = \new_[33972]_  & \new_[33959]_ ;
  assign \new_[2015]_  = \new_[33948]_  & \new_[33935]_ ;
  assign \new_[2016]_  = \new_[33924]_  & \new_[33911]_ ;
  assign \new_[2017]_  = \new_[33900]_  & \new_[33887]_ ;
  assign \new_[2018]_  = \new_[33876]_  & \new_[33863]_ ;
  assign \new_[2019]_  = \new_[33852]_  & \new_[33839]_ ;
  assign \new_[2020]_  = \new_[33828]_  & \new_[33815]_ ;
  assign \new_[2021]_  = \new_[33804]_  & \new_[33791]_ ;
  assign \new_[2022]_  = \new_[33780]_  & \new_[33767]_ ;
  assign \new_[2023]_  = \new_[33756]_  & \new_[33743]_ ;
  assign \new_[2024]_  = \new_[33732]_  & \new_[33719]_ ;
  assign \new_[2025]_  = \new_[33708]_  & \new_[33695]_ ;
  assign \new_[2026]_  = \new_[33684]_  & \new_[33671]_ ;
  assign \new_[2027]_  = \new_[33660]_  & \new_[33647]_ ;
  assign \new_[2028]_  = \new_[33636]_  & \new_[33623]_ ;
  assign \new_[2029]_  = \new_[33612]_  & \new_[33599]_ ;
  assign \new_[2030]_  = \new_[33588]_  & \new_[33575]_ ;
  assign \new_[2031]_  = \new_[33564]_  & \new_[33551]_ ;
  assign \new_[2032]_  = \new_[33540]_  & \new_[33527]_ ;
  assign \new_[2033]_  = \new_[33516]_  & \new_[33503]_ ;
  assign \new_[2034]_  = \new_[33492]_  & \new_[33479]_ ;
  assign \new_[2035]_  = \new_[33468]_  & \new_[33455]_ ;
  assign \new_[2036]_  = \new_[33444]_  & \new_[33431]_ ;
  assign \new_[2037]_  = \new_[33420]_  & \new_[33407]_ ;
  assign \new_[2038]_  = \new_[33396]_  & \new_[33383]_ ;
  assign \new_[2039]_  = \new_[33372]_  & \new_[33359]_ ;
  assign \new_[2040]_  = \new_[33348]_  & \new_[33335]_ ;
  assign \new_[2041]_  = \new_[33324]_  & \new_[33311]_ ;
  assign \new_[2042]_  = \new_[33300]_  & \new_[33287]_ ;
  assign \new_[2043]_  = \new_[33276]_  & \new_[33263]_ ;
  assign \new_[2044]_  = \new_[33252]_  & \new_[33239]_ ;
  assign \new_[2045]_  = \new_[33228]_  & \new_[33215]_ ;
  assign \new_[2046]_  = \new_[33204]_  & \new_[33191]_ ;
  assign \new_[2047]_  = \new_[33180]_  & \new_[33167]_ ;
  assign \new_[2048]_  = \new_[33156]_  & \new_[33143]_ ;
  assign \new_[2049]_  = \new_[33132]_  & \new_[33119]_ ;
  assign \new_[2050]_  = \new_[33108]_  & \new_[33095]_ ;
  assign \new_[2051]_  = \new_[33084]_  & \new_[33071]_ ;
  assign \new_[2052]_  = \new_[33060]_  & \new_[33047]_ ;
  assign \new_[2053]_  = \new_[33036]_  & \new_[33023]_ ;
  assign \new_[2054]_  = \new_[33012]_  & \new_[32999]_ ;
  assign \new_[2055]_  = \new_[32988]_  & \new_[32975]_ ;
  assign \new_[2056]_  = \new_[32964]_  & \new_[32951]_ ;
  assign \new_[2057]_  = \new_[32940]_  & \new_[32927]_ ;
  assign \new_[2058]_  = \new_[32916]_  & \new_[32903]_ ;
  assign \new_[2059]_  = \new_[32892]_  & \new_[32879]_ ;
  assign \new_[2060]_  = \new_[32868]_  & \new_[32855]_ ;
  assign \new_[2061]_  = \new_[32844]_  & \new_[32831]_ ;
  assign \new_[2062]_  = \new_[32820]_  & \new_[32807]_ ;
  assign \new_[2063]_  = \new_[32796]_  & \new_[32783]_ ;
  assign \new_[2064]_  = \new_[32772]_  & \new_[32759]_ ;
  assign \new_[2065]_  = \new_[32748]_  & \new_[32735]_ ;
  assign \new_[2066]_  = \new_[32724]_  & \new_[32711]_ ;
  assign \new_[2067]_  = \new_[32700]_  & \new_[32687]_ ;
  assign \new_[2068]_  = \new_[32676]_  & \new_[32663]_ ;
  assign \new_[2069]_  = \new_[32652]_  & \new_[32639]_ ;
  assign \new_[2070]_  = \new_[32628]_  & \new_[32615]_ ;
  assign \new_[2071]_  = \new_[32604]_  & \new_[32591]_ ;
  assign \new_[2072]_  = \new_[32580]_  & \new_[32567]_ ;
  assign \new_[2073]_  = \new_[32556]_  & \new_[32543]_ ;
  assign \new_[2074]_  = \new_[32532]_  & \new_[32519]_ ;
  assign \new_[2075]_  = \new_[32508]_  & \new_[32495]_ ;
  assign \new_[2076]_  = \new_[32484]_  & \new_[32471]_ ;
  assign \new_[2077]_  = \new_[32460]_  & \new_[32447]_ ;
  assign \new_[2078]_  = \new_[32436]_  & \new_[32423]_ ;
  assign \new_[2079]_  = \new_[32412]_  & \new_[32399]_ ;
  assign \new_[2080]_  = \new_[32388]_  & \new_[32375]_ ;
  assign \new_[2081]_  = \new_[32364]_  & \new_[32351]_ ;
  assign \new_[2082]_  = \new_[32340]_  & \new_[32327]_ ;
  assign \new_[2083]_  = \new_[32316]_  & \new_[32303]_ ;
  assign \new_[2084]_  = \new_[32292]_  & \new_[32279]_ ;
  assign \new_[2085]_  = \new_[32268]_  & \new_[32255]_ ;
  assign \new_[2086]_  = \new_[32244]_  & \new_[32231]_ ;
  assign \new_[2087]_  = \new_[32220]_  & \new_[32207]_ ;
  assign \new_[2088]_  = \new_[32196]_  & \new_[32183]_ ;
  assign \new_[2089]_  = \new_[32172]_  & \new_[32159]_ ;
  assign \new_[2090]_  = \new_[32148]_  & \new_[32135]_ ;
  assign \new_[2091]_  = \new_[32124]_  & \new_[32111]_ ;
  assign \new_[2092]_  = \new_[32100]_  & \new_[32087]_ ;
  assign \new_[2093]_  = \new_[32076]_  & \new_[32063]_ ;
  assign \new_[2094]_  = \new_[32052]_  & \new_[32039]_ ;
  assign \new_[2095]_  = \new_[32028]_  & \new_[32015]_ ;
  assign \new_[2096]_  = \new_[32004]_  & \new_[31991]_ ;
  assign \new_[2097]_  = \new_[31980]_  & \new_[31967]_ ;
  assign \new_[2098]_  = \new_[31956]_  & \new_[31943]_ ;
  assign \new_[2099]_  = \new_[31932]_  & \new_[31919]_ ;
  assign \new_[2100]_  = \new_[31908]_  & \new_[31895]_ ;
  assign \new_[2101]_  = \new_[31884]_  & \new_[31871]_ ;
  assign \new_[2102]_  = \new_[31860]_  & \new_[31847]_ ;
  assign \new_[2103]_  = \new_[31836]_  & \new_[31823]_ ;
  assign \new_[2104]_  = \new_[31812]_  & \new_[31799]_ ;
  assign \new_[2105]_  = \new_[31788]_  & \new_[31775]_ ;
  assign \new_[2106]_  = \new_[31764]_  & \new_[31751]_ ;
  assign \new_[2107]_  = \new_[31740]_  & \new_[31727]_ ;
  assign \new_[2108]_  = \new_[31716]_  & \new_[31703]_ ;
  assign \new_[2109]_  = \new_[31692]_  & \new_[31679]_ ;
  assign \new_[2110]_  = \new_[31668]_  & \new_[31655]_ ;
  assign \new_[2111]_  = \new_[31644]_  & \new_[31631]_ ;
  assign \new_[2112]_  = \new_[31620]_  & \new_[31607]_ ;
  assign \new_[2113]_  = \new_[31596]_  & \new_[31583]_ ;
  assign \new_[2114]_  = \new_[31572]_  & \new_[31559]_ ;
  assign \new_[2115]_  = \new_[31548]_  & \new_[31535]_ ;
  assign \new_[2116]_  = \new_[31524]_  & \new_[31511]_ ;
  assign \new_[2117]_  = \new_[31500]_  & \new_[31487]_ ;
  assign \new_[2118]_  = \new_[31476]_  & \new_[31463]_ ;
  assign \new_[2119]_  = \new_[31452]_  & \new_[31439]_ ;
  assign \new_[2120]_  = \new_[31428]_  & \new_[31415]_ ;
  assign \new_[2121]_  = \new_[31404]_  & \new_[31391]_ ;
  assign \new_[2122]_  = \new_[31380]_  & \new_[31367]_ ;
  assign \new_[2123]_  = \new_[31356]_  & \new_[31343]_ ;
  assign \new_[2124]_  = \new_[31332]_  & \new_[31319]_ ;
  assign \new_[2125]_  = \new_[31308]_  & \new_[31295]_ ;
  assign \new_[2126]_  = \new_[31284]_  & \new_[31271]_ ;
  assign \new_[2127]_  = \new_[31260]_  & \new_[31247]_ ;
  assign \new_[2128]_  = \new_[31236]_  & \new_[31223]_ ;
  assign \new_[2129]_  = \new_[31212]_  & \new_[31199]_ ;
  assign \new_[2130]_  = \new_[31188]_  & \new_[31175]_ ;
  assign \new_[2131]_  = \new_[31164]_  & \new_[31151]_ ;
  assign \new_[2132]_  = \new_[31140]_  & \new_[31127]_ ;
  assign \new_[2133]_  = \new_[31116]_  & \new_[31103]_ ;
  assign \new_[2134]_  = \new_[31092]_  & \new_[31079]_ ;
  assign \new_[2135]_  = \new_[31068]_  & \new_[31055]_ ;
  assign \new_[2136]_  = \new_[31044]_  & \new_[31031]_ ;
  assign \new_[2137]_  = \new_[31020]_  & \new_[31007]_ ;
  assign \new_[2138]_  = \new_[30996]_  & \new_[30983]_ ;
  assign \new_[2139]_  = \new_[30972]_  & \new_[30959]_ ;
  assign \new_[2140]_  = \new_[30948]_  & \new_[30935]_ ;
  assign \new_[2141]_  = \new_[30924]_  & \new_[30911]_ ;
  assign \new_[2142]_  = \new_[30900]_  & \new_[30887]_ ;
  assign \new_[2143]_  = \new_[30876]_  & \new_[30863]_ ;
  assign \new_[2144]_  = \new_[30852]_  & \new_[30839]_ ;
  assign \new_[2145]_  = \new_[30828]_  & \new_[30815]_ ;
  assign \new_[2146]_  = \new_[30804]_  & \new_[30791]_ ;
  assign \new_[2147]_  = \new_[30780]_  & \new_[30767]_ ;
  assign \new_[2148]_  = \new_[30756]_  & \new_[30743]_ ;
  assign \new_[2149]_  = \new_[30732]_  & \new_[30719]_ ;
  assign \new_[2150]_  = \new_[30708]_  & \new_[30695]_ ;
  assign \new_[2151]_  = \new_[30684]_  & \new_[30671]_ ;
  assign \new_[2152]_  = \new_[30660]_  & \new_[30647]_ ;
  assign \new_[2153]_  = \new_[30636]_  & \new_[30623]_ ;
  assign \new_[2154]_  = \new_[30612]_  & \new_[30599]_ ;
  assign \new_[2155]_  = \new_[30588]_  & \new_[30575]_ ;
  assign \new_[2156]_  = \new_[30564]_  & \new_[30551]_ ;
  assign \new_[2157]_  = \new_[30540]_  & \new_[30527]_ ;
  assign \new_[2158]_  = \new_[30516]_  & \new_[30503]_ ;
  assign \new_[2159]_  = \new_[30492]_  & \new_[30479]_ ;
  assign \new_[2160]_  = \new_[30468]_  & \new_[30455]_ ;
  assign \new_[2161]_  = \new_[30444]_  & \new_[30431]_ ;
  assign \new_[2162]_  = \new_[30420]_  & \new_[30407]_ ;
  assign \new_[2163]_  = \new_[30396]_  & \new_[30383]_ ;
  assign \new_[2164]_  = \new_[30372]_  & \new_[30359]_ ;
  assign \new_[2165]_  = \new_[30348]_  & \new_[30335]_ ;
  assign \new_[2166]_  = \new_[30324]_  & \new_[30311]_ ;
  assign \new_[2167]_  = \new_[30300]_  & \new_[30287]_ ;
  assign \new_[2168]_  = \new_[30276]_  & \new_[30263]_ ;
  assign \new_[2169]_  = \new_[30252]_  & \new_[30239]_ ;
  assign \new_[2170]_  = \new_[30228]_  & \new_[30215]_ ;
  assign \new_[2171]_  = \new_[30204]_  & \new_[30191]_ ;
  assign \new_[2172]_  = \new_[30180]_  & \new_[30167]_ ;
  assign \new_[2173]_  = \new_[30156]_  & \new_[30143]_ ;
  assign \new_[2174]_  = \new_[30132]_  & \new_[30119]_ ;
  assign \new_[2175]_  = \new_[30108]_  & \new_[30095]_ ;
  assign \new_[2176]_  = \new_[30084]_  & \new_[30071]_ ;
  assign \new_[2177]_  = \new_[30060]_  & \new_[30047]_ ;
  assign \new_[2178]_  = \new_[30036]_  & \new_[30023]_ ;
  assign \new_[2179]_  = \new_[30012]_  & \new_[29999]_ ;
  assign \new_[2180]_  = \new_[29988]_  & \new_[29975]_ ;
  assign \new_[2181]_  = \new_[29964]_  & \new_[29951]_ ;
  assign \new_[2182]_  = \new_[29940]_  & \new_[29927]_ ;
  assign \new_[2183]_  = \new_[29916]_  & \new_[29903]_ ;
  assign \new_[2184]_  = \new_[29892]_  & \new_[29879]_ ;
  assign \new_[2185]_  = \new_[29868]_  & \new_[29855]_ ;
  assign \new_[2186]_  = \new_[29844]_  & \new_[29831]_ ;
  assign \new_[2187]_  = \new_[29820]_  & \new_[29807]_ ;
  assign \new_[2188]_  = \new_[29796]_  & \new_[29783]_ ;
  assign \new_[2189]_  = \new_[29772]_  & \new_[29759]_ ;
  assign \new_[2190]_  = \new_[29748]_  & \new_[29735]_ ;
  assign \new_[2191]_  = \new_[29724]_  & \new_[29711]_ ;
  assign \new_[2192]_  = \new_[29700]_  & \new_[29687]_ ;
  assign \new_[2193]_  = \new_[29676]_  & \new_[29663]_ ;
  assign \new_[2194]_  = \new_[29652]_  & \new_[29639]_ ;
  assign \new_[2195]_  = \new_[29628]_  & \new_[29615]_ ;
  assign \new_[2196]_  = \new_[29604]_  & \new_[29591]_ ;
  assign \new_[2197]_  = \new_[29580]_  & \new_[29567]_ ;
  assign \new_[2198]_  = \new_[29556]_  & \new_[29543]_ ;
  assign \new_[2199]_  = \new_[29532]_  & \new_[29519]_ ;
  assign \new_[2200]_  = \new_[29508]_  & \new_[29495]_ ;
  assign \new_[2201]_  = \new_[29484]_  & \new_[29473]_ ;
  assign \new_[2202]_  = \new_[29462]_  & \new_[29451]_ ;
  assign \new_[2203]_  = \new_[29440]_  & \new_[29429]_ ;
  assign \new_[2204]_  = \new_[29418]_  & \new_[29407]_ ;
  assign \new_[2205]_  = \new_[29396]_  & \new_[29385]_ ;
  assign \new_[2206]_  = \new_[29374]_  & \new_[29363]_ ;
  assign \new_[2207]_  = \new_[29352]_  & \new_[29341]_ ;
  assign \new_[2208]_  = \new_[29330]_  & \new_[29319]_ ;
  assign \new_[2209]_  = \new_[29308]_  & \new_[29297]_ ;
  assign \new_[2210]_  = \new_[29286]_  & \new_[29275]_ ;
  assign \new_[2211]_  = \new_[29264]_  & \new_[29253]_ ;
  assign \new_[2212]_  = \new_[29242]_  & \new_[29231]_ ;
  assign \new_[2213]_  = \new_[29220]_  & \new_[29209]_ ;
  assign \new_[2214]_  = \new_[29198]_  & \new_[29187]_ ;
  assign \new_[2215]_  = \new_[29176]_  & \new_[29165]_ ;
  assign \new_[2216]_  = \new_[29154]_  & \new_[29143]_ ;
  assign \new_[2217]_  = \new_[29132]_  & \new_[29121]_ ;
  assign \new_[2218]_  = \new_[29110]_  & \new_[29099]_ ;
  assign \new_[2219]_  = \new_[29088]_  & \new_[29077]_ ;
  assign \new_[2220]_  = \new_[29066]_  & \new_[29055]_ ;
  assign \new_[2221]_  = \new_[29044]_  & \new_[29033]_ ;
  assign \new_[2222]_  = \new_[29022]_  & \new_[29011]_ ;
  assign \new_[2223]_  = \new_[29000]_  & \new_[28989]_ ;
  assign \new_[2224]_  = \new_[28978]_  & \new_[28967]_ ;
  assign \new_[2225]_  = \new_[28956]_  & \new_[28945]_ ;
  assign \new_[2226]_  = \new_[28934]_  & \new_[28923]_ ;
  assign \new_[2227]_  = \new_[28912]_  & \new_[28901]_ ;
  assign \new_[2228]_  = \new_[28890]_  & \new_[28879]_ ;
  assign \new_[2229]_  = \new_[28868]_  & \new_[28857]_ ;
  assign \new_[2230]_  = \new_[28846]_  & \new_[28835]_ ;
  assign \new_[2231]_  = \new_[28824]_  & \new_[28813]_ ;
  assign \new_[2232]_  = \new_[28802]_  & \new_[28791]_ ;
  assign \new_[2233]_  = \new_[28780]_  & \new_[28769]_ ;
  assign \new_[2234]_  = \new_[28758]_  & \new_[28747]_ ;
  assign \new_[2235]_  = \new_[28736]_  & \new_[28725]_ ;
  assign \new_[2236]_  = \new_[28714]_  & \new_[28703]_ ;
  assign \new_[2237]_  = \new_[28692]_  & \new_[28681]_ ;
  assign \new_[2238]_  = \new_[28670]_  & \new_[28659]_ ;
  assign \new_[2239]_  = \new_[28648]_  & \new_[28637]_ ;
  assign \new_[2240]_  = \new_[28626]_  & \new_[28615]_ ;
  assign \new_[2241]_  = \new_[28604]_  & \new_[28593]_ ;
  assign \new_[2242]_  = \new_[28582]_  & \new_[28571]_ ;
  assign \new_[2243]_  = \new_[28560]_  & \new_[28549]_ ;
  assign \new_[2244]_  = \new_[28538]_  & \new_[28527]_ ;
  assign \new_[2245]_  = \new_[28516]_  & \new_[28505]_ ;
  assign \new_[2246]_  = \new_[28494]_  & \new_[28483]_ ;
  assign \new_[2247]_  = \new_[28472]_  & \new_[28461]_ ;
  assign \new_[2248]_  = \new_[28450]_  & \new_[28439]_ ;
  assign \new_[2249]_  = \new_[28428]_  & \new_[28417]_ ;
  assign \new_[2250]_  = \new_[28406]_  & \new_[28395]_ ;
  assign \new_[2251]_  = \new_[28384]_  & \new_[28373]_ ;
  assign \new_[2252]_  = \new_[28362]_  & \new_[28351]_ ;
  assign \new_[2253]_  = \new_[28340]_  & \new_[28329]_ ;
  assign \new_[2254]_  = \new_[28318]_  & \new_[28307]_ ;
  assign \new_[2255]_  = \new_[28296]_  & \new_[28285]_ ;
  assign \new_[2256]_  = \new_[28274]_  & \new_[28263]_ ;
  assign \new_[2257]_  = \new_[28252]_  & \new_[28241]_ ;
  assign \new_[2258]_  = \new_[28230]_  & \new_[28219]_ ;
  assign \new_[2259]_  = \new_[28208]_  & \new_[28197]_ ;
  assign \new_[2260]_  = \new_[28186]_  & \new_[28175]_ ;
  assign \new_[2261]_  = \new_[28164]_  & \new_[28153]_ ;
  assign \new_[2262]_  = \new_[28142]_  & \new_[28131]_ ;
  assign \new_[2263]_  = \new_[28120]_  & \new_[28109]_ ;
  assign \new_[2264]_  = \new_[28098]_  & \new_[28087]_ ;
  assign \new_[2265]_  = \new_[28076]_  & \new_[28065]_ ;
  assign \new_[2266]_  = \new_[28054]_  & \new_[28043]_ ;
  assign \new_[2267]_  = \new_[28032]_  & \new_[28021]_ ;
  assign \new_[2268]_  = \new_[28010]_  & \new_[27999]_ ;
  assign \new_[2269]_  = \new_[27988]_  & \new_[27977]_ ;
  assign \new_[2270]_  = \new_[27966]_  & \new_[27955]_ ;
  assign \new_[2271]_  = \new_[27944]_  & \new_[27933]_ ;
  assign \new_[2272]_  = \new_[27922]_  & \new_[27911]_ ;
  assign \new_[2273]_  = \new_[27900]_  & \new_[27889]_ ;
  assign \new_[2274]_  = \new_[27878]_  & \new_[27867]_ ;
  assign \new_[2275]_  = \new_[27856]_  & \new_[27845]_ ;
  assign \new_[2276]_  = \new_[27834]_  & \new_[27823]_ ;
  assign \new_[2277]_  = \new_[27812]_  & \new_[27801]_ ;
  assign \new_[2278]_  = \new_[27790]_  & \new_[27779]_ ;
  assign \new_[2279]_  = \new_[27768]_  & \new_[27757]_ ;
  assign \new_[2280]_  = \new_[27746]_  & \new_[27735]_ ;
  assign \new_[2281]_  = \new_[27724]_  & \new_[27713]_ ;
  assign \new_[2282]_  = \new_[27702]_  & \new_[27691]_ ;
  assign \new_[2283]_  = \new_[27680]_  & \new_[27669]_ ;
  assign \new_[2284]_  = \new_[27658]_  & \new_[27647]_ ;
  assign \new_[2285]_  = \new_[27636]_  & \new_[27625]_ ;
  assign \new_[2286]_  = \new_[27614]_  & \new_[27603]_ ;
  assign \new_[2287]_  = \new_[27592]_  & \new_[27581]_ ;
  assign \new_[2288]_  = \new_[27570]_  & \new_[27559]_ ;
  assign \new_[2289]_  = \new_[27548]_  & \new_[27537]_ ;
  assign \new_[2290]_  = \new_[27526]_  & \new_[27515]_ ;
  assign \new_[2291]_  = \new_[27504]_  & \new_[27493]_ ;
  assign \new_[2292]_  = \new_[27482]_  & \new_[27471]_ ;
  assign \new_[2293]_  = \new_[27460]_  & \new_[27449]_ ;
  assign \new_[2294]_  = \new_[27438]_  & \new_[27427]_ ;
  assign \new_[2295]_  = \new_[27416]_  & \new_[27405]_ ;
  assign \new_[2296]_  = \new_[27394]_  & \new_[27383]_ ;
  assign \new_[2297]_  = \new_[27372]_  & \new_[27361]_ ;
  assign \new_[2298]_  = \new_[27350]_  & \new_[27339]_ ;
  assign \new_[2299]_  = \new_[27328]_  & \new_[27317]_ ;
  assign \new_[2300]_  = \new_[27306]_  & \new_[27295]_ ;
  assign \new_[2301]_  = \new_[27284]_  & \new_[27273]_ ;
  assign \new_[2302]_  = \new_[27262]_  & \new_[27251]_ ;
  assign \new_[2303]_  = \new_[27240]_  & \new_[27229]_ ;
  assign \new_[2304]_  = \new_[27218]_  & \new_[27207]_ ;
  assign \new_[2305]_  = \new_[27196]_  & \new_[27185]_ ;
  assign \new_[2306]_  = \new_[27174]_  & \new_[27163]_ ;
  assign \new_[2307]_  = \new_[27152]_  & \new_[27141]_ ;
  assign \new_[2308]_  = \new_[27130]_  & \new_[27119]_ ;
  assign \new_[2309]_  = \new_[27108]_  & \new_[27097]_ ;
  assign \new_[2310]_  = \new_[27086]_  & \new_[27075]_ ;
  assign \new_[2311]_  = \new_[27064]_  & \new_[27053]_ ;
  assign \new_[2312]_  = \new_[27042]_  & \new_[27031]_ ;
  assign \new_[2313]_  = \new_[27020]_  & \new_[27009]_ ;
  assign \new_[2314]_  = \new_[26998]_  & \new_[26987]_ ;
  assign \new_[2315]_  = \new_[26976]_  & \new_[26965]_ ;
  assign \new_[2316]_  = \new_[26954]_  & \new_[26943]_ ;
  assign \new_[2317]_  = \new_[26932]_  & \new_[26921]_ ;
  assign \new_[2318]_  = \new_[26910]_  & \new_[26899]_ ;
  assign \new_[2319]_  = \new_[26888]_  & \new_[26877]_ ;
  assign \new_[2320]_  = \new_[26866]_  & \new_[26855]_ ;
  assign \new_[2321]_  = \new_[26844]_  & \new_[26833]_ ;
  assign \new_[2322]_  = \new_[26822]_  & \new_[26811]_ ;
  assign \new_[2323]_  = \new_[26800]_  & \new_[26789]_ ;
  assign \new_[2324]_  = \new_[26778]_  & \new_[26767]_ ;
  assign \new_[2325]_  = \new_[26756]_  & \new_[26745]_ ;
  assign \new_[2326]_  = \new_[26734]_  & \new_[26723]_ ;
  assign \new_[2327]_  = \new_[26712]_  & \new_[26701]_ ;
  assign \new_[2328]_  = \new_[26690]_  & \new_[26679]_ ;
  assign \new_[2329]_  = \new_[26668]_  & \new_[26657]_ ;
  assign \new_[2330]_  = \new_[26646]_  & \new_[26635]_ ;
  assign \new_[2331]_  = \new_[26624]_  & \new_[26613]_ ;
  assign \new_[2332]_  = \new_[26602]_  & \new_[26591]_ ;
  assign \new_[2333]_  = \new_[26580]_  & \new_[26569]_ ;
  assign \new_[2334]_  = \new_[26558]_  & \new_[26547]_ ;
  assign \new_[2335]_  = \new_[26536]_  & \new_[26525]_ ;
  assign \new_[2336]_  = \new_[26514]_  & \new_[26503]_ ;
  assign \new_[2337]_  = \new_[26492]_  & \new_[26481]_ ;
  assign \new_[2338]_  = \new_[26470]_  & \new_[26459]_ ;
  assign \new_[2339]_  = \new_[26448]_  & \new_[26437]_ ;
  assign \new_[2340]_  = \new_[26426]_  & \new_[26415]_ ;
  assign \new_[2341]_  = \new_[26404]_  & \new_[26393]_ ;
  assign \new_[2342]_  = \new_[26382]_  & \new_[26371]_ ;
  assign \new_[2343]_  = \new_[26360]_  & \new_[26349]_ ;
  assign \new_[2344]_  = \new_[26338]_  & \new_[26327]_ ;
  assign \new_[2345]_  = \new_[26316]_  & \new_[26305]_ ;
  assign \new_[2346]_  = \new_[26294]_  & \new_[26283]_ ;
  assign \new_[2347]_  = \new_[26272]_  & \new_[26261]_ ;
  assign \new_[2348]_  = \new_[26250]_  & \new_[26239]_ ;
  assign \new_[2349]_  = \new_[26228]_  & \new_[26217]_ ;
  assign \new_[2350]_  = \new_[26206]_  & \new_[26195]_ ;
  assign \new_[2351]_  = \new_[26184]_  & \new_[26173]_ ;
  assign \new_[2352]_  = \new_[26162]_  & \new_[26151]_ ;
  assign \new_[2353]_  = \new_[26140]_  & \new_[26129]_ ;
  assign \new_[2354]_  = \new_[26118]_  & \new_[26107]_ ;
  assign \new_[2355]_  = \new_[26096]_  & \new_[26085]_ ;
  assign \new_[2356]_  = \new_[26074]_  & \new_[26063]_ ;
  assign \new_[2357]_  = \new_[26052]_  & \new_[26041]_ ;
  assign \new_[2358]_  = \new_[26030]_  & \new_[26019]_ ;
  assign \new_[2359]_  = \new_[26008]_  & \new_[25997]_ ;
  assign \new_[2360]_  = \new_[25986]_  & \new_[25975]_ ;
  assign \new_[2361]_  = \new_[25964]_  & \new_[25953]_ ;
  assign \new_[2362]_  = \new_[25942]_  & \new_[25931]_ ;
  assign \new_[2363]_  = \new_[25920]_  & \new_[25909]_ ;
  assign \new_[2364]_  = \new_[25898]_  & \new_[25887]_ ;
  assign \new_[2365]_  = \new_[25876]_  & \new_[25865]_ ;
  assign \new_[2366]_  = \new_[25854]_  & \new_[25843]_ ;
  assign \new_[2367]_  = \new_[25832]_  & \new_[25821]_ ;
  assign \new_[2368]_  = \new_[25810]_  & \new_[25799]_ ;
  assign \new_[2369]_  = \new_[25788]_  & \new_[25777]_ ;
  assign \new_[2370]_  = \new_[25766]_  & \new_[25755]_ ;
  assign \new_[2371]_  = \new_[25744]_  & \new_[25733]_ ;
  assign \new_[2372]_  = \new_[25722]_  & \new_[25711]_ ;
  assign \new_[2373]_  = \new_[25700]_  & \new_[25689]_ ;
  assign \new_[2374]_  = \new_[25678]_  & \new_[25667]_ ;
  assign \new_[2375]_  = \new_[25656]_  & \new_[25645]_ ;
  assign \new_[2376]_  = \new_[25634]_  & \new_[25623]_ ;
  assign \new_[2377]_  = \new_[25612]_  & \new_[25601]_ ;
  assign \new_[2378]_  = \new_[25590]_  & \new_[25579]_ ;
  assign \new_[2379]_  = \new_[25568]_  & \new_[25557]_ ;
  assign \new_[2380]_  = \new_[25546]_  & \new_[25535]_ ;
  assign \new_[2381]_  = \new_[25524]_  & \new_[25513]_ ;
  assign \new_[2382]_  = \new_[25502]_  & \new_[25491]_ ;
  assign \new_[2383]_  = \new_[25480]_  & \new_[25469]_ ;
  assign \new_[2384]_  = \new_[25458]_  & \new_[25447]_ ;
  assign \new_[2385]_  = \new_[25436]_  & \new_[25425]_ ;
  assign \new_[2386]_  = \new_[25414]_  & \new_[25403]_ ;
  assign \new_[2387]_  = \new_[25392]_  & \new_[25381]_ ;
  assign \new_[2388]_  = \new_[25370]_  & \new_[25359]_ ;
  assign \new_[2389]_  = \new_[25348]_  & \new_[25337]_ ;
  assign \new_[2390]_  = \new_[25326]_  & \new_[25315]_ ;
  assign \new_[2391]_  = \new_[25304]_  & \new_[25293]_ ;
  assign \new_[2392]_  = \new_[25282]_  & \new_[25271]_ ;
  assign \new_[2393]_  = \new_[25260]_  & \new_[25249]_ ;
  assign \new_[2394]_  = \new_[25238]_  & \new_[25227]_ ;
  assign \new_[2395]_  = \new_[25216]_  & \new_[25205]_ ;
  assign \new_[2396]_  = \new_[25194]_  & \new_[25183]_ ;
  assign \new_[2397]_  = \new_[25172]_  & \new_[25161]_ ;
  assign \new_[2398]_  = \new_[25150]_  & \new_[25139]_ ;
  assign \new_[2399]_  = \new_[25128]_  & \new_[25117]_ ;
  assign \new_[2400]_  = \new_[25106]_  & \new_[25095]_ ;
  assign \new_[2401]_  = \new_[25084]_  & \new_[25073]_ ;
  assign \new_[2402]_  = \new_[25062]_  & \new_[25051]_ ;
  assign \new_[2403]_  = \new_[25040]_  & \new_[25029]_ ;
  assign \new_[2404]_  = \new_[25018]_  & \new_[25007]_ ;
  assign \new_[2405]_  = \new_[24996]_  & \new_[24985]_ ;
  assign \new_[2406]_  = \new_[24974]_  & \new_[24963]_ ;
  assign \new_[2407]_  = \new_[24952]_  & \new_[24941]_ ;
  assign \new_[2408]_  = \new_[24930]_  & \new_[24919]_ ;
  assign \new_[2409]_  = \new_[24908]_  & \new_[24897]_ ;
  assign \new_[2410]_  = \new_[24886]_  & \new_[24875]_ ;
  assign \new_[2411]_  = \new_[24864]_  & \new_[24853]_ ;
  assign \new_[2412]_  = \new_[24842]_  & \new_[24831]_ ;
  assign \new_[2413]_  = \new_[24820]_  & \new_[24809]_ ;
  assign \new_[2414]_  = \new_[24798]_  & \new_[24787]_ ;
  assign \new_[2415]_  = \new_[24776]_  & \new_[24765]_ ;
  assign \new_[2416]_  = \new_[24754]_  & \new_[24743]_ ;
  assign \new_[2417]_  = \new_[24732]_  & \new_[24721]_ ;
  assign \new_[2418]_  = \new_[24710]_  & \new_[24699]_ ;
  assign \new_[2419]_  = \new_[24688]_  & \new_[24677]_ ;
  assign \new_[2420]_  = \new_[24666]_  & \new_[24655]_ ;
  assign \new_[2421]_  = \new_[24644]_  & \new_[24633]_ ;
  assign \new_[2422]_  = \new_[24622]_  & \new_[24611]_ ;
  assign \new_[2423]_  = \new_[24600]_  & \new_[24589]_ ;
  assign \new_[2424]_  = \new_[24578]_  & \new_[24567]_ ;
  assign \new_[2425]_  = \new_[24556]_  & \new_[24545]_ ;
  assign \new_[2426]_  = \new_[24534]_  & \new_[24523]_ ;
  assign \new_[2427]_  = \new_[24512]_  & \new_[24501]_ ;
  assign \new_[2428]_  = \new_[24490]_  & \new_[24479]_ ;
  assign \new_[2429]_  = \new_[24468]_  & \new_[24457]_ ;
  assign \new_[2430]_  = \new_[24446]_  & \new_[24435]_ ;
  assign \new_[2431]_  = \new_[24424]_  & \new_[24413]_ ;
  assign \new_[2432]_  = \new_[24402]_  & \new_[24391]_ ;
  assign \new_[2433]_  = \new_[24380]_  & \new_[24369]_ ;
  assign \new_[2434]_  = \new_[24358]_  & \new_[24347]_ ;
  assign \new_[2435]_  = \new_[24336]_  & \new_[24325]_ ;
  assign \new_[2436]_  = \new_[24314]_  & \new_[24303]_ ;
  assign \new_[2437]_  = \new_[24292]_  & \new_[24281]_ ;
  assign \new_[2438]_  = \new_[24270]_  & \new_[24259]_ ;
  assign \new_[2439]_  = \new_[24248]_  & \new_[24237]_ ;
  assign \new_[2440]_  = \new_[24226]_  & \new_[24215]_ ;
  assign \new_[2441]_  = \new_[24204]_  & \new_[24193]_ ;
  assign \new_[2442]_  = \new_[24182]_  & \new_[24171]_ ;
  assign \new_[2443]_  = \new_[24160]_  & \new_[24149]_ ;
  assign \new_[2444]_  = \new_[24138]_  & \new_[24127]_ ;
  assign \new_[2445]_  = \new_[24116]_  & \new_[24105]_ ;
  assign \new_[2446]_  = \new_[24094]_  & \new_[24083]_ ;
  assign \new_[2447]_  = \new_[24072]_  & \new_[24061]_ ;
  assign \new_[2448]_  = \new_[24050]_  & \new_[24039]_ ;
  assign \new_[2449]_  = \new_[24028]_  & \new_[24017]_ ;
  assign \new_[2450]_  = \new_[24006]_  & \new_[23995]_ ;
  assign \new_[2451]_  = \new_[23984]_  & \new_[23973]_ ;
  assign \new_[2452]_  = \new_[23962]_  & \new_[23951]_ ;
  assign \new_[2453]_  = \new_[23940]_  & \new_[23929]_ ;
  assign \new_[2454]_  = \new_[23918]_  & \new_[23907]_ ;
  assign \new_[2455]_  = \new_[23896]_  & \new_[23885]_ ;
  assign \new_[2456]_  = \new_[23874]_  & \new_[23863]_ ;
  assign \new_[2457]_  = \new_[23852]_  & \new_[23841]_ ;
  assign \new_[2458]_  = \new_[23830]_  & \new_[23819]_ ;
  assign \new_[2459]_  = \new_[23808]_  & \new_[23797]_ ;
  assign \new_[2460]_  = \new_[23786]_  & \new_[23775]_ ;
  assign \new_[2461]_  = \new_[23764]_  & \new_[23753]_ ;
  assign \new_[2462]_  = \new_[23742]_  & \new_[23731]_ ;
  assign \new_[2463]_  = \new_[23720]_  & \new_[23709]_ ;
  assign \new_[2464]_  = \new_[23698]_  & \new_[23687]_ ;
  assign \new_[2465]_  = \new_[23676]_  & \new_[23665]_ ;
  assign \new_[2466]_  = \new_[23654]_  & \new_[23643]_ ;
  assign \new_[2467]_  = \new_[23632]_  & \new_[23621]_ ;
  assign \new_[2468]_  = \new_[23610]_  & \new_[23599]_ ;
  assign \new_[2469]_  = \new_[23588]_  & \new_[23577]_ ;
  assign \new_[2470]_  = \new_[23566]_  & \new_[23555]_ ;
  assign \new_[2471]_  = \new_[23544]_  & \new_[23533]_ ;
  assign \new_[2472]_  = \new_[23522]_  & \new_[23511]_ ;
  assign \new_[2473]_  = \new_[23500]_  & \new_[23489]_ ;
  assign \new_[2474]_  = \new_[23478]_  & \new_[23467]_ ;
  assign \new_[2475]_  = \new_[23456]_  & \new_[23445]_ ;
  assign \new_[2476]_  = \new_[23434]_  & \new_[23423]_ ;
  assign \new_[2477]_  = \new_[23412]_  & \new_[23401]_ ;
  assign \new_[2478]_  = \new_[23390]_  & \new_[23379]_ ;
  assign \new_[2479]_  = \new_[23368]_  & \new_[23357]_ ;
  assign \new_[2480]_  = \new_[23346]_  & \new_[23335]_ ;
  assign \new_[2481]_  = \new_[23324]_  & \new_[23313]_ ;
  assign \new_[2482]_  = \new_[23302]_  & \new_[23291]_ ;
  assign \new_[2483]_  = \new_[23280]_  & \new_[23269]_ ;
  assign \new_[2484]_  = \new_[23258]_  & \new_[23247]_ ;
  assign \new_[2485]_  = \new_[23236]_  & \new_[23225]_ ;
  assign \new_[2486]_  = \new_[23214]_  & \new_[23203]_ ;
  assign \new_[2487]_  = \new_[23192]_  & \new_[23181]_ ;
  assign \new_[2488]_  = \new_[23170]_  & \new_[23159]_ ;
  assign \new_[2489]_  = \new_[23148]_  & \new_[23137]_ ;
  assign \new_[2490]_  = \new_[23126]_  & \new_[23115]_ ;
  assign \new_[2491]_  = \new_[23104]_  & \new_[23093]_ ;
  assign \new_[2492]_  = \new_[23082]_  & \new_[23071]_ ;
  assign \new_[2493]_  = \new_[23060]_  & \new_[23049]_ ;
  assign \new_[2494]_  = \new_[23038]_  & \new_[23027]_ ;
  assign \new_[2495]_  = \new_[23016]_  & \new_[23005]_ ;
  assign \new_[2496]_  = \new_[22994]_  & \new_[22983]_ ;
  assign \new_[2497]_  = \new_[22972]_  & \new_[22961]_ ;
  assign \new_[2498]_  = \new_[22950]_  & \new_[22939]_ ;
  assign \new_[2499]_  = \new_[22928]_  & \new_[22917]_ ;
  assign \new_[2500]_  = \new_[22906]_  & \new_[22895]_ ;
  assign \new_[2501]_  = \new_[22884]_  & \new_[22873]_ ;
  assign \new_[2502]_  = \new_[22862]_  & \new_[22851]_ ;
  assign \new_[2503]_  = \new_[22840]_  & \new_[22829]_ ;
  assign \new_[2504]_  = \new_[22818]_  & \new_[22807]_ ;
  assign \new_[2505]_  = \new_[22796]_  & \new_[22785]_ ;
  assign \new_[2506]_  = \new_[22774]_  & \new_[22763]_ ;
  assign \new_[2507]_  = \new_[22752]_  & \new_[22741]_ ;
  assign \new_[2508]_  = \new_[22730]_  & \new_[22719]_ ;
  assign \new_[2509]_  = \new_[22708]_  & \new_[22697]_ ;
  assign \new_[2510]_  = \new_[22686]_  & \new_[22675]_ ;
  assign \new_[2511]_  = \new_[22664]_  & \new_[22653]_ ;
  assign \new_[2512]_  = \new_[22642]_  & \new_[22631]_ ;
  assign \new_[2513]_  = \new_[22620]_  & \new_[22609]_ ;
  assign \new_[2514]_  = \new_[22598]_  & \new_[22587]_ ;
  assign \new_[2515]_  = \new_[22576]_  & \new_[22565]_ ;
  assign \new_[2516]_  = \new_[22554]_  & \new_[22543]_ ;
  assign \new_[2517]_  = \new_[22532]_  & \new_[22521]_ ;
  assign \new_[2518]_  = \new_[22510]_  & \new_[22499]_ ;
  assign \new_[2519]_  = \new_[22488]_  & \new_[22477]_ ;
  assign \new_[2520]_  = \new_[22466]_  & \new_[22455]_ ;
  assign \new_[2521]_  = \new_[22444]_  & \new_[22433]_ ;
  assign \new_[2522]_  = \new_[22422]_  & \new_[22411]_ ;
  assign \new_[2523]_  = \new_[22400]_  & \new_[22389]_ ;
  assign \new_[2524]_  = \new_[22378]_  & \new_[22367]_ ;
  assign \new_[2525]_  = \new_[22356]_  & \new_[22345]_ ;
  assign \new_[2526]_  = \new_[22334]_  & \new_[22323]_ ;
  assign \new_[2527]_  = \new_[22312]_  & \new_[22301]_ ;
  assign \new_[2528]_  = \new_[22290]_  & \new_[22279]_ ;
  assign \new_[2529]_  = \new_[22268]_  & \new_[22257]_ ;
  assign \new_[2530]_  = \new_[22246]_  & \new_[22235]_ ;
  assign \new_[2531]_  = \new_[22224]_  & \new_[22213]_ ;
  assign \new_[2532]_  = \new_[22202]_  & \new_[22191]_ ;
  assign \new_[2533]_  = \new_[22180]_  & \new_[22169]_ ;
  assign \new_[2534]_  = \new_[22158]_  & \new_[22147]_ ;
  assign \new_[2535]_  = \new_[22136]_  & \new_[22125]_ ;
  assign \new_[2536]_  = \new_[22114]_  & \new_[22103]_ ;
  assign \new_[2537]_  = \new_[22092]_  & \new_[22081]_ ;
  assign \new_[2538]_  = \new_[22070]_  & \new_[22059]_ ;
  assign \new_[2539]_  = \new_[22048]_  & \new_[22037]_ ;
  assign \new_[2540]_  = \new_[22026]_  & \new_[22015]_ ;
  assign \new_[2541]_  = \new_[22004]_  & \new_[21993]_ ;
  assign \new_[2542]_  = \new_[21982]_  & \new_[21971]_ ;
  assign \new_[2543]_  = \new_[21960]_  & \new_[21949]_ ;
  assign \new_[2544]_  = \new_[21938]_  & \new_[21927]_ ;
  assign \new_[2545]_  = \new_[21916]_  & \new_[21905]_ ;
  assign \new_[2546]_  = \new_[21894]_  & \new_[21883]_ ;
  assign \new_[2547]_  = \new_[21872]_  & \new_[21861]_ ;
  assign \new_[2548]_  = \new_[21850]_  & \new_[21839]_ ;
  assign \new_[2549]_  = \new_[21828]_  & \new_[21817]_ ;
  assign \new_[2550]_  = \new_[21806]_  & \new_[21795]_ ;
  assign \new_[2551]_  = \new_[21784]_  & \new_[21773]_ ;
  assign \new_[2552]_  = \new_[21762]_  & \new_[21751]_ ;
  assign \new_[2553]_  = \new_[21740]_  & \new_[21729]_ ;
  assign \new_[2554]_  = \new_[21718]_  & \new_[21707]_ ;
  assign \new_[2555]_  = \new_[21696]_  & \new_[21685]_ ;
  assign \new_[2556]_  = \new_[21674]_  & \new_[21663]_ ;
  assign \new_[2557]_  = \new_[21652]_  & \new_[21641]_ ;
  assign \new_[2558]_  = \new_[21630]_  & \new_[21619]_ ;
  assign \new_[2559]_  = \new_[21608]_  & \new_[21597]_ ;
  assign \new_[2560]_  = \new_[21586]_  & \new_[21575]_ ;
  assign \new_[2561]_  = \new_[21564]_  & \new_[21553]_ ;
  assign \new_[2562]_  = \new_[21542]_  & \new_[21531]_ ;
  assign \new_[2563]_  = \new_[21520]_  & \new_[21509]_ ;
  assign \new_[2564]_  = \new_[21498]_  & \new_[21487]_ ;
  assign \new_[2565]_  = \new_[21476]_  & \new_[21465]_ ;
  assign \new_[2566]_  = \new_[21454]_  & \new_[21443]_ ;
  assign \new_[2567]_  = \new_[21432]_  & \new_[21421]_ ;
  assign \new_[2568]_  = \new_[21410]_  & \new_[21399]_ ;
  assign \new_[2569]_  = \new_[21388]_  & \new_[21377]_ ;
  assign \new_[2570]_  = \new_[21366]_  & \new_[21355]_ ;
  assign \new_[2571]_  = \new_[21344]_  & \new_[21333]_ ;
  assign \new_[2572]_  = \new_[21322]_  & \new_[21311]_ ;
  assign \new_[2573]_  = \new_[21300]_  & \new_[21289]_ ;
  assign \new_[2574]_  = \new_[21278]_  & \new_[21267]_ ;
  assign \new_[2575]_  = \new_[21256]_  & \new_[21245]_ ;
  assign \new_[2576]_  = \new_[21234]_  & \new_[21223]_ ;
  assign \new_[2577]_  = \new_[21212]_  & \new_[21201]_ ;
  assign \new_[2578]_  = \new_[21190]_  & \new_[21179]_ ;
  assign \new_[2579]_  = \new_[21168]_  & \new_[21157]_ ;
  assign \new_[2580]_  = \new_[21146]_  & \new_[21135]_ ;
  assign \new_[2581]_  = \new_[21124]_  & \new_[21113]_ ;
  assign \new_[2582]_  = \new_[21102]_  & \new_[21091]_ ;
  assign \new_[2583]_  = \new_[21080]_  & \new_[21069]_ ;
  assign \new_[2584]_  = \new_[21058]_  & \new_[21047]_ ;
  assign \new_[2585]_  = \new_[21036]_  & \new_[21025]_ ;
  assign \new_[2586]_  = \new_[21014]_  & \new_[21003]_ ;
  assign \new_[2587]_  = \new_[20992]_  & \new_[20981]_ ;
  assign \new_[2588]_  = \new_[20970]_  & \new_[20959]_ ;
  assign \new_[2589]_  = \new_[20948]_  & \new_[20937]_ ;
  assign \new_[2590]_  = \new_[20926]_  & \new_[20915]_ ;
  assign \new_[2591]_  = \new_[20904]_  & \new_[20893]_ ;
  assign \new_[2592]_  = \new_[20882]_  & \new_[20871]_ ;
  assign \new_[2593]_  = \new_[20860]_  & \new_[20849]_ ;
  assign \new_[2594]_  = \new_[20838]_  & \new_[20827]_ ;
  assign \new_[2595]_  = \new_[20816]_  & \new_[20805]_ ;
  assign \new_[2596]_  = \new_[20794]_  & \new_[20783]_ ;
  assign \new_[2597]_  = \new_[20772]_  & \new_[20761]_ ;
  assign \new_[2598]_  = \new_[20750]_  & \new_[20739]_ ;
  assign \new_[2599]_  = \new_[20728]_  & \new_[20717]_ ;
  assign \new_[2600]_  = \new_[20706]_  & \new_[20695]_ ;
  assign \new_[2601]_  = \new_[20684]_  & \new_[20673]_ ;
  assign \new_[2602]_  = \new_[20662]_  & \new_[20651]_ ;
  assign \new_[2603]_  = \new_[20640]_  & \new_[20629]_ ;
  assign \new_[2604]_  = \new_[20618]_  & \new_[20607]_ ;
  assign \new_[2605]_  = \new_[20596]_  & \new_[20585]_ ;
  assign \new_[2606]_  = \new_[20574]_  & \new_[20563]_ ;
  assign \new_[2607]_  = \new_[20552]_  & \new_[20541]_ ;
  assign \new_[2608]_  = \new_[20530]_  & \new_[20519]_ ;
  assign \new_[2609]_  = \new_[20508]_  & \new_[20497]_ ;
  assign \new_[2610]_  = \new_[20486]_  & \new_[20475]_ ;
  assign \new_[2611]_  = \new_[20464]_  & \new_[20453]_ ;
  assign \new_[2612]_  = \new_[20442]_  & \new_[20431]_ ;
  assign \new_[2613]_  = \new_[20420]_  & \new_[20409]_ ;
  assign \new_[2614]_  = \new_[20398]_  & \new_[20387]_ ;
  assign \new_[2615]_  = \new_[20376]_  & \new_[20365]_ ;
  assign \new_[2616]_  = \new_[20354]_  & \new_[20343]_ ;
  assign \new_[2617]_  = \new_[20332]_  & \new_[20321]_ ;
  assign \new_[2618]_  = \new_[20310]_  & \new_[20299]_ ;
  assign \new_[2619]_  = \new_[20288]_  & \new_[20277]_ ;
  assign \new_[2620]_  = \new_[20266]_  & \new_[20255]_ ;
  assign \new_[2621]_  = \new_[20244]_  & \new_[20233]_ ;
  assign \new_[2622]_  = \new_[20222]_  & \new_[20211]_ ;
  assign \new_[2623]_  = \new_[20200]_  & \new_[20189]_ ;
  assign \new_[2624]_  = \new_[20178]_  & \new_[20167]_ ;
  assign \new_[2625]_  = \new_[20156]_  & \new_[20145]_ ;
  assign \new_[2626]_  = \new_[20134]_  & \new_[20123]_ ;
  assign \new_[2627]_  = \new_[20112]_  & \new_[20101]_ ;
  assign \new_[2628]_  = \new_[20090]_  & \new_[20079]_ ;
  assign \new_[2629]_  = \new_[20068]_  & \new_[20057]_ ;
  assign \new_[2630]_  = \new_[20046]_  & \new_[20035]_ ;
  assign \new_[2631]_  = \new_[20024]_  & \new_[20013]_ ;
  assign \new_[2632]_  = \new_[20002]_  & \new_[19991]_ ;
  assign \new_[2633]_  = \new_[19980]_  & \new_[19969]_ ;
  assign \new_[2634]_  = \new_[19958]_  & \new_[19947]_ ;
  assign \new_[2635]_  = \new_[19936]_  & \new_[19925]_ ;
  assign \new_[2636]_  = \new_[19914]_  & \new_[19903]_ ;
  assign \new_[2637]_  = \new_[19892]_  & \new_[19881]_ ;
  assign \new_[2638]_  = \new_[19870]_  & \new_[19859]_ ;
  assign \new_[2639]_  = \new_[19848]_  & \new_[19837]_ ;
  assign \new_[2640]_  = \new_[19826]_  & \new_[19815]_ ;
  assign \new_[2641]_  = \new_[19804]_  & \new_[19793]_ ;
  assign \new_[2642]_  = \new_[19782]_  & \new_[19771]_ ;
  assign \new_[2643]_  = \new_[19760]_  & \new_[19749]_ ;
  assign \new_[2644]_  = \new_[19738]_  & \new_[19727]_ ;
  assign \new_[2645]_  = \new_[19716]_  & \new_[19705]_ ;
  assign \new_[2646]_  = \new_[19694]_  & \new_[19683]_ ;
  assign \new_[2647]_  = \new_[19672]_  & \new_[19661]_ ;
  assign \new_[2648]_  = \new_[19650]_  & \new_[19639]_ ;
  assign \new_[2649]_  = \new_[19628]_  & \new_[19617]_ ;
  assign \new_[2650]_  = \new_[19606]_  & \new_[19595]_ ;
  assign \new_[2651]_  = \new_[19584]_  & \new_[19573]_ ;
  assign \new_[2652]_  = \new_[19562]_  & \new_[19551]_ ;
  assign \new_[2653]_  = \new_[19540]_  & \new_[19529]_ ;
  assign \new_[2654]_  = \new_[19518]_  & \new_[19507]_ ;
  assign \new_[2655]_  = \new_[19496]_  & \new_[19485]_ ;
  assign \new_[2656]_  = \new_[19474]_  & \new_[19463]_ ;
  assign \new_[2657]_  = \new_[19452]_  & \new_[19441]_ ;
  assign \new_[2658]_  = \new_[19430]_  & \new_[19419]_ ;
  assign \new_[2659]_  = \new_[19408]_  & \new_[19397]_ ;
  assign \new_[2660]_  = \new_[19386]_  & \new_[19375]_ ;
  assign \new_[2661]_  = \new_[19364]_  & \new_[19353]_ ;
  assign \new_[2662]_  = \new_[19342]_  & \new_[19331]_ ;
  assign \new_[2663]_  = \new_[19320]_  & \new_[19309]_ ;
  assign \new_[2664]_  = \new_[19298]_  & \new_[19287]_ ;
  assign \new_[2665]_  = \new_[19276]_  & \new_[19265]_ ;
  assign \new_[2666]_  = \new_[19254]_  & \new_[19243]_ ;
  assign \new_[2667]_  = \new_[19232]_  & \new_[19221]_ ;
  assign \new_[2668]_  = \new_[19210]_  & \new_[19199]_ ;
  assign \new_[2669]_  = \new_[19188]_  & \new_[19177]_ ;
  assign \new_[2670]_  = \new_[19166]_  & \new_[19155]_ ;
  assign \new_[2671]_  = \new_[19144]_  & \new_[19133]_ ;
  assign \new_[2672]_  = \new_[19122]_  & \new_[19111]_ ;
  assign \new_[2673]_  = \new_[19100]_  & \new_[19089]_ ;
  assign \new_[2674]_  = \new_[19078]_  & \new_[19067]_ ;
  assign \new_[2675]_  = \new_[19056]_  & \new_[19045]_ ;
  assign \new_[2676]_  = \new_[19034]_  & \new_[19023]_ ;
  assign \new_[2677]_  = \new_[19012]_  & \new_[19001]_ ;
  assign \new_[2678]_  = \new_[18990]_  & \new_[18979]_ ;
  assign \new_[2679]_  = \new_[18968]_  & \new_[18957]_ ;
  assign \new_[2680]_  = \new_[18946]_  & \new_[18935]_ ;
  assign \new_[2681]_  = \new_[18924]_  & \new_[18913]_ ;
  assign \new_[2682]_  = \new_[18902]_  & \new_[18891]_ ;
  assign \new_[2683]_  = \new_[18880]_  & \new_[18869]_ ;
  assign \new_[2684]_  = \new_[18858]_  & \new_[18847]_ ;
  assign \new_[2685]_  = \new_[18836]_  & \new_[18825]_ ;
  assign \new_[2686]_  = \new_[18814]_  & \new_[18803]_ ;
  assign \new_[2687]_  = \new_[18792]_  & \new_[18781]_ ;
  assign \new_[2688]_  = \new_[18770]_  & \new_[18759]_ ;
  assign \new_[2689]_  = \new_[18748]_  & \new_[18737]_ ;
  assign \new_[2690]_  = \new_[18726]_  & \new_[18715]_ ;
  assign \new_[2691]_  = \new_[18704]_  & \new_[18693]_ ;
  assign \new_[2692]_  = \new_[18682]_  & \new_[18671]_ ;
  assign \new_[2693]_  = \new_[18660]_  & \new_[18649]_ ;
  assign \new_[2694]_  = \new_[18638]_  & \new_[18627]_ ;
  assign \new_[2695]_  = \new_[18616]_  & \new_[18605]_ ;
  assign \new_[2696]_  = \new_[18594]_  & \new_[18583]_ ;
  assign \new_[2697]_  = \new_[18572]_  & \new_[18561]_ ;
  assign \new_[2698]_  = \new_[18550]_  & \new_[18539]_ ;
  assign \new_[2699]_  = \new_[18528]_  & \new_[18517]_ ;
  assign \new_[2700]_  = \new_[18506]_  & \new_[18495]_ ;
  assign \new_[2701]_  = \new_[18484]_  & \new_[18473]_ ;
  assign \new_[2702]_  = \new_[18462]_  & \new_[18451]_ ;
  assign \new_[2703]_  = \new_[18440]_  & \new_[18429]_ ;
  assign \new_[2704]_  = \new_[18418]_  & \new_[18407]_ ;
  assign \new_[2705]_  = \new_[18396]_  & \new_[18385]_ ;
  assign \new_[2706]_  = \new_[18374]_  & \new_[18363]_ ;
  assign \new_[2707]_  = \new_[18352]_  & \new_[18341]_ ;
  assign \new_[2708]_  = \new_[18330]_  & \new_[18319]_ ;
  assign \new_[2709]_  = \new_[18308]_  & \new_[18297]_ ;
  assign \new_[2710]_  = \new_[18286]_  & \new_[18275]_ ;
  assign \new_[2711]_  = \new_[18264]_  & \new_[18253]_ ;
  assign \new_[2712]_  = \new_[18242]_  & \new_[18231]_ ;
  assign \new_[2713]_  = \new_[18220]_  & \new_[18209]_ ;
  assign \new_[2714]_  = \new_[18198]_  & \new_[18187]_ ;
  assign \new_[2715]_  = \new_[18176]_  & \new_[18165]_ ;
  assign \new_[2716]_  = \new_[18154]_  & \new_[18143]_ ;
  assign \new_[2717]_  = \new_[18132]_  & \new_[18121]_ ;
  assign \new_[2718]_  = \new_[18110]_  & \new_[18099]_ ;
  assign \new_[2719]_  = \new_[18088]_  & \new_[18077]_ ;
  assign \new_[2720]_  = \new_[18066]_  & \new_[18055]_ ;
  assign \new_[2721]_  = \new_[18044]_  & \new_[18033]_ ;
  assign \new_[2722]_  = \new_[18022]_  & \new_[18011]_ ;
  assign \new_[2723]_  = \new_[18000]_  & \new_[17989]_ ;
  assign \new_[2724]_  = \new_[17978]_  & \new_[17967]_ ;
  assign \new_[2725]_  = \new_[17956]_  & \new_[17945]_ ;
  assign \new_[2726]_  = \new_[17934]_  & \new_[17923]_ ;
  assign \new_[2727]_  = \new_[17912]_  & \new_[17901]_ ;
  assign \new_[2728]_  = \new_[17890]_  & \new_[17879]_ ;
  assign \new_[2729]_  = \new_[17868]_  & \new_[17857]_ ;
  assign \new_[2730]_  = \new_[17846]_  & \new_[17835]_ ;
  assign \new_[2731]_  = \new_[17824]_  & \new_[17813]_ ;
  assign \new_[2732]_  = \new_[17802]_  & \new_[17791]_ ;
  assign \new_[2733]_  = \new_[17780]_  & \new_[17769]_ ;
  assign \new_[2734]_  = \new_[17758]_  & \new_[17747]_ ;
  assign \new_[2735]_  = \new_[17736]_  & \new_[17725]_ ;
  assign \new_[2736]_  = \new_[17714]_  & \new_[17703]_ ;
  assign \new_[2737]_  = \new_[17692]_  & \new_[17681]_ ;
  assign \new_[2738]_  = \new_[17670]_  & \new_[17659]_ ;
  assign \new_[2739]_  = \new_[17648]_  & \new_[17637]_ ;
  assign \new_[2740]_  = \new_[17626]_  & \new_[17615]_ ;
  assign \new_[2741]_  = \new_[17604]_  & \new_[17593]_ ;
  assign \new_[2742]_  = \new_[17582]_  & \new_[17571]_ ;
  assign \new_[2743]_  = \new_[17560]_  & \new_[17549]_ ;
  assign \new_[2744]_  = \new_[17538]_  & \new_[17527]_ ;
  assign \new_[2745]_  = \new_[17516]_  & \new_[17505]_ ;
  assign \new_[2746]_  = \new_[17494]_  & \new_[17483]_ ;
  assign \new_[2747]_  = \new_[17472]_  & \new_[17461]_ ;
  assign \new_[2748]_  = \new_[17450]_  & \new_[17439]_ ;
  assign \new_[2749]_  = \new_[17428]_  & \new_[17417]_ ;
  assign \new_[2750]_  = \new_[17408]_  & \new_[17397]_ ;
  assign \new_[2751]_  = \new_[17388]_  & \new_[17377]_ ;
  assign \new_[2752]_  = \new_[17368]_  & \new_[17357]_ ;
  assign \new_[2753]_  = \new_[17348]_  & \new_[17337]_ ;
  assign \new_[2754]_  = \new_[17328]_  & \new_[17317]_ ;
  assign \new_[2755]_  = \new_[17308]_  & \new_[17297]_ ;
  assign \new_[2756]_  = \new_[17288]_  & \new_[17277]_ ;
  assign \new_[2757]_  = \new_[17268]_  & \new_[17257]_ ;
  assign \new_[2758]_  = \new_[17248]_  & \new_[17237]_ ;
  assign \new_[2759]_  = \new_[17228]_  & \new_[17217]_ ;
  assign \new_[2760]_  = \new_[17208]_  & \new_[17197]_ ;
  assign \new_[2761]_  = \new_[17188]_  & \new_[17177]_ ;
  assign \new_[2762]_  = \new_[17168]_  & \new_[17157]_ ;
  assign \new_[2763]_  = \new_[17148]_  & \new_[17137]_ ;
  assign \new_[2764]_  = \new_[17128]_  & \new_[17117]_ ;
  assign \new_[2765]_  = \new_[17108]_  & \new_[17097]_ ;
  assign \new_[2766]_  = \new_[17088]_  & \new_[17077]_ ;
  assign \new_[2767]_  = \new_[17068]_  & \new_[17057]_ ;
  assign \new_[2768]_  = \new_[17048]_  & \new_[17037]_ ;
  assign \new_[2769]_  = \new_[17028]_  & \new_[17017]_ ;
  assign \new_[2770]_  = \new_[17008]_  & \new_[16997]_ ;
  assign \new_[2771]_  = \new_[16988]_  & \new_[16977]_ ;
  assign \new_[2772]_  = \new_[16968]_  & \new_[16957]_ ;
  assign \new_[2773]_  = \new_[16948]_  & \new_[16937]_ ;
  assign \new_[2774]_  = \new_[16928]_  & \new_[16917]_ ;
  assign \new_[2775]_  = \new_[16908]_  & \new_[16897]_ ;
  assign \new_[2776]_  = \new_[16888]_  & \new_[16877]_ ;
  assign \new_[2777]_  = \new_[16868]_  & \new_[16857]_ ;
  assign \new_[2778]_  = \new_[16848]_  & \new_[16837]_ ;
  assign \new_[2779]_  = \new_[16828]_  & \new_[16817]_ ;
  assign \new_[2780]_  = \new_[16808]_  & \new_[16797]_ ;
  assign \new_[2781]_  = \new_[16788]_  & \new_[16777]_ ;
  assign \new_[2782]_  = \new_[16768]_  & \new_[16757]_ ;
  assign \new_[2783]_  = \new_[16748]_  & \new_[16737]_ ;
  assign \new_[2784]_  = \new_[16728]_  & \new_[16717]_ ;
  assign \new_[2785]_  = \new_[16708]_  & \new_[16697]_ ;
  assign \new_[2786]_  = \new_[16688]_  & \new_[16677]_ ;
  assign \new_[2787]_  = \new_[16668]_  & \new_[16657]_ ;
  assign \new_[2788]_  = \new_[16648]_  & \new_[16637]_ ;
  assign \new_[2789]_  = \new_[16628]_  & \new_[16617]_ ;
  assign \new_[2790]_  = \new_[16608]_  & \new_[16597]_ ;
  assign \new_[2791]_  = \new_[16588]_  & \new_[16577]_ ;
  assign \new_[2792]_  = \new_[16568]_  & \new_[16557]_ ;
  assign \new_[2793]_  = \new_[16548]_  & \new_[16537]_ ;
  assign \new_[2794]_  = \new_[16528]_  & \new_[16517]_ ;
  assign \new_[2795]_  = \new_[16508]_  & \new_[16497]_ ;
  assign \new_[2796]_  = \new_[16488]_  & \new_[16477]_ ;
  assign \new_[2797]_  = \new_[16468]_  & \new_[16457]_ ;
  assign \new_[2798]_  = \new_[16448]_  & \new_[16437]_ ;
  assign \new_[2799]_  = \new_[16428]_  & \new_[16417]_ ;
  assign \new_[2800]_  = \new_[16408]_  & \new_[16397]_ ;
  assign \new_[2801]_  = \new_[16388]_  & \new_[16377]_ ;
  assign \new_[2802]_  = \new_[16368]_  & \new_[16357]_ ;
  assign \new_[2803]_  = \new_[16348]_  & \new_[16337]_ ;
  assign \new_[2804]_  = \new_[16328]_  & \new_[16317]_ ;
  assign \new_[2805]_  = \new_[16308]_  & \new_[16297]_ ;
  assign \new_[2806]_  = \new_[16288]_  & \new_[16277]_ ;
  assign \new_[2807]_  = \new_[16268]_  & \new_[16257]_ ;
  assign \new_[2808]_  = \new_[16248]_  & \new_[16237]_ ;
  assign \new_[2809]_  = \new_[16228]_  & \new_[16217]_ ;
  assign \new_[2810]_  = \new_[16208]_  & \new_[16197]_ ;
  assign \new_[2811]_  = \new_[16188]_  & \new_[16177]_ ;
  assign \new_[2812]_  = \new_[16168]_  & \new_[16157]_ ;
  assign \new_[2813]_  = \new_[16148]_  & \new_[16137]_ ;
  assign \new_[2814]_  = \new_[16128]_  & \new_[16117]_ ;
  assign \new_[2815]_  = \new_[16108]_  & \new_[16097]_ ;
  assign \new_[2816]_  = \new_[16088]_  & \new_[16077]_ ;
  assign \new_[2817]_  = \new_[16068]_  & \new_[16057]_ ;
  assign \new_[2818]_  = \new_[16048]_  & \new_[16037]_ ;
  assign \new_[2819]_  = \new_[16028]_  & \new_[16017]_ ;
  assign \new_[2820]_  = \new_[16008]_  & \new_[15997]_ ;
  assign \new_[2821]_  = \new_[15988]_  & \new_[15977]_ ;
  assign \new_[2822]_  = \new_[15968]_  & \new_[15957]_ ;
  assign \new_[2823]_  = \new_[15948]_  & \new_[15937]_ ;
  assign \new_[2824]_  = \new_[15928]_  & \new_[15917]_ ;
  assign \new_[2825]_  = \new_[15908]_  & \new_[15897]_ ;
  assign \new_[2826]_  = \new_[15888]_  & \new_[15877]_ ;
  assign \new_[2827]_  = \new_[15868]_  & \new_[15857]_ ;
  assign \new_[2828]_  = \new_[15848]_  & \new_[15837]_ ;
  assign \new_[2829]_  = \new_[15828]_  & \new_[15817]_ ;
  assign \new_[2830]_  = \new_[15808]_  & \new_[15797]_ ;
  assign \new_[2831]_  = \new_[15788]_  & \new_[15777]_ ;
  assign \new_[2832]_  = \new_[15768]_  & \new_[15757]_ ;
  assign \new_[2833]_  = \new_[15748]_  & \new_[15737]_ ;
  assign \new_[2834]_  = \new_[15728]_  & \new_[15717]_ ;
  assign \new_[2835]_  = \new_[15708]_  & \new_[15697]_ ;
  assign \new_[2836]_  = \new_[15688]_  & \new_[15677]_ ;
  assign \new_[2837]_  = \new_[15668]_  & \new_[15657]_ ;
  assign \new_[2838]_  = \new_[15648]_  & \new_[15637]_ ;
  assign \new_[2839]_  = \new_[15628]_  & \new_[15617]_ ;
  assign \new_[2840]_  = \new_[15608]_  & \new_[15597]_ ;
  assign \new_[2841]_  = \new_[15588]_  & \new_[15577]_ ;
  assign \new_[2842]_  = \new_[15568]_  & \new_[15557]_ ;
  assign \new_[2843]_  = \new_[15548]_  & \new_[15537]_ ;
  assign \new_[2844]_  = \new_[15528]_  & \new_[15517]_ ;
  assign \new_[2845]_  = \new_[15508]_  & \new_[15497]_ ;
  assign \new_[2846]_  = \new_[15488]_  & \new_[15477]_ ;
  assign \new_[2847]_  = \new_[15468]_  & \new_[15457]_ ;
  assign \new_[2848]_  = \new_[15448]_  & \new_[15437]_ ;
  assign \new_[2849]_  = \new_[15428]_  & \new_[15417]_ ;
  assign \new_[2850]_  = \new_[15408]_  & \new_[15397]_ ;
  assign \new_[2851]_  = \new_[15388]_  & \new_[15377]_ ;
  assign \new_[2852]_  = \new_[15368]_  & \new_[15357]_ ;
  assign \new_[2853]_  = \new_[15348]_  & \new_[15337]_ ;
  assign \new_[2854]_  = \new_[15328]_  & \new_[15317]_ ;
  assign \new_[2855]_  = \new_[15308]_  & \new_[15297]_ ;
  assign \new_[2856]_  = \new_[15288]_  & \new_[15277]_ ;
  assign \new_[2857]_  = \new_[15268]_  & \new_[15257]_ ;
  assign \new_[2858]_  = \new_[15248]_  & \new_[15237]_ ;
  assign \new_[2859]_  = \new_[15228]_  & \new_[15217]_ ;
  assign \new_[2860]_  = \new_[15208]_  & \new_[15197]_ ;
  assign \new_[2861]_  = \new_[15188]_  & \new_[15177]_ ;
  assign \new_[2862]_  = \new_[15168]_  & \new_[15157]_ ;
  assign \new_[2863]_  = \new_[15148]_  & \new_[15137]_ ;
  assign \new_[2864]_  = \new_[15128]_  & \new_[15117]_ ;
  assign \new_[2865]_  = \new_[15108]_  & \new_[15097]_ ;
  assign \new_[2866]_  = \new_[15088]_  & \new_[15077]_ ;
  assign \new_[2867]_  = \new_[15068]_  & \new_[15057]_ ;
  assign \new_[2868]_  = \new_[15048]_  & \new_[15037]_ ;
  assign \new_[2869]_  = \new_[15028]_  & \new_[15017]_ ;
  assign \new_[2870]_  = \new_[15008]_  & \new_[14997]_ ;
  assign \new_[2871]_  = \new_[14988]_  & \new_[14977]_ ;
  assign \new_[2872]_  = \new_[14968]_  & \new_[14957]_ ;
  assign \new_[2873]_  = \new_[14948]_  & \new_[14937]_ ;
  assign \new_[2874]_  = \new_[14928]_  & \new_[14917]_ ;
  assign \new_[2875]_  = \new_[14908]_  & \new_[14897]_ ;
  assign \new_[2876]_  = \new_[14888]_  & \new_[14877]_ ;
  assign \new_[2877]_  = \new_[14868]_  & \new_[14857]_ ;
  assign \new_[2878]_  = \new_[14848]_  & \new_[14837]_ ;
  assign \new_[2879]_  = \new_[14828]_  & \new_[14817]_ ;
  assign \new_[2880]_  = \new_[14808]_  & \new_[14797]_ ;
  assign \new_[2881]_  = \new_[14788]_  & \new_[14777]_ ;
  assign \new_[2882]_  = \new_[14768]_  & \new_[14757]_ ;
  assign \new_[2883]_  = \new_[14748]_  & \new_[14737]_ ;
  assign \new_[2884]_  = \new_[14728]_  & \new_[14717]_ ;
  assign \new_[2885]_  = \new_[14708]_  & \new_[14697]_ ;
  assign \new_[2886]_  = \new_[14688]_  & \new_[14677]_ ;
  assign \new_[2887]_  = \new_[14668]_  & \new_[14657]_ ;
  assign \new_[2888]_  = \new_[14648]_  & \new_[14637]_ ;
  assign \new_[2889]_  = \new_[14628]_  & \new_[14617]_ ;
  assign \new_[2890]_  = \new_[14608]_  & \new_[14597]_ ;
  assign \new_[2891]_  = \new_[14588]_  & \new_[14577]_ ;
  assign \new_[2892]_  = \new_[14568]_  & \new_[14557]_ ;
  assign \new_[2893]_  = \new_[14548]_  & \new_[14537]_ ;
  assign \new_[2894]_  = \new_[14528]_  & \new_[14517]_ ;
  assign \new_[2895]_  = \new_[14508]_  & \new_[14497]_ ;
  assign \new_[2896]_  = \new_[14488]_  & \new_[14477]_ ;
  assign \new_[2897]_  = \new_[14468]_  & \new_[14457]_ ;
  assign \new_[2898]_  = \new_[14448]_  & \new_[14437]_ ;
  assign \new_[2899]_  = \new_[14428]_  & \new_[14417]_ ;
  assign \new_[2900]_  = \new_[14408]_  & \new_[14397]_ ;
  assign \new_[2901]_  = \new_[14388]_  & \new_[14377]_ ;
  assign \new_[2902]_  = \new_[14368]_  & \new_[14357]_ ;
  assign \new_[2903]_  = \new_[14348]_  & \new_[14337]_ ;
  assign \new_[2904]_  = \new_[14328]_  & \new_[14317]_ ;
  assign \new_[2905]_  = \new_[14308]_  & \new_[14297]_ ;
  assign \new_[2906]_  = \new_[14288]_  & \new_[14277]_ ;
  assign \new_[2907]_  = \new_[14268]_  & \new_[14257]_ ;
  assign \new_[2908]_  = \new_[14248]_  & \new_[14237]_ ;
  assign \new_[2909]_  = \new_[14228]_  & \new_[14217]_ ;
  assign \new_[2910]_  = \new_[14208]_  & \new_[14197]_ ;
  assign \new_[2911]_  = \new_[14188]_  & \new_[14177]_ ;
  assign \new_[2912]_  = \new_[14168]_  & \new_[14157]_ ;
  assign \new_[2913]_  = \new_[14148]_  & \new_[14137]_ ;
  assign \new_[2914]_  = \new_[14128]_  & \new_[14117]_ ;
  assign \new_[2915]_  = \new_[14108]_  & \new_[14097]_ ;
  assign \new_[2916]_  = \new_[14088]_  & \new_[14077]_ ;
  assign \new_[2917]_  = \new_[14068]_  & \new_[14057]_ ;
  assign \new_[2918]_  = \new_[14048]_  & \new_[14037]_ ;
  assign \new_[2919]_  = \new_[14028]_  & \new_[14017]_ ;
  assign \new_[2920]_  = \new_[14008]_  & \new_[13997]_ ;
  assign \new_[2921]_  = \new_[13988]_  & \new_[13977]_ ;
  assign \new_[2922]_  = \new_[13968]_  & \new_[13957]_ ;
  assign \new_[2923]_  = \new_[13948]_  & \new_[13937]_ ;
  assign \new_[2924]_  = \new_[13928]_  & \new_[13917]_ ;
  assign \new_[2925]_  = \new_[13908]_  & \new_[13897]_ ;
  assign \new_[2926]_  = \new_[13888]_  & \new_[13877]_ ;
  assign \new_[2927]_  = \new_[13868]_  & \new_[13857]_ ;
  assign \new_[2928]_  = \new_[13848]_  & \new_[13837]_ ;
  assign \new_[2929]_  = \new_[13828]_  & \new_[13817]_ ;
  assign \new_[2930]_  = \new_[13808]_  & \new_[13797]_ ;
  assign \new_[2931]_  = \new_[13788]_  & \new_[13777]_ ;
  assign \new_[2932]_  = \new_[13768]_  & \new_[13757]_ ;
  assign \new_[2933]_  = \new_[13748]_  & \new_[13737]_ ;
  assign \new_[2934]_  = \new_[13728]_  & \new_[13717]_ ;
  assign \new_[2935]_  = \new_[13708]_  & \new_[13697]_ ;
  assign \new_[2936]_  = \new_[13688]_  & \new_[13677]_ ;
  assign \new_[2937]_  = \new_[13668]_  & \new_[13657]_ ;
  assign \new_[2938]_  = \new_[13648]_  & \new_[13637]_ ;
  assign \new_[2939]_  = \new_[13628]_  & \new_[13619]_ ;
  assign \new_[2940]_  = \new_[13610]_  & \new_[13601]_ ;
  assign \new_[2941]_  = \new_[13592]_  & \new_[13583]_ ;
  assign \new_[2942]_  = \new_[13574]_  & \new_[13565]_ ;
  assign \new_[2943]_  = \new_[13556]_  & \new_[13547]_ ;
  assign \new_[2944]_  = \new_[13538]_  & \new_[13529]_ ;
  assign \new_[2945]_  = \new_[13520]_  & \new_[13511]_ ;
  assign \new_[2946]_  = \new_[13502]_  & \new_[13493]_ ;
  assign \new_[2947]_  = \new_[13484]_  & \new_[13475]_ ;
  assign \new_[2948]_  = \new_[13466]_  & \new_[13457]_ ;
  assign \new_[2949]_  = \new_[13448]_  & \new_[13439]_ ;
  assign \new_[2950]_  = \new_[13430]_  & \new_[13421]_ ;
  assign \new_[2951]_  = \new_[13412]_  & \new_[13403]_ ;
  assign \new_[2952]_  = \new_[13394]_  & \new_[13385]_ ;
  assign \new_[2953]_  = \new_[13376]_  & \new_[13367]_ ;
  assign \new_[2954]_  = \new_[13358]_  & \new_[13349]_ ;
  assign \new_[2955]_  = \new_[13340]_  & \new_[13331]_ ;
  assign \new_[2956]_  = \new_[13322]_  & \new_[13313]_ ;
  assign \new_[2957]_  = \new_[13304]_  & \new_[13295]_ ;
  assign \new_[2958]_  = \new_[13286]_  & \new_[13277]_ ;
  assign \new_[2959]_  = \new_[13268]_  & \new_[13259]_ ;
  assign \new_[2960]_  = \new_[13250]_  & \new_[13241]_ ;
  assign \new_[2961]_  = \new_[13232]_  & \new_[13223]_ ;
  assign \new_[2962]_  = \new_[13214]_  & \new_[13205]_ ;
  assign \new_[2963]_  = \new_[13196]_  & \new_[13187]_ ;
  assign \new_[2964]_  = \new_[13178]_  & \new_[13169]_ ;
  assign \new_[2965]_  = \new_[13160]_  & \new_[13151]_ ;
  assign \new_[2966]_  = \new_[13142]_  & \new_[13133]_ ;
  assign \new_[2967]_  = \new_[13124]_  & \new_[13115]_ ;
  assign \new_[2968]_  = \new_[13106]_  & \new_[13097]_ ;
  assign \new_[2969]_  = \new_[13088]_  & \new_[13079]_ ;
  assign \new_[2970]_  = \new_[13070]_  & \new_[13061]_ ;
  assign \new_[2971]_  = \new_[13052]_  & \new_[13043]_ ;
  assign \new_[2972]_  = \new_[13034]_  & \new_[13025]_ ;
  assign \new_[2973]_  = \new_[13016]_  & \new_[13007]_ ;
  assign \new_[2974]_  = \new_[12998]_  & \new_[12989]_ ;
  assign \new_[2975]_  = \new_[12980]_  & \new_[12971]_ ;
  assign \new_[2976]_  = \new_[12962]_  & \new_[12953]_ ;
  assign \new_[2977]_  = \new_[12944]_  & \new_[12935]_ ;
  assign \new_[2978]_  = \new_[12926]_  & \new_[12917]_ ;
  assign \new_[2979]_  = \new_[12908]_  & \new_[12899]_ ;
  assign \new_[2980]_  = \new_[12890]_  & \new_[12881]_ ;
  assign \new_[2981]_  = \new_[12872]_  & \new_[12863]_ ;
  assign \new_[2982]_  = \new_[12854]_  & \new_[12845]_ ;
  assign \new_[2983]_  = \new_[12836]_  & \new_[12827]_ ;
  assign \new_[2984]_  = \new_[12818]_  & \new_[12809]_ ;
  assign \new_[2985]_  = \new_[12800]_  & \new_[12791]_ ;
  assign \new_[2986]_  = \new_[12782]_  & \new_[12773]_ ;
  assign \new_[2987]_  = \new_[12764]_  & \new_[12755]_ ;
  assign \new_[2988]_  = \new_[12746]_  & \new_[12737]_ ;
  assign \new_[2989]_  = \new_[12728]_  & \new_[12719]_ ;
  assign \new_[2990]_  = \new_[12710]_  & \new_[12701]_ ;
  assign \new_[2991]_  = \new_[12692]_  & \new_[12683]_ ;
  assign \new_[2992]_  = \new_[12674]_  & \new_[12665]_ ;
  assign \new_[2993]_  = \new_[12656]_  & \new_[12647]_ ;
  assign \new_[2994]_  = \new_[12638]_  & \new_[12629]_ ;
  assign \new_[2995]_  = \new_[12620]_  & \new_[12611]_ ;
  assign \new_[2996]_  = \new_[12602]_  & \new_[12593]_ ;
  assign \new_[2997]_  = \new_[12584]_  & \new_[12575]_ ;
  assign \new_[2998]_  = \new_[12566]_  & \new_[12557]_ ;
  assign \new_[2999]_  = \new_[12548]_  & \new_[12539]_ ;
  assign \new_[3000]_  = \new_[12530]_  & \new_[12521]_ ;
  assign \new_[3001]_  = \new_[12512]_  & \new_[12503]_ ;
  assign \new_[3002]_  = \new_[12494]_  & \new_[12485]_ ;
  assign \new_[3003]_  = \new_[12476]_  & \new_[12467]_ ;
  assign \new_[3004]_  = \new_[12458]_  & \new_[12449]_ ;
  assign \new_[3005]_  = \new_[12440]_  & \new_[12431]_ ;
  assign \new_[3006]_  = \new_[12422]_  & \new_[12413]_ ;
  assign \new_[3007]_  = \new_[12404]_  & \new_[12395]_ ;
  assign \new_[3008]_  = \new_[12386]_  & \new_[12377]_ ;
  assign \new_[3009]_  = \new_[12368]_  & \new_[12359]_ ;
  assign \new_[3010]_  = \new_[12350]_  & \new_[12341]_ ;
  assign \new_[3011]_  = \new_[12332]_  & \new_[12323]_ ;
  assign \new_[3012]_  = \new_[12314]_  & \new_[12305]_ ;
  assign \new_[3013]_  = \new_[12296]_  & \new_[12287]_ ;
  assign \new_[3014]_  = \new_[12278]_  & \new_[12269]_ ;
  assign \new_[3015]_  = \new_[12260]_  & \new_[12251]_ ;
  assign \new_[3016]_  = \new_[12242]_  & \new_[12233]_ ;
  assign \new_[3017]_  = \new_[12224]_  & \new_[12215]_ ;
  assign \new_[3018]_  = \new_[12206]_  & \new_[12197]_ ;
  assign \new_[3019]_  = \new_[12188]_  & \new_[12179]_ ;
  assign \new_[3020]_  = \new_[12170]_  & \new_[12161]_ ;
  assign \new_[3021]_  = \new_[12152]_  & \new_[12143]_ ;
  assign \new_[3022]_  = \new_[12134]_  & \new_[12125]_ ;
  assign \new_[3023]_  = \new_[12116]_  & \new_[12107]_ ;
  assign \new_[3024]_  = \new_[12098]_  & \new_[12089]_ ;
  assign \new_[3025]_  = \new_[12080]_  & \new_[12071]_ ;
  assign \new_[3026]_  = \new_[12062]_  & \new_[12053]_ ;
  assign \new_[3027]_  = \new_[12044]_  & \new_[12035]_ ;
  assign \new_[3028]_  = \new_[12026]_  & \new_[12017]_ ;
  assign \new_[3029]_  = \new_[12008]_  & \new_[11999]_ ;
  assign \new_[3030]_  = \new_[11990]_  & \new_[11981]_ ;
  assign \new_[3031]_  = \new_[11972]_  & \new_[11963]_ ;
  assign \new_[3032]_  = \new_[11954]_  & \new_[11945]_ ;
  assign \new_[3033]_  = \new_[11936]_  & \new_[11927]_ ;
  assign \new_[3034]_  = \new_[11918]_  & \new_[11909]_ ;
  assign \new_[3035]_  = \new_[11900]_  & \new_[11891]_ ;
  assign \new_[3036]_  = \new_[11882]_  & \new_[11873]_ ;
  assign \new_[3037]_  = \new_[11864]_  & \new_[11855]_ ;
  assign \new_[3038]_  = \new_[11846]_  & \new_[11837]_ ;
  assign \new_[3039]_  = \new_[11828]_  & \new_[11819]_ ;
  assign \new_[3040]_  = \new_[11810]_  & \new_[11801]_ ;
  assign \new_[3041]_  = \new_[11792]_  & \new_[11783]_ ;
  assign \new_[3042]_  = \new_[11774]_  & \new_[11765]_ ;
  assign \new_[3043]_  = \new_[11756]_  & \new_[11747]_ ;
  assign \new_[3044]_  = \new_[11738]_  & \new_[11729]_ ;
  assign \new_[3045]_  = \new_[11720]_  & \new_[11711]_ ;
  assign \new_[3046]_  = \new_[11702]_  & \new_[11693]_ ;
  assign \new_[3047]_  = \new_[11684]_  & \new_[11675]_ ;
  assign \new_[3048]_  = \new_[11666]_  & \new_[11657]_ ;
  assign \new_[3049]_  = \new_[11648]_  & \new_[11639]_ ;
  assign \new_[3050]_  = \new_[11630]_  & \new_[11621]_ ;
  assign \new_[3051]_  = \new_[11612]_  & \new_[11603]_ ;
  assign \new_[3052]_  = \new_[11594]_  & \new_[11585]_ ;
  assign \new_[3053]_  = \new_[11576]_  & \new_[11567]_ ;
  assign \new_[3054]_  = \new_[11558]_  & \new_[11549]_ ;
  assign \new_[3055]_  = \new_[11540]_  & \new_[11531]_ ;
  assign \new_[3056]_  = \new_[11522]_  & \new_[11513]_ ;
  assign \new_[3057]_  = \new_[11504]_  & \new_[11495]_ ;
  assign \new_[3058]_  = \new_[11486]_  & \new_[11477]_ ;
  assign \new_[3059]_  = \new_[11468]_  & \new_[11459]_ ;
  assign \new_[3060]_  = \new_[11450]_  & \new_[11441]_ ;
  assign \new_[3061]_  = \new_[11432]_  & \new_[11423]_ ;
  assign \new_[3062]_  = \new_[11414]_  & \new_[11405]_ ;
  assign \new_[3063]_  = \new_[11396]_  & \new_[11387]_ ;
  assign \new_[3064]_  = \new_[11378]_  & \new_[11369]_ ;
  assign \new_[3065]_  = \new_[11360]_  & \new_[11351]_ ;
  assign \new_[3066]_  = \new_[11342]_  & \new_[11333]_ ;
  assign \new_[3067]_  = \new_[11324]_  & \new_[11315]_ ;
  assign \new_[3068]_  = \new_[11306]_  & \new_[11297]_ ;
  assign \new_[3069]_  = \new_[11288]_  & \new_[11279]_ ;
  assign \new_[3070]_  = \new_[11270]_  & \new_[11261]_ ;
  assign \new_[3071]_  = \new_[11252]_  & \new_[11243]_ ;
  assign \new_[3072]_  = \new_[11234]_  & \new_[11225]_ ;
  assign \new_[3073]_  = \new_[11216]_  & \new_[11207]_ ;
  assign \new_[3074]_  = \new_[11198]_  & \new_[11189]_ ;
  assign \new_[3075]_  = \new_[11180]_  & \new_[11171]_ ;
  assign \new_[3076]_  = \new_[11162]_  & \new_[11153]_ ;
  assign \new_[3077]_  = \new_[11144]_  & \new_[11135]_ ;
  assign \new_[3078]_  = \new_[11126]_  & \new_[11117]_ ;
  assign \new_[3079]_  = \new_[11108]_  & \new_[11099]_ ;
  assign \new_[3080]_  = \new_[11090]_  & \new_[11081]_ ;
  assign \new_[3081]_  = \new_[11072]_  & \new_[11063]_ ;
  assign \new_[3082]_  = \new_[11054]_  & \new_[11045]_ ;
  assign \new_[3083]_  = \new_[11036]_  & \new_[11027]_ ;
  assign \new_[3084]_  = \new_[11018]_  & \new_[11009]_ ;
  assign \new_[3085]_  = \new_[11000]_  & \new_[10991]_ ;
  assign \new_[3086]_  = \new_[10982]_  & \new_[10973]_ ;
  assign \new_[3087]_  = \new_[10964]_  & \new_[10955]_ ;
  assign \new_[3088]_  = \new_[10946]_  & \new_[10937]_ ;
  assign \new_[3089]_  = \new_[10928]_  & \new_[10919]_ ;
  assign \new_[3090]_  = \new_[10910]_  & \new_[10901]_ ;
  assign \new_[3091]_  = \new_[10892]_  & \new_[10883]_ ;
  assign \new_[3092]_  = \new_[10874]_  & \new_[10865]_ ;
  assign \new_[3093]_  = \new_[10856]_  & \new_[10847]_ ;
  assign \new_[3094]_  = \new_[10838]_  & \new_[10829]_ ;
  assign \new_[3095]_  = \new_[10820]_  & \new_[10811]_ ;
  assign \new_[3096]_  = \new_[10802]_  & \new_[10793]_ ;
  assign \new_[3097]_  = \new_[10784]_  & \new_[10775]_ ;
  assign \new_[3098]_  = \new_[10766]_  & \new_[10757]_ ;
  assign \new_[3099]_  = \new_[10748]_  & \new_[10739]_ ;
  assign \new_[3100]_  = \new_[10730]_  & \new_[10721]_ ;
  assign \new_[3101]_  = \new_[10712]_  & \new_[10703]_ ;
  assign \new_[3102]_  = \new_[10694]_  & \new_[10685]_ ;
  assign \new_[3103]_  = \new_[10676]_  & \new_[10667]_ ;
  assign \new_[3104]_  = \new_[10658]_  & \new_[10649]_ ;
  assign \new_[3105]_  = \new_[10640]_  & \new_[10631]_ ;
  assign \new_[3106]_  = \new_[10622]_  & \new_[10613]_ ;
  assign \new_[3107]_  = \new_[10604]_  & \new_[10595]_ ;
  assign \new_[3108]_  = \new_[10586]_  & \new_[10577]_ ;
  assign \new_[3109]_  = \new_[10568]_  & \new_[10559]_ ;
  assign \new_[3110]_  = \new_[10550]_  & \new_[10541]_ ;
  assign \new_[3111]_  = \new_[10532]_  & \new_[10523]_ ;
  assign \new_[3112]_  = \new_[10514]_  & \new_[10505]_ ;
  assign \new_[3113]_  = \new_[10496]_  & \new_[10487]_ ;
  assign \new_[3114]_  = \new_[10478]_  & \new_[10469]_ ;
  assign \new_[3115]_  = \new_[10460]_  & \new_[10451]_ ;
  assign \new_[3116]_  = \new_[10442]_  & \new_[10433]_ ;
  assign \new_[3117]_  = \new_[10424]_  & \new_[10415]_ ;
  assign \new_[3118]_  = \new_[10406]_  & \new_[10397]_ ;
  assign \new_[3119]_  = \new_[10388]_  & \new_[10379]_ ;
  assign \new_[3120]_  = \new_[10370]_  & \new_[10361]_ ;
  assign \new_[3121]_  = \new_[10352]_  & \new_[10343]_ ;
  assign \new_[3122]_  = \new_[10334]_  & \new_[10325]_ ;
  assign \new_[3123]_  = \new_[10316]_  & \new_[10307]_ ;
  assign \new_[3124]_  = \new_[10298]_  & \new_[10289]_ ;
  assign \new_[3125]_  = \new_[10280]_  & \new_[10271]_ ;
  assign \new_[3126]_  = \new_[10262]_  & \new_[10253]_ ;
  assign \new_[3127]_  = \new_[10244]_  & \new_[10235]_ ;
  assign \new_[3128]_  = \new_[10226]_  & \new_[10217]_ ;
  assign \new_[3129]_  = \new_[10208]_  & \new_[10199]_ ;
  assign \new_[3130]_  = \new_[10192]_  & \new_[10183]_ ;
  assign \new_[3131]_  = \new_[10176]_  & \new_[10167]_ ;
  assign \new_[3132]_  = \new_[10160]_  & \new_[10151]_ ;
  assign \new_[3133]_  = \new_[10144]_  & \new_[10135]_ ;
  assign \new_[3134]_  = \new_[10128]_  & \new_[10119]_ ;
  assign \new_[3135]_  = \new_[10112]_  & \new_[10103]_ ;
  assign \new_[3136]_  = \new_[10096]_  & \new_[10087]_ ;
  assign \new_[3137]_  = \new_[10080]_  & \new_[10071]_ ;
  assign \new_[3138]_  = \new_[10064]_  & \new_[10055]_ ;
  assign \new_[3139]_  = \new_[10048]_  & \new_[10039]_ ;
  assign \new_[3140]_  = \new_[10032]_  & \new_[10023]_ ;
  assign \new_[3141]_  = \new_[10016]_  & \new_[10007]_ ;
  assign \new_[3142]_  = \new_[10000]_  & \new_[9991]_ ;
  assign \new_[3143]_  = \new_[9984]_  & \new_[9975]_ ;
  assign \new_[3144]_  = \new_[9968]_  & \new_[9959]_ ;
  assign \new_[3145]_  = \new_[9952]_  & \new_[9943]_ ;
  assign \new_[3146]_  = \new_[9936]_  & \new_[9927]_ ;
  assign \new_[3147]_  = \new_[9920]_  & \new_[9911]_ ;
  assign \new_[3148]_  = \new_[9904]_  & \new_[9895]_ ;
  assign \new_[3149]_  = \new_[9888]_  & \new_[9879]_ ;
  assign \new_[3150]_  = \new_[9872]_  & \new_[9863]_ ;
  assign \new_[3151]_  = \new_[9856]_  & \new_[9849]_ ;
  assign \new_[3152]_  = \new_[9842]_  & \new_[9835]_ ;
  assign \new_[3153]_  = \new_[9828]_  & \new_[9821]_ ;
  assign \new_[3154]_  = \new_[9814]_  & \new_[9807]_ ;
  assign \new_[3155]_  = \new_[9800]_  & \new_[9793]_ ;
  assign \new_[3156]_  = \new_[9786]_  & \new_[9779]_ ;
  assign \new_[3157]_  = \new_[9772]_  & \new_[9765]_ ;
  assign \new_[3158]_  = \new_[9758]_  & \new_[9751]_ ;
  assign \new_[3159]_  = \new_[9744]_  & \new_[9737]_ ;
  assign \new_[3160]_  = \new_[9730]_  & \new_[9723]_ ;
  assign \new_[3161]_  = \new_[9716]_  & \new_[9709]_ ;
  assign \new_[3162]_  = \new_[9702]_  & \new_[9695]_ ;
  assign \new_[3163]_  = \new_[9688]_  & \new_[9681]_ ;
  assign \new_[3164]_  = \new_[9674]_  & \new_[9667]_ ;
  assign \new_[3165]_  = \new_[9660]_  & \new_[9653]_ ;
  assign \new_[3166]_  = \new_[9646]_  & \new_[9639]_ ;
  assign \new_[3167]_  = \new_[9632]_  & \new_[9625]_ ;
  assign \new_[3168]_  = \new_[9618]_  & \new_[9611]_ ;
  assign \new_[3169]_  = \new_[9604]_  & \new_[9597]_ ;
  assign \new_[3170]_  = \new_[9590]_  & \new_[9583]_ ;
  assign \new_[3171]_  = \new_[9576]_  & \new_[9569]_ ;
  assign \new_[3172]_  = \new_[9562]_  & \new_[9555]_ ;
  assign \new_[3173]_  = \new_[9548]_  & \new_[9541]_ ;
  assign \new_[3174]_  = \new_[9534]_  & \new_[9527]_ ;
  assign \new_[3178]_  = \new_[3172]_  | \new_[3173]_ ;
  assign \new_[3179]_  = \new_[3174]_  | \new_[3178]_ ;
  assign \new_[3183]_  = \new_[3169]_  | \new_[3170]_ ;
  assign \new_[3184]_  = \new_[3171]_  | \new_[3183]_ ;
  assign \new_[3185]_  = \new_[3184]_  | \new_[3179]_ ;
  assign \new_[3189]_  = \new_[3166]_  | \new_[3167]_ ;
  assign \new_[3190]_  = \new_[3168]_  | \new_[3189]_ ;
  assign \new_[3194]_  = \new_[3163]_  | \new_[3164]_ ;
  assign \new_[3195]_  = \new_[3165]_  | \new_[3194]_ ;
  assign \new_[3196]_  = \new_[3195]_  | \new_[3190]_ ;
  assign \new_[3197]_  = \new_[3196]_  | \new_[3185]_ ;
  assign \new_[3201]_  = \new_[3160]_  | \new_[3161]_ ;
  assign \new_[3202]_  = \new_[3162]_  | \new_[3201]_ ;
  assign \new_[3206]_  = \new_[3157]_  | \new_[3158]_ ;
  assign \new_[3207]_  = \new_[3159]_  | \new_[3206]_ ;
  assign \new_[3208]_  = \new_[3207]_  | \new_[3202]_ ;
  assign \new_[3212]_  = \new_[3154]_  | \new_[3155]_ ;
  assign \new_[3213]_  = \new_[3156]_  | \new_[3212]_ ;
  assign \new_[3217]_  = \new_[3151]_  | \new_[3152]_ ;
  assign \new_[3218]_  = \new_[3153]_  | \new_[3217]_ ;
  assign \new_[3219]_  = \new_[3218]_  | \new_[3213]_ ;
  assign \new_[3220]_  = \new_[3219]_  | \new_[3208]_ ;
  assign \new_[3221]_  = \new_[3220]_  | \new_[3197]_ ;
  assign \new_[3225]_  = \new_[3148]_  | \new_[3149]_ ;
  assign \new_[3226]_  = \new_[3150]_  | \new_[3225]_ ;
  assign \new_[3230]_  = \new_[3145]_  | \new_[3146]_ ;
  assign \new_[3231]_  = \new_[3147]_  | \new_[3230]_ ;
  assign \new_[3232]_  = \new_[3231]_  | \new_[3226]_ ;
  assign \new_[3236]_  = \new_[3142]_  | \new_[3143]_ ;
  assign \new_[3237]_  = \new_[3144]_  | \new_[3236]_ ;
  assign \new_[3241]_  = \new_[3139]_  | \new_[3140]_ ;
  assign \new_[3242]_  = \new_[3141]_  | \new_[3241]_ ;
  assign \new_[3243]_  = \new_[3242]_  | \new_[3237]_ ;
  assign \new_[3244]_  = \new_[3243]_  | \new_[3232]_ ;
  assign \new_[3248]_  = \new_[3136]_  | \new_[3137]_ ;
  assign \new_[3249]_  = \new_[3138]_  | \new_[3248]_ ;
  assign \new_[3253]_  = \new_[3133]_  | \new_[3134]_ ;
  assign \new_[3254]_  = \new_[3135]_  | \new_[3253]_ ;
  assign \new_[3255]_  = \new_[3254]_  | \new_[3249]_ ;
  assign \new_[3259]_  = \new_[3130]_  | \new_[3131]_ ;
  assign \new_[3260]_  = \new_[3132]_  | \new_[3259]_ ;
  assign \new_[3263]_  = \new_[3128]_  | \new_[3129]_ ;
  assign \new_[3266]_  = \new_[3126]_  | \new_[3127]_ ;
  assign \new_[3267]_  = \new_[3266]_  | \new_[3263]_ ;
  assign \new_[3268]_  = \new_[3267]_  | \new_[3260]_ ;
  assign \new_[3269]_  = \new_[3268]_  | \new_[3255]_ ;
  assign \new_[3270]_  = \new_[3269]_  | \new_[3244]_ ;
  assign \new_[3271]_  = \new_[3270]_  | \new_[3221]_ ;
  assign \new_[3275]_  = \new_[3123]_  | \new_[3124]_ ;
  assign \new_[3276]_  = \new_[3125]_  | \new_[3275]_ ;
  assign \new_[3280]_  = \new_[3120]_  | \new_[3121]_ ;
  assign \new_[3281]_  = \new_[3122]_  | \new_[3280]_ ;
  assign \new_[3282]_  = \new_[3281]_  | \new_[3276]_ ;
  assign \new_[3286]_  = \new_[3117]_  | \new_[3118]_ ;
  assign \new_[3287]_  = \new_[3119]_  | \new_[3286]_ ;
  assign \new_[3291]_  = \new_[3114]_  | \new_[3115]_ ;
  assign \new_[3292]_  = \new_[3116]_  | \new_[3291]_ ;
  assign \new_[3293]_  = \new_[3292]_  | \new_[3287]_ ;
  assign \new_[3294]_  = \new_[3293]_  | \new_[3282]_ ;
  assign \new_[3298]_  = \new_[3111]_  | \new_[3112]_ ;
  assign \new_[3299]_  = \new_[3113]_  | \new_[3298]_ ;
  assign \new_[3303]_  = \new_[3108]_  | \new_[3109]_ ;
  assign \new_[3304]_  = \new_[3110]_  | \new_[3303]_ ;
  assign \new_[3305]_  = \new_[3304]_  | \new_[3299]_ ;
  assign \new_[3309]_  = \new_[3105]_  | \new_[3106]_ ;
  assign \new_[3310]_  = \new_[3107]_  | \new_[3309]_ ;
  assign \new_[3313]_  = \new_[3103]_  | \new_[3104]_ ;
  assign \new_[3316]_  = \new_[3101]_  | \new_[3102]_ ;
  assign \new_[3317]_  = \new_[3316]_  | \new_[3313]_ ;
  assign \new_[3318]_  = \new_[3317]_  | \new_[3310]_ ;
  assign \new_[3319]_  = \new_[3318]_  | \new_[3305]_ ;
  assign \new_[3320]_  = \new_[3319]_  | \new_[3294]_ ;
  assign \new_[3324]_  = \new_[3098]_  | \new_[3099]_ ;
  assign \new_[3325]_  = \new_[3100]_  | \new_[3324]_ ;
  assign \new_[3329]_  = \new_[3095]_  | \new_[3096]_ ;
  assign \new_[3330]_  = \new_[3097]_  | \new_[3329]_ ;
  assign \new_[3331]_  = \new_[3330]_  | \new_[3325]_ ;
  assign \new_[3335]_  = \new_[3092]_  | \new_[3093]_ ;
  assign \new_[3336]_  = \new_[3094]_  | \new_[3335]_ ;
  assign \new_[3340]_  = \new_[3089]_  | \new_[3090]_ ;
  assign \new_[3341]_  = \new_[3091]_  | \new_[3340]_ ;
  assign \new_[3342]_  = \new_[3341]_  | \new_[3336]_ ;
  assign \new_[3343]_  = \new_[3342]_  | \new_[3331]_ ;
  assign \new_[3347]_  = \new_[3086]_  | \new_[3087]_ ;
  assign \new_[3348]_  = \new_[3088]_  | \new_[3347]_ ;
  assign \new_[3352]_  = \new_[3083]_  | \new_[3084]_ ;
  assign \new_[3353]_  = \new_[3085]_  | \new_[3352]_ ;
  assign \new_[3354]_  = \new_[3353]_  | \new_[3348]_ ;
  assign \new_[3358]_  = \new_[3080]_  | \new_[3081]_ ;
  assign \new_[3359]_  = \new_[3082]_  | \new_[3358]_ ;
  assign \new_[3362]_  = \new_[3078]_  | \new_[3079]_ ;
  assign \new_[3365]_  = \new_[3076]_  | \new_[3077]_ ;
  assign \new_[3366]_  = \new_[3365]_  | \new_[3362]_ ;
  assign \new_[3367]_  = \new_[3366]_  | \new_[3359]_ ;
  assign \new_[3368]_  = \new_[3367]_  | \new_[3354]_ ;
  assign \new_[3369]_  = \new_[3368]_  | \new_[3343]_ ;
  assign \new_[3370]_  = \new_[3369]_  | \new_[3320]_ ;
  assign \new_[3371]_  = \new_[3370]_  | \new_[3271]_ ;
  assign \new_[3375]_  = \new_[3073]_  | \new_[3074]_ ;
  assign \new_[3376]_  = \new_[3075]_  | \new_[3375]_ ;
  assign \new_[3380]_  = \new_[3070]_  | \new_[3071]_ ;
  assign \new_[3381]_  = \new_[3072]_  | \new_[3380]_ ;
  assign \new_[3382]_  = \new_[3381]_  | \new_[3376]_ ;
  assign \new_[3386]_  = \new_[3067]_  | \new_[3068]_ ;
  assign \new_[3387]_  = \new_[3069]_  | \new_[3386]_ ;
  assign \new_[3391]_  = \new_[3064]_  | \new_[3065]_ ;
  assign \new_[3392]_  = \new_[3066]_  | \new_[3391]_ ;
  assign \new_[3393]_  = \new_[3392]_  | \new_[3387]_ ;
  assign \new_[3394]_  = \new_[3393]_  | \new_[3382]_ ;
  assign \new_[3398]_  = \new_[3061]_  | \new_[3062]_ ;
  assign \new_[3399]_  = \new_[3063]_  | \new_[3398]_ ;
  assign \new_[3403]_  = \new_[3058]_  | \new_[3059]_ ;
  assign \new_[3404]_  = \new_[3060]_  | \new_[3403]_ ;
  assign \new_[3405]_  = \new_[3404]_  | \new_[3399]_ ;
  assign \new_[3409]_  = \new_[3055]_  | \new_[3056]_ ;
  assign \new_[3410]_  = \new_[3057]_  | \new_[3409]_ ;
  assign \new_[3414]_  = \new_[3052]_  | \new_[3053]_ ;
  assign \new_[3415]_  = \new_[3054]_  | \new_[3414]_ ;
  assign \new_[3416]_  = \new_[3415]_  | \new_[3410]_ ;
  assign \new_[3417]_  = \new_[3416]_  | \new_[3405]_ ;
  assign \new_[3418]_  = \new_[3417]_  | \new_[3394]_ ;
  assign \new_[3422]_  = \new_[3049]_  | \new_[3050]_ ;
  assign \new_[3423]_  = \new_[3051]_  | \new_[3422]_ ;
  assign \new_[3427]_  = \new_[3046]_  | \new_[3047]_ ;
  assign \new_[3428]_  = \new_[3048]_  | \new_[3427]_ ;
  assign \new_[3429]_  = \new_[3428]_  | \new_[3423]_ ;
  assign \new_[3433]_  = \new_[3043]_  | \new_[3044]_ ;
  assign \new_[3434]_  = \new_[3045]_  | \new_[3433]_ ;
  assign \new_[3438]_  = \new_[3040]_  | \new_[3041]_ ;
  assign \new_[3439]_  = \new_[3042]_  | \new_[3438]_ ;
  assign \new_[3440]_  = \new_[3439]_  | \new_[3434]_ ;
  assign \new_[3441]_  = \new_[3440]_  | \new_[3429]_ ;
  assign \new_[3445]_  = \new_[3037]_  | \new_[3038]_ ;
  assign \new_[3446]_  = \new_[3039]_  | \new_[3445]_ ;
  assign \new_[3450]_  = \new_[3034]_  | \new_[3035]_ ;
  assign \new_[3451]_  = \new_[3036]_  | \new_[3450]_ ;
  assign \new_[3452]_  = \new_[3451]_  | \new_[3446]_ ;
  assign \new_[3456]_  = \new_[3031]_  | \new_[3032]_ ;
  assign \new_[3457]_  = \new_[3033]_  | \new_[3456]_ ;
  assign \new_[3460]_  = \new_[3029]_  | \new_[3030]_ ;
  assign \new_[3463]_  = \new_[3027]_  | \new_[3028]_ ;
  assign \new_[3464]_  = \new_[3463]_  | \new_[3460]_ ;
  assign \new_[3465]_  = \new_[3464]_  | \new_[3457]_ ;
  assign \new_[3466]_  = \new_[3465]_  | \new_[3452]_ ;
  assign \new_[3467]_  = \new_[3466]_  | \new_[3441]_ ;
  assign \new_[3468]_  = \new_[3467]_  | \new_[3418]_ ;
  assign \new_[3472]_  = \new_[3024]_  | \new_[3025]_ ;
  assign \new_[3473]_  = \new_[3026]_  | \new_[3472]_ ;
  assign \new_[3477]_  = \new_[3021]_  | \new_[3022]_ ;
  assign \new_[3478]_  = \new_[3023]_  | \new_[3477]_ ;
  assign \new_[3479]_  = \new_[3478]_  | \new_[3473]_ ;
  assign \new_[3483]_  = \new_[3018]_  | \new_[3019]_ ;
  assign \new_[3484]_  = \new_[3020]_  | \new_[3483]_ ;
  assign \new_[3488]_  = \new_[3015]_  | \new_[3016]_ ;
  assign \new_[3489]_  = \new_[3017]_  | \new_[3488]_ ;
  assign \new_[3490]_  = \new_[3489]_  | \new_[3484]_ ;
  assign \new_[3491]_  = \new_[3490]_  | \new_[3479]_ ;
  assign \new_[3495]_  = \new_[3012]_  | \new_[3013]_ ;
  assign \new_[3496]_  = \new_[3014]_  | \new_[3495]_ ;
  assign \new_[3500]_  = \new_[3009]_  | \new_[3010]_ ;
  assign \new_[3501]_  = \new_[3011]_  | \new_[3500]_ ;
  assign \new_[3502]_  = \new_[3501]_  | \new_[3496]_ ;
  assign \new_[3506]_  = \new_[3006]_  | \new_[3007]_ ;
  assign \new_[3507]_  = \new_[3008]_  | \new_[3506]_ ;
  assign \new_[3510]_  = \new_[3004]_  | \new_[3005]_ ;
  assign \new_[3513]_  = \new_[3002]_  | \new_[3003]_ ;
  assign \new_[3514]_  = \new_[3513]_  | \new_[3510]_ ;
  assign \new_[3515]_  = \new_[3514]_  | \new_[3507]_ ;
  assign \new_[3516]_  = \new_[3515]_  | \new_[3502]_ ;
  assign \new_[3517]_  = \new_[3516]_  | \new_[3491]_ ;
  assign \new_[3521]_  = \new_[2999]_  | \new_[3000]_ ;
  assign \new_[3522]_  = \new_[3001]_  | \new_[3521]_ ;
  assign \new_[3526]_  = \new_[2996]_  | \new_[2997]_ ;
  assign \new_[3527]_  = \new_[2998]_  | \new_[3526]_ ;
  assign \new_[3528]_  = \new_[3527]_  | \new_[3522]_ ;
  assign \new_[3532]_  = \new_[2993]_  | \new_[2994]_ ;
  assign \new_[3533]_  = \new_[2995]_  | \new_[3532]_ ;
  assign \new_[3537]_  = \new_[2990]_  | \new_[2991]_ ;
  assign \new_[3538]_  = \new_[2992]_  | \new_[3537]_ ;
  assign \new_[3539]_  = \new_[3538]_  | \new_[3533]_ ;
  assign \new_[3540]_  = \new_[3539]_  | \new_[3528]_ ;
  assign \new_[3544]_  = \new_[2987]_  | \new_[2988]_ ;
  assign \new_[3545]_  = \new_[2989]_  | \new_[3544]_ ;
  assign \new_[3549]_  = \new_[2984]_  | \new_[2985]_ ;
  assign \new_[3550]_  = \new_[2986]_  | \new_[3549]_ ;
  assign \new_[3551]_  = \new_[3550]_  | \new_[3545]_ ;
  assign \new_[3555]_  = \new_[2981]_  | \new_[2982]_ ;
  assign \new_[3556]_  = \new_[2983]_  | \new_[3555]_ ;
  assign \new_[3559]_  = \new_[2979]_  | \new_[2980]_ ;
  assign \new_[3562]_  = \new_[2977]_  | \new_[2978]_ ;
  assign \new_[3563]_  = \new_[3562]_  | \new_[3559]_ ;
  assign \new_[3564]_  = \new_[3563]_  | \new_[3556]_ ;
  assign \new_[3565]_  = \new_[3564]_  | \new_[3551]_ ;
  assign \new_[3566]_  = \new_[3565]_  | \new_[3540]_ ;
  assign \new_[3567]_  = \new_[3566]_  | \new_[3517]_ ;
  assign \new_[3568]_  = \new_[3567]_  | \new_[3468]_ ;
  assign \new_[3569]_  = \new_[3568]_  | \new_[3371]_ ;
  assign \new_[3573]_  = \new_[2974]_  | \new_[2975]_ ;
  assign \new_[3574]_  = \new_[2976]_  | \new_[3573]_ ;
  assign \new_[3578]_  = \new_[2971]_  | \new_[2972]_ ;
  assign \new_[3579]_  = \new_[2973]_  | \new_[3578]_ ;
  assign \new_[3580]_  = \new_[3579]_  | \new_[3574]_ ;
  assign \new_[3584]_  = \new_[2968]_  | \new_[2969]_ ;
  assign \new_[3585]_  = \new_[2970]_  | \new_[3584]_ ;
  assign \new_[3589]_  = \new_[2965]_  | \new_[2966]_ ;
  assign \new_[3590]_  = \new_[2967]_  | \new_[3589]_ ;
  assign \new_[3591]_  = \new_[3590]_  | \new_[3585]_ ;
  assign \new_[3592]_  = \new_[3591]_  | \new_[3580]_ ;
  assign \new_[3596]_  = \new_[2962]_  | \new_[2963]_ ;
  assign \new_[3597]_  = \new_[2964]_  | \new_[3596]_ ;
  assign \new_[3601]_  = \new_[2959]_  | \new_[2960]_ ;
  assign \new_[3602]_  = \new_[2961]_  | \new_[3601]_ ;
  assign \new_[3603]_  = \new_[3602]_  | \new_[3597]_ ;
  assign \new_[3607]_  = \new_[2956]_  | \new_[2957]_ ;
  assign \new_[3608]_  = \new_[2958]_  | \new_[3607]_ ;
  assign \new_[3612]_  = \new_[2953]_  | \new_[2954]_ ;
  assign \new_[3613]_  = \new_[2955]_  | \new_[3612]_ ;
  assign \new_[3614]_  = \new_[3613]_  | \new_[3608]_ ;
  assign \new_[3615]_  = \new_[3614]_  | \new_[3603]_ ;
  assign \new_[3616]_  = \new_[3615]_  | \new_[3592]_ ;
  assign \new_[3620]_  = \new_[2950]_  | \new_[2951]_ ;
  assign \new_[3621]_  = \new_[2952]_  | \new_[3620]_ ;
  assign \new_[3625]_  = \new_[2947]_  | \new_[2948]_ ;
  assign \new_[3626]_  = \new_[2949]_  | \new_[3625]_ ;
  assign \new_[3627]_  = \new_[3626]_  | \new_[3621]_ ;
  assign \new_[3631]_  = \new_[2944]_  | \new_[2945]_ ;
  assign \new_[3632]_  = \new_[2946]_  | \new_[3631]_ ;
  assign \new_[3636]_  = \new_[2941]_  | \new_[2942]_ ;
  assign \new_[3637]_  = \new_[2943]_  | \new_[3636]_ ;
  assign \new_[3638]_  = \new_[3637]_  | \new_[3632]_ ;
  assign \new_[3639]_  = \new_[3638]_  | \new_[3627]_ ;
  assign \new_[3643]_  = \new_[2938]_  | \new_[2939]_ ;
  assign \new_[3644]_  = \new_[2940]_  | \new_[3643]_ ;
  assign \new_[3648]_  = \new_[2935]_  | \new_[2936]_ ;
  assign \new_[3649]_  = \new_[2937]_  | \new_[3648]_ ;
  assign \new_[3650]_  = \new_[3649]_  | \new_[3644]_ ;
  assign \new_[3654]_  = \new_[2932]_  | \new_[2933]_ ;
  assign \new_[3655]_  = \new_[2934]_  | \new_[3654]_ ;
  assign \new_[3658]_  = \new_[2930]_  | \new_[2931]_ ;
  assign \new_[3661]_  = \new_[2928]_  | \new_[2929]_ ;
  assign \new_[3662]_  = \new_[3661]_  | \new_[3658]_ ;
  assign \new_[3663]_  = \new_[3662]_  | \new_[3655]_ ;
  assign \new_[3664]_  = \new_[3663]_  | \new_[3650]_ ;
  assign \new_[3665]_  = \new_[3664]_  | \new_[3639]_ ;
  assign \new_[3666]_  = \new_[3665]_  | \new_[3616]_ ;
  assign \new_[3670]_  = \new_[2925]_  | \new_[2926]_ ;
  assign \new_[3671]_  = \new_[2927]_  | \new_[3670]_ ;
  assign \new_[3675]_  = \new_[2922]_  | \new_[2923]_ ;
  assign \new_[3676]_  = \new_[2924]_  | \new_[3675]_ ;
  assign \new_[3677]_  = \new_[3676]_  | \new_[3671]_ ;
  assign \new_[3681]_  = \new_[2919]_  | \new_[2920]_ ;
  assign \new_[3682]_  = \new_[2921]_  | \new_[3681]_ ;
  assign \new_[3686]_  = \new_[2916]_  | \new_[2917]_ ;
  assign \new_[3687]_  = \new_[2918]_  | \new_[3686]_ ;
  assign \new_[3688]_  = \new_[3687]_  | \new_[3682]_ ;
  assign \new_[3689]_  = \new_[3688]_  | \new_[3677]_ ;
  assign \new_[3693]_  = \new_[2913]_  | \new_[2914]_ ;
  assign \new_[3694]_  = \new_[2915]_  | \new_[3693]_ ;
  assign \new_[3698]_  = \new_[2910]_  | \new_[2911]_ ;
  assign \new_[3699]_  = \new_[2912]_  | \new_[3698]_ ;
  assign \new_[3700]_  = \new_[3699]_  | \new_[3694]_ ;
  assign \new_[3704]_  = \new_[2907]_  | \new_[2908]_ ;
  assign \new_[3705]_  = \new_[2909]_  | \new_[3704]_ ;
  assign \new_[3708]_  = \new_[2905]_  | \new_[2906]_ ;
  assign \new_[3711]_  = \new_[2903]_  | \new_[2904]_ ;
  assign \new_[3712]_  = \new_[3711]_  | \new_[3708]_ ;
  assign \new_[3713]_  = \new_[3712]_  | \new_[3705]_ ;
  assign \new_[3714]_  = \new_[3713]_  | \new_[3700]_ ;
  assign \new_[3715]_  = \new_[3714]_  | \new_[3689]_ ;
  assign \new_[3719]_  = \new_[2900]_  | \new_[2901]_ ;
  assign \new_[3720]_  = \new_[2902]_  | \new_[3719]_ ;
  assign \new_[3724]_  = \new_[2897]_  | \new_[2898]_ ;
  assign \new_[3725]_  = \new_[2899]_  | \new_[3724]_ ;
  assign \new_[3726]_  = \new_[3725]_  | \new_[3720]_ ;
  assign \new_[3730]_  = \new_[2894]_  | \new_[2895]_ ;
  assign \new_[3731]_  = \new_[2896]_  | \new_[3730]_ ;
  assign \new_[3735]_  = \new_[2891]_  | \new_[2892]_ ;
  assign \new_[3736]_  = \new_[2893]_  | \new_[3735]_ ;
  assign \new_[3737]_  = \new_[3736]_  | \new_[3731]_ ;
  assign \new_[3738]_  = \new_[3737]_  | \new_[3726]_ ;
  assign \new_[3742]_  = \new_[2888]_  | \new_[2889]_ ;
  assign \new_[3743]_  = \new_[2890]_  | \new_[3742]_ ;
  assign \new_[3747]_  = \new_[2885]_  | \new_[2886]_ ;
  assign \new_[3748]_  = \new_[2887]_  | \new_[3747]_ ;
  assign \new_[3749]_  = \new_[3748]_  | \new_[3743]_ ;
  assign \new_[3753]_  = \new_[2882]_  | \new_[2883]_ ;
  assign \new_[3754]_  = \new_[2884]_  | \new_[3753]_ ;
  assign \new_[3757]_  = \new_[2880]_  | \new_[2881]_ ;
  assign \new_[3760]_  = \new_[2878]_  | \new_[2879]_ ;
  assign \new_[3761]_  = \new_[3760]_  | \new_[3757]_ ;
  assign \new_[3762]_  = \new_[3761]_  | \new_[3754]_ ;
  assign \new_[3763]_  = \new_[3762]_  | \new_[3749]_ ;
  assign \new_[3764]_  = \new_[3763]_  | \new_[3738]_ ;
  assign \new_[3765]_  = \new_[3764]_  | \new_[3715]_ ;
  assign \new_[3766]_  = \new_[3765]_  | \new_[3666]_ ;
  assign \new_[3770]_  = \new_[2875]_  | \new_[2876]_ ;
  assign \new_[3771]_  = \new_[2877]_  | \new_[3770]_ ;
  assign \new_[3775]_  = \new_[2872]_  | \new_[2873]_ ;
  assign \new_[3776]_  = \new_[2874]_  | \new_[3775]_ ;
  assign \new_[3777]_  = \new_[3776]_  | \new_[3771]_ ;
  assign \new_[3781]_  = \new_[2869]_  | \new_[2870]_ ;
  assign \new_[3782]_  = \new_[2871]_  | \new_[3781]_ ;
  assign \new_[3786]_  = \new_[2866]_  | \new_[2867]_ ;
  assign \new_[3787]_  = \new_[2868]_  | \new_[3786]_ ;
  assign \new_[3788]_  = \new_[3787]_  | \new_[3782]_ ;
  assign \new_[3789]_  = \new_[3788]_  | \new_[3777]_ ;
  assign \new_[3793]_  = \new_[2863]_  | \new_[2864]_ ;
  assign \new_[3794]_  = \new_[2865]_  | \new_[3793]_ ;
  assign \new_[3798]_  = \new_[2860]_  | \new_[2861]_ ;
  assign \new_[3799]_  = \new_[2862]_  | \new_[3798]_ ;
  assign \new_[3800]_  = \new_[3799]_  | \new_[3794]_ ;
  assign \new_[3804]_  = \new_[2857]_  | \new_[2858]_ ;
  assign \new_[3805]_  = \new_[2859]_  | \new_[3804]_ ;
  assign \new_[3809]_  = \new_[2854]_  | \new_[2855]_ ;
  assign \new_[3810]_  = \new_[2856]_  | \new_[3809]_ ;
  assign \new_[3811]_  = \new_[3810]_  | \new_[3805]_ ;
  assign \new_[3812]_  = \new_[3811]_  | \new_[3800]_ ;
  assign \new_[3813]_  = \new_[3812]_  | \new_[3789]_ ;
  assign \new_[3817]_  = \new_[2851]_  | \new_[2852]_ ;
  assign \new_[3818]_  = \new_[2853]_  | \new_[3817]_ ;
  assign \new_[3822]_  = \new_[2848]_  | \new_[2849]_ ;
  assign \new_[3823]_  = \new_[2850]_  | \new_[3822]_ ;
  assign \new_[3824]_  = \new_[3823]_  | \new_[3818]_ ;
  assign \new_[3828]_  = \new_[2845]_  | \new_[2846]_ ;
  assign \new_[3829]_  = \new_[2847]_  | \new_[3828]_ ;
  assign \new_[3833]_  = \new_[2842]_  | \new_[2843]_ ;
  assign \new_[3834]_  = \new_[2844]_  | \new_[3833]_ ;
  assign \new_[3835]_  = \new_[3834]_  | \new_[3829]_ ;
  assign \new_[3836]_  = \new_[3835]_  | \new_[3824]_ ;
  assign \new_[3840]_  = \new_[2839]_  | \new_[2840]_ ;
  assign \new_[3841]_  = \new_[2841]_  | \new_[3840]_ ;
  assign \new_[3845]_  = \new_[2836]_  | \new_[2837]_ ;
  assign \new_[3846]_  = \new_[2838]_  | \new_[3845]_ ;
  assign \new_[3847]_  = \new_[3846]_  | \new_[3841]_ ;
  assign \new_[3851]_  = \new_[2833]_  | \new_[2834]_ ;
  assign \new_[3852]_  = \new_[2835]_  | \new_[3851]_ ;
  assign \new_[3855]_  = \new_[2831]_  | \new_[2832]_ ;
  assign \new_[3858]_  = \new_[2829]_  | \new_[2830]_ ;
  assign \new_[3859]_  = \new_[3858]_  | \new_[3855]_ ;
  assign \new_[3860]_  = \new_[3859]_  | \new_[3852]_ ;
  assign \new_[3861]_  = \new_[3860]_  | \new_[3847]_ ;
  assign \new_[3862]_  = \new_[3861]_  | \new_[3836]_ ;
  assign \new_[3863]_  = \new_[3862]_  | \new_[3813]_ ;
  assign \new_[3867]_  = \new_[2826]_  | \new_[2827]_ ;
  assign \new_[3868]_  = \new_[2828]_  | \new_[3867]_ ;
  assign \new_[3872]_  = \new_[2823]_  | \new_[2824]_ ;
  assign \new_[3873]_  = \new_[2825]_  | \new_[3872]_ ;
  assign \new_[3874]_  = \new_[3873]_  | \new_[3868]_ ;
  assign \new_[3878]_  = \new_[2820]_  | \new_[2821]_ ;
  assign \new_[3879]_  = \new_[2822]_  | \new_[3878]_ ;
  assign \new_[3883]_  = \new_[2817]_  | \new_[2818]_ ;
  assign \new_[3884]_  = \new_[2819]_  | \new_[3883]_ ;
  assign \new_[3885]_  = \new_[3884]_  | \new_[3879]_ ;
  assign \new_[3886]_  = \new_[3885]_  | \new_[3874]_ ;
  assign \new_[3890]_  = \new_[2814]_  | \new_[2815]_ ;
  assign \new_[3891]_  = \new_[2816]_  | \new_[3890]_ ;
  assign \new_[3895]_  = \new_[2811]_  | \new_[2812]_ ;
  assign \new_[3896]_  = \new_[2813]_  | \new_[3895]_ ;
  assign \new_[3897]_  = \new_[3896]_  | \new_[3891]_ ;
  assign \new_[3901]_  = \new_[2808]_  | \new_[2809]_ ;
  assign \new_[3902]_  = \new_[2810]_  | \new_[3901]_ ;
  assign \new_[3905]_  = \new_[2806]_  | \new_[2807]_ ;
  assign \new_[3908]_  = \new_[2804]_  | \new_[2805]_ ;
  assign \new_[3909]_  = \new_[3908]_  | \new_[3905]_ ;
  assign \new_[3910]_  = \new_[3909]_  | \new_[3902]_ ;
  assign \new_[3911]_  = \new_[3910]_  | \new_[3897]_ ;
  assign \new_[3912]_  = \new_[3911]_  | \new_[3886]_ ;
  assign \new_[3916]_  = \new_[2801]_  | \new_[2802]_ ;
  assign \new_[3917]_  = \new_[2803]_  | \new_[3916]_ ;
  assign \new_[3921]_  = \new_[2798]_  | \new_[2799]_ ;
  assign \new_[3922]_  = \new_[2800]_  | \new_[3921]_ ;
  assign \new_[3923]_  = \new_[3922]_  | \new_[3917]_ ;
  assign \new_[3927]_  = \new_[2795]_  | \new_[2796]_ ;
  assign \new_[3928]_  = \new_[2797]_  | \new_[3927]_ ;
  assign \new_[3932]_  = \new_[2792]_  | \new_[2793]_ ;
  assign \new_[3933]_  = \new_[2794]_  | \new_[3932]_ ;
  assign \new_[3934]_  = \new_[3933]_  | \new_[3928]_ ;
  assign \new_[3935]_  = \new_[3934]_  | \new_[3923]_ ;
  assign \new_[3939]_  = \new_[2789]_  | \new_[2790]_ ;
  assign \new_[3940]_  = \new_[2791]_  | \new_[3939]_ ;
  assign \new_[3944]_  = \new_[2786]_  | \new_[2787]_ ;
  assign \new_[3945]_  = \new_[2788]_  | \new_[3944]_ ;
  assign \new_[3946]_  = \new_[3945]_  | \new_[3940]_ ;
  assign \new_[3950]_  = \new_[2783]_  | \new_[2784]_ ;
  assign \new_[3951]_  = \new_[2785]_  | \new_[3950]_ ;
  assign \new_[3954]_  = \new_[2781]_  | \new_[2782]_ ;
  assign \new_[3957]_  = \new_[2779]_  | \new_[2780]_ ;
  assign \new_[3958]_  = \new_[3957]_  | \new_[3954]_ ;
  assign \new_[3959]_  = \new_[3958]_  | \new_[3951]_ ;
  assign \new_[3960]_  = \new_[3959]_  | \new_[3946]_ ;
  assign \new_[3961]_  = \new_[3960]_  | \new_[3935]_ ;
  assign \new_[3962]_  = \new_[3961]_  | \new_[3912]_ ;
  assign \new_[3963]_  = \new_[3962]_  | \new_[3863]_ ;
  assign \new_[3964]_  = \new_[3963]_  | \new_[3766]_ ;
  assign \new_[3965]_  = \new_[3964]_  | \new_[3569]_ ;
  assign \new_[3969]_  = \new_[2776]_  | \new_[2777]_ ;
  assign \new_[3970]_  = \new_[2778]_  | \new_[3969]_ ;
  assign \new_[3974]_  = \new_[2773]_  | \new_[2774]_ ;
  assign \new_[3975]_  = \new_[2775]_  | \new_[3974]_ ;
  assign \new_[3976]_  = \new_[3975]_  | \new_[3970]_ ;
  assign \new_[3980]_  = \new_[2770]_  | \new_[2771]_ ;
  assign \new_[3981]_  = \new_[2772]_  | \new_[3980]_ ;
  assign \new_[3985]_  = \new_[2767]_  | \new_[2768]_ ;
  assign \new_[3986]_  = \new_[2769]_  | \new_[3985]_ ;
  assign \new_[3987]_  = \new_[3986]_  | \new_[3981]_ ;
  assign \new_[3988]_  = \new_[3987]_  | \new_[3976]_ ;
  assign \new_[3992]_  = \new_[2764]_  | \new_[2765]_ ;
  assign \new_[3993]_  = \new_[2766]_  | \new_[3992]_ ;
  assign \new_[3997]_  = \new_[2761]_  | \new_[2762]_ ;
  assign \new_[3998]_  = \new_[2763]_  | \new_[3997]_ ;
  assign \new_[3999]_  = \new_[3998]_  | \new_[3993]_ ;
  assign \new_[4003]_  = \new_[2758]_  | \new_[2759]_ ;
  assign \new_[4004]_  = \new_[2760]_  | \new_[4003]_ ;
  assign \new_[4008]_  = \new_[2755]_  | \new_[2756]_ ;
  assign \new_[4009]_  = \new_[2757]_  | \new_[4008]_ ;
  assign \new_[4010]_  = \new_[4009]_  | \new_[4004]_ ;
  assign \new_[4011]_  = \new_[4010]_  | \new_[3999]_ ;
  assign \new_[4012]_  = \new_[4011]_  | \new_[3988]_ ;
  assign \new_[4016]_  = \new_[2752]_  | \new_[2753]_ ;
  assign \new_[4017]_  = \new_[2754]_  | \new_[4016]_ ;
  assign \new_[4021]_  = \new_[2749]_  | \new_[2750]_ ;
  assign \new_[4022]_  = \new_[2751]_  | \new_[4021]_ ;
  assign \new_[4023]_  = \new_[4022]_  | \new_[4017]_ ;
  assign \new_[4027]_  = \new_[2746]_  | \new_[2747]_ ;
  assign \new_[4028]_  = \new_[2748]_  | \new_[4027]_ ;
  assign \new_[4032]_  = \new_[2743]_  | \new_[2744]_ ;
  assign \new_[4033]_  = \new_[2745]_  | \new_[4032]_ ;
  assign \new_[4034]_  = \new_[4033]_  | \new_[4028]_ ;
  assign \new_[4035]_  = \new_[4034]_  | \new_[4023]_ ;
  assign \new_[4039]_  = \new_[2740]_  | \new_[2741]_ ;
  assign \new_[4040]_  = \new_[2742]_  | \new_[4039]_ ;
  assign \new_[4044]_  = \new_[2737]_  | \new_[2738]_ ;
  assign \new_[4045]_  = \new_[2739]_  | \new_[4044]_ ;
  assign \new_[4046]_  = \new_[4045]_  | \new_[4040]_ ;
  assign \new_[4050]_  = \new_[2734]_  | \new_[2735]_ ;
  assign \new_[4051]_  = \new_[2736]_  | \new_[4050]_ ;
  assign \new_[4054]_  = \new_[2732]_  | \new_[2733]_ ;
  assign \new_[4057]_  = \new_[2730]_  | \new_[2731]_ ;
  assign \new_[4058]_  = \new_[4057]_  | \new_[4054]_ ;
  assign \new_[4059]_  = \new_[4058]_  | \new_[4051]_ ;
  assign \new_[4060]_  = \new_[4059]_  | \new_[4046]_ ;
  assign \new_[4061]_  = \new_[4060]_  | \new_[4035]_ ;
  assign \new_[4062]_  = \new_[4061]_  | \new_[4012]_ ;
  assign \new_[4066]_  = \new_[2727]_  | \new_[2728]_ ;
  assign \new_[4067]_  = \new_[2729]_  | \new_[4066]_ ;
  assign \new_[4071]_  = \new_[2724]_  | \new_[2725]_ ;
  assign \new_[4072]_  = \new_[2726]_  | \new_[4071]_ ;
  assign \new_[4073]_  = \new_[4072]_  | \new_[4067]_ ;
  assign \new_[4077]_  = \new_[2721]_  | \new_[2722]_ ;
  assign \new_[4078]_  = \new_[2723]_  | \new_[4077]_ ;
  assign \new_[4082]_  = \new_[2718]_  | \new_[2719]_ ;
  assign \new_[4083]_  = \new_[2720]_  | \new_[4082]_ ;
  assign \new_[4084]_  = \new_[4083]_  | \new_[4078]_ ;
  assign \new_[4085]_  = \new_[4084]_  | \new_[4073]_ ;
  assign \new_[4089]_  = \new_[2715]_  | \new_[2716]_ ;
  assign \new_[4090]_  = \new_[2717]_  | \new_[4089]_ ;
  assign \new_[4094]_  = \new_[2712]_  | \new_[2713]_ ;
  assign \new_[4095]_  = \new_[2714]_  | \new_[4094]_ ;
  assign \new_[4096]_  = \new_[4095]_  | \new_[4090]_ ;
  assign \new_[4100]_  = \new_[2709]_  | \new_[2710]_ ;
  assign \new_[4101]_  = \new_[2711]_  | \new_[4100]_ ;
  assign \new_[4104]_  = \new_[2707]_  | \new_[2708]_ ;
  assign \new_[4107]_  = \new_[2705]_  | \new_[2706]_ ;
  assign \new_[4108]_  = \new_[4107]_  | \new_[4104]_ ;
  assign \new_[4109]_  = \new_[4108]_  | \new_[4101]_ ;
  assign \new_[4110]_  = \new_[4109]_  | \new_[4096]_ ;
  assign \new_[4111]_  = \new_[4110]_  | \new_[4085]_ ;
  assign \new_[4115]_  = \new_[2702]_  | \new_[2703]_ ;
  assign \new_[4116]_  = \new_[2704]_  | \new_[4115]_ ;
  assign \new_[4120]_  = \new_[2699]_  | \new_[2700]_ ;
  assign \new_[4121]_  = \new_[2701]_  | \new_[4120]_ ;
  assign \new_[4122]_  = \new_[4121]_  | \new_[4116]_ ;
  assign \new_[4126]_  = \new_[2696]_  | \new_[2697]_ ;
  assign \new_[4127]_  = \new_[2698]_  | \new_[4126]_ ;
  assign \new_[4131]_  = \new_[2693]_  | \new_[2694]_ ;
  assign \new_[4132]_  = \new_[2695]_  | \new_[4131]_ ;
  assign \new_[4133]_  = \new_[4132]_  | \new_[4127]_ ;
  assign \new_[4134]_  = \new_[4133]_  | \new_[4122]_ ;
  assign \new_[4138]_  = \new_[2690]_  | \new_[2691]_ ;
  assign \new_[4139]_  = \new_[2692]_  | \new_[4138]_ ;
  assign \new_[4143]_  = \new_[2687]_  | \new_[2688]_ ;
  assign \new_[4144]_  = \new_[2689]_  | \new_[4143]_ ;
  assign \new_[4145]_  = \new_[4144]_  | \new_[4139]_ ;
  assign \new_[4149]_  = \new_[2684]_  | \new_[2685]_ ;
  assign \new_[4150]_  = \new_[2686]_  | \new_[4149]_ ;
  assign \new_[4153]_  = \new_[2682]_  | \new_[2683]_ ;
  assign \new_[4156]_  = \new_[2680]_  | \new_[2681]_ ;
  assign \new_[4157]_  = \new_[4156]_  | \new_[4153]_ ;
  assign \new_[4158]_  = \new_[4157]_  | \new_[4150]_ ;
  assign \new_[4159]_  = \new_[4158]_  | \new_[4145]_ ;
  assign \new_[4160]_  = \new_[4159]_  | \new_[4134]_ ;
  assign \new_[4161]_  = \new_[4160]_  | \new_[4111]_ ;
  assign \new_[4162]_  = \new_[4161]_  | \new_[4062]_ ;
  assign \new_[4166]_  = \new_[2677]_  | \new_[2678]_ ;
  assign \new_[4167]_  = \new_[2679]_  | \new_[4166]_ ;
  assign \new_[4171]_  = \new_[2674]_  | \new_[2675]_ ;
  assign \new_[4172]_  = \new_[2676]_  | \new_[4171]_ ;
  assign \new_[4173]_  = \new_[4172]_  | \new_[4167]_ ;
  assign \new_[4177]_  = \new_[2671]_  | \new_[2672]_ ;
  assign \new_[4178]_  = \new_[2673]_  | \new_[4177]_ ;
  assign \new_[4182]_  = \new_[2668]_  | \new_[2669]_ ;
  assign \new_[4183]_  = \new_[2670]_  | \new_[4182]_ ;
  assign \new_[4184]_  = \new_[4183]_  | \new_[4178]_ ;
  assign \new_[4185]_  = \new_[4184]_  | \new_[4173]_ ;
  assign \new_[4189]_  = \new_[2665]_  | \new_[2666]_ ;
  assign \new_[4190]_  = \new_[2667]_  | \new_[4189]_ ;
  assign \new_[4194]_  = \new_[2662]_  | \new_[2663]_ ;
  assign \new_[4195]_  = \new_[2664]_  | \new_[4194]_ ;
  assign \new_[4196]_  = \new_[4195]_  | \new_[4190]_ ;
  assign \new_[4200]_  = \new_[2659]_  | \new_[2660]_ ;
  assign \new_[4201]_  = \new_[2661]_  | \new_[4200]_ ;
  assign \new_[4205]_  = \new_[2656]_  | \new_[2657]_ ;
  assign \new_[4206]_  = \new_[2658]_  | \new_[4205]_ ;
  assign \new_[4207]_  = \new_[4206]_  | \new_[4201]_ ;
  assign \new_[4208]_  = \new_[4207]_  | \new_[4196]_ ;
  assign \new_[4209]_  = \new_[4208]_  | \new_[4185]_ ;
  assign \new_[4213]_  = \new_[2653]_  | \new_[2654]_ ;
  assign \new_[4214]_  = \new_[2655]_  | \new_[4213]_ ;
  assign \new_[4218]_  = \new_[2650]_  | \new_[2651]_ ;
  assign \new_[4219]_  = \new_[2652]_  | \new_[4218]_ ;
  assign \new_[4220]_  = \new_[4219]_  | \new_[4214]_ ;
  assign \new_[4224]_  = \new_[2647]_  | \new_[2648]_ ;
  assign \new_[4225]_  = \new_[2649]_  | \new_[4224]_ ;
  assign \new_[4229]_  = \new_[2644]_  | \new_[2645]_ ;
  assign \new_[4230]_  = \new_[2646]_  | \new_[4229]_ ;
  assign \new_[4231]_  = \new_[4230]_  | \new_[4225]_ ;
  assign \new_[4232]_  = \new_[4231]_  | \new_[4220]_ ;
  assign \new_[4236]_  = \new_[2641]_  | \new_[2642]_ ;
  assign \new_[4237]_  = \new_[2643]_  | \new_[4236]_ ;
  assign \new_[4241]_  = \new_[2638]_  | \new_[2639]_ ;
  assign \new_[4242]_  = \new_[2640]_  | \new_[4241]_ ;
  assign \new_[4243]_  = \new_[4242]_  | \new_[4237]_ ;
  assign \new_[4247]_  = \new_[2635]_  | \new_[2636]_ ;
  assign \new_[4248]_  = \new_[2637]_  | \new_[4247]_ ;
  assign \new_[4251]_  = \new_[2633]_  | \new_[2634]_ ;
  assign \new_[4254]_  = \new_[2631]_  | \new_[2632]_ ;
  assign \new_[4255]_  = \new_[4254]_  | \new_[4251]_ ;
  assign \new_[4256]_  = \new_[4255]_  | \new_[4248]_ ;
  assign \new_[4257]_  = \new_[4256]_  | \new_[4243]_ ;
  assign \new_[4258]_  = \new_[4257]_  | \new_[4232]_ ;
  assign \new_[4259]_  = \new_[4258]_  | \new_[4209]_ ;
  assign \new_[4263]_  = \new_[2628]_  | \new_[2629]_ ;
  assign \new_[4264]_  = \new_[2630]_  | \new_[4263]_ ;
  assign \new_[4268]_  = \new_[2625]_  | \new_[2626]_ ;
  assign \new_[4269]_  = \new_[2627]_  | \new_[4268]_ ;
  assign \new_[4270]_  = \new_[4269]_  | \new_[4264]_ ;
  assign \new_[4274]_  = \new_[2622]_  | \new_[2623]_ ;
  assign \new_[4275]_  = \new_[2624]_  | \new_[4274]_ ;
  assign \new_[4279]_  = \new_[2619]_  | \new_[2620]_ ;
  assign \new_[4280]_  = \new_[2621]_  | \new_[4279]_ ;
  assign \new_[4281]_  = \new_[4280]_  | \new_[4275]_ ;
  assign \new_[4282]_  = \new_[4281]_  | \new_[4270]_ ;
  assign \new_[4286]_  = \new_[2616]_  | \new_[2617]_ ;
  assign \new_[4287]_  = \new_[2618]_  | \new_[4286]_ ;
  assign \new_[4291]_  = \new_[2613]_  | \new_[2614]_ ;
  assign \new_[4292]_  = \new_[2615]_  | \new_[4291]_ ;
  assign \new_[4293]_  = \new_[4292]_  | \new_[4287]_ ;
  assign \new_[4297]_  = \new_[2610]_  | \new_[2611]_ ;
  assign \new_[4298]_  = \new_[2612]_  | \new_[4297]_ ;
  assign \new_[4301]_  = \new_[2608]_  | \new_[2609]_ ;
  assign \new_[4304]_  = \new_[2606]_  | \new_[2607]_ ;
  assign \new_[4305]_  = \new_[4304]_  | \new_[4301]_ ;
  assign \new_[4306]_  = \new_[4305]_  | \new_[4298]_ ;
  assign \new_[4307]_  = \new_[4306]_  | \new_[4293]_ ;
  assign \new_[4308]_  = \new_[4307]_  | \new_[4282]_ ;
  assign \new_[4312]_  = \new_[2603]_  | \new_[2604]_ ;
  assign \new_[4313]_  = \new_[2605]_  | \new_[4312]_ ;
  assign \new_[4317]_  = \new_[2600]_  | \new_[2601]_ ;
  assign \new_[4318]_  = \new_[2602]_  | \new_[4317]_ ;
  assign \new_[4319]_  = \new_[4318]_  | \new_[4313]_ ;
  assign \new_[4323]_  = \new_[2597]_  | \new_[2598]_ ;
  assign \new_[4324]_  = \new_[2599]_  | \new_[4323]_ ;
  assign \new_[4328]_  = \new_[2594]_  | \new_[2595]_ ;
  assign \new_[4329]_  = \new_[2596]_  | \new_[4328]_ ;
  assign \new_[4330]_  = \new_[4329]_  | \new_[4324]_ ;
  assign \new_[4331]_  = \new_[4330]_  | \new_[4319]_ ;
  assign \new_[4335]_  = \new_[2591]_  | \new_[2592]_ ;
  assign \new_[4336]_  = \new_[2593]_  | \new_[4335]_ ;
  assign \new_[4340]_  = \new_[2588]_  | \new_[2589]_ ;
  assign \new_[4341]_  = \new_[2590]_  | \new_[4340]_ ;
  assign \new_[4342]_  = \new_[4341]_  | \new_[4336]_ ;
  assign \new_[4346]_  = \new_[2585]_  | \new_[2586]_ ;
  assign \new_[4347]_  = \new_[2587]_  | \new_[4346]_ ;
  assign \new_[4350]_  = \new_[2583]_  | \new_[2584]_ ;
  assign \new_[4353]_  = \new_[2581]_  | \new_[2582]_ ;
  assign \new_[4354]_  = \new_[4353]_  | \new_[4350]_ ;
  assign \new_[4355]_  = \new_[4354]_  | \new_[4347]_ ;
  assign \new_[4356]_  = \new_[4355]_  | \new_[4342]_ ;
  assign \new_[4357]_  = \new_[4356]_  | \new_[4331]_ ;
  assign \new_[4358]_  = \new_[4357]_  | \new_[4308]_ ;
  assign \new_[4359]_  = \new_[4358]_  | \new_[4259]_ ;
  assign \new_[4360]_  = \new_[4359]_  | \new_[4162]_ ;
  assign \new_[4364]_  = \new_[2578]_  | \new_[2579]_ ;
  assign \new_[4365]_  = \new_[2580]_  | \new_[4364]_ ;
  assign \new_[4369]_  = \new_[2575]_  | \new_[2576]_ ;
  assign \new_[4370]_  = \new_[2577]_  | \new_[4369]_ ;
  assign \new_[4371]_  = \new_[4370]_  | \new_[4365]_ ;
  assign \new_[4375]_  = \new_[2572]_  | \new_[2573]_ ;
  assign \new_[4376]_  = \new_[2574]_  | \new_[4375]_ ;
  assign \new_[4380]_  = \new_[2569]_  | \new_[2570]_ ;
  assign \new_[4381]_  = \new_[2571]_  | \new_[4380]_ ;
  assign \new_[4382]_  = \new_[4381]_  | \new_[4376]_ ;
  assign \new_[4383]_  = \new_[4382]_  | \new_[4371]_ ;
  assign \new_[4387]_  = \new_[2566]_  | \new_[2567]_ ;
  assign \new_[4388]_  = \new_[2568]_  | \new_[4387]_ ;
  assign \new_[4392]_  = \new_[2563]_  | \new_[2564]_ ;
  assign \new_[4393]_  = \new_[2565]_  | \new_[4392]_ ;
  assign \new_[4394]_  = \new_[4393]_  | \new_[4388]_ ;
  assign \new_[4398]_  = \new_[2560]_  | \new_[2561]_ ;
  assign \new_[4399]_  = \new_[2562]_  | \new_[4398]_ ;
  assign \new_[4403]_  = \new_[2557]_  | \new_[2558]_ ;
  assign \new_[4404]_  = \new_[2559]_  | \new_[4403]_ ;
  assign \new_[4405]_  = \new_[4404]_  | \new_[4399]_ ;
  assign \new_[4406]_  = \new_[4405]_  | \new_[4394]_ ;
  assign \new_[4407]_  = \new_[4406]_  | \new_[4383]_ ;
  assign \new_[4411]_  = \new_[2554]_  | \new_[2555]_ ;
  assign \new_[4412]_  = \new_[2556]_  | \new_[4411]_ ;
  assign \new_[4416]_  = \new_[2551]_  | \new_[2552]_ ;
  assign \new_[4417]_  = \new_[2553]_  | \new_[4416]_ ;
  assign \new_[4418]_  = \new_[4417]_  | \new_[4412]_ ;
  assign \new_[4422]_  = \new_[2548]_  | \new_[2549]_ ;
  assign \new_[4423]_  = \new_[2550]_  | \new_[4422]_ ;
  assign \new_[4427]_  = \new_[2545]_  | \new_[2546]_ ;
  assign \new_[4428]_  = \new_[2547]_  | \new_[4427]_ ;
  assign \new_[4429]_  = \new_[4428]_  | \new_[4423]_ ;
  assign \new_[4430]_  = \new_[4429]_  | \new_[4418]_ ;
  assign \new_[4434]_  = \new_[2542]_  | \new_[2543]_ ;
  assign \new_[4435]_  = \new_[2544]_  | \new_[4434]_ ;
  assign \new_[4439]_  = \new_[2539]_  | \new_[2540]_ ;
  assign \new_[4440]_  = \new_[2541]_  | \new_[4439]_ ;
  assign \new_[4441]_  = \new_[4440]_  | \new_[4435]_ ;
  assign \new_[4445]_  = \new_[2536]_  | \new_[2537]_ ;
  assign \new_[4446]_  = \new_[2538]_  | \new_[4445]_ ;
  assign \new_[4449]_  = \new_[2534]_  | \new_[2535]_ ;
  assign \new_[4452]_  = \new_[2532]_  | \new_[2533]_ ;
  assign \new_[4453]_  = \new_[4452]_  | \new_[4449]_ ;
  assign \new_[4454]_  = \new_[4453]_  | \new_[4446]_ ;
  assign \new_[4455]_  = \new_[4454]_  | \new_[4441]_ ;
  assign \new_[4456]_  = \new_[4455]_  | \new_[4430]_ ;
  assign \new_[4457]_  = \new_[4456]_  | \new_[4407]_ ;
  assign \new_[4461]_  = \new_[2529]_  | \new_[2530]_ ;
  assign \new_[4462]_  = \new_[2531]_  | \new_[4461]_ ;
  assign \new_[4466]_  = \new_[2526]_  | \new_[2527]_ ;
  assign \new_[4467]_  = \new_[2528]_  | \new_[4466]_ ;
  assign \new_[4468]_  = \new_[4467]_  | \new_[4462]_ ;
  assign \new_[4472]_  = \new_[2523]_  | \new_[2524]_ ;
  assign \new_[4473]_  = \new_[2525]_  | \new_[4472]_ ;
  assign \new_[4477]_  = \new_[2520]_  | \new_[2521]_ ;
  assign \new_[4478]_  = \new_[2522]_  | \new_[4477]_ ;
  assign \new_[4479]_  = \new_[4478]_  | \new_[4473]_ ;
  assign \new_[4480]_  = \new_[4479]_  | \new_[4468]_ ;
  assign \new_[4484]_  = \new_[2517]_  | \new_[2518]_ ;
  assign \new_[4485]_  = \new_[2519]_  | \new_[4484]_ ;
  assign \new_[4489]_  = \new_[2514]_  | \new_[2515]_ ;
  assign \new_[4490]_  = \new_[2516]_  | \new_[4489]_ ;
  assign \new_[4491]_  = \new_[4490]_  | \new_[4485]_ ;
  assign \new_[4495]_  = \new_[2511]_  | \new_[2512]_ ;
  assign \new_[4496]_  = \new_[2513]_  | \new_[4495]_ ;
  assign \new_[4499]_  = \new_[2509]_  | \new_[2510]_ ;
  assign \new_[4502]_  = \new_[2507]_  | \new_[2508]_ ;
  assign \new_[4503]_  = \new_[4502]_  | \new_[4499]_ ;
  assign \new_[4504]_  = \new_[4503]_  | \new_[4496]_ ;
  assign \new_[4505]_  = \new_[4504]_  | \new_[4491]_ ;
  assign \new_[4506]_  = \new_[4505]_  | \new_[4480]_ ;
  assign \new_[4510]_  = \new_[2504]_  | \new_[2505]_ ;
  assign \new_[4511]_  = \new_[2506]_  | \new_[4510]_ ;
  assign \new_[4515]_  = \new_[2501]_  | \new_[2502]_ ;
  assign \new_[4516]_  = \new_[2503]_  | \new_[4515]_ ;
  assign \new_[4517]_  = \new_[4516]_  | \new_[4511]_ ;
  assign \new_[4521]_  = \new_[2498]_  | \new_[2499]_ ;
  assign \new_[4522]_  = \new_[2500]_  | \new_[4521]_ ;
  assign \new_[4526]_  = \new_[2495]_  | \new_[2496]_ ;
  assign \new_[4527]_  = \new_[2497]_  | \new_[4526]_ ;
  assign \new_[4528]_  = \new_[4527]_  | \new_[4522]_ ;
  assign \new_[4529]_  = \new_[4528]_  | \new_[4517]_ ;
  assign \new_[4533]_  = \new_[2492]_  | \new_[2493]_ ;
  assign \new_[4534]_  = \new_[2494]_  | \new_[4533]_ ;
  assign \new_[4538]_  = \new_[2489]_  | \new_[2490]_ ;
  assign \new_[4539]_  = \new_[2491]_  | \new_[4538]_ ;
  assign \new_[4540]_  = \new_[4539]_  | \new_[4534]_ ;
  assign \new_[4544]_  = \new_[2486]_  | \new_[2487]_ ;
  assign \new_[4545]_  = \new_[2488]_  | \new_[4544]_ ;
  assign \new_[4548]_  = \new_[2484]_  | \new_[2485]_ ;
  assign \new_[4551]_  = \new_[2482]_  | \new_[2483]_ ;
  assign \new_[4552]_  = \new_[4551]_  | \new_[4548]_ ;
  assign \new_[4553]_  = \new_[4552]_  | \new_[4545]_ ;
  assign \new_[4554]_  = \new_[4553]_  | \new_[4540]_ ;
  assign \new_[4555]_  = \new_[4554]_  | \new_[4529]_ ;
  assign \new_[4556]_  = \new_[4555]_  | \new_[4506]_ ;
  assign \new_[4557]_  = \new_[4556]_  | \new_[4457]_ ;
  assign \new_[4561]_  = \new_[2479]_  | \new_[2480]_ ;
  assign \new_[4562]_  = \new_[2481]_  | \new_[4561]_ ;
  assign \new_[4566]_  = \new_[2476]_  | \new_[2477]_ ;
  assign \new_[4567]_  = \new_[2478]_  | \new_[4566]_ ;
  assign \new_[4568]_  = \new_[4567]_  | \new_[4562]_ ;
  assign \new_[4572]_  = \new_[2473]_  | \new_[2474]_ ;
  assign \new_[4573]_  = \new_[2475]_  | \new_[4572]_ ;
  assign \new_[4577]_  = \new_[2470]_  | \new_[2471]_ ;
  assign \new_[4578]_  = \new_[2472]_  | \new_[4577]_ ;
  assign \new_[4579]_  = \new_[4578]_  | \new_[4573]_ ;
  assign \new_[4580]_  = \new_[4579]_  | \new_[4568]_ ;
  assign \new_[4584]_  = \new_[2467]_  | \new_[2468]_ ;
  assign \new_[4585]_  = \new_[2469]_  | \new_[4584]_ ;
  assign \new_[4589]_  = \new_[2464]_  | \new_[2465]_ ;
  assign \new_[4590]_  = \new_[2466]_  | \new_[4589]_ ;
  assign \new_[4591]_  = \new_[4590]_  | \new_[4585]_ ;
  assign \new_[4595]_  = \new_[2461]_  | \new_[2462]_ ;
  assign \new_[4596]_  = \new_[2463]_  | \new_[4595]_ ;
  assign \new_[4599]_  = \new_[2459]_  | \new_[2460]_ ;
  assign \new_[4602]_  = \new_[2457]_  | \new_[2458]_ ;
  assign \new_[4603]_  = \new_[4602]_  | \new_[4599]_ ;
  assign \new_[4604]_  = \new_[4603]_  | \new_[4596]_ ;
  assign \new_[4605]_  = \new_[4604]_  | \new_[4591]_ ;
  assign \new_[4606]_  = \new_[4605]_  | \new_[4580]_ ;
  assign \new_[4610]_  = \new_[2454]_  | \new_[2455]_ ;
  assign \new_[4611]_  = \new_[2456]_  | \new_[4610]_ ;
  assign \new_[4615]_  = \new_[2451]_  | \new_[2452]_ ;
  assign \new_[4616]_  = \new_[2453]_  | \new_[4615]_ ;
  assign \new_[4617]_  = \new_[4616]_  | \new_[4611]_ ;
  assign \new_[4621]_  = \new_[2448]_  | \new_[2449]_ ;
  assign \new_[4622]_  = \new_[2450]_  | \new_[4621]_ ;
  assign \new_[4626]_  = \new_[2445]_  | \new_[2446]_ ;
  assign \new_[4627]_  = \new_[2447]_  | \new_[4626]_ ;
  assign \new_[4628]_  = \new_[4627]_  | \new_[4622]_ ;
  assign \new_[4629]_  = \new_[4628]_  | \new_[4617]_ ;
  assign \new_[4633]_  = \new_[2442]_  | \new_[2443]_ ;
  assign \new_[4634]_  = \new_[2444]_  | \new_[4633]_ ;
  assign \new_[4638]_  = \new_[2439]_  | \new_[2440]_ ;
  assign \new_[4639]_  = \new_[2441]_  | \new_[4638]_ ;
  assign \new_[4640]_  = \new_[4639]_  | \new_[4634]_ ;
  assign \new_[4644]_  = \new_[2436]_  | \new_[2437]_ ;
  assign \new_[4645]_  = \new_[2438]_  | \new_[4644]_ ;
  assign \new_[4648]_  = \new_[2434]_  | \new_[2435]_ ;
  assign \new_[4651]_  = \new_[2432]_  | \new_[2433]_ ;
  assign \new_[4652]_  = \new_[4651]_  | \new_[4648]_ ;
  assign \new_[4653]_  = \new_[4652]_  | \new_[4645]_ ;
  assign \new_[4654]_  = \new_[4653]_  | \new_[4640]_ ;
  assign \new_[4655]_  = \new_[4654]_  | \new_[4629]_ ;
  assign \new_[4656]_  = \new_[4655]_  | \new_[4606]_ ;
  assign \new_[4660]_  = \new_[2429]_  | \new_[2430]_ ;
  assign \new_[4661]_  = \new_[2431]_  | \new_[4660]_ ;
  assign \new_[4665]_  = \new_[2426]_  | \new_[2427]_ ;
  assign \new_[4666]_  = \new_[2428]_  | \new_[4665]_ ;
  assign \new_[4667]_  = \new_[4666]_  | \new_[4661]_ ;
  assign \new_[4671]_  = \new_[2423]_  | \new_[2424]_ ;
  assign \new_[4672]_  = \new_[2425]_  | \new_[4671]_ ;
  assign \new_[4676]_  = \new_[2420]_  | \new_[2421]_ ;
  assign \new_[4677]_  = \new_[2422]_  | \new_[4676]_ ;
  assign \new_[4678]_  = \new_[4677]_  | \new_[4672]_ ;
  assign \new_[4679]_  = \new_[4678]_  | \new_[4667]_ ;
  assign \new_[4683]_  = \new_[2417]_  | \new_[2418]_ ;
  assign \new_[4684]_  = \new_[2419]_  | \new_[4683]_ ;
  assign \new_[4688]_  = \new_[2414]_  | \new_[2415]_ ;
  assign \new_[4689]_  = \new_[2416]_  | \new_[4688]_ ;
  assign \new_[4690]_  = \new_[4689]_  | \new_[4684]_ ;
  assign \new_[4694]_  = \new_[2411]_  | \new_[2412]_ ;
  assign \new_[4695]_  = \new_[2413]_  | \new_[4694]_ ;
  assign \new_[4698]_  = \new_[2409]_  | \new_[2410]_ ;
  assign \new_[4701]_  = \new_[2407]_  | \new_[2408]_ ;
  assign \new_[4702]_  = \new_[4701]_  | \new_[4698]_ ;
  assign \new_[4703]_  = \new_[4702]_  | \new_[4695]_ ;
  assign \new_[4704]_  = \new_[4703]_  | \new_[4690]_ ;
  assign \new_[4705]_  = \new_[4704]_  | \new_[4679]_ ;
  assign \new_[4709]_  = \new_[2404]_  | \new_[2405]_ ;
  assign \new_[4710]_  = \new_[2406]_  | \new_[4709]_ ;
  assign \new_[4714]_  = \new_[2401]_  | \new_[2402]_ ;
  assign \new_[4715]_  = \new_[2403]_  | \new_[4714]_ ;
  assign \new_[4716]_  = \new_[4715]_  | \new_[4710]_ ;
  assign \new_[4720]_  = \new_[2398]_  | \new_[2399]_ ;
  assign \new_[4721]_  = \new_[2400]_  | \new_[4720]_ ;
  assign \new_[4725]_  = \new_[2395]_  | \new_[2396]_ ;
  assign \new_[4726]_  = \new_[2397]_  | \new_[4725]_ ;
  assign \new_[4727]_  = \new_[4726]_  | \new_[4721]_ ;
  assign \new_[4728]_  = \new_[4727]_  | \new_[4716]_ ;
  assign \new_[4732]_  = \new_[2392]_  | \new_[2393]_ ;
  assign \new_[4733]_  = \new_[2394]_  | \new_[4732]_ ;
  assign \new_[4737]_  = \new_[2389]_  | \new_[2390]_ ;
  assign \new_[4738]_  = \new_[2391]_  | \new_[4737]_ ;
  assign \new_[4739]_  = \new_[4738]_  | \new_[4733]_ ;
  assign \new_[4743]_  = \new_[2386]_  | \new_[2387]_ ;
  assign \new_[4744]_  = \new_[2388]_  | \new_[4743]_ ;
  assign \new_[4747]_  = \new_[2384]_  | \new_[2385]_ ;
  assign \new_[4750]_  = \new_[2382]_  | \new_[2383]_ ;
  assign \new_[4751]_  = \new_[4750]_  | \new_[4747]_ ;
  assign \new_[4752]_  = \new_[4751]_  | \new_[4744]_ ;
  assign \new_[4753]_  = \new_[4752]_  | \new_[4739]_ ;
  assign \new_[4754]_  = \new_[4753]_  | \new_[4728]_ ;
  assign \new_[4755]_  = \new_[4754]_  | \new_[4705]_ ;
  assign \new_[4756]_  = \new_[4755]_  | \new_[4656]_ ;
  assign \new_[4757]_  = \new_[4756]_  | \new_[4557]_ ;
  assign \new_[4758]_  = \new_[4757]_  | \new_[4360]_ ;
  assign \new_[4759]_  = \new_[4758]_  | \new_[3965]_ ;
  assign \new_[4763]_  = \new_[2379]_  | \new_[2380]_ ;
  assign \new_[4764]_  = \new_[2381]_  | \new_[4763]_ ;
  assign \new_[4768]_  = \new_[2376]_  | \new_[2377]_ ;
  assign \new_[4769]_  = \new_[2378]_  | \new_[4768]_ ;
  assign \new_[4770]_  = \new_[4769]_  | \new_[4764]_ ;
  assign \new_[4774]_  = \new_[2373]_  | \new_[2374]_ ;
  assign \new_[4775]_  = \new_[2375]_  | \new_[4774]_ ;
  assign \new_[4779]_  = \new_[2370]_  | \new_[2371]_ ;
  assign \new_[4780]_  = \new_[2372]_  | \new_[4779]_ ;
  assign \new_[4781]_  = \new_[4780]_  | \new_[4775]_ ;
  assign \new_[4782]_  = \new_[4781]_  | \new_[4770]_ ;
  assign \new_[4786]_  = \new_[2367]_  | \new_[2368]_ ;
  assign \new_[4787]_  = \new_[2369]_  | \new_[4786]_ ;
  assign \new_[4791]_  = \new_[2364]_  | \new_[2365]_ ;
  assign \new_[4792]_  = \new_[2366]_  | \new_[4791]_ ;
  assign \new_[4793]_  = \new_[4792]_  | \new_[4787]_ ;
  assign \new_[4797]_  = \new_[2361]_  | \new_[2362]_ ;
  assign \new_[4798]_  = \new_[2363]_  | \new_[4797]_ ;
  assign \new_[4802]_  = \new_[2358]_  | \new_[2359]_ ;
  assign \new_[4803]_  = \new_[2360]_  | \new_[4802]_ ;
  assign \new_[4804]_  = \new_[4803]_  | \new_[4798]_ ;
  assign \new_[4805]_  = \new_[4804]_  | \new_[4793]_ ;
  assign \new_[4806]_  = \new_[4805]_  | \new_[4782]_ ;
  assign \new_[4810]_  = \new_[2355]_  | \new_[2356]_ ;
  assign \new_[4811]_  = \new_[2357]_  | \new_[4810]_ ;
  assign \new_[4815]_  = \new_[2352]_  | \new_[2353]_ ;
  assign \new_[4816]_  = \new_[2354]_  | \new_[4815]_ ;
  assign \new_[4817]_  = \new_[4816]_  | \new_[4811]_ ;
  assign \new_[4821]_  = \new_[2349]_  | \new_[2350]_ ;
  assign \new_[4822]_  = \new_[2351]_  | \new_[4821]_ ;
  assign \new_[4826]_  = \new_[2346]_  | \new_[2347]_ ;
  assign \new_[4827]_  = \new_[2348]_  | \new_[4826]_ ;
  assign \new_[4828]_  = \new_[4827]_  | \new_[4822]_ ;
  assign \new_[4829]_  = \new_[4828]_  | \new_[4817]_ ;
  assign \new_[4833]_  = \new_[2343]_  | \new_[2344]_ ;
  assign \new_[4834]_  = \new_[2345]_  | \new_[4833]_ ;
  assign \new_[4838]_  = \new_[2340]_  | \new_[2341]_ ;
  assign \new_[4839]_  = \new_[2342]_  | \new_[4838]_ ;
  assign \new_[4840]_  = \new_[4839]_  | \new_[4834]_ ;
  assign \new_[4844]_  = \new_[2337]_  | \new_[2338]_ ;
  assign \new_[4845]_  = \new_[2339]_  | \new_[4844]_ ;
  assign \new_[4848]_  = \new_[2335]_  | \new_[2336]_ ;
  assign \new_[4851]_  = \new_[2333]_  | \new_[2334]_ ;
  assign \new_[4852]_  = \new_[4851]_  | \new_[4848]_ ;
  assign \new_[4853]_  = \new_[4852]_  | \new_[4845]_ ;
  assign \new_[4854]_  = \new_[4853]_  | \new_[4840]_ ;
  assign \new_[4855]_  = \new_[4854]_  | \new_[4829]_ ;
  assign \new_[4856]_  = \new_[4855]_  | \new_[4806]_ ;
  assign \new_[4860]_  = \new_[2330]_  | \new_[2331]_ ;
  assign \new_[4861]_  = \new_[2332]_  | \new_[4860]_ ;
  assign \new_[4865]_  = \new_[2327]_  | \new_[2328]_ ;
  assign \new_[4866]_  = \new_[2329]_  | \new_[4865]_ ;
  assign \new_[4867]_  = \new_[4866]_  | \new_[4861]_ ;
  assign \new_[4871]_  = \new_[2324]_  | \new_[2325]_ ;
  assign \new_[4872]_  = \new_[2326]_  | \new_[4871]_ ;
  assign \new_[4876]_  = \new_[2321]_  | \new_[2322]_ ;
  assign \new_[4877]_  = \new_[2323]_  | \new_[4876]_ ;
  assign \new_[4878]_  = \new_[4877]_  | \new_[4872]_ ;
  assign \new_[4879]_  = \new_[4878]_  | \new_[4867]_ ;
  assign \new_[4883]_  = \new_[2318]_  | \new_[2319]_ ;
  assign \new_[4884]_  = \new_[2320]_  | \new_[4883]_ ;
  assign \new_[4888]_  = \new_[2315]_  | \new_[2316]_ ;
  assign \new_[4889]_  = \new_[2317]_  | \new_[4888]_ ;
  assign \new_[4890]_  = \new_[4889]_  | \new_[4884]_ ;
  assign \new_[4894]_  = \new_[2312]_  | \new_[2313]_ ;
  assign \new_[4895]_  = \new_[2314]_  | \new_[4894]_ ;
  assign \new_[4898]_  = \new_[2310]_  | \new_[2311]_ ;
  assign \new_[4901]_  = \new_[2308]_  | \new_[2309]_ ;
  assign \new_[4902]_  = \new_[4901]_  | \new_[4898]_ ;
  assign \new_[4903]_  = \new_[4902]_  | \new_[4895]_ ;
  assign \new_[4904]_  = \new_[4903]_  | \new_[4890]_ ;
  assign \new_[4905]_  = \new_[4904]_  | \new_[4879]_ ;
  assign \new_[4909]_  = \new_[2305]_  | \new_[2306]_ ;
  assign \new_[4910]_  = \new_[2307]_  | \new_[4909]_ ;
  assign \new_[4914]_  = \new_[2302]_  | \new_[2303]_ ;
  assign \new_[4915]_  = \new_[2304]_  | \new_[4914]_ ;
  assign \new_[4916]_  = \new_[4915]_  | \new_[4910]_ ;
  assign \new_[4920]_  = \new_[2299]_  | \new_[2300]_ ;
  assign \new_[4921]_  = \new_[2301]_  | \new_[4920]_ ;
  assign \new_[4925]_  = \new_[2296]_  | \new_[2297]_ ;
  assign \new_[4926]_  = \new_[2298]_  | \new_[4925]_ ;
  assign \new_[4927]_  = \new_[4926]_  | \new_[4921]_ ;
  assign \new_[4928]_  = \new_[4927]_  | \new_[4916]_ ;
  assign \new_[4932]_  = \new_[2293]_  | \new_[2294]_ ;
  assign \new_[4933]_  = \new_[2295]_  | \new_[4932]_ ;
  assign \new_[4937]_  = \new_[2290]_  | \new_[2291]_ ;
  assign \new_[4938]_  = \new_[2292]_  | \new_[4937]_ ;
  assign \new_[4939]_  = \new_[4938]_  | \new_[4933]_ ;
  assign \new_[4943]_  = \new_[2287]_  | \new_[2288]_ ;
  assign \new_[4944]_  = \new_[2289]_  | \new_[4943]_ ;
  assign \new_[4947]_  = \new_[2285]_  | \new_[2286]_ ;
  assign \new_[4950]_  = \new_[2283]_  | \new_[2284]_ ;
  assign \new_[4951]_  = \new_[4950]_  | \new_[4947]_ ;
  assign \new_[4952]_  = \new_[4951]_  | \new_[4944]_ ;
  assign \new_[4953]_  = \new_[4952]_  | \new_[4939]_ ;
  assign \new_[4954]_  = \new_[4953]_  | \new_[4928]_ ;
  assign \new_[4955]_  = \new_[4954]_  | \new_[4905]_ ;
  assign \new_[4956]_  = \new_[4955]_  | \new_[4856]_ ;
  assign \new_[4960]_  = \new_[2280]_  | \new_[2281]_ ;
  assign \new_[4961]_  = \new_[2282]_  | \new_[4960]_ ;
  assign \new_[4965]_  = \new_[2277]_  | \new_[2278]_ ;
  assign \new_[4966]_  = \new_[2279]_  | \new_[4965]_ ;
  assign \new_[4967]_  = \new_[4966]_  | \new_[4961]_ ;
  assign \new_[4971]_  = \new_[2274]_  | \new_[2275]_ ;
  assign \new_[4972]_  = \new_[2276]_  | \new_[4971]_ ;
  assign \new_[4976]_  = \new_[2271]_  | \new_[2272]_ ;
  assign \new_[4977]_  = \new_[2273]_  | \new_[4976]_ ;
  assign \new_[4978]_  = \new_[4977]_  | \new_[4972]_ ;
  assign \new_[4979]_  = \new_[4978]_  | \new_[4967]_ ;
  assign \new_[4983]_  = \new_[2268]_  | \new_[2269]_ ;
  assign \new_[4984]_  = \new_[2270]_  | \new_[4983]_ ;
  assign \new_[4988]_  = \new_[2265]_  | \new_[2266]_ ;
  assign \new_[4989]_  = \new_[2267]_  | \new_[4988]_ ;
  assign \new_[4990]_  = \new_[4989]_  | \new_[4984]_ ;
  assign \new_[4994]_  = \new_[2262]_  | \new_[2263]_ ;
  assign \new_[4995]_  = \new_[2264]_  | \new_[4994]_ ;
  assign \new_[4999]_  = \new_[2259]_  | \new_[2260]_ ;
  assign \new_[5000]_  = \new_[2261]_  | \new_[4999]_ ;
  assign \new_[5001]_  = \new_[5000]_  | \new_[4995]_ ;
  assign \new_[5002]_  = \new_[5001]_  | \new_[4990]_ ;
  assign \new_[5003]_  = \new_[5002]_  | \new_[4979]_ ;
  assign \new_[5007]_  = \new_[2256]_  | \new_[2257]_ ;
  assign \new_[5008]_  = \new_[2258]_  | \new_[5007]_ ;
  assign \new_[5012]_  = \new_[2253]_  | \new_[2254]_ ;
  assign \new_[5013]_  = \new_[2255]_  | \new_[5012]_ ;
  assign \new_[5014]_  = \new_[5013]_  | \new_[5008]_ ;
  assign \new_[5018]_  = \new_[2250]_  | \new_[2251]_ ;
  assign \new_[5019]_  = \new_[2252]_  | \new_[5018]_ ;
  assign \new_[5023]_  = \new_[2247]_  | \new_[2248]_ ;
  assign \new_[5024]_  = \new_[2249]_  | \new_[5023]_ ;
  assign \new_[5025]_  = \new_[5024]_  | \new_[5019]_ ;
  assign \new_[5026]_  = \new_[5025]_  | \new_[5014]_ ;
  assign \new_[5030]_  = \new_[2244]_  | \new_[2245]_ ;
  assign \new_[5031]_  = \new_[2246]_  | \new_[5030]_ ;
  assign \new_[5035]_  = \new_[2241]_  | \new_[2242]_ ;
  assign \new_[5036]_  = \new_[2243]_  | \new_[5035]_ ;
  assign \new_[5037]_  = \new_[5036]_  | \new_[5031]_ ;
  assign \new_[5041]_  = \new_[2238]_  | \new_[2239]_ ;
  assign \new_[5042]_  = \new_[2240]_  | \new_[5041]_ ;
  assign \new_[5045]_  = \new_[2236]_  | \new_[2237]_ ;
  assign \new_[5048]_  = \new_[2234]_  | \new_[2235]_ ;
  assign \new_[5049]_  = \new_[5048]_  | \new_[5045]_ ;
  assign \new_[5050]_  = \new_[5049]_  | \new_[5042]_ ;
  assign \new_[5051]_  = \new_[5050]_  | \new_[5037]_ ;
  assign \new_[5052]_  = \new_[5051]_  | \new_[5026]_ ;
  assign \new_[5053]_  = \new_[5052]_  | \new_[5003]_ ;
  assign \new_[5057]_  = \new_[2231]_  | \new_[2232]_ ;
  assign \new_[5058]_  = \new_[2233]_  | \new_[5057]_ ;
  assign \new_[5062]_  = \new_[2228]_  | \new_[2229]_ ;
  assign \new_[5063]_  = \new_[2230]_  | \new_[5062]_ ;
  assign \new_[5064]_  = \new_[5063]_  | \new_[5058]_ ;
  assign \new_[5068]_  = \new_[2225]_  | \new_[2226]_ ;
  assign \new_[5069]_  = \new_[2227]_  | \new_[5068]_ ;
  assign \new_[5073]_  = \new_[2222]_  | \new_[2223]_ ;
  assign \new_[5074]_  = \new_[2224]_  | \new_[5073]_ ;
  assign \new_[5075]_  = \new_[5074]_  | \new_[5069]_ ;
  assign \new_[5076]_  = \new_[5075]_  | \new_[5064]_ ;
  assign \new_[5080]_  = \new_[2219]_  | \new_[2220]_ ;
  assign \new_[5081]_  = \new_[2221]_  | \new_[5080]_ ;
  assign \new_[5085]_  = \new_[2216]_  | \new_[2217]_ ;
  assign \new_[5086]_  = \new_[2218]_  | \new_[5085]_ ;
  assign \new_[5087]_  = \new_[5086]_  | \new_[5081]_ ;
  assign \new_[5091]_  = \new_[2213]_  | \new_[2214]_ ;
  assign \new_[5092]_  = \new_[2215]_  | \new_[5091]_ ;
  assign \new_[5095]_  = \new_[2211]_  | \new_[2212]_ ;
  assign \new_[5098]_  = \new_[2209]_  | \new_[2210]_ ;
  assign \new_[5099]_  = \new_[5098]_  | \new_[5095]_ ;
  assign \new_[5100]_  = \new_[5099]_  | \new_[5092]_ ;
  assign \new_[5101]_  = \new_[5100]_  | \new_[5087]_ ;
  assign \new_[5102]_  = \new_[5101]_  | \new_[5076]_ ;
  assign \new_[5106]_  = \new_[2206]_  | \new_[2207]_ ;
  assign \new_[5107]_  = \new_[2208]_  | \new_[5106]_ ;
  assign \new_[5111]_  = \new_[2203]_  | \new_[2204]_ ;
  assign \new_[5112]_  = \new_[2205]_  | \new_[5111]_ ;
  assign \new_[5113]_  = \new_[5112]_  | \new_[5107]_ ;
  assign \new_[5117]_  = \new_[2200]_  | \new_[2201]_ ;
  assign \new_[5118]_  = \new_[2202]_  | \new_[5117]_ ;
  assign \new_[5122]_  = \new_[2197]_  | \new_[2198]_ ;
  assign \new_[5123]_  = \new_[2199]_  | \new_[5122]_ ;
  assign \new_[5124]_  = \new_[5123]_  | \new_[5118]_ ;
  assign \new_[5125]_  = \new_[5124]_  | \new_[5113]_ ;
  assign \new_[5129]_  = \new_[2194]_  | \new_[2195]_ ;
  assign \new_[5130]_  = \new_[2196]_  | \new_[5129]_ ;
  assign \new_[5134]_  = \new_[2191]_  | \new_[2192]_ ;
  assign \new_[5135]_  = \new_[2193]_  | \new_[5134]_ ;
  assign \new_[5136]_  = \new_[5135]_  | \new_[5130]_ ;
  assign \new_[5140]_  = \new_[2188]_  | \new_[2189]_ ;
  assign \new_[5141]_  = \new_[2190]_  | \new_[5140]_ ;
  assign \new_[5144]_  = \new_[2186]_  | \new_[2187]_ ;
  assign \new_[5147]_  = \new_[2184]_  | \new_[2185]_ ;
  assign \new_[5148]_  = \new_[5147]_  | \new_[5144]_ ;
  assign \new_[5149]_  = \new_[5148]_  | \new_[5141]_ ;
  assign \new_[5150]_  = \new_[5149]_  | \new_[5136]_ ;
  assign \new_[5151]_  = \new_[5150]_  | \new_[5125]_ ;
  assign \new_[5152]_  = \new_[5151]_  | \new_[5102]_ ;
  assign \new_[5153]_  = \new_[5152]_  | \new_[5053]_ ;
  assign \new_[5154]_  = \new_[5153]_  | \new_[4956]_ ;
  assign \new_[5158]_  = \new_[2181]_  | \new_[2182]_ ;
  assign \new_[5159]_  = \new_[2183]_  | \new_[5158]_ ;
  assign \new_[5163]_  = \new_[2178]_  | \new_[2179]_ ;
  assign \new_[5164]_  = \new_[2180]_  | \new_[5163]_ ;
  assign \new_[5165]_  = \new_[5164]_  | \new_[5159]_ ;
  assign \new_[5169]_  = \new_[2175]_  | \new_[2176]_ ;
  assign \new_[5170]_  = \new_[2177]_  | \new_[5169]_ ;
  assign \new_[5174]_  = \new_[2172]_  | \new_[2173]_ ;
  assign \new_[5175]_  = \new_[2174]_  | \new_[5174]_ ;
  assign \new_[5176]_  = \new_[5175]_  | \new_[5170]_ ;
  assign \new_[5177]_  = \new_[5176]_  | \new_[5165]_ ;
  assign \new_[5181]_  = \new_[2169]_  | \new_[2170]_ ;
  assign \new_[5182]_  = \new_[2171]_  | \new_[5181]_ ;
  assign \new_[5186]_  = \new_[2166]_  | \new_[2167]_ ;
  assign \new_[5187]_  = \new_[2168]_  | \new_[5186]_ ;
  assign \new_[5188]_  = \new_[5187]_  | \new_[5182]_ ;
  assign \new_[5192]_  = \new_[2163]_  | \new_[2164]_ ;
  assign \new_[5193]_  = \new_[2165]_  | \new_[5192]_ ;
  assign \new_[5197]_  = \new_[2160]_  | \new_[2161]_ ;
  assign \new_[5198]_  = \new_[2162]_  | \new_[5197]_ ;
  assign \new_[5199]_  = \new_[5198]_  | \new_[5193]_ ;
  assign \new_[5200]_  = \new_[5199]_  | \new_[5188]_ ;
  assign \new_[5201]_  = \new_[5200]_  | \new_[5177]_ ;
  assign \new_[5205]_  = \new_[2157]_  | \new_[2158]_ ;
  assign \new_[5206]_  = \new_[2159]_  | \new_[5205]_ ;
  assign \new_[5210]_  = \new_[2154]_  | \new_[2155]_ ;
  assign \new_[5211]_  = \new_[2156]_  | \new_[5210]_ ;
  assign \new_[5212]_  = \new_[5211]_  | \new_[5206]_ ;
  assign \new_[5216]_  = \new_[2151]_  | \new_[2152]_ ;
  assign \new_[5217]_  = \new_[2153]_  | \new_[5216]_ ;
  assign \new_[5221]_  = \new_[2148]_  | \new_[2149]_ ;
  assign \new_[5222]_  = \new_[2150]_  | \new_[5221]_ ;
  assign \new_[5223]_  = \new_[5222]_  | \new_[5217]_ ;
  assign \new_[5224]_  = \new_[5223]_  | \new_[5212]_ ;
  assign \new_[5228]_  = \new_[2145]_  | \new_[2146]_ ;
  assign \new_[5229]_  = \new_[2147]_  | \new_[5228]_ ;
  assign \new_[5233]_  = \new_[2142]_  | \new_[2143]_ ;
  assign \new_[5234]_  = \new_[2144]_  | \new_[5233]_ ;
  assign \new_[5235]_  = \new_[5234]_  | \new_[5229]_ ;
  assign \new_[5239]_  = \new_[2139]_  | \new_[2140]_ ;
  assign \new_[5240]_  = \new_[2141]_  | \new_[5239]_ ;
  assign \new_[5243]_  = \new_[2137]_  | \new_[2138]_ ;
  assign \new_[5246]_  = \new_[2135]_  | \new_[2136]_ ;
  assign \new_[5247]_  = \new_[5246]_  | \new_[5243]_ ;
  assign \new_[5248]_  = \new_[5247]_  | \new_[5240]_ ;
  assign \new_[5249]_  = \new_[5248]_  | \new_[5235]_ ;
  assign \new_[5250]_  = \new_[5249]_  | \new_[5224]_ ;
  assign \new_[5251]_  = \new_[5250]_  | \new_[5201]_ ;
  assign \new_[5255]_  = \new_[2132]_  | \new_[2133]_ ;
  assign \new_[5256]_  = \new_[2134]_  | \new_[5255]_ ;
  assign \new_[5260]_  = \new_[2129]_  | \new_[2130]_ ;
  assign \new_[5261]_  = \new_[2131]_  | \new_[5260]_ ;
  assign \new_[5262]_  = \new_[5261]_  | \new_[5256]_ ;
  assign \new_[5266]_  = \new_[2126]_  | \new_[2127]_ ;
  assign \new_[5267]_  = \new_[2128]_  | \new_[5266]_ ;
  assign \new_[5271]_  = \new_[2123]_  | \new_[2124]_ ;
  assign \new_[5272]_  = \new_[2125]_  | \new_[5271]_ ;
  assign \new_[5273]_  = \new_[5272]_  | \new_[5267]_ ;
  assign \new_[5274]_  = \new_[5273]_  | \new_[5262]_ ;
  assign \new_[5278]_  = \new_[2120]_  | \new_[2121]_ ;
  assign \new_[5279]_  = \new_[2122]_  | \new_[5278]_ ;
  assign \new_[5283]_  = \new_[2117]_  | \new_[2118]_ ;
  assign \new_[5284]_  = \new_[2119]_  | \new_[5283]_ ;
  assign \new_[5285]_  = \new_[5284]_  | \new_[5279]_ ;
  assign \new_[5289]_  = \new_[2114]_  | \new_[2115]_ ;
  assign \new_[5290]_  = \new_[2116]_  | \new_[5289]_ ;
  assign \new_[5293]_  = \new_[2112]_  | \new_[2113]_ ;
  assign \new_[5296]_  = \new_[2110]_  | \new_[2111]_ ;
  assign \new_[5297]_  = \new_[5296]_  | \new_[5293]_ ;
  assign \new_[5298]_  = \new_[5297]_  | \new_[5290]_ ;
  assign \new_[5299]_  = \new_[5298]_  | \new_[5285]_ ;
  assign \new_[5300]_  = \new_[5299]_  | \new_[5274]_ ;
  assign \new_[5304]_  = \new_[2107]_  | \new_[2108]_ ;
  assign \new_[5305]_  = \new_[2109]_  | \new_[5304]_ ;
  assign \new_[5309]_  = \new_[2104]_  | \new_[2105]_ ;
  assign \new_[5310]_  = \new_[2106]_  | \new_[5309]_ ;
  assign \new_[5311]_  = \new_[5310]_  | \new_[5305]_ ;
  assign \new_[5315]_  = \new_[2101]_  | \new_[2102]_ ;
  assign \new_[5316]_  = \new_[2103]_  | \new_[5315]_ ;
  assign \new_[5320]_  = \new_[2098]_  | \new_[2099]_ ;
  assign \new_[5321]_  = \new_[2100]_  | \new_[5320]_ ;
  assign \new_[5322]_  = \new_[5321]_  | \new_[5316]_ ;
  assign \new_[5323]_  = \new_[5322]_  | \new_[5311]_ ;
  assign \new_[5327]_  = \new_[2095]_  | \new_[2096]_ ;
  assign \new_[5328]_  = \new_[2097]_  | \new_[5327]_ ;
  assign \new_[5332]_  = \new_[2092]_  | \new_[2093]_ ;
  assign \new_[5333]_  = \new_[2094]_  | \new_[5332]_ ;
  assign \new_[5334]_  = \new_[5333]_  | \new_[5328]_ ;
  assign \new_[5338]_  = \new_[2089]_  | \new_[2090]_ ;
  assign \new_[5339]_  = \new_[2091]_  | \new_[5338]_ ;
  assign \new_[5342]_  = \new_[2087]_  | \new_[2088]_ ;
  assign \new_[5345]_  = \new_[2085]_  | \new_[2086]_ ;
  assign \new_[5346]_  = \new_[5345]_  | \new_[5342]_ ;
  assign \new_[5347]_  = \new_[5346]_  | \new_[5339]_ ;
  assign \new_[5348]_  = \new_[5347]_  | \new_[5334]_ ;
  assign \new_[5349]_  = \new_[5348]_  | \new_[5323]_ ;
  assign \new_[5350]_  = \new_[5349]_  | \new_[5300]_ ;
  assign \new_[5351]_  = \new_[5350]_  | \new_[5251]_ ;
  assign \new_[5355]_  = \new_[2082]_  | \new_[2083]_ ;
  assign \new_[5356]_  = \new_[2084]_  | \new_[5355]_ ;
  assign \new_[5360]_  = \new_[2079]_  | \new_[2080]_ ;
  assign \new_[5361]_  = \new_[2081]_  | \new_[5360]_ ;
  assign \new_[5362]_  = \new_[5361]_  | \new_[5356]_ ;
  assign \new_[5366]_  = \new_[2076]_  | \new_[2077]_ ;
  assign \new_[5367]_  = \new_[2078]_  | \new_[5366]_ ;
  assign \new_[5371]_  = \new_[2073]_  | \new_[2074]_ ;
  assign \new_[5372]_  = \new_[2075]_  | \new_[5371]_ ;
  assign \new_[5373]_  = \new_[5372]_  | \new_[5367]_ ;
  assign \new_[5374]_  = \new_[5373]_  | \new_[5362]_ ;
  assign \new_[5378]_  = \new_[2070]_  | \new_[2071]_ ;
  assign \new_[5379]_  = \new_[2072]_  | \new_[5378]_ ;
  assign \new_[5383]_  = \new_[2067]_  | \new_[2068]_ ;
  assign \new_[5384]_  = \new_[2069]_  | \new_[5383]_ ;
  assign \new_[5385]_  = \new_[5384]_  | \new_[5379]_ ;
  assign \new_[5389]_  = \new_[2064]_  | \new_[2065]_ ;
  assign \new_[5390]_  = \new_[2066]_  | \new_[5389]_ ;
  assign \new_[5393]_  = \new_[2062]_  | \new_[2063]_ ;
  assign \new_[5396]_  = \new_[2060]_  | \new_[2061]_ ;
  assign \new_[5397]_  = \new_[5396]_  | \new_[5393]_ ;
  assign \new_[5398]_  = \new_[5397]_  | \new_[5390]_ ;
  assign \new_[5399]_  = \new_[5398]_  | \new_[5385]_ ;
  assign \new_[5400]_  = \new_[5399]_  | \new_[5374]_ ;
  assign \new_[5404]_  = \new_[2057]_  | \new_[2058]_ ;
  assign \new_[5405]_  = \new_[2059]_  | \new_[5404]_ ;
  assign \new_[5409]_  = \new_[2054]_  | \new_[2055]_ ;
  assign \new_[5410]_  = \new_[2056]_  | \new_[5409]_ ;
  assign \new_[5411]_  = \new_[5410]_  | \new_[5405]_ ;
  assign \new_[5415]_  = \new_[2051]_  | \new_[2052]_ ;
  assign \new_[5416]_  = \new_[2053]_  | \new_[5415]_ ;
  assign \new_[5420]_  = \new_[2048]_  | \new_[2049]_ ;
  assign \new_[5421]_  = \new_[2050]_  | \new_[5420]_ ;
  assign \new_[5422]_  = \new_[5421]_  | \new_[5416]_ ;
  assign \new_[5423]_  = \new_[5422]_  | \new_[5411]_ ;
  assign \new_[5427]_  = \new_[2045]_  | \new_[2046]_ ;
  assign \new_[5428]_  = \new_[2047]_  | \new_[5427]_ ;
  assign \new_[5432]_  = \new_[2042]_  | \new_[2043]_ ;
  assign \new_[5433]_  = \new_[2044]_  | \new_[5432]_ ;
  assign \new_[5434]_  = \new_[5433]_  | \new_[5428]_ ;
  assign \new_[5438]_  = \new_[2039]_  | \new_[2040]_ ;
  assign \new_[5439]_  = \new_[2041]_  | \new_[5438]_ ;
  assign \new_[5442]_  = \new_[2037]_  | \new_[2038]_ ;
  assign \new_[5445]_  = \new_[2035]_  | \new_[2036]_ ;
  assign \new_[5446]_  = \new_[5445]_  | \new_[5442]_ ;
  assign \new_[5447]_  = \new_[5446]_  | \new_[5439]_ ;
  assign \new_[5448]_  = \new_[5447]_  | \new_[5434]_ ;
  assign \new_[5449]_  = \new_[5448]_  | \new_[5423]_ ;
  assign \new_[5450]_  = \new_[5449]_  | \new_[5400]_ ;
  assign \new_[5454]_  = \new_[2032]_  | \new_[2033]_ ;
  assign \new_[5455]_  = \new_[2034]_  | \new_[5454]_ ;
  assign \new_[5459]_  = \new_[2029]_  | \new_[2030]_ ;
  assign \new_[5460]_  = \new_[2031]_  | \new_[5459]_ ;
  assign \new_[5461]_  = \new_[5460]_  | \new_[5455]_ ;
  assign \new_[5465]_  = \new_[2026]_  | \new_[2027]_ ;
  assign \new_[5466]_  = \new_[2028]_  | \new_[5465]_ ;
  assign \new_[5470]_  = \new_[2023]_  | \new_[2024]_ ;
  assign \new_[5471]_  = \new_[2025]_  | \new_[5470]_ ;
  assign \new_[5472]_  = \new_[5471]_  | \new_[5466]_ ;
  assign \new_[5473]_  = \new_[5472]_  | \new_[5461]_ ;
  assign \new_[5477]_  = \new_[2020]_  | \new_[2021]_ ;
  assign \new_[5478]_  = \new_[2022]_  | \new_[5477]_ ;
  assign \new_[5482]_  = \new_[2017]_  | \new_[2018]_ ;
  assign \new_[5483]_  = \new_[2019]_  | \new_[5482]_ ;
  assign \new_[5484]_  = \new_[5483]_  | \new_[5478]_ ;
  assign \new_[5488]_  = \new_[2014]_  | \new_[2015]_ ;
  assign \new_[5489]_  = \new_[2016]_  | \new_[5488]_ ;
  assign \new_[5492]_  = \new_[2012]_  | \new_[2013]_ ;
  assign \new_[5495]_  = \new_[2010]_  | \new_[2011]_ ;
  assign \new_[5496]_  = \new_[5495]_  | \new_[5492]_ ;
  assign \new_[5497]_  = \new_[5496]_  | \new_[5489]_ ;
  assign \new_[5498]_  = \new_[5497]_  | \new_[5484]_ ;
  assign \new_[5499]_  = \new_[5498]_  | \new_[5473]_ ;
  assign \new_[5503]_  = \new_[2007]_  | \new_[2008]_ ;
  assign \new_[5504]_  = \new_[2009]_  | \new_[5503]_ ;
  assign \new_[5508]_  = \new_[2004]_  | \new_[2005]_ ;
  assign \new_[5509]_  = \new_[2006]_  | \new_[5508]_ ;
  assign \new_[5510]_  = \new_[5509]_  | \new_[5504]_ ;
  assign \new_[5514]_  = \new_[2001]_  | \new_[2002]_ ;
  assign \new_[5515]_  = \new_[2003]_  | \new_[5514]_ ;
  assign \new_[5519]_  = \new_[1998]_  | \new_[1999]_ ;
  assign \new_[5520]_  = \new_[2000]_  | \new_[5519]_ ;
  assign \new_[5521]_  = \new_[5520]_  | \new_[5515]_ ;
  assign \new_[5522]_  = \new_[5521]_  | \new_[5510]_ ;
  assign \new_[5526]_  = \new_[1995]_  | \new_[1996]_ ;
  assign \new_[5527]_  = \new_[1997]_  | \new_[5526]_ ;
  assign \new_[5531]_  = \new_[1992]_  | \new_[1993]_ ;
  assign \new_[5532]_  = \new_[1994]_  | \new_[5531]_ ;
  assign \new_[5533]_  = \new_[5532]_  | \new_[5527]_ ;
  assign \new_[5537]_  = \new_[1989]_  | \new_[1990]_ ;
  assign \new_[5538]_  = \new_[1991]_  | \new_[5537]_ ;
  assign \new_[5541]_  = \new_[1987]_  | \new_[1988]_ ;
  assign \new_[5544]_  = \new_[1985]_  | \new_[1986]_ ;
  assign \new_[5545]_  = \new_[5544]_  | \new_[5541]_ ;
  assign \new_[5546]_  = \new_[5545]_  | \new_[5538]_ ;
  assign \new_[5547]_  = \new_[5546]_  | \new_[5533]_ ;
  assign \new_[5548]_  = \new_[5547]_  | \new_[5522]_ ;
  assign \new_[5549]_  = \new_[5548]_  | \new_[5499]_ ;
  assign \new_[5550]_  = \new_[5549]_  | \new_[5450]_ ;
  assign \new_[5551]_  = \new_[5550]_  | \new_[5351]_ ;
  assign \new_[5552]_  = \new_[5551]_  | \new_[5154]_ ;
  assign \new_[5556]_  = \new_[1982]_  | \new_[1983]_ ;
  assign \new_[5557]_  = \new_[1984]_  | \new_[5556]_ ;
  assign \new_[5561]_  = \new_[1979]_  | \new_[1980]_ ;
  assign \new_[5562]_  = \new_[1981]_  | \new_[5561]_ ;
  assign \new_[5563]_  = \new_[5562]_  | \new_[5557]_ ;
  assign \new_[5567]_  = \new_[1976]_  | \new_[1977]_ ;
  assign \new_[5568]_  = \new_[1978]_  | \new_[5567]_ ;
  assign \new_[5572]_  = \new_[1973]_  | \new_[1974]_ ;
  assign \new_[5573]_  = \new_[1975]_  | \new_[5572]_ ;
  assign \new_[5574]_  = \new_[5573]_  | \new_[5568]_ ;
  assign \new_[5575]_  = \new_[5574]_  | \new_[5563]_ ;
  assign \new_[5579]_  = \new_[1970]_  | \new_[1971]_ ;
  assign \new_[5580]_  = \new_[1972]_  | \new_[5579]_ ;
  assign \new_[5584]_  = \new_[1967]_  | \new_[1968]_ ;
  assign \new_[5585]_  = \new_[1969]_  | \new_[5584]_ ;
  assign \new_[5586]_  = \new_[5585]_  | \new_[5580]_ ;
  assign \new_[5590]_  = \new_[1964]_  | \new_[1965]_ ;
  assign \new_[5591]_  = \new_[1966]_  | \new_[5590]_ ;
  assign \new_[5595]_  = \new_[1961]_  | \new_[1962]_ ;
  assign \new_[5596]_  = \new_[1963]_  | \new_[5595]_ ;
  assign \new_[5597]_  = \new_[5596]_  | \new_[5591]_ ;
  assign \new_[5598]_  = \new_[5597]_  | \new_[5586]_ ;
  assign \new_[5599]_  = \new_[5598]_  | \new_[5575]_ ;
  assign \new_[5603]_  = \new_[1958]_  | \new_[1959]_ ;
  assign \new_[5604]_  = \new_[1960]_  | \new_[5603]_ ;
  assign \new_[5608]_  = \new_[1955]_  | \new_[1956]_ ;
  assign \new_[5609]_  = \new_[1957]_  | \new_[5608]_ ;
  assign \new_[5610]_  = \new_[5609]_  | \new_[5604]_ ;
  assign \new_[5614]_  = \new_[1952]_  | \new_[1953]_ ;
  assign \new_[5615]_  = \new_[1954]_  | \new_[5614]_ ;
  assign \new_[5619]_  = \new_[1949]_  | \new_[1950]_ ;
  assign \new_[5620]_  = \new_[1951]_  | \new_[5619]_ ;
  assign \new_[5621]_  = \new_[5620]_  | \new_[5615]_ ;
  assign \new_[5622]_  = \new_[5621]_  | \new_[5610]_ ;
  assign \new_[5626]_  = \new_[1946]_  | \new_[1947]_ ;
  assign \new_[5627]_  = \new_[1948]_  | \new_[5626]_ ;
  assign \new_[5631]_  = \new_[1943]_  | \new_[1944]_ ;
  assign \new_[5632]_  = \new_[1945]_  | \new_[5631]_ ;
  assign \new_[5633]_  = \new_[5632]_  | \new_[5627]_ ;
  assign \new_[5637]_  = \new_[1940]_  | \new_[1941]_ ;
  assign \new_[5638]_  = \new_[1942]_  | \new_[5637]_ ;
  assign \new_[5641]_  = \new_[1938]_  | \new_[1939]_ ;
  assign \new_[5644]_  = \new_[1936]_  | \new_[1937]_ ;
  assign \new_[5645]_  = \new_[5644]_  | \new_[5641]_ ;
  assign \new_[5646]_  = \new_[5645]_  | \new_[5638]_ ;
  assign \new_[5647]_  = \new_[5646]_  | \new_[5633]_ ;
  assign \new_[5648]_  = \new_[5647]_  | \new_[5622]_ ;
  assign \new_[5649]_  = \new_[5648]_  | \new_[5599]_ ;
  assign \new_[5653]_  = \new_[1933]_  | \new_[1934]_ ;
  assign \new_[5654]_  = \new_[1935]_  | \new_[5653]_ ;
  assign \new_[5658]_  = \new_[1930]_  | \new_[1931]_ ;
  assign \new_[5659]_  = \new_[1932]_  | \new_[5658]_ ;
  assign \new_[5660]_  = \new_[5659]_  | \new_[5654]_ ;
  assign \new_[5664]_  = \new_[1927]_  | \new_[1928]_ ;
  assign \new_[5665]_  = \new_[1929]_  | \new_[5664]_ ;
  assign \new_[5669]_  = \new_[1924]_  | \new_[1925]_ ;
  assign \new_[5670]_  = \new_[1926]_  | \new_[5669]_ ;
  assign \new_[5671]_  = \new_[5670]_  | \new_[5665]_ ;
  assign \new_[5672]_  = \new_[5671]_  | \new_[5660]_ ;
  assign \new_[5676]_  = \new_[1921]_  | \new_[1922]_ ;
  assign \new_[5677]_  = \new_[1923]_  | \new_[5676]_ ;
  assign \new_[5681]_  = \new_[1918]_  | \new_[1919]_ ;
  assign \new_[5682]_  = \new_[1920]_  | \new_[5681]_ ;
  assign \new_[5683]_  = \new_[5682]_  | \new_[5677]_ ;
  assign \new_[5687]_  = \new_[1915]_  | \new_[1916]_ ;
  assign \new_[5688]_  = \new_[1917]_  | \new_[5687]_ ;
  assign \new_[5691]_  = \new_[1913]_  | \new_[1914]_ ;
  assign \new_[5694]_  = \new_[1911]_  | \new_[1912]_ ;
  assign \new_[5695]_  = \new_[5694]_  | \new_[5691]_ ;
  assign \new_[5696]_  = \new_[5695]_  | \new_[5688]_ ;
  assign \new_[5697]_  = \new_[5696]_  | \new_[5683]_ ;
  assign \new_[5698]_  = \new_[5697]_  | \new_[5672]_ ;
  assign \new_[5702]_  = \new_[1908]_  | \new_[1909]_ ;
  assign \new_[5703]_  = \new_[1910]_  | \new_[5702]_ ;
  assign \new_[5707]_  = \new_[1905]_  | \new_[1906]_ ;
  assign \new_[5708]_  = \new_[1907]_  | \new_[5707]_ ;
  assign \new_[5709]_  = \new_[5708]_  | \new_[5703]_ ;
  assign \new_[5713]_  = \new_[1902]_  | \new_[1903]_ ;
  assign \new_[5714]_  = \new_[1904]_  | \new_[5713]_ ;
  assign \new_[5718]_  = \new_[1899]_  | \new_[1900]_ ;
  assign \new_[5719]_  = \new_[1901]_  | \new_[5718]_ ;
  assign \new_[5720]_  = \new_[5719]_  | \new_[5714]_ ;
  assign \new_[5721]_  = \new_[5720]_  | \new_[5709]_ ;
  assign \new_[5725]_  = \new_[1896]_  | \new_[1897]_ ;
  assign \new_[5726]_  = \new_[1898]_  | \new_[5725]_ ;
  assign \new_[5730]_  = \new_[1893]_  | \new_[1894]_ ;
  assign \new_[5731]_  = \new_[1895]_  | \new_[5730]_ ;
  assign \new_[5732]_  = \new_[5731]_  | \new_[5726]_ ;
  assign \new_[5736]_  = \new_[1890]_  | \new_[1891]_ ;
  assign \new_[5737]_  = \new_[1892]_  | \new_[5736]_ ;
  assign \new_[5740]_  = \new_[1888]_  | \new_[1889]_ ;
  assign \new_[5743]_  = \new_[1886]_  | \new_[1887]_ ;
  assign \new_[5744]_  = \new_[5743]_  | \new_[5740]_ ;
  assign \new_[5745]_  = \new_[5744]_  | \new_[5737]_ ;
  assign \new_[5746]_  = \new_[5745]_  | \new_[5732]_ ;
  assign \new_[5747]_  = \new_[5746]_  | \new_[5721]_ ;
  assign \new_[5748]_  = \new_[5747]_  | \new_[5698]_ ;
  assign \new_[5749]_  = \new_[5748]_  | \new_[5649]_ ;
  assign \new_[5753]_  = \new_[1883]_  | \new_[1884]_ ;
  assign \new_[5754]_  = \new_[1885]_  | \new_[5753]_ ;
  assign \new_[5758]_  = \new_[1880]_  | \new_[1881]_ ;
  assign \new_[5759]_  = \new_[1882]_  | \new_[5758]_ ;
  assign \new_[5760]_  = \new_[5759]_  | \new_[5754]_ ;
  assign \new_[5764]_  = \new_[1877]_  | \new_[1878]_ ;
  assign \new_[5765]_  = \new_[1879]_  | \new_[5764]_ ;
  assign \new_[5769]_  = \new_[1874]_  | \new_[1875]_ ;
  assign \new_[5770]_  = \new_[1876]_  | \new_[5769]_ ;
  assign \new_[5771]_  = \new_[5770]_  | \new_[5765]_ ;
  assign \new_[5772]_  = \new_[5771]_  | \new_[5760]_ ;
  assign \new_[5776]_  = \new_[1871]_  | \new_[1872]_ ;
  assign \new_[5777]_  = \new_[1873]_  | \new_[5776]_ ;
  assign \new_[5781]_  = \new_[1868]_  | \new_[1869]_ ;
  assign \new_[5782]_  = \new_[1870]_  | \new_[5781]_ ;
  assign \new_[5783]_  = \new_[5782]_  | \new_[5777]_ ;
  assign \new_[5787]_  = \new_[1865]_  | \new_[1866]_ ;
  assign \new_[5788]_  = \new_[1867]_  | \new_[5787]_ ;
  assign \new_[5792]_  = \new_[1862]_  | \new_[1863]_ ;
  assign \new_[5793]_  = \new_[1864]_  | \new_[5792]_ ;
  assign \new_[5794]_  = \new_[5793]_  | \new_[5788]_ ;
  assign \new_[5795]_  = \new_[5794]_  | \new_[5783]_ ;
  assign \new_[5796]_  = \new_[5795]_  | \new_[5772]_ ;
  assign \new_[5800]_  = \new_[1859]_  | \new_[1860]_ ;
  assign \new_[5801]_  = \new_[1861]_  | \new_[5800]_ ;
  assign \new_[5805]_  = \new_[1856]_  | \new_[1857]_ ;
  assign \new_[5806]_  = \new_[1858]_  | \new_[5805]_ ;
  assign \new_[5807]_  = \new_[5806]_  | \new_[5801]_ ;
  assign \new_[5811]_  = \new_[1853]_  | \new_[1854]_ ;
  assign \new_[5812]_  = \new_[1855]_  | \new_[5811]_ ;
  assign \new_[5816]_  = \new_[1850]_  | \new_[1851]_ ;
  assign \new_[5817]_  = \new_[1852]_  | \new_[5816]_ ;
  assign \new_[5818]_  = \new_[5817]_  | \new_[5812]_ ;
  assign \new_[5819]_  = \new_[5818]_  | \new_[5807]_ ;
  assign \new_[5823]_  = \new_[1847]_  | \new_[1848]_ ;
  assign \new_[5824]_  = \new_[1849]_  | \new_[5823]_ ;
  assign \new_[5828]_  = \new_[1844]_  | \new_[1845]_ ;
  assign \new_[5829]_  = \new_[1846]_  | \new_[5828]_ ;
  assign \new_[5830]_  = \new_[5829]_  | \new_[5824]_ ;
  assign \new_[5834]_  = \new_[1841]_  | \new_[1842]_ ;
  assign \new_[5835]_  = \new_[1843]_  | \new_[5834]_ ;
  assign \new_[5838]_  = \new_[1839]_  | \new_[1840]_ ;
  assign \new_[5841]_  = \new_[1837]_  | \new_[1838]_ ;
  assign \new_[5842]_  = \new_[5841]_  | \new_[5838]_ ;
  assign \new_[5843]_  = \new_[5842]_  | \new_[5835]_ ;
  assign \new_[5844]_  = \new_[5843]_  | \new_[5830]_ ;
  assign \new_[5845]_  = \new_[5844]_  | \new_[5819]_ ;
  assign \new_[5846]_  = \new_[5845]_  | \new_[5796]_ ;
  assign \new_[5850]_  = \new_[1834]_  | \new_[1835]_ ;
  assign \new_[5851]_  = \new_[1836]_  | \new_[5850]_ ;
  assign \new_[5855]_  = \new_[1831]_  | \new_[1832]_ ;
  assign \new_[5856]_  = \new_[1833]_  | \new_[5855]_ ;
  assign \new_[5857]_  = \new_[5856]_  | \new_[5851]_ ;
  assign \new_[5861]_  = \new_[1828]_  | \new_[1829]_ ;
  assign \new_[5862]_  = \new_[1830]_  | \new_[5861]_ ;
  assign \new_[5866]_  = \new_[1825]_  | \new_[1826]_ ;
  assign \new_[5867]_  = \new_[1827]_  | \new_[5866]_ ;
  assign \new_[5868]_  = \new_[5867]_  | \new_[5862]_ ;
  assign \new_[5869]_  = \new_[5868]_  | \new_[5857]_ ;
  assign \new_[5873]_  = \new_[1822]_  | \new_[1823]_ ;
  assign \new_[5874]_  = \new_[1824]_  | \new_[5873]_ ;
  assign \new_[5878]_  = \new_[1819]_  | \new_[1820]_ ;
  assign \new_[5879]_  = \new_[1821]_  | \new_[5878]_ ;
  assign \new_[5880]_  = \new_[5879]_  | \new_[5874]_ ;
  assign \new_[5884]_  = \new_[1816]_  | \new_[1817]_ ;
  assign \new_[5885]_  = \new_[1818]_  | \new_[5884]_ ;
  assign \new_[5888]_  = \new_[1814]_  | \new_[1815]_ ;
  assign \new_[5891]_  = \new_[1812]_  | \new_[1813]_ ;
  assign \new_[5892]_  = \new_[5891]_  | \new_[5888]_ ;
  assign \new_[5893]_  = \new_[5892]_  | \new_[5885]_ ;
  assign \new_[5894]_  = \new_[5893]_  | \new_[5880]_ ;
  assign \new_[5895]_  = \new_[5894]_  | \new_[5869]_ ;
  assign \new_[5899]_  = \new_[1809]_  | \new_[1810]_ ;
  assign \new_[5900]_  = \new_[1811]_  | \new_[5899]_ ;
  assign \new_[5904]_  = \new_[1806]_  | \new_[1807]_ ;
  assign \new_[5905]_  = \new_[1808]_  | \new_[5904]_ ;
  assign \new_[5906]_  = \new_[5905]_  | \new_[5900]_ ;
  assign \new_[5910]_  = \new_[1803]_  | \new_[1804]_ ;
  assign \new_[5911]_  = \new_[1805]_  | \new_[5910]_ ;
  assign \new_[5915]_  = \new_[1800]_  | \new_[1801]_ ;
  assign \new_[5916]_  = \new_[1802]_  | \new_[5915]_ ;
  assign \new_[5917]_  = \new_[5916]_  | \new_[5911]_ ;
  assign \new_[5918]_  = \new_[5917]_  | \new_[5906]_ ;
  assign \new_[5922]_  = \new_[1797]_  | \new_[1798]_ ;
  assign \new_[5923]_  = \new_[1799]_  | \new_[5922]_ ;
  assign \new_[5927]_  = \new_[1794]_  | \new_[1795]_ ;
  assign \new_[5928]_  = \new_[1796]_  | \new_[5927]_ ;
  assign \new_[5929]_  = \new_[5928]_  | \new_[5923]_ ;
  assign \new_[5933]_  = \new_[1791]_  | \new_[1792]_ ;
  assign \new_[5934]_  = \new_[1793]_  | \new_[5933]_ ;
  assign \new_[5937]_  = \new_[1789]_  | \new_[1790]_ ;
  assign \new_[5940]_  = \new_[1787]_  | \new_[1788]_ ;
  assign \new_[5941]_  = \new_[5940]_  | \new_[5937]_ ;
  assign \new_[5942]_  = \new_[5941]_  | \new_[5934]_ ;
  assign \new_[5943]_  = \new_[5942]_  | \new_[5929]_ ;
  assign \new_[5944]_  = \new_[5943]_  | \new_[5918]_ ;
  assign \new_[5945]_  = \new_[5944]_  | \new_[5895]_ ;
  assign \new_[5946]_  = \new_[5945]_  | \new_[5846]_ ;
  assign \new_[5947]_  = \new_[5946]_  | \new_[5749]_ ;
  assign \new_[5951]_  = \new_[1784]_  | \new_[1785]_ ;
  assign \new_[5952]_  = \new_[1786]_  | \new_[5951]_ ;
  assign \new_[5956]_  = \new_[1781]_  | \new_[1782]_ ;
  assign \new_[5957]_  = \new_[1783]_  | \new_[5956]_ ;
  assign \new_[5958]_  = \new_[5957]_  | \new_[5952]_ ;
  assign \new_[5962]_  = \new_[1778]_  | \new_[1779]_ ;
  assign \new_[5963]_  = \new_[1780]_  | \new_[5962]_ ;
  assign \new_[5967]_  = \new_[1775]_  | \new_[1776]_ ;
  assign \new_[5968]_  = \new_[1777]_  | \new_[5967]_ ;
  assign \new_[5969]_  = \new_[5968]_  | \new_[5963]_ ;
  assign \new_[5970]_  = \new_[5969]_  | \new_[5958]_ ;
  assign \new_[5974]_  = \new_[1772]_  | \new_[1773]_ ;
  assign \new_[5975]_  = \new_[1774]_  | \new_[5974]_ ;
  assign \new_[5979]_  = \new_[1769]_  | \new_[1770]_ ;
  assign \new_[5980]_  = \new_[1771]_  | \new_[5979]_ ;
  assign \new_[5981]_  = \new_[5980]_  | \new_[5975]_ ;
  assign \new_[5985]_  = \new_[1766]_  | \new_[1767]_ ;
  assign \new_[5986]_  = \new_[1768]_  | \new_[5985]_ ;
  assign \new_[5990]_  = \new_[1763]_  | \new_[1764]_ ;
  assign \new_[5991]_  = \new_[1765]_  | \new_[5990]_ ;
  assign \new_[5992]_  = \new_[5991]_  | \new_[5986]_ ;
  assign \new_[5993]_  = \new_[5992]_  | \new_[5981]_ ;
  assign \new_[5994]_  = \new_[5993]_  | \new_[5970]_ ;
  assign \new_[5998]_  = \new_[1760]_  | \new_[1761]_ ;
  assign \new_[5999]_  = \new_[1762]_  | \new_[5998]_ ;
  assign \new_[6003]_  = \new_[1757]_  | \new_[1758]_ ;
  assign \new_[6004]_  = \new_[1759]_  | \new_[6003]_ ;
  assign \new_[6005]_  = \new_[6004]_  | \new_[5999]_ ;
  assign \new_[6009]_  = \new_[1754]_  | \new_[1755]_ ;
  assign \new_[6010]_  = \new_[1756]_  | \new_[6009]_ ;
  assign \new_[6014]_  = \new_[1751]_  | \new_[1752]_ ;
  assign \new_[6015]_  = \new_[1753]_  | \new_[6014]_ ;
  assign \new_[6016]_  = \new_[6015]_  | \new_[6010]_ ;
  assign \new_[6017]_  = \new_[6016]_  | \new_[6005]_ ;
  assign \new_[6021]_  = \new_[1748]_  | \new_[1749]_ ;
  assign \new_[6022]_  = \new_[1750]_  | \new_[6021]_ ;
  assign \new_[6026]_  = \new_[1745]_  | \new_[1746]_ ;
  assign \new_[6027]_  = \new_[1747]_  | \new_[6026]_ ;
  assign \new_[6028]_  = \new_[6027]_  | \new_[6022]_ ;
  assign \new_[6032]_  = \new_[1742]_  | \new_[1743]_ ;
  assign \new_[6033]_  = \new_[1744]_  | \new_[6032]_ ;
  assign \new_[6036]_  = \new_[1740]_  | \new_[1741]_ ;
  assign \new_[6039]_  = \new_[1738]_  | \new_[1739]_ ;
  assign \new_[6040]_  = \new_[6039]_  | \new_[6036]_ ;
  assign \new_[6041]_  = \new_[6040]_  | \new_[6033]_ ;
  assign \new_[6042]_  = \new_[6041]_  | \new_[6028]_ ;
  assign \new_[6043]_  = \new_[6042]_  | \new_[6017]_ ;
  assign \new_[6044]_  = \new_[6043]_  | \new_[5994]_ ;
  assign \new_[6048]_  = \new_[1735]_  | \new_[1736]_ ;
  assign \new_[6049]_  = \new_[1737]_  | \new_[6048]_ ;
  assign \new_[6053]_  = \new_[1732]_  | \new_[1733]_ ;
  assign \new_[6054]_  = \new_[1734]_  | \new_[6053]_ ;
  assign \new_[6055]_  = \new_[6054]_  | \new_[6049]_ ;
  assign \new_[6059]_  = \new_[1729]_  | \new_[1730]_ ;
  assign \new_[6060]_  = \new_[1731]_  | \new_[6059]_ ;
  assign \new_[6064]_  = \new_[1726]_  | \new_[1727]_ ;
  assign \new_[6065]_  = \new_[1728]_  | \new_[6064]_ ;
  assign \new_[6066]_  = \new_[6065]_  | \new_[6060]_ ;
  assign \new_[6067]_  = \new_[6066]_  | \new_[6055]_ ;
  assign \new_[6071]_  = \new_[1723]_  | \new_[1724]_ ;
  assign \new_[6072]_  = \new_[1725]_  | \new_[6071]_ ;
  assign \new_[6076]_  = \new_[1720]_  | \new_[1721]_ ;
  assign \new_[6077]_  = \new_[1722]_  | \new_[6076]_ ;
  assign \new_[6078]_  = \new_[6077]_  | \new_[6072]_ ;
  assign \new_[6082]_  = \new_[1717]_  | \new_[1718]_ ;
  assign \new_[6083]_  = \new_[1719]_  | \new_[6082]_ ;
  assign \new_[6086]_  = \new_[1715]_  | \new_[1716]_ ;
  assign \new_[6089]_  = \new_[1713]_  | \new_[1714]_ ;
  assign \new_[6090]_  = \new_[6089]_  | \new_[6086]_ ;
  assign \new_[6091]_  = \new_[6090]_  | \new_[6083]_ ;
  assign \new_[6092]_  = \new_[6091]_  | \new_[6078]_ ;
  assign \new_[6093]_  = \new_[6092]_  | \new_[6067]_ ;
  assign \new_[6097]_  = \new_[1710]_  | \new_[1711]_ ;
  assign \new_[6098]_  = \new_[1712]_  | \new_[6097]_ ;
  assign \new_[6102]_  = \new_[1707]_  | \new_[1708]_ ;
  assign \new_[6103]_  = \new_[1709]_  | \new_[6102]_ ;
  assign \new_[6104]_  = \new_[6103]_  | \new_[6098]_ ;
  assign \new_[6108]_  = \new_[1704]_  | \new_[1705]_ ;
  assign \new_[6109]_  = \new_[1706]_  | \new_[6108]_ ;
  assign \new_[6113]_  = \new_[1701]_  | \new_[1702]_ ;
  assign \new_[6114]_  = \new_[1703]_  | \new_[6113]_ ;
  assign \new_[6115]_  = \new_[6114]_  | \new_[6109]_ ;
  assign \new_[6116]_  = \new_[6115]_  | \new_[6104]_ ;
  assign \new_[6120]_  = \new_[1698]_  | \new_[1699]_ ;
  assign \new_[6121]_  = \new_[1700]_  | \new_[6120]_ ;
  assign \new_[6125]_  = \new_[1695]_  | \new_[1696]_ ;
  assign \new_[6126]_  = \new_[1697]_  | \new_[6125]_ ;
  assign \new_[6127]_  = \new_[6126]_  | \new_[6121]_ ;
  assign \new_[6131]_  = \new_[1692]_  | \new_[1693]_ ;
  assign \new_[6132]_  = \new_[1694]_  | \new_[6131]_ ;
  assign \new_[6135]_  = \new_[1690]_  | \new_[1691]_ ;
  assign \new_[6138]_  = \new_[1688]_  | \new_[1689]_ ;
  assign \new_[6139]_  = \new_[6138]_  | \new_[6135]_ ;
  assign \new_[6140]_  = \new_[6139]_  | \new_[6132]_ ;
  assign \new_[6141]_  = \new_[6140]_  | \new_[6127]_ ;
  assign \new_[6142]_  = \new_[6141]_  | \new_[6116]_ ;
  assign \new_[6143]_  = \new_[6142]_  | \new_[6093]_ ;
  assign \new_[6144]_  = \new_[6143]_  | \new_[6044]_ ;
  assign \new_[6148]_  = \new_[1685]_  | \new_[1686]_ ;
  assign \new_[6149]_  = \new_[1687]_  | \new_[6148]_ ;
  assign \new_[6153]_  = \new_[1682]_  | \new_[1683]_ ;
  assign \new_[6154]_  = \new_[1684]_  | \new_[6153]_ ;
  assign \new_[6155]_  = \new_[6154]_  | \new_[6149]_ ;
  assign \new_[6159]_  = \new_[1679]_  | \new_[1680]_ ;
  assign \new_[6160]_  = \new_[1681]_  | \new_[6159]_ ;
  assign \new_[6164]_  = \new_[1676]_  | \new_[1677]_ ;
  assign \new_[6165]_  = \new_[1678]_  | \new_[6164]_ ;
  assign \new_[6166]_  = \new_[6165]_  | \new_[6160]_ ;
  assign \new_[6167]_  = \new_[6166]_  | \new_[6155]_ ;
  assign \new_[6171]_  = \new_[1673]_  | \new_[1674]_ ;
  assign \new_[6172]_  = \new_[1675]_  | \new_[6171]_ ;
  assign \new_[6176]_  = \new_[1670]_  | \new_[1671]_ ;
  assign \new_[6177]_  = \new_[1672]_  | \new_[6176]_ ;
  assign \new_[6178]_  = \new_[6177]_  | \new_[6172]_ ;
  assign \new_[6182]_  = \new_[1667]_  | \new_[1668]_ ;
  assign \new_[6183]_  = \new_[1669]_  | \new_[6182]_ ;
  assign \new_[6186]_  = \new_[1665]_  | \new_[1666]_ ;
  assign \new_[6189]_  = \new_[1663]_  | \new_[1664]_ ;
  assign \new_[6190]_  = \new_[6189]_  | \new_[6186]_ ;
  assign \new_[6191]_  = \new_[6190]_  | \new_[6183]_ ;
  assign \new_[6192]_  = \new_[6191]_  | \new_[6178]_ ;
  assign \new_[6193]_  = \new_[6192]_  | \new_[6167]_ ;
  assign \new_[6197]_  = \new_[1660]_  | \new_[1661]_ ;
  assign \new_[6198]_  = \new_[1662]_  | \new_[6197]_ ;
  assign \new_[6202]_  = \new_[1657]_  | \new_[1658]_ ;
  assign \new_[6203]_  = \new_[1659]_  | \new_[6202]_ ;
  assign \new_[6204]_  = \new_[6203]_  | \new_[6198]_ ;
  assign \new_[6208]_  = \new_[1654]_  | \new_[1655]_ ;
  assign \new_[6209]_  = \new_[1656]_  | \new_[6208]_ ;
  assign \new_[6213]_  = \new_[1651]_  | \new_[1652]_ ;
  assign \new_[6214]_  = \new_[1653]_  | \new_[6213]_ ;
  assign \new_[6215]_  = \new_[6214]_  | \new_[6209]_ ;
  assign \new_[6216]_  = \new_[6215]_  | \new_[6204]_ ;
  assign \new_[6220]_  = \new_[1648]_  | \new_[1649]_ ;
  assign \new_[6221]_  = \new_[1650]_  | \new_[6220]_ ;
  assign \new_[6225]_  = \new_[1645]_  | \new_[1646]_ ;
  assign \new_[6226]_  = \new_[1647]_  | \new_[6225]_ ;
  assign \new_[6227]_  = \new_[6226]_  | \new_[6221]_ ;
  assign \new_[6231]_  = \new_[1642]_  | \new_[1643]_ ;
  assign \new_[6232]_  = \new_[1644]_  | \new_[6231]_ ;
  assign \new_[6235]_  = \new_[1640]_  | \new_[1641]_ ;
  assign \new_[6238]_  = \new_[1638]_  | \new_[1639]_ ;
  assign \new_[6239]_  = \new_[6238]_  | \new_[6235]_ ;
  assign \new_[6240]_  = \new_[6239]_  | \new_[6232]_ ;
  assign \new_[6241]_  = \new_[6240]_  | \new_[6227]_ ;
  assign \new_[6242]_  = \new_[6241]_  | \new_[6216]_ ;
  assign \new_[6243]_  = \new_[6242]_  | \new_[6193]_ ;
  assign \new_[6247]_  = \new_[1635]_  | \new_[1636]_ ;
  assign \new_[6248]_  = \new_[1637]_  | \new_[6247]_ ;
  assign \new_[6252]_  = \new_[1632]_  | \new_[1633]_ ;
  assign \new_[6253]_  = \new_[1634]_  | \new_[6252]_ ;
  assign \new_[6254]_  = \new_[6253]_  | \new_[6248]_ ;
  assign \new_[6258]_  = \new_[1629]_  | \new_[1630]_ ;
  assign \new_[6259]_  = \new_[1631]_  | \new_[6258]_ ;
  assign \new_[6263]_  = \new_[1626]_  | \new_[1627]_ ;
  assign \new_[6264]_  = \new_[1628]_  | \new_[6263]_ ;
  assign \new_[6265]_  = \new_[6264]_  | \new_[6259]_ ;
  assign \new_[6266]_  = \new_[6265]_  | \new_[6254]_ ;
  assign \new_[6270]_  = \new_[1623]_  | \new_[1624]_ ;
  assign \new_[6271]_  = \new_[1625]_  | \new_[6270]_ ;
  assign \new_[6275]_  = \new_[1620]_  | \new_[1621]_ ;
  assign \new_[6276]_  = \new_[1622]_  | \new_[6275]_ ;
  assign \new_[6277]_  = \new_[6276]_  | \new_[6271]_ ;
  assign \new_[6281]_  = \new_[1617]_  | \new_[1618]_ ;
  assign \new_[6282]_  = \new_[1619]_  | \new_[6281]_ ;
  assign \new_[6285]_  = \new_[1615]_  | \new_[1616]_ ;
  assign \new_[6288]_  = \new_[1613]_  | \new_[1614]_ ;
  assign \new_[6289]_  = \new_[6288]_  | \new_[6285]_ ;
  assign \new_[6290]_  = \new_[6289]_  | \new_[6282]_ ;
  assign \new_[6291]_  = \new_[6290]_  | \new_[6277]_ ;
  assign \new_[6292]_  = \new_[6291]_  | \new_[6266]_ ;
  assign \new_[6296]_  = \new_[1610]_  | \new_[1611]_ ;
  assign \new_[6297]_  = \new_[1612]_  | \new_[6296]_ ;
  assign \new_[6301]_  = \new_[1607]_  | \new_[1608]_ ;
  assign \new_[6302]_  = \new_[1609]_  | \new_[6301]_ ;
  assign \new_[6303]_  = \new_[6302]_  | \new_[6297]_ ;
  assign \new_[6307]_  = \new_[1604]_  | \new_[1605]_ ;
  assign \new_[6308]_  = \new_[1606]_  | \new_[6307]_ ;
  assign \new_[6312]_  = \new_[1601]_  | \new_[1602]_ ;
  assign \new_[6313]_  = \new_[1603]_  | \new_[6312]_ ;
  assign \new_[6314]_  = \new_[6313]_  | \new_[6308]_ ;
  assign \new_[6315]_  = \new_[6314]_  | \new_[6303]_ ;
  assign \new_[6319]_  = \new_[1598]_  | \new_[1599]_ ;
  assign \new_[6320]_  = \new_[1600]_  | \new_[6319]_ ;
  assign \new_[6324]_  = \new_[1595]_  | \new_[1596]_ ;
  assign \new_[6325]_  = \new_[1597]_  | \new_[6324]_ ;
  assign \new_[6326]_  = \new_[6325]_  | \new_[6320]_ ;
  assign \new_[6330]_  = \new_[1592]_  | \new_[1593]_ ;
  assign \new_[6331]_  = \new_[1594]_  | \new_[6330]_ ;
  assign \new_[6334]_  = \new_[1590]_  | \new_[1591]_ ;
  assign \new_[6337]_  = \new_[1588]_  | \new_[1589]_ ;
  assign \new_[6338]_  = \new_[6337]_  | \new_[6334]_ ;
  assign \new_[6339]_  = \new_[6338]_  | \new_[6331]_ ;
  assign \new_[6340]_  = \new_[6339]_  | \new_[6326]_ ;
  assign \new_[6341]_  = \new_[6340]_  | \new_[6315]_ ;
  assign \new_[6342]_  = \new_[6341]_  | \new_[6292]_ ;
  assign \new_[6343]_  = \new_[6342]_  | \new_[6243]_ ;
  assign \new_[6344]_  = \new_[6343]_  | \new_[6144]_ ;
  assign \new_[6345]_  = \new_[6344]_  | \new_[5947]_ ;
  assign \new_[6346]_  = \new_[6345]_  | \new_[5552]_ ;
  assign \new_[6347]_  = \new_[6346]_  | \new_[4759]_ ;
  assign \new_[6351]_  = \new_[1585]_  | \new_[1586]_ ;
  assign \new_[6352]_  = \new_[1587]_  | \new_[6351]_ ;
  assign \new_[6356]_  = \new_[1582]_  | \new_[1583]_ ;
  assign \new_[6357]_  = \new_[1584]_  | \new_[6356]_ ;
  assign \new_[6358]_  = \new_[6357]_  | \new_[6352]_ ;
  assign \new_[6362]_  = \new_[1579]_  | \new_[1580]_ ;
  assign \new_[6363]_  = \new_[1581]_  | \new_[6362]_ ;
  assign \new_[6367]_  = \new_[1576]_  | \new_[1577]_ ;
  assign \new_[6368]_  = \new_[1578]_  | \new_[6367]_ ;
  assign \new_[6369]_  = \new_[6368]_  | \new_[6363]_ ;
  assign \new_[6370]_  = \new_[6369]_  | \new_[6358]_ ;
  assign \new_[6374]_  = \new_[1573]_  | \new_[1574]_ ;
  assign \new_[6375]_  = \new_[1575]_  | \new_[6374]_ ;
  assign \new_[6379]_  = \new_[1570]_  | \new_[1571]_ ;
  assign \new_[6380]_  = \new_[1572]_  | \new_[6379]_ ;
  assign \new_[6381]_  = \new_[6380]_  | \new_[6375]_ ;
  assign \new_[6385]_  = \new_[1567]_  | \new_[1568]_ ;
  assign \new_[6386]_  = \new_[1569]_  | \new_[6385]_ ;
  assign \new_[6390]_  = \new_[1564]_  | \new_[1565]_ ;
  assign \new_[6391]_  = \new_[1566]_  | \new_[6390]_ ;
  assign \new_[6392]_  = \new_[6391]_  | \new_[6386]_ ;
  assign \new_[6393]_  = \new_[6392]_  | \new_[6381]_ ;
  assign \new_[6394]_  = \new_[6393]_  | \new_[6370]_ ;
  assign \new_[6398]_  = \new_[1561]_  | \new_[1562]_ ;
  assign \new_[6399]_  = \new_[1563]_  | \new_[6398]_ ;
  assign \new_[6403]_  = \new_[1558]_  | \new_[1559]_ ;
  assign \new_[6404]_  = \new_[1560]_  | \new_[6403]_ ;
  assign \new_[6405]_  = \new_[6404]_  | \new_[6399]_ ;
  assign \new_[6409]_  = \new_[1555]_  | \new_[1556]_ ;
  assign \new_[6410]_  = \new_[1557]_  | \new_[6409]_ ;
  assign \new_[6414]_  = \new_[1552]_  | \new_[1553]_ ;
  assign \new_[6415]_  = \new_[1554]_  | \new_[6414]_ ;
  assign \new_[6416]_  = \new_[6415]_  | \new_[6410]_ ;
  assign \new_[6417]_  = \new_[6416]_  | \new_[6405]_ ;
  assign \new_[6421]_  = \new_[1549]_  | \new_[1550]_ ;
  assign \new_[6422]_  = \new_[1551]_  | \new_[6421]_ ;
  assign \new_[6426]_  = \new_[1546]_  | \new_[1547]_ ;
  assign \new_[6427]_  = \new_[1548]_  | \new_[6426]_ ;
  assign \new_[6428]_  = \new_[6427]_  | \new_[6422]_ ;
  assign \new_[6432]_  = \new_[1543]_  | \new_[1544]_ ;
  assign \new_[6433]_  = \new_[1545]_  | \new_[6432]_ ;
  assign \new_[6436]_  = \new_[1541]_  | \new_[1542]_ ;
  assign \new_[6439]_  = \new_[1539]_  | \new_[1540]_ ;
  assign \new_[6440]_  = \new_[6439]_  | \new_[6436]_ ;
  assign \new_[6441]_  = \new_[6440]_  | \new_[6433]_ ;
  assign \new_[6442]_  = \new_[6441]_  | \new_[6428]_ ;
  assign \new_[6443]_  = \new_[6442]_  | \new_[6417]_ ;
  assign \new_[6444]_  = \new_[6443]_  | \new_[6394]_ ;
  assign \new_[6448]_  = \new_[1536]_  | \new_[1537]_ ;
  assign \new_[6449]_  = \new_[1538]_  | \new_[6448]_ ;
  assign \new_[6453]_  = \new_[1533]_  | \new_[1534]_ ;
  assign \new_[6454]_  = \new_[1535]_  | \new_[6453]_ ;
  assign \new_[6455]_  = \new_[6454]_  | \new_[6449]_ ;
  assign \new_[6459]_  = \new_[1530]_  | \new_[1531]_ ;
  assign \new_[6460]_  = \new_[1532]_  | \new_[6459]_ ;
  assign \new_[6464]_  = \new_[1527]_  | \new_[1528]_ ;
  assign \new_[6465]_  = \new_[1529]_  | \new_[6464]_ ;
  assign \new_[6466]_  = \new_[6465]_  | \new_[6460]_ ;
  assign \new_[6467]_  = \new_[6466]_  | \new_[6455]_ ;
  assign \new_[6471]_  = \new_[1524]_  | \new_[1525]_ ;
  assign \new_[6472]_  = \new_[1526]_  | \new_[6471]_ ;
  assign \new_[6476]_  = \new_[1521]_  | \new_[1522]_ ;
  assign \new_[6477]_  = \new_[1523]_  | \new_[6476]_ ;
  assign \new_[6478]_  = \new_[6477]_  | \new_[6472]_ ;
  assign \new_[6482]_  = \new_[1518]_  | \new_[1519]_ ;
  assign \new_[6483]_  = \new_[1520]_  | \new_[6482]_ ;
  assign \new_[6486]_  = \new_[1516]_  | \new_[1517]_ ;
  assign \new_[6489]_  = \new_[1514]_  | \new_[1515]_ ;
  assign \new_[6490]_  = \new_[6489]_  | \new_[6486]_ ;
  assign \new_[6491]_  = \new_[6490]_  | \new_[6483]_ ;
  assign \new_[6492]_  = \new_[6491]_  | \new_[6478]_ ;
  assign \new_[6493]_  = \new_[6492]_  | \new_[6467]_ ;
  assign \new_[6497]_  = \new_[1511]_  | \new_[1512]_ ;
  assign \new_[6498]_  = \new_[1513]_  | \new_[6497]_ ;
  assign \new_[6502]_  = \new_[1508]_  | \new_[1509]_ ;
  assign \new_[6503]_  = \new_[1510]_  | \new_[6502]_ ;
  assign \new_[6504]_  = \new_[6503]_  | \new_[6498]_ ;
  assign \new_[6508]_  = \new_[1505]_  | \new_[1506]_ ;
  assign \new_[6509]_  = \new_[1507]_  | \new_[6508]_ ;
  assign \new_[6513]_  = \new_[1502]_  | \new_[1503]_ ;
  assign \new_[6514]_  = \new_[1504]_  | \new_[6513]_ ;
  assign \new_[6515]_  = \new_[6514]_  | \new_[6509]_ ;
  assign \new_[6516]_  = \new_[6515]_  | \new_[6504]_ ;
  assign \new_[6520]_  = \new_[1499]_  | \new_[1500]_ ;
  assign \new_[6521]_  = \new_[1501]_  | \new_[6520]_ ;
  assign \new_[6525]_  = \new_[1496]_  | \new_[1497]_ ;
  assign \new_[6526]_  = \new_[1498]_  | \new_[6525]_ ;
  assign \new_[6527]_  = \new_[6526]_  | \new_[6521]_ ;
  assign \new_[6531]_  = \new_[1493]_  | \new_[1494]_ ;
  assign \new_[6532]_  = \new_[1495]_  | \new_[6531]_ ;
  assign \new_[6535]_  = \new_[1491]_  | \new_[1492]_ ;
  assign \new_[6538]_  = \new_[1489]_  | \new_[1490]_ ;
  assign \new_[6539]_  = \new_[6538]_  | \new_[6535]_ ;
  assign \new_[6540]_  = \new_[6539]_  | \new_[6532]_ ;
  assign \new_[6541]_  = \new_[6540]_  | \new_[6527]_ ;
  assign \new_[6542]_  = \new_[6541]_  | \new_[6516]_ ;
  assign \new_[6543]_  = \new_[6542]_  | \new_[6493]_ ;
  assign \new_[6544]_  = \new_[6543]_  | \new_[6444]_ ;
  assign \new_[6548]_  = \new_[1486]_  | \new_[1487]_ ;
  assign \new_[6549]_  = \new_[1488]_  | \new_[6548]_ ;
  assign \new_[6553]_  = \new_[1483]_  | \new_[1484]_ ;
  assign \new_[6554]_  = \new_[1485]_  | \new_[6553]_ ;
  assign \new_[6555]_  = \new_[6554]_  | \new_[6549]_ ;
  assign \new_[6559]_  = \new_[1480]_  | \new_[1481]_ ;
  assign \new_[6560]_  = \new_[1482]_  | \new_[6559]_ ;
  assign \new_[6564]_  = \new_[1477]_  | \new_[1478]_ ;
  assign \new_[6565]_  = \new_[1479]_  | \new_[6564]_ ;
  assign \new_[6566]_  = \new_[6565]_  | \new_[6560]_ ;
  assign \new_[6567]_  = \new_[6566]_  | \new_[6555]_ ;
  assign \new_[6571]_  = \new_[1474]_  | \new_[1475]_ ;
  assign \new_[6572]_  = \new_[1476]_  | \new_[6571]_ ;
  assign \new_[6576]_  = \new_[1471]_  | \new_[1472]_ ;
  assign \new_[6577]_  = \new_[1473]_  | \new_[6576]_ ;
  assign \new_[6578]_  = \new_[6577]_  | \new_[6572]_ ;
  assign \new_[6582]_  = \new_[1468]_  | \new_[1469]_ ;
  assign \new_[6583]_  = \new_[1470]_  | \new_[6582]_ ;
  assign \new_[6587]_  = \new_[1465]_  | \new_[1466]_ ;
  assign \new_[6588]_  = \new_[1467]_  | \new_[6587]_ ;
  assign \new_[6589]_  = \new_[6588]_  | \new_[6583]_ ;
  assign \new_[6590]_  = \new_[6589]_  | \new_[6578]_ ;
  assign \new_[6591]_  = \new_[6590]_  | \new_[6567]_ ;
  assign \new_[6595]_  = \new_[1462]_  | \new_[1463]_ ;
  assign \new_[6596]_  = \new_[1464]_  | \new_[6595]_ ;
  assign \new_[6600]_  = \new_[1459]_  | \new_[1460]_ ;
  assign \new_[6601]_  = \new_[1461]_  | \new_[6600]_ ;
  assign \new_[6602]_  = \new_[6601]_  | \new_[6596]_ ;
  assign \new_[6606]_  = \new_[1456]_  | \new_[1457]_ ;
  assign \new_[6607]_  = \new_[1458]_  | \new_[6606]_ ;
  assign \new_[6611]_  = \new_[1453]_  | \new_[1454]_ ;
  assign \new_[6612]_  = \new_[1455]_  | \new_[6611]_ ;
  assign \new_[6613]_  = \new_[6612]_  | \new_[6607]_ ;
  assign \new_[6614]_  = \new_[6613]_  | \new_[6602]_ ;
  assign \new_[6618]_  = \new_[1450]_  | \new_[1451]_ ;
  assign \new_[6619]_  = \new_[1452]_  | \new_[6618]_ ;
  assign \new_[6623]_  = \new_[1447]_  | \new_[1448]_ ;
  assign \new_[6624]_  = \new_[1449]_  | \new_[6623]_ ;
  assign \new_[6625]_  = \new_[6624]_  | \new_[6619]_ ;
  assign \new_[6629]_  = \new_[1444]_  | \new_[1445]_ ;
  assign \new_[6630]_  = \new_[1446]_  | \new_[6629]_ ;
  assign \new_[6633]_  = \new_[1442]_  | \new_[1443]_ ;
  assign \new_[6636]_  = \new_[1440]_  | \new_[1441]_ ;
  assign \new_[6637]_  = \new_[6636]_  | \new_[6633]_ ;
  assign \new_[6638]_  = \new_[6637]_  | \new_[6630]_ ;
  assign \new_[6639]_  = \new_[6638]_  | \new_[6625]_ ;
  assign \new_[6640]_  = \new_[6639]_  | \new_[6614]_ ;
  assign \new_[6641]_  = \new_[6640]_  | \new_[6591]_ ;
  assign \new_[6645]_  = \new_[1437]_  | \new_[1438]_ ;
  assign \new_[6646]_  = \new_[1439]_  | \new_[6645]_ ;
  assign \new_[6650]_  = \new_[1434]_  | \new_[1435]_ ;
  assign \new_[6651]_  = \new_[1436]_  | \new_[6650]_ ;
  assign \new_[6652]_  = \new_[6651]_  | \new_[6646]_ ;
  assign \new_[6656]_  = \new_[1431]_  | \new_[1432]_ ;
  assign \new_[6657]_  = \new_[1433]_  | \new_[6656]_ ;
  assign \new_[6661]_  = \new_[1428]_  | \new_[1429]_ ;
  assign \new_[6662]_  = \new_[1430]_  | \new_[6661]_ ;
  assign \new_[6663]_  = \new_[6662]_  | \new_[6657]_ ;
  assign \new_[6664]_  = \new_[6663]_  | \new_[6652]_ ;
  assign \new_[6668]_  = \new_[1425]_  | \new_[1426]_ ;
  assign \new_[6669]_  = \new_[1427]_  | \new_[6668]_ ;
  assign \new_[6673]_  = \new_[1422]_  | \new_[1423]_ ;
  assign \new_[6674]_  = \new_[1424]_  | \new_[6673]_ ;
  assign \new_[6675]_  = \new_[6674]_  | \new_[6669]_ ;
  assign \new_[6679]_  = \new_[1419]_  | \new_[1420]_ ;
  assign \new_[6680]_  = \new_[1421]_  | \new_[6679]_ ;
  assign \new_[6683]_  = \new_[1417]_  | \new_[1418]_ ;
  assign \new_[6686]_  = \new_[1415]_  | \new_[1416]_ ;
  assign \new_[6687]_  = \new_[6686]_  | \new_[6683]_ ;
  assign \new_[6688]_  = \new_[6687]_  | \new_[6680]_ ;
  assign \new_[6689]_  = \new_[6688]_  | \new_[6675]_ ;
  assign \new_[6690]_  = \new_[6689]_  | \new_[6664]_ ;
  assign \new_[6694]_  = \new_[1412]_  | \new_[1413]_ ;
  assign \new_[6695]_  = \new_[1414]_  | \new_[6694]_ ;
  assign \new_[6699]_  = \new_[1409]_  | \new_[1410]_ ;
  assign \new_[6700]_  = \new_[1411]_  | \new_[6699]_ ;
  assign \new_[6701]_  = \new_[6700]_  | \new_[6695]_ ;
  assign \new_[6705]_  = \new_[1406]_  | \new_[1407]_ ;
  assign \new_[6706]_  = \new_[1408]_  | \new_[6705]_ ;
  assign \new_[6710]_  = \new_[1403]_  | \new_[1404]_ ;
  assign \new_[6711]_  = \new_[1405]_  | \new_[6710]_ ;
  assign \new_[6712]_  = \new_[6711]_  | \new_[6706]_ ;
  assign \new_[6713]_  = \new_[6712]_  | \new_[6701]_ ;
  assign \new_[6717]_  = \new_[1400]_  | \new_[1401]_ ;
  assign \new_[6718]_  = \new_[1402]_  | \new_[6717]_ ;
  assign \new_[6722]_  = \new_[1397]_  | \new_[1398]_ ;
  assign \new_[6723]_  = \new_[1399]_  | \new_[6722]_ ;
  assign \new_[6724]_  = \new_[6723]_  | \new_[6718]_ ;
  assign \new_[6728]_  = \new_[1394]_  | \new_[1395]_ ;
  assign \new_[6729]_  = \new_[1396]_  | \new_[6728]_ ;
  assign \new_[6732]_  = \new_[1392]_  | \new_[1393]_ ;
  assign \new_[6735]_  = \new_[1390]_  | \new_[1391]_ ;
  assign \new_[6736]_  = \new_[6735]_  | \new_[6732]_ ;
  assign \new_[6737]_  = \new_[6736]_  | \new_[6729]_ ;
  assign \new_[6738]_  = \new_[6737]_  | \new_[6724]_ ;
  assign \new_[6739]_  = \new_[6738]_  | \new_[6713]_ ;
  assign \new_[6740]_  = \new_[6739]_  | \new_[6690]_ ;
  assign \new_[6741]_  = \new_[6740]_  | \new_[6641]_ ;
  assign \new_[6742]_  = \new_[6741]_  | \new_[6544]_ ;
  assign \new_[6746]_  = \new_[1387]_  | \new_[1388]_ ;
  assign \new_[6747]_  = \new_[1389]_  | \new_[6746]_ ;
  assign \new_[6751]_  = \new_[1384]_  | \new_[1385]_ ;
  assign \new_[6752]_  = \new_[1386]_  | \new_[6751]_ ;
  assign \new_[6753]_  = \new_[6752]_  | \new_[6747]_ ;
  assign \new_[6757]_  = \new_[1381]_  | \new_[1382]_ ;
  assign \new_[6758]_  = \new_[1383]_  | \new_[6757]_ ;
  assign \new_[6762]_  = \new_[1378]_  | \new_[1379]_ ;
  assign \new_[6763]_  = \new_[1380]_  | \new_[6762]_ ;
  assign \new_[6764]_  = \new_[6763]_  | \new_[6758]_ ;
  assign \new_[6765]_  = \new_[6764]_  | \new_[6753]_ ;
  assign \new_[6769]_  = \new_[1375]_  | \new_[1376]_ ;
  assign \new_[6770]_  = \new_[1377]_  | \new_[6769]_ ;
  assign \new_[6774]_  = \new_[1372]_  | \new_[1373]_ ;
  assign \new_[6775]_  = \new_[1374]_  | \new_[6774]_ ;
  assign \new_[6776]_  = \new_[6775]_  | \new_[6770]_ ;
  assign \new_[6780]_  = \new_[1369]_  | \new_[1370]_ ;
  assign \new_[6781]_  = \new_[1371]_  | \new_[6780]_ ;
  assign \new_[6785]_  = \new_[1366]_  | \new_[1367]_ ;
  assign \new_[6786]_  = \new_[1368]_  | \new_[6785]_ ;
  assign \new_[6787]_  = \new_[6786]_  | \new_[6781]_ ;
  assign \new_[6788]_  = \new_[6787]_  | \new_[6776]_ ;
  assign \new_[6789]_  = \new_[6788]_  | \new_[6765]_ ;
  assign \new_[6793]_  = \new_[1363]_  | \new_[1364]_ ;
  assign \new_[6794]_  = \new_[1365]_  | \new_[6793]_ ;
  assign \new_[6798]_  = \new_[1360]_  | \new_[1361]_ ;
  assign \new_[6799]_  = \new_[1362]_  | \new_[6798]_ ;
  assign \new_[6800]_  = \new_[6799]_  | \new_[6794]_ ;
  assign \new_[6804]_  = \new_[1357]_  | \new_[1358]_ ;
  assign \new_[6805]_  = \new_[1359]_  | \new_[6804]_ ;
  assign \new_[6809]_  = \new_[1354]_  | \new_[1355]_ ;
  assign \new_[6810]_  = \new_[1356]_  | \new_[6809]_ ;
  assign \new_[6811]_  = \new_[6810]_  | \new_[6805]_ ;
  assign \new_[6812]_  = \new_[6811]_  | \new_[6800]_ ;
  assign \new_[6816]_  = \new_[1351]_  | \new_[1352]_ ;
  assign \new_[6817]_  = \new_[1353]_  | \new_[6816]_ ;
  assign \new_[6821]_  = \new_[1348]_  | \new_[1349]_ ;
  assign \new_[6822]_  = \new_[1350]_  | \new_[6821]_ ;
  assign \new_[6823]_  = \new_[6822]_  | \new_[6817]_ ;
  assign \new_[6827]_  = \new_[1345]_  | \new_[1346]_ ;
  assign \new_[6828]_  = \new_[1347]_  | \new_[6827]_ ;
  assign \new_[6831]_  = \new_[1343]_  | \new_[1344]_ ;
  assign \new_[6834]_  = \new_[1341]_  | \new_[1342]_ ;
  assign \new_[6835]_  = \new_[6834]_  | \new_[6831]_ ;
  assign \new_[6836]_  = \new_[6835]_  | \new_[6828]_ ;
  assign \new_[6837]_  = \new_[6836]_  | \new_[6823]_ ;
  assign \new_[6838]_  = \new_[6837]_  | \new_[6812]_ ;
  assign \new_[6839]_  = \new_[6838]_  | \new_[6789]_ ;
  assign \new_[6843]_  = \new_[1338]_  | \new_[1339]_ ;
  assign \new_[6844]_  = \new_[1340]_  | \new_[6843]_ ;
  assign \new_[6848]_  = \new_[1335]_  | \new_[1336]_ ;
  assign \new_[6849]_  = \new_[1337]_  | \new_[6848]_ ;
  assign \new_[6850]_  = \new_[6849]_  | \new_[6844]_ ;
  assign \new_[6854]_  = \new_[1332]_  | \new_[1333]_ ;
  assign \new_[6855]_  = \new_[1334]_  | \new_[6854]_ ;
  assign \new_[6859]_  = \new_[1329]_  | \new_[1330]_ ;
  assign \new_[6860]_  = \new_[1331]_  | \new_[6859]_ ;
  assign \new_[6861]_  = \new_[6860]_  | \new_[6855]_ ;
  assign \new_[6862]_  = \new_[6861]_  | \new_[6850]_ ;
  assign \new_[6866]_  = \new_[1326]_  | \new_[1327]_ ;
  assign \new_[6867]_  = \new_[1328]_  | \new_[6866]_ ;
  assign \new_[6871]_  = \new_[1323]_  | \new_[1324]_ ;
  assign \new_[6872]_  = \new_[1325]_  | \new_[6871]_ ;
  assign \new_[6873]_  = \new_[6872]_  | \new_[6867]_ ;
  assign \new_[6877]_  = \new_[1320]_  | \new_[1321]_ ;
  assign \new_[6878]_  = \new_[1322]_  | \new_[6877]_ ;
  assign \new_[6881]_  = \new_[1318]_  | \new_[1319]_ ;
  assign \new_[6884]_  = \new_[1316]_  | \new_[1317]_ ;
  assign \new_[6885]_  = \new_[6884]_  | \new_[6881]_ ;
  assign \new_[6886]_  = \new_[6885]_  | \new_[6878]_ ;
  assign \new_[6887]_  = \new_[6886]_  | \new_[6873]_ ;
  assign \new_[6888]_  = \new_[6887]_  | \new_[6862]_ ;
  assign \new_[6892]_  = \new_[1313]_  | \new_[1314]_ ;
  assign \new_[6893]_  = \new_[1315]_  | \new_[6892]_ ;
  assign \new_[6897]_  = \new_[1310]_  | \new_[1311]_ ;
  assign \new_[6898]_  = \new_[1312]_  | \new_[6897]_ ;
  assign \new_[6899]_  = \new_[6898]_  | \new_[6893]_ ;
  assign \new_[6903]_  = \new_[1307]_  | \new_[1308]_ ;
  assign \new_[6904]_  = \new_[1309]_  | \new_[6903]_ ;
  assign \new_[6908]_  = \new_[1304]_  | \new_[1305]_ ;
  assign \new_[6909]_  = \new_[1306]_  | \new_[6908]_ ;
  assign \new_[6910]_  = \new_[6909]_  | \new_[6904]_ ;
  assign \new_[6911]_  = \new_[6910]_  | \new_[6899]_ ;
  assign \new_[6915]_  = \new_[1301]_  | \new_[1302]_ ;
  assign \new_[6916]_  = \new_[1303]_  | \new_[6915]_ ;
  assign \new_[6920]_  = \new_[1298]_  | \new_[1299]_ ;
  assign \new_[6921]_  = \new_[1300]_  | \new_[6920]_ ;
  assign \new_[6922]_  = \new_[6921]_  | \new_[6916]_ ;
  assign \new_[6926]_  = \new_[1295]_  | \new_[1296]_ ;
  assign \new_[6927]_  = \new_[1297]_  | \new_[6926]_ ;
  assign \new_[6930]_  = \new_[1293]_  | \new_[1294]_ ;
  assign \new_[6933]_  = \new_[1291]_  | \new_[1292]_ ;
  assign \new_[6934]_  = \new_[6933]_  | \new_[6930]_ ;
  assign \new_[6935]_  = \new_[6934]_  | \new_[6927]_ ;
  assign \new_[6936]_  = \new_[6935]_  | \new_[6922]_ ;
  assign \new_[6937]_  = \new_[6936]_  | \new_[6911]_ ;
  assign \new_[6938]_  = \new_[6937]_  | \new_[6888]_ ;
  assign \new_[6939]_  = \new_[6938]_  | \new_[6839]_ ;
  assign \new_[6943]_  = \new_[1288]_  | \new_[1289]_ ;
  assign \new_[6944]_  = \new_[1290]_  | \new_[6943]_ ;
  assign \new_[6948]_  = \new_[1285]_  | \new_[1286]_ ;
  assign \new_[6949]_  = \new_[1287]_  | \new_[6948]_ ;
  assign \new_[6950]_  = \new_[6949]_  | \new_[6944]_ ;
  assign \new_[6954]_  = \new_[1282]_  | \new_[1283]_ ;
  assign \new_[6955]_  = \new_[1284]_  | \new_[6954]_ ;
  assign \new_[6959]_  = \new_[1279]_  | \new_[1280]_ ;
  assign \new_[6960]_  = \new_[1281]_  | \new_[6959]_ ;
  assign \new_[6961]_  = \new_[6960]_  | \new_[6955]_ ;
  assign \new_[6962]_  = \new_[6961]_  | \new_[6950]_ ;
  assign \new_[6966]_  = \new_[1276]_  | \new_[1277]_ ;
  assign \new_[6967]_  = \new_[1278]_  | \new_[6966]_ ;
  assign \new_[6971]_  = \new_[1273]_  | \new_[1274]_ ;
  assign \new_[6972]_  = \new_[1275]_  | \new_[6971]_ ;
  assign \new_[6973]_  = \new_[6972]_  | \new_[6967]_ ;
  assign \new_[6977]_  = \new_[1270]_  | \new_[1271]_ ;
  assign \new_[6978]_  = \new_[1272]_  | \new_[6977]_ ;
  assign \new_[6982]_  = \new_[1267]_  | \new_[1268]_ ;
  assign \new_[6983]_  = \new_[1269]_  | \new_[6982]_ ;
  assign \new_[6984]_  = \new_[6983]_  | \new_[6978]_ ;
  assign \new_[6985]_  = \new_[6984]_  | \new_[6973]_ ;
  assign \new_[6986]_  = \new_[6985]_  | \new_[6962]_ ;
  assign \new_[6990]_  = \new_[1264]_  | \new_[1265]_ ;
  assign \new_[6991]_  = \new_[1266]_  | \new_[6990]_ ;
  assign \new_[6995]_  = \new_[1261]_  | \new_[1262]_ ;
  assign \new_[6996]_  = \new_[1263]_  | \new_[6995]_ ;
  assign \new_[6997]_  = \new_[6996]_  | \new_[6991]_ ;
  assign \new_[7001]_  = \new_[1258]_  | \new_[1259]_ ;
  assign \new_[7002]_  = \new_[1260]_  | \new_[7001]_ ;
  assign \new_[7006]_  = \new_[1255]_  | \new_[1256]_ ;
  assign \new_[7007]_  = \new_[1257]_  | \new_[7006]_ ;
  assign \new_[7008]_  = \new_[7007]_  | \new_[7002]_ ;
  assign \new_[7009]_  = \new_[7008]_  | \new_[6997]_ ;
  assign \new_[7013]_  = \new_[1252]_  | \new_[1253]_ ;
  assign \new_[7014]_  = \new_[1254]_  | \new_[7013]_ ;
  assign \new_[7018]_  = \new_[1249]_  | \new_[1250]_ ;
  assign \new_[7019]_  = \new_[1251]_  | \new_[7018]_ ;
  assign \new_[7020]_  = \new_[7019]_  | \new_[7014]_ ;
  assign \new_[7024]_  = \new_[1246]_  | \new_[1247]_ ;
  assign \new_[7025]_  = \new_[1248]_  | \new_[7024]_ ;
  assign \new_[7028]_  = \new_[1244]_  | \new_[1245]_ ;
  assign \new_[7031]_  = \new_[1242]_  | \new_[1243]_ ;
  assign \new_[7032]_  = \new_[7031]_  | \new_[7028]_ ;
  assign \new_[7033]_  = \new_[7032]_  | \new_[7025]_ ;
  assign \new_[7034]_  = \new_[7033]_  | \new_[7020]_ ;
  assign \new_[7035]_  = \new_[7034]_  | \new_[7009]_ ;
  assign \new_[7036]_  = \new_[7035]_  | \new_[6986]_ ;
  assign \new_[7040]_  = \new_[1239]_  | \new_[1240]_ ;
  assign \new_[7041]_  = \new_[1241]_  | \new_[7040]_ ;
  assign \new_[7045]_  = \new_[1236]_  | \new_[1237]_ ;
  assign \new_[7046]_  = \new_[1238]_  | \new_[7045]_ ;
  assign \new_[7047]_  = \new_[7046]_  | \new_[7041]_ ;
  assign \new_[7051]_  = \new_[1233]_  | \new_[1234]_ ;
  assign \new_[7052]_  = \new_[1235]_  | \new_[7051]_ ;
  assign \new_[7056]_  = \new_[1230]_  | \new_[1231]_ ;
  assign \new_[7057]_  = \new_[1232]_  | \new_[7056]_ ;
  assign \new_[7058]_  = \new_[7057]_  | \new_[7052]_ ;
  assign \new_[7059]_  = \new_[7058]_  | \new_[7047]_ ;
  assign \new_[7063]_  = \new_[1227]_  | \new_[1228]_ ;
  assign \new_[7064]_  = \new_[1229]_  | \new_[7063]_ ;
  assign \new_[7068]_  = \new_[1224]_  | \new_[1225]_ ;
  assign \new_[7069]_  = \new_[1226]_  | \new_[7068]_ ;
  assign \new_[7070]_  = \new_[7069]_  | \new_[7064]_ ;
  assign \new_[7074]_  = \new_[1221]_  | \new_[1222]_ ;
  assign \new_[7075]_  = \new_[1223]_  | \new_[7074]_ ;
  assign \new_[7078]_  = \new_[1219]_  | \new_[1220]_ ;
  assign \new_[7081]_  = \new_[1217]_  | \new_[1218]_ ;
  assign \new_[7082]_  = \new_[7081]_  | \new_[7078]_ ;
  assign \new_[7083]_  = \new_[7082]_  | \new_[7075]_ ;
  assign \new_[7084]_  = \new_[7083]_  | \new_[7070]_ ;
  assign \new_[7085]_  = \new_[7084]_  | \new_[7059]_ ;
  assign \new_[7089]_  = \new_[1214]_  | \new_[1215]_ ;
  assign \new_[7090]_  = \new_[1216]_  | \new_[7089]_ ;
  assign \new_[7094]_  = \new_[1211]_  | \new_[1212]_ ;
  assign \new_[7095]_  = \new_[1213]_  | \new_[7094]_ ;
  assign \new_[7096]_  = \new_[7095]_  | \new_[7090]_ ;
  assign \new_[7100]_  = \new_[1208]_  | \new_[1209]_ ;
  assign \new_[7101]_  = \new_[1210]_  | \new_[7100]_ ;
  assign \new_[7105]_  = \new_[1205]_  | \new_[1206]_ ;
  assign \new_[7106]_  = \new_[1207]_  | \new_[7105]_ ;
  assign \new_[7107]_  = \new_[7106]_  | \new_[7101]_ ;
  assign \new_[7108]_  = \new_[7107]_  | \new_[7096]_ ;
  assign \new_[7112]_  = \new_[1202]_  | \new_[1203]_ ;
  assign \new_[7113]_  = \new_[1204]_  | \new_[7112]_ ;
  assign \new_[7117]_  = \new_[1199]_  | \new_[1200]_ ;
  assign \new_[7118]_  = \new_[1201]_  | \new_[7117]_ ;
  assign \new_[7119]_  = \new_[7118]_  | \new_[7113]_ ;
  assign \new_[7123]_  = \new_[1196]_  | \new_[1197]_ ;
  assign \new_[7124]_  = \new_[1198]_  | \new_[7123]_ ;
  assign \new_[7127]_  = \new_[1194]_  | \new_[1195]_ ;
  assign \new_[7130]_  = \new_[1192]_  | \new_[1193]_ ;
  assign \new_[7131]_  = \new_[7130]_  | \new_[7127]_ ;
  assign \new_[7132]_  = \new_[7131]_  | \new_[7124]_ ;
  assign \new_[7133]_  = \new_[7132]_  | \new_[7119]_ ;
  assign \new_[7134]_  = \new_[7133]_  | \new_[7108]_ ;
  assign \new_[7135]_  = \new_[7134]_  | \new_[7085]_ ;
  assign \new_[7136]_  = \new_[7135]_  | \new_[7036]_ ;
  assign \new_[7137]_  = \new_[7136]_  | \new_[6939]_ ;
  assign \new_[7138]_  = \new_[7137]_  | \new_[6742]_ ;
  assign \new_[7142]_  = \new_[1189]_  | \new_[1190]_ ;
  assign \new_[7143]_  = \new_[1191]_  | \new_[7142]_ ;
  assign \new_[7147]_  = \new_[1186]_  | \new_[1187]_ ;
  assign \new_[7148]_  = \new_[1188]_  | \new_[7147]_ ;
  assign \new_[7149]_  = \new_[7148]_  | \new_[7143]_ ;
  assign \new_[7153]_  = \new_[1183]_  | \new_[1184]_ ;
  assign \new_[7154]_  = \new_[1185]_  | \new_[7153]_ ;
  assign \new_[7158]_  = \new_[1180]_  | \new_[1181]_ ;
  assign \new_[7159]_  = \new_[1182]_  | \new_[7158]_ ;
  assign \new_[7160]_  = \new_[7159]_  | \new_[7154]_ ;
  assign \new_[7161]_  = \new_[7160]_  | \new_[7149]_ ;
  assign \new_[7165]_  = \new_[1177]_  | \new_[1178]_ ;
  assign \new_[7166]_  = \new_[1179]_  | \new_[7165]_ ;
  assign \new_[7170]_  = \new_[1174]_  | \new_[1175]_ ;
  assign \new_[7171]_  = \new_[1176]_  | \new_[7170]_ ;
  assign \new_[7172]_  = \new_[7171]_  | \new_[7166]_ ;
  assign \new_[7176]_  = \new_[1171]_  | \new_[1172]_ ;
  assign \new_[7177]_  = \new_[1173]_  | \new_[7176]_ ;
  assign \new_[7181]_  = \new_[1168]_  | \new_[1169]_ ;
  assign \new_[7182]_  = \new_[1170]_  | \new_[7181]_ ;
  assign \new_[7183]_  = \new_[7182]_  | \new_[7177]_ ;
  assign \new_[7184]_  = \new_[7183]_  | \new_[7172]_ ;
  assign \new_[7185]_  = \new_[7184]_  | \new_[7161]_ ;
  assign \new_[7189]_  = \new_[1165]_  | \new_[1166]_ ;
  assign \new_[7190]_  = \new_[1167]_  | \new_[7189]_ ;
  assign \new_[7194]_  = \new_[1162]_  | \new_[1163]_ ;
  assign \new_[7195]_  = \new_[1164]_  | \new_[7194]_ ;
  assign \new_[7196]_  = \new_[7195]_  | \new_[7190]_ ;
  assign \new_[7200]_  = \new_[1159]_  | \new_[1160]_ ;
  assign \new_[7201]_  = \new_[1161]_  | \new_[7200]_ ;
  assign \new_[7205]_  = \new_[1156]_  | \new_[1157]_ ;
  assign \new_[7206]_  = \new_[1158]_  | \new_[7205]_ ;
  assign \new_[7207]_  = \new_[7206]_  | \new_[7201]_ ;
  assign \new_[7208]_  = \new_[7207]_  | \new_[7196]_ ;
  assign \new_[7212]_  = \new_[1153]_  | \new_[1154]_ ;
  assign \new_[7213]_  = \new_[1155]_  | \new_[7212]_ ;
  assign \new_[7217]_  = \new_[1150]_  | \new_[1151]_ ;
  assign \new_[7218]_  = \new_[1152]_  | \new_[7217]_ ;
  assign \new_[7219]_  = \new_[7218]_  | \new_[7213]_ ;
  assign \new_[7223]_  = \new_[1147]_  | \new_[1148]_ ;
  assign \new_[7224]_  = \new_[1149]_  | \new_[7223]_ ;
  assign \new_[7227]_  = \new_[1145]_  | \new_[1146]_ ;
  assign \new_[7230]_  = \new_[1143]_  | \new_[1144]_ ;
  assign \new_[7231]_  = \new_[7230]_  | \new_[7227]_ ;
  assign \new_[7232]_  = \new_[7231]_  | \new_[7224]_ ;
  assign \new_[7233]_  = \new_[7232]_  | \new_[7219]_ ;
  assign \new_[7234]_  = \new_[7233]_  | \new_[7208]_ ;
  assign \new_[7235]_  = \new_[7234]_  | \new_[7185]_ ;
  assign \new_[7239]_  = \new_[1140]_  | \new_[1141]_ ;
  assign \new_[7240]_  = \new_[1142]_  | \new_[7239]_ ;
  assign \new_[7244]_  = \new_[1137]_  | \new_[1138]_ ;
  assign \new_[7245]_  = \new_[1139]_  | \new_[7244]_ ;
  assign \new_[7246]_  = \new_[7245]_  | \new_[7240]_ ;
  assign \new_[7250]_  = \new_[1134]_  | \new_[1135]_ ;
  assign \new_[7251]_  = \new_[1136]_  | \new_[7250]_ ;
  assign \new_[7255]_  = \new_[1131]_  | \new_[1132]_ ;
  assign \new_[7256]_  = \new_[1133]_  | \new_[7255]_ ;
  assign \new_[7257]_  = \new_[7256]_  | \new_[7251]_ ;
  assign \new_[7258]_  = \new_[7257]_  | \new_[7246]_ ;
  assign \new_[7262]_  = \new_[1128]_  | \new_[1129]_ ;
  assign \new_[7263]_  = \new_[1130]_  | \new_[7262]_ ;
  assign \new_[7267]_  = \new_[1125]_  | \new_[1126]_ ;
  assign \new_[7268]_  = \new_[1127]_  | \new_[7267]_ ;
  assign \new_[7269]_  = \new_[7268]_  | \new_[7263]_ ;
  assign \new_[7273]_  = \new_[1122]_  | \new_[1123]_ ;
  assign \new_[7274]_  = \new_[1124]_  | \new_[7273]_ ;
  assign \new_[7277]_  = \new_[1120]_  | \new_[1121]_ ;
  assign \new_[7280]_  = \new_[1118]_  | \new_[1119]_ ;
  assign \new_[7281]_  = \new_[7280]_  | \new_[7277]_ ;
  assign \new_[7282]_  = \new_[7281]_  | \new_[7274]_ ;
  assign \new_[7283]_  = \new_[7282]_  | \new_[7269]_ ;
  assign \new_[7284]_  = \new_[7283]_  | \new_[7258]_ ;
  assign \new_[7288]_  = \new_[1115]_  | \new_[1116]_ ;
  assign \new_[7289]_  = \new_[1117]_  | \new_[7288]_ ;
  assign \new_[7293]_  = \new_[1112]_  | \new_[1113]_ ;
  assign \new_[7294]_  = \new_[1114]_  | \new_[7293]_ ;
  assign \new_[7295]_  = \new_[7294]_  | \new_[7289]_ ;
  assign \new_[7299]_  = \new_[1109]_  | \new_[1110]_ ;
  assign \new_[7300]_  = \new_[1111]_  | \new_[7299]_ ;
  assign \new_[7304]_  = \new_[1106]_  | \new_[1107]_ ;
  assign \new_[7305]_  = \new_[1108]_  | \new_[7304]_ ;
  assign \new_[7306]_  = \new_[7305]_  | \new_[7300]_ ;
  assign \new_[7307]_  = \new_[7306]_  | \new_[7295]_ ;
  assign \new_[7311]_  = \new_[1103]_  | \new_[1104]_ ;
  assign \new_[7312]_  = \new_[1105]_  | \new_[7311]_ ;
  assign \new_[7316]_  = \new_[1100]_  | \new_[1101]_ ;
  assign \new_[7317]_  = \new_[1102]_  | \new_[7316]_ ;
  assign \new_[7318]_  = \new_[7317]_  | \new_[7312]_ ;
  assign \new_[7322]_  = \new_[1097]_  | \new_[1098]_ ;
  assign \new_[7323]_  = \new_[1099]_  | \new_[7322]_ ;
  assign \new_[7326]_  = \new_[1095]_  | \new_[1096]_ ;
  assign \new_[7329]_  = \new_[1093]_  | \new_[1094]_ ;
  assign \new_[7330]_  = \new_[7329]_  | \new_[7326]_ ;
  assign \new_[7331]_  = \new_[7330]_  | \new_[7323]_ ;
  assign \new_[7332]_  = \new_[7331]_  | \new_[7318]_ ;
  assign \new_[7333]_  = \new_[7332]_  | \new_[7307]_ ;
  assign \new_[7334]_  = \new_[7333]_  | \new_[7284]_ ;
  assign \new_[7335]_  = \new_[7334]_  | \new_[7235]_ ;
  assign \new_[7339]_  = \new_[1090]_  | \new_[1091]_ ;
  assign \new_[7340]_  = \new_[1092]_  | \new_[7339]_ ;
  assign \new_[7344]_  = \new_[1087]_  | \new_[1088]_ ;
  assign \new_[7345]_  = \new_[1089]_  | \new_[7344]_ ;
  assign \new_[7346]_  = \new_[7345]_  | \new_[7340]_ ;
  assign \new_[7350]_  = \new_[1084]_  | \new_[1085]_ ;
  assign \new_[7351]_  = \new_[1086]_  | \new_[7350]_ ;
  assign \new_[7355]_  = \new_[1081]_  | \new_[1082]_ ;
  assign \new_[7356]_  = \new_[1083]_  | \new_[7355]_ ;
  assign \new_[7357]_  = \new_[7356]_  | \new_[7351]_ ;
  assign \new_[7358]_  = \new_[7357]_  | \new_[7346]_ ;
  assign \new_[7362]_  = \new_[1078]_  | \new_[1079]_ ;
  assign \new_[7363]_  = \new_[1080]_  | \new_[7362]_ ;
  assign \new_[7367]_  = \new_[1075]_  | \new_[1076]_ ;
  assign \new_[7368]_  = \new_[1077]_  | \new_[7367]_ ;
  assign \new_[7369]_  = \new_[7368]_  | \new_[7363]_ ;
  assign \new_[7373]_  = \new_[1072]_  | \new_[1073]_ ;
  assign \new_[7374]_  = \new_[1074]_  | \new_[7373]_ ;
  assign \new_[7378]_  = \new_[1069]_  | \new_[1070]_ ;
  assign \new_[7379]_  = \new_[1071]_  | \new_[7378]_ ;
  assign \new_[7380]_  = \new_[7379]_  | \new_[7374]_ ;
  assign \new_[7381]_  = \new_[7380]_  | \new_[7369]_ ;
  assign \new_[7382]_  = \new_[7381]_  | \new_[7358]_ ;
  assign \new_[7386]_  = \new_[1066]_  | \new_[1067]_ ;
  assign \new_[7387]_  = \new_[1068]_  | \new_[7386]_ ;
  assign \new_[7391]_  = \new_[1063]_  | \new_[1064]_ ;
  assign \new_[7392]_  = \new_[1065]_  | \new_[7391]_ ;
  assign \new_[7393]_  = \new_[7392]_  | \new_[7387]_ ;
  assign \new_[7397]_  = \new_[1060]_  | \new_[1061]_ ;
  assign \new_[7398]_  = \new_[1062]_  | \new_[7397]_ ;
  assign \new_[7402]_  = \new_[1057]_  | \new_[1058]_ ;
  assign \new_[7403]_  = \new_[1059]_  | \new_[7402]_ ;
  assign \new_[7404]_  = \new_[7403]_  | \new_[7398]_ ;
  assign \new_[7405]_  = \new_[7404]_  | \new_[7393]_ ;
  assign \new_[7409]_  = \new_[1054]_  | \new_[1055]_ ;
  assign \new_[7410]_  = \new_[1056]_  | \new_[7409]_ ;
  assign \new_[7414]_  = \new_[1051]_  | \new_[1052]_ ;
  assign \new_[7415]_  = \new_[1053]_  | \new_[7414]_ ;
  assign \new_[7416]_  = \new_[7415]_  | \new_[7410]_ ;
  assign \new_[7420]_  = \new_[1048]_  | \new_[1049]_ ;
  assign \new_[7421]_  = \new_[1050]_  | \new_[7420]_ ;
  assign \new_[7424]_  = \new_[1046]_  | \new_[1047]_ ;
  assign \new_[7427]_  = \new_[1044]_  | \new_[1045]_ ;
  assign \new_[7428]_  = \new_[7427]_  | \new_[7424]_ ;
  assign \new_[7429]_  = \new_[7428]_  | \new_[7421]_ ;
  assign \new_[7430]_  = \new_[7429]_  | \new_[7416]_ ;
  assign \new_[7431]_  = \new_[7430]_  | \new_[7405]_ ;
  assign \new_[7432]_  = \new_[7431]_  | \new_[7382]_ ;
  assign \new_[7436]_  = \new_[1041]_  | \new_[1042]_ ;
  assign \new_[7437]_  = \new_[1043]_  | \new_[7436]_ ;
  assign \new_[7441]_  = \new_[1038]_  | \new_[1039]_ ;
  assign \new_[7442]_  = \new_[1040]_  | \new_[7441]_ ;
  assign \new_[7443]_  = \new_[7442]_  | \new_[7437]_ ;
  assign \new_[7447]_  = \new_[1035]_  | \new_[1036]_ ;
  assign \new_[7448]_  = \new_[1037]_  | \new_[7447]_ ;
  assign \new_[7452]_  = \new_[1032]_  | \new_[1033]_ ;
  assign \new_[7453]_  = \new_[1034]_  | \new_[7452]_ ;
  assign \new_[7454]_  = \new_[7453]_  | \new_[7448]_ ;
  assign \new_[7455]_  = \new_[7454]_  | \new_[7443]_ ;
  assign \new_[7459]_  = \new_[1029]_  | \new_[1030]_ ;
  assign \new_[7460]_  = \new_[1031]_  | \new_[7459]_ ;
  assign \new_[7464]_  = \new_[1026]_  | \new_[1027]_ ;
  assign \new_[7465]_  = \new_[1028]_  | \new_[7464]_ ;
  assign \new_[7466]_  = \new_[7465]_  | \new_[7460]_ ;
  assign \new_[7470]_  = \new_[1023]_  | \new_[1024]_ ;
  assign \new_[7471]_  = \new_[1025]_  | \new_[7470]_ ;
  assign \new_[7474]_  = \new_[1021]_  | \new_[1022]_ ;
  assign \new_[7477]_  = \new_[1019]_  | \new_[1020]_ ;
  assign \new_[7478]_  = \new_[7477]_  | \new_[7474]_ ;
  assign \new_[7479]_  = \new_[7478]_  | \new_[7471]_ ;
  assign \new_[7480]_  = \new_[7479]_  | \new_[7466]_ ;
  assign \new_[7481]_  = \new_[7480]_  | \new_[7455]_ ;
  assign \new_[7485]_  = \new_[1016]_  | \new_[1017]_ ;
  assign \new_[7486]_  = \new_[1018]_  | \new_[7485]_ ;
  assign \new_[7490]_  = \new_[1013]_  | \new_[1014]_ ;
  assign \new_[7491]_  = \new_[1015]_  | \new_[7490]_ ;
  assign \new_[7492]_  = \new_[7491]_  | \new_[7486]_ ;
  assign \new_[7496]_  = \new_[1010]_  | \new_[1011]_ ;
  assign \new_[7497]_  = \new_[1012]_  | \new_[7496]_ ;
  assign \new_[7501]_  = \new_[1007]_  | \new_[1008]_ ;
  assign \new_[7502]_  = \new_[1009]_  | \new_[7501]_ ;
  assign \new_[7503]_  = \new_[7502]_  | \new_[7497]_ ;
  assign \new_[7504]_  = \new_[7503]_  | \new_[7492]_ ;
  assign \new_[7508]_  = \new_[1004]_  | \new_[1005]_ ;
  assign \new_[7509]_  = \new_[1006]_  | \new_[7508]_ ;
  assign \new_[7513]_  = \new_[1001]_  | \new_[1002]_ ;
  assign \new_[7514]_  = \new_[1003]_  | \new_[7513]_ ;
  assign \new_[7515]_  = \new_[7514]_  | \new_[7509]_ ;
  assign \new_[7519]_  = \new_[998]_  | \new_[999]_ ;
  assign \new_[7520]_  = \new_[1000]_  | \new_[7519]_ ;
  assign \new_[7523]_  = \new_[996]_  | \new_[997]_ ;
  assign \new_[7526]_  = \new_[994]_  | \new_[995]_ ;
  assign \new_[7527]_  = \new_[7526]_  | \new_[7523]_ ;
  assign \new_[7528]_  = \new_[7527]_  | \new_[7520]_ ;
  assign \new_[7529]_  = \new_[7528]_  | \new_[7515]_ ;
  assign \new_[7530]_  = \new_[7529]_  | \new_[7504]_ ;
  assign \new_[7531]_  = \new_[7530]_  | \new_[7481]_ ;
  assign \new_[7532]_  = \new_[7531]_  | \new_[7432]_ ;
  assign \new_[7533]_  = \new_[7532]_  | \new_[7335]_ ;
  assign \new_[7537]_  = \new_[991]_  | \new_[992]_ ;
  assign \new_[7538]_  = \new_[993]_  | \new_[7537]_ ;
  assign \new_[7542]_  = \new_[988]_  | \new_[989]_ ;
  assign \new_[7543]_  = \new_[990]_  | \new_[7542]_ ;
  assign \new_[7544]_  = \new_[7543]_  | \new_[7538]_ ;
  assign \new_[7548]_  = \new_[985]_  | \new_[986]_ ;
  assign \new_[7549]_  = \new_[987]_  | \new_[7548]_ ;
  assign \new_[7553]_  = \new_[982]_  | \new_[983]_ ;
  assign \new_[7554]_  = \new_[984]_  | \new_[7553]_ ;
  assign \new_[7555]_  = \new_[7554]_  | \new_[7549]_ ;
  assign \new_[7556]_  = \new_[7555]_  | \new_[7544]_ ;
  assign \new_[7560]_  = \new_[979]_  | \new_[980]_ ;
  assign \new_[7561]_  = \new_[981]_  | \new_[7560]_ ;
  assign \new_[7565]_  = \new_[976]_  | \new_[977]_ ;
  assign \new_[7566]_  = \new_[978]_  | \new_[7565]_ ;
  assign \new_[7567]_  = \new_[7566]_  | \new_[7561]_ ;
  assign \new_[7571]_  = \new_[973]_  | \new_[974]_ ;
  assign \new_[7572]_  = \new_[975]_  | \new_[7571]_ ;
  assign \new_[7576]_  = \new_[970]_  | \new_[971]_ ;
  assign \new_[7577]_  = \new_[972]_  | \new_[7576]_ ;
  assign \new_[7578]_  = \new_[7577]_  | \new_[7572]_ ;
  assign \new_[7579]_  = \new_[7578]_  | \new_[7567]_ ;
  assign \new_[7580]_  = \new_[7579]_  | \new_[7556]_ ;
  assign \new_[7584]_  = \new_[967]_  | \new_[968]_ ;
  assign \new_[7585]_  = \new_[969]_  | \new_[7584]_ ;
  assign \new_[7589]_  = \new_[964]_  | \new_[965]_ ;
  assign \new_[7590]_  = \new_[966]_  | \new_[7589]_ ;
  assign \new_[7591]_  = \new_[7590]_  | \new_[7585]_ ;
  assign \new_[7595]_  = \new_[961]_  | \new_[962]_ ;
  assign \new_[7596]_  = \new_[963]_  | \new_[7595]_ ;
  assign \new_[7600]_  = \new_[958]_  | \new_[959]_ ;
  assign \new_[7601]_  = \new_[960]_  | \new_[7600]_ ;
  assign \new_[7602]_  = \new_[7601]_  | \new_[7596]_ ;
  assign \new_[7603]_  = \new_[7602]_  | \new_[7591]_ ;
  assign \new_[7607]_  = \new_[955]_  | \new_[956]_ ;
  assign \new_[7608]_  = \new_[957]_  | \new_[7607]_ ;
  assign \new_[7612]_  = \new_[952]_  | \new_[953]_ ;
  assign \new_[7613]_  = \new_[954]_  | \new_[7612]_ ;
  assign \new_[7614]_  = \new_[7613]_  | \new_[7608]_ ;
  assign \new_[7618]_  = \new_[949]_  | \new_[950]_ ;
  assign \new_[7619]_  = \new_[951]_  | \new_[7618]_ ;
  assign \new_[7622]_  = \new_[947]_  | \new_[948]_ ;
  assign \new_[7625]_  = \new_[945]_  | \new_[946]_ ;
  assign \new_[7626]_  = \new_[7625]_  | \new_[7622]_ ;
  assign \new_[7627]_  = \new_[7626]_  | \new_[7619]_ ;
  assign \new_[7628]_  = \new_[7627]_  | \new_[7614]_ ;
  assign \new_[7629]_  = \new_[7628]_  | \new_[7603]_ ;
  assign \new_[7630]_  = \new_[7629]_  | \new_[7580]_ ;
  assign \new_[7634]_  = \new_[942]_  | \new_[943]_ ;
  assign \new_[7635]_  = \new_[944]_  | \new_[7634]_ ;
  assign \new_[7639]_  = \new_[939]_  | \new_[940]_ ;
  assign \new_[7640]_  = \new_[941]_  | \new_[7639]_ ;
  assign \new_[7641]_  = \new_[7640]_  | \new_[7635]_ ;
  assign \new_[7645]_  = \new_[936]_  | \new_[937]_ ;
  assign \new_[7646]_  = \new_[938]_  | \new_[7645]_ ;
  assign \new_[7650]_  = \new_[933]_  | \new_[934]_ ;
  assign \new_[7651]_  = \new_[935]_  | \new_[7650]_ ;
  assign \new_[7652]_  = \new_[7651]_  | \new_[7646]_ ;
  assign \new_[7653]_  = \new_[7652]_  | \new_[7641]_ ;
  assign \new_[7657]_  = \new_[930]_  | \new_[931]_ ;
  assign \new_[7658]_  = \new_[932]_  | \new_[7657]_ ;
  assign \new_[7662]_  = \new_[927]_  | \new_[928]_ ;
  assign \new_[7663]_  = \new_[929]_  | \new_[7662]_ ;
  assign \new_[7664]_  = \new_[7663]_  | \new_[7658]_ ;
  assign \new_[7668]_  = \new_[924]_  | \new_[925]_ ;
  assign \new_[7669]_  = \new_[926]_  | \new_[7668]_ ;
  assign \new_[7672]_  = \new_[922]_  | \new_[923]_ ;
  assign \new_[7675]_  = \new_[920]_  | \new_[921]_ ;
  assign \new_[7676]_  = \new_[7675]_  | \new_[7672]_ ;
  assign \new_[7677]_  = \new_[7676]_  | \new_[7669]_ ;
  assign \new_[7678]_  = \new_[7677]_  | \new_[7664]_ ;
  assign \new_[7679]_  = \new_[7678]_  | \new_[7653]_ ;
  assign \new_[7683]_  = \new_[917]_  | \new_[918]_ ;
  assign \new_[7684]_  = \new_[919]_  | \new_[7683]_ ;
  assign \new_[7688]_  = \new_[914]_  | \new_[915]_ ;
  assign \new_[7689]_  = \new_[916]_  | \new_[7688]_ ;
  assign \new_[7690]_  = \new_[7689]_  | \new_[7684]_ ;
  assign \new_[7694]_  = \new_[911]_  | \new_[912]_ ;
  assign \new_[7695]_  = \new_[913]_  | \new_[7694]_ ;
  assign \new_[7699]_  = \new_[908]_  | \new_[909]_ ;
  assign \new_[7700]_  = \new_[910]_  | \new_[7699]_ ;
  assign \new_[7701]_  = \new_[7700]_  | \new_[7695]_ ;
  assign \new_[7702]_  = \new_[7701]_  | \new_[7690]_ ;
  assign \new_[7706]_  = \new_[905]_  | \new_[906]_ ;
  assign \new_[7707]_  = \new_[907]_  | \new_[7706]_ ;
  assign \new_[7711]_  = \new_[902]_  | \new_[903]_ ;
  assign \new_[7712]_  = \new_[904]_  | \new_[7711]_ ;
  assign \new_[7713]_  = \new_[7712]_  | \new_[7707]_ ;
  assign \new_[7717]_  = \new_[899]_  | \new_[900]_ ;
  assign \new_[7718]_  = \new_[901]_  | \new_[7717]_ ;
  assign \new_[7721]_  = \new_[897]_  | \new_[898]_ ;
  assign \new_[7724]_  = \new_[895]_  | \new_[896]_ ;
  assign \new_[7725]_  = \new_[7724]_  | \new_[7721]_ ;
  assign \new_[7726]_  = \new_[7725]_  | \new_[7718]_ ;
  assign \new_[7727]_  = \new_[7726]_  | \new_[7713]_ ;
  assign \new_[7728]_  = \new_[7727]_  | \new_[7702]_ ;
  assign \new_[7729]_  = \new_[7728]_  | \new_[7679]_ ;
  assign \new_[7730]_  = \new_[7729]_  | \new_[7630]_ ;
  assign \new_[7734]_  = \new_[892]_  | \new_[893]_ ;
  assign \new_[7735]_  = \new_[894]_  | \new_[7734]_ ;
  assign \new_[7739]_  = \new_[889]_  | \new_[890]_ ;
  assign \new_[7740]_  = \new_[891]_  | \new_[7739]_ ;
  assign \new_[7741]_  = \new_[7740]_  | \new_[7735]_ ;
  assign \new_[7745]_  = \new_[886]_  | \new_[887]_ ;
  assign \new_[7746]_  = \new_[888]_  | \new_[7745]_ ;
  assign \new_[7750]_  = \new_[883]_  | \new_[884]_ ;
  assign \new_[7751]_  = \new_[885]_  | \new_[7750]_ ;
  assign \new_[7752]_  = \new_[7751]_  | \new_[7746]_ ;
  assign \new_[7753]_  = \new_[7752]_  | \new_[7741]_ ;
  assign \new_[7757]_  = \new_[880]_  | \new_[881]_ ;
  assign \new_[7758]_  = \new_[882]_  | \new_[7757]_ ;
  assign \new_[7762]_  = \new_[877]_  | \new_[878]_ ;
  assign \new_[7763]_  = \new_[879]_  | \new_[7762]_ ;
  assign \new_[7764]_  = \new_[7763]_  | \new_[7758]_ ;
  assign \new_[7768]_  = \new_[874]_  | \new_[875]_ ;
  assign \new_[7769]_  = \new_[876]_  | \new_[7768]_ ;
  assign \new_[7772]_  = \new_[872]_  | \new_[873]_ ;
  assign \new_[7775]_  = \new_[870]_  | \new_[871]_ ;
  assign \new_[7776]_  = \new_[7775]_  | \new_[7772]_ ;
  assign \new_[7777]_  = \new_[7776]_  | \new_[7769]_ ;
  assign \new_[7778]_  = \new_[7777]_  | \new_[7764]_ ;
  assign \new_[7779]_  = \new_[7778]_  | \new_[7753]_ ;
  assign \new_[7783]_  = \new_[867]_  | \new_[868]_ ;
  assign \new_[7784]_  = \new_[869]_  | \new_[7783]_ ;
  assign \new_[7788]_  = \new_[864]_  | \new_[865]_ ;
  assign \new_[7789]_  = \new_[866]_  | \new_[7788]_ ;
  assign \new_[7790]_  = \new_[7789]_  | \new_[7784]_ ;
  assign \new_[7794]_  = \new_[861]_  | \new_[862]_ ;
  assign \new_[7795]_  = \new_[863]_  | \new_[7794]_ ;
  assign \new_[7799]_  = \new_[858]_  | \new_[859]_ ;
  assign \new_[7800]_  = \new_[860]_  | \new_[7799]_ ;
  assign \new_[7801]_  = \new_[7800]_  | \new_[7795]_ ;
  assign \new_[7802]_  = \new_[7801]_  | \new_[7790]_ ;
  assign \new_[7806]_  = \new_[855]_  | \new_[856]_ ;
  assign \new_[7807]_  = \new_[857]_  | \new_[7806]_ ;
  assign \new_[7811]_  = \new_[852]_  | \new_[853]_ ;
  assign \new_[7812]_  = \new_[854]_  | \new_[7811]_ ;
  assign \new_[7813]_  = \new_[7812]_  | \new_[7807]_ ;
  assign \new_[7817]_  = \new_[849]_  | \new_[850]_ ;
  assign \new_[7818]_  = \new_[851]_  | \new_[7817]_ ;
  assign \new_[7821]_  = \new_[847]_  | \new_[848]_ ;
  assign \new_[7824]_  = \new_[845]_  | \new_[846]_ ;
  assign \new_[7825]_  = \new_[7824]_  | \new_[7821]_ ;
  assign \new_[7826]_  = \new_[7825]_  | \new_[7818]_ ;
  assign \new_[7827]_  = \new_[7826]_  | \new_[7813]_ ;
  assign \new_[7828]_  = \new_[7827]_  | \new_[7802]_ ;
  assign \new_[7829]_  = \new_[7828]_  | \new_[7779]_ ;
  assign \new_[7833]_  = \new_[842]_  | \new_[843]_ ;
  assign \new_[7834]_  = \new_[844]_  | \new_[7833]_ ;
  assign \new_[7838]_  = \new_[839]_  | \new_[840]_ ;
  assign \new_[7839]_  = \new_[841]_  | \new_[7838]_ ;
  assign \new_[7840]_  = \new_[7839]_  | \new_[7834]_ ;
  assign \new_[7844]_  = \new_[836]_  | \new_[837]_ ;
  assign \new_[7845]_  = \new_[838]_  | \new_[7844]_ ;
  assign \new_[7849]_  = \new_[833]_  | \new_[834]_ ;
  assign \new_[7850]_  = \new_[835]_  | \new_[7849]_ ;
  assign \new_[7851]_  = \new_[7850]_  | \new_[7845]_ ;
  assign \new_[7852]_  = \new_[7851]_  | \new_[7840]_ ;
  assign \new_[7856]_  = \new_[830]_  | \new_[831]_ ;
  assign \new_[7857]_  = \new_[832]_  | \new_[7856]_ ;
  assign \new_[7861]_  = \new_[827]_  | \new_[828]_ ;
  assign \new_[7862]_  = \new_[829]_  | \new_[7861]_ ;
  assign \new_[7863]_  = \new_[7862]_  | \new_[7857]_ ;
  assign \new_[7867]_  = \new_[824]_  | \new_[825]_ ;
  assign \new_[7868]_  = \new_[826]_  | \new_[7867]_ ;
  assign \new_[7871]_  = \new_[822]_  | \new_[823]_ ;
  assign \new_[7874]_  = \new_[820]_  | \new_[821]_ ;
  assign \new_[7875]_  = \new_[7874]_  | \new_[7871]_ ;
  assign \new_[7876]_  = \new_[7875]_  | \new_[7868]_ ;
  assign \new_[7877]_  = \new_[7876]_  | \new_[7863]_ ;
  assign \new_[7878]_  = \new_[7877]_  | \new_[7852]_ ;
  assign \new_[7882]_  = \new_[817]_  | \new_[818]_ ;
  assign \new_[7883]_  = \new_[819]_  | \new_[7882]_ ;
  assign \new_[7887]_  = \new_[814]_  | \new_[815]_ ;
  assign \new_[7888]_  = \new_[816]_  | \new_[7887]_ ;
  assign \new_[7889]_  = \new_[7888]_  | \new_[7883]_ ;
  assign \new_[7893]_  = \new_[811]_  | \new_[812]_ ;
  assign \new_[7894]_  = \new_[813]_  | \new_[7893]_ ;
  assign \new_[7898]_  = \new_[808]_  | \new_[809]_ ;
  assign \new_[7899]_  = \new_[810]_  | \new_[7898]_ ;
  assign \new_[7900]_  = \new_[7899]_  | \new_[7894]_ ;
  assign \new_[7901]_  = \new_[7900]_  | \new_[7889]_ ;
  assign \new_[7905]_  = \new_[805]_  | \new_[806]_ ;
  assign \new_[7906]_  = \new_[807]_  | \new_[7905]_ ;
  assign \new_[7910]_  = \new_[802]_  | \new_[803]_ ;
  assign \new_[7911]_  = \new_[804]_  | \new_[7910]_ ;
  assign \new_[7912]_  = \new_[7911]_  | \new_[7906]_ ;
  assign \new_[7916]_  = \new_[799]_  | \new_[800]_ ;
  assign \new_[7917]_  = \new_[801]_  | \new_[7916]_ ;
  assign \new_[7920]_  = \new_[797]_  | \new_[798]_ ;
  assign \new_[7923]_  = \new_[795]_  | \new_[796]_ ;
  assign \new_[7924]_  = \new_[7923]_  | \new_[7920]_ ;
  assign \new_[7925]_  = \new_[7924]_  | \new_[7917]_ ;
  assign \new_[7926]_  = \new_[7925]_  | \new_[7912]_ ;
  assign \new_[7927]_  = \new_[7926]_  | \new_[7901]_ ;
  assign \new_[7928]_  = \new_[7927]_  | \new_[7878]_ ;
  assign \new_[7929]_  = \new_[7928]_  | \new_[7829]_ ;
  assign \new_[7930]_  = \new_[7929]_  | \new_[7730]_ ;
  assign \new_[7931]_  = \new_[7930]_  | \new_[7533]_ ;
  assign \new_[7932]_  = \new_[7931]_  | \new_[7138]_ ;
  assign \new_[7936]_  = \new_[792]_  | \new_[793]_ ;
  assign \new_[7937]_  = \new_[794]_  | \new_[7936]_ ;
  assign \new_[7941]_  = \new_[789]_  | \new_[790]_ ;
  assign \new_[7942]_  = \new_[791]_  | \new_[7941]_ ;
  assign \new_[7943]_  = \new_[7942]_  | \new_[7937]_ ;
  assign \new_[7947]_  = \new_[786]_  | \new_[787]_ ;
  assign \new_[7948]_  = \new_[788]_  | \new_[7947]_ ;
  assign \new_[7952]_  = \new_[783]_  | \new_[784]_ ;
  assign \new_[7953]_  = \new_[785]_  | \new_[7952]_ ;
  assign \new_[7954]_  = \new_[7953]_  | \new_[7948]_ ;
  assign \new_[7955]_  = \new_[7954]_  | \new_[7943]_ ;
  assign \new_[7959]_  = \new_[780]_  | \new_[781]_ ;
  assign \new_[7960]_  = \new_[782]_  | \new_[7959]_ ;
  assign \new_[7964]_  = \new_[777]_  | \new_[778]_ ;
  assign \new_[7965]_  = \new_[779]_  | \new_[7964]_ ;
  assign \new_[7966]_  = \new_[7965]_  | \new_[7960]_ ;
  assign \new_[7970]_  = \new_[774]_  | \new_[775]_ ;
  assign \new_[7971]_  = \new_[776]_  | \new_[7970]_ ;
  assign \new_[7975]_  = \new_[771]_  | \new_[772]_ ;
  assign \new_[7976]_  = \new_[773]_  | \new_[7975]_ ;
  assign \new_[7977]_  = \new_[7976]_  | \new_[7971]_ ;
  assign \new_[7978]_  = \new_[7977]_  | \new_[7966]_ ;
  assign \new_[7979]_  = \new_[7978]_  | \new_[7955]_ ;
  assign \new_[7983]_  = \new_[768]_  | \new_[769]_ ;
  assign \new_[7984]_  = \new_[770]_  | \new_[7983]_ ;
  assign \new_[7988]_  = \new_[765]_  | \new_[766]_ ;
  assign \new_[7989]_  = \new_[767]_  | \new_[7988]_ ;
  assign \new_[7990]_  = \new_[7989]_  | \new_[7984]_ ;
  assign \new_[7994]_  = \new_[762]_  | \new_[763]_ ;
  assign \new_[7995]_  = \new_[764]_  | \new_[7994]_ ;
  assign \new_[7999]_  = \new_[759]_  | \new_[760]_ ;
  assign \new_[8000]_  = \new_[761]_  | \new_[7999]_ ;
  assign \new_[8001]_  = \new_[8000]_  | \new_[7995]_ ;
  assign \new_[8002]_  = \new_[8001]_  | \new_[7990]_ ;
  assign \new_[8006]_  = \new_[756]_  | \new_[757]_ ;
  assign \new_[8007]_  = \new_[758]_  | \new_[8006]_ ;
  assign \new_[8011]_  = \new_[753]_  | \new_[754]_ ;
  assign \new_[8012]_  = \new_[755]_  | \new_[8011]_ ;
  assign \new_[8013]_  = \new_[8012]_  | \new_[8007]_ ;
  assign \new_[8017]_  = \new_[750]_  | \new_[751]_ ;
  assign \new_[8018]_  = \new_[752]_  | \new_[8017]_ ;
  assign \new_[8021]_  = \new_[748]_  | \new_[749]_ ;
  assign \new_[8024]_  = \new_[746]_  | \new_[747]_ ;
  assign \new_[8025]_  = \new_[8024]_  | \new_[8021]_ ;
  assign \new_[8026]_  = \new_[8025]_  | \new_[8018]_ ;
  assign \new_[8027]_  = \new_[8026]_  | \new_[8013]_ ;
  assign \new_[8028]_  = \new_[8027]_  | \new_[8002]_ ;
  assign \new_[8029]_  = \new_[8028]_  | \new_[7979]_ ;
  assign \new_[8033]_  = \new_[743]_  | \new_[744]_ ;
  assign \new_[8034]_  = \new_[745]_  | \new_[8033]_ ;
  assign \new_[8038]_  = \new_[740]_  | \new_[741]_ ;
  assign \new_[8039]_  = \new_[742]_  | \new_[8038]_ ;
  assign \new_[8040]_  = \new_[8039]_  | \new_[8034]_ ;
  assign \new_[8044]_  = \new_[737]_  | \new_[738]_ ;
  assign \new_[8045]_  = \new_[739]_  | \new_[8044]_ ;
  assign \new_[8049]_  = \new_[734]_  | \new_[735]_ ;
  assign \new_[8050]_  = \new_[736]_  | \new_[8049]_ ;
  assign \new_[8051]_  = \new_[8050]_  | \new_[8045]_ ;
  assign \new_[8052]_  = \new_[8051]_  | \new_[8040]_ ;
  assign \new_[8056]_  = \new_[731]_  | \new_[732]_ ;
  assign \new_[8057]_  = \new_[733]_  | \new_[8056]_ ;
  assign \new_[8061]_  = \new_[728]_  | \new_[729]_ ;
  assign \new_[8062]_  = \new_[730]_  | \new_[8061]_ ;
  assign \new_[8063]_  = \new_[8062]_  | \new_[8057]_ ;
  assign \new_[8067]_  = \new_[725]_  | \new_[726]_ ;
  assign \new_[8068]_  = \new_[727]_  | \new_[8067]_ ;
  assign \new_[8071]_  = \new_[723]_  | \new_[724]_ ;
  assign \new_[8074]_  = \new_[721]_  | \new_[722]_ ;
  assign \new_[8075]_  = \new_[8074]_  | \new_[8071]_ ;
  assign \new_[8076]_  = \new_[8075]_  | \new_[8068]_ ;
  assign \new_[8077]_  = \new_[8076]_  | \new_[8063]_ ;
  assign \new_[8078]_  = \new_[8077]_  | \new_[8052]_ ;
  assign \new_[8082]_  = \new_[718]_  | \new_[719]_ ;
  assign \new_[8083]_  = \new_[720]_  | \new_[8082]_ ;
  assign \new_[8087]_  = \new_[715]_  | \new_[716]_ ;
  assign \new_[8088]_  = \new_[717]_  | \new_[8087]_ ;
  assign \new_[8089]_  = \new_[8088]_  | \new_[8083]_ ;
  assign \new_[8093]_  = \new_[712]_  | \new_[713]_ ;
  assign \new_[8094]_  = \new_[714]_  | \new_[8093]_ ;
  assign \new_[8098]_  = \new_[709]_  | \new_[710]_ ;
  assign \new_[8099]_  = \new_[711]_  | \new_[8098]_ ;
  assign \new_[8100]_  = \new_[8099]_  | \new_[8094]_ ;
  assign \new_[8101]_  = \new_[8100]_  | \new_[8089]_ ;
  assign \new_[8105]_  = \new_[706]_  | \new_[707]_ ;
  assign \new_[8106]_  = \new_[708]_  | \new_[8105]_ ;
  assign \new_[8110]_  = \new_[703]_  | \new_[704]_ ;
  assign \new_[8111]_  = \new_[705]_  | \new_[8110]_ ;
  assign \new_[8112]_  = \new_[8111]_  | \new_[8106]_ ;
  assign \new_[8116]_  = \new_[700]_  | \new_[701]_ ;
  assign \new_[8117]_  = \new_[702]_  | \new_[8116]_ ;
  assign \new_[8120]_  = \new_[698]_  | \new_[699]_ ;
  assign \new_[8123]_  = \new_[696]_  | \new_[697]_ ;
  assign \new_[8124]_  = \new_[8123]_  | \new_[8120]_ ;
  assign \new_[8125]_  = \new_[8124]_  | \new_[8117]_ ;
  assign \new_[8126]_  = \new_[8125]_  | \new_[8112]_ ;
  assign \new_[8127]_  = \new_[8126]_  | \new_[8101]_ ;
  assign \new_[8128]_  = \new_[8127]_  | \new_[8078]_ ;
  assign \new_[8129]_  = \new_[8128]_  | \new_[8029]_ ;
  assign \new_[8133]_  = \new_[693]_  | \new_[694]_ ;
  assign \new_[8134]_  = \new_[695]_  | \new_[8133]_ ;
  assign \new_[8138]_  = \new_[690]_  | \new_[691]_ ;
  assign \new_[8139]_  = \new_[692]_  | \new_[8138]_ ;
  assign \new_[8140]_  = \new_[8139]_  | \new_[8134]_ ;
  assign \new_[8144]_  = \new_[687]_  | \new_[688]_ ;
  assign \new_[8145]_  = \new_[689]_  | \new_[8144]_ ;
  assign \new_[8149]_  = \new_[684]_  | \new_[685]_ ;
  assign \new_[8150]_  = \new_[686]_  | \new_[8149]_ ;
  assign \new_[8151]_  = \new_[8150]_  | \new_[8145]_ ;
  assign \new_[8152]_  = \new_[8151]_  | \new_[8140]_ ;
  assign \new_[8156]_  = \new_[681]_  | \new_[682]_ ;
  assign \new_[8157]_  = \new_[683]_  | \new_[8156]_ ;
  assign \new_[8161]_  = \new_[678]_  | \new_[679]_ ;
  assign \new_[8162]_  = \new_[680]_  | \new_[8161]_ ;
  assign \new_[8163]_  = \new_[8162]_  | \new_[8157]_ ;
  assign \new_[8167]_  = \new_[675]_  | \new_[676]_ ;
  assign \new_[8168]_  = \new_[677]_  | \new_[8167]_ ;
  assign \new_[8172]_  = \new_[672]_  | \new_[673]_ ;
  assign \new_[8173]_  = \new_[674]_  | \new_[8172]_ ;
  assign \new_[8174]_  = \new_[8173]_  | \new_[8168]_ ;
  assign \new_[8175]_  = \new_[8174]_  | \new_[8163]_ ;
  assign \new_[8176]_  = \new_[8175]_  | \new_[8152]_ ;
  assign \new_[8180]_  = \new_[669]_  | \new_[670]_ ;
  assign \new_[8181]_  = \new_[671]_  | \new_[8180]_ ;
  assign \new_[8185]_  = \new_[666]_  | \new_[667]_ ;
  assign \new_[8186]_  = \new_[668]_  | \new_[8185]_ ;
  assign \new_[8187]_  = \new_[8186]_  | \new_[8181]_ ;
  assign \new_[8191]_  = \new_[663]_  | \new_[664]_ ;
  assign \new_[8192]_  = \new_[665]_  | \new_[8191]_ ;
  assign \new_[8196]_  = \new_[660]_  | \new_[661]_ ;
  assign \new_[8197]_  = \new_[662]_  | \new_[8196]_ ;
  assign \new_[8198]_  = \new_[8197]_  | \new_[8192]_ ;
  assign \new_[8199]_  = \new_[8198]_  | \new_[8187]_ ;
  assign \new_[8203]_  = \new_[657]_  | \new_[658]_ ;
  assign \new_[8204]_  = \new_[659]_  | \new_[8203]_ ;
  assign \new_[8208]_  = \new_[654]_  | \new_[655]_ ;
  assign \new_[8209]_  = \new_[656]_  | \new_[8208]_ ;
  assign \new_[8210]_  = \new_[8209]_  | \new_[8204]_ ;
  assign \new_[8214]_  = \new_[651]_  | \new_[652]_ ;
  assign \new_[8215]_  = \new_[653]_  | \new_[8214]_ ;
  assign \new_[8218]_  = \new_[649]_  | \new_[650]_ ;
  assign \new_[8221]_  = \new_[647]_  | \new_[648]_ ;
  assign \new_[8222]_  = \new_[8221]_  | \new_[8218]_ ;
  assign \new_[8223]_  = \new_[8222]_  | \new_[8215]_ ;
  assign \new_[8224]_  = \new_[8223]_  | \new_[8210]_ ;
  assign \new_[8225]_  = \new_[8224]_  | \new_[8199]_ ;
  assign \new_[8226]_  = \new_[8225]_  | \new_[8176]_ ;
  assign \new_[8230]_  = \new_[644]_  | \new_[645]_ ;
  assign \new_[8231]_  = \new_[646]_  | \new_[8230]_ ;
  assign \new_[8235]_  = \new_[641]_  | \new_[642]_ ;
  assign \new_[8236]_  = \new_[643]_  | \new_[8235]_ ;
  assign \new_[8237]_  = \new_[8236]_  | \new_[8231]_ ;
  assign \new_[8241]_  = \new_[638]_  | \new_[639]_ ;
  assign \new_[8242]_  = \new_[640]_  | \new_[8241]_ ;
  assign \new_[8246]_  = \new_[635]_  | \new_[636]_ ;
  assign \new_[8247]_  = \new_[637]_  | \new_[8246]_ ;
  assign \new_[8248]_  = \new_[8247]_  | \new_[8242]_ ;
  assign \new_[8249]_  = \new_[8248]_  | \new_[8237]_ ;
  assign \new_[8253]_  = \new_[632]_  | \new_[633]_ ;
  assign \new_[8254]_  = \new_[634]_  | \new_[8253]_ ;
  assign \new_[8258]_  = \new_[629]_  | \new_[630]_ ;
  assign \new_[8259]_  = \new_[631]_  | \new_[8258]_ ;
  assign \new_[8260]_  = \new_[8259]_  | \new_[8254]_ ;
  assign \new_[8264]_  = \new_[626]_  | \new_[627]_ ;
  assign \new_[8265]_  = \new_[628]_  | \new_[8264]_ ;
  assign \new_[8268]_  = \new_[624]_  | \new_[625]_ ;
  assign \new_[8271]_  = \new_[622]_  | \new_[623]_ ;
  assign \new_[8272]_  = \new_[8271]_  | \new_[8268]_ ;
  assign \new_[8273]_  = \new_[8272]_  | \new_[8265]_ ;
  assign \new_[8274]_  = \new_[8273]_  | \new_[8260]_ ;
  assign \new_[8275]_  = \new_[8274]_  | \new_[8249]_ ;
  assign \new_[8279]_  = \new_[619]_  | \new_[620]_ ;
  assign \new_[8280]_  = \new_[621]_  | \new_[8279]_ ;
  assign \new_[8284]_  = \new_[616]_  | \new_[617]_ ;
  assign \new_[8285]_  = \new_[618]_  | \new_[8284]_ ;
  assign \new_[8286]_  = \new_[8285]_  | \new_[8280]_ ;
  assign \new_[8290]_  = \new_[613]_  | \new_[614]_ ;
  assign \new_[8291]_  = \new_[615]_  | \new_[8290]_ ;
  assign \new_[8295]_  = \new_[610]_  | \new_[611]_ ;
  assign \new_[8296]_  = \new_[612]_  | \new_[8295]_ ;
  assign \new_[8297]_  = \new_[8296]_  | \new_[8291]_ ;
  assign \new_[8298]_  = \new_[8297]_  | \new_[8286]_ ;
  assign \new_[8302]_  = \new_[607]_  | \new_[608]_ ;
  assign \new_[8303]_  = \new_[609]_  | \new_[8302]_ ;
  assign \new_[8307]_  = \new_[604]_  | \new_[605]_ ;
  assign \new_[8308]_  = \new_[606]_  | \new_[8307]_ ;
  assign \new_[8309]_  = \new_[8308]_  | \new_[8303]_ ;
  assign \new_[8313]_  = \new_[601]_  | \new_[602]_ ;
  assign \new_[8314]_  = \new_[603]_  | \new_[8313]_ ;
  assign \new_[8317]_  = \new_[599]_  | \new_[600]_ ;
  assign \new_[8320]_  = \new_[597]_  | \new_[598]_ ;
  assign \new_[8321]_  = \new_[8320]_  | \new_[8317]_ ;
  assign \new_[8322]_  = \new_[8321]_  | \new_[8314]_ ;
  assign \new_[8323]_  = \new_[8322]_  | \new_[8309]_ ;
  assign \new_[8324]_  = \new_[8323]_  | \new_[8298]_ ;
  assign \new_[8325]_  = \new_[8324]_  | \new_[8275]_ ;
  assign \new_[8326]_  = \new_[8325]_  | \new_[8226]_ ;
  assign \new_[8327]_  = \new_[8326]_  | \new_[8129]_ ;
  assign \new_[8331]_  = \new_[594]_  | \new_[595]_ ;
  assign \new_[8332]_  = \new_[596]_  | \new_[8331]_ ;
  assign \new_[8336]_  = \new_[591]_  | \new_[592]_ ;
  assign \new_[8337]_  = \new_[593]_  | \new_[8336]_ ;
  assign \new_[8338]_  = \new_[8337]_  | \new_[8332]_ ;
  assign \new_[8342]_  = \new_[588]_  | \new_[589]_ ;
  assign \new_[8343]_  = \new_[590]_  | \new_[8342]_ ;
  assign \new_[8347]_  = \new_[585]_  | \new_[586]_ ;
  assign \new_[8348]_  = \new_[587]_  | \new_[8347]_ ;
  assign \new_[8349]_  = \new_[8348]_  | \new_[8343]_ ;
  assign \new_[8350]_  = \new_[8349]_  | \new_[8338]_ ;
  assign \new_[8354]_  = \new_[582]_  | \new_[583]_ ;
  assign \new_[8355]_  = \new_[584]_  | \new_[8354]_ ;
  assign \new_[8359]_  = \new_[579]_  | \new_[580]_ ;
  assign \new_[8360]_  = \new_[581]_  | \new_[8359]_ ;
  assign \new_[8361]_  = \new_[8360]_  | \new_[8355]_ ;
  assign \new_[8365]_  = \new_[576]_  | \new_[577]_ ;
  assign \new_[8366]_  = \new_[578]_  | \new_[8365]_ ;
  assign \new_[8370]_  = \new_[573]_  | \new_[574]_ ;
  assign \new_[8371]_  = \new_[575]_  | \new_[8370]_ ;
  assign \new_[8372]_  = \new_[8371]_  | \new_[8366]_ ;
  assign \new_[8373]_  = \new_[8372]_  | \new_[8361]_ ;
  assign \new_[8374]_  = \new_[8373]_  | \new_[8350]_ ;
  assign \new_[8378]_  = \new_[570]_  | \new_[571]_ ;
  assign \new_[8379]_  = \new_[572]_  | \new_[8378]_ ;
  assign \new_[8383]_  = \new_[567]_  | \new_[568]_ ;
  assign \new_[8384]_  = \new_[569]_  | \new_[8383]_ ;
  assign \new_[8385]_  = \new_[8384]_  | \new_[8379]_ ;
  assign \new_[8389]_  = \new_[564]_  | \new_[565]_ ;
  assign \new_[8390]_  = \new_[566]_  | \new_[8389]_ ;
  assign \new_[8394]_  = \new_[561]_  | \new_[562]_ ;
  assign \new_[8395]_  = \new_[563]_  | \new_[8394]_ ;
  assign \new_[8396]_  = \new_[8395]_  | \new_[8390]_ ;
  assign \new_[8397]_  = \new_[8396]_  | \new_[8385]_ ;
  assign \new_[8401]_  = \new_[558]_  | \new_[559]_ ;
  assign \new_[8402]_  = \new_[560]_  | \new_[8401]_ ;
  assign \new_[8406]_  = \new_[555]_  | \new_[556]_ ;
  assign \new_[8407]_  = \new_[557]_  | \new_[8406]_ ;
  assign \new_[8408]_  = \new_[8407]_  | \new_[8402]_ ;
  assign \new_[8412]_  = \new_[552]_  | \new_[553]_ ;
  assign \new_[8413]_  = \new_[554]_  | \new_[8412]_ ;
  assign \new_[8416]_  = \new_[550]_  | \new_[551]_ ;
  assign \new_[8419]_  = \new_[548]_  | \new_[549]_ ;
  assign \new_[8420]_  = \new_[8419]_  | \new_[8416]_ ;
  assign \new_[8421]_  = \new_[8420]_  | \new_[8413]_ ;
  assign \new_[8422]_  = \new_[8421]_  | \new_[8408]_ ;
  assign \new_[8423]_  = \new_[8422]_  | \new_[8397]_ ;
  assign \new_[8424]_  = \new_[8423]_  | \new_[8374]_ ;
  assign \new_[8428]_  = \new_[545]_  | \new_[546]_ ;
  assign \new_[8429]_  = \new_[547]_  | \new_[8428]_ ;
  assign \new_[8433]_  = \new_[542]_  | \new_[543]_ ;
  assign \new_[8434]_  = \new_[544]_  | \new_[8433]_ ;
  assign \new_[8435]_  = \new_[8434]_  | \new_[8429]_ ;
  assign \new_[8439]_  = \new_[539]_  | \new_[540]_ ;
  assign \new_[8440]_  = \new_[541]_  | \new_[8439]_ ;
  assign \new_[8444]_  = \new_[536]_  | \new_[537]_ ;
  assign \new_[8445]_  = \new_[538]_  | \new_[8444]_ ;
  assign \new_[8446]_  = \new_[8445]_  | \new_[8440]_ ;
  assign \new_[8447]_  = \new_[8446]_  | \new_[8435]_ ;
  assign \new_[8451]_  = \new_[533]_  | \new_[534]_ ;
  assign \new_[8452]_  = \new_[535]_  | \new_[8451]_ ;
  assign \new_[8456]_  = \new_[530]_  | \new_[531]_ ;
  assign \new_[8457]_  = \new_[532]_  | \new_[8456]_ ;
  assign \new_[8458]_  = \new_[8457]_  | \new_[8452]_ ;
  assign \new_[8462]_  = \new_[527]_  | \new_[528]_ ;
  assign \new_[8463]_  = \new_[529]_  | \new_[8462]_ ;
  assign \new_[8466]_  = \new_[525]_  | \new_[526]_ ;
  assign \new_[8469]_  = \new_[523]_  | \new_[524]_ ;
  assign \new_[8470]_  = \new_[8469]_  | \new_[8466]_ ;
  assign \new_[8471]_  = \new_[8470]_  | \new_[8463]_ ;
  assign \new_[8472]_  = \new_[8471]_  | \new_[8458]_ ;
  assign \new_[8473]_  = \new_[8472]_  | \new_[8447]_ ;
  assign \new_[8477]_  = \new_[520]_  | \new_[521]_ ;
  assign \new_[8478]_  = \new_[522]_  | \new_[8477]_ ;
  assign \new_[8482]_  = \new_[517]_  | \new_[518]_ ;
  assign \new_[8483]_  = \new_[519]_  | \new_[8482]_ ;
  assign \new_[8484]_  = \new_[8483]_  | \new_[8478]_ ;
  assign \new_[8488]_  = \new_[514]_  | \new_[515]_ ;
  assign \new_[8489]_  = \new_[516]_  | \new_[8488]_ ;
  assign \new_[8493]_  = \new_[511]_  | \new_[512]_ ;
  assign \new_[8494]_  = \new_[513]_  | \new_[8493]_ ;
  assign \new_[8495]_  = \new_[8494]_  | \new_[8489]_ ;
  assign \new_[8496]_  = \new_[8495]_  | \new_[8484]_ ;
  assign \new_[8500]_  = \new_[508]_  | \new_[509]_ ;
  assign \new_[8501]_  = \new_[510]_  | \new_[8500]_ ;
  assign \new_[8505]_  = \new_[505]_  | \new_[506]_ ;
  assign \new_[8506]_  = \new_[507]_  | \new_[8505]_ ;
  assign \new_[8507]_  = \new_[8506]_  | \new_[8501]_ ;
  assign \new_[8511]_  = \new_[502]_  | \new_[503]_ ;
  assign \new_[8512]_  = \new_[504]_  | \new_[8511]_ ;
  assign \new_[8515]_  = \new_[500]_  | \new_[501]_ ;
  assign \new_[8518]_  = \new_[498]_  | \new_[499]_ ;
  assign \new_[8519]_  = \new_[8518]_  | \new_[8515]_ ;
  assign \new_[8520]_  = \new_[8519]_  | \new_[8512]_ ;
  assign \new_[8521]_  = \new_[8520]_  | \new_[8507]_ ;
  assign \new_[8522]_  = \new_[8521]_  | \new_[8496]_ ;
  assign \new_[8523]_  = \new_[8522]_  | \new_[8473]_ ;
  assign \new_[8524]_  = \new_[8523]_  | \new_[8424]_ ;
  assign \new_[8528]_  = \new_[495]_  | \new_[496]_ ;
  assign \new_[8529]_  = \new_[497]_  | \new_[8528]_ ;
  assign \new_[8533]_  = \new_[492]_  | \new_[493]_ ;
  assign \new_[8534]_  = \new_[494]_  | \new_[8533]_ ;
  assign \new_[8535]_  = \new_[8534]_  | \new_[8529]_ ;
  assign \new_[8539]_  = \new_[489]_  | \new_[490]_ ;
  assign \new_[8540]_  = \new_[491]_  | \new_[8539]_ ;
  assign \new_[8544]_  = \new_[486]_  | \new_[487]_ ;
  assign \new_[8545]_  = \new_[488]_  | \new_[8544]_ ;
  assign \new_[8546]_  = \new_[8545]_  | \new_[8540]_ ;
  assign \new_[8547]_  = \new_[8546]_  | \new_[8535]_ ;
  assign \new_[8551]_  = \new_[483]_  | \new_[484]_ ;
  assign \new_[8552]_  = \new_[485]_  | \new_[8551]_ ;
  assign \new_[8556]_  = \new_[480]_  | \new_[481]_ ;
  assign \new_[8557]_  = \new_[482]_  | \new_[8556]_ ;
  assign \new_[8558]_  = \new_[8557]_  | \new_[8552]_ ;
  assign \new_[8562]_  = \new_[477]_  | \new_[478]_ ;
  assign \new_[8563]_  = \new_[479]_  | \new_[8562]_ ;
  assign \new_[8566]_  = \new_[475]_  | \new_[476]_ ;
  assign \new_[8569]_  = \new_[473]_  | \new_[474]_ ;
  assign \new_[8570]_  = \new_[8569]_  | \new_[8566]_ ;
  assign \new_[8571]_  = \new_[8570]_  | \new_[8563]_ ;
  assign \new_[8572]_  = \new_[8571]_  | \new_[8558]_ ;
  assign \new_[8573]_  = \new_[8572]_  | \new_[8547]_ ;
  assign \new_[8577]_  = \new_[470]_  | \new_[471]_ ;
  assign \new_[8578]_  = \new_[472]_  | \new_[8577]_ ;
  assign \new_[8582]_  = \new_[467]_  | \new_[468]_ ;
  assign \new_[8583]_  = \new_[469]_  | \new_[8582]_ ;
  assign \new_[8584]_  = \new_[8583]_  | \new_[8578]_ ;
  assign \new_[8588]_  = \new_[464]_  | \new_[465]_ ;
  assign \new_[8589]_  = \new_[466]_  | \new_[8588]_ ;
  assign \new_[8593]_  = \new_[461]_  | \new_[462]_ ;
  assign \new_[8594]_  = \new_[463]_  | \new_[8593]_ ;
  assign \new_[8595]_  = \new_[8594]_  | \new_[8589]_ ;
  assign \new_[8596]_  = \new_[8595]_  | \new_[8584]_ ;
  assign \new_[8600]_  = \new_[458]_  | \new_[459]_ ;
  assign \new_[8601]_  = \new_[460]_  | \new_[8600]_ ;
  assign \new_[8605]_  = \new_[455]_  | \new_[456]_ ;
  assign \new_[8606]_  = \new_[457]_  | \new_[8605]_ ;
  assign \new_[8607]_  = \new_[8606]_  | \new_[8601]_ ;
  assign \new_[8611]_  = \new_[452]_  | \new_[453]_ ;
  assign \new_[8612]_  = \new_[454]_  | \new_[8611]_ ;
  assign \new_[8615]_  = \new_[450]_  | \new_[451]_ ;
  assign \new_[8618]_  = \new_[448]_  | \new_[449]_ ;
  assign \new_[8619]_  = \new_[8618]_  | \new_[8615]_ ;
  assign \new_[8620]_  = \new_[8619]_  | \new_[8612]_ ;
  assign \new_[8621]_  = \new_[8620]_  | \new_[8607]_ ;
  assign \new_[8622]_  = \new_[8621]_  | \new_[8596]_ ;
  assign \new_[8623]_  = \new_[8622]_  | \new_[8573]_ ;
  assign \new_[8627]_  = \new_[445]_  | \new_[446]_ ;
  assign \new_[8628]_  = \new_[447]_  | \new_[8627]_ ;
  assign \new_[8632]_  = \new_[442]_  | \new_[443]_ ;
  assign \new_[8633]_  = \new_[444]_  | \new_[8632]_ ;
  assign \new_[8634]_  = \new_[8633]_  | \new_[8628]_ ;
  assign \new_[8638]_  = \new_[439]_  | \new_[440]_ ;
  assign \new_[8639]_  = \new_[441]_  | \new_[8638]_ ;
  assign \new_[8643]_  = \new_[436]_  | \new_[437]_ ;
  assign \new_[8644]_  = \new_[438]_  | \new_[8643]_ ;
  assign \new_[8645]_  = \new_[8644]_  | \new_[8639]_ ;
  assign \new_[8646]_  = \new_[8645]_  | \new_[8634]_ ;
  assign \new_[8650]_  = \new_[433]_  | \new_[434]_ ;
  assign \new_[8651]_  = \new_[435]_  | \new_[8650]_ ;
  assign \new_[8655]_  = \new_[430]_  | \new_[431]_ ;
  assign \new_[8656]_  = \new_[432]_  | \new_[8655]_ ;
  assign \new_[8657]_  = \new_[8656]_  | \new_[8651]_ ;
  assign \new_[8661]_  = \new_[427]_  | \new_[428]_ ;
  assign \new_[8662]_  = \new_[429]_  | \new_[8661]_ ;
  assign \new_[8665]_  = \new_[425]_  | \new_[426]_ ;
  assign \new_[8668]_  = \new_[423]_  | \new_[424]_ ;
  assign \new_[8669]_  = \new_[8668]_  | \new_[8665]_ ;
  assign \new_[8670]_  = \new_[8669]_  | \new_[8662]_ ;
  assign \new_[8671]_  = \new_[8670]_  | \new_[8657]_ ;
  assign \new_[8672]_  = \new_[8671]_  | \new_[8646]_ ;
  assign \new_[8676]_  = \new_[420]_  | \new_[421]_ ;
  assign \new_[8677]_  = \new_[422]_  | \new_[8676]_ ;
  assign \new_[8681]_  = \new_[417]_  | \new_[418]_ ;
  assign \new_[8682]_  = \new_[419]_  | \new_[8681]_ ;
  assign \new_[8683]_  = \new_[8682]_  | \new_[8677]_ ;
  assign \new_[8687]_  = \new_[414]_  | \new_[415]_ ;
  assign \new_[8688]_  = \new_[416]_  | \new_[8687]_ ;
  assign \new_[8692]_  = \new_[411]_  | \new_[412]_ ;
  assign \new_[8693]_  = \new_[413]_  | \new_[8692]_ ;
  assign \new_[8694]_  = \new_[8693]_  | \new_[8688]_ ;
  assign \new_[8695]_  = \new_[8694]_  | \new_[8683]_ ;
  assign \new_[8699]_  = \new_[408]_  | \new_[409]_ ;
  assign \new_[8700]_  = \new_[410]_  | \new_[8699]_ ;
  assign \new_[8704]_  = \new_[405]_  | \new_[406]_ ;
  assign \new_[8705]_  = \new_[407]_  | \new_[8704]_ ;
  assign \new_[8706]_  = \new_[8705]_  | \new_[8700]_ ;
  assign \new_[8710]_  = \new_[402]_  | \new_[403]_ ;
  assign \new_[8711]_  = \new_[404]_  | \new_[8710]_ ;
  assign \new_[8714]_  = \new_[400]_  | \new_[401]_ ;
  assign \new_[8717]_  = \new_[398]_  | \new_[399]_ ;
  assign \new_[8718]_  = \new_[8717]_  | \new_[8714]_ ;
  assign \new_[8719]_  = \new_[8718]_  | \new_[8711]_ ;
  assign \new_[8720]_  = \new_[8719]_  | \new_[8706]_ ;
  assign \new_[8721]_  = \new_[8720]_  | \new_[8695]_ ;
  assign \new_[8722]_  = \new_[8721]_  | \new_[8672]_ ;
  assign \new_[8723]_  = \new_[8722]_  | \new_[8623]_ ;
  assign \new_[8724]_  = \new_[8723]_  | \new_[8524]_ ;
  assign \new_[8725]_  = \new_[8724]_  | \new_[8327]_ ;
  assign \new_[8729]_  = \new_[395]_  | \new_[396]_ ;
  assign \new_[8730]_  = \new_[397]_  | \new_[8729]_ ;
  assign \new_[8734]_  = \new_[392]_  | \new_[393]_ ;
  assign \new_[8735]_  = \new_[394]_  | \new_[8734]_ ;
  assign \new_[8736]_  = \new_[8735]_  | \new_[8730]_ ;
  assign \new_[8740]_  = \new_[389]_  | \new_[390]_ ;
  assign \new_[8741]_  = \new_[391]_  | \new_[8740]_ ;
  assign \new_[8745]_  = \new_[386]_  | \new_[387]_ ;
  assign \new_[8746]_  = \new_[388]_  | \new_[8745]_ ;
  assign \new_[8747]_  = \new_[8746]_  | \new_[8741]_ ;
  assign \new_[8748]_  = \new_[8747]_  | \new_[8736]_ ;
  assign \new_[8752]_  = \new_[383]_  | \new_[384]_ ;
  assign \new_[8753]_  = \new_[385]_  | \new_[8752]_ ;
  assign \new_[8757]_  = \new_[380]_  | \new_[381]_ ;
  assign \new_[8758]_  = \new_[382]_  | \new_[8757]_ ;
  assign \new_[8759]_  = \new_[8758]_  | \new_[8753]_ ;
  assign \new_[8763]_  = \new_[377]_  | \new_[378]_ ;
  assign \new_[8764]_  = \new_[379]_  | \new_[8763]_ ;
  assign \new_[8768]_  = \new_[374]_  | \new_[375]_ ;
  assign \new_[8769]_  = \new_[376]_  | \new_[8768]_ ;
  assign \new_[8770]_  = \new_[8769]_  | \new_[8764]_ ;
  assign \new_[8771]_  = \new_[8770]_  | \new_[8759]_ ;
  assign \new_[8772]_  = \new_[8771]_  | \new_[8748]_ ;
  assign \new_[8776]_  = \new_[371]_  | \new_[372]_ ;
  assign \new_[8777]_  = \new_[373]_  | \new_[8776]_ ;
  assign \new_[8781]_  = \new_[368]_  | \new_[369]_ ;
  assign \new_[8782]_  = \new_[370]_  | \new_[8781]_ ;
  assign \new_[8783]_  = \new_[8782]_  | \new_[8777]_ ;
  assign \new_[8787]_  = \new_[365]_  | \new_[366]_ ;
  assign \new_[8788]_  = \new_[367]_  | \new_[8787]_ ;
  assign \new_[8792]_  = \new_[362]_  | \new_[363]_ ;
  assign \new_[8793]_  = \new_[364]_  | \new_[8792]_ ;
  assign \new_[8794]_  = \new_[8793]_  | \new_[8788]_ ;
  assign \new_[8795]_  = \new_[8794]_  | \new_[8783]_ ;
  assign \new_[8799]_  = \new_[359]_  | \new_[360]_ ;
  assign \new_[8800]_  = \new_[361]_  | \new_[8799]_ ;
  assign \new_[8804]_  = \new_[356]_  | \new_[357]_ ;
  assign \new_[8805]_  = \new_[358]_  | \new_[8804]_ ;
  assign \new_[8806]_  = \new_[8805]_  | \new_[8800]_ ;
  assign \new_[8810]_  = \new_[353]_  | \new_[354]_ ;
  assign \new_[8811]_  = \new_[355]_  | \new_[8810]_ ;
  assign \new_[8814]_  = \new_[351]_  | \new_[352]_ ;
  assign \new_[8817]_  = \new_[349]_  | \new_[350]_ ;
  assign \new_[8818]_  = \new_[8817]_  | \new_[8814]_ ;
  assign \new_[8819]_  = \new_[8818]_  | \new_[8811]_ ;
  assign \new_[8820]_  = \new_[8819]_  | \new_[8806]_ ;
  assign \new_[8821]_  = \new_[8820]_  | \new_[8795]_ ;
  assign \new_[8822]_  = \new_[8821]_  | \new_[8772]_ ;
  assign \new_[8826]_  = \new_[346]_  | \new_[347]_ ;
  assign \new_[8827]_  = \new_[348]_  | \new_[8826]_ ;
  assign \new_[8831]_  = \new_[343]_  | \new_[344]_ ;
  assign \new_[8832]_  = \new_[345]_  | \new_[8831]_ ;
  assign \new_[8833]_  = \new_[8832]_  | \new_[8827]_ ;
  assign \new_[8837]_  = \new_[340]_  | \new_[341]_ ;
  assign \new_[8838]_  = \new_[342]_  | \new_[8837]_ ;
  assign \new_[8842]_  = \new_[337]_  | \new_[338]_ ;
  assign \new_[8843]_  = \new_[339]_  | \new_[8842]_ ;
  assign \new_[8844]_  = \new_[8843]_  | \new_[8838]_ ;
  assign \new_[8845]_  = \new_[8844]_  | \new_[8833]_ ;
  assign \new_[8849]_  = \new_[334]_  | \new_[335]_ ;
  assign \new_[8850]_  = \new_[336]_  | \new_[8849]_ ;
  assign \new_[8854]_  = \new_[331]_  | \new_[332]_ ;
  assign \new_[8855]_  = \new_[333]_  | \new_[8854]_ ;
  assign \new_[8856]_  = \new_[8855]_  | \new_[8850]_ ;
  assign \new_[8860]_  = \new_[328]_  | \new_[329]_ ;
  assign \new_[8861]_  = \new_[330]_  | \new_[8860]_ ;
  assign \new_[8864]_  = \new_[326]_  | \new_[327]_ ;
  assign \new_[8867]_  = \new_[324]_  | \new_[325]_ ;
  assign \new_[8868]_  = \new_[8867]_  | \new_[8864]_ ;
  assign \new_[8869]_  = \new_[8868]_  | \new_[8861]_ ;
  assign \new_[8870]_  = \new_[8869]_  | \new_[8856]_ ;
  assign \new_[8871]_  = \new_[8870]_  | \new_[8845]_ ;
  assign \new_[8875]_  = \new_[321]_  | \new_[322]_ ;
  assign \new_[8876]_  = \new_[323]_  | \new_[8875]_ ;
  assign \new_[8880]_  = \new_[318]_  | \new_[319]_ ;
  assign \new_[8881]_  = \new_[320]_  | \new_[8880]_ ;
  assign \new_[8882]_  = \new_[8881]_  | \new_[8876]_ ;
  assign \new_[8886]_  = \new_[315]_  | \new_[316]_ ;
  assign \new_[8887]_  = \new_[317]_  | \new_[8886]_ ;
  assign \new_[8891]_  = \new_[312]_  | \new_[313]_ ;
  assign \new_[8892]_  = \new_[314]_  | \new_[8891]_ ;
  assign \new_[8893]_  = \new_[8892]_  | \new_[8887]_ ;
  assign \new_[8894]_  = \new_[8893]_  | \new_[8882]_ ;
  assign \new_[8898]_  = \new_[309]_  | \new_[310]_ ;
  assign \new_[8899]_  = \new_[311]_  | \new_[8898]_ ;
  assign \new_[8903]_  = \new_[306]_  | \new_[307]_ ;
  assign \new_[8904]_  = \new_[308]_  | \new_[8903]_ ;
  assign \new_[8905]_  = \new_[8904]_  | \new_[8899]_ ;
  assign \new_[8909]_  = \new_[303]_  | \new_[304]_ ;
  assign \new_[8910]_  = \new_[305]_  | \new_[8909]_ ;
  assign \new_[8913]_  = \new_[301]_  | \new_[302]_ ;
  assign \new_[8916]_  = \new_[299]_  | \new_[300]_ ;
  assign \new_[8917]_  = \new_[8916]_  | \new_[8913]_ ;
  assign \new_[8918]_  = \new_[8917]_  | \new_[8910]_ ;
  assign \new_[8919]_  = \new_[8918]_  | \new_[8905]_ ;
  assign \new_[8920]_  = \new_[8919]_  | \new_[8894]_ ;
  assign \new_[8921]_  = \new_[8920]_  | \new_[8871]_ ;
  assign \new_[8922]_  = \new_[8921]_  | \new_[8822]_ ;
  assign \new_[8926]_  = \new_[296]_  | \new_[297]_ ;
  assign \new_[8927]_  = \new_[298]_  | \new_[8926]_ ;
  assign \new_[8931]_  = \new_[293]_  | \new_[294]_ ;
  assign \new_[8932]_  = \new_[295]_  | \new_[8931]_ ;
  assign \new_[8933]_  = \new_[8932]_  | \new_[8927]_ ;
  assign \new_[8937]_  = \new_[290]_  | \new_[291]_ ;
  assign \new_[8938]_  = \new_[292]_  | \new_[8937]_ ;
  assign \new_[8942]_  = \new_[287]_  | \new_[288]_ ;
  assign \new_[8943]_  = \new_[289]_  | \new_[8942]_ ;
  assign \new_[8944]_  = \new_[8943]_  | \new_[8938]_ ;
  assign \new_[8945]_  = \new_[8944]_  | \new_[8933]_ ;
  assign \new_[8949]_  = \new_[284]_  | \new_[285]_ ;
  assign \new_[8950]_  = \new_[286]_  | \new_[8949]_ ;
  assign \new_[8954]_  = \new_[281]_  | \new_[282]_ ;
  assign \new_[8955]_  = \new_[283]_  | \new_[8954]_ ;
  assign \new_[8956]_  = \new_[8955]_  | \new_[8950]_ ;
  assign \new_[8960]_  = \new_[278]_  | \new_[279]_ ;
  assign \new_[8961]_  = \new_[280]_  | \new_[8960]_ ;
  assign \new_[8965]_  = \new_[275]_  | \new_[276]_ ;
  assign \new_[8966]_  = \new_[277]_  | \new_[8965]_ ;
  assign \new_[8967]_  = \new_[8966]_  | \new_[8961]_ ;
  assign \new_[8968]_  = \new_[8967]_  | \new_[8956]_ ;
  assign \new_[8969]_  = \new_[8968]_  | \new_[8945]_ ;
  assign \new_[8973]_  = \new_[272]_  | \new_[273]_ ;
  assign \new_[8974]_  = \new_[274]_  | \new_[8973]_ ;
  assign \new_[8978]_  = \new_[269]_  | \new_[270]_ ;
  assign \new_[8979]_  = \new_[271]_  | \new_[8978]_ ;
  assign \new_[8980]_  = \new_[8979]_  | \new_[8974]_ ;
  assign \new_[8984]_  = \new_[266]_  | \new_[267]_ ;
  assign \new_[8985]_  = \new_[268]_  | \new_[8984]_ ;
  assign \new_[8989]_  = \new_[263]_  | \new_[264]_ ;
  assign \new_[8990]_  = \new_[265]_  | \new_[8989]_ ;
  assign \new_[8991]_  = \new_[8990]_  | \new_[8985]_ ;
  assign \new_[8992]_  = \new_[8991]_  | \new_[8980]_ ;
  assign \new_[8996]_  = \new_[260]_  | \new_[261]_ ;
  assign \new_[8997]_  = \new_[262]_  | \new_[8996]_ ;
  assign \new_[9001]_  = \new_[257]_  | \new_[258]_ ;
  assign \new_[9002]_  = \new_[259]_  | \new_[9001]_ ;
  assign \new_[9003]_  = \new_[9002]_  | \new_[8997]_ ;
  assign \new_[9007]_  = \new_[254]_  | \new_[255]_ ;
  assign \new_[9008]_  = \new_[256]_  | \new_[9007]_ ;
  assign \new_[9011]_  = \new_[252]_  | \new_[253]_ ;
  assign \new_[9014]_  = \new_[250]_  | \new_[251]_ ;
  assign \new_[9015]_  = \new_[9014]_  | \new_[9011]_ ;
  assign \new_[9016]_  = \new_[9015]_  | \new_[9008]_ ;
  assign \new_[9017]_  = \new_[9016]_  | \new_[9003]_ ;
  assign \new_[9018]_  = \new_[9017]_  | \new_[8992]_ ;
  assign \new_[9019]_  = \new_[9018]_  | \new_[8969]_ ;
  assign \new_[9023]_  = \new_[247]_  | \new_[248]_ ;
  assign \new_[9024]_  = \new_[249]_  | \new_[9023]_ ;
  assign \new_[9028]_  = \new_[244]_  | \new_[245]_ ;
  assign \new_[9029]_  = \new_[246]_  | \new_[9028]_ ;
  assign \new_[9030]_  = \new_[9029]_  | \new_[9024]_ ;
  assign \new_[9034]_  = \new_[241]_  | \new_[242]_ ;
  assign \new_[9035]_  = \new_[243]_  | \new_[9034]_ ;
  assign \new_[9039]_  = \new_[238]_  | \new_[239]_ ;
  assign \new_[9040]_  = \new_[240]_  | \new_[9039]_ ;
  assign \new_[9041]_  = \new_[9040]_  | \new_[9035]_ ;
  assign \new_[9042]_  = \new_[9041]_  | \new_[9030]_ ;
  assign \new_[9046]_  = \new_[235]_  | \new_[236]_ ;
  assign \new_[9047]_  = \new_[237]_  | \new_[9046]_ ;
  assign \new_[9051]_  = \new_[232]_  | \new_[233]_ ;
  assign \new_[9052]_  = \new_[234]_  | \new_[9051]_ ;
  assign \new_[9053]_  = \new_[9052]_  | \new_[9047]_ ;
  assign \new_[9057]_  = \new_[229]_  | \new_[230]_ ;
  assign \new_[9058]_  = \new_[231]_  | \new_[9057]_ ;
  assign \new_[9061]_  = \new_[227]_  | \new_[228]_ ;
  assign \new_[9064]_  = \new_[225]_  | \new_[226]_ ;
  assign \new_[9065]_  = \new_[9064]_  | \new_[9061]_ ;
  assign \new_[9066]_  = \new_[9065]_  | \new_[9058]_ ;
  assign \new_[9067]_  = \new_[9066]_  | \new_[9053]_ ;
  assign \new_[9068]_  = \new_[9067]_  | \new_[9042]_ ;
  assign \new_[9072]_  = \new_[222]_  | \new_[223]_ ;
  assign \new_[9073]_  = \new_[224]_  | \new_[9072]_ ;
  assign \new_[9077]_  = \new_[219]_  | \new_[220]_ ;
  assign \new_[9078]_  = \new_[221]_  | \new_[9077]_ ;
  assign \new_[9079]_  = \new_[9078]_  | \new_[9073]_ ;
  assign \new_[9083]_  = \new_[216]_  | \new_[217]_ ;
  assign \new_[9084]_  = \new_[218]_  | \new_[9083]_ ;
  assign \new_[9088]_  = \new_[213]_  | \new_[214]_ ;
  assign \new_[9089]_  = \new_[215]_  | \new_[9088]_ ;
  assign \new_[9090]_  = \new_[9089]_  | \new_[9084]_ ;
  assign \new_[9091]_  = \new_[9090]_  | \new_[9079]_ ;
  assign \new_[9095]_  = \new_[210]_  | \new_[211]_ ;
  assign \new_[9096]_  = \new_[212]_  | \new_[9095]_ ;
  assign \new_[9100]_  = \new_[207]_  | \new_[208]_ ;
  assign \new_[9101]_  = \new_[209]_  | \new_[9100]_ ;
  assign \new_[9102]_  = \new_[9101]_  | \new_[9096]_ ;
  assign \new_[9106]_  = \new_[204]_  | \new_[205]_ ;
  assign \new_[9107]_  = \new_[206]_  | \new_[9106]_ ;
  assign \new_[9110]_  = \new_[202]_  | \new_[203]_ ;
  assign \new_[9113]_  = \new_[200]_  | \new_[201]_ ;
  assign \new_[9114]_  = \new_[9113]_  | \new_[9110]_ ;
  assign \new_[9115]_  = \new_[9114]_  | \new_[9107]_ ;
  assign \new_[9116]_  = \new_[9115]_  | \new_[9102]_ ;
  assign \new_[9117]_  = \new_[9116]_  | \new_[9091]_ ;
  assign \new_[9118]_  = \new_[9117]_  | \new_[9068]_ ;
  assign \new_[9119]_  = \new_[9118]_  | \new_[9019]_ ;
  assign \new_[9120]_  = \new_[9119]_  | \new_[8922]_ ;
  assign \new_[9124]_  = \new_[197]_  | \new_[198]_ ;
  assign \new_[9125]_  = \new_[199]_  | \new_[9124]_ ;
  assign \new_[9129]_  = \new_[194]_  | \new_[195]_ ;
  assign \new_[9130]_  = \new_[196]_  | \new_[9129]_ ;
  assign \new_[9131]_  = \new_[9130]_  | \new_[9125]_ ;
  assign \new_[9135]_  = \new_[191]_  | \new_[192]_ ;
  assign \new_[9136]_  = \new_[193]_  | \new_[9135]_ ;
  assign \new_[9140]_  = \new_[188]_  | \new_[189]_ ;
  assign \new_[9141]_  = \new_[190]_  | \new_[9140]_ ;
  assign \new_[9142]_  = \new_[9141]_  | \new_[9136]_ ;
  assign \new_[9143]_  = \new_[9142]_  | \new_[9131]_ ;
  assign \new_[9147]_  = \new_[185]_  | \new_[186]_ ;
  assign \new_[9148]_  = \new_[187]_  | \new_[9147]_ ;
  assign \new_[9152]_  = \new_[182]_  | \new_[183]_ ;
  assign \new_[9153]_  = \new_[184]_  | \new_[9152]_ ;
  assign \new_[9154]_  = \new_[9153]_  | \new_[9148]_ ;
  assign \new_[9158]_  = \new_[179]_  | \new_[180]_ ;
  assign \new_[9159]_  = \new_[181]_  | \new_[9158]_ ;
  assign \new_[9163]_  = \new_[176]_  | \new_[177]_ ;
  assign \new_[9164]_  = \new_[178]_  | \new_[9163]_ ;
  assign \new_[9165]_  = \new_[9164]_  | \new_[9159]_ ;
  assign \new_[9166]_  = \new_[9165]_  | \new_[9154]_ ;
  assign \new_[9167]_  = \new_[9166]_  | \new_[9143]_ ;
  assign \new_[9171]_  = \new_[173]_  | \new_[174]_ ;
  assign \new_[9172]_  = \new_[175]_  | \new_[9171]_ ;
  assign \new_[9176]_  = \new_[170]_  | \new_[171]_ ;
  assign \new_[9177]_  = \new_[172]_  | \new_[9176]_ ;
  assign \new_[9178]_  = \new_[9177]_  | \new_[9172]_ ;
  assign \new_[9182]_  = \new_[167]_  | \new_[168]_ ;
  assign \new_[9183]_  = \new_[169]_  | \new_[9182]_ ;
  assign \new_[9187]_  = \new_[164]_  | \new_[165]_ ;
  assign \new_[9188]_  = \new_[166]_  | \new_[9187]_ ;
  assign \new_[9189]_  = \new_[9188]_  | \new_[9183]_ ;
  assign \new_[9190]_  = \new_[9189]_  | \new_[9178]_ ;
  assign \new_[9194]_  = \new_[161]_  | \new_[162]_ ;
  assign \new_[9195]_  = \new_[163]_  | \new_[9194]_ ;
  assign \new_[9199]_  = \new_[158]_  | \new_[159]_ ;
  assign \new_[9200]_  = \new_[160]_  | \new_[9199]_ ;
  assign \new_[9201]_  = \new_[9200]_  | \new_[9195]_ ;
  assign \new_[9205]_  = \new_[155]_  | \new_[156]_ ;
  assign \new_[9206]_  = \new_[157]_  | \new_[9205]_ ;
  assign \new_[9209]_  = \new_[153]_  | \new_[154]_ ;
  assign \new_[9212]_  = \new_[151]_  | \new_[152]_ ;
  assign \new_[9213]_  = \new_[9212]_  | \new_[9209]_ ;
  assign \new_[9214]_  = \new_[9213]_  | \new_[9206]_ ;
  assign \new_[9215]_  = \new_[9214]_  | \new_[9201]_ ;
  assign \new_[9216]_  = \new_[9215]_  | \new_[9190]_ ;
  assign \new_[9217]_  = \new_[9216]_  | \new_[9167]_ ;
  assign \new_[9221]_  = \new_[148]_  | \new_[149]_ ;
  assign \new_[9222]_  = \new_[150]_  | \new_[9221]_ ;
  assign \new_[9226]_  = \new_[145]_  | \new_[146]_ ;
  assign \new_[9227]_  = \new_[147]_  | \new_[9226]_ ;
  assign \new_[9228]_  = \new_[9227]_  | \new_[9222]_ ;
  assign \new_[9232]_  = \new_[142]_  | \new_[143]_ ;
  assign \new_[9233]_  = \new_[144]_  | \new_[9232]_ ;
  assign \new_[9237]_  = \new_[139]_  | \new_[140]_ ;
  assign \new_[9238]_  = \new_[141]_  | \new_[9237]_ ;
  assign \new_[9239]_  = \new_[9238]_  | \new_[9233]_ ;
  assign \new_[9240]_  = \new_[9239]_  | \new_[9228]_ ;
  assign \new_[9244]_  = \new_[136]_  | \new_[137]_ ;
  assign \new_[9245]_  = \new_[138]_  | \new_[9244]_ ;
  assign \new_[9249]_  = \new_[133]_  | \new_[134]_ ;
  assign \new_[9250]_  = \new_[135]_  | \new_[9249]_ ;
  assign \new_[9251]_  = \new_[9250]_  | \new_[9245]_ ;
  assign \new_[9255]_  = \new_[130]_  | \new_[131]_ ;
  assign \new_[9256]_  = \new_[132]_  | \new_[9255]_ ;
  assign \new_[9259]_  = \new_[128]_  | \new_[129]_ ;
  assign \new_[9262]_  = \new_[126]_  | \new_[127]_ ;
  assign \new_[9263]_  = \new_[9262]_  | \new_[9259]_ ;
  assign \new_[9264]_  = \new_[9263]_  | \new_[9256]_ ;
  assign \new_[9265]_  = \new_[9264]_  | \new_[9251]_ ;
  assign \new_[9266]_  = \new_[9265]_  | \new_[9240]_ ;
  assign \new_[9270]_  = \new_[123]_  | \new_[124]_ ;
  assign \new_[9271]_  = \new_[125]_  | \new_[9270]_ ;
  assign \new_[9275]_  = \new_[120]_  | \new_[121]_ ;
  assign \new_[9276]_  = \new_[122]_  | \new_[9275]_ ;
  assign \new_[9277]_  = \new_[9276]_  | \new_[9271]_ ;
  assign \new_[9281]_  = \new_[117]_  | \new_[118]_ ;
  assign \new_[9282]_  = \new_[119]_  | \new_[9281]_ ;
  assign \new_[9286]_  = \new_[114]_  | \new_[115]_ ;
  assign \new_[9287]_  = \new_[116]_  | \new_[9286]_ ;
  assign \new_[9288]_  = \new_[9287]_  | \new_[9282]_ ;
  assign \new_[9289]_  = \new_[9288]_  | \new_[9277]_ ;
  assign \new_[9293]_  = \new_[111]_  | \new_[112]_ ;
  assign \new_[9294]_  = \new_[113]_  | \new_[9293]_ ;
  assign \new_[9298]_  = \new_[108]_  | \new_[109]_ ;
  assign \new_[9299]_  = \new_[110]_  | \new_[9298]_ ;
  assign \new_[9300]_  = \new_[9299]_  | \new_[9294]_ ;
  assign \new_[9304]_  = \new_[105]_  | \new_[106]_ ;
  assign \new_[9305]_  = \new_[107]_  | \new_[9304]_ ;
  assign \new_[9308]_  = \new_[103]_  | \new_[104]_ ;
  assign \new_[9311]_  = \new_[101]_  | \new_[102]_ ;
  assign \new_[9312]_  = \new_[9311]_  | \new_[9308]_ ;
  assign \new_[9313]_  = \new_[9312]_  | \new_[9305]_ ;
  assign \new_[9314]_  = \new_[9313]_  | \new_[9300]_ ;
  assign \new_[9315]_  = \new_[9314]_  | \new_[9289]_ ;
  assign \new_[9316]_  = \new_[9315]_  | \new_[9266]_ ;
  assign \new_[9317]_  = \new_[9316]_  | \new_[9217]_ ;
  assign \new_[9321]_  = \new_[98]_  | \new_[99]_ ;
  assign \new_[9322]_  = \new_[100]_  | \new_[9321]_ ;
  assign \new_[9326]_  = \new_[95]_  | \new_[96]_ ;
  assign \new_[9327]_  = \new_[97]_  | \new_[9326]_ ;
  assign \new_[9328]_  = \new_[9327]_  | \new_[9322]_ ;
  assign \new_[9332]_  = \new_[92]_  | \new_[93]_ ;
  assign \new_[9333]_  = \new_[94]_  | \new_[9332]_ ;
  assign \new_[9337]_  = \new_[89]_  | \new_[90]_ ;
  assign \new_[9338]_  = \new_[91]_  | \new_[9337]_ ;
  assign \new_[9339]_  = \new_[9338]_  | \new_[9333]_ ;
  assign \new_[9340]_  = \new_[9339]_  | \new_[9328]_ ;
  assign \new_[9344]_  = \new_[86]_  | \new_[87]_ ;
  assign \new_[9345]_  = \new_[88]_  | \new_[9344]_ ;
  assign \new_[9349]_  = \new_[83]_  | \new_[84]_ ;
  assign \new_[9350]_  = \new_[85]_  | \new_[9349]_ ;
  assign \new_[9351]_  = \new_[9350]_  | \new_[9345]_ ;
  assign \new_[9355]_  = \new_[80]_  | \new_[81]_ ;
  assign \new_[9356]_  = \new_[82]_  | \new_[9355]_ ;
  assign \new_[9359]_  = \new_[78]_  | \new_[79]_ ;
  assign \new_[9362]_  = \new_[76]_  | \new_[77]_ ;
  assign \new_[9363]_  = \new_[9362]_  | \new_[9359]_ ;
  assign \new_[9364]_  = \new_[9363]_  | \new_[9356]_ ;
  assign \new_[9365]_  = \new_[9364]_  | \new_[9351]_ ;
  assign \new_[9366]_  = \new_[9365]_  | \new_[9340]_ ;
  assign \new_[9370]_  = \new_[73]_  | \new_[74]_ ;
  assign \new_[9371]_  = \new_[75]_  | \new_[9370]_ ;
  assign \new_[9375]_  = \new_[70]_  | \new_[71]_ ;
  assign \new_[9376]_  = \new_[72]_  | \new_[9375]_ ;
  assign \new_[9377]_  = \new_[9376]_  | \new_[9371]_ ;
  assign \new_[9381]_  = \new_[67]_  | \new_[68]_ ;
  assign \new_[9382]_  = \new_[69]_  | \new_[9381]_ ;
  assign \new_[9386]_  = \new_[64]_  | \new_[65]_ ;
  assign \new_[9387]_  = \new_[66]_  | \new_[9386]_ ;
  assign \new_[9388]_  = \new_[9387]_  | \new_[9382]_ ;
  assign \new_[9389]_  = \new_[9388]_  | \new_[9377]_ ;
  assign \new_[9393]_  = \new_[61]_  | \new_[62]_ ;
  assign \new_[9394]_  = \new_[63]_  | \new_[9393]_ ;
  assign \new_[9398]_  = \new_[58]_  | \new_[59]_ ;
  assign \new_[9399]_  = \new_[60]_  | \new_[9398]_ ;
  assign \new_[9400]_  = \new_[9399]_  | \new_[9394]_ ;
  assign \new_[9404]_  = \new_[55]_  | \new_[56]_ ;
  assign \new_[9405]_  = \new_[57]_  | \new_[9404]_ ;
  assign \new_[9408]_  = \new_[53]_  | \new_[54]_ ;
  assign \new_[9411]_  = \new_[51]_  | \new_[52]_ ;
  assign \new_[9412]_  = \new_[9411]_  | \new_[9408]_ ;
  assign \new_[9413]_  = \new_[9412]_  | \new_[9405]_ ;
  assign \new_[9414]_  = \new_[9413]_  | \new_[9400]_ ;
  assign \new_[9415]_  = \new_[9414]_  | \new_[9389]_ ;
  assign \new_[9416]_  = \new_[9415]_  | \new_[9366]_ ;
  assign \new_[9420]_  = \new_[48]_  | \new_[49]_ ;
  assign \new_[9421]_  = \new_[50]_  | \new_[9420]_ ;
  assign \new_[9425]_  = \new_[45]_  | \new_[46]_ ;
  assign \new_[9426]_  = \new_[47]_  | \new_[9425]_ ;
  assign \new_[9427]_  = \new_[9426]_  | \new_[9421]_ ;
  assign \new_[9431]_  = \new_[42]_  | \new_[43]_ ;
  assign \new_[9432]_  = \new_[44]_  | \new_[9431]_ ;
  assign \new_[9436]_  = \new_[39]_  | \new_[40]_ ;
  assign \new_[9437]_  = \new_[41]_  | \new_[9436]_ ;
  assign \new_[9438]_  = \new_[9437]_  | \new_[9432]_ ;
  assign \new_[9439]_  = \new_[9438]_  | \new_[9427]_ ;
  assign \new_[9443]_  = \new_[36]_  | \new_[37]_ ;
  assign \new_[9444]_  = \new_[38]_  | \new_[9443]_ ;
  assign \new_[9448]_  = \new_[33]_  | \new_[34]_ ;
  assign \new_[9449]_  = \new_[35]_  | \new_[9448]_ ;
  assign \new_[9450]_  = \new_[9449]_  | \new_[9444]_ ;
  assign \new_[9454]_  = \new_[30]_  | \new_[31]_ ;
  assign \new_[9455]_  = \new_[32]_  | \new_[9454]_ ;
  assign \new_[9458]_  = \new_[28]_  | \new_[29]_ ;
  assign \new_[9461]_  = \new_[26]_  | \new_[27]_ ;
  assign \new_[9462]_  = \new_[9461]_  | \new_[9458]_ ;
  assign \new_[9463]_  = \new_[9462]_  | \new_[9455]_ ;
  assign \new_[9464]_  = \new_[9463]_  | \new_[9450]_ ;
  assign \new_[9465]_  = \new_[9464]_  | \new_[9439]_ ;
  assign \new_[9469]_  = \new_[23]_  | \new_[24]_ ;
  assign \new_[9470]_  = \new_[25]_  | \new_[9469]_ ;
  assign \new_[9474]_  = \new_[20]_  | \new_[21]_ ;
  assign \new_[9475]_  = \new_[22]_  | \new_[9474]_ ;
  assign \new_[9476]_  = \new_[9475]_  | \new_[9470]_ ;
  assign \new_[9480]_  = \new_[17]_  | \new_[18]_ ;
  assign \new_[9481]_  = \new_[19]_  | \new_[9480]_ ;
  assign \new_[9485]_  = \new_[14]_  | \new_[15]_ ;
  assign \new_[9486]_  = \new_[16]_  | \new_[9485]_ ;
  assign \new_[9487]_  = \new_[9486]_  | \new_[9481]_ ;
  assign \new_[9488]_  = \new_[9487]_  | \new_[9476]_ ;
  assign \new_[9492]_  = \new_[11]_  | \new_[12]_ ;
  assign \new_[9493]_  = \new_[13]_  | \new_[9492]_ ;
  assign \new_[9497]_  = \new_[8]_  | \new_[9]_ ;
  assign \new_[9498]_  = \new_[10]_  | \new_[9497]_ ;
  assign \new_[9499]_  = \new_[9498]_  | \new_[9493]_ ;
  assign \new_[9503]_  = \new_[5]_  | \new_[6]_ ;
  assign \new_[9504]_  = \new_[7]_  | \new_[9503]_ ;
  assign \new_[9507]_  = \new_[3]_  | \new_[4]_ ;
  assign \new_[9510]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[9511]_  = \new_[9510]_  | \new_[9507]_ ;
  assign \new_[9512]_  = \new_[9511]_  | \new_[9504]_ ;
  assign \new_[9513]_  = \new_[9512]_  | \new_[9499]_ ;
  assign \new_[9514]_  = \new_[9513]_  | \new_[9488]_ ;
  assign \new_[9515]_  = \new_[9514]_  | \new_[9465]_ ;
  assign \new_[9516]_  = \new_[9515]_  | \new_[9416]_ ;
  assign \new_[9517]_  = \new_[9516]_  | \new_[9317]_ ;
  assign \new_[9518]_  = \new_[9517]_  | \new_[9120]_ ;
  assign \new_[9519]_  = \new_[9518]_  | \new_[8725]_ ;
  assign \new_[9520]_  = \new_[9519]_  | \new_[7932]_ ;
  assign \new_[9523]_  = A166 & A168;
  assign \new_[9526]_  = A200 & A199;
  assign \new_[9527]_  = \new_[9526]_  & \new_[9523]_ ;
  assign \new_[9530]_  = A233 & ~A232;
  assign \new_[9533]_  = ~A300 & ~A299;
  assign \new_[9534]_  = \new_[9533]_  & \new_[9530]_ ;
  assign \new_[9537]_  = A166 & A168;
  assign \new_[9540]_  = A200 & A199;
  assign \new_[9541]_  = \new_[9540]_  & \new_[9537]_ ;
  assign \new_[9544]_  = A233 & ~A232;
  assign \new_[9547]_  = A299 & A298;
  assign \new_[9548]_  = \new_[9547]_  & \new_[9544]_ ;
  assign \new_[9551]_  = A166 & A168;
  assign \new_[9554]_  = A200 & A199;
  assign \new_[9555]_  = \new_[9554]_  & \new_[9551]_ ;
  assign \new_[9558]_  = A233 & ~A232;
  assign \new_[9561]_  = ~A299 & ~A298;
  assign \new_[9562]_  = \new_[9561]_  & \new_[9558]_ ;
  assign \new_[9565]_  = A166 & A168;
  assign \new_[9568]_  = A200 & A199;
  assign \new_[9569]_  = \new_[9568]_  & \new_[9565]_ ;
  assign \new_[9572]_  = A233 & ~A232;
  assign \new_[9575]_  = A266 & ~A265;
  assign \new_[9576]_  = \new_[9575]_  & \new_[9572]_ ;
  assign \new_[9579]_  = A166 & A168;
  assign \new_[9582]_  = ~A201 & ~A200;
  assign \new_[9583]_  = \new_[9582]_  & \new_[9579]_ ;
  assign \new_[9586]_  = A233 & ~A232;
  assign \new_[9589]_  = ~A300 & ~A299;
  assign \new_[9590]_  = \new_[9589]_  & \new_[9586]_ ;
  assign \new_[9593]_  = A166 & A168;
  assign \new_[9596]_  = ~A201 & ~A200;
  assign \new_[9597]_  = \new_[9596]_  & \new_[9593]_ ;
  assign \new_[9600]_  = A233 & ~A232;
  assign \new_[9603]_  = A299 & A298;
  assign \new_[9604]_  = \new_[9603]_  & \new_[9600]_ ;
  assign \new_[9607]_  = A166 & A168;
  assign \new_[9610]_  = ~A201 & ~A200;
  assign \new_[9611]_  = \new_[9610]_  & \new_[9607]_ ;
  assign \new_[9614]_  = A233 & ~A232;
  assign \new_[9617]_  = ~A299 & ~A298;
  assign \new_[9618]_  = \new_[9617]_  & \new_[9614]_ ;
  assign \new_[9621]_  = A166 & A168;
  assign \new_[9624]_  = ~A201 & ~A200;
  assign \new_[9625]_  = \new_[9624]_  & \new_[9621]_ ;
  assign \new_[9628]_  = A233 & ~A232;
  assign \new_[9631]_  = A266 & ~A265;
  assign \new_[9632]_  = \new_[9631]_  & \new_[9628]_ ;
  assign \new_[9635]_  = A166 & A168;
  assign \new_[9638]_  = ~A200 & ~A199;
  assign \new_[9639]_  = \new_[9638]_  & \new_[9635]_ ;
  assign \new_[9642]_  = A233 & ~A232;
  assign \new_[9645]_  = ~A300 & ~A299;
  assign \new_[9646]_  = \new_[9645]_  & \new_[9642]_ ;
  assign \new_[9649]_  = A166 & A168;
  assign \new_[9652]_  = ~A200 & ~A199;
  assign \new_[9653]_  = \new_[9652]_  & \new_[9649]_ ;
  assign \new_[9656]_  = A233 & ~A232;
  assign \new_[9659]_  = A299 & A298;
  assign \new_[9660]_  = \new_[9659]_  & \new_[9656]_ ;
  assign \new_[9663]_  = A166 & A168;
  assign \new_[9666]_  = ~A200 & ~A199;
  assign \new_[9667]_  = \new_[9666]_  & \new_[9663]_ ;
  assign \new_[9670]_  = A233 & ~A232;
  assign \new_[9673]_  = ~A299 & ~A298;
  assign \new_[9674]_  = \new_[9673]_  & \new_[9670]_ ;
  assign \new_[9677]_  = A166 & A168;
  assign \new_[9680]_  = ~A200 & ~A199;
  assign \new_[9681]_  = \new_[9680]_  & \new_[9677]_ ;
  assign \new_[9684]_  = A233 & ~A232;
  assign \new_[9687]_  = A266 & ~A265;
  assign \new_[9688]_  = \new_[9687]_  & \new_[9684]_ ;
  assign \new_[9691]_  = A167 & A168;
  assign \new_[9694]_  = A200 & A199;
  assign \new_[9695]_  = \new_[9694]_  & \new_[9691]_ ;
  assign \new_[9698]_  = A233 & ~A232;
  assign \new_[9701]_  = ~A300 & ~A299;
  assign \new_[9702]_  = \new_[9701]_  & \new_[9698]_ ;
  assign \new_[9705]_  = A167 & A168;
  assign \new_[9708]_  = A200 & A199;
  assign \new_[9709]_  = \new_[9708]_  & \new_[9705]_ ;
  assign \new_[9712]_  = A233 & ~A232;
  assign \new_[9715]_  = A299 & A298;
  assign \new_[9716]_  = \new_[9715]_  & \new_[9712]_ ;
  assign \new_[9719]_  = A167 & A168;
  assign \new_[9722]_  = A200 & A199;
  assign \new_[9723]_  = \new_[9722]_  & \new_[9719]_ ;
  assign \new_[9726]_  = A233 & ~A232;
  assign \new_[9729]_  = ~A299 & ~A298;
  assign \new_[9730]_  = \new_[9729]_  & \new_[9726]_ ;
  assign \new_[9733]_  = A167 & A168;
  assign \new_[9736]_  = A200 & A199;
  assign \new_[9737]_  = \new_[9736]_  & \new_[9733]_ ;
  assign \new_[9740]_  = A233 & ~A232;
  assign \new_[9743]_  = A266 & ~A265;
  assign \new_[9744]_  = \new_[9743]_  & \new_[9740]_ ;
  assign \new_[9747]_  = A167 & A168;
  assign \new_[9750]_  = ~A201 & ~A200;
  assign \new_[9751]_  = \new_[9750]_  & \new_[9747]_ ;
  assign \new_[9754]_  = A233 & ~A232;
  assign \new_[9757]_  = ~A300 & ~A299;
  assign \new_[9758]_  = \new_[9757]_  & \new_[9754]_ ;
  assign \new_[9761]_  = A167 & A168;
  assign \new_[9764]_  = ~A201 & ~A200;
  assign \new_[9765]_  = \new_[9764]_  & \new_[9761]_ ;
  assign \new_[9768]_  = A233 & ~A232;
  assign \new_[9771]_  = A299 & A298;
  assign \new_[9772]_  = \new_[9771]_  & \new_[9768]_ ;
  assign \new_[9775]_  = A167 & A168;
  assign \new_[9778]_  = ~A201 & ~A200;
  assign \new_[9779]_  = \new_[9778]_  & \new_[9775]_ ;
  assign \new_[9782]_  = A233 & ~A232;
  assign \new_[9785]_  = ~A299 & ~A298;
  assign \new_[9786]_  = \new_[9785]_  & \new_[9782]_ ;
  assign \new_[9789]_  = A167 & A168;
  assign \new_[9792]_  = ~A201 & ~A200;
  assign \new_[9793]_  = \new_[9792]_  & \new_[9789]_ ;
  assign \new_[9796]_  = A233 & ~A232;
  assign \new_[9799]_  = A266 & ~A265;
  assign \new_[9800]_  = \new_[9799]_  & \new_[9796]_ ;
  assign \new_[9803]_  = A167 & A168;
  assign \new_[9806]_  = ~A200 & ~A199;
  assign \new_[9807]_  = \new_[9806]_  & \new_[9803]_ ;
  assign \new_[9810]_  = A233 & ~A232;
  assign \new_[9813]_  = ~A300 & ~A299;
  assign \new_[9814]_  = \new_[9813]_  & \new_[9810]_ ;
  assign \new_[9817]_  = A167 & A168;
  assign \new_[9820]_  = ~A200 & ~A199;
  assign \new_[9821]_  = \new_[9820]_  & \new_[9817]_ ;
  assign \new_[9824]_  = A233 & ~A232;
  assign \new_[9827]_  = A299 & A298;
  assign \new_[9828]_  = \new_[9827]_  & \new_[9824]_ ;
  assign \new_[9831]_  = A167 & A168;
  assign \new_[9834]_  = ~A200 & ~A199;
  assign \new_[9835]_  = \new_[9834]_  & \new_[9831]_ ;
  assign \new_[9838]_  = A233 & ~A232;
  assign \new_[9841]_  = ~A299 & ~A298;
  assign \new_[9842]_  = \new_[9841]_  & \new_[9838]_ ;
  assign \new_[9845]_  = A167 & A168;
  assign \new_[9848]_  = ~A200 & ~A199;
  assign \new_[9849]_  = \new_[9848]_  & \new_[9845]_ ;
  assign \new_[9852]_  = A233 & ~A232;
  assign \new_[9855]_  = A266 & ~A265;
  assign \new_[9856]_  = \new_[9855]_  & \new_[9852]_ ;
  assign \new_[9859]_  = A166 & A168;
  assign \new_[9862]_  = A200 & A199;
  assign \new_[9863]_  = \new_[9862]_  & \new_[9859]_ ;
  assign \new_[9866]_  = A233 & ~A232;
  assign \new_[9870]_  = ~A302 & ~A301;
  assign \new_[9871]_  = ~A299 & \new_[9870]_ ;
  assign \new_[9872]_  = \new_[9871]_  & \new_[9866]_ ;
  assign \new_[9875]_  = A166 & A168;
  assign \new_[9878]_  = ~A202 & ~A200;
  assign \new_[9879]_  = \new_[9878]_  & \new_[9875]_ ;
  assign \new_[9882]_  = ~A232 & ~A203;
  assign \new_[9886]_  = ~A300 & ~A299;
  assign \new_[9887]_  = A233 & \new_[9886]_ ;
  assign \new_[9888]_  = \new_[9887]_  & \new_[9882]_ ;
  assign \new_[9891]_  = A166 & A168;
  assign \new_[9894]_  = ~A202 & ~A200;
  assign \new_[9895]_  = \new_[9894]_  & \new_[9891]_ ;
  assign \new_[9898]_  = ~A232 & ~A203;
  assign \new_[9902]_  = A299 & A298;
  assign \new_[9903]_  = A233 & \new_[9902]_ ;
  assign \new_[9904]_  = \new_[9903]_  & \new_[9898]_ ;
  assign \new_[9907]_  = A166 & A168;
  assign \new_[9910]_  = ~A202 & ~A200;
  assign \new_[9911]_  = \new_[9910]_  & \new_[9907]_ ;
  assign \new_[9914]_  = ~A232 & ~A203;
  assign \new_[9918]_  = ~A299 & ~A298;
  assign \new_[9919]_  = A233 & \new_[9918]_ ;
  assign \new_[9920]_  = \new_[9919]_  & \new_[9914]_ ;
  assign \new_[9923]_  = A166 & A168;
  assign \new_[9926]_  = ~A202 & ~A200;
  assign \new_[9927]_  = \new_[9926]_  & \new_[9923]_ ;
  assign \new_[9930]_  = ~A232 & ~A203;
  assign \new_[9934]_  = A266 & ~A265;
  assign \new_[9935]_  = A233 & \new_[9934]_ ;
  assign \new_[9936]_  = \new_[9935]_  & \new_[9930]_ ;
  assign \new_[9939]_  = A166 & A168;
  assign \new_[9942]_  = ~A201 & ~A200;
  assign \new_[9943]_  = \new_[9942]_  & \new_[9939]_ ;
  assign \new_[9946]_  = A233 & ~A232;
  assign \new_[9950]_  = ~A302 & ~A301;
  assign \new_[9951]_  = ~A299 & \new_[9950]_ ;
  assign \new_[9952]_  = \new_[9951]_  & \new_[9946]_ ;
  assign \new_[9955]_  = A166 & A168;
  assign \new_[9958]_  = ~A200 & ~A199;
  assign \new_[9959]_  = \new_[9958]_  & \new_[9955]_ ;
  assign \new_[9962]_  = A233 & ~A232;
  assign \new_[9966]_  = ~A302 & ~A301;
  assign \new_[9967]_  = ~A299 & \new_[9966]_ ;
  assign \new_[9968]_  = \new_[9967]_  & \new_[9962]_ ;
  assign \new_[9971]_  = A167 & A168;
  assign \new_[9974]_  = A200 & A199;
  assign \new_[9975]_  = \new_[9974]_  & \new_[9971]_ ;
  assign \new_[9978]_  = A233 & ~A232;
  assign \new_[9982]_  = ~A302 & ~A301;
  assign \new_[9983]_  = ~A299 & \new_[9982]_ ;
  assign \new_[9984]_  = \new_[9983]_  & \new_[9978]_ ;
  assign \new_[9987]_  = A167 & A168;
  assign \new_[9990]_  = ~A202 & ~A200;
  assign \new_[9991]_  = \new_[9990]_  & \new_[9987]_ ;
  assign \new_[9994]_  = ~A232 & ~A203;
  assign \new_[9998]_  = ~A300 & ~A299;
  assign \new_[9999]_  = A233 & \new_[9998]_ ;
  assign \new_[10000]_  = \new_[9999]_  & \new_[9994]_ ;
  assign \new_[10003]_  = A167 & A168;
  assign \new_[10006]_  = ~A202 & ~A200;
  assign \new_[10007]_  = \new_[10006]_  & \new_[10003]_ ;
  assign \new_[10010]_  = ~A232 & ~A203;
  assign \new_[10014]_  = A299 & A298;
  assign \new_[10015]_  = A233 & \new_[10014]_ ;
  assign \new_[10016]_  = \new_[10015]_  & \new_[10010]_ ;
  assign \new_[10019]_  = A167 & A168;
  assign \new_[10022]_  = ~A202 & ~A200;
  assign \new_[10023]_  = \new_[10022]_  & \new_[10019]_ ;
  assign \new_[10026]_  = ~A232 & ~A203;
  assign \new_[10030]_  = ~A299 & ~A298;
  assign \new_[10031]_  = A233 & \new_[10030]_ ;
  assign \new_[10032]_  = \new_[10031]_  & \new_[10026]_ ;
  assign \new_[10035]_  = A167 & A168;
  assign \new_[10038]_  = ~A202 & ~A200;
  assign \new_[10039]_  = \new_[10038]_  & \new_[10035]_ ;
  assign \new_[10042]_  = ~A232 & ~A203;
  assign \new_[10046]_  = A266 & ~A265;
  assign \new_[10047]_  = A233 & \new_[10046]_ ;
  assign \new_[10048]_  = \new_[10047]_  & \new_[10042]_ ;
  assign \new_[10051]_  = A167 & A168;
  assign \new_[10054]_  = ~A201 & ~A200;
  assign \new_[10055]_  = \new_[10054]_  & \new_[10051]_ ;
  assign \new_[10058]_  = A233 & ~A232;
  assign \new_[10062]_  = ~A302 & ~A301;
  assign \new_[10063]_  = ~A299 & \new_[10062]_ ;
  assign \new_[10064]_  = \new_[10063]_  & \new_[10058]_ ;
  assign \new_[10067]_  = A167 & A168;
  assign \new_[10070]_  = ~A200 & ~A199;
  assign \new_[10071]_  = \new_[10070]_  & \new_[10067]_ ;
  assign \new_[10074]_  = A233 & ~A232;
  assign \new_[10078]_  = ~A302 & ~A301;
  assign \new_[10079]_  = ~A299 & \new_[10078]_ ;
  assign \new_[10080]_  = \new_[10079]_  & \new_[10074]_ ;
  assign \new_[10083]_  = ~A167 & A170;
  assign \new_[10086]_  = ~A199 & ~A166;
  assign \new_[10087]_  = \new_[10086]_  & \new_[10083]_ ;
  assign \new_[10090]_  = ~A232 & A200;
  assign \new_[10094]_  = ~A300 & ~A299;
  assign \new_[10095]_  = A233 & \new_[10094]_ ;
  assign \new_[10096]_  = \new_[10095]_  & \new_[10090]_ ;
  assign \new_[10099]_  = ~A167 & A170;
  assign \new_[10102]_  = ~A199 & ~A166;
  assign \new_[10103]_  = \new_[10102]_  & \new_[10099]_ ;
  assign \new_[10106]_  = ~A232 & A200;
  assign \new_[10110]_  = A299 & A298;
  assign \new_[10111]_  = A233 & \new_[10110]_ ;
  assign \new_[10112]_  = \new_[10111]_  & \new_[10106]_ ;
  assign \new_[10115]_  = ~A167 & A170;
  assign \new_[10118]_  = ~A199 & ~A166;
  assign \new_[10119]_  = \new_[10118]_  & \new_[10115]_ ;
  assign \new_[10122]_  = ~A232 & A200;
  assign \new_[10126]_  = ~A299 & ~A298;
  assign \new_[10127]_  = A233 & \new_[10126]_ ;
  assign \new_[10128]_  = \new_[10127]_  & \new_[10122]_ ;
  assign \new_[10131]_  = ~A167 & A170;
  assign \new_[10134]_  = ~A199 & ~A166;
  assign \new_[10135]_  = \new_[10134]_  & \new_[10131]_ ;
  assign \new_[10138]_  = ~A232 & A200;
  assign \new_[10142]_  = A266 & ~A265;
  assign \new_[10143]_  = A233 & \new_[10142]_ ;
  assign \new_[10144]_  = \new_[10143]_  & \new_[10138]_ ;
  assign \new_[10147]_  = ~A167 & ~A169;
  assign \new_[10150]_  = ~A199 & ~A166;
  assign \new_[10151]_  = \new_[10150]_  & \new_[10147]_ ;
  assign \new_[10154]_  = ~A232 & A200;
  assign \new_[10158]_  = ~A300 & ~A299;
  assign \new_[10159]_  = A233 & \new_[10158]_ ;
  assign \new_[10160]_  = \new_[10159]_  & \new_[10154]_ ;
  assign \new_[10163]_  = ~A167 & ~A169;
  assign \new_[10166]_  = ~A199 & ~A166;
  assign \new_[10167]_  = \new_[10166]_  & \new_[10163]_ ;
  assign \new_[10170]_  = ~A232 & A200;
  assign \new_[10174]_  = A299 & A298;
  assign \new_[10175]_  = A233 & \new_[10174]_ ;
  assign \new_[10176]_  = \new_[10175]_  & \new_[10170]_ ;
  assign \new_[10179]_  = ~A167 & ~A169;
  assign \new_[10182]_  = ~A199 & ~A166;
  assign \new_[10183]_  = \new_[10182]_  & \new_[10179]_ ;
  assign \new_[10186]_  = ~A232 & A200;
  assign \new_[10190]_  = ~A299 & ~A298;
  assign \new_[10191]_  = A233 & \new_[10190]_ ;
  assign \new_[10192]_  = \new_[10191]_  & \new_[10186]_ ;
  assign \new_[10195]_  = ~A167 & ~A169;
  assign \new_[10198]_  = ~A199 & ~A166;
  assign \new_[10199]_  = \new_[10198]_  & \new_[10195]_ ;
  assign \new_[10202]_  = ~A232 & A200;
  assign \new_[10206]_  = A266 & ~A265;
  assign \new_[10207]_  = A233 & \new_[10206]_ ;
  assign \new_[10208]_  = \new_[10207]_  & \new_[10202]_ ;
  assign \new_[10211]_  = A166 & A168;
  assign \new_[10215]_  = A232 & A200;
  assign \new_[10216]_  = A199 & \new_[10215]_ ;
  assign \new_[10217]_  = \new_[10216]_  & \new_[10211]_ ;
  assign \new_[10220]_  = A265 & A233;
  assign \new_[10224]_  = A299 & ~A298;
  assign \new_[10225]_  = ~A267 & \new_[10224]_ ;
  assign \new_[10226]_  = \new_[10225]_  & \new_[10220]_ ;
  assign \new_[10229]_  = A166 & A168;
  assign \new_[10233]_  = A232 & A200;
  assign \new_[10234]_  = A199 & \new_[10233]_ ;
  assign \new_[10235]_  = \new_[10234]_  & \new_[10229]_ ;
  assign \new_[10238]_  = A265 & A233;
  assign \new_[10242]_  = A299 & ~A298;
  assign \new_[10243]_  = A266 & \new_[10242]_ ;
  assign \new_[10244]_  = \new_[10243]_  & \new_[10238]_ ;
  assign \new_[10247]_  = A166 & A168;
  assign \new_[10251]_  = A232 & A200;
  assign \new_[10252]_  = A199 & \new_[10251]_ ;
  assign \new_[10253]_  = \new_[10252]_  & \new_[10247]_ ;
  assign \new_[10256]_  = ~A265 & A233;
  assign \new_[10260]_  = A299 & ~A298;
  assign \new_[10261]_  = ~A266 & \new_[10260]_ ;
  assign \new_[10262]_  = \new_[10261]_  & \new_[10256]_ ;
  assign \new_[10265]_  = A166 & A168;
  assign \new_[10269]_  = ~A232 & A200;
  assign \new_[10270]_  = A199 & \new_[10269]_ ;
  assign \new_[10271]_  = \new_[10270]_  & \new_[10265]_ ;
  assign \new_[10274]_  = A265 & A233;
  assign \new_[10278]_  = A268 & A267;
  assign \new_[10279]_  = ~A266 & \new_[10278]_ ;
  assign \new_[10280]_  = \new_[10279]_  & \new_[10274]_ ;
  assign \new_[10283]_  = A166 & A168;
  assign \new_[10287]_  = ~A232 & A200;
  assign \new_[10288]_  = A199 & \new_[10287]_ ;
  assign \new_[10289]_  = \new_[10288]_  & \new_[10283]_ ;
  assign \new_[10292]_  = A265 & A233;
  assign \new_[10296]_  = A269 & A267;
  assign \new_[10297]_  = ~A266 & \new_[10296]_ ;
  assign \new_[10298]_  = \new_[10297]_  & \new_[10292]_ ;
  assign \new_[10301]_  = A166 & A168;
  assign \new_[10305]_  = ~A233 & A200;
  assign \new_[10306]_  = A199 & \new_[10305]_ ;
  assign \new_[10307]_  = \new_[10306]_  & \new_[10301]_ ;
  assign \new_[10310]_  = A265 & ~A234;
  assign \new_[10314]_  = A299 & ~A298;
  assign \new_[10315]_  = A266 & \new_[10314]_ ;
  assign \new_[10316]_  = \new_[10315]_  & \new_[10310]_ ;
  assign \new_[10319]_  = A166 & A168;
  assign \new_[10323]_  = ~A233 & A200;
  assign \new_[10324]_  = A199 & \new_[10323]_ ;
  assign \new_[10325]_  = \new_[10324]_  & \new_[10319]_ ;
  assign \new_[10328]_  = ~A266 & ~A234;
  assign \new_[10332]_  = A299 & ~A298;
  assign \new_[10333]_  = ~A267 & \new_[10332]_ ;
  assign \new_[10334]_  = \new_[10333]_  & \new_[10328]_ ;
  assign \new_[10337]_  = A166 & A168;
  assign \new_[10341]_  = ~A233 & A200;
  assign \new_[10342]_  = A199 & \new_[10341]_ ;
  assign \new_[10343]_  = \new_[10342]_  & \new_[10337]_ ;
  assign \new_[10346]_  = ~A265 & ~A234;
  assign \new_[10350]_  = A299 & ~A298;
  assign \new_[10351]_  = ~A266 & \new_[10350]_ ;
  assign \new_[10352]_  = \new_[10351]_  & \new_[10346]_ ;
  assign \new_[10355]_  = A166 & A168;
  assign \new_[10359]_  = A232 & A200;
  assign \new_[10360]_  = A199 & \new_[10359]_ ;
  assign \new_[10361]_  = \new_[10360]_  & \new_[10355]_ ;
  assign \new_[10364]_  = A234 & ~A233;
  assign \new_[10368]_  = ~A300 & A298;
  assign \new_[10369]_  = A235 & \new_[10368]_ ;
  assign \new_[10370]_  = \new_[10369]_  & \new_[10364]_ ;
  assign \new_[10373]_  = A166 & A168;
  assign \new_[10377]_  = A232 & A200;
  assign \new_[10378]_  = A199 & \new_[10377]_ ;
  assign \new_[10379]_  = \new_[10378]_  & \new_[10373]_ ;
  assign \new_[10382]_  = A234 & ~A233;
  assign \new_[10386]_  = A299 & A298;
  assign \new_[10387]_  = A235 & \new_[10386]_ ;
  assign \new_[10388]_  = \new_[10387]_  & \new_[10382]_ ;
  assign \new_[10391]_  = A166 & A168;
  assign \new_[10395]_  = A232 & A200;
  assign \new_[10396]_  = A199 & \new_[10395]_ ;
  assign \new_[10397]_  = \new_[10396]_  & \new_[10391]_ ;
  assign \new_[10400]_  = A234 & ~A233;
  assign \new_[10404]_  = ~A299 & ~A298;
  assign \new_[10405]_  = A235 & \new_[10404]_ ;
  assign \new_[10406]_  = \new_[10405]_  & \new_[10400]_ ;
  assign \new_[10409]_  = A166 & A168;
  assign \new_[10413]_  = A232 & A200;
  assign \new_[10414]_  = A199 & \new_[10413]_ ;
  assign \new_[10415]_  = \new_[10414]_  & \new_[10409]_ ;
  assign \new_[10418]_  = A234 & ~A233;
  assign \new_[10422]_  = A266 & ~A265;
  assign \new_[10423]_  = A235 & \new_[10422]_ ;
  assign \new_[10424]_  = \new_[10423]_  & \new_[10418]_ ;
  assign \new_[10427]_  = A166 & A168;
  assign \new_[10431]_  = A232 & A200;
  assign \new_[10432]_  = A199 & \new_[10431]_ ;
  assign \new_[10433]_  = \new_[10432]_  & \new_[10427]_ ;
  assign \new_[10436]_  = A234 & ~A233;
  assign \new_[10440]_  = ~A300 & A298;
  assign \new_[10441]_  = A236 & \new_[10440]_ ;
  assign \new_[10442]_  = \new_[10441]_  & \new_[10436]_ ;
  assign \new_[10445]_  = A166 & A168;
  assign \new_[10449]_  = A232 & A200;
  assign \new_[10450]_  = A199 & \new_[10449]_ ;
  assign \new_[10451]_  = \new_[10450]_  & \new_[10445]_ ;
  assign \new_[10454]_  = A234 & ~A233;
  assign \new_[10458]_  = A299 & A298;
  assign \new_[10459]_  = A236 & \new_[10458]_ ;
  assign \new_[10460]_  = \new_[10459]_  & \new_[10454]_ ;
  assign \new_[10463]_  = A166 & A168;
  assign \new_[10467]_  = A232 & A200;
  assign \new_[10468]_  = A199 & \new_[10467]_ ;
  assign \new_[10469]_  = \new_[10468]_  & \new_[10463]_ ;
  assign \new_[10472]_  = A234 & ~A233;
  assign \new_[10476]_  = ~A299 & ~A298;
  assign \new_[10477]_  = A236 & \new_[10476]_ ;
  assign \new_[10478]_  = \new_[10477]_  & \new_[10472]_ ;
  assign \new_[10481]_  = A166 & A168;
  assign \new_[10485]_  = A232 & A200;
  assign \new_[10486]_  = A199 & \new_[10485]_ ;
  assign \new_[10487]_  = \new_[10486]_  & \new_[10481]_ ;
  assign \new_[10490]_  = A234 & ~A233;
  assign \new_[10494]_  = A266 & ~A265;
  assign \new_[10495]_  = A236 & \new_[10494]_ ;
  assign \new_[10496]_  = \new_[10495]_  & \new_[10490]_ ;
  assign \new_[10499]_  = A166 & A168;
  assign \new_[10503]_  = ~A232 & A200;
  assign \new_[10504]_  = A199 & \new_[10503]_ ;
  assign \new_[10505]_  = \new_[10504]_  & \new_[10499]_ ;
  assign \new_[10508]_  = A265 & ~A233;
  assign \new_[10512]_  = A299 & ~A298;
  assign \new_[10513]_  = A266 & \new_[10512]_ ;
  assign \new_[10514]_  = \new_[10513]_  & \new_[10508]_ ;
  assign \new_[10517]_  = A166 & A168;
  assign \new_[10521]_  = ~A232 & A200;
  assign \new_[10522]_  = A199 & \new_[10521]_ ;
  assign \new_[10523]_  = \new_[10522]_  & \new_[10517]_ ;
  assign \new_[10526]_  = ~A266 & ~A233;
  assign \new_[10530]_  = A299 & ~A298;
  assign \new_[10531]_  = ~A267 & \new_[10530]_ ;
  assign \new_[10532]_  = \new_[10531]_  & \new_[10526]_ ;
  assign \new_[10535]_  = A166 & A168;
  assign \new_[10539]_  = ~A232 & A200;
  assign \new_[10540]_  = A199 & \new_[10539]_ ;
  assign \new_[10541]_  = \new_[10540]_  & \new_[10535]_ ;
  assign \new_[10544]_  = ~A265 & ~A233;
  assign \new_[10548]_  = A299 & ~A298;
  assign \new_[10549]_  = ~A266 & \new_[10548]_ ;
  assign \new_[10550]_  = \new_[10549]_  & \new_[10544]_ ;
  assign \new_[10553]_  = A166 & A168;
  assign \new_[10557]_  = ~A203 & ~A202;
  assign \new_[10558]_  = ~A200 & \new_[10557]_ ;
  assign \new_[10559]_  = \new_[10558]_  & \new_[10553]_ ;
  assign \new_[10562]_  = A233 & ~A232;
  assign \new_[10566]_  = ~A302 & ~A301;
  assign \new_[10567]_  = ~A299 & \new_[10566]_ ;
  assign \new_[10568]_  = \new_[10567]_  & \new_[10562]_ ;
  assign \new_[10571]_  = A166 & A168;
  assign \new_[10575]_  = A232 & ~A201;
  assign \new_[10576]_  = ~A200 & \new_[10575]_ ;
  assign \new_[10577]_  = \new_[10576]_  & \new_[10571]_ ;
  assign \new_[10580]_  = A265 & A233;
  assign \new_[10584]_  = A299 & ~A298;
  assign \new_[10585]_  = ~A267 & \new_[10584]_ ;
  assign \new_[10586]_  = \new_[10585]_  & \new_[10580]_ ;
  assign \new_[10589]_  = A166 & A168;
  assign \new_[10593]_  = A232 & ~A201;
  assign \new_[10594]_  = ~A200 & \new_[10593]_ ;
  assign \new_[10595]_  = \new_[10594]_  & \new_[10589]_ ;
  assign \new_[10598]_  = A265 & A233;
  assign \new_[10602]_  = A299 & ~A298;
  assign \new_[10603]_  = A266 & \new_[10602]_ ;
  assign \new_[10604]_  = \new_[10603]_  & \new_[10598]_ ;
  assign \new_[10607]_  = A166 & A168;
  assign \new_[10611]_  = A232 & ~A201;
  assign \new_[10612]_  = ~A200 & \new_[10611]_ ;
  assign \new_[10613]_  = \new_[10612]_  & \new_[10607]_ ;
  assign \new_[10616]_  = ~A265 & A233;
  assign \new_[10620]_  = A299 & ~A298;
  assign \new_[10621]_  = ~A266 & \new_[10620]_ ;
  assign \new_[10622]_  = \new_[10621]_  & \new_[10616]_ ;
  assign \new_[10625]_  = A166 & A168;
  assign \new_[10629]_  = ~A232 & ~A201;
  assign \new_[10630]_  = ~A200 & \new_[10629]_ ;
  assign \new_[10631]_  = \new_[10630]_  & \new_[10625]_ ;
  assign \new_[10634]_  = A265 & A233;
  assign \new_[10638]_  = A268 & A267;
  assign \new_[10639]_  = ~A266 & \new_[10638]_ ;
  assign \new_[10640]_  = \new_[10639]_  & \new_[10634]_ ;
  assign \new_[10643]_  = A166 & A168;
  assign \new_[10647]_  = ~A232 & ~A201;
  assign \new_[10648]_  = ~A200 & \new_[10647]_ ;
  assign \new_[10649]_  = \new_[10648]_  & \new_[10643]_ ;
  assign \new_[10652]_  = A265 & A233;
  assign \new_[10656]_  = A269 & A267;
  assign \new_[10657]_  = ~A266 & \new_[10656]_ ;
  assign \new_[10658]_  = \new_[10657]_  & \new_[10652]_ ;
  assign \new_[10661]_  = A166 & A168;
  assign \new_[10665]_  = ~A233 & ~A201;
  assign \new_[10666]_  = ~A200 & \new_[10665]_ ;
  assign \new_[10667]_  = \new_[10666]_  & \new_[10661]_ ;
  assign \new_[10670]_  = A265 & ~A234;
  assign \new_[10674]_  = A299 & ~A298;
  assign \new_[10675]_  = A266 & \new_[10674]_ ;
  assign \new_[10676]_  = \new_[10675]_  & \new_[10670]_ ;
  assign \new_[10679]_  = A166 & A168;
  assign \new_[10683]_  = ~A233 & ~A201;
  assign \new_[10684]_  = ~A200 & \new_[10683]_ ;
  assign \new_[10685]_  = \new_[10684]_  & \new_[10679]_ ;
  assign \new_[10688]_  = ~A266 & ~A234;
  assign \new_[10692]_  = A299 & ~A298;
  assign \new_[10693]_  = ~A267 & \new_[10692]_ ;
  assign \new_[10694]_  = \new_[10693]_  & \new_[10688]_ ;
  assign \new_[10697]_  = A166 & A168;
  assign \new_[10701]_  = ~A233 & ~A201;
  assign \new_[10702]_  = ~A200 & \new_[10701]_ ;
  assign \new_[10703]_  = \new_[10702]_  & \new_[10697]_ ;
  assign \new_[10706]_  = ~A265 & ~A234;
  assign \new_[10710]_  = A299 & ~A298;
  assign \new_[10711]_  = ~A266 & \new_[10710]_ ;
  assign \new_[10712]_  = \new_[10711]_  & \new_[10706]_ ;
  assign \new_[10715]_  = A166 & A168;
  assign \new_[10719]_  = A232 & ~A201;
  assign \new_[10720]_  = ~A200 & \new_[10719]_ ;
  assign \new_[10721]_  = \new_[10720]_  & \new_[10715]_ ;
  assign \new_[10724]_  = A234 & ~A233;
  assign \new_[10728]_  = ~A300 & A298;
  assign \new_[10729]_  = A235 & \new_[10728]_ ;
  assign \new_[10730]_  = \new_[10729]_  & \new_[10724]_ ;
  assign \new_[10733]_  = A166 & A168;
  assign \new_[10737]_  = A232 & ~A201;
  assign \new_[10738]_  = ~A200 & \new_[10737]_ ;
  assign \new_[10739]_  = \new_[10738]_  & \new_[10733]_ ;
  assign \new_[10742]_  = A234 & ~A233;
  assign \new_[10746]_  = A299 & A298;
  assign \new_[10747]_  = A235 & \new_[10746]_ ;
  assign \new_[10748]_  = \new_[10747]_  & \new_[10742]_ ;
  assign \new_[10751]_  = A166 & A168;
  assign \new_[10755]_  = A232 & ~A201;
  assign \new_[10756]_  = ~A200 & \new_[10755]_ ;
  assign \new_[10757]_  = \new_[10756]_  & \new_[10751]_ ;
  assign \new_[10760]_  = A234 & ~A233;
  assign \new_[10764]_  = ~A299 & ~A298;
  assign \new_[10765]_  = A235 & \new_[10764]_ ;
  assign \new_[10766]_  = \new_[10765]_  & \new_[10760]_ ;
  assign \new_[10769]_  = A166 & A168;
  assign \new_[10773]_  = A232 & ~A201;
  assign \new_[10774]_  = ~A200 & \new_[10773]_ ;
  assign \new_[10775]_  = \new_[10774]_  & \new_[10769]_ ;
  assign \new_[10778]_  = A234 & ~A233;
  assign \new_[10782]_  = A266 & ~A265;
  assign \new_[10783]_  = A235 & \new_[10782]_ ;
  assign \new_[10784]_  = \new_[10783]_  & \new_[10778]_ ;
  assign \new_[10787]_  = A166 & A168;
  assign \new_[10791]_  = A232 & ~A201;
  assign \new_[10792]_  = ~A200 & \new_[10791]_ ;
  assign \new_[10793]_  = \new_[10792]_  & \new_[10787]_ ;
  assign \new_[10796]_  = A234 & ~A233;
  assign \new_[10800]_  = ~A300 & A298;
  assign \new_[10801]_  = A236 & \new_[10800]_ ;
  assign \new_[10802]_  = \new_[10801]_  & \new_[10796]_ ;
  assign \new_[10805]_  = A166 & A168;
  assign \new_[10809]_  = A232 & ~A201;
  assign \new_[10810]_  = ~A200 & \new_[10809]_ ;
  assign \new_[10811]_  = \new_[10810]_  & \new_[10805]_ ;
  assign \new_[10814]_  = A234 & ~A233;
  assign \new_[10818]_  = A299 & A298;
  assign \new_[10819]_  = A236 & \new_[10818]_ ;
  assign \new_[10820]_  = \new_[10819]_  & \new_[10814]_ ;
  assign \new_[10823]_  = A166 & A168;
  assign \new_[10827]_  = A232 & ~A201;
  assign \new_[10828]_  = ~A200 & \new_[10827]_ ;
  assign \new_[10829]_  = \new_[10828]_  & \new_[10823]_ ;
  assign \new_[10832]_  = A234 & ~A233;
  assign \new_[10836]_  = ~A299 & ~A298;
  assign \new_[10837]_  = A236 & \new_[10836]_ ;
  assign \new_[10838]_  = \new_[10837]_  & \new_[10832]_ ;
  assign \new_[10841]_  = A166 & A168;
  assign \new_[10845]_  = A232 & ~A201;
  assign \new_[10846]_  = ~A200 & \new_[10845]_ ;
  assign \new_[10847]_  = \new_[10846]_  & \new_[10841]_ ;
  assign \new_[10850]_  = A234 & ~A233;
  assign \new_[10854]_  = A266 & ~A265;
  assign \new_[10855]_  = A236 & \new_[10854]_ ;
  assign \new_[10856]_  = \new_[10855]_  & \new_[10850]_ ;
  assign \new_[10859]_  = A166 & A168;
  assign \new_[10863]_  = ~A232 & ~A201;
  assign \new_[10864]_  = ~A200 & \new_[10863]_ ;
  assign \new_[10865]_  = \new_[10864]_  & \new_[10859]_ ;
  assign \new_[10868]_  = A265 & ~A233;
  assign \new_[10872]_  = A299 & ~A298;
  assign \new_[10873]_  = A266 & \new_[10872]_ ;
  assign \new_[10874]_  = \new_[10873]_  & \new_[10868]_ ;
  assign \new_[10877]_  = A166 & A168;
  assign \new_[10881]_  = ~A232 & ~A201;
  assign \new_[10882]_  = ~A200 & \new_[10881]_ ;
  assign \new_[10883]_  = \new_[10882]_  & \new_[10877]_ ;
  assign \new_[10886]_  = ~A266 & ~A233;
  assign \new_[10890]_  = A299 & ~A298;
  assign \new_[10891]_  = ~A267 & \new_[10890]_ ;
  assign \new_[10892]_  = \new_[10891]_  & \new_[10886]_ ;
  assign \new_[10895]_  = A166 & A168;
  assign \new_[10899]_  = ~A232 & ~A201;
  assign \new_[10900]_  = ~A200 & \new_[10899]_ ;
  assign \new_[10901]_  = \new_[10900]_  & \new_[10895]_ ;
  assign \new_[10904]_  = ~A265 & ~A233;
  assign \new_[10908]_  = A299 & ~A298;
  assign \new_[10909]_  = ~A266 & \new_[10908]_ ;
  assign \new_[10910]_  = \new_[10909]_  & \new_[10904]_ ;
  assign \new_[10913]_  = A166 & A168;
  assign \new_[10917]_  = A232 & ~A200;
  assign \new_[10918]_  = ~A199 & \new_[10917]_ ;
  assign \new_[10919]_  = \new_[10918]_  & \new_[10913]_ ;
  assign \new_[10922]_  = A265 & A233;
  assign \new_[10926]_  = A299 & ~A298;
  assign \new_[10927]_  = ~A267 & \new_[10926]_ ;
  assign \new_[10928]_  = \new_[10927]_  & \new_[10922]_ ;
  assign \new_[10931]_  = A166 & A168;
  assign \new_[10935]_  = A232 & ~A200;
  assign \new_[10936]_  = ~A199 & \new_[10935]_ ;
  assign \new_[10937]_  = \new_[10936]_  & \new_[10931]_ ;
  assign \new_[10940]_  = A265 & A233;
  assign \new_[10944]_  = A299 & ~A298;
  assign \new_[10945]_  = A266 & \new_[10944]_ ;
  assign \new_[10946]_  = \new_[10945]_  & \new_[10940]_ ;
  assign \new_[10949]_  = A166 & A168;
  assign \new_[10953]_  = A232 & ~A200;
  assign \new_[10954]_  = ~A199 & \new_[10953]_ ;
  assign \new_[10955]_  = \new_[10954]_  & \new_[10949]_ ;
  assign \new_[10958]_  = ~A265 & A233;
  assign \new_[10962]_  = A299 & ~A298;
  assign \new_[10963]_  = ~A266 & \new_[10962]_ ;
  assign \new_[10964]_  = \new_[10963]_  & \new_[10958]_ ;
  assign \new_[10967]_  = A166 & A168;
  assign \new_[10971]_  = ~A232 & ~A200;
  assign \new_[10972]_  = ~A199 & \new_[10971]_ ;
  assign \new_[10973]_  = \new_[10972]_  & \new_[10967]_ ;
  assign \new_[10976]_  = A265 & A233;
  assign \new_[10980]_  = A268 & A267;
  assign \new_[10981]_  = ~A266 & \new_[10980]_ ;
  assign \new_[10982]_  = \new_[10981]_  & \new_[10976]_ ;
  assign \new_[10985]_  = A166 & A168;
  assign \new_[10989]_  = ~A232 & ~A200;
  assign \new_[10990]_  = ~A199 & \new_[10989]_ ;
  assign \new_[10991]_  = \new_[10990]_  & \new_[10985]_ ;
  assign \new_[10994]_  = A265 & A233;
  assign \new_[10998]_  = A269 & A267;
  assign \new_[10999]_  = ~A266 & \new_[10998]_ ;
  assign \new_[11000]_  = \new_[10999]_  & \new_[10994]_ ;
  assign \new_[11003]_  = A166 & A168;
  assign \new_[11007]_  = ~A233 & ~A200;
  assign \new_[11008]_  = ~A199 & \new_[11007]_ ;
  assign \new_[11009]_  = \new_[11008]_  & \new_[11003]_ ;
  assign \new_[11012]_  = A265 & ~A234;
  assign \new_[11016]_  = A299 & ~A298;
  assign \new_[11017]_  = A266 & \new_[11016]_ ;
  assign \new_[11018]_  = \new_[11017]_  & \new_[11012]_ ;
  assign \new_[11021]_  = A166 & A168;
  assign \new_[11025]_  = ~A233 & ~A200;
  assign \new_[11026]_  = ~A199 & \new_[11025]_ ;
  assign \new_[11027]_  = \new_[11026]_  & \new_[11021]_ ;
  assign \new_[11030]_  = ~A266 & ~A234;
  assign \new_[11034]_  = A299 & ~A298;
  assign \new_[11035]_  = ~A267 & \new_[11034]_ ;
  assign \new_[11036]_  = \new_[11035]_  & \new_[11030]_ ;
  assign \new_[11039]_  = A166 & A168;
  assign \new_[11043]_  = ~A233 & ~A200;
  assign \new_[11044]_  = ~A199 & \new_[11043]_ ;
  assign \new_[11045]_  = \new_[11044]_  & \new_[11039]_ ;
  assign \new_[11048]_  = ~A265 & ~A234;
  assign \new_[11052]_  = A299 & ~A298;
  assign \new_[11053]_  = ~A266 & \new_[11052]_ ;
  assign \new_[11054]_  = \new_[11053]_  & \new_[11048]_ ;
  assign \new_[11057]_  = A166 & A168;
  assign \new_[11061]_  = A232 & ~A200;
  assign \new_[11062]_  = ~A199 & \new_[11061]_ ;
  assign \new_[11063]_  = \new_[11062]_  & \new_[11057]_ ;
  assign \new_[11066]_  = A234 & ~A233;
  assign \new_[11070]_  = ~A300 & A298;
  assign \new_[11071]_  = A235 & \new_[11070]_ ;
  assign \new_[11072]_  = \new_[11071]_  & \new_[11066]_ ;
  assign \new_[11075]_  = A166 & A168;
  assign \new_[11079]_  = A232 & ~A200;
  assign \new_[11080]_  = ~A199 & \new_[11079]_ ;
  assign \new_[11081]_  = \new_[11080]_  & \new_[11075]_ ;
  assign \new_[11084]_  = A234 & ~A233;
  assign \new_[11088]_  = A299 & A298;
  assign \new_[11089]_  = A235 & \new_[11088]_ ;
  assign \new_[11090]_  = \new_[11089]_  & \new_[11084]_ ;
  assign \new_[11093]_  = A166 & A168;
  assign \new_[11097]_  = A232 & ~A200;
  assign \new_[11098]_  = ~A199 & \new_[11097]_ ;
  assign \new_[11099]_  = \new_[11098]_  & \new_[11093]_ ;
  assign \new_[11102]_  = A234 & ~A233;
  assign \new_[11106]_  = ~A299 & ~A298;
  assign \new_[11107]_  = A235 & \new_[11106]_ ;
  assign \new_[11108]_  = \new_[11107]_  & \new_[11102]_ ;
  assign \new_[11111]_  = A166 & A168;
  assign \new_[11115]_  = A232 & ~A200;
  assign \new_[11116]_  = ~A199 & \new_[11115]_ ;
  assign \new_[11117]_  = \new_[11116]_  & \new_[11111]_ ;
  assign \new_[11120]_  = A234 & ~A233;
  assign \new_[11124]_  = A266 & ~A265;
  assign \new_[11125]_  = A235 & \new_[11124]_ ;
  assign \new_[11126]_  = \new_[11125]_  & \new_[11120]_ ;
  assign \new_[11129]_  = A166 & A168;
  assign \new_[11133]_  = A232 & ~A200;
  assign \new_[11134]_  = ~A199 & \new_[11133]_ ;
  assign \new_[11135]_  = \new_[11134]_  & \new_[11129]_ ;
  assign \new_[11138]_  = A234 & ~A233;
  assign \new_[11142]_  = ~A300 & A298;
  assign \new_[11143]_  = A236 & \new_[11142]_ ;
  assign \new_[11144]_  = \new_[11143]_  & \new_[11138]_ ;
  assign \new_[11147]_  = A166 & A168;
  assign \new_[11151]_  = A232 & ~A200;
  assign \new_[11152]_  = ~A199 & \new_[11151]_ ;
  assign \new_[11153]_  = \new_[11152]_  & \new_[11147]_ ;
  assign \new_[11156]_  = A234 & ~A233;
  assign \new_[11160]_  = A299 & A298;
  assign \new_[11161]_  = A236 & \new_[11160]_ ;
  assign \new_[11162]_  = \new_[11161]_  & \new_[11156]_ ;
  assign \new_[11165]_  = A166 & A168;
  assign \new_[11169]_  = A232 & ~A200;
  assign \new_[11170]_  = ~A199 & \new_[11169]_ ;
  assign \new_[11171]_  = \new_[11170]_  & \new_[11165]_ ;
  assign \new_[11174]_  = A234 & ~A233;
  assign \new_[11178]_  = ~A299 & ~A298;
  assign \new_[11179]_  = A236 & \new_[11178]_ ;
  assign \new_[11180]_  = \new_[11179]_  & \new_[11174]_ ;
  assign \new_[11183]_  = A166 & A168;
  assign \new_[11187]_  = A232 & ~A200;
  assign \new_[11188]_  = ~A199 & \new_[11187]_ ;
  assign \new_[11189]_  = \new_[11188]_  & \new_[11183]_ ;
  assign \new_[11192]_  = A234 & ~A233;
  assign \new_[11196]_  = A266 & ~A265;
  assign \new_[11197]_  = A236 & \new_[11196]_ ;
  assign \new_[11198]_  = \new_[11197]_  & \new_[11192]_ ;
  assign \new_[11201]_  = A166 & A168;
  assign \new_[11205]_  = ~A232 & ~A200;
  assign \new_[11206]_  = ~A199 & \new_[11205]_ ;
  assign \new_[11207]_  = \new_[11206]_  & \new_[11201]_ ;
  assign \new_[11210]_  = A265 & ~A233;
  assign \new_[11214]_  = A299 & ~A298;
  assign \new_[11215]_  = A266 & \new_[11214]_ ;
  assign \new_[11216]_  = \new_[11215]_  & \new_[11210]_ ;
  assign \new_[11219]_  = A166 & A168;
  assign \new_[11223]_  = ~A232 & ~A200;
  assign \new_[11224]_  = ~A199 & \new_[11223]_ ;
  assign \new_[11225]_  = \new_[11224]_  & \new_[11219]_ ;
  assign \new_[11228]_  = ~A266 & ~A233;
  assign \new_[11232]_  = A299 & ~A298;
  assign \new_[11233]_  = ~A267 & \new_[11232]_ ;
  assign \new_[11234]_  = \new_[11233]_  & \new_[11228]_ ;
  assign \new_[11237]_  = A166 & A168;
  assign \new_[11241]_  = ~A232 & ~A200;
  assign \new_[11242]_  = ~A199 & \new_[11241]_ ;
  assign \new_[11243]_  = \new_[11242]_  & \new_[11237]_ ;
  assign \new_[11246]_  = ~A265 & ~A233;
  assign \new_[11250]_  = A299 & ~A298;
  assign \new_[11251]_  = ~A266 & \new_[11250]_ ;
  assign \new_[11252]_  = \new_[11251]_  & \new_[11246]_ ;
  assign \new_[11255]_  = A167 & A168;
  assign \new_[11259]_  = A232 & A200;
  assign \new_[11260]_  = A199 & \new_[11259]_ ;
  assign \new_[11261]_  = \new_[11260]_  & \new_[11255]_ ;
  assign \new_[11264]_  = A265 & A233;
  assign \new_[11268]_  = A299 & ~A298;
  assign \new_[11269]_  = ~A267 & \new_[11268]_ ;
  assign \new_[11270]_  = \new_[11269]_  & \new_[11264]_ ;
  assign \new_[11273]_  = A167 & A168;
  assign \new_[11277]_  = A232 & A200;
  assign \new_[11278]_  = A199 & \new_[11277]_ ;
  assign \new_[11279]_  = \new_[11278]_  & \new_[11273]_ ;
  assign \new_[11282]_  = A265 & A233;
  assign \new_[11286]_  = A299 & ~A298;
  assign \new_[11287]_  = A266 & \new_[11286]_ ;
  assign \new_[11288]_  = \new_[11287]_  & \new_[11282]_ ;
  assign \new_[11291]_  = A167 & A168;
  assign \new_[11295]_  = A232 & A200;
  assign \new_[11296]_  = A199 & \new_[11295]_ ;
  assign \new_[11297]_  = \new_[11296]_  & \new_[11291]_ ;
  assign \new_[11300]_  = ~A265 & A233;
  assign \new_[11304]_  = A299 & ~A298;
  assign \new_[11305]_  = ~A266 & \new_[11304]_ ;
  assign \new_[11306]_  = \new_[11305]_  & \new_[11300]_ ;
  assign \new_[11309]_  = A167 & A168;
  assign \new_[11313]_  = ~A232 & A200;
  assign \new_[11314]_  = A199 & \new_[11313]_ ;
  assign \new_[11315]_  = \new_[11314]_  & \new_[11309]_ ;
  assign \new_[11318]_  = A265 & A233;
  assign \new_[11322]_  = A268 & A267;
  assign \new_[11323]_  = ~A266 & \new_[11322]_ ;
  assign \new_[11324]_  = \new_[11323]_  & \new_[11318]_ ;
  assign \new_[11327]_  = A167 & A168;
  assign \new_[11331]_  = ~A232 & A200;
  assign \new_[11332]_  = A199 & \new_[11331]_ ;
  assign \new_[11333]_  = \new_[11332]_  & \new_[11327]_ ;
  assign \new_[11336]_  = A265 & A233;
  assign \new_[11340]_  = A269 & A267;
  assign \new_[11341]_  = ~A266 & \new_[11340]_ ;
  assign \new_[11342]_  = \new_[11341]_  & \new_[11336]_ ;
  assign \new_[11345]_  = A167 & A168;
  assign \new_[11349]_  = ~A233 & A200;
  assign \new_[11350]_  = A199 & \new_[11349]_ ;
  assign \new_[11351]_  = \new_[11350]_  & \new_[11345]_ ;
  assign \new_[11354]_  = A265 & ~A234;
  assign \new_[11358]_  = A299 & ~A298;
  assign \new_[11359]_  = A266 & \new_[11358]_ ;
  assign \new_[11360]_  = \new_[11359]_  & \new_[11354]_ ;
  assign \new_[11363]_  = A167 & A168;
  assign \new_[11367]_  = ~A233 & A200;
  assign \new_[11368]_  = A199 & \new_[11367]_ ;
  assign \new_[11369]_  = \new_[11368]_  & \new_[11363]_ ;
  assign \new_[11372]_  = ~A266 & ~A234;
  assign \new_[11376]_  = A299 & ~A298;
  assign \new_[11377]_  = ~A267 & \new_[11376]_ ;
  assign \new_[11378]_  = \new_[11377]_  & \new_[11372]_ ;
  assign \new_[11381]_  = A167 & A168;
  assign \new_[11385]_  = ~A233 & A200;
  assign \new_[11386]_  = A199 & \new_[11385]_ ;
  assign \new_[11387]_  = \new_[11386]_  & \new_[11381]_ ;
  assign \new_[11390]_  = ~A265 & ~A234;
  assign \new_[11394]_  = A299 & ~A298;
  assign \new_[11395]_  = ~A266 & \new_[11394]_ ;
  assign \new_[11396]_  = \new_[11395]_  & \new_[11390]_ ;
  assign \new_[11399]_  = A167 & A168;
  assign \new_[11403]_  = A232 & A200;
  assign \new_[11404]_  = A199 & \new_[11403]_ ;
  assign \new_[11405]_  = \new_[11404]_  & \new_[11399]_ ;
  assign \new_[11408]_  = A234 & ~A233;
  assign \new_[11412]_  = ~A300 & A298;
  assign \new_[11413]_  = A235 & \new_[11412]_ ;
  assign \new_[11414]_  = \new_[11413]_  & \new_[11408]_ ;
  assign \new_[11417]_  = A167 & A168;
  assign \new_[11421]_  = A232 & A200;
  assign \new_[11422]_  = A199 & \new_[11421]_ ;
  assign \new_[11423]_  = \new_[11422]_  & \new_[11417]_ ;
  assign \new_[11426]_  = A234 & ~A233;
  assign \new_[11430]_  = A299 & A298;
  assign \new_[11431]_  = A235 & \new_[11430]_ ;
  assign \new_[11432]_  = \new_[11431]_  & \new_[11426]_ ;
  assign \new_[11435]_  = A167 & A168;
  assign \new_[11439]_  = A232 & A200;
  assign \new_[11440]_  = A199 & \new_[11439]_ ;
  assign \new_[11441]_  = \new_[11440]_  & \new_[11435]_ ;
  assign \new_[11444]_  = A234 & ~A233;
  assign \new_[11448]_  = ~A299 & ~A298;
  assign \new_[11449]_  = A235 & \new_[11448]_ ;
  assign \new_[11450]_  = \new_[11449]_  & \new_[11444]_ ;
  assign \new_[11453]_  = A167 & A168;
  assign \new_[11457]_  = A232 & A200;
  assign \new_[11458]_  = A199 & \new_[11457]_ ;
  assign \new_[11459]_  = \new_[11458]_  & \new_[11453]_ ;
  assign \new_[11462]_  = A234 & ~A233;
  assign \new_[11466]_  = A266 & ~A265;
  assign \new_[11467]_  = A235 & \new_[11466]_ ;
  assign \new_[11468]_  = \new_[11467]_  & \new_[11462]_ ;
  assign \new_[11471]_  = A167 & A168;
  assign \new_[11475]_  = A232 & A200;
  assign \new_[11476]_  = A199 & \new_[11475]_ ;
  assign \new_[11477]_  = \new_[11476]_  & \new_[11471]_ ;
  assign \new_[11480]_  = A234 & ~A233;
  assign \new_[11484]_  = ~A300 & A298;
  assign \new_[11485]_  = A236 & \new_[11484]_ ;
  assign \new_[11486]_  = \new_[11485]_  & \new_[11480]_ ;
  assign \new_[11489]_  = A167 & A168;
  assign \new_[11493]_  = A232 & A200;
  assign \new_[11494]_  = A199 & \new_[11493]_ ;
  assign \new_[11495]_  = \new_[11494]_  & \new_[11489]_ ;
  assign \new_[11498]_  = A234 & ~A233;
  assign \new_[11502]_  = A299 & A298;
  assign \new_[11503]_  = A236 & \new_[11502]_ ;
  assign \new_[11504]_  = \new_[11503]_  & \new_[11498]_ ;
  assign \new_[11507]_  = A167 & A168;
  assign \new_[11511]_  = A232 & A200;
  assign \new_[11512]_  = A199 & \new_[11511]_ ;
  assign \new_[11513]_  = \new_[11512]_  & \new_[11507]_ ;
  assign \new_[11516]_  = A234 & ~A233;
  assign \new_[11520]_  = ~A299 & ~A298;
  assign \new_[11521]_  = A236 & \new_[11520]_ ;
  assign \new_[11522]_  = \new_[11521]_  & \new_[11516]_ ;
  assign \new_[11525]_  = A167 & A168;
  assign \new_[11529]_  = A232 & A200;
  assign \new_[11530]_  = A199 & \new_[11529]_ ;
  assign \new_[11531]_  = \new_[11530]_  & \new_[11525]_ ;
  assign \new_[11534]_  = A234 & ~A233;
  assign \new_[11538]_  = A266 & ~A265;
  assign \new_[11539]_  = A236 & \new_[11538]_ ;
  assign \new_[11540]_  = \new_[11539]_  & \new_[11534]_ ;
  assign \new_[11543]_  = A167 & A168;
  assign \new_[11547]_  = ~A232 & A200;
  assign \new_[11548]_  = A199 & \new_[11547]_ ;
  assign \new_[11549]_  = \new_[11548]_  & \new_[11543]_ ;
  assign \new_[11552]_  = A265 & ~A233;
  assign \new_[11556]_  = A299 & ~A298;
  assign \new_[11557]_  = A266 & \new_[11556]_ ;
  assign \new_[11558]_  = \new_[11557]_  & \new_[11552]_ ;
  assign \new_[11561]_  = A167 & A168;
  assign \new_[11565]_  = ~A232 & A200;
  assign \new_[11566]_  = A199 & \new_[11565]_ ;
  assign \new_[11567]_  = \new_[11566]_  & \new_[11561]_ ;
  assign \new_[11570]_  = ~A266 & ~A233;
  assign \new_[11574]_  = A299 & ~A298;
  assign \new_[11575]_  = ~A267 & \new_[11574]_ ;
  assign \new_[11576]_  = \new_[11575]_  & \new_[11570]_ ;
  assign \new_[11579]_  = A167 & A168;
  assign \new_[11583]_  = ~A232 & A200;
  assign \new_[11584]_  = A199 & \new_[11583]_ ;
  assign \new_[11585]_  = \new_[11584]_  & \new_[11579]_ ;
  assign \new_[11588]_  = ~A265 & ~A233;
  assign \new_[11592]_  = A299 & ~A298;
  assign \new_[11593]_  = ~A266 & \new_[11592]_ ;
  assign \new_[11594]_  = \new_[11593]_  & \new_[11588]_ ;
  assign \new_[11597]_  = A167 & A168;
  assign \new_[11601]_  = ~A203 & ~A202;
  assign \new_[11602]_  = ~A200 & \new_[11601]_ ;
  assign \new_[11603]_  = \new_[11602]_  & \new_[11597]_ ;
  assign \new_[11606]_  = A233 & ~A232;
  assign \new_[11610]_  = ~A302 & ~A301;
  assign \new_[11611]_  = ~A299 & \new_[11610]_ ;
  assign \new_[11612]_  = \new_[11611]_  & \new_[11606]_ ;
  assign \new_[11615]_  = A167 & A168;
  assign \new_[11619]_  = A232 & ~A201;
  assign \new_[11620]_  = ~A200 & \new_[11619]_ ;
  assign \new_[11621]_  = \new_[11620]_  & \new_[11615]_ ;
  assign \new_[11624]_  = A265 & A233;
  assign \new_[11628]_  = A299 & ~A298;
  assign \new_[11629]_  = ~A267 & \new_[11628]_ ;
  assign \new_[11630]_  = \new_[11629]_  & \new_[11624]_ ;
  assign \new_[11633]_  = A167 & A168;
  assign \new_[11637]_  = A232 & ~A201;
  assign \new_[11638]_  = ~A200 & \new_[11637]_ ;
  assign \new_[11639]_  = \new_[11638]_  & \new_[11633]_ ;
  assign \new_[11642]_  = A265 & A233;
  assign \new_[11646]_  = A299 & ~A298;
  assign \new_[11647]_  = A266 & \new_[11646]_ ;
  assign \new_[11648]_  = \new_[11647]_  & \new_[11642]_ ;
  assign \new_[11651]_  = A167 & A168;
  assign \new_[11655]_  = A232 & ~A201;
  assign \new_[11656]_  = ~A200 & \new_[11655]_ ;
  assign \new_[11657]_  = \new_[11656]_  & \new_[11651]_ ;
  assign \new_[11660]_  = ~A265 & A233;
  assign \new_[11664]_  = A299 & ~A298;
  assign \new_[11665]_  = ~A266 & \new_[11664]_ ;
  assign \new_[11666]_  = \new_[11665]_  & \new_[11660]_ ;
  assign \new_[11669]_  = A167 & A168;
  assign \new_[11673]_  = ~A232 & ~A201;
  assign \new_[11674]_  = ~A200 & \new_[11673]_ ;
  assign \new_[11675]_  = \new_[11674]_  & \new_[11669]_ ;
  assign \new_[11678]_  = A265 & A233;
  assign \new_[11682]_  = A268 & A267;
  assign \new_[11683]_  = ~A266 & \new_[11682]_ ;
  assign \new_[11684]_  = \new_[11683]_  & \new_[11678]_ ;
  assign \new_[11687]_  = A167 & A168;
  assign \new_[11691]_  = ~A232 & ~A201;
  assign \new_[11692]_  = ~A200 & \new_[11691]_ ;
  assign \new_[11693]_  = \new_[11692]_  & \new_[11687]_ ;
  assign \new_[11696]_  = A265 & A233;
  assign \new_[11700]_  = A269 & A267;
  assign \new_[11701]_  = ~A266 & \new_[11700]_ ;
  assign \new_[11702]_  = \new_[11701]_  & \new_[11696]_ ;
  assign \new_[11705]_  = A167 & A168;
  assign \new_[11709]_  = ~A233 & ~A201;
  assign \new_[11710]_  = ~A200 & \new_[11709]_ ;
  assign \new_[11711]_  = \new_[11710]_  & \new_[11705]_ ;
  assign \new_[11714]_  = A265 & ~A234;
  assign \new_[11718]_  = A299 & ~A298;
  assign \new_[11719]_  = A266 & \new_[11718]_ ;
  assign \new_[11720]_  = \new_[11719]_  & \new_[11714]_ ;
  assign \new_[11723]_  = A167 & A168;
  assign \new_[11727]_  = ~A233 & ~A201;
  assign \new_[11728]_  = ~A200 & \new_[11727]_ ;
  assign \new_[11729]_  = \new_[11728]_  & \new_[11723]_ ;
  assign \new_[11732]_  = ~A266 & ~A234;
  assign \new_[11736]_  = A299 & ~A298;
  assign \new_[11737]_  = ~A267 & \new_[11736]_ ;
  assign \new_[11738]_  = \new_[11737]_  & \new_[11732]_ ;
  assign \new_[11741]_  = A167 & A168;
  assign \new_[11745]_  = ~A233 & ~A201;
  assign \new_[11746]_  = ~A200 & \new_[11745]_ ;
  assign \new_[11747]_  = \new_[11746]_  & \new_[11741]_ ;
  assign \new_[11750]_  = ~A265 & ~A234;
  assign \new_[11754]_  = A299 & ~A298;
  assign \new_[11755]_  = ~A266 & \new_[11754]_ ;
  assign \new_[11756]_  = \new_[11755]_  & \new_[11750]_ ;
  assign \new_[11759]_  = A167 & A168;
  assign \new_[11763]_  = A232 & ~A201;
  assign \new_[11764]_  = ~A200 & \new_[11763]_ ;
  assign \new_[11765]_  = \new_[11764]_  & \new_[11759]_ ;
  assign \new_[11768]_  = A234 & ~A233;
  assign \new_[11772]_  = ~A300 & A298;
  assign \new_[11773]_  = A235 & \new_[11772]_ ;
  assign \new_[11774]_  = \new_[11773]_  & \new_[11768]_ ;
  assign \new_[11777]_  = A167 & A168;
  assign \new_[11781]_  = A232 & ~A201;
  assign \new_[11782]_  = ~A200 & \new_[11781]_ ;
  assign \new_[11783]_  = \new_[11782]_  & \new_[11777]_ ;
  assign \new_[11786]_  = A234 & ~A233;
  assign \new_[11790]_  = A299 & A298;
  assign \new_[11791]_  = A235 & \new_[11790]_ ;
  assign \new_[11792]_  = \new_[11791]_  & \new_[11786]_ ;
  assign \new_[11795]_  = A167 & A168;
  assign \new_[11799]_  = A232 & ~A201;
  assign \new_[11800]_  = ~A200 & \new_[11799]_ ;
  assign \new_[11801]_  = \new_[11800]_  & \new_[11795]_ ;
  assign \new_[11804]_  = A234 & ~A233;
  assign \new_[11808]_  = ~A299 & ~A298;
  assign \new_[11809]_  = A235 & \new_[11808]_ ;
  assign \new_[11810]_  = \new_[11809]_  & \new_[11804]_ ;
  assign \new_[11813]_  = A167 & A168;
  assign \new_[11817]_  = A232 & ~A201;
  assign \new_[11818]_  = ~A200 & \new_[11817]_ ;
  assign \new_[11819]_  = \new_[11818]_  & \new_[11813]_ ;
  assign \new_[11822]_  = A234 & ~A233;
  assign \new_[11826]_  = A266 & ~A265;
  assign \new_[11827]_  = A235 & \new_[11826]_ ;
  assign \new_[11828]_  = \new_[11827]_  & \new_[11822]_ ;
  assign \new_[11831]_  = A167 & A168;
  assign \new_[11835]_  = A232 & ~A201;
  assign \new_[11836]_  = ~A200 & \new_[11835]_ ;
  assign \new_[11837]_  = \new_[11836]_  & \new_[11831]_ ;
  assign \new_[11840]_  = A234 & ~A233;
  assign \new_[11844]_  = ~A300 & A298;
  assign \new_[11845]_  = A236 & \new_[11844]_ ;
  assign \new_[11846]_  = \new_[11845]_  & \new_[11840]_ ;
  assign \new_[11849]_  = A167 & A168;
  assign \new_[11853]_  = A232 & ~A201;
  assign \new_[11854]_  = ~A200 & \new_[11853]_ ;
  assign \new_[11855]_  = \new_[11854]_  & \new_[11849]_ ;
  assign \new_[11858]_  = A234 & ~A233;
  assign \new_[11862]_  = A299 & A298;
  assign \new_[11863]_  = A236 & \new_[11862]_ ;
  assign \new_[11864]_  = \new_[11863]_  & \new_[11858]_ ;
  assign \new_[11867]_  = A167 & A168;
  assign \new_[11871]_  = A232 & ~A201;
  assign \new_[11872]_  = ~A200 & \new_[11871]_ ;
  assign \new_[11873]_  = \new_[11872]_  & \new_[11867]_ ;
  assign \new_[11876]_  = A234 & ~A233;
  assign \new_[11880]_  = ~A299 & ~A298;
  assign \new_[11881]_  = A236 & \new_[11880]_ ;
  assign \new_[11882]_  = \new_[11881]_  & \new_[11876]_ ;
  assign \new_[11885]_  = A167 & A168;
  assign \new_[11889]_  = A232 & ~A201;
  assign \new_[11890]_  = ~A200 & \new_[11889]_ ;
  assign \new_[11891]_  = \new_[11890]_  & \new_[11885]_ ;
  assign \new_[11894]_  = A234 & ~A233;
  assign \new_[11898]_  = A266 & ~A265;
  assign \new_[11899]_  = A236 & \new_[11898]_ ;
  assign \new_[11900]_  = \new_[11899]_  & \new_[11894]_ ;
  assign \new_[11903]_  = A167 & A168;
  assign \new_[11907]_  = ~A232 & ~A201;
  assign \new_[11908]_  = ~A200 & \new_[11907]_ ;
  assign \new_[11909]_  = \new_[11908]_  & \new_[11903]_ ;
  assign \new_[11912]_  = A265 & ~A233;
  assign \new_[11916]_  = A299 & ~A298;
  assign \new_[11917]_  = A266 & \new_[11916]_ ;
  assign \new_[11918]_  = \new_[11917]_  & \new_[11912]_ ;
  assign \new_[11921]_  = A167 & A168;
  assign \new_[11925]_  = ~A232 & ~A201;
  assign \new_[11926]_  = ~A200 & \new_[11925]_ ;
  assign \new_[11927]_  = \new_[11926]_  & \new_[11921]_ ;
  assign \new_[11930]_  = ~A266 & ~A233;
  assign \new_[11934]_  = A299 & ~A298;
  assign \new_[11935]_  = ~A267 & \new_[11934]_ ;
  assign \new_[11936]_  = \new_[11935]_  & \new_[11930]_ ;
  assign \new_[11939]_  = A167 & A168;
  assign \new_[11943]_  = ~A232 & ~A201;
  assign \new_[11944]_  = ~A200 & \new_[11943]_ ;
  assign \new_[11945]_  = \new_[11944]_  & \new_[11939]_ ;
  assign \new_[11948]_  = ~A265 & ~A233;
  assign \new_[11952]_  = A299 & ~A298;
  assign \new_[11953]_  = ~A266 & \new_[11952]_ ;
  assign \new_[11954]_  = \new_[11953]_  & \new_[11948]_ ;
  assign \new_[11957]_  = A167 & A168;
  assign \new_[11961]_  = A232 & ~A200;
  assign \new_[11962]_  = ~A199 & \new_[11961]_ ;
  assign \new_[11963]_  = \new_[11962]_  & \new_[11957]_ ;
  assign \new_[11966]_  = A265 & A233;
  assign \new_[11970]_  = A299 & ~A298;
  assign \new_[11971]_  = ~A267 & \new_[11970]_ ;
  assign \new_[11972]_  = \new_[11971]_  & \new_[11966]_ ;
  assign \new_[11975]_  = A167 & A168;
  assign \new_[11979]_  = A232 & ~A200;
  assign \new_[11980]_  = ~A199 & \new_[11979]_ ;
  assign \new_[11981]_  = \new_[11980]_  & \new_[11975]_ ;
  assign \new_[11984]_  = A265 & A233;
  assign \new_[11988]_  = A299 & ~A298;
  assign \new_[11989]_  = A266 & \new_[11988]_ ;
  assign \new_[11990]_  = \new_[11989]_  & \new_[11984]_ ;
  assign \new_[11993]_  = A167 & A168;
  assign \new_[11997]_  = A232 & ~A200;
  assign \new_[11998]_  = ~A199 & \new_[11997]_ ;
  assign \new_[11999]_  = \new_[11998]_  & \new_[11993]_ ;
  assign \new_[12002]_  = ~A265 & A233;
  assign \new_[12006]_  = A299 & ~A298;
  assign \new_[12007]_  = ~A266 & \new_[12006]_ ;
  assign \new_[12008]_  = \new_[12007]_  & \new_[12002]_ ;
  assign \new_[12011]_  = A167 & A168;
  assign \new_[12015]_  = ~A232 & ~A200;
  assign \new_[12016]_  = ~A199 & \new_[12015]_ ;
  assign \new_[12017]_  = \new_[12016]_  & \new_[12011]_ ;
  assign \new_[12020]_  = A265 & A233;
  assign \new_[12024]_  = A268 & A267;
  assign \new_[12025]_  = ~A266 & \new_[12024]_ ;
  assign \new_[12026]_  = \new_[12025]_  & \new_[12020]_ ;
  assign \new_[12029]_  = A167 & A168;
  assign \new_[12033]_  = ~A232 & ~A200;
  assign \new_[12034]_  = ~A199 & \new_[12033]_ ;
  assign \new_[12035]_  = \new_[12034]_  & \new_[12029]_ ;
  assign \new_[12038]_  = A265 & A233;
  assign \new_[12042]_  = A269 & A267;
  assign \new_[12043]_  = ~A266 & \new_[12042]_ ;
  assign \new_[12044]_  = \new_[12043]_  & \new_[12038]_ ;
  assign \new_[12047]_  = A167 & A168;
  assign \new_[12051]_  = ~A233 & ~A200;
  assign \new_[12052]_  = ~A199 & \new_[12051]_ ;
  assign \new_[12053]_  = \new_[12052]_  & \new_[12047]_ ;
  assign \new_[12056]_  = A265 & ~A234;
  assign \new_[12060]_  = A299 & ~A298;
  assign \new_[12061]_  = A266 & \new_[12060]_ ;
  assign \new_[12062]_  = \new_[12061]_  & \new_[12056]_ ;
  assign \new_[12065]_  = A167 & A168;
  assign \new_[12069]_  = ~A233 & ~A200;
  assign \new_[12070]_  = ~A199 & \new_[12069]_ ;
  assign \new_[12071]_  = \new_[12070]_  & \new_[12065]_ ;
  assign \new_[12074]_  = ~A266 & ~A234;
  assign \new_[12078]_  = A299 & ~A298;
  assign \new_[12079]_  = ~A267 & \new_[12078]_ ;
  assign \new_[12080]_  = \new_[12079]_  & \new_[12074]_ ;
  assign \new_[12083]_  = A167 & A168;
  assign \new_[12087]_  = ~A233 & ~A200;
  assign \new_[12088]_  = ~A199 & \new_[12087]_ ;
  assign \new_[12089]_  = \new_[12088]_  & \new_[12083]_ ;
  assign \new_[12092]_  = ~A265 & ~A234;
  assign \new_[12096]_  = A299 & ~A298;
  assign \new_[12097]_  = ~A266 & \new_[12096]_ ;
  assign \new_[12098]_  = \new_[12097]_  & \new_[12092]_ ;
  assign \new_[12101]_  = A167 & A168;
  assign \new_[12105]_  = A232 & ~A200;
  assign \new_[12106]_  = ~A199 & \new_[12105]_ ;
  assign \new_[12107]_  = \new_[12106]_  & \new_[12101]_ ;
  assign \new_[12110]_  = A234 & ~A233;
  assign \new_[12114]_  = ~A300 & A298;
  assign \new_[12115]_  = A235 & \new_[12114]_ ;
  assign \new_[12116]_  = \new_[12115]_  & \new_[12110]_ ;
  assign \new_[12119]_  = A167 & A168;
  assign \new_[12123]_  = A232 & ~A200;
  assign \new_[12124]_  = ~A199 & \new_[12123]_ ;
  assign \new_[12125]_  = \new_[12124]_  & \new_[12119]_ ;
  assign \new_[12128]_  = A234 & ~A233;
  assign \new_[12132]_  = A299 & A298;
  assign \new_[12133]_  = A235 & \new_[12132]_ ;
  assign \new_[12134]_  = \new_[12133]_  & \new_[12128]_ ;
  assign \new_[12137]_  = A167 & A168;
  assign \new_[12141]_  = A232 & ~A200;
  assign \new_[12142]_  = ~A199 & \new_[12141]_ ;
  assign \new_[12143]_  = \new_[12142]_  & \new_[12137]_ ;
  assign \new_[12146]_  = A234 & ~A233;
  assign \new_[12150]_  = ~A299 & ~A298;
  assign \new_[12151]_  = A235 & \new_[12150]_ ;
  assign \new_[12152]_  = \new_[12151]_  & \new_[12146]_ ;
  assign \new_[12155]_  = A167 & A168;
  assign \new_[12159]_  = A232 & ~A200;
  assign \new_[12160]_  = ~A199 & \new_[12159]_ ;
  assign \new_[12161]_  = \new_[12160]_  & \new_[12155]_ ;
  assign \new_[12164]_  = A234 & ~A233;
  assign \new_[12168]_  = A266 & ~A265;
  assign \new_[12169]_  = A235 & \new_[12168]_ ;
  assign \new_[12170]_  = \new_[12169]_  & \new_[12164]_ ;
  assign \new_[12173]_  = A167 & A168;
  assign \new_[12177]_  = A232 & ~A200;
  assign \new_[12178]_  = ~A199 & \new_[12177]_ ;
  assign \new_[12179]_  = \new_[12178]_  & \new_[12173]_ ;
  assign \new_[12182]_  = A234 & ~A233;
  assign \new_[12186]_  = ~A300 & A298;
  assign \new_[12187]_  = A236 & \new_[12186]_ ;
  assign \new_[12188]_  = \new_[12187]_  & \new_[12182]_ ;
  assign \new_[12191]_  = A167 & A168;
  assign \new_[12195]_  = A232 & ~A200;
  assign \new_[12196]_  = ~A199 & \new_[12195]_ ;
  assign \new_[12197]_  = \new_[12196]_  & \new_[12191]_ ;
  assign \new_[12200]_  = A234 & ~A233;
  assign \new_[12204]_  = A299 & A298;
  assign \new_[12205]_  = A236 & \new_[12204]_ ;
  assign \new_[12206]_  = \new_[12205]_  & \new_[12200]_ ;
  assign \new_[12209]_  = A167 & A168;
  assign \new_[12213]_  = A232 & ~A200;
  assign \new_[12214]_  = ~A199 & \new_[12213]_ ;
  assign \new_[12215]_  = \new_[12214]_  & \new_[12209]_ ;
  assign \new_[12218]_  = A234 & ~A233;
  assign \new_[12222]_  = ~A299 & ~A298;
  assign \new_[12223]_  = A236 & \new_[12222]_ ;
  assign \new_[12224]_  = \new_[12223]_  & \new_[12218]_ ;
  assign \new_[12227]_  = A167 & A168;
  assign \new_[12231]_  = A232 & ~A200;
  assign \new_[12232]_  = ~A199 & \new_[12231]_ ;
  assign \new_[12233]_  = \new_[12232]_  & \new_[12227]_ ;
  assign \new_[12236]_  = A234 & ~A233;
  assign \new_[12240]_  = A266 & ~A265;
  assign \new_[12241]_  = A236 & \new_[12240]_ ;
  assign \new_[12242]_  = \new_[12241]_  & \new_[12236]_ ;
  assign \new_[12245]_  = A167 & A168;
  assign \new_[12249]_  = ~A232 & ~A200;
  assign \new_[12250]_  = ~A199 & \new_[12249]_ ;
  assign \new_[12251]_  = \new_[12250]_  & \new_[12245]_ ;
  assign \new_[12254]_  = A265 & ~A233;
  assign \new_[12258]_  = A299 & ~A298;
  assign \new_[12259]_  = A266 & \new_[12258]_ ;
  assign \new_[12260]_  = \new_[12259]_  & \new_[12254]_ ;
  assign \new_[12263]_  = A167 & A168;
  assign \new_[12267]_  = ~A232 & ~A200;
  assign \new_[12268]_  = ~A199 & \new_[12267]_ ;
  assign \new_[12269]_  = \new_[12268]_  & \new_[12263]_ ;
  assign \new_[12272]_  = ~A266 & ~A233;
  assign \new_[12276]_  = A299 & ~A298;
  assign \new_[12277]_  = ~A267 & \new_[12276]_ ;
  assign \new_[12278]_  = \new_[12277]_  & \new_[12272]_ ;
  assign \new_[12281]_  = A167 & A168;
  assign \new_[12285]_  = ~A232 & ~A200;
  assign \new_[12286]_  = ~A199 & \new_[12285]_ ;
  assign \new_[12287]_  = \new_[12286]_  & \new_[12281]_ ;
  assign \new_[12290]_  = ~A265 & ~A233;
  assign \new_[12294]_  = A299 & ~A298;
  assign \new_[12295]_  = ~A266 & \new_[12294]_ ;
  assign \new_[12296]_  = \new_[12295]_  & \new_[12290]_ ;
  assign \new_[12299]_  = ~A167 & A170;
  assign \new_[12303]_  = A200 & ~A199;
  assign \new_[12304]_  = ~A166 & \new_[12303]_ ;
  assign \new_[12305]_  = \new_[12304]_  & \new_[12299]_ ;
  assign \new_[12308]_  = A233 & ~A232;
  assign \new_[12312]_  = ~A302 & ~A301;
  assign \new_[12313]_  = ~A299 & \new_[12312]_ ;
  assign \new_[12314]_  = \new_[12313]_  & \new_[12308]_ ;
  assign \new_[12317]_  = ~A168 & A170;
  assign \new_[12321]_  = ~A199 & A166;
  assign \new_[12322]_  = A167 & \new_[12321]_ ;
  assign \new_[12323]_  = \new_[12322]_  & \new_[12317]_ ;
  assign \new_[12326]_  = ~A232 & A200;
  assign \new_[12330]_  = ~A300 & ~A299;
  assign \new_[12331]_  = A233 & \new_[12330]_ ;
  assign \new_[12332]_  = \new_[12331]_  & \new_[12326]_ ;
  assign \new_[12335]_  = ~A168 & A170;
  assign \new_[12339]_  = ~A199 & A166;
  assign \new_[12340]_  = A167 & \new_[12339]_ ;
  assign \new_[12341]_  = \new_[12340]_  & \new_[12335]_ ;
  assign \new_[12344]_  = ~A232 & A200;
  assign \new_[12348]_  = A299 & A298;
  assign \new_[12349]_  = A233 & \new_[12348]_ ;
  assign \new_[12350]_  = \new_[12349]_  & \new_[12344]_ ;
  assign \new_[12353]_  = ~A168 & A170;
  assign \new_[12357]_  = ~A199 & A166;
  assign \new_[12358]_  = A167 & \new_[12357]_ ;
  assign \new_[12359]_  = \new_[12358]_  & \new_[12353]_ ;
  assign \new_[12362]_  = ~A232 & A200;
  assign \new_[12366]_  = ~A299 & ~A298;
  assign \new_[12367]_  = A233 & \new_[12366]_ ;
  assign \new_[12368]_  = \new_[12367]_  & \new_[12362]_ ;
  assign \new_[12371]_  = ~A168 & A170;
  assign \new_[12375]_  = ~A199 & A166;
  assign \new_[12376]_  = A167 & \new_[12375]_ ;
  assign \new_[12377]_  = \new_[12376]_  & \new_[12371]_ ;
  assign \new_[12380]_  = ~A232 & A200;
  assign \new_[12384]_  = A266 & ~A265;
  assign \new_[12385]_  = A233 & \new_[12384]_ ;
  assign \new_[12386]_  = \new_[12385]_  & \new_[12380]_ ;
  assign \new_[12389]_  = ~A168 & ~A170;
  assign \new_[12393]_  = ~A199 & ~A166;
  assign \new_[12394]_  = A167 & \new_[12393]_ ;
  assign \new_[12395]_  = \new_[12394]_  & \new_[12389]_ ;
  assign \new_[12398]_  = ~A232 & A200;
  assign \new_[12402]_  = ~A300 & ~A299;
  assign \new_[12403]_  = A233 & \new_[12402]_ ;
  assign \new_[12404]_  = \new_[12403]_  & \new_[12398]_ ;
  assign \new_[12407]_  = ~A168 & ~A170;
  assign \new_[12411]_  = ~A199 & ~A166;
  assign \new_[12412]_  = A167 & \new_[12411]_ ;
  assign \new_[12413]_  = \new_[12412]_  & \new_[12407]_ ;
  assign \new_[12416]_  = ~A232 & A200;
  assign \new_[12420]_  = A299 & A298;
  assign \new_[12421]_  = A233 & \new_[12420]_ ;
  assign \new_[12422]_  = \new_[12421]_  & \new_[12416]_ ;
  assign \new_[12425]_  = ~A168 & ~A170;
  assign \new_[12429]_  = ~A199 & ~A166;
  assign \new_[12430]_  = A167 & \new_[12429]_ ;
  assign \new_[12431]_  = \new_[12430]_  & \new_[12425]_ ;
  assign \new_[12434]_  = ~A232 & A200;
  assign \new_[12438]_  = ~A299 & ~A298;
  assign \new_[12439]_  = A233 & \new_[12438]_ ;
  assign \new_[12440]_  = \new_[12439]_  & \new_[12434]_ ;
  assign \new_[12443]_  = ~A168 & ~A170;
  assign \new_[12447]_  = ~A199 & ~A166;
  assign \new_[12448]_  = A167 & \new_[12447]_ ;
  assign \new_[12449]_  = \new_[12448]_  & \new_[12443]_ ;
  assign \new_[12452]_  = ~A232 & A200;
  assign \new_[12456]_  = A266 & ~A265;
  assign \new_[12457]_  = A233 & \new_[12456]_ ;
  assign \new_[12458]_  = \new_[12457]_  & \new_[12452]_ ;
  assign \new_[12461]_  = ~A168 & ~A170;
  assign \new_[12465]_  = ~A199 & A166;
  assign \new_[12466]_  = ~A167 & \new_[12465]_ ;
  assign \new_[12467]_  = \new_[12466]_  & \new_[12461]_ ;
  assign \new_[12470]_  = ~A232 & A200;
  assign \new_[12474]_  = ~A300 & ~A299;
  assign \new_[12475]_  = A233 & \new_[12474]_ ;
  assign \new_[12476]_  = \new_[12475]_  & \new_[12470]_ ;
  assign \new_[12479]_  = ~A168 & ~A170;
  assign \new_[12483]_  = ~A199 & A166;
  assign \new_[12484]_  = ~A167 & \new_[12483]_ ;
  assign \new_[12485]_  = \new_[12484]_  & \new_[12479]_ ;
  assign \new_[12488]_  = ~A232 & A200;
  assign \new_[12492]_  = A299 & A298;
  assign \new_[12493]_  = A233 & \new_[12492]_ ;
  assign \new_[12494]_  = \new_[12493]_  & \new_[12488]_ ;
  assign \new_[12497]_  = ~A168 & ~A170;
  assign \new_[12501]_  = ~A199 & A166;
  assign \new_[12502]_  = ~A167 & \new_[12501]_ ;
  assign \new_[12503]_  = \new_[12502]_  & \new_[12497]_ ;
  assign \new_[12506]_  = ~A232 & A200;
  assign \new_[12510]_  = ~A299 & ~A298;
  assign \new_[12511]_  = A233 & \new_[12510]_ ;
  assign \new_[12512]_  = \new_[12511]_  & \new_[12506]_ ;
  assign \new_[12515]_  = ~A168 & ~A170;
  assign \new_[12519]_  = ~A199 & A166;
  assign \new_[12520]_  = ~A167 & \new_[12519]_ ;
  assign \new_[12521]_  = \new_[12520]_  & \new_[12515]_ ;
  assign \new_[12524]_  = ~A232 & A200;
  assign \new_[12528]_  = A266 & ~A265;
  assign \new_[12529]_  = A233 & \new_[12528]_ ;
  assign \new_[12530]_  = \new_[12529]_  & \new_[12524]_ ;
  assign \new_[12533]_  = ~A168 & A169;
  assign \new_[12537]_  = ~A199 & ~A166;
  assign \new_[12538]_  = A167 & \new_[12537]_ ;
  assign \new_[12539]_  = \new_[12538]_  & \new_[12533]_ ;
  assign \new_[12542]_  = ~A232 & A200;
  assign \new_[12546]_  = ~A300 & ~A299;
  assign \new_[12547]_  = A233 & \new_[12546]_ ;
  assign \new_[12548]_  = \new_[12547]_  & \new_[12542]_ ;
  assign \new_[12551]_  = ~A168 & A169;
  assign \new_[12555]_  = ~A199 & ~A166;
  assign \new_[12556]_  = A167 & \new_[12555]_ ;
  assign \new_[12557]_  = \new_[12556]_  & \new_[12551]_ ;
  assign \new_[12560]_  = ~A232 & A200;
  assign \new_[12564]_  = A299 & A298;
  assign \new_[12565]_  = A233 & \new_[12564]_ ;
  assign \new_[12566]_  = \new_[12565]_  & \new_[12560]_ ;
  assign \new_[12569]_  = ~A168 & A169;
  assign \new_[12573]_  = ~A199 & ~A166;
  assign \new_[12574]_  = A167 & \new_[12573]_ ;
  assign \new_[12575]_  = \new_[12574]_  & \new_[12569]_ ;
  assign \new_[12578]_  = ~A232 & A200;
  assign \new_[12582]_  = ~A299 & ~A298;
  assign \new_[12583]_  = A233 & \new_[12582]_ ;
  assign \new_[12584]_  = \new_[12583]_  & \new_[12578]_ ;
  assign \new_[12587]_  = ~A168 & A169;
  assign \new_[12591]_  = ~A199 & ~A166;
  assign \new_[12592]_  = A167 & \new_[12591]_ ;
  assign \new_[12593]_  = \new_[12592]_  & \new_[12587]_ ;
  assign \new_[12596]_  = ~A232 & A200;
  assign \new_[12600]_  = A266 & ~A265;
  assign \new_[12601]_  = A233 & \new_[12600]_ ;
  assign \new_[12602]_  = \new_[12601]_  & \new_[12596]_ ;
  assign \new_[12605]_  = ~A168 & A169;
  assign \new_[12609]_  = ~A199 & A166;
  assign \new_[12610]_  = ~A167 & \new_[12609]_ ;
  assign \new_[12611]_  = \new_[12610]_  & \new_[12605]_ ;
  assign \new_[12614]_  = ~A232 & A200;
  assign \new_[12618]_  = ~A300 & ~A299;
  assign \new_[12619]_  = A233 & \new_[12618]_ ;
  assign \new_[12620]_  = \new_[12619]_  & \new_[12614]_ ;
  assign \new_[12623]_  = ~A168 & A169;
  assign \new_[12627]_  = ~A199 & A166;
  assign \new_[12628]_  = ~A167 & \new_[12627]_ ;
  assign \new_[12629]_  = \new_[12628]_  & \new_[12623]_ ;
  assign \new_[12632]_  = ~A232 & A200;
  assign \new_[12636]_  = A299 & A298;
  assign \new_[12637]_  = A233 & \new_[12636]_ ;
  assign \new_[12638]_  = \new_[12637]_  & \new_[12632]_ ;
  assign \new_[12641]_  = ~A168 & A169;
  assign \new_[12645]_  = ~A199 & A166;
  assign \new_[12646]_  = ~A167 & \new_[12645]_ ;
  assign \new_[12647]_  = \new_[12646]_  & \new_[12641]_ ;
  assign \new_[12650]_  = ~A232 & A200;
  assign \new_[12654]_  = ~A299 & ~A298;
  assign \new_[12655]_  = A233 & \new_[12654]_ ;
  assign \new_[12656]_  = \new_[12655]_  & \new_[12650]_ ;
  assign \new_[12659]_  = ~A168 & A169;
  assign \new_[12663]_  = ~A199 & A166;
  assign \new_[12664]_  = ~A167 & \new_[12663]_ ;
  assign \new_[12665]_  = \new_[12664]_  & \new_[12659]_ ;
  assign \new_[12668]_  = ~A232 & A200;
  assign \new_[12672]_  = A266 & ~A265;
  assign \new_[12673]_  = A233 & \new_[12672]_ ;
  assign \new_[12674]_  = \new_[12673]_  & \new_[12668]_ ;
  assign \new_[12677]_  = A169 & ~A170;
  assign \new_[12681]_  = A199 & A166;
  assign \new_[12682]_  = A167 & \new_[12681]_ ;
  assign \new_[12683]_  = \new_[12682]_  & \new_[12677]_ ;
  assign \new_[12686]_  = ~A232 & A200;
  assign \new_[12690]_  = ~A300 & ~A299;
  assign \new_[12691]_  = A233 & \new_[12690]_ ;
  assign \new_[12692]_  = \new_[12691]_  & \new_[12686]_ ;
  assign \new_[12695]_  = A169 & ~A170;
  assign \new_[12699]_  = A199 & A166;
  assign \new_[12700]_  = A167 & \new_[12699]_ ;
  assign \new_[12701]_  = \new_[12700]_  & \new_[12695]_ ;
  assign \new_[12704]_  = ~A232 & A200;
  assign \new_[12708]_  = A299 & A298;
  assign \new_[12709]_  = A233 & \new_[12708]_ ;
  assign \new_[12710]_  = \new_[12709]_  & \new_[12704]_ ;
  assign \new_[12713]_  = A169 & ~A170;
  assign \new_[12717]_  = A199 & A166;
  assign \new_[12718]_  = A167 & \new_[12717]_ ;
  assign \new_[12719]_  = \new_[12718]_  & \new_[12713]_ ;
  assign \new_[12722]_  = ~A232 & A200;
  assign \new_[12726]_  = ~A299 & ~A298;
  assign \new_[12727]_  = A233 & \new_[12726]_ ;
  assign \new_[12728]_  = \new_[12727]_  & \new_[12722]_ ;
  assign \new_[12731]_  = A169 & ~A170;
  assign \new_[12735]_  = A199 & A166;
  assign \new_[12736]_  = A167 & \new_[12735]_ ;
  assign \new_[12737]_  = \new_[12736]_  & \new_[12731]_ ;
  assign \new_[12740]_  = ~A232 & A200;
  assign \new_[12744]_  = A266 & ~A265;
  assign \new_[12745]_  = A233 & \new_[12744]_ ;
  assign \new_[12746]_  = \new_[12745]_  & \new_[12740]_ ;
  assign \new_[12749]_  = A169 & ~A170;
  assign \new_[12753]_  = ~A200 & A166;
  assign \new_[12754]_  = A167 & \new_[12753]_ ;
  assign \new_[12755]_  = \new_[12754]_  & \new_[12749]_ ;
  assign \new_[12758]_  = ~A232 & ~A201;
  assign \new_[12762]_  = ~A300 & ~A299;
  assign \new_[12763]_  = A233 & \new_[12762]_ ;
  assign \new_[12764]_  = \new_[12763]_  & \new_[12758]_ ;
  assign \new_[12767]_  = A169 & ~A170;
  assign \new_[12771]_  = ~A200 & A166;
  assign \new_[12772]_  = A167 & \new_[12771]_ ;
  assign \new_[12773]_  = \new_[12772]_  & \new_[12767]_ ;
  assign \new_[12776]_  = ~A232 & ~A201;
  assign \new_[12780]_  = A299 & A298;
  assign \new_[12781]_  = A233 & \new_[12780]_ ;
  assign \new_[12782]_  = \new_[12781]_  & \new_[12776]_ ;
  assign \new_[12785]_  = A169 & ~A170;
  assign \new_[12789]_  = ~A200 & A166;
  assign \new_[12790]_  = A167 & \new_[12789]_ ;
  assign \new_[12791]_  = \new_[12790]_  & \new_[12785]_ ;
  assign \new_[12794]_  = ~A232 & ~A201;
  assign \new_[12798]_  = ~A299 & ~A298;
  assign \new_[12799]_  = A233 & \new_[12798]_ ;
  assign \new_[12800]_  = \new_[12799]_  & \new_[12794]_ ;
  assign \new_[12803]_  = A169 & ~A170;
  assign \new_[12807]_  = ~A200 & A166;
  assign \new_[12808]_  = A167 & \new_[12807]_ ;
  assign \new_[12809]_  = \new_[12808]_  & \new_[12803]_ ;
  assign \new_[12812]_  = ~A232 & ~A201;
  assign \new_[12816]_  = A266 & ~A265;
  assign \new_[12817]_  = A233 & \new_[12816]_ ;
  assign \new_[12818]_  = \new_[12817]_  & \new_[12812]_ ;
  assign \new_[12821]_  = A169 & ~A170;
  assign \new_[12825]_  = ~A199 & A166;
  assign \new_[12826]_  = A167 & \new_[12825]_ ;
  assign \new_[12827]_  = \new_[12826]_  & \new_[12821]_ ;
  assign \new_[12830]_  = ~A232 & ~A200;
  assign \new_[12834]_  = ~A300 & ~A299;
  assign \new_[12835]_  = A233 & \new_[12834]_ ;
  assign \new_[12836]_  = \new_[12835]_  & \new_[12830]_ ;
  assign \new_[12839]_  = A169 & ~A170;
  assign \new_[12843]_  = ~A199 & A166;
  assign \new_[12844]_  = A167 & \new_[12843]_ ;
  assign \new_[12845]_  = \new_[12844]_  & \new_[12839]_ ;
  assign \new_[12848]_  = ~A232 & ~A200;
  assign \new_[12852]_  = A299 & A298;
  assign \new_[12853]_  = A233 & \new_[12852]_ ;
  assign \new_[12854]_  = \new_[12853]_  & \new_[12848]_ ;
  assign \new_[12857]_  = A169 & ~A170;
  assign \new_[12861]_  = ~A199 & A166;
  assign \new_[12862]_  = A167 & \new_[12861]_ ;
  assign \new_[12863]_  = \new_[12862]_  & \new_[12857]_ ;
  assign \new_[12866]_  = ~A232 & ~A200;
  assign \new_[12870]_  = ~A299 & ~A298;
  assign \new_[12871]_  = A233 & \new_[12870]_ ;
  assign \new_[12872]_  = \new_[12871]_  & \new_[12866]_ ;
  assign \new_[12875]_  = A169 & ~A170;
  assign \new_[12879]_  = ~A199 & A166;
  assign \new_[12880]_  = A167 & \new_[12879]_ ;
  assign \new_[12881]_  = \new_[12880]_  & \new_[12875]_ ;
  assign \new_[12884]_  = ~A232 & ~A200;
  assign \new_[12888]_  = A266 & ~A265;
  assign \new_[12889]_  = A233 & \new_[12888]_ ;
  assign \new_[12890]_  = \new_[12889]_  & \new_[12884]_ ;
  assign \new_[12893]_  = A169 & ~A170;
  assign \new_[12897]_  = A199 & ~A166;
  assign \new_[12898]_  = ~A167 & \new_[12897]_ ;
  assign \new_[12899]_  = \new_[12898]_  & \new_[12893]_ ;
  assign \new_[12902]_  = ~A232 & A200;
  assign \new_[12906]_  = ~A300 & ~A299;
  assign \new_[12907]_  = A233 & \new_[12906]_ ;
  assign \new_[12908]_  = \new_[12907]_  & \new_[12902]_ ;
  assign \new_[12911]_  = A169 & ~A170;
  assign \new_[12915]_  = A199 & ~A166;
  assign \new_[12916]_  = ~A167 & \new_[12915]_ ;
  assign \new_[12917]_  = \new_[12916]_  & \new_[12911]_ ;
  assign \new_[12920]_  = ~A232 & A200;
  assign \new_[12924]_  = A299 & A298;
  assign \new_[12925]_  = A233 & \new_[12924]_ ;
  assign \new_[12926]_  = \new_[12925]_  & \new_[12920]_ ;
  assign \new_[12929]_  = A169 & ~A170;
  assign \new_[12933]_  = A199 & ~A166;
  assign \new_[12934]_  = ~A167 & \new_[12933]_ ;
  assign \new_[12935]_  = \new_[12934]_  & \new_[12929]_ ;
  assign \new_[12938]_  = ~A232 & A200;
  assign \new_[12942]_  = ~A299 & ~A298;
  assign \new_[12943]_  = A233 & \new_[12942]_ ;
  assign \new_[12944]_  = \new_[12943]_  & \new_[12938]_ ;
  assign \new_[12947]_  = A169 & ~A170;
  assign \new_[12951]_  = A199 & ~A166;
  assign \new_[12952]_  = ~A167 & \new_[12951]_ ;
  assign \new_[12953]_  = \new_[12952]_  & \new_[12947]_ ;
  assign \new_[12956]_  = ~A232 & A200;
  assign \new_[12960]_  = A266 & ~A265;
  assign \new_[12961]_  = A233 & \new_[12960]_ ;
  assign \new_[12962]_  = \new_[12961]_  & \new_[12956]_ ;
  assign \new_[12965]_  = A169 & ~A170;
  assign \new_[12969]_  = ~A200 & ~A166;
  assign \new_[12970]_  = ~A167 & \new_[12969]_ ;
  assign \new_[12971]_  = \new_[12970]_  & \new_[12965]_ ;
  assign \new_[12974]_  = ~A232 & ~A201;
  assign \new_[12978]_  = ~A300 & ~A299;
  assign \new_[12979]_  = A233 & \new_[12978]_ ;
  assign \new_[12980]_  = \new_[12979]_  & \new_[12974]_ ;
  assign \new_[12983]_  = A169 & ~A170;
  assign \new_[12987]_  = ~A200 & ~A166;
  assign \new_[12988]_  = ~A167 & \new_[12987]_ ;
  assign \new_[12989]_  = \new_[12988]_  & \new_[12983]_ ;
  assign \new_[12992]_  = ~A232 & ~A201;
  assign \new_[12996]_  = A299 & A298;
  assign \new_[12997]_  = A233 & \new_[12996]_ ;
  assign \new_[12998]_  = \new_[12997]_  & \new_[12992]_ ;
  assign \new_[13001]_  = A169 & ~A170;
  assign \new_[13005]_  = ~A200 & ~A166;
  assign \new_[13006]_  = ~A167 & \new_[13005]_ ;
  assign \new_[13007]_  = \new_[13006]_  & \new_[13001]_ ;
  assign \new_[13010]_  = ~A232 & ~A201;
  assign \new_[13014]_  = ~A299 & ~A298;
  assign \new_[13015]_  = A233 & \new_[13014]_ ;
  assign \new_[13016]_  = \new_[13015]_  & \new_[13010]_ ;
  assign \new_[13019]_  = A169 & ~A170;
  assign \new_[13023]_  = ~A200 & ~A166;
  assign \new_[13024]_  = ~A167 & \new_[13023]_ ;
  assign \new_[13025]_  = \new_[13024]_  & \new_[13019]_ ;
  assign \new_[13028]_  = ~A232 & ~A201;
  assign \new_[13032]_  = A266 & ~A265;
  assign \new_[13033]_  = A233 & \new_[13032]_ ;
  assign \new_[13034]_  = \new_[13033]_  & \new_[13028]_ ;
  assign \new_[13037]_  = A169 & ~A170;
  assign \new_[13041]_  = ~A199 & ~A166;
  assign \new_[13042]_  = ~A167 & \new_[13041]_ ;
  assign \new_[13043]_  = \new_[13042]_  & \new_[13037]_ ;
  assign \new_[13046]_  = ~A232 & ~A200;
  assign \new_[13050]_  = ~A300 & ~A299;
  assign \new_[13051]_  = A233 & \new_[13050]_ ;
  assign \new_[13052]_  = \new_[13051]_  & \new_[13046]_ ;
  assign \new_[13055]_  = A169 & ~A170;
  assign \new_[13059]_  = ~A199 & ~A166;
  assign \new_[13060]_  = ~A167 & \new_[13059]_ ;
  assign \new_[13061]_  = \new_[13060]_  & \new_[13055]_ ;
  assign \new_[13064]_  = ~A232 & ~A200;
  assign \new_[13068]_  = A299 & A298;
  assign \new_[13069]_  = A233 & \new_[13068]_ ;
  assign \new_[13070]_  = \new_[13069]_  & \new_[13064]_ ;
  assign \new_[13073]_  = A169 & ~A170;
  assign \new_[13077]_  = ~A199 & ~A166;
  assign \new_[13078]_  = ~A167 & \new_[13077]_ ;
  assign \new_[13079]_  = \new_[13078]_  & \new_[13073]_ ;
  assign \new_[13082]_  = ~A232 & ~A200;
  assign \new_[13086]_  = ~A299 & ~A298;
  assign \new_[13087]_  = A233 & \new_[13086]_ ;
  assign \new_[13088]_  = \new_[13087]_  & \new_[13082]_ ;
  assign \new_[13091]_  = A169 & ~A170;
  assign \new_[13095]_  = ~A199 & ~A166;
  assign \new_[13096]_  = ~A167 & \new_[13095]_ ;
  assign \new_[13097]_  = \new_[13096]_  & \new_[13091]_ ;
  assign \new_[13100]_  = ~A232 & ~A200;
  assign \new_[13104]_  = A266 & ~A265;
  assign \new_[13105]_  = A233 & \new_[13104]_ ;
  assign \new_[13106]_  = \new_[13105]_  & \new_[13100]_ ;
  assign \new_[13109]_  = ~A167 & ~A169;
  assign \new_[13113]_  = A200 & ~A199;
  assign \new_[13114]_  = ~A166 & \new_[13113]_ ;
  assign \new_[13115]_  = \new_[13114]_  & \new_[13109]_ ;
  assign \new_[13118]_  = A233 & ~A232;
  assign \new_[13122]_  = ~A302 & ~A301;
  assign \new_[13123]_  = ~A299 & \new_[13122]_ ;
  assign \new_[13124]_  = \new_[13123]_  & \new_[13118]_ ;
  assign \new_[13127]_  = ~A168 & ~A169;
  assign \new_[13131]_  = ~A199 & A166;
  assign \new_[13132]_  = A167 & \new_[13131]_ ;
  assign \new_[13133]_  = \new_[13132]_  & \new_[13127]_ ;
  assign \new_[13136]_  = ~A232 & A200;
  assign \new_[13140]_  = ~A300 & ~A299;
  assign \new_[13141]_  = A233 & \new_[13140]_ ;
  assign \new_[13142]_  = \new_[13141]_  & \new_[13136]_ ;
  assign \new_[13145]_  = ~A168 & ~A169;
  assign \new_[13149]_  = ~A199 & A166;
  assign \new_[13150]_  = A167 & \new_[13149]_ ;
  assign \new_[13151]_  = \new_[13150]_  & \new_[13145]_ ;
  assign \new_[13154]_  = ~A232 & A200;
  assign \new_[13158]_  = A299 & A298;
  assign \new_[13159]_  = A233 & \new_[13158]_ ;
  assign \new_[13160]_  = \new_[13159]_  & \new_[13154]_ ;
  assign \new_[13163]_  = ~A168 & ~A169;
  assign \new_[13167]_  = ~A199 & A166;
  assign \new_[13168]_  = A167 & \new_[13167]_ ;
  assign \new_[13169]_  = \new_[13168]_  & \new_[13163]_ ;
  assign \new_[13172]_  = ~A232 & A200;
  assign \new_[13176]_  = ~A299 & ~A298;
  assign \new_[13177]_  = A233 & \new_[13176]_ ;
  assign \new_[13178]_  = \new_[13177]_  & \new_[13172]_ ;
  assign \new_[13181]_  = ~A168 & ~A169;
  assign \new_[13185]_  = ~A199 & A166;
  assign \new_[13186]_  = A167 & \new_[13185]_ ;
  assign \new_[13187]_  = \new_[13186]_  & \new_[13181]_ ;
  assign \new_[13190]_  = ~A232 & A200;
  assign \new_[13194]_  = A266 & ~A265;
  assign \new_[13195]_  = A233 & \new_[13194]_ ;
  assign \new_[13196]_  = \new_[13195]_  & \new_[13190]_ ;
  assign \new_[13199]_  = ~A169 & A170;
  assign \new_[13203]_  = A199 & ~A166;
  assign \new_[13204]_  = A167 & \new_[13203]_ ;
  assign \new_[13205]_  = \new_[13204]_  & \new_[13199]_ ;
  assign \new_[13208]_  = ~A232 & A200;
  assign \new_[13212]_  = ~A300 & ~A299;
  assign \new_[13213]_  = A233 & \new_[13212]_ ;
  assign \new_[13214]_  = \new_[13213]_  & \new_[13208]_ ;
  assign \new_[13217]_  = ~A169 & A170;
  assign \new_[13221]_  = A199 & ~A166;
  assign \new_[13222]_  = A167 & \new_[13221]_ ;
  assign \new_[13223]_  = \new_[13222]_  & \new_[13217]_ ;
  assign \new_[13226]_  = ~A232 & A200;
  assign \new_[13230]_  = A299 & A298;
  assign \new_[13231]_  = A233 & \new_[13230]_ ;
  assign \new_[13232]_  = \new_[13231]_  & \new_[13226]_ ;
  assign \new_[13235]_  = ~A169 & A170;
  assign \new_[13239]_  = A199 & ~A166;
  assign \new_[13240]_  = A167 & \new_[13239]_ ;
  assign \new_[13241]_  = \new_[13240]_  & \new_[13235]_ ;
  assign \new_[13244]_  = ~A232 & A200;
  assign \new_[13248]_  = ~A299 & ~A298;
  assign \new_[13249]_  = A233 & \new_[13248]_ ;
  assign \new_[13250]_  = \new_[13249]_  & \new_[13244]_ ;
  assign \new_[13253]_  = ~A169 & A170;
  assign \new_[13257]_  = A199 & ~A166;
  assign \new_[13258]_  = A167 & \new_[13257]_ ;
  assign \new_[13259]_  = \new_[13258]_  & \new_[13253]_ ;
  assign \new_[13262]_  = ~A232 & A200;
  assign \new_[13266]_  = A266 & ~A265;
  assign \new_[13267]_  = A233 & \new_[13266]_ ;
  assign \new_[13268]_  = \new_[13267]_  & \new_[13262]_ ;
  assign \new_[13271]_  = ~A169 & A170;
  assign \new_[13275]_  = ~A200 & ~A166;
  assign \new_[13276]_  = A167 & \new_[13275]_ ;
  assign \new_[13277]_  = \new_[13276]_  & \new_[13271]_ ;
  assign \new_[13280]_  = ~A232 & ~A201;
  assign \new_[13284]_  = ~A300 & ~A299;
  assign \new_[13285]_  = A233 & \new_[13284]_ ;
  assign \new_[13286]_  = \new_[13285]_  & \new_[13280]_ ;
  assign \new_[13289]_  = ~A169 & A170;
  assign \new_[13293]_  = ~A200 & ~A166;
  assign \new_[13294]_  = A167 & \new_[13293]_ ;
  assign \new_[13295]_  = \new_[13294]_  & \new_[13289]_ ;
  assign \new_[13298]_  = ~A232 & ~A201;
  assign \new_[13302]_  = A299 & A298;
  assign \new_[13303]_  = A233 & \new_[13302]_ ;
  assign \new_[13304]_  = \new_[13303]_  & \new_[13298]_ ;
  assign \new_[13307]_  = ~A169 & A170;
  assign \new_[13311]_  = ~A200 & ~A166;
  assign \new_[13312]_  = A167 & \new_[13311]_ ;
  assign \new_[13313]_  = \new_[13312]_  & \new_[13307]_ ;
  assign \new_[13316]_  = ~A232 & ~A201;
  assign \new_[13320]_  = ~A299 & ~A298;
  assign \new_[13321]_  = A233 & \new_[13320]_ ;
  assign \new_[13322]_  = \new_[13321]_  & \new_[13316]_ ;
  assign \new_[13325]_  = ~A169 & A170;
  assign \new_[13329]_  = ~A200 & ~A166;
  assign \new_[13330]_  = A167 & \new_[13329]_ ;
  assign \new_[13331]_  = \new_[13330]_  & \new_[13325]_ ;
  assign \new_[13334]_  = ~A232 & ~A201;
  assign \new_[13338]_  = A266 & ~A265;
  assign \new_[13339]_  = A233 & \new_[13338]_ ;
  assign \new_[13340]_  = \new_[13339]_  & \new_[13334]_ ;
  assign \new_[13343]_  = ~A169 & A170;
  assign \new_[13347]_  = ~A199 & ~A166;
  assign \new_[13348]_  = A167 & \new_[13347]_ ;
  assign \new_[13349]_  = \new_[13348]_  & \new_[13343]_ ;
  assign \new_[13352]_  = ~A232 & ~A200;
  assign \new_[13356]_  = ~A300 & ~A299;
  assign \new_[13357]_  = A233 & \new_[13356]_ ;
  assign \new_[13358]_  = \new_[13357]_  & \new_[13352]_ ;
  assign \new_[13361]_  = ~A169 & A170;
  assign \new_[13365]_  = ~A199 & ~A166;
  assign \new_[13366]_  = A167 & \new_[13365]_ ;
  assign \new_[13367]_  = \new_[13366]_  & \new_[13361]_ ;
  assign \new_[13370]_  = ~A232 & ~A200;
  assign \new_[13374]_  = A299 & A298;
  assign \new_[13375]_  = A233 & \new_[13374]_ ;
  assign \new_[13376]_  = \new_[13375]_  & \new_[13370]_ ;
  assign \new_[13379]_  = ~A169 & A170;
  assign \new_[13383]_  = ~A199 & ~A166;
  assign \new_[13384]_  = A167 & \new_[13383]_ ;
  assign \new_[13385]_  = \new_[13384]_  & \new_[13379]_ ;
  assign \new_[13388]_  = ~A232 & ~A200;
  assign \new_[13392]_  = ~A299 & ~A298;
  assign \new_[13393]_  = A233 & \new_[13392]_ ;
  assign \new_[13394]_  = \new_[13393]_  & \new_[13388]_ ;
  assign \new_[13397]_  = ~A169 & A170;
  assign \new_[13401]_  = ~A199 & ~A166;
  assign \new_[13402]_  = A167 & \new_[13401]_ ;
  assign \new_[13403]_  = \new_[13402]_  & \new_[13397]_ ;
  assign \new_[13406]_  = ~A232 & ~A200;
  assign \new_[13410]_  = A266 & ~A265;
  assign \new_[13411]_  = A233 & \new_[13410]_ ;
  assign \new_[13412]_  = \new_[13411]_  & \new_[13406]_ ;
  assign \new_[13415]_  = ~A169 & A170;
  assign \new_[13419]_  = A199 & A166;
  assign \new_[13420]_  = ~A167 & \new_[13419]_ ;
  assign \new_[13421]_  = \new_[13420]_  & \new_[13415]_ ;
  assign \new_[13424]_  = ~A232 & A200;
  assign \new_[13428]_  = ~A300 & ~A299;
  assign \new_[13429]_  = A233 & \new_[13428]_ ;
  assign \new_[13430]_  = \new_[13429]_  & \new_[13424]_ ;
  assign \new_[13433]_  = ~A169 & A170;
  assign \new_[13437]_  = A199 & A166;
  assign \new_[13438]_  = ~A167 & \new_[13437]_ ;
  assign \new_[13439]_  = \new_[13438]_  & \new_[13433]_ ;
  assign \new_[13442]_  = ~A232 & A200;
  assign \new_[13446]_  = A299 & A298;
  assign \new_[13447]_  = A233 & \new_[13446]_ ;
  assign \new_[13448]_  = \new_[13447]_  & \new_[13442]_ ;
  assign \new_[13451]_  = ~A169 & A170;
  assign \new_[13455]_  = A199 & A166;
  assign \new_[13456]_  = ~A167 & \new_[13455]_ ;
  assign \new_[13457]_  = \new_[13456]_  & \new_[13451]_ ;
  assign \new_[13460]_  = ~A232 & A200;
  assign \new_[13464]_  = ~A299 & ~A298;
  assign \new_[13465]_  = A233 & \new_[13464]_ ;
  assign \new_[13466]_  = \new_[13465]_  & \new_[13460]_ ;
  assign \new_[13469]_  = ~A169 & A170;
  assign \new_[13473]_  = A199 & A166;
  assign \new_[13474]_  = ~A167 & \new_[13473]_ ;
  assign \new_[13475]_  = \new_[13474]_  & \new_[13469]_ ;
  assign \new_[13478]_  = ~A232 & A200;
  assign \new_[13482]_  = A266 & ~A265;
  assign \new_[13483]_  = A233 & \new_[13482]_ ;
  assign \new_[13484]_  = \new_[13483]_  & \new_[13478]_ ;
  assign \new_[13487]_  = ~A169 & A170;
  assign \new_[13491]_  = ~A200 & A166;
  assign \new_[13492]_  = ~A167 & \new_[13491]_ ;
  assign \new_[13493]_  = \new_[13492]_  & \new_[13487]_ ;
  assign \new_[13496]_  = ~A232 & ~A201;
  assign \new_[13500]_  = ~A300 & ~A299;
  assign \new_[13501]_  = A233 & \new_[13500]_ ;
  assign \new_[13502]_  = \new_[13501]_  & \new_[13496]_ ;
  assign \new_[13505]_  = ~A169 & A170;
  assign \new_[13509]_  = ~A200 & A166;
  assign \new_[13510]_  = ~A167 & \new_[13509]_ ;
  assign \new_[13511]_  = \new_[13510]_  & \new_[13505]_ ;
  assign \new_[13514]_  = ~A232 & ~A201;
  assign \new_[13518]_  = A299 & A298;
  assign \new_[13519]_  = A233 & \new_[13518]_ ;
  assign \new_[13520]_  = \new_[13519]_  & \new_[13514]_ ;
  assign \new_[13523]_  = ~A169 & A170;
  assign \new_[13527]_  = ~A200 & A166;
  assign \new_[13528]_  = ~A167 & \new_[13527]_ ;
  assign \new_[13529]_  = \new_[13528]_  & \new_[13523]_ ;
  assign \new_[13532]_  = ~A232 & ~A201;
  assign \new_[13536]_  = ~A299 & ~A298;
  assign \new_[13537]_  = A233 & \new_[13536]_ ;
  assign \new_[13538]_  = \new_[13537]_  & \new_[13532]_ ;
  assign \new_[13541]_  = ~A169 & A170;
  assign \new_[13545]_  = ~A200 & A166;
  assign \new_[13546]_  = ~A167 & \new_[13545]_ ;
  assign \new_[13547]_  = \new_[13546]_  & \new_[13541]_ ;
  assign \new_[13550]_  = ~A232 & ~A201;
  assign \new_[13554]_  = A266 & ~A265;
  assign \new_[13555]_  = A233 & \new_[13554]_ ;
  assign \new_[13556]_  = \new_[13555]_  & \new_[13550]_ ;
  assign \new_[13559]_  = ~A169 & A170;
  assign \new_[13563]_  = ~A199 & A166;
  assign \new_[13564]_  = ~A167 & \new_[13563]_ ;
  assign \new_[13565]_  = \new_[13564]_  & \new_[13559]_ ;
  assign \new_[13568]_  = ~A232 & ~A200;
  assign \new_[13572]_  = ~A300 & ~A299;
  assign \new_[13573]_  = A233 & \new_[13572]_ ;
  assign \new_[13574]_  = \new_[13573]_  & \new_[13568]_ ;
  assign \new_[13577]_  = ~A169 & A170;
  assign \new_[13581]_  = ~A199 & A166;
  assign \new_[13582]_  = ~A167 & \new_[13581]_ ;
  assign \new_[13583]_  = \new_[13582]_  & \new_[13577]_ ;
  assign \new_[13586]_  = ~A232 & ~A200;
  assign \new_[13590]_  = A299 & A298;
  assign \new_[13591]_  = A233 & \new_[13590]_ ;
  assign \new_[13592]_  = \new_[13591]_  & \new_[13586]_ ;
  assign \new_[13595]_  = ~A169 & A170;
  assign \new_[13599]_  = ~A199 & A166;
  assign \new_[13600]_  = ~A167 & \new_[13599]_ ;
  assign \new_[13601]_  = \new_[13600]_  & \new_[13595]_ ;
  assign \new_[13604]_  = ~A232 & ~A200;
  assign \new_[13608]_  = ~A299 & ~A298;
  assign \new_[13609]_  = A233 & \new_[13608]_ ;
  assign \new_[13610]_  = \new_[13609]_  & \new_[13604]_ ;
  assign \new_[13613]_  = ~A169 & A170;
  assign \new_[13617]_  = ~A199 & A166;
  assign \new_[13618]_  = ~A167 & \new_[13617]_ ;
  assign \new_[13619]_  = \new_[13618]_  & \new_[13613]_ ;
  assign \new_[13622]_  = ~A232 & ~A200;
  assign \new_[13626]_  = A266 & ~A265;
  assign \new_[13627]_  = A233 & \new_[13626]_ ;
  assign \new_[13628]_  = \new_[13627]_  & \new_[13622]_ ;
  assign \new_[13631]_  = A166 & A168;
  assign \new_[13635]_  = A232 & A200;
  assign \new_[13636]_  = A199 & \new_[13635]_ ;
  assign \new_[13637]_  = \new_[13636]_  & \new_[13631]_ ;
  assign \new_[13641]_  = ~A268 & A265;
  assign \new_[13642]_  = A233 & \new_[13641]_ ;
  assign \new_[13646]_  = A299 & ~A298;
  assign \new_[13647]_  = ~A269 & \new_[13646]_ ;
  assign \new_[13648]_  = \new_[13647]_  & \new_[13642]_ ;
  assign \new_[13651]_  = A166 & A168;
  assign \new_[13655]_  = ~A233 & A200;
  assign \new_[13656]_  = A199 & \new_[13655]_ ;
  assign \new_[13657]_  = \new_[13656]_  & \new_[13651]_ ;
  assign \new_[13661]_  = A265 & ~A236;
  assign \new_[13662]_  = ~A235 & \new_[13661]_ ;
  assign \new_[13666]_  = A299 & ~A298;
  assign \new_[13667]_  = A266 & \new_[13666]_ ;
  assign \new_[13668]_  = \new_[13667]_  & \new_[13662]_ ;
  assign \new_[13671]_  = A166 & A168;
  assign \new_[13675]_  = ~A233 & A200;
  assign \new_[13676]_  = A199 & \new_[13675]_ ;
  assign \new_[13677]_  = \new_[13676]_  & \new_[13671]_ ;
  assign \new_[13681]_  = ~A266 & ~A236;
  assign \new_[13682]_  = ~A235 & \new_[13681]_ ;
  assign \new_[13686]_  = A299 & ~A298;
  assign \new_[13687]_  = ~A267 & \new_[13686]_ ;
  assign \new_[13688]_  = \new_[13687]_  & \new_[13682]_ ;
  assign \new_[13691]_  = A166 & A168;
  assign \new_[13695]_  = ~A233 & A200;
  assign \new_[13696]_  = A199 & \new_[13695]_ ;
  assign \new_[13697]_  = \new_[13696]_  & \new_[13691]_ ;
  assign \new_[13701]_  = ~A265 & ~A236;
  assign \new_[13702]_  = ~A235 & \new_[13701]_ ;
  assign \new_[13706]_  = A299 & ~A298;
  assign \new_[13707]_  = ~A266 & \new_[13706]_ ;
  assign \new_[13708]_  = \new_[13707]_  & \new_[13702]_ ;
  assign \new_[13711]_  = A166 & A168;
  assign \new_[13715]_  = ~A233 & A200;
  assign \new_[13716]_  = A199 & \new_[13715]_ ;
  assign \new_[13717]_  = \new_[13716]_  & \new_[13711]_ ;
  assign \new_[13721]_  = ~A268 & ~A266;
  assign \new_[13722]_  = ~A234 & \new_[13721]_ ;
  assign \new_[13726]_  = A299 & ~A298;
  assign \new_[13727]_  = ~A269 & \new_[13726]_ ;
  assign \new_[13728]_  = \new_[13727]_  & \new_[13722]_ ;
  assign \new_[13731]_  = A166 & A168;
  assign \new_[13735]_  = A232 & A200;
  assign \new_[13736]_  = A199 & \new_[13735]_ ;
  assign \new_[13737]_  = \new_[13736]_  & \new_[13731]_ ;
  assign \new_[13741]_  = A235 & A234;
  assign \new_[13742]_  = ~A233 & \new_[13741]_ ;
  assign \new_[13746]_  = ~A302 & ~A301;
  assign \new_[13747]_  = A298 & \new_[13746]_ ;
  assign \new_[13748]_  = \new_[13747]_  & \new_[13742]_ ;
  assign \new_[13751]_  = A166 & A168;
  assign \new_[13755]_  = A232 & A200;
  assign \new_[13756]_  = A199 & \new_[13755]_ ;
  assign \new_[13757]_  = \new_[13756]_  & \new_[13751]_ ;
  assign \new_[13761]_  = A236 & A234;
  assign \new_[13762]_  = ~A233 & \new_[13761]_ ;
  assign \new_[13766]_  = ~A302 & ~A301;
  assign \new_[13767]_  = A298 & \new_[13766]_ ;
  assign \new_[13768]_  = \new_[13767]_  & \new_[13762]_ ;
  assign \new_[13771]_  = A166 & A168;
  assign \new_[13775]_  = ~A232 & A200;
  assign \new_[13776]_  = A199 & \new_[13775]_ ;
  assign \new_[13777]_  = \new_[13776]_  & \new_[13771]_ ;
  assign \new_[13781]_  = ~A268 & ~A266;
  assign \new_[13782]_  = ~A233 & \new_[13781]_ ;
  assign \new_[13786]_  = A299 & ~A298;
  assign \new_[13787]_  = ~A269 & \new_[13786]_ ;
  assign \new_[13788]_  = \new_[13787]_  & \new_[13782]_ ;
  assign \new_[13791]_  = A166 & A168;
  assign \new_[13795]_  = ~A203 & ~A202;
  assign \new_[13796]_  = ~A200 & \new_[13795]_ ;
  assign \new_[13797]_  = \new_[13796]_  & \new_[13791]_ ;
  assign \new_[13801]_  = A265 & A233;
  assign \new_[13802]_  = A232 & \new_[13801]_ ;
  assign \new_[13806]_  = A299 & ~A298;
  assign \new_[13807]_  = ~A267 & \new_[13806]_ ;
  assign \new_[13808]_  = \new_[13807]_  & \new_[13802]_ ;
  assign \new_[13811]_  = A166 & A168;
  assign \new_[13815]_  = ~A203 & ~A202;
  assign \new_[13816]_  = ~A200 & \new_[13815]_ ;
  assign \new_[13817]_  = \new_[13816]_  & \new_[13811]_ ;
  assign \new_[13821]_  = A265 & A233;
  assign \new_[13822]_  = A232 & \new_[13821]_ ;
  assign \new_[13826]_  = A299 & ~A298;
  assign \new_[13827]_  = A266 & \new_[13826]_ ;
  assign \new_[13828]_  = \new_[13827]_  & \new_[13822]_ ;
  assign \new_[13831]_  = A166 & A168;
  assign \new_[13835]_  = ~A203 & ~A202;
  assign \new_[13836]_  = ~A200 & \new_[13835]_ ;
  assign \new_[13837]_  = \new_[13836]_  & \new_[13831]_ ;
  assign \new_[13841]_  = ~A265 & A233;
  assign \new_[13842]_  = A232 & \new_[13841]_ ;
  assign \new_[13846]_  = A299 & ~A298;
  assign \new_[13847]_  = ~A266 & \new_[13846]_ ;
  assign \new_[13848]_  = \new_[13847]_  & \new_[13842]_ ;
  assign \new_[13851]_  = A166 & A168;
  assign \new_[13855]_  = ~A203 & ~A202;
  assign \new_[13856]_  = ~A200 & \new_[13855]_ ;
  assign \new_[13857]_  = \new_[13856]_  & \new_[13851]_ ;
  assign \new_[13861]_  = A265 & A233;
  assign \new_[13862]_  = ~A232 & \new_[13861]_ ;
  assign \new_[13866]_  = A268 & A267;
  assign \new_[13867]_  = ~A266 & \new_[13866]_ ;
  assign \new_[13868]_  = \new_[13867]_  & \new_[13862]_ ;
  assign \new_[13871]_  = A166 & A168;
  assign \new_[13875]_  = ~A203 & ~A202;
  assign \new_[13876]_  = ~A200 & \new_[13875]_ ;
  assign \new_[13877]_  = \new_[13876]_  & \new_[13871]_ ;
  assign \new_[13881]_  = A265 & A233;
  assign \new_[13882]_  = ~A232 & \new_[13881]_ ;
  assign \new_[13886]_  = A269 & A267;
  assign \new_[13887]_  = ~A266 & \new_[13886]_ ;
  assign \new_[13888]_  = \new_[13887]_  & \new_[13882]_ ;
  assign \new_[13891]_  = A166 & A168;
  assign \new_[13895]_  = ~A203 & ~A202;
  assign \new_[13896]_  = ~A200 & \new_[13895]_ ;
  assign \new_[13897]_  = \new_[13896]_  & \new_[13891]_ ;
  assign \new_[13901]_  = A265 & ~A234;
  assign \new_[13902]_  = ~A233 & \new_[13901]_ ;
  assign \new_[13906]_  = A299 & ~A298;
  assign \new_[13907]_  = A266 & \new_[13906]_ ;
  assign \new_[13908]_  = \new_[13907]_  & \new_[13902]_ ;
  assign \new_[13911]_  = A166 & A168;
  assign \new_[13915]_  = ~A203 & ~A202;
  assign \new_[13916]_  = ~A200 & \new_[13915]_ ;
  assign \new_[13917]_  = \new_[13916]_  & \new_[13911]_ ;
  assign \new_[13921]_  = ~A266 & ~A234;
  assign \new_[13922]_  = ~A233 & \new_[13921]_ ;
  assign \new_[13926]_  = A299 & ~A298;
  assign \new_[13927]_  = ~A267 & \new_[13926]_ ;
  assign \new_[13928]_  = \new_[13927]_  & \new_[13922]_ ;
  assign \new_[13931]_  = A166 & A168;
  assign \new_[13935]_  = ~A203 & ~A202;
  assign \new_[13936]_  = ~A200 & \new_[13935]_ ;
  assign \new_[13937]_  = \new_[13936]_  & \new_[13931]_ ;
  assign \new_[13941]_  = ~A265 & ~A234;
  assign \new_[13942]_  = ~A233 & \new_[13941]_ ;
  assign \new_[13946]_  = A299 & ~A298;
  assign \new_[13947]_  = ~A266 & \new_[13946]_ ;
  assign \new_[13948]_  = \new_[13947]_  & \new_[13942]_ ;
  assign \new_[13951]_  = A166 & A168;
  assign \new_[13955]_  = ~A203 & ~A202;
  assign \new_[13956]_  = ~A200 & \new_[13955]_ ;
  assign \new_[13957]_  = \new_[13956]_  & \new_[13951]_ ;
  assign \new_[13961]_  = A234 & ~A233;
  assign \new_[13962]_  = A232 & \new_[13961]_ ;
  assign \new_[13966]_  = ~A300 & A298;
  assign \new_[13967]_  = A235 & \new_[13966]_ ;
  assign \new_[13968]_  = \new_[13967]_  & \new_[13962]_ ;
  assign \new_[13971]_  = A166 & A168;
  assign \new_[13975]_  = ~A203 & ~A202;
  assign \new_[13976]_  = ~A200 & \new_[13975]_ ;
  assign \new_[13977]_  = \new_[13976]_  & \new_[13971]_ ;
  assign \new_[13981]_  = A234 & ~A233;
  assign \new_[13982]_  = A232 & \new_[13981]_ ;
  assign \new_[13986]_  = A299 & A298;
  assign \new_[13987]_  = A235 & \new_[13986]_ ;
  assign \new_[13988]_  = \new_[13987]_  & \new_[13982]_ ;
  assign \new_[13991]_  = A166 & A168;
  assign \new_[13995]_  = ~A203 & ~A202;
  assign \new_[13996]_  = ~A200 & \new_[13995]_ ;
  assign \new_[13997]_  = \new_[13996]_  & \new_[13991]_ ;
  assign \new_[14001]_  = A234 & ~A233;
  assign \new_[14002]_  = A232 & \new_[14001]_ ;
  assign \new_[14006]_  = ~A299 & ~A298;
  assign \new_[14007]_  = A235 & \new_[14006]_ ;
  assign \new_[14008]_  = \new_[14007]_  & \new_[14002]_ ;
  assign \new_[14011]_  = A166 & A168;
  assign \new_[14015]_  = ~A203 & ~A202;
  assign \new_[14016]_  = ~A200 & \new_[14015]_ ;
  assign \new_[14017]_  = \new_[14016]_  & \new_[14011]_ ;
  assign \new_[14021]_  = A234 & ~A233;
  assign \new_[14022]_  = A232 & \new_[14021]_ ;
  assign \new_[14026]_  = A266 & ~A265;
  assign \new_[14027]_  = A235 & \new_[14026]_ ;
  assign \new_[14028]_  = \new_[14027]_  & \new_[14022]_ ;
  assign \new_[14031]_  = A166 & A168;
  assign \new_[14035]_  = ~A203 & ~A202;
  assign \new_[14036]_  = ~A200 & \new_[14035]_ ;
  assign \new_[14037]_  = \new_[14036]_  & \new_[14031]_ ;
  assign \new_[14041]_  = A234 & ~A233;
  assign \new_[14042]_  = A232 & \new_[14041]_ ;
  assign \new_[14046]_  = ~A300 & A298;
  assign \new_[14047]_  = A236 & \new_[14046]_ ;
  assign \new_[14048]_  = \new_[14047]_  & \new_[14042]_ ;
  assign \new_[14051]_  = A166 & A168;
  assign \new_[14055]_  = ~A203 & ~A202;
  assign \new_[14056]_  = ~A200 & \new_[14055]_ ;
  assign \new_[14057]_  = \new_[14056]_  & \new_[14051]_ ;
  assign \new_[14061]_  = A234 & ~A233;
  assign \new_[14062]_  = A232 & \new_[14061]_ ;
  assign \new_[14066]_  = A299 & A298;
  assign \new_[14067]_  = A236 & \new_[14066]_ ;
  assign \new_[14068]_  = \new_[14067]_  & \new_[14062]_ ;
  assign \new_[14071]_  = A166 & A168;
  assign \new_[14075]_  = ~A203 & ~A202;
  assign \new_[14076]_  = ~A200 & \new_[14075]_ ;
  assign \new_[14077]_  = \new_[14076]_  & \new_[14071]_ ;
  assign \new_[14081]_  = A234 & ~A233;
  assign \new_[14082]_  = A232 & \new_[14081]_ ;
  assign \new_[14086]_  = ~A299 & ~A298;
  assign \new_[14087]_  = A236 & \new_[14086]_ ;
  assign \new_[14088]_  = \new_[14087]_  & \new_[14082]_ ;
  assign \new_[14091]_  = A166 & A168;
  assign \new_[14095]_  = ~A203 & ~A202;
  assign \new_[14096]_  = ~A200 & \new_[14095]_ ;
  assign \new_[14097]_  = \new_[14096]_  & \new_[14091]_ ;
  assign \new_[14101]_  = A234 & ~A233;
  assign \new_[14102]_  = A232 & \new_[14101]_ ;
  assign \new_[14106]_  = A266 & ~A265;
  assign \new_[14107]_  = A236 & \new_[14106]_ ;
  assign \new_[14108]_  = \new_[14107]_  & \new_[14102]_ ;
  assign \new_[14111]_  = A166 & A168;
  assign \new_[14115]_  = ~A203 & ~A202;
  assign \new_[14116]_  = ~A200 & \new_[14115]_ ;
  assign \new_[14117]_  = \new_[14116]_  & \new_[14111]_ ;
  assign \new_[14121]_  = A265 & ~A233;
  assign \new_[14122]_  = ~A232 & \new_[14121]_ ;
  assign \new_[14126]_  = A299 & ~A298;
  assign \new_[14127]_  = A266 & \new_[14126]_ ;
  assign \new_[14128]_  = \new_[14127]_  & \new_[14122]_ ;
  assign \new_[14131]_  = A166 & A168;
  assign \new_[14135]_  = ~A203 & ~A202;
  assign \new_[14136]_  = ~A200 & \new_[14135]_ ;
  assign \new_[14137]_  = \new_[14136]_  & \new_[14131]_ ;
  assign \new_[14141]_  = ~A266 & ~A233;
  assign \new_[14142]_  = ~A232 & \new_[14141]_ ;
  assign \new_[14146]_  = A299 & ~A298;
  assign \new_[14147]_  = ~A267 & \new_[14146]_ ;
  assign \new_[14148]_  = \new_[14147]_  & \new_[14142]_ ;
  assign \new_[14151]_  = A166 & A168;
  assign \new_[14155]_  = ~A203 & ~A202;
  assign \new_[14156]_  = ~A200 & \new_[14155]_ ;
  assign \new_[14157]_  = \new_[14156]_  & \new_[14151]_ ;
  assign \new_[14161]_  = ~A265 & ~A233;
  assign \new_[14162]_  = ~A232 & \new_[14161]_ ;
  assign \new_[14166]_  = A299 & ~A298;
  assign \new_[14167]_  = ~A266 & \new_[14166]_ ;
  assign \new_[14168]_  = \new_[14167]_  & \new_[14162]_ ;
  assign \new_[14171]_  = A166 & A168;
  assign \new_[14175]_  = A232 & ~A201;
  assign \new_[14176]_  = ~A200 & \new_[14175]_ ;
  assign \new_[14177]_  = \new_[14176]_  & \new_[14171]_ ;
  assign \new_[14181]_  = ~A268 & A265;
  assign \new_[14182]_  = A233 & \new_[14181]_ ;
  assign \new_[14186]_  = A299 & ~A298;
  assign \new_[14187]_  = ~A269 & \new_[14186]_ ;
  assign \new_[14188]_  = \new_[14187]_  & \new_[14182]_ ;
  assign \new_[14191]_  = A166 & A168;
  assign \new_[14195]_  = ~A233 & ~A201;
  assign \new_[14196]_  = ~A200 & \new_[14195]_ ;
  assign \new_[14197]_  = \new_[14196]_  & \new_[14191]_ ;
  assign \new_[14201]_  = A265 & ~A236;
  assign \new_[14202]_  = ~A235 & \new_[14201]_ ;
  assign \new_[14206]_  = A299 & ~A298;
  assign \new_[14207]_  = A266 & \new_[14206]_ ;
  assign \new_[14208]_  = \new_[14207]_  & \new_[14202]_ ;
  assign \new_[14211]_  = A166 & A168;
  assign \new_[14215]_  = ~A233 & ~A201;
  assign \new_[14216]_  = ~A200 & \new_[14215]_ ;
  assign \new_[14217]_  = \new_[14216]_  & \new_[14211]_ ;
  assign \new_[14221]_  = ~A266 & ~A236;
  assign \new_[14222]_  = ~A235 & \new_[14221]_ ;
  assign \new_[14226]_  = A299 & ~A298;
  assign \new_[14227]_  = ~A267 & \new_[14226]_ ;
  assign \new_[14228]_  = \new_[14227]_  & \new_[14222]_ ;
  assign \new_[14231]_  = A166 & A168;
  assign \new_[14235]_  = ~A233 & ~A201;
  assign \new_[14236]_  = ~A200 & \new_[14235]_ ;
  assign \new_[14237]_  = \new_[14236]_  & \new_[14231]_ ;
  assign \new_[14241]_  = ~A265 & ~A236;
  assign \new_[14242]_  = ~A235 & \new_[14241]_ ;
  assign \new_[14246]_  = A299 & ~A298;
  assign \new_[14247]_  = ~A266 & \new_[14246]_ ;
  assign \new_[14248]_  = \new_[14247]_  & \new_[14242]_ ;
  assign \new_[14251]_  = A166 & A168;
  assign \new_[14255]_  = ~A233 & ~A201;
  assign \new_[14256]_  = ~A200 & \new_[14255]_ ;
  assign \new_[14257]_  = \new_[14256]_  & \new_[14251]_ ;
  assign \new_[14261]_  = ~A268 & ~A266;
  assign \new_[14262]_  = ~A234 & \new_[14261]_ ;
  assign \new_[14266]_  = A299 & ~A298;
  assign \new_[14267]_  = ~A269 & \new_[14266]_ ;
  assign \new_[14268]_  = \new_[14267]_  & \new_[14262]_ ;
  assign \new_[14271]_  = A166 & A168;
  assign \new_[14275]_  = A232 & ~A201;
  assign \new_[14276]_  = ~A200 & \new_[14275]_ ;
  assign \new_[14277]_  = \new_[14276]_  & \new_[14271]_ ;
  assign \new_[14281]_  = A235 & A234;
  assign \new_[14282]_  = ~A233 & \new_[14281]_ ;
  assign \new_[14286]_  = ~A302 & ~A301;
  assign \new_[14287]_  = A298 & \new_[14286]_ ;
  assign \new_[14288]_  = \new_[14287]_  & \new_[14282]_ ;
  assign \new_[14291]_  = A166 & A168;
  assign \new_[14295]_  = A232 & ~A201;
  assign \new_[14296]_  = ~A200 & \new_[14295]_ ;
  assign \new_[14297]_  = \new_[14296]_  & \new_[14291]_ ;
  assign \new_[14301]_  = A236 & A234;
  assign \new_[14302]_  = ~A233 & \new_[14301]_ ;
  assign \new_[14306]_  = ~A302 & ~A301;
  assign \new_[14307]_  = A298 & \new_[14306]_ ;
  assign \new_[14308]_  = \new_[14307]_  & \new_[14302]_ ;
  assign \new_[14311]_  = A166 & A168;
  assign \new_[14315]_  = ~A232 & ~A201;
  assign \new_[14316]_  = ~A200 & \new_[14315]_ ;
  assign \new_[14317]_  = \new_[14316]_  & \new_[14311]_ ;
  assign \new_[14321]_  = ~A268 & ~A266;
  assign \new_[14322]_  = ~A233 & \new_[14321]_ ;
  assign \new_[14326]_  = A299 & ~A298;
  assign \new_[14327]_  = ~A269 & \new_[14326]_ ;
  assign \new_[14328]_  = \new_[14327]_  & \new_[14322]_ ;
  assign \new_[14331]_  = A166 & A168;
  assign \new_[14335]_  = A232 & ~A200;
  assign \new_[14336]_  = ~A199 & \new_[14335]_ ;
  assign \new_[14337]_  = \new_[14336]_  & \new_[14331]_ ;
  assign \new_[14341]_  = ~A268 & A265;
  assign \new_[14342]_  = A233 & \new_[14341]_ ;
  assign \new_[14346]_  = A299 & ~A298;
  assign \new_[14347]_  = ~A269 & \new_[14346]_ ;
  assign \new_[14348]_  = \new_[14347]_  & \new_[14342]_ ;
  assign \new_[14351]_  = A166 & A168;
  assign \new_[14355]_  = ~A233 & ~A200;
  assign \new_[14356]_  = ~A199 & \new_[14355]_ ;
  assign \new_[14357]_  = \new_[14356]_  & \new_[14351]_ ;
  assign \new_[14361]_  = A265 & ~A236;
  assign \new_[14362]_  = ~A235 & \new_[14361]_ ;
  assign \new_[14366]_  = A299 & ~A298;
  assign \new_[14367]_  = A266 & \new_[14366]_ ;
  assign \new_[14368]_  = \new_[14367]_  & \new_[14362]_ ;
  assign \new_[14371]_  = A166 & A168;
  assign \new_[14375]_  = ~A233 & ~A200;
  assign \new_[14376]_  = ~A199 & \new_[14375]_ ;
  assign \new_[14377]_  = \new_[14376]_  & \new_[14371]_ ;
  assign \new_[14381]_  = ~A266 & ~A236;
  assign \new_[14382]_  = ~A235 & \new_[14381]_ ;
  assign \new_[14386]_  = A299 & ~A298;
  assign \new_[14387]_  = ~A267 & \new_[14386]_ ;
  assign \new_[14388]_  = \new_[14387]_  & \new_[14382]_ ;
  assign \new_[14391]_  = A166 & A168;
  assign \new_[14395]_  = ~A233 & ~A200;
  assign \new_[14396]_  = ~A199 & \new_[14395]_ ;
  assign \new_[14397]_  = \new_[14396]_  & \new_[14391]_ ;
  assign \new_[14401]_  = ~A265 & ~A236;
  assign \new_[14402]_  = ~A235 & \new_[14401]_ ;
  assign \new_[14406]_  = A299 & ~A298;
  assign \new_[14407]_  = ~A266 & \new_[14406]_ ;
  assign \new_[14408]_  = \new_[14407]_  & \new_[14402]_ ;
  assign \new_[14411]_  = A166 & A168;
  assign \new_[14415]_  = ~A233 & ~A200;
  assign \new_[14416]_  = ~A199 & \new_[14415]_ ;
  assign \new_[14417]_  = \new_[14416]_  & \new_[14411]_ ;
  assign \new_[14421]_  = ~A268 & ~A266;
  assign \new_[14422]_  = ~A234 & \new_[14421]_ ;
  assign \new_[14426]_  = A299 & ~A298;
  assign \new_[14427]_  = ~A269 & \new_[14426]_ ;
  assign \new_[14428]_  = \new_[14427]_  & \new_[14422]_ ;
  assign \new_[14431]_  = A166 & A168;
  assign \new_[14435]_  = A232 & ~A200;
  assign \new_[14436]_  = ~A199 & \new_[14435]_ ;
  assign \new_[14437]_  = \new_[14436]_  & \new_[14431]_ ;
  assign \new_[14441]_  = A235 & A234;
  assign \new_[14442]_  = ~A233 & \new_[14441]_ ;
  assign \new_[14446]_  = ~A302 & ~A301;
  assign \new_[14447]_  = A298 & \new_[14446]_ ;
  assign \new_[14448]_  = \new_[14447]_  & \new_[14442]_ ;
  assign \new_[14451]_  = A166 & A168;
  assign \new_[14455]_  = A232 & ~A200;
  assign \new_[14456]_  = ~A199 & \new_[14455]_ ;
  assign \new_[14457]_  = \new_[14456]_  & \new_[14451]_ ;
  assign \new_[14461]_  = A236 & A234;
  assign \new_[14462]_  = ~A233 & \new_[14461]_ ;
  assign \new_[14466]_  = ~A302 & ~A301;
  assign \new_[14467]_  = A298 & \new_[14466]_ ;
  assign \new_[14468]_  = \new_[14467]_  & \new_[14462]_ ;
  assign \new_[14471]_  = A166 & A168;
  assign \new_[14475]_  = ~A232 & ~A200;
  assign \new_[14476]_  = ~A199 & \new_[14475]_ ;
  assign \new_[14477]_  = \new_[14476]_  & \new_[14471]_ ;
  assign \new_[14481]_  = ~A268 & ~A266;
  assign \new_[14482]_  = ~A233 & \new_[14481]_ ;
  assign \new_[14486]_  = A299 & ~A298;
  assign \new_[14487]_  = ~A269 & \new_[14486]_ ;
  assign \new_[14488]_  = \new_[14487]_  & \new_[14482]_ ;
  assign \new_[14491]_  = A167 & A168;
  assign \new_[14495]_  = A232 & A200;
  assign \new_[14496]_  = A199 & \new_[14495]_ ;
  assign \new_[14497]_  = \new_[14496]_  & \new_[14491]_ ;
  assign \new_[14501]_  = ~A268 & A265;
  assign \new_[14502]_  = A233 & \new_[14501]_ ;
  assign \new_[14506]_  = A299 & ~A298;
  assign \new_[14507]_  = ~A269 & \new_[14506]_ ;
  assign \new_[14508]_  = \new_[14507]_  & \new_[14502]_ ;
  assign \new_[14511]_  = A167 & A168;
  assign \new_[14515]_  = ~A233 & A200;
  assign \new_[14516]_  = A199 & \new_[14515]_ ;
  assign \new_[14517]_  = \new_[14516]_  & \new_[14511]_ ;
  assign \new_[14521]_  = A265 & ~A236;
  assign \new_[14522]_  = ~A235 & \new_[14521]_ ;
  assign \new_[14526]_  = A299 & ~A298;
  assign \new_[14527]_  = A266 & \new_[14526]_ ;
  assign \new_[14528]_  = \new_[14527]_  & \new_[14522]_ ;
  assign \new_[14531]_  = A167 & A168;
  assign \new_[14535]_  = ~A233 & A200;
  assign \new_[14536]_  = A199 & \new_[14535]_ ;
  assign \new_[14537]_  = \new_[14536]_  & \new_[14531]_ ;
  assign \new_[14541]_  = ~A266 & ~A236;
  assign \new_[14542]_  = ~A235 & \new_[14541]_ ;
  assign \new_[14546]_  = A299 & ~A298;
  assign \new_[14547]_  = ~A267 & \new_[14546]_ ;
  assign \new_[14548]_  = \new_[14547]_  & \new_[14542]_ ;
  assign \new_[14551]_  = A167 & A168;
  assign \new_[14555]_  = ~A233 & A200;
  assign \new_[14556]_  = A199 & \new_[14555]_ ;
  assign \new_[14557]_  = \new_[14556]_  & \new_[14551]_ ;
  assign \new_[14561]_  = ~A265 & ~A236;
  assign \new_[14562]_  = ~A235 & \new_[14561]_ ;
  assign \new_[14566]_  = A299 & ~A298;
  assign \new_[14567]_  = ~A266 & \new_[14566]_ ;
  assign \new_[14568]_  = \new_[14567]_  & \new_[14562]_ ;
  assign \new_[14571]_  = A167 & A168;
  assign \new_[14575]_  = ~A233 & A200;
  assign \new_[14576]_  = A199 & \new_[14575]_ ;
  assign \new_[14577]_  = \new_[14576]_  & \new_[14571]_ ;
  assign \new_[14581]_  = ~A268 & ~A266;
  assign \new_[14582]_  = ~A234 & \new_[14581]_ ;
  assign \new_[14586]_  = A299 & ~A298;
  assign \new_[14587]_  = ~A269 & \new_[14586]_ ;
  assign \new_[14588]_  = \new_[14587]_  & \new_[14582]_ ;
  assign \new_[14591]_  = A167 & A168;
  assign \new_[14595]_  = A232 & A200;
  assign \new_[14596]_  = A199 & \new_[14595]_ ;
  assign \new_[14597]_  = \new_[14596]_  & \new_[14591]_ ;
  assign \new_[14601]_  = A235 & A234;
  assign \new_[14602]_  = ~A233 & \new_[14601]_ ;
  assign \new_[14606]_  = ~A302 & ~A301;
  assign \new_[14607]_  = A298 & \new_[14606]_ ;
  assign \new_[14608]_  = \new_[14607]_  & \new_[14602]_ ;
  assign \new_[14611]_  = A167 & A168;
  assign \new_[14615]_  = A232 & A200;
  assign \new_[14616]_  = A199 & \new_[14615]_ ;
  assign \new_[14617]_  = \new_[14616]_  & \new_[14611]_ ;
  assign \new_[14621]_  = A236 & A234;
  assign \new_[14622]_  = ~A233 & \new_[14621]_ ;
  assign \new_[14626]_  = ~A302 & ~A301;
  assign \new_[14627]_  = A298 & \new_[14626]_ ;
  assign \new_[14628]_  = \new_[14627]_  & \new_[14622]_ ;
  assign \new_[14631]_  = A167 & A168;
  assign \new_[14635]_  = ~A232 & A200;
  assign \new_[14636]_  = A199 & \new_[14635]_ ;
  assign \new_[14637]_  = \new_[14636]_  & \new_[14631]_ ;
  assign \new_[14641]_  = ~A268 & ~A266;
  assign \new_[14642]_  = ~A233 & \new_[14641]_ ;
  assign \new_[14646]_  = A299 & ~A298;
  assign \new_[14647]_  = ~A269 & \new_[14646]_ ;
  assign \new_[14648]_  = \new_[14647]_  & \new_[14642]_ ;
  assign \new_[14651]_  = A167 & A168;
  assign \new_[14655]_  = ~A203 & ~A202;
  assign \new_[14656]_  = ~A200 & \new_[14655]_ ;
  assign \new_[14657]_  = \new_[14656]_  & \new_[14651]_ ;
  assign \new_[14661]_  = A265 & A233;
  assign \new_[14662]_  = A232 & \new_[14661]_ ;
  assign \new_[14666]_  = A299 & ~A298;
  assign \new_[14667]_  = ~A267 & \new_[14666]_ ;
  assign \new_[14668]_  = \new_[14667]_  & \new_[14662]_ ;
  assign \new_[14671]_  = A167 & A168;
  assign \new_[14675]_  = ~A203 & ~A202;
  assign \new_[14676]_  = ~A200 & \new_[14675]_ ;
  assign \new_[14677]_  = \new_[14676]_  & \new_[14671]_ ;
  assign \new_[14681]_  = A265 & A233;
  assign \new_[14682]_  = A232 & \new_[14681]_ ;
  assign \new_[14686]_  = A299 & ~A298;
  assign \new_[14687]_  = A266 & \new_[14686]_ ;
  assign \new_[14688]_  = \new_[14687]_  & \new_[14682]_ ;
  assign \new_[14691]_  = A167 & A168;
  assign \new_[14695]_  = ~A203 & ~A202;
  assign \new_[14696]_  = ~A200 & \new_[14695]_ ;
  assign \new_[14697]_  = \new_[14696]_  & \new_[14691]_ ;
  assign \new_[14701]_  = ~A265 & A233;
  assign \new_[14702]_  = A232 & \new_[14701]_ ;
  assign \new_[14706]_  = A299 & ~A298;
  assign \new_[14707]_  = ~A266 & \new_[14706]_ ;
  assign \new_[14708]_  = \new_[14707]_  & \new_[14702]_ ;
  assign \new_[14711]_  = A167 & A168;
  assign \new_[14715]_  = ~A203 & ~A202;
  assign \new_[14716]_  = ~A200 & \new_[14715]_ ;
  assign \new_[14717]_  = \new_[14716]_  & \new_[14711]_ ;
  assign \new_[14721]_  = A265 & A233;
  assign \new_[14722]_  = ~A232 & \new_[14721]_ ;
  assign \new_[14726]_  = A268 & A267;
  assign \new_[14727]_  = ~A266 & \new_[14726]_ ;
  assign \new_[14728]_  = \new_[14727]_  & \new_[14722]_ ;
  assign \new_[14731]_  = A167 & A168;
  assign \new_[14735]_  = ~A203 & ~A202;
  assign \new_[14736]_  = ~A200 & \new_[14735]_ ;
  assign \new_[14737]_  = \new_[14736]_  & \new_[14731]_ ;
  assign \new_[14741]_  = A265 & A233;
  assign \new_[14742]_  = ~A232 & \new_[14741]_ ;
  assign \new_[14746]_  = A269 & A267;
  assign \new_[14747]_  = ~A266 & \new_[14746]_ ;
  assign \new_[14748]_  = \new_[14747]_  & \new_[14742]_ ;
  assign \new_[14751]_  = A167 & A168;
  assign \new_[14755]_  = ~A203 & ~A202;
  assign \new_[14756]_  = ~A200 & \new_[14755]_ ;
  assign \new_[14757]_  = \new_[14756]_  & \new_[14751]_ ;
  assign \new_[14761]_  = A265 & ~A234;
  assign \new_[14762]_  = ~A233 & \new_[14761]_ ;
  assign \new_[14766]_  = A299 & ~A298;
  assign \new_[14767]_  = A266 & \new_[14766]_ ;
  assign \new_[14768]_  = \new_[14767]_  & \new_[14762]_ ;
  assign \new_[14771]_  = A167 & A168;
  assign \new_[14775]_  = ~A203 & ~A202;
  assign \new_[14776]_  = ~A200 & \new_[14775]_ ;
  assign \new_[14777]_  = \new_[14776]_  & \new_[14771]_ ;
  assign \new_[14781]_  = ~A266 & ~A234;
  assign \new_[14782]_  = ~A233 & \new_[14781]_ ;
  assign \new_[14786]_  = A299 & ~A298;
  assign \new_[14787]_  = ~A267 & \new_[14786]_ ;
  assign \new_[14788]_  = \new_[14787]_  & \new_[14782]_ ;
  assign \new_[14791]_  = A167 & A168;
  assign \new_[14795]_  = ~A203 & ~A202;
  assign \new_[14796]_  = ~A200 & \new_[14795]_ ;
  assign \new_[14797]_  = \new_[14796]_  & \new_[14791]_ ;
  assign \new_[14801]_  = ~A265 & ~A234;
  assign \new_[14802]_  = ~A233 & \new_[14801]_ ;
  assign \new_[14806]_  = A299 & ~A298;
  assign \new_[14807]_  = ~A266 & \new_[14806]_ ;
  assign \new_[14808]_  = \new_[14807]_  & \new_[14802]_ ;
  assign \new_[14811]_  = A167 & A168;
  assign \new_[14815]_  = ~A203 & ~A202;
  assign \new_[14816]_  = ~A200 & \new_[14815]_ ;
  assign \new_[14817]_  = \new_[14816]_  & \new_[14811]_ ;
  assign \new_[14821]_  = A234 & ~A233;
  assign \new_[14822]_  = A232 & \new_[14821]_ ;
  assign \new_[14826]_  = ~A300 & A298;
  assign \new_[14827]_  = A235 & \new_[14826]_ ;
  assign \new_[14828]_  = \new_[14827]_  & \new_[14822]_ ;
  assign \new_[14831]_  = A167 & A168;
  assign \new_[14835]_  = ~A203 & ~A202;
  assign \new_[14836]_  = ~A200 & \new_[14835]_ ;
  assign \new_[14837]_  = \new_[14836]_  & \new_[14831]_ ;
  assign \new_[14841]_  = A234 & ~A233;
  assign \new_[14842]_  = A232 & \new_[14841]_ ;
  assign \new_[14846]_  = A299 & A298;
  assign \new_[14847]_  = A235 & \new_[14846]_ ;
  assign \new_[14848]_  = \new_[14847]_  & \new_[14842]_ ;
  assign \new_[14851]_  = A167 & A168;
  assign \new_[14855]_  = ~A203 & ~A202;
  assign \new_[14856]_  = ~A200 & \new_[14855]_ ;
  assign \new_[14857]_  = \new_[14856]_  & \new_[14851]_ ;
  assign \new_[14861]_  = A234 & ~A233;
  assign \new_[14862]_  = A232 & \new_[14861]_ ;
  assign \new_[14866]_  = ~A299 & ~A298;
  assign \new_[14867]_  = A235 & \new_[14866]_ ;
  assign \new_[14868]_  = \new_[14867]_  & \new_[14862]_ ;
  assign \new_[14871]_  = A167 & A168;
  assign \new_[14875]_  = ~A203 & ~A202;
  assign \new_[14876]_  = ~A200 & \new_[14875]_ ;
  assign \new_[14877]_  = \new_[14876]_  & \new_[14871]_ ;
  assign \new_[14881]_  = A234 & ~A233;
  assign \new_[14882]_  = A232 & \new_[14881]_ ;
  assign \new_[14886]_  = A266 & ~A265;
  assign \new_[14887]_  = A235 & \new_[14886]_ ;
  assign \new_[14888]_  = \new_[14887]_  & \new_[14882]_ ;
  assign \new_[14891]_  = A167 & A168;
  assign \new_[14895]_  = ~A203 & ~A202;
  assign \new_[14896]_  = ~A200 & \new_[14895]_ ;
  assign \new_[14897]_  = \new_[14896]_  & \new_[14891]_ ;
  assign \new_[14901]_  = A234 & ~A233;
  assign \new_[14902]_  = A232 & \new_[14901]_ ;
  assign \new_[14906]_  = ~A300 & A298;
  assign \new_[14907]_  = A236 & \new_[14906]_ ;
  assign \new_[14908]_  = \new_[14907]_  & \new_[14902]_ ;
  assign \new_[14911]_  = A167 & A168;
  assign \new_[14915]_  = ~A203 & ~A202;
  assign \new_[14916]_  = ~A200 & \new_[14915]_ ;
  assign \new_[14917]_  = \new_[14916]_  & \new_[14911]_ ;
  assign \new_[14921]_  = A234 & ~A233;
  assign \new_[14922]_  = A232 & \new_[14921]_ ;
  assign \new_[14926]_  = A299 & A298;
  assign \new_[14927]_  = A236 & \new_[14926]_ ;
  assign \new_[14928]_  = \new_[14927]_  & \new_[14922]_ ;
  assign \new_[14931]_  = A167 & A168;
  assign \new_[14935]_  = ~A203 & ~A202;
  assign \new_[14936]_  = ~A200 & \new_[14935]_ ;
  assign \new_[14937]_  = \new_[14936]_  & \new_[14931]_ ;
  assign \new_[14941]_  = A234 & ~A233;
  assign \new_[14942]_  = A232 & \new_[14941]_ ;
  assign \new_[14946]_  = ~A299 & ~A298;
  assign \new_[14947]_  = A236 & \new_[14946]_ ;
  assign \new_[14948]_  = \new_[14947]_  & \new_[14942]_ ;
  assign \new_[14951]_  = A167 & A168;
  assign \new_[14955]_  = ~A203 & ~A202;
  assign \new_[14956]_  = ~A200 & \new_[14955]_ ;
  assign \new_[14957]_  = \new_[14956]_  & \new_[14951]_ ;
  assign \new_[14961]_  = A234 & ~A233;
  assign \new_[14962]_  = A232 & \new_[14961]_ ;
  assign \new_[14966]_  = A266 & ~A265;
  assign \new_[14967]_  = A236 & \new_[14966]_ ;
  assign \new_[14968]_  = \new_[14967]_  & \new_[14962]_ ;
  assign \new_[14971]_  = A167 & A168;
  assign \new_[14975]_  = ~A203 & ~A202;
  assign \new_[14976]_  = ~A200 & \new_[14975]_ ;
  assign \new_[14977]_  = \new_[14976]_  & \new_[14971]_ ;
  assign \new_[14981]_  = A265 & ~A233;
  assign \new_[14982]_  = ~A232 & \new_[14981]_ ;
  assign \new_[14986]_  = A299 & ~A298;
  assign \new_[14987]_  = A266 & \new_[14986]_ ;
  assign \new_[14988]_  = \new_[14987]_  & \new_[14982]_ ;
  assign \new_[14991]_  = A167 & A168;
  assign \new_[14995]_  = ~A203 & ~A202;
  assign \new_[14996]_  = ~A200 & \new_[14995]_ ;
  assign \new_[14997]_  = \new_[14996]_  & \new_[14991]_ ;
  assign \new_[15001]_  = ~A266 & ~A233;
  assign \new_[15002]_  = ~A232 & \new_[15001]_ ;
  assign \new_[15006]_  = A299 & ~A298;
  assign \new_[15007]_  = ~A267 & \new_[15006]_ ;
  assign \new_[15008]_  = \new_[15007]_  & \new_[15002]_ ;
  assign \new_[15011]_  = A167 & A168;
  assign \new_[15015]_  = ~A203 & ~A202;
  assign \new_[15016]_  = ~A200 & \new_[15015]_ ;
  assign \new_[15017]_  = \new_[15016]_  & \new_[15011]_ ;
  assign \new_[15021]_  = ~A265 & ~A233;
  assign \new_[15022]_  = ~A232 & \new_[15021]_ ;
  assign \new_[15026]_  = A299 & ~A298;
  assign \new_[15027]_  = ~A266 & \new_[15026]_ ;
  assign \new_[15028]_  = \new_[15027]_  & \new_[15022]_ ;
  assign \new_[15031]_  = A167 & A168;
  assign \new_[15035]_  = A232 & ~A201;
  assign \new_[15036]_  = ~A200 & \new_[15035]_ ;
  assign \new_[15037]_  = \new_[15036]_  & \new_[15031]_ ;
  assign \new_[15041]_  = ~A268 & A265;
  assign \new_[15042]_  = A233 & \new_[15041]_ ;
  assign \new_[15046]_  = A299 & ~A298;
  assign \new_[15047]_  = ~A269 & \new_[15046]_ ;
  assign \new_[15048]_  = \new_[15047]_  & \new_[15042]_ ;
  assign \new_[15051]_  = A167 & A168;
  assign \new_[15055]_  = ~A233 & ~A201;
  assign \new_[15056]_  = ~A200 & \new_[15055]_ ;
  assign \new_[15057]_  = \new_[15056]_  & \new_[15051]_ ;
  assign \new_[15061]_  = A265 & ~A236;
  assign \new_[15062]_  = ~A235 & \new_[15061]_ ;
  assign \new_[15066]_  = A299 & ~A298;
  assign \new_[15067]_  = A266 & \new_[15066]_ ;
  assign \new_[15068]_  = \new_[15067]_  & \new_[15062]_ ;
  assign \new_[15071]_  = A167 & A168;
  assign \new_[15075]_  = ~A233 & ~A201;
  assign \new_[15076]_  = ~A200 & \new_[15075]_ ;
  assign \new_[15077]_  = \new_[15076]_  & \new_[15071]_ ;
  assign \new_[15081]_  = ~A266 & ~A236;
  assign \new_[15082]_  = ~A235 & \new_[15081]_ ;
  assign \new_[15086]_  = A299 & ~A298;
  assign \new_[15087]_  = ~A267 & \new_[15086]_ ;
  assign \new_[15088]_  = \new_[15087]_  & \new_[15082]_ ;
  assign \new_[15091]_  = A167 & A168;
  assign \new_[15095]_  = ~A233 & ~A201;
  assign \new_[15096]_  = ~A200 & \new_[15095]_ ;
  assign \new_[15097]_  = \new_[15096]_  & \new_[15091]_ ;
  assign \new_[15101]_  = ~A265 & ~A236;
  assign \new_[15102]_  = ~A235 & \new_[15101]_ ;
  assign \new_[15106]_  = A299 & ~A298;
  assign \new_[15107]_  = ~A266 & \new_[15106]_ ;
  assign \new_[15108]_  = \new_[15107]_  & \new_[15102]_ ;
  assign \new_[15111]_  = A167 & A168;
  assign \new_[15115]_  = ~A233 & ~A201;
  assign \new_[15116]_  = ~A200 & \new_[15115]_ ;
  assign \new_[15117]_  = \new_[15116]_  & \new_[15111]_ ;
  assign \new_[15121]_  = ~A268 & ~A266;
  assign \new_[15122]_  = ~A234 & \new_[15121]_ ;
  assign \new_[15126]_  = A299 & ~A298;
  assign \new_[15127]_  = ~A269 & \new_[15126]_ ;
  assign \new_[15128]_  = \new_[15127]_  & \new_[15122]_ ;
  assign \new_[15131]_  = A167 & A168;
  assign \new_[15135]_  = A232 & ~A201;
  assign \new_[15136]_  = ~A200 & \new_[15135]_ ;
  assign \new_[15137]_  = \new_[15136]_  & \new_[15131]_ ;
  assign \new_[15141]_  = A235 & A234;
  assign \new_[15142]_  = ~A233 & \new_[15141]_ ;
  assign \new_[15146]_  = ~A302 & ~A301;
  assign \new_[15147]_  = A298 & \new_[15146]_ ;
  assign \new_[15148]_  = \new_[15147]_  & \new_[15142]_ ;
  assign \new_[15151]_  = A167 & A168;
  assign \new_[15155]_  = A232 & ~A201;
  assign \new_[15156]_  = ~A200 & \new_[15155]_ ;
  assign \new_[15157]_  = \new_[15156]_  & \new_[15151]_ ;
  assign \new_[15161]_  = A236 & A234;
  assign \new_[15162]_  = ~A233 & \new_[15161]_ ;
  assign \new_[15166]_  = ~A302 & ~A301;
  assign \new_[15167]_  = A298 & \new_[15166]_ ;
  assign \new_[15168]_  = \new_[15167]_  & \new_[15162]_ ;
  assign \new_[15171]_  = A167 & A168;
  assign \new_[15175]_  = ~A232 & ~A201;
  assign \new_[15176]_  = ~A200 & \new_[15175]_ ;
  assign \new_[15177]_  = \new_[15176]_  & \new_[15171]_ ;
  assign \new_[15181]_  = ~A268 & ~A266;
  assign \new_[15182]_  = ~A233 & \new_[15181]_ ;
  assign \new_[15186]_  = A299 & ~A298;
  assign \new_[15187]_  = ~A269 & \new_[15186]_ ;
  assign \new_[15188]_  = \new_[15187]_  & \new_[15182]_ ;
  assign \new_[15191]_  = A167 & A168;
  assign \new_[15195]_  = A232 & ~A200;
  assign \new_[15196]_  = ~A199 & \new_[15195]_ ;
  assign \new_[15197]_  = \new_[15196]_  & \new_[15191]_ ;
  assign \new_[15201]_  = ~A268 & A265;
  assign \new_[15202]_  = A233 & \new_[15201]_ ;
  assign \new_[15206]_  = A299 & ~A298;
  assign \new_[15207]_  = ~A269 & \new_[15206]_ ;
  assign \new_[15208]_  = \new_[15207]_  & \new_[15202]_ ;
  assign \new_[15211]_  = A167 & A168;
  assign \new_[15215]_  = ~A233 & ~A200;
  assign \new_[15216]_  = ~A199 & \new_[15215]_ ;
  assign \new_[15217]_  = \new_[15216]_  & \new_[15211]_ ;
  assign \new_[15221]_  = A265 & ~A236;
  assign \new_[15222]_  = ~A235 & \new_[15221]_ ;
  assign \new_[15226]_  = A299 & ~A298;
  assign \new_[15227]_  = A266 & \new_[15226]_ ;
  assign \new_[15228]_  = \new_[15227]_  & \new_[15222]_ ;
  assign \new_[15231]_  = A167 & A168;
  assign \new_[15235]_  = ~A233 & ~A200;
  assign \new_[15236]_  = ~A199 & \new_[15235]_ ;
  assign \new_[15237]_  = \new_[15236]_  & \new_[15231]_ ;
  assign \new_[15241]_  = ~A266 & ~A236;
  assign \new_[15242]_  = ~A235 & \new_[15241]_ ;
  assign \new_[15246]_  = A299 & ~A298;
  assign \new_[15247]_  = ~A267 & \new_[15246]_ ;
  assign \new_[15248]_  = \new_[15247]_  & \new_[15242]_ ;
  assign \new_[15251]_  = A167 & A168;
  assign \new_[15255]_  = ~A233 & ~A200;
  assign \new_[15256]_  = ~A199 & \new_[15255]_ ;
  assign \new_[15257]_  = \new_[15256]_  & \new_[15251]_ ;
  assign \new_[15261]_  = ~A265 & ~A236;
  assign \new_[15262]_  = ~A235 & \new_[15261]_ ;
  assign \new_[15266]_  = A299 & ~A298;
  assign \new_[15267]_  = ~A266 & \new_[15266]_ ;
  assign \new_[15268]_  = \new_[15267]_  & \new_[15262]_ ;
  assign \new_[15271]_  = A167 & A168;
  assign \new_[15275]_  = ~A233 & ~A200;
  assign \new_[15276]_  = ~A199 & \new_[15275]_ ;
  assign \new_[15277]_  = \new_[15276]_  & \new_[15271]_ ;
  assign \new_[15281]_  = ~A268 & ~A266;
  assign \new_[15282]_  = ~A234 & \new_[15281]_ ;
  assign \new_[15286]_  = A299 & ~A298;
  assign \new_[15287]_  = ~A269 & \new_[15286]_ ;
  assign \new_[15288]_  = \new_[15287]_  & \new_[15282]_ ;
  assign \new_[15291]_  = A167 & A168;
  assign \new_[15295]_  = A232 & ~A200;
  assign \new_[15296]_  = ~A199 & \new_[15295]_ ;
  assign \new_[15297]_  = \new_[15296]_  & \new_[15291]_ ;
  assign \new_[15301]_  = A235 & A234;
  assign \new_[15302]_  = ~A233 & \new_[15301]_ ;
  assign \new_[15306]_  = ~A302 & ~A301;
  assign \new_[15307]_  = A298 & \new_[15306]_ ;
  assign \new_[15308]_  = \new_[15307]_  & \new_[15302]_ ;
  assign \new_[15311]_  = A167 & A168;
  assign \new_[15315]_  = A232 & ~A200;
  assign \new_[15316]_  = ~A199 & \new_[15315]_ ;
  assign \new_[15317]_  = \new_[15316]_  & \new_[15311]_ ;
  assign \new_[15321]_  = A236 & A234;
  assign \new_[15322]_  = ~A233 & \new_[15321]_ ;
  assign \new_[15326]_  = ~A302 & ~A301;
  assign \new_[15327]_  = A298 & \new_[15326]_ ;
  assign \new_[15328]_  = \new_[15327]_  & \new_[15322]_ ;
  assign \new_[15331]_  = A167 & A168;
  assign \new_[15335]_  = ~A232 & ~A200;
  assign \new_[15336]_  = ~A199 & \new_[15335]_ ;
  assign \new_[15337]_  = \new_[15336]_  & \new_[15331]_ ;
  assign \new_[15341]_  = ~A268 & ~A266;
  assign \new_[15342]_  = ~A233 & \new_[15341]_ ;
  assign \new_[15346]_  = A299 & ~A298;
  assign \new_[15347]_  = ~A269 & \new_[15346]_ ;
  assign \new_[15348]_  = \new_[15347]_  & \new_[15342]_ ;
  assign \new_[15351]_  = ~A167 & A170;
  assign \new_[15355]_  = A200 & ~A199;
  assign \new_[15356]_  = ~A166 & \new_[15355]_ ;
  assign \new_[15357]_  = \new_[15356]_  & \new_[15351]_ ;
  assign \new_[15361]_  = A265 & A233;
  assign \new_[15362]_  = A232 & \new_[15361]_ ;
  assign \new_[15366]_  = A299 & ~A298;
  assign \new_[15367]_  = ~A267 & \new_[15366]_ ;
  assign \new_[15368]_  = \new_[15367]_  & \new_[15362]_ ;
  assign \new_[15371]_  = ~A167 & A170;
  assign \new_[15375]_  = A200 & ~A199;
  assign \new_[15376]_  = ~A166 & \new_[15375]_ ;
  assign \new_[15377]_  = \new_[15376]_  & \new_[15371]_ ;
  assign \new_[15381]_  = A265 & A233;
  assign \new_[15382]_  = A232 & \new_[15381]_ ;
  assign \new_[15386]_  = A299 & ~A298;
  assign \new_[15387]_  = A266 & \new_[15386]_ ;
  assign \new_[15388]_  = \new_[15387]_  & \new_[15382]_ ;
  assign \new_[15391]_  = ~A167 & A170;
  assign \new_[15395]_  = A200 & ~A199;
  assign \new_[15396]_  = ~A166 & \new_[15395]_ ;
  assign \new_[15397]_  = \new_[15396]_  & \new_[15391]_ ;
  assign \new_[15401]_  = ~A265 & A233;
  assign \new_[15402]_  = A232 & \new_[15401]_ ;
  assign \new_[15406]_  = A299 & ~A298;
  assign \new_[15407]_  = ~A266 & \new_[15406]_ ;
  assign \new_[15408]_  = \new_[15407]_  & \new_[15402]_ ;
  assign \new_[15411]_  = ~A167 & A170;
  assign \new_[15415]_  = A200 & ~A199;
  assign \new_[15416]_  = ~A166 & \new_[15415]_ ;
  assign \new_[15417]_  = \new_[15416]_  & \new_[15411]_ ;
  assign \new_[15421]_  = A265 & A233;
  assign \new_[15422]_  = ~A232 & \new_[15421]_ ;
  assign \new_[15426]_  = A268 & A267;
  assign \new_[15427]_  = ~A266 & \new_[15426]_ ;
  assign \new_[15428]_  = \new_[15427]_  & \new_[15422]_ ;
  assign \new_[15431]_  = ~A167 & A170;
  assign \new_[15435]_  = A200 & ~A199;
  assign \new_[15436]_  = ~A166 & \new_[15435]_ ;
  assign \new_[15437]_  = \new_[15436]_  & \new_[15431]_ ;
  assign \new_[15441]_  = A265 & A233;
  assign \new_[15442]_  = ~A232 & \new_[15441]_ ;
  assign \new_[15446]_  = A269 & A267;
  assign \new_[15447]_  = ~A266 & \new_[15446]_ ;
  assign \new_[15448]_  = \new_[15447]_  & \new_[15442]_ ;
  assign \new_[15451]_  = ~A167 & A170;
  assign \new_[15455]_  = A200 & ~A199;
  assign \new_[15456]_  = ~A166 & \new_[15455]_ ;
  assign \new_[15457]_  = \new_[15456]_  & \new_[15451]_ ;
  assign \new_[15461]_  = A265 & ~A234;
  assign \new_[15462]_  = ~A233 & \new_[15461]_ ;
  assign \new_[15466]_  = A299 & ~A298;
  assign \new_[15467]_  = A266 & \new_[15466]_ ;
  assign \new_[15468]_  = \new_[15467]_  & \new_[15462]_ ;
  assign \new_[15471]_  = ~A167 & A170;
  assign \new_[15475]_  = A200 & ~A199;
  assign \new_[15476]_  = ~A166 & \new_[15475]_ ;
  assign \new_[15477]_  = \new_[15476]_  & \new_[15471]_ ;
  assign \new_[15481]_  = ~A266 & ~A234;
  assign \new_[15482]_  = ~A233 & \new_[15481]_ ;
  assign \new_[15486]_  = A299 & ~A298;
  assign \new_[15487]_  = ~A267 & \new_[15486]_ ;
  assign \new_[15488]_  = \new_[15487]_  & \new_[15482]_ ;
  assign \new_[15491]_  = ~A167 & A170;
  assign \new_[15495]_  = A200 & ~A199;
  assign \new_[15496]_  = ~A166 & \new_[15495]_ ;
  assign \new_[15497]_  = \new_[15496]_  & \new_[15491]_ ;
  assign \new_[15501]_  = ~A265 & ~A234;
  assign \new_[15502]_  = ~A233 & \new_[15501]_ ;
  assign \new_[15506]_  = A299 & ~A298;
  assign \new_[15507]_  = ~A266 & \new_[15506]_ ;
  assign \new_[15508]_  = \new_[15507]_  & \new_[15502]_ ;
  assign \new_[15511]_  = ~A167 & A170;
  assign \new_[15515]_  = A200 & ~A199;
  assign \new_[15516]_  = ~A166 & \new_[15515]_ ;
  assign \new_[15517]_  = \new_[15516]_  & \new_[15511]_ ;
  assign \new_[15521]_  = A234 & ~A233;
  assign \new_[15522]_  = A232 & \new_[15521]_ ;
  assign \new_[15526]_  = ~A300 & A298;
  assign \new_[15527]_  = A235 & \new_[15526]_ ;
  assign \new_[15528]_  = \new_[15527]_  & \new_[15522]_ ;
  assign \new_[15531]_  = ~A167 & A170;
  assign \new_[15535]_  = A200 & ~A199;
  assign \new_[15536]_  = ~A166 & \new_[15535]_ ;
  assign \new_[15537]_  = \new_[15536]_  & \new_[15531]_ ;
  assign \new_[15541]_  = A234 & ~A233;
  assign \new_[15542]_  = A232 & \new_[15541]_ ;
  assign \new_[15546]_  = A299 & A298;
  assign \new_[15547]_  = A235 & \new_[15546]_ ;
  assign \new_[15548]_  = \new_[15547]_  & \new_[15542]_ ;
  assign \new_[15551]_  = ~A167 & A170;
  assign \new_[15555]_  = A200 & ~A199;
  assign \new_[15556]_  = ~A166 & \new_[15555]_ ;
  assign \new_[15557]_  = \new_[15556]_  & \new_[15551]_ ;
  assign \new_[15561]_  = A234 & ~A233;
  assign \new_[15562]_  = A232 & \new_[15561]_ ;
  assign \new_[15566]_  = ~A299 & ~A298;
  assign \new_[15567]_  = A235 & \new_[15566]_ ;
  assign \new_[15568]_  = \new_[15567]_  & \new_[15562]_ ;
  assign \new_[15571]_  = ~A167 & A170;
  assign \new_[15575]_  = A200 & ~A199;
  assign \new_[15576]_  = ~A166 & \new_[15575]_ ;
  assign \new_[15577]_  = \new_[15576]_  & \new_[15571]_ ;
  assign \new_[15581]_  = A234 & ~A233;
  assign \new_[15582]_  = A232 & \new_[15581]_ ;
  assign \new_[15586]_  = A266 & ~A265;
  assign \new_[15587]_  = A235 & \new_[15586]_ ;
  assign \new_[15588]_  = \new_[15587]_  & \new_[15582]_ ;
  assign \new_[15591]_  = ~A167 & A170;
  assign \new_[15595]_  = A200 & ~A199;
  assign \new_[15596]_  = ~A166 & \new_[15595]_ ;
  assign \new_[15597]_  = \new_[15596]_  & \new_[15591]_ ;
  assign \new_[15601]_  = A234 & ~A233;
  assign \new_[15602]_  = A232 & \new_[15601]_ ;
  assign \new_[15606]_  = ~A300 & A298;
  assign \new_[15607]_  = A236 & \new_[15606]_ ;
  assign \new_[15608]_  = \new_[15607]_  & \new_[15602]_ ;
  assign \new_[15611]_  = ~A167 & A170;
  assign \new_[15615]_  = A200 & ~A199;
  assign \new_[15616]_  = ~A166 & \new_[15615]_ ;
  assign \new_[15617]_  = \new_[15616]_  & \new_[15611]_ ;
  assign \new_[15621]_  = A234 & ~A233;
  assign \new_[15622]_  = A232 & \new_[15621]_ ;
  assign \new_[15626]_  = A299 & A298;
  assign \new_[15627]_  = A236 & \new_[15626]_ ;
  assign \new_[15628]_  = \new_[15627]_  & \new_[15622]_ ;
  assign \new_[15631]_  = ~A167 & A170;
  assign \new_[15635]_  = A200 & ~A199;
  assign \new_[15636]_  = ~A166 & \new_[15635]_ ;
  assign \new_[15637]_  = \new_[15636]_  & \new_[15631]_ ;
  assign \new_[15641]_  = A234 & ~A233;
  assign \new_[15642]_  = A232 & \new_[15641]_ ;
  assign \new_[15646]_  = ~A299 & ~A298;
  assign \new_[15647]_  = A236 & \new_[15646]_ ;
  assign \new_[15648]_  = \new_[15647]_  & \new_[15642]_ ;
  assign \new_[15651]_  = ~A167 & A170;
  assign \new_[15655]_  = A200 & ~A199;
  assign \new_[15656]_  = ~A166 & \new_[15655]_ ;
  assign \new_[15657]_  = \new_[15656]_  & \new_[15651]_ ;
  assign \new_[15661]_  = A234 & ~A233;
  assign \new_[15662]_  = A232 & \new_[15661]_ ;
  assign \new_[15666]_  = A266 & ~A265;
  assign \new_[15667]_  = A236 & \new_[15666]_ ;
  assign \new_[15668]_  = \new_[15667]_  & \new_[15662]_ ;
  assign \new_[15671]_  = ~A167 & A170;
  assign \new_[15675]_  = A200 & ~A199;
  assign \new_[15676]_  = ~A166 & \new_[15675]_ ;
  assign \new_[15677]_  = \new_[15676]_  & \new_[15671]_ ;
  assign \new_[15681]_  = A265 & ~A233;
  assign \new_[15682]_  = ~A232 & \new_[15681]_ ;
  assign \new_[15686]_  = A299 & ~A298;
  assign \new_[15687]_  = A266 & \new_[15686]_ ;
  assign \new_[15688]_  = \new_[15687]_  & \new_[15682]_ ;
  assign \new_[15691]_  = ~A167 & A170;
  assign \new_[15695]_  = A200 & ~A199;
  assign \new_[15696]_  = ~A166 & \new_[15695]_ ;
  assign \new_[15697]_  = \new_[15696]_  & \new_[15691]_ ;
  assign \new_[15701]_  = ~A266 & ~A233;
  assign \new_[15702]_  = ~A232 & \new_[15701]_ ;
  assign \new_[15706]_  = A299 & ~A298;
  assign \new_[15707]_  = ~A267 & \new_[15706]_ ;
  assign \new_[15708]_  = \new_[15707]_  & \new_[15702]_ ;
  assign \new_[15711]_  = ~A167 & A170;
  assign \new_[15715]_  = A200 & ~A199;
  assign \new_[15716]_  = ~A166 & \new_[15715]_ ;
  assign \new_[15717]_  = \new_[15716]_  & \new_[15711]_ ;
  assign \new_[15721]_  = ~A265 & ~A233;
  assign \new_[15722]_  = ~A232 & \new_[15721]_ ;
  assign \new_[15726]_  = A299 & ~A298;
  assign \new_[15727]_  = ~A266 & \new_[15726]_ ;
  assign \new_[15728]_  = \new_[15727]_  & \new_[15722]_ ;
  assign \new_[15731]_  = ~A167 & A170;
  assign \new_[15735]_  = ~A200 & A199;
  assign \new_[15736]_  = ~A166 & \new_[15735]_ ;
  assign \new_[15737]_  = \new_[15736]_  & \new_[15731]_ ;
  assign \new_[15741]_  = ~A232 & A202;
  assign \new_[15742]_  = A201 & \new_[15741]_ ;
  assign \new_[15746]_  = ~A300 & ~A299;
  assign \new_[15747]_  = A233 & \new_[15746]_ ;
  assign \new_[15748]_  = \new_[15747]_  & \new_[15742]_ ;
  assign \new_[15751]_  = ~A167 & A170;
  assign \new_[15755]_  = ~A200 & A199;
  assign \new_[15756]_  = ~A166 & \new_[15755]_ ;
  assign \new_[15757]_  = \new_[15756]_  & \new_[15751]_ ;
  assign \new_[15761]_  = ~A232 & A202;
  assign \new_[15762]_  = A201 & \new_[15761]_ ;
  assign \new_[15766]_  = A299 & A298;
  assign \new_[15767]_  = A233 & \new_[15766]_ ;
  assign \new_[15768]_  = \new_[15767]_  & \new_[15762]_ ;
  assign \new_[15771]_  = ~A167 & A170;
  assign \new_[15775]_  = ~A200 & A199;
  assign \new_[15776]_  = ~A166 & \new_[15775]_ ;
  assign \new_[15777]_  = \new_[15776]_  & \new_[15771]_ ;
  assign \new_[15781]_  = ~A232 & A202;
  assign \new_[15782]_  = A201 & \new_[15781]_ ;
  assign \new_[15786]_  = ~A299 & ~A298;
  assign \new_[15787]_  = A233 & \new_[15786]_ ;
  assign \new_[15788]_  = \new_[15787]_  & \new_[15782]_ ;
  assign \new_[15791]_  = ~A167 & A170;
  assign \new_[15795]_  = ~A200 & A199;
  assign \new_[15796]_  = ~A166 & \new_[15795]_ ;
  assign \new_[15797]_  = \new_[15796]_  & \new_[15791]_ ;
  assign \new_[15801]_  = ~A232 & A202;
  assign \new_[15802]_  = A201 & \new_[15801]_ ;
  assign \new_[15806]_  = A266 & ~A265;
  assign \new_[15807]_  = A233 & \new_[15806]_ ;
  assign \new_[15808]_  = \new_[15807]_  & \new_[15802]_ ;
  assign \new_[15811]_  = ~A167 & A170;
  assign \new_[15815]_  = ~A200 & A199;
  assign \new_[15816]_  = ~A166 & \new_[15815]_ ;
  assign \new_[15817]_  = \new_[15816]_  & \new_[15811]_ ;
  assign \new_[15821]_  = ~A232 & A203;
  assign \new_[15822]_  = A201 & \new_[15821]_ ;
  assign \new_[15826]_  = ~A300 & ~A299;
  assign \new_[15827]_  = A233 & \new_[15826]_ ;
  assign \new_[15828]_  = \new_[15827]_  & \new_[15822]_ ;
  assign \new_[15831]_  = ~A167 & A170;
  assign \new_[15835]_  = ~A200 & A199;
  assign \new_[15836]_  = ~A166 & \new_[15835]_ ;
  assign \new_[15837]_  = \new_[15836]_  & \new_[15831]_ ;
  assign \new_[15841]_  = ~A232 & A203;
  assign \new_[15842]_  = A201 & \new_[15841]_ ;
  assign \new_[15846]_  = A299 & A298;
  assign \new_[15847]_  = A233 & \new_[15846]_ ;
  assign \new_[15848]_  = \new_[15847]_  & \new_[15842]_ ;
  assign \new_[15851]_  = ~A167 & A170;
  assign \new_[15855]_  = ~A200 & A199;
  assign \new_[15856]_  = ~A166 & \new_[15855]_ ;
  assign \new_[15857]_  = \new_[15856]_  & \new_[15851]_ ;
  assign \new_[15861]_  = ~A232 & A203;
  assign \new_[15862]_  = A201 & \new_[15861]_ ;
  assign \new_[15866]_  = ~A299 & ~A298;
  assign \new_[15867]_  = A233 & \new_[15866]_ ;
  assign \new_[15868]_  = \new_[15867]_  & \new_[15862]_ ;
  assign \new_[15871]_  = ~A167 & A170;
  assign \new_[15875]_  = ~A200 & A199;
  assign \new_[15876]_  = ~A166 & \new_[15875]_ ;
  assign \new_[15877]_  = \new_[15876]_  & \new_[15871]_ ;
  assign \new_[15881]_  = ~A232 & A203;
  assign \new_[15882]_  = A201 & \new_[15881]_ ;
  assign \new_[15886]_  = A266 & ~A265;
  assign \new_[15887]_  = A233 & \new_[15886]_ ;
  assign \new_[15888]_  = \new_[15887]_  & \new_[15882]_ ;
  assign \new_[15891]_  = ~A168 & A170;
  assign \new_[15895]_  = ~A199 & A166;
  assign \new_[15896]_  = A167 & \new_[15895]_ ;
  assign \new_[15897]_  = \new_[15896]_  & \new_[15891]_ ;
  assign \new_[15901]_  = A233 & ~A232;
  assign \new_[15902]_  = A200 & \new_[15901]_ ;
  assign \new_[15906]_  = ~A302 & ~A301;
  assign \new_[15907]_  = ~A299 & \new_[15906]_ ;
  assign \new_[15908]_  = \new_[15907]_  & \new_[15902]_ ;
  assign \new_[15911]_  = ~A168 & ~A170;
  assign \new_[15915]_  = ~A199 & ~A166;
  assign \new_[15916]_  = A167 & \new_[15915]_ ;
  assign \new_[15917]_  = \new_[15916]_  & \new_[15911]_ ;
  assign \new_[15921]_  = A233 & ~A232;
  assign \new_[15922]_  = A200 & \new_[15921]_ ;
  assign \new_[15926]_  = ~A302 & ~A301;
  assign \new_[15927]_  = ~A299 & \new_[15926]_ ;
  assign \new_[15928]_  = \new_[15927]_  & \new_[15922]_ ;
  assign \new_[15931]_  = ~A168 & ~A170;
  assign \new_[15935]_  = ~A199 & A166;
  assign \new_[15936]_  = ~A167 & \new_[15935]_ ;
  assign \new_[15937]_  = \new_[15936]_  & \new_[15931]_ ;
  assign \new_[15941]_  = A233 & ~A232;
  assign \new_[15942]_  = A200 & \new_[15941]_ ;
  assign \new_[15946]_  = ~A302 & ~A301;
  assign \new_[15947]_  = ~A299 & \new_[15946]_ ;
  assign \new_[15948]_  = \new_[15947]_  & \new_[15942]_ ;
  assign \new_[15951]_  = ~A168 & A169;
  assign \new_[15955]_  = ~A199 & ~A166;
  assign \new_[15956]_  = A167 & \new_[15955]_ ;
  assign \new_[15957]_  = \new_[15956]_  & \new_[15951]_ ;
  assign \new_[15961]_  = A233 & ~A232;
  assign \new_[15962]_  = A200 & \new_[15961]_ ;
  assign \new_[15966]_  = ~A302 & ~A301;
  assign \new_[15967]_  = ~A299 & \new_[15966]_ ;
  assign \new_[15968]_  = \new_[15967]_  & \new_[15962]_ ;
  assign \new_[15971]_  = ~A168 & A169;
  assign \new_[15975]_  = ~A199 & A166;
  assign \new_[15976]_  = ~A167 & \new_[15975]_ ;
  assign \new_[15977]_  = \new_[15976]_  & \new_[15971]_ ;
  assign \new_[15981]_  = A233 & ~A232;
  assign \new_[15982]_  = A200 & \new_[15981]_ ;
  assign \new_[15986]_  = ~A302 & ~A301;
  assign \new_[15987]_  = ~A299 & \new_[15986]_ ;
  assign \new_[15988]_  = \new_[15987]_  & \new_[15982]_ ;
  assign \new_[15991]_  = A169 & A170;
  assign \new_[15995]_  = ~A200 & A199;
  assign \new_[15996]_  = ~A168 & \new_[15995]_ ;
  assign \new_[15997]_  = \new_[15996]_  & \new_[15991]_ ;
  assign \new_[16001]_  = ~A232 & A202;
  assign \new_[16002]_  = A201 & \new_[16001]_ ;
  assign \new_[16006]_  = ~A300 & ~A299;
  assign \new_[16007]_  = A233 & \new_[16006]_ ;
  assign \new_[16008]_  = \new_[16007]_  & \new_[16002]_ ;
  assign \new_[16011]_  = A169 & A170;
  assign \new_[16015]_  = ~A200 & A199;
  assign \new_[16016]_  = ~A168 & \new_[16015]_ ;
  assign \new_[16017]_  = \new_[16016]_  & \new_[16011]_ ;
  assign \new_[16021]_  = ~A232 & A202;
  assign \new_[16022]_  = A201 & \new_[16021]_ ;
  assign \new_[16026]_  = A299 & A298;
  assign \new_[16027]_  = A233 & \new_[16026]_ ;
  assign \new_[16028]_  = \new_[16027]_  & \new_[16022]_ ;
  assign \new_[16031]_  = A169 & A170;
  assign \new_[16035]_  = ~A200 & A199;
  assign \new_[16036]_  = ~A168 & \new_[16035]_ ;
  assign \new_[16037]_  = \new_[16036]_  & \new_[16031]_ ;
  assign \new_[16041]_  = ~A232 & A202;
  assign \new_[16042]_  = A201 & \new_[16041]_ ;
  assign \new_[16046]_  = ~A299 & ~A298;
  assign \new_[16047]_  = A233 & \new_[16046]_ ;
  assign \new_[16048]_  = \new_[16047]_  & \new_[16042]_ ;
  assign \new_[16051]_  = A169 & A170;
  assign \new_[16055]_  = ~A200 & A199;
  assign \new_[16056]_  = ~A168 & \new_[16055]_ ;
  assign \new_[16057]_  = \new_[16056]_  & \new_[16051]_ ;
  assign \new_[16061]_  = ~A232 & A202;
  assign \new_[16062]_  = A201 & \new_[16061]_ ;
  assign \new_[16066]_  = A266 & ~A265;
  assign \new_[16067]_  = A233 & \new_[16066]_ ;
  assign \new_[16068]_  = \new_[16067]_  & \new_[16062]_ ;
  assign \new_[16071]_  = A169 & A170;
  assign \new_[16075]_  = ~A200 & A199;
  assign \new_[16076]_  = ~A168 & \new_[16075]_ ;
  assign \new_[16077]_  = \new_[16076]_  & \new_[16071]_ ;
  assign \new_[16081]_  = ~A232 & A203;
  assign \new_[16082]_  = A201 & \new_[16081]_ ;
  assign \new_[16086]_  = ~A300 & ~A299;
  assign \new_[16087]_  = A233 & \new_[16086]_ ;
  assign \new_[16088]_  = \new_[16087]_  & \new_[16082]_ ;
  assign \new_[16091]_  = A169 & A170;
  assign \new_[16095]_  = ~A200 & A199;
  assign \new_[16096]_  = ~A168 & \new_[16095]_ ;
  assign \new_[16097]_  = \new_[16096]_  & \new_[16091]_ ;
  assign \new_[16101]_  = ~A232 & A203;
  assign \new_[16102]_  = A201 & \new_[16101]_ ;
  assign \new_[16106]_  = A299 & A298;
  assign \new_[16107]_  = A233 & \new_[16106]_ ;
  assign \new_[16108]_  = \new_[16107]_  & \new_[16102]_ ;
  assign \new_[16111]_  = A169 & A170;
  assign \new_[16115]_  = ~A200 & A199;
  assign \new_[16116]_  = ~A168 & \new_[16115]_ ;
  assign \new_[16117]_  = \new_[16116]_  & \new_[16111]_ ;
  assign \new_[16121]_  = ~A232 & A203;
  assign \new_[16122]_  = A201 & \new_[16121]_ ;
  assign \new_[16126]_  = ~A299 & ~A298;
  assign \new_[16127]_  = A233 & \new_[16126]_ ;
  assign \new_[16128]_  = \new_[16127]_  & \new_[16122]_ ;
  assign \new_[16131]_  = A169 & A170;
  assign \new_[16135]_  = ~A200 & A199;
  assign \new_[16136]_  = ~A168 & \new_[16135]_ ;
  assign \new_[16137]_  = \new_[16136]_  & \new_[16131]_ ;
  assign \new_[16141]_  = ~A232 & A203;
  assign \new_[16142]_  = A201 & \new_[16141]_ ;
  assign \new_[16146]_  = A266 & ~A265;
  assign \new_[16147]_  = A233 & \new_[16146]_ ;
  assign \new_[16148]_  = \new_[16147]_  & \new_[16142]_ ;
  assign \new_[16151]_  = A169 & ~A170;
  assign \new_[16155]_  = A199 & A166;
  assign \new_[16156]_  = A167 & \new_[16155]_ ;
  assign \new_[16157]_  = \new_[16156]_  & \new_[16151]_ ;
  assign \new_[16161]_  = A233 & ~A232;
  assign \new_[16162]_  = A200 & \new_[16161]_ ;
  assign \new_[16166]_  = ~A302 & ~A301;
  assign \new_[16167]_  = ~A299 & \new_[16166]_ ;
  assign \new_[16168]_  = \new_[16167]_  & \new_[16162]_ ;
  assign \new_[16171]_  = A169 & ~A170;
  assign \new_[16175]_  = ~A200 & A166;
  assign \new_[16176]_  = A167 & \new_[16175]_ ;
  assign \new_[16177]_  = \new_[16176]_  & \new_[16171]_ ;
  assign \new_[16181]_  = ~A232 & ~A203;
  assign \new_[16182]_  = ~A202 & \new_[16181]_ ;
  assign \new_[16186]_  = ~A300 & ~A299;
  assign \new_[16187]_  = A233 & \new_[16186]_ ;
  assign \new_[16188]_  = \new_[16187]_  & \new_[16182]_ ;
  assign \new_[16191]_  = A169 & ~A170;
  assign \new_[16195]_  = ~A200 & A166;
  assign \new_[16196]_  = A167 & \new_[16195]_ ;
  assign \new_[16197]_  = \new_[16196]_  & \new_[16191]_ ;
  assign \new_[16201]_  = ~A232 & ~A203;
  assign \new_[16202]_  = ~A202 & \new_[16201]_ ;
  assign \new_[16206]_  = A299 & A298;
  assign \new_[16207]_  = A233 & \new_[16206]_ ;
  assign \new_[16208]_  = \new_[16207]_  & \new_[16202]_ ;
  assign \new_[16211]_  = A169 & ~A170;
  assign \new_[16215]_  = ~A200 & A166;
  assign \new_[16216]_  = A167 & \new_[16215]_ ;
  assign \new_[16217]_  = \new_[16216]_  & \new_[16211]_ ;
  assign \new_[16221]_  = ~A232 & ~A203;
  assign \new_[16222]_  = ~A202 & \new_[16221]_ ;
  assign \new_[16226]_  = ~A299 & ~A298;
  assign \new_[16227]_  = A233 & \new_[16226]_ ;
  assign \new_[16228]_  = \new_[16227]_  & \new_[16222]_ ;
  assign \new_[16231]_  = A169 & ~A170;
  assign \new_[16235]_  = ~A200 & A166;
  assign \new_[16236]_  = A167 & \new_[16235]_ ;
  assign \new_[16237]_  = \new_[16236]_  & \new_[16231]_ ;
  assign \new_[16241]_  = ~A232 & ~A203;
  assign \new_[16242]_  = ~A202 & \new_[16241]_ ;
  assign \new_[16246]_  = A266 & ~A265;
  assign \new_[16247]_  = A233 & \new_[16246]_ ;
  assign \new_[16248]_  = \new_[16247]_  & \new_[16242]_ ;
  assign \new_[16251]_  = A169 & ~A170;
  assign \new_[16255]_  = ~A200 & A166;
  assign \new_[16256]_  = A167 & \new_[16255]_ ;
  assign \new_[16257]_  = \new_[16256]_  & \new_[16251]_ ;
  assign \new_[16261]_  = A233 & ~A232;
  assign \new_[16262]_  = ~A201 & \new_[16261]_ ;
  assign \new_[16266]_  = ~A302 & ~A301;
  assign \new_[16267]_  = ~A299 & \new_[16266]_ ;
  assign \new_[16268]_  = \new_[16267]_  & \new_[16262]_ ;
  assign \new_[16271]_  = A169 & ~A170;
  assign \new_[16275]_  = ~A199 & A166;
  assign \new_[16276]_  = A167 & \new_[16275]_ ;
  assign \new_[16277]_  = \new_[16276]_  & \new_[16271]_ ;
  assign \new_[16281]_  = A233 & ~A232;
  assign \new_[16282]_  = ~A200 & \new_[16281]_ ;
  assign \new_[16286]_  = ~A302 & ~A301;
  assign \new_[16287]_  = ~A299 & \new_[16286]_ ;
  assign \new_[16288]_  = \new_[16287]_  & \new_[16282]_ ;
  assign \new_[16291]_  = A169 & ~A170;
  assign \new_[16295]_  = A199 & ~A166;
  assign \new_[16296]_  = ~A167 & \new_[16295]_ ;
  assign \new_[16297]_  = \new_[16296]_  & \new_[16291]_ ;
  assign \new_[16301]_  = A233 & ~A232;
  assign \new_[16302]_  = A200 & \new_[16301]_ ;
  assign \new_[16306]_  = ~A302 & ~A301;
  assign \new_[16307]_  = ~A299 & \new_[16306]_ ;
  assign \new_[16308]_  = \new_[16307]_  & \new_[16302]_ ;
  assign \new_[16311]_  = A169 & ~A170;
  assign \new_[16315]_  = ~A200 & ~A166;
  assign \new_[16316]_  = ~A167 & \new_[16315]_ ;
  assign \new_[16317]_  = \new_[16316]_  & \new_[16311]_ ;
  assign \new_[16321]_  = ~A232 & ~A203;
  assign \new_[16322]_  = ~A202 & \new_[16321]_ ;
  assign \new_[16326]_  = ~A300 & ~A299;
  assign \new_[16327]_  = A233 & \new_[16326]_ ;
  assign \new_[16328]_  = \new_[16327]_  & \new_[16322]_ ;
  assign \new_[16331]_  = A169 & ~A170;
  assign \new_[16335]_  = ~A200 & ~A166;
  assign \new_[16336]_  = ~A167 & \new_[16335]_ ;
  assign \new_[16337]_  = \new_[16336]_  & \new_[16331]_ ;
  assign \new_[16341]_  = ~A232 & ~A203;
  assign \new_[16342]_  = ~A202 & \new_[16341]_ ;
  assign \new_[16346]_  = A299 & A298;
  assign \new_[16347]_  = A233 & \new_[16346]_ ;
  assign \new_[16348]_  = \new_[16347]_  & \new_[16342]_ ;
  assign \new_[16351]_  = A169 & ~A170;
  assign \new_[16355]_  = ~A200 & ~A166;
  assign \new_[16356]_  = ~A167 & \new_[16355]_ ;
  assign \new_[16357]_  = \new_[16356]_  & \new_[16351]_ ;
  assign \new_[16361]_  = ~A232 & ~A203;
  assign \new_[16362]_  = ~A202 & \new_[16361]_ ;
  assign \new_[16366]_  = ~A299 & ~A298;
  assign \new_[16367]_  = A233 & \new_[16366]_ ;
  assign \new_[16368]_  = \new_[16367]_  & \new_[16362]_ ;
  assign \new_[16371]_  = A169 & ~A170;
  assign \new_[16375]_  = ~A200 & ~A166;
  assign \new_[16376]_  = ~A167 & \new_[16375]_ ;
  assign \new_[16377]_  = \new_[16376]_  & \new_[16371]_ ;
  assign \new_[16381]_  = ~A232 & ~A203;
  assign \new_[16382]_  = ~A202 & \new_[16381]_ ;
  assign \new_[16386]_  = A266 & ~A265;
  assign \new_[16387]_  = A233 & \new_[16386]_ ;
  assign \new_[16388]_  = \new_[16387]_  & \new_[16382]_ ;
  assign \new_[16391]_  = A169 & ~A170;
  assign \new_[16395]_  = ~A200 & ~A166;
  assign \new_[16396]_  = ~A167 & \new_[16395]_ ;
  assign \new_[16397]_  = \new_[16396]_  & \new_[16391]_ ;
  assign \new_[16401]_  = A233 & ~A232;
  assign \new_[16402]_  = ~A201 & \new_[16401]_ ;
  assign \new_[16406]_  = ~A302 & ~A301;
  assign \new_[16407]_  = ~A299 & \new_[16406]_ ;
  assign \new_[16408]_  = \new_[16407]_  & \new_[16402]_ ;
  assign \new_[16411]_  = A169 & ~A170;
  assign \new_[16415]_  = ~A199 & ~A166;
  assign \new_[16416]_  = ~A167 & \new_[16415]_ ;
  assign \new_[16417]_  = \new_[16416]_  & \new_[16411]_ ;
  assign \new_[16421]_  = A233 & ~A232;
  assign \new_[16422]_  = ~A200 & \new_[16421]_ ;
  assign \new_[16426]_  = ~A302 & ~A301;
  assign \new_[16427]_  = ~A299 & \new_[16426]_ ;
  assign \new_[16428]_  = \new_[16427]_  & \new_[16422]_ ;
  assign \new_[16431]_  = ~A167 & ~A169;
  assign \new_[16435]_  = A200 & ~A199;
  assign \new_[16436]_  = ~A166 & \new_[16435]_ ;
  assign \new_[16437]_  = \new_[16436]_  & \new_[16431]_ ;
  assign \new_[16441]_  = A265 & A233;
  assign \new_[16442]_  = A232 & \new_[16441]_ ;
  assign \new_[16446]_  = A299 & ~A298;
  assign \new_[16447]_  = ~A267 & \new_[16446]_ ;
  assign \new_[16448]_  = \new_[16447]_  & \new_[16442]_ ;
  assign \new_[16451]_  = ~A167 & ~A169;
  assign \new_[16455]_  = A200 & ~A199;
  assign \new_[16456]_  = ~A166 & \new_[16455]_ ;
  assign \new_[16457]_  = \new_[16456]_  & \new_[16451]_ ;
  assign \new_[16461]_  = A265 & A233;
  assign \new_[16462]_  = A232 & \new_[16461]_ ;
  assign \new_[16466]_  = A299 & ~A298;
  assign \new_[16467]_  = A266 & \new_[16466]_ ;
  assign \new_[16468]_  = \new_[16467]_  & \new_[16462]_ ;
  assign \new_[16471]_  = ~A167 & ~A169;
  assign \new_[16475]_  = A200 & ~A199;
  assign \new_[16476]_  = ~A166 & \new_[16475]_ ;
  assign \new_[16477]_  = \new_[16476]_  & \new_[16471]_ ;
  assign \new_[16481]_  = ~A265 & A233;
  assign \new_[16482]_  = A232 & \new_[16481]_ ;
  assign \new_[16486]_  = A299 & ~A298;
  assign \new_[16487]_  = ~A266 & \new_[16486]_ ;
  assign \new_[16488]_  = \new_[16487]_  & \new_[16482]_ ;
  assign \new_[16491]_  = ~A167 & ~A169;
  assign \new_[16495]_  = A200 & ~A199;
  assign \new_[16496]_  = ~A166 & \new_[16495]_ ;
  assign \new_[16497]_  = \new_[16496]_  & \new_[16491]_ ;
  assign \new_[16501]_  = A265 & A233;
  assign \new_[16502]_  = ~A232 & \new_[16501]_ ;
  assign \new_[16506]_  = A268 & A267;
  assign \new_[16507]_  = ~A266 & \new_[16506]_ ;
  assign \new_[16508]_  = \new_[16507]_  & \new_[16502]_ ;
  assign \new_[16511]_  = ~A167 & ~A169;
  assign \new_[16515]_  = A200 & ~A199;
  assign \new_[16516]_  = ~A166 & \new_[16515]_ ;
  assign \new_[16517]_  = \new_[16516]_  & \new_[16511]_ ;
  assign \new_[16521]_  = A265 & A233;
  assign \new_[16522]_  = ~A232 & \new_[16521]_ ;
  assign \new_[16526]_  = A269 & A267;
  assign \new_[16527]_  = ~A266 & \new_[16526]_ ;
  assign \new_[16528]_  = \new_[16527]_  & \new_[16522]_ ;
  assign \new_[16531]_  = ~A167 & ~A169;
  assign \new_[16535]_  = A200 & ~A199;
  assign \new_[16536]_  = ~A166 & \new_[16535]_ ;
  assign \new_[16537]_  = \new_[16536]_  & \new_[16531]_ ;
  assign \new_[16541]_  = A265 & ~A234;
  assign \new_[16542]_  = ~A233 & \new_[16541]_ ;
  assign \new_[16546]_  = A299 & ~A298;
  assign \new_[16547]_  = A266 & \new_[16546]_ ;
  assign \new_[16548]_  = \new_[16547]_  & \new_[16542]_ ;
  assign \new_[16551]_  = ~A167 & ~A169;
  assign \new_[16555]_  = A200 & ~A199;
  assign \new_[16556]_  = ~A166 & \new_[16555]_ ;
  assign \new_[16557]_  = \new_[16556]_  & \new_[16551]_ ;
  assign \new_[16561]_  = ~A266 & ~A234;
  assign \new_[16562]_  = ~A233 & \new_[16561]_ ;
  assign \new_[16566]_  = A299 & ~A298;
  assign \new_[16567]_  = ~A267 & \new_[16566]_ ;
  assign \new_[16568]_  = \new_[16567]_  & \new_[16562]_ ;
  assign \new_[16571]_  = ~A167 & ~A169;
  assign \new_[16575]_  = A200 & ~A199;
  assign \new_[16576]_  = ~A166 & \new_[16575]_ ;
  assign \new_[16577]_  = \new_[16576]_  & \new_[16571]_ ;
  assign \new_[16581]_  = ~A265 & ~A234;
  assign \new_[16582]_  = ~A233 & \new_[16581]_ ;
  assign \new_[16586]_  = A299 & ~A298;
  assign \new_[16587]_  = ~A266 & \new_[16586]_ ;
  assign \new_[16588]_  = \new_[16587]_  & \new_[16582]_ ;
  assign \new_[16591]_  = ~A167 & ~A169;
  assign \new_[16595]_  = A200 & ~A199;
  assign \new_[16596]_  = ~A166 & \new_[16595]_ ;
  assign \new_[16597]_  = \new_[16596]_  & \new_[16591]_ ;
  assign \new_[16601]_  = A234 & ~A233;
  assign \new_[16602]_  = A232 & \new_[16601]_ ;
  assign \new_[16606]_  = ~A300 & A298;
  assign \new_[16607]_  = A235 & \new_[16606]_ ;
  assign \new_[16608]_  = \new_[16607]_  & \new_[16602]_ ;
  assign \new_[16611]_  = ~A167 & ~A169;
  assign \new_[16615]_  = A200 & ~A199;
  assign \new_[16616]_  = ~A166 & \new_[16615]_ ;
  assign \new_[16617]_  = \new_[16616]_  & \new_[16611]_ ;
  assign \new_[16621]_  = A234 & ~A233;
  assign \new_[16622]_  = A232 & \new_[16621]_ ;
  assign \new_[16626]_  = A299 & A298;
  assign \new_[16627]_  = A235 & \new_[16626]_ ;
  assign \new_[16628]_  = \new_[16627]_  & \new_[16622]_ ;
  assign \new_[16631]_  = ~A167 & ~A169;
  assign \new_[16635]_  = A200 & ~A199;
  assign \new_[16636]_  = ~A166 & \new_[16635]_ ;
  assign \new_[16637]_  = \new_[16636]_  & \new_[16631]_ ;
  assign \new_[16641]_  = A234 & ~A233;
  assign \new_[16642]_  = A232 & \new_[16641]_ ;
  assign \new_[16646]_  = ~A299 & ~A298;
  assign \new_[16647]_  = A235 & \new_[16646]_ ;
  assign \new_[16648]_  = \new_[16647]_  & \new_[16642]_ ;
  assign \new_[16651]_  = ~A167 & ~A169;
  assign \new_[16655]_  = A200 & ~A199;
  assign \new_[16656]_  = ~A166 & \new_[16655]_ ;
  assign \new_[16657]_  = \new_[16656]_  & \new_[16651]_ ;
  assign \new_[16661]_  = A234 & ~A233;
  assign \new_[16662]_  = A232 & \new_[16661]_ ;
  assign \new_[16666]_  = A266 & ~A265;
  assign \new_[16667]_  = A235 & \new_[16666]_ ;
  assign \new_[16668]_  = \new_[16667]_  & \new_[16662]_ ;
  assign \new_[16671]_  = ~A167 & ~A169;
  assign \new_[16675]_  = A200 & ~A199;
  assign \new_[16676]_  = ~A166 & \new_[16675]_ ;
  assign \new_[16677]_  = \new_[16676]_  & \new_[16671]_ ;
  assign \new_[16681]_  = A234 & ~A233;
  assign \new_[16682]_  = A232 & \new_[16681]_ ;
  assign \new_[16686]_  = ~A300 & A298;
  assign \new_[16687]_  = A236 & \new_[16686]_ ;
  assign \new_[16688]_  = \new_[16687]_  & \new_[16682]_ ;
  assign \new_[16691]_  = ~A167 & ~A169;
  assign \new_[16695]_  = A200 & ~A199;
  assign \new_[16696]_  = ~A166 & \new_[16695]_ ;
  assign \new_[16697]_  = \new_[16696]_  & \new_[16691]_ ;
  assign \new_[16701]_  = A234 & ~A233;
  assign \new_[16702]_  = A232 & \new_[16701]_ ;
  assign \new_[16706]_  = A299 & A298;
  assign \new_[16707]_  = A236 & \new_[16706]_ ;
  assign \new_[16708]_  = \new_[16707]_  & \new_[16702]_ ;
  assign \new_[16711]_  = ~A167 & ~A169;
  assign \new_[16715]_  = A200 & ~A199;
  assign \new_[16716]_  = ~A166 & \new_[16715]_ ;
  assign \new_[16717]_  = \new_[16716]_  & \new_[16711]_ ;
  assign \new_[16721]_  = A234 & ~A233;
  assign \new_[16722]_  = A232 & \new_[16721]_ ;
  assign \new_[16726]_  = ~A299 & ~A298;
  assign \new_[16727]_  = A236 & \new_[16726]_ ;
  assign \new_[16728]_  = \new_[16727]_  & \new_[16722]_ ;
  assign \new_[16731]_  = ~A167 & ~A169;
  assign \new_[16735]_  = A200 & ~A199;
  assign \new_[16736]_  = ~A166 & \new_[16735]_ ;
  assign \new_[16737]_  = \new_[16736]_  & \new_[16731]_ ;
  assign \new_[16741]_  = A234 & ~A233;
  assign \new_[16742]_  = A232 & \new_[16741]_ ;
  assign \new_[16746]_  = A266 & ~A265;
  assign \new_[16747]_  = A236 & \new_[16746]_ ;
  assign \new_[16748]_  = \new_[16747]_  & \new_[16742]_ ;
  assign \new_[16751]_  = ~A167 & ~A169;
  assign \new_[16755]_  = A200 & ~A199;
  assign \new_[16756]_  = ~A166 & \new_[16755]_ ;
  assign \new_[16757]_  = \new_[16756]_  & \new_[16751]_ ;
  assign \new_[16761]_  = A265 & ~A233;
  assign \new_[16762]_  = ~A232 & \new_[16761]_ ;
  assign \new_[16766]_  = A299 & ~A298;
  assign \new_[16767]_  = A266 & \new_[16766]_ ;
  assign \new_[16768]_  = \new_[16767]_  & \new_[16762]_ ;
  assign \new_[16771]_  = ~A167 & ~A169;
  assign \new_[16775]_  = A200 & ~A199;
  assign \new_[16776]_  = ~A166 & \new_[16775]_ ;
  assign \new_[16777]_  = \new_[16776]_  & \new_[16771]_ ;
  assign \new_[16781]_  = ~A266 & ~A233;
  assign \new_[16782]_  = ~A232 & \new_[16781]_ ;
  assign \new_[16786]_  = A299 & ~A298;
  assign \new_[16787]_  = ~A267 & \new_[16786]_ ;
  assign \new_[16788]_  = \new_[16787]_  & \new_[16782]_ ;
  assign \new_[16791]_  = ~A167 & ~A169;
  assign \new_[16795]_  = A200 & ~A199;
  assign \new_[16796]_  = ~A166 & \new_[16795]_ ;
  assign \new_[16797]_  = \new_[16796]_  & \new_[16791]_ ;
  assign \new_[16801]_  = ~A265 & ~A233;
  assign \new_[16802]_  = ~A232 & \new_[16801]_ ;
  assign \new_[16806]_  = A299 & ~A298;
  assign \new_[16807]_  = ~A266 & \new_[16806]_ ;
  assign \new_[16808]_  = \new_[16807]_  & \new_[16802]_ ;
  assign \new_[16811]_  = ~A167 & ~A169;
  assign \new_[16815]_  = ~A200 & A199;
  assign \new_[16816]_  = ~A166 & \new_[16815]_ ;
  assign \new_[16817]_  = \new_[16816]_  & \new_[16811]_ ;
  assign \new_[16821]_  = ~A232 & A202;
  assign \new_[16822]_  = A201 & \new_[16821]_ ;
  assign \new_[16826]_  = ~A300 & ~A299;
  assign \new_[16827]_  = A233 & \new_[16826]_ ;
  assign \new_[16828]_  = \new_[16827]_  & \new_[16822]_ ;
  assign \new_[16831]_  = ~A167 & ~A169;
  assign \new_[16835]_  = ~A200 & A199;
  assign \new_[16836]_  = ~A166 & \new_[16835]_ ;
  assign \new_[16837]_  = \new_[16836]_  & \new_[16831]_ ;
  assign \new_[16841]_  = ~A232 & A202;
  assign \new_[16842]_  = A201 & \new_[16841]_ ;
  assign \new_[16846]_  = A299 & A298;
  assign \new_[16847]_  = A233 & \new_[16846]_ ;
  assign \new_[16848]_  = \new_[16847]_  & \new_[16842]_ ;
  assign \new_[16851]_  = ~A167 & ~A169;
  assign \new_[16855]_  = ~A200 & A199;
  assign \new_[16856]_  = ~A166 & \new_[16855]_ ;
  assign \new_[16857]_  = \new_[16856]_  & \new_[16851]_ ;
  assign \new_[16861]_  = ~A232 & A202;
  assign \new_[16862]_  = A201 & \new_[16861]_ ;
  assign \new_[16866]_  = ~A299 & ~A298;
  assign \new_[16867]_  = A233 & \new_[16866]_ ;
  assign \new_[16868]_  = \new_[16867]_  & \new_[16862]_ ;
  assign \new_[16871]_  = ~A167 & ~A169;
  assign \new_[16875]_  = ~A200 & A199;
  assign \new_[16876]_  = ~A166 & \new_[16875]_ ;
  assign \new_[16877]_  = \new_[16876]_  & \new_[16871]_ ;
  assign \new_[16881]_  = ~A232 & A202;
  assign \new_[16882]_  = A201 & \new_[16881]_ ;
  assign \new_[16886]_  = A266 & ~A265;
  assign \new_[16887]_  = A233 & \new_[16886]_ ;
  assign \new_[16888]_  = \new_[16887]_  & \new_[16882]_ ;
  assign \new_[16891]_  = ~A167 & ~A169;
  assign \new_[16895]_  = ~A200 & A199;
  assign \new_[16896]_  = ~A166 & \new_[16895]_ ;
  assign \new_[16897]_  = \new_[16896]_  & \new_[16891]_ ;
  assign \new_[16901]_  = ~A232 & A203;
  assign \new_[16902]_  = A201 & \new_[16901]_ ;
  assign \new_[16906]_  = ~A300 & ~A299;
  assign \new_[16907]_  = A233 & \new_[16906]_ ;
  assign \new_[16908]_  = \new_[16907]_  & \new_[16902]_ ;
  assign \new_[16911]_  = ~A167 & ~A169;
  assign \new_[16915]_  = ~A200 & A199;
  assign \new_[16916]_  = ~A166 & \new_[16915]_ ;
  assign \new_[16917]_  = \new_[16916]_  & \new_[16911]_ ;
  assign \new_[16921]_  = ~A232 & A203;
  assign \new_[16922]_  = A201 & \new_[16921]_ ;
  assign \new_[16926]_  = A299 & A298;
  assign \new_[16927]_  = A233 & \new_[16926]_ ;
  assign \new_[16928]_  = \new_[16927]_  & \new_[16922]_ ;
  assign \new_[16931]_  = ~A167 & ~A169;
  assign \new_[16935]_  = ~A200 & A199;
  assign \new_[16936]_  = ~A166 & \new_[16935]_ ;
  assign \new_[16937]_  = \new_[16936]_  & \new_[16931]_ ;
  assign \new_[16941]_  = ~A232 & A203;
  assign \new_[16942]_  = A201 & \new_[16941]_ ;
  assign \new_[16946]_  = ~A299 & ~A298;
  assign \new_[16947]_  = A233 & \new_[16946]_ ;
  assign \new_[16948]_  = \new_[16947]_  & \new_[16942]_ ;
  assign \new_[16951]_  = ~A167 & ~A169;
  assign \new_[16955]_  = ~A200 & A199;
  assign \new_[16956]_  = ~A166 & \new_[16955]_ ;
  assign \new_[16957]_  = \new_[16956]_  & \new_[16951]_ ;
  assign \new_[16961]_  = ~A232 & A203;
  assign \new_[16962]_  = A201 & \new_[16961]_ ;
  assign \new_[16966]_  = A266 & ~A265;
  assign \new_[16967]_  = A233 & \new_[16966]_ ;
  assign \new_[16968]_  = \new_[16967]_  & \new_[16962]_ ;
  assign \new_[16971]_  = ~A168 & ~A169;
  assign \new_[16975]_  = ~A199 & A166;
  assign \new_[16976]_  = A167 & \new_[16975]_ ;
  assign \new_[16977]_  = \new_[16976]_  & \new_[16971]_ ;
  assign \new_[16981]_  = A233 & ~A232;
  assign \new_[16982]_  = A200 & \new_[16981]_ ;
  assign \new_[16986]_  = ~A302 & ~A301;
  assign \new_[16987]_  = ~A299 & \new_[16986]_ ;
  assign \new_[16988]_  = \new_[16987]_  & \new_[16982]_ ;
  assign \new_[16991]_  = ~A169 & A170;
  assign \new_[16995]_  = A199 & ~A166;
  assign \new_[16996]_  = A167 & \new_[16995]_ ;
  assign \new_[16997]_  = \new_[16996]_  & \new_[16991]_ ;
  assign \new_[17001]_  = A233 & ~A232;
  assign \new_[17002]_  = A200 & \new_[17001]_ ;
  assign \new_[17006]_  = ~A302 & ~A301;
  assign \new_[17007]_  = ~A299 & \new_[17006]_ ;
  assign \new_[17008]_  = \new_[17007]_  & \new_[17002]_ ;
  assign \new_[17011]_  = ~A169 & A170;
  assign \new_[17015]_  = ~A200 & ~A166;
  assign \new_[17016]_  = A167 & \new_[17015]_ ;
  assign \new_[17017]_  = \new_[17016]_  & \new_[17011]_ ;
  assign \new_[17021]_  = ~A232 & ~A203;
  assign \new_[17022]_  = ~A202 & \new_[17021]_ ;
  assign \new_[17026]_  = ~A300 & ~A299;
  assign \new_[17027]_  = A233 & \new_[17026]_ ;
  assign \new_[17028]_  = \new_[17027]_  & \new_[17022]_ ;
  assign \new_[17031]_  = ~A169 & A170;
  assign \new_[17035]_  = ~A200 & ~A166;
  assign \new_[17036]_  = A167 & \new_[17035]_ ;
  assign \new_[17037]_  = \new_[17036]_  & \new_[17031]_ ;
  assign \new_[17041]_  = ~A232 & ~A203;
  assign \new_[17042]_  = ~A202 & \new_[17041]_ ;
  assign \new_[17046]_  = A299 & A298;
  assign \new_[17047]_  = A233 & \new_[17046]_ ;
  assign \new_[17048]_  = \new_[17047]_  & \new_[17042]_ ;
  assign \new_[17051]_  = ~A169 & A170;
  assign \new_[17055]_  = ~A200 & ~A166;
  assign \new_[17056]_  = A167 & \new_[17055]_ ;
  assign \new_[17057]_  = \new_[17056]_  & \new_[17051]_ ;
  assign \new_[17061]_  = ~A232 & ~A203;
  assign \new_[17062]_  = ~A202 & \new_[17061]_ ;
  assign \new_[17066]_  = ~A299 & ~A298;
  assign \new_[17067]_  = A233 & \new_[17066]_ ;
  assign \new_[17068]_  = \new_[17067]_  & \new_[17062]_ ;
  assign \new_[17071]_  = ~A169 & A170;
  assign \new_[17075]_  = ~A200 & ~A166;
  assign \new_[17076]_  = A167 & \new_[17075]_ ;
  assign \new_[17077]_  = \new_[17076]_  & \new_[17071]_ ;
  assign \new_[17081]_  = ~A232 & ~A203;
  assign \new_[17082]_  = ~A202 & \new_[17081]_ ;
  assign \new_[17086]_  = A266 & ~A265;
  assign \new_[17087]_  = A233 & \new_[17086]_ ;
  assign \new_[17088]_  = \new_[17087]_  & \new_[17082]_ ;
  assign \new_[17091]_  = ~A169 & A170;
  assign \new_[17095]_  = ~A200 & ~A166;
  assign \new_[17096]_  = A167 & \new_[17095]_ ;
  assign \new_[17097]_  = \new_[17096]_  & \new_[17091]_ ;
  assign \new_[17101]_  = A233 & ~A232;
  assign \new_[17102]_  = ~A201 & \new_[17101]_ ;
  assign \new_[17106]_  = ~A302 & ~A301;
  assign \new_[17107]_  = ~A299 & \new_[17106]_ ;
  assign \new_[17108]_  = \new_[17107]_  & \new_[17102]_ ;
  assign \new_[17111]_  = ~A169 & A170;
  assign \new_[17115]_  = ~A199 & ~A166;
  assign \new_[17116]_  = A167 & \new_[17115]_ ;
  assign \new_[17117]_  = \new_[17116]_  & \new_[17111]_ ;
  assign \new_[17121]_  = A233 & ~A232;
  assign \new_[17122]_  = ~A200 & \new_[17121]_ ;
  assign \new_[17126]_  = ~A302 & ~A301;
  assign \new_[17127]_  = ~A299 & \new_[17126]_ ;
  assign \new_[17128]_  = \new_[17127]_  & \new_[17122]_ ;
  assign \new_[17131]_  = ~A169 & A170;
  assign \new_[17135]_  = A199 & A166;
  assign \new_[17136]_  = ~A167 & \new_[17135]_ ;
  assign \new_[17137]_  = \new_[17136]_  & \new_[17131]_ ;
  assign \new_[17141]_  = A233 & ~A232;
  assign \new_[17142]_  = A200 & \new_[17141]_ ;
  assign \new_[17146]_  = ~A302 & ~A301;
  assign \new_[17147]_  = ~A299 & \new_[17146]_ ;
  assign \new_[17148]_  = \new_[17147]_  & \new_[17142]_ ;
  assign \new_[17151]_  = ~A169 & A170;
  assign \new_[17155]_  = ~A200 & A166;
  assign \new_[17156]_  = ~A167 & \new_[17155]_ ;
  assign \new_[17157]_  = \new_[17156]_  & \new_[17151]_ ;
  assign \new_[17161]_  = ~A232 & ~A203;
  assign \new_[17162]_  = ~A202 & \new_[17161]_ ;
  assign \new_[17166]_  = ~A300 & ~A299;
  assign \new_[17167]_  = A233 & \new_[17166]_ ;
  assign \new_[17168]_  = \new_[17167]_  & \new_[17162]_ ;
  assign \new_[17171]_  = ~A169 & A170;
  assign \new_[17175]_  = ~A200 & A166;
  assign \new_[17176]_  = ~A167 & \new_[17175]_ ;
  assign \new_[17177]_  = \new_[17176]_  & \new_[17171]_ ;
  assign \new_[17181]_  = ~A232 & ~A203;
  assign \new_[17182]_  = ~A202 & \new_[17181]_ ;
  assign \new_[17186]_  = A299 & A298;
  assign \new_[17187]_  = A233 & \new_[17186]_ ;
  assign \new_[17188]_  = \new_[17187]_  & \new_[17182]_ ;
  assign \new_[17191]_  = ~A169 & A170;
  assign \new_[17195]_  = ~A200 & A166;
  assign \new_[17196]_  = ~A167 & \new_[17195]_ ;
  assign \new_[17197]_  = \new_[17196]_  & \new_[17191]_ ;
  assign \new_[17201]_  = ~A232 & ~A203;
  assign \new_[17202]_  = ~A202 & \new_[17201]_ ;
  assign \new_[17206]_  = ~A299 & ~A298;
  assign \new_[17207]_  = A233 & \new_[17206]_ ;
  assign \new_[17208]_  = \new_[17207]_  & \new_[17202]_ ;
  assign \new_[17211]_  = ~A169 & A170;
  assign \new_[17215]_  = ~A200 & A166;
  assign \new_[17216]_  = ~A167 & \new_[17215]_ ;
  assign \new_[17217]_  = \new_[17216]_  & \new_[17211]_ ;
  assign \new_[17221]_  = ~A232 & ~A203;
  assign \new_[17222]_  = ~A202 & \new_[17221]_ ;
  assign \new_[17226]_  = A266 & ~A265;
  assign \new_[17227]_  = A233 & \new_[17226]_ ;
  assign \new_[17228]_  = \new_[17227]_  & \new_[17222]_ ;
  assign \new_[17231]_  = ~A169 & A170;
  assign \new_[17235]_  = ~A200 & A166;
  assign \new_[17236]_  = ~A167 & \new_[17235]_ ;
  assign \new_[17237]_  = \new_[17236]_  & \new_[17231]_ ;
  assign \new_[17241]_  = A233 & ~A232;
  assign \new_[17242]_  = ~A201 & \new_[17241]_ ;
  assign \new_[17246]_  = ~A302 & ~A301;
  assign \new_[17247]_  = ~A299 & \new_[17246]_ ;
  assign \new_[17248]_  = \new_[17247]_  & \new_[17242]_ ;
  assign \new_[17251]_  = ~A169 & A170;
  assign \new_[17255]_  = ~A199 & A166;
  assign \new_[17256]_  = ~A167 & \new_[17255]_ ;
  assign \new_[17257]_  = \new_[17256]_  & \new_[17251]_ ;
  assign \new_[17261]_  = A233 & ~A232;
  assign \new_[17262]_  = ~A200 & \new_[17261]_ ;
  assign \new_[17266]_  = ~A302 & ~A301;
  assign \new_[17267]_  = ~A299 & \new_[17266]_ ;
  assign \new_[17268]_  = \new_[17267]_  & \new_[17262]_ ;
  assign \new_[17271]_  = ~A169 & ~A170;
  assign \new_[17275]_  = ~A200 & A199;
  assign \new_[17276]_  = ~A168 & \new_[17275]_ ;
  assign \new_[17277]_  = \new_[17276]_  & \new_[17271]_ ;
  assign \new_[17281]_  = ~A232 & A202;
  assign \new_[17282]_  = A201 & \new_[17281]_ ;
  assign \new_[17286]_  = ~A300 & ~A299;
  assign \new_[17287]_  = A233 & \new_[17286]_ ;
  assign \new_[17288]_  = \new_[17287]_  & \new_[17282]_ ;
  assign \new_[17291]_  = ~A169 & ~A170;
  assign \new_[17295]_  = ~A200 & A199;
  assign \new_[17296]_  = ~A168 & \new_[17295]_ ;
  assign \new_[17297]_  = \new_[17296]_  & \new_[17291]_ ;
  assign \new_[17301]_  = ~A232 & A202;
  assign \new_[17302]_  = A201 & \new_[17301]_ ;
  assign \new_[17306]_  = A299 & A298;
  assign \new_[17307]_  = A233 & \new_[17306]_ ;
  assign \new_[17308]_  = \new_[17307]_  & \new_[17302]_ ;
  assign \new_[17311]_  = ~A169 & ~A170;
  assign \new_[17315]_  = ~A200 & A199;
  assign \new_[17316]_  = ~A168 & \new_[17315]_ ;
  assign \new_[17317]_  = \new_[17316]_  & \new_[17311]_ ;
  assign \new_[17321]_  = ~A232 & A202;
  assign \new_[17322]_  = A201 & \new_[17321]_ ;
  assign \new_[17326]_  = ~A299 & ~A298;
  assign \new_[17327]_  = A233 & \new_[17326]_ ;
  assign \new_[17328]_  = \new_[17327]_  & \new_[17322]_ ;
  assign \new_[17331]_  = ~A169 & ~A170;
  assign \new_[17335]_  = ~A200 & A199;
  assign \new_[17336]_  = ~A168 & \new_[17335]_ ;
  assign \new_[17337]_  = \new_[17336]_  & \new_[17331]_ ;
  assign \new_[17341]_  = ~A232 & A202;
  assign \new_[17342]_  = A201 & \new_[17341]_ ;
  assign \new_[17346]_  = A266 & ~A265;
  assign \new_[17347]_  = A233 & \new_[17346]_ ;
  assign \new_[17348]_  = \new_[17347]_  & \new_[17342]_ ;
  assign \new_[17351]_  = ~A169 & ~A170;
  assign \new_[17355]_  = ~A200 & A199;
  assign \new_[17356]_  = ~A168 & \new_[17355]_ ;
  assign \new_[17357]_  = \new_[17356]_  & \new_[17351]_ ;
  assign \new_[17361]_  = ~A232 & A203;
  assign \new_[17362]_  = A201 & \new_[17361]_ ;
  assign \new_[17366]_  = ~A300 & ~A299;
  assign \new_[17367]_  = A233 & \new_[17366]_ ;
  assign \new_[17368]_  = \new_[17367]_  & \new_[17362]_ ;
  assign \new_[17371]_  = ~A169 & ~A170;
  assign \new_[17375]_  = ~A200 & A199;
  assign \new_[17376]_  = ~A168 & \new_[17375]_ ;
  assign \new_[17377]_  = \new_[17376]_  & \new_[17371]_ ;
  assign \new_[17381]_  = ~A232 & A203;
  assign \new_[17382]_  = A201 & \new_[17381]_ ;
  assign \new_[17386]_  = A299 & A298;
  assign \new_[17387]_  = A233 & \new_[17386]_ ;
  assign \new_[17388]_  = \new_[17387]_  & \new_[17382]_ ;
  assign \new_[17391]_  = ~A169 & ~A170;
  assign \new_[17395]_  = ~A200 & A199;
  assign \new_[17396]_  = ~A168 & \new_[17395]_ ;
  assign \new_[17397]_  = \new_[17396]_  & \new_[17391]_ ;
  assign \new_[17401]_  = ~A232 & A203;
  assign \new_[17402]_  = A201 & \new_[17401]_ ;
  assign \new_[17406]_  = ~A299 & ~A298;
  assign \new_[17407]_  = A233 & \new_[17406]_ ;
  assign \new_[17408]_  = \new_[17407]_  & \new_[17402]_ ;
  assign \new_[17411]_  = ~A169 & ~A170;
  assign \new_[17415]_  = ~A200 & A199;
  assign \new_[17416]_  = ~A168 & \new_[17415]_ ;
  assign \new_[17417]_  = \new_[17416]_  & \new_[17411]_ ;
  assign \new_[17421]_  = ~A232 & A203;
  assign \new_[17422]_  = A201 & \new_[17421]_ ;
  assign \new_[17426]_  = A266 & ~A265;
  assign \new_[17427]_  = A233 & \new_[17426]_ ;
  assign \new_[17428]_  = \new_[17427]_  & \new_[17422]_ ;
  assign \new_[17432]_  = A199 & A166;
  assign \new_[17433]_  = A168 & \new_[17432]_ ;
  assign \new_[17437]_  = A233 & A232;
  assign \new_[17438]_  = A200 & \new_[17437]_ ;
  assign \new_[17439]_  = \new_[17438]_  & \new_[17433]_ ;
  assign \new_[17443]_  = A298 & ~A267;
  assign \new_[17444]_  = A265 & \new_[17443]_ ;
  assign \new_[17448]_  = A301 & A300;
  assign \new_[17449]_  = ~A299 & \new_[17448]_ ;
  assign \new_[17450]_  = \new_[17449]_  & \new_[17444]_ ;
  assign \new_[17454]_  = A199 & A166;
  assign \new_[17455]_  = A168 & \new_[17454]_ ;
  assign \new_[17459]_  = A233 & A232;
  assign \new_[17460]_  = A200 & \new_[17459]_ ;
  assign \new_[17461]_  = \new_[17460]_  & \new_[17455]_ ;
  assign \new_[17465]_  = A298 & ~A267;
  assign \new_[17466]_  = A265 & \new_[17465]_ ;
  assign \new_[17470]_  = A302 & A300;
  assign \new_[17471]_  = ~A299 & \new_[17470]_ ;
  assign \new_[17472]_  = \new_[17471]_  & \new_[17466]_ ;
  assign \new_[17476]_  = A199 & A166;
  assign \new_[17477]_  = A168 & \new_[17476]_ ;
  assign \new_[17481]_  = A233 & A232;
  assign \new_[17482]_  = A200 & \new_[17481]_ ;
  assign \new_[17483]_  = \new_[17482]_  & \new_[17477]_ ;
  assign \new_[17487]_  = A298 & A266;
  assign \new_[17488]_  = A265 & \new_[17487]_ ;
  assign \new_[17492]_  = A301 & A300;
  assign \new_[17493]_  = ~A299 & \new_[17492]_ ;
  assign \new_[17494]_  = \new_[17493]_  & \new_[17488]_ ;
  assign \new_[17498]_  = A199 & A166;
  assign \new_[17499]_  = A168 & \new_[17498]_ ;
  assign \new_[17503]_  = A233 & A232;
  assign \new_[17504]_  = A200 & \new_[17503]_ ;
  assign \new_[17505]_  = \new_[17504]_  & \new_[17499]_ ;
  assign \new_[17509]_  = A298 & A266;
  assign \new_[17510]_  = A265 & \new_[17509]_ ;
  assign \new_[17514]_  = A302 & A300;
  assign \new_[17515]_  = ~A299 & \new_[17514]_ ;
  assign \new_[17516]_  = \new_[17515]_  & \new_[17510]_ ;
  assign \new_[17520]_  = A199 & A166;
  assign \new_[17521]_  = A168 & \new_[17520]_ ;
  assign \new_[17525]_  = A233 & A232;
  assign \new_[17526]_  = A200 & \new_[17525]_ ;
  assign \new_[17527]_  = \new_[17526]_  & \new_[17521]_ ;
  assign \new_[17531]_  = A298 & ~A266;
  assign \new_[17532]_  = ~A265 & \new_[17531]_ ;
  assign \new_[17536]_  = A301 & A300;
  assign \new_[17537]_  = ~A299 & \new_[17536]_ ;
  assign \new_[17538]_  = \new_[17537]_  & \new_[17532]_ ;
  assign \new_[17542]_  = A199 & A166;
  assign \new_[17543]_  = A168 & \new_[17542]_ ;
  assign \new_[17547]_  = A233 & A232;
  assign \new_[17548]_  = A200 & \new_[17547]_ ;
  assign \new_[17549]_  = \new_[17548]_  & \new_[17543]_ ;
  assign \new_[17553]_  = A298 & ~A266;
  assign \new_[17554]_  = ~A265 & \new_[17553]_ ;
  assign \new_[17558]_  = A302 & A300;
  assign \new_[17559]_  = ~A299 & \new_[17558]_ ;
  assign \new_[17560]_  = \new_[17559]_  & \new_[17554]_ ;
  assign \new_[17564]_  = A199 & A166;
  assign \new_[17565]_  = A168 & \new_[17564]_ ;
  assign \new_[17569]_  = ~A235 & ~A233;
  assign \new_[17570]_  = A200 & \new_[17569]_ ;
  assign \new_[17571]_  = \new_[17570]_  & \new_[17565]_ ;
  assign \new_[17575]_  = ~A268 & ~A266;
  assign \new_[17576]_  = ~A236 & \new_[17575]_ ;
  assign \new_[17580]_  = A299 & ~A298;
  assign \new_[17581]_  = ~A269 & \new_[17580]_ ;
  assign \new_[17582]_  = \new_[17581]_  & \new_[17576]_ ;
  assign \new_[17586]_  = A199 & A166;
  assign \new_[17587]_  = A168 & \new_[17586]_ ;
  assign \new_[17591]_  = ~A234 & ~A233;
  assign \new_[17592]_  = A200 & \new_[17591]_ ;
  assign \new_[17593]_  = \new_[17592]_  & \new_[17587]_ ;
  assign \new_[17597]_  = A298 & A266;
  assign \new_[17598]_  = A265 & \new_[17597]_ ;
  assign \new_[17602]_  = A301 & A300;
  assign \new_[17603]_  = ~A299 & \new_[17602]_ ;
  assign \new_[17604]_  = \new_[17603]_  & \new_[17598]_ ;
  assign \new_[17608]_  = A199 & A166;
  assign \new_[17609]_  = A168 & \new_[17608]_ ;
  assign \new_[17613]_  = ~A234 & ~A233;
  assign \new_[17614]_  = A200 & \new_[17613]_ ;
  assign \new_[17615]_  = \new_[17614]_  & \new_[17609]_ ;
  assign \new_[17619]_  = A298 & A266;
  assign \new_[17620]_  = A265 & \new_[17619]_ ;
  assign \new_[17624]_  = A302 & A300;
  assign \new_[17625]_  = ~A299 & \new_[17624]_ ;
  assign \new_[17626]_  = \new_[17625]_  & \new_[17620]_ ;
  assign \new_[17630]_  = A199 & A166;
  assign \new_[17631]_  = A168 & \new_[17630]_ ;
  assign \new_[17635]_  = ~A234 & ~A233;
  assign \new_[17636]_  = A200 & \new_[17635]_ ;
  assign \new_[17637]_  = \new_[17636]_  & \new_[17631]_ ;
  assign \new_[17641]_  = A298 & ~A267;
  assign \new_[17642]_  = ~A266 & \new_[17641]_ ;
  assign \new_[17646]_  = A301 & A300;
  assign \new_[17647]_  = ~A299 & \new_[17646]_ ;
  assign \new_[17648]_  = \new_[17647]_  & \new_[17642]_ ;
  assign \new_[17652]_  = A199 & A166;
  assign \new_[17653]_  = A168 & \new_[17652]_ ;
  assign \new_[17657]_  = ~A234 & ~A233;
  assign \new_[17658]_  = A200 & \new_[17657]_ ;
  assign \new_[17659]_  = \new_[17658]_  & \new_[17653]_ ;
  assign \new_[17663]_  = A298 & ~A267;
  assign \new_[17664]_  = ~A266 & \new_[17663]_ ;
  assign \new_[17668]_  = A302 & A300;
  assign \new_[17669]_  = ~A299 & \new_[17668]_ ;
  assign \new_[17670]_  = \new_[17669]_  & \new_[17664]_ ;
  assign \new_[17674]_  = A199 & A166;
  assign \new_[17675]_  = A168 & \new_[17674]_ ;
  assign \new_[17679]_  = ~A234 & ~A233;
  assign \new_[17680]_  = A200 & \new_[17679]_ ;
  assign \new_[17681]_  = \new_[17680]_  & \new_[17675]_ ;
  assign \new_[17685]_  = A298 & ~A266;
  assign \new_[17686]_  = ~A265 & \new_[17685]_ ;
  assign \new_[17690]_  = A301 & A300;
  assign \new_[17691]_  = ~A299 & \new_[17690]_ ;
  assign \new_[17692]_  = \new_[17691]_  & \new_[17686]_ ;
  assign \new_[17696]_  = A199 & A166;
  assign \new_[17697]_  = A168 & \new_[17696]_ ;
  assign \new_[17701]_  = ~A234 & ~A233;
  assign \new_[17702]_  = A200 & \new_[17701]_ ;
  assign \new_[17703]_  = \new_[17702]_  & \new_[17697]_ ;
  assign \new_[17707]_  = A298 & ~A266;
  assign \new_[17708]_  = ~A265 & \new_[17707]_ ;
  assign \new_[17712]_  = A302 & A300;
  assign \new_[17713]_  = ~A299 & \new_[17712]_ ;
  assign \new_[17714]_  = \new_[17713]_  & \new_[17708]_ ;
  assign \new_[17718]_  = A199 & A166;
  assign \new_[17719]_  = A168 & \new_[17718]_ ;
  assign \new_[17723]_  = ~A233 & A232;
  assign \new_[17724]_  = A200 & \new_[17723]_ ;
  assign \new_[17725]_  = \new_[17724]_  & \new_[17719]_ ;
  assign \new_[17729]_  = A265 & A235;
  assign \new_[17730]_  = A234 & \new_[17729]_ ;
  assign \new_[17734]_  = A268 & A267;
  assign \new_[17735]_  = ~A266 & \new_[17734]_ ;
  assign \new_[17736]_  = \new_[17735]_  & \new_[17730]_ ;
  assign \new_[17740]_  = A199 & A166;
  assign \new_[17741]_  = A168 & \new_[17740]_ ;
  assign \new_[17745]_  = ~A233 & A232;
  assign \new_[17746]_  = A200 & \new_[17745]_ ;
  assign \new_[17747]_  = \new_[17746]_  & \new_[17741]_ ;
  assign \new_[17751]_  = A265 & A235;
  assign \new_[17752]_  = A234 & \new_[17751]_ ;
  assign \new_[17756]_  = A269 & A267;
  assign \new_[17757]_  = ~A266 & \new_[17756]_ ;
  assign \new_[17758]_  = \new_[17757]_  & \new_[17752]_ ;
  assign \new_[17762]_  = A199 & A166;
  assign \new_[17763]_  = A168 & \new_[17762]_ ;
  assign \new_[17767]_  = ~A233 & A232;
  assign \new_[17768]_  = A200 & \new_[17767]_ ;
  assign \new_[17769]_  = \new_[17768]_  & \new_[17763]_ ;
  assign \new_[17773]_  = A265 & A236;
  assign \new_[17774]_  = A234 & \new_[17773]_ ;
  assign \new_[17778]_  = A268 & A267;
  assign \new_[17779]_  = ~A266 & \new_[17778]_ ;
  assign \new_[17780]_  = \new_[17779]_  & \new_[17774]_ ;
  assign \new_[17784]_  = A199 & A166;
  assign \new_[17785]_  = A168 & \new_[17784]_ ;
  assign \new_[17789]_  = ~A233 & A232;
  assign \new_[17790]_  = A200 & \new_[17789]_ ;
  assign \new_[17791]_  = \new_[17790]_  & \new_[17785]_ ;
  assign \new_[17795]_  = A265 & A236;
  assign \new_[17796]_  = A234 & \new_[17795]_ ;
  assign \new_[17800]_  = A269 & A267;
  assign \new_[17801]_  = ~A266 & \new_[17800]_ ;
  assign \new_[17802]_  = \new_[17801]_  & \new_[17796]_ ;
  assign \new_[17806]_  = A199 & A166;
  assign \new_[17807]_  = A168 & \new_[17806]_ ;
  assign \new_[17811]_  = ~A233 & ~A232;
  assign \new_[17812]_  = A200 & \new_[17811]_ ;
  assign \new_[17813]_  = \new_[17812]_  & \new_[17807]_ ;
  assign \new_[17817]_  = A298 & A266;
  assign \new_[17818]_  = A265 & \new_[17817]_ ;
  assign \new_[17822]_  = A301 & A300;
  assign \new_[17823]_  = ~A299 & \new_[17822]_ ;
  assign \new_[17824]_  = \new_[17823]_  & \new_[17818]_ ;
  assign \new_[17828]_  = A199 & A166;
  assign \new_[17829]_  = A168 & \new_[17828]_ ;
  assign \new_[17833]_  = ~A233 & ~A232;
  assign \new_[17834]_  = A200 & \new_[17833]_ ;
  assign \new_[17835]_  = \new_[17834]_  & \new_[17829]_ ;
  assign \new_[17839]_  = A298 & A266;
  assign \new_[17840]_  = A265 & \new_[17839]_ ;
  assign \new_[17844]_  = A302 & A300;
  assign \new_[17845]_  = ~A299 & \new_[17844]_ ;
  assign \new_[17846]_  = \new_[17845]_  & \new_[17840]_ ;
  assign \new_[17850]_  = A199 & A166;
  assign \new_[17851]_  = A168 & \new_[17850]_ ;
  assign \new_[17855]_  = ~A233 & ~A232;
  assign \new_[17856]_  = A200 & \new_[17855]_ ;
  assign \new_[17857]_  = \new_[17856]_  & \new_[17851]_ ;
  assign \new_[17861]_  = A298 & ~A267;
  assign \new_[17862]_  = ~A266 & \new_[17861]_ ;
  assign \new_[17866]_  = A301 & A300;
  assign \new_[17867]_  = ~A299 & \new_[17866]_ ;
  assign \new_[17868]_  = \new_[17867]_  & \new_[17862]_ ;
  assign \new_[17872]_  = A199 & A166;
  assign \new_[17873]_  = A168 & \new_[17872]_ ;
  assign \new_[17877]_  = ~A233 & ~A232;
  assign \new_[17878]_  = A200 & \new_[17877]_ ;
  assign \new_[17879]_  = \new_[17878]_  & \new_[17873]_ ;
  assign \new_[17883]_  = A298 & ~A267;
  assign \new_[17884]_  = ~A266 & \new_[17883]_ ;
  assign \new_[17888]_  = A302 & A300;
  assign \new_[17889]_  = ~A299 & \new_[17888]_ ;
  assign \new_[17890]_  = \new_[17889]_  & \new_[17884]_ ;
  assign \new_[17894]_  = A199 & A166;
  assign \new_[17895]_  = A168 & \new_[17894]_ ;
  assign \new_[17899]_  = ~A233 & ~A232;
  assign \new_[17900]_  = A200 & \new_[17899]_ ;
  assign \new_[17901]_  = \new_[17900]_  & \new_[17895]_ ;
  assign \new_[17905]_  = A298 & ~A266;
  assign \new_[17906]_  = ~A265 & \new_[17905]_ ;
  assign \new_[17910]_  = A301 & A300;
  assign \new_[17911]_  = ~A299 & \new_[17910]_ ;
  assign \new_[17912]_  = \new_[17911]_  & \new_[17906]_ ;
  assign \new_[17916]_  = A199 & A166;
  assign \new_[17917]_  = A168 & \new_[17916]_ ;
  assign \new_[17921]_  = ~A233 & ~A232;
  assign \new_[17922]_  = A200 & \new_[17921]_ ;
  assign \new_[17923]_  = \new_[17922]_  & \new_[17917]_ ;
  assign \new_[17927]_  = A298 & ~A266;
  assign \new_[17928]_  = ~A265 & \new_[17927]_ ;
  assign \new_[17932]_  = A302 & A300;
  assign \new_[17933]_  = ~A299 & \new_[17932]_ ;
  assign \new_[17934]_  = \new_[17933]_  & \new_[17928]_ ;
  assign \new_[17938]_  = ~A200 & A166;
  assign \new_[17939]_  = A168 & \new_[17938]_ ;
  assign \new_[17943]_  = A232 & ~A203;
  assign \new_[17944]_  = ~A202 & \new_[17943]_ ;
  assign \new_[17945]_  = \new_[17944]_  & \new_[17939]_ ;
  assign \new_[17949]_  = ~A268 & A265;
  assign \new_[17950]_  = A233 & \new_[17949]_ ;
  assign \new_[17954]_  = A299 & ~A298;
  assign \new_[17955]_  = ~A269 & \new_[17954]_ ;
  assign \new_[17956]_  = \new_[17955]_  & \new_[17950]_ ;
  assign \new_[17960]_  = ~A200 & A166;
  assign \new_[17961]_  = A168 & \new_[17960]_ ;
  assign \new_[17965]_  = ~A233 & ~A203;
  assign \new_[17966]_  = ~A202 & \new_[17965]_ ;
  assign \new_[17967]_  = \new_[17966]_  & \new_[17961]_ ;
  assign \new_[17971]_  = A265 & ~A236;
  assign \new_[17972]_  = ~A235 & \new_[17971]_ ;
  assign \new_[17976]_  = A299 & ~A298;
  assign \new_[17977]_  = A266 & \new_[17976]_ ;
  assign \new_[17978]_  = \new_[17977]_  & \new_[17972]_ ;
  assign \new_[17982]_  = ~A200 & A166;
  assign \new_[17983]_  = A168 & \new_[17982]_ ;
  assign \new_[17987]_  = ~A233 & ~A203;
  assign \new_[17988]_  = ~A202 & \new_[17987]_ ;
  assign \new_[17989]_  = \new_[17988]_  & \new_[17983]_ ;
  assign \new_[17993]_  = ~A266 & ~A236;
  assign \new_[17994]_  = ~A235 & \new_[17993]_ ;
  assign \new_[17998]_  = A299 & ~A298;
  assign \new_[17999]_  = ~A267 & \new_[17998]_ ;
  assign \new_[18000]_  = \new_[17999]_  & \new_[17994]_ ;
  assign \new_[18004]_  = ~A200 & A166;
  assign \new_[18005]_  = A168 & \new_[18004]_ ;
  assign \new_[18009]_  = ~A233 & ~A203;
  assign \new_[18010]_  = ~A202 & \new_[18009]_ ;
  assign \new_[18011]_  = \new_[18010]_  & \new_[18005]_ ;
  assign \new_[18015]_  = ~A265 & ~A236;
  assign \new_[18016]_  = ~A235 & \new_[18015]_ ;
  assign \new_[18020]_  = A299 & ~A298;
  assign \new_[18021]_  = ~A266 & \new_[18020]_ ;
  assign \new_[18022]_  = \new_[18021]_  & \new_[18016]_ ;
  assign \new_[18026]_  = ~A200 & A166;
  assign \new_[18027]_  = A168 & \new_[18026]_ ;
  assign \new_[18031]_  = ~A233 & ~A203;
  assign \new_[18032]_  = ~A202 & \new_[18031]_ ;
  assign \new_[18033]_  = \new_[18032]_  & \new_[18027]_ ;
  assign \new_[18037]_  = ~A268 & ~A266;
  assign \new_[18038]_  = ~A234 & \new_[18037]_ ;
  assign \new_[18042]_  = A299 & ~A298;
  assign \new_[18043]_  = ~A269 & \new_[18042]_ ;
  assign \new_[18044]_  = \new_[18043]_  & \new_[18038]_ ;
  assign \new_[18048]_  = ~A200 & A166;
  assign \new_[18049]_  = A168 & \new_[18048]_ ;
  assign \new_[18053]_  = A232 & ~A203;
  assign \new_[18054]_  = ~A202 & \new_[18053]_ ;
  assign \new_[18055]_  = \new_[18054]_  & \new_[18049]_ ;
  assign \new_[18059]_  = A235 & A234;
  assign \new_[18060]_  = ~A233 & \new_[18059]_ ;
  assign \new_[18064]_  = ~A302 & ~A301;
  assign \new_[18065]_  = A298 & \new_[18064]_ ;
  assign \new_[18066]_  = \new_[18065]_  & \new_[18060]_ ;
  assign \new_[18070]_  = ~A200 & A166;
  assign \new_[18071]_  = A168 & \new_[18070]_ ;
  assign \new_[18075]_  = A232 & ~A203;
  assign \new_[18076]_  = ~A202 & \new_[18075]_ ;
  assign \new_[18077]_  = \new_[18076]_  & \new_[18071]_ ;
  assign \new_[18081]_  = A236 & A234;
  assign \new_[18082]_  = ~A233 & \new_[18081]_ ;
  assign \new_[18086]_  = ~A302 & ~A301;
  assign \new_[18087]_  = A298 & \new_[18086]_ ;
  assign \new_[18088]_  = \new_[18087]_  & \new_[18082]_ ;
  assign \new_[18092]_  = ~A200 & A166;
  assign \new_[18093]_  = A168 & \new_[18092]_ ;
  assign \new_[18097]_  = ~A232 & ~A203;
  assign \new_[18098]_  = ~A202 & \new_[18097]_ ;
  assign \new_[18099]_  = \new_[18098]_  & \new_[18093]_ ;
  assign \new_[18103]_  = ~A268 & ~A266;
  assign \new_[18104]_  = ~A233 & \new_[18103]_ ;
  assign \new_[18108]_  = A299 & ~A298;
  assign \new_[18109]_  = ~A269 & \new_[18108]_ ;
  assign \new_[18110]_  = \new_[18109]_  & \new_[18104]_ ;
  assign \new_[18114]_  = ~A200 & A166;
  assign \new_[18115]_  = A168 & \new_[18114]_ ;
  assign \new_[18119]_  = A233 & A232;
  assign \new_[18120]_  = ~A201 & \new_[18119]_ ;
  assign \new_[18121]_  = \new_[18120]_  & \new_[18115]_ ;
  assign \new_[18125]_  = A298 & ~A267;
  assign \new_[18126]_  = A265 & \new_[18125]_ ;
  assign \new_[18130]_  = A301 & A300;
  assign \new_[18131]_  = ~A299 & \new_[18130]_ ;
  assign \new_[18132]_  = \new_[18131]_  & \new_[18126]_ ;
  assign \new_[18136]_  = ~A200 & A166;
  assign \new_[18137]_  = A168 & \new_[18136]_ ;
  assign \new_[18141]_  = A233 & A232;
  assign \new_[18142]_  = ~A201 & \new_[18141]_ ;
  assign \new_[18143]_  = \new_[18142]_  & \new_[18137]_ ;
  assign \new_[18147]_  = A298 & ~A267;
  assign \new_[18148]_  = A265 & \new_[18147]_ ;
  assign \new_[18152]_  = A302 & A300;
  assign \new_[18153]_  = ~A299 & \new_[18152]_ ;
  assign \new_[18154]_  = \new_[18153]_  & \new_[18148]_ ;
  assign \new_[18158]_  = ~A200 & A166;
  assign \new_[18159]_  = A168 & \new_[18158]_ ;
  assign \new_[18163]_  = A233 & A232;
  assign \new_[18164]_  = ~A201 & \new_[18163]_ ;
  assign \new_[18165]_  = \new_[18164]_  & \new_[18159]_ ;
  assign \new_[18169]_  = A298 & A266;
  assign \new_[18170]_  = A265 & \new_[18169]_ ;
  assign \new_[18174]_  = A301 & A300;
  assign \new_[18175]_  = ~A299 & \new_[18174]_ ;
  assign \new_[18176]_  = \new_[18175]_  & \new_[18170]_ ;
  assign \new_[18180]_  = ~A200 & A166;
  assign \new_[18181]_  = A168 & \new_[18180]_ ;
  assign \new_[18185]_  = A233 & A232;
  assign \new_[18186]_  = ~A201 & \new_[18185]_ ;
  assign \new_[18187]_  = \new_[18186]_  & \new_[18181]_ ;
  assign \new_[18191]_  = A298 & A266;
  assign \new_[18192]_  = A265 & \new_[18191]_ ;
  assign \new_[18196]_  = A302 & A300;
  assign \new_[18197]_  = ~A299 & \new_[18196]_ ;
  assign \new_[18198]_  = \new_[18197]_  & \new_[18192]_ ;
  assign \new_[18202]_  = ~A200 & A166;
  assign \new_[18203]_  = A168 & \new_[18202]_ ;
  assign \new_[18207]_  = A233 & A232;
  assign \new_[18208]_  = ~A201 & \new_[18207]_ ;
  assign \new_[18209]_  = \new_[18208]_  & \new_[18203]_ ;
  assign \new_[18213]_  = A298 & ~A266;
  assign \new_[18214]_  = ~A265 & \new_[18213]_ ;
  assign \new_[18218]_  = A301 & A300;
  assign \new_[18219]_  = ~A299 & \new_[18218]_ ;
  assign \new_[18220]_  = \new_[18219]_  & \new_[18214]_ ;
  assign \new_[18224]_  = ~A200 & A166;
  assign \new_[18225]_  = A168 & \new_[18224]_ ;
  assign \new_[18229]_  = A233 & A232;
  assign \new_[18230]_  = ~A201 & \new_[18229]_ ;
  assign \new_[18231]_  = \new_[18230]_  & \new_[18225]_ ;
  assign \new_[18235]_  = A298 & ~A266;
  assign \new_[18236]_  = ~A265 & \new_[18235]_ ;
  assign \new_[18240]_  = A302 & A300;
  assign \new_[18241]_  = ~A299 & \new_[18240]_ ;
  assign \new_[18242]_  = \new_[18241]_  & \new_[18236]_ ;
  assign \new_[18246]_  = ~A200 & A166;
  assign \new_[18247]_  = A168 & \new_[18246]_ ;
  assign \new_[18251]_  = ~A235 & ~A233;
  assign \new_[18252]_  = ~A201 & \new_[18251]_ ;
  assign \new_[18253]_  = \new_[18252]_  & \new_[18247]_ ;
  assign \new_[18257]_  = ~A268 & ~A266;
  assign \new_[18258]_  = ~A236 & \new_[18257]_ ;
  assign \new_[18262]_  = A299 & ~A298;
  assign \new_[18263]_  = ~A269 & \new_[18262]_ ;
  assign \new_[18264]_  = \new_[18263]_  & \new_[18258]_ ;
  assign \new_[18268]_  = ~A200 & A166;
  assign \new_[18269]_  = A168 & \new_[18268]_ ;
  assign \new_[18273]_  = ~A234 & ~A233;
  assign \new_[18274]_  = ~A201 & \new_[18273]_ ;
  assign \new_[18275]_  = \new_[18274]_  & \new_[18269]_ ;
  assign \new_[18279]_  = A298 & A266;
  assign \new_[18280]_  = A265 & \new_[18279]_ ;
  assign \new_[18284]_  = A301 & A300;
  assign \new_[18285]_  = ~A299 & \new_[18284]_ ;
  assign \new_[18286]_  = \new_[18285]_  & \new_[18280]_ ;
  assign \new_[18290]_  = ~A200 & A166;
  assign \new_[18291]_  = A168 & \new_[18290]_ ;
  assign \new_[18295]_  = ~A234 & ~A233;
  assign \new_[18296]_  = ~A201 & \new_[18295]_ ;
  assign \new_[18297]_  = \new_[18296]_  & \new_[18291]_ ;
  assign \new_[18301]_  = A298 & A266;
  assign \new_[18302]_  = A265 & \new_[18301]_ ;
  assign \new_[18306]_  = A302 & A300;
  assign \new_[18307]_  = ~A299 & \new_[18306]_ ;
  assign \new_[18308]_  = \new_[18307]_  & \new_[18302]_ ;
  assign \new_[18312]_  = ~A200 & A166;
  assign \new_[18313]_  = A168 & \new_[18312]_ ;
  assign \new_[18317]_  = ~A234 & ~A233;
  assign \new_[18318]_  = ~A201 & \new_[18317]_ ;
  assign \new_[18319]_  = \new_[18318]_  & \new_[18313]_ ;
  assign \new_[18323]_  = A298 & ~A267;
  assign \new_[18324]_  = ~A266 & \new_[18323]_ ;
  assign \new_[18328]_  = A301 & A300;
  assign \new_[18329]_  = ~A299 & \new_[18328]_ ;
  assign \new_[18330]_  = \new_[18329]_  & \new_[18324]_ ;
  assign \new_[18334]_  = ~A200 & A166;
  assign \new_[18335]_  = A168 & \new_[18334]_ ;
  assign \new_[18339]_  = ~A234 & ~A233;
  assign \new_[18340]_  = ~A201 & \new_[18339]_ ;
  assign \new_[18341]_  = \new_[18340]_  & \new_[18335]_ ;
  assign \new_[18345]_  = A298 & ~A267;
  assign \new_[18346]_  = ~A266 & \new_[18345]_ ;
  assign \new_[18350]_  = A302 & A300;
  assign \new_[18351]_  = ~A299 & \new_[18350]_ ;
  assign \new_[18352]_  = \new_[18351]_  & \new_[18346]_ ;
  assign \new_[18356]_  = ~A200 & A166;
  assign \new_[18357]_  = A168 & \new_[18356]_ ;
  assign \new_[18361]_  = ~A234 & ~A233;
  assign \new_[18362]_  = ~A201 & \new_[18361]_ ;
  assign \new_[18363]_  = \new_[18362]_  & \new_[18357]_ ;
  assign \new_[18367]_  = A298 & ~A266;
  assign \new_[18368]_  = ~A265 & \new_[18367]_ ;
  assign \new_[18372]_  = A301 & A300;
  assign \new_[18373]_  = ~A299 & \new_[18372]_ ;
  assign \new_[18374]_  = \new_[18373]_  & \new_[18368]_ ;
  assign \new_[18378]_  = ~A200 & A166;
  assign \new_[18379]_  = A168 & \new_[18378]_ ;
  assign \new_[18383]_  = ~A234 & ~A233;
  assign \new_[18384]_  = ~A201 & \new_[18383]_ ;
  assign \new_[18385]_  = \new_[18384]_  & \new_[18379]_ ;
  assign \new_[18389]_  = A298 & ~A266;
  assign \new_[18390]_  = ~A265 & \new_[18389]_ ;
  assign \new_[18394]_  = A302 & A300;
  assign \new_[18395]_  = ~A299 & \new_[18394]_ ;
  assign \new_[18396]_  = \new_[18395]_  & \new_[18390]_ ;
  assign \new_[18400]_  = ~A200 & A166;
  assign \new_[18401]_  = A168 & \new_[18400]_ ;
  assign \new_[18405]_  = ~A233 & A232;
  assign \new_[18406]_  = ~A201 & \new_[18405]_ ;
  assign \new_[18407]_  = \new_[18406]_  & \new_[18401]_ ;
  assign \new_[18411]_  = A265 & A235;
  assign \new_[18412]_  = A234 & \new_[18411]_ ;
  assign \new_[18416]_  = A268 & A267;
  assign \new_[18417]_  = ~A266 & \new_[18416]_ ;
  assign \new_[18418]_  = \new_[18417]_  & \new_[18412]_ ;
  assign \new_[18422]_  = ~A200 & A166;
  assign \new_[18423]_  = A168 & \new_[18422]_ ;
  assign \new_[18427]_  = ~A233 & A232;
  assign \new_[18428]_  = ~A201 & \new_[18427]_ ;
  assign \new_[18429]_  = \new_[18428]_  & \new_[18423]_ ;
  assign \new_[18433]_  = A265 & A235;
  assign \new_[18434]_  = A234 & \new_[18433]_ ;
  assign \new_[18438]_  = A269 & A267;
  assign \new_[18439]_  = ~A266 & \new_[18438]_ ;
  assign \new_[18440]_  = \new_[18439]_  & \new_[18434]_ ;
  assign \new_[18444]_  = ~A200 & A166;
  assign \new_[18445]_  = A168 & \new_[18444]_ ;
  assign \new_[18449]_  = ~A233 & A232;
  assign \new_[18450]_  = ~A201 & \new_[18449]_ ;
  assign \new_[18451]_  = \new_[18450]_  & \new_[18445]_ ;
  assign \new_[18455]_  = A265 & A236;
  assign \new_[18456]_  = A234 & \new_[18455]_ ;
  assign \new_[18460]_  = A268 & A267;
  assign \new_[18461]_  = ~A266 & \new_[18460]_ ;
  assign \new_[18462]_  = \new_[18461]_  & \new_[18456]_ ;
  assign \new_[18466]_  = ~A200 & A166;
  assign \new_[18467]_  = A168 & \new_[18466]_ ;
  assign \new_[18471]_  = ~A233 & A232;
  assign \new_[18472]_  = ~A201 & \new_[18471]_ ;
  assign \new_[18473]_  = \new_[18472]_  & \new_[18467]_ ;
  assign \new_[18477]_  = A265 & A236;
  assign \new_[18478]_  = A234 & \new_[18477]_ ;
  assign \new_[18482]_  = A269 & A267;
  assign \new_[18483]_  = ~A266 & \new_[18482]_ ;
  assign \new_[18484]_  = \new_[18483]_  & \new_[18478]_ ;
  assign \new_[18488]_  = ~A200 & A166;
  assign \new_[18489]_  = A168 & \new_[18488]_ ;
  assign \new_[18493]_  = ~A233 & ~A232;
  assign \new_[18494]_  = ~A201 & \new_[18493]_ ;
  assign \new_[18495]_  = \new_[18494]_  & \new_[18489]_ ;
  assign \new_[18499]_  = A298 & A266;
  assign \new_[18500]_  = A265 & \new_[18499]_ ;
  assign \new_[18504]_  = A301 & A300;
  assign \new_[18505]_  = ~A299 & \new_[18504]_ ;
  assign \new_[18506]_  = \new_[18505]_  & \new_[18500]_ ;
  assign \new_[18510]_  = ~A200 & A166;
  assign \new_[18511]_  = A168 & \new_[18510]_ ;
  assign \new_[18515]_  = ~A233 & ~A232;
  assign \new_[18516]_  = ~A201 & \new_[18515]_ ;
  assign \new_[18517]_  = \new_[18516]_  & \new_[18511]_ ;
  assign \new_[18521]_  = A298 & A266;
  assign \new_[18522]_  = A265 & \new_[18521]_ ;
  assign \new_[18526]_  = A302 & A300;
  assign \new_[18527]_  = ~A299 & \new_[18526]_ ;
  assign \new_[18528]_  = \new_[18527]_  & \new_[18522]_ ;
  assign \new_[18532]_  = ~A200 & A166;
  assign \new_[18533]_  = A168 & \new_[18532]_ ;
  assign \new_[18537]_  = ~A233 & ~A232;
  assign \new_[18538]_  = ~A201 & \new_[18537]_ ;
  assign \new_[18539]_  = \new_[18538]_  & \new_[18533]_ ;
  assign \new_[18543]_  = A298 & ~A267;
  assign \new_[18544]_  = ~A266 & \new_[18543]_ ;
  assign \new_[18548]_  = A301 & A300;
  assign \new_[18549]_  = ~A299 & \new_[18548]_ ;
  assign \new_[18550]_  = \new_[18549]_  & \new_[18544]_ ;
  assign \new_[18554]_  = ~A200 & A166;
  assign \new_[18555]_  = A168 & \new_[18554]_ ;
  assign \new_[18559]_  = ~A233 & ~A232;
  assign \new_[18560]_  = ~A201 & \new_[18559]_ ;
  assign \new_[18561]_  = \new_[18560]_  & \new_[18555]_ ;
  assign \new_[18565]_  = A298 & ~A267;
  assign \new_[18566]_  = ~A266 & \new_[18565]_ ;
  assign \new_[18570]_  = A302 & A300;
  assign \new_[18571]_  = ~A299 & \new_[18570]_ ;
  assign \new_[18572]_  = \new_[18571]_  & \new_[18566]_ ;
  assign \new_[18576]_  = ~A200 & A166;
  assign \new_[18577]_  = A168 & \new_[18576]_ ;
  assign \new_[18581]_  = ~A233 & ~A232;
  assign \new_[18582]_  = ~A201 & \new_[18581]_ ;
  assign \new_[18583]_  = \new_[18582]_  & \new_[18577]_ ;
  assign \new_[18587]_  = A298 & ~A266;
  assign \new_[18588]_  = ~A265 & \new_[18587]_ ;
  assign \new_[18592]_  = A301 & A300;
  assign \new_[18593]_  = ~A299 & \new_[18592]_ ;
  assign \new_[18594]_  = \new_[18593]_  & \new_[18588]_ ;
  assign \new_[18598]_  = ~A200 & A166;
  assign \new_[18599]_  = A168 & \new_[18598]_ ;
  assign \new_[18603]_  = ~A233 & ~A232;
  assign \new_[18604]_  = ~A201 & \new_[18603]_ ;
  assign \new_[18605]_  = \new_[18604]_  & \new_[18599]_ ;
  assign \new_[18609]_  = A298 & ~A266;
  assign \new_[18610]_  = ~A265 & \new_[18609]_ ;
  assign \new_[18614]_  = A302 & A300;
  assign \new_[18615]_  = ~A299 & \new_[18614]_ ;
  assign \new_[18616]_  = \new_[18615]_  & \new_[18610]_ ;
  assign \new_[18620]_  = ~A199 & A166;
  assign \new_[18621]_  = A168 & \new_[18620]_ ;
  assign \new_[18625]_  = A233 & A232;
  assign \new_[18626]_  = ~A200 & \new_[18625]_ ;
  assign \new_[18627]_  = \new_[18626]_  & \new_[18621]_ ;
  assign \new_[18631]_  = A298 & ~A267;
  assign \new_[18632]_  = A265 & \new_[18631]_ ;
  assign \new_[18636]_  = A301 & A300;
  assign \new_[18637]_  = ~A299 & \new_[18636]_ ;
  assign \new_[18638]_  = \new_[18637]_  & \new_[18632]_ ;
  assign \new_[18642]_  = ~A199 & A166;
  assign \new_[18643]_  = A168 & \new_[18642]_ ;
  assign \new_[18647]_  = A233 & A232;
  assign \new_[18648]_  = ~A200 & \new_[18647]_ ;
  assign \new_[18649]_  = \new_[18648]_  & \new_[18643]_ ;
  assign \new_[18653]_  = A298 & ~A267;
  assign \new_[18654]_  = A265 & \new_[18653]_ ;
  assign \new_[18658]_  = A302 & A300;
  assign \new_[18659]_  = ~A299 & \new_[18658]_ ;
  assign \new_[18660]_  = \new_[18659]_  & \new_[18654]_ ;
  assign \new_[18664]_  = ~A199 & A166;
  assign \new_[18665]_  = A168 & \new_[18664]_ ;
  assign \new_[18669]_  = A233 & A232;
  assign \new_[18670]_  = ~A200 & \new_[18669]_ ;
  assign \new_[18671]_  = \new_[18670]_  & \new_[18665]_ ;
  assign \new_[18675]_  = A298 & A266;
  assign \new_[18676]_  = A265 & \new_[18675]_ ;
  assign \new_[18680]_  = A301 & A300;
  assign \new_[18681]_  = ~A299 & \new_[18680]_ ;
  assign \new_[18682]_  = \new_[18681]_  & \new_[18676]_ ;
  assign \new_[18686]_  = ~A199 & A166;
  assign \new_[18687]_  = A168 & \new_[18686]_ ;
  assign \new_[18691]_  = A233 & A232;
  assign \new_[18692]_  = ~A200 & \new_[18691]_ ;
  assign \new_[18693]_  = \new_[18692]_  & \new_[18687]_ ;
  assign \new_[18697]_  = A298 & A266;
  assign \new_[18698]_  = A265 & \new_[18697]_ ;
  assign \new_[18702]_  = A302 & A300;
  assign \new_[18703]_  = ~A299 & \new_[18702]_ ;
  assign \new_[18704]_  = \new_[18703]_  & \new_[18698]_ ;
  assign \new_[18708]_  = ~A199 & A166;
  assign \new_[18709]_  = A168 & \new_[18708]_ ;
  assign \new_[18713]_  = A233 & A232;
  assign \new_[18714]_  = ~A200 & \new_[18713]_ ;
  assign \new_[18715]_  = \new_[18714]_  & \new_[18709]_ ;
  assign \new_[18719]_  = A298 & ~A266;
  assign \new_[18720]_  = ~A265 & \new_[18719]_ ;
  assign \new_[18724]_  = A301 & A300;
  assign \new_[18725]_  = ~A299 & \new_[18724]_ ;
  assign \new_[18726]_  = \new_[18725]_  & \new_[18720]_ ;
  assign \new_[18730]_  = ~A199 & A166;
  assign \new_[18731]_  = A168 & \new_[18730]_ ;
  assign \new_[18735]_  = A233 & A232;
  assign \new_[18736]_  = ~A200 & \new_[18735]_ ;
  assign \new_[18737]_  = \new_[18736]_  & \new_[18731]_ ;
  assign \new_[18741]_  = A298 & ~A266;
  assign \new_[18742]_  = ~A265 & \new_[18741]_ ;
  assign \new_[18746]_  = A302 & A300;
  assign \new_[18747]_  = ~A299 & \new_[18746]_ ;
  assign \new_[18748]_  = \new_[18747]_  & \new_[18742]_ ;
  assign \new_[18752]_  = ~A199 & A166;
  assign \new_[18753]_  = A168 & \new_[18752]_ ;
  assign \new_[18757]_  = ~A235 & ~A233;
  assign \new_[18758]_  = ~A200 & \new_[18757]_ ;
  assign \new_[18759]_  = \new_[18758]_  & \new_[18753]_ ;
  assign \new_[18763]_  = ~A268 & ~A266;
  assign \new_[18764]_  = ~A236 & \new_[18763]_ ;
  assign \new_[18768]_  = A299 & ~A298;
  assign \new_[18769]_  = ~A269 & \new_[18768]_ ;
  assign \new_[18770]_  = \new_[18769]_  & \new_[18764]_ ;
  assign \new_[18774]_  = ~A199 & A166;
  assign \new_[18775]_  = A168 & \new_[18774]_ ;
  assign \new_[18779]_  = ~A234 & ~A233;
  assign \new_[18780]_  = ~A200 & \new_[18779]_ ;
  assign \new_[18781]_  = \new_[18780]_  & \new_[18775]_ ;
  assign \new_[18785]_  = A298 & A266;
  assign \new_[18786]_  = A265 & \new_[18785]_ ;
  assign \new_[18790]_  = A301 & A300;
  assign \new_[18791]_  = ~A299 & \new_[18790]_ ;
  assign \new_[18792]_  = \new_[18791]_  & \new_[18786]_ ;
  assign \new_[18796]_  = ~A199 & A166;
  assign \new_[18797]_  = A168 & \new_[18796]_ ;
  assign \new_[18801]_  = ~A234 & ~A233;
  assign \new_[18802]_  = ~A200 & \new_[18801]_ ;
  assign \new_[18803]_  = \new_[18802]_  & \new_[18797]_ ;
  assign \new_[18807]_  = A298 & A266;
  assign \new_[18808]_  = A265 & \new_[18807]_ ;
  assign \new_[18812]_  = A302 & A300;
  assign \new_[18813]_  = ~A299 & \new_[18812]_ ;
  assign \new_[18814]_  = \new_[18813]_  & \new_[18808]_ ;
  assign \new_[18818]_  = ~A199 & A166;
  assign \new_[18819]_  = A168 & \new_[18818]_ ;
  assign \new_[18823]_  = ~A234 & ~A233;
  assign \new_[18824]_  = ~A200 & \new_[18823]_ ;
  assign \new_[18825]_  = \new_[18824]_  & \new_[18819]_ ;
  assign \new_[18829]_  = A298 & ~A267;
  assign \new_[18830]_  = ~A266 & \new_[18829]_ ;
  assign \new_[18834]_  = A301 & A300;
  assign \new_[18835]_  = ~A299 & \new_[18834]_ ;
  assign \new_[18836]_  = \new_[18835]_  & \new_[18830]_ ;
  assign \new_[18840]_  = ~A199 & A166;
  assign \new_[18841]_  = A168 & \new_[18840]_ ;
  assign \new_[18845]_  = ~A234 & ~A233;
  assign \new_[18846]_  = ~A200 & \new_[18845]_ ;
  assign \new_[18847]_  = \new_[18846]_  & \new_[18841]_ ;
  assign \new_[18851]_  = A298 & ~A267;
  assign \new_[18852]_  = ~A266 & \new_[18851]_ ;
  assign \new_[18856]_  = A302 & A300;
  assign \new_[18857]_  = ~A299 & \new_[18856]_ ;
  assign \new_[18858]_  = \new_[18857]_  & \new_[18852]_ ;
  assign \new_[18862]_  = ~A199 & A166;
  assign \new_[18863]_  = A168 & \new_[18862]_ ;
  assign \new_[18867]_  = ~A234 & ~A233;
  assign \new_[18868]_  = ~A200 & \new_[18867]_ ;
  assign \new_[18869]_  = \new_[18868]_  & \new_[18863]_ ;
  assign \new_[18873]_  = A298 & ~A266;
  assign \new_[18874]_  = ~A265 & \new_[18873]_ ;
  assign \new_[18878]_  = A301 & A300;
  assign \new_[18879]_  = ~A299 & \new_[18878]_ ;
  assign \new_[18880]_  = \new_[18879]_  & \new_[18874]_ ;
  assign \new_[18884]_  = ~A199 & A166;
  assign \new_[18885]_  = A168 & \new_[18884]_ ;
  assign \new_[18889]_  = ~A234 & ~A233;
  assign \new_[18890]_  = ~A200 & \new_[18889]_ ;
  assign \new_[18891]_  = \new_[18890]_  & \new_[18885]_ ;
  assign \new_[18895]_  = A298 & ~A266;
  assign \new_[18896]_  = ~A265 & \new_[18895]_ ;
  assign \new_[18900]_  = A302 & A300;
  assign \new_[18901]_  = ~A299 & \new_[18900]_ ;
  assign \new_[18902]_  = \new_[18901]_  & \new_[18896]_ ;
  assign \new_[18906]_  = ~A199 & A166;
  assign \new_[18907]_  = A168 & \new_[18906]_ ;
  assign \new_[18911]_  = ~A233 & A232;
  assign \new_[18912]_  = ~A200 & \new_[18911]_ ;
  assign \new_[18913]_  = \new_[18912]_  & \new_[18907]_ ;
  assign \new_[18917]_  = A265 & A235;
  assign \new_[18918]_  = A234 & \new_[18917]_ ;
  assign \new_[18922]_  = A268 & A267;
  assign \new_[18923]_  = ~A266 & \new_[18922]_ ;
  assign \new_[18924]_  = \new_[18923]_  & \new_[18918]_ ;
  assign \new_[18928]_  = ~A199 & A166;
  assign \new_[18929]_  = A168 & \new_[18928]_ ;
  assign \new_[18933]_  = ~A233 & A232;
  assign \new_[18934]_  = ~A200 & \new_[18933]_ ;
  assign \new_[18935]_  = \new_[18934]_  & \new_[18929]_ ;
  assign \new_[18939]_  = A265 & A235;
  assign \new_[18940]_  = A234 & \new_[18939]_ ;
  assign \new_[18944]_  = A269 & A267;
  assign \new_[18945]_  = ~A266 & \new_[18944]_ ;
  assign \new_[18946]_  = \new_[18945]_  & \new_[18940]_ ;
  assign \new_[18950]_  = ~A199 & A166;
  assign \new_[18951]_  = A168 & \new_[18950]_ ;
  assign \new_[18955]_  = ~A233 & A232;
  assign \new_[18956]_  = ~A200 & \new_[18955]_ ;
  assign \new_[18957]_  = \new_[18956]_  & \new_[18951]_ ;
  assign \new_[18961]_  = A265 & A236;
  assign \new_[18962]_  = A234 & \new_[18961]_ ;
  assign \new_[18966]_  = A268 & A267;
  assign \new_[18967]_  = ~A266 & \new_[18966]_ ;
  assign \new_[18968]_  = \new_[18967]_  & \new_[18962]_ ;
  assign \new_[18972]_  = ~A199 & A166;
  assign \new_[18973]_  = A168 & \new_[18972]_ ;
  assign \new_[18977]_  = ~A233 & A232;
  assign \new_[18978]_  = ~A200 & \new_[18977]_ ;
  assign \new_[18979]_  = \new_[18978]_  & \new_[18973]_ ;
  assign \new_[18983]_  = A265 & A236;
  assign \new_[18984]_  = A234 & \new_[18983]_ ;
  assign \new_[18988]_  = A269 & A267;
  assign \new_[18989]_  = ~A266 & \new_[18988]_ ;
  assign \new_[18990]_  = \new_[18989]_  & \new_[18984]_ ;
  assign \new_[18994]_  = ~A199 & A166;
  assign \new_[18995]_  = A168 & \new_[18994]_ ;
  assign \new_[18999]_  = ~A233 & ~A232;
  assign \new_[19000]_  = ~A200 & \new_[18999]_ ;
  assign \new_[19001]_  = \new_[19000]_  & \new_[18995]_ ;
  assign \new_[19005]_  = A298 & A266;
  assign \new_[19006]_  = A265 & \new_[19005]_ ;
  assign \new_[19010]_  = A301 & A300;
  assign \new_[19011]_  = ~A299 & \new_[19010]_ ;
  assign \new_[19012]_  = \new_[19011]_  & \new_[19006]_ ;
  assign \new_[19016]_  = ~A199 & A166;
  assign \new_[19017]_  = A168 & \new_[19016]_ ;
  assign \new_[19021]_  = ~A233 & ~A232;
  assign \new_[19022]_  = ~A200 & \new_[19021]_ ;
  assign \new_[19023]_  = \new_[19022]_  & \new_[19017]_ ;
  assign \new_[19027]_  = A298 & A266;
  assign \new_[19028]_  = A265 & \new_[19027]_ ;
  assign \new_[19032]_  = A302 & A300;
  assign \new_[19033]_  = ~A299 & \new_[19032]_ ;
  assign \new_[19034]_  = \new_[19033]_  & \new_[19028]_ ;
  assign \new_[19038]_  = ~A199 & A166;
  assign \new_[19039]_  = A168 & \new_[19038]_ ;
  assign \new_[19043]_  = ~A233 & ~A232;
  assign \new_[19044]_  = ~A200 & \new_[19043]_ ;
  assign \new_[19045]_  = \new_[19044]_  & \new_[19039]_ ;
  assign \new_[19049]_  = A298 & ~A267;
  assign \new_[19050]_  = ~A266 & \new_[19049]_ ;
  assign \new_[19054]_  = A301 & A300;
  assign \new_[19055]_  = ~A299 & \new_[19054]_ ;
  assign \new_[19056]_  = \new_[19055]_  & \new_[19050]_ ;
  assign \new_[19060]_  = ~A199 & A166;
  assign \new_[19061]_  = A168 & \new_[19060]_ ;
  assign \new_[19065]_  = ~A233 & ~A232;
  assign \new_[19066]_  = ~A200 & \new_[19065]_ ;
  assign \new_[19067]_  = \new_[19066]_  & \new_[19061]_ ;
  assign \new_[19071]_  = A298 & ~A267;
  assign \new_[19072]_  = ~A266 & \new_[19071]_ ;
  assign \new_[19076]_  = A302 & A300;
  assign \new_[19077]_  = ~A299 & \new_[19076]_ ;
  assign \new_[19078]_  = \new_[19077]_  & \new_[19072]_ ;
  assign \new_[19082]_  = ~A199 & A166;
  assign \new_[19083]_  = A168 & \new_[19082]_ ;
  assign \new_[19087]_  = ~A233 & ~A232;
  assign \new_[19088]_  = ~A200 & \new_[19087]_ ;
  assign \new_[19089]_  = \new_[19088]_  & \new_[19083]_ ;
  assign \new_[19093]_  = A298 & ~A266;
  assign \new_[19094]_  = ~A265 & \new_[19093]_ ;
  assign \new_[19098]_  = A301 & A300;
  assign \new_[19099]_  = ~A299 & \new_[19098]_ ;
  assign \new_[19100]_  = \new_[19099]_  & \new_[19094]_ ;
  assign \new_[19104]_  = ~A199 & A166;
  assign \new_[19105]_  = A168 & \new_[19104]_ ;
  assign \new_[19109]_  = ~A233 & ~A232;
  assign \new_[19110]_  = ~A200 & \new_[19109]_ ;
  assign \new_[19111]_  = \new_[19110]_  & \new_[19105]_ ;
  assign \new_[19115]_  = A298 & ~A266;
  assign \new_[19116]_  = ~A265 & \new_[19115]_ ;
  assign \new_[19120]_  = A302 & A300;
  assign \new_[19121]_  = ~A299 & \new_[19120]_ ;
  assign \new_[19122]_  = \new_[19121]_  & \new_[19116]_ ;
  assign \new_[19126]_  = A199 & A167;
  assign \new_[19127]_  = A168 & \new_[19126]_ ;
  assign \new_[19131]_  = A233 & A232;
  assign \new_[19132]_  = A200 & \new_[19131]_ ;
  assign \new_[19133]_  = \new_[19132]_  & \new_[19127]_ ;
  assign \new_[19137]_  = A298 & ~A267;
  assign \new_[19138]_  = A265 & \new_[19137]_ ;
  assign \new_[19142]_  = A301 & A300;
  assign \new_[19143]_  = ~A299 & \new_[19142]_ ;
  assign \new_[19144]_  = \new_[19143]_  & \new_[19138]_ ;
  assign \new_[19148]_  = A199 & A167;
  assign \new_[19149]_  = A168 & \new_[19148]_ ;
  assign \new_[19153]_  = A233 & A232;
  assign \new_[19154]_  = A200 & \new_[19153]_ ;
  assign \new_[19155]_  = \new_[19154]_  & \new_[19149]_ ;
  assign \new_[19159]_  = A298 & ~A267;
  assign \new_[19160]_  = A265 & \new_[19159]_ ;
  assign \new_[19164]_  = A302 & A300;
  assign \new_[19165]_  = ~A299 & \new_[19164]_ ;
  assign \new_[19166]_  = \new_[19165]_  & \new_[19160]_ ;
  assign \new_[19170]_  = A199 & A167;
  assign \new_[19171]_  = A168 & \new_[19170]_ ;
  assign \new_[19175]_  = A233 & A232;
  assign \new_[19176]_  = A200 & \new_[19175]_ ;
  assign \new_[19177]_  = \new_[19176]_  & \new_[19171]_ ;
  assign \new_[19181]_  = A298 & A266;
  assign \new_[19182]_  = A265 & \new_[19181]_ ;
  assign \new_[19186]_  = A301 & A300;
  assign \new_[19187]_  = ~A299 & \new_[19186]_ ;
  assign \new_[19188]_  = \new_[19187]_  & \new_[19182]_ ;
  assign \new_[19192]_  = A199 & A167;
  assign \new_[19193]_  = A168 & \new_[19192]_ ;
  assign \new_[19197]_  = A233 & A232;
  assign \new_[19198]_  = A200 & \new_[19197]_ ;
  assign \new_[19199]_  = \new_[19198]_  & \new_[19193]_ ;
  assign \new_[19203]_  = A298 & A266;
  assign \new_[19204]_  = A265 & \new_[19203]_ ;
  assign \new_[19208]_  = A302 & A300;
  assign \new_[19209]_  = ~A299 & \new_[19208]_ ;
  assign \new_[19210]_  = \new_[19209]_  & \new_[19204]_ ;
  assign \new_[19214]_  = A199 & A167;
  assign \new_[19215]_  = A168 & \new_[19214]_ ;
  assign \new_[19219]_  = A233 & A232;
  assign \new_[19220]_  = A200 & \new_[19219]_ ;
  assign \new_[19221]_  = \new_[19220]_  & \new_[19215]_ ;
  assign \new_[19225]_  = A298 & ~A266;
  assign \new_[19226]_  = ~A265 & \new_[19225]_ ;
  assign \new_[19230]_  = A301 & A300;
  assign \new_[19231]_  = ~A299 & \new_[19230]_ ;
  assign \new_[19232]_  = \new_[19231]_  & \new_[19226]_ ;
  assign \new_[19236]_  = A199 & A167;
  assign \new_[19237]_  = A168 & \new_[19236]_ ;
  assign \new_[19241]_  = A233 & A232;
  assign \new_[19242]_  = A200 & \new_[19241]_ ;
  assign \new_[19243]_  = \new_[19242]_  & \new_[19237]_ ;
  assign \new_[19247]_  = A298 & ~A266;
  assign \new_[19248]_  = ~A265 & \new_[19247]_ ;
  assign \new_[19252]_  = A302 & A300;
  assign \new_[19253]_  = ~A299 & \new_[19252]_ ;
  assign \new_[19254]_  = \new_[19253]_  & \new_[19248]_ ;
  assign \new_[19258]_  = A199 & A167;
  assign \new_[19259]_  = A168 & \new_[19258]_ ;
  assign \new_[19263]_  = ~A235 & ~A233;
  assign \new_[19264]_  = A200 & \new_[19263]_ ;
  assign \new_[19265]_  = \new_[19264]_  & \new_[19259]_ ;
  assign \new_[19269]_  = ~A268 & ~A266;
  assign \new_[19270]_  = ~A236 & \new_[19269]_ ;
  assign \new_[19274]_  = A299 & ~A298;
  assign \new_[19275]_  = ~A269 & \new_[19274]_ ;
  assign \new_[19276]_  = \new_[19275]_  & \new_[19270]_ ;
  assign \new_[19280]_  = A199 & A167;
  assign \new_[19281]_  = A168 & \new_[19280]_ ;
  assign \new_[19285]_  = ~A234 & ~A233;
  assign \new_[19286]_  = A200 & \new_[19285]_ ;
  assign \new_[19287]_  = \new_[19286]_  & \new_[19281]_ ;
  assign \new_[19291]_  = A298 & A266;
  assign \new_[19292]_  = A265 & \new_[19291]_ ;
  assign \new_[19296]_  = A301 & A300;
  assign \new_[19297]_  = ~A299 & \new_[19296]_ ;
  assign \new_[19298]_  = \new_[19297]_  & \new_[19292]_ ;
  assign \new_[19302]_  = A199 & A167;
  assign \new_[19303]_  = A168 & \new_[19302]_ ;
  assign \new_[19307]_  = ~A234 & ~A233;
  assign \new_[19308]_  = A200 & \new_[19307]_ ;
  assign \new_[19309]_  = \new_[19308]_  & \new_[19303]_ ;
  assign \new_[19313]_  = A298 & A266;
  assign \new_[19314]_  = A265 & \new_[19313]_ ;
  assign \new_[19318]_  = A302 & A300;
  assign \new_[19319]_  = ~A299 & \new_[19318]_ ;
  assign \new_[19320]_  = \new_[19319]_  & \new_[19314]_ ;
  assign \new_[19324]_  = A199 & A167;
  assign \new_[19325]_  = A168 & \new_[19324]_ ;
  assign \new_[19329]_  = ~A234 & ~A233;
  assign \new_[19330]_  = A200 & \new_[19329]_ ;
  assign \new_[19331]_  = \new_[19330]_  & \new_[19325]_ ;
  assign \new_[19335]_  = A298 & ~A267;
  assign \new_[19336]_  = ~A266 & \new_[19335]_ ;
  assign \new_[19340]_  = A301 & A300;
  assign \new_[19341]_  = ~A299 & \new_[19340]_ ;
  assign \new_[19342]_  = \new_[19341]_  & \new_[19336]_ ;
  assign \new_[19346]_  = A199 & A167;
  assign \new_[19347]_  = A168 & \new_[19346]_ ;
  assign \new_[19351]_  = ~A234 & ~A233;
  assign \new_[19352]_  = A200 & \new_[19351]_ ;
  assign \new_[19353]_  = \new_[19352]_  & \new_[19347]_ ;
  assign \new_[19357]_  = A298 & ~A267;
  assign \new_[19358]_  = ~A266 & \new_[19357]_ ;
  assign \new_[19362]_  = A302 & A300;
  assign \new_[19363]_  = ~A299 & \new_[19362]_ ;
  assign \new_[19364]_  = \new_[19363]_  & \new_[19358]_ ;
  assign \new_[19368]_  = A199 & A167;
  assign \new_[19369]_  = A168 & \new_[19368]_ ;
  assign \new_[19373]_  = ~A234 & ~A233;
  assign \new_[19374]_  = A200 & \new_[19373]_ ;
  assign \new_[19375]_  = \new_[19374]_  & \new_[19369]_ ;
  assign \new_[19379]_  = A298 & ~A266;
  assign \new_[19380]_  = ~A265 & \new_[19379]_ ;
  assign \new_[19384]_  = A301 & A300;
  assign \new_[19385]_  = ~A299 & \new_[19384]_ ;
  assign \new_[19386]_  = \new_[19385]_  & \new_[19380]_ ;
  assign \new_[19390]_  = A199 & A167;
  assign \new_[19391]_  = A168 & \new_[19390]_ ;
  assign \new_[19395]_  = ~A234 & ~A233;
  assign \new_[19396]_  = A200 & \new_[19395]_ ;
  assign \new_[19397]_  = \new_[19396]_  & \new_[19391]_ ;
  assign \new_[19401]_  = A298 & ~A266;
  assign \new_[19402]_  = ~A265 & \new_[19401]_ ;
  assign \new_[19406]_  = A302 & A300;
  assign \new_[19407]_  = ~A299 & \new_[19406]_ ;
  assign \new_[19408]_  = \new_[19407]_  & \new_[19402]_ ;
  assign \new_[19412]_  = A199 & A167;
  assign \new_[19413]_  = A168 & \new_[19412]_ ;
  assign \new_[19417]_  = ~A233 & A232;
  assign \new_[19418]_  = A200 & \new_[19417]_ ;
  assign \new_[19419]_  = \new_[19418]_  & \new_[19413]_ ;
  assign \new_[19423]_  = A265 & A235;
  assign \new_[19424]_  = A234 & \new_[19423]_ ;
  assign \new_[19428]_  = A268 & A267;
  assign \new_[19429]_  = ~A266 & \new_[19428]_ ;
  assign \new_[19430]_  = \new_[19429]_  & \new_[19424]_ ;
  assign \new_[19434]_  = A199 & A167;
  assign \new_[19435]_  = A168 & \new_[19434]_ ;
  assign \new_[19439]_  = ~A233 & A232;
  assign \new_[19440]_  = A200 & \new_[19439]_ ;
  assign \new_[19441]_  = \new_[19440]_  & \new_[19435]_ ;
  assign \new_[19445]_  = A265 & A235;
  assign \new_[19446]_  = A234 & \new_[19445]_ ;
  assign \new_[19450]_  = A269 & A267;
  assign \new_[19451]_  = ~A266 & \new_[19450]_ ;
  assign \new_[19452]_  = \new_[19451]_  & \new_[19446]_ ;
  assign \new_[19456]_  = A199 & A167;
  assign \new_[19457]_  = A168 & \new_[19456]_ ;
  assign \new_[19461]_  = ~A233 & A232;
  assign \new_[19462]_  = A200 & \new_[19461]_ ;
  assign \new_[19463]_  = \new_[19462]_  & \new_[19457]_ ;
  assign \new_[19467]_  = A265 & A236;
  assign \new_[19468]_  = A234 & \new_[19467]_ ;
  assign \new_[19472]_  = A268 & A267;
  assign \new_[19473]_  = ~A266 & \new_[19472]_ ;
  assign \new_[19474]_  = \new_[19473]_  & \new_[19468]_ ;
  assign \new_[19478]_  = A199 & A167;
  assign \new_[19479]_  = A168 & \new_[19478]_ ;
  assign \new_[19483]_  = ~A233 & A232;
  assign \new_[19484]_  = A200 & \new_[19483]_ ;
  assign \new_[19485]_  = \new_[19484]_  & \new_[19479]_ ;
  assign \new_[19489]_  = A265 & A236;
  assign \new_[19490]_  = A234 & \new_[19489]_ ;
  assign \new_[19494]_  = A269 & A267;
  assign \new_[19495]_  = ~A266 & \new_[19494]_ ;
  assign \new_[19496]_  = \new_[19495]_  & \new_[19490]_ ;
  assign \new_[19500]_  = A199 & A167;
  assign \new_[19501]_  = A168 & \new_[19500]_ ;
  assign \new_[19505]_  = ~A233 & ~A232;
  assign \new_[19506]_  = A200 & \new_[19505]_ ;
  assign \new_[19507]_  = \new_[19506]_  & \new_[19501]_ ;
  assign \new_[19511]_  = A298 & A266;
  assign \new_[19512]_  = A265 & \new_[19511]_ ;
  assign \new_[19516]_  = A301 & A300;
  assign \new_[19517]_  = ~A299 & \new_[19516]_ ;
  assign \new_[19518]_  = \new_[19517]_  & \new_[19512]_ ;
  assign \new_[19522]_  = A199 & A167;
  assign \new_[19523]_  = A168 & \new_[19522]_ ;
  assign \new_[19527]_  = ~A233 & ~A232;
  assign \new_[19528]_  = A200 & \new_[19527]_ ;
  assign \new_[19529]_  = \new_[19528]_  & \new_[19523]_ ;
  assign \new_[19533]_  = A298 & A266;
  assign \new_[19534]_  = A265 & \new_[19533]_ ;
  assign \new_[19538]_  = A302 & A300;
  assign \new_[19539]_  = ~A299 & \new_[19538]_ ;
  assign \new_[19540]_  = \new_[19539]_  & \new_[19534]_ ;
  assign \new_[19544]_  = A199 & A167;
  assign \new_[19545]_  = A168 & \new_[19544]_ ;
  assign \new_[19549]_  = ~A233 & ~A232;
  assign \new_[19550]_  = A200 & \new_[19549]_ ;
  assign \new_[19551]_  = \new_[19550]_  & \new_[19545]_ ;
  assign \new_[19555]_  = A298 & ~A267;
  assign \new_[19556]_  = ~A266 & \new_[19555]_ ;
  assign \new_[19560]_  = A301 & A300;
  assign \new_[19561]_  = ~A299 & \new_[19560]_ ;
  assign \new_[19562]_  = \new_[19561]_  & \new_[19556]_ ;
  assign \new_[19566]_  = A199 & A167;
  assign \new_[19567]_  = A168 & \new_[19566]_ ;
  assign \new_[19571]_  = ~A233 & ~A232;
  assign \new_[19572]_  = A200 & \new_[19571]_ ;
  assign \new_[19573]_  = \new_[19572]_  & \new_[19567]_ ;
  assign \new_[19577]_  = A298 & ~A267;
  assign \new_[19578]_  = ~A266 & \new_[19577]_ ;
  assign \new_[19582]_  = A302 & A300;
  assign \new_[19583]_  = ~A299 & \new_[19582]_ ;
  assign \new_[19584]_  = \new_[19583]_  & \new_[19578]_ ;
  assign \new_[19588]_  = A199 & A167;
  assign \new_[19589]_  = A168 & \new_[19588]_ ;
  assign \new_[19593]_  = ~A233 & ~A232;
  assign \new_[19594]_  = A200 & \new_[19593]_ ;
  assign \new_[19595]_  = \new_[19594]_  & \new_[19589]_ ;
  assign \new_[19599]_  = A298 & ~A266;
  assign \new_[19600]_  = ~A265 & \new_[19599]_ ;
  assign \new_[19604]_  = A301 & A300;
  assign \new_[19605]_  = ~A299 & \new_[19604]_ ;
  assign \new_[19606]_  = \new_[19605]_  & \new_[19600]_ ;
  assign \new_[19610]_  = A199 & A167;
  assign \new_[19611]_  = A168 & \new_[19610]_ ;
  assign \new_[19615]_  = ~A233 & ~A232;
  assign \new_[19616]_  = A200 & \new_[19615]_ ;
  assign \new_[19617]_  = \new_[19616]_  & \new_[19611]_ ;
  assign \new_[19621]_  = A298 & ~A266;
  assign \new_[19622]_  = ~A265 & \new_[19621]_ ;
  assign \new_[19626]_  = A302 & A300;
  assign \new_[19627]_  = ~A299 & \new_[19626]_ ;
  assign \new_[19628]_  = \new_[19627]_  & \new_[19622]_ ;
  assign \new_[19632]_  = ~A200 & A167;
  assign \new_[19633]_  = A168 & \new_[19632]_ ;
  assign \new_[19637]_  = A232 & ~A203;
  assign \new_[19638]_  = ~A202 & \new_[19637]_ ;
  assign \new_[19639]_  = \new_[19638]_  & \new_[19633]_ ;
  assign \new_[19643]_  = ~A268 & A265;
  assign \new_[19644]_  = A233 & \new_[19643]_ ;
  assign \new_[19648]_  = A299 & ~A298;
  assign \new_[19649]_  = ~A269 & \new_[19648]_ ;
  assign \new_[19650]_  = \new_[19649]_  & \new_[19644]_ ;
  assign \new_[19654]_  = ~A200 & A167;
  assign \new_[19655]_  = A168 & \new_[19654]_ ;
  assign \new_[19659]_  = ~A233 & ~A203;
  assign \new_[19660]_  = ~A202 & \new_[19659]_ ;
  assign \new_[19661]_  = \new_[19660]_  & \new_[19655]_ ;
  assign \new_[19665]_  = A265 & ~A236;
  assign \new_[19666]_  = ~A235 & \new_[19665]_ ;
  assign \new_[19670]_  = A299 & ~A298;
  assign \new_[19671]_  = A266 & \new_[19670]_ ;
  assign \new_[19672]_  = \new_[19671]_  & \new_[19666]_ ;
  assign \new_[19676]_  = ~A200 & A167;
  assign \new_[19677]_  = A168 & \new_[19676]_ ;
  assign \new_[19681]_  = ~A233 & ~A203;
  assign \new_[19682]_  = ~A202 & \new_[19681]_ ;
  assign \new_[19683]_  = \new_[19682]_  & \new_[19677]_ ;
  assign \new_[19687]_  = ~A266 & ~A236;
  assign \new_[19688]_  = ~A235 & \new_[19687]_ ;
  assign \new_[19692]_  = A299 & ~A298;
  assign \new_[19693]_  = ~A267 & \new_[19692]_ ;
  assign \new_[19694]_  = \new_[19693]_  & \new_[19688]_ ;
  assign \new_[19698]_  = ~A200 & A167;
  assign \new_[19699]_  = A168 & \new_[19698]_ ;
  assign \new_[19703]_  = ~A233 & ~A203;
  assign \new_[19704]_  = ~A202 & \new_[19703]_ ;
  assign \new_[19705]_  = \new_[19704]_  & \new_[19699]_ ;
  assign \new_[19709]_  = ~A265 & ~A236;
  assign \new_[19710]_  = ~A235 & \new_[19709]_ ;
  assign \new_[19714]_  = A299 & ~A298;
  assign \new_[19715]_  = ~A266 & \new_[19714]_ ;
  assign \new_[19716]_  = \new_[19715]_  & \new_[19710]_ ;
  assign \new_[19720]_  = ~A200 & A167;
  assign \new_[19721]_  = A168 & \new_[19720]_ ;
  assign \new_[19725]_  = ~A233 & ~A203;
  assign \new_[19726]_  = ~A202 & \new_[19725]_ ;
  assign \new_[19727]_  = \new_[19726]_  & \new_[19721]_ ;
  assign \new_[19731]_  = ~A268 & ~A266;
  assign \new_[19732]_  = ~A234 & \new_[19731]_ ;
  assign \new_[19736]_  = A299 & ~A298;
  assign \new_[19737]_  = ~A269 & \new_[19736]_ ;
  assign \new_[19738]_  = \new_[19737]_  & \new_[19732]_ ;
  assign \new_[19742]_  = ~A200 & A167;
  assign \new_[19743]_  = A168 & \new_[19742]_ ;
  assign \new_[19747]_  = A232 & ~A203;
  assign \new_[19748]_  = ~A202 & \new_[19747]_ ;
  assign \new_[19749]_  = \new_[19748]_  & \new_[19743]_ ;
  assign \new_[19753]_  = A235 & A234;
  assign \new_[19754]_  = ~A233 & \new_[19753]_ ;
  assign \new_[19758]_  = ~A302 & ~A301;
  assign \new_[19759]_  = A298 & \new_[19758]_ ;
  assign \new_[19760]_  = \new_[19759]_  & \new_[19754]_ ;
  assign \new_[19764]_  = ~A200 & A167;
  assign \new_[19765]_  = A168 & \new_[19764]_ ;
  assign \new_[19769]_  = A232 & ~A203;
  assign \new_[19770]_  = ~A202 & \new_[19769]_ ;
  assign \new_[19771]_  = \new_[19770]_  & \new_[19765]_ ;
  assign \new_[19775]_  = A236 & A234;
  assign \new_[19776]_  = ~A233 & \new_[19775]_ ;
  assign \new_[19780]_  = ~A302 & ~A301;
  assign \new_[19781]_  = A298 & \new_[19780]_ ;
  assign \new_[19782]_  = \new_[19781]_  & \new_[19776]_ ;
  assign \new_[19786]_  = ~A200 & A167;
  assign \new_[19787]_  = A168 & \new_[19786]_ ;
  assign \new_[19791]_  = ~A232 & ~A203;
  assign \new_[19792]_  = ~A202 & \new_[19791]_ ;
  assign \new_[19793]_  = \new_[19792]_  & \new_[19787]_ ;
  assign \new_[19797]_  = ~A268 & ~A266;
  assign \new_[19798]_  = ~A233 & \new_[19797]_ ;
  assign \new_[19802]_  = A299 & ~A298;
  assign \new_[19803]_  = ~A269 & \new_[19802]_ ;
  assign \new_[19804]_  = \new_[19803]_  & \new_[19798]_ ;
  assign \new_[19808]_  = ~A200 & A167;
  assign \new_[19809]_  = A168 & \new_[19808]_ ;
  assign \new_[19813]_  = A233 & A232;
  assign \new_[19814]_  = ~A201 & \new_[19813]_ ;
  assign \new_[19815]_  = \new_[19814]_  & \new_[19809]_ ;
  assign \new_[19819]_  = A298 & ~A267;
  assign \new_[19820]_  = A265 & \new_[19819]_ ;
  assign \new_[19824]_  = A301 & A300;
  assign \new_[19825]_  = ~A299 & \new_[19824]_ ;
  assign \new_[19826]_  = \new_[19825]_  & \new_[19820]_ ;
  assign \new_[19830]_  = ~A200 & A167;
  assign \new_[19831]_  = A168 & \new_[19830]_ ;
  assign \new_[19835]_  = A233 & A232;
  assign \new_[19836]_  = ~A201 & \new_[19835]_ ;
  assign \new_[19837]_  = \new_[19836]_  & \new_[19831]_ ;
  assign \new_[19841]_  = A298 & ~A267;
  assign \new_[19842]_  = A265 & \new_[19841]_ ;
  assign \new_[19846]_  = A302 & A300;
  assign \new_[19847]_  = ~A299 & \new_[19846]_ ;
  assign \new_[19848]_  = \new_[19847]_  & \new_[19842]_ ;
  assign \new_[19852]_  = ~A200 & A167;
  assign \new_[19853]_  = A168 & \new_[19852]_ ;
  assign \new_[19857]_  = A233 & A232;
  assign \new_[19858]_  = ~A201 & \new_[19857]_ ;
  assign \new_[19859]_  = \new_[19858]_  & \new_[19853]_ ;
  assign \new_[19863]_  = A298 & A266;
  assign \new_[19864]_  = A265 & \new_[19863]_ ;
  assign \new_[19868]_  = A301 & A300;
  assign \new_[19869]_  = ~A299 & \new_[19868]_ ;
  assign \new_[19870]_  = \new_[19869]_  & \new_[19864]_ ;
  assign \new_[19874]_  = ~A200 & A167;
  assign \new_[19875]_  = A168 & \new_[19874]_ ;
  assign \new_[19879]_  = A233 & A232;
  assign \new_[19880]_  = ~A201 & \new_[19879]_ ;
  assign \new_[19881]_  = \new_[19880]_  & \new_[19875]_ ;
  assign \new_[19885]_  = A298 & A266;
  assign \new_[19886]_  = A265 & \new_[19885]_ ;
  assign \new_[19890]_  = A302 & A300;
  assign \new_[19891]_  = ~A299 & \new_[19890]_ ;
  assign \new_[19892]_  = \new_[19891]_  & \new_[19886]_ ;
  assign \new_[19896]_  = ~A200 & A167;
  assign \new_[19897]_  = A168 & \new_[19896]_ ;
  assign \new_[19901]_  = A233 & A232;
  assign \new_[19902]_  = ~A201 & \new_[19901]_ ;
  assign \new_[19903]_  = \new_[19902]_  & \new_[19897]_ ;
  assign \new_[19907]_  = A298 & ~A266;
  assign \new_[19908]_  = ~A265 & \new_[19907]_ ;
  assign \new_[19912]_  = A301 & A300;
  assign \new_[19913]_  = ~A299 & \new_[19912]_ ;
  assign \new_[19914]_  = \new_[19913]_  & \new_[19908]_ ;
  assign \new_[19918]_  = ~A200 & A167;
  assign \new_[19919]_  = A168 & \new_[19918]_ ;
  assign \new_[19923]_  = A233 & A232;
  assign \new_[19924]_  = ~A201 & \new_[19923]_ ;
  assign \new_[19925]_  = \new_[19924]_  & \new_[19919]_ ;
  assign \new_[19929]_  = A298 & ~A266;
  assign \new_[19930]_  = ~A265 & \new_[19929]_ ;
  assign \new_[19934]_  = A302 & A300;
  assign \new_[19935]_  = ~A299 & \new_[19934]_ ;
  assign \new_[19936]_  = \new_[19935]_  & \new_[19930]_ ;
  assign \new_[19940]_  = ~A200 & A167;
  assign \new_[19941]_  = A168 & \new_[19940]_ ;
  assign \new_[19945]_  = ~A235 & ~A233;
  assign \new_[19946]_  = ~A201 & \new_[19945]_ ;
  assign \new_[19947]_  = \new_[19946]_  & \new_[19941]_ ;
  assign \new_[19951]_  = ~A268 & ~A266;
  assign \new_[19952]_  = ~A236 & \new_[19951]_ ;
  assign \new_[19956]_  = A299 & ~A298;
  assign \new_[19957]_  = ~A269 & \new_[19956]_ ;
  assign \new_[19958]_  = \new_[19957]_  & \new_[19952]_ ;
  assign \new_[19962]_  = ~A200 & A167;
  assign \new_[19963]_  = A168 & \new_[19962]_ ;
  assign \new_[19967]_  = ~A234 & ~A233;
  assign \new_[19968]_  = ~A201 & \new_[19967]_ ;
  assign \new_[19969]_  = \new_[19968]_  & \new_[19963]_ ;
  assign \new_[19973]_  = A298 & A266;
  assign \new_[19974]_  = A265 & \new_[19973]_ ;
  assign \new_[19978]_  = A301 & A300;
  assign \new_[19979]_  = ~A299 & \new_[19978]_ ;
  assign \new_[19980]_  = \new_[19979]_  & \new_[19974]_ ;
  assign \new_[19984]_  = ~A200 & A167;
  assign \new_[19985]_  = A168 & \new_[19984]_ ;
  assign \new_[19989]_  = ~A234 & ~A233;
  assign \new_[19990]_  = ~A201 & \new_[19989]_ ;
  assign \new_[19991]_  = \new_[19990]_  & \new_[19985]_ ;
  assign \new_[19995]_  = A298 & A266;
  assign \new_[19996]_  = A265 & \new_[19995]_ ;
  assign \new_[20000]_  = A302 & A300;
  assign \new_[20001]_  = ~A299 & \new_[20000]_ ;
  assign \new_[20002]_  = \new_[20001]_  & \new_[19996]_ ;
  assign \new_[20006]_  = ~A200 & A167;
  assign \new_[20007]_  = A168 & \new_[20006]_ ;
  assign \new_[20011]_  = ~A234 & ~A233;
  assign \new_[20012]_  = ~A201 & \new_[20011]_ ;
  assign \new_[20013]_  = \new_[20012]_  & \new_[20007]_ ;
  assign \new_[20017]_  = A298 & ~A267;
  assign \new_[20018]_  = ~A266 & \new_[20017]_ ;
  assign \new_[20022]_  = A301 & A300;
  assign \new_[20023]_  = ~A299 & \new_[20022]_ ;
  assign \new_[20024]_  = \new_[20023]_  & \new_[20018]_ ;
  assign \new_[20028]_  = ~A200 & A167;
  assign \new_[20029]_  = A168 & \new_[20028]_ ;
  assign \new_[20033]_  = ~A234 & ~A233;
  assign \new_[20034]_  = ~A201 & \new_[20033]_ ;
  assign \new_[20035]_  = \new_[20034]_  & \new_[20029]_ ;
  assign \new_[20039]_  = A298 & ~A267;
  assign \new_[20040]_  = ~A266 & \new_[20039]_ ;
  assign \new_[20044]_  = A302 & A300;
  assign \new_[20045]_  = ~A299 & \new_[20044]_ ;
  assign \new_[20046]_  = \new_[20045]_  & \new_[20040]_ ;
  assign \new_[20050]_  = ~A200 & A167;
  assign \new_[20051]_  = A168 & \new_[20050]_ ;
  assign \new_[20055]_  = ~A234 & ~A233;
  assign \new_[20056]_  = ~A201 & \new_[20055]_ ;
  assign \new_[20057]_  = \new_[20056]_  & \new_[20051]_ ;
  assign \new_[20061]_  = A298 & ~A266;
  assign \new_[20062]_  = ~A265 & \new_[20061]_ ;
  assign \new_[20066]_  = A301 & A300;
  assign \new_[20067]_  = ~A299 & \new_[20066]_ ;
  assign \new_[20068]_  = \new_[20067]_  & \new_[20062]_ ;
  assign \new_[20072]_  = ~A200 & A167;
  assign \new_[20073]_  = A168 & \new_[20072]_ ;
  assign \new_[20077]_  = ~A234 & ~A233;
  assign \new_[20078]_  = ~A201 & \new_[20077]_ ;
  assign \new_[20079]_  = \new_[20078]_  & \new_[20073]_ ;
  assign \new_[20083]_  = A298 & ~A266;
  assign \new_[20084]_  = ~A265 & \new_[20083]_ ;
  assign \new_[20088]_  = A302 & A300;
  assign \new_[20089]_  = ~A299 & \new_[20088]_ ;
  assign \new_[20090]_  = \new_[20089]_  & \new_[20084]_ ;
  assign \new_[20094]_  = ~A200 & A167;
  assign \new_[20095]_  = A168 & \new_[20094]_ ;
  assign \new_[20099]_  = ~A233 & A232;
  assign \new_[20100]_  = ~A201 & \new_[20099]_ ;
  assign \new_[20101]_  = \new_[20100]_  & \new_[20095]_ ;
  assign \new_[20105]_  = A265 & A235;
  assign \new_[20106]_  = A234 & \new_[20105]_ ;
  assign \new_[20110]_  = A268 & A267;
  assign \new_[20111]_  = ~A266 & \new_[20110]_ ;
  assign \new_[20112]_  = \new_[20111]_  & \new_[20106]_ ;
  assign \new_[20116]_  = ~A200 & A167;
  assign \new_[20117]_  = A168 & \new_[20116]_ ;
  assign \new_[20121]_  = ~A233 & A232;
  assign \new_[20122]_  = ~A201 & \new_[20121]_ ;
  assign \new_[20123]_  = \new_[20122]_  & \new_[20117]_ ;
  assign \new_[20127]_  = A265 & A235;
  assign \new_[20128]_  = A234 & \new_[20127]_ ;
  assign \new_[20132]_  = A269 & A267;
  assign \new_[20133]_  = ~A266 & \new_[20132]_ ;
  assign \new_[20134]_  = \new_[20133]_  & \new_[20128]_ ;
  assign \new_[20138]_  = ~A200 & A167;
  assign \new_[20139]_  = A168 & \new_[20138]_ ;
  assign \new_[20143]_  = ~A233 & A232;
  assign \new_[20144]_  = ~A201 & \new_[20143]_ ;
  assign \new_[20145]_  = \new_[20144]_  & \new_[20139]_ ;
  assign \new_[20149]_  = A265 & A236;
  assign \new_[20150]_  = A234 & \new_[20149]_ ;
  assign \new_[20154]_  = A268 & A267;
  assign \new_[20155]_  = ~A266 & \new_[20154]_ ;
  assign \new_[20156]_  = \new_[20155]_  & \new_[20150]_ ;
  assign \new_[20160]_  = ~A200 & A167;
  assign \new_[20161]_  = A168 & \new_[20160]_ ;
  assign \new_[20165]_  = ~A233 & A232;
  assign \new_[20166]_  = ~A201 & \new_[20165]_ ;
  assign \new_[20167]_  = \new_[20166]_  & \new_[20161]_ ;
  assign \new_[20171]_  = A265 & A236;
  assign \new_[20172]_  = A234 & \new_[20171]_ ;
  assign \new_[20176]_  = A269 & A267;
  assign \new_[20177]_  = ~A266 & \new_[20176]_ ;
  assign \new_[20178]_  = \new_[20177]_  & \new_[20172]_ ;
  assign \new_[20182]_  = ~A200 & A167;
  assign \new_[20183]_  = A168 & \new_[20182]_ ;
  assign \new_[20187]_  = ~A233 & ~A232;
  assign \new_[20188]_  = ~A201 & \new_[20187]_ ;
  assign \new_[20189]_  = \new_[20188]_  & \new_[20183]_ ;
  assign \new_[20193]_  = A298 & A266;
  assign \new_[20194]_  = A265 & \new_[20193]_ ;
  assign \new_[20198]_  = A301 & A300;
  assign \new_[20199]_  = ~A299 & \new_[20198]_ ;
  assign \new_[20200]_  = \new_[20199]_  & \new_[20194]_ ;
  assign \new_[20204]_  = ~A200 & A167;
  assign \new_[20205]_  = A168 & \new_[20204]_ ;
  assign \new_[20209]_  = ~A233 & ~A232;
  assign \new_[20210]_  = ~A201 & \new_[20209]_ ;
  assign \new_[20211]_  = \new_[20210]_  & \new_[20205]_ ;
  assign \new_[20215]_  = A298 & A266;
  assign \new_[20216]_  = A265 & \new_[20215]_ ;
  assign \new_[20220]_  = A302 & A300;
  assign \new_[20221]_  = ~A299 & \new_[20220]_ ;
  assign \new_[20222]_  = \new_[20221]_  & \new_[20216]_ ;
  assign \new_[20226]_  = ~A200 & A167;
  assign \new_[20227]_  = A168 & \new_[20226]_ ;
  assign \new_[20231]_  = ~A233 & ~A232;
  assign \new_[20232]_  = ~A201 & \new_[20231]_ ;
  assign \new_[20233]_  = \new_[20232]_  & \new_[20227]_ ;
  assign \new_[20237]_  = A298 & ~A267;
  assign \new_[20238]_  = ~A266 & \new_[20237]_ ;
  assign \new_[20242]_  = A301 & A300;
  assign \new_[20243]_  = ~A299 & \new_[20242]_ ;
  assign \new_[20244]_  = \new_[20243]_  & \new_[20238]_ ;
  assign \new_[20248]_  = ~A200 & A167;
  assign \new_[20249]_  = A168 & \new_[20248]_ ;
  assign \new_[20253]_  = ~A233 & ~A232;
  assign \new_[20254]_  = ~A201 & \new_[20253]_ ;
  assign \new_[20255]_  = \new_[20254]_  & \new_[20249]_ ;
  assign \new_[20259]_  = A298 & ~A267;
  assign \new_[20260]_  = ~A266 & \new_[20259]_ ;
  assign \new_[20264]_  = A302 & A300;
  assign \new_[20265]_  = ~A299 & \new_[20264]_ ;
  assign \new_[20266]_  = \new_[20265]_  & \new_[20260]_ ;
  assign \new_[20270]_  = ~A200 & A167;
  assign \new_[20271]_  = A168 & \new_[20270]_ ;
  assign \new_[20275]_  = ~A233 & ~A232;
  assign \new_[20276]_  = ~A201 & \new_[20275]_ ;
  assign \new_[20277]_  = \new_[20276]_  & \new_[20271]_ ;
  assign \new_[20281]_  = A298 & ~A266;
  assign \new_[20282]_  = ~A265 & \new_[20281]_ ;
  assign \new_[20286]_  = A301 & A300;
  assign \new_[20287]_  = ~A299 & \new_[20286]_ ;
  assign \new_[20288]_  = \new_[20287]_  & \new_[20282]_ ;
  assign \new_[20292]_  = ~A200 & A167;
  assign \new_[20293]_  = A168 & \new_[20292]_ ;
  assign \new_[20297]_  = ~A233 & ~A232;
  assign \new_[20298]_  = ~A201 & \new_[20297]_ ;
  assign \new_[20299]_  = \new_[20298]_  & \new_[20293]_ ;
  assign \new_[20303]_  = A298 & ~A266;
  assign \new_[20304]_  = ~A265 & \new_[20303]_ ;
  assign \new_[20308]_  = A302 & A300;
  assign \new_[20309]_  = ~A299 & \new_[20308]_ ;
  assign \new_[20310]_  = \new_[20309]_  & \new_[20304]_ ;
  assign \new_[20314]_  = ~A199 & A167;
  assign \new_[20315]_  = A168 & \new_[20314]_ ;
  assign \new_[20319]_  = A233 & A232;
  assign \new_[20320]_  = ~A200 & \new_[20319]_ ;
  assign \new_[20321]_  = \new_[20320]_  & \new_[20315]_ ;
  assign \new_[20325]_  = A298 & ~A267;
  assign \new_[20326]_  = A265 & \new_[20325]_ ;
  assign \new_[20330]_  = A301 & A300;
  assign \new_[20331]_  = ~A299 & \new_[20330]_ ;
  assign \new_[20332]_  = \new_[20331]_  & \new_[20326]_ ;
  assign \new_[20336]_  = ~A199 & A167;
  assign \new_[20337]_  = A168 & \new_[20336]_ ;
  assign \new_[20341]_  = A233 & A232;
  assign \new_[20342]_  = ~A200 & \new_[20341]_ ;
  assign \new_[20343]_  = \new_[20342]_  & \new_[20337]_ ;
  assign \new_[20347]_  = A298 & ~A267;
  assign \new_[20348]_  = A265 & \new_[20347]_ ;
  assign \new_[20352]_  = A302 & A300;
  assign \new_[20353]_  = ~A299 & \new_[20352]_ ;
  assign \new_[20354]_  = \new_[20353]_  & \new_[20348]_ ;
  assign \new_[20358]_  = ~A199 & A167;
  assign \new_[20359]_  = A168 & \new_[20358]_ ;
  assign \new_[20363]_  = A233 & A232;
  assign \new_[20364]_  = ~A200 & \new_[20363]_ ;
  assign \new_[20365]_  = \new_[20364]_  & \new_[20359]_ ;
  assign \new_[20369]_  = A298 & A266;
  assign \new_[20370]_  = A265 & \new_[20369]_ ;
  assign \new_[20374]_  = A301 & A300;
  assign \new_[20375]_  = ~A299 & \new_[20374]_ ;
  assign \new_[20376]_  = \new_[20375]_  & \new_[20370]_ ;
  assign \new_[20380]_  = ~A199 & A167;
  assign \new_[20381]_  = A168 & \new_[20380]_ ;
  assign \new_[20385]_  = A233 & A232;
  assign \new_[20386]_  = ~A200 & \new_[20385]_ ;
  assign \new_[20387]_  = \new_[20386]_  & \new_[20381]_ ;
  assign \new_[20391]_  = A298 & A266;
  assign \new_[20392]_  = A265 & \new_[20391]_ ;
  assign \new_[20396]_  = A302 & A300;
  assign \new_[20397]_  = ~A299 & \new_[20396]_ ;
  assign \new_[20398]_  = \new_[20397]_  & \new_[20392]_ ;
  assign \new_[20402]_  = ~A199 & A167;
  assign \new_[20403]_  = A168 & \new_[20402]_ ;
  assign \new_[20407]_  = A233 & A232;
  assign \new_[20408]_  = ~A200 & \new_[20407]_ ;
  assign \new_[20409]_  = \new_[20408]_  & \new_[20403]_ ;
  assign \new_[20413]_  = A298 & ~A266;
  assign \new_[20414]_  = ~A265 & \new_[20413]_ ;
  assign \new_[20418]_  = A301 & A300;
  assign \new_[20419]_  = ~A299 & \new_[20418]_ ;
  assign \new_[20420]_  = \new_[20419]_  & \new_[20414]_ ;
  assign \new_[20424]_  = ~A199 & A167;
  assign \new_[20425]_  = A168 & \new_[20424]_ ;
  assign \new_[20429]_  = A233 & A232;
  assign \new_[20430]_  = ~A200 & \new_[20429]_ ;
  assign \new_[20431]_  = \new_[20430]_  & \new_[20425]_ ;
  assign \new_[20435]_  = A298 & ~A266;
  assign \new_[20436]_  = ~A265 & \new_[20435]_ ;
  assign \new_[20440]_  = A302 & A300;
  assign \new_[20441]_  = ~A299 & \new_[20440]_ ;
  assign \new_[20442]_  = \new_[20441]_  & \new_[20436]_ ;
  assign \new_[20446]_  = ~A199 & A167;
  assign \new_[20447]_  = A168 & \new_[20446]_ ;
  assign \new_[20451]_  = ~A235 & ~A233;
  assign \new_[20452]_  = ~A200 & \new_[20451]_ ;
  assign \new_[20453]_  = \new_[20452]_  & \new_[20447]_ ;
  assign \new_[20457]_  = ~A268 & ~A266;
  assign \new_[20458]_  = ~A236 & \new_[20457]_ ;
  assign \new_[20462]_  = A299 & ~A298;
  assign \new_[20463]_  = ~A269 & \new_[20462]_ ;
  assign \new_[20464]_  = \new_[20463]_  & \new_[20458]_ ;
  assign \new_[20468]_  = ~A199 & A167;
  assign \new_[20469]_  = A168 & \new_[20468]_ ;
  assign \new_[20473]_  = ~A234 & ~A233;
  assign \new_[20474]_  = ~A200 & \new_[20473]_ ;
  assign \new_[20475]_  = \new_[20474]_  & \new_[20469]_ ;
  assign \new_[20479]_  = A298 & A266;
  assign \new_[20480]_  = A265 & \new_[20479]_ ;
  assign \new_[20484]_  = A301 & A300;
  assign \new_[20485]_  = ~A299 & \new_[20484]_ ;
  assign \new_[20486]_  = \new_[20485]_  & \new_[20480]_ ;
  assign \new_[20490]_  = ~A199 & A167;
  assign \new_[20491]_  = A168 & \new_[20490]_ ;
  assign \new_[20495]_  = ~A234 & ~A233;
  assign \new_[20496]_  = ~A200 & \new_[20495]_ ;
  assign \new_[20497]_  = \new_[20496]_  & \new_[20491]_ ;
  assign \new_[20501]_  = A298 & A266;
  assign \new_[20502]_  = A265 & \new_[20501]_ ;
  assign \new_[20506]_  = A302 & A300;
  assign \new_[20507]_  = ~A299 & \new_[20506]_ ;
  assign \new_[20508]_  = \new_[20507]_  & \new_[20502]_ ;
  assign \new_[20512]_  = ~A199 & A167;
  assign \new_[20513]_  = A168 & \new_[20512]_ ;
  assign \new_[20517]_  = ~A234 & ~A233;
  assign \new_[20518]_  = ~A200 & \new_[20517]_ ;
  assign \new_[20519]_  = \new_[20518]_  & \new_[20513]_ ;
  assign \new_[20523]_  = A298 & ~A267;
  assign \new_[20524]_  = ~A266 & \new_[20523]_ ;
  assign \new_[20528]_  = A301 & A300;
  assign \new_[20529]_  = ~A299 & \new_[20528]_ ;
  assign \new_[20530]_  = \new_[20529]_  & \new_[20524]_ ;
  assign \new_[20534]_  = ~A199 & A167;
  assign \new_[20535]_  = A168 & \new_[20534]_ ;
  assign \new_[20539]_  = ~A234 & ~A233;
  assign \new_[20540]_  = ~A200 & \new_[20539]_ ;
  assign \new_[20541]_  = \new_[20540]_  & \new_[20535]_ ;
  assign \new_[20545]_  = A298 & ~A267;
  assign \new_[20546]_  = ~A266 & \new_[20545]_ ;
  assign \new_[20550]_  = A302 & A300;
  assign \new_[20551]_  = ~A299 & \new_[20550]_ ;
  assign \new_[20552]_  = \new_[20551]_  & \new_[20546]_ ;
  assign \new_[20556]_  = ~A199 & A167;
  assign \new_[20557]_  = A168 & \new_[20556]_ ;
  assign \new_[20561]_  = ~A234 & ~A233;
  assign \new_[20562]_  = ~A200 & \new_[20561]_ ;
  assign \new_[20563]_  = \new_[20562]_  & \new_[20557]_ ;
  assign \new_[20567]_  = A298 & ~A266;
  assign \new_[20568]_  = ~A265 & \new_[20567]_ ;
  assign \new_[20572]_  = A301 & A300;
  assign \new_[20573]_  = ~A299 & \new_[20572]_ ;
  assign \new_[20574]_  = \new_[20573]_  & \new_[20568]_ ;
  assign \new_[20578]_  = ~A199 & A167;
  assign \new_[20579]_  = A168 & \new_[20578]_ ;
  assign \new_[20583]_  = ~A234 & ~A233;
  assign \new_[20584]_  = ~A200 & \new_[20583]_ ;
  assign \new_[20585]_  = \new_[20584]_  & \new_[20579]_ ;
  assign \new_[20589]_  = A298 & ~A266;
  assign \new_[20590]_  = ~A265 & \new_[20589]_ ;
  assign \new_[20594]_  = A302 & A300;
  assign \new_[20595]_  = ~A299 & \new_[20594]_ ;
  assign \new_[20596]_  = \new_[20595]_  & \new_[20590]_ ;
  assign \new_[20600]_  = ~A199 & A167;
  assign \new_[20601]_  = A168 & \new_[20600]_ ;
  assign \new_[20605]_  = ~A233 & A232;
  assign \new_[20606]_  = ~A200 & \new_[20605]_ ;
  assign \new_[20607]_  = \new_[20606]_  & \new_[20601]_ ;
  assign \new_[20611]_  = A265 & A235;
  assign \new_[20612]_  = A234 & \new_[20611]_ ;
  assign \new_[20616]_  = A268 & A267;
  assign \new_[20617]_  = ~A266 & \new_[20616]_ ;
  assign \new_[20618]_  = \new_[20617]_  & \new_[20612]_ ;
  assign \new_[20622]_  = ~A199 & A167;
  assign \new_[20623]_  = A168 & \new_[20622]_ ;
  assign \new_[20627]_  = ~A233 & A232;
  assign \new_[20628]_  = ~A200 & \new_[20627]_ ;
  assign \new_[20629]_  = \new_[20628]_  & \new_[20623]_ ;
  assign \new_[20633]_  = A265 & A235;
  assign \new_[20634]_  = A234 & \new_[20633]_ ;
  assign \new_[20638]_  = A269 & A267;
  assign \new_[20639]_  = ~A266 & \new_[20638]_ ;
  assign \new_[20640]_  = \new_[20639]_  & \new_[20634]_ ;
  assign \new_[20644]_  = ~A199 & A167;
  assign \new_[20645]_  = A168 & \new_[20644]_ ;
  assign \new_[20649]_  = ~A233 & A232;
  assign \new_[20650]_  = ~A200 & \new_[20649]_ ;
  assign \new_[20651]_  = \new_[20650]_  & \new_[20645]_ ;
  assign \new_[20655]_  = A265 & A236;
  assign \new_[20656]_  = A234 & \new_[20655]_ ;
  assign \new_[20660]_  = A268 & A267;
  assign \new_[20661]_  = ~A266 & \new_[20660]_ ;
  assign \new_[20662]_  = \new_[20661]_  & \new_[20656]_ ;
  assign \new_[20666]_  = ~A199 & A167;
  assign \new_[20667]_  = A168 & \new_[20666]_ ;
  assign \new_[20671]_  = ~A233 & A232;
  assign \new_[20672]_  = ~A200 & \new_[20671]_ ;
  assign \new_[20673]_  = \new_[20672]_  & \new_[20667]_ ;
  assign \new_[20677]_  = A265 & A236;
  assign \new_[20678]_  = A234 & \new_[20677]_ ;
  assign \new_[20682]_  = A269 & A267;
  assign \new_[20683]_  = ~A266 & \new_[20682]_ ;
  assign \new_[20684]_  = \new_[20683]_  & \new_[20678]_ ;
  assign \new_[20688]_  = ~A199 & A167;
  assign \new_[20689]_  = A168 & \new_[20688]_ ;
  assign \new_[20693]_  = ~A233 & ~A232;
  assign \new_[20694]_  = ~A200 & \new_[20693]_ ;
  assign \new_[20695]_  = \new_[20694]_  & \new_[20689]_ ;
  assign \new_[20699]_  = A298 & A266;
  assign \new_[20700]_  = A265 & \new_[20699]_ ;
  assign \new_[20704]_  = A301 & A300;
  assign \new_[20705]_  = ~A299 & \new_[20704]_ ;
  assign \new_[20706]_  = \new_[20705]_  & \new_[20700]_ ;
  assign \new_[20710]_  = ~A199 & A167;
  assign \new_[20711]_  = A168 & \new_[20710]_ ;
  assign \new_[20715]_  = ~A233 & ~A232;
  assign \new_[20716]_  = ~A200 & \new_[20715]_ ;
  assign \new_[20717]_  = \new_[20716]_  & \new_[20711]_ ;
  assign \new_[20721]_  = A298 & A266;
  assign \new_[20722]_  = A265 & \new_[20721]_ ;
  assign \new_[20726]_  = A302 & A300;
  assign \new_[20727]_  = ~A299 & \new_[20726]_ ;
  assign \new_[20728]_  = \new_[20727]_  & \new_[20722]_ ;
  assign \new_[20732]_  = ~A199 & A167;
  assign \new_[20733]_  = A168 & \new_[20732]_ ;
  assign \new_[20737]_  = ~A233 & ~A232;
  assign \new_[20738]_  = ~A200 & \new_[20737]_ ;
  assign \new_[20739]_  = \new_[20738]_  & \new_[20733]_ ;
  assign \new_[20743]_  = A298 & ~A267;
  assign \new_[20744]_  = ~A266 & \new_[20743]_ ;
  assign \new_[20748]_  = A301 & A300;
  assign \new_[20749]_  = ~A299 & \new_[20748]_ ;
  assign \new_[20750]_  = \new_[20749]_  & \new_[20744]_ ;
  assign \new_[20754]_  = ~A199 & A167;
  assign \new_[20755]_  = A168 & \new_[20754]_ ;
  assign \new_[20759]_  = ~A233 & ~A232;
  assign \new_[20760]_  = ~A200 & \new_[20759]_ ;
  assign \new_[20761]_  = \new_[20760]_  & \new_[20755]_ ;
  assign \new_[20765]_  = A298 & ~A267;
  assign \new_[20766]_  = ~A266 & \new_[20765]_ ;
  assign \new_[20770]_  = A302 & A300;
  assign \new_[20771]_  = ~A299 & \new_[20770]_ ;
  assign \new_[20772]_  = \new_[20771]_  & \new_[20766]_ ;
  assign \new_[20776]_  = ~A199 & A167;
  assign \new_[20777]_  = A168 & \new_[20776]_ ;
  assign \new_[20781]_  = ~A233 & ~A232;
  assign \new_[20782]_  = ~A200 & \new_[20781]_ ;
  assign \new_[20783]_  = \new_[20782]_  & \new_[20777]_ ;
  assign \new_[20787]_  = A298 & ~A266;
  assign \new_[20788]_  = ~A265 & \new_[20787]_ ;
  assign \new_[20792]_  = A301 & A300;
  assign \new_[20793]_  = ~A299 & \new_[20792]_ ;
  assign \new_[20794]_  = \new_[20793]_  & \new_[20788]_ ;
  assign \new_[20798]_  = ~A199 & A167;
  assign \new_[20799]_  = A168 & \new_[20798]_ ;
  assign \new_[20803]_  = ~A233 & ~A232;
  assign \new_[20804]_  = ~A200 & \new_[20803]_ ;
  assign \new_[20805]_  = \new_[20804]_  & \new_[20799]_ ;
  assign \new_[20809]_  = A298 & ~A266;
  assign \new_[20810]_  = ~A265 & \new_[20809]_ ;
  assign \new_[20814]_  = A302 & A300;
  assign \new_[20815]_  = ~A299 & \new_[20814]_ ;
  assign \new_[20816]_  = \new_[20815]_  & \new_[20810]_ ;
  assign \new_[20820]_  = ~A166 & ~A167;
  assign \new_[20821]_  = A170 & \new_[20820]_ ;
  assign \new_[20825]_  = A232 & A200;
  assign \new_[20826]_  = ~A199 & \new_[20825]_ ;
  assign \new_[20827]_  = \new_[20826]_  & \new_[20821]_ ;
  assign \new_[20831]_  = ~A268 & A265;
  assign \new_[20832]_  = A233 & \new_[20831]_ ;
  assign \new_[20836]_  = A299 & ~A298;
  assign \new_[20837]_  = ~A269 & \new_[20836]_ ;
  assign \new_[20838]_  = \new_[20837]_  & \new_[20832]_ ;
  assign \new_[20842]_  = ~A166 & ~A167;
  assign \new_[20843]_  = A170 & \new_[20842]_ ;
  assign \new_[20847]_  = ~A233 & A200;
  assign \new_[20848]_  = ~A199 & \new_[20847]_ ;
  assign \new_[20849]_  = \new_[20848]_  & \new_[20843]_ ;
  assign \new_[20853]_  = A265 & ~A236;
  assign \new_[20854]_  = ~A235 & \new_[20853]_ ;
  assign \new_[20858]_  = A299 & ~A298;
  assign \new_[20859]_  = A266 & \new_[20858]_ ;
  assign \new_[20860]_  = \new_[20859]_  & \new_[20854]_ ;
  assign \new_[20864]_  = ~A166 & ~A167;
  assign \new_[20865]_  = A170 & \new_[20864]_ ;
  assign \new_[20869]_  = ~A233 & A200;
  assign \new_[20870]_  = ~A199 & \new_[20869]_ ;
  assign \new_[20871]_  = \new_[20870]_  & \new_[20865]_ ;
  assign \new_[20875]_  = ~A266 & ~A236;
  assign \new_[20876]_  = ~A235 & \new_[20875]_ ;
  assign \new_[20880]_  = A299 & ~A298;
  assign \new_[20881]_  = ~A267 & \new_[20880]_ ;
  assign \new_[20882]_  = \new_[20881]_  & \new_[20876]_ ;
  assign \new_[20886]_  = ~A166 & ~A167;
  assign \new_[20887]_  = A170 & \new_[20886]_ ;
  assign \new_[20891]_  = ~A233 & A200;
  assign \new_[20892]_  = ~A199 & \new_[20891]_ ;
  assign \new_[20893]_  = \new_[20892]_  & \new_[20887]_ ;
  assign \new_[20897]_  = ~A265 & ~A236;
  assign \new_[20898]_  = ~A235 & \new_[20897]_ ;
  assign \new_[20902]_  = A299 & ~A298;
  assign \new_[20903]_  = ~A266 & \new_[20902]_ ;
  assign \new_[20904]_  = \new_[20903]_  & \new_[20898]_ ;
  assign \new_[20908]_  = ~A166 & ~A167;
  assign \new_[20909]_  = A170 & \new_[20908]_ ;
  assign \new_[20913]_  = ~A233 & A200;
  assign \new_[20914]_  = ~A199 & \new_[20913]_ ;
  assign \new_[20915]_  = \new_[20914]_  & \new_[20909]_ ;
  assign \new_[20919]_  = ~A268 & ~A266;
  assign \new_[20920]_  = ~A234 & \new_[20919]_ ;
  assign \new_[20924]_  = A299 & ~A298;
  assign \new_[20925]_  = ~A269 & \new_[20924]_ ;
  assign \new_[20926]_  = \new_[20925]_  & \new_[20920]_ ;
  assign \new_[20930]_  = ~A166 & ~A167;
  assign \new_[20931]_  = A170 & \new_[20930]_ ;
  assign \new_[20935]_  = A232 & A200;
  assign \new_[20936]_  = ~A199 & \new_[20935]_ ;
  assign \new_[20937]_  = \new_[20936]_  & \new_[20931]_ ;
  assign \new_[20941]_  = A235 & A234;
  assign \new_[20942]_  = ~A233 & \new_[20941]_ ;
  assign \new_[20946]_  = ~A302 & ~A301;
  assign \new_[20947]_  = A298 & \new_[20946]_ ;
  assign \new_[20948]_  = \new_[20947]_  & \new_[20942]_ ;
  assign \new_[20952]_  = ~A166 & ~A167;
  assign \new_[20953]_  = A170 & \new_[20952]_ ;
  assign \new_[20957]_  = A232 & A200;
  assign \new_[20958]_  = ~A199 & \new_[20957]_ ;
  assign \new_[20959]_  = \new_[20958]_  & \new_[20953]_ ;
  assign \new_[20963]_  = A236 & A234;
  assign \new_[20964]_  = ~A233 & \new_[20963]_ ;
  assign \new_[20968]_  = ~A302 & ~A301;
  assign \new_[20969]_  = A298 & \new_[20968]_ ;
  assign \new_[20970]_  = \new_[20969]_  & \new_[20964]_ ;
  assign \new_[20974]_  = ~A166 & ~A167;
  assign \new_[20975]_  = A170 & \new_[20974]_ ;
  assign \new_[20979]_  = ~A232 & A200;
  assign \new_[20980]_  = ~A199 & \new_[20979]_ ;
  assign \new_[20981]_  = \new_[20980]_  & \new_[20975]_ ;
  assign \new_[20985]_  = ~A268 & ~A266;
  assign \new_[20986]_  = ~A233 & \new_[20985]_ ;
  assign \new_[20990]_  = A299 & ~A298;
  assign \new_[20991]_  = ~A269 & \new_[20990]_ ;
  assign \new_[20992]_  = \new_[20991]_  & \new_[20986]_ ;
  assign \new_[20996]_  = ~A166 & ~A167;
  assign \new_[20997]_  = A170 & \new_[20996]_ ;
  assign \new_[21001]_  = A201 & ~A200;
  assign \new_[21002]_  = A199 & \new_[21001]_ ;
  assign \new_[21003]_  = \new_[21002]_  & \new_[20997]_ ;
  assign \new_[21007]_  = A233 & ~A232;
  assign \new_[21008]_  = A202 & \new_[21007]_ ;
  assign \new_[21012]_  = ~A302 & ~A301;
  assign \new_[21013]_  = ~A299 & \new_[21012]_ ;
  assign \new_[21014]_  = \new_[21013]_  & \new_[21008]_ ;
  assign \new_[21018]_  = ~A166 & ~A167;
  assign \new_[21019]_  = A170 & \new_[21018]_ ;
  assign \new_[21023]_  = A201 & ~A200;
  assign \new_[21024]_  = A199 & \new_[21023]_ ;
  assign \new_[21025]_  = \new_[21024]_  & \new_[21019]_ ;
  assign \new_[21029]_  = A233 & ~A232;
  assign \new_[21030]_  = A203 & \new_[21029]_ ;
  assign \new_[21034]_  = ~A302 & ~A301;
  assign \new_[21035]_  = ~A299 & \new_[21034]_ ;
  assign \new_[21036]_  = \new_[21035]_  & \new_[21030]_ ;
  assign \new_[21040]_  = A167 & ~A168;
  assign \new_[21041]_  = A170 & \new_[21040]_ ;
  assign \new_[21045]_  = A200 & ~A199;
  assign \new_[21046]_  = A166 & \new_[21045]_ ;
  assign \new_[21047]_  = \new_[21046]_  & \new_[21041]_ ;
  assign \new_[21051]_  = A265 & A233;
  assign \new_[21052]_  = A232 & \new_[21051]_ ;
  assign \new_[21056]_  = A299 & ~A298;
  assign \new_[21057]_  = ~A267 & \new_[21056]_ ;
  assign \new_[21058]_  = \new_[21057]_  & \new_[21052]_ ;
  assign \new_[21062]_  = A167 & ~A168;
  assign \new_[21063]_  = A170 & \new_[21062]_ ;
  assign \new_[21067]_  = A200 & ~A199;
  assign \new_[21068]_  = A166 & \new_[21067]_ ;
  assign \new_[21069]_  = \new_[21068]_  & \new_[21063]_ ;
  assign \new_[21073]_  = A265 & A233;
  assign \new_[21074]_  = A232 & \new_[21073]_ ;
  assign \new_[21078]_  = A299 & ~A298;
  assign \new_[21079]_  = A266 & \new_[21078]_ ;
  assign \new_[21080]_  = \new_[21079]_  & \new_[21074]_ ;
  assign \new_[21084]_  = A167 & ~A168;
  assign \new_[21085]_  = A170 & \new_[21084]_ ;
  assign \new_[21089]_  = A200 & ~A199;
  assign \new_[21090]_  = A166 & \new_[21089]_ ;
  assign \new_[21091]_  = \new_[21090]_  & \new_[21085]_ ;
  assign \new_[21095]_  = ~A265 & A233;
  assign \new_[21096]_  = A232 & \new_[21095]_ ;
  assign \new_[21100]_  = A299 & ~A298;
  assign \new_[21101]_  = ~A266 & \new_[21100]_ ;
  assign \new_[21102]_  = \new_[21101]_  & \new_[21096]_ ;
  assign \new_[21106]_  = A167 & ~A168;
  assign \new_[21107]_  = A170 & \new_[21106]_ ;
  assign \new_[21111]_  = A200 & ~A199;
  assign \new_[21112]_  = A166 & \new_[21111]_ ;
  assign \new_[21113]_  = \new_[21112]_  & \new_[21107]_ ;
  assign \new_[21117]_  = A265 & A233;
  assign \new_[21118]_  = ~A232 & \new_[21117]_ ;
  assign \new_[21122]_  = A268 & A267;
  assign \new_[21123]_  = ~A266 & \new_[21122]_ ;
  assign \new_[21124]_  = \new_[21123]_  & \new_[21118]_ ;
  assign \new_[21128]_  = A167 & ~A168;
  assign \new_[21129]_  = A170 & \new_[21128]_ ;
  assign \new_[21133]_  = A200 & ~A199;
  assign \new_[21134]_  = A166 & \new_[21133]_ ;
  assign \new_[21135]_  = \new_[21134]_  & \new_[21129]_ ;
  assign \new_[21139]_  = A265 & A233;
  assign \new_[21140]_  = ~A232 & \new_[21139]_ ;
  assign \new_[21144]_  = A269 & A267;
  assign \new_[21145]_  = ~A266 & \new_[21144]_ ;
  assign \new_[21146]_  = \new_[21145]_  & \new_[21140]_ ;
  assign \new_[21150]_  = A167 & ~A168;
  assign \new_[21151]_  = A170 & \new_[21150]_ ;
  assign \new_[21155]_  = A200 & ~A199;
  assign \new_[21156]_  = A166 & \new_[21155]_ ;
  assign \new_[21157]_  = \new_[21156]_  & \new_[21151]_ ;
  assign \new_[21161]_  = A265 & ~A234;
  assign \new_[21162]_  = ~A233 & \new_[21161]_ ;
  assign \new_[21166]_  = A299 & ~A298;
  assign \new_[21167]_  = A266 & \new_[21166]_ ;
  assign \new_[21168]_  = \new_[21167]_  & \new_[21162]_ ;
  assign \new_[21172]_  = A167 & ~A168;
  assign \new_[21173]_  = A170 & \new_[21172]_ ;
  assign \new_[21177]_  = A200 & ~A199;
  assign \new_[21178]_  = A166 & \new_[21177]_ ;
  assign \new_[21179]_  = \new_[21178]_  & \new_[21173]_ ;
  assign \new_[21183]_  = ~A266 & ~A234;
  assign \new_[21184]_  = ~A233 & \new_[21183]_ ;
  assign \new_[21188]_  = A299 & ~A298;
  assign \new_[21189]_  = ~A267 & \new_[21188]_ ;
  assign \new_[21190]_  = \new_[21189]_  & \new_[21184]_ ;
  assign \new_[21194]_  = A167 & ~A168;
  assign \new_[21195]_  = A170 & \new_[21194]_ ;
  assign \new_[21199]_  = A200 & ~A199;
  assign \new_[21200]_  = A166 & \new_[21199]_ ;
  assign \new_[21201]_  = \new_[21200]_  & \new_[21195]_ ;
  assign \new_[21205]_  = ~A265 & ~A234;
  assign \new_[21206]_  = ~A233 & \new_[21205]_ ;
  assign \new_[21210]_  = A299 & ~A298;
  assign \new_[21211]_  = ~A266 & \new_[21210]_ ;
  assign \new_[21212]_  = \new_[21211]_  & \new_[21206]_ ;
  assign \new_[21216]_  = A167 & ~A168;
  assign \new_[21217]_  = A170 & \new_[21216]_ ;
  assign \new_[21221]_  = A200 & ~A199;
  assign \new_[21222]_  = A166 & \new_[21221]_ ;
  assign \new_[21223]_  = \new_[21222]_  & \new_[21217]_ ;
  assign \new_[21227]_  = A234 & ~A233;
  assign \new_[21228]_  = A232 & \new_[21227]_ ;
  assign \new_[21232]_  = ~A300 & A298;
  assign \new_[21233]_  = A235 & \new_[21232]_ ;
  assign \new_[21234]_  = \new_[21233]_  & \new_[21228]_ ;
  assign \new_[21238]_  = A167 & ~A168;
  assign \new_[21239]_  = A170 & \new_[21238]_ ;
  assign \new_[21243]_  = A200 & ~A199;
  assign \new_[21244]_  = A166 & \new_[21243]_ ;
  assign \new_[21245]_  = \new_[21244]_  & \new_[21239]_ ;
  assign \new_[21249]_  = A234 & ~A233;
  assign \new_[21250]_  = A232 & \new_[21249]_ ;
  assign \new_[21254]_  = A299 & A298;
  assign \new_[21255]_  = A235 & \new_[21254]_ ;
  assign \new_[21256]_  = \new_[21255]_  & \new_[21250]_ ;
  assign \new_[21260]_  = A167 & ~A168;
  assign \new_[21261]_  = A170 & \new_[21260]_ ;
  assign \new_[21265]_  = A200 & ~A199;
  assign \new_[21266]_  = A166 & \new_[21265]_ ;
  assign \new_[21267]_  = \new_[21266]_  & \new_[21261]_ ;
  assign \new_[21271]_  = A234 & ~A233;
  assign \new_[21272]_  = A232 & \new_[21271]_ ;
  assign \new_[21276]_  = ~A299 & ~A298;
  assign \new_[21277]_  = A235 & \new_[21276]_ ;
  assign \new_[21278]_  = \new_[21277]_  & \new_[21272]_ ;
  assign \new_[21282]_  = A167 & ~A168;
  assign \new_[21283]_  = A170 & \new_[21282]_ ;
  assign \new_[21287]_  = A200 & ~A199;
  assign \new_[21288]_  = A166 & \new_[21287]_ ;
  assign \new_[21289]_  = \new_[21288]_  & \new_[21283]_ ;
  assign \new_[21293]_  = A234 & ~A233;
  assign \new_[21294]_  = A232 & \new_[21293]_ ;
  assign \new_[21298]_  = A266 & ~A265;
  assign \new_[21299]_  = A235 & \new_[21298]_ ;
  assign \new_[21300]_  = \new_[21299]_  & \new_[21294]_ ;
  assign \new_[21304]_  = A167 & ~A168;
  assign \new_[21305]_  = A170 & \new_[21304]_ ;
  assign \new_[21309]_  = A200 & ~A199;
  assign \new_[21310]_  = A166 & \new_[21309]_ ;
  assign \new_[21311]_  = \new_[21310]_  & \new_[21305]_ ;
  assign \new_[21315]_  = A234 & ~A233;
  assign \new_[21316]_  = A232 & \new_[21315]_ ;
  assign \new_[21320]_  = ~A300 & A298;
  assign \new_[21321]_  = A236 & \new_[21320]_ ;
  assign \new_[21322]_  = \new_[21321]_  & \new_[21316]_ ;
  assign \new_[21326]_  = A167 & ~A168;
  assign \new_[21327]_  = A170 & \new_[21326]_ ;
  assign \new_[21331]_  = A200 & ~A199;
  assign \new_[21332]_  = A166 & \new_[21331]_ ;
  assign \new_[21333]_  = \new_[21332]_  & \new_[21327]_ ;
  assign \new_[21337]_  = A234 & ~A233;
  assign \new_[21338]_  = A232 & \new_[21337]_ ;
  assign \new_[21342]_  = A299 & A298;
  assign \new_[21343]_  = A236 & \new_[21342]_ ;
  assign \new_[21344]_  = \new_[21343]_  & \new_[21338]_ ;
  assign \new_[21348]_  = A167 & ~A168;
  assign \new_[21349]_  = A170 & \new_[21348]_ ;
  assign \new_[21353]_  = A200 & ~A199;
  assign \new_[21354]_  = A166 & \new_[21353]_ ;
  assign \new_[21355]_  = \new_[21354]_  & \new_[21349]_ ;
  assign \new_[21359]_  = A234 & ~A233;
  assign \new_[21360]_  = A232 & \new_[21359]_ ;
  assign \new_[21364]_  = ~A299 & ~A298;
  assign \new_[21365]_  = A236 & \new_[21364]_ ;
  assign \new_[21366]_  = \new_[21365]_  & \new_[21360]_ ;
  assign \new_[21370]_  = A167 & ~A168;
  assign \new_[21371]_  = A170 & \new_[21370]_ ;
  assign \new_[21375]_  = A200 & ~A199;
  assign \new_[21376]_  = A166 & \new_[21375]_ ;
  assign \new_[21377]_  = \new_[21376]_  & \new_[21371]_ ;
  assign \new_[21381]_  = A234 & ~A233;
  assign \new_[21382]_  = A232 & \new_[21381]_ ;
  assign \new_[21386]_  = A266 & ~A265;
  assign \new_[21387]_  = A236 & \new_[21386]_ ;
  assign \new_[21388]_  = \new_[21387]_  & \new_[21382]_ ;
  assign \new_[21392]_  = A167 & ~A168;
  assign \new_[21393]_  = A170 & \new_[21392]_ ;
  assign \new_[21397]_  = A200 & ~A199;
  assign \new_[21398]_  = A166 & \new_[21397]_ ;
  assign \new_[21399]_  = \new_[21398]_  & \new_[21393]_ ;
  assign \new_[21403]_  = A265 & ~A233;
  assign \new_[21404]_  = ~A232 & \new_[21403]_ ;
  assign \new_[21408]_  = A299 & ~A298;
  assign \new_[21409]_  = A266 & \new_[21408]_ ;
  assign \new_[21410]_  = \new_[21409]_  & \new_[21404]_ ;
  assign \new_[21414]_  = A167 & ~A168;
  assign \new_[21415]_  = A170 & \new_[21414]_ ;
  assign \new_[21419]_  = A200 & ~A199;
  assign \new_[21420]_  = A166 & \new_[21419]_ ;
  assign \new_[21421]_  = \new_[21420]_  & \new_[21415]_ ;
  assign \new_[21425]_  = ~A266 & ~A233;
  assign \new_[21426]_  = ~A232 & \new_[21425]_ ;
  assign \new_[21430]_  = A299 & ~A298;
  assign \new_[21431]_  = ~A267 & \new_[21430]_ ;
  assign \new_[21432]_  = \new_[21431]_  & \new_[21426]_ ;
  assign \new_[21436]_  = A167 & ~A168;
  assign \new_[21437]_  = A170 & \new_[21436]_ ;
  assign \new_[21441]_  = A200 & ~A199;
  assign \new_[21442]_  = A166 & \new_[21441]_ ;
  assign \new_[21443]_  = \new_[21442]_  & \new_[21437]_ ;
  assign \new_[21447]_  = ~A265 & ~A233;
  assign \new_[21448]_  = ~A232 & \new_[21447]_ ;
  assign \new_[21452]_  = A299 & ~A298;
  assign \new_[21453]_  = ~A266 & \new_[21452]_ ;
  assign \new_[21454]_  = \new_[21453]_  & \new_[21448]_ ;
  assign \new_[21458]_  = A167 & ~A168;
  assign \new_[21459]_  = ~A170 & \new_[21458]_ ;
  assign \new_[21463]_  = A200 & ~A199;
  assign \new_[21464]_  = ~A166 & \new_[21463]_ ;
  assign \new_[21465]_  = \new_[21464]_  & \new_[21459]_ ;
  assign \new_[21469]_  = A265 & A233;
  assign \new_[21470]_  = A232 & \new_[21469]_ ;
  assign \new_[21474]_  = A299 & ~A298;
  assign \new_[21475]_  = ~A267 & \new_[21474]_ ;
  assign \new_[21476]_  = \new_[21475]_  & \new_[21470]_ ;
  assign \new_[21480]_  = A167 & ~A168;
  assign \new_[21481]_  = ~A170 & \new_[21480]_ ;
  assign \new_[21485]_  = A200 & ~A199;
  assign \new_[21486]_  = ~A166 & \new_[21485]_ ;
  assign \new_[21487]_  = \new_[21486]_  & \new_[21481]_ ;
  assign \new_[21491]_  = A265 & A233;
  assign \new_[21492]_  = A232 & \new_[21491]_ ;
  assign \new_[21496]_  = A299 & ~A298;
  assign \new_[21497]_  = A266 & \new_[21496]_ ;
  assign \new_[21498]_  = \new_[21497]_  & \new_[21492]_ ;
  assign \new_[21502]_  = A167 & ~A168;
  assign \new_[21503]_  = ~A170 & \new_[21502]_ ;
  assign \new_[21507]_  = A200 & ~A199;
  assign \new_[21508]_  = ~A166 & \new_[21507]_ ;
  assign \new_[21509]_  = \new_[21508]_  & \new_[21503]_ ;
  assign \new_[21513]_  = ~A265 & A233;
  assign \new_[21514]_  = A232 & \new_[21513]_ ;
  assign \new_[21518]_  = A299 & ~A298;
  assign \new_[21519]_  = ~A266 & \new_[21518]_ ;
  assign \new_[21520]_  = \new_[21519]_  & \new_[21514]_ ;
  assign \new_[21524]_  = A167 & ~A168;
  assign \new_[21525]_  = ~A170 & \new_[21524]_ ;
  assign \new_[21529]_  = A200 & ~A199;
  assign \new_[21530]_  = ~A166 & \new_[21529]_ ;
  assign \new_[21531]_  = \new_[21530]_  & \new_[21525]_ ;
  assign \new_[21535]_  = A265 & A233;
  assign \new_[21536]_  = ~A232 & \new_[21535]_ ;
  assign \new_[21540]_  = A268 & A267;
  assign \new_[21541]_  = ~A266 & \new_[21540]_ ;
  assign \new_[21542]_  = \new_[21541]_  & \new_[21536]_ ;
  assign \new_[21546]_  = A167 & ~A168;
  assign \new_[21547]_  = ~A170 & \new_[21546]_ ;
  assign \new_[21551]_  = A200 & ~A199;
  assign \new_[21552]_  = ~A166 & \new_[21551]_ ;
  assign \new_[21553]_  = \new_[21552]_  & \new_[21547]_ ;
  assign \new_[21557]_  = A265 & A233;
  assign \new_[21558]_  = ~A232 & \new_[21557]_ ;
  assign \new_[21562]_  = A269 & A267;
  assign \new_[21563]_  = ~A266 & \new_[21562]_ ;
  assign \new_[21564]_  = \new_[21563]_  & \new_[21558]_ ;
  assign \new_[21568]_  = A167 & ~A168;
  assign \new_[21569]_  = ~A170 & \new_[21568]_ ;
  assign \new_[21573]_  = A200 & ~A199;
  assign \new_[21574]_  = ~A166 & \new_[21573]_ ;
  assign \new_[21575]_  = \new_[21574]_  & \new_[21569]_ ;
  assign \new_[21579]_  = A265 & ~A234;
  assign \new_[21580]_  = ~A233 & \new_[21579]_ ;
  assign \new_[21584]_  = A299 & ~A298;
  assign \new_[21585]_  = A266 & \new_[21584]_ ;
  assign \new_[21586]_  = \new_[21585]_  & \new_[21580]_ ;
  assign \new_[21590]_  = A167 & ~A168;
  assign \new_[21591]_  = ~A170 & \new_[21590]_ ;
  assign \new_[21595]_  = A200 & ~A199;
  assign \new_[21596]_  = ~A166 & \new_[21595]_ ;
  assign \new_[21597]_  = \new_[21596]_  & \new_[21591]_ ;
  assign \new_[21601]_  = ~A266 & ~A234;
  assign \new_[21602]_  = ~A233 & \new_[21601]_ ;
  assign \new_[21606]_  = A299 & ~A298;
  assign \new_[21607]_  = ~A267 & \new_[21606]_ ;
  assign \new_[21608]_  = \new_[21607]_  & \new_[21602]_ ;
  assign \new_[21612]_  = A167 & ~A168;
  assign \new_[21613]_  = ~A170 & \new_[21612]_ ;
  assign \new_[21617]_  = A200 & ~A199;
  assign \new_[21618]_  = ~A166 & \new_[21617]_ ;
  assign \new_[21619]_  = \new_[21618]_  & \new_[21613]_ ;
  assign \new_[21623]_  = ~A265 & ~A234;
  assign \new_[21624]_  = ~A233 & \new_[21623]_ ;
  assign \new_[21628]_  = A299 & ~A298;
  assign \new_[21629]_  = ~A266 & \new_[21628]_ ;
  assign \new_[21630]_  = \new_[21629]_  & \new_[21624]_ ;
  assign \new_[21634]_  = A167 & ~A168;
  assign \new_[21635]_  = ~A170 & \new_[21634]_ ;
  assign \new_[21639]_  = A200 & ~A199;
  assign \new_[21640]_  = ~A166 & \new_[21639]_ ;
  assign \new_[21641]_  = \new_[21640]_  & \new_[21635]_ ;
  assign \new_[21645]_  = A234 & ~A233;
  assign \new_[21646]_  = A232 & \new_[21645]_ ;
  assign \new_[21650]_  = ~A300 & A298;
  assign \new_[21651]_  = A235 & \new_[21650]_ ;
  assign \new_[21652]_  = \new_[21651]_  & \new_[21646]_ ;
  assign \new_[21656]_  = A167 & ~A168;
  assign \new_[21657]_  = ~A170 & \new_[21656]_ ;
  assign \new_[21661]_  = A200 & ~A199;
  assign \new_[21662]_  = ~A166 & \new_[21661]_ ;
  assign \new_[21663]_  = \new_[21662]_  & \new_[21657]_ ;
  assign \new_[21667]_  = A234 & ~A233;
  assign \new_[21668]_  = A232 & \new_[21667]_ ;
  assign \new_[21672]_  = A299 & A298;
  assign \new_[21673]_  = A235 & \new_[21672]_ ;
  assign \new_[21674]_  = \new_[21673]_  & \new_[21668]_ ;
  assign \new_[21678]_  = A167 & ~A168;
  assign \new_[21679]_  = ~A170 & \new_[21678]_ ;
  assign \new_[21683]_  = A200 & ~A199;
  assign \new_[21684]_  = ~A166 & \new_[21683]_ ;
  assign \new_[21685]_  = \new_[21684]_  & \new_[21679]_ ;
  assign \new_[21689]_  = A234 & ~A233;
  assign \new_[21690]_  = A232 & \new_[21689]_ ;
  assign \new_[21694]_  = ~A299 & ~A298;
  assign \new_[21695]_  = A235 & \new_[21694]_ ;
  assign \new_[21696]_  = \new_[21695]_  & \new_[21690]_ ;
  assign \new_[21700]_  = A167 & ~A168;
  assign \new_[21701]_  = ~A170 & \new_[21700]_ ;
  assign \new_[21705]_  = A200 & ~A199;
  assign \new_[21706]_  = ~A166 & \new_[21705]_ ;
  assign \new_[21707]_  = \new_[21706]_  & \new_[21701]_ ;
  assign \new_[21711]_  = A234 & ~A233;
  assign \new_[21712]_  = A232 & \new_[21711]_ ;
  assign \new_[21716]_  = A266 & ~A265;
  assign \new_[21717]_  = A235 & \new_[21716]_ ;
  assign \new_[21718]_  = \new_[21717]_  & \new_[21712]_ ;
  assign \new_[21722]_  = A167 & ~A168;
  assign \new_[21723]_  = ~A170 & \new_[21722]_ ;
  assign \new_[21727]_  = A200 & ~A199;
  assign \new_[21728]_  = ~A166 & \new_[21727]_ ;
  assign \new_[21729]_  = \new_[21728]_  & \new_[21723]_ ;
  assign \new_[21733]_  = A234 & ~A233;
  assign \new_[21734]_  = A232 & \new_[21733]_ ;
  assign \new_[21738]_  = ~A300 & A298;
  assign \new_[21739]_  = A236 & \new_[21738]_ ;
  assign \new_[21740]_  = \new_[21739]_  & \new_[21734]_ ;
  assign \new_[21744]_  = A167 & ~A168;
  assign \new_[21745]_  = ~A170 & \new_[21744]_ ;
  assign \new_[21749]_  = A200 & ~A199;
  assign \new_[21750]_  = ~A166 & \new_[21749]_ ;
  assign \new_[21751]_  = \new_[21750]_  & \new_[21745]_ ;
  assign \new_[21755]_  = A234 & ~A233;
  assign \new_[21756]_  = A232 & \new_[21755]_ ;
  assign \new_[21760]_  = A299 & A298;
  assign \new_[21761]_  = A236 & \new_[21760]_ ;
  assign \new_[21762]_  = \new_[21761]_  & \new_[21756]_ ;
  assign \new_[21766]_  = A167 & ~A168;
  assign \new_[21767]_  = ~A170 & \new_[21766]_ ;
  assign \new_[21771]_  = A200 & ~A199;
  assign \new_[21772]_  = ~A166 & \new_[21771]_ ;
  assign \new_[21773]_  = \new_[21772]_  & \new_[21767]_ ;
  assign \new_[21777]_  = A234 & ~A233;
  assign \new_[21778]_  = A232 & \new_[21777]_ ;
  assign \new_[21782]_  = ~A299 & ~A298;
  assign \new_[21783]_  = A236 & \new_[21782]_ ;
  assign \new_[21784]_  = \new_[21783]_  & \new_[21778]_ ;
  assign \new_[21788]_  = A167 & ~A168;
  assign \new_[21789]_  = ~A170 & \new_[21788]_ ;
  assign \new_[21793]_  = A200 & ~A199;
  assign \new_[21794]_  = ~A166 & \new_[21793]_ ;
  assign \new_[21795]_  = \new_[21794]_  & \new_[21789]_ ;
  assign \new_[21799]_  = A234 & ~A233;
  assign \new_[21800]_  = A232 & \new_[21799]_ ;
  assign \new_[21804]_  = A266 & ~A265;
  assign \new_[21805]_  = A236 & \new_[21804]_ ;
  assign \new_[21806]_  = \new_[21805]_  & \new_[21800]_ ;
  assign \new_[21810]_  = A167 & ~A168;
  assign \new_[21811]_  = ~A170 & \new_[21810]_ ;
  assign \new_[21815]_  = A200 & ~A199;
  assign \new_[21816]_  = ~A166 & \new_[21815]_ ;
  assign \new_[21817]_  = \new_[21816]_  & \new_[21811]_ ;
  assign \new_[21821]_  = A265 & ~A233;
  assign \new_[21822]_  = ~A232 & \new_[21821]_ ;
  assign \new_[21826]_  = A299 & ~A298;
  assign \new_[21827]_  = A266 & \new_[21826]_ ;
  assign \new_[21828]_  = \new_[21827]_  & \new_[21822]_ ;
  assign \new_[21832]_  = A167 & ~A168;
  assign \new_[21833]_  = ~A170 & \new_[21832]_ ;
  assign \new_[21837]_  = A200 & ~A199;
  assign \new_[21838]_  = ~A166 & \new_[21837]_ ;
  assign \new_[21839]_  = \new_[21838]_  & \new_[21833]_ ;
  assign \new_[21843]_  = ~A266 & ~A233;
  assign \new_[21844]_  = ~A232 & \new_[21843]_ ;
  assign \new_[21848]_  = A299 & ~A298;
  assign \new_[21849]_  = ~A267 & \new_[21848]_ ;
  assign \new_[21850]_  = \new_[21849]_  & \new_[21844]_ ;
  assign \new_[21854]_  = A167 & ~A168;
  assign \new_[21855]_  = ~A170 & \new_[21854]_ ;
  assign \new_[21859]_  = A200 & ~A199;
  assign \new_[21860]_  = ~A166 & \new_[21859]_ ;
  assign \new_[21861]_  = \new_[21860]_  & \new_[21855]_ ;
  assign \new_[21865]_  = ~A265 & ~A233;
  assign \new_[21866]_  = ~A232 & \new_[21865]_ ;
  assign \new_[21870]_  = A299 & ~A298;
  assign \new_[21871]_  = ~A266 & \new_[21870]_ ;
  assign \new_[21872]_  = \new_[21871]_  & \new_[21866]_ ;
  assign \new_[21876]_  = ~A167 & ~A168;
  assign \new_[21877]_  = ~A170 & \new_[21876]_ ;
  assign \new_[21881]_  = A200 & ~A199;
  assign \new_[21882]_  = A166 & \new_[21881]_ ;
  assign \new_[21883]_  = \new_[21882]_  & \new_[21877]_ ;
  assign \new_[21887]_  = A265 & A233;
  assign \new_[21888]_  = A232 & \new_[21887]_ ;
  assign \new_[21892]_  = A299 & ~A298;
  assign \new_[21893]_  = ~A267 & \new_[21892]_ ;
  assign \new_[21894]_  = \new_[21893]_  & \new_[21888]_ ;
  assign \new_[21898]_  = ~A167 & ~A168;
  assign \new_[21899]_  = ~A170 & \new_[21898]_ ;
  assign \new_[21903]_  = A200 & ~A199;
  assign \new_[21904]_  = A166 & \new_[21903]_ ;
  assign \new_[21905]_  = \new_[21904]_  & \new_[21899]_ ;
  assign \new_[21909]_  = A265 & A233;
  assign \new_[21910]_  = A232 & \new_[21909]_ ;
  assign \new_[21914]_  = A299 & ~A298;
  assign \new_[21915]_  = A266 & \new_[21914]_ ;
  assign \new_[21916]_  = \new_[21915]_  & \new_[21910]_ ;
  assign \new_[21920]_  = ~A167 & ~A168;
  assign \new_[21921]_  = ~A170 & \new_[21920]_ ;
  assign \new_[21925]_  = A200 & ~A199;
  assign \new_[21926]_  = A166 & \new_[21925]_ ;
  assign \new_[21927]_  = \new_[21926]_  & \new_[21921]_ ;
  assign \new_[21931]_  = ~A265 & A233;
  assign \new_[21932]_  = A232 & \new_[21931]_ ;
  assign \new_[21936]_  = A299 & ~A298;
  assign \new_[21937]_  = ~A266 & \new_[21936]_ ;
  assign \new_[21938]_  = \new_[21937]_  & \new_[21932]_ ;
  assign \new_[21942]_  = ~A167 & ~A168;
  assign \new_[21943]_  = ~A170 & \new_[21942]_ ;
  assign \new_[21947]_  = A200 & ~A199;
  assign \new_[21948]_  = A166 & \new_[21947]_ ;
  assign \new_[21949]_  = \new_[21948]_  & \new_[21943]_ ;
  assign \new_[21953]_  = A265 & A233;
  assign \new_[21954]_  = ~A232 & \new_[21953]_ ;
  assign \new_[21958]_  = A268 & A267;
  assign \new_[21959]_  = ~A266 & \new_[21958]_ ;
  assign \new_[21960]_  = \new_[21959]_  & \new_[21954]_ ;
  assign \new_[21964]_  = ~A167 & ~A168;
  assign \new_[21965]_  = ~A170 & \new_[21964]_ ;
  assign \new_[21969]_  = A200 & ~A199;
  assign \new_[21970]_  = A166 & \new_[21969]_ ;
  assign \new_[21971]_  = \new_[21970]_  & \new_[21965]_ ;
  assign \new_[21975]_  = A265 & A233;
  assign \new_[21976]_  = ~A232 & \new_[21975]_ ;
  assign \new_[21980]_  = A269 & A267;
  assign \new_[21981]_  = ~A266 & \new_[21980]_ ;
  assign \new_[21982]_  = \new_[21981]_  & \new_[21976]_ ;
  assign \new_[21986]_  = ~A167 & ~A168;
  assign \new_[21987]_  = ~A170 & \new_[21986]_ ;
  assign \new_[21991]_  = A200 & ~A199;
  assign \new_[21992]_  = A166 & \new_[21991]_ ;
  assign \new_[21993]_  = \new_[21992]_  & \new_[21987]_ ;
  assign \new_[21997]_  = A265 & ~A234;
  assign \new_[21998]_  = ~A233 & \new_[21997]_ ;
  assign \new_[22002]_  = A299 & ~A298;
  assign \new_[22003]_  = A266 & \new_[22002]_ ;
  assign \new_[22004]_  = \new_[22003]_  & \new_[21998]_ ;
  assign \new_[22008]_  = ~A167 & ~A168;
  assign \new_[22009]_  = ~A170 & \new_[22008]_ ;
  assign \new_[22013]_  = A200 & ~A199;
  assign \new_[22014]_  = A166 & \new_[22013]_ ;
  assign \new_[22015]_  = \new_[22014]_  & \new_[22009]_ ;
  assign \new_[22019]_  = ~A266 & ~A234;
  assign \new_[22020]_  = ~A233 & \new_[22019]_ ;
  assign \new_[22024]_  = A299 & ~A298;
  assign \new_[22025]_  = ~A267 & \new_[22024]_ ;
  assign \new_[22026]_  = \new_[22025]_  & \new_[22020]_ ;
  assign \new_[22030]_  = ~A167 & ~A168;
  assign \new_[22031]_  = ~A170 & \new_[22030]_ ;
  assign \new_[22035]_  = A200 & ~A199;
  assign \new_[22036]_  = A166 & \new_[22035]_ ;
  assign \new_[22037]_  = \new_[22036]_  & \new_[22031]_ ;
  assign \new_[22041]_  = ~A265 & ~A234;
  assign \new_[22042]_  = ~A233 & \new_[22041]_ ;
  assign \new_[22046]_  = A299 & ~A298;
  assign \new_[22047]_  = ~A266 & \new_[22046]_ ;
  assign \new_[22048]_  = \new_[22047]_  & \new_[22042]_ ;
  assign \new_[22052]_  = ~A167 & ~A168;
  assign \new_[22053]_  = ~A170 & \new_[22052]_ ;
  assign \new_[22057]_  = A200 & ~A199;
  assign \new_[22058]_  = A166 & \new_[22057]_ ;
  assign \new_[22059]_  = \new_[22058]_  & \new_[22053]_ ;
  assign \new_[22063]_  = A234 & ~A233;
  assign \new_[22064]_  = A232 & \new_[22063]_ ;
  assign \new_[22068]_  = ~A300 & A298;
  assign \new_[22069]_  = A235 & \new_[22068]_ ;
  assign \new_[22070]_  = \new_[22069]_  & \new_[22064]_ ;
  assign \new_[22074]_  = ~A167 & ~A168;
  assign \new_[22075]_  = ~A170 & \new_[22074]_ ;
  assign \new_[22079]_  = A200 & ~A199;
  assign \new_[22080]_  = A166 & \new_[22079]_ ;
  assign \new_[22081]_  = \new_[22080]_  & \new_[22075]_ ;
  assign \new_[22085]_  = A234 & ~A233;
  assign \new_[22086]_  = A232 & \new_[22085]_ ;
  assign \new_[22090]_  = A299 & A298;
  assign \new_[22091]_  = A235 & \new_[22090]_ ;
  assign \new_[22092]_  = \new_[22091]_  & \new_[22086]_ ;
  assign \new_[22096]_  = ~A167 & ~A168;
  assign \new_[22097]_  = ~A170 & \new_[22096]_ ;
  assign \new_[22101]_  = A200 & ~A199;
  assign \new_[22102]_  = A166 & \new_[22101]_ ;
  assign \new_[22103]_  = \new_[22102]_  & \new_[22097]_ ;
  assign \new_[22107]_  = A234 & ~A233;
  assign \new_[22108]_  = A232 & \new_[22107]_ ;
  assign \new_[22112]_  = ~A299 & ~A298;
  assign \new_[22113]_  = A235 & \new_[22112]_ ;
  assign \new_[22114]_  = \new_[22113]_  & \new_[22108]_ ;
  assign \new_[22118]_  = ~A167 & ~A168;
  assign \new_[22119]_  = ~A170 & \new_[22118]_ ;
  assign \new_[22123]_  = A200 & ~A199;
  assign \new_[22124]_  = A166 & \new_[22123]_ ;
  assign \new_[22125]_  = \new_[22124]_  & \new_[22119]_ ;
  assign \new_[22129]_  = A234 & ~A233;
  assign \new_[22130]_  = A232 & \new_[22129]_ ;
  assign \new_[22134]_  = A266 & ~A265;
  assign \new_[22135]_  = A235 & \new_[22134]_ ;
  assign \new_[22136]_  = \new_[22135]_  & \new_[22130]_ ;
  assign \new_[22140]_  = ~A167 & ~A168;
  assign \new_[22141]_  = ~A170 & \new_[22140]_ ;
  assign \new_[22145]_  = A200 & ~A199;
  assign \new_[22146]_  = A166 & \new_[22145]_ ;
  assign \new_[22147]_  = \new_[22146]_  & \new_[22141]_ ;
  assign \new_[22151]_  = A234 & ~A233;
  assign \new_[22152]_  = A232 & \new_[22151]_ ;
  assign \new_[22156]_  = ~A300 & A298;
  assign \new_[22157]_  = A236 & \new_[22156]_ ;
  assign \new_[22158]_  = \new_[22157]_  & \new_[22152]_ ;
  assign \new_[22162]_  = ~A167 & ~A168;
  assign \new_[22163]_  = ~A170 & \new_[22162]_ ;
  assign \new_[22167]_  = A200 & ~A199;
  assign \new_[22168]_  = A166 & \new_[22167]_ ;
  assign \new_[22169]_  = \new_[22168]_  & \new_[22163]_ ;
  assign \new_[22173]_  = A234 & ~A233;
  assign \new_[22174]_  = A232 & \new_[22173]_ ;
  assign \new_[22178]_  = A299 & A298;
  assign \new_[22179]_  = A236 & \new_[22178]_ ;
  assign \new_[22180]_  = \new_[22179]_  & \new_[22174]_ ;
  assign \new_[22184]_  = ~A167 & ~A168;
  assign \new_[22185]_  = ~A170 & \new_[22184]_ ;
  assign \new_[22189]_  = A200 & ~A199;
  assign \new_[22190]_  = A166 & \new_[22189]_ ;
  assign \new_[22191]_  = \new_[22190]_  & \new_[22185]_ ;
  assign \new_[22195]_  = A234 & ~A233;
  assign \new_[22196]_  = A232 & \new_[22195]_ ;
  assign \new_[22200]_  = ~A299 & ~A298;
  assign \new_[22201]_  = A236 & \new_[22200]_ ;
  assign \new_[22202]_  = \new_[22201]_  & \new_[22196]_ ;
  assign \new_[22206]_  = ~A167 & ~A168;
  assign \new_[22207]_  = ~A170 & \new_[22206]_ ;
  assign \new_[22211]_  = A200 & ~A199;
  assign \new_[22212]_  = A166 & \new_[22211]_ ;
  assign \new_[22213]_  = \new_[22212]_  & \new_[22207]_ ;
  assign \new_[22217]_  = A234 & ~A233;
  assign \new_[22218]_  = A232 & \new_[22217]_ ;
  assign \new_[22222]_  = A266 & ~A265;
  assign \new_[22223]_  = A236 & \new_[22222]_ ;
  assign \new_[22224]_  = \new_[22223]_  & \new_[22218]_ ;
  assign \new_[22228]_  = ~A167 & ~A168;
  assign \new_[22229]_  = ~A170 & \new_[22228]_ ;
  assign \new_[22233]_  = A200 & ~A199;
  assign \new_[22234]_  = A166 & \new_[22233]_ ;
  assign \new_[22235]_  = \new_[22234]_  & \new_[22229]_ ;
  assign \new_[22239]_  = A265 & ~A233;
  assign \new_[22240]_  = ~A232 & \new_[22239]_ ;
  assign \new_[22244]_  = A299 & ~A298;
  assign \new_[22245]_  = A266 & \new_[22244]_ ;
  assign \new_[22246]_  = \new_[22245]_  & \new_[22240]_ ;
  assign \new_[22250]_  = ~A167 & ~A168;
  assign \new_[22251]_  = ~A170 & \new_[22250]_ ;
  assign \new_[22255]_  = A200 & ~A199;
  assign \new_[22256]_  = A166 & \new_[22255]_ ;
  assign \new_[22257]_  = \new_[22256]_  & \new_[22251]_ ;
  assign \new_[22261]_  = ~A266 & ~A233;
  assign \new_[22262]_  = ~A232 & \new_[22261]_ ;
  assign \new_[22266]_  = A299 & ~A298;
  assign \new_[22267]_  = ~A267 & \new_[22266]_ ;
  assign \new_[22268]_  = \new_[22267]_  & \new_[22262]_ ;
  assign \new_[22272]_  = ~A167 & ~A168;
  assign \new_[22273]_  = ~A170 & \new_[22272]_ ;
  assign \new_[22277]_  = A200 & ~A199;
  assign \new_[22278]_  = A166 & \new_[22277]_ ;
  assign \new_[22279]_  = \new_[22278]_  & \new_[22273]_ ;
  assign \new_[22283]_  = ~A265 & ~A233;
  assign \new_[22284]_  = ~A232 & \new_[22283]_ ;
  assign \new_[22288]_  = A299 & ~A298;
  assign \new_[22289]_  = ~A266 & \new_[22288]_ ;
  assign \new_[22290]_  = \new_[22289]_  & \new_[22284]_ ;
  assign \new_[22294]_  = A167 & ~A168;
  assign \new_[22295]_  = A169 & \new_[22294]_ ;
  assign \new_[22299]_  = A200 & ~A199;
  assign \new_[22300]_  = ~A166 & \new_[22299]_ ;
  assign \new_[22301]_  = \new_[22300]_  & \new_[22295]_ ;
  assign \new_[22305]_  = A265 & A233;
  assign \new_[22306]_  = A232 & \new_[22305]_ ;
  assign \new_[22310]_  = A299 & ~A298;
  assign \new_[22311]_  = ~A267 & \new_[22310]_ ;
  assign \new_[22312]_  = \new_[22311]_  & \new_[22306]_ ;
  assign \new_[22316]_  = A167 & ~A168;
  assign \new_[22317]_  = A169 & \new_[22316]_ ;
  assign \new_[22321]_  = A200 & ~A199;
  assign \new_[22322]_  = ~A166 & \new_[22321]_ ;
  assign \new_[22323]_  = \new_[22322]_  & \new_[22317]_ ;
  assign \new_[22327]_  = A265 & A233;
  assign \new_[22328]_  = A232 & \new_[22327]_ ;
  assign \new_[22332]_  = A299 & ~A298;
  assign \new_[22333]_  = A266 & \new_[22332]_ ;
  assign \new_[22334]_  = \new_[22333]_  & \new_[22328]_ ;
  assign \new_[22338]_  = A167 & ~A168;
  assign \new_[22339]_  = A169 & \new_[22338]_ ;
  assign \new_[22343]_  = A200 & ~A199;
  assign \new_[22344]_  = ~A166 & \new_[22343]_ ;
  assign \new_[22345]_  = \new_[22344]_  & \new_[22339]_ ;
  assign \new_[22349]_  = ~A265 & A233;
  assign \new_[22350]_  = A232 & \new_[22349]_ ;
  assign \new_[22354]_  = A299 & ~A298;
  assign \new_[22355]_  = ~A266 & \new_[22354]_ ;
  assign \new_[22356]_  = \new_[22355]_  & \new_[22350]_ ;
  assign \new_[22360]_  = A167 & ~A168;
  assign \new_[22361]_  = A169 & \new_[22360]_ ;
  assign \new_[22365]_  = A200 & ~A199;
  assign \new_[22366]_  = ~A166 & \new_[22365]_ ;
  assign \new_[22367]_  = \new_[22366]_  & \new_[22361]_ ;
  assign \new_[22371]_  = A265 & A233;
  assign \new_[22372]_  = ~A232 & \new_[22371]_ ;
  assign \new_[22376]_  = A268 & A267;
  assign \new_[22377]_  = ~A266 & \new_[22376]_ ;
  assign \new_[22378]_  = \new_[22377]_  & \new_[22372]_ ;
  assign \new_[22382]_  = A167 & ~A168;
  assign \new_[22383]_  = A169 & \new_[22382]_ ;
  assign \new_[22387]_  = A200 & ~A199;
  assign \new_[22388]_  = ~A166 & \new_[22387]_ ;
  assign \new_[22389]_  = \new_[22388]_  & \new_[22383]_ ;
  assign \new_[22393]_  = A265 & A233;
  assign \new_[22394]_  = ~A232 & \new_[22393]_ ;
  assign \new_[22398]_  = A269 & A267;
  assign \new_[22399]_  = ~A266 & \new_[22398]_ ;
  assign \new_[22400]_  = \new_[22399]_  & \new_[22394]_ ;
  assign \new_[22404]_  = A167 & ~A168;
  assign \new_[22405]_  = A169 & \new_[22404]_ ;
  assign \new_[22409]_  = A200 & ~A199;
  assign \new_[22410]_  = ~A166 & \new_[22409]_ ;
  assign \new_[22411]_  = \new_[22410]_  & \new_[22405]_ ;
  assign \new_[22415]_  = A265 & ~A234;
  assign \new_[22416]_  = ~A233 & \new_[22415]_ ;
  assign \new_[22420]_  = A299 & ~A298;
  assign \new_[22421]_  = A266 & \new_[22420]_ ;
  assign \new_[22422]_  = \new_[22421]_  & \new_[22416]_ ;
  assign \new_[22426]_  = A167 & ~A168;
  assign \new_[22427]_  = A169 & \new_[22426]_ ;
  assign \new_[22431]_  = A200 & ~A199;
  assign \new_[22432]_  = ~A166 & \new_[22431]_ ;
  assign \new_[22433]_  = \new_[22432]_  & \new_[22427]_ ;
  assign \new_[22437]_  = ~A266 & ~A234;
  assign \new_[22438]_  = ~A233 & \new_[22437]_ ;
  assign \new_[22442]_  = A299 & ~A298;
  assign \new_[22443]_  = ~A267 & \new_[22442]_ ;
  assign \new_[22444]_  = \new_[22443]_  & \new_[22438]_ ;
  assign \new_[22448]_  = A167 & ~A168;
  assign \new_[22449]_  = A169 & \new_[22448]_ ;
  assign \new_[22453]_  = A200 & ~A199;
  assign \new_[22454]_  = ~A166 & \new_[22453]_ ;
  assign \new_[22455]_  = \new_[22454]_  & \new_[22449]_ ;
  assign \new_[22459]_  = ~A265 & ~A234;
  assign \new_[22460]_  = ~A233 & \new_[22459]_ ;
  assign \new_[22464]_  = A299 & ~A298;
  assign \new_[22465]_  = ~A266 & \new_[22464]_ ;
  assign \new_[22466]_  = \new_[22465]_  & \new_[22460]_ ;
  assign \new_[22470]_  = A167 & ~A168;
  assign \new_[22471]_  = A169 & \new_[22470]_ ;
  assign \new_[22475]_  = A200 & ~A199;
  assign \new_[22476]_  = ~A166 & \new_[22475]_ ;
  assign \new_[22477]_  = \new_[22476]_  & \new_[22471]_ ;
  assign \new_[22481]_  = A234 & ~A233;
  assign \new_[22482]_  = A232 & \new_[22481]_ ;
  assign \new_[22486]_  = ~A300 & A298;
  assign \new_[22487]_  = A235 & \new_[22486]_ ;
  assign \new_[22488]_  = \new_[22487]_  & \new_[22482]_ ;
  assign \new_[22492]_  = A167 & ~A168;
  assign \new_[22493]_  = A169 & \new_[22492]_ ;
  assign \new_[22497]_  = A200 & ~A199;
  assign \new_[22498]_  = ~A166 & \new_[22497]_ ;
  assign \new_[22499]_  = \new_[22498]_  & \new_[22493]_ ;
  assign \new_[22503]_  = A234 & ~A233;
  assign \new_[22504]_  = A232 & \new_[22503]_ ;
  assign \new_[22508]_  = A299 & A298;
  assign \new_[22509]_  = A235 & \new_[22508]_ ;
  assign \new_[22510]_  = \new_[22509]_  & \new_[22504]_ ;
  assign \new_[22514]_  = A167 & ~A168;
  assign \new_[22515]_  = A169 & \new_[22514]_ ;
  assign \new_[22519]_  = A200 & ~A199;
  assign \new_[22520]_  = ~A166 & \new_[22519]_ ;
  assign \new_[22521]_  = \new_[22520]_  & \new_[22515]_ ;
  assign \new_[22525]_  = A234 & ~A233;
  assign \new_[22526]_  = A232 & \new_[22525]_ ;
  assign \new_[22530]_  = ~A299 & ~A298;
  assign \new_[22531]_  = A235 & \new_[22530]_ ;
  assign \new_[22532]_  = \new_[22531]_  & \new_[22526]_ ;
  assign \new_[22536]_  = A167 & ~A168;
  assign \new_[22537]_  = A169 & \new_[22536]_ ;
  assign \new_[22541]_  = A200 & ~A199;
  assign \new_[22542]_  = ~A166 & \new_[22541]_ ;
  assign \new_[22543]_  = \new_[22542]_  & \new_[22537]_ ;
  assign \new_[22547]_  = A234 & ~A233;
  assign \new_[22548]_  = A232 & \new_[22547]_ ;
  assign \new_[22552]_  = A266 & ~A265;
  assign \new_[22553]_  = A235 & \new_[22552]_ ;
  assign \new_[22554]_  = \new_[22553]_  & \new_[22548]_ ;
  assign \new_[22558]_  = A167 & ~A168;
  assign \new_[22559]_  = A169 & \new_[22558]_ ;
  assign \new_[22563]_  = A200 & ~A199;
  assign \new_[22564]_  = ~A166 & \new_[22563]_ ;
  assign \new_[22565]_  = \new_[22564]_  & \new_[22559]_ ;
  assign \new_[22569]_  = A234 & ~A233;
  assign \new_[22570]_  = A232 & \new_[22569]_ ;
  assign \new_[22574]_  = ~A300 & A298;
  assign \new_[22575]_  = A236 & \new_[22574]_ ;
  assign \new_[22576]_  = \new_[22575]_  & \new_[22570]_ ;
  assign \new_[22580]_  = A167 & ~A168;
  assign \new_[22581]_  = A169 & \new_[22580]_ ;
  assign \new_[22585]_  = A200 & ~A199;
  assign \new_[22586]_  = ~A166 & \new_[22585]_ ;
  assign \new_[22587]_  = \new_[22586]_  & \new_[22581]_ ;
  assign \new_[22591]_  = A234 & ~A233;
  assign \new_[22592]_  = A232 & \new_[22591]_ ;
  assign \new_[22596]_  = A299 & A298;
  assign \new_[22597]_  = A236 & \new_[22596]_ ;
  assign \new_[22598]_  = \new_[22597]_  & \new_[22592]_ ;
  assign \new_[22602]_  = A167 & ~A168;
  assign \new_[22603]_  = A169 & \new_[22602]_ ;
  assign \new_[22607]_  = A200 & ~A199;
  assign \new_[22608]_  = ~A166 & \new_[22607]_ ;
  assign \new_[22609]_  = \new_[22608]_  & \new_[22603]_ ;
  assign \new_[22613]_  = A234 & ~A233;
  assign \new_[22614]_  = A232 & \new_[22613]_ ;
  assign \new_[22618]_  = ~A299 & ~A298;
  assign \new_[22619]_  = A236 & \new_[22618]_ ;
  assign \new_[22620]_  = \new_[22619]_  & \new_[22614]_ ;
  assign \new_[22624]_  = A167 & ~A168;
  assign \new_[22625]_  = A169 & \new_[22624]_ ;
  assign \new_[22629]_  = A200 & ~A199;
  assign \new_[22630]_  = ~A166 & \new_[22629]_ ;
  assign \new_[22631]_  = \new_[22630]_  & \new_[22625]_ ;
  assign \new_[22635]_  = A234 & ~A233;
  assign \new_[22636]_  = A232 & \new_[22635]_ ;
  assign \new_[22640]_  = A266 & ~A265;
  assign \new_[22641]_  = A236 & \new_[22640]_ ;
  assign \new_[22642]_  = \new_[22641]_  & \new_[22636]_ ;
  assign \new_[22646]_  = A167 & ~A168;
  assign \new_[22647]_  = A169 & \new_[22646]_ ;
  assign \new_[22651]_  = A200 & ~A199;
  assign \new_[22652]_  = ~A166 & \new_[22651]_ ;
  assign \new_[22653]_  = \new_[22652]_  & \new_[22647]_ ;
  assign \new_[22657]_  = A265 & ~A233;
  assign \new_[22658]_  = ~A232 & \new_[22657]_ ;
  assign \new_[22662]_  = A299 & ~A298;
  assign \new_[22663]_  = A266 & \new_[22662]_ ;
  assign \new_[22664]_  = \new_[22663]_  & \new_[22658]_ ;
  assign \new_[22668]_  = A167 & ~A168;
  assign \new_[22669]_  = A169 & \new_[22668]_ ;
  assign \new_[22673]_  = A200 & ~A199;
  assign \new_[22674]_  = ~A166 & \new_[22673]_ ;
  assign \new_[22675]_  = \new_[22674]_  & \new_[22669]_ ;
  assign \new_[22679]_  = ~A266 & ~A233;
  assign \new_[22680]_  = ~A232 & \new_[22679]_ ;
  assign \new_[22684]_  = A299 & ~A298;
  assign \new_[22685]_  = ~A267 & \new_[22684]_ ;
  assign \new_[22686]_  = \new_[22685]_  & \new_[22680]_ ;
  assign \new_[22690]_  = A167 & ~A168;
  assign \new_[22691]_  = A169 & \new_[22690]_ ;
  assign \new_[22695]_  = A200 & ~A199;
  assign \new_[22696]_  = ~A166 & \new_[22695]_ ;
  assign \new_[22697]_  = \new_[22696]_  & \new_[22691]_ ;
  assign \new_[22701]_  = ~A265 & ~A233;
  assign \new_[22702]_  = ~A232 & \new_[22701]_ ;
  assign \new_[22706]_  = A299 & ~A298;
  assign \new_[22707]_  = ~A266 & \new_[22706]_ ;
  assign \new_[22708]_  = \new_[22707]_  & \new_[22702]_ ;
  assign \new_[22712]_  = A167 & ~A168;
  assign \new_[22713]_  = A169 & \new_[22712]_ ;
  assign \new_[22717]_  = ~A200 & A199;
  assign \new_[22718]_  = ~A166 & \new_[22717]_ ;
  assign \new_[22719]_  = \new_[22718]_  & \new_[22713]_ ;
  assign \new_[22723]_  = ~A232 & A202;
  assign \new_[22724]_  = A201 & \new_[22723]_ ;
  assign \new_[22728]_  = ~A300 & ~A299;
  assign \new_[22729]_  = A233 & \new_[22728]_ ;
  assign \new_[22730]_  = \new_[22729]_  & \new_[22724]_ ;
  assign \new_[22734]_  = A167 & ~A168;
  assign \new_[22735]_  = A169 & \new_[22734]_ ;
  assign \new_[22739]_  = ~A200 & A199;
  assign \new_[22740]_  = ~A166 & \new_[22739]_ ;
  assign \new_[22741]_  = \new_[22740]_  & \new_[22735]_ ;
  assign \new_[22745]_  = ~A232 & A202;
  assign \new_[22746]_  = A201 & \new_[22745]_ ;
  assign \new_[22750]_  = A299 & A298;
  assign \new_[22751]_  = A233 & \new_[22750]_ ;
  assign \new_[22752]_  = \new_[22751]_  & \new_[22746]_ ;
  assign \new_[22756]_  = A167 & ~A168;
  assign \new_[22757]_  = A169 & \new_[22756]_ ;
  assign \new_[22761]_  = ~A200 & A199;
  assign \new_[22762]_  = ~A166 & \new_[22761]_ ;
  assign \new_[22763]_  = \new_[22762]_  & \new_[22757]_ ;
  assign \new_[22767]_  = ~A232 & A202;
  assign \new_[22768]_  = A201 & \new_[22767]_ ;
  assign \new_[22772]_  = ~A299 & ~A298;
  assign \new_[22773]_  = A233 & \new_[22772]_ ;
  assign \new_[22774]_  = \new_[22773]_  & \new_[22768]_ ;
  assign \new_[22778]_  = A167 & ~A168;
  assign \new_[22779]_  = A169 & \new_[22778]_ ;
  assign \new_[22783]_  = ~A200 & A199;
  assign \new_[22784]_  = ~A166 & \new_[22783]_ ;
  assign \new_[22785]_  = \new_[22784]_  & \new_[22779]_ ;
  assign \new_[22789]_  = ~A232 & A202;
  assign \new_[22790]_  = A201 & \new_[22789]_ ;
  assign \new_[22794]_  = A266 & ~A265;
  assign \new_[22795]_  = A233 & \new_[22794]_ ;
  assign \new_[22796]_  = \new_[22795]_  & \new_[22790]_ ;
  assign \new_[22800]_  = A167 & ~A168;
  assign \new_[22801]_  = A169 & \new_[22800]_ ;
  assign \new_[22805]_  = ~A200 & A199;
  assign \new_[22806]_  = ~A166 & \new_[22805]_ ;
  assign \new_[22807]_  = \new_[22806]_  & \new_[22801]_ ;
  assign \new_[22811]_  = ~A232 & A203;
  assign \new_[22812]_  = A201 & \new_[22811]_ ;
  assign \new_[22816]_  = ~A300 & ~A299;
  assign \new_[22817]_  = A233 & \new_[22816]_ ;
  assign \new_[22818]_  = \new_[22817]_  & \new_[22812]_ ;
  assign \new_[22822]_  = A167 & ~A168;
  assign \new_[22823]_  = A169 & \new_[22822]_ ;
  assign \new_[22827]_  = ~A200 & A199;
  assign \new_[22828]_  = ~A166 & \new_[22827]_ ;
  assign \new_[22829]_  = \new_[22828]_  & \new_[22823]_ ;
  assign \new_[22833]_  = ~A232 & A203;
  assign \new_[22834]_  = A201 & \new_[22833]_ ;
  assign \new_[22838]_  = A299 & A298;
  assign \new_[22839]_  = A233 & \new_[22838]_ ;
  assign \new_[22840]_  = \new_[22839]_  & \new_[22834]_ ;
  assign \new_[22844]_  = A167 & ~A168;
  assign \new_[22845]_  = A169 & \new_[22844]_ ;
  assign \new_[22849]_  = ~A200 & A199;
  assign \new_[22850]_  = ~A166 & \new_[22849]_ ;
  assign \new_[22851]_  = \new_[22850]_  & \new_[22845]_ ;
  assign \new_[22855]_  = ~A232 & A203;
  assign \new_[22856]_  = A201 & \new_[22855]_ ;
  assign \new_[22860]_  = ~A299 & ~A298;
  assign \new_[22861]_  = A233 & \new_[22860]_ ;
  assign \new_[22862]_  = \new_[22861]_  & \new_[22856]_ ;
  assign \new_[22866]_  = A167 & ~A168;
  assign \new_[22867]_  = A169 & \new_[22866]_ ;
  assign \new_[22871]_  = ~A200 & A199;
  assign \new_[22872]_  = ~A166 & \new_[22871]_ ;
  assign \new_[22873]_  = \new_[22872]_  & \new_[22867]_ ;
  assign \new_[22877]_  = ~A232 & A203;
  assign \new_[22878]_  = A201 & \new_[22877]_ ;
  assign \new_[22882]_  = A266 & ~A265;
  assign \new_[22883]_  = A233 & \new_[22882]_ ;
  assign \new_[22884]_  = \new_[22883]_  & \new_[22878]_ ;
  assign \new_[22888]_  = ~A167 & ~A168;
  assign \new_[22889]_  = A169 & \new_[22888]_ ;
  assign \new_[22893]_  = A200 & ~A199;
  assign \new_[22894]_  = A166 & \new_[22893]_ ;
  assign \new_[22895]_  = \new_[22894]_  & \new_[22889]_ ;
  assign \new_[22899]_  = A265 & A233;
  assign \new_[22900]_  = A232 & \new_[22899]_ ;
  assign \new_[22904]_  = A299 & ~A298;
  assign \new_[22905]_  = ~A267 & \new_[22904]_ ;
  assign \new_[22906]_  = \new_[22905]_  & \new_[22900]_ ;
  assign \new_[22910]_  = ~A167 & ~A168;
  assign \new_[22911]_  = A169 & \new_[22910]_ ;
  assign \new_[22915]_  = A200 & ~A199;
  assign \new_[22916]_  = A166 & \new_[22915]_ ;
  assign \new_[22917]_  = \new_[22916]_  & \new_[22911]_ ;
  assign \new_[22921]_  = A265 & A233;
  assign \new_[22922]_  = A232 & \new_[22921]_ ;
  assign \new_[22926]_  = A299 & ~A298;
  assign \new_[22927]_  = A266 & \new_[22926]_ ;
  assign \new_[22928]_  = \new_[22927]_  & \new_[22922]_ ;
  assign \new_[22932]_  = ~A167 & ~A168;
  assign \new_[22933]_  = A169 & \new_[22932]_ ;
  assign \new_[22937]_  = A200 & ~A199;
  assign \new_[22938]_  = A166 & \new_[22937]_ ;
  assign \new_[22939]_  = \new_[22938]_  & \new_[22933]_ ;
  assign \new_[22943]_  = ~A265 & A233;
  assign \new_[22944]_  = A232 & \new_[22943]_ ;
  assign \new_[22948]_  = A299 & ~A298;
  assign \new_[22949]_  = ~A266 & \new_[22948]_ ;
  assign \new_[22950]_  = \new_[22949]_  & \new_[22944]_ ;
  assign \new_[22954]_  = ~A167 & ~A168;
  assign \new_[22955]_  = A169 & \new_[22954]_ ;
  assign \new_[22959]_  = A200 & ~A199;
  assign \new_[22960]_  = A166 & \new_[22959]_ ;
  assign \new_[22961]_  = \new_[22960]_  & \new_[22955]_ ;
  assign \new_[22965]_  = A265 & A233;
  assign \new_[22966]_  = ~A232 & \new_[22965]_ ;
  assign \new_[22970]_  = A268 & A267;
  assign \new_[22971]_  = ~A266 & \new_[22970]_ ;
  assign \new_[22972]_  = \new_[22971]_  & \new_[22966]_ ;
  assign \new_[22976]_  = ~A167 & ~A168;
  assign \new_[22977]_  = A169 & \new_[22976]_ ;
  assign \new_[22981]_  = A200 & ~A199;
  assign \new_[22982]_  = A166 & \new_[22981]_ ;
  assign \new_[22983]_  = \new_[22982]_  & \new_[22977]_ ;
  assign \new_[22987]_  = A265 & A233;
  assign \new_[22988]_  = ~A232 & \new_[22987]_ ;
  assign \new_[22992]_  = A269 & A267;
  assign \new_[22993]_  = ~A266 & \new_[22992]_ ;
  assign \new_[22994]_  = \new_[22993]_  & \new_[22988]_ ;
  assign \new_[22998]_  = ~A167 & ~A168;
  assign \new_[22999]_  = A169 & \new_[22998]_ ;
  assign \new_[23003]_  = A200 & ~A199;
  assign \new_[23004]_  = A166 & \new_[23003]_ ;
  assign \new_[23005]_  = \new_[23004]_  & \new_[22999]_ ;
  assign \new_[23009]_  = A265 & ~A234;
  assign \new_[23010]_  = ~A233 & \new_[23009]_ ;
  assign \new_[23014]_  = A299 & ~A298;
  assign \new_[23015]_  = A266 & \new_[23014]_ ;
  assign \new_[23016]_  = \new_[23015]_  & \new_[23010]_ ;
  assign \new_[23020]_  = ~A167 & ~A168;
  assign \new_[23021]_  = A169 & \new_[23020]_ ;
  assign \new_[23025]_  = A200 & ~A199;
  assign \new_[23026]_  = A166 & \new_[23025]_ ;
  assign \new_[23027]_  = \new_[23026]_  & \new_[23021]_ ;
  assign \new_[23031]_  = ~A266 & ~A234;
  assign \new_[23032]_  = ~A233 & \new_[23031]_ ;
  assign \new_[23036]_  = A299 & ~A298;
  assign \new_[23037]_  = ~A267 & \new_[23036]_ ;
  assign \new_[23038]_  = \new_[23037]_  & \new_[23032]_ ;
  assign \new_[23042]_  = ~A167 & ~A168;
  assign \new_[23043]_  = A169 & \new_[23042]_ ;
  assign \new_[23047]_  = A200 & ~A199;
  assign \new_[23048]_  = A166 & \new_[23047]_ ;
  assign \new_[23049]_  = \new_[23048]_  & \new_[23043]_ ;
  assign \new_[23053]_  = ~A265 & ~A234;
  assign \new_[23054]_  = ~A233 & \new_[23053]_ ;
  assign \new_[23058]_  = A299 & ~A298;
  assign \new_[23059]_  = ~A266 & \new_[23058]_ ;
  assign \new_[23060]_  = \new_[23059]_  & \new_[23054]_ ;
  assign \new_[23064]_  = ~A167 & ~A168;
  assign \new_[23065]_  = A169 & \new_[23064]_ ;
  assign \new_[23069]_  = A200 & ~A199;
  assign \new_[23070]_  = A166 & \new_[23069]_ ;
  assign \new_[23071]_  = \new_[23070]_  & \new_[23065]_ ;
  assign \new_[23075]_  = A234 & ~A233;
  assign \new_[23076]_  = A232 & \new_[23075]_ ;
  assign \new_[23080]_  = ~A300 & A298;
  assign \new_[23081]_  = A235 & \new_[23080]_ ;
  assign \new_[23082]_  = \new_[23081]_  & \new_[23076]_ ;
  assign \new_[23086]_  = ~A167 & ~A168;
  assign \new_[23087]_  = A169 & \new_[23086]_ ;
  assign \new_[23091]_  = A200 & ~A199;
  assign \new_[23092]_  = A166 & \new_[23091]_ ;
  assign \new_[23093]_  = \new_[23092]_  & \new_[23087]_ ;
  assign \new_[23097]_  = A234 & ~A233;
  assign \new_[23098]_  = A232 & \new_[23097]_ ;
  assign \new_[23102]_  = A299 & A298;
  assign \new_[23103]_  = A235 & \new_[23102]_ ;
  assign \new_[23104]_  = \new_[23103]_  & \new_[23098]_ ;
  assign \new_[23108]_  = ~A167 & ~A168;
  assign \new_[23109]_  = A169 & \new_[23108]_ ;
  assign \new_[23113]_  = A200 & ~A199;
  assign \new_[23114]_  = A166 & \new_[23113]_ ;
  assign \new_[23115]_  = \new_[23114]_  & \new_[23109]_ ;
  assign \new_[23119]_  = A234 & ~A233;
  assign \new_[23120]_  = A232 & \new_[23119]_ ;
  assign \new_[23124]_  = ~A299 & ~A298;
  assign \new_[23125]_  = A235 & \new_[23124]_ ;
  assign \new_[23126]_  = \new_[23125]_  & \new_[23120]_ ;
  assign \new_[23130]_  = ~A167 & ~A168;
  assign \new_[23131]_  = A169 & \new_[23130]_ ;
  assign \new_[23135]_  = A200 & ~A199;
  assign \new_[23136]_  = A166 & \new_[23135]_ ;
  assign \new_[23137]_  = \new_[23136]_  & \new_[23131]_ ;
  assign \new_[23141]_  = A234 & ~A233;
  assign \new_[23142]_  = A232 & \new_[23141]_ ;
  assign \new_[23146]_  = A266 & ~A265;
  assign \new_[23147]_  = A235 & \new_[23146]_ ;
  assign \new_[23148]_  = \new_[23147]_  & \new_[23142]_ ;
  assign \new_[23152]_  = ~A167 & ~A168;
  assign \new_[23153]_  = A169 & \new_[23152]_ ;
  assign \new_[23157]_  = A200 & ~A199;
  assign \new_[23158]_  = A166 & \new_[23157]_ ;
  assign \new_[23159]_  = \new_[23158]_  & \new_[23153]_ ;
  assign \new_[23163]_  = A234 & ~A233;
  assign \new_[23164]_  = A232 & \new_[23163]_ ;
  assign \new_[23168]_  = ~A300 & A298;
  assign \new_[23169]_  = A236 & \new_[23168]_ ;
  assign \new_[23170]_  = \new_[23169]_  & \new_[23164]_ ;
  assign \new_[23174]_  = ~A167 & ~A168;
  assign \new_[23175]_  = A169 & \new_[23174]_ ;
  assign \new_[23179]_  = A200 & ~A199;
  assign \new_[23180]_  = A166 & \new_[23179]_ ;
  assign \new_[23181]_  = \new_[23180]_  & \new_[23175]_ ;
  assign \new_[23185]_  = A234 & ~A233;
  assign \new_[23186]_  = A232 & \new_[23185]_ ;
  assign \new_[23190]_  = A299 & A298;
  assign \new_[23191]_  = A236 & \new_[23190]_ ;
  assign \new_[23192]_  = \new_[23191]_  & \new_[23186]_ ;
  assign \new_[23196]_  = ~A167 & ~A168;
  assign \new_[23197]_  = A169 & \new_[23196]_ ;
  assign \new_[23201]_  = A200 & ~A199;
  assign \new_[23202]_  = A166 & \new_[23201]_ ;
  assign \new_[23203]_  = \new_[23202]_  & \new_[23197]_ ;
  assign \new_[23207]_  = A234 & ~A233;
  assign \new_[23208]_  = A232 & \new_[23207]_ ;
  assign \new_[23212]_  = ~A299 & ~A298;
  assign \new_[23213]_  = A236 & \new_[23212]_ ;
  assign \new_[23214]_  = \new_[23213]_  & \new_[23208]_ ;
  assign \new_[23218]_  = ~A167 & ~A168;
  assign \new_[23219]_  = A169 & \new_[23218]_ ;
  assign \new_[23223]_  = A200 & ~A199;
  assign \new_[23224]_  = A166 & \new_[23223]_ ;
  assign \new_[23225]_  = \new_[23224]_  & \new_[23219]_ ;
  assign \new_[23229]_  = A234 & ~A233;
  assign \new_[23230]_  = A232 & \new_[23229]_ ;
  assign \new_[23234]_  = A266 & ~A265;
  assign \new_[23235]_  = A236 & \new_[23234]_ ;
  assign \new_[23236]_  = \new_[23235]_  & \new_[23230]_ ;
  assign \new_[23240]_  = ~A167 & ~A168;
  assign \new_[23241]_  = A169 & \new_[23240]_ ;
  assign \new_[23245]_  = A200 & ~A199;
  assign \new_[23246]_  = A166 & \new_[23245]_ ;
  assign \new_[23247]_  = \new_[23246]_  & \new_[23241]_ ;
  assign \new_[23251]_  = A265 & ~A233;
  assign \new_[23252]_  = ~A232 & \new_[23251]_ ;
  assign \new_[23256]_  = A299 & ~A298;
  assign \new_[23257]_  = A266 & \new_[23256]_ ;
  assign \new_[23258]_  = \new_[23257]_  & \new_[23252]_ ;
  assign \new_[23262]_  = ~A167 & ~A168;
  assign \new_[23263]_  = A169 & \new_[23262]_ ;
  assign \new_[23267]_  = A200 & ~A199;
  assign \new_[23268]_  = A166 & \new_[23267]_ ;
  assign \new_[23269]_  = \new_[23268]_  & \new_[23263]_ ;
  assign \new_[23273]_  = ~A266 & ~A233;
  assign \new_[23274]_  = ~A232 & \new_[23273]_ ;
  assign \new_[23278]_  = A299 & ~A298;
  assign \new_[23279]_  = ~A267 & \new_[23278]_ ;
  assign \new_[23280]_  = \new_[23279]_  & \new_[23274]_ ;
  assign \new_[23284]_  = ~A167 & ~A168;
  assign \new_[23285]_  = A169 & \new_[23284]_ ;
  assign \new_[23289]_  = A200 & ~A199;
  assign \new_[23290]_  = A166 & \new_[23289]_ ;
  assign \new_[23291]_  = \new_[23290]_  & \new_[23285]_ ;
  assign \new_[23295]_  = ~A265 & ~A233;
  assign \new_[23296]_  = ~A232 & \new_[23295]_ ;
  assign \new_[23300]_  = A299 & ~A298;
  assign \new_[23301]_  = ~A266 & \new_[23300]_ ;
  assign \new_[23302]_  = \new_[23301]_  & \new_[23296]_ ;
  assign \new_[23306]_  = ~A167 & ~A168;
  assign \new_[23307]_  = A169 & \new_[23306]_ ;
  assign \new_[23311]_  = ~A200 & A199;
  assign \new_[23312]_  = A166 & \new_[23311]_ ;
  assign \new_[23313]_  = \new_[23312]_  & \new_[23307]_ ;
  assign \new_[23317]_  = ~A232 & A202;
  assign \new_[23318]_  = A201 & \new_[23317]_ ;
  assign \new_[23322]_  = ~A300 & ~A299;
  assign \new_[23323]_  = A233 & \new_[23322]_ ;
  assign \new_[23324]_  = \new_[23323]_  & \new_[23318]_ ;
  assign \new_[23328]_  = ~A167 & ~A168;
  assign \new_[23329]_  = A169 & \new_[23328]_ ;
  assign \new_[23333]_  = ~A200 & A199;
  assign \new_[23334]_  = A166 & \new_[23333]_ ;
  assign \new_[23335]_  = \new_[23334]_  & \new_[23329]_ ;
  assign \new_[23339]_  = ~A232 & A202;
  assign \new_[23340]_  = A201 & \new_[23339]_ ;
  assign \new_[23344]_  = A299 & A298;
  assign \new_[23345]_  = A233 & \new_[23344]_ ;
  assign \new_[23346]_  = \new_[23345]_  & \new_[23340]_ ;
  assign \new_[23350]_  = ~A167 & ~A168;
  assign \new_[23351]_  = A169 & \new_[23350]_ ;
  assign \new_[23355]_  = ~A200 & A199;
  assign \new_[23356]_  = A166 & \new_[23355]_ ;
  assign \new_[23357]_  = \new_[23356]_  & \new_[23351]_ ;
  assign \new_[23361]_  = ~A232 & A202;
  assign \new_[23362]_  = A201 & \new_[23361]_ ;
  assign \new_[23366]_  = ~A299 & ~A298;
  assign \new_[23367]_  = A233 & \new_[23366]_ ;
  assign \new_[23368]_  = \new_[23367]_  & \new_[23362]_ ;
  assign \new_[23372]_  = ~A167 & ~A168;
  assign \new_[23373]_  = A169 & \new_[23372]_ ;
  assign \new_[23377]_  = ~A200 & A199;
  assign \new_[23378]_  = A166 & \new_[23377]_ ;
  assign \new_[23379]_  = \new_[23378]_  & \new_[23373]_ ;
  assign \new_[23383]_  = ~A232 & A202;
  assign \new_[23384]_  = A201 & \new_[23383]_ ;
  assign \new_[23388]_  = A266 & ~A265;
  assign \new_[23389]_  = A233 & \new_[23388]_ ;
  assign \new_[23390]_  = \new_[23389]_  & \new_[23384]_ ;
  assign \new_[23394]_  = ~A167 & ~A168;
  assign \new_[23395]_  = A169 & \new_[23394]_ ;
  assign \new_[23399]_  = ~A200 & A199;
  assign \new_[23400]_  = A166 & \new_[23399]_ ;
  assign \new_[23401]_  = \new_[23400]_  & \new_[23395]_ ;
  assign \new_[23405]_  = ~A232 & A203;
  assign \new_[23406]_  = A201 & \new_[23405]_ ;
  assign \new_[23410]_  = ~A300 & ~A299;
  assign \new_[23411]_  = A233 & \new_[23410]_ ;
  assign \new_[23412]_  = \new_[23411]_  & \new_[23406]_ ;
  assign \new_[23416]_  = ~A167 & ~A168;
  assign \new_[23417]_  = A169 & \new_[23416]_ ;
  assign \new_[23421]_  = ~A200 & A199;
  assign \new_[23422]_  = A166 & \new_[23421]_ ;
  assign \new_[23423]_  = \new_[23422]_  & \new_[23417]_ ;
  assign \new_[23427]_  = ~A232 & A203;
  assign \new_[23428]_  = A201 & \new_[23427]_ ;
  assign \new_[23432]_  = A299 & A298;
  assign \new_[23433]_  = A233 & \new_[23432]_ ;
  assign \new_[23434]_  = \new_[23433]_  & \new_[23428]_ ;
  assign \new_[23438]_  = ~A167 & ~A168;
  assign \new_[23439]_  = A169 & \new_[23438]_ ;
  assign \new_[23443]_  = ~A200 & A199;
  assign \new_[23444]_  = A166 & \new_[23443]_ ;
  assign \new_[23445]_  = \new_[23444]_  & \new_[23439]_ ;
  assign \new_[23449]_  = ~A232 & A203;
  assign \new_[23450]_  = A201 & \new_[23449]_ ;
  assign \new_[23454]_  = ~A299 & ~A298;
  assign \new_[23455]_  = A233 & \new_[23454]_ ;
  assign \new_[23456]_  = \new_[23455]_  & \new_[23450]_ ;
  assign \new_[23460]_  = ~A167 & ~A168;
  assign \new_[23461]_  = A169 & \new_[23460]_ ;
  assign \new_[23465]_  = ~A200 & A199;
  assign \new_[23466]_  = A166 & \new_[23465]_ ;
  assign \new_[23467]_  = \new_[23466]_  & \new_[23461]_ ;
  assign \new_[23471]_  = ~A232 & A203;
  assign \new_[23472]_  = A201 & \new_[23471]_ ;
  assign \new_[23476]_  = A266 & ~A265;
  assign \new_[23477]_  = A233 & \new_[23476]_ ;
  assign \new_[23478]_  = \new_[23477]_  & \new_[23472]_ ;
  assign \new_[23482]_  = ~A168 & A169;
  assign \new_[23483]_  = A170 & \new_[23482]_ ;
  assign \new_[23487]_  = A201 & ~A200;
  assign \new_[23488]_  = A199 & \new_[23487]_ ;
  assign \new_[23489]_  = \new_[23488]_  & \new_[23483]_ ;
  assign \new_[23493]_  = A233 & ~A232;
  assign \new_[23494]_  = A202 & \new_[23493]_ ;
  assign \new_[23498]_  = ~A302 & ~A301;
  assign \new_[23499]_  = ~A299 & \new_[23498]_ ;
  assign \new_[23500]_  = \new_[23499]_  & \new_[23494]_ ;
  assign \new_[23504]_  = ~A168 & A169;
  assign \new_[23505]_  = A170 & \new_[23504]_ ;
  assign \new_[23509]_  = A201 & ~A200;
  assign \new_[23510]_  = A199 & \new_[23509]_ ;
  assign \new_[23511]_  = \new_[23510]_  & \new_[23505]_ ;
  assign \new_[23515]_  = A233 & ~A232;
  assign \new_[23516]_  = A203 & \new_[23515]_ ;
  assign \new_[23520]_  = ~A302 & ~A301;
  assign \new_[23521]_  = ~A299 & \new_[23520]_ ;
  assign \new_[23522]_  = \new_[23521]_  & \new_[23516]_ ;
  assign \new_[23526]_  = A167 & A169;
  assign \new_[23527]_  = ~A170 & \new_[23526]_ ;
  assign \new_[23531]_  = A200 & A199;
  assign \new_[23532]_  = A166 & \new_[23531]_ ;
  assign \new_[23533]_  = \new_[23532]_  & \new_[23527]_ ;
  assign \new_[23537]_  = A265 & A233;
  assign \new_[23538]_  = A232 & \new_[23537]_ ;
  assign \new_[23542]_  = A299 & ~A298;
  assign \new_[23543]_  = ~A267 & \new_[23542]_ ;
  assign \new_[23544]_  = \new_[23543]_  & \new_[23538]_ ;
  assign \new_[23548]_  = A167 & A169;
  assign \new_[23549]_  = ~A170 & \new_[23548]_ ;
  assign \new_[23553]_  = A200 & A199;
  assign \new_[23554]_  = A166 & \new_[23553]_ ;
  assign \new_[23555]_  = \new_[23554]_  & \new_[23549]_ ;
  assign \new_[23559]_  = A265 & A233;
  assign \new_[23560]_  = A232 & \new_[23559]_ ;
  assign \new_[23564]_  = A299 & ~A298;
  assign \new_[23565]_  = A266 & \new_[23564]_ ;
  assign \new_[23566]_  = \new_[23565]_  & \new_[23560]_ ;
  assign \new_[23570]_  = A167 & A169;
  assign \new_[23571]_  = ~A170 & \new_[23570]_ ;
  assign \new_[23575]_  = A200 & A199;
  assign \new_[23576]_  = A166 & \new_[23575]_ ;
  assign \new_[23577]_  = \new_[23576]_  & \new_[23571]_ ;
  assign \new_[23581]_  = ~A265 & A233;
  assign \new_[23582]_  = A232 & \new_[23581]_ ;
  assign \new_[23586]_  = A299 & ~A298;
  assign \new_[23587]_  = ~A266 & \new_[23586]_ ;
  assign \new_[23588]_  = \new_[23587]_  & \new_[23582]_ ;
  assign \new_[23592]_  = A167 & A169;
  assign \new_[23593]_  = ~A170 & \new_[23592]_ ;
  assign \new_[23597]_  = A200 & A199;
  assign \new_[23598]_  = A166 & \new_[23597]_ ;
  assign \new_[23599]_  = \new_[23598]_  & \new_[23593]_ ;
  assign \new_[23603]_  = A265 & A233;
  assign \new_[23604]_  = ~A232 & \new_[23603]_ ;
  assign \new_[23608]_  = A268 & A267;
  assign \new_[23609]_  = ~A266 & \new_[23608]_ ;
  assign \new_[23610]_  = \new_[23609]_  & \new_[23604]_ ;
  assign \new_[23614]_  = A167 & A169;
  assign \new_[23615]_  = ~A170 & \new_[23614]_ ;
  assign \new_[23619]_  = A200 & A199;
  assign \new_[23620]_  = A166 & \new_[23619]_ ;
  assign \new_[23621]_  = \new_[23620]_  & \new_[23615]_ ;
  assign \new_[23625]_  = A265 & A233;
  assign \new_[23626]_  = ~A232 & \new_[23625]_ ;
  assign \new_[23630]_  = A269 & A267;
  assign \new_[23631]_  = ~A266 & \new_[23630]_ ;
  assign \new_[23632]_  = \new_[23631]_  & \new_[23626]_ ;
  assign \new_[23636]_  = A167 & A169;
  assign \new_[23637]_  = ~A170 & \new_[23636]_ ;
  assign \new_[23641]_  = A200 & A199;
  assign \new_[23642]_  = A166 & \new_[23641]_ ;
  assign \new_[23643]_  = \new_[23642]_  & \new_[23637]_ ;
  assign \new_[23647]_  = A265 & ~A234;
  assign \new_[23648]_  = ~A233 & \new_[23647]_ ;
  assign \new_[23652]_  = A299 & ~A298;
  assign \new_[23653]_  = A266 & \new_[23652]_ ;
  assign \new_[23654]_  = \new_[23653]_  & \new_[23648]_ ;
  assign \new_[23658]_  = A167 & A169;
  assign \new_[23659]_  = ~A170 & \new_[23658]_ ;
  assign \new_[23663]_  = A200 & A199;
  assign \new_[23664]_  = A166 & \new_[23663]_ ;
  assign \new_[23665]_  = \new_[23664]_  & \new_[23659]_ ;
  assign \new_[23669]_  = ~A266 & ~A234;
  assign \new_[23670]_  = ~A233 & \new_[23669]_ ;
  assign \new_[23674]_  = A299 & ~A298;
  assign \new_[23675]_  = ~A267 & \new_[23674]_ ;
  assign \new_[23676]_  = \new_[23675]_  & \new_[23670]_ ;
  assign \new_[23680]_  = A167 & A169;
  assign \new_[23681]_  = ~A170 & \new_[23680]_ ;
  assign \new_[23685]_  = A200 & A199;
  assign \new_[23686]_  = A166 & \new_[23685]_ ;
  assign \new_[23687]_  = \new_[23686]_  & \new_[23681]_ ;
  assign \new_[23691]_  = ~A265 & ~A234;
  assign \new_[23692]_  = ~A233 & \new_[23691]_ ;
  assign \new_[23696]_  = A299 & ~A298;
  assign \new_[23697]_  = ~A266 & \new_[23696]_ ;
  assign \new_[23698]_  = \new_[23697]_  & \new_[23692]_ ;
  assign \new_[23702]_  = A167 & A169;
  assign \new_[23703]_  = ~A170 & \new_[23702]_ ;
  assign \new_[23707]_  = A200 & A199;
  assign \new_[23708]_  = A166 & \new_[23707]_ ;
  assign \new_[23709]_  = \new_[23708]_  & \new_[23703]_ ;
  assign \new_[23713]_  = A234 & ~A233;
  assign \new_[23714]_  = A232 & \new_[23713]_ ;
  assign \new_[23718]_  = ~A300 & A298;
  assign \new_[23719]_  = A235 & \new_[23718]_ ;
  assign \new_[23720]_  = \new_[23719]_  & \new_[23714]_ ;
  assign \new_[23724]_  = A167 & A169;
  assign \new_[23725]_  = ~A170 & \new_[23724]_ ;
  assign \new_[23729]_  = A200 & A199;
  assign \new_[23730]_  = A166 & \new_[23729]_ ;
  assign \new_[23731]_  = \new_[23730]_  & \new_[23725]_ ;
  assign \new_[23735]_  = A234 & ~A233;
  assign \new_[23736]_  = A232 & \new_[23735]_ ;
  assign \new_[23740]_  = A299 & A298;
  assign \new_[23741]_  = A235 & \new_[23740]_ ;
  assign \new_[23742]_  = \new_[23741]_  & \new_[23736]_ ;
  assign \new_[23746]_  = A167 & A169;
  assign \new_[23747]_  = ~A170 & \new_[23746]_ ;
  assign \new_[23751]_  = A200 & A199;
  assign \new_[23752]_  = A166 & \new_[23751]_ ;
  assign \new_[23753]_  = \new_[23752]_  & \new_[23747]_ ;
  assign \new_[23757]_  = A234 & ~A233;
  assign \new_[23758]_  = A232 & \new_[23757]_ ;
  assign \new_[23762]_  = ~A299 & ~A298;
  assign \new_[23763]_  = A235 & \new_[23762]_ ;
  assign \new_[23764]_  = \new_[23763]_  & \new_[23758]_ ;
  assign \new_[23768]_  = A167 & A169;
  assign \new_[23769]_  = ~A170 & \new_[23768]_ ;
  assign \new_[23773]_  = A200 & A199;
  assign \new_[23774]_  = A166 & \new_[23773]_ ;
  assign \new_[23775]_  = \new_[23774]_  & \new_[23769]_ ;
  assign \new_[23779]_  = A234 & ~A233;
  assign \new_[23780]_  = A232 & \new_[23779]_ ;
  assign \new_[23784]_  = A266 & ~A265;
  assign \new_[23785]_  = A235 & \new_[23784]_ ;
  assign \new_[23786]_  = \new_[23785]_  & \new_[23780]_ ;
  assign \new_[23790]_  = A167 & A169;
  assign \new_[23791]_  = ~A170 & \new_[23790]_ ;
  assign \new_[23795]_  = A200 & A199;
  assign \new_[23796]_  = A166 & \new_[23795]_ ;
  assign \new_[23797]_  = \new_[23796]_  & \new_[23791]_ ;
  assign \new_[23801]_  = A234 & ~A233;
  assign \new_[23802]_  = A232 & \new_[23801]_ ;
  assign \new_[23806]_  = ~A300 & A298;
  assign \new_[23807]_  = A236 & \new_[23806]_ ;
  assign \new_[23808]_  = \new_[23807]_  & \new_[23802]_ ;
  assign \new_[23812]_  = A167 & A169;
  assign \new_[23813]_  = ~A170 & \new_[23812]_ ;
  assign \new_[23817]_  = A200 & A199;
  assign \new_[23818]_  = A166 & \new_[23817]_ ;
  assign \new_[23819]_  = \new_[23818]_  & \new_[23813]_ ;
  assign \new_[23823]_  = A234 & ~A233;
  assign \new_[23824]_  = A232 & \new_[23823]_ ;
  assign \new_[23828]_  = A299 & A298;
  assign \new_[23829]_  = A236 & \new_[23828]_ ;
  assign \new_[23830]_  = \new_[23829]_  & \new_[23824]_ ;
  assign \new_[23834]_  = A167 & A169;
  assign \new_[23835]_  = ~A170 & \new_[23834]_ ;
  assign \new_[23839]_  = A200 & A199;
  assign \new_[23840]_  = A166 & \new_[23839]_ ;
  assign \new_[23841]_  = \new_[23840]_  & \new_[23835]_ ;
  assign \new_[23845]_  = A234 & ~A233;
  assign \new_[23846]_  = A232 & \new_[23845]_ ;
  assign \new_[23850]_  = ~A299 & ~A298;
  assign \new_[23851]_  = A236 & \new_[23850]_ ;
  assign \new_[23852]_  = \new_[23851]_  & \new_[23846]_ ;
  assign \new_[23856]_  = A167 & A169;
  assign \new_[23857]_  = ~A170 & \new_[23856]_ ;
  assign \new_[23861]_  = A200 & A199;
  assign \new_[23862]_  = A166 & \new_[23861]_ ;
  assign \new_[23863]_  = \new_[23862]_  & \new_[23857]_ ;
  assign \new_[23867]_  = A234 & ~A233;
  assign \new_[23868]_  = A232 & \new_[23867]_ ;
  assign \new_[23872]_  = A266 & ~A265;
  assign \new_[23873]_  = A236 & \new_[23872]_ ;
  assign \new_[23874]_  = \new_[23873]_  & \new_[23868]_ ;
  assign \new_[23878]_  = A167 & A169;
  assign \new_[23879]_  = ~A170 & \new_[23878]_ ;
  assign \new_[23883]_  = A200 & A199;
  assign \new_[23884]_  = A166 & \new_[23883]_ ;
  assign \new_[23885]_  = \new_[23884]_  & \new_[23879]_ ;
  assign \new_[23889]_  = A265 & ~A233;
  assign \new_[23890]_  = ~A232 & \new_[23889]_ ;
  assign \new_[23894]_  = A299 & ~A298;
  assign \new_[23895]_  = A266 & \new_[23894]_ ;
  assign \new_[23896]_  = \new_[23895]_  & \new_[23890]_ ;
  assign \new_[23900]_  = A167 & A169;
  assign \new_[23901]_  = ~A170 & \new_[23900]_ ;
  assign \new_[23905]_  = A200 & A199;
  assign \new_[23906]_  = A166 & \new_[23905]_ ;
  assign \new_[23907]_  = \new_[23906]_  & \new_[23901]_ ;
  assign \new_[23911]_  = ~A266 & ~A233;
  assign \new_[23912]_  = ~A232 & \new_[23911]_ ;
  assign \new_[23916]_  = A299 & ~A298;
  assign \new_[23917]_  = ~A267 & \new_[23916]_ ;
  assign \new_[23918]_  = \new_[23917]_  & \new_[23912]_ ;
  assign \new_[23922]_  = A167 & A169;
  assign \new_[23923]_  = ~A170 & \new_[23922]_ ;
  assign \new_[23927]_  = A200 & A199;
  assign \new_[23928]_  = A166 & \new_[23927]_ ;
  assign \new_[23929]_  = \new_[23928]_  & \new_[23923]_ ;
  assign \new_[23933]_  = ~A265 & ~A233;
  assign \new_[23934]_  = ~A232 & \new_[23933]_ ;
  assign \new_[23938]_  = A299 & ~A298;
  assign \new_[23939]_  = ~A266 & \new_[23938]_ ;
  assign \new_[23940]_  = \new_[23939]_  & \new_[23934]_ ;
  assign \new_[23944]_  = A167 & A169;
  assign \new_[23945]_  = ~A170 & \new_[23944]_ ;
  assign \new_[23949]_  = ~A202 & ~A200;
  assign \new_[23950]_  = A166 & \new_[23949]_ ;
  assign \new_[23951]_  = \new_[23950]_  & \new_[23945]_ ;
  assign \new_[23955]_  = A233 & ~A232;
  assign \new_[23956]_  = ~A203 & \new_[23955]_ ;
  assign \new_[23960]_  = ~A302 & ~A301;
  assign \new_[23961]_  = ~A299 & \new_[23960]_ ;
  assign \new_[23962]_  = \new_[23961]_  & \new_[23956]_ ;
  assign \new_[23966]_  = A167 & A169;
  assign \new_[23967]_  = ~A170 & \new_[23966]_ ;
  assign \new_[23971]_  = ~A201 & ~A200;
  assign \new_[23972]_  = A166 & \new_[23971]_ ;
  assign \new_[23973]_  = \new_[23972]_  & \new_[23967]_ ;
  assign \new_[23977]_  = A265 & A233;
  assign \new_[23978]_  = A232 & \new_[23977]_ ;
  assign \new_[23982]_  = A299 & ~A298;
  assign \new_[23983]_  = ~A267 & \new_[23982]_ ;
  assign \new_[23984]_  = \new_[23983]_  & \new_[23978]_ ;
  assign \new_[23988]_  = A167 & A169;
  assign \new_[23989]_  = ~A170 & \new_[23988]_ ;
  assign \new_[23993]_  = ~A201 & ~A200;
  assign \new_[23994]_  = A166 & \new_[23993]_ ;
  assign \new_[23995]_  = \new_[23994]_  & \new_[23989]_ ;
  assign \new_[23999]_  = A265 & A233;
  assign \new_[24000]_  = A232 & \new_[23999]_ ;
  assign \new_[24004]_  = A299 & ~A298;
  assign \new_[24005]_  = A266 & \new_[24004]_ ;
  assign \new_[24006]_  = \new_[24005]_  & \new_[24000]_ ;
  assign \new_[24010]_  = A167 & A169;
  assign \new_[24011]_  = ~A170 & \new_[24010]_ ;
  assign \new_[24015]_  = ~A201 & ~A200;
  assign \new_[24016]_  = A166 & \new_[24015]_ ;
  assign \new_[24017]_  = \new_[24016]_  & \new_[24011]_ ;
  assign \new_[24021]_  = ~A265 & A233;
  assign \new_[24022]_  = A232 & \new_[24021]_ ;
  assign \new_[24026]_  = A299 & ~A298;
  assign \new_[24027]_  = ~A266 & \new_[24026]_ ;
  assign \new_[24028]_  = \new_[24027]_  & \new_[24022]_ ;
  assign \new_[24032]_  = A167 & A169;
  assign \new_[24033]_  = ~A170 & \new_[24032]_ ;
  assign \new_[24037]_  = ~A201 & ~A200;
  assign \new_[24038]_  = A166 & \new_[24037]_ ;
  assign \new_[24039]_  = \new_[24038]_  & \new_[24033]_ ;
  assign \new_[24043]_  = A265 & A233;
  assign \new_[24044]_  = ~A232 & \new_[24043]_ ;
  assign \new_[24048]_  = A268 & A267;
  assign \new_[24049]_  = ~A266 & \new_[24048]_ ;
  assign \new_[24050]_  = \new_[24049]_  & \new_[24044]_ ;
  assign \new_[24054]_  = A167 & A169;
  assign \new_[24055]_  = ~A170 & \new_[24054]_ ;
  assign \new_[24059]_  = ~A201 & ~A200;
  assign \new_[24060]_  = A166 & \new_[24059]_ ;
  assign \new_[24061]_  = \new_[24060]_  & \new_[24055]_ ;
  assign \new_[24065]_  = A265 & A233;
  assign \new_[24066]_  = ~A232 & \new_[24065]_ ;
  assign \new_[24070]_  = A269 & A267;
  assign \new_[24071]_  = ~A266 & \new_[24070]_ ;
  assign \new_[24072]_  = \new_[24071]_  & \new_[24066]_ ;
  assign \new_[24076]_  = A167 & A169;
  assign \new_[24077]_  = ~A170 & \new_[24076]_ ;
  assign \new_[24081]_  = ~A201 & ~A200;
  assign \new_[24082]_  = A166 & \new_[24081]_ ;
  assign \new_[24083]_  = \new_[24082]_  & \new_[24077]_ ;
  assign \new_[24087]_  = A265 & ~A234;
  assign \new_[24088]_  = ~A233 & \new_[24087]_ ;
  assign \new_[24092]_  = A299 & ~A298;
  assign \new_[24093]_  = A266 & \new_[24092]_ ;
  assign \new_[24094]_  = \new_[24093]_  & \new_[24088]_ ;
  assign \new_[24098]_  = A167 & A169;
  assign \new_[24099]_  = ~A170 & \new_[24098]_ ;
  assign \new_[24103]_  = ~A201 & ~A200;
  assign \new_[24104]_  = A166 & \new_[24103]_ ;
  assign \new_[24105]_  = \new_[24104]_  & \new_[24099]_ ;
  assign \new_[24109]_  = ~A266 & ~A234;
  assign \new_[24110]_  = ~A233 & \new_[24109]_ ;
  assign \new_[24114]_  = A299 & ~A298;
  assign \new_[24115]_  = ~A267 & \new_[24114]_ ;
  assign \new_[24116]_  = \new_[24115]_  & \new_[24110]_ ;
  assign \new_[24120]_  = A167 & A169;
  assign \new_[24121]_  = ~A170 & \new_[24120]_ ;
  assign \new_[24125]_  = ~A201 & ~A200;
  assign \new_[24126]_  = A166 & \new_[24125]_ ;
  assign \new_[24127]_  = \new_[24126]_  & \new_[24121]_ ;
  assign \new_[24131]_  = ~A265 & ~A234;
  assign \new_[24132]_  = ~A233 & \new_[24131]_ ;
  assign \new_[24136]_  = A299 & ~A298;
  assign \new_[24137]_  = ~A266 & \new_[24136]_ ;
  assign \new_[24138]_  = \new_[24137]_  & \new_[24132]_ ;
  assign \new_[24142]_  = A167 & A169;
  assign \new_[24143]_  = ~A170 & \new_[24142]_ ;
  assign \new_[24147]_  = ~A201 & ~A200;
  assign \new_[24148]_  = A166 & \new_[24147]_ ;
  assign \new_[24149]_  = \new_[24148]_  & \new_[24143]_ ;
  assign \new_[24153]_  = A234 & ~A233;
  assign \new_[24154]_  = A232 & \new_[24153]_ ;
  assign \new_[24158]_  = ~A300 & A298;
  assign \new_[24159]_  = A235 & \new_[24158]_ ;
  assign \new_[24160]_  = \new_[24159]_  & \new_[24154]_ ;
  assign \new_[24164]_  = A167 & A169;
  assign \new_[24165]_  = ~A170 & \new_[24164]_ ;
  assign \new_[24169]_  = ~A201 & ~A200;
  assign \new_[24170]_  = A166 & \new_[24169]_ ;
  assign \new_[24171]_  = \new_[24170]_  & \new_[24165]_ ;
  assign \new_[24175]_  = A234 & ~A233;
  assign \new_[24176]_  = A232 & \new_[24175]_ ;
  assign \new_[24180]_  = A299 & A298;
  assign \new_[24181]_  = A235 & \new_[24180]_ ;
  assign \new_[24182]_  = \new_[24181]_  & \new_[24176]_ ;
  assign \new_[24186]_  = A167 & A169;
  assign \new_[24187]_  = ~A170 & \new_[24186]_ ;
  assign \new_[24191]_  = ~A201 & ~A200;
  assign \new_[24192]_  = A166 & \new_[24191]_ ;
  assign \new_[24193]_  = \new_[24192]_  & \new_[24187]_ ;
  assign \new_[24197]_  = A234 & ~A233;
  assign \new_[24198]_  = A232 & \new_[24197]_ ;
  assign \new_[24202]_  = ~A299 & ~A298;
  assign \new_[24203]_  = A235 & \new_[24202]_ ;
  assign \new_[24204]_  = \new_[24203]_  & \new_[24198]_ ;
  assign \new_[24208]_  = A167 & A169;
  assign \new_[24209]_  = ~A170 & \new_[24208]_ ;
  assign \new_[24213]_  = ~A201 & ~A200;
  assign \new_[24214]_  = A166 & \new_[24213]_ ;
  assign \new_[24215]_  = \new_[24214]_  & \new_[24209]_ ;
  assign \new_[24219]_  = A234 & ~A233;
  assign \new_[24220]_  = A232 & \new_[24219]_ ;
  assign \new_[24224]_  = A266 & ~A265;
  assign \new_[24225]_  = A235 & \new_[24224]_ ;
  assign \new_[24226]_  = \new_[24225]_  & \new_[24220]_ ;
  assign \new_[24230]_  = A167 & A169;
  assign \new_[24231]_  = ~A170 & \new_[24230]_ ;
  assign \new_[24235]_  = ~A201 & ~A200;
  assign \new_[24236]_  = A166 & \new_[24235]_ ;
  assign \new_[24237]_  = \new_[24236]_  & \new_[24231]_ ;
  assign \new_[24241]_  = A234 & ~A233;
  assign \new_[24242]_  = A232 & \new_[24241]_ ;
  assign \new_[24246]_  = ~A300 & A298;
  assign \new_[24247]_  = A236 & \new_[24246]_ ;
  assign \new_[24248]_  = \new_[24247]_  & \new_[24242]_ ;
  assign \new_[24252]_  = A167 & A169;
  assign \new_[24253]_  = ~A170 & \new_[24252]_ ;
  assign \new_[24257]_  = ~A201 & ~A200;
  assign \new_[24258]_  = A166 & \new_[24257]_ ;
  assign \new_[24259]_  = \new_[24258]_  & \new_[24253]_ ;
  assign \new_[24263]_  = A234 & ~A233;
  assign \new_[24264]_  = A232 & \new_[24263]_ ;
  assign \new_[24268]_  = A299 & A298;
  assign \new_[24269]_  = A236 & \new_[24268]_ ;
  assign \new_[24270]_  = \new_[24269]_  & \new_[24264]_ ;
  assign \new_[24274]_  = A167 & A169;
  assign \new_[24275]_  = ~A170 & \new_[24274]_ ;
  assign \new_[24279]_  = ~A201 & ~A200;
  assign \new_[24280]_  = A166 & \new_[24279]_ ;
  assign \new_[24281]_  = \new_[24280]_  & \new_[24275]_ ;
  assign \new_[24285]_  = A234 & ~A233;
  assign \new_[24286]_  = A232 & \new_[24285]_ ;
  assign \new_[24290]_  = ~A299 & ~A298;
  assign \new_[24291]_  = A236 & \new_[24290]_ ;
  assign \new_[24292]_  = \new_[24291]_  & \new_[24286]_ ;
  assign \new_[24296]_  = A167 & A169;
  assign \new_[24297]_  = ~A170 & \new_[24296]_ ;
  assign \new_[24301]_  = ~A201 & ~A200;
  assign \new_[24302]_  = A166 & \new_[24301]_ ;
  assign \new_[24303]_  = \new_[24302]_  & \new_[24297]_ ;
  assign \new_[24307]_  = A234 & ~A233;
  assign \new_[24308]_  = A232 & \new_[24307]_ ;
  assign \new_[24312]_  = A266 & ~A265;
  assign \new_[24313]_  = A236 & \new_[24312]_ ;
  assign \new_[24314]_  = \new_[24313]_  & \new_[24308]_ ;
  assign \new_[24318]_  = A167 & A169;
  assign \new_[24319]_  = ~A170 & \new_[24318]_ ;
  assign \new_[24323]_  = ~A201 & ~A200;
  assign \new_[24324]_  = A166 & \new_[24323]_ ;
  assign \new_[24325]_  = \new_[24324]_  & \new_[24319]_ ;
  assign \new_[24329]_  = A265 & ~A233;
  assign \new_[24330]_  = ~A232 & \new_[24329]_ ;
  assign \new_[24334]_  = A299 & ~A298;
  assign \new_[24335]_  = A266 & \new_[24334]_ ;
  assign \new_[24336]_  = \new_[24335]_  & \new_[24330]_ ;
  assign \new_[24340]_  = A167 & A169;
  assign \new_[24341]_  = ~A170 & \new_[24340]_ ;
  assign \new_[24345]_  = ~A201 & ~A200;
  assign \new_[24346]_  = A166 & \new_[24345]_ ;
  assign \new_[24347]_  = \new_[24346]_  & \new_[24341]_ ;
  assign \new_[24351]_  = ~A266 & ~A233;
  assign \new_[24352]_  = ~A232 & \new_[24351]_ ;
  assign \new_[24356]_  = A299 & ~A298;
  assign \new_[24357]_  = ~A267 & \new_[24356]_ ;
  assign \new_[24358]_  = \new_[24357]_  & \new_[24352]_ ;
  assign \new_[24362]_  = A167 & A169;
  assign \new_[24363]_  = ~A170 & \new_[24362]_ ;
  assign \new_[24367]_  = ~A201 & ~A200;
  assign \new_[24368]_  = A166 & \new_[24367]_ ;
  assign \new_[24369]_  = \new_[24368]_  & \new_[24363]_ ;
  assign \new_[24373]_  = ~A265 & ~A233;
  assign \new_[24374]_  = ~A232 & \new_[24373]_ ;
  assign \new_[24378]_  = A299 & ~A298;
  assign \new_[24379]_  = ~A266 & \new_[24378]_ ;
  assign \new_[24380]_  = \new_[24379]_  & \new_[24374]_ ;
  assign \new_[24384]_  = A167 & A169;
  assign \new_[24385]_  = ~A170 & \new_[24384]_ ;
  assign \new_[24389]_  = ~A200 & ~A199;
  assign \new_[24390]_  = A166 & \new_[24389]_ ;
  assign \new_[24391]_  = \new_[24390]_  & \new_[24385]_ ;
  assign \new_[24395]_  = A265 & A233;
  assign \new_[24396]_  = A232 & \new_[24395]_ ;
  assign \new_[24400]_  = A299 & ~A298;
  assign \new_[24401]_  = ~A267 & \new_[24400]_ ;
  assign \new_[24402]_  = \new_[24401]_  & \new_[24396]_ ;
  assign \new_[24406]_  = A167 & A169;
  assign \new_[24407]_  = ~A170 & \new_[24406]_ ;
  assign \new_[24411]_  = ~A200 & ~A199;
  assign \new_[24412]_  = A166 & \new_[24411]_ ;
  assign \new_[24413]_  = \new_[24412]_  & \new_[24407]_ ;
  assign \new_[24417]_  = A265 & A233;
  assign \new_[24418]_  = A232 & \new_[24417]_ ;
  assign \new_[24422]_  = A299 & ~A298;
  assign \new_[24423]_  = A266 & \new_[24422]_ ;
  assign \new_[24424]_  = \new_[24423]_  & \new_[24418]_ ;
  assign \new_[24428]_  = A167 & A169;
  assign \new_[24429]_  = ~A170 & \new_[24428]_ ;
  assign \new_[24433]_  = ~A200 & ~A199;
  assign \new_[24434]_  = A166 & \new_[24433]_ ;
  assign \new_[24435]_  = \new_[24434]_  & \new_[24429]_ ;
  assign \new_[24439]_  = ~A265 & A233;
  assign \new_[24440]_  = A232 & \new_[24439]_ ;
  assign \new_[24444]_  = A299 & ~A298;
  assign \new_[24445]_  = ~A266 & \new_[24444]_ ;
  assign \new_[24446]_  = \new_[24445]_  & \new_[24440]_ ;
  assign \new_[24450]_  = A167 & A169;
  assign \new_[24451]_  = ~A170 & \new_[24450]_ ;
  assign \new_[24455]_  = ~A200 & ~A199;
  assign \new_[24456]_  = A166 & \new_[24455]_ ;
  assign \new_[24457]_  = \new_[24456]_  & \new_[24451]_ ;
  assign \new_[24461]_  = A265 & A233;
  assign \new_[24462]_  = ~A232 & \new_[24461]_ ;
  assign \new_[24466]_  = A268 & A267;
  assign \new_[24467]_  = ~A266 & \new_[24466]_ ;
  assign \new_[24468]_  = \new_[24467]_  & \new_[24462]_ ;
  assign \new_[24472]_  = A167 & A169;
  assign \new_[24473]_  = ~A170 & \new_[24472]_ ;
  assign \new_[24477]_  = ~A200 & ~A199;
  assign \new_[24478]_  = A166 & \new_[24477]_ ;
  assign \new_[24479]_  = \new_[24478]_  & \new_[24473]_ ;
  assign \new_[24483]_  = A265 & A233;
  assign \new_[24484]_  = ~A232 & \new_[24483]_ ;
  assign \new_[24488]_  = A269 & A267;
  assign \new_[24489]_  = ~A266 & \new_[24488]_ ;
  assign \new_[24490]_  = \new_[24489]_  & \new_[24484]_ ;
  assign \new_[24494]_  = A167 & A169;
  assign \new_[24495]_  = ~A170 & \new_[24494]_ ;
  assign \new_[24499]_  = ~A200 & ~A199;
  assign \new_[24500]_  = A166 & \new_[24499]_ ;
  assign \new_[24501]_  = \new_[24500]_  & \new_[24495]_ ;
  assign \new_[24505]_  = A265 & ~A234;
  assign \new_[24506]_  = ~A233 & \new_[24505]_ ;
  assign \new_[24510]_  = A299 & ~A298;
  assign \new_[24511]_  = A266 & \new_[24510]_ ;
  assign \new_[24512]_  = \new_[24511]_  & \new_[24506]_ ;
  assign \new_[24516]_  = A167 & A169;
  assign \new_[24517]_  = ~A170 & \new_[24516]_ ;
  assign \new_[24521]_  = ~A200 & ~A199;
  assign \new_[24522]_  = A166 & \new_[24521]_ ;
  assign \new_[24523]_  = \new_[24522]_  & \new_[24517]_ ;
  assign \new_[24527]_  = ~A266 & ~A234;
  assign \new_[24528]_  = ~A233 & \new_[24527]_ ;
  assign \new_[24532]_  = A299 & ~A298;
  assign \new_[24533]_  = ~A267 & \new_[24532]_ ;
  assign \new_[24534]_  = \new_[24533]_  & \new_[24528]_ ;
  assign \new_[24538]_  = A167 & A169;
  assign \new_[24539]_  = ~A170 & \new_[24538]_ ;
  assign \new_[24543]_  = ~A200 & ~A199;
  assign \new_[24544]_  = A166 & \new_[24543]_ ;
  assign \new_[24545]_  = \new_[24544]_  & \new_[24539]_ ;
  assign \new_[24549]_  = ~A265 & ~A234;
  assign \new_[24550]_  = ~A233 & \new_[24549]_ ;
  assign \new_[24554]_  = A299 & ~A298;
  assign \new_[24555]_  = ~A266 & \new_[24554]_ ;
  assign \new_[24556]_  = \new_[24555]_  & \new_[24550]_ ;
  assign \new_[24560]_  = A167 & A169;
  assign \new_[24561]_  = ~A170 & \new_[24560]_ ;
  assign \new_[24565]_  = ~A200 & ~A199;
  assign \new_[24566]_  = A166 & \new_[24565]_ ;
  assign \new_[24567]_  = \new_[24566]_  & \new_[24561]_ ;
  assign \new_[24571]_  = A234 & ~A233;
  assign \new_[24572]_  = A232 & \new_[24571]_ ;
  assign \new_[24576]_  = ~A300 & A298;
  assign \new_[24577]_  = A235 & \new_[24576]_ ;
  assign \new_[24578]_  = \new_[24577]_  & \new_[24572]_ ;
  assign \new_[24582]_  = A167 & A169;
  assign \new_[24583]_  = ~A170 & \new_[24582]_ ;
  assign \new_[24587]_  = ~A200 & ~A199;
  assign \new_[24588]_  = A166 & \new_[24587]_ ;
  assign \new_[24589]_  = \new_[24588]_  & \new_[24583]_ ;
  assign \new_[24593]_  = A234 & ~A233;
  assign \new_[24594]_  = A232 & \new_[24593]_ ;
  assign \new_[24598]_  = A299 & A298;
  assign \new_[24599]_  = A235 & \new_[24598]_ ;
  assign \new_[24600]_  = \new_[24599]_  & \new_[24594]_ ;
  assign \new_[24604]_  = A167 & A169;
  assign \new_[24605]_  = ~A170 & \new_[24604]_ ;
  assign \new_[24609]_  = ~A200 & ~A199;
  assign \new_[24610]_  = A166 & \new_[24609]_ ;
  assign \new_[24611]_  = \new_[24610]_  & \new_[24605]_ ;
  assign \new_[24615]_  = A234 & ~A233;
  assign \new_[24616]_  = A232 & \new_[24615]_ ;
  assign \new_[24620]_  = ~A299 & ~A298;
  assign \new_[24621]_  = A235 & \new_[24620]_ ;
  assign \new_[24622]_  = \new_[24621]_  & \new_[24616]_ ;
  assign \new_[24626]_  = A167 & A169;
  assign \new_[24627]_  = ~A170 & \new_[24626]_ ;
  assign \new_[24631]_  = ~A200 & ~A199;
  assign \new_[24632]_  = A166 & \new_[24631]_ ;
  assign \new_[24633]_  = \new_[24632]_  & \new_[24627]_ ;
  assign \new_[24637]_  = A234 & ~A233;
  assign \new_[24638]_  = A232 & \new_[24637]_ ;
  assign \new_[24642]_  = A266 & ~A265;
  assign \new_[24643]_  = A235 & \new_[24642]_ ;
  assign \new_[24644]_  = \new_[24643]_  & \new_[24638]_ ;
  assign \new_[24648]_  = A167 & A169;
  assign \new_[24649]_  = ~A170 & \new_[24648]_ ;
  assign \new_[24653]_  = ~A200 & ~A199;
  assign \new_[24654]_  = A166 & \new_[24653]_ ;
  assign \new_[24655]_  = \new_[24654]_  & \new_[24649]_ ;
  assign \new_[24659]_  = A234 & ~A233;
  assign \new_[24660]_  = A232 & \new_[24659]_ ;
  assign \new_[24664]_  = ~A300 & A298;
  assign \new_[24665]_  = A236 & \new_[24664]_ ;
  assign \new_[24666]_  = \new_[24665]_  & \new_[24660]_ ;
  assign \new_[24670]_  = A167 & A169;
  assign \new_[24671]_  = ~A170 & \new_[24670]_ ;
  assign \new_[24675]_  = ~A200 & ~A199;
  assign \new_[24676]_  = A166 & \new_[24675]_ ;
  assign \new_[24677]_  = \new_[24676]_  & \new_[24671]_ ;
  assign \new_[24681]_  = A234 & ~A233;
  assign \new_[24682]_  = A232 & \new_[24681]_ ;
  assign \new_[24686]_  = A299 & A298;
  assign \new_[24687]_  = A236 & \new_[24686]_ ;
  assign \new_[24688]_  = \new_[24687]_  & \new_[24682]_ ;
  assign \new_[24692]_  = A167 & A169;
  assign \new_[24693]_  = ~A170 & \new_[24692]_ ;
  assign \new_[24697]_  = ~A200 & ~A199;
  assign \new_[24698]_  = A166 & \new_[24697]_ ;
  assign \new_[24699]_  = \new_[24698]_  & \new_[24693]_ ;
  assign \new_[24703]_  = A234 & ~A233;
  assign \new_[24704]_  = A232 & \new_[24703]_ ;
  assign \new_[24708]_  = ~A299 & ~A298;
  assign \new_[24709]_  = A236 & \new_[24708]_ ;
  assign \new_[24710]_  = \new_[24709]_  & \new_[24704]_ ;
  assign \new_[24714]_  = A167 & A169;
  assign \new_[24715]_  = ~A170 & \new_[24714]_ ;
  assign \new_[24719]_  = ~A200 & ~A199;
  assign \new_[24720]_  = A166 & \new_[24719]_ ;
  assign \new_[24721]_  = \new_[24720]_  & \new_[24715]_ ;
  assign \new_[24725]_  = A234 & ~A233;
  assign \new_[24726]_  = A232 & \new_[24725]_ ;
  assign \new_[24730]_  = A266 & ~A265;
  assign \new_[24731]_  = A236 & \new_[24730]_ ;
  assign \new_[24732]_  = \new_[24731]_  & \new_[24726]_ ;
  assign \new_[24736]_  = A167 & A169;
  assign \new_[24737]_  = ~A170 & \new_[24736]_ ;
  assign \new_[24741]_  = ~A200 & ~A199;
  assign \new_[24742]_  = A166 & \new_[24741]_ ;
  assign \new_[24743]_  = \new_[24742]_  & \new_[24737]_ ;
  assign \new_[24747]_  = A265 & ~A233;
  assign \new_[24748]_  = ~A232 & \new_[24747]_ ;
  assign \new_[24752]_  = A299 & ~A298;
  assign \new_[24753]_  = A266 & \new_[24752]_ ;
  assign \new_[24754]_  = \new_[24753]_  & \new_[24748]_ ;
  assign \new_[24758]_  = A167 & A169;
  assign \new_[24759]_  = ~A170 & \new_[24758]_ ;
  assign \new_[24763]_  = ~A200 & ~A199;
  assign \new_[24764]_  = A166 & \new_[24763]_ ;
  assign \new_[24765]_  = \new_[24764]_  & \new_[24759]_ ;
  assign \new_[24769]_  = ~A266 & ~A233;
  assign \new_[24770]_  = ~A232 & \new_[24769]_ ;
  assign \new_[24774]_  = A299 & ~A298;
  assign \new_[24775]_  = ~A267 & \new_[24774]_ ;
  assign \new_[24776]_  = \new_[24775]_  & \new_[24770]_ ;
  assign \new_[24780]_  = A167 & A169;
  assign \new_[24781]_  = ~A170 & \new_[24780]_ ;
  assign \new_[24785]_  = ~A200 & ~A199;
  assign \new_[24786]_  = A166 & \new_[24785]_ ;
  assign \new_[24787]_  = \new_[24786]_  & \new_[24781]_ ;
  assign \new_[24791]_  = ~A265 & ~A233;
  assign \new_[24792]_  = ~A232 & \new_[24791]_ ;
  assign \new_[24796]_  = A299 & ~A298;
  assign \new_[24797]_  = ~A266 & \new_[24796]_ ;
  assign \new_[24798]_  = \new_[24797]_  & \new_[24792]_ ;
  assign \new_[24802]_  = ~A167 & A169;
  assign \new_[24803]_  = ~A170 & \new_[24802]_ ;
  assign \new_[24807]_  = A200 & A199;
  assign \new_[24808]_  = ~A166 & \new_[24807]_ ;
  assign \new_[24809]_  = \new_[24808]_  & \new_[24803]_ ;
  assign \new_[24813]_  = A265 & A233;
  assign \new_[24814]_  = A232 & \new_[24813]_ ;
  assign \new_[24818]_  = A299 & ~A298;
  assign \new_[24819]_  = ~A267 & \new_[24818]_ ;
  assign \new_[24820]_  = \new_[24819]_  & \new_[24814]_ ;
  assign \new_[24824]_  = ~A167 & A169;
  assign \new_[24825]_  = ~A170 & \new_[24824]_ ;
  assign \new_[24829]_  = A200 & A199;
  assign \new_[24830]_  = ~A166 & \new_[24829]_ ;
  assign \new_[24831]_  = \new_[24830]_  & \new_[24825]_ ;
  assign \new_[24835]_  = A265 & A233;
  assign \new_[24836]_  = A232 & \new_[24835]_ ;
  assign \new_[24840]_  = A299 & ~A298;
  assign \new_[24841]_  = A266 & \new_[24840]_ ;
  assign \new_[24842]_  = \new_[24841]_  & \new_[24836]_ ;
  assign \new_[24846]_  = ~A167 & A169;
  assign \new_[24847]_  = ~A170 & \new_[24846]_ ;
  assign \new_[24851]_  = A200 & A199;
  assign \new_[24852]_  = ~A166 & \new_[24851]_ ;
  assign \new_[24853]_  = \new_[24852]_  & \new_[24847]_ ;
  assign \new_[24857]_  = ~A265 & A233;
  assign \new_[24858]_  = A232 & \new_[24857]_ ;
  assign \new_[24862]_  = A299 & ~A298;
  assign \new_[24863]_  = ~A266 & \new_[24862]_ ;
  assign \new_[24864]_  = \new_[24863]_  & \new_[24858]_ ;
  assign \new_[24868]_  = ~A167 & A169;
  assign \new_[24869]_  = ~A170 & \new_[24868]_ ;
  assign \new_[24873]_  = A200 & A199;
  assign \new_[24874]_  = ~A166 & \new_[24873]_ ;
  assign \new_[24875]_  = \new_[24874]_  & \new_[24869]_ ;
  assign \new_[24879]_  = A265 & A233;
  assign \new_[24880]_  = ~A232 & \new_[24879]_ ;
  assign \new_[24884]_  = A268 & A267;
  assign \new_[24885]_  = ~A266 & \new_[24884]_ ;
  assign \new_[24886]_  = \new_[24885]_  & \new_[24880]_ ;
  assign \new_[24890]_  = ~A167 & A169;
  assign \new_[24891]_  = ~A170 & \new_[24890]_ ;
  assign \new_[24895]_  = A200 & A199;
  assign \new_[24896]_  = ~A166 & \new_[24895]_ ;
  assign \new_[24897]_  = \new_[24896]_  & \new_[24891]_ ;
  assign \new_[24901]_  = A265 & A233;
  assign \new_[24902]_  = ~A232 & \new_[24901]_ ;
  assign \new_[24906]_  = A269 & A267;
  assign \new_[24907]_  = ~A266 & \new_[24906]_ ;
  assign \new_[24908]_  = \new_[24907]_  & \new_[24902]_ ;
  assign \new_[24912]_  = ~A167 & A169;
  assign \new_[24913]_  = ~A170 & \new_[24912]_ ;
  assign \new_[24917]_  = A200 & A199;
  assign \new_[24918]_  = ~A166 & \new_[24917]_ ;
  assign \new_[24919]_  = \new_[24918]_  & \new_[24913]_ ;
  assign \new_[24923]_  = A265 & ~A234;
  assign \new_[24924]_  = ~A233 & \new_[24923]_ ;
  assign \new_[24928]_  = A299 & ~A298;
  assign \new_[24929]_  = A266 & \new_[24928]_ ;
  assign \new_[24930]_  = \new_[24929]_  & \new_[24924]_ ;
  assign \new_[24934]_  = ~A167 & A169;
  assign \new_[24935]_  = ~A170 & \new_[24934]_ ;
  assign \new_[24939]_  = A200 & A199;
  assign \new_[24940]_  = ~A166 & \new_[24939]_ ;
  assign \new_[24941]_  = \new_[24940]_  & \new_[24935]_ ;
  assign \new_[24945]_  = ~A266 & ~A234;
  assign \new_[24946]_  = ~A233 & \new_[24945]_ ;
  assign \new_[24950]_  = A299 & ~A298;
  assign \new_[24951]_  = ~A267 & \new_[24950]_ ;
  assign \new_[24952]_  = \new_[24951]_  & \new_[24946]_ ;
  assign \new_[24956]_  = ~A167 & A169;
  assign \new_[24957]_  = ~A170 & \new_[24956]_ ;
  assign \new_[24961]_  = A200 & A199;
  assign \new_[24962]_  = ~A166 & \new_[24961]_ ;
  assign \new_[24963]_  = \new_[24962]_  & \new_[24957]_ ;
  assign \new_[24967]_  = ~A265 & ~A234;
  assign \new_[24968]_  = ~A233 & \new_[24967]_ ;
  assign \new_[24972]_  = A299 & ~A298;
  assign \new_[24973]_  = ~A266 & \new_[24972]_ ;
  assign \new_[24974]_  = \new_[24973]_  & \new_[24968]_ ;
  assign \new_[24978]_  = ~A167 & A169;
  assign \new_[24979]_  = ~A170 & \new_[24978]_ ;
  assign \new_[24983]_  = A200 & A199;
  assign \new_[24984]_  = ~A166 & \new_[24983]_ ;
  assign \new_[24985]_  = \new_[24984]_  & \new_[24979]_ ;
  assign \new_[24989]_  = A234 & ~A233;
  assign \new_[24990]_  = A232 & \new_[24989]_ ;
  assign \new_[24994]_  = ~A300 & A298;
  assign \new_[24995]_  = A235 & \new_[24994]_ ;
  assign \new_[24996]_  = \new_[24995]_  & \new_[24990]_ ;
  assign \new_[25000]_  = ~A167 & A169;
  assign \new_[25001]_  = ~A170 & \new_[25000]_ ;
  assign \new_[25005]_  = A200 & A199;
  assign \new_[25006]_  = ~A166 & \new_[25005]_ ;
  assign \new_[25007]_  = \new_[25006]_  & \new_[25001]_ ;
  assign \new_[25011]_  = A234 & ~A233;
  assign \new_[25012]_  = A232 & \new_[25011]_ ;
  assign \new_[25016]_  = A299 & A298;
  assign \new_[25017]_  = A235 & \new_[25016]_ ;
  assign \new_[25018]_  = \new_[25017]_  & \new_[25012]_ ;
  assign \new_[25022]_  = ~A167 & A169;
  assign \new_[25023]_  = ~A170 & \new_[25022]_ ;
  assign \new_[25027]_  = A200 & A199;
  assign \new_[25028]_  = ~A166 & \new_[25027]_ ;
  assign \new_[25029]_  = \new_[25028]_  & \new_[25023]_ ;
  assign \new_[25033]_  = A234 & ~A233;
  assign \new_[25034]_  = A232 & \new_[25033]_ ;
  assign \new_[25038]_  = ~A299 & ~A298;
  assign \new_[25039]_  = A235 & \new_[25038]_ ;
  assign \new_[25040]_  = \new_[25039]_  & \new_[25034]_ ;
  assign \new_[25044]_  = ~A167 & A169;
  assign \new_[25045]_  = ~A170 & \new_[25044]_ ;
  assign \new_[25049]_  = A200 & A199;
  assign \new_[25050]_  = ~A166 & \new_[25049]_ ;
  assign \new_[25051]_  = \new_[25050]_  & \new_[25045]_ ;
  assign \new_[25055]_  = A234 & ~A233;
  assign \new_[25056]_  = A232 & \new_[25055]_ ;
  assign \new_[25060]_  = A266 & ~A265;
  assign \new_[25061]_  = A235 & \new_[25060]_ ;
  assign \new_[25062]_  = \new_[25061]_  & \new_[25056]_ ;
  assign \new_[25066]_  = ~A167 & A169;
  assign \new_[25067]_  = ~A170 & \new_[25066]_ ;
  assign \new_[25071]_  = A200 & A199;
  assign \new_[25072]_  = ~A166 & \new_[25071]_ ;
  assign \new_[25073]_  = \new_[25072]_  & \new_[25067]_ ;
  assign \new_[25077]_  = A234 & ~A233;
  assign \new_[25078]_  = A232 & \new_[25077]_ ;
  assign \new_[25082]_  = ~A300 & A298;
  assign \new_[25083]_  = A236 & \new_[25082]_ ;
  assign \new_[25084]_  = \new_[25083]_  & \new_[25078]_ ;
  assign \new_[25088]_  = ~A167 & A169;
  assign \new_[25089]_  = ~A170 & \new_[25088]_ ;
  assign \new_[25093]_  = A200 & A199;
  assign \new_[25094]_  = ~A166 & \new_[25093]_ ;
  assign \new_[25095]_  = \new_[25094]_  & \new_[25089]_ ;
  assign \new_[25099]_  = A234 & ~A233;
  assign \new_[25100]_  = A232 & \new_[25099]_ ;
  assign \new_[25104]_  = A299 & A298;
  assign \new_[25105]_  = A236 & \new_[25104]_ ;
  assign \new_[25106]_  = \new_[25105]_  & \new_[25100]_ ;
  assign \new_[25110]_  = ~A167 & A169;
  assign \new_[25111]_  = ~A170 & \new_[25110]_ ;
  assign \new_[25115]_  = A200 & A199;
  assign \new_[25116]_  = ~A166 & \new_[25115]_ ;
  assign \new_[25117]_  = \new_[25116]_  & \new_[25111]_ ;
  assign \new_[25121]_  = A234 & ~A233;
  assign \new_[25122]_  = A232 & \new_[25121]_ ;
  assign \new_[25126]_  = ~A299 & ~A298;
  assign \new_[25127]_  = A236 & \new_[25126]_ ;
  assign \new_[25128]_  = \new_[25127]_  & \new_[25122]_ ;
  assign \new_[25132]_  = ~A167 & A169;
  assign \new_[25133]_  = ~A170 & \new_[25132]_ ;
  assign \new_[25137]_  = A200 & A199;
  assign \new_[25138]_  = ~A166 & \new_[25137]_ ;
  assign \new_[25139]_  = \new_[25138]_  & \new_[25133]_ ;
  assign \new_[25143]_  = A234 & ~A233;
  assign \new_[25144]_  = A232 & \new_[25143]_ ;
  assign \new_[25148]_  = A266 & ~A265;
  assign \new_[25149]_  = A236 & \new_[25148]_ ;
  assign \new_[25150]_  = \new_[25149]_  & \new_[25144]_ ;
  assign \new_[25154]_  = ~A167 & A169;
  assign \new_[25155]_  = ~A170 & \new_[25154]_ ;
  assign \new_[25159]_  = A200 & A199;
  assign \new_[25160]_  = ~A166 & \new_[25159]_ ;
  assign \new_[25161]_  = \new_[25160]_  & \new_[25155]_ ;
  assign \new_[25165]_  = A265 & ~A233;
  assign \new_[25166]_  = ~A232 & \new_[25165]_ ;
  assign \new_[25170]_  = A299 & ~A298;
  assign \new_[25171]_  = A266 & \new_[25170]_ ;
  assign \new_[25172]_  = \new_[25171]_  & \new_[25166]_ ;
  assign \new_[25176]_  = ~A167 & A169;
  assign \new_[25177]_  = ~A170 & \new_[25176]_ ;
  assign \new_[25181]_  = A200 & A199;
  assign \new_[25182]_  = ~A166 & \new_[25181]_ ;
  assign \new_[25183]_  = \new_[25182]_  & \new_[25177]_ ;
  assign \new_[25187]_  = ~A266 & ~A233;
  assign \new_[25188]_  = ~A232 & \new_[25187]_ ;
  assign \new_[25192]_  = A299 & ~A298;
  assign \new_[25193]_  = ~A267 & \new_[25192]_ ;
  assign \new_[25194]_  = \new_[25193]_  & \new_[25188]_ ;
  assign \new_[25198]_  = ~A167 & A169;
  assign \new_[25199]_  = ~A170 & \new_[25198]_ ;
  assign \new_[25203]_  = A200 & A199;
  assign \new_[25204]_  = ~A166 & \new_[25203]_ ;
  assign \new_[25205]_  = \new_[25204]_  & \new_[25199]_ ;
  assign \new_[25209]_  = ~A265 & ~A233;
  assign \new_[25210]_  = ~A232 & \new_[25209]_ ;
  assign \new_[25214]_  = A299 & ~A298;
  assign \new_[25215]_  = ~A266 & \new_[25214]_ ;
  assign \new_[25216]_  = \new_[25215]_  & \new_[25210]_ ;
  assign \new_[25220]_  = ~A167 & A169;
  assign \new_[25221]_  = ~A170 & \new_[25220]_ ;
  assign \new_[25225]_  = ~A202 & ~A200;
  assign \new_[25226]_  = ~A166 & \new_[25225]_ ;
  assign \new_[25227]_  = \new_[25226]_  & \new_[25221]_ ;
  assign \new_[25231]_  = A233 & ~A232;
  assign \new_[25232]_  = ~A203 & \new_[25231]_ ;
  assign \new_[25236]_  = ~A302 & ~A301;
  assign \new_[25237]_  = ~A299 & \new_[25236]_ ;
  assign \new_[25238]_  = \new_[25237]_  & \new_[25232]_ ;
  assign \new_[25242]_  = ~A167 & A169;
  assign \new_[25243]_  = ~A170 & \new_[25242]_ ;
  assign \new_[25247]_  = ~A201 & ~A200;
  assign \new_[25248]_  = ~A166 & \new_[25247]_ ;
  assign \new_[25249]_  = \new_[25248]_  & \new_[25243]_ ;
  assign \new_[25253]_  = A265 & A233;
  assign \new_[25254]_  = A232 & \new_[25253]_ ;
  assign \new_[25258]_  = A299 & ~A298;
  assign \new_[25259]_  = ~A267 & \new_[25258]_ ;
  assign \new_[25260]_  = \new_[25259]_  & \new_[25254]_ ;
  assign \new_[25264]_  = ~A167 & A169;
  assign \new_[25265]_  = ~A170 & \new_[25264]_ ;
  assign \new_[25269]_  = ~A201 & ~A200;
  assign \new_[25270]_  = ~A166 & \new_[25269]_ ;
  assign \new_[25271]_  = \new_[25270]_  & \new_[25265]_ ;
  assign \new_[25275]_  = A265 & A233;
  assign \new_[25276]_  = A232 & \new_[25275]_ ;
  assign \new_[25280]_  = A299 & ~A298;
  assign \new_[25281]_  = A266 & \new_[25280]_ ;
  assign \new_[25282]_  = \new_[25281]_  & \new_[25276]_ ;
  assign \new_[25286]_  = ~A167 & A169;
  assign \new_[25287]_  = ~A170 & \new_[25286]_ ;
  assign \new_[25291]_  = ~A201 & ~A200;
  assign \new_[25292]_  = ~A166 & \new_[25291]_ ;
  assign \new_[25293]_  = \new_[25292]_  & \new_[25287]_ ;
  assign \new_[25297]_  = ~A265 & A233;
  assign \new_[25298]_  = A232 & \new_[25297]_ ;
  assign \new_[25302]_  = A299 & ~A298;
  assign \new_[25303]_  = ~A266 & \new_[25302]_ ;
  assign \new_[25304]_  = \new_[25303]_  & \new_[25298]_ ;
  assign \new_[25308]_  = ~A167 & A169;
  assign \new_[25309]_  = ~A170 & \new_[25308]_ ;
  assign \new_[25313]_  = ~A201 & ~A200;
  assign \new_[25314]_  = ~A166 & \new_[25313]_ ;
  assign \new_[25315]_  = \new_[25314]_  & \new_[25309]_ ;
  assign \new_[25319]_  = A265 & A233;
  assign \new_[25320]_  = ~A232 & \new_[25319]_ ;
  assign \new_[25324]_  = A268 & A267;
  assign \new_[25325]_  = ~A266 & \new_[25324]_ ;
  assign \new_[25326]_  = \new_[25325]_  & \new_[25320]_ ;
  assign \new_[25330]_  = ~A167 & A169;
  assign \new_[25331]_  = ~A170 & \new_[25330]_ ;
  assign \new_[25335]_  = ~A201 & ~A200;
  assign \new_[25336]_  = ~A166 & \new_[25335]_ ;
  assign \new_[25337]_  = \new_[25336]_  & \new_[25331]_ ;
  assign \new_[25341]_  = A265 & A233;
  assign \new_[25342]_  = ~A232 & \new_[25341]_ ;
  assign \new_[25346]_  = A269 & A267;
  assign \new_[25347]_  = ~A266 & \new_[25346]_ ;
  assign \new_[25348]_  = \new_[25347]_  & \new_[25342]_ ;
  assign \new_[25352]_  = ~A167 & A169;
  assign \new_[25353]_  = ~A170 & \new_[25352]_ ;
  assign \new_[25357]_  = ~A201 & ~A200;
  assign \new_[25358]_  = ~A166 & \new_[25357]_ ;
  assign \new_[25359]_  = \new_[25358]_  & \new_[25353]_ ;
  assign \new_[25363]_  = A265 & ~A234;
  assign \new_[25364]_  = ~A233 & \new_[25363]_ ;
  assign \new_[25368]_  = A299 & ~A298;
  assign \new_[25369]_  = A266 & \new_[25368]_ ;
  assign \new_[25370]_  = \new_[25369]_  & \new_[25364]_ ;
  assign \new_[25374]_  = ~A167 & A169;
  assign \new_[25375]_  = ~A170 & \new_[25374]_ ;
  assign \new_[25379]_  = ~A201 & ~A200;
  assign \new_[25380]_  = ~A166 & \new_[25379]_ ;
  assign \new_[25381]_  = \new_[25380]_  & \new_[25375]_ ;
  assign \new_[25385]_  = ~A266 & ~A234;
  assign \new_[25386]_  = ~A233 & \new_[25385]_ ;
  assign \new_[25390]_  = A299 & ~A298;
  assign \new_[25391]_  = ~A267 & \new_[25390]_ ;
  assign \new_[25392]_  = \new_[25391]_  & \new_[25386]_ ;
  assign \new_[25396]_  = ~A167 & A169;
  assign \new_[25397]_  = ~A170 & \new_[25396]_ ;
  assign \new_[25401]_  = ~A201 & ~A200;
  assign \new_[25402]_  = ~A166 & \new_[25401]_ ;
  assign \new_[25403]_  = \new_[25402]_  & \new_[25397]_ ;
  assign \new_[25407]_  = ~A265 & ~A234;
  assign \new_[25408]_  = ~A233 & \new_[25407]_ ;
  assign \new_[25412]_  = A299 & ~A298;
  assign \new_[25413]_  = ~A266 & \new_[25412]_ ;
  assign \new_[25414]_  = \new_[25413]_  & \new_[25408]_ ;
  assign \new_[25418]_  = ~A167 & A169;
  assign \new_[25419]_  = ~A170 & \new_[25418]_ ;
  assign \new_[25423]_  = ~A201 & ~A200;
  assign \new_[25424]_  = ~A166 & \new_[25423]_ ;
  assign \new_[25425]_  = \new_[25424]_  & \new_[25419]_ ;
  assign \new_[25429]_  = A234 & ~A233;
  assign \new_[25430]_  = A232 & \new_[25429]_ ;
  assign \new_[25434]_  = ~A300 & A298;
  assign \new_[25435]_  = A235 & \new_[25434]_ ;
  assign \new_[25436]_  = \new_[25435]_  & \new_[25430]_ ;
  assign \new_[25440]_  = ~A167 & A169;
  assign \new_[25441]_  = ~A170 & \new_[25440]_ ;
  assign \new_[25445]_  = ~A201 & ~A200;
  assign \new_[25446]_  = ~A166 & \new_[25445]_ ;
  assign \new_[25447]_  = \new_[25446]_  & \new_[25441]_ ;
  assign \new_[25451]_  = A234 & ~A233;
  assign \new_[25452]_  = A232 & \new_[25451]_ ;
  assign \new_[25456]_  = A299 & A298;
  assign \new_[25457]_  = A235 & \new_[25456]_ ;
  assign \new_[25458]_  = \new_[25457]_  & \new_[25452]_ ;
  assign \new_[25462]_  = ~A167 & A169;
  assign \new_[25463]_  = ~A170 & \new_[25462]_ ;
  assign \new_[25467]_  = ~A201 & ~A200;
  assign \new_[25468]_  = ~A166 & \new_[25467]_ ;
  assign \new_[25469]_  = \new_[25468]_  & \new_[25463]_ ;
  assign \new_[25473]_  = A234 & ~A233;
  assign \new_[25474]_  = A232 & \new_[25473]_ ;
  assign \new_[25478]_  = ~A299 & ~A298;
  assign \new_[25479]_  = A235 & \new_[25478]_ ;
  assign \new_[25480]_  = \new_[25479]_  & \new_[25474]_ ;
  assign \new_[25484]_  = ~A167 & A169;
  assign \new_[25485]_  = ~A170 & \new_[25484]_ ;
  assign \new_[25489]_  = ~A201 & ~A200;
  assign \new_[25490]_  = ~A166 & \new_[25489]_ ;
  assign \new_[25491]_  = \new_[25490]_  & \new_[25485]_ ;
  assign \new_[25495]_  = A234 & ~A233;
  assign \new_[25496]_  = A232 & \new_[25495]_ ;
  assign \new_[25500]_  = A266 & ~A265;
  assign \new_[25501]_  = A235 & \new_[25500]_ ;
  assign \new_[25502]_  = \new_[25501]_  & \new_[25496]_ ;
  assign \new_[25506]_  = ~A167 & A169;
  assign \new_[25507]_  = ~A170 & \new_[25506]_ ;
  assign \new_[25511]_  = ~A201 & ~A200;
  assign \new_[25512]_  = ~A166 & \new_[25511]_ ;
  assign \new_[25513]_  = \new_[25512]_  & \new_[25507]_ ;
  assign \new_[25517]_  = A234 & ~A233;
  assign \new_[25518]_  = A232 & \new_[25517]_ ;
  assign \new_[25522]_  = ~A300 & A298;
  assign \new_[25523]_  = A236 & \new_[25522]_ ;
  assign \new_[25524]_  = \new_[25523]_  & \new_[25518]_ ;
  assign \new_[25528]_  = ~A167 & A169;
  assign \new_[25529]_  = ~A170 & \new_[25528]_ ;
  assign \new_[25533]_  = ~A201 & ~A200;
  assign \new_[25534]_  = ~A166 & \new_[25533]_ ;
  assign \new_[25535]_  = \new_[25534]_  & \new_[25529]_ ;
  assign \new_[25539]_  = A234 & ~A233;
  assign \new_[25540]_  = A232 & \new_[25539]_ ;
  assign \new_[25544]_  = A299 & A298;
  assign \new_[25545]_  = A236 & \new_[25544]_ ;
  assign \new_[25546]_  = \new_[25545]_  & \new_[25540]_ ;
  assign \new_[25550]_  = ~A167 & A169;
  assign \new_[25551]_  = ~A170 & \new_[25550]_ ;
  assign \new_[25555]_  = ~A201 & ~A200;
  assign \new_[25556]_  = ~A166 & \new_[25555]_ ;
  assign \new_[25557]_  = \new_[25556]_  & \new_[25551]_ ;
  assign \new_[25561]_  = A234 & ~A233;
  assign \new_[25562]_  = A232 & \new_[25561]_ ;
  assign \new_[25566]_  = ~A299 & ~A298;
  assign \new_[25567]_  = A236 & \new_[25566]_ ;
  assign \new_[25568]_  = \new_[25567]_  & \new_[25562]_ ;
  assign \new_[25572]_  = ~A167 & A169;
  assign \new_[25573]_  = ~A170 & \new_[25572]_ ;
  assign \new_[25577]_  = ~A201 & ~A200;
  assign \new_[25578]_  = ~A166 & \new_[25577]_ ;
  assign \new_[25579]_  = \new_[25578]_  & \new_[25573]_ ;
  assign \new_[25583]_  = A234 & ~A233;
  assign \new_[25584]_  = A232 & \new_[25583]_ ;
  assign \new_[25588]_  = A266 & ~A265;
  assign \new_[25589]_  = A236 & \new_[25588]_ ;
  assign \new_[25590]_  = \new_[25589]_  & \new_[25584]_ ;
  assign \new_[25594]_  = ~A167 & A169;
  assign \new_[25595]_  = ~A170 & \new_[25594]_ ;
  assign \new_[25599]_  = ~A201 & ~A200;
  assign \new_[25600]_  = ~A166 & \new_[25599]_ ;
  assign \new_[25601]_  = \new_[25600]_  & \new_[25595]_ ;
  assign \new_[25605]_  = A265 & ~A233;
  assign \new_[25606]_  = ~A232 & \new_[25605]_ ;
  assign \new_[25610]_  = A299 & ~A298;
  assign \new_[25611]_  = A266 & \new_[25610]_ ;
  assign \new_[25612]_  = \new_[25611]_  & \new_[25606]_ ;
  assign \new_[25616]_  = ~A167 & A169;
  assign \new_[25617]_  = ~A170 & \new_[25616]_ ;
  assign \new_[25621]_  = ~A201 & ~A200;
  assign \new_[25622]_  = ~A166 & \new_[25621]_ ;
  assign \new_[25623]_  = \new_[25622]_  & \new_[25617]_ ;
  assign \new_[25627]_  = ~A266 & ~A233;
  assign \new_[25628]_  = ~A232 & \new_[25627]_ ;
  assign \new_[25632]_  = A299 & ~A298;
  assign \new_[25633]_  = ~A267 & \new_[25632]_ ;
  assign \new_[25634]_  = \new_[25633]_  & \new_[25628]_ ;
  assign \new_[25638]_  = ~A167 & A169;
  assign \new_[25639]_  = ~A170 & \new_[25638]_ ;
  assign \new_[25643]_  = ~A201 & ~A200;
  assign \new_[25644]_  = ~A166 & \new_[25643]_ ;
  assign \new_[25645]_  = \new_[25644]_  & \new_[25639]_ ;
  assign \new_[25649]_  = ~A265 & ~A233;
  assign \new_[25650]_  = ~A232 & \new_[25649]_ ;
  assign \new_[25654]_  = A299 & ~A298;
  assign \new_[25655]_  = ~A266 & \new_[25654]_ ;
  assign \new_[25656]_  = \new_[25655]_  & \new_[25650]_ ;
  assign \new_[25660]_  = ~A167 & A169;
  assign \new_[25661]_  = ~A170 & \new_[25660]_ ;
  assign \new_[25665]_  = ~A200 & ~A199;
  assign \new_[25666]_  = ~A166 & \new_[25665]_ ;
  assign \new_[25667]_  = \new_[25666]_  & \new_[25661]_ ;
  assign \new_[25671]_  = A265 & A233;
  assign \new_[25672]_  = A232 & \new_[25671]_ ;
  assign \new_[25676]_  = A299 & ~A298;
  assign \new_[25677]_  = ~A267 & \new_[25676]_ ;
  assign \new_[25678]_  = \new_[25677]_  & \new_[25672]_ ;
  assign \new_[25682]_  = ~A167 & A169;
  assign \new_[25683]_  = ~A170 & \new_[25682]_ ;
  assign \new_[25687]_  = ~A200 & ~A199;
  assign \new_[25688]_  = ~A166 & \new_[25687]_ ;
  assign \new_[25689]_  = \new_[25688]_  & \new_[25683]_ ;
  assign \new_[25693]_  = A265 & A233;
  assign \new_[25694]_  = A232 & \new_[25693]_ ;
  assign \new_[25698]_  = A299 & ~A298;
  assign \new_[25699]_  = A266 & \new_[25698]_ ;
  assign \new_[25700]_  = \new_[25699]_  & \new_[25694]_ ;
  assign \new_[25704]_  = ~A167 & A169;
  assign \new_[25705]_  = ~A170 & \new_[25704]_ ;
  assign \new_[25709]_  = ~A200 & ~A199;
  assign \new_[25710]_  = ~A166 & \new_[25709]_ ;
  assign \new_[25711]_  = \new_[25710]_  & \new_[25705]_ ;
  assign \new_[25715]_  = ~A265 & A233;
  assign \new_[25716]_  = A232 & \new_[25715]_ ;
  assign \new_[25720]_  = A299 & ~A298;
  assign \new_[25721]_  = ~A266 & \new_[25720]_ ;
  assign \new_[25722]_  = \new_[25721]_  & \new_[25716]_ ;
  assign \new_[25726]_  = ~A167 & A169;
  assign \new_[25727]_  = ~A170 & \new_[25726]_ ;
  assign \new_[25731]_  = ~A200 & ~A199;
  assign \new_[25732]_  = ~A166 & \new_[25731]_ ;
  assign \new_[25733]_  = \new_[25732]_  & \new_[25727]_ ;
  assign \new_[25737]_  = A265 & A233;
  assign \new_[25738]_  = ~A232 & \new_[25737]_ ;
  assign \new_[25742]_  = A268 & A267;
  assign \new_[25743]_  = ~A266 & \new_[25742]_ ;
  assign \new_[25744]_  = \new_[25743]_  & \new_[25738]_ ;
  assign \new_[25748]_  = ~A167 & A169;
  assign \new_[25749]_  = ~A170 & \new_[25748]_ ;
  assign \new_[25753]_  = ~A200 & ~A199;
  assign \new_[25754]_  = ~A166 & \new_[25753]_ ;
  assign \new_[25755]_  = \new_[25754]_  & \new_[25749]_ ;
  assign \new_[25759]_  = A265 & A233;
  assign \new_[25760]_  = ~A232 & \new_[25759]_ ;
  assign \new_[25764]_  = A269 & A267;
  assign \new_[25765]_  = ~A266 & \new_[25764]_ ;
  assign \new_[25766]_  = \new_[25765]_  & \new_[25760]_ ;
  assign \new_[25770]_  = ~A167 & A169;
  assign \new_[25771]_  = ~A170 & \new_[25770]_ ;
  assign \new_[25775]_  = ~A200 & ~A199;
  assign \new_[25776]_  = ~A166 & \new_[25775]_ ;
  assign \new_[25777]_  = \new_[25776]_  & \new_[25771]_ ;
  assign \new_[25781]_  = A265 & ~A234;
  assign \new_[25782]_  = ~A233 & \new_[25781]_ ;
  assign \new_[25786]_  = A299 & ~A298;
  assign \new_[25787]_  = A266 & \new_[25786]_ ;
  assign \new_[25788]_  = \new_[25787]_  & \new_[25782]_ ;
  assign \new_[25792]_  = ~A167 & A169;
  assign \new_[25793]_  = ~A170 & \new_[25792]_ ;
  assign \new_[25797]_  = ~A200 & ~A199;
  assign \new_[25798]_  = ~A166 & \new_[25797]_ ;
  assign \new_[25799]_  = \new_[25798]_  & \new_[25793]_ ;
  assign \new_[25803]_  = ~A266 & ~A234;
  assign \new_[25804]_  = ~A233 & \new_[25803]_ ;
  assign \new_[25808]_  = A299 & ~A298;
  assign \new_[25809]_  = ~A267 & \new_[25808]_ ;
  assign \new_[25810]_  = \new_[25809]_  & \new_[25804]_ ;
  assign \new_[25814]_  = ~A167 & A169;
  assign \new_[25815]_  = ~A170 & \new_[25814]_ ;
  assign \new_[25819]_  = ~A200 & ~A199;
  assign \new_[25820]_  = ~A166 & \new_[25819]_ ;
  assign \new_[25821]_  = \new_[25820]_  & \new_[25815]_ ;
  assign \new_[25825]_  = ~A265 & ~A234;
  assign \new_[25826]_  = ~A233 & \new_[25825]_ ;
  assign \new_[25830]_  = A299 & ~A298;
  assign \new_[25831]_  = ~A266 & \new_[25830]_ ;
  assign \new_[25832]_  = \new_[25831]_  & \new_[25826]_ ;
  assign \new_[25836]_  = ~A167 & A169;
  assign \new_[25837]_  = ~A170 & \new_[25836]_ ;
  assign \new_[25841]_  = ~A200 & ~A199;
  assign \new_[25842]_  = ~A166 & \new_[25841]_ ;
  assign \new_[25843]_  = \new_[25842]_  & \new_[25837]_ ;
  assign \new_[25847]_  = A234 & ~A233;
  assign \new_[25848]_  = A232 & \new_[25847]_ ;
  assign \new_[25852]_  = ~A300 & A298;
  assign \new_[25853]_  = A235 & \new_[25852]_ ;
  assign \new_[25854]_  = \new_[25853]_  & \new_[25848]_ ;
  assign \new_[25858]_  = ~A167 & A169;
  assign \new_[25859]_  = ~A170 & \new_[25858]_ ;
  assign \new_[25863]_  = ~A200 & ~A199;
  assign \new_[25864]_  = ~A166 & \new_[25863]_ ;
  assign \new_[25865]_  = \new_[25864]_  & \new_[25859]_ ;
  assign \new_[25869]_  = A234 & ~A233;
  assign \new_[25870]_  = A232 & \new_[25869]_ ;
  assign \new_[25874]_  = A299 & A298;
  assign \new_[25875]_  = A235 & \new_[25874]_ ;
  assign \new_[25876]_  = \new_[25875]_  & \new_[25870]_ ;
  assign \new_[25880]_  = ~A167 & A169;
  assign \new_[25881]_  = ~A170 & \new_[25880]_ ;
  assign \new_[25885]_  = ~A200 & ~A199;
  assign \new_[25886]_  = ~A166 & \new_[25885]_ ;
  assign \new_[25887]_  = \new_[25886]_  & \new_[25881]_ ;
  assign \new_[25891]_  = A234 & ~A233;
  assign \new_[25892]_  = A232 & \new_[25891]_ ;
  assign \new_[25896]_  = ~A299 & ~A298;
  assign \new_[25897]_  = A235 & \new_[25896]_ ;
  assign \new_[25898]_  = \new_[25897]_  & \new_[25892]_ ;
  assign \new_[25902]_  = ~A167 & A169;
  assign \new_[25903]_  = ~A170 & \new_[25902]_ ;
  assign \new_[25907]_  = ~A200 & ~A199;
  assign \new_[25908]_  = ~A166 & \new_[25907]_ ;
  assign \new_[25909]_  = \new_[25908]_  & \new_[25903]_ ;
  assign \new_[25913]_  = A234 & ~A233;
  assign \new_[25914]_  = A232 & \new_[25913]_ ;
  assign \new_[25918]_  = A266 & ~A265;
  assign \new_[25919]_  = A235 & \new_[25918]_ ;
  assign \new_[25920]_  = \new_[25919]_  & \new_[25914]_ ;
  assign \new_[25924]_  = ~A167 & A169;
  assign \new_[25925]_  = ~A170 & \new_[25924]_ ;
  assign \new_[25929]_  = ~A200 & ~A199;
  assign \new_[25930]_  = ~A166 & \new_[25929]_ ;
  assign \new_[25931]_  = \new_[25930]_  & \new_[25925]_ ;
  assign \new_[25935]_  = A234 & ~A233;
  assign \new_[25936]_  = A232 & \new_[25935]_ ;
  assign \new_[25940]_  = ~A300 & A298;
  assign \new_[25941]_  = A236 & \new_[25940]_ ;
  assign \new_[25942]_  = \new_[25941]_  & \new_[25936]_ ;
  assign \new_[25946]_  = ~A167 & A169;
  assign \new_[25947]_  = ~A170 & \new_[25946]_ ;
  assign \new_[25951]_  = ~A200 & ~A199;
  assign \new_[25952]_  = ~A166 & \new_[25951]_ ;
  assign \new_[25953]_  = \new_[25952]_  & \new_[25947]_ ;
  assign \new_[25957]_  = A234 & ~A233;
  assign \new_[25958]_  = A232 & \new_[25957]_ ;
  assign \new_[25962]_  = A299 & A298;
  assign \new_[25963]_  = A236 & \new_[25962]_ ;
  assign \new_[25964]_  = \new_[25963]_  & \new_[25958]_ ;
  assign \new_[25968]_  = ~A167 & A169;
  assign \new_[25969]_  = ~A170 & \new_[25968]_ ;
  assign \new_[25973]_  = ~A200 & ~A199;
  assign \new_[25974]_  = ~A166 & \new_[25973]_ ;
  assign \new_[25975]_  = \new_[25974]_  & \new_[25969]_ ;
  assign \new_[25979]_  = A234 & ~A233;
  assign \new_[25980]_  = A232 & \new_[25979]_ ;
  assign \new_[25984]_  = ~A299 & ~A298;
  assign \new_[25985]_  = A236 & \new_[25984]_ ;
  assign \new_[25986]_  = \new_[25985]_  & \new_[25980]_ ;
  assign \new_[25990]_  = ~A167 & A169;
  assign \new_[25991]_  = ~A170 & \new_[25990]_ ;
  assign \new_[25995]_  = ~A200 & ~A199;
  assign \new_[25996]_  = ~A166 & \new_[25995]_ ;
  assign \new_[25997]_  = \new_[25996]_  & \new_[25991]_ ;
  assign \new_[26001]_  = A234 & ~A233;
  assign \new_[26002]_  = A232 & \new_[26001]_ ;
  assign \new_[26006]_  = A266 & ~A265;
  assign \new_[26007]_  = A236 & \new_[26006]_ ;
  assign \new_[26008]_  = \new_[26007]_  & \new_[26002]_ ;
  assign \new_[26012]_  = ~A167 & A169;
  assign \new_[26013]_  = ~A170 & \new_[26012]_ ;
  assign \new_[26017]_  = ~A200 & ~A199;
  assign \new_[26018]_  = ~A166 & \new_[26017]_ ;
  assign \new_[26019]_  = \new_[26018]_  & \new_[26013]_ ;
  assign \new_[26023]_  = A265 & ~A233;
  assign \new_[26024]_  = ~A232 & \new_[26023]_ ;
  assign \new_[26028]_  = A299 & ~A298;
  assign \new_[26029]_  = A266 & \new_[26028]_ ;
  assign \new_[26030]_  = \new_[26029]_  & \new_[26024]_ ;
  assign \new_[26034]_  = ~A167 & A169;
  assign \new_[26035]_  = ~A170 & \new_[26034]_ ;
  assign \new_[26039]_  = ~A200 & ~A199;
  assign \new_[26040]_  = ~A166 & \new_[26039]_ ;
  assign \new_[26041]_  = \new_[26040]_  & \new_[26035]_ ;
  assign \new_[26045]_  = ~A266 & ~A233;
  assign \new_[26046]_  = ~A232 & \new_[26045]_ ;
  assign \new_[26050]_  = A299 & ~A298;
  assign \new_[26051]_  = ~A267 & \new_[26050]_ ;
  assign \new_[26052]_  = \new_[26051]_  & \new_[26046]_ ;
  assign \new_[26056]_  = ~A167 & A169;
  assign \new_[26057]_  = ~A170 & \new_[26056]_ ;
  assign \new_[26061]_  = ~A200 & ~A199;
  assign \new_[26062]_  = ~A166 & \new_[26061]_ ;
  assign \new_[26063]_  = \new_[26062]_  & \new_[26057]_ ;
  assign \new_[26067]_  = ~A265 & ~A233;
  assign \new_[26068]_  = ~A232 & \new_[26067]_ ;
  assign \new_[26072]_  = A299 & ~A298;
  assign \new_[26073]_  = ~A266 & \new_[26072]_ ;
  assign \new_[26074]_  = \new_[26073]_  & \new_[26068]_ ;
  assign \new_[26078]_  = ~A166 & ~A167;
  assign \new_[26079]_  = ~A169 & \new_[26078]_ ;
  assign \new_[26083]_  = A232 & A200;
  assign \new_[26084]_  = ~A199 & \new_[26083]_ ;
  assign \new_[26085]_  = \new_[26084]_  & \new_[26079]_ ;
  assign \new_[26089]_  = ~A268 & A265;
  assign \new_[26090]_  = A233 & \new_[26089]_ ;
  assign \new_[26094]_  = A299 & ~A298;
  assign \new_[26095]_  = ~A269 & \new_[26094]_ ;
  assign \new_[26096]_  = \new_[26095]_  & \new_[26090]_ ;
  assign \new_[26100]_  = ~A166 & ~A167;
  assign \new_[26101]_  = ~A169 & \new_[26100]_ ;
  assign \new_[26105]_  = ~A233 & A200;
  assign \new_[26106]_  = ~A199 & \new_[26105]_ ;
  assign \new_[26107]_  = \new_[26106]_  & \new_[26101]_ ;
  assign \new_[26111]_  = A265 & ~A236;
  assign \new_[26112]_  = ~A235 & \new_[26111]_ ;
  assign \new_[26116]_  = A299 & ~A298;
  assign \new_[26117]_  = A266 & \new_[26116]_ ;
  assign \new_[26118]_  = \new_[26117]_  & \new_[26112]_ ;
  assign \new_[26122]_  = ~A166 & ~A167;
  assign \new_[26123]_  = ~A169 & \new_[26122]_ ;
  assign \new_[26127]_  = ~A233 & A200;
  assign \new_[26128]_  = ~A199 & \new_[26127]_ ;
  assign \new_[26129]_  = \new_[26128]_  & \new_[26123]_ ;
  assign \new_[26133]_  = ~A266 & ~A236;
  assign \new_[26134]_  = ~A235 & \new_[26133]_ ;
  assign \new_[26138]_  = A299 & ~A298;
  assign \new_[26139]_  = ~A267 & \new_[26138]_ ;
  assign \new_[26140]_  = \new_[26139]_  & \new_[26134]_ ;
  assign \new_[26144]_  = ~A166 & ~A167;
  assign \new_[26145]_  = ~A169 & \new_[26144]_ ;
  assign \new_[26149]_  = ~A233 & A200;
  assign \new_[26150]_  = ~A199 & \new_[26149]_ ;
  assign \new_[26151]_  = \new_[26150]_  & \new_[26145]_ ;
  assign \new_[26155]_  = ~A265 & ~A236;
  assign \new_[26156]_  = ~A235 & \new_[26155]_ ;
  assign \new_[26160]_  = A299 & ~A298;
  assign \new_[26161]_  = ~A266 & \new_[26160]_ ;
  assign \new_[26162]_  = \new_[26161]_  & \new_[26156]_ ;
  assign \new_[26166]_  = ~A166 & ~A167;
  assign \new_[26167]_  = ~A169 & \new_[26166]_ ;
  assign \new_[26171]_  = ~A233 & A200;
  assign \new_[26172]_  = ~A199 & \new_[26171]_ ;
  assign \new_[26173]_  = \new_[26172]_  & \new_[26167]_ ;
  assign \new_[26177]_  = ~A268 & ~A266;
  assign \new_[26178]_  = ~A234 & \new_[26177]_ ;
  assign \new_[26182]_  = A299 & ~A298;
  assign \new_[26183]_  = ~A269 & \new_[26182]_ ;
  assign \new_[26184]_  = \new_[26183]_  & \new_[26178]_ ;
  assign \new_[26188]_  = ~A166 & ~A167;
  assign \new_[26189]_  = ~A169 & \new_[26188]_ ;
  assign \new_[26193]_  = A232 & A200;
  assign \new_[26194]_  = ~A199 & \new_[26193]_ ;
  assign \new_[26195]_  = \new_[26194]_  & \new_[26189]_ ;
  assign \new_[26199]_  = A235 & A234;
  assign \new_[26200]_  = ~A233 & \new_[26199]_ ;
  assign \new_[26204]_  = ~A302 & ~A301;
  assign \new_[26205]_  = A298 & \new_[26204]_ ;
  assign \new_[26206]_  = \new_[26205]_  & \new_[26200]_ ;
  assign \new_[26210]_  = ~A166 & ~A167;
  assign \new_[26211]_  = ~A169 & \new_[26210]_ ;
  assign \new_[26215]_  = A232 & A200;
  assign \new_[26216]_  = ~A199 & \new_[26215]_ ;
  assign \new_[26217]_  = \new_[26216]_  & \new_[26211]_ ;
  assign \new_[26221]_  = A236 & A234;
  assign \new_[26222]_  = ~A233 & \new_[26221]_ ;
  assign \new_[26226]_  = ~A302 & ~A301;
  assign \new_[26227]_  = A298 & \new_[26226]_ ;
  assign \new_[26228]_  = \new_[26227]_  & \new_[26222]_ ;
  assign \new_[26232]_  = ~A166 & ~A167;
  assign \new_[26233]_  = ~A169 & \new_[26232]_ ;
  assign \new_[26237]_  = ~A232 & A200;
  assign \new_[26238]_  = ~A199 & \new_[26237]_ ;
  assign \new_[26239]_  = \new_[26238]_  & \new_[26233]_ ;
  assign \new_[26243]_  = ~A268 & ~A266;
  assign \new_[26244]_  = ~A233 & \new_[26243]_ ;
  assign \new_[26248]_  = A299 & ~A298;
  assign \new_[26249]_  = ~A269 & \new_[26248]_ ;
  assign \new_[26250]_  = \new_[26249]_  & \new_[26244]_ ;
  assign \new_[26254]_  = ~A166 & ~A167;
  assign \new_[26255]_  = ~A169 & \new_[26254]_ ;
  assign \new_[26259]_  = A201 & ~A200;
  assign \new_[26260]_  = A199 & \new_[26259]_ ;
  assign \new_[26261]_  = \new_[26260]_  & \new_[26255]_ ;
  assign \new_[26265]_  = A233 & ~A232;
  assign \new_[26266]_  = A202 & \new_[26265]_ ;
  assign \new_[26270]_  = ~A302 & ~A301;
  assign \new_[26271]_  = ~A299 & \new_[26270]_ ;
  assign \new_[26272]_  = \new_[26271]_  & \new_[26266]_ ;
  assign \new_[26276]_  = ~A166 & ~A167;
  assign \new_[26277]_  = ~A169 & \new_[26276]_ ;
  assign \new_[26281]_  = A201 & ~A200;
  assign \new_[26282]_  = A199 & \new_[26281]_ ;
  assign \new_[26283]_  = \new_[26282]_  & \new_[26277]_ ;
  assign \new_[26287]_  = A233 & ~A232;
  assign \new_[26288]_  = A203 & \new_[26287]_ ;
  assign \new_[26292]_  = ~A302 & ~A301;
  assign \new_[26293]_  = ~A299 & \new_[26292]_ ;
  assign \new_[26294]_  = \new_[26293]_  & \new_[26288]_ ;
  assign \new_[26298]_  = A167 & ~A168;
  assign \new_[26299]_  = ~A169 & \new_[26298]_ ;
  assign \new_[26303]_  = A200 & ~A199;
  assign \new_[26304]_  = A166 & \new_[26303]_ ;
  assign \new_[26305]_  = \new_[26304]_  & \new_[26299]_ ;
  assign \new_[26309]_  = A265 & A233;
  assign \new_[26310]_  = A232 & \new_[26309]_ ;
  assign \new_[26314]_  = A299 & ~A298;
  assign \new_[26315]_  = ~A267 & \new_[26314]_ ;
  assign \new_[26316]_  = \new_[26315]_  & \new_[26310]_ ;
  assign \new_[26320]_  = A167 & ~A168;
  assign \new_[26321]_  = ~A169 & \new_[26320]_ ;
  assign \new_[26325]_  = A200 & ~A199;
  assign \new_[26326]_  = A166 & \new_[26325]_ ;
  assign \new_[26327]_  = \new_[26326]_  & \new_[26321]_ ;
  assign \new_[26331]_  = A265 & A233;
  assign \new_[26332]_  = A232 & \new_[26331]_ ;
  assign \new_[26336]_  = A299 & ~A298;
  assign \new_[26337]_  = A266 & \new_[26336]_ ;
  assign \new_[26338]_  = \new_[26337]_  & \new_[26332]_ ;
  assign \new_[26342]_  = A167 & ~A168;
  assign \new_[26343]_  = ~A169 & \new_[26342]_ ;
  assign \new_[26347]_  = A200 & ~A199;
  assign \new_[26348]_  = A166 & \new_[26347]_ ;
  assign \new_[26349]_  = \new_[26348]_  & \new_[26343]_ ;
  assign \new_[26353]_  = ~A265 & A233;
  assign \new_[26354]_  = A232 & \new_[26353]_ ;
  assign \new_[26358]_  = A299 & ~A298;
  assign \new_[26359]_  = ~A266 & \new_[26358]_ ;
  assign \new_[26360]_  = \new_[26359]_  & \new_[26354]_ ;
  assign \new_[26364]_  = A167 & ~A168;
  assign \new_[26365]_  = ~A169 & \new_[26364]_ ;
  assign \new_[26369]_  = A200 & ~A199;
  assign \new_[26370]_  = A166 & \new_[26369]_ ;
  assign \new_[26371]_  = \new_[26370]_  & \new_[26365]_ ;
  assign \new_[26375]_  = A265 & A233;
  assign \new_[26376]_  = ~A232 & \new_[26375]_ ;
  assign \new_[26380]_  = A268 & A267;
  assign \new_[26381]_  = ~A266 & \new_[26380]_ ;
  assign \new_[26382]_  = \new_[26381]_  & \new_[26376]_ ;
  assign \new_[26386]_  = A167 & ~A168;
  assign \new_[26387]_  = ~A169 & \new_[26386]_ ;
  assign \new_[26391]_  = A200 & ~A199;
  assign \new_[26392]_  = A166 & \new_[26391]_ ;
  assign \new_[26393]_  = \new_[26392]_  & \new_[26387]_ ;
  assign \new_[26397]_  = A265 & A233;
  assign \new_[26398]_  = ~A232 & \new_[26397]_ ;
  assign \new_[26402]_  = A269 & A267;
  assign \new_[26403]_  = ~A266 & \new_[26402]_ ;
  assign \new_[26404]_  = \new_[26403]_  & \new_[26398]_ ;
  assign \new_[26408]_  = A167 & ~A168;
  assign \new_[26409]_  = ~A169 & \new_[26408]_ ;
  assign \new_[26413]_  = A200 & ~A199;
  assign \new_[26414]_  = A166 & \new_[26413]_ ;
  assign \new_[26415]_  = \new_[26414]_  & \new_[26409]_ ;
  assign \new_[26419]_  = A265 & ~A234;
  assign \new_[26420]_  = ~A233 & \new_[26419]_ ;
  assign \new_[26424]_  = A299 & ~A298;
  assign \new_[26425]_  = A266 & \new_[26424]_ ;
  assign \new_[26426]_  = \new_[26425]_  & \new_[26420]_ ;
  assign \new_[26430]_  = A167 & ~A168;
  assign \new_[26431]_  = ~A169 & \new_[26430]_ ;
  assign \new_[26435]_  = A200 & ~A199;
  assign \new_[26436]_  = A166 & \new_[26435]_ ;
  assign \new_[26437]_  = \new_[26436]_  & \new_[26431]_ ;
  assign \new_[26441]_  = ~A266 & ~A234;
  assign \new_[26442]_  = ~A233 & \new_[26441]_ ;
  assign \new_[26446]_  = A299 & ~A298;
  assign \new_[26447]_  = ~A267 & \new_[26446]_ ;
  assign \new_[26448]_  = \new_[26447]_  & \new_[26442]_ ;
  assign \new_[26452]_  = A167 & ~A168;
  assign \new_[26453]_  = ~A169 & \new_[26452]_ ;
  assign \new_[26457]_  = A200 & ~A199;
  assign \new_[26458]_  = A166 & \new_[26457]_ ;
  assign \new_[26459]_  = \new_[26458]_  & \new_[26453]_ ;
  assign \new_[26463]_  = ~A265 & ~A234;
  assign \new_[26464]_  = ~A233 & \new_[26463]_ ;
  assign \new_[26468]_  = A299 & ~A298;
  assign \new_[26469]_  = ~A266 & \new_[26468]_ ;
  assign \new_[26470]_  = \new_[26469]_  & \new_[26464]_ ;
  assign \new_[26474]_  = A167 & ~A168;
  assign \new_[26475]_  = ~A169 & \new_[26474]_ ;
  assign \new_[26479]_  = A200 & ~A199;
  assign \new_[26480]_  = A166 & \new_[26479]_ ;
  assign \new_[26481]_  = \new_[26480]_  & \new_[26475]_ ;
  assign \new_[26485]_  = A234 & ~A233;
  assign \new_[26486]_  = A232 & \new_[26485]_ ;
  assign \new_[26490]_  = ~A300 & A298;
  assign \new_[26491]_  = A235 & \new_[26490]_ ;
  assign \new_[26492]_  = \new_[26491]_  & \new_[26486]_ ;
  assign \new_[26496]_  = A167 & ~A168;
  assign \new_[26497]_  = ~A169 & \new_[26496]_ ;
  assign \new_[26501]_  = A200 & ~A199;
  assign \new_[26502]_  = A166 & \new_[26501]_ ;
  assign \new_[26503]_  = \new_[26502]_  & \new_[26497]_ ;
  assign \new_[26507]_  = A234 & ~A233;
  assign \new_[26508]_  = A232 & \new_[26507]_ ;
  assign \new_[26512]_  = A299 & A298;
  assign \new_[26513]_  = A235 & \new_[26512]_ ;
  assign \new_[26514]_  = \new_[26513]_  & \new_[26508]_ ;
  assign \new_[26518]_  = A167 & ~A168;
  assign \new_[26519]_  = ~A169 & \new_[26518]_ ;
  assign \new_[26523]_  = A200 & ~A199;
  assign \new_[26524]_  = A166 & \new_[26523]_ ;
  assign \new_[26525]_  = \new_[26524]_  & \new_[26519]_ ;
  assign \new_[26529]_  = A234 & ~A233;
  assign \new_[26530]_  = A232 & \new_[26529]_ ;
  assign \new_[26534]_  = ~A299 & ~A298;
  assign \new_[26535]_  = A235 & \new_[26534]_ ;
  assign \new_[26536]_  = \new_[26535]_  & \new_[26530]_ ;
  assign \new_[26540]_  = A167 & ~A168;
  assign \new_[26541]_  = ~A169 & \new_[26540]_ ;
  assign \new_[26545]_  = A200 & ~A199;
  assign \new_[26546]_  = A166 & \new_[26545]_ ;
  assign \new_[26547]_  = \new_[26546]_  & \new_[26541]_ ;
  assign \new_[26551]_  = A234 & ~A233;
  assign \new_[26552]_  = A232 & \new_[26551]_ ;
  assign \new_[26556]_  = A266 & ~A265;
  assign \new_[26557]_  = A235 & \new_[26556]_ ;
  assign \new_[26558]_  = \new_[26557]_  & \new_[26552]_ ;
  assign \new_[26562]_  = A167 & ~A168;
  assign \new_[26563]_  = ~A169 & \new_[26562]_ ;
  assign \new_[26567]_  = A200 & ~A199;
  assign \new_[26568]_  = A166 & \new_[26567]_ ;
  assign \new_[26569]_  = \new_[26568]_  & \new_[26563]_ ;
  assign \new_[26573]_  = A234 & ~A233;
  assign \new_[26574]_  = A232 & \new_[26573]_ ;
  assign \new_[26578]_  = ~A300 & A298;
  assign \new_[26579]_  = A236 & \new_[26578]_ ;
  assign \new_[26580]_  = \new_[26579]_  & \new_[26574]_ ;
  assign \new_[26584]_  = A167 & ~A168;
  assign \new_[26585]_  = ~A169 & \new_[26584]_ ;
  assign \new_[26589]_  = A200 & ~A199;
  assign \new_[26590]_  = A166 & \new_[26589]_ ;
  assign \new_[26591]_  = \new_[26590]_  & \new_[26585]_ ;
  assign \new_[26595]_  = A234 & ~A233;
  assign \new_[26596]_  = A232 & \new_[26595]_ ;
  assign \new_[26600]_  = A299 & A298;
  assign \new_[26601]_  = A236 & \new_[26600]_ ;
  assign \new_[26602]_  = \new_[26601]_  & \new_[26596]_ ;
  assign \new_[26606]_  = A167 & ~A168;
  assign \new_[26607]_  = ~A169 & \new_[26606]_ ;
  assign \new_[26611]_  = A200 & ~A199;
  assign \new_[26612]_  = A166 & \new_[26611]_ ;
  assign \new_[26613]_  = \new_[26612]_  & \new_[26607]_ ;
  assign \new_[26617]_  = A234 & ~A233;
  assign \new_[26618]_  = A232 & \new_[26617]_ ;
  assign \new_[26622]_  = ~A299 & ~A298;
  assign \new_[26623]_  = A236 & \new_[26622]_ ;
  assign \new_[26624]_  = \new_[26623]_  & \new_[26618]_ ;
  assign \new_[26628]_  = A167 & ~A168;
  assign \new_[26629]_  = ~A169 & \new_[26628]_ ;
  assign \new_[26633]_  = A200 & ~A199;
  assign \new_[26634]_  = A166 & \new_[26633]_ ;
  assign \new_[26635]_  = \new_[26634]_  & \new_[26629]_ ;
  assign \new_[26639]_  = A234 & ~A233;
  assign \new_[26640]_  = A232 & \new_[26639]_ ;
  assign \new_[26644]_  = A266 & ~A265;
  assign \new_[26645]_  = A236 & \new_[26644]_ ;
  assign \new_[26646]_  = \new_[26645]_  & \new_[26640]_ ;
  assign \new_[26650]_  = A167 & ~A168;
  assign \new_[26651]_  = ~A169 & \new_[26650]_ ;
  assign \new_[26655]_  = A200 & ~A199;
  assign \new_[26656]_  = A166 & \new_[26655]_ ;
  assign \new_[26657]_  = \new_[26656]_  & \new_[26651]_ ;
  assign \new_[26661]_  = A265 & ~A233;
  assign \new_[26662]_  = ~A232 & \new_[26661]_ ;
  assign \new_[26666]_  = A299 & ~A298;
  assign \new_[26667]_  = A266 & \new_[26666]_ ;
  assign \new_[26668]_  = \new_[26667]_  & \new_[26662]_ ;
  assign \new_[26672]_  = A167 & ~A168;
  assign \new_[26673]_  = ~A169 & \new_[26672]_ ;
  assign \new_[26677]_  = A200 & ~A199;
  assign \new_[26678]_  = A166 & \new_[26677]_ ;
  assign \new_[26679]_  = \new_[26678]_  & \new_[26673]_ ;
  assign \new_[26683]_  = ~A266 & ~A233;
  assign \new_[26684]_  = ~A232 & \new_[26683]_ ;
  assign \new_[26688]_  = A299 & ~A298;
  assign \new_[26689]_  = ~A267 & \new_[26688]_ ;
  assign \new_[26690]_  = \new_[26689]_  & \new_[26684]_ ;
  assign \new_[26694]_  = A167 & ~A168;
  assign \new_[26695]_  = ~A169 & \new_[26694]_ ;
  assign \new_[26699]_  = A200 & ~A199;
  assign \new_[26700]_  = A166 & \new_[26699]_ ;
  assign \new_[26701]_  = \new_[26700]_  & \new_[26695]_ ;
  assign \new_[26705]_  = ~A265 & ~A233;
  assign \new_[26706]_  = ~A232 & \new_[26705]_ ;
  assign \new_[26710]_  = A299 & ~A298;
  assign \new_[26711]_  = ~A266 & \new_[26710]_ ;
  assign \new_[26712]_  = \new_[26711]_  & \new_[26706]_ ;
  assign \new_[26716]_  = A167 & ~A168;
  assign \new_[26717]_  = ~A169 & \new_[26716]_ ;
  assign \new_[26721]_  = ~A200 & A199;
  assign \new_[26722]_  = A166 & \new_[26721]_ ;
  assign \new_[26723]_  = \new_[26722]_  & \new_[26717]_ ;
  assign \new_[26727]_  = ~A232 & A202;
  assign \new_[26728]_  = A201 & \new_[26727]_ ;
  assign \new_[26732]_  = ~A300 & ~A299;
  assign \new_[26733]_  = A233 & \new_[26732]_ ;
  assign \new_[26734]_  = \new_[26733]_  & \new_[26728]_ ;
  assign \new_[26738]_  = A167 & ~A168;
  assign \new_[26739]_  = ~A169 & \new_[26738]_ ;
  assign \new_[26743]_  = ~A200 & A199;
  assign \new_[26744]_  = A166 & \new_[26743]_ ;
  assign \new_[26745]_  = \new_[26744]_  & \new_[26739]_ ;
  assign \new_[26749]_  = ~A232 & A202;
  assign \new_[26750]_  = A201 & \new_[26749]_ ;
  assign \new_[26754]_  = A299 & A298;
  assign \new_[26755]_  = A233 & \new_[26754]_ ;
  assign \new_[26756]_  = \new_[26755]_  & \new_[26750]_ ;
  assign \new_[26760]_  = A167 & ~A168;
  assign \new_[26761]_  = ~A169 & \new_[26760]_ ;
  assign \new_[26765]_  = ~A200 & A199;
  assign \new_[26766]_  = A166 & \new_[26765]_ ;
  assign \new_[26767]_  = \new_[26766]_  & \new_[26761]_ ;
  assign \new_[26771]_  = ~A232 & A202;
  assign \new_[26772]_  = A201 & \new_[26771]_ ;
  assign \new_[26776]_  = ~A299 & ~A298;
  assign \new_[26777]_  = A233 & \new_[26776]_ ;
  assign \new_[26778]_  = \new_[26777]_  & \new_[26772]_ ;
  assign \new_[26782]_  = A167 & ~A168;
  assign \new_[26783]_  = ~A169 & \new_[26782]_ ;
  assign \new_[26787]_  = ~A200 & A199;
  assign \new_[26788]_  = A166 & \new_[26787]_ ;
  assign \new_[26789]_  = \new_[26788]_  & \new_[26783]_ ;
  assign \new_[26793]_  = ~A232 & A202;
  assign \new_[26794]_  = A201 & \new_[26793]_ ;
  assign \new_[26798]_  = A266 & ~A265;
  assign \new_[26799]_  = A233 & \new_[26798]_ ;
  assign \new_[26800]_  = \new_[26799]_  & \new_[26794]_ ;
  assign \new_[26804]_  = A167 & ~A168;
  assign \new_[26805]_  = ~A169 & \new_[26804]_ ;
  assign \new_[26809]_  = ~A200 & A199;
  assign \new_[26810]_  = A166 & \new_[26809]_ ;
  assign \new_[26811]_  = \new_[26810]_  & \new_[26805]_ ;
  assign \new_[26815]_  = ~A232 & A203;
  assign \new_[26816]_  = A201 & \new_[26815]_ ;
  assign \new_[26820]_  = ~A300 & ~A299;
  assign \new_[26821]_  = A233 & \new_[26820]_ ;
  assign \new_[26822]_  = \new_[26821]_  & \new_[26816]_ ;
  assign \new_[26826]_  = A167 & ~A168;
  assign \new_[26827]_  = ~A169 & \new_[26826]_ ;
  assign \new_[26831]_  = ~A200 & A199;
  assign \new_[26832]_  = A166 & \new_[26831]_ ;
  assign \new_[26833]_  = \new_[26832]_  & \new_[26827]_ ;
  assign \new_[26837]_  = ~A232 & A203;
  assign \new_[26838]_  = A201 & \new_[26837]_ ;
  assign \new_[26842]_  = A299 & A298;
  assign \new_[26843]_  = A233 & \new_[26842]_ ;
  assign \new_[26844]_  = \new_[26843]_  & \new_[26838]_ ;
  assign \new_[26848]_  = A167 & ~A168;
  assign \new_[26849]_  = ~A169 & \new_[26848]_ ;
  assign \new_[26853]_  = ~A200 & A199;
  assign \new_[26854]_  = A166 & \new_[26853]_ ;
  assign \new_[26855]_  = \new_[26854]_  & \new_[26849]_ ;
  assign \new_[26859]_  = ~A232 & A203;
  assign \new_[26860]_  = A201 & \new_[26859]_ ;
  assign \new_[26864]_  = ~A299 & ~A298;
  assign \new_[26865]_  = A233 & \new_[26864]_ ;
  assign \new_[26866]_  = \new_[26865]_  & \new_[26860]_ ;
  assign \new_[26870]_  = A167 & ~A168;
  assign \new_[26871]_  = ~A169 & \new_[26870]_ ;
  assign \new_[26875]_  = ~A200 & A199;
  assign \new_[26876]_  = A166 & \new_[26875]_ ;
  assign \new_[26877]_  = \new_[26876]_  & \new_[26871]_ ;
  assign \new_[26881]_  = ~A232 & A203;
  assign \new_[26882]_  = A201 & \new_[26881]_ ;
  assign \new_[26886]_  = A266 & ~A265;
  assign \new_[26887]_  = A233 & \new_[26886]_ ;
  assign \new_[26888]_  = \new_[26887]_  & \new_[26882]_ ;
  assign \new_[26892]_  = A167 & ~A169;
  assign \new_[26893]_  = A170 & \new_[26892]_ ;
  assign \new_[26897]_  = A200 & A199;
  assign \new_[26898]_  = ~A166 & \new_[26897]_ ;
  assign \new_[26899]_  = \new_[26898]_  & \new_[26893]_ ;
  assign \new_[26903]_  = A265 & A233;
  assign \new_[26904]_  = A232 & \new_[26903]_ ;
  assign \new_[26908]_  = A299 & ~A298;
  assign \new_[26909]_  = ~A267 & \new_[26908]_ ;
  assign \new_[26910]_  = \new_[26909]_  & \new_[26904]_ ;
  assign \new_[26914]_  = A167 & ~A169;
  assign \new_[26915]_  = A170 & \new_[26914]_ ;
  assign \new_[26919]_  = A200 & A199;
  assign \new_[26920]_  = ~A166 & \new_[26919]_ ;
  assign \new_[26921]_  = \new_[26920]_  & \new_[26915]_ ;
  assign \new_[26925]_  = A265 & A233;
  assign \new_[26926]_  = A232 & \new_[26925]_ ;
  assign \new_[26930]_  = A299 & ~A298;
  assign \new_[26931]_  = A266 & \new_[26930]_ ;
  assign \new_[26932]_  = \new_[26931]_  & \new_[26926]_ ;
  assign \new_[26936]_  = A167 & ~A169;
  assign \new_[26937]_  = A170 & \new_[26936]_ ;
  assign \new_[26941]_  = A200 & A199;
  assign \new_[26942]_  = ~A166 & \new_[26941]_ ;
  assign \new_[26943]_  = \new_[26942]_  & \new_[26937]_ ;
  assign \new_[26947]_  = ~A265 & A233;
  assign \new_[26948]_  = A232 & \new_[26947]_ ;
  assign \new_[26952]_  = A299 & ~A298;
  assign \new_[26953]_  = ~A266 & \new_[26952]_ ;
  assign \new_[26954]_  = \new_[26953]_  & \new_[26948]_ ;
  assign \new_[26958]_  = A167 & ~A169;
  assign \new_[26959]_  = A170 & \new_[26958]_ ;
  assign \new_[26963]_  = A200 & A199;
  assign \new_[26964]_  = ~A166 & \new_[26963]_ ;
  assign \new_[26965]_  = \new_[26964]_  & \new_[26959]_ ;
  assign \new_[26969]_  = A265 & A233;
  assign \new_[26970]_  = ~A232 & \new_[26969]_ ;
  assign \new_[26974]_  = A268 & A267;
  assign \new_[26975]_  = ~A266 & \new_[26974]_ ;
  assign \new_[26976]_  = \new_[26975]_  & \new_[26970]_ ;
  assign \new_[26980]_  = A167 & ~A169;
  assign \new_[26981]_  = A170 & \new_[26980]_ ;
  assign \new_[26985]_  = A200 & A199;
  assign \new_[26986]_  = ~A166 & \new_[26985]_ ;
  assign \new_[26987]_  = \new_[26986]_  & \new_[26981]_ ;
  assign \new_[26991]_  = A265 & A233;
  assign \new_[26992]_  = ~A232 & \new_[26991]_ ;
  assign \new_[26996]_  = A269 & A267;
  assign \new_[26997]_  = ~A266 & \new_[26996]_ ;
  assign \new_[26998]_  = \new_[26997]_  & \new_[26992]_ ;
  assign \new_[27002]_  = A167 & ~A169;
  assign \new_[27003]_  = A170 & \new_[27002]_ ;
  assign \new_[27007]_  = A200 & A199;
  assign \new_[27008]_  = ~A166 & \new_[27007]_ ;
  assign \new_[27009]_  = \new_[27008]_  & \new_[27003]_ ;
  assign \new_[27013]_  = A265 & ~A234;
  assign \new_[27014]_  = ~A233 & \new_[27013]_ ;
  assign \new_[27018]_  = A299 & ~A298;
  assign \new_[27019]_  = A266 & \new_[27018]_ ;
  assign \new_[27020]_  = \new_[27019]_  & \new_[27014]_ ;
  assign \new_[27024]_  = A167 & ~A169;
  assign \new_[27025]_  = A170 & \new_[27024]_ ;
  assign \new_[27029]_  = A200 & A199;
  assign \new_[27030]_  = ~A166 & \new_[27029]_ ;
  assign \new_[27031]_  = \new_[27030]_  & \new_[27025]_ ;
  assign \new_[27035]_  = ~A266 & ~A234;
  assign \new_[27036]_  = ~A233 & \new_[27035]_ ;
  assign \new_[27040]_  = A299 & ~A298;
  assign \new_[27041]_  = ~A267 & \new_[27040]_ ;
  assign \new_[27042]_  = \new_[27041]_  & \new_[27036]_ ;
  assign \new_[27046]_  = A167 & ~A169;
  assign \new_[27047]_  = A170 & \new_[27046]_ ;
  assign \new_[27051]_  = A200 & A199;
  assign \new_[27052]_  = ~A166 & \new_[27051]_ ;
  assign \new_[27053]_  = \new_[27052]_  & \new_[27047]_ ;
  assign \new_[27057]_  = ~A265 & ~A234;
  assign \new_[27058]_  = ~A233 & \new_[27057]_ ;
  assign \new_[27062]_  = A299 & ~A298;
  assign \new_[27063]_  = ~A266 & \new_[27062]_ ;
  assign \new_[27064]_  = \new_[27063]_  & \new_[27058]_ ;
  assign \new_[27068]_  = A167 & ~A169;
  assign \new_[27069]_  = A170 & \new_[27068]_ ;
  assign \new_[27073]_  = A200 & A199;
  assign \new_[27074]_  = ~A166 & \new_[27073]_ ;
  assign \new_[27075]_  = \new_[27074]_  & \new_[27069]_ ;
  assign \new_[27079]_  = A234 & ~A233;
  assign \new_[27080]_  = A232 & \new_[27079]_ ;
  assign \new_[27084]_  = ~A300 & A298;
  assign \new_[27085]_  = A235 & \new_[27084]_ ;
  assign \new_[27086]_  = \new_[27085]_  & \new_[27080]_ ;
  assign \new_[27090]_  = A167 & ~A169;
  assign \new_[27091]_  = A170 & \new_[27090]_ ;
  assign \new_[27095]_  = A200 & A199;
  assign \new_[27096]_  = ~A166 & \new_[27095]_ ;
  assign \new_[27097]_  = \new_[27096]_  & \new_[27091]_ ;
  assign \new_[27101]_  = A234 & ~A233;
  assign \new_[27102]_  = A232 & \new_[27101]_ ;
  assign \new_[27106]_  = A299 & A298;
  assign \new_[27107]_  = A235 & \new_[27106]_ ;
  assign \new_[27108]_  = \new_[27107]_  & \new_[27102]_ ;
  assign \new_[27112]_  = A167 & ~A169;
  assign \new_[27113]_  = A170 & \new_[27112]_ ;
  assign \new_[27117]_  = A200 & A199;
  assign \new_[27118]_  = ~A166 & \new_[27117]_ ;
  assign \new_[27119]_  = \new_[27118]_  & \new_[27113]_ ;
  assign \new_[27123]_  = A234 & ~A233;
  assign \new_[27124]_  = A232 & \new_[27123]_ ;
  assign \new_[27128]_  = ~A299 & ~A298;
  assign \new_[27129]_  = A235 & \new_[27128]_ ;
  assign \new_[27130]_  = \new_[27129]_  & \new_[27124]_ ;
  assign \new_[27134]_  = A167 & ~A169;
  assign \new_[27135]_  = A170 & \new_[27134]_ ;
  assign \new_[27139]_  = A200 & A199;
  assign \new_[27140]_  = ~A166 & \new_[27139]_ ;
  assign \new_[27141]_  = \new_[27140]_  & \new_[27135]_ ;
  assign \new_[27145]_  = A234 & ~A233;
  assign \new_[27146]_  = A232 & \new_[27145]_ ;
  assign \new_[27150]_  = A266 & ~A265;
  assign \new_[27151]_  = A235 & \new_[27150]_ ;
  assign \new_[27152]_  = \new_[27151]_  & \new_[27146]_ ;
  assign \new_[27156]_  = A167 & ~A169;
  assign \new_[27157]_  = A170 & \new_[27156]_ ;
  assign \new_[27161]_  = A200 & A199;
  assign \new_[27162]_  = ~A166 & \new_[27161]_ ;
  assign \new_[27163]_  = \new_[27162]_  & \new_[27157]_ ;
  assign \new_[27167]_  = A234 & ~A233;
  assign \new_[27168]_  = A232 & \new_[27167]_ ;
  assign \new_[27172]_  = ~A300 & A298;
  assign \new_[27173]_  = A236 & \new_[27172]_ ;
  assign \new_[27174]_  = \new_[27173]_  & \new_[27168]_ ;
  assign \new_[27178]_  = A167 & ~A169;
  assign \new_[27179]_  = A170 & \new_[27178]_ ;
  assign \new_[27183]_  = A200 & A199;
  assign \new_[27184]_  = ~A166 & \new_[27183]_ ;
  assign \new_[27185]_  = \new_[27184]_  & \new_[27179]_ ;
  assign \new_[27189]_  = A234 & ~A233;
  assign \new_[27190]_  = A232 & \new_[27189]_ ;
  assign \new_[27194]_  = A299 & A298;
  assign \new_[27195]_  = A236 & \new_[27194]_ ;
  assign \new_[27196]_  = \new_[27195]_  & \new_[27190]_ ;
  assign \new_[27200]_  = A167 & ~A169;
  assign \new_[27201]_  = A170 & \new_[27200]_ ;
  assign \new_[27205]_  = A200 & A199;
  assign \new_[27206]_  = ~A166 & \new_[27205]_ ;
  assign \new_[27207]_  = \new_[27206]_  & \new_[27201]_ ;
  assign \new_[27211]_  = A234 & ~A233;
  assign \new_[27212]_  = A232 & \new_[27211]_ ;
  assign \new_[27216]_  = ~A299 & ~A298;
  assign \new_[27217]_  = A236 & \new_[27216]_ ;
  assign \new_[27218]_  = \new_[27217]_  & \new_[27212]_ ;
  assign \new_[27222]_  = A167 & ~A169;
  assign \new_[27223]_  = A170 & \new_[27222]_ ;
  assign \new_[27227]_  = A200 & A199;
  assign \new_[27228]_  = ~A166 & \new_[27227]_ ;
  assign \new_[27229]_  = \new_[27228]_  & \new_[27223]_ ;
  assign \new_[27233]_  = A234 & ~A233;
  assign \new_[27234]_  = A232 & \new_[27233]_ ;
  assign \new_[27238]_  = A266 & ~A265;
  assign \new_[27239]_  = A236 & \new_[27238]_ ;
  assign \new_[27240]_  = \new_[27239]_  & \new_[27234]_ ;
  assign \new_[27244]_  = A167 & ~A169;
  assign \new_[27245]_  = A170 & \new_[27244]_ ;
  assign \new_[27249]_  = A200 & A199;
  assign \new_[27250]_  = ~A166 & \new_[27249]_ ;
  assign \new_[27251]_  = \new_[27250]_  & \new_[27245]_ ;
  assign \new_[27255]_  = A265 & ~A233;
  assign \new_[27256]_  = ~A232 & \new_[27255]_ ;
  assign \new_[27260]_  = A299 & ~A298;
  assign \new_[27261]_  = A266 & \new_[27260]_ ;
  assign \new_[27262]_  = \new_[27261]_  & \new_[27256]_ ;
  assign \new_[27266]_  = A167 & ~A169;
  assign \new_[27267]_  = A170 & \new_[27266]_ ;
  assign \new_[27271]_  = A200 & A199;
  assign \new_[27272]_  = ~A166 & \new_[27271]_ ;
  assign \new_[27273]_  = \new_[27272]_  & \new_[27267]_ ;
  assign \new_[27277]_  = ~A266 & ~A233;
  assign \new_[27278]_  = ~A232 & \new_[27277]_ ;
  assign \new_[27282]_  = A299 & ~A298;
  assign \new_[27283]_  = ~A267 & \new_[27282]_ ;
  assign \new_[27284]_  = \new_[27283]_  & \new_[27278]_ ;
  assign \new_[27288]_  = A167 & ~A169;
  assign \new_[27289]_  = A170 & \new_[27288]_ ;
  assign \new_[27293]_  = A200 & A199;
  assign \new_[27294]_  = ~A166 & \new_[27293]_ ;
  assign \new_[27295]_  = \new_[27294]_  & \new_[27289]_ ;
  assign \new_[27299]_  = ~A265 & ~A233;
  assign \new_[27300]_  = ~A232 & \new_[27299]_ ;
  assign \new_[27304]_  = A299 & ~A298;
  assign \new_[27305]_  = ~A266 & \new_[27304]_ ;
  assign \new_[27306]_  = \new_[27305]_  & \new_[27300]_ ;
  assign \new_[27310]_  = A167 & ~A169;
  assign \new_[27311]_  = A170 & \new_[27310]_ ;
  assign \new_[27315]_  = ~A202 & ~A200;
  assign \new_[27316]_  = ~A166 & \new_[27315]_ ;
  assign \new_[27317]_  = \new_[27316]_  & \new_[27311]_ ;
  assign \new_[27321]_  = A233 & ~A232;
  assign \new_[27322]_  = ~A203 & \new_[27321]_ ;
  assign \new_[27326]_  = ~A302 & ~A301;
  assign \new_[27327]_  = ~A299 & \new_[27326]_ ;
  assign \new_[27328]_  = \new_[27327]_  & \new_[27322]_ ;
  assign \new_[27332]_  = A167 & ~A169;
  assign \new_[27333]_  = A170 & \new_[27332]_ ;
  assign \new_[27337]_  = ~A201 & ~A200;
  assign \new_[27338]_  = ~A166 & \new_[27337]_ ;
  assign \new_[27339]_  = \new_[27338]_  & \new_[27333]_ ;
  assign \new_[27343]_  = A265 & A233;
  assign \new_[27344]_  = A232 & \new_[27343]_ ;
  assign \new_[27348]_  = A299 & ~A298;
  assign \new_[27349]_  = ~A267 & \new_[27348]_ ;
  assign \new_[27350]_  = \new_[27349]_  & \new_[27344]_ ;
  assign \new_[27354]_  = A167 & ~A169;
  assign \new_[27355]_  = A170 & \new_[27354]_ ;
  assign \new_[27359]_  = ~A201 & ~A200;
  assign \new_[27360]_  = ~A166 & \new_[27359]_ ;
  assign \new_[27361]_  = \new_[27360]_  & \new_[27355]_ ;
  assign \new_[27365]_  = A265 & A233;
  assign \new_[27366]_  = A232 & \new_[27365]_ ;
  assign \new_[27370]_  = A299 & ~A298;
  assign \new_[27371]_  = A266 & \new_[27370]_ ;
  assign \new_[27372]_  = \new_[27371]_  & \new_[27366]_ ;
  assign \new_[27376]_  = A167 & ~A169;
  assign \new_[27377]_  = A170 & \new_[27376]_ ;
  assign \new_[27381]_  = ~A201 & ~A200;
  assign \new_[27382]_  = ~A166 & \new_[27381]_ ;
  assign \new_[27383]_  = \new_[27382]_  & \new_[27377]_ ;
  assign \new_[27387]_  = ~A265 & A233;
  assign \new_[27388]_  = A232 & \new_[27387]_ ;
  assign \new_[27392]_  = A299 & ~A298;
  assign \new_[27393]_  = ~A266 & \new_[27392]_ ;
  assign \new_[27394]_  = \new_[27393]_  & \new_[27388]_ ;
  assign \new_[27398]_  = A167 & ~A169;
  assign \new_[27399]_  = A170 & \new_[27398]_ ;
  assign \new_[27403]_  = ~A201 & ~A200;
  assign \new_[27404]_  = ~A166 & \new_[27403]_ ;
  assign \new_[27405]_  = \new_[27404]_  & \new_[27399]_ ;
  assign \new_[27409]_  = A265 & A233;
  assign \new_[27410]_  = ~A232 & \new_[27409]_ ;
  assign \new_[27414]_  = A268 & A267;
  assign \new_[27415]_  = ~A266 & \new_[27414]_ ;
  assign \new_[27416]_  = \new_[27415]_  & \new_[27410]_ ;
  assign \new_[27420]_  = A167 & ~A169;
  assign \new_[27421]_  = A170 & \new_[27420]_ ;
  assign \new_[27425]_  = ~A201 & ~A200;
  assign \new_[27426]_  = ~A166 & \new_[27425]_ ;
  assign \new_[27427]_  = \new_[27426]_  & \new_[27421]_ ;
  assign \new_[27431]_  = A265 & A233;
  assign \new_[27432]_  = ~A232 & \new_[27431]_ ;
  assign \new_[27436]_  = A269 & A267;
  assign \new_[27437]_  = ~A266 & \new_[27436]_ ;
  assign \new_[27438]_  = \new_[27437]_  & \new_[27432]_ ;
  assign \new_[27442]_  = A167 & ~A169;
  assign \new_[27443]_  = A170 & \new_[27442]_ ;
  assign \new_[27447]_  = ~A201 & ~A200;
  assign \new_[27448]_  = ~A166 & \new_[27447]_ ;
  assign \new_[27449]_  = \new_[27448]_  & \new_[27443]_ ;
  assign \new_[27453]_  = A265 & ~A234;
  assign \new_[27454]_  = ~A233 & \new_[27453]_ ;
  assign \new_[27458]_  = A299 & ~A298;
  assign \new_[27459]_  = A266 & \new_[27458]_ ;
  assign \new_[27460]_  = \new_[27459]_  & \new_[27454]_ ;
  assign \new_[27464]_  = A167 & ~A169;
  assign \new_[27465]_  = A170 & \new_[27464]_ ;
  assign \new_[27469]_  = ~A201 & ~A200;
  assign \new_[27470]_  = ~A166 & \new_[27469]_ ;
  assign \new_[27471]_  = \new_[27470]_  & \new_[27465]_ ;
  assign \new_[27475]_  = ~A266 & ~A234;
  assign \new_[27476]_  = ~A233 & \new_[27475]_ ;
  assign \new_[27480]_  = A299 & ~A298;
  assign \new_[27481]_  = ~A267 & \new_[27480]_ ;
  assign \new_[27482]_  = \new_[27481]_  & \new_[27476]_ ;
  assign \new_[27486]_  = A167 & ~A169;
  assign \new_[27487]_  = A170 & \new_[27486]_ ;
  assign \new_[27491]_  = ~A201 & ~A200;
  assign \new_[27492]_  = ~A166 & \new_[27491]_ ;
  assign \new_[27493]_  = \new_[27492]_  & \new_[27487]_ ;
  assign \new_[27497]_  = ~A265 & ~A234;
  assign \new_[27498]_  = ~A233 & \new_[27497]_ ;
  assign \new_[27502]_  = A299 & ~A298;
  assign \new_[27503]_  = ~A266 & \new_[27502]_ ;
  assign \new_[27504]_  = \new_[27503]_  & \new_[27498]_ ;
  assign \new_[27508]_  = A167 & ~A169;
  assign \new_[27509]_  = A170 & \new_[27508]_ ;
  assign \new_[27513]_  = ~A201 & ~A200;
  assign \new_[27514]_  = ~A166 & \new_[27513]_ ;
  assign \new_[27515]_  = \new_[27514]_  & \new_[27509]_ ;
  assign \new_[27519]_  = A234 & ~A233;
  assign \new_[27520]_  = A232 & \new_[27519]_ ;
  assign \new_[27524]_  = ~A300 & A298;
  assign \new_[27525]_  = A235 & \new_[27524]_ ;
  assign \new_[27526]_  = \new_[27525]_  & \new_[27520]_ ;
  assign \new_[27530]_  = A167 & ~A169;
  assign \new_[27531]_  = A170 & \new_[27530]_ ;
  assign \new_[27535]_  = ~A201 & ~A200;
  assign \new_[27536]_  = ~A166 & \new_[27535]_ ;
  assign \new_[27537]_  = \new_[27536]_  & \new_[27531]_ ;
  assign \new_[27541]_  = A234 & ~A233;
  assign \new_[27542]_  = A232 & \new_[27541]_ ;
  assign \new_[27546]_  = A299 & A298;
  assign \new_[27547]_  = A235 & \new_[27546]_ ;
  assign \new_[27548]_  = \new_[27547]_  & \new_[27542]_ ;
  assign \new_[27552]_  = A167 & ~A169;
  assign \new_[27553]_  = A170 & \new_[27552]_ ;
  assign \new_[27557]_  = ~A201 & ~A200;
  assign \new_[27558]_  = ~A166 & \new_[27557]_ ;
  assign \new_[27559]_  = \new_[27558]_  & \new_[27553]_ ;
  assign \new_[27563]_  = A234 & ~A233;
  assign \new_[27564]_  = A232 & \new_[27563]_ ;
  assign \new_[27568]_  = ~A299 & ~A298;
  assign \new_[27569]_  = A235 & \new_[27568]_ ;
  assign \new_[27570]_  = \new_[27569]_  & \new_[27564]_ ;
  assign \new_[27574]_  = A167 & ~A169;
  assign \new_[27575]_  = A170 & \new_[27574]_ ;
  assign \new_[27579]_  = ~A201 & ~A200;
  assign \new_[27580]_  = ~A166 & \new_[27579]_ ;
  assign \new_[27581]_  = \new_[27580]_  & \new_[27575]_ ;
  assign \new_[27585]_  = A234 & ~A233;
  assign \new_[27586]_  = A232 & \new_[27585]_ ;
  assign \new_[27590]_  = A266 & ~A265;
  assign \new_[27591]_  = A235 & \new_[27590]_ ;
  assign \new_[27592]_  = \new_[27591]_  & \new_[27586]_ ;
  assign \new_[27596]_  = A167 & ~A169;
  assign \new_[27597]_  = A170 & \new_[27596]_ ;
  assign \new_[27601]_  = ~A201 & ~A200;
  assign \new_[27602]_  = ~A166 & \new_[27601]_ ;
  assign \new_[27603]_  = \new_[27602]_  & \new_[27597]_ ;
  assign \new_[27607]_  = A234 & ~A233;
  assign \new_[27608]_  = A232 & \new_[27607]_ ;
  assign \new_[27612]_  = ~A300 & A298;
  assign \new_[27613]_  = A236 & \new_[27612]_ ;
  assign \new_[27614]_  = \new_[27613]_  & \new_[27608]_ ;
  assign \new_[27618]_  = A167 & ~A169;
  assign \new_[27619]_  = A170 & \new_[27618]_ ;
  assign \new_[27623]_  = ~A201 & ~A200;
  assign \new_[27624]_  = ~A166 & \new_[27623]_ ;
  assign \new_[27625]_  = \new_[27624]_  & \new_[27619]_ ;
  assign \new_[27629]_  = A234 & ~A233;
  assign \new_[27630]_  = A232 & \new_[27629]_ ;
  assign \new_[27634]_  = A299 & A298;
  assign \new_[27635]_  = A236 & \new_[27634]_ ;
  assign \new_[27636]_  = \new_[27635]_  & \new_[27630]_ ;
  assign \new_[27640]_  = A167 & ~A169;
  assign \new_[27641]_  = A170 & \new_[27640]_ ;
  assign \new_[27645]_  = ~A201 & ~A200;
  assign \new_[27646]_  = ~A166 & \new_[27645]_ ;
  assign \new_[27647]_  = \new_[27646]_  & \new_[27641]_ ;
  assign \new_[27651]_  = A234 & ~A233;
  assign \new_[27652]_  = A232 & \new_[27651]_ ;
  assign \new_[27656]_  = ~A299 & ~A298;
  assign \new_[27657]_  = A236 & \new_[27656]_ ;
  assign \new_[27658]_  = \new_[27657]_  & \new_[27652]_ ;
  assign \new_[27662]_  = A167 & ~A169;
  assign \new_[27663]_  = A170 & \new_[27662]_ ;
  assign \new_[27667]_  = ~A201 & ~A200;
  assign \new_[27668]_  = ~A166 & \new_[27667]_ ;
  assign \new_[27669]_  = \new_[27668]_  & \new_[27663]_ ;
  assign \new_[27673]_  = A234 & ~A233;
  assign \new_[27674]_  = A232 & \new_[27673]_ ;
  assign \new_[27678]_  = A266 & ~A265;
  assign \new_[27679]_  = A236 & \new_[27678]_ ;
  assign \new_[27680]_  = \new_[27679]_  & \new_[27674]_ ;
  assign \new_[27684]_  = A167 & ~A169;
  assign \new_[27685]_  = A170 & \new_[27684]_ ;
  assign \new_[27689]_  = ~A201 & ~A200;
  assign \new_[27690]_  = ~A166 & \new_[27689]_ ;
  assign \new_[27691]_  = \new_[27690]_  & \new_[27685]_ ;
  assign \new_[27695]_  = A265 & ~A233;
  assign \new_[27696]_  = ~A232 & \new_[27695]_ ;
  assign \new_[27700]_  = A299 & ~A298;
  assign \new_[27701]_  = A266 & \new_[27700]_ ;
  assign \new_[27702]_  = \new_[27701]_  & \new_[27696]_ ;
  assign \new_[27706]_  = A167 & ~A169;
  assign \new_[27707]_  = A170 & \new_[27706]_ ;
  assign \new_[27711]_  = ~A201 & ~A200;
  assign \new_[27712]_  = ~A166 & \new_[27711]_ ;
  assign \new_[27713]_  = \new_[27712]_  & \new_[27707]_ ;
  assign \new_[27717]_  = ~A266 & ~A233;
  assign \new_[27718]_  = ~A232 & \new_[27717]_ ;
  assign \new_[27722]_  = A299 & ~A298;
  assign \new_[27723]_  = ~A267 & \new_[27722]_ ;
  assign \new_[27724]_  = \new_[27723]_  & \new_[27718]_ ;
  assign \new_[27728]_  = A167 & ~A169;
  assign \new_[27729]_  = A170 & \new_[27728]_ ;
  assign \new_[27733]_  = ~A201 & ~A200;
  assign \new_[27734]_  = ~A166 & \new_[27733]_ ;
  assign \new_[27735]_  = \new_[27734]_  & \new_[27729]_ ;
  assign \new_[27739]_  = ~A265 & ~A233;
  assign \new_[27740]_  = ~A232 & \new_[27739]_ ;
  assign \new_[27744]_  = A299 & ~A298;
  assign \new_[27745]_  = ~A266 & \new_[27744]_ ;
  assign \new_[27746]_  = \new_[27745]_  & \new_[27740]_ ;
  assign \new_[27750]_  = A167 & ~A169;
  assign \new_[27751]_  = A170 & \new_[27750]_ ;
  assign \new_[27755]_  = ~A200 & ~A199;
  assign \new_[27756]_  = ~A166 & \new_[27755]_ ;
  assign \new_[27757]_  = \new_[27756]_  & \new_[27751]_ ;
  assign \new_[27761]_  = A265 & A233;
  assign \new_[27762]_  = A232 & \new_[27761]_ ;
  assign \new_[27766]_  = A299 & ~A298;
  assign \new_[27767]_  = ~A267 & \new_[27766]_ ;
  assign \new_[27768]_  = \new_[27767]_  & \new_[27762]_ ;
  assign \new_[27772]_  = A167 & ~A169;
  assign \new_[27773]_  = A170 & \new_[27772]_ ;
  assign \new_[27777]_  = ~A200 & ~A199;
  assign \new_[27778]_  = ~A166 & \new_[27777]_ ;
  assign \new_[27779]_  = \new_[27778]_  & \new_[27773]_ ;
  assign \new_[27783]_  = A265 & A233;
  assign \new_[27784]_  = A232 & \new_[27783]_ ;
  assign \new_[27788]_  = A299 & ~A298;
  assign \new_[27789]_  = A266 & \new_[27788]_ ;
  assign \new_[27790]_  = \new_[27789]_  & \new_[27784]_ ;
  assign \new_[27794]_  = A167 & ~A169;
  assign \new_[27795]_  = A170 & \new_[27794]_ ;
  assign \new_[27799]_  = ~A200 & ~A199;
  assign \new_[27800]_  = ~A166 & \new_[27799]_ ;
  assign \new_[27801]_  = \new_[27800]_  & \new_[27795]_ ;
  assign \new_[27805]_  = ~A265 & A233;
  assign \new_[27806]_  = A232 & \new_[27805]_ ;
  assign \new_[27810]_  = A299 & ~A298;
  assign \new_[27811]_  = ~A266 & \new_[27810]_ ;
  assign \new_[27812]_  = \new_[27811]_  & \new_[27806]_ ;
  assign \new_[27816]_  = A167 & ~A169;
  assign \new_[27817]_  = A170 & \new_[27816]_ ;
  assign \new_[27821]_  = ~A200 & ~A199;
  assign \new_[27822]_  = ~A166 & \new_[27821]_ ;
  assign \new_[27823]_  = \new_[27822]_  & \new_[27817]_ ;
  assign \new_[27827]_  = A265 & A233;
  assign \new_[27828]_  = ~A232 & \new_[27827]_ ;
  assign \new_[27832]_  = A268 & A267;
  assign \new_[27833]_  = ~A266 & \new_[27832]_ ;
  assign \new_[27834]_  = \new_[27833]_  & \new_[27828]_ ;
  assign \new_[27838]_  = A167 & ~A169;
  assign \new_[27839]_  = A170 & \new_[27838]_ ;
  assign \new_[27843]_  = ~A200 & ~A199;
  assign \new_[27844]_  = ~A166 & \new_[27843]_ ;
  assign \new_[27845]_  = \new_[27844]_  & \new_[27839]_ ;
  assign \new_[27849]_  = A265 & A233;
  assign \new_[27850]_  = ~A232 & \new_[27849]_ ;
  assign \new_[27854]_  = A269 & A267;
  assign \new_[27855]_  = ~A266 & \new_[27854]_ ;
  assign \new_[27856]_  = \new_[27855]_  & \new_[27850]_ ;
  assign \new_[27860]_  = A167 & ~A169;
  assign \new_[27861]_  = A170 & \new_[27860]_ ;
  assign \new_[27865]_  = ~A200 & ~A199;
  assign \new_[27866]_  = ~A166 & \new_[27865]_ ;
  assign \new_[27867]_  = \new_[27866]_  & \new_[27861]_ ;
  assign \new_[27871]_  = A265 & ~A234;
  assign \new_[27872]_  = ~A233 & \new_[27871]_ ;
  assign \new_[27876]_  = A299 & ~A298;
  assign \new_[27877]_  = A266 & \new_[27876]_ ;
  assign \new_[27878]_  = \new_[27877]_  & \new_[27872]_ ;
  assign \new_[27882]_  = A167 & ~A169;
  assign \new_[27883]_  = A170 & \new_[27882]_ ;
  assign \new_[27887]_  = ~A200 & ~A199;
  assign \new_[27888]_  = ~A166 & \new_[27887]_ ;
  assign \new_[27889]_  = \new_[27888]_  & \new_[27883]_ ;
  assign \new_[27893]_  = ~A266 & ~A234;
  assign \new_[27894]_  = ~A233 & \new_[27893]_ ;
  assign \new_[27898]_  = A299 & ~A298;
  assign \new_[27899]_  = ~A267 & \new_[27898]_ ;
  assign \new_[27900]_  = \new_[27899]_  & \new_[27894]_ ;
  assign \new_[27904]_  = A167 & ~A169;
  assign \new_[27905]_  = A170 & \new_[27904]_ ;
  assign \new_[27909]_  = ~A200 & ~A199;
  assign \new_[27910]_  = ~A166 & \new_[27909]_ ;
  assign \new_[27911]_  = \new_[27910]_  & \new_[27905]_ ;
  assign \new_[27915]_  = ~A265 & ~A234;
  assign \new_[27916]_  = ~A233 & \new_[27915]_ ;
  assign \new_[27920]_  = A299 & ~A298;
  assign \new_[27921]_  = ~A266 & \new_[27920]_ ;
  assign \new_[27922]_  = \new_[27921]_  & \new_[27916]_ ;
  assign \new_[27926]_  = A167 & ~A169;
  assign \new_[27927]_  = A170 & \new_[27926]_ ;
  assign \new_[27931]_  = ~A200 & ~A199;
  assign \new_[27932]_  = ~A166 & \new_[27931]_ ;
  assign \new_[27933]_  = \new_[27932]_  & \new_[27927]_ ;
  assign \new_[27937]_  = A234 & ~A233;
  assign \new_[27938]_  = A232 & \new_[27937]_ ;
  assign \new_[27942]_  = ~A300 & A298;
  assign \new_[27943]_  = A235 & \new_[27942]_ ;
  assign \new_[27944]_  = \new_[27943]_  & \new_[27938]_ ;
  assign \new_[27948]_  = A167 & ~A169;
  assign \new_[27949]_  = A170 & \new_[27948]_ ;
  assign \new_[27953]_  = ~A200 & ~A199;
  assign \new_[27954]_  = ~A166 & \new_[27953]_ ;
  assign \new_[27955]_  = \new_[27954]_  & \new_[27949]_ ;
  assign \new_[27959]_  = A234 & ~A233;
  assign \new_[27960]_  = A232 & \new_[27959]_ ;
  assign \new_[27964]_  = A299 & A298;
  assign \new_[27965]_  = A235 & \new_[27964]_ ;
  assign \new_[27966]_  = \new_[27965]_  & \new_[27960]_ ;
  assign \new_[27970]_  = A167 & ~A169;
  assign \new_[27971]_  = A170 & \new_[27970]_ ;
  assign \new_[27975]_  = ~A200 & ~A199;
  assign \new_[27976]_  = ~A166 & \new_[27975]_ ;
  assign \new_[27977]_  = \new_[27976]_  & \new_[27971]_ ;
  assign \new_[27981]_  = A234 & ~A233;
  assign \new_[27982]_  = A232 & \new_[27981]_ ;
  assign \new_[27986]_  = ~A299 & ~A298;
  assign \new_[27987]_  = A235 & \new_[27986]_ ;
  assign \new_[27988]_  = \new_[27987]_  & \new_[27982]_ ;
  assign \new_[27992]_  = A167 & ~A169;
  assign \new_[27993]_  = A170 & \new_[27992]_ ;
  assign \new_[27997]_  = ~A200 & ~A199;
  assign \new_[27998]_  = ~A166 & \new_[27997]_ ;
  assign \new_[27999]_  = \new_[27998]_  & \new_[27993]_ ;
  assign \new_[28003]_  = A234 & ~A233;
  assign \new_[28004]_  = A232 & \new_[28003]_ ;
  assign \new_[28008]_  = A266 & ~A265;
  assign \new_[28009]_  = A235 & \new_[28008]_ ;
  assign \new_[28010]_  = \new_[28009]_  & \new_[28004]_ ;
  assign \new_[28014]_  = A167 & ~A169;
  assign \new_[28015]_  = A170 & \new_[28014]_ ;
  assign \new_[28019]_  = ~A200 & ~A199;
  assign \new_[28020]_  = ~A166 & \new_[28019]_ ;
  assign \new_[28021]_  = \new_[28020]_  & \new_[28015]_ ;
  assign \new_[28025]_  = A234 & ~A233;
  assign \new_[28026]_  = A232 & \new_[28025]_ ;
  assign \new_[28030]_  = ~A300 & A298;
  assign \new_[28031]_  = A236 & \new_[28030]_ ;
  assign \new_[28032]_  = \new_[28031]_  & \new_[28026]_ ;
  assign \new_[28036]_  = A167 & ~A169;
  assign \new_[28037]_  = A170 & \new_[28036]_ ;
  assign \new_[28041]_  = ~A200 & ~A199;
  assign \new_[28042]_  = ~A166 & \new_[28041]_ ;
  assign \new_[28043]_  = \new_[28042]_  & \new_[28037]_ ;
  assign \new_[28047]_  = A234 & ~A233;
  assign \new_[28048]_  = A232 & \new_[28047]_ ;
  assign \new_[28052]_  = A299 & A298;
  assign \new_[28053]_  = A236 & \new_[28052]_ ;
  assign \new_[28054]_  = \new_[28053]_  & \new_[28048]_ ;
  assign \new_[28058]_  = A167 & ~A169;
  assign \new_[28059]_  = A170 & \new_[28058]_ ;
  assign \new_[28063]_  = ~A200 & ~A199;
  assign \new_[28064]_  = ~A166 & \new_[28063]_ ;
  assign \new_[28065]_  = \new_[28064]_  & \new_[28059]_ ;
  assign \new_[28069]_  = A234 & ~A233;
  assign \new_[28070]_  = A232 & \new_[28069]_ ;
  assign \new_[28074]_  = ~A299 & ~A298;
  assign \new_[28075]_  = A236 & \new_[28074]_ ;
  assign \new_[28076]_  = \new_[28075]_  & \new_[28070]_ ;
  assign \new_[28080]_  = A167 & ~A169;
  assign \new_[28081]_  = A170 & \new_[28080]_ ;
  assign \new_[28085]_  = ~A200 & ~A199;
  assign \new_[28086]_  = ~A166 & \new_[28085]_ ;
  assign \new_[28087]_  = \new_[28086]_  & \new_[28081]_ ;
  assign \new_[28091]_  = A234 & ~A233;
  assign \new_[28092]_  = A232 & \new_[28091]_ ;
  assign \new_[28096]_  = A266 & ~A265;
  assign \new_[28097]_  = A236 & \new_[28096]_ ;
  assign \new_[28098]_  = \new_[28097]_  & \new_[28092]_ ;
  assign \new_[28102]_  = A167 & ~A169;
  assign \new_[28103]_  = A170 & \new_[28102]_ ;
  assign \new_[28107]_  = ~A200 & ~A199;
  assign \new_[28108]_  = ~A166 & \new_[28107]_ ;
  assign \new_[28109]_  = \new_[28108]_  & \new_[28103]_ ;
  assign \new_[28113]_  = A265 & ~A233;
  assign \new_[28114]_  = ~A232 & \new_[28113]_ ;
  assign \new_[28118]_  = A299 & ~A298;
  assign \new_[28119]_  = A266 & \new_[28118]_ ;
  assign \new_[28120]_  = \new_[28119]_  & \new_[28114]_ ;
  assign \new_[28124]_  = A167 & ~A169;
  assign \new_[28125]_  = A170 & \new_[28124]_ ;
  assign \new_[28129]_  = ~A200 & ~A199;
  assign \new_[28130]_  = ~A166 & \new_[28129]_ ;
  assign \new_[28131]_  = \new_[28130]_  & \new_[28125]_ ;
  assign \new_[28135]_  = ~A266 & ~A233;
  assign \new_[28136]_  = ~A232 & \new_[28135]_ ;
  assign \new_[28140]_  = A299 & ~A298;
  assign \new_[28141]_  = ~A267 & \new_[28140]_ ;
  assign \new_[28142]_  = \new_[28141]_  & \new_[28136]_ ;
  assign \new_[28146]_  = A167 & ~A169;
  assign \new_[28147]_  = A170 & \new_[28146]_ ;
  assign \new_[28151]_  = ~A200 & ~A199;
  assign \new_[28152]_  = ~A166 & \new_[28151]_ ;
  assign \new_[28153]_  = \new_[28152]_  & \new_[28147]_ ;
  assign \new_[28157]_  = ~A265 & ~A233;
  assign \new_[28158]_  = ~A232 & \new_[28157]_ ;
  assign \new_[28162]_  = A299 & ~A298;
  assign \new_[28163]_  = ~A266 & \new_[28162]_ ;
  assign \new_[28164]_  = \new_[28163]_  & \new_[28158]_ ;
  assign \new_[28168]_  = ~A167 & ~A169;
  assign \new_[28169]_  = A170 & \new_[28168]_ ;
  assign \new_[28173]_  = A200 & A199;
  assign \new_[28174]_  = A166 & \new_[28173]_ ;
  assign \new_[28175]_  = \new_[28174]_  & \new_[28169]_ ;
  assign \new_[28179]_  = A265 & A233;
  assign \new_[28180]_  = A232 & \new_[28179]_ ;
  assign \new_[28184]_  = A299 & ~A298;
  assign \new_[28185]_  = ~A267 & \new_[28184]_ ;
  assign \new_[28186]_  = \new_[28185]_  & \new_[28180]_ ;
  assign \new_[28190]_  = ~A167 & ~A169;
  assign \new_[28191]_  = A170 & \new_[28190]_ ;
  assign \new_[28195]_  = A200 & A199;
  assign \new_[28196]_  = A166 & \new_[28195]_ ;
  assign \new_[28197]_  = \new_[28196]_  & \new_[28191]_ ;
  assign \new_[28201]_  = A265 & A233;
  assign \new_[28202]_  = A232 & \new_[28201]_ ;
  assign \new_[28206]_  = A299 & ~A298;
  assign \new_[28207]_  = A266 & \new_[28206]_ ;
  assign \new_[28208]_  = \new_[28207]_  & \new_[28202]_ ;
  assign \new_[28212]_  = ~A167 & ~A169;
  assign \new_[28213]_  = A170 & \new_[28212]_ ;
  assign \new_[28217]_  = A200 & A199;
  assign \new_[28218]_  = A166 & \new_[28217]_ ;
  assign \new_[28219]_  = \new_[28218]_  & \new_[28213]_ ;
  assign \new_[28223]_  = ~A265 & A233;
  assign \new_[28224]_  = A232 & \new_[28223]_ ;
  assign \new_[28228]_  = A299 & ~A298;
  assign \new_[28229]_  = ~A266 & \new_[28228]_ ;
  assign \new_[28230]_  = \new_[28229]_  & \new_[28224]_ ;
  assign \new_[28234]_  = ~A167 & ~A169;
  assign \new_[28235]_  = A170 & \new_[28234]_ ;
  assign \new_[28239]_  = A200 & A199;
  assign \new_[28240]_  = A166 & \new_[28239]_ ;
  assign \new_[28241]_  = \new_[28240]_  & \new_[28235]_ ;
  assign \new_[28245]_  = A265 & A233;
  assign \new_[28246]_  = ~A232 & \new_[28245]_ ;
  assign \new_[28250]_  = A268 & A267;
  assign \new_[28251]_  = ~A266 & \new_[28250]_ ;
  assign \new_[28252]_  = \new_[28251]_  & \new_[28246]_ ;
  assign \new_[28256]_  = ~A167 & ~A169;
  assign \new_[28257]_  = A170 & \new_[28256]_ ;
  assign \new_[28261]_  = A200 & A199;
  assign \new_[28262]_  = A166 & \new_[28261]_ ;
  assign \new_[28263]_  = \new_[28262]_  & \new_[28257]_ ;
  assign \new_[28267]_  = A265 & A233;
  assign \new_[28268]_  = ~A232 & \new_[28267]_ ;
  assign \new_[28272]_  = A269 & A267;
  assign \new_[28273]_  = ~A266 & \new_[28272]_ ;
  assign \new_[28274]_  = \new_[28273]_  & \new_[28268]_ ;
  assign \new_[28278]_  = ~A167 & ~A169;
  assign \new_[28279]_  = A170 & \new_[28278]_ ;
  assign \new_[28283]_  = A200 & A199;
  assign \new_[28284]_  = A166 & \new_[28283]_ ;
  assign \new_[28285]_  = \new_[28284]_  & \new_[28279]_ ;
  assign \new_[28289]_  = A265 & ~A234;
  assign \new_[28290]_  = ~A233 & \new_[28289]_ ;
  assign \new_[28294]_  = A299 & ~A298;
  assign \new_[28295]_  = A266 & \new_[28294]_ ;
  assign \new_[28296]_  = \new_[28295]_  & \new_[28290]_ ;
  assign \new_[28300]_  = ~A167 & ~A169;
  assign \new_[28301]_  = A170 & \new_[28300]_ ;
  assign \new_[28305]_  = A200 & A199;
  assign \new_[28306]_  = A166 & \new_[28305]_ ;
  assign \new_[28307]_  = \new_[28306]_  & \new_[28301]_ ;
  assign \new_[28311]_  = ~A266 & ~A234;
  assign \new_[28312]_  = ~A233 & \new_[28311]_ ;
  assign \new_[28316]_  = A299 & ~A298;
  assign \new_[28317]_  = ~A267 & \new_[28316]_ ;
  assign \new_[28318]_  = \new_[28317]_  & \new_[28312]_ ;
  assign \new_[28322]_  = ~A167 & ~A169;
  assign \new_[28323]_  = A170 & \new_[28322]_ ;
  assign \new_[28327]_  = A200 & A199;
  assign \new_[28328]_  = A166 & \new_[28327]_ ;
  assign \new_[28329]_  = \new_[28328]_  & \new_[28323]_ ;
  assign \new_[28333]_  = ~A265 & ~A234;
  assign \new_[28334]_  = ~A233 & \new_[28333]_ ;
  assign \new_[28338]_  = A299 & ~A298;
  assign \new_[28339]_  = ~A266 & \new_[28338]_ ;
  assign \new_[28340]_  = \new_[28339]_  & \new_[28334]_ ;
  assign \new_[28344]_  = ~A167 & ~A169;
  assign \new_[28345]_  = A170 & \new_[28344]_ ;
  assign \new_[28349]_  = A200 & A199;
  assign \new_[28350]_  = A166 & \new_[28349]_ ;
  assign \new_[28351]_  = \new_[28350]_  & \new_[28345]_ ;
  assign \new_[28355]_  = A234 & ~A233;
  assign \new_[28356]_  = A232 & \new_[28355]_ ;
  assign \new_[28360]_  = ~A300 & A298;
  assign \new_[28361]_  = A235 & \new_[28360]_ ;
  assign \new_[28362]_  = \new_[28361]_  & \new_[28356]_ ;
  assign \new_[28366]_  = ~A167 & ~A169;
  assign \new_[28367]_  = A170 & \new_[28366]_ ;
  assign \new_[28371]_  = A200 & A199;
  assign \new_[28372]_  = A166 & \new_[28371]_ ;
  assign \new_[28373]_  = \new_[28372]_  & \new_[28367]_ ;
  assign \new_[28377]_  = A234 & ~A233;
  assign \new_[28378]_  = A232 & \new_[28377]_ ;
  assign \new_[28382]_  = A299 & A298;
  assign \new_[28383]_  = A235 & \new_[28382]_ ;
  assign \new_[28384]_  = \new_[28383]_  & \new_[28378]_ ;
  assign \new_[28388]_  = ~A167 & ~A169;
  assign \new_[28389]_  = A170 & \new_[28388]_ ;
  assign \new_[28393]_  = A200 & A199;
  assign \new_[28394]_  = A166 & \new_[28393]_ ;
  assign \new_[28395]_  = \new_[28394]_  & \new_[28389]_ ;
  assign \new_[28399]_  = A234 & ~A233;
  assign \new_[28400]_  = A232 & \new_[28399]_ ;
  assign \new_[28404]_  = ~A299 & ~A298;
  assign \new_[28405]_  = A235 & \new_[28404]_ ;
  assign \new_[28406]_  = \new_[28405]_  & \new_[28400]_ ;
  assign \new_[28410]_  = ~A167 & ~A169;
  assign \new_[28411]_  = A170 & \new_[28410]_ ;
  assign \new_[28415]_  = A200 & A199;
  assign \new_[28416]_  = A166 & \new_[28415]_ ;
  assign \new_[28417]_  = \new_[28416]_  & \new_[28411]_ ;
  assign \new_[28421]_  = A234 & ~A233;
  assign \new_[28422]_  = A232 & \new_[28421]_ ;
  assign \new_[28426]_  = A266 & ~A265;
  assign \new_[28427]_  = A235 & \new_[28426]_ ;
  assign \new_[28428]_  = \new_[28427]_  & \new_[28422]_ ;
  assign \new_[28432]_  = ~A167 & ~A169;
  assign \new_[28433]_  = A170 & \new_[28432]_ ;
  assign \new_[28437]_  = A200 & A199;
  assign \new_[28438]_  = A166 & \new_[28437]_ ;
  assign \new_[28439]_  = \new_[28438]_  & \new_[28433]_ ;
  assign \new_[28443]_  = A234 & ~A233;
  assign \new_[28444]_  = A232 & \new_[28443]_ ;
  assign \new_[28448]_  = ~A300 & A298;
  assign \new_[28449]_  = A236 & \new_[28448]_ ;
  assign \new_[28450]_  = \new_[28449]_  & \new_[28444]_ ;
  assign \new_[28454]_  = ~A167 & ~A169;
  assign \new_[28455]_  = A170 & \new_[28454]_ ;
  assign \new_[28459]_  = A200 & A199;
  assign \new_[28460]_  = A166 & \new_[28459]_ ;
  assign \new_[28461]_  = \new_[28460]_  & \new_[28455]_ ;
  assign \new_[28465]_  = A234 & ~A233;
  assign \new_[28466]_  = A232 & \new_[28465]_ ;
  assign \new_[28470]_  = A299 & A298;
  assign \new_[28471]_  = A236 & \new_[28470]_ ;
  assign \new_[28472]_  = \new_[28471]_  & \new_[28466]_ ;
  assign \new_[28476]_  = ~A167 & ~A169;
  assign \new_[28477]_  = A170 & \new_[28476]_ ;
  assign \new_[28481]_  = A200 & A199;
  assign \new_[28482]_  = A166 & \new_[28481]_ ;
  assign \new_[28483]_  = \new_[28482]_  & \new_[28477]_ ;
  assign \new_[28487]_  = A234 & ~A233;
  assign \new_[28488]_  = A232 & \new_[28487]_ ;
  assign \new_[28492]_  = ~A299 & ~A298;
  assign \new_[28493]_  = A236 & \new_[28492]_ ;
  assign \new_[28494]_  = \new_[28493]_  & \new_[28488]_ ;
  assign \new_[28498]_  = ~A167 & ~A169;
  assign \new_[28499]_  = A170 & \new_[28498]_ ;
  assign \new_[28503]_  = A200 & A199;
  assign \new_[28504]_  = A166 & \new_[28503]_ ;
  assign \new_[28505]_  = \new_[28504]_  & \new_[28499]_ ;
  assign \new_[28509]_  = A234 & ~A233;
  assign \new_[28510]_  = A232 & \new_[28509]_ ;
  assign \new_[28514]_  = A266 & ~A265;
  assign \new_[28515]_  = A236 & \new_[28514]_ ;
  assign \new_[28516]_  = \new_[28515]_  & \new_[28510]_ ;
  assign \new_[28520]_  = ~A167 & ~A169;
  assign \new_[28521]_  = A170 & \new_[28520]_ ;
  assign \new_[28525]_  = A200 & A199;
  assign \new_[28526]_  = A166 & \new_[28525]_ ;
  assign \new_[28527]_  = \new_[28526]_  & \new_[28521]_ ;
  assign \new_[28531]_  = A265 & ~A233;
  assign \new_[28532]_  = ~A232 & \new_[28531]_ ;
  assign \new_[28536]_  = A299 & ~A298;
  assign \new_[28537]_  = A266 & \new_[28536]_ ;
  assign \new_[28538]_  = \new_[28537]_  & \new_[28532]_ ;
  assign \new_[28542]_  = ~A167 & ~A169;
  assign \new_[28543]_  = A170 & \new_[28542]_ ;
  assign \new_[28547]_  = A200 & A199;
  assign \new_[28548]_  = A166 & \new_[28547]_ ;
  assign \new_[28549]_  = \new_[28548]_  & \new_[28543]_ ;
  assign \new_[28553]_  = ~A266 & ~A233;
  assign \new_[28554]_  = ~A232 & \new_[28553]_ ;
  assign \new_[28558]_  = A299 & ~A298;
  assign \new_[28559]_  = ~A267 & \new_[28558]_ ;
  assign \new_[28560]_  = \new_[28559]_  & \new_[28554]_ ;
  assign \new_[28564]_  = ~A167 & ~A169;
  assign \new_[28565]_  = A170 & \new_[28564]_ ;
  assign \new_[28569]_  = A200 & A199;
  assign \new_[28570]_  = A166 & \new_[28569]_ ;
  assign \new_[28571]_  = \new_[28570]_  & \new_[28565]_ ;
  assign \new_[28575]_  = ~A265 & ~A233;
  assign \new_[28576]_  = ~A232 & \new_[28575]_ ;
  assign \new_[28580]_  = A299 & ~A298;
  assign \new_[28581]_  = ~A266 & \new_[28580]_ ;
  assign \new_[28582]_  = \new_[28581]_  & \new_[28576]_ ;
  assign \new_[28586]_  = ~A167 & ~A169;
  assign \new_[28587]_  = A170 & \new_[28586]_ ;
  assign \new_[28591]_  = ~A202 & ~A200;
  assign \new_[28592]_  = A166 & \new_[28591]_ ;
  assign \new_[28593]_  = \new_[28592]_  & \new_[28587]_ ;
  assign \new_[28597]_  = A233 & ~A232;
  assign \new_[28598]_  = ~A203 & \new_[28597]_ ;
  assign \new_[28602]_  = ~A302 & ~A301;
  assign \new_[28603]_  = ~A299 & \new_[28602]_ ;
  assign \new_[28604]_  = \new_[28603]_  & \new_[28598]_ ;
  assign \new_[28608]_  = ~A167 & ~A169;
  assign \new_[28609]_  = A170 & \new_[28608]_ ;
  assign \new_[28613]_  = ~A201 & ~A200;
  assign \new_[28614]_  = A166 & \new_[28613]_ ;
  assign \new_[28615]_  = \new_[28614]_  & \new_[28609]_ ;
  assign \new_[28619]_  = A265 & A233;
  assign \new_[28620]_  = A232 & \new_[28619]_ ;
  assign \new_[28624]_  = A299 & ~A298;
  assign \new_[28625]_  = ~A267 & \new_[28624]_ ;
  assign \new_[28626]_  = \new_[28625]_  & \new_[28620]_ ;
  assign \new_[28630]_  = ~A167 & ~A169;
  assign \new_[28631]_  = A170 & \new_[28630]_ ;
  assign \new_[28635]_  = ~A201 & ~A200;
  assign \new_[28636]_  = A166 & \new_[28635]_ ;
  assign \new_[28637]_  = \new_[28636]_  & \new_[28631]_ ;
  assign \new_[28641]_  = A265 & A233;
  assign \new_[28642]_  = A232 & \new_[28641]_ ;
  assign \new_[28646]_  = A299 & ~A298;
  assign \new_[28647]_  = A266 & \new_[28646]_ ;
  assign \new_[28648]_  = \new_[28647]_  & \new_[28642]_ ;
  assign \new_[28652]_  = ~A167 & ~A169;
  assign \new_[28653]_  = A170 & \new_[28652]_ ;
  assign \new_[28657]_  = ~A201 & ~A200;
  assign \new_[28658]_  = A166 & \new_[28657]_ ;
  assign \new_[28659]_  = \new_[28658]_  & \new_[28653]_ ;
  assign \new_[28663]_  = ~A265 & A233;
  assign \new_[28664]_  = A232 & \new_[28663]_ ;
  assign \new_[28668]_  = A299 & ~A298;
  assign \new_[28669]_  = ~A266 & \new_[28668]_ ;
  assign \new_[28670]_  = \new_[28669]_  & \new_[28664]_ ;
  assign \new_[28674]_  = ~A167 & ~A169;
  assign \new_[28675]_  = A170 & \new_[28674]_ ;
  assign \new_[28679]_  = ~A201 & ~A200;
  assign \new_[28680]_  = A166 & \new_[28679]_ ;
  assign \new_[28681]_  = \new_[28680]_  & \new_[28675]_ ;
  assign \new_[28685]_  = A265 & A233;
  assign \new_[28686]_  = ~A232 & \new_[28685]_ ;
  assign \new_[28690]_  = A268 & A267;
  assign \new_[28691]_  = ~A266 & \new_[28690]_ ;
  assign \new_[28692]_  = \new_[28691]_  & \new_[28686]_ ;
  assign \new_[28696]_  = ~A167 & ~A169;
  assign \new_[28697]_  = A170 & \new_[28696]_ ;
  assign \new_[28701]_  = ~A201 & ~A200;
  assign \new_[28702]_  = A166 & \new_[28701]_ ;
  assign \new_[28703]_  = \new_[28702]_  & \new_[28697]_ ;
  assign \new_[28707]_  = A265 & A233;
  assign \new_[28708]_  = ~A232 & \new_[28707]_ ;
  assign \new_[28712]_  = A269 & A267;
  assign \new_[28713]_  = ~A266 & \new_[28712]_ ;
  assign \new_[28714]_  = \new_[28713]_  & \new_[28708]_ ;
  assign \new_[28718]_  = ~A167 & ~A169;
  assign \new_[28719]_  = A170 & \new_[28718]_ ;
  assign \new_[28723]_  = ~A201 & ~A200;
  assign \new_[28724]_  = A166 & \new_[28723]_ ;
  assign \new_[28725]_  = \new_[28724]_  & \new_[28719]_ ;
  assign \new_[28729]_  = A265 & ~A234;
  assign \new_[28730]_  = ~A233 & \new_[28729]_ ;
  assign \new_[28734]_  = A299 & ~A298;
  assign \new_[28735]_  = A266 & \new_[28734]_ ;
  assign \new_[28736]_  = \new_[28735]_  & \new_[28730]_ ;
  assign \new_[28740]_  = ~A167 & ~A169;
  assign \new_[28741]_  = A170 & \new_[28740]_ ;
  assign \new_[28745]_  = ~A201 & ~A200;
  assign \new_[28746]_  = A166 & \new_[28745]_ ;
  assign \new_[28747]_  = \new_[28746]_  & \new_[28741]_ ;
  assign \new_[28751]_  = ~A266 & ~A234;
  assign \new_[28752]_  = ~A233 & \new_[28751]_ ;
  assign \new_[28756]_  = A299 & ~A298;
  assign \new_[28757]_  = ~A267 & \new_[28756]_ ;
  assign \new_[28758]_  = \new_[28757]_  & \new_[28752]_ ;
  assign \new_[28762]_  = ~A167 & ~A169;
  assign \new_[28763]_  = A170 & \new_[28762]_ ;
  assign \new_[28767]_  = ~A201 & ~A200;
  assign \new_[28768]_  = A166 & \new_[28767]_ ;
  assign \new_[28769]_  = \new_[28768]_  & \new_[28763]_ ;
  assign \new_[28773]_  = ~A265 & ~A234;
  assign \new_[28774]_  = ~A233 & \new_[28773]_ ;
  assign \new_[28778]_  = A299 & ~A298;
  assign \new_[28779]_  = ~A266 & \new_[28778]_ ;
  assign \new_[28780]_  = \new_[28779]_  & \new_[28774]_ ;
  assign \new_[28784]_  = ~A167 & ~A169;
  assign \new_[28785]_  = A170 & \new_[28784]_ ;
  assign \new_[28789]_  = ~A201 & ~A200;
  assign \new_[28790]_  = A166 & \new_[28789]_ ;
  assign \new_[28791]_  = \new_[28790]_  & \new_[28785]_ ;
  assign \new_[28795]_  = A234 & ~A233;
  assign \new_[28796]_  = A232 & \new_[28795]_ ;
  assign \new_[28800]_  = ~A300 & A298;
  assign \new_[28801]_  = A235 & \new_[28800]_ ;
  assign \new_[28802]_  = \new_[28801]_  & \new_[28796]_ ;
  assign \new_[28806]_  = ~A167 & ~A169;
  assign \new_[28807]_  = A170 & \new_[28806]_ ;
  assign \new_[28811]_  = ~A201 & ~A200;
  assign \new_[28812]_  = A166 & \new_[28811]_ ;
  assign \new_[28813]_  = \new_[28812]_  & \new_[28807]_ ;
  assign \new_[28817]_  = A234 & ~A233;
  assign \new_[28818]_  = A232 & \new_[28817]_ ;
  assign \new_[28822]_  = A299 & A298;
  assign \new_[28823]_  = A235 & \new_[28822]_ ;
  assign \new_[28824]_  = \new_[28823]_  & \new_[28818]_ ;
  assign \new_[28828]_  = ~A167 & ~A169;
  assign \new_[28829]_  = A170 & \new_[28828]_ ;
  assign \new_[28833]_  = ~A201 & ~A200;
  assign \new_[28834]_  = A166 & \new_[28833]_ ;
  assign \new_[28835]_  = \new_[28834]_  & \new_[28829]_ ;
  assign \new_[28839]_  = A234 & ~A233;
  assign \new_[28840]_  = A232 & \new_[28839]_ ;
  assign \new_[28844]_  = ~A299 & ~A298;
  assign \new_[28845]_  = A235 & \new_[28844]_ ;
  assign \new_[28846]_  = \new_[28845]_  & \new_[28840]_ ;
  assign \new_[28850]_  = ~A167 & ~A169;
  assign \new_[28851]_  = A170 & \new_[28850]_ ;
  assign \new_[28855]_  = ~A201 & ~A200;
  assign \new_[28856]_  = A166 & \new_[28855]_ ;
  assign \new_[28857]_  = \new_[28856]_  & \new_[28851]_ ;
  assign \new_[28861]_  = A234 & ~A233;
  assign \new_[28862]_  = A232 & \new_[28861]_ ;
  assign \new_[28866]_  = A266 & ~A265;
  assign \new_[28867]_  = A235 & \new_[28866]_ ;
  assign \new_[28868]_  = \new_[28867]_  & \new_[28862]_ ;
  assign \new_[28872]_  = ~A167 & ~A169;
  assign \new_[28873]_  = A170 & \new_[28872]_ ;
  assign \new_[28877]_  = ~A201 & ~A200;
  assign \new_[28878]_  = A166 & \new_[28877]_ ;
  assign \new_[28879]_  = \new_[28878]_  & \new_[28873]_ ;
  assign \new_[28883]_  = A234 & ~A233;
  assign \new_[28884]_  = A232 & \new_[28883]_ ;
  assign \new_[28888]_  = ~A300 & A298;
  assign \new_[28889]_  = A236 & \new_[28888]_ ;
  assign \new_[28890]_  = \new_[28889]_  & \new_[28884]_ ;
  assign \new_[28894]_  = ~A167 & ~A169;
  assign \new_[28895]_  = A170 & \new_[28894]_ ;
  assign \new_[28899]_  = ~A201 & ~A200;
  assign \new_[28900]_  = A166 & \new_[28899]_ ;
  assign \new_[28901]_  = \new_[28900]_  & \new_[28895]_ ;
  assign \new_[28905]_  = A234 & ~A233;
  assign \new_[28906]_  = A232 & \new_[28905]_ ;
  assign \new_[28910]_  = A299 & A298;
  assign \new_[28911]_  = A236 & \new_[28910]_ ;
  assign \new_[28912]_  = \new_[28911]_  & \new_[28906]_ ;
  assign \new_[28916]_  = ~A167 & ~A169;
  assign \new_[28917]_  = A170 & \new_[28916]_ ;
  assign \new_[28921]_  = ~A201 & ~A200;
  assign \new_[28922]_  = A166 & \new_[28921]_ ;
  assign \new_[28923]_  = \new_[28922]_  & \new_[28917]_ ;
  assign \new_[28927]_  = A234 & ~A233;
  assign \new_[28928]_  = A232 & \new_[28927]_ ;
  assign \new_[28932]_  = ~A299 & ~A298;
  assign \new_[28933]_  = A236 & \new_[28932]_ ;
  assign \new_[28934]_  = \new_[28933]_  & \new_[28928]_ ;
  assign \new_[28938]_  = ~A167 & ~A169;
  assign \new_[28939]_  = A170 & \new_[28938]_ ;
  assign \new_[28943]_  = ~A201 & ~A200;
  assign \new_[28944]_  = A166 & \new_[28943]_ ;
  assign \new_[28945]_  = \new_[28944]_  & \new_[28939]_ ;
  assign \new_[28949]_  = A234 & ~A233;
  assign \new_[28950]_  = A232 & \new_[28949]_ ;
  assign \new_[28954]_  = A266 & ~A265;
  assign \new_[28955]_  = A236 & \new_[28954]_ ;
  assign \new_[28956]_  = \new_[28955]_  & \new_[28950]_ ;
  assign \new_[28960]_  = ~A167 & ~A169;
  assign \new_[28961]_  = A170 & \new_[28960]_ ;
  assign \new_[28965]_  = ~A201 & ~A200;
  assign \new_[28966]_  = A166 & \new_[28965]_ ;
  assign \new_[28967]_  = \new_[28966]_  & \new_[28961]_ ;
  assign \new_[28971]_  = A265 & ~A233;
  assign \new_[28972]_  = ~A232 & \new_[28971]_ ;
  assign \new_[28976]_  = A299 & ~A298;
  assign \new_[28977]_  = A266 & \new_[28976]_ ;
  assign \new_[28978]_  = \new_[28977]_  & \new_[28972]_ ;
  assign \new_[28982]_  = ~A167 & ~A169;
  assign \new_[28983]_  = A170 & \new_[28982]_ ;
  assign \new_[28987]_  = ~A201 & ~A200;
  assign \new_[28988]_  = A166 & \new_[28987]_ ;
  assign \new_[28989]_  = \new_[28988]_  & \new_[28983]_ ;
  assign \new_[28993]_  = ~A266 & ~A233;
  assign \new_[28994]_  = ~A232 & \new_[28993]_ ;
  assign \new_[28998]_  = A299 & ~A298;
  assign \new_[28999]_  = ~A267 & \new_[28998]_ ;
  assign \new_[29000]_  = \new_[28999]_  & \new_[28994]_ ;
  assign \new_[29004]_  = ~A167 & ~A169;
  assign \new_[29005]_  = A170 & \new_[29004]_ ;
  assign \new_[29009]_  = ~A201 & ~A200;
  assign \new_[29010]_  = A166 & \new_[29009]_ ;
  assign \new_[29011]_  = \new_[29010]_  & \new_[29005]_ ;
  assign \new_[29015]_  = ~A265 & ~A233;
  assign \new_[29016]_  = ~A232 & \new_[29015]_ ;
  assign \new_[29020]_  = A299 & ~A298;
  assign \new_[29021]_  = ~A266 & \new_[29020]_ ;
  assign \new_[29022]_  = \new_[29021]_  & \new_[29016]_ ;
  assign \new_[29026]_  = ~A167 & ~A169;
  assign \new_[29027]_  = A170 & \new_[29026]_ ;
  assign \new_[29031]_  = ~A200 & ~A199;
  assign \new_[29032]_  = A166 & \new_[29031]_ ;
  assign \new_[29033]_  = \new_[29032]_  & \new_[29027]_ ;
  assign \new_[29037]_  = A265 & A233;
  assign \new_[29038]_  = A232 & \new_[29037]_ ;
  assign \new_[29042]_  = A299 & ~A298;
  assign \new_[29043]_  = ~A267 & \new_[29042]_ ;
  assign \new_[29044]_  = \new_[29043]_  & \new_[29038]_ ;
  assign \new_[29048]_  = ~A167 & ~A169;
  assign \new_[29049]_  = A170 & \new_[29048]_ ;
  assign \new_[29053]_  = ~A200 & ~A199;
  assign \new_[29054]_  = A166 & \new_[29053]_ ;
  assign \new_[29055]_  = \new_[29054]_  & \new_[29049]_ ;
  assign \new_[29059]_  = A265 & A233;
  assign \new_[29060]_  = A232 & \new_[29059]_ ;
  assign \new_[29064]_  = A299 & ~A298;
  assign \new_[29065]_  = A266 & \new_[29064]_ ;
  assign \new_[29066]_  = \new_[29065]_  & \new_[29060]_ ;
  assign \new_[29070]_  = ~A167 & ~A169;
  assign \new_[29071]_  = A170 & \new_[29070]_ ;
  assign \new_[29075]_  = ~A200 & ~A199;
  assign \new_[29076]_  = A166 & \new_[29075]_ ;
  assign \new_[29077]_  = \new_[29076]_  & \new_[29071]_ ;
  assign \new_[29081]_  = ~A265 & A233;
  assign \new_[29082]_  = A232 & \new_[29081]_ ;
  assign \new_[29086]_  = A299 & ~A298;
  assign \new_[29087]_  = ~A266 & \new_[29086]_ ;
  assign \new_[29088]_  = \new_[29087]_  & \new_[29082]_ ;
  assign \new_[29092]_  = ~A167 & ~A169;
  assign \new_[29093]_  = A170 & \new_[29092]_ ;
  assign \new_[29097]_  = ~A200 & ~A199;
  assign \new_[29098]_  = A166 & \new_[29097]_ ;
  assign \new_[29099]_  = \new_[29098]_  & \new_[29093]_ ;
  assign \new_[29103]_  = A265 & A233;
  assign \new_[29104]_  = ~A232 & \new_[29103]_ ;
  assign \new_[29108]_  = A268 & A267;
  assign \new_[29109]_  = ~A266 & \new_[29108]_ ;
  assign \new_[29110]_  = \new_[29109]_  & \new_[29104]_ ;
  assign \new_[29114]_  = ~A167 & ~A169;
  assign \new_[29115]_  = A170 & \new_[29114]_ ;
  assign \new_[29119]_  = ~A200 & ~A199;
  assign \new_[29120]_  = A166 & \new_[29119]_ ;
  assign \new_[29121]_  = \new_[29120]_  & \new_[29115]_ ;
  assign \new_[29125]_  = A265 & A233;
  assign \new_[29126]_  = ~A232 & \new_[29125]_ ;
  assign \new_[29130]_  = A269 & A267;
  assign \new_[29131]_  = ~A266 & \new_[29130]_ ;
  assign \new_[29132]_  = \new_[29131]_  & \new_[29126]_ ;
  assign \new_[29136]_  = ~A167 & ~A169;
  assign \new_[29137]_  = A170 & \new_[29136]_ ;
  assign \new_[29141]_  = ~A200 & ~A199;
  assign \new_[29142]_  = A166 & \new_[29141]_ ;
  assign \new_[29143]_  = \new_[29142]_  & \new_[29137]_ ;
  assign \new_[29147]_  = A265 & ~A234;
  assign \new_[29148]_  = ~A233 & \new_[29147]_ ;
  assign \new_[29152]_  = A299 & ~A298;
  assign \new_[29153]_  = A266 & \new_[29152]_ ;
  assign \new_[29154]_  = \new_[29153]_  & \new_[29148]_ ;
  assign \new_[29158]_  = ~A167 & ~A169;
  assign \new_[29159]_  = A170 & \new_[29158]_ ;
  assign \new_[29163]_  = ~A200 & ~A199;
  assign \new_[29164]_  = A166 & \new_[29163]_ ;
  assign \new_[29165]_  = \new_[29164]_  & \new_[29159]_ ;
  assign \new_[29169]_  = ~A266 & ~A234;
  assign \new_[29170]_  = ~A233 & \new_[29169]_ ;
  assign \new_[29174]_  = A299 & ~A298;
  assign \new_[29175]_  = ~A267 & \new_[29174]_ ;
  assign \new_[29176]_  = \new_[29175]_  & \new_[29170]_ ;
  assign \new_[29180]_  = ~A167 & ~A169;
  assign \new_[29181]_  = A170 & \new_[29180]_ ;
  assign \new_[29185]_  = ~A200 & ~A199;
  assign \new_[29186]_  = A166 & \new_[29185]_ ;
  assign \new_[29187]_  = \new_[29186]_  & \new_[29181]_ ;
  assign \new_[29191]_  = ~A265 & ~A234;
  assign \new_[29192]_  = ~A233 & \new_[29191]_ ;
  assign \new_[29196]_  = A299 & ~A298;
  assign \new_[29197]_  = ~A266 & \new_[29196]_ ;
  assign \new_[29198]_  = \new_[29197]_  & \new_[29192]_ ;
  assign \new_[29202]_  = ~A167 & ~A169;
  assign \new_[29203]_  = A170 & \new_[29202]_ ;
  assign \new_[29207]_  = ~A200 & ~A199;
  assign \new_[29208]_  = A166 & \new_[29207]_ ;
  assign \new_[29209]_  = \new_[29208]_  & \new_[29203]_ ;
  assign \new_[29213]_  = A234 & ~A233;
  assign \new_[29214]_  = A232 & \new_[29213]_ ;
  assign \new_[29218]_  = ~A300 & A298;
  assign \new_[29219]_  = A235 & \new_[29218]_ ;
  assign \new_[29220]_  = \new_[29219]_  & \new_[29214]_ ;
  assign \new_[29224]_  = ~A167 & ~A169;
  assign \new_[29225]_  = A170 & \new_[29224]_ ;
  assign \new_[29229]_  = ~A200 & ~A199;
  assign \new_[29230]_  = A166 & \new_[29229]_ ;
  assign \new_[29231]_  = \new_[29230]_  & \new_[29225]_ ;
  assign \new_[29235]_  = A234 & ~A233;
  assign \new_[29236]_  = A232 & \new_[29235]_ ;
  assign \new_[29240]_  = A299 & A298;
  assign \new_[29241]_  = A235 & \new_[29240]_ ;
  assign \new_[29242]_  = \new_[29241]_  & \new_[29236]_ ;
  assign \new_[29246]_  = ~A167 & ~A169;
  assign \new_[29247]_  = A170 & \new_[29246]_ ;
  assign \new_[29251]_  = ~A200 & ~A199;
  assign \new_[29252]_  = A166 & \new_[29251]_ ;
  assign \new_[29253]_  = \new_[29252]_  & \new_[29247]_ ;
  assign \new_[29257]_  = A234 & ~A233;
  assign \new_[29258]_  = A232 & \new_[29257]_ ;
  assign \new_[29262]_  = ~A299 & ~A298;
  assign \new_[29263]_  = A235 & \new_[29262]_ ;
  assign \new_[29264]_  = \new_[29263]_  & \new_[29258]_ ;
  assign \new_[29268]_  = ~A167 & ~A169;
  assign \new_[29269]_  = A170 & \new_[29268]_ ;
  assign \new_[29273]_  = ~A200 & ~A199;
  assign \new_[29274]_  = A166 & \new_[29273]_ ;
  assign \new_[29275]_  = \new_[29274]_  & \new_[29269]_ ;
  assign \new_[29279]_  = A234 & ~A233;
  assign \new_[29280]_  = A232 & \new_[29279]_ ;
  assign \new_[29284]_  = A266 & ~A265;
  assign \new_[29285]_  = A235 & \new_[29284]_ ;
  assign \new_[29286]_  = \new_[29285]_  & \new_[29280]_ ;
  assign \new_[29290]_  = ~A167 & ~A169;
  assign \new_[29291]_  = A170 & \new_[29290]_ ;
  assign \new_[29295]_  = ~A200 & ~A199;
  assign \new_[29296]_  = A166 & \new_[29295]_ ;
  assign \new_[29297]_  = \new_[29296]_  & \new_[29291]_ ;
  assign \new_[29301]_  = A234 & ~A233;
  assign \new_[29302]_  = A232 & \new_[29301]_ ;
  assign \new_[29306]_  = ~A300 & A298;
  assign \new_[29307]_  = A236 & \new_[29306]_ ;
  assign \new_[29308]_  = \new_[29307]_  & \new_[29302]_ ;
  assign \new_[29312]_  = ~A167 & ~A169;
  assign \new_[29313]_  = A170 & \new_[29312]_ ;
  assign \new_[29317]_  = ~A200 & ~A199;
  assign \new_[29318]_  = A166 & \new_[29317]_ ;
  assign \new_[29319]_  = \new_[29318]_  & \new_[29313]_ ;
  assign \new_[29323]_  = A234 & ~A233;
  assign \new_[29324]_  = A232 & \new_[29323]_ ;
  assign \new_[29328]_  = A299 & A298;
  assign \new_[29329]_  = A236 & \new_[29328]_ ;
  assign \new_[29330]_  = \new_[29329]_  & \new_[29324]_ ;
  assign \new_[29334]_  = ~A167 & ~A169;
  assign \new_[29335]_  = A170 & \new_[29334]_ ;
  assign \new_[29339]_  = ~A200 & ~A199;
  assign \new_[29340]_  = A166 & \new_[29339]_ ;
  assign \new_[29341]_  = \new_[29340]_  & \new_[29335]_ ;
  assign \new_[29345]_  = A234 & ~A233;
  assign \new_[29346]_  = A232 & \new_[29345]_ ;
  assign \new_[29350]_  = ~A299 & ~A298;
  assign \new_[29351]_  = A236 & \new_[29350]_ ;
  assign \new_[29352]_  = \new_[29351]_  & \new_[29346]_ ;
  assign \new_[29356]_  = ~A167 & ~A169;
  assign \new_[29357]_  = A170 & \new_[29356]_ ;
  assign \new_[29361]_  = ~A200 & ~A199;
  assign \new_[29362]_  = A166 & \new_[29361]_ ;
  assign \new_[29363]_  = \new_[29362]_  & \new_[29357]_ ;
  assign \new_[29367]_  = A234 & ~A233;
  assign \new_[29368]_  = A232 & \new_[29367]_ ;
  assign \new_[29372]_  = A266 & ~A265;
  assign \new_[29373]_  = A236 & \new_[29372]_ ;
  assign \new_[29374]_  = \new_[29373]_  & \new_[29368]_ ;
  assign \new_[29378]_  = ~A167 & ~A169;
  assign \new_[29379]_  = A170 & \new_[29378]_ ;
  assign \new_[29383]_  = ~A200 & ~A199;
  assign \new_[29384]_  = A166 & \new_[29383]_ ;
  assign \new_[29385]_  = \new_[29384]_  & \new_[29379]_ ;
  assign \new_[29389]_  = A265 & ~A233;
  assign \new_[29390]_  = ~A232 & \new_[29389]_ ;
  assign \new_[29394]_  = A299 & ~A298;
  assign \new_[29395]_  = A266 & \new_[29394]_ ;
  assign \new_[29396]_  = \new_[29395]_  & \new_[29390]_ ;
  assign \new_[29400]_  = ~A167 & ~A169;
  assign \new_[29401]_  = A170 & \new_[29400]_ ;
  assign \new_[29405]_  = ~A200 & ~A199;
  assign \new_[29406]_  = A166 & \new_[29405]_ ;
  assign \new_[29407]_  = \new_[29406]_  & \new_[29401]_ ;
  assign \new_[29411]_  = ~A266 & ~A233;
  assign \new_[29412]_  = ~A232 & \new_[29411]_ ;
  assign \new_[29416]_  = A299 & ~A298;
  assign \new_[29417]_  = ~A267 & \new_[29416]_ ;
  assign \new_[29418]_  = \new_[29417]_  & \new_[29412]_ ;
  assign \new_[29422]_  = ~A167 & ~A169;
  assign \new_[29423]_  = A170 & \new_[29422]_ ;
  assign \new_[29427]_  = ~A200 & ~A199;
  assign \new_[29428]_  = A166 & \new_[29427]_ ;
  assign \new_[29429]_  = \new_[29428]_  & \new_[29423]_ ;
  assign \new_[29433]_  = ~A265 & ~A233;
  assign \new_[29434]_  = ~A232 & \new_[29433]_ ;
  assign \new_[29438]_  = A299 & ~A298;
  assign \new_[29439]_  = ~A266 & \new_[29438]_ ;
  assign \new_[29440]_  = \new_[29439]_  & \new_[29434]_ ;
  assign \new_[29444]_  = ~A168 & ~A169;
  assign \new_[29445]_  = ~A170 & \new_[29444]_ ;
  assign \new_[29449]_  = A201 & ~A200;
  assign \new_[29450]_  = A199 & \new_[29449]_ ;
  assign \new_[29451]_  = \new_[29450]_  & \new_[29445]_ ;
  assign \new_[29455]_  = A233 & ~A232;
  assign \new_[29456]_  = A202 & \new_[29455]_ ;
  assign \new_[29460]_  = ~A302 & ~A301;
  assign \new_[29461]_  = ~A299 & \new_[29460]_ ;
  assign \new_[29462]_  = \new_[29461]_  & \new_[29456]_ ;
  assign \new_[29466]_  = ~A168 & ~A169;
  assign \new_[29467]_  = ~A170 & \new_[29466]_ ;
  assign \new_[29471]_  = A201 & ~A200;
  assign \new_[29472]_  = A199 & \new_[29471]_ ;
  assign \new_[29473]_  = \new_[29472]_  & \new_[29467]_ ;
  assign \new_[29477]_  = A233 & ~A232;
  assign \new_[29478]_  = A203 & \new_[29477]_ ;
  assign \new_[29482]_  = ~A302 & ~A301;
  assign \new_[29483]_  = ~A299 & \new_[29482]_ ;
  assign \new_[29484]_  = \new_[29483]_  & \new_[29478]_ ;
  assign \new_[29488]_  = A199 & A166;
  assign \new_[29489]_  = A168 & \new_[29488]_ ;
  assign \new_[29493]_  = A233 & A232;
  assign \new_[29494]_  = A200 & \new_[29493]_ ;
  assign \new_[29495]_  = \new_[29494]_  & \new_[29489]_ ;
  assign \new_[29499]_  = ~A269 & ~A268;
  assign \new_[29500]_  = A265 & \new_[29499]_ ;
  assign \new_[29503]_  = ~A299 & A298;
  assign \new_[29506]_  = A301 & A300;
  assign \new_[29507]_  = \new_[29506]_  & \new_[29503]_ ;
  assign \new_[29508]_  = \new_[29507]_  & \new_[29500]_ ;
  assign \new_[29512]_  = A199 & A166;
  assign \new_[29513]_  = A168 & \new_[29512]_ ;
  assign \new_[29517]_  = A233 & A232;
  assign \new_[29518]_  = A200 & \new_[29517]_ ;
  assign \new_[29519]_  = \new_[29518]_  & \new_[29513]_ ;
  assign \new_[29523]_  = ~A269 & ~A268;
  assign \new_[29524]_  = A265 & \new_[29523]_ ;
  assign \new_[29527]_  = ~A299 & A298;
  assign \new_[29530]_  = A302 & A300;
  assign \new_[29531]_  = \new_[29530]_  & \new_[29527]_ ;
  assign \new_[29532]_  = \new_[29531]_  & \new_[29524]_ ;
  assign \new_[29536]_  = A199 & A166;
  assign \new_[29537]_  = A168 & \new_[29536]_ ;
  assign \new_[29541]_  = ~A235 & ~A233;
  assign \new_[29542]_  = A200 & \new_[29541]_ ;
  assign \new_[29543]_  = \new_[29542]_  & \new_[29537]_ ;
  assign \new_[29547]_  = A266 & A265;
  assign \new_[29548]_  = ~A236 & \new_[29547]_ ;
  assign \new_[29551]_  = ~A299 & A298;
  assign \new_[29554]_  = A301 & A300;
  assign \new_[29555]_  = \new_[29554]_  & \new_[29551]_ ;
  assign \new_[29556]_  = \new_[29555]_  & \new_[29548]_ ;
  assign \new_[29560]_  = A199 & A166;
  assign \new_[29561]_  = A168 & \new_[29560]_ ;
  assign \new_[29565]_  = ~A235 & ~A233;
  assign \new_[29566]_  = A200 & \new_[29565]_ ;
  assign \new_[29567]_  = \new_[29566]_  & \new_[29561]_ ;
  assign \new_[29571]_  = A266 & A265;
  assign \new_[29572]_  = ~A236 & \new_[29571]_ ;
  assign \new_[29575]_  = ~A299 & A298;
  assign \new_[29578]_  = A302 & A300;
  assign \new_[29579]_  = \new_[29578]_  & \new_[29575]_ ;
  assign \new_[29580]_  = \new_[29579]_  & \new_[29572]_ ;
  assign \new_[29584]_  = A199 & A166;
  assign \new_[29585]_  = A168 & \new_[29584]_ ;
  assign \new_[29589]_  = ~A235 & ~A233;
  assign \new_[29590]_  = A200 & \new_[29589]_ ;
  assign \new_[29591]_  = \new_[29590]_  & \new_[29585]_ ;
  assign \new_[29595]_  = ~A267 & ~A266;
  assign \new_[29596]_  = ~A236 & \new_[29595]_ ;
  assign \new_[29599]_  = ~A299 & A298;
  assign \new_[29602]_  = A301 & A300;
  assign \new_[29603]_  = \new_[29602]_  & \new_[29599]_ ;
  assign \new_[29604]_  = \new_[29603]_  & \new_[29596]_ ;
  assign \new_[29608]_  = A199 & A166;
  assign \new_[29609]_  = A168 & \new_[29608]_ ;
  assign \new_[29613]_  = ~A235 & ~A233;
  assign \new_[29614]_  = A200 & \new_[29613]_ ;
  assign \new_[29615]_  = \new_[29614]_  & \new_[29609]_ ;
  assign \new_[29619]_  = ~A267 & ~A266;
  assign \new_[29620]_  = ~A236 & \new_[29619]_ ;
  assign \new_[29623]_  = ~A299 & A298;
  assign \new_[29626]_  = A302 & A300;
  assign \new_[29627]_  = \new_[29626]_  & \new_[29623]_ ;
  assign \new_[29628]_  = \new_[29627]_  & \new_[29620]_ ;
  assign \new_[29632]_  = A199 & A166;
  assign \new_[29633]_  = A168 & \new_[29632]_ ;
  assign \new_[29637]_  = ~A235 & ~A233;
  assign \new_[29638]_  = A200 & \new_[29637]_ ;
  assign \new_[29639]_  = \new_[29638]_  & \new_[29633]_ ;
  assign \new_[29643]_  = ~A266 & ~A265;
  assign \new_[29644]_  = ~A236 & \new_[29643]_ ;
  assign \new_[29647]_  = ~A299 & A298;
  assign \new_[29650]_  = A301 & A300;
  assign \new_[29651]_  = \new_[29650]_  & \new_[29647]_ ;
  assign \new_[29652]_  = \new_[29651]_  & \new_[29644]_ ;
  assign \new_[29656]_  = A199 & A166;
  assign \new_[29657]_  = A168 & \new_[29656]_ ;
  assign \new_[29661]_  = ~A235 & ~A233;
  assign \new_[29662]_  = A200 & \new_[29661]_ ;
  assign \new_[29663]_  = \new_[29662]_  & \new_[29657]_ ;
  assign \new_[29667]_  = ~A266 & ~A265;
  assign \new_[29668]_  = ~A236 & \new_[29667]_ ;
  assign \new_[29671]_  = ~A299 & A298;
  assign \new_[29674]_  = A302 & A300;
  assign \new_[29675]_  = \new_[29674]_  & \new_[29671]_ ;
  assign \new_[29676]_  = \new_[29675]_  & \new_[29668]_ ;
  assign \new_[29680]_  = A199 & A166;
  assign \new_[29681]_  = A168 & \new_[29680]_ ;
  assign \new_[29685]_  = ~A234 & ~A233;
  assign \new_[29686]_  = A200 & \new_[29685]_ ;
  assign \new_[29687]_  = \new_[29686]_  & \new_[29681]_ ;
  assign \new_[29691]_  = ~A269 & ~A268;
  assign \new_[29692]_  = ~A266 & \new_[29691]_ ;
  assign \new_[29695]_  = ~A299 & A298;
  assign \new_[29698]_  = A301 & A300;
  assign \new_[29699]_  = \new_[29698]_  & \new_[29695]_ ;
  assign \new_[29700]_  = \new_[29699]_  & \new_[29692]_ ;
  assign \new_[29704]_  = A199 & A166;
  assign \new_[29705]_  = A168 & \new_[29704]_ ;
  assign \new_[29709]_  = ~A234 & ~A233;
  assign \new_[29710]_  = A200 & \new_[29709]_ ;
  assign \new_[29711]_  = \new_[29710]_  & \new_[29705]_ ;
  assign \new_[29715]_  = ~A269 & ~A268;
  assign \new_[29716]_  = ~A266 & \new_[29715]_ ;
  assign \new_[29719]_  = ~A299 & A298;
  assign \new_[29722]_  = A302 & A300;
  assign \new_[29723]_  = \new_[29722]_  & \new_[29719]_ ;
  assign \new_[29724]_  = \new_[29723]_  & \new_[29716]_ ;
  assign \new_[29728]_  = A199 & A166;
  assign \new_[29729]_  = A168 & \new_[29728]_ ;
  assign \new_[29733]_  = ~A233 & ~A232;
  assign \new_[29734]_  = A200 & \new_[29733]_ ;
  assign \new_[29735]_  = \new_[29734]_  & \new_[29729]_ ;
  assign \new_[29739]_  = ~A269 & ~A268;
  assign \new_[29740]_  = ~A266 & \new_[29739]_ ;
  assign \new_[29743]_  = ~A299 & A298;
  assign \new_[29746]_  = A301 & A300;
  assign \new_[29747]_  = \new_[29746]_  & \new_[29743]_ ;
  assign \new_[29748]_  = \new_[29747]_  & \new_[29740]_ ;
  assign \new_[29752]_  = A199 & A166;
  assign \new_[29753]_  = A168 & \new_[29752]_ ;
  assign \new_[29757]_  = ~A233 & ~A232;
  assign \new_[29758]_  = A200 & \new_[29757]_ ;
  assign \new_[29759]_  = \new_[29758]_  & \new_[29753]_ ;
  assign \new_[29763]_  = ~A269 & ~A268;
  assign \new_[29764]_  = ~A266 & \new_[29763]_ ;
  assign \new_[29767]_  = ~A299 & A298;
  assign \new_[29770]_  = A302 & A300;
  assign \new_[29771]_  = \new_[29770]_  & \new_[29767]_ ;
  assign \new_[29772]_  = \new_[29771]_  & \new_[29764]_ ;
  assign \new_[29776]_  = ~A200 & A166;
  assign \new_[29777]_  = A168 & \new_[29776]_ ;
  assign \new_[29781]_  = A232 & ~A203;
  assign \new_[29782]_  = ~A202 & \new_[29781]_ ;
  assign \new_[29783]_  = \new_[29782]_  & \new_[29777]_ ;
  assign \new_[29787]_  = ~A267 & A265;
  assign \new_[29788]_  = A233 & \new_[29787]_ ;
  assign \new_[29791]_  = ~A299 & A298;
  assign \new_[29794]_  = A301 & A300;
  assign \new_[29795]_  = \new_[29794]_  & \new_[29791]_ ;
  assign \new_[29796]_  = \new_[29795]_  & \new_[29788]_ ;
  assign \new_[29800]_  = ~A200 & A166;
  assign \new_[29801]_  = A168 & \new_[29800]_ ;
  assign \new_[29805]_  = A232 & ~A203;
  assign \new_[29806]_  = ~A202 & \new_[29805]_ ;
  assign \new_[29807]_  = \new_[29806]_  & \new_[29801]_ ;
  assign \new_[29811]_  = ~A267 & A265;
  assign \new_[29812]_  = A233 & \new_[29811]_ ;
  assign \new_[29815]_  = ~A299 & A298;
  assign \new_[29818]_  = A302 & A300;
  assign \new_[29819]_  = \new_[29818]_  & \new_[29815]_ ;
  assign \new_[29820]_  = \new_[29819]_  & \new_[29812]_ ;
  assign \new_[29824]_  = ~A200 & A166;
  assign \new_[29825]_  = A168 & \new_[29824]_ ;
  assign \new_[29829]_  = A232 & ~A203;
  assign \new_[29830]_  = ~A202 & \new_[29829]_ ;
  assign \new_[29831]_  = \new_[29830]_  & \new_[29825]_ ;
  assign \new_[29835]_  = A266 & A265;
  assign \new_[29836]_  = A233 & \new_[29835]_ ;
  assign \new_[29839]_  = ~A299 & A298;
  assign \new_[29842]_  = A301 & A300;
  assign \new_[29843]_  = \new_[29842]_  & \new_[29839]_ ;
  assign \new_[29844]_  = \new_[29843]_  & \new_[29836]_ ;
  assign \new_[29848]_  = ~A200 & A166;
  assign \new_[29849]_  = A168 & \new_[29848]_ ;
  assign \new_[29853]_  = A232 & ~A203;
  assign \new_[29854]_  = ~A202 & \new_[29853]_ ;
  assign \new_[29855]_  = \new_[29854]_  & \new_[29849]_ ;
  assign \new_[29859]_  = A266 & A265;
  assign \new_[29860]_  = A233 & \new_[29859]_ ;
  assign \new_[29863]_  = ~A299 & A298;
  assign \new_[29866]_  = A302 & A300;
  assign \new_[29867]_  = \new_[29866]_  & \new_[29863]_ ;
  assign \new_[29868]_  = \new_[29867]_  & \new_[29860]_ ;
  assign \new_[29872]_  = ~A200 & A166;
  assign \new_[29873]_  = A168 & \new_[29872]_ ;
  assign \new_[29877]_  = A232 & ~A203;
  assign \new_[29878]_  = ~A202 & \new_[29877]_ ;
  assign \new_[29879]_  = \new_[29878]_  & \new_[29873]_ ;
  assign \new_[29883]_  = ~A266 & ~A265;
  assign \new_[29884]_  = A233 & \new_[29883]_ ;
  assign \new_[29887]_  = ~A299 & A298;
  assign \new_[29890]_  = A301 & A300;
  assign \new_[29891]_  = \new_[29890]_  & \new_[29887]_ ;
  assign \new_[29892]_  = \new_[29891]_  & \new_[29884]_ ;
  assign \new_[29896]_  = ~A200 & A166;
  assign \new_[29897]_  = A168 & \new_[29896]_ ;
  assign \new_[29901]_  = A232 & ~A203;
  assign \new_[29902]_  = ~A202 & \new_[29901]_ ;
  assign \new_[29903]_  = \new_[29902]_  & \new_[29897]_ ;
  assign \new_[29907]_  = ~A266 & ~A265;
  assign \new_[29908]_  = A233 & \new_[29907]_ ;
  assign \new_[29911]_  = ~A299 & A298;
  assign \new_[29914]_  = A302 & A300;
  assign \new_[29915]_  = \new_[29914]_  & \new_[29911]_ ;
  assign \new_[29916]_  = \new_[29915]_  & \new_[29908]_ ;
  assign \new_[29920]_  = ~A200 & A166;
  assign \new_[29921]_  = A168 & \new_[29920]_ ;
  assign \new_[29925]_  = ~A233 & ~A203;
  assign \new_[29926]_  = ~A202 & \new_[29925]_ ;
  assign \new_[29927]_  = \new_[29926]_  & \new_[29921]_ ;
  assign \new_[29931]_  = ~A266 & ~A236;
  assign \new_[29932]_  = ~A235 & \new_[29931]_ ;
  assign \new_[29935]_  = ~A269 & ~A268;
  assign \new_[29938]_  = A299 & ~A298;
  assign \new_[29939]_  = \new_[29938]_  & \new_[29935]_ ;
  assign \new_[29940]_  = \new_[29939]_  & \new_[29932]_ ;
  assign \new_[29944]_  = ~A200 & A166;
  assign \new_[29945]_  = A168 & \new_[29944]_ ;
  assign \new_[29949]_  = ~A233 & ~A203;
  assign \new_[29950]_  = ~A202 & \new_[29949]_ ;
  assign \new_[29951]_  = \new_[29950]_  & \new_[29945]_ ;
  assign \new_[29955]_  = A266 & A265;
  assign \new_[29956]_  = ~A234 & \new_[29955]_ ;
  assign \new_[29959]_  = ~A299 & A298;
  assign \new_[29962]_  = A301 & A300;
  assign \new_[29963]_  = \new_[29962]_  & \new_[29959]_ ;
  assign \new_[29964]_  = \new_[29963]_  & \new_[29956]_ ;
  assign \new_[29968]_  = ~A200 & A166;
  assign \new_[29969]_  = A168 & \new_[29968]_ ;
  assign \new_[29973]_  = ~A233 & ~A203;
  assign \new_[29974]_  = ~A202 & \new_[29973]_ ;
  assign \new_[29975]_  = \new_[29974]_  & \new_[29969]_ ;
  assign \new_[29979]_  = A266 & A265;
  assign \new_[29980]_  = ~A234 & \new_[29979]_ ;
  assign \new_[29983]_  = ~A299 & A298;
  assign \new_[29986]_  = A302 & A300;
  assign \new_[29987]_  = \new_[29986]_  & \new_[29983]_ ;
  assign \new_[29988]_  = \new_[29987]_  & \new_[29980]_ ;
  assign \new_[29992]_  = ~A200 & A166;
  assign \new_[29993]_  = A168 & \new_[29992]_ ;
  assign \new_[29997]_  = ~A233 & ~A203;
  assign \new_[29998]_  = ~A202 & \new_[29997]_ ;
  assign \new_[29999]_  = \new_[29998]_  & \new_[29993]_ ;
  assign \new_[30003]_  = ~A267 & ~A266;
  assign \new_[30004]_  = ~A234 & \new_[30003]_ ;
  assign \new_[30007]_  = ~A299 & A298;
  assign \new_[30010]_  = A301 & A300;
  assign \new_[30011]_  = \new_[30010]_  & \new_[30007]_ ;
  assign \new_[30012]_  = \new_[30011]_  & \new_[30004]_ ;
  assign \new_[30016]_  = ~A200 & A166;
  assign \new_[30017]_  = A168 & \new_[30016]_ ;
  assign \new_[30021]_  = ~A233 & ~A203;
  assign \new_[30022]_  = ~A202 & \new_[30021]_ ;
  assign \new_[30023]_  = \new_[30022]_  & \new_[30017]_ ;
  assign \new_[30027]_  = ~A267 & ~A266;
  assign \new_[30028]_  = ~A234 & \new_[30027]_ ;
  assign \new_[30031]_  = ~A299 & A298;
  assign \new_[30034]_  = A302 & A300;
  assign \new_[30035]_  = \new_[30034]_  & \new_[30031]_ ;
  assign \new_[30036]_  = \new_[30035]_  & \new_[30028]_ ;
  assign \new_[30040]_  = ~A200 & A166;
  assign \new_[30041]_  = A168 & \new_[30040]_ ;
  assign \new_[30045]_  = ~A233 & ~A203;
  assign \new_[30046]_  = ~A202 & \new_[30045]_ ;
  assign \new_[30047]_  = \new_[30046]_  & \new_[30041]_ ;
  assign \new_[30051]_  = ~A266 & ~A265;
  assign \new_[30052]_  = ~A234 & \new_[30051]_ ;
  assign \new_[30055]_  = ~A299 & A298;
  assign \new_[30058]_  = A301 & A300;
  assign \new_[30059]_  = \new_[30058]_  & \new_[30055]_ ;
  assign \new_[30060]_  = \new_[30059]_  & \new_[30052]_ ;
  assign \new_[30064]_  = ~A200 & A166;
  assign \new_[30065]_  = A168 & \new_[30064]_ ;
  assign \new_[30069]_  = ~A233 & ~A203;
  assign \new_[30070]_  = ~A202 & \new_[30069]_ ;
  assign \new_[30071]_  = \new_[30070]_  & \new_[30065]_ ;
  assign \new_[30075]_  = ~A266 & ~A265;
  assign \new_[30076]_  = ~A234 & \new_[30075]_ ;
  assign \new_[30079]_  = ~A299 & A298;
  assign \new_[30082]_  = A302 & A300;
  assign \new_[30083]_  = \new_[30082]_  & \new_[30079]_ ;
  assign \new_[30084]_  = \new_[30083]_  & \new_[30076]_ ;
  assign \new_[30088]_  = ~A200 & A166;
  assign \new_[30089]_  = A168 & \new_[30088]_ ;
  assign \new_[30093]_  = A232 & ~A203;
  assign \new_[30094]_  = ~A202 & \new_[30093]_ ;
  assign \new_[30095]_  = \new_[30094]_  & \new_[30089]_ ;
  assign \new_[30099]_  = A235 & A234;
  assign \new_[30100]_  = ~A233 & \new_[30099]_ ;
  assign \new_[30103]_  = ~A266 & A265;
  assign \new_[30106]_  = A268 & A267;
  assign \new_[30107]_  = \new_[30106]_  & \new_[30103]_ ;
  assign \new_[30108]_  = \new_[30107]_  & \new_[30100]_ ;
  assign \new_[30112]_  = ~A200 & A166;
  assign \new_[30113]_  = A168 & \new_[30112]_ ;
  assign \new_[30117]_  = A232 & ~A203;
  assign \new_[30118]_  = ~A202 & \new_[30117]_ ;
  assign \new_[30119]_  = \new_[30118]_  & \new_[30113]_ ;
  assign \new_[30123]_  = A235 & A234;
  assign \new_[30124]_  = ~A233 & \new_[30123]_ ;
  assign \new_[30127]_  = ~A266 & A265;
  assign \new_[30130]_  = A269 & A267;
  assign \new_[30131]_  = \new_[30130]_  & \new_[30127]_ ;
  assign \new_[30132]_  = \new_[30131]_  & \new_[30124]_ ;
  assign \new_[30136]_  = ~A200 & A166;
  assign \new_[30137]_  = A168 & \new_[30136]_ ;
  assign \new_[30141]_  = A232 & ~A203;
  assign \new_[30142]_  = ~A202 & \new_[30141]_ ;
  assign \new_[30143]_  = \new_[30142]_  & \new_[30137]_ ;
  assign \new_[30147]_  = A236 & A234;
  assign \new_[30148]_  = ~A233 & \new_[30147]_ ;
  assign \new_[30151]_  = ~A266 & A265;
  assign \new_[30154]_  = A268 & A267;
  assign \new_[30155]_  = \new_[30154]_  & \new_[30151]_ ;
  assign \new_[30156]_  = \new_[30155]_  & \new_[30148]_ ;
  assign \new_[30160]_  = ~A200 & A166;
  assign \new_[30161]_  = A168 & \new_[30160]_ ;
  assign \new_[30165]_  = A232 & ~A203;
  assign \new_[30166]_  = ~A202 & \new_[30165]_ ;
  assign \new_[30167]_  = \new_[30166]_  & \new_[30161]_ ;
  assign \new_[30171]_  = A236 & A234;
  assign \new_[30172]_  = ~A233 & \new_[30171]_ ;
  assign \new_[30175]_  = ~A266 & A265;
  assign \new_[30178]_  = A269 & A267;
  assign \new_[30179]_  = \new_[30178]_  & \new_[30175]_ ;
  assign \new_[30180]_  = \new_[30179]_  & \new_[30172]_ ;
  assign \new_[30184]_  = ~A200 & A166;
  assign \new_[30185]_  = A168 & \new_[30184]_ ;
  assign \new_[30189]_  = ~A232 & ~A203;
  assign \new_[30190]_  = ~A202 & \new_[30189]_ ;
  assign \new_[30191]_  = \new_[30190]_  & \new_[30185]_ ;
  assign \new_[30195]_  = A266 & A265;
  assign \new_[30196]_  = ~A233 & \new_[30195]_ ;
  assign \new_[30199]_  = ~A299 & A298;
  assign \new_[30202]_  = A301 & A300;
  assign \new_[30203]_  = \new_[30202]_  & \new_[30199]_ ;
  assign \new_[30204]_  = \new_[30203]_  & \new_[30196]_ ;
  assign \new_[30208]_  = ~A200 & A166;
  assign \new_[30209]_  = A168 & \new_[30208]_ ;
  assign \new_[30213]_  = ~A232 & ~A203;
  assign \new_[30214]_  = ~A202 & \new_[30213]_ ;
  assign \new_[30215]_  = \new_[30214]_  & \new_[30209]_ ;
  assign \new_[30219]_  = A266 & A265;
  assign \new_[30220]_  = ~A233 & \new_[30219]_ ;
  assign \new_[30223]_  = ~A299 & A298;
  assign \new_[30226]_  = A302 & A300;
  assign \new_[30227]_  = \new_[30226]_  & \new_[30223]_ ;
  assign \new_[30228]_  = \new_[30227]_  & \new_[30220]_ ;
  assign \new_[30232]_  = ~A200 & A166;
  assign \new_[30233]_  = A168 & \new_[30232]_ ;
  assign \new_[30237]_  = ~A232 & ~A203;
  assign \new_[30238]_  = ~A202 & \new_[30237]_ ;
  assign \new_[30239]_  = \new_[30238]_  & \new_[30233]_ ;
  assign \new_[30243]_  = ~A267 & ~A266;
  assign \new_[30244]_  = ~A233 & \new_[30243]_ ;
  assign \new_[30247]_  = ~A299 & A298;
  assign \new_[30250]_  = A301 & A300;
  assign \new_[30251]_  = \new_[30250]_  & \new_[30247]_ ;
  assign \new_[30252]_  = \new_[30251]_  & \new_[30244]_ ;
  assign \new_[30256]_  = ~A200 & A166;
  assign \new_[30257]_  = A168 & \new_[30256]_ ;
  assign \new_[30261]_  = ~A232 & ~A203;
  assign \new_[30262]_  = ~A202 & \new_[30261]_ ;
  assign \new_[30263]_  = \new_[30262]_  & \new_[30257]_ ;
  assign \new_[30267]_  = ~A267 & ~A266;
  assign \new_[30268]_  = ~A233 & \new_[30267]_ ;
  assign \new_[30271]_  = ~A299 & A298;
  assign \new_[30274]_  = A302 & A300;
  assign \new_[30275]_  = \new_[30274]_  & \new_[30271]_ ;
  assign \new_[30276]_  = \new_[30275]_  & \new_[30268]_ ;
  assign \new_[30280]_  = ~A200 & A166;
  assign \new_[30281]_  = A168 & \new_[30280]_ ;
  assign \new_[30285]_  = ~A232 & ~A203;
  assign \new_[30286]_  = ~A202 & \new_[30285]_ ;
  assign \new_[30287]_  = \new_[30286]_  & \new_[30281]_ ;
  assign \new_[30291]_  = ~A266 & ~A265;
  assign \new_[30292]_  = ~A233 & \new_[30291]_ ;
  assign \new_[30295]_  = ~A299 & A298;
  assign \new_[30298]_  = A301 & A300;
  assign \new_[30299]_  = \new_[30298]_  & \new_[30295]_ ;
  assign \new_[30300]_  = \new_[30299]_  & \new_[30292]_ ;
  assign \new_[30304]_  = ~A200 & A166;
  assign \new_[30305]_  = A168 & \new_[30304]_ ;
  assign \new_[30309]_  = ~A232 & ~A203;
  assign \new_[30310]_  = ~A202 & \new_[30309]_ ;
  assign \new_[30311]_  = \new_[30310]_  & \new_[30305]_ ;
  assign \new_[30315]_  = ~A266 & ~A265;
  assign \new_[30316]_  = ~A233 & \new_[30315]_ ;
  assign \new_[30319]_  = ~A299 & A298;
  assign \new_[30322]_  = A302 & A300;
  assign \new_[30323]_  = \new_[30322]_  & \new_[30319]_ ;
  assign \new_[30324]_  = \new_[30323]_  & \new_[30316]_ ;
  assign \new_[30328]_  = ~A200 & A166;
  assign \new_[30329]_  = A168 & \new_[30328]_ ;
  assign \new_[30333]_  = A233 & A232;
  assign \new_[30334]_  = ~A201 & \new_[30333]_ ;
  assign \new_[30335]_  = \new_[30334]_  & \new_[30329]_ ;
  assign \new_[30339]_  = ~A269 & ~A268;
  assign \new_[30340]_  = A265 & \new_[30339]_ ;
  assign \new_[30343]_  = ~A299 & A298;
  assign \new_[30346]_  = A301 & A300;
  assign \new_[30347]_  = \new_[30346]_  & \new_[30343]_ ;
  assign \new_[30348]_  = \new_[30347]_  & \new_[30340]_ ;
  assign \new_[30352]_  = ~A200 & A166;
  assign \new_[30353]_  = A168 & \new_[30352]_ ;
  assign \new_[30357]_  = A233 & A232;
  assign \new_[30358]_  = ~A201 & \new_[30357]_ ;
  assign \new_[30359]_  = \new_[30358]_  & \new_[30353]_ ;
  assign \new_[30363]_  = ~A269 & ~A268;
  assign \new_[30364]_  = A265 & \new_[30363]_ ;
  assign \new_[30367]_  = ~A299 & A298;
  assign \new_[30370]_  = A302 & A300;
  assign \new_[30371]_  = \new_[30370]_  & \new_[30367]_ ;
  assign \new_[30372]_  = \new_[30371]_  & \new_[30364]_ ;
  assign \new_[30376]_  = ~A200 & A166;
  assign \new_[30377]_  = A168 & \new_[30376]_ ;
  assign \new_[30381]_  = ~A235 & ~A233;
  assign \new_[30382]_  = ~A201 & \new_[30381]_ ;
  assign \new_[30383]_  = \new_[30382]_  & \new_[30377]_ ;
  assign \new_[30387]_  = A266 & A265;
  assign \new_[30388]_  = ~A236 & \new_[30387]_ ;
  assign \new_[30391]_  = ~A299 & A298;
  assign \new_[30394]_  = A301 & A300;
  assign \new_[30395]_  = \new_[30394]_  & \new_[30391]_ ;
  assign \new_[30396]_  = \new_[30395]_  & \new_[30388]_ ;
  assign \new_[30400]_  = ~A200 & A166;
  assign \new_[30401]_  = A168 & \new_[30400]_ ;
  assign \new_[30405]_  = ~A235 & ~A233;
  assign \new_[30406]_  = ~A201 & \new_[30405]_ ;
  assign \new_[30407]_  = \new_[30406]_  & \new_[30401]_ ;
  assign \new_[30411]_  = A266 & A265;
  assign \new_[30412]_  = ~A236 & \new_[30411]_ ;
  assign \new_[30415]_  = ~A299 & A298;
  assign \new_[30418]_  = A302 & A300;
  assign \new_[30419]_  = \new_[30418]_  & \new_[30415]_ ;
  assign \new_[30420]_  = \new_[30419]_  & \new_[30412]_ ;
  assign \new_[30424]_  = ~A200 & A166;
  assign \new_[30425]_  = A168 & \new_[30424]_ ;
  assign \new_[30429]_  = ~A235 & ~A233;
  assign \new_[30430]_  = ~A201 & \new_[30429]_ ;
  assign \new_[30431]_  = \new_[30430]_  & \new_[30425]_ ;
  assign \new_[30435]_  = ~A267 & ~A266;
  assign \new_[30436]_  = ~A236 & \new_[30435]_ ;
  assign \new_[30439]_  = ~A299 & A298;
  assign \new_[30442]_  = A301 & A300;
  assign \new_[30443]_  = \new_[30442]_  & \new_[30439]_ ;
  assign \new_[30444]_  = \new_[30443]_  & \new_[30436]_ ;
  assign \new_[30448]_  = ~A200 & A166;
  assign \new_[30449]_  = A168 & \new_[30448]_ ;
  assign \new_[30453]_  = ~A235 & ~A233;
  assign \new_[30454]_  = ~A201 & \new_[30453]_ ;
  assign \new_[30455]_  = \new_[30454]_  & \new_[30449]_ ;
  assign \new_[30459]_  = ~A267 & ~A266;
  assign \new_[30460]_  = ~A236 & \new_[30459]_ ;
  assign \new_[30463]_  = ~A299 & A298;
  assign \new_[30466]_  = A302 & A300;
  assign \new_[30467]_  = \new_[30466]_  & \new_[30463]_ ;
  assign \new_[30468]_  = \new_[30467]_  & \new_[30460]_ ;
  assign \new_[30472]_  = ~A200 & A166;
  assign \new_[30473]_  = A168 & \new_[30472]_ ;
  assign \new_[30477]_  = ~A235 & ~A233;
  assign \new_[30478]_  = ~A201 & \new_[30477]_ ;
  assign \new_[30479]_  = \new_[30478]_  & \new_[30473]_ ;
  assign \new_[30483]_  = ~A266 & ~A265;
  assign \new_[30484]_  = ~A236 & \new_[30483]_ ;
  assign \new_[30487]_  = ~A299 & A298;
  assign \new_[30490]_  = A301 & A300;
  assign \new_[30491]_  = \new_[30490]_  & \new_[30487]_ ;
  assign \new_[30492]_  = \new_[30491]_  & \new_[30484]_ ;
  assign \new_[30496]_  = ~A200 & A166;
  assign \new_[30497]_  = A168 & \new_[30496]_ ;
  assign \new_[30501]_  = ~A235 & ~A233;
  assign \new_[30502]_  = ~A201 & \new_[30501]_ ;
  assign \new_[30503]_  = \new_[30502]_  & \new_[30497]_ ;
  assign \new_[30507]_  = ~A266 & ~A265;
  assign \new_[30508]_  = ~A236 & \new_[30507]_ ;
  assign \new_[30511]_  = ~A299 & A298;
  assign \new_[30514]_  = A302 & A300;
  assign \new_[30515]_  = \new_[30514]_  & \new_[30511]_ ;
  assign \new_[30516]_  = \new_[30515]_  & \new_[30508]_ ;
  assign \new_[30520]_  = ~A200 & A166;
  assign \new_[30521]_  = A168 & \new_[30520]_ ;
  assign \new_[30525]_  = ~A234 & ~A233;
  assign \new_[30526]_  = ~A201 & \new_[30525]_ ;
  assign \new_[30527]_  = \new_[30526]_  & \new_[30521]_ ;
  assign \new_[30531]_  = ~A269 & ~A268;
  assign \new_[30532]_  = ~A266 & \new_[30531]_ ;
  assign \new_[30535]_  = ~A299 & A298;
  assign \new_[30538]_  = A301 & A300;
  assign \new_[30539]_  = \new_[30538]_  & \new_[30535]_ ;
  assign \new_[30540]_  = \new_[30539]_  & \new_[30532]_ ;
  assign \new_[30544]_  = ~A200 & A166;
  assign \new_[30545]_  = A168 & \new_[30544]_ ;
  assign \new_[30549]_  = ~A234 & ~A233;
  assign \new_[30550]_  = ~A201 & \new_[30549]_ ;
  assign \new_[30551]_  = \new_[30550]_  & \new_[30545]_ ;
  assign \new_[30555]_  = ~A269 & ~A268;
  assign \new_[30556]_  = ~A266 & \new_[30555]_ ;
  assign \new_[30559]_  = ~A299 & A298;
  assign \new_[30562]_  = A302 & A300;
  assign \new_[30563]_  = \new_[30562]_  & \new_[30559]_ ;
  assign \new_[30564]_  = \new_[30563]_  & \new_[30556]_ ;
  assign \new_[30568]_  = ~A200 & A166;
  assign \new_[30569]_  = A168 & \new_[30568]_ ;
  assign \new_[30573]_  = ~A233 & ~A232;
  assign \new_[30574]_  = ~A201 & \new_[30573]_ ;
  assign \new_[30575]_  = \new_[30574]_  & \new_[30569]_ ;
  assign \new_[30579]_  = ~A269 & ~A268;
  assign \new_[30580]_  = ~A266 & \new_[30579]_ ;
  assign \new_[30583]_  = ~A299 & A298;
  assign \new_[30586]_  = A301 & A300;
  assign \new_[30587]_  = \new_[30586]_  & \new_[30583]_ ;
  assign \new_[30588]_  = \new_[30587]_  & \new_[30580]_ ;
  assign \new_[30592]_  = ~A200 & A166;
  assign \new_[30593]_  = A168 & \new_[30592]_ ;
  assign \new_[30597]_  = ~A233 & ~A232;
  assign \new_[30598]_  = ~A201 & \new_[30597]_ ;
  assign \new_[30599]_  = \new_[30598]_  & \new_[30593]_ ;
  assign \new_[30603]_  = ~A269 & ~A268;
  assign \new_[30604]_  = ~A266 & \new_[30603]_ ;
  assign \new_[30607]_  = ~A299 & A298;
  assign \new_[30610]_  = A302 & A300;
  assign \new_[30611]_  = \new_[30610]_  & \new_[30607]_ ;
  assign \new_[30612]_  = \new_[30611]_  & \new_[30604]_ ;
  assign \new_[30616]_  = ~A199 & A166;
  assign \new_[30617]_  = A168 & \new_[30616]_ ;
  assign \new_[30621]_  = A233 & A232;
  assign \new_[30622]_  = ~A200 & \new_[30621]_ ;
  assign \new_[30623]_  = \new_[30622]_  & \new_[30617]_ ;
  assign \new_[30627]_  = ~A269 & ~A268;
  assign \new_[30628]_  = A265 & \new_[30627]_ ;
  assign \new_[30631]_  = ~A299 & A298;
  assign \new_[30634]_  = A301 & A300;
  assign \new_[30635]_  = \new_[30634]_  & \new_[30631]_ ;
  assign \new_[30636]_  = \new_[30635]_  & \new_[30628]_ ;
  assign \new_[30640]_  = ~A199 & A166;
  assign \new_[30641]_  = A168 & \new_[30640]_ ;
  assign \new_[30645]_  = A233 & A232;
  assign \new_[30646]_  = ~A200 & \new_[30645]_ ;
  assign \new_[30647]_  = \new_[30646]_  & \new_[30641]_ ;
  assign \new_[30651]_  = ~A269 & ~A268;
  assign \new_[30652]_  = A265 & \new_[30651]_ ;
  assign \new_[30655]_  = ~A299 & A298;
  assign \new_[30658]_  = A302 & A300;
  assign \new_[30659]_  = \new_[30658]_  & \new_[30655]_ ;
  assign \new_[30660]_  = \new_[30659]_  & \new_[30652]_ ;
  assign \new_[30664]_  = ~A199 & A166;
  assign \new_[30665]_  = A168 & \new_[30664]_ ;
  assign \new_[30669]_  = ~A235 & ~A233;
  assign \new_[30670]_  = ~A200 & \new_[30669]_ ;
  assign \new_[30671]_  = \new_[30670]_  & \new_[30665]_ ;
  assign \new_[30675]_  = A266 & A265;
  assign \new_[30676]_  = ~A236 & \new_[30675]_ ;
  assign \new_[30679]_  = ~A299 & A298;
  assign \new_[30682]_  = A301 & A300;
  assign \new_[30683]_  = \new_[30682]_  & \new_[30679]_ ;
  assign \new_[30684]_  = \new_[30683]_  & \new_[30676]_ ;
  assign \new_[30688]_  = ~A199 & A166;
  assign \new_[30689]_  = A168 & \new_[30688]_ ;
  assign \new_[30693]_  = ~A235 & ~A233;
  assign \new_[30694]_  = ~A200 & \new_[30693]_ ;
  assign \new_[30695]_  = \new_[30694]_  & \new_[30689]_ ;
  assign \new_[30699]_  = A266 & A265;
  assign \new_[30700]_  = ~A236 & \new_[30699]_ ;
  assign \new_[30703]_  = ~A299 & A298;
  assign \new_[30706]_  = A302 & A300;
  assign \new_[30707]_  = \new_[30706]_  & \new_[30703]_ ;
  assign \new_[30708]_  = \new_[30707]_  & \new_[30700]_ ;
  assign \new_[30712]_  = ~A199 & A166;
  assign \new_[30713]_  = A168 & \new_[30712]_ ;
  assign \new_[30717]_  = ~A235 & ~A233;
  assign \new_[30718]_  = ~A200 & \new_[30717]_ ;
  assign \new_[30719]_  = \new_[30718]_  & \new_[30713]_ ;
  assign \new_[30723]_  = ~A267 & ~A266;
  assign \new_[30724]_  = ~A236 & \new_[30723]_ ;
  assign \new_[30727]_  = ~A299 & A298;
  assign \new_[30730]_  = A301 & A300;
  assign \new_[30731]_  = \new_[30730]_  & \new_[30727]_ ;
  assign \new_[30732]_  = \new_[30731]_  & \new_[30724]_ ;
  assign \new_[30736]_  = ~A199 & A166;
  assign \new_[30737]_  = A168 & \new_[30736]_ ;
  assign \new_[30741]_  = ~A235 & ~A233;
  assign \new_[30742]_  = ~A200 & \new_[30741]_ ;
  assign \new_[30743]_  = \new_[30742]_  & \new_[30737]_ ;
  assign \new_[30747]_  = ~A267 & ~A266;
  assign \new_[30748]_  = ~A236 & \new_[30747]_ ;
  assign \new_[30751]_  = ~A299 & A298;
  assign \new_[30754]_  = A302 & A300;
  assign \new_[30755]_  = \new_[30754]_  & \new_[30751]_ ;
  assign \new_[30756]_  = \new_[30755]_  & \new_[30748]_ ;
  assign \new_[30760]_  = ~A199 & A166;
  assign \new_[30761]_  = A168 & \new_[30760]_ ;
  assign \new_[30765]_  = ~A235 & ~A233;
  assign \new_[30766]_  = ~A200 & \new_[30765]_ ;
  assign \new_[30767]_  = \new_[30766]_  & \new_[30761]_ ;
  assign \new_[30771]_  = ~A266 & ~A265;
  assign \new_[30772]_  = ~A236 & \new_[30771]_ ;
  assign \new_[30775]_  = ~A299 & A298;
  assign \new_[30778]_  = A301 & A300;
  assign \new_[30779]_  = \new_[30778]_  & \new_[30775]_ ;
  assign \new_[30780]_  = \new_[30779]_  & \new_[30772]_ ;
  assign \new_[30784]_  = ~A199 & A166;
  assign \new_[30785]_  = A168 & \new_[30784]_ ;
  assign \new_[30789]_  = ~A235 & ~A233;
  assign \new_[30790]_  = ~A200 & \new_[30789]_ ;
  assign \new_[30791]_  = \new_[30790]_  & \new_[30785]_ ;
  assign \new_[30795]_  = ~A266 & ~A265;
  assign \new_[30796]_  = ~A236 & \new_[30795]_ ;
  assign \new_[30799]_  = ~A299 & A298;
  assign \new_[30802]_  = A302 & A300;
  assign \new_[30803]_  = \new_[30802]_  & \new_[30799]_ ;
  assign \new_[30804]_  = \new_[30803]_  & \new_[30796]_ ;
  assign \new_[30808]_  = ~A199 & A166;
  assign \new_[30809]_  = A168 & \new_[30808]_ ;
  assign \new_[30813]_  = ~A234 & ~A233;
  assign \new_[30814]_  = ~A200 & \new_[30813]_ ;
  assign \new_[30815]_  = \new_[30814]_  & \new_[30809]_ ;
  assign \new_[30819]_  = ~A269 & ~A268;
  assign \new_[30820]_  = ~A266 & \new_[30819]_ ;
  assign \new_[30823]_  = ~A299 & A298;
  assign \new_[30826]_  = A301 & A300;
  assign \new_[30827]_  = \new_[30826]_  & \new_[30823]_ ;
  assign \new_[30828]_  = \new_[30827]_  & \new_[30820]_ ;
  assign \new_[30832]_  = ~A199 & A166;
  assign \new_[30833]_  = A168 & \new_[30832]_ ;
  assign \new_[30837]_  = ~A234 & ~A233;
  assign \new_[30838]_  = ~A200 & \new_[30837]_ ;
  assign \new_[30839]_  = \new_[30838]_  & \new_[30833]_ ;
  assign \new_[30843]_  = ~A269 & ~A268;
  assign \new_[30844]_  = ~A266 & \new_[30843]_ ;
  assign \new_[30847]_  = ~A299 & A298;
  assign \new_[30850]_  = A302 & A300;
  assign \new_[30851]_  = \new_[30850]_  & \new_[30847]_ ;
  assign \new_[30852]_  = \new_[30851]_  & \new_[30844]_ ;
  assign \new_[30856]_  = ~A199 & A166;
  assign \new_[30857]_  = A168 & \new_[30856]_ ;
  assign \new_[30861]_  = ~A233 & ~A232;
  assign \new_[30862]_  = ~A200 & \new_[30861]_ ;
  assign \new_[30863]_  = \new_[30862]_  & \new_[30857]_ ;
  assign \new_[30867]_  = ~A269 & ~A268;
  assign \new_[30868]_  = ~A266 & \new_[30867]_ ;
  assign \new_[30871]_  = ~A299 & A298;
  assign \new_[30874]_  = A301 & A300;
  assign \new_[30875]_  = \new_[30874]_  & \new_[30871]_ ;
  assign \new_[30876]_  = \new_[30875]_  & \new_[30868]_ ;
  assign \new_[30880]_  = ~A199 & A166;
  assign \new_[30881]_  = A168 & \new_[30880]_ ;
  assign \new_[30885]_  = ~A233 & ~A232;
  assign \new_[30886]_  = ~A200 & \new_[30885]_ ;
  assign \new_[30887]_  = \new_[30886]_  & \new_[30881]_ ;
  assign \new_[30891]_  = ~A269 & ~A268;
  assign \new_[30892]_  = ~A266 & \new_[30891]_ ;
  assign \new_[30895]_  = ~A299 & A298;
  assign \new_[30898]_  = A302 & A300;
  assign \new_[30899]_  = \new_[30898]_  & \new_[30895]_ ;
  assign \new_[30900]_  = \new_[30899]_  & \new_[30892]_ ;
  assign \new_[30904]_  = A199 & A167;
  assign \new_[30905]_  = A168 & \new_[30904]_ ;
  assign \new_[30909]_  = A233 & A232;
  assign \new_[30910]_  = A200 & \new_[30909]_ ;
  assign \new_[30911]_  = \new_[30910]_  & \new_[30905]_ ;
  assign \new_[30915]_  = ~A269 & ~A268;
  assign \new_[30916]_  = A265 & \new_[30915]_ ;
  assign \new_[30919]_  = ~A299 & A298;
  assign \new_[30922]_  = A301 & A300;
  assign \new_[30923]_  = \new_[30922]_  & \new_[30919]_ ;
  assign \new_[30924]_  = \new_[30923]_  & \new_[30916]_ ;
  assign \new_[30928]_  = A199 & A167;
  assign \new_[30929]_  = A168 & \new_[30928]_ ;
  assign \new_[30933]_  = A233 & A232;
  assign \new_[30934]_  = A200 & \new_[30933]_ ;
  assign \new_[30935]_  = \new_[30934]_  & \new_[30929]_ ;
  assign \new_[30939]_  = ~A269 & ~A268;
  assign \new_[30940]_  = A265 & \new_[30939]_ ;
  assign \new_[30943]_  = ~A299 & A298;
  assign \new_[30946]_  = A302 & A300;
  assign \new_[30947]_  = \new_[30946]_  & \new_[30943]_ ;
  assign \new_[30948]_  = \new_[30947]_  & \new_[30940]_ ;
  assign \new_[30952]_  = A199 & A167;
  assign \new_[30953]_  = A168 & \new_[30952]_ ;
  assign \new_[30957]_  = ~A235 & ~A233;
  assign \new_[30958]_  = A200 & \new_[30957]_ ;
  assign \new_[30959]_  = \new_[30958]_  & \new_[30953]_ ;
  assign \new_[30963]_  = A266 & A265;
  assign \new_[30964]_  = ~A236 & \new_[30963]_ ;
  assign \new_[30967]_  = ~A299 & A298;
  assign \new_[30970]_  = A301 & A300;
  assign \new_[30971]_  = \new_[30970]_  & \new_[30967]_ ;
  assign \new_[30972]_  = \new_[30971]_  & \new_[30964]_ ;
  assign \new_[30976]_  = A199 & A167;
  assign \new_[30977]_  = A168 & \new_[30976]_ ;
  assign \new_[30981]_  = ~A235 & ~A233;
  assign \new_[30982]_  = A200 & \new_[30981]_ ;
  assign \new_[30983]_  = \new_[30982]_  & \new_[30977]_ ;
  assign \new_[30987]_  = A266 & A265;
  assign \new_[30988]_  = ~A236 & \new_[30987]_ ;
  assign \new_[30991]_  = ~A299 & A298;
  assign \new_[30994]_  = A302 & A300;
  assign \new_[30995]_  = \new_[30994]_  & \new_[30991]_ ;
  assign \new_[30996]_  = \new_[30995]_  & \new_[30988]_ ;
  assign \new_[31000]_  = A199 & A167;
  assign \new_[31001]_  = A168 & \new_[31000]_ ;
  assign \new_[31005]_  = ~A235 & ~A233;
  assign \new_[31006]_  = A200 & \new_[31005]_ ;
  assign \new_[31007]_  = \new_[31006]_  & \new_[31001]_ ;
  assign \new_[31011]_  = ~A267 & ~A266;
  assign \new_[31012]_  = ~A236 & \new_[31011]_ ;
  assign \new_[31015]_  = ~A299 & A298;
  assign \new_[31018]_  = A301 & A300;
  assign \new_[31019]_  = \new_[31018]_  & \new_[31015]_ ;
  assign \new_[31020]_  = \new_[31019]_  & \new_[31012]_ ;
  assign \new_[31024]_  = A199 & A167;
  assign \new_[31025]_  = A168 & \new_[31024]_ ;
  assign \new_[31029]_  = ~A235 & ~A233;
  assign \new_[31030]_  = A200 & \new_[31029]_ ;
  assign \new_[31031]_  = \new_[31030]_  & \new_[31025]_ ;
  assign \new_[31035]_  = ~A267 & ~A266;
  assign \new_[31036]_  = ~A236 & \new_[31035]_ ;
  assign \new_[31039]_  = ~A299 & A298;
  assign \new_[31042]_  = A302 & A300;
  assign \new_[31043]_  = \new_[31042]_  & \new_[31039]_ ;
  assign \new_[31044]_  = \new_[31043]_  & \new_[31036]_ ;
  assign \new_[31048]_  = A199 & A167;
  assign \new_[31049]_  = A168 & \new_[31048]_ ;
  assign \new_[31053]_  = ~A235 & ~A233;
  assign \new_[31054]_  = A200 & \new_[31053]_ ;
  assign \new_[31055]_  = \new_[31054]_  & \new_[31049]_ ;
  assign \new_[31059]_  = ~A266 & ~A265;
  assign \new_[31060]_  = ~A236 & \new_[31059]_ ;
  assign \new_[31063]_  = ~A299 & A298;
  assign \new_[31066]_  = A301 & A300;
  assign \new_[31067]_  = \new_[31066]_  & \new_[31063]_ ;
  assign \new_[31068]_  = \new_[31067]_  & \new_[31060]_ ;
  assign \new_[31072]_  = A199 & A167;
  assign \new_[31073]_  = A168 & \new_[31072]_ ;
  assign \new_[31077]_  = ~A235 & ~A233;
  assign \new_[31078]_  = A200 & \new_[31077]_ ;
  assign \new_[31079]_  = \new_[31078]_  & \new_[31073]_ ;
  assign \new_[31083]_  = ~A266 & ~A265;
  assign \new_[31084]_  = ~A236 & \new_[31083]_ ;
  assign \new_[31087]_  = ~A299 & A298;
  assign \new_[31090]_  = A302 & A300;
  assign \new_[31091]_  = \new_[31090]_  & \new_[31087]_ ;
  assign \new_[31092]_  = \new_[31091]_  & \new_[31084]_ ;
  assign \new_[31096]_  = A199 & A167;
  assign \new_[31097]_  = A168 & \new_[31096]_ ;
  assign \new_[31101]_  = ~A234 & ~A233;
  assign \new_[31102]_  = A200 & \new_[31101]_ ;
  assign \new_[31103]_  = \new_[31102]_  & \new_[31097]_ ;
  assign \new_[31107]_  = ~A269 & ~A268;
  assign \new_[31108]_  = ~A266 & \new_[31107]_ ;
  assign \new_[31111]_  = ~A299 & A298;
  assign \new_[31114]_  = A301 & A300;
  assign \new_[31115]_  = \new_[31114]_  & \new_[31111]_ ;
  assign \new_[31116]_  = \new_[31115]_  & \new_[31108]_ ;
  assign \new_[31120]_  = A199 & A167;
  assign \new_[31121]_  = A168 & \new_[31120]_ ;
  assign \new_[31125]_  = ~A234 & ~A233;
  assign \new_[31126]_  = A200 & \new_[31125]_ ;
  assign \new_[31127]_  = \new_[31126]_  & \new_[31121]_ ;
  assign \new_[31131]_  = ~A269 & ~A268;
  assign \new_[31132]_  = ~A266 & \new_[31131]_ ;
  assign \new_[31135]_  = ~A299 & A298;
  assign \new_[31138]_  = A302 & A300;
  assign \new_[31139]_  = \new_[31138]_  & \new_[31135]_ ;
  assign \new_[31140]_  = \new_[31139]_  & \new_[31132]_ ;
  assign \new_[31144]_  = A199 & A167;
  assign \new_[31145]_  = A168 & \new_[31144]_ ;
  assign \new_[31149]_  = ~A233 & ~A232;
  assign \new_[31150]_  = A200 & \new_[31149]_ ;
  assign \new_[31151]_  = \new_[31150]_  & \new_[31145]_ ;
  assign \new_[31155]_  = ~A269 & ~A268;
  assign \new_[31156]_  = ~A266 & \new_[31155]_ ;
  assign \new_[31159]_  = ~A299 & A298;
  assign \new_[31162]_  = A301 & A300;
  assign \new_[31163]_  = \new_[31162]_  & \new_[31159]_ ;
  assign \new_[31164]_  = \new_[31163]_  & \new_[31156]_ ;
  assign \new_[31168]_  = A199 & A167;
  assign \new_[31169]_  = A168 & \new_[31168]_ ;
  assign \new_[31173]_  = ~A233 & ~A232;
  assign \new_[31174]_  = A200 & \new_[31173]_ ;
  assign \new_[31175]_  = \new_[31174]_  & \new_[31169]_ ;
  assign \new_[31179]_  = ~A269 & ~A268;
  assign \new_[31180]_  = ~A266 & \new_[31179]_ ;
  assign \new_[31183]_  = ~A299 & A298;
  assign \new_[31186]_  = A302 & A300;
  assign \new_[31187]_  = \new_[31186]_  & \new_[31183]_ ;
  assign \new_[31188]_  = \new_[31187]_  & \new_[31180]_ ;
  assign \new_[31192]_  = ~A200 & A167;
  assign \new_[31193]_  = A168 & \new_[31192]_ ;
  assign \new_[31197]_  = A232 & ~A203;
  assign \new_[31198]_  = ~A202 & \new_[31197]_ ;
  assign \new_[31199]_  = \new_[31198]_  & \new_[31193]_ ;
  assign \new_[31203]_  = ~A267 & A265;
  assign \new_[31204]_  = A233 & \new_[31203]_ ;
  assign \new_[31207]_  = ~A299 & A298;
  assign \new_[31210]_  = A301 & A300;
  assign \new_[31211]_  = \new_[31210]_  & \new_[31207]_ ;
  assign \new_[31212]_  = \new_[31211]_  & \new_[31204]_ ;
  assign \new_[31216]_  = ~A200 & A167;
  assign \new_[31217]_  = A168 & \new_[31216]_ ;
  assign \new_[31221]_  = A232 & ~A203;
  assign \new_[31222]_  = ~A202 & \new_[31221]_ ;
  assign \new_[31223]_  = \new_[31222]_  & \new_[31217]_ ;
  assign \new_[31227]_  = ~A267 & A265;
  assign \new_[31228]_  = A233 & \new_[31227]_ ;
  assign \new_[31231]_  = ~A299 & A298;
  assign \new_[31234]_  = A302 & A300;
  assign \new_[31235]_  = \new_[31234]_  & \new_[31231]_ ;
  assign \new_[31236]_  = \new_[31235]_  & \new_[31228]_ ;
  assign \new_[31240]_  = ~A200 & A167;
  assign \new_[31241]_  = A168 & \new_[31240]_ ;
  assign \new_[31245]_  = A232 & ~A203;
  assign \new_[31246]_  = ~A202 & \new_[31245]_ ;
  assign \new_[31247]_  = \new_[31246]_  & \new_[31241]_ ;
  assign \new_[31251]_  = A266 & A265;
  assign \new_[31252]_  = A233 & \new_[31251]_ ;
  assign \new_[31255]_  = ~A299 & A298;
  assign \new_[31258]_  = A301 & A300;
  assign \new_[31259]_  = \new_[31258]_  & \new_[31255]_ ;
  assign \new_[31260]_  = \new_[31259]_  & \new_[31252]_ ;
  assign \new_[31264]_  = ~A200 & A167;
  assign \new_[31265]_  = A168 & \new_[31264]_ ;
  assign \new_[31269]_  = A232 & ~A203;
  assign \new_[31270]_  = ~A202 & \new_[31269]_ ;
  assign \new_[31271]_  = \new_[31270]_  & \new_[31265]_ ;
  assign \new_[31275]_  = A266 & A265;
  assign \new_[31276]_  = A233 & \new_[31275]_ ;
  assign \new_[31279]_  = ~A299 & A298;
  assign \new_[31282]_  = A302 & A300;
  assign \new_[31283]_  = \new_[31282]_  & \new_[31279]_ ;
  assign \new_[31284]_  = \new_[31283]_  & \new_[31276]_ ;
  assign \new_[31288]_  = ~A200 & A167;
  assign \new_[31289]_  = A168 & \new_[31288]_ ;
  assign \new_[31293]_  = A232 & ~A203;
  assign \new_[31294]_  = ~A202 & \new_[31293]_ ;
  assign \new_[31295]_  = \new_[31294]_  & \new_[31289]_ ;
  assign \new_[31299]_  = ~A266 & ~A265;
  assign \new_[31300]_  = A233 & \new_[31299]_ ;
  assign \new_[31303]_  = ~A299 & A298;
  assign \new_[31306]_  = A301 & A300;
  assign \new_[31307]_  = \new_[31306]_  & \new_[31303]_ ;
  assign \new_[31308]_  = \new_[31307]_  & \new_[31300]_ ;
  assign \new_[31312]_  = ~A200 & A167;
  assign \new_[31313]_  = A168 & \new_[31312]_ ;
  assign \new_[31317]_  = A232 & ~A203;
  assign \new_[31318]_  = ~A202 & \new_[31317]_ ;
  assign \new_[31319]_  = \new_[31318]_  & \new_[31313]_ ;
  assign \new_[31323]_  = ~A266 & ~A265;
  assign \new_[31324]_  = A233 & \new_[31323]_ ;
  assign \new_[31327]_  = ~A299 & A298;
  assign \new_[31330]_  = A302 & A300;
  assign \new_[31331]_  = \new_[31330]_  & \new_[31327]_ ;
  assign \new_[31332]_  = \new_[31331]_  & \new_[31324]_ ;
  assign \new_[31336]_  = ~A200 & A167;
  assign \new_[31337]_  = A168 & \new_[31336]_ ;
  assign \new_[31341]_  = ~A233 & ~A203;
  assign \new_[31342]_  = ~A202 & \new_[31341]_ ;
  assign \new_[31343]_  = \new_[31342]_  & \new_[31337]_ ;
  assign \new_[31347]_  = ~A266 & ~A236;
  assign \new_[31348]_  = ~A235 & \new_[31347]_ ;
  assign \new_[31351]_  = ~A269 & ~A268;
  assign \new_[31354]_  = A299 & ~A298;
  assign \new_[31355]_  = \new_[31354]_  & \new_[31351]_ ;
  assign \new_[31356]_  = \new_[31355]_  & \new_[31348]_ ;
  assign \new_[31360]_  = ~A200 & A167;
  assign \new_[31361]_  = A168 & \new_[31360]_ ;
  assign \new_[31365]_  = ~A233 & ~A203;
  assign \new_[31366]_  = ~A202 & \new_[31365]_ ;
  assign \new_[31367]_  = \new_[31366]_  & \new_[31361]_ ;
  assign \new_[31371]_  = A266 & A265;
  assign \new_[31372]_  = ~A234 & \new_[31371]_ ;
  assign \new_[31375]_  = ~A299 & A298;
  assign \new_[31378]_  = A301 & A300;
  assign \new_[31379]_  = \new_[31378]_  & \new_[31375]_ ;
  assign \new_[31380]_  = \new_[31379]_  & \new_[31372]_ ;
  assign \new_[31384]_  = ~A200 & A167;
  assign \new_[31385]_  = A168 & \new_[31384]_ ;
  assign \new_[31389]_  = ~A233 & ~A203;
  assign \new_[31390]_  = ~A202 & \new_[31389]_ ;
  assign \new_[31391]_  = \new_[31390]_  & \new_[31385]_ ;
  assign \new_[31395]_  = A266 & A265;
  assign \new_[31396]_  = ~A234 & \new_[31395]_ ;
  assign \new_[31399]_  = ~A299 & A298;
  assign \new_[31402]_  = A302 & A300;
  assign \new_[31403]_  = \new_[31402]_  & \new_[31399]_ ;
  assign \new_[31404]_  = \new_[31403]_  & \new_[31396]_ ;
  assign \new_[31408]_  = ~A200 & A167;
  assign \new_[31409]_  = A168 & \new_[31408]_ ;
  assign \new_[31413]_  = ~A233 & ~A203;
  assign \new_[31414]_  = ~A202 & \new_[31413]_ ;
  assign \new_[31415]_  = \new_[31414]_  & \new_[31409]_ ;
  assign \new_[31419]_  = ~A267 & ~A266;
  assign \new_[31420]_  = ~A234 & \new_[31419]_ ;
  assign \new_[31423]_  = ~A299 & A298;
  assign \new_[31426]_  = A301 & A300;
  assign \new_[31427]_  = \new_[31426]_  & \new_[31423]_ ;
  assign \new_[31428]_  = \new_[31427]_  & \new_[31420]_ ;
  assign \new_[31432]_  = ~A200 & A167;
  assign \new_[31433]_  = A168 & \new_[31432]_ ;
  assign \new_[31437]_  = ~A233 & ~A203;
  assign \new_[31438]_  = ~A202 & \new_[31437]_ ;
  assign \new_[31439]_  = \new_[31438]_  & \new_[31433]_ ;
  assign \new_[31443]_  = ~A267 & ~A266;
  assign \new_[31444]_  = ~A234 & \new_[31443]_ ;
  assign \new_[31447]_  = ~A299 & A298;
  assign \new_[31450]_  = A302 & A300;
  assign \new_[31451]_  = \new_[31450]_  & \new_[31447]_ ;
  assign \new_[31452]_  = \new_[31451]_  & \new_[31444]_ ;
  assign \new_[31456]_  = ~A200 & A167;
  assign \new_[31457]_  = A168 & \new_[31456]_ ;
  assign \new_[31461]_  = ~A233 & ~A203;
  assign \new_[31462]_  = ~A202 & \new_[31461]_ ;
  assign \new_[31463]_  = \new_[31462]_  & \new_[31457]_ ;
  assign \new_[31467]_  = ~A266 & ~A265;
  assign \new_[31468]_  = ~A234 & \new_[31467]_ ;
  assign \new_[31471]_  = ~A299 & A298;
  assign \new_[31474]_  = A301 & A300;
  assign \new_[31475]_  = \new_[31474]_  & \new_[31471]_ ;
  assign \new_[31476]_  = \new_[31475]_  & \new_[31468]_ ;
  assign \new_[31480]_  = ~A200 & A167;
  assign \new_[31481]_  = A168 & \new_[31480]_ ;
  assign \new_[31485]_  = ~A233 & ~A203;
  assign \new_[31486]_  = ~A202 & \new_[31485]_ ;
  assign \new_[31487]_  = \new_[31486]_  & \new_[31481]_ ;
  assign \new_[31491]_  = ~A266 & ~A265;
  assign \new_[31492]_  = ~A234 & \new_[31491]_ ;
  assign \new_[31495]_  = ~A299 & A298;
  assign \new_[31498]_  = A302 & A300;
  assign \new_[31499]_  = \new_[31498]_  & \new_[31495]_ ;
  assign \new_[31500]_  = \new_[31499]_  & \new_[31492]_ ;
  assign \new_[31504]_  = ~A200 & A167;
  assign \new_[31505]_  = A168 & \new_[31504]_ ;
  assign \new_[31509]_  = A232 & ~A203;
  assign \new_[31510]_  = ~A202 & \new_[31509]_ ;
  assign \new_[31511]_  = \new_[31510]_  & \new_[31505]_ ;
  assign \new_[31515]_  = A235 & A234;
  assign \new_[31516]_  = ~A233 & \new_[31515]_ ;
  assign \new_[31519]_  = ~A266 & A265;
  assign \new_[31522]_  = A268 & A267;
  assign \new_[31523]_  = \new_[31522]_  & \new_[31519]_ ;
  assign \new_[31524]_  = \new_[31523]_  & \new_[31516]_ ;
  assign \new_[31528]_  = ~A200 & A167;
  assign \new_[31529]_  = A168 & \new_[31528]_ ;
  assign \new_[31533]_  = A232 & ~A203;
  assign \new_[31534]_  = ~A202 & \new_[31533]_ ;
  assign \new_[31535]_  = \new_[31534]_  & \new_[31529]_ ;
  assign \new_[31539]_  = A235 & A234;
  assign \new_[31540]_  = ~A233 & \new_[31539]_ ;
  assign \new_[31543]_  = ~A266 & A265;
  assign \new_[31546]_  = A269 & A267;
  assign \new_[31547]_  = \new_[31546]_  & \new_[31543]_ ;
  assign \new_[31548]_  = \new_[31547]_  & \new_[31540]_ ;
  assign \new_[31552]_  = ~A200 & A167;
  assign \new_[31553]_  = A168 & \new_[31552]_ ;
  assign \new_[31557]_  = A232 & ~A203;
  assign \new_[31558]_  = ~A202 & \new_[31557]_ ;
  assign \new_[31559]_  = \new_[31558]_  & \new_[31553]_ ;
  assign \new_[31563]_  = A236 & A234;
  assign \new_[31564]_  = ~A233 & \new_[31563]_ ;
  assign \new_[31567]_  = ~A266 & A265;
  assign \new_[31570]_  = A268 & A267;
  assign \new_[31571]_  = \new_[31570]_  & \new_[31567]_ ;
  assign \new_[31572]_  = \new_[31571]_  & \new_[31564]_ ;
  assign \new_[31576]_  = ~A200 & A167;
  assign \new_[31577]_  = A168 & \new_[31576]_ ;
  assign \new_[31581]_  = A232 & ~A203;
  assign \new_[31582]_  = ~A202 & \new_[31581]_ ;
  assign \new_[31583]_  = \new_[31582]_  & \new_[31577]_ ;
  assign \new_[31587]_  = A236 & A234;
  assign \new_[31588]_  = ~A233 & \new_[31587]_ ;
  assign \new_[31591]_  = ~A266 & A265;
  assign \new_[31594]_  = A269 & A267;
  assign \new_[31595]_  = \new_[31594]_  & \new_[31591]_ ;
  assign \new_[31596]_  = \new_[31595]_  & \new_[31588]_ ;
  assign \new_[31600]_  = ~A200 & A167;
  assign \new_[31601]_  = A168 & \new_[31600]_ ;
  assign \new_[31605]_  = ~A232 & ~A203;
  assign \new_[31606]_  = ~A202 & \new_[31605]_ ;
  assign \new_[31607]_  = \new_[31606]_  & \new_[31601]_ ;
  assign \new_[31611]_  = A266 & A265;
  assign \new_[31612]_  = ~A233 & \new_[31611]_ ;
  assign \new_[31615]_  = ~A299 & A298;
  assign \new_[31618]_  = A301 & A300;
  assign \new_[31619]_  = \new_[31618]_  & \new_[31615]_ ;
  assign \new_[31620]_  = \new_[31619]_  & \new_[31612]_ ;
  assign \new_[31624]_  = ~A200 & A167;
  assign \new_[31625]_  = A168 & \new_[31624]_ ;
  assign \new_[31629]_  = ~A232 & ~A203;
  assign \new_[31630]_  = ~A202 & \new_[31629]_ ;
  assign \new_[31631]_  = \new_[31630]_  & \new_[31625]_ ;
  assign \new_[31635]_  = A266 & A265;
  assign \new_[31636]_  = ~A233 & \new_[31635]_ ;
  assign \new_[31639]_  = ~A299 & A298;
  assign \new_[31642]_  = A302 & A300;
  assign \new_[31643]_  = \new_[31642]_  & \new_[31639]_ ;
  assign \new_[31644]_  = \new_[31643]_  & \new_[31636]_ ;
  assign \new_[31648]_  = ~A200 & A167;
  assign \new_[31649]_  = A168 & \new_[31648]_ ;
  assign \new_[31653]_  = ~A232 & ~A203;
  assign \new_[31654]_  = ~A202 & \new_[31653]_ ;
  assign \new_[31655]_  = \new_[31654]_  & \new_[31649]_ ;
  assign \new_[31659]_  = ~A267 & ~A266;
  assign \new_[31660]_  = ~A233 & \new_[31659]_ ;
  assign \new_[31663]_  = ~A299 & A298;
  assign \new_[31666]_  = A301 & A300;
  assign \new_[31667]_  = \new_[31666]_  & \new_[31663]_ ;
  assign \new_[31668]_  = \new_[31667]_  & \new_[31660]_ ;
  assign \new_[31672]_  = ~A200 & A167;
  assign \new_[31673]_  = A168 & \new_[31672]_ ;
  assign \new_[31677]_  = ~A232 & ~A203;
  assign \new_[31678]_  = ~A202 & \new_[31677]_ ;
  assign \new_[31679]_  = \new_[31678]_  & \new_[31673]_ ;
  assign \new_[31683]_  = ~A267 & ~A266;
  assign \new_[31684]_  = ~A233 & \new_[31683]_ ;
  assign \new_[31687]_  = ~A299 & A298;
  assign \new_[31690]_  = A302 & A300;
  assign \new_[31691]_  = \new_[31690]_  & \new_[31687]_ ;
  assign \new_[31692]_  = \new_[31691]_  & \new_[31684]_ ;
  assign \new_[31696]_  = ~A200 & A167;
  assign \new_[31697]_  = A168 & \new_[31696]_ ;
  assign \new_[31701]_  = ~A232 & ~A203;
  assign \new_[31702]_  = ~A202 & \new_[31701]_ ;
  assign \new_[31703]_  = \new_[31702]_  & \new_[31697]_ ;
  assign \new_[31707]_  = ~A266 & ~A265;
  assign \new_[31708]_  = ~A233 & \new_[31707]_ ;
  assign \new_[31711]_  = ~A299 & A298;
  assign \new_[31714]_  = A301 & A300;
  assign \new_[31715]_  = \new_[31714]_  & \new_[31711]_ ;
  assign \new_[31716]_  = \new_[31715]_  & \new_[31708]_ ;
  assign \new_[31720]_  = ~A200 & A167;
  assign \new_[31721]_  = A168 & \new_[31720]_ ;
  assign \new_[31725]_  = ~A232 & ~A203;
  assign \new_[31726]_  = ~A202 & \new_[31725]_ ;
  assign \new_[31727]_  = \new_[31726]_  & \new_[31721]_ ;
  assign \new_[31731]_  = ~A266 & ~A265;
  assign \new_[31732]_  = ~A233 & \new_[31731]_ ;
  assign \new_[31735]_  = ~A299 & A298;
  assign \new_[31738]_  = A302 & A300;
  assign \new_[31739]_  = \new_[31738]_  & \new_[31735]_ ;
  assign \new_[31740]_  = \new_[31739]_  & \new_[31732]_ ;
  assign \new_[31744]_  = ~A200 & A167;
  assign \new_[31745]_  = A168 & \new_[31744]_ ;
  assign \new_[31749]_  = A233 & A232;
  assign \new_[31750]_  = ~A201 & \new_[31749]_ ;
  assign \new_[31751]_  = \new_[31750]_  & \new_[31745]_ ;
  assign \new_[31755]_  = ~A269 & ~A268;
  assign \new_[31756]_  = A265 & \new_[31755]_ ;
  assign \new_[31759]_  = ~A299 & A298;
  assign \new_[31762]_  = A301 & A300;
  assign \new_[31763]_  = \new_[31762]_  & \new_[31759]_ ;
  assign \new_[31764]_  = \new_[31763]_  & \new_[31756]_ ;
  assign \new_[31768]_  = ~A200 & A167;
  assign \new_[31769]_  = A168 & \new_[31768]_ ;
  assign \new_[31773]_  = A233 & A232;
  assign \new_[31774]_  = ~A201 & \new_[31773]_ ;
  assign \new_[31775]_  = \new_[31774]_  & \new_[31769]_ ;
  assign \new_[31779]_  = ~A269 & ~A268;
  assign \new_[31780]_  = A265 & \new_[31779]_ ;
  assign \new_[31783]_  = ~A299 & A298;
  assign \new_[31786]_  = A302 & A300;
  assign \new_[31787]_  = \new_[31786]_  & \new_[31783]_ ;
  assign \new_[31788]_  = \new_[31787]_  & \new_[31780]_ ;
  assign \new_[31792]_  = ~A200 & A167;
  assign \new_[31793]_  = A168 & \new_[31792]_ ;
  assign \new_[31797]_  = ~A235 & ~A233;
  assign \new_[31798]_  = ~A201 & \new_[31797]_ ;
  assign \new_[31799]_  = \new_[31798]_  & \new_[31793]_ ;
  assign \new_[31803]_  = A266 & A265;
  assign \new_[31804]_  = ~A236 & \new_[31803]_ ;
  assign \new_[31807]_  = ~A299 & A298;
  assign \new_[31810]_  = A301 & A300;
  assign \new_[31811]_  = \new_[31810]_  & \new_[31807]_ ;
  assign \new_[31812]_  = \new_[31811]_  & \new_[31804]_ ;
  assign \new_[31816]_  = ~A200 & A167;
  assign \new_[31817]_  = A168 & \new_[31816]_ ;
  assign \new_[31821]_  = ~A235 & ~A233;
  assign \new_[31822]_  = ~A201 & \new_[31821]_ ;
  assign \new_[31823]_  = \new_[31822]_  & \new_[31817]_ ;
  assign \new_[31827]_  = A266 & A265;
  assign \new_[31828]_  = ~A236 & \new_[31827]_ ;
  assign \new_[31831]_  = ~A299 & A298;
  assign \new_[31834]_  = A302 & A300;
  assign \new_[31835]_  = \new_[31834]_  & \new_[31831]_ ;
  assign \new_[31836]_  = \new_[31835]_  & \new_[31828]_ ;
  assign \new_[31840]_  = ~A200 & A167;
  assign \new_[31841]_  = A168 & \new_[31840]_ ;
  assign \new_[31845]_  = ~A235 & ~A233;
  assign \new_[31846]_  = ~A201 & \new_[31845]_ ;
  assign \new_[31847]_  = \new_[31846]_  & \new_[31841]_ ;
  assign \new_[31851]_  = ~A267 & ~A266;
  assign \new_[31852]_  = ~A236 & \new_[31851]_ ;
  assign \new_[31855]_  = ~A299 & A298;
  assign \new_[31858]_  = A301 & A300;
  assign \new_[31859]_  = \new_[31858]_  & \new_[31855]_ ;
  assign \new_[31860]_  = \new_[31859]_  & \new_[31852]_ ;
  assign \new_[31864]_  = ~A200 & A167;
  assign \new_[31865]_  = A168 & \new_[31864]_ ;
  assign \new_[31869]_  = ~A235 & ~A233;
  assign \new_[31870]_  = ~A201 & \new_[31869]_ ;
  assign \new_[31871]_  = \new_[31870]_  & \new_[31865]_ ;
  assign \new_[31875]_  = ~A267 & ~A266;
  assign \new_[31876]_  = ~A236 & \new_[31875]_ ;
  assign \new_[31879]_  = ~A299 & A298;
  assign \new_[31882]_  = A302 & A300;
  assign \new_[31883]_  = \new_[31882]_  & \new_[31879]_ ;
  assign \new_[31884]_  = \new_[31883]_  & \new_[31876]_ ;
  assign \new_[31888]_  = ~A200 & A167;
  assign \new_[31889]_  = A168 & \new_[31888]_ ;
  assign \new_[31893]_  = ~A235 & ~A233;
  assign \new_[31894]_  = ~A201 & \new_[31893]_ ;
  assign \new_[31895]_  = \new_[31894]_  & \new_[31889]_ ;
  assign \new_[31899]_  = ~A266 & ~A265;
  assign \new_[31900]_  = ~A236 & \new_[31899]_ ;
  assign \new_[31903]_  = ~A299 & A298;
  assign \new_[31906]_  = A301 & A300;
  assign \new_[31907]_  = \new_[31906]_  & \new_[31903]_ ;
  assign \new_[31908]_  = \new_[31907]_  & \new_[31900]_ ;
  assign \new_[31912]_  = ~A200 & A167;
  assign \new_[31913]_  = A168 & \new_[31912]_ ;
  assign \new_[31917]_  = ~A235 & ~A233;
  assign \new_[31918]_  = ~A201 & \new_[31917]_ ;
  assign \new_[31919]_  = \new_[31918]_  & \new_[31913]_ ;
  assign \new_[31923]_  = ~A266 & ~A265;
  assign \new_[31924]_  = ~A236 & \new_[31923]_ ;
  assign \new_[31927]_  = ~A299 & A298;
  assign \new_[31930]_  = A302 & A300;
  assign \new_[31931]_  = \new_[31930]_  & \new_[31927]_ ;
  assign \new_[31932]_  = \new_[31931]_  & \new_[31924]_ ;
  assign \new_[31936]_  = ~A200 & A167;
  assign \new_[31937]_  = A168 & \new_[31936]_ ;
  assign \new_[31941]_  = ~A234 & ~A233;
  assign \new_[31942]_  = ~A201 & \new_[31941]_ ;
  assign \new_[31943]_  = \new_[31942]_  & \new_[31937]_ ;
  assign \new_[31947]_  = ~A269 & ~A268;
  assign \new_[31948]_  = ~A266 & \new_[31947]_ ;
  assign \new_[31951]_  = ~A299 & A298;
  assign \new_[31954]_  = A301 & A300;
  assign \new_[31955]_  = \new_[31954]_  & \new_[31951]_ ;
  assign \new_[31956]_  = \new_[31955]_  & \new_[31948]_ ;
  assign \new_[31960]_  = ~A200 & A167;
  assign \new_[31961]_  = A168 & \new_[31960]_ ;
  assign \new_[31965]_  = ~A234 & ~A233;
  assign \new_[31966]_  = ~A201 & \new_[31965]_ ;
  assign \new_[31967]_  = \new_[31966]_  & \new_[31961]_ ;
  assign \new_[31971]_  = ~A269 & ~A268;
  assign \new_[31972]_  = ~A266 & \new_[31971]_ ;
  assign \new_[31975]_  = ~A299 & A298;
  assign \new_[31978]_  = A302 & A300;
  assign \new_[31979]_  = \new_[31978]_  & \new_[31975]_ ;
  assign \new_[31980]_  = \new_[31979]_  & \new_[31972]_ ;
  assign \new_[31984]_  = ~A200 & A167;
  assign \new_[31985]_  = A168 & \new_[31984]_ ;
  assign \new_[31989]_  = ~A233 & ~A232;
  assign \new_[31990]_  = ~A201 & \new_[31989]_ ;
  assign \new_[31991]_  = \new_[31990]_  & \new_[31985]_ ;
  assign \new_[31995]_  = ~A269 & ~A268;
  assign \new_[31996]_  = ~A266 & \new_[31995]_ ;
  assign \new_[31999]_  = ~A299 & A298;
  assign \new_[32002]_  = A301 & A300;
  assign \new_[32003]_  = \new_[32002]_  & \new_[31999]_ ;
  assign \new_[32004]_  = \new_[32003]_  & \new_[31996]_ ;
  assign \new_[32008]_  = ~A200 & A167;
  assign \new_[32009]_  = A168 & \new_[32008]_ ;
  assign \new_[32013]_  = ~A233 & ~A232;
  assign \new_[32014]_  = ~A201 & \new_[32013]_ ;
  assign \new_[32015]_  = \new_[32014]_  & \new_[32009]_ ;
  assign \new_[32019]_  = ~A269 & ~A268;
  assign \new_[32020]_  = ~A266 & \new_[32019]_ ;
  assign \new_[32023]_  = ~A299 & A298;
  assign \new_[32026]_  = A302 & A300;
  assign \new_[32027]_  = \new_[32026]_  & \new_[32023]_ ;
  assign \new_[32028]_  = \new_[32027]_  & \new_[32020]_ ;
  assign \new_[32032]_  = ~A199 & A167;
  assign \new_[32033]_  = A168 & \new_[32032]_ ;
  assign \new_[32037]_  = A233 & A232;
  assign \new_[32038]_  = ~A200 & \new_[32037]_ ;
  assign \new_[32039]_  = \new_[32038]_  & \new_[32033]_ ;
  assign \new_[32043]_  = ~A269 & ~A268;
  assign \new_[32044]_  = A265 & \new_[32043]_ ;
  assign \new_[32047]_  = ~A299 & A298;
  assign \new_[32050]_  = A301 & A300;
  assign \new_[32051]_  = \new_[32050]_  & \new_[32047]_ ;
  assign \new_[32052]_  = \new_[32051]_  & \new_[32044]_ ;
  assign \new_[32056]_  = ~A199 & A167;
  assign \new_[32057]_  = A168 & \new_[32056]_ ;
  assign \new_[32061]_  = A233 & A232;
  assign \new_[32062]_  = ~A200 & \new_[32061]_ ;
  assign \new_[32063]_  = \new_[32062]_  & \new_[32057]_ ;
  assign \new_[32067]_  = ~A269 & ~A268;
  assign \new_[32068]_  = A265 & \new_[32067]_ ;
  assign \new_[32071]_  = ~A299 & A298;
  assign \new_[32074]_  = A302 & A300;
  assign \new_[32075]_  = \new_[32074]_  & \new_[32071]_ ;
  assign \new_[32076]_  = \new_[32075]_  & \new_[32068]_ ;
  assign \new_[32080]_  = ~A199 & A167;
  assign \new_[32081]_  = A168 & \new_[32080]_ ;
  assign \new_[32085]_  = ~A235 & ~A233;
  assign \new_[32086]_  = ~A200 & \new_[32085]_ ;
  assign \new_[32087]_  = \new_[32086]_  & \new_[32081]_ ;
  assign \new_[32091]_  = A266 & A265;
  assign \new_[32092]_  = ~A236 & \new_[32091]_ ;
  assign \new_[32095]_  = ~A299 & A298;
  assign \new_[32098]_  = A301 & A300;
  assign \new_[32099]_  = \new_[32098]_  & \new_[32095]_ ;
  assign \new_[32100]_  = \new_[32099]_  & \new_[32092]_ ;
  assign \new_[32104]_  = ~A199 & A167;
  assign \new_[32105]_  = A168 & \new_[32104]_ ;
  assign \new_[32109]_  = ~A235 & ~A233;
  assign \new_[32110]_  = ~A200 & \new_[32109]_ ;
  assign \new_[32111]_  = \new_[32110]_  & \new_[32105]_ ;
  assign \new_[32115]_  = A266 & A265;
  assign \new_[32116]_  = ~A236 & \new_[32115]_ ;
  assign \new_[32119]_  = ~A299 & A298;
  assign \new_[32122]_  = A302 & A300;
  assign \new_[32123]_  = \new_[32122]_  & \new_[32119]_ ;
  assign \new_[32124]_  = \new_[32123]_  & \new_[32116]_ ;
  assign \new_[32128]_  = ~A199 & A167;
  assign \new_[32129]_  = A168 & \new_[32128]_ ;
  assign \new_[32133]_  = ~A235 & ~A233;
  assign \new_[32134]_  = ~A200 & \new_[32133]_ ;
  assign \new_[32135]_  = \new_[32134]_  & \new_[32129]_ ;
  assign \new_[32139]_  = ~A267 & ~A266;
  assign \new_[32140]_  = ~A236 & \new_[32139]_ ;
  assign \new_[32143]_  = ~A299 & A298;
  assign \new_[32146]_  = A301 & A300;
  assign \new_[32147]_  = \new_[32146]_  & \new_[32143]_ ;
  assign \new_[32148]_  = \new_[32147]_  & \new_[32140]_ ;
  assign \new_[32152]_  = ~A199 & A167;
  assign \new_[32153]_  = A168 & \new_[32152]_ ;
  assign \new_[32157]_  = ~A235 & ~A233;
  assign \new_[32158]_  = ~A200 & \new_[32157]_ ;
  assign \new_[32159]_  = \new_[32158]_  & \new_[32153]_ ;
  assign \new_[32163]_  = ~A267 & ~A266;
  assign \new_[32164]_  = ~A236 & \new_[32163]_ ;
  assign \new_[32167]_  = ~A299 & A298;
  assign \new_[32170]_  = A302 & A300;
  assign \new_[32171]_  = \new_[32170]_  & \new_[32167]_ ;
  assign \new_[32172]_  = \new_[32171]_  & \new_[32164]_ ;
  assign \new_[32176]_  = ~A199 & A167;
  assign \new_[32177]_  = A168 & \new_[32176]_ ;
  assign \new_[32181]_  = ~A235 & ~A233;
  assign \new_[32182]_  = ~A200 & \new_[32181]_ ;
  assign \new_[32183]_  = \new_[32182]_  & \new_[32177]_ ;
  assign \new_[32187]_  = ~A266 & ~A265;
  assign \new_[32188]_  = ~A236 & \new_[32187]_ ;
  assign \new_[32191]_  = ~A299 & A298;
  assign \new_[32194]_  = A301 & A300;
  assign \new_[32195]_  = \new_[32194]_  & \new_[32191]_ ;
  assign \new_[32196]_  = \new_[32195]_  & \new_[32188]_ ;
  assign \new_[32200]_  = ~A199 & A167;
  assign \new_[32201]_  = A168 & \new_[32200]_ ;
  assign \new_[32205]_  = ~A235 & ~A233;
  assign \new_[32206]_  = ~A200 & \new_[32205]_ ;
  assign \new_[32207]_  = \new_[32206]_  & \new_[32201]_ ;
  assign \new_[32211]_  = ~A266 & ~A265;
  assign \new_[32212]_  = ~A236 & \new_[32211]_ ;
  assign \new_[32215]_  = ~A299 & A298;
  assign \new_[32218]_  = A302 & A300;
  assign \new_[32219]_  = \new_[32218]_  & \new_[32215]_ ;
  assign \new_[32220]_  = \new_[32219]_  & \new_[32212]_ ;
  assign \new_[32224]_  = ~A199 & A167;
  assign \new_[32225]_  = A168 & \new_[32224]_ ;
  assign \new_[32229]_  = ~A234 & ~A233;
  assign \new_[32230]_  = ~A200 & \new_[32229]_ ;
  assign \new_[32231]_  = \new_[32230]_  & \new_[32225]_ ;
  assign \new_[32235]_  = ~A269 & ~A268;
  assign \new_[32236]_  = ~A266 & \new_[32235]_ ;
  assign \new_[32239]_  = ~A299 & A298;
  assign \new_[32242]_  = A301 & A300;
  assign \new_[32243]_  = \new_[32242]_  & \new_[32239]_ ;
  assign \new_[32244]_  = \new_[32243]_  & \new_[32236]_ ;
  assign \new_[32248]_  = ~A199 & A167;
  assign \new_[32249]_  = A168 & \new_[32248]_ ;
  assign \new_[32253]_  = ~A234 & ~A233;
  assign \new_[32254]_  = ~A200 & \new_[32253]_ ;
  assign \new_[32255]_  = \new_[32254]_  & \new_[32249]_ ;
  assign \new_[32259]_  = ~A269 & ~A268;
  assign \new_[32260]_  = ~A266 & \new_[32259]_ ;
  assign \new_[32263]_  = ~A299 & A298;
  assign \new_[32266]_  = A302 & A300;
  assign \new_[32267]_  = \new_[32266]_  & \new_[32263]_ ;
  assign \new_[32268]_  = \new_[32267]_  & \new_[32260]_ ;
  assign \new_[32272]_  = ~A199 & A167;
  assign \new_[32273]_  = A168 & \new_[32272]_ ;
  assign \new_[32277]_  = ~A233 & ~A232;
  assign \new_[32278]_  = ~A200 & \new_[32277]_ ;
  assign \new_[32279]_  = \new_[32278]_  & \new_[32273]_ ;
  assign \new_[32283]_  = ~A269 & ~A268;
  assign \new_[32284]_  = ~A266 & \new_[32283]_ ;
  assign \new_[32287]_  = ~A299 & A298;
  assign \new_[32290]_  = A301 & A300;
  assign \new_[32291]_  = \new_[32290]_  & \new_[32287]_ ;
  assign \new_[32292]_  = \new_[32291]_  & \new_[32284]_ ;
  assign \new_[32296]_  = ~A199 & A167;
  assign \new_[32297]_  = A168 & \new_[32296]_ ;
  assign \new_[32301]_  = ~A233 & ~A232;
  assign \new_[32302]_  = ~A200 & \new_[32301]_ ;
  assign \new_[32303]_  = \new_[32302]_  & \new_[32297]_ ;
  assign \new_[32307]_  = ~A269 & ~A268;
  assign \new_[32308]_  = ~A266 & \new_[32307]_ ;
  assign \new_[32311]_  = ~A299 & A298;
  assign \new_[32314]_  = A302 & A300;
  assign \new_[32315]_  = \new_[32314]_  & \new_[32311]_ ;
  assign \new_[32316]_  = \new_[32315]_  & \new_[32308]_ ;
  assign \new_[32320]_  = ~A166 & ~A167;
  assign \new_[32321]_  = A170 & \new_[32320]_ ;
  assign \new_[32325]_  = A232 & A200;
  assign \new_[32326]_  = ~A199 & \new_[32325]_ ;
  assign \new_[32327]_  = \new_[32326]_  & \new_[32321]_ ;
  assign \new_[32331]_  = ~A267 & A265;
  assign \new_[32332]_  = A233 & \new_[32331]_ ;
  assign \new_[32335]_  = ~A299 & A298;
  assign \new_[32338]_  = A301 & A300;
  assign \new_[32339]_  = \new_[32338]_  & \new_[32335]_ ;
  assign \new_[32340]_  = \new_[32339]_  & \new_[32332]_ ;
  assign \new_[32344]_  = ~A166 & ~A167;
  assign \new_[32345]_  = A170 & \new_[32344]_ ;
  assign \new_[32349]_  = A232 & A200;
  assign \new_[32350]_  = ~A199 & \new_[32349]_ ;
  assign \new_[32351]_  = \new_[32350]_  & \new_[32345]_ ;
  assign \new_[32355]_  = ~A267 & A265;
  assign \new_[32356]_  = A233 & \new_[32355]_ ;
  assign \new_[32359]_  = ~A299 & A298;
  assign \new_[32362]_  = A302 & A300;
  assign \new_[32363]_  = \new_[32362]_  & \new_[32359]_ ;
  assign \new_[32364]_  = \new_[32363]_  & \new_[32356]_ ;
  assign \new_[32368]_  = ~A166 & ~A167;
  assign \new_[32369]_  = A170 & \new_[32368]_ ;
  assign \new_[32373]_  = A232 & A200;
  assign \new_[32374]_  = ~A199 & \new_[32373]_ ;
  assign \new_[32375]_  = \new_[32374]_  & \new_[32369]_ ;
  assign \new_[32379]_  = A266 & A265;
  assign \new_[32380]_  = A233 & \new_[32379]_ ;
  assign \new_[32383]_  = ~A299 & A298;
  assign \new_[32386]_  = A301 & A300;
  assign \new_[32387]_  = \new_[32386]_  & \new_[32383]_ ;
  assign \new_[32388]_  = \new_[32387]_  & \new_[32380]_ ;
  assign \new_[32392]_  = ~A166 & ~A167;
  assign \new_[32393]_  = A170 & \new_[32392]_ ;
  assign \new_[32397]_  = A232 & A200;
  assign \new_[32398]_  = ~A199 & \new_[32397]_ ;
  assign \new_[32399]_  = \new_[32398]_  & \new_[32393]_ ;
  assign \new_[32403]_  = A266 & A265;
  assign \new_[32404]_  = A233 & \new_[32403]_ ;
  assign \new_[32407]_  = ~A299 & A298;
  assign \new_[32410]_  = A302 & A300;
  assign \new_[32411]_  = \new_[32410]_  & \new_[32407]_ ;
  assign \new_[32412]_  = \new_[32411]_  & \new_[32404]_ ;
  assign \new_[32416]_  = ~A166 & ~A167;
  assign \new_[32417]_  = A170 & \new_[32416]_ ;
  assign \new_[32421]_  = A232 & A200;
  assign \new_[32422]_  = ~A199 & \new_[32421]_ ;
  assign \new_[32423]_  = \new_[32422]_  & \new_[32417]_ ;
  assign \new_[32427]_  = ~A266 & ~A265;
  assign \new_[32428]_  = A233 & \new_[32427]_ ;
  assign \new_[32431]_  = ~A299 & A298;
  assign \new_[32434]_  = A301 & A300;
  assign \new_[32435]_  = \new_[32434]_  & \new_[32431]_ ;
  assign \new_[32436]_  = \new_[32435]_  & \new_[32428]_ ;
  assign \new_[32440]_  = ~A166 & ~A167;
  assign \new_[32441]_  = A170 & \new_[32440]_ ;
  assign \new_[32445]_  = A232 & A200;
  assign \new_[32446]_  = ~A199 & \new_[32445]_ ;
  assign \new_[32447]_  = \new_[32446]_  & \new_[32441]_ ;
  assign \new_[32451]_  = ~A266 & ~A265;
  assign \new_[32452]_  = A233 & \new_[32451]_ ;
  assign \new_[32455]_  = ~A299 & A298;
  assign \new_[32458]_  = A302 & A300;
  assign \new_[32459]_  = \new_[32458]_  & \new_[32455]_ ;
  assign \new_[32460]_  = \new_[32459]_  & \new_[32452]_ ;
  assign \new_[32464]_  = ~A166 & ~A167;
  assign \new_[32465]_  = A170 & \new_[32464]_ ;
  assign \new_[32469]_  = ~A233 & A200;
  assign \new_[32470]_  = ~A199 & \new_[32469]_ ;
  assign \new_[32471]_  = \new_[32470]_  & \new_[32465]_ ;
  assign \new_[32475]_  = ~A266 & ~A236;
  assign \new_[32476]_  = ~A235 & \new_[32475]_ ;
  assign \new_[32479]_  = ~A269 & ~A268;
  assign \new_[32482]_  = A299 & ~A298;
  assign \new_[32483]_  = \new_[32482]_  & \new_[32479]_ ;
  assign \new_[32484]_  = \new_[32483]_  & \new_[32476]_ ;
  assign \new_[32488]_  = ~A166 & ~A167;
  assign \new_[32489]_  = A170 & \new_[32488]_ ;
  assign \new_[32493]_  = ~A233 & A200;
  assign \new_[32494]_  = ~A199 & \new_[32493]_ ;
  assign \new_[32495]_  = \new_[32494]_  & \new_[32489]_ ;
  assign \new_[32499]_  = A266 & A265;
  assign \new_[32500]_  = ~A234 & \new_[32499]_ ;
  assign \new_[32503]_  = ~A299 & A298;
  assign \new_[32506]_  = A301 & A300;
  assign \new_[32507]_  = \new_[32506]_  & \new_[32503]_ ;
  assign \new_[32508]_  = \new_[32507]_  & \new_[32500]_ ;
  assign \new_[32512]_  = ~A166 & ~A167;
  assign \new_[32513]_  = A170 & \new_[32512]_ ;
  assign \new_[32517]_  = ~A233 & A200;
  assign \new_[32518]_  = ~A199 & \new_[32517]_ ;
  assign \new_[32519]_  = \new_[32518]_  & \new_[32513]_ ;
  assign \new_[32523]_  = A266 & A265;
  assign \new_[32524]_  = ~A234 & \new_[32523]_ ;
  assign \new_[32527]_  = ~A299 & A298;
  assign \new_[32530]_  = A302 & A300;
  assign \new_[32531]_  = \new_[32530]_  & \new_[32527]_ ;
  assign \new_[32532]_  = \new_[32531]_  & \new_[32524]_ ;
  assign \new_[32536]_  = ~A166 & ~A167;
  assign \new_[32537]_  = A170 & \new_[32536]_ ;
  assign \new_[32541]_  = ~A233 & A200;
  assign \new_[32542]_  = ~A199 & \new_[32541]_ ;
  assign \new_[32543]_  = \new_[32542]_  & \new_[32537]_ ;
  assign \new_[32547]_  = ~A267 & ~A266;
  assign \new_[32548]_  = ~A234 & \new_[32547]_ ;
  assign \new_[32551]_  = ~A299 & A298;
  assign \new_[32554]_  = A301 & A300;
  assign \new_[32555]_  = \new_[32554]_  & \new_[32551]_ ;
  assign \new_[32556]_  = \new_[32555]_  & \new_[32548]_ ;
  assign \new_[32560]_  = ~A166 & ~A167;
  assign \new_[32561]_  = A170 & \new_[32560]_ ;
  assign \new_[32565]_  = ~A233 & A200;
  assign \new_[32566]_  = ~A199 & \new_[32565]_ ;
  assign \new_[32567]_  = \new_[32566]_  & \new_[32561]_ ;
  assign \new_[32571]_  = ~A267 & ~A266;
  assign \new_[32572]_  = ~A234 & \new_[32571]_ ;
  assign \new_[32575]_  = ~A299 & A298;
  assign \new_[32578]_  = A302 & A300;
  assign \new_[32579]_  = \new_[32578]_  & \new_[32575]_ ;
  assign \new_[32580]_  = \new_[32579]_  & \new_[32572]_ ;
  assign \new_[32584]_  = ~A166 & ~A167;
  assign \new_[32585]_  = A170 & \new_[32584]_ ;
  assign \new_[32589]_  = ~A233 & A200;
  assign \new_[32590]_  = ~A199 & \new_[32589]_ ;
  assign \new_[32591]_  = \new_[32590]_  & \new_[32585]_ ;
  assign \new_[32595]_  = ~A266 & ~A265;
  assign \new_[32596]_  = ~A234 & \new_[32595]_ ;
  assign \new_[32599]_  = ~A299 & A298;
  assign \new_[32602]_  = A301 & A300;
  assign \new_[32603]_  = \new_[32602]_  & \new_[32599]_ ;
  assign \new_[32604]_  = \new_[32603]_  & \new_[32596]_ ;
  assign \new_[32608]_  = ~A166 & ~A167;
  assign \new_[32609]_  = A170 & \new_[32608]_ ;
  assign \new_[32613]_  = ~A233 & A200;
  assign \new_[32614]_  = ~A199 & \new_[32613]_ ;
  assign \new_[32615]_  = \new_[32614]_  & \new_[32609]_ ;
  assign \new_[32619]_  = ~A266 & ~A265;
  assign \new_[32620]_  = ~A234 & \new_[32619]_ ;
  assign \new_[32623]_  = ~A299 & A298;
  assign \new_[32626]_  = A302 & A300;
  assign \new_[32627]_  = \new_[32626]_  & \new_[32623]_ ;
  assign \new_[32628]_  = \new_[32627]_  & \new_[32620]_ ;
  assign \new_[32632]_  = ~A166 & ~A167;
  assign \new_[32633]_  = A170 & \new_[32632]_ ;
  assign \new_[32637]_  = A232 & A200;
  assign \new_[32638]_  = ~A199 & \new_[32637]_ ;
  assign \new_[32639]_  = \new_[32638]_  & \new_[32633]_ ;
  assign \new_[32643]_  = A235 & A234;
  assign \new_[32644]_  = ~A233 & \new_[32643]_ ;
  assign \new_[32647]_  = ~A266 & A265;
  assign \new_[32650]_  = A268 & A267;
  assign \new_[32651]_  = \new_[32650]_  & \new_[32647]_ ;
  assign \new_[32652]_  = \new_[32651]_  & \new_[32644]_ ;
  assign \new_[32656]_  = ~A166 & ~A167;
  assign \new_[32657]_  = A170 & \new_[32656]_ ;
  assign \new_[32661]_  = A232 & A200;
  assign \new_[32662]_  = ~A199 & \new_[32661]_ ;
  assign \new_[32663]_  = \new_[32662]_  & \new_[32657]_ ;
  assign \new_[32667]_  = A235 & A234;
  assign \new_[32668]_  = ~A233 & \new_[32667]_ ;
  assign \new_[32671]_  = ~A266 & A265;
  assign \new_[32674]_  = A269 & A267;
  assign \new_[32675]_  = \new_[32674]_  & \new_[32671]_ ;
  assign \new_[32676]_  = \new_[32675]_  & \new_[32668]_ ;
  assign \new_[32680]_  = ~A166 & ~A167;
  assign \new_[32681]_  = A170 & \new_[32680]_ ;
  assign \new_[32685]_  = A232 & A200;
  assign \new_[32686]_  = ~A199 & \new_[32685]_ ;
  assign \new_[32687]_  = \new_[32686]_  & \new_[32681]_ ;
  assign \new_[32691]_  = A236 & A234;
  assign \new_[32692]_  = ~A233 & \new_[32691]_ ;
  assign \new_[32695]_  = ~A266 & A265;
  assign \new_[32698]_  = A268 & A267;
  assign \new_[32699]_  = \new_[32698]_  & \new_[32695]_ ;
  assign \new_[32700]_  = \new_[32699]_  & \new_[32692]_ ;
  assign \new_[32704]_  = ~A166 & ~A167;
  assign \new_[32705]_  = A170 & \new_[32704]_ ;
  assign \new_[32709]_  = A232 & A200;
  assign \new_[32710]_  = ~A199 & \new_[32709]_ ;
  assign \new_[32711]_  = \new_[32710]_  & \new_[32705]_ ;
  assign \new_[32715]_  = A236 & A234;
  assign \new_[32716]_  = ~A233 & \new_[32715]_ ;
  assign \new_[32719]_  = ~A266 & A265;
  assign \new_[32722]_  = A269 & A267;
  assign \new_[32723]_  = \new_[32722]_  & \new_[32719]_ ;
  assign \new_[32724]_  = \new_[32723]_  & \new_[32716]_ ;
  assign \new_[32728]_  = ~A166 & ~A167;
  assign \new_[32729]_  = A170 & \new_[32728]_ ;
  assign \new_[32733]_  = ~A232 & A200;
  assign \new_[32734]_  = ~A199 & \new_[32733]_ ;
  assign \new_[32735]_  = \new_[32734]_  & \new_[32729]_ ;
  assign \new_[32739]_  = A266 & A265;
  assign \new_[32740]_  = ~A233 & \new_[32739]_ ;
  assign \new_[32743]_  = ~A299 & A298;
  assign \new_[32746]_  = A301 & A300;
  assign \new_[32747]_  = \new_[32746]_  & \new_[32743]_ ;
  assign \new_[32748]_  = \new_[32747]_  & \new_[32740]_ ;
  assign \new_[32752]_  = ~A166 & ~A167;
  assign \new_[32753]_  = A170 & \new_[32752]_ ;
  assign \new_[32757]_  = ~A232 & A200;
  assign \new_[32758]_  = ~A199 & \new_[32757]_ ;
  assign \new_[32759]_  = \new_[32758]_  & \new_[32753]_ ;
  assign \new_[32763]_  = A266 & A265;
  assign \new_[32764]_  = ~A233 & \new_[32763]_ ;
  assign \new_[32767]_  = ~A299 & A298;
  assign \new_[32770]_  = A302 & A300;
  assign \new_[32771]_  = \new_[32770]_  & \new_[32767]_ ;
  assign \new_[32772]_  = \new_[32771]_  & \new_[32764]_ ;
  assign \new_[32776]_  = ~A166 & ~A167;
  assign \new_[32777]_  = A170 & \new_[32776]_ ;
  assign \new_[32781]_  = ~A232 & A200;
  assign \new_[32782]_  = ~A199 & \new_[32781]_ ;
  assign \new_[32783]_  = \new_[32782]_  & \new_[32777]_ ;
  assign \new_[32787]_  = ~A267 & ~A266;
  assign \new_[32788]_  = ~A233 & \new_[32787]_ ;
  assign \new_[32791]_  = ~A299 & A298;
  assign \new_[32794]_  = A301 & A300;
  assign \new_[32795]_  = \new_[32794]_  & \new_[32791]_ ;
  assign \new_[32796]_  = \new_[32795]_  & \new_[32788]_ ;
  assign \new_[32800]_  = ~A166 & ~A167;
  assign \new_[32801]_  = A170 & \new_[32800]_ ;
  assign \new_[32805]_  = ~A232 & A200;
  assign \new_[32806]_  = ~A199 & \new_[32805]_ ;
  assign \new_[32807]_  = \new_[32806]_  & \new_[32801]_ ;
  assign \new_[32811]_  = ~A267 & ~A266;
  assign \new_[32812]_  = ~A233 & \new_[32811]_ ;
  assign \new_[32815]_  = ~A299 & A298;
  assign \new_[32818]_  = A302 & A300;
  assign \new_[32819]_  = \new_[32818]_  & \new_[32815]_ ;
  assign \new_[32820]_  = \new_[32819]_  & \new_[32812]_ ;
  assign \new_[32824]_  = ~A166 & ~A167;
  assign \new_[32825]_  = A170 & \new_[32824]_ ;
  assign \new_[32829]_  = ~A232 & A200;
  assign \new_[32830]_  = ~A199 & \new_[32829]_ ;
  assign \new_[32831]_  = \new_[32830]_  & \new_[32825]_ ;
  assign \new_[32835]_  = ~A266 & ~A265;
  assign \new_[32836]_  = ~A233 & \new_[32835]_ ;
  assign \new_[32839]_  = ~A299 & A298;
  assign \new_[32842]_  = A301 & A300;
  assign \new_[32843]_  = \new_[32842]_  & \new_[32839]_ ;
  assign \new_[32844]_  = \new_[32843]_  & \new_[32836]_ ;
  assign \new_[32848]_  = ~A166 & ~A167;
  assign \new_[32849]_  = A170 & \new_[32848]_ ;
  assign \new_[32853]_  = ~A232 & A200;
  assign \new_[32854]_  = ~A199 & \new_[32853]_ ;
  assign \new_[32855]_  = \new_[32854]_  & \new_[32849]_ ;
  assign \new_[32859]_  = ~A266 & ~A265;
  assign \new_[32860]_  = ~A233 & \new_[32859]_ ;
  assign \new_[32863]_  = ~A299 & A298;
  assign \new_[32866]_  = A302 & A300;
  assign \new_[32867]_  = \new_[32866]_  & \new_[32863]_ ;
  assign \new_[32868]_  = \new_[32867]_  & \new_[32860]_ ;
  assign \new_[32872]_  = ~A166 & ~A167;
  assign \new_[32873]_  = A170 & \new_[32872]_ ;
  assign \new_[32877]_  = A201 & ~A200;
  assign \new_[32878]_  = A199 & \new_[32877]_ ;
  assign \new_[32879]_  = \new_[32878]_  & \new_[32873]_ ;
  assign \new_[32883]_  = A233 & A232;
  assign \new_[32884]_  = A202 & \new_[32883]_ ;
  assign \new_[32887]_  = ~A267 & A265;
  assign \new_[32890]_  = A299 & ~A298;
  assign \new_[32891]_  = \new_[32890]_  & \new_[32887]_ ;
  assign \new_[32892]_  = \new_[32891]_  & \new_[32884]_ ;
  assign \new_[32896]_  = ~A166 & ~A167;
  assign \new_[32897]_  = A170 & \new_[32896]_ ;
  assign \new_[32901]_  = A201 & ~A200;
  assign \new_[32902]_  = A199 & \new_[32901]_ ;
  assign \new_[32903]_  = \new_[32902]_  & \new_[32897]_ ;
  assign \new_[32907]_  = A233 & A232;
  assign \new_[32908]_  = A202 & \new_[32907]_ ;
  assign \new_[32911]_  = A266 & A265;
  assign \new_[32914]_  = A299 & ~A298;
  assign \new_[32915]_  = \new_[32914]_  & \new_[32911]_ ;
  assign \new_[32916]_  = \new_[32915]_  & \new_[32908]_ ;
  assign \new_[32920]_  = ~A166 & ~A167;
  assign \new_[32921]_  = A170 & \new_[32920]_ ;
  assign \new_[32925]_  = A201 & ~A200;
  assign \new_[32926]_  = A199 & \new_[32925]_ ;
  assign \new_[32927]_  = \new_[32926]_  & \new_[32921]_ ;
  assign \new_[32931]_  = A233 & A232;
  assign \new_[32932]_  = A202 & \new_[32931]_ ;
  assign \new_[32935]_  = ~A266 & ~A265;
  assign \new_[32938]_  = A299 & ~A298;
  assign \new_[32939]_  = \new_[32938]_  & \new_[32935]_ ;
  assign \new_[32940]_  = \new_[32939]_  & \new_[32932]_ ;
  assign \new_[32944]_  = ~A166 & ~A167;
  assign \new_[32945]_  = A170 & \new_[32944]_ ;
  assign \new_[32949]_  = A201 & ~A200;
  assign \new_[32950]_  = A199 & \new_[32949]_ ;
  assign \new_[32951]_  = \new_[32950]_  & \new_[32945]_ ;
  assign \new_[32955]_  = A233 & ~A232;
  assign \new_[32956]_  = A202 & \new_[32955]_ ;
  assign \new_[32959]_  = ~A266 & A265;
  assign \new_[32962]_  = A268 & A267;
  assign \new_[32963]_  = \new_[32962]_  & \new_[32959]_ ;
  assign \new_[32964]_  = \new_[32963]_  & \new_[32956]_ ;
  assign \new_[32968]_  = ~A166 & ~A167;
  assign \new_[32969]_  = A170 & \new_[32968]_ ;
  assign \new_[32973]_  = A201 & ~A200;
  assign \new_[32974]_  = A199 & \new_[32973]_ ;
  assign \new_[32975]_  = \new_[32974]_  & \new_[32969]_ ;
  assign \new_[32979]_  = A233 & ~A232;
  assign \new_[32980]_  = A202 & \new_[32979]_ ;
  assign \new_[32983]_  = ~A266 & A265;
  assign \new_[32986]_  = A269 & A267;
  assign \new_[32987]_  = \new_[32986]_  & \new_[32983]_ ;
  assign \new_[32988]_  = \new_[32987]_  & \new_[32980]_ ;
  assign \new_[32992]_  = ~A166 & ~A167;
  assign \new_[32993]_  = A170 & \new_[32992]_ ;
  assign \new_[32997]_  = A201 & ~A200;
  assign \new_[32998]_  = A199 & \new_[32997]_ ;
  assign \new_[32999]_  = \new_[32998]_  & \new_[32993]_ ;
  assign \new_[33003]_  = ~A234 & ~A233;
  assign \new_[33004]_  = A202 & \new_[33003]_ ;
  assign \new_[33007]_  = A266 & A265;
  assign \new_[33010]_  = A299 & ~A298;
  assign \new_[33011]_  = \new_[33010]_  & \new_[33007]_ ;
  assign \new_[33012]_  = \new_[33011]_  & \new_[33004]_ ;
  assign \new_[33016]_  = ~A166 & ~A167;
  assign \new_[33017]_  = A170 & \new_[33016]_ ;
  assign \new_[33021]_  = A201 & ~A200;
  assign \new_[33022]_  = A199 & \new_[33021]_ ;
  assign \new_[33023]_  = \new_[33022]_  & \new_[33017]_ ;
  assign \new_[33027]_  = ~A234 & ~A233;
  assign \new_[33028]_  = A202 & \new_[33027]_ ;
  assign \new_[33031]_  = ~A267 & ~A266;
  assign \new_[33034]_  = A299 & ~A298;
  assign \new_[33035]_  = \new_[33034]_  & \new_[33031]_ ;
  assign \new_[33036]_  = \new_[33035]_  & \new_[33028]_ ;
  assign \new_[33040]_  = ~A166 & ~A167;
  assign \new_[33041]_  = A170 & \new_[33040]_ ;
  assign \new_[33045]_  = A201 & ~A200;
  assign \new_[33046]_  = A199 & \new_[33045]_ ;
  assign \new_[33047]_  = \new_[33046]_  & \new_[33041]_ ;
  assign \new_[33051]_  = ~A234 & ~A233;
  assign \new_[33052]_  = A202 & \new_[33051]_ ;
  assign \new_[33055]_  = ~A266 & ~A265;
  assign \new_[33058]_  = A299 & ~A298;
  assign \new_[33059]_  = \new_[33058]_  & \new_[33055]_ ;
  assign \new_[33060]_  = \new_[33059]_  & \new_[33052]_ ;
  assign \new_[33064]_  = ~A166 & ~A167;
  assign \new_[33065]_  = A170 & \new_[33064]_ ;
  assign \new_[33069]_  = A201 & ~A200;
  assign \new_[33070]_  = A199 & \new_[33069]_ ;
  assign \new_[33071]_  = \new_[33070]_  & \new_[33065]_ ;
  assign \new_[33075]_  = ~A233 & A232;
  assign \new_[33076]_  = A202 & \new_[33075]_ ;
  assign \new_[33079]_  = A235 & A234;
  assign \new_[33082]_  = ~A300 & A298;
  assign \new_[33083]_  = \new_[33082]_  & \new_[33079]_ ;
  assign \new_[33084]_  = \new_[33083]_  & \new_[33076]_ ;
  assign \new_[33088]_  = ~A166 & ~A167;
  assign \new_[33089]_  = A170 & \new_[33088]_ ;
  assign \new_[33093]_  = A201 & ~A200;
  assign \new_[33094]_  = A199 & \new_[33093]_ ;
  assign \new_[33095]_  = \new_[33094]_  & \new_[33089]_ ;
  assign \new_[33099]_  = ~A233 & A232;
  assign \new_[33100]_  = A202 & \new_[33099]_ ;
  assign \new_[33103]_  = A235 & A234;
  assign \new_[33106]_  = A299 & A298;
  assign \new_[33107]_  = \new_[33106]_  & \new_[33103]_ ;
  assign \new_[33108]_  = \new_[33107]_  & \new_[33100]_ ;
  assign \new_[33112]_  = ~A166 & ~A167;
  assign \new_[33113]_  = A170 & \new_[33112]_ ;
  assign \new_[33117]_  = A201 & ~A200;
  assign \new_[33118]_  = A199 & \new_[33117]_ ;
  assign \new_[33119]_  = \new_[33118]_  & \new_[33113]_ ;
  assign \new_[33123]_  = ~A233 & A232;
  assign \new_[33124]_  = A202 & \new_[33123]_ ;
  assign \new_[33127]_  = A235 & A234;
  assign \new_[33130]_  = ~A299 & ~A298;
  assign \new_[33131]_  = \new_[33130]_  & \new_[33127]_ ;
  assign \new_[33132]_  = \new_[33131]_  & \new_[33124]_ ;
  assign \new_[33136]_  = ~A166 & ~A167;
  assign \new_[33137]_  = A170 & \new_[33136]_ ;
  assign \new_[33141]_  = A201 & ~A200;
  assign \new_[33142]_  = A199 & \new_[33141]_ ;
  assign \new_[33143]_  = \new_[33142]_  & \new_[33137]_ ;
  assign \new_[33147]_  = ~A233 & A232;
  assign \new_[33148]_  = A202 & \new_[33147]_ ;
  assign \new_[33151]_  = A235 & A234;
  assign \new_[33154]_  = A266 & ~A265;
  assign \new_[33155]_  = \new_[33154]_  & \new_[33151]_ ;
  assign \new_[33156]_  = \new_[33155]_  & \new_[33148]_ ;
  assign \new_[33160]_  = ~A166 & ~A167;
  assign \new_[33161]_  = A170 & \new_[33160]_ ;
  assign \new_[33165]_  = A201 & ~A200;
  assign \new_[33166]_  = A199 & \new_[33165]_ ;
  assign \new_[33167]_  = \new_[33166]_  & \new_[33161]_ ;
  assign \new_[33171]_  = ~A233 & A232;
  assign \new_[33172]_  = A202 & \new_[33171]_ ;
  assign \new_[33175]_  = A236 & A234;
  assign \new_[33178]_  = ~A300 & A298;
  assign \new_[33179]_  = \new_[33178]_  & \new_[33175]_ ;
  assign \new_[33180]_  = \new_[33179]_  & \new_[33172]_ ;
  assign \new_[33184]_  = ~A166 & ~A167;
  assign \new_[33185]_  = A170 & \new_[33184]_ ;
  assign \new_[33189]_  = A201 & ~A200;
  assign \new_[33190]_  = A199 & \new_[33189]_ ;
  assign \new_[33191]_  = \new_[33190]_  & \new_[33185]_ ;
  assign \new_[33195]_  = ~A233 & A232;
  assign \new_[33196]_  = A202 & \new_[33195]_ ;
  assign \new_[33199]_  = A236 & A234;
  assign \new_[33202]_  = A299 & A298;
  assign \new_[33203]_  = \new_[33202]_  & \new_[33199]_ ;
  assign \new_[33204]_  = \new_[33203]_  & \new_[33196]_ ;
  assign \new_[33208]_  = ~A166 & ~A167;
  assign \new_[33209]_  = A170 & \new_[33208]_ ;
  assign \new_[33213]_  = A201 & ~A200;
  assign \new_[33214]_  = A199 & \new_[33213]_ ;
  assign \new_[33215]_  = \new_[33214]_  & \new_[33209]_ ;
  assign \new_[33219]_  = ~A233 & A232;
  assign \new_[33220]_  = A202 & \new_[33219]_ ;
  assign \new_[33223]_  = A236 & A234;
  assign \new_[33226]_  = ~A299 & ~A298;
  assign \new_[33227]_  = \new_[33226]_  & \new_[33223]_ ;
  assign \new_[33228]_  = \new_[33227]_  & \new_[33220]_ ;
  assign \new_[33232]_  = ~A166 & ~A167;
  assign \new_[33233]_  = A170 & \new_[33232]_ ;
  assign \new_[33237]_  = A201 & ~A200;
  assign \new_[33238]_  = A199 & \new_[33237]_ ;
  assign \new_[33239]_  = \new_[33238]_  & \new_[33233]_ ;
  assign \new_[33243]_  = ~A233 & A232;
  assign \new_[33244]_  = A202 & \new_[33243]_ ;
  assign \new_[33247]_  = A236 & A234;
  assign \new_[33250]_  = A266 & ~A265;
  assign \new_[33251]_  = \new_[33250]_  & \new_[33247]_ ;
  assign \new_[33252]_  = \new_[33251]_  & \new_[33244]_ ;
  assign \new_[33256]_  = ~A166 & ~A167;
  assign \new_[33257]_  = A170 & \new_[33256]_ ;
  assign \new_[33261]_  = A201 & ~A200;
  assign \new_[33262]_  = A199 & \new_[33261]_ ;
  assign \new_[33263]_  = \new_[33262]_  & \new_[33257]_ ;
  assign \new_[33267]_  = ~A233 & ~A232;
  assign \new_[33268]_  = A202 & \new_[33267]_ ;
  assign \new_[33271]_  = A266 & A265;
  assign \new_[33274]_  = A299 & ~A298;
  assign \new_[33275]_  = \new_[33274]_  & \new_[33271]_ ;
  assign \new_[33276]_  = \new_[33275]_  & \new_[33268]_ ;
  assign \new_[33280]_  = ~A166 & ~A167;
  assign \new_[33281]_  = A170 & \new_[33280]_ ;
  assign \new_[33285]_  = A201 & ~A200;
  assign \new_[33286]_  = A199 & \new_[33285]_ ;
  assign \new_[33287]_  = \new_[33286]_  & \new_[33281]_ ;
  assign \new_[33291]_  = ~A233 & ~A232;
  assign \new_[33292]_  = A202 & \new_[33291]_ ;
  assign \new_[33295]_  = ~A267 & ~A266;
  assign \new_[33298]_  = A299 & ~A298;
  assign \new_[33299]_  = \new_[33298]_  & \new_[33295]_ ;
  assign \new_[33300]_  = \new_[33299]_  & \new_[33292]_ ;
  assign \new_[33304]_  = ~A166 & ~A167;
  assign \new_[33305]_  = A170 & \new_[33304]_ ;
  assign \new_[33309]_  = A201 & ~A200;
  assign \new_[33310]_  = A199 & \new_[33309]_ ;
  assign \new_[33311]_  = \new_[33310]_  & \new_[33305]_ ;
  assign \new_[33315]_  = ~A233 & ~A232;
  assign \new_[33316]_  = A202 & \new_[33315]_ ;
  assign \new_[33319]_  = ~A266 & ~A265;
  assign \new_[33322]_  = A299 & ~A298;
  assign \new_[33323]_  = \new_[33322]_  & \new_[33319]_ ;
  assign \new_[33324]_  = \new_[33323]_  & \new_[33316]_ ;
  assign \new_[33328]_  = ~A166 & ~A167;
  assign \new_[33329]_  = A170 & \new_[33328]_ ;
  assign \new_[33333]_  = A201 & ~A200;
  assign \new_[33334]_  = A199 & \new_[33333]_ ;
  assign \new_[33335]_  = \new_[33334]_  & \new_[33329]_ ;
  assign \new_[33339]_  = A233 & A232;
  assign \new_[33340]_  = A203 & \new_[33339]_ ;
  assign \new_[33343]_  = ~A267 & A265;
  assign \new_[33346]_  = A299 & ~A298;
  assign \new_[33347]_  = \new_[33346]_  & \new_[33343]_ ;
  assign \new_[33348]_  = \new_[33347]_  & \new_[33340]_ ;
  assign \new_[33352]_  = ~A166 & ~A167;
  assign \new_[33353]_  = A170 & \new_[33352]_ ;
  assign \new_[33357]_  = A201 & ~A200;
  assign \new_[33358]_  = A199 & \new_[33357]_ ;
  assign \new_[33359]_  = \new_[33358]_  & \new_[33353]_ ;
  assign \new_[33363]_  = A233 & A232;
  assign \new_[33364]_  = A203 & \new_[33363]_ ;
  assign \new_[33367]_  = A266 & A265;
  assign \new_[33370]_  = A299 & ~A298;
  assign \new_[33371]_  = \new_[33370]_  & \new_[33367]_ ;
  assign \new_[33372]_  = \new_[33371]_  & \new_[33364]_ ;
  assign \new_[33376]_  = ~A166 & ~A167;
  assign \new_[33377]_  = A170 & \new_[33376]_ ;
  assign \new_[33381]_  = A201 & ~A200;
  assign \new_[33382]_  = A199 & \new_[33381]_ ;
  assign \new_[33383]_  = \new_[33382]_  & \new_[33377]_ ;
  assign \new_[33387]_  = A233 & A232;
  assign \new_[33388]_  = A203 & \new_[33387]_ ;
  assign \new_[33391]_  = ~A266 & ~A265;
  assign \new_[33394]_  = A299 & ~A298;
  assign \new_[33395]_  = \new_[33394]_  & \new_[33391]_ ;
  assign \new_[33396]_  = \new_[33395]_  & \new_[33388]_ ;
  assign \new_[33400]_  = ~A166 & ~A167;
  assign \new_[33401]_  = A170 & \new_[33400]_ ;
  assign \new_[33405]_  = A201 & ~A200;
  assign \new_[33406]_  = A199 & \new_[33405]_ ;
  assign \new_[33407]_  = \new_[33406]_  & \new_[33401]_ ;
  assign \new_[33411]_  = A233 & ~A232;
  assign \new_[33412]_  = A203 & \new_[33411]_ ;
  assign \new_[33415]_  = ~A266 & A265;
  assign \new_[33418]_  = A268 & A267;
  assign \new_[33419]_  = \new_[33418]_  & \new_[33415]_ ;
  assign \new_[33420]_  = \new_[33419]_  & \new_[33412]_ ;
  assign \new_[33424]_  = ~A166 & ~A167;
  assign \new_[33425]_  = A170 & \new_[33424]_ ;
  assign \new_[33429]_  = A201 & ~A200;
  assign \new_[33430]_  = A199 & \new_[33429]_ ;
  assign \new_[33431]_  = \new_[33430]_  & \new_[33425]_ ;
  assign \new_[33435]_  = A233 & ~A232;
  assign \new_[33436]_  = A203 & \new_[33435]_ ;
  assign \new_[33439]_  = ~A266 & A265;
  assign \new_[33442]_  = A269 & A267;
  assign \new_[33443]_  = \new_[33442]_  & \new_[33439]_ ;
  assign \new_[33444]_  = \new_[33443]_  & \new_[33436]_ ;
  assign \new_[33448]_  = ~A166 & ~A167;
  assign \new_[33449]_  = A170 & \new_[33448]_ ;
  assign \new_[33453]_  = A201 & ~A200;
  assign \new_[33454]_  = A199 & \new_[33453]_ ;
  assign \new_[33455]_  = \new_[33454]_  & \new_[33449]_ ;
  assign \new_[33459]_  = ~A234 & ~A233;
  assign \new_[33460]_  = A203 & \new_[33459]_ ;
  assign \new_[33463]_  = A266 & A265;
  assign \new_[33466]_  = A299 & ~A298;
  assign \new_[33467]_  = \new_[33466]_  & \new_[33463]_ ;
  assign \new_[33468]_  = \new_[33467]_  & \new_[33460]_ ;
  assign \new_[33472]_  = ~A166 & ~A167;
  assign \new_[33473]_  = A170 & \new_[33472]_ ;
  assign \new_[33477]_  = A201 & ~A200;
  assign \new_[33478]_  = A199 & \new_[33477]_ ;
  assign \new_[33479]_  = \new_[33478]_  & \new_[33473]_ ;
  assign \new_[33483]_  = ~A234 & ~A233;
  assign \new_[33484]_  = A203 & \new_[33483]_ ;
  assign \new_[33487]_  = ~A267 & ~A266;
  assign \new_[33490]_  = A299 & ~A298;
  assign \new_[33491]_  = \new_[33490]_  & \new_[33487]_ ;
  assign \new_[33492]_  = \new_[33491]_  & \new_[33484]_ ;
  assign \new_[33496]_  = ~A166 & ~A167;
  assign \new_[33497]_  = A170 & \new_[33496]_ ;
  assign \new_[33501]_  = A201 & ~A200;
  assign \new_[33502]_  = A199 & \new_[33501]_ ;
  assign \new_[33503]_  = \new_[33502]_  & \new_[33497]_ ;
  assign \new_[33507]_  = ~A234 & ~A233;
  assign \new_[33508]_  = A203 & \new_[33507]_ ;
  assign \new_[33511]_  = ~A266 & ~A265;
  assign \new_[33514]_  = A299 & ~A298;
  assign \new_[33515]_  = \new_[33514]_  & \new_[33511]_ ;
  assign \new_[33516]_  = \new_[33515]_  & \new_[33508]_ ;
  assign \new_[33520]_  = ~A166 & ~A167;
  assign \new_[33521]_  = A170 & \new_[33520]_ ;
  assign \new_[33525]_  = A201 & ~A200;
  assign \new_[33526]_  = A199 & \new_[33525]_ ;
  assign \new_[33527]_  = \new_[33526]_  & \new_[33521]_ ;
  assign \new_[33531]_  = ~A233 & A232;
  assign \new_[33532]_  = A203 & \new_[33531]_ ;
  assign \new_[33535]_  = A235 & A234;
  assign \new_[33538]_  = ~A300 & A298;
  assign \new_[33539]_  = \new_[33538]_  & \new_[33535]_ ;
  assign \new_[33540]_  = \new_[33539]_  & \new_[33532]_ ;
  assign \new_[33544]_  = ~A166 & ~A167;
  assign \new_[33545]_  = A170 & \new_[33544]_ ;
  assign \new_[33549]_  = A201 & ~A200;
  assign \new_[33550]_  = A199 & \new_[33549]_ ;
  assign \new_[33551]_  = \new_[33550]_  & \new_[33545]_ ;
  assign \new_[33555]_  = ~A233 & A232;
  assign \new_[33556]_  = A203 & \new_[33555]_ ;
  assign \new_[33559]_  = A235 & A234;
  assign \new_[33562]_  = A299 & A298;
  assign \new_[33563]_  = \new_[33562]_  & \new_[33559]_ ;
  assign \new_[33564]_  = \new_[33563]_  & \new_[33556]_ ;
  assign \new_[33568]_  = ~A166 & ~A167;
  assign \new_[33569]_  = A170 & \new_[33568]_ ;
  assign \new_[33573]_  = A201 & ~A200;
  assign \new_[33574]_  = A199 & \new_[33573]_ ;
  assign \new_[33575]_  = \new_[33574]_  & \new_[33569]_ ;
  assign \new_[33579]_  = ~A233 & A232;
  assign \new_[33580]_  = A203 & \new_[33579]_ ;
  assign \new_[33583]_  = A235 & A234;
  assign \new_[33586]_  = ~A299 & ~A298;
  assign \new_[33587]_  = \new_[33586]_  & \new_[33583]_ ;
  assign \new_[33588]_  = \new_[33587]_  & \new_[33580]_ ;
  assign \new_[33592]_  = ~A166 & ~A167;
  assign \new_[33593]_  = A170 & \new_[33592]_ ;
  assign \new_[33597]_  = A201 & ~A200;
  assign \new_[33598]_  = A199 & \new_[33597]_ ;
  assign \new_[33599]_  = \new_[33598]_  & \new_[33593]_ ;
  assign \new_[33603]_  = ~A233 & A232;
  assign \new_[33604]_  = A203 & \new_[33603]_ ;
  assign \new_[33607]_  = A235 & A234;
  assign \new_[33610]_  = A266 & ~A265;
  assign \new_[33611]_  = \new_[33610]_  & \new_[33607]_ ;
  assign \new_[33612]_  = \new_[33611]_  & \new_[33604]_ ;
  assign \new_[33616]_  = ~A166 & ~A167;
  assign \new_[33617]_  = A170 & \new_[33616]_ ;
  assign \new_[33621]_  = A201 & ~A200;
  assign \new_[33622]_  = A199 & \new_[33621]_ ;
  assign \new_[33623]_  = \new_[33622]_  & \new_[33617]_ ;
  assign \new_[33627]_  = ~A233 & A232;
  assign \new_[33628]_  = A203 & \new_[33627]_ ;
  assign \new_[33631]_  = A236 & A234;
  assign \new_[33634]_  = ~A300 & A298;
  assign \new_[33635]_  = \new_[33634]_  & \new_[33631]_ ;
  assign \new_[33636]_  = \new_[33635]_  & \new_[33628]_ ;
  assign \new_[33640]_  = ~A166 & ~A167;
  assign \new_[33641]_  = A170 & \new_[33640]_ ;
  assign \new_[33645]_  = A201 & ~A200;
  assign \new_[33646]_  = A199 & \new_[33645]_ ;
  assign \new_[33647]_  = \new_[33646]_  & \new_[33641]_ ;
  assign \new_[33651]_  = ~A233 & A232;
  assign \new_[33652]_  = A203 & \new_[33651]_ ;
  assign \new_[33655]_  = A236 & A234;
  assign \new_[33658]_  = A299 & A298;
  assign \new_[33659]_  = \new_[33658]_  & \new_[33655]_ ;
  assign \new_[33660]_  = \new_[33659]_  & \new_[33652]_ ;
  assign \new_[33664]_  = ~A166 & ~A167;
  assign \new_[33665]_  = A170 & \new_[33664]_ ;
  assign \new_[33669]_  = A201 & ~A200;
  assign \new_[33670]_  = A199 & \new_[33669]_ ;
  assign \new_[33671]_  = \new_[33670]_  & \new_[33665]_ ;
  assign \new_[33675]_  = ~A233 & A232;
  assign \new_[33676]_  = A203 & \new_[33675]_ ;
  assign \new_[33679]_  = A236 & A234;
  assign \new_[33682]_  = ~A299 & ~A298;
  assign \new_[33683]_  = \new_[33682]_  & \new_[33679]_ ;
  assign \new_[33684]_  = \new_[33683]_  & \new_[33676]_ ;
  assign \new_[33688]_  = ~A166 & ~A167;
  assign \new_[33689]_  = A170 & \new_[33688]_ ;
  assign \new_[33693]_  = A201 & ~A200;
  assign \new_[33694]_  = A199 & \new_[33693]_ ;
  assign \new_[33695]_  = \new_[33694]_  & \new_[33689]_ ;
  assign \new_[33699]_  = ~A233 & A232;
  assign \new_[33700]_  = A203 & \new_[33699]_ ;
  assign \new_[33703]_  = A236 & A234;
  assign \new_[33706]_  = A266 & ~A265;
  assign \new_[33707]_  = \new_[33706]_  & \new_[33703]_ ;
  assign \new_[33708]_  = \new_[33707]_  & \new_[33700]_ ;
  assign \new_[33712]_  = ~A166 & ~A167;
  assign \new_[33713]_  = A170 & \new_[33712]_ ;
  assign \new_[33717]_  = A201 & ~A200;
  assign \new_[33718]_  = A199 & \new_[33717]_ ;
  assign \new_[33719]_  = \new_[33718]_  & \new_[33713]_ ;
  assign \new_[33723]_  = ~A233 & ~A232;
  assign \new_[33724]_  = A203 & \new_[33723]_ ;
  assign \new_[33727]_  = A266 & A265;
  assign \new_[33730]_  = A299 & ~A298;
  assign \new_[33731]_  = \new_[33730]_  & \new_[33727]_ ;
  assign \new_[33732]_  = \new_[33731]_  & \new_[33724]_ ;
  assign \new_[33736]_  = ~A166 & ~A167;
  assign \new_[33737]_  = A170 & \new_[33736]_ ;
  assign \new_[33741]_  = A201 & ~A200;
  assign \new_[33742]_  = A199 & \new_[33741]_ ;
  assign \new_[33743]_  = \new_[33742]_  & \new_[33737]_ ;
  assign \new_[33747]_  = ~A233 & ~A232;
  assign \new_[33748]_  = A203 & \new_[33747]_ ;
  assign \new_[33751]_  = ~A267 & ~A266;
  assign \new_[33754]_  = A299 & ~A298;
  assign \new_[33755]_  = \new_[33754]_  & \new_[33751]_ ;
  assign \new_[33756]_  = \new_[33755]_  & \new_[33748]_ ;
  assign \new_[33760]_  = ~A166 & ~A167;
  assign \new_[33761]_  = A170 & \new_[33760]_ ;
  assign \new_[33765]_  = A201 & ~A200;
  assign \new_[33766]_  = A199 & \new_[33765]_ ;
  assign \new_[33767]_  = \new_[33766]_  & \new_[33761]_ ;
  assign \new_[33771]_  = ~A233 & ~A232;
  assign \new_[33772]_  = A203 & \new_[33771]_ ;
  assign \new_[33775]_  = ~A266 & ~A265;
  assign \new_[33778]_  = A299 & ~A298;
  assign \new_[33779]_  = \new_[33778]_  & \new_[33775]_ ;
  assign \new_[33780]_  = \new_[33779]_  & \new_[33772]_ ;
  assign \new_[33784]_  = A167 & ~A168;
  assign \new_[33785]_  = A170 & \new_[33784]_ ;
  assign \new_[33789]_  = A200 & ~A199;
  assign \new_[33790]_  = A166 & \new_[33789]_ ;
  assign \new_[33791]_  = \new_[33790]_  & \new_[33785]_ ;
  assign \new_[33795]_  = A265 & A233;
  assign \new_[33796]_  = A232 & \new_[33795]_ ;
  assign \new_[33799]_  = ~A269 & ~A268;
  assign \new_[33802]_  = A299 & ~A298;
  assign \new_[33803]_  = \new_[33802]_  & \new_[33799]_ ;
  assign \new_[33804]_  = \new_[33803]_  & \new_[33796]_ ;
  assign \new_[33808]_  = A167 & ~A168;
  assign \new_[33809]_  = A170 & \new_[33808]_ ;
  assign \new_[33813]_  = A200 & ~A199;
  assign \new_[33814]_  = A166 & \new_[33813]_ ;
  assign \new_[33815]_  = \new_[33814]_  & \new_[33809]_ ;
  assign \new_[33819]_  = ~A236 & ~A235;
  assign \new_[33820]_  = ~A233 & \new_[33819]_ ;
  assign \new_[33823]_  = A266 & A265;
  assign \new_[33826]_  = A299 & ~A298;
  assign \new_[33827]_  = \new_[33826]_  & \new_[33823]_ ;
  assign \new_[33828]_  = \new_[33827]_  & \new_[33820]_ ;
  assign \new_[33832]_  = A167 & ~A168;
  assign \new_[33833]_  = A170 & \new_[33832]_ ;
  assign \new_[33837]_  = A200 & ~A199;
  assign \new_[33838]_  = A166 & \new_[33837]_ ;
  assign \new_[33839]_  = \new_[33838]_  & \new_[33833]_ ;
  assign \new_[33843]_  = ~A236 & ~A235;
  assign \new_[33844]_  = ~A233 & \new_[33843]_ ;
  assign \new_[33847]_  = ~A267 & ~A266;
  assign \new_[33850]_  = A299 & ~A298;
  assign \new_[33851]_  = \new_[33850]_  & \new_[33847]_ ;
  assign \new_[33852]_  = \new_[33851]_  & \new_[33844]_ ;
  assign \new_[33856]_  = A167 & ~A168;
  assign \new_[33857]_  = A170 & \new_[33856]_ ;
  assign \new_[33861]_  = A200 & ~A199;
  assign \new_[33862]_  = A166 & \new_[33861]_ ;
  assign \new_[33863]_  = \new_[33862]_  & \new_[33857]_ ;
  assign \new_[33867]_  = ~A236 & ~A235;
  assign \new_[33868]_  = ~A233 & \new_[33867]_ ;
  assign \new_[33871]_  = ~A266 & ~A265;
  assign \new_[33874]_  = A299 & ~A298;
  assign \new_[33875]_  = \new_[33874]_  & \new_[33871]_ ;
  assign \new_[33876]_  = \new_[33875]_  & \new_[33868]_ ;
  assign \new_[33880]_  = A167 & ~A168;
  assign \new_[33881]_  = A170 & \new_[33880]_ ;
  assign \new_[33885]_  = A200 & ~A199;
  assign \new_[33886]_  = A166 & \new_[33885]_ ;
  assign \new_[33887]_  = \new_[33886]_  & \new_[33881]_ ;
  assign \new_[33891]_  = ~A266 & ~A234;
  assign \new_[33892]_  = ~A233 & \new_[33891]_ ;
  assign \new_[33895]_  = ~A269 & ~A268;
  assign \new_[33898]_  = A299 & ~A298;
  assign \new_[33899]_  = \new_[33898]_  & \new_[33895]_ ;
  assign \new_[33900]_  = \new_[33899]_  & \new_[33892]_ ;
  assign \new_[33904]_  = A167 & ~A168;
  assign \new_[33905]_  = A170 & \new_[33904]_ ;
  assign \new_[33909]_  = A200 & ~A199;
  assign \new_[33910]_  = A166 & \new_[33909]_ ;
  assign \new_[33911]_  = \new_[33910]_  & \new_[33905]_ ;
  assign \new_[33915]_  = A234 & ~A233;
  assign \new_[33916]_  = A232 & \new_[33915]_ ;
  assign \new_[33919]_  = A298 & A235;
  assign \new_[33922]_  = ~A302 & ~A301;
  assign \new_[33923]_  = \new_[33922]_  & \new_[33919]_ ;
  assign \new_[33924]_  = \new_[33923]_  & \new_[33916]_ ;
  assign \new_[33928]_  = A167 & ~A168;
  assign \new_[33929]_  = A170 & \new_[33928]_ ;
  assign \new_[33933]_  = A200 & ~A199;
  assign \new_[33934]_  = A166 & \new_[33933]_ ;
  assign \new_[33935]_  = \new_[33934]_  & \new_[33929]_ ;
  assign \new_[33939]_  = A234 & ~A233;
  assign \new_[33940]_  = A232 & \new_[33939]_ ;
  assign \new_[33943]_  = A298 & A236;
  assign \new_[33946]_  = ~A302 & ~A301;
  assign \new_[33947]_  = \new_[33946]_  & \new_[33943]_ ;
  assign \new_[33948]_  = \new_[33947]_  & \new_[33940]_ ;
  assign \new_[33952]_  = A167 & ~A168;
  assign \new_[33953]_  = A170 & \new_[33952]_ ;
  assign \new_[33957]_  = A200 & ~A199;
  assign \new_[33958]_  = A166 & \new_[33957]_ ;
  assign \new_[33959]_  = \new_[33958]_  & \new_[33953]_ ;
  assign \new_[33963]_  = ~A266 & ~A233;
  assign \new_[33964]_  = ~A232 & \new_[33963]_ ;
  assign \new_[33967]_  = ~A269 & ~A268;
  assign \new_[33970]_  = A299 & ~A298;
  assign \new_[33971]_  = \new_[33970]_  & \new_[33967]_ ;
  assign \new_[33972]_  = \new_[33971]_  & \new_[33964]_ ;
  assign \new_[33976]_  = A167 & ~A168;
  assign \new_[33977]_  = ~A170 & \new_[33976]_ ;
  assign \new_[33981]_  = A200 & ~A199;
  assign \new_[33982]_  = ~A166 & \new_[33981]_ ;
  assign \new_[33983]_  = \new_[33982]_  & \new_[33977]_ ;
  assign \new_[33987]_  = A265 & A233;
  assign \new_[33988]_  = A232 & \new_[33987]_ ;
  assign \new_[33991]_  = ~A269 & ~A268;
  assign \new_[33994]_  = A299 & ~A298;
  assign \new_[33995]_  = \new_[33994]_  & \new_[33991]_ ;
  assign \new_[33996]_  = \new_[33995]_  & \new_[33988]_ ;
  assign \new_[34000]_  = A167 & ~A168;
  assign \new_[34001]_  = ~A170 & \new_[34000]_ ;
  assign \new_[34005]_  = A200 & ~A199;
  assign \new_[34006]_  = ~A166 & \new_[34005]_ ;
  assign \new_[34007]_  = \new_[34006]_  & \new_[34001]_ ;
  assign \new_[34011]_  = ~A236 & ~A235;
  assign \new_[34012]_  = ~A233 & \new_[34011]_ ;
  assign \new_[34015]_  = A266 & A265;
  assign \new_[34018]_  = A299 & ~A298;
  assign \new_[34019]_  = \new_[34018]_  & \new_[34015]_ ;
  assign \new_[34020]_  = \new_[34019]_  & \new_[34012]_ ;
  assign \new_[34024]_  = A167 & ~A168;
  assign \new_[34025]_  = ~A170 & \new_[34024]_ ;
  assign \new_[34029]_  = A200 & ~A199;
  assign \new_[34030]_  = ~A166 & \new_[34029]_ ;
  assign \new_[34031]_  = \new_[34030]_  & \new_[34025]_ ;
  assign \new_[34035]_  = ~A236 & ~A235;
  assign \new_[34036]_  = ~A233 & \new_[34035]_ ;
  assign \new_[34039]_  = ~A267 & ~A266;
  assign \new_[34042]_  = A299 & ~A298;
  assign \new_[34043]_  = \new_[34042]_  & \new_[34039]_ ;
  assign \new_[34044]_  = \new_[34043]_  & \new_[34036]_ ;
  assign \new_[34048]_  = A167 & ~A168;
  assign \new_[34049]_  = ~A170 & \new_[34048]_ ;
  assign \new_[34053]_  = A200 & ~A199;
  assign \new_[34054]_  = ~A166 & \new_[34053]_ ;
  assign \new_[34055]_  = \new_[34054]_  & \new_[34049]_ ;
  assign \new_[34059]_  = ~A236 & ~A235;
  assign \new_[34060]_  = ~A233 & \new_[34059]_ ;
  assign \new_[34063]_  = ~A266 & ~A265;
  assign \new_[34066]_  = A299 & ~A298;
  assign \new_[34067]_  = \new_[34066]_  & \new_[34063]_ ;
  assign \new_[34068]_  = \new_[34067]_  & \new_[34060]_ ;
  assign \new_[34072]_  = A167 & ~A168;
  assign \new_[34073]_  = ~A170 & \new_[34072]_ ;
  assign \new_[34077]_  = A200 & ~A199;
  assign \new_[34078]_  = ~A166 & \new_[34077]_ ;
  assign \new_[34079]_  = \new_[34078]_  & \new_[34073]_ ;
  assign \new_[34083]_  = ~A266 & ~A234;
  assign \new_[34084]_  = ~A233 & \new_[34083]_ ;
  assign \new_[34087]_  = ~A269 & ~A268;
  assign \new_[34090]_  = A299 & ~A298;
  assign \new_[34091]_  = \new_[34090]_  & \new_[34087]_ ;
  assign \new_[34092]_  = \new_[34091]_  & \new_[34084]_ ;
  assign \new_[34096]_  = A167 & ~A168;
  assign \new_[34097]_  = ~A170 & \new_[34096]_ ;
  assign \new_[34101]_  = A200 & ~A199;
  assign \new_[34102]_  = ~A166 & \new_[34101]_ ;
  assign \new_[34103]_  = \new_[34102]_  & \new_[34097]_ ;
  assign \new_[34107]_  = A234 & ~A233;
  assign \new_[34108]_  = A232 & \new_[34107]_ ;
  assign \new_[34111]_  = A298 & A235;
  assign \new_[34114]_  = ~A302 & ~A301;
  assign \new_[34115]_  = \new_[34114]_  & \new_[34111]_ ;
  assign \new_[34116]_  = \new_[34115]_  & \new_[34108]_ ;
  assign \new_[34120]_  = A167 & ~A168;
  assign \new_[34121]_  = ~A170 & \new_[34120]_ ;
  assign \new_[34125]_  = A200 & ~A199;
  assign \new_[34126]_  = ~A166 & \new_[34125]_ ;
  assign \new_[34127]_  = \new_[34126]_  & \new_[34121]_ ;
  assign \new_[34131]_  = A234 & ~A233;
  assign \new_[34132]_  = A232 & \new_[34131]_ ;
  assign \new_[34135]_  = A298 & A236;
  assign \new_[34138]_  = ~A302 & ~A301;
  assign \new_[34139]_  = \new_[34138]_  & \new_[34135]_ ;
  assign \new_[34140]_  = \new_[34139]_  & \new_[34132]_ ;
  assign \new_[34144]_  = A167 & ~A168;
  assign \new_[34145]_  = ~A170 & \new_[34144]_ ;
  assign \new_[34149]_  = A200 & ~A199;
  assign \new_[34150]_  = ~A166 & \new_[34149]_ ;
  assign \new_[34151]_  = \new_[34150]_  & \new_[34145]_ ;
  assign \new_[34155]_  = ~A266 & ~A233;
  assign \new_[34156]_  = ~A232 & \new_[34155]_ ;
  assign \new_[34159]_  = ~A269 & ~A268;
  assign \new_[34162]_  = A299 & ~A298;
  assign \new_[34163]_  = \new_[34162]_  & \new_[34159]_ ;
  assign \new_[34164]_  = \new_[34163]_  & \new_[34156]_ ;
  assign \new_[34168]_  = ~A167 & ~A168;
  assign \new_[34169]_  = ~A170 & \new_[34168]_ ;
  assign \new_[34173]_  = A200 & ~A199;
  assign \new_[34174]_  = A166 & \new_[34173]_ ;
  assign \new_[34175]_  = \new_[34174]_  & \new_[34169]_ ;
  assign \new_[34179]_  = A265 & A233;
  assign \new_[34180]_  = A232 & \new_[34179]_ ;
  assign \new_[34183]_  = ~A269 & ~A268;
  assign \new_[34186]_  = A299 & ~A298;
  assign \new_[34187]_  = \new_[34186]_  & \new_[34183]_ ;
  assign \new_[34188]_  = \new_[34187]_  & \new_[34180]_ ;
  assign \new_[34192]_  = ~A167 & ~A168;
  assign \new_[34193]_  = ~A170 & \new_[34192]_ ;
  assign \new_[34197]_  = A200 & ~A199;
  assign \new_[34198]_  = A166 & \new_[34197]_ ;
  assign \new_[34199]_  = \new_[34198]_  & \new_[34193]_ ;
  assign \new_[34203]_  = ~A236 & ~A235;
  assign \new_[34204]_  = ~A233 & \new_[34203]_ ;
  assign \new_[34207]_  = A266 & A265;
  assign \new_[34210]_  = A299 & ~A298;
  assign \new_[34211]_  = \new_[34210]_  & \new_[34207]_ ;
  assign \new_[34212]_  = \new_[34211]_  & \new_[34204]_ ;
  assign \new_[34216]_  = ~A167 & ~A168;
  assign \new_[34217]_  = ~A170 & \new_[34216]_ ;
  assign \new_[34221]_  = A200 & ~A199;
  assign \new_[34222]_  = A166 & \new_[34221]_ ;
  assign \new_[34223]_  = \new_[34222]_  & \new_[34217]_ ;
  assign \new_[34227]_  = ~A236 & ~A235;
  assign \new_[34228]_  = ~A233 & \new_[34227]_ ;
  assign \new_[34231]_  = ~A267 & ~A266;
  assign \new_[34234]_  = A299 & ~A298;
  assign \new_[34235]_  = \new_[34234]_  & \new_[34231]_ ;
  assign \new_[34236]_  = \new_[34235]_  & \new_[34228]_ ;
  assign \new_[34240]_  = ~A167 & ~A168;
  assign \new_[34241]_  = ~A170 & \new_[34240]_ ;
  assign \new_[34245]_  = A200 & ~A199;
  assign \new_[34246]_  = A166 & \new_[34245]_ ;
  assign \new_[34247]_  = \new_[34246]_  & \new_[34241]_ ;
  assign \new_[34251]_  = ~A236 & ~A235;
  assign \new_[34252]_  = ~A233 & \new_[34251]_ ;
  assign \new_[34255]_  = ~A266 & ~A265;
  assign \new_[34258]_  = A299 & ~A298;
  assign \new_[34259]_  = \new_[34258]_  & \new_[34255]_ ;
  assign \new_[34260]_  = \new_[34259]_  & \new_[34252]_ ;
  assign \new_[34264]_  = ~A167 & ~A168;
  assign \new_[34265]_  = ~A170 & \new_[34264]_ ;
  assign \new_[34269]_  = A200 & ~A199;
  assign \new_[34270]_  = A166 & \new_[34269]_ ;
  assign \new_[34271]_  = \new_[34270]_  & \new_[34265]_ ;
  assign \new_[34275]_  = ~A266 & ~A234;
  assign \new_[34276]_  = ~A233 & \new_[34275]_ ;
  assign \new_[34279]_  = ~A269 & ~A268;
  assign \new_[34282]_  = A299 & ~A298;
  assign \new_[34283]_  = \new_[34282]_  & \new_[34279]_ ;
  assign \new_[34284]_  = \new_[34283]_  & \new_[34276]_ ;
  assign \new_[34288]_  = ~A167 & ~A168;
  assign \new_[34289]_  = ~A170 & \new_[34288]_ ;
  assign \new_[34293]_  = A200 & ~A199;
  assign \new_[34294]_  = A166 & \new_[34293]_ ;
  assign \new_[34295]_  = \new_[34294]_  & \new_[34289]_ ;
  assign \new_[34299]_  = A234 & ~A233;
  assign \new_[34300]_  = A232 & \new_[34299]_ ;
  assign \new_[34303]_  = A298 & A235;
  assign \new_[34306]_  = ~A302 & ~A301;
  assign \new_[34307]_  = \new_[34306]_  & \new_[34303]_ ;
  assign \new_[34308]_  = \new_[34307]_  & \new_[34300]_ ;
  assign \new_[34312]_  = ~A167 & ~A168;
  assign \new_[34313]_  = ~A170 & \new_[34312]_ ;
  assign \new_[34317]_  = A200 & ~A199;
  assign \new_[34318]_  = A166 & \new_[34317]_ ;
  assign \new_[34319]_  = \new_[34318]_  & \new_[34313]_ ;
  assign \new_[34323]_  = A234 & ~A233;
  assign \new_[34324]_  = A232 & \new_[34323]_ ;
  assign \new_[34327]_  = A298 & A236;
  assign \new_[34330]_  = ~A302 & ~A301;
  assign \new_[34331]_  = \new_[34330]_  & \new_[34327]_ ;
  assign \new_[34332]_  = \new_[34331]_  & \new_[34324]_ ;
  assign \new_[34336]_  = ~A167 & ~A168;
  assign \new_[34337]_  = ~A170 & \new_[34336]_ ;
  assign \new_[34341]_  = A200 & ~A199;
  assign \new_[34342]_  = A166 & \new_[34341]_ ;
  assign \new_[34343]_  = \new_[34342]_  & \new_[34337]_ ;
  assign \new_[34347]_  = ~A266 & ~A233;
  assign \new_[34348]_  = ~A232 & \new_[34347]_ ;
  assign \new_[34351]_  = ~A269 & ~A268;
  assign \new_[34354]_  = A299 & ~A298;
  assign \new_[34355]_  = \new_[34354]_  & \new_[34351]_ ;
  assign \new_[34356]_  = \new_[34355]_  & \new_[34348]_ ;
  assign \new_[34360]_  = A167 & ~A168;
  assign \new_[34361]_  = A169 & \new_[34360]_ ;
  assign \new_[34365]_  = A200 & ~A199;
  assign \new_[34366]_  = ~A166 & \new_[34365]_ ;
  assign \new_[34367]_  = \new_[34366]_  & \new_[34361]_ ;
  assign \new_[34371]_  = A265 & A233;
  assign \new_[34372]_  = A232 & \new_[34371]_ ;
  assign \new_[34375]_  = ~A269 & ~A268;
  assign \new_[34378]_  = A299 & ~A298;
  assign \new_[34379]_  = \new_[34378]_  & \new_[34375]_ ;
  assign \new_[34380]_  = \new_[34379]_  & \new_[34372]_ ;
  assign \new_[34384]_  = A167 & ~A168;
  assign \new_[34385]_  = A169 & \new_[34384]_ ;
  assign \new_[34389]_  = A200 & ~A199;
  assign \new_[34390]_  = ~A166 & \new_[34389]_ ;
  assign \new_[34391]_  = \new_[34390]_  & \new_[34385]_ ;
  assign \new_[34395]_  = ~A236 & ~A235;
  assign \new_[34396]_  = ~A233 & \new_[34395]_ ;
  assign \new_[34399]_  = A266 & A265;
  assign \new_[34402]_  = A299 & ~A298;
  assign \new_[34403]_  = \new_[34402]_  & \new_[34399]_ ;
  assign \new_[34404]_  = \new_[34403]_  & \new_[34396]_ ;
  assign \new_[34408]_  = A167 & ~A168;
  assign \new_[34409]_  = A169 & \new_[34408]_ ;
  assign \new_[34413]_  = A200 & ~A199;
  assign \new_[34414]_  = ~A166 & \new_[34413]_ ;
  assign \new_[34415]_  = \new_[34414]_  & \new_[34409]_ ;
  assign \new_[34419]_  = ~A236 & ~A235;
  assign \new_[34420]_  = ~A233 & \new_[34419]_ ;
  assign \new_[34423]_  = ~A267 & ~A266;
  assign \new_[34426]_  = A299 & ~A298;
  assign \new_[34427]_  = \new_[34426]_  & \new_[34423]_ ;
  assign \new_[34428]_  = \new_[34427]_  & \new_[34420]_ ;
  assign \new_[34432]_  = A167 & ~A168;
  assign \new_[34433]_  = A169 & \new_[34432]_ ;
  assign \new_[34437]_  = A200 & ~A199;
  assign \new_[34438]_  = ~A166 & \new_[34437]_ ;
  assign \new_[34439]_  = \new_[34438]_  & \new_[34433]_ ;
  assign \new_[34443]_  = ~A236 & ~A235;
  assign \new_[34444]_  = ~A233 & \new_[34443]_ ;
  assign \new_[34447]_  = ~A266 & ~A265;
  assign \new_[34450]_  = A299 & ~A298;
  assign \new_[34451]_  = \new_[34450]_  & \new_[34447]_ ;
  assign \new_[34452]_  = \new_[34451]_  & \new_[34444]_ ;
  assign \new_[34456]_  = A167 & ~A168;
  assign \new_[34457]_  = A169 & \new_[34456]_ ;
  assign \new_[34461]_  = A200 & ~A199;
  assign \new_[34462]_  = ~A166 & \new_[34461]_ ;
  assign \new_[34463]_  = \new_[34462]_  & \new_[34457]_ ;
  assign \new_[34467]_  = ~A266 & ~A234;
  assign \new_[34468]_  = ~A233 & \new_[34467]_ ;
  assign \new_[34471]_  = ~A269 & ~A268;
  assign \new_[34474]_  = A299 & ~A298;
  assign \new_[34475]_  = \new_[34474]_  & \new_[34471]_ ;
  assign \new_[34476]_  = \new_[34475]_  & \new_[34468]_ ;
  assign \new_[34480]_  = A167 & ~A168;
  assign \new_[34481]_  = A169 & \new_[34480]_ ;
  assign \new_[34485]_  = A200 & ~A199;
  assign \new_[34486]_  = ~A166 & \new_[34485]_ ;
  assign \new_[34487]_  = \new_[34486]_  & \new_[34481]_ ;
  assign \new_[34491]_  = A234 & ~A233;
  assign \new_[34492]_  = A232 & \new_[34491]_ ;
  assign \new_[34495]_  = A298 & A235;
  assign \new_[34498]_  = ~A302 & ~A301;
  assign \new_[34499]_  = \new_[34498]_  & \new_[34495]_ ;
  assign \new_[34500]_  = \new_[34499]_  & \new_[34492]_ ;
  assign \new_[34504]_  = A167 & ~A168;
  assign \new_[34505]_  = A169 & \new_[34504]_ ;
  assign \new_[34509]_  = A200 & ~A199;
  assign \new_[34510]_  = ~A166 & \new_[34509]_ ;
  assign \new_[34511]_  = \new_[34510]_  & \new_[34505]_ ;
  assign \new_[34515]_  = A234 & ~A233;
  assign \new_[34516]_  = A232 & \new_[34515]_ ;
  assign \new_[34519]_  = A298 & A236;
  assign \new_[34522]_  = ~A302 & ~A301;
  assign \new_[34523]_  = \new_[34522]_  & \new_[34519]_ ;
  assign \new_[34524]_  = \new_[34523]_  & \new_[34516]_ ;
  assign \new_[34528]_  = A167 & ~A168;
  assign \new_[34529]_  = A169 & \new_[34528]_ ;
  assign \new_[34533]_  = A200 & ~A199;
  assign \new_[34534]_  = ~A166 & \new_[34533]_ ;
  assign \new_[34535]_  = \new_[34534]_  & \new_[34529]_ ;
  assign \new_[34539]_  = ~A266 & ~A233;
  assign \new_[34540]_  = ~A232 & \new_[34539]_ ;
  assign \new_[34543]_  = ~A269 & ~A268;
  assign \new_[34546]_  = A299 & ~A298;
  assign \new_[34547]_  = \new_[34546]_  & \new_[34543]_ ;
  assign \new_[34548]_  = \new_[34547]_  & \new_[34540]_ ;
  assign \new_[34552]_  = A167 & ~A168;
  assign \new_[34553]_  = A169 & \new_[34552]_ ;
  assign \new_[34557]_  = ~A200 & A199;
  assign \new_[34558]_  = ~A166 & \new_[34557]_ ;
  assign \new_[34559]_  = \new_[34558]_  & \new_[34553]_ ;
  assign \new_[34563]_  = ~A232 & A202;
  assign \new_[34564]_  = A201 & \new_[34563]_ ;
  assign \new_[34567]_  = ~A299 & A233;
  assign \new_[34570]_  = ~A302 & ~A301;
  assign \new_[34571]_  = \new_[34570]_  & \new_[34567]_ ;
  assign \new_[34572]_  = \new_[34571]_  & \new_[34564]_ ;
  assign \new_[34576]_  = A167 & ~A168;
  assign \new_[34577]_  = A169 & \new_[34576]_ ;
  assign \new_[34581]_  = ~A200 & A199;
  assign \new_[34582]_  = ~A166 & \new_[34581]_ ;
  assign \new_[34583]_  = \new_[34582]_  & \new_[34577]_ ;
  assign \new_[34587]_  = ~A232 & A203;
  assign \new_[34588]_  = A201 & \new_[34587]_ ;
  assign \new_[34591]_  = ~A299 & A233;
  assign \new_[34594]_  = ~A302 & ~A301;
  assign \new_[34595]_  = \new_[34594]_  & \new_[34591]_ ;
  assign \new_[34596]_  = \new_[34595]_  & \new_[34588]_ ;
  assign \new_[34600]_  = ~A167 & ~A168;
  assign \new_[34601]_  = A169 & \new_[34600]_ ;
  assign \new_[34605]_  = A200 & ~A199;
  assign \new_[34606]_  = A166 & \new_[34605]_ ;
  assign \new_[34607]_  = \new_[34606]_  & \new_[34601]_ ;
  assign \new_[34611]_  = A265 & A233;
  assign \new_[34612]_  = A232 & \new_[34611]_ ;
  assign \new_[34615]_  = ~A269 & ~A268;
  assign \new_[34618]_  = A299 & ~A298;
  assign \new_[34619]_  = \new_[34618]_  & \new_[34615]_ ;
  assign \new_[34620]_  = \new_[34619]_  & \new_[34612]_ ;
  assign \new_[34624]_  = ~A167 & ~A168;
  assign \new_[34625]_  = A169 & \new_[34624]_ ;
  assign \new_[34629]_  = A200 & ~A199;
  assign \new_[34630]_  = A166 & \new_[34629]_ ;
  assign \new_[34631]_  = \new_[34630]_  & \new_[34625]_ ;
  assign \new_[34635]_  = ~A236 & ~A235;
  assign \new_[34636]_  = ~A233 & \new_[34635]_ ;
  assign \new_[34639]_  = A266 & A265;
  assign \new_[34642]_  = A299 & ~A298;
  assign \new_[34643]_  = \new_[34642]_  & \new_[34639]_ ;
  assign \new_[34644]_  = \new_[34643]_  & \new_[34636]_ ;
  assign \new_[34648]_  = ~A167 & ~A168;
  assign \new_[34649]_  = A169 & \new_[34648]_ ;
  assign \new_[34653]_  = A200 & ~A199;
  assign \new_[34654]_  = A166 & \new_[34653]_ ;
  assign \new_[34655]_  = \new_[34654]_  & \new_[34649]_ ;
  assign \new_[34659]_  = ~A236 & ~A235;
  assign \new_[34660]_  = ~A233 & \new_[34659]_ ;
  assign \new_[34663]_  = ~A267 & ~A266;
  assign \new_[34666]_  = A299 & ~A298;
  assign \new_[34667]_  = \new_[34666]_  & \new_[34663]_ ;
  assign \new_[34668]_  = \new_[34667]_  & \new_[34660]_ ;
  assign \new_[34672]_  = ~A167 & ~A168;
  assign \new_[34673]_  = A169 & \new_[34672]_ ;
  assign \new_[34677]_  = A200 & ~A199;
  assign \new_[34678]_  = A166 & \new_[34677]_ ;
  assign \new_[34679]_  = \new_[34678]_  & \new_[34673]_ ;
  assign \new_[34683]_  = ~A236 & ~A235;
  assign \new_[34684]_  = ~A233 & \new_[34683]_ ;
  assign \new_[34687]_  = ~A266 & ~A265;
  assign \new_[34690]_  = A299 & ~A298;
  assign \new_[34691]_  = \new_[34690]_  & \new_[34687]_ ;
  assign \new_[34692]_  = \new_[34691]_  & \new_[34684]_ ;
  assign \new_[34696]_  = ~A167 & ~A168;
  assign \new_[34697]_  = A169 & \new_[34696]_ ;
  assign \new_[34701]_  = A200 & ~A199;
  assign \new_[34702]_  = A166 & \new_[34701]_ ;
  assign \new_[34703]_  = \new_[34702]_  & \new_[34697]_ ;
  assign \new_[34707]_  = ~A266 & ~A234;
  assign \new_[34708]_  = ~A233 & \new_[34707]_ ;
  assign \new_[34711]_  = ~A269 & ~A268;
  assign \new_[34714]_  = A299 & ~A298;
  assign \new_[34715]_  = \new_[34714]_  & \new_[34711]_ ;
  assign \new_[34716]_  = \new_[34715]_  & \new_[34708]_ ;
  assign \new_[34720]_  = ~A167 & ~A168;
  assign \new_[34721]_  = A169 & \new_[34720]_ ;
  assign \new_[34725]_  = A200 & ~A199;
  assign \new_[34726]_  = A166 & \new_[34725]_ ;
  assign \new_[34727]_  = \new_[34726]_  & \new_[34721]_ ;
  assign \new_[34731]_  = A234 & ~A233;
  assign \new_[34732]_  = A232 & \new_[34731]_ ;
  assign \new_[34735]_  = A298 & A235;
  assign \new_[34738]_  = ~A302 & ~A301;
  assign \new_[34739]_  = \new_[34738]_  & \new_[34735]_ ;
  assign \new_[34740]_  = \new_[34739]_  & \new_[34732]_ ;
  assign \new_[34744]_  = ~A167 & ~A168;
  assign \new_[34745]_  = A169 & \new_[34744]_ ;
  assign \new_[34749]_  = A200 & ~A199;
  assign \new_[34750]_  = A166 & \new_[34749]_ ;
  assign \new_[34751]_  = \new_[34750]_  & \new_[34745]_ ;
  assign \new_[34755]_  = A234 & ~A233;
  assign \new_[34756]_  = A232 & \new_[34755]_ ;
  assign \new_[34759]_  = A298 & A236;
  assign \new_[34762]_  = ~A302 & ~A301;
  assign \new_[34763]_  = \new_[34762]_  & \new_[34759]_ ;
  assign \new_[34764]_  = \new_[34763]_  & \new_[34756]_ ;
  assign \new_[34768]_  = ~A167 & ~A168;
  assign \new_[34769]_  = A169 & \new_[34768]_ ;
  assign \new_[34773]_  = A200 & ~A199;
  assign \new_[34774]_  = A166 & \new_[34773]_ ;
  assign \new_[34775]_  = \new_[34774]_  & \new_[34769]_ ;
  assign \new_[34779]_  = ~A266 & ~A233;
  assign \new_[34780]_  = ~A232 & \new_[34779]_ ;
  assign \new_[34783]_  = ~A269 & ~A268;
  assign \new_[34786]_  = A299 & ~A298;
  assign \new_[34787]_  = \new_[34786]_  & \new_[34783]_ ;
  assign \new_[34788]_  = \new_[34787]_  & \new_[34780]_ ;
  assign \new_[34792]_  = ~A167 & ~A168;
  assign \new_[34793]_  = A169 & \new_[34792]_ ;
  assign \new_[34797]_  = ~A200 & A199;
  assign \new_[34798]_  = A166 & \new_[34797]_ ;
  assign \new_[34799]_  = \new_[34798]_  & \new_[34793]_ ;
  assign \new_[34803]_  = ~A232 & A202;
  assign \new_[34804]_  = A201 & \new_[34803]_ ;
  assign \new_[34807]_  = ~A299 & A233;
  assign \new_[34810]_  = ~A302 & ~A301;
  assign \new_[34811]_  = \new_[34810]_  & \new_[34807]_ ;
  assign \new_[34812]_  = \new_[34811]_  & \new_[34804]_ ;
  assign \new_[34816]_  = ~A167 & ~A168;
  assign \new_[34817]_  = A169 & \new_[34816]_ ;
  assign \new_[34821]_  = ~A200 & A199;
  assign \new_[34822]_  = A166 & \new_[34821]_ ;
  assign \new_[34823]_  = \new_[34822]_  & \new_[34817]_ ;
  assign \new_[34827]_  = ~A232 & A203;
  assign \new_[34828]_  = A201 & \new_[34827]_ ;
  assign \new_[34831]_  = ~A299 & A233;
  assign \new_[34834]_  = ~A302 & ~A301;
  assign \new_[34835]_  = \new_[34834]_  & \new_[34831]_ ;
  assign \new_[34836]_  = \new_[34835]_  & \new_[34828]_ ;
  assign \new_[34840]_  = ~A168 & A169;
  assign \new_[34841]_  = A170 & \new_[34840]_ ;
  assign \new_[34845]_  = A201 & ~A200;
  assign \new_[34846]_  = A199 & \new_[34845]_ ;
  assign \new_[34847]_  = \new_[34846]_  & \new_[34841]_ ;
  assign \new_[34851]_  = A233 & A232;
  assign \new_[34852]_  = A202 & \new_[34851]_ ;
  assign \new_[34855]_  = ~A267 & A265;
  assign \new_[34858]_  = A299 & ~A298;
  assign \new_[34859]_  = \new_[34858]_  & \new_[34855]_ ;
  assign \new_[34860]_  = \new_[34859]_  & \new_[34852]_ ;
  assign \new_[34864]_  = ~A168 & A169;
  assign \new_[34865]_  = A170 & \new_[34864]_ ;
  assign \new_[34869]_  = A201 & ~A200;
  assign \new_[34870]_  = A199 & \new_[34869]_ ;
  assign \new_[34871]_  = \new_[34870]_  & \new_[34865]_ ;
  assign \new_[34875]_  = A233 & A232;
  assign \new_[34876]_  = A202 & \new_[34875]_ ;
  assign \new_[34879]_  = A266 & A265;
  assign \new_[34882]_  = A299 & ~A298;
  assign \new_[34883]_  = \new_[34882]_  & \new_[34879]_ ;
  assign \new_[34884]_  = \new_[34883]_  & \new_[34876]_ ;
  assign \new_[34888]_  = ~A168 & A169;
  assign \new_[34889]_  = A170 & \new_[34888]_ ;
  assign \new_[34893]_  = A201 & ~A200;
  assign \new_[34894]_  = A199 & \new_[34893]_ ;
  assign \new_[34895]_  = \new_[34894]_  & \new_[34889]_ ;
  assign \new_[34899]_  = A233 & A232;
  assign \new_[34900]_  = A202 & \new_[34899]_ ;
  assign \new_[34903]_  = ~A266 & ~A265;
  assign \new_[34906]_  = A299 & ~A298;
  assign \new_[34907]_  = \new_[34906]_  & \new_[34903]_ ;
  assign \new_[34908]_  = \new_[34907]_  & \new_[34900]_ ;
  assign \new_[34912]_  = ~A168 & A169;
  assign \new_[34913]_  = A170 & \new_[34912]_ ;
  assign \new_[34917]_  = A201 & ~A200;
  assign \new_[34918]_  = A199 & \new_[34917]_ ;
  assign \new_[34919]_  = \new_[34918]_  & \new_[34913]_ ;
  assign \new_[34923]_  = A233 & ~A232;
  assign \new_[34924]_  = A202 & \new_[34923]_ ;
  assign \new_[34927]_  = ~A266 & A265;
  assign \new_[34930]_  = A268 & A267;
  assign \new_[34931]_  = \new_[34930]_  & \new_[34927]_ ;
  assign \new_[34932]_  = \new_[34931]_  & \new_[34924]_ ;
  assign \new_[34936]_  = ~A168 & A169;
  assign \new_[34937]_  = A170 & \new_[34936]_ ;
  assign \new_[34941]_  = A201 & ~A200;
  assign \new_[34942]_  = A199 & \new_[34941]_ ;
  assign \new_[34943]_  = \new_[34942]_  & \new_[34937]_ ;
  assign \new_[34947]_  = A233 & ~A232;
  assign \new_[34948]_  = A202 & \new_[34947]_ ;
  assign \new_[34951]_  = ~A266 & A265;
  assign \new_[34954]_  = A269 & A267;
  assign \new_[34955]_  = \new_[34954]_  & \new_[34951]_ ;
  assign \new_[34956]_  = \new_[34955]_  & \new_[34948]_ ;
  assign \new_[34960]_  = ~A168 & A169;
  assign \new_[34961]_  = A170 & \new_[34960]_ ;
  assign \new_[34965]_  = A201 & ~A200;
  assign \new_[34966]_  = A199 & \new_[34965]_ ;
  assign \new_[34967]_  = \new_[34966]_  & \new_[34961]_ ;
  assign \new_[34971]_  = ~A234 & ~A233;
  assign \new_[34972]_  = A202 & \new_[34971]_ ;
  assign \new_[34975]_  = A266 & A265;
  assign \new_[34978]_  = A299 & ~A298;
  assign \new_[34979]_  = \new_[34978]_  & \new_[34975]_ ;
  assign \new_[34980]_  = \new_[34979]_  & \new_[34972]_ ;
  assign \new_[34984]_  = ~A168 & A169;
  assign \new_[34985]_  = A170 & \new_[34984]_ ;
  assign \new_[34989]_  = A201 & ~A200;
  assign \new_[34990]_  = A199 & \new_[34989]_ ;
  assign \new_[34991]_  = \new_[34990]_  & \new_[34985]_ ;
  assign \new_[34995]_  = ~A234 & ~A233;
  assign \new_[34996]_  = A202 & \new_[34995]_ ;
  assign \new_[34999]_  = ~A267 & ~A266;
  assign \new_[35002]_  = A299 & ~A298;
  assign \new_[35003]_  = \new_[35002]_  & \new_[34999]_ ;
  assign \new_[35004]_  = \new_[35003]_  & \new_[34996]_ ;
  assign \new_[35008]_  = ~A168 & A169;
  assign \new_[35009]_  = A170 & \new_[35008]_ ;
  assign \new_[35013]_  = A201 & ~A200;
  assign \new_[35014]_  = A199 & \new_[35013]_ ;
  assign \new_[35015]_  = \new_[35014]_  & \new_[35009]_ ;
  assign \new_[35019]_  = ~A234 & ~A233;
  assign \new_[35020]_  = A202 & \new_[35019]_ ;
  assign \new_[35023]_  = ~A266 & ~A265;
  assign \new_[35026]_  = A299 & ~A298;
  assign \new_[35027]_  = \new_[35026]_  & \new_[35023]_ ;
  assign \new_[35028]_  = \new_[35027]_  & \new_[35020]_ ;
  assign \new_[35032]_  = ~A168 & A169;
  assign \new_[35033]_  = A170 & \new_[35032]_ ;
  assign \new_[35037]_  = A201 & ~A200;
  assign \new_[35038]_  = A199 & \new_[35037]_ ;
  assign \new_[35039]_  = \new_[35038]_  & \new_[35033]_ ;
  assign \new_[35043]_  = ~A233 & A232;
  assign \new_[35044]_  = A202 & \new_[35043]_ ;
  assign \new_[35047]_  = A235 & A234;
  assign \new_[35050]_  = ~A300 & A298;
  assign \new_[35051]_  = \new_[35050]_  & \new_[35047]_ ;
  assign \new_[35052]_  = \new_[35051]_  & \new_[35044]_ ;
  assign \new_[35056]_  = ~A168 & A169;
  assign \new_[35057]_  = A170 & \new_[35056]_ ;
  assign \new_[35061]_  = A201 & ~A200;
  assign \new_[35062]_  = A199 & \new_[35061]_ ;
  assign \new_[35063]_  = \new_[35062]_  & \new_[35057]_ ;
  assign \new_[35067]_  = ~A233 & A232;
  assign \new_[35068]_  = A202 & \new_[35067]_ ;
  assign \new_[35071]_  = A235 & A234;
  assign \new_[35074]_  = A299 & A298;
  assign \new_[35075]_  = \new_[35074]_  & \new_[35071]_ ;
  assign \new_[35076]_  = \new_[35075]_  & \new_[35068]_ ;
  assign \new_[35080]_  = ~A168 & A169;
  assign \new_[35081]_  = A170 & \new_[35080]_ ;
  assign \new_[35085]_  = A201 & ~A200;
  assign \new_[35086]_  = A199 & \new_[35085]_ ;
  assign \new_[35087]_  = \new_[35086]_  & \new_[35081]_ ;
  assign \new_[35091]_  = ~A233 & A232;
  assign \new_[35092]_  = A202 & \new_[35091]_ ;
  assign \new_[35095]_  = A235 & A234;
  assign \new_[35098]_  = ~A299 & ~A298;
  assign \new_[35099]_  = \new_[35098]_  & \new_[35095]_ ;
  assign \new_[35100]_  = \new_[35099]_  & \new_[35092]_ ;
  assign \new_[35104]_  = ~A168 & A169;
  assign \new_[35105]_  = A170 & \new_[35104]_ ;
  assign \new_[35109]_  = A201 & ~A200;
  assign \new_[35110]_  = A199 & \new_[35109]_ ;
  assign \new_[35111]_  = \new_[35110]_  & \new_[35105]_ ;
  assign \new_[35115]_  = ~A233 & A232;
  assign \new_[35116]_  = A202 & \new_[35115]_ ;
  assign \new_[35119]_  = A235 & A234;
  assign \new_[35122]_  = A266 & ~A265;
  assign \new_[35123]_  = \new_[35122]_  & \new_[35119]_ ;
  assign \new_[35124]_  = \new_[35123]_  & \new_[35116]_ ;
  assign \new_[35128]_  = ~A168 & A169;
  assign \new_[35129]_  = A170 & \new_[35128]_ ;
  assign \new_[35133]_  = A201 & ~A200;
  assign \new_[35134]_  = A199 & \new_[35133]_ ;
  assign \new_[35135]_  = \new_[35134]_  & \new_[35129]_ ;
  assign \new_[35139]_  = ~A233 & A232;
  assign \new_[35140]_  = A202 & \new_[35139]_ ;
  assign \new_[35143]_  = A236 & A234;
  assign \new_[35146]_  = ~A300 & A298;
  assign \new_[35147]_  = \new_[35146]_  & \new_[35143]_ ;
  assign \new_[35148]_  = \new_[35147]_  & \new_[35140]_ ;
  assign \new_[35152]_  = ~A168 & A169;
  assign \new_[35153]_  = A170 & \new_[35152]_ ;
  assign \new_[35157]_  = A201 & ~A200;
  assign \new_[35158]_  = A199 & \new_[35157]_ ;
  assign \new_[35159]_  = \new_[35158]_  & \new_[35153]_ ;
  assign \new_[35163]_  = ~A233 & A232;
  assign \new_[35164]_  = A202 & \new_[35163]_ ;
  assign \new_[35167]_  = A236 & A234;
  assign \new_[35170]_  = A299 & A298;
  assign \new_[35171]_  = \new_[35170]_  & \new_[35167]_ ;
  assign \new_[35172]_  = \new_[35171]_  & \new_[35164]_ ;
  assign \new_[35176]_  = ~A168 & A169;
  assign \new_[35177]_  = A170 & \new_[35176]_ ;
  assign \new_[35181]_  = A201 & ~A200;
  assign \new_[35182]_  = A199 & \new_[35181]_ ;
  assign \new_[35183]_  = \new_[35182]_  & \new_[35177]_ ;
  assign \new_[35187]_  = ~A233 & A232;
  assign \new_[35188]_  = A202 & \new_[35187]_ ;
  assign \new_[35191]_  = A236 & A234;
  assign \new_[35194]_  = ~A299 & ~A298;
  assign \new_[35195]_  = \new_[35194]_  & \new_[35191]_ ;
  assign \new_[35196]_  = \new_[35195]_  & \new_[35188]_ ;
  assign \new_[35200]_  = ~A168 & A169;
  assign \new_[35201]_  = A170 & \new_[35200]_ ;
  assign \new_[35205]_  = A201 & ~A200;
  assign \new_[35206]_  = A199 & \new_[35205]_ ;
  assign \new_[35207]_  = \new_[35206]_  & \new_[35201]_ ;
  assign \new_[35211]_  = ~A233 & A232;
  assign \new_[35212]_  = A202 & \new_[35211]_ ;
  assign \new_[35215]_  = A236 & A234;
  assign \new_[35218]_  = A266 & ~A265;
  assign \new_[35219]_  = \new_[35218]_  & \new_[35215]_ ;
  assign \new_[35220]_  = \new_[35219]_  & \new_[35212]_ ;
  assign \new_[35224]_  = ~A168 & A169;
  assign \new_[35225]_  = A170 & \new_[35224]_ ;
  assign \new_[35229]_  = A201 & ~A200;
  assign \new_[35230]_  = A199 & \new_[35229]_ ;
  assign \new_[35231]_  = \new_[35230]_  & \new_[35225]_ ;
  assign \new_[35235]_  = ~A233 & ~A232;
  assign \new_[35236]_  = A202 & \new_[35235]_ ;
  assign \new_[35239]_  = A266 & A265;
  assign \new_[35242]_  = A299 & ~A298;
  assign \new_[35243]_  = \new_[35242]_  & \new_[35239]_ ;
  assign \new_[35244]_  = \new_[35243]_  & \new_[35236]_ ;
  assign \new_[35248]_  = ~A168 & A169;
  assign \new_[35249]_  = A170 & \new_[35248]_ ;
  assign \new_[35253]_  = A201 & ~A200;
  assign \new_[35254]_  = A199 & \new_[35253]_ ;
  assign \new_[35255]_  = \new_[35254]_  & \new_[35249]_ ;
  assign \new_[35259]_  = ~A233 & ~A232;
  assign \new_[35260]_  = A202 & \new_[35259]_ ;
  assign \new_[35263]_  = ~A267 & ~A266;
  assign \new_[35266]_  = A299 & ~A298;
  assign \new_[35267]_  = \new_[35266]_  & \new_[35263]_ ;
  assign \new_[35268]_  = \new_[35267]_  & \new_[35260]_ ;
  assign \new_[35272]_  = ~A168 & A169;
  assign \new_[35273]_  = A170 & \new_[35272]_ ;
  assign \new_[35277]_  = A201 & ~A200;
  assign \new_[35278]_  = A199 & \new_[35277]_ ;
  assign \new_[35279]_  = \new_[35278]_  & \new_[35273]_ ;
  assign \new_[35283]_  = ~A233 & ~A232;
  assign \new_[35284]_  = A202 & \new_[35283]_ ;
  assign \new_[35287]_  = ~A266 & ~A265;
  assign \new_[35290]_  = A299 & ~A298;
  assign \new_[35291]_  = \new_[35290]_  & \new_[35287]_ ;
  assign \new_[35292]_  = \new_[35291]_  & \new_[35284]_ ;
  assign \new_[35296]_  = ~A168 & A169;
  assign \new_[35297]_  = A170 & \new_[35296]_ ;
  assign \new_[35301]_  = A201 & ~A200;
  assign \new_[35302]_  = A199 & \new_[35301]_ ;
  assign \new_[35303]_  = \new_[35302]_  & \new_[35297]_ ;
  assign \new_[35307]_  = A233 & A232;
  assign \new_[35308]_  = A203 & \new_[35307]_ ;
  assign \new_[35311]_  = ~A267 & A265;
  assign \new_[35314]_  = A299 & ~A298;
  assign \new_[35315]_  = \new_[35314]_  & \new_[35311]_ ;
  assign \new_[35316]_  = \new_[35315]_  & \new_[35308]_ ;
  assign \new_[35320]_  = ~A168 & A169;
  assign \new_[35321]_  = A170 & \new_[35320]_ ;
  assign \new_[35325]_  = A201 & ~A200;
  assign \new_[35326]_  = A199 & \new_[35325]_ ;
  assign \new_[35327]_  = \new_[35326]_  & \new_[35321]_ ;
  assign \new_[35331]_  = A233 & A232;
  assign \new_[35332]_  = A203 & \new_[35331]_ ;
  assign \new_[35335]_  = A266 & A265;
  assign \new_[35338]_  = A299 & ~A298;
  assign \new_[35339]_  = \new_[35338]_  & \new_[35335]_ ;
  assign \new_[35340]_  = \new_[35339]_  & \new_[35332]_ ;
  assign \new_[35344]_  = ~A168 & A169;
  assign \new_[35345]_  = A170 & \new_[35344]_ ;
  assign \new_[35349]_  = A201 & ~A200;
  assign \new_[35350]_  = A199 & \new_[35349]_ ;
  assign \new_[35351]_  = \new_[35350]_  & \new_[35345]_ ;
  assign \new_[35355]_  = A233 & A232;
  assign \new_[35356]_  = A203 & \new_[35355]_ ;
  assign \new_[35359]_  = ~A266 & ~A265;
  assign \new_[35362]_  = A299 & ~A298;
  assign \new_[35363]_  = \new_[35362]_  & \new_[35359]_ ;
  assign \new_[35364]_  = \new_[35363]_  & \new_[35356]_ ;
  assign \new_[35368]_  = ~A168 & A169;
  assign \new_[35369]_  = A170 & \new_[35368]_ ;
  assign \new_[35373]_  = A201 & ~A200;
  assign \new_[35374]_  = A199 & \new_[35373]_ ;
  assign \new_[35375]_  = \new_[35374]_  & \new_[35369]_ ;
  assign \new_[35379]_  = A233 & ~A232;
  assign \new_[35380]_  = A203 & \new_[35379]_ ;
  assign \new_[35383]_  = ~A266 & A265;
  assign \new_[35386]_  = A268 & A267;
  assign \new_[35387]_  = \new_[35386]_  & \new_[35383]_ ;
  assign \new_[35388]_  = \new_[35387]_  & \new_[35380]_ ;
  assign \new_[35392]_  = ~A168 & A169;
  assign \new_[35393]_  = A170 & \new_[35392]_ ;
  assign \new_[35397]_  = A201 & ~A200;
  assign \new_[35398]_  = A199 & \new_[35397]_ ;
  assign \new_[35399]_  = \new_[35398]_  & \new_[35393]_ ;
  assign \new_[35403]_  = A233 & ~A232;
  assign \new_[35404]_  = A203 & \new_[35403]_ ;
  assign \new_[35407]_  = ~A266 & A265;
  assign \new_[35410]_  = A269 & A267;
  assign \new_[35411]_  = \new_[35410]_  & \new_[35407]_ ;
  assign \new_[35412]_  = \new_[35411]_  & \new_[35404]_ ;
  assign \new_[35416]_  = ~A168 & A169;
  assign \new_[35417]_  = A170 & \new_[35416]_ ;
  assign \new_[35421]_  = A201 & ~A200;
  assign \new_[35422]_  = A199 & \new_[35421]_ ;
  assign \new_[35423]_  = \new_[35422]_  & \new_[35417]_ ;
  assign \new_[35427]_  = ~A234 & ~A233;
  assign \new_[35428]_  = A203 & \new_[35427]_ ;
  assign \new_[35431]_  = A266 & A265;
  assign \new_[35434]_  = A299 & ~A298;
  assign \new_[35435]_  = \new_[35434]_  & \new_[35431]_ ;
  assign \new_[35436]_  = \new_[35435]_  & \new_[35428]_ ;
  assign \new_[35440]_  = ~A168 & A169;
  assign \new_[35441]_  = A170 & \new_[35440]_ ;
  assign \new_[35445]_  = A201 & ~A200;
  assign \new_[35446]_  = A199 & \new_[35445]_ ;
  assign \new_[35447]_  = \new_[35446]_  & \new_[35441]_ ;
  assign \new_[35451]_  = ~A234 & ~A233;
  assign \new_[35452]_  = A203 & \new_[35451]_ ;
  assign \new_[35455]_  = ~A267 & ~A266;
  assign \new_[35458]_  = A299 & ~A298;
  assign \new_[35459]_  = \new_[35458]_  & \new_[35455]_ ;
  assign \new_[35460]_  = \new_[35459]_  & \new_[35452]_ ;
  assign \new_[35464]_  = ~A168 & A169;
  assign \new_[35465]_  = A170 & \new_[35464]_ ;
  assign \new_[35469]_  = A201 & ~A200;
  assign \new_[35470]_  = A199 & \new_[35469]_ ;
  assign \new_[35471]_  = \new_[35470]_  & \new_[35465]_ ;
  assign \new_[35475]_  = ~A234 & ~A233;
  assign \new_[35476]_  = A203 & \new_[35475]_ ;
  assign \new_[35479]_  = ~A266 & ~A265;
  assign \new_[35482]_  = A299 & ~A298;
  assign \new_[35483]_  = \new_[35482]_  & \new_[35479]_ ;
  assign \new_[35484]_  = \new_[35483]_  & \new_[35476]_ ;
  assign \new_[35488]_  = ~A168 & A169;
  assign \new_[35489]_  = A170 & \new_[35488]_ ;
  assign \new_[35493]_  = A201 & ~A200;
  assign \new_[35494]_  = A199 & \new_[35493]_ ;
  assign \new_[35495]_  = \new_[35494]_  & \new_[35489]_ ;
  assign \new_[35499]_  = ~A233 & A232;
  assign \new_[35500]_  = A203 & \new_[35499]_ ;
  assign \new_[35503]_  = A235 & A234;
  assign \new_[35506]_  = ~A300 & A298;
  assign \new_[35507]_  = \new_[35506]_  & \new_[35503]_ ;
  assign \new_[35508]_  = \new_[35507]_  & \new_[35500]_ ;
  assign \new_[35512]_  = ~A168 & A169;
  assign \new_[35513]_  = A170 & \new_[35512]_ ;
  assign \new_[35517]_  = A201 & ~A200;
  assign \new_[35518]_  = A199 & \new_[35517]_ ;
  assign \new_[35519]_  = \new_[35518]_  & \new_[35513]_ ;
  assign \new_[35523]_  = ~A233 & A232;
  assign \new_[35524]_  = A203 & \new_[35523]_ ;
  assign \new_[35527]_  = A235 & A234;
  assign \new_[35530]_  = A299 & A298;
  assign \new_[35531]_  = \new_[35530]_  & \new_[35527]_ ;
  assign \new_[35532]_  = \new_[35531]_  & \new_[35524]_ ;
  assign \new_[35536]_  = ~A168 & A169;
  assign \new_[35537]_  = A170 & \new_[35536]_ ;
  assign \new_[35541]_  = A201 & ~A200;
  assign \new_[35542]_  = A199 & \new_[35541]_ ;
  assign \new_[35543]_  = \new_[35542]_  & \new_[35537]_ ;
  assign \new_[35547]_  = ~A233 & A232;
  assign \new_[35548]_  = A203 & \new_[35547]_ ;
  assign \new_[35551]_  = A235 & A234;
  assign \new_[35554]_  = ~A299 & ~A298;
  assign \new_[35555]_  = \new_[35554]_  & \new_[35551]_ ;
  assign \new_[35556]_  = \new_[35555]_  & \new_[35548]_ ;
  assign \new_[35560]_  = ~A168 & A169;
  assign \new_[35561]_  = A170 & \new_[35560]_ ;
  assign \new_[35565]_  = A201 & ~A200;
  assign \new_[35566]_  = A199 & \new_[35565]_ ;
  assign \new_[35567]_  = \new_[35566]_  & \new_[35561]_ ;
  assign \new_[35571]_  = ~A233 & A232;
  assign \new_[35572]_  = A203 & \new_[35571]_ ;
  assign \new_[35575]_  = A235 & A234;
  assign \new_[35578]_  = A266 & ~A265;
  assign \new_[35579]_  = \new_[35578]_  & \new_[35575]_ ;
  assign \new_[35580]_  = \new_[35579]_  & \new_[35572]_ ;
  assign \new_[35584]_  = ~A168 & A169;
  assign \new_[35585]_  = A170 & \new_[35584]_ ;
  assign \new_[35589]_  = A201 & ~A200;
  assign \new_[35590]_  = A199 & \new_[35589]_ ;
  assign \new_[35591]_  = \new_[35590]_  & \new_[35585]_ ;
  assign \new_[35595]_  = ~A233 & A232;
  assign \new_[35596]_  = A203 & \new_[35595]_ ;
  assign \new_[35599]_  = A236 & A234;
  assign \new_[35602]_  = ~A300 & A298;
  assign \new_[35603]_  = \new_[35602]_  & \new_[35599]_ ;
  assign \new_[35604]_  = \new_[35603]_  & \new_[35596]_ ;
  assign \new_[35608]_  = ~A168 & A169;
  assign \new_[35609]_  = A170 & \new_[35608]_ ;
  assign \new_[35613]_  = A201 & ~A200;
  assign \new_[35614]_  = A199 & \new_[35613]_ ;
  assign \new_[35615]_  = \new_[35614]_  & \new_[35609]_ ;
  assign \new_[35619]_  = ~A233 & A232;
  assign \new_[35620]_  = A203 & \new_[35619]_ ;
  assign \new_[35623]_  = A236 & A234;
  assign \new_[35626]_  = A299 & A298;
  assign \new_[35627]_  = \new_[35626]_  & \new_[35623]_ ;
  assign \new_[35628]_  = \new_[35627]_  & \new_[35620]_ ;
  assign \new_[35632]_  = ~A168 & A169;
  assign \new_[35633]_  = A170 & \new_[35632]_ ;
  assign \new_[35637]_  = A201 & ~A200;
  assign \new_[35638]_  = A199 & \new_[35637]_ ;
  assign \new_[35639]_  = \new_[35638]_  & \new_[35633]_ ;
  assign \new_[35643]_  = ~A233 & A232;
  assign \new_[35644]_  = A203 & \new_[35643]_ ;
  assign \new_[35647]_  = A236 & A234;
  assign \new_[35650]_  = ~A299 & ~A298;
  assign \new_[35651]_  = \new_[35650]_  & \new_[35647]_ ;
  assign \new_[35652]_  = \new_[35651]_  & \new_[35644]_ ;
  assign \new_[35656]_  = ~A168 & A169;
  assign \new_[35657]_  = A170 & \new_[35656]_ ;
  assign \new_[35661]_  = A201 & ~A200;
  assign \new_[35662]_  = A199 & \new_[35661]_ ;
  assign \new_[35663]_  = \new_[35662]_  & \new_[35657]_ ;
  assign \new_[35667]_  = ~A233 & A232;
  assign \new_[35668]_  = A203 & \new_[35667]_ ;
  assign \new_[35671]_  = A236 & A234;
  assign \new_[35674]_  = A266 & ~A265;
  assign \new_[35675]_  = \new_[35674]_  & \new_[35671]_ ;
  assign \new_[35676]_  = \new_[35675]_  & \new_[35668]_ ;
  assign \new_[35680]_  = ~A168 & A169;
  assign \new_[35681]_  = A170 & \new_[35680]_ ;
  assign \new_[35685]_  = A201 & ~A200;
  assign \new_[35686]_  = A199 & \new_[35685]_ ;
  assign \new_[35687]_  = \new_[35686]_  & \new_[35681]_ ;
  assign \new_[35691]_  = ~A233 & ~A232;
  assign \new_[35692]_  = A203 & \new_[35691]_ ;
  assign \new_[35695]_  = A266 & A265;
  assign \new_[35698]_  = A299 & ~A298;
  assign \new_[35699]_  = \new_[35698]_  & \new_[35695]_ ;
  assign \new_[35700]_  = \new_[35699]_  & \new_[35692]_ ;
  assign \new_[35704]_  = ~A168 & A169;
  assign \new_[35705]_  = A170 & \new_[35704]_ ;
  assign \new_[35709]_  = A201 & ~A200;
  assign \new_[35710]_  = A199 & \new_[35709]_ ;
  assign \new_[35711]_  = \new_[35710]_  & \new_[35705]_ ;
  assign \new_[35715]_  = ~A233 & ~A232;
  assign \new_[35716]_  = A203 & \new_[35715]_ ;
  assign \new_[35719]_  = ~A267 & ~A266;
  assign \new_[35722]_  = A299 & ~A298;
  assign \new_[35723]_  = \new_[35722]_  & \new_[35719]_ ;
  assign \new_[35724]_  = \new_[35723]_  & \new_[35716]_ ;
  assign \new_[35728]_  = ~A168 & A169;
  assign \new_[35729]_  = A170 & \new_[35728]_ ;
  assign \new_[35733]_  = A201 & ~A200;
  assign \new_[35734]_  = A199 & \new_[35733]_ ;
  assign \new_[35735]_  = \new_[35734]_  & \new_[35729]_ ;
  assign \new_[35739]_  = ~A233 & ~A232;
  assign \new_[35740]_  = A203 & \new_[35739]_ ;
  assign \new_[35743]_  = ~A266 & ~A265;
  assign \new_[35746]_  = A299 & ~A298;
  assign \new_[35747]_  = \new_[35746]_  & \new_[35743]_ ;
  assign \new_[35748]_  = \new_[35747]_  & \new_[35740]_ ;
  assign \new_[35752]_  = A167 & A169;
  assign \new_[35753]_  = ~A170 & \new_[35752]_ ;
  assign \new_[35757]_  = A200 & A199;
  assign \new_[35758]_  = A166 & \new_[35757]_ ;
  assign \new_[35759]_  = \new_[35758]_  & \new_[35753]_ ;
  assign \new_[35763]_  = A265 & A233;
  assign \new_[35764]_  = A232 & \new_[35763]_ ;
  assign \new_[35767]_  = ~A269 & ~A268;
  assign \new_[35770]_  = A299 & ~A298;
  assign \new_[35771]_  = \new_[35770]_  & \new_[35767]_ ;
  assign \new_[35772]_  = \new_[35771]_  & \new_[35764]_ ;
  assign \new_[35776]_  = A167 & A169;
  assign \new_[35777]_  = ~A170 & \new_[35776]_ ;
  assign \new_[35781]_  = A200 & A199;
  assign \new_[35782]_  = A166 & \new_[35781]_ ;
  assign \new_[35783]_  = \new_[35782]_  & \new_[35777]_ ;
  assign \new_[35787]_  = ~A236 & ~A235;
  assign \new_[35788]_  = ~A233 & \new_[35787]_ ;
  assign \new_[35791]_  = A266 & A265;
  assign \new_[35794]_  = A299 & ~A298;
  assign \new_[35795]_  = \new_[35794]_  & \new_[35791]_ ;
  assign \new_[35796]_  = \new_[35795]_  & \new_[35788]_ ;
  assign \new_[35800]_  = A167 & A169;
  assign \new_[35801]_  = ~A170 & \new_[35800]_ ;
  assign \new_[35805]_  = A200 & A199;
  assign \new_[35806]_  = A166 & \new_[35805]_ ;
  assign \new_[35807]_  = \new_[35806]_  & \new_[35801]_ ;
  assign \new_[35811]_  = ~A236 & ~A235;
  assign \new_[35812]_  = ~A233 & \new_[35811]_ ;
  assign \new_[35815]_  = ~A267 & ~A266;
  assign \new_[35818]_  = A299 & ~A298;
  assign \new_[35819]_  = \new_[35818]_  & \new_[35815]_ ;
  assign \new_[35820]_  = \new_[35819]_  & \new_[35812]_ ;
  assign \new_[35824]_  = A167 & A169;
  assign \new_[35825]_  = ~A170 & \new_[35824]_ ;
  assign \new_[35829]_  = A200 & A199;
  assign \new_[35830]_  = A166 & \new_[35829]_ ;
  assign \new_[35831]_  = \new_[35830]_  & \new_[35825]_ ;
  assign \new_[35835]_  = ~A236 & ~A235;
  assign \new_[35836]_  = ~A233 & \new_[35835]_ ;
  assign \new_[35839]_  = ~A266 & ~A265;
  assign \new_[35842]_  = A299 & ~A298;
  assign \new_[35843]_  = \new_[35842]_  & \new_[35839]_ ;
  assign \new_[35844]_  = \new_[35843]_  & \new_[35836]_ ;
  assign \new_[35848]_  = A167 & A169;
  assign \new_[35849]_  = ~A170 & \new_[35848]_ ;
  assign \new_[35853]_  = A200 & A199;
  assign \new_[35854]_  = A166 & \new_[35853]_ ;
  assign \new_[35855]_  = \new_[35854]_  & \new_[35849]_ ;
  assign \new_[35859]_  = ~A266 & ~A234;
  assign \new_[35860]_  = ~A233 & \new_[35859]_ ;
  assign \new_[35863]_  = ~A269 & ~A268;
  assign \new_[35866]_  = A299 & ~A298;
  assign \new_[35867]_  = \new_[35866]_  & \new_[35863]_ ;
  assign \new_[35868]_  = \new_[35867]_  & \new_[35860]_ ;
  assign \new_[35872]_  = A167 & A169;
  assign \new_[35873]_  = ~A170 & \new_[35872]_ ;
  assign \new_[35877]_  = A200 & A199;
  assign \new_[35878]_  = A166 & \new_[35877]_ ;
  assign \new_[35879]_  = \new_[35878]_  & \new_[35873]_ ;
  assign \new_[35883]_  = A234 & ~A233;
  assign \new_[35884]_  = A232 & \new_[35883]_ ;
  assign \new_[35887]_  = A298 & A235;
  assign \new_[35890]_  = ~A302 & ~A301;
  assign \new_[35891]_  = \new_[35890]_  & \new_[35887]_ ;
  assign \new_[35892]_  = \new_[35891]_  & \new_[35884]_ ;
  assign \new_[35896]_  = A167 & A169;
  assign \new_[35897]_  = ~A170 & \new_[35896]_ ;
  assign \new_[35901]_  = A200 & A199;
  assign \new_[35902]_  = A166 & \new_[35901]_ ;
  assign \new_[35903]_  = \new_[35902]_  & \new_[35897]_ ;
  assign \new_[35907]_  = A234 & ~A233;
  assign \new_[35908]_  = A232 & \new_[35907]_ ;
  assign \new_[35911]_  = A298 & A236;
  assign \new_[35914]_  = ~A302 & ~A301;
  assign \new_[35915]_  = \new_[35914]_  & \new_[35911]_ ;
  assign \new_[35916]_  = \new_[35915]_  & \new_[35908]_ ;
  assign \new_[35920]_  = A167 & A169;
  assign \new_[35921]_  = ~A170 & \new_[35920]_ ;
  assign \new_[35925]_  = A200 & A199;
  assign \new_[35926]_  = A166 & \new_[35925]_ ;
  assign \new_[35927]_  = \new_[35926]_  & \new_[35921]_ ;
  assign \new_[35931]_  = ~A266 & ~A233;
  assign \new_[35932]_  = ~A232 & \new_[35931]_ ;
  assign \new_[35935]_  = ~A269 & ~A268;
  assign \new_[35938]_  = A299 & ~A298;
  assign \new_[35939]_  = \new_[35938]_  & \new_[35935]_ ;
  assign \new_[35940]_  = \new_[35939]_  & \new_[35932]_ ;
  assign \new_[35944]_  = A167 & A169;
  assign \new_[35945]_  = ~A170 & \new_[35944]_ ;
  assign \new_[35949]_  = ~A202 & ~A200;
  assign \new_[35950]_  = A166 & \new_[35949]_ ;
  assign \new_[35951]_  = \new_[35950]_  & \new_[35945]_ ;
  assign \new_[35955]_  = A233 & A232;
  assign \new_[35956]_  = ~A203 & \new_[35955]_ ;
  assign \new_[35959]_  = ~A267 & A265;
  assign \new_[35962]_  = A299 & ~A298;
  assign \new_[35963]_  = \new_[35962]_  & \new_[35959]_ ;
  assign \new_[35964]_  = \new_[35963]_  & \new_[35956]_ ;
  assign \new_[35968]_  = A167 & A169;
  assign \new_[35969]_  = ~A170 & \new_[35968]_ ;
  assign \new_[35973]_  = ~A202 & ~A200;
  assign \new_[35974]_  = A166 & \new_[35973]_ ;
  assign \new_[35975]_  = \new_[35974]_  & \new_[35969]_ ;
  assign \new_[35979]_  = A233 & A232;
  assign \new_[35980]_  = ~A203 & \new_[35979]_ ;
  assign \new_[35983]_  = A266 & A265;
  assign \new_[35986]_  = A299 & ~A298;
  assign \new_[35987]_  = \new_[35986]_  & \new_[35983]_ ;
  assign \new_[35988]_  = \new_[35987]_  & \new_[35980]_ ;
  assign \new_[35992]_  = A167 & A169;
  assign \new_[35993]_  = ~A170 & \new_[35992]_ ;
  assign \new_[35997]_  = ~A202 & ~A200;
  assign \new_[35998]_  = A166 & \new_[35997]_ ;
  assign \new_[35999]_  = \new_[35998]_  & \new_[35993]_ ;
  assign \new_[36003]_  = A233 & A232;
  assign \new_[36004]_  = ~A203 & \new_[36003]_ ;
  assign \new_[36007]_  = ~A266 & ~A265;
  assign \new_[36010]_  = A299 & ~A298;
  assign \new_[36011]_  = \new_[36010]_  & \new_[36007]_ ;
  assign \new_[36012]_  = \new_[36011]_  & \new_[36004]_ ;
  assign \new_[36016]_  = A167 & A169;
  assign \new_[36017]_  = ~A170 & \new_[36016]_ ;
  assign \new_[36021]_  = ~A202 & ~A200;
  assign \new_[36022]_  = A166 & \new_[36021]_ ;
  assign \new_[36023]_  = \new_[36022]_  & \new_[36017]_ ;
  assign \new_[36027]_  = A233 & ~A232;
  assign \new_[36028]_  = ~A203 & \new_[36027]_ ;
  assign \new_[36031]_  = ~A266 & A265;
  assign \new_[36034]_  = A268 & A267;
  assign \new_[36035]_  = \new_[36034]_  & \new_[36031]_ ;
  assign \new_[36036]_  = \new_[36035]_  & \new_[36028]_ ;
  assign \new_[36040]_  = A167 & A169;
  assign \new_[36041]_  = ~A170 & \new_[36040]_ ;
  assign \new_[36045]_  = ~A202 & ~A200;
  assign \new_[36046]_  = A166 & \new_[36045]_ ;
  assign \new_[36047]_  = \new_[36046]_  & \new_[36041]_ ;
  assign \new_[36051]_  = A233 & ~A232;
  assign \new_[36052]_  = ~A203 & \new_[36051]_ ;
  assign \new_[36055]_  = ~A266 & A265;
  assign \new_[36058]_  = A269 & A267;
  assign \new_[36059]_  = \new_[36058]_  & \new_[36055]_ ;
  assign \new_[36060]_  = \new_[36059]_  & \new_[36052]_ ;
  assign \new_[36064]_  = A167 & A169;
  assign \new_[36065]_  = ~A170 & \new_[36064]_ ;
  assign \new_[36069]_  = ~A202 & ~A200;
  assign \new_[36070]_  = A166 & \new_[36069]_ ;
  assign \new_[36071]_  = \new_[36070]_  & \new_[36065]_ ;
  assign \new_[36075]_  = ~A234 & ~A233;
  assign \new_[36076]_  = ~A203 & \new_[36075]_ ;
  assign \new_[36079]_  = A266 & A265;
  assign \new_[36082]_  = A299 & ~A298;
  assign \new_[36083]_  = \new_[36082]_  & \new_[36079]_ ;
  assign \new_[36084]_  = \new_[36083]_  & \new_[36076]_ ;
  assign \new_[36088]_  = A167 & A169;
  assign \new_[36089]_  = ~A170 & \new_[36088]_ ;
  assign \new_[36093]_  = ~A202 & ~A200;
  assign \new_[36094]_  = A166 & \new_[36093]_ ;
  assign \new_[36095]_  = \new_[36094]_  & \new_[36089]_ ;
  assign \new_[36099]_  = ~A234 & ~A233;
  assign \new_[36100]_  = ~A203 & \new_[36099]_ ;
  assign \new_[36103]_  = ~A267 & ~A266;
  assign \new_[36106]_  = A299 & ~A298;
  assign \new_[36107]_  = \new_[36106]_  & \new_[36103]_ ;
  assign \new_[36108]_  = \new_[36107]_  & \new_[36100]_ ;
  assign \new_[36112]_  = A167 & A169;
  assign \new_[36113]_  = ~A170 & \new_[36112]_ ;
  assign \new_[36117]_  = ~A202 & ~A200;
  assign \new_[36118]_  = A166 & \new_[36117]_ ;
  assign \new_[36119]_  = \new_[36118]_  & \new_[36113]_ ;
  assign \new_[36123]_  = ~A234 & ~A233;
  assign \new_[36124]_  = ~A203 & \new_[36123]_ ;
  assign \new_[36127]_  = ~A266 & ~A265;
  assign \new_[36130]_  = A299 & ~A298;
  assign \new_[36131]_  = \new_[36130]_  & \new_[36127]_ ;
  assign \new_[36132]_  = \new_[36131]_  & \new_[36124]_ ;
  assign \new_[36136]_  = A167 & A169;
  assign \new_[36137]_  = ~A170 & \new_[36136]_ ;
  assign \new_[36141]_  = ~A202 & ~A200;
  assign \new_[36142]_  = A166 & \new_[36141]_ ;
  assign \new_[36143]_  = \new_[36142]_  & \new_[36137]_ ;
  assign \new_[36147]_  = ~A233 & A232;
  assign \new_[36148]_  = ~A203 & \new_[36147]_ ;
  assign \new_[36151]_  = A235 & A234;
  assign \new_[36154]_  = ~A300 & A298;
  assign \new_[36155]_  = \new_[36154]_  & \new_[36151]_ ;
  assign \new_[36156]_  = \new_[36155]_  & \new_[36148]_ ;
  assign \new_[36160]_  = A167 & A169;
  assign \new_[36161]_  = ~A170 & \new_[36160]_ ;
  assign \new_[36165]_  = ~A202 & ~A200;
  assign \new_[36166]_  = A166 & \new_[36165]_ ;
  assign \new_[36167]_  = \new_[36166]_  & \new_[36161]_ ;
  assign \new_[36171]_  = ~A233 & A232;
  assign \new_[36172]_  = ~A203 & \new_[36171]_ ;
  assign \new_[36175]_  = A235 & A234;
  assign \new_[36178]_  = A299 & A298;
  assign \new_[36179]_  = \new_[36178]_  & \new_[36175]_ ;
  assign \new_[36180]_  = \new_[36179]_  & \new_[36172]_ ;
  assign \new_[36184]_  = A167 & A169;
  assign \new_[36185]_  = ~A170 & \new_[36184]_ ;
  assign \new_[36189]_  = ~A202 & ~A200;
  assign \new_[36190]_  = A166 & \new_[36189]_ ;
  assign \new_[36191]_  = \new_[36190]_  & \new_[36185]_ ;
  assign \new_[36195]_  = ~A233 & A232;
  assign \new_[36196]_  = ~A203 & \new_[36195]_ ;
  assign \new_[36199]_  = A235 & A234;
  assign \new_[36202]_  = ~A299 & ~A298;
  assign \new_[36203]_  = \new_[36202]_  & \new_[36199]_ ;
  assign \new_[36204]_  = \new_[36203]_  & \new_[36196]_ ;
  assign \new_[36208]_  = A167 & A169;
  assign \new_[36209]_  = ~A170 & \new_[36208]_ ;
  assign \new_[36213]_  = ~A202 & ~A200;
  assign \new_[36214]_  = A166 & \new_[36213]_ ;
  assign \new_[36215]_  = \new_[36214]_  & \new_[36209]_ ;
  assign \new_[36219]_  = ~A233 & A232;
  assign \new_[36220]_  = ~A203 & \new_[36219]_ ;
  assign \new_[36223]_  = A235 & A234;
  assign \new_[36226]_  = A266 & ~A265;
  assign \new_[36227]_  = \new_[36226]_  & \new_[36223]_ ;
  assign \new_[36228]_  = \new_[36227]_  & \new_[36220]_ ;
  assign \new_[36232]_  = A167 & A169;
  assign \new_[36233]_  = ~A170 & \new_[36232]_ ;
  assign \new_[36237]_  = ~A202 & ~A200;
  assign \new_[36238]_  = A166 & \new_[36237]_ ;
  assign \new_[36239]_  = \new_[36238]_  & \new_[36233]_ ;
  assign \new_[36243]_  = ~A233 & A232;
  assign \new_[36244]_  = ~A203 & \new_[36243]_ ;
  assign \new_[36247]_  = A236 & A234;
  assign \new_[36250]_  = ~A300 & A298;
  assign \new_[36251]_  = \new_[36250]_  & \new_[36247]_ ;
  assign \new_[36252]_  = \new_[36251]_  & \new_[36244]_ ;
  assign \new_[36256]_  = A167 & A169;
  assign \new_[36257]_  = ~A170 & \new_[36256]_ ;
  assign \new_[36261]_  = ~A202 & ~A200;
  assign \new_[36262]_  = A166 & \new_[36261]_ ;
  assign \new_[36263]_  = \new_[36262]_  & \new_[36257]_ ;
  assign \new_[36267]_  = ~A233 & A232;
  assign \new_[36268]_  = ~A203 & \new_[36267]_ ;
  assign \new_[36271]_  = A236 & A234;
  assign \new_[36274]_  = A299 & A298;
  assign \new_[36275]_  = \new_[36274]_  & \new_[36271]_ ;
  assign \new_[36276]_  = \new_[36275]_  & \new_[36268]_ ;
  assign \new_[36280]_  = A167 & A169;
  assign \new_[36281]_  = ~A170 & \new_[36280]_ ;
  assign \new_[36285]_  = ~A202 & ~A200;
  assign \new_[36286]_  = A166 & \new_[36285]_ ;
  assign \new_[36287]_  = \new_[36286]_  & \new_[36281]_ ;
  assign \new_[36291]_  = ~A233 & A232;
  assign \new_[36292]_  = ~A203 & \new_[36291]_ ;
  assign \new_[36295]_  = A236 & A234;
  assign \new_[36298]_  = ~A299 & ~A298;
  assign \new_[36299]_  = \new_[36298]_  & \new_[36295]_ ;
  assign \new_[36300]_  = \new_[36299]_  & \new_[36292]_ ;
  assign \new_[36304]_  = A167 & A169;
  assign \new_[36305]_  = ~A170 & \new_[36304]_ ;
  assign \new_[36309]_  = ~A202 & ~A200;
  assign \new_[36310]_  = A166 & \new_[36309]_ ;
  assign \new_[36311]_  = \new_[36310]_  & \new_[36305]_ ;
  assign \new_[36315]_  = ~A233 & A232;
  assign \new_[36316]_  = ~A203 & \new_[36315]_ ;
  assign \new_[36319]_  = A236 & A234;
  assign \new_[36322]_  = A266 & ~A265;
  assign \new_[36323]_  = \new_[36322]_  & \new_[36319]_ ;
  assign \new_[36324]_  = \new_[36323]_  & \new_[36316]_ ;
  assign \new_[36328]_  = A167 & A169;
  assign \new_[36329]_  = ~A170 & \new_[36328]_ ;
  assign \new_[36333]_  = ~A202 & ~A200;
  assign \new_[36334]_  = A166 & \new_[36333]_ ;
  assign \new_[36335]_  = \new_[36334]_  & \new_[36329]_ ;
  assign \new_[36339]_  = ~A233 & ~A232;
  assign \new_[36340]_  = ~A203 & \new_[36339]_ ;
  assign \new_[36343]_  = A266 & A265;
  assign \new_[36346]_  = A299 & ~A298;
  assign \new_[36347]_  = \new_[36346]_  & \new_[36343]_ ;
  assign \new_[36348]_  = \new_[36347]_  & \new_[36340]_ ;
  assign \new_[36352]_  = A167 & A169;
  assign \new_[36353]_  = ~A170 & \new_[36352]_ ;
  assign \new_[36357]_  = ~A202 & ~A200;
  assign \new_[36358]_  = A166 & \new_[36357]_ ;
  assign \new_[36359]_  = \new_[36358]_  & \new_[36353]_ ;
  assign \new_[36363]_  = ~A233 & ~A232;
  assign \new_[36364]_  = ~A203 & \new_[36363]_ ;
  assign \new_[36367]_  = ~A267 & ~A266;
  assign \new_[36370]_  = A299 & ~A298;
  assign \new_[36371]_  = \new_[36370]_  & \new_[36367]_ ;
  assign \new_[36372]_  = \new_[36371]_  & \new_[36364]_ ;
  assign \new_[36376]_  = A167 & A169;
  assign \new_[36377]_  = ~A170 & \new_[36376]_ ;
  assign \new_[36381]_  = ~A202 & ~A200;
  assign \new_[36382]_  = A166 & \new_[36381]_ ;
  assign \new_[36383]_  = \new_[36382]_  & \new_[36377]_ ;
  assign \new_[36387]_  = ~A233 & ~A232;
  assign \new_[36388]_  = ~A203 & \new_[36387]_ ;
  assign \new_[36391]_  = ~A266 & ~A265;
  assign \new_[36394]_  = A299 & ~A298;
  assign \new_[36395]_  = \new_[36394]_  & \new_[36391]_ ;
  assign \new_[36396]_  = \new_[36395]_  & \new_[36388]_ ;
  assign \new_[36400]_  = A167 & A169;
  assign \new_[36401]_  = ~A170 & \new_[36400]_ ;
  assign \new_[36405]_  = ~A201 & ~A200;
  assign \new_[36406]_  = A166 & \new_[36405]_ ;
  assign \new_[36407]_  = \new_[36406]_  & \new_[36401]_ ;
  assign \new_[36411]_  = A265 & A233;
  assign \new_[36412]_  = A232 & \new_[36411]_ ;
  assign \new_[36415]_  = ~A269 & ~A268;
  assign \new_[36418]_  = A299 & ~A298;
  assign \new_[36419]_  = \new_[36418]_  & \new_[36415]_ ;
  assign \new_[36420]_  = \new_[36419]_  & \new_[36412]_ ;
  assign \new_[36424]_  = A167 & A169;
  assign \new_[36425]_  = ~A170 & \new_[36424]_ ;
  assign \new_[36429]_  = ~A201 & ~A200;
  assign \new_[36430]_  = A166 & \new_[36429]_ ;
  assign \new_[36431]_  = \new_[36430]_  & \new_[36425]_ ;
  assign \new_[36435]_  = ~A236 & ~A235;
  assign \new_[36436]_  = ~A233 & \new_[36435]_ ;
  assign \new_[36439]_  = A266 & A265;
  assign \new_[36442]_  = A299 & ~A298;
  assign \new_[36443]_  = \new_[36442]_  & \new_[36439]_ ;
  assign \new_[36444]_  = \new_[36443]_  & \new_[36436]_ ;
  assign \new_[36448]_  = A167 & A169;
  assign \new_[36449]_  = ~A170 & \new_[36448]_ ;
  assign \new_[36453]_  = ~A201 & ~A200;
  assign \new_[36454]_  = A166 & \new_[36453]_ ;
  assign \new_[36455]_  = \new_[36454]_  & \new_[36449]_ ;
  assign \new_[36459]_  = ~A236 & ~A235;
  assign \new_[36460]_  = ~A233 & \new_[36459]_ ;
  assign \new_[36463]_  = ~A267 & ~A266;
  assign \new_[36466]_  = A299 & ~A298;
  assign \new_[36467]_  = \new_[36466]_  & \new_[36463]_ ;
  assign \new_[36468]_  = \new_[36467]_  & \new_[36460]_ ;
  assign \new_[36472]_  = A167 & A169;
  assign \new_[36473]_  = ~A170 & \new_[36472]_ ;
  assign \new_[36477]_  = ~A201 & ~A200;
  assign \new_[36478]_  = A166 & \new_[36477]_ ;
  assign \new_[36479]_  = \new_[36478]_  & \new_[36473]_ ;
  assign \new_[36483]_  = ~A236 & ~A235;
  assign \new_[36484]_  = ~A233 & \new_[36483]_ ;
  assign \new_[36487]_  = ~A266 & ~A265;
  assign \new_[36490]_  = A299 & ~A298;
  assign \new_[36491]_  = \new_[36490]_  & \new_[36487]_ ;
  assign \new_[36492]_  = \new_[36491]_  & \new_[36484]_ ;
  assign \new_[36496]_  = A167 & A169;
  assign \new_[36497]_  = ~A170 & \new_[36496]_ ;
  assign \new_[36501]_  = ~A201 & ~A200;
  assign \new_[36502]_  = A166 & \new_[36501]_ ;
  assign \new_[36503]_  = \new_[36502]_  & \new_[36497]_ ;
  assign \new_[36507]_  = ~A266 & ~A234;
  assign \new_[36508]_  = ~A233 & \new_[36507]_ ;
  assign \new_[36511]_  = ~A269 & ~A268;
  assign \new_[36514]_  = A299 & ~A298;
  assign \new_[36515]_  = \new_[36514]_  & \new_[36511]_ ;
  assign \new_[36516]_  = \new_[36515]_  & \new_[36508]_ ;
  assign \new_[36520]_  = A167 & A169;
  assign \new_[36521]_  = ~A170 & \new_[36520]_ ;
  assign \new_[36525]_  = ~A201 & ~A200;
  assign \new_[36526]_  = A166 & \new_[36525]_ ;
  assign \new_[36527]_  = \new_[36526]_  & \new_[36521]_ ;
  assign \new_[36531]_  = A234 & ~A233;
  assign \new_[36532]_  = A232 & \new_[36531]_ ;
  assign \new_[36535]_  = A298 & A235;
  assign \new_[36538]_  = ~A302 & ~A301;
  assign \new_[36539]_  = \new_[36538]_  & \new_[36535]_ ;
  assign \new_[36540]_  = \new_[36539]_  & \new_[36532]_ ;
  assign \new_[36544]_  = A167 & A169;
  assign \new_[36545]_  = ~A170 & \new_[36544]_ ;
  assign \new_[36549]_  = ~A201 & ~A200;
  assign \new_[36550]_  = A166 & \new_[36549]_ ;
  assign \new_[36551]_  = \new_[36550]_  & \new_[36545]_ ;
  assign \new_[36555]_  = A234 & ~A233;
  assign \new_[36556]_  = A232 & \new_[36555]_ ;
  assign \new_[36559]_  = A298 & A236;
  assign \new_[36562]_  = ~A302 & ~A301;
  assign \new_[36563]_  = \new_[36562]_  & \new_[36559]_ ;
  assign \new_[36564]_  = \new_[36563]_  & \new_[36556]_ ;
  assign \new_[36568]_  = A167 & A169;
  assign \new_[36569]_  = ~A170 & \new_[36568]_ ;
  assign \new_[36573]_  = ~A201 & ~A200;
  assign \new_[36574]_  = A166 & \new_[36573]_ ;
  assign \new_[36575]_  = \new_[36574]_  & \new_[36569]_ ;
  assign \new_[36579]_  = ~A266 & ~A233;
  assign \new_[36580]_  = ~A232 & \new_[36579]_ ;
  assign \new_[36583]_  = ~A269 & ~A268;
  assign \new_[36586]_  = A299 & ~A298;
  assign \new_[36587]_  = \new_[36586]_  & \new_[36583]_ ;
  assign \new_[36588]_  = \new_[36587]_  & \new_[36580]_ ;
  assign \new_[36592]_  = A167 & A169;
  assign \new_[36593]_  = ~A170 & \new_[36592]_ ;
  assign \new_[36597]_  = ~A200 & ~A199;
  assign \new_[36598]_  = A166 & \new_[36597]_ ;
  assign \new_[36599]_  = \new_[36598]_  & \new_[36593]_ ;
  assign \new_[36603]_  = A265 & A233;
  assign \new_[36604]_  = A232 & \new_[36603]_ ;
  assign \new_[36607]_  = ~A269 & ~A268;
  assign \new_[36610]_  = A299 & ~A298;
  assign \new_[36611]_  = \new_[36610]_  & \new_[36607]_ ;
  assign \new_[36612]_  = \new_[36611]_  & \new_[36604]_ ;
  assign \new_[36616]_  = A167 & A169;
  assign \new_[36617]_  = ~A170 & \new_[36616]_ ;
  assign \new_[36621]_  = ~A200 & ~A199;
  assign \new_[36622]_  = A166 & \new_[36621]_ ;
  assign \new_[36623]_  = \new_[36622]_  & \new_[36617]_ ;
  assign \new_[36627]_  = ~A236 & ~A235;
  assign \new_[36628]_  = ~A233 & \new_[36627]_ ;
  assign \new_[36631]_  = A266 & A265;
  assign \new_[36634]_  = A299 & ~A298;
  assign \new_[36635]_  = \new_[36634]_  & \new_[36631]_ ;
  assign \new_[36636]_  = \new_[36635]_  & \new_[36628]_ ;
  assign \new_[36640]_  = A167 & A169;
  assign \new_[36641]_  = ~A170 & \new_[36640]_ ;
  assign \new_[36645]_  = ~A200 & ~A199;
  assign \new_[36646]_  = A166 & \new_[36645]_ ;
  assign \new_[36647]_  = \new_[36646]_  & \new_[36641]_ ;
  assign \new_[36651]_  = ~A236 & ~A235;
  assign \new_[36652]_  = ~A233 & \new_[36651]_ ;
  assign \new_[36655]_  = ~A267 & ~A266;
  assign \new_[36658]_  = A299 & ~A298;
  assign \new_[36659]_  = \new_[36658]_  & \new_[36655]_ ;
  assign \new_[36660]_  = \new_[36659]_  & \new_[36652]_ ;
  assign \new_[36664]_  = A167 & A169;
  assign \new_[36665]_  = ~A170 & \new_[36664]_ ;
  assign \new_[36669]_  = ~A200 & ~A199;
  assign \new_[36670]_  = A166 & \new_[36669]_ ;
  assign \new_[36671]_  = \new_[36670]_  & \new_[36665]_ ;
  assign \new_[36675]_  = ~A236 & ~A235;
  assign \new_[36676]_  = ~A233 & \new_[36675]_ ;
  assign \new_[36679]_  = ~A266 & ~A265;
  assign \new_[36682]_  = A299 & ~A298;
  assign \new_[36683]_  = \new_[36682]_  & \new_[36679]_ ;
  assign \new_[36684]_  = \new_[36683]_  & \new_[36676]_ ;
  assign \new_[36688]_  = A167 & A169;
  assign \new_[36689]_  = ~A170 & \new_[36688]_ ;
  assign \new_[36693]_  = ~A200 & ~A199;
  assign \new_[36694]_  = A166 & \new_[36693]_ ;
  assign \new_[36695]_  = \new_[36694]_  & \new_[36689]_ ;
  assign \new_[36699]_  = ~A266 & ~A234;
  assign \new_[36700]_  = ~A233 & \new_[36699]_ ;
  assign \new_[36703]_  = ~A269 & ~A268;
  assign \new_[36706]_  = A299 & ~A298;
  assign \new_[36707]_  = \new_[36706]_  & \new_[36703]_ ;
  assign \new_[36708]_  = \new_[36707]_  & \new_[36700]_ ;
  assign \new_[36712]_  = A167 & A169;
  assign \new_[36713]_  = ~A170 & \new_[36712]_ ;
  assign \new_[36717]_  = ~A200 & ~A199;
  assign \new_[36718]_  = A166 & \new_[36717]_ ;
  assign \new_[36719]_  = \new_[36718]_  & \new_[36713]_ ;
  assign \new_[36723]_  = A234 & ~A233;
  assign \new_[36724]_  = A232 & \new_[36723]_ ;
  assign \new_[36727]_  = A298 & A235;
  assign \new_[36730]_  = ~A302 & ~A301;
  assign \new_[36731]_  = \new_[36730]_  & \new_[36727]_ ;
  assign \new_[36732]_  = \new_[36731]_  & \new_[36724]_ ;
  assign \new_[36736]_  = A167 & A169;
  assign \new_[36737]_  = ~A170 & \new_[36736]_ ;
  assign \new_[36741]_  = ~A200 & ~A199;
  assign \new_[36742]_  = A166 & \new_[36741]_ ;
  assign \new_[36743]_  = \new_[36742]_  & \new_[36737]_ ;
  assign \new_[36747]_  = A234 & ~A233;
  assign \new_[36748]_  = A232 & \new_[36747]_ ;
  assign \new_[36751]_  = A298 & A236;
  assign \new_[36754]_  = ~A302 & ~A301;
  assign \new_[36755]_  = \new_[36754]_  & \new_[36751]_ ;
  assign \new_[36756]_  = \new_[36755]_  & \new_[36748]_ ;
  assign \new_[36760]_  = A167 & A169;
  assign \new_[36761]_  = ~A170 & \new_[36760]_ ;
  assign \new_[36765]_  = ~A200 & ~A199;
  assign \new_[36766]_  = A166 & \new_[36765]_ ;
  assign \new_[36767]_  = \new_[36766]_  & \new_[36761]_ ;
  assign \new_[36771]_  = ~A266 & ~A233;
  assign \new_[36772]_  = ~A232 & \new_[36771]_ ;
  assign \new_[36775]_  = ~A269 & ~A268;
  assign \new_[36778]_  = A299 & ~A298;
  assign \new_[36779]_  = \new_[36778]_  & \new_[36775]_ ;
  assign \new_[36780]_  = \new_[36779]_  & \new_[36772]_ ;
  assign \new_[36784]_  = ~A167 & A169;
  assign \new_[36785]_  = ~A170 & \new_[36784]_ ;
  assign \new_[36789]_  = A200 & A199;
  assign \new_[36790]_  = ~A166 & \new_[36789]_ ;
  assign \new_[36791]_  = \new_[36790]_  & \new_[36785]_ ;
  assign \new_[36795]_  = A265 & A233;
  assign \new_[36796]_  = A232 & \new_[36795]_ ;
  assign \new_[36799]_  = ~A269 & ~A268;
  assign \new_[36802]_  = A299 & ~A298;
  assign \new_[36803]_  = \new_[36802]_  & \new_[36799]_ ;
  assign \new_[36804]_  = \new_[36803]_  & \new_[36796]_ ;
  assign \new_[36808]_  = ~A167 & A169;
  assign \new_[36809]_  = ~A170 & \new_[36808]_ ;
  assign \new_[36813]_  = A200 & A199;
  assign \new_[36814]_  = ~A166 & \new_[36813]_ ;
  assign \new_[36815]_  = \new_[36814]_  & \new_[36809]_ ;
  assign \new_[36819]_  = ~A236 & ~A235;
  assign \new_[36820]_  = ~A233 & \new_[36819]_ ;
  assign \new_[36823]_  = A266 & A265;
  assign \new_[36826]_  = A299 & ~A298;
  assign \new_[36827]_  = \new_[36826]_  & \new_[36823]_ ;
  assign \new_[36828]_  = \new_[36827]_  & \new_[36820]_ ;
  assign \new_[36832]_  = ~A167 & A169;
  assign \new_[36833]_  = ~A170 & \new_[36832]_ ;
  assign \new_[36837]_  = A200 & A199;
  assign \new_[36838]_  = ~A166 & \new_[36837]_ ;
  assign \new_[36839]_  = \new_[36838]_  & \new_[36833]_ ;
  assign \new_[36843]_  = ~A236 & ~A235;
  assign \new_[36844]_  = ~A233 & \new_[36843]_ ;
  assign \new_[36847]_  = ~A267 & ~A266;
  assign \new_[36850]_  = A299 & ~A298;
  assign \new_[36851]_  = \new_[36850]_  & \new_[36847]_ ;
  assign \new_[36852]_  = \new_[36851]_  & \new_[36844]_ ;
  assign \new_[36856]_  = ~A167 & A169;
  assign \new_[36857]_  = ~A170 & \new_[36856]_ ;
  assign \new_[36861]_  = A200 & A199;
  assign \new_[36862]_  = ~A166 & \new_[36861]_ ;
  assign \new_[36863]_  = \new_[36862]_  & \new_[36857]_ ;
  assign \new_[36867]_  = ~A236 & ~A235;
  assign \new_[36868]_  = ~A233 & \new_[36867]_ ;
  assign \new_[36871]_  = ~A266 & ~A265;
  assign \new_[36874]_  = A299 & ~A298;
  assign \new_[36875]_  = \new_[36874]_  & \new_[36871]_ ;
  assign \new_[36876]_  = \new_[36875]_  & \new_[36868]_ ;
  assign \new_[36880]_  = ~A167 & A169;
  assign \new_[36881]_  = ~A170 & \new_[36880]_ ;
  assign \new_[36885]_  = A200 & A199;
  assign \new_[36886]_  = ~A166 & \new_[36885]_ ;
  assign \new_[36887]_  = \new_[36886]_  & \new_[36881]_ ;
  assign \new_[36891]_  = ~A266 & ~A234;
  assign \new_[36892]_  = ~A233 & \new_[36891]_ ;
  assign \new_[36895]_  = ~A269 & ~A268;
  assign \new_[36898]_  = A299 & ~A298;
  assign \new_[36899]_  = \new_[36898]_  & \new_[36895]_ ;
  assign \new_[36900]_  = \new_[36899]_  & \new_[36892]_ ;
  assign \new_[36904]_  = ~A167 & A169;
  assign \new_[36905]_  = ~A170 & \new_[36904]_ ;
  assign \new_[36909]_  = A200 & A199;
  assign \new_[36910]_  = ~A166 & \new_[36909]_ ;
  assign \new_[36911]_  = \new_[36910]_  & \new_[36905]_ ;
  assign \new_[36915]_  = A234 & ~A233;
  assign \new_[36916]_  = A232 & \new_[36915]_ ;
  assign \new_[36919]_  = A298 & A235;
  assign \new_[36922]_  = ~A302 & ~A301;
  assign \new_[36923]_  = \new_[36922]_  & \new_[36919]_ ;
  assign \new_[36924]_  = \new_[36923]_  & \new_[36916]_ ;
  assign \new_[36928]_  = ~A167 & A169;
  assign \new_[36929]_  = ~A170 & \new_[36928]_ ;
  assign \new_[36933]_  = A200 & A199;
  assign \new_[36934]_  = ~A166 & \new_[36933]_ ;
  assign \new_[36935]_  = \new_[36934]_  & \new_[36929]_ ;
  assign \new_[36939]_  = A234 & ~A233;
  assign \new_[36940]_  = A232 & \new_[36939]_ ;
  assign \new_[36943]_  = A298 & A236;
  assign \new_[36946]_  = ~A302 & ~A301;
  assign \new_[36947]_  = \new_[36946]_  & \new_[36943]_ ;
  assign \new_[36948]_  = \new_[36947]_  & \new_[36940]_ ;
  assign \new_[36952]_  = ~A167 & A169;
  assign \new_[36953]_  = ~A170 & \new_[36952]_ ;
  assign \new_[36957]_  = A200 & A199;
  assign \new_[36958]_  = ~A166 & \new_[36957]_ ;
  assign \new_[36959]_  = \new_[36958]_  & \new_[36953]_ ;
  assign \new_[36963]_  = ~A266 & ~A233;
  assign \new_[36964]_  = ~A232 & \new_[36963]_ ;
  assign \new_[36967]_  = ~A269 & ~A268;
  assign \new_[36970]_  = A299 & ~A298;
  assign \new_[36971]_  = \new_[36970]_  & \new_[36967]_ ;
  assign \new_[36972]_  = \new_[36971]_  & \new_[36964]_ ;
  assign \new_[36976]_  = ~A167 & A169;
  assign \new_[36977]_  = ~A170 & \new_[36976]_ ;
  assign \new_[36981]_  = ~A202 & ~A200;
  assign \new_[36982]_  = ~A166 & \new_[36981]_ ;
  assign \new_[36983]_  = \new_[36982]_  & \new_[36977]_ ;
  assign \new_[36987]_  = A233 & A232;
  assign \new_[36988]_  = ~A203 & \new_[36987]_ ;
  assign \new_[36991]_  = ~A267 & A265;
  assign \new_[36994]_  = A299 & ~A298;
  assign \new_[36995]_  = \new_[36994]_  & \new_[36991]_ ;
  assign \new_[36996]_  = \new_[36995]_  & \new_[36988]_ ;
  assign \new_[37000]_  = ~A167 & A169;
  assign \new_[37001]_  = ~A170 & \new_[37000]_ ;
  assign \new_[37005]_  = ~A202 & ~A200;
  assign \new_[37006]_  = ~A166 & \new_[37005]_ ;
  assign \new_[37007]_  = \new_[37006]_  & \new_[37001]_ ;
  assign \new_[37011]_  = A233 & A232;
  assign \new_[37012]_  = ~A203 & \new_[37011]_ ;
  assign \new_[37015]_  = A266 & A265;
  assign \new_[37018]_  = A299 & ~A298;
  assign \new_[37019]_  = \new_[37018]_  & \new_[37015]_ ;
  assign \new_[37020]_  = \new_[37019]_  & \new_[37012]_ ;
  assign \new_[37024]_  = ~A167 & A169;
  assign \new_[37025]_  = ~A170 & \new_[37024]_ ;
  assign \new_[37029]_  = ~A202 & ~A200;
  assign \new_[37030]_  = ~A166 & \new_[37029]_ ;
  assign \new_[37031]_  = \new_[37030]_  & \new_[37025]_ ;
  assign \new_[37035]_  = A233 & A232;
  assign \new_[37036]_  = ~A203 & \new_[37035]_ ;
  assign \new_[37039]_  = ~A266 & ~A265;
  assign \new_[37042]_  = A299 & ~A298;
  assign \new_[37043]_  = \new_[37042]_  & \new_[37039]_ ;
  assign \new_[37044]_  = \new_[37043]_  & \new_[37036]_ ;
  assign \new_[37048]_  = ~A167 & A169;
  assign \new_[37049]_  = ~A170 & \new_[37048]_ ;
  assign \new_[37053]_  = ~A202 & ~A200;
  assign \new_[37054]_  = ~A166 & \new_[37053]_ ;
  assign \new_[37055]_  = \new_[37054]_  & \new_[37049]_ ;
  assign \new_[37059]_  = A233 & ~A232;
  assign \new_[37060]_  = ~A203 & \new_[37059]_ ;
  assign \new_[37063]_  = ~A266 & A265;
  assign \new_[37066]_  = A268 & A267;
  assign \new_[37067]_  = \new_[37066]_  & \new_[37063]_ ;
  assign \new_[37068]_  = \new_[37067]_  & \new_[37060]_ ;
  assign \new_[37072]_  = ~A167 & A169;
  assign \new_[37073]_  = ~A170 & \new_[37072]_ ;
  assign \new_[37077]_  = ~A202 & ~A200;
  assign \new_[37078]_  = ~A166 & \new_[37077]_ ;
  assign \new_[37079]_  = \new_[37078]_  & \new_[37073]_ ;
  assign \new_[37083]_  = A233 & ~A232;
  assign \new_[37084]_  = ~A203 & \new_[37083]_ ;
  assign \new_[37087]_  = ~A266 & A265;
  assign \new_[37090]_  = A269 & A267;
  assign \new_[37091]_  = \new_[37090]_  & \new_[37087]_ ;
  assign \new_[37092]_  = \new_[37091]_  & \new_[37084]_ ;
  assign \new_[37096]_  = ~A167 & A169;
  assign \new_[37097]_  = ~A170 & \new_[37096]_ ;
  assign \new_[37101]_  = ~A202 & ~A200;
  assign \new_[37102]_  = ~A166 & \new_[37101]_ ;
  assign \new_[37103]_  = \new_[37102]_  & \new_[37097]_ ;
  assign \new_[37107]_  = ~A234 & ~A233;
  assign \new_[37108]_  = ~A203 & \new_[37107]_ ;
  assign \new_[37111]_  = A266 & A265;
  assign \new_[37114]_  = A299 & ~A298;
  assign \new_[37115]_  = \new_[37114]_  & \new_[37111]_ ;
  assign \new_[37116]_  = \new_[37115]_  & \new_[37108]_ ;
  assign \new_[37120]_  = ~A167 & A169;
  assign \new_[37121]_  = ~A170 & \new_[37120]_ ;
  assign \new_[37125]_  = ~A202 & ~A200;
  assign \new_[37126]_  = ~A166 & \new_[37125]_ ;
  assign \new_[37127]_  = \new_[37126]_  & \new_[37121]_ ;
  assign \new_[37131]_  = ~A234 & ~A233;
  assign \new_[37132]_  = ~A203 & \new_[37131]_ ;
  assign \new_[37135]_  = ~A267 & ~A266;
  assign \new_[37138]_  = A299 & ~A298;
  assign \new_[37139]_  = \new_[37138]_  & \new_[37135]_ ;
  assign \new_[37140]_  = \new_[37139]_  & \new_[37132]_ ;
  assign \new_[37144]_  = ~A167 & A169;
  assign \new_[37145]_  = ~A170 & \new_[37144]_ ;
  assign \new_[37149]_  = ~A202 & ~A200;
  assign \new_[37150]_  = ~A166 & \new_[37149]_ ;
  assign \new_[37151]_  = \new_[37150]_  & \new_[37145]_ ;
  assign \new_[37155]_  = ~A234 & ~A233;
  assign \new_[37156]_  = ~A203 & \new_[37155]_ ;
  assign \new_[37159]_  = ~A266 & ~A265;
  assign \new_[37162]_  = A299 & ~A298;
  assign \new_[37163]_  = \new_[37162]_  & \new_[37159]_ ;
  assign \new_[37164]_  = \new_[37163]_  & \new_[37156]_ ;
  assign \new_[37168]_  = ~A167 & A169;
  assign \new_[37169]_  = ~A170 & \new_[37168]_ ;
  assign \new_[37173]_  = ~A202 & ~A200;
  assign \new_[37174]_  = ~A166 & \new_[37173]_ ;
  assign \new_[37175]_  = \new_[37174]_  & \new_[37169]_ ;
  assign \new_[37179]_  = ~A233 & A232;
  assign \new_[37180]_  = ~A203 & \new_[37179]_ ;
  assign \new_[37183]_  = A235 & A234;
  assign \new_[37186]_  = ~A300 & A298;
  assign \new_[37187]_  = \new_[37186]_  & \new_[37183]_ ;
  assign \new_[37188]_  = \new_[37187]_  & \new_[37180]_ ;
  assign \new_[37192]_  = ~A167 & A169;
  assign \new_[37193]_  = ~A170 & \new_[37192]_ ;
  assign \new_[37197]_  = ~A202 & ~A200;
  assign \new_[37198]_  = ~A166 & \new_[37197]_ ;
  assign \new_[37199]_  = \new_[37198]_  & \new_[37193]_ ;
  assign \new_[37203]_  = ~A233 & A232;
  assign \new_[37204]_  = ~A203 & \new_[37203]_ ;
  assign \new_[37207]_  = A235 & A234;
  assign \new_[37210]_  = A299 & A298;
  assign \new_[37211]_  = \new_[37210]_  & \new_[37207]_ ;
  assign \new_[37212]_  = \new_[37211]_  & \new_[37204]_ ;
  assign \new_[37216]_  = ~A167 & A169;
  assign \new_[37217]_  = ~A170 & \new_[37216]_ ;
  assign \new_[37221]_  = ~A202 & ~A200;
  assign \new_[37222]_  = ~A166 & \new_[37221]_ ;
  assign \new_[37223]_  = \new_[37222]_  & \new_[37217]_ ;
  assign \new_[37227]_  = ~A233 & A232;
  assign \new_[37228]_  = ~A203 & \new_[37227]_ ;
  assign \new_[37231]_  = A235 & A234;
  assign \new_[37234]_  = ~A299 & ~A298;
  assign \new_[37235]_  = \new_[37234]_  & \new_[37231]_ ;
  assign \new_[37236]_  = \new_[37235]_  & \new_[37228]_ ;
  assign \new_[37240]_  = ~A167 & A169;
  assign \new_[37241]_  = ~A170 & \new_[37240]_ ;
  assign \new_[37245]_  = ~A202 & ~A200;
  assign \new_[37246]_  = ~A166 & \new_[37245]_ ;
  assign \new_[37247]_  = \new_[37246]_  & \new_[37241]_ ;
  assign \new_[37251]_  = ~A233 & A232;
  assign \new_[37252]_  = ~A203 & \new_[37251]_ ;
  assign \new_[37255]_  = A235 & A234;
  assign \new_[37258]_  = A266 & ~A265;
  assign \new_[37259]_  = \new_[37258]_  & \new_[37255]_ ;
  assign \new_[37260]_  = \new_[37259]_  & \new_[37252]_ ;
  assign \new_[37264]_  = ~A167 & A169;
  assign \new_[37265]_  = ~A170 & \new_[37264]_ ;
  assign \new_[37269]_  = ~A202 & ~A200;
  assign \new_[37270]_  = ~A166 & \new_[37269]_ ;
  assign \new_[37271]_  = \new_[37270]_  & \new_[37265]_ ;
  assign \new_[37275]_  = ~A233 & A232;
  assign \new_[37276]_  = ~A203 & \new_[37275]_ ;
  assign \new_[37279]_  = A236 & A234;
  assign \new_[37282]_  = ~A300 & A298;
  assign \new_[37283]_  = \new_[37282]_  & \new_[37279]_ ;
  assign \new_[37284]_  = \new_[37283]_  & \new_[37276]_ ;
  assign \new_[37288]_  = ~A167 & A169;
  assign \new_[37289]_  = ~A170 & \new_[37288]_ ;
  assign \new_[37293]_  = ~A202 & ~A200;
  assign \new_[37294]_  = ~A166 & \new_[37293]_ ;
  assign \new_[37295]_  = \new_[37294]_  & \new_[37289]_ ;
  assign \new_[37299]_  = ~A233 & A232;
  assign \new_[37300]_  = ~A203 & \new_[37299]_ ;
  assign \new_[37303]_  = A236 & A234;
  assign \new_[37306]_  = A299 & A298;
  assign \new_[37307]_  = \new_[37306]_  & \new_[37303]_ ;
  assign \new_[37308]_  = \new_[37307]_  & \new_[37300]_ ;
  assign \new_[37312]_  = ~A167 & A169;
  assign \new_[37313]_  = ~A170 & \new_[37312]_ ;
  assign \new_[37317]_  = ~A202 & ~A200;
  assign \new_[37318]_  = ~A166 & \new_[37317]_ ;
  assign \new_[37319]_  = \new_[37318]_  & \new_[37313]_ ;
  assign \new_[37323]_  = ~A233 & A232;
  assign \new_[37324]_  = ~A203 & \new_[37323]_ ;
  assign \new_[37327]_  = A236 & A234;
  assign \new_[37330]_  = ~A299 & ~A298;
  assign \new_[37331]_  = \new_[37330]_  & \new_[37327]_ ;
  assign \new_[37332]_  = \new_[37331]_  & \new_[37324]_ ;
  assign \new_[37336]_  = ~A167 & A169;
  assign \new_[37337]_  = ~A170 & \new_[37336]_ ;
  assign \new_[37341]_  = ~A202 & ~A200;
  assign \new_[37342]_  = ~A166 & \new_[37341]_ ;
  assign \new_[37343]_  = \new_[37342]_  & \new_[37337]_ ;
  assign \new_[37347]_  = ~A233 & A232;
  assign \new_[37348]_  = ~A203 & \new_[37347]_ ;
  assign \new_[37351]_  = A236 & A234;
  assign \new_[37354]_  = A266 & ~A265;
  assign \new_[37355]_  = \new_[37354]_  & \new_[37351]_ ;
  assign \new_[37356]_  = \new_[37355]_  & \new_[37348]_ ;
  assign \new_[37360]_  = ~A167 & A169;
  assign \new_[37361]_  = ~A170 & \new_[37360]_ ;
  assign \new_[37365]_  = ~A202 & ~A200;
  assign \new_[37366]_  = ~A166 & \new_[37365]_ ;
  assign \new_[37367]_  = \new_[37366]_  & \new_[37361]_ ;
  assign \new_[37371]_  = ~A233 & ~A232;
  assign \new_[37372]_  = ~A203 & \new_[37371]_ ;
  assign \new_[37375]_  = A266 & A265;
  assign \new_[37378]_  = A299 & ~A298;
  assign \new_[37379]_  = \new_[37378]_  & \new_[37375]_ ;
  assign \new_[37380]_  = \new_[37379]_  & \new_[37372]_ ;
  assign \new_[37384]_  = ~A167 & A169;
  assign \new_[37385]_  = ~A170 & \new_[37384]_ ;
  assign \new_[37389]_  = ~A202 & ~A200;
  assign \new_[37390]_  = ~A166 & \new_[37389]_ ;
  assign \new_[37391]_  = \new_[37390]_  & \new_[37385]_ ;
  assign \new_[37395]_  = ~A233 & ~A232;
  assign \new_[37396]_  = ~A203 & \new_[37395]_ ;
  assign \new_[37399]_  = ~A267 & ~A266;
  assign \new_[37402]_  = A299 & ~A298;
  assign \new_[37403]_  = \new_[37402]_  & \new_[37399]_ ;
  assign \new_[37404]_  = \new_[37403]_  & \new_[37396]_ ;
  assign \new_[37408]_  = ~A167 & A169;
  assign \new_[37409]_  = ~A170 & \new_[37408]_ ;
  assign \new_[37413]_  = ~A202 & ~A200;
  assign \new_[37414]_  = ~A166 & \new_[37413]_ ;
  assign \new_[37415]_  = \new_[37414]_  & \new_[37409]_ ;
  assign \new_[37419]_  = ~A233 & ~A232;
  assign \new_[37420]_  = ~A203 & \new_[37419]_ ;
  assign \new_[37423]_  = ~A266 & ~A265;
  assign \new_[37426]_  = A299 & ~A298;
  assign \new_[37427]_  = \new_[37426]_  & \new_[37423]_ ;
  assign \new_[37428]_  = \new_[37427]_  & \new_[37420]_ ;
  assign \new_[37432]_  = ~A167 & A169;
  assign \new_[37433]_  = ~A170 & \new_[37432]_ ;
  assign \new_[37437]_  = ~A201 & ~A200;
  assign \new_[37438]_  = ~A166 & \new_[37437]_ ;
  assign \new_[37439]_  = \new_[37438]_  & \new_[37433]_ ;
  assign \new_[37443]_  = A265 & A233;
  assign \new_[37444]_  = A232 & \new_[37443]_ ;
  assign \new_[37447]_  = ~A269 & ~A268;
  assign \new_[37450]_  = A299 & ~A298;
  assign \new_[37451]_  = \new_[37450]_  & \new_[37447]_ ;
  assign \new_[37452]_  = \new_[37451]_  & \new_[37444]_ ;
  assign \new_[37456]_  = ~A167 & A169;
  assign \new_[37457]_  = ~A170 & \new_[37456]_ ;
  assign \new_[37461]_  = ~A201 & ~A200;
  assign \new_[37462]_  = ~A166 & \new_[37461]_ ;
  assign \new_[37463]_  = \new_[37462]_  & \new_[37457]_ ;
  assign \new_[37467]_  = ~A236 & ~A235;
  assign \new_[37468]_  = ~A233 & \new_[37467]_ ;
  assign \new_[37471]_  = A266 & A265;
  assign \new_[37474]_  = A299 & ~A298;
  assign \new_[37475]_  = \new_[37474]_  & \new_[37471]_ ;
  assign \new_[37476]_  = \new_[37475]_  & \new_[37468]_ ;
  assign \new_[37480]_  = ~A167 & A169;
  assign \new_[37481]_  = ~A170 & \new_[37480]_ ;
  assign \new_[37485]_  = ~A201 & ~A200;
  assign \new_[37486]_  = ~A166 & \new_[37485]_ ;
  assign \new_[37487]_  = \new_[37486]_  & \new_[37481]_ ;
  assign \new_[37491]_  = ~A236 & ~A235;
  assign \new_[37492]_  = ~A233 & \new_[37491]_ ;
  assign \new_[37495]_  = ~A267 & ~A266;
  assign \new_[37498]_  = A299 & ~A298;
  assign \new_[37499]_  = \new_[37498]_  & \new_[37495]_ ;
  assign \new_[37500]_  = \new_[37499]_  & \new_[37492]_ ;
  assign \new_[37504]_  = ~A167 & A169;
  assign \new_[37505]_  = ~A170 & \new_[37504]_ ;
  assign \new_[37509]_  = ~A201 & ~A200;
  assign \new_[37510]_  = ~A166 & \new_[37509]_ ;
  assign \new_[37511]_  = \new_[37510]_  & \new_[37505]_ ;
  assign \new_[37515]_  = ~A236 & ~A235;
  assign \new_[37516]_  = ~A233 & \new_[37515]_ ;
  assign \new_[37519]_  = ~A266 & ~A265;
  assign \new_[37522]_  = A299 & ~A298;
  assign \new_[37523]_  = \new_[37522]_  & \new_[37519]_ ;
  assign \new_[37524]_  = \new_[37523]_  & \new_[37516]_ ;
  assign \new_[37528]_  = ~A167 & A169;
  assign \new_[37529]_  = ~A170 & \new_[37528]_ ;
  assign \new_[37533]_  = ~A201 & ~A200;
  assign \new_[37534]_  = ~A166 & \new_[37533]_ ;
  assign \new_[37535]_  = \new_[37534]_  & \new_[37529]_ ;
  assign \new_[37539]_  = ~A266 & ~A234;
  assign \new_[37540]_  = ~A233 & \new_[37539]_ ;
  assign \new_[37543]_  = ~A269 & ~A268;
  assign \new_[37546]_  = A299 & ~A298;
  assign \new_[37547]_  = \new_[37546]_  & \new_[37543]_ ;
  assign \new_[37548]_  = \new_[37547]_  & \new_[37540]_ ;
  assign \new_[37552]_  = ~A167 & A169;
  assign \new_[37553]_  = ~A170 & \new_[37552]_ ;
  assign \new_[37557]_  = ~A201 & ~A200;
  assign \new_[37558]_  = ~A166 & \new_[37557]_ ;
  assign \new_[37559]_  = \new_[37558]_  & \new_[37553]_ ;
  assign \new_[37563]_  = A234 & ~A233;
  assign \new_[37564]_  = A232 & \new_[37563]_ ;
  assign \new_[37567]_  = A298 & A235;
  assign \new_[37570]_  = ~A302 & ~A301;
  assign \new_[37571]_  = \new_[37570]_  & \new_[37567]_ ;
  assign \new_[37572]_  = \new_[37571]_  & \new_[37564]_ ;
  assign \new_[37576]_  = ~A167 & A169;
  assign \new_[37577]_  = ~A170 & \new_[37576]_ ;
  assign \new_[37581]_  = ~A201 & ~A200;
  assign \new_[37582]_  = ~A166 & \new_[37581]_ ;
  assign \new_[37583]_  = \new_[37582]_  & \new_[37577]_ ;
  assign \new_[37587]_  = A234 & ~A233;
  assign \new_[37588]_  = A232 & \new_[37587]_ ;
  assign \new_[37591]_  = A298 & A236;
  assign \new_[37594]_  = ~A302 & ~A301;
  assign \new_[37595]_  = \new_[37594]_  & \new_[37591]_ ;
  assign \new_[37596]_  = \new_[37595]_  & \new_[37588]_ ;
  assign \new_[37600]_  = ~A167 & A169;
  assign \new_[37601]_  = ~A170 & \new_[37600]_ ;
  assign \new_[37605]_  = ~A201 & ~A200;
  assign \new_[37606]_  = ~A166 & \new_[37605]_ ;
  assign \new_[37607]_  = \new_[37606]_  & \new_[37601]_ ;
  assign \new_[37611]_  = ~A266 & ~A233;
  assign \new_[37612]_  = ~A232 & \new_[37611]_ ;
  assign \new_[37615]_  = ~A269 & ~A268;
  assign \new_[37618]_  = A299 & ~A298;
  assign \new_[37619]_  = \new_[37618]_  & \new_[37615]_ ;
  assign \new_[37620]_  = \new_[37619]_  & \new_[37612]_ ;
  assign \new_[37624]_  = ~A167 & A169;
  assign \new_[37625]_  = ~A170 & \new_[37624]_ ;
  assign \new_[37629]_  = ~A200 & ~A199;
  assign \new_[37630]_  = ~A166 & \new_[37629]_ ;
  assign \new_[37631]_  = \new_[37630]_  & \new_[37625]_ ;
  assign \new_[37635]_  = A265 & A233;
  assign \new_[37636]_  = A232 & \new_[37635]_ ;
  assign \new_[37639]_  = ~A269 & ~A268;
  assign \new_[37642]_  = A299 & ~A298;
  assign \new_[37643]_  = \new_[37642]_  & \new_[37639]_ ;
  assign \new_[37644]_  = \new_[37643]_  & \new_[37636]_ ;
  assign \new_[37648]_  = ~A167 & A169;
  assign \new_[37649]_  = ~A170 & \new_[37648]_ ;
  assign \new_[37653]_  = ~A200 & ~A199;
  assign \new_[37654]_  = ~A166 & \new_[37653]_ ;
  assign \new_[37655]_  = \new_[37654]_  & \new_[37649]_ ;
  assign \new_[37659]_  = ~A236 & ~A235;
  assign \new_[37660]_  = ~A233 & \new_[37659]_ ;
  assign \new_[37663]_  = A266 & A265;
  assign \new_[37666]_  = A299 & ~A298;
  assign \new_[37667]_  = \new_[37666]_  & \new_[37663]_ ;
  assign \new_[37668]_  = \new_[37667]_  & \new_[37660]_ ;
  assign \new_[37672]_  = ~A167 & A169;
  assign \new_[37673]_  = ~A170 & \new_[37672]_ ;
  assign \new_[37677]_  = ~A200 & ~A199;
  assign \new_[37678]_  = ~A166 & \new_[37677]_ ;
  assign \new_[37679]_  = \new_[37678]_  & \new_[37673]_ ;
  assign \new_[37683]_  = ~A236 & ~A235;
  assign \new_[37684]_  = ~A233 & \new_[37683]_ ;
  assign \new_[37687]_  = ~A267 & ~A266;
  assign \new_[37690]_  = A299 & ~A298;
  assign \new_[37691]_  = \new_[37690]_  & \new_[37687]_ ;
  assign \new_[37692]_  = \new_[37691]_  & \new_[37684]_ ;
  assign \new_[37696]_  = ~A167 & A169;
  assign \new_[37697]_  = ~A170 & \new_[37696]_ ;
  assign \new_[37701]_  = ~A200 & ~A199;
  assign \new_[37702]_  = ~A166 & \new_[37701]_ ;
  assign \new_[37703]_  = \new_[37702]_  & \new_[37697]_ ;
  assign \new_[37707]_  = ~A236 & ~A235;
  assign \new_[37708]_  = ~A233 & \new_[37707]_ ;
  assign \new_[37711]_  = ~A266 & ~A265;
  assign \new_[37714]_  = A299 & ~A298;
  assign \new_[37715]_  = \new_[37714]_  & \new_[37711]_ ;
  assign \new_[37716]_  = \new_[37715]_  & \new_[37708]_ ;
  assign \new_[37720]_  = ~A167 & A169;
  assign \new_[37721]_  = ~A170 & \new_[37720]_ ;
  assign \new_[37725]_  = ~A200 & ~A199;
  assign \new_[37726]_  = ~A166 & \new_[37725]_ ;
  assign \new_[37727]_  = \new_[37726]_  & \new_[37721]_ ;
  assign \new_[37731]_  = ~A266 & ~A234;
  assign \new_[37732]_  = ~A233 & \new_[37731]_ ;
  assign \new_[37735]_  = ~A269 & ~A268;
  assign \new_[37738]_  = A299 & ~A298;
  assign \new_[37739]_  = \new_[37738]_  & \new_[37735]_ ;
  assign \new_[37740]_  = \new_[37739]_  & \new_[37732]_ ;
  assign \new_[37744]_  = ~A167 & A169;
  assign \new_[37745]_  = ~A170 & \new_[37744]_ ;
  assign \new_[37749]_  = ~A200 & ~A199;
  assign \new_[37750]_  = ~A166 & \new_[37749]_ ;
  assign \new_[37751]_  = \new_[37750]_  & \new_[37745]_ ;
  assign \new_[37755]_  = A234 & ~A233;
  assign \new_[37756]_  = A232 & \new_[37755]_ ;
  assign \new_[37759]_  = A298 & A235;
  assign \new_[37762]_  = ~A302 & ~A301;
  assign \new_[37763]_  = \new_[37762]_  & \new_[37759]_ ;
  assign \new_[37764]_  = \new_[37763]_  & \new_[37756]_ ;
  assign \new_[37768]_  = ~A167 & A169;
  assign \new_[37769]_  = ~A170 & \new_[37768]_ ;
  assign \new_[37773]_  = ~A200 & ~A199;
  assign \new_[37774]_  = ~A166 & \new_[37773]_ ;
  assign \new_[37775]_  = \new_[37774]_  & \new_[37769]_ ;
  assign \new_[37779]_  = A234 & ~A233;
  assign \new_[37780]_  = A232 & \new_[37779]_ ;
  assign \new_[37783]_  = A298 & A236;
  assign \new_[37786]_  = ~A302 & ~A301;
  assign \new_[37787]_  = \new_[37786]_  & \new_[37783]_ ;
  assign \new_[37788]_  = \new_[37787]_  & \new_[37780]_ ;
  assign \new_[37792]_  = ~A167 & A169;
  assign \new_[37793]_  = ~A170 & \new_[37792]_ ;
  assign \new_[37797]_  = ~A200 & ~A199;
  assign \new_[37798]_  = ~A166 & \new_[37797]_ ;
  assign \new_[37799]_  = \new_[37798]_  & \new_[37793]_ ;
  assign \new_[37803]_  = ~A266 & ~A233;
  assign \new_[37804]_  = ~A232 & \new_[37803]_ ;
  assign \new_[37807]_  = ~A269 & ~A268;
  assign \new_[37810]_  = A299 & ~A298;
  assign \new_[37811]_  = \new_[37810]_  & \new_[37807]_ ;
  assign \new_[37812]_  = \new_[37811]_  & \new_[37804]_ ;
  assign \new_[37816]_  = ~A166 & ~A167;
  assign \new_[37817]_  = ~A169 & \new_[37816]_ ;
  assign \new_[37821]_  = A232 & A200;
  assign \new_[37822]_  = ~A199 & \new_[37821]_ ;
  assign \new_[37823]_  = \new_[37822]_  & \new_[37817]_ ;
  assign \new_[37827]_  = ~A267 & A265;
  assign \new_[37828]_  = A233 & \new_[37827]_ ;
  assign \new_[37831]_  = ~A299 & A298;
  assign \new_[37834]_  = A301 & A300;
  assign \new_[37835]_  = \new_[37834]_  & \new_[37831]_ ;
  assign \new_[37836]_  = \new_[37835]_  & \new_[37828]_ ;
  assign \new_[37840]_  = ~A166 & ~A167;
  assign \new_[37841]_  = ~A169 & \new_[37840]_ ;
  assign \new_[37845]_  = A232 & A200;
  assign \new_[37846]_  = ~A199 & \new_[37845]_ ;
  assign \new_[37847]_  = \new_[37846]_  & \new_[37841]_ ;
  assign \new_[37851]_  = ~A267 & A265;
  assign \new_[37852]_  = A233 & \new_[37851]_ ;
  assign \new_[37855]_  = ~A299 & A298;
  assign \new_[37858]_  = A302 & A300;
  assign \new_[37859]_  = \new_[37858]_  & \new_[37855]_ ;
  assign \new_[37860]_  = \new_[37859]_  & \new_[37852]_ ;
  assign \new_[37864]_  = ~A166 & ~A167;
  assign \new_[37865]_  = ~A169 & \new_[37864]_ ;
  assign \new_[37869]_  = A232 & A200;
  assign \new_[37870]_  = ~A199 & \new_[37869]_ ;
  assign \new_[37871]_  = \new_[37870]_  & \new_[37865]_ ;
  assign \new_[37875]_  = A266 & A265;
  assign \new_[37876]_  = A233 & \new_[37875]_ ;
  assign \new_[37879]_  = ~A299 & A298;
  assign \new_[37882]_  = A301 & A300;
  assign \new_[37883]_  = \new_[37882]_  & \new_[37879]_ ;
  assign \new_[37884]_  = \new_[37883]_  & \new_[37876]_ ;
  assign \new_[37888]_  = ~A166 & ~A167;
  assign \new_[37889]_  = ~A169 & \new_[37888]_ ;
  assign \new_[37893]_  = A232 & A200;
  assign \new_[37894]_  = ~A199 & \new_[37893]_ ;
  assign \new_[37895]_  = \new_[37894]_  & \new_[37889]_ ;
  assign \new_[37899]_  = A266 & A265;
  assign \new_[37900]_  = A233 & \new_[37899]_ ;
  assign \new_[37903]_  = ~A299 & A298;
  assign \new_[37906]_  = A302 & A300;
  assign \new_[37907]_  = \new_[37906]_  & \new_[37903]_ ;
  assign \new_[37908]_  = \new_[37907]_  & \new_[37900]_ ;
  assign \new_[37912]_  = ~A166 & ~A167;
  assign \new_[37913]_  = ~A169 & \new_[37912]_ ;
  assign \new_[37917]_  = A232 & A200;
  assign \new_[37918]_  = ~A199 & \new_[37917]_ ;
  assign \new_[37919]_  = \new_[37918]_  & \new_[37913]_ ;
  assign \new_[37923]_  = ~A266 & ~A265;
  assign \new_[37924]_  = A233 & \new_[37923]_ ;
  assign \new_[37927]_  = ~A299 & A298;
  assign \new_[37930]_  = A301 & A300;
  assign \new_[37931]_  = \new_[37930]_  & \new_[37927]_ ;
  assign \new_[37932]_  = \new_[37931]_  & \new_[37924]_ ;
  assign \new_[37936]_  = ~A166 & ~A167;
  assign \new_[37937]_  = ~A169 & \new_[37936]_ ;
  assign \new_[37941]_  = A232 & A200;
  assign \new_[37942]_  = ~A199 & \new_[37941]_ ;
  assign \new_[37943]_  = \new_[37942]_  & \new_[37937]_ ;
  assign \new_[37947]_  = ~A266 & ~A265;
  assign \new_[37948]_  = A233 & \new_[37947]_ ;
  assign \new_[37951]_  = ~A299 & A298;
  assign \new_[37954]_  = A302 & A300;
  assign \new_[37955]_  = \new_[37954]_  & \new_[37951]_ ;
  assign \new_[37956]_  = \new_[37955]_  & \new_[37948]_ ;
  assign \new_[37960]_  = ~A166 & ~A167;
  assign \new_[37961]_  = ~A169 & \new_[37960]_ ;
  assign \new_[37965]_  = ~A233 & A200;
  assign \new_[37966]_  = ~A199 & \new_[37965]_ ;
  assign \new_[37967]_  = \new_[37966]_  & \new_[37961]_ ;
  assign \new_[37971]_  = ~A266 & ~A236;
  assign \new_[37972]_  = ~A235 & \new_[37971]_ ;
  assign \new_[37975]_  = ~A269 & ~A268;
  assign \new_[37978]_  = A299 & ~A298;
  assign \new_[37979]_  = \new_[37978]_  & \new_[37975]_ ;
  assign \new_[37980]_  = \new_[37979]_  & \new_[37972]_ ;
  assign \new_[37984]_  = ~A166 & ~A167;
  assign \new_[37985]_  = ~A169 & \new_[37984]_ ;
  assign \new_[37989]_  = ~A233 & A200;
  assign \new_[37990]_  = ~A199 & \new_[37989]_ ;
  assign \new_[37991]_  = \new_[37990]_  & \new_[37985]_ ;
  assign \new_[37995]_  = A266 & A265;
  assign \new_[37996]_  = ~A234 & \new_[37995]_ ;
  assign \new_[37999]_  = ~A299 & A298;
  assign \new_[38002]_  = A301 & A300;
  assign \new_[38003]_  = \new_[38002]_  & \new_[37999]_ ;
  assign \new_[38004]_  = \new_[38003]_  & \new_[37996]_ ;
  assign \new_[38008]_  = ~A166 & ~A167;
  assign \new_[38009]_  = ~A169 & \new_[38008]_ ;
  assign \new_[38013]_  = ~A233 & A200;
  assign \new_[38014]_  = ~A199 & \new_[38013]_ ;
  assign \new_[38015]_  = \new_[38014]_  & \new_[38009]_ ;
  assign \new_[38019]_  = A266 & A265;
  assign \new_[38020]_  = ~A234 & \new_[38019]_ ;
  assign \new_[38023]_  = ~A299 & A298;
  assign \new_[38026]_  = A302 & A300;
  assign \new_[38027]_  = \new_[38026]_  & \new_[38023]_ ;
  assign \new_[38028]_  = \new_[38027]_  & \new_[38020]_ ;
  assign \new_[38032]_  = ~A166 & ~A167;
  assign \new_[38033]_  = ~A169 & \new_[38032]_ ;
  assign \new_[38037]_  = ~A233 & A200;
  assign \new_[38038]_  = ~A199 & \new_[38037]_ ;
  assign \new_[38039]_  = \new_[38038]_  & \new_[38033]_ ;
  assign \new_[38043]_  = ~A267 & ~A266;
  assign \new_[38044]_  = ~A234 & \new_[38043]_ ;
  assign \new_[38047]_  = ~A299 & A298;
  assign \new_[38050]_  = A301 & A300;
  assign \new_[38051]_  = \new_[38050]_  & \new_[38047]_ ;
  assign \new_[38052]_  = \new_[38051]_  & \new_[38044]_ ;
  assign \new_[38056]_  = ~A166 & ~A167;
  assign \new_[38057]_  = ~A169 & \new_[38056]_ ;
  assign \new_[38061]_  = ~A233 & A200;
  assign \new_[38062]_  = ~A199 & \new_[38061]_ ;
  assign \new_[38063]_  = \new_[38062]_  & \new_[38057]_ ;
  assign \new_[38067]_  = ~A267 & ~A266;
  assign \new_[38068]_  = ~A234 & \new_[38067]_ ;
  assign \new_[38071]_  = ~A299 & A298;
  assign \new_[38074]_  = A302 & A300;
  assign \new_[38075]_  = \new_[38074]_  & \new_[38071]_ ;
  assign \new_[38076]_  = \new_[38075]_  & \new_[38068]_ ;
  assign \new_[38080]_  = ~A166 & ~A167;
  assign \new_[38081]_  = ~A169 & \new_[38080]_ ;
  assign \new_[38085]_  = ~A233 & A200;
  assign \new_[38086]_  = ~A199 & \new_[38085]_ ;
  assign \new_[38087]_  = \new_[38086]_  & \new_[38081]_ ;
  assign \new_[38091]_  = ~A266 & ~A265;
  assign \new_[38092]_  = ~A234 & \new_[38091]_ ;
  assign \new_[38095]_  = ~A299 & A298;
  assign \new_[38098]_  = A301 & A300;
  assign \new_[38099]_  = \new_[38098]_  & \new_[38095]_ ;
  assign \new_[38100]_  = \new_[38099]_  & \new_[38092]_ ;
  assign \new_[38104]_  = ~A166 & ~A167;
  assign \new_[38105]_  = ~A169 & \new_[38104]_ ;
  assign \new_[38109]_  = ~A233 & A200;
  assign \new_[38110]_  = ~A199 & \new_[38109]_ ;
  assign \new_[38111]_  = \new_[38110]_  & \new_[38105]_ ;
  assign \new_[38115]_  = ~A266 & ~A265;
  assign \new_[38116]_  = ~A234 & \new_[38115]_ ;
  assign \new_[38119]_  = ~A299 & A298;
  assign \new_[38122]_  = A302 & A300;
  assign \new_[38123]_  = \new_[38122]_  & \new_[38119]_ ;
  assign \new_[38124]_  = \new_[38123]_  & \new_[38116]_ ;
  assign \new_[38128]_  = ~A166 & ~A167;
  assign \new_[38129]_  = ~A169 & \new_[38128]_ ;
  assign \new_[38133]_  = A232 & A200;
  assign \new_[38134]_  = ~A199 & \new_[38133]_ ;
  assign \new_[38135]_  = \new_[38134]_  & \new_[38129]_ ;
  assign \new_[38139]_  = A235 & A234;
  assign \new_[38140]_  = ~A233 & \new_[38139]_ ;
  assign \new_[38143]_  = ~A266 & A265;
  assign \new_[38146]_  = A268 & A267;
  assign \new_[38147]_  = \new_[38146]_  & \new_[38143]_ ;
  assign \new_[38148]_  = \new_[38147]_  & \new_[38140]_ ;
  assign \new_[38152]_  = ~A166 & ~A167;
  assign \new_[38153]_  = ~A169 & \new_[38152]_ ;
  assign \new_[38157]_  = A232 & A200;
  assign \new_[38158]_  = ~A199 & \new_[38157]_ ;
  assign \new_[38159]_  = \new_[38158]_  & \new_[38153]_ ;
  assign \new_[38163]_  = A235 & A234;
  assign \new_[38164]_  = ~A233 & \new_[38163]_ ;
  assign \new_[38167]_  = ~A266 & A265;
  assign \new_[38170]_  = A269 & A267;
  assign \new_[38171]_  = \new_[38170]_  & \new_[38167]_ ;
  assign \new_[38172]_  = \new_[38171]_  & \new_[38164]_ ;
  assign \new_[38176]_  = ~A166 & ~A167;
  assign \new_[38177]_  = ~A169 & \new_[38176]_ ;
  assign \new_[38181]_  = A232 & A200;
  assign \new_[38182]_  = ~A199 & \new_[38181]_ ;
  assign \new_[38183]_  = \new_[38182]_  & \new_[38177]_ ;
  assign \new_[38187]_  = A236 & A234;
  assign \new_[38188]_  = ~A233 & \new_[38187]_ ;
  assign \new_[38191]_  = ~A266 & A265;
  assign \new_[38194]_  = A268 & A267;
  assign \new_[38195]_  = \new_[38194]_  & \new_[38191]_ ;
  assign \new_[38196]_  = \new_[38195]_  & \new_[38188]_ ;
  assign \new_[38200]_  = ~A166 & ~A167;
  assign \new_[38201]_  = ~A169 & \new_[38200]_ ;
  assign \new_[38205]_  = A232 & A200;
  assign \new_[38206]_  = ~A199 & \new_[38205]_ ;
  assign \new_[38207]_  = \new_[38206]_  & \new_[38201]_ ;
  assign \new_[38211]_  = A236 & A234;
  assign \new_[38212]_  = ~A233 & \new_[38211]_ ;
  assign \new_[38215]_  = ~A266 & A265;
  assign \new_[38218]_  = A269 & A267;
  assign \new_[38219]_  = \new_[38218]_  & \new_[38215]_ ;
  assign \new_[38220]_  = \new_[38219]_  & \new_[38212]_ ;
  assign \new_[38224]_  = ~A166 & ~A167;
  assign \new_[38225]_  = ~A169 & \new_[38224]_ ;
  assign \new_[38229]_  = ~A232 & A200;
  assign \new_[38230]_  = ~A199 & \new_[38229]_ ;
  assign \new_[38231]_  = \new_[38230]_  & \new_[38225]_ ;
  assign \new_[38235]_  = A266 & A265;
  assign \new_[38236]_  = ~A233 & \new_[38235]_ ;
  assign \new_[38239]_  = ~A299 & A298;
  assign \new_[38242]_  = A301 & A300;
  assign \new_[38243]_  = \new_[38242]_  & \new_[38239]_ ;
  assign \new_[38244]_  = \new_[38243]_  & \new_[38236]_ ;
  assign \new_[38248]_  = ~A166 & ~A167;
  assign \new_[38249]_  = ~A169 & \new_[38248]_ ;
  assign \new_[38253]_  = ~A232 & A200;
  assign \new_[38254]_  = ~A199 & \new_[38253]_ ;
  assign \new_[38255]_  = \new_[38254]_  & \new_[38249]_ ;
  assign \new_[38259]_  = A266 & A265;
  assign \new_[38260]_  = ~A233 & \new_[38259]_ ;
  assign \new_[38263]_  = ~A299 & A298;
  assign \new_[38266]_  = A302 & A300;
  assign \new_[38267]_  = \new_[38266]_  & \new_[38263]_ ;
  assign \new_[38268]_  = \new_[38267]_  & \new_[38260]_ ;
  assign \new_[38272]_  = ~A166 & ~A167;
  assign \new_[38273]_  = ~A169 & \new_[38272]_ ;
  assign \new_[38277]_  = ~A232 & A200;
  assign \new_[38278]_  = ~A199 & \new_[38277]_ ;
  assign \new_[38279]_  = \new_[38278]_  & \new_[38273]_ ;
  assign \new_[38283]_  = ~A267 & ~A266;
  assign \new_[38284]_  = ~A233 & \new_[38283]_ ;
  assign \new_[38287]_  = ~A299 & A298;
  assign \new_[38290]_  = A301 & A300;
  assign \new_[38291]_  = \new_[38290]_  & \new_[38287]_ ;
  assign \new_[38292]_  = \new_[38291]_  & \new_[38284]_ ;
  assign \new_[38296]_  = ~A166 & ~A167;
  assign \new_[38297]_  = ~A169 & \new_[38296]_ ;
  assign \new_[38301]_  = ~A232 & A200;
  assign \new_[38302]_  = ~A199 & \new_[38301]_ ;
  assign \new_[38303]_  = \new_[38302]_  & \new_[38297]_ ;
  assign \new_[38307]_  = ~A267 & ~A266;
  assign \new_[38308]_  = ~A233 & \new_[38307]_ ;
  assign \new_[38311]_  = ~A299 & A298;
  assign \new_[38314]_  = A302 & A300;
  assign \new_[38315]_  = \new_[38314]_  & \new_[38311]_ ;
  assign \new_[38316]_  = \new_[38315]_  & \new_[38308]_ ;
  assign \new_[38320]_  = ~A166 & ~A167;
  assign \new_[38321]_  = ~A169 & \new_[38320]_ ;
  assign \new_[38325]_  = ~A232 & A200;
  assign \new_[38326]_  = ~A199 & \new_[38325]_ ;
  assign \new_[38327]_  = \new_[38326]_  & \new_[38321]_ ;
  assign \new_[38331]_  = ~A266 & ~A265;
  assign \new_[38332]_  = ~A233 & \new_[38331]_ ;
  assign \new_[38335]_  = ~A299 & A298;
  assign \new_[38338]_  = A301 & A300;
  assign \new_[38339]_  = \new_[38338]_  & \new_[38335]_ ;
  assign \new_[38340]_  = \new_[38339]_  & \new_[38332]_ ;
  assign \new_[38344]_  = ~A166 & ~A167;
  assign \new_[38345]_  = ~A169 & \new_[38344]_ ;
  assign \new_[38349]_  = ~A232 & A200;
  assign \new_[38350]_  = ~A199 & \new_[38349]_ ;
  assign \new_[38351]_  = \new_[38350]_  & \new_[38345]_ ;
  assign \new_[38355]_  = ~A266 & ~A265;
  assign \new_[38356]_  = ~A233 & \new_[38355]_ ;
  assign \new_[38359]_  = ~A299 & A298;
  assign \new_[38362]_  = A302 & A300;
  assign \new_[38363]_  = \new_[38362]_  & \new_[38359]_ ;
  assign \new_[38364]_  = \new_[38363]_  & \new_[38356]_ ;
  assign \new_[38368]_  = ~A166 & ~A167;
  assign \new_[38369]_  = ~A169 & \new_[38368]_ ;
  assign \new_[38373]_  = A201 & ~A200;
  assign \new_[38374]_  = A199 & \new_[38373]_ ;
  assign \new_[38375]_  = \new_[38374]_  & \new_[38369]_ ;
  assign \new_[38379]_  = A233 & A232;
  assign \new_[38380]_  = A202 & \new_[38379]_ ;
  assign \new_[38383]_  = ~A267 & A265;
  assign \new_[38386]_  = A299 & ~A298;
  assign \new_[38387]_  = \new_[38386]_  & \new_[38383]_ ;
  assign \new_[38388]_  = \new_[38387]_  & \new_[38380]_ ;
  assign \new_[38392]_  = ~A166 & ~A167;
  assign \new_[38393]_  = ~A169 & \new_[38392]_ ;
  assign \new_[38397]_  = A201 & ~A200;
  assign \new_[38398]_  = A199 & \new_[38397]_ ;
  assign \new_[38399]_  = \new_[38398]_  & \new_[38393]_ ;
  assign \new_[38403]_  = A233 & A232;
  assign \new_[38404]_  = A202 & \new_[38403]_ ;
  assign \new_[38407]_  = A266 & A265;
  assign \new_[38410]_  = A299 & ~A298;
  assign \new_[38411]_  = \new_[38410]_  & \new_[38407]_ ;
  assign \new_[38412]_  = \new_[38411]_  & \new_[38404]_ ;
  assign \new_[38416]_  = ~A166 & ~A167;
  assign \new_[38417]_  = ~A169 & \new_[38416]_ ;
  assign \new_[38421]_  = A201 & ~A200;
  assign \new_[38422]_  = A199 & \new_[38421]_ ;
  assign \new_[38423]_  = \new_[38422]_  & \new_[38417]_ ;
  assign \new_[38427]_  = A233 & A232;
  assign \new_[38428]_  = A202 & \new_[38427]_ ;
  assign \new_[38431]_  = ~A266 & ~A265;
  assign \new_[38434]_  = A299 & ~A298;
  assign \new_[38435]_  = \new_[38434]_  & \new_[38431]_ ;
  assign \new_[38436]_  = \new_[38435]_  & \new_[38428]_ ;
  assign \new_[38440]_  = ~A166 & ~A167;
  assign \new_[38441]_  = ~A169 & \new_[38440]_ ;
  assign \new_[38445]_  = A201 & ~A200;
  assign \new_[38446]_  = A199 & \new_[38445]_ ;
  assign \new_[38447]_  = \new_[38446]_  & \new_[38441]_ ;
  assign \new_[38451]_  = A233 & ~A232;
  assign \new_[38452]_  = A202 & \new_[38451]_ ;
  assign \new_[38455]_  = ~A266 & A265;
  assign \new_[38458]_  = A268 & A267;
  assign \new_[38459]_  = \new_[38458]_  & \new_[38455]_ ;
  assign \new_[38460]_  = \new_[38459]_  & \new_[38452]_ ;
  assign \new_[38464]_  = ~A166 & ~A167;
  assign \new_[38465]_  = ~A169 & \new_[38464]_ ;
  assign \new_[38469]_  = A201 & ~A200;
  assign \new_[38470]_  = A199 & \new_[38469]_ ;
  assign \new_[38471]_  = \new_[38470]_  & \new_[38465]_ ;
  assign \new_[38475]_  = A233 & ~A232;
  assign \new_[38476]_  = A202 & \new_[38475]_ ;
  assign \new_[38479]_  = ~A266 & A265;
  assign \new_[38482]_  = A269 & A267;
  assign \new_[38483]_  = \new_[38482]_  & \new_[38479]_ ;
  assign \new_[38484]_  = \new_[38483]_  & \new_[38476]_ ;
  assign \new_[38488]_  = ~A166 & ~A167;
  assign \new_[38489]_  = ~A169 & \new_[38488]_ ;
  assign \new_[38493]_  = A201 & ~A200;
  assign \new_[38494]_  = A199 & \new_[38493]_ ;
  assign \new_[38495]_  = \new_[38494]_  & \new_[38489]_ ;
  assign \new_[38499]_  = ~A234 & ~A233;
  assign \new_[38500]_  = A202 & \new_[38499]_ ;
  assign \new_[38503]_  = A266 & A265;
  assign \new_[38506]_  = A299 & ~A298;
  assign \new_[38507]_  = \new_[38506]_  & \new_[38503]_ ;
  assign \new_[38508]_  = \new_[38507]_  & \new_[38500]_ ;
  assign \new_[38512]_  = ~A166 & ~A167;
  assign \new_[38513]_  = ~A169 & \new_[38512]_ ;
  assign \new_[38517]_  = A201 & ~A200;
  assign \new_[38518]_  = A199 & \new_[38517]_ ;
  assign \new_[38519]_  = \new_[38518]_  & \new_[38513]_ ;
  assign \new_[38523]_  = ~A234 & ~A233;
  assign \new_[38524]_  = A202 & \new_[38523]_ ;
  assign \new_[38527]_  = ~A267 & ~A266;
  assign \new_[38530]_  = A299 & ~A298;
  assign \new_[38531]_  = \new_[38530]_  & \new_[38527]_ ;
  assign \new_[38532]_  = \new_[38531]_  & \new_[38524]_ ;
  assign \new_[38536]_  = ~A166 & ~A167;
  assign \new_[38537]_  = ~A169 & \new_[38536]_ ;
  assign \new_[38541]_  = A201 & ~A200;
  assign \new_[38542]_  = A199 & \new_[38541]_ ;
  assign \new_[38543]_  = \new_[38542]_  & \new_[38537]_ ;
  assign \new_[38547]_  = ~A234 & ~A233;
  assign \new_[38548]_  = A202 & \new_[38547]_ ;
  assign \new_[38551]_  = ~A266 & ~A265;
  assign \new_[38554]_  = A299 & ~A298;
  assign \new_[38555]_  = \new_[38554]_  & \new_[38551]_ ;
  assign \new_[38556]_  = \new_[38555]_  & \new_[38548]_ ;
  assign \new_[38560]_  = ~A166 & ~A167;
  assign \new_[38561]_  = ~A169 & \new_[38560]_ ;
  assign \new_[38565]_  = A201 & ~A200;
  assign \new_[38566]_  = A199 & \new_[38565]_ ;
  assign \new_[38567]_  = \new_[38566]_  & \new_[38561]_ ;
  assign \new_[38571]_  = ~A233 & A232;
  assign \new_[38572]_  = A202 & \new_[38571]_ ;
  assign \new_[38575]_  = A235 & A234;
  assign \new_[38578]_  = ~A300 & A298;
  assign \new_[38579]_  = \new_[38578]_  & \new_[38575]_ ;
  assign \new_[38580]_  = \new_[38579]_  & \new_[38572]_ ;
  assign \new_[38584]_  = ~A166 & ~A167;
  assign \new_[38585]_  = ~A169 & \new_[38584]_ ;
  assign \new_[38589]_  = A201 & ~A200;
  assign \new_[38590]_  = A199 & \new_[38589]_ ;
  assign \new_[38591]_  = \new_[38590]_  & \new_[38585]_ ;
  assign \new_[38595]_  = ~A233 & A232;
  assign \new_[38596]_  = A202 & \new_[38595]_ ;
  assign \new_[38599]_  = A235 & A234;
  assign \new_[38602]_  = A299 & A298;
  assign \new_[38603]_  = \new_[38602]_  & \new_[38599]_ ;
  assign \new_[38604]_  = \new_[38603]_  & \new_[38596]_ ;
  assign \new_[38608]_  = ~A166 & ~A167;
  assign \new_[38609]_  = ~A169 & \new_[38608]_ ;
  assign \new_[38613]_  = A201 & ~A200;
  assign \new_[38614]_  = A199 & \new_[38613]_ ;
  assign \new_[38615]_  = \new_[38614]_  & \new_[38609]_ ;
  assign \new_[38619]_  = ~A233 & A232;
  assign \new_[38620]_  = A202 & \new_[38619]_ ;
  assign \new_[38623]_  = A235 & A234;
  assign \new_[38626]_  = ~A299 & ~A298;
  assign \new_[38627]_  = \new_[38626]_  & \new_[38623]_ ;
  assign \new_[38628]_  = \new_[38627]_  & \new_[38620]_ ;
  assign \new_[38632]_  = ~A166 & ~A167;
  assign \new_[38633]_  = ~A169 & \new_[38632]_ ;
  assign \new_[38637]_  = A201 & ~A200;
  assign \new_[38638]_  = A199 & \new_[38637]_ ;
  assign \new_[38639]_  = \new_[38638]_  & \new_[38633]_ ;
  assign \new_[38643]_  = ~A233 & A232;
  assign \new_[38644]_  = A202 & \new_[38643]_ ;
  assign \new_[38647]_  = A235 & A234;
  assign \new_[38650]_  = A266 & ~A265;
  assign \new_[38651]_  = \new_[38650]_  & \new_[38647]_ ;
  assign \new_[38652]_  = \new_[38651]_  & \new_[38644]_ ;
  assign \new_[38656]_  = ~A166 & ~A167;
  assign \new_[38657]_  = ~A169 & \new_[38656]_ ;
  assign \new_[38661]_  = A201 & ~A200;
  assign \new_[38662]_  = A199 & \new_[38661]_ ;
  assign \new_[38663]_  = \new_[38662]_  & \new_[38657]_ ;
  assign \new_[38667]_  = ~A233 & A232;
  assign \new_[38668]_  = A202 & \new_[38667]_ ;
  assign \new_[38671]_  = A236 & A234;
  assign \new_[38674]_  = ~A300 & A298;
  assign \new_[38675]_  = \new_[38674]_  & \new_[38671]_ ;
  assign \new_[38676]_  = \new_[38675]_  & \new_[38668]_ ;
  assign \new_[38680]_  = ~A166 & ~A167;
  assign \new_[38681]_  = ~A169 & \new_[38680]_ ;
  assign \new_[38685]_  = A201 & ~A200;
  assign \new_[38686]_  = A199 & \new_[38685]_ ;
  assign \new_[38687]_  = \new_[38686]_  & \new_[38681]_ ;
  assign \new_[38691]_  = ~A233 & A232;
  assign \new_[38692]_  = A202 & \new_[38691]_ ;
  assign \new_[38695]_  = A236 & A234;
  assign \new_[38698]_  = A299 & A298;
  assign \new_[38699]_  = \new_[38698]_  & \new_[38695]_ ;
  assign \new_[38700]_  = \new_[38699]_  & \new_[38692]_ ;
  assign \new_[38704]_  = ~A166 & ~A167;
  assign \new_[38705]_  = ~A169 & \new_[38704]_ ;
  assign \new_[38709]_  = A201 & ~A200;
  assign \new_[38710]_  = A199 & \new_[38709]_ ;
  assign \new_[38711]_  = \new_[38710]_  & \new_[38705]_ ;
  assign \new_[38715]_  = ~A233 & A232;
  assign \new_[38716]_  = A202 & \new_[38715]_ ;
  assign \new_[38719]_  = A236 & A234;
  assign \new_[38722]_  = ~A299 & ~A298;
  assign \new_[38723]_  = \new_[38722]_  & \new_[38719]_ ;
  assign \new_[38724]_  = \new_[38723]_  & \new_[38716]_ ;
  assign \new_[38728]_  = ~A166 & ~A167;
  assign \new_[38729]_  = ~A169 & \new_[38728]_ ;
  assign \new_[38733]_  = A201 & ~A200;
  assign \new_[38734]_  = A199 & \new_[38733]_ ;
  assign \new_[38735]_  = \new_[38734]_  & \new_[38729]_ ;
  assign \new_[38739]_  = ~A233 & A232;
  assign \new_[38740]_  = A202 & \new_[38739]_ ;
  assign \new_[38743]_  = A236 & A234;
  assign \new_[38746]_  = A266 & ~A265;
  assign \new_[38747]_  = \new_[38746]_  & \new_[38743]_ ;
  assign \new_[38748]_  = \new_[38747]_  & \new_[38740]_ ;
  assign \new_[38752]_  = ~A166 & ~A167;
  assign \new_[38753]_  = ~A169 & \new_[38752]_ ;
  assign \new_[38757]_  = A201 & ~A200;
  assign \new_[38758]_  = A199 & \new_[38757]_ ;
  assign \new_[38759]_  = \new_[38758]_  & \new_[38753]_ ;
  assign \new_[38763]_  = ~A233 & ~A232;
  assign \new_[38764]_  = A202 & \new_[38763]_ ;
  assign \new_[38767]_  = A266 & A265;
  assign \new_[38770]_  = A299 & ~A298;
  assign \new_[38771]_  = \new_[38770]_  & \new_[38767]_ ;
  assign \new_[38772]_  = \new_[38771]_  & \new_[38764]_ ;
  assign \new_[38776]_  = ~A166 & ~A167;
  assign \new_[38777]_  = ~A169 & \new_[38776]_ ;
  assign \new_[38781]_  = A201 & ~A200;
  assign \new_[38782]_  = A199 & \new_[38781]_ ;
  assign \new_[38783]_  = \new_[38782]_  & \new_[38777]_ ;
  assign \new_[38787]_  = ~A233 & ~A232;
  assign \new_[38788]_  = A202 & \new_[38787]_ ;
  assign \new_[38791]_  = ~A267 & ~A266;
  assign \new_[38794]_  = A299 & ~A298;
  assign \new_[38795]_  = \new_[38794]_  & \new_[38791]_ ;
  assign \new_[38796]_  = \new_[38795]_  & \new_[38788]_ ;
  assign \new_[38800]_  = ~A166 & ~A167;
  assign \new_[38801]_  = ~A169 & \new_[38800]_ ;
  assign \new_[38805]_  = A201 & ~A200;
  assign \new_[38806]_  = A199 & \new_[38805]_ ;
  assign \new_[38807]_  = \new_[38806]_  & \new_[38801]_ ;
  assign \new_[38811]_  = ~A233 & ~A232;
  assign \new_[38812]_  = A202 & \new_[38811]_ ;
  assign \new_[38815]_  = ~A266 & ~A265;
  assign \new_[38818]_  = A299 & ~A298;
  assign \new_[38819]_  = \new_[38818]_  & \new_[38815]_ ;
  assign \new_[38820]_  = \new_[38819]_  & \new_[38812]_ ;
  assign \new_[38824]_  = ~A166 & ~A167;
  assign \new_[38825]_  = ~A169 & \new_[38824]_ ;
  assign \new_[38829]_  = A201 & ~A200;
  assign \new_[38830]_  = A199 & \new_[38829]_ ;
  assign \new_[38831]_  = \new_[38830]_  & \new_[38825]_ ;
  assign \new_[38835]_  = A233 & A232;
  assign \new_[38836]_  = A203 & \new_[38835]_ ;
  assign \new_[38839]_  = ~A267 & A265;
  assign \new_[38842]_  = A299 & ~A298;
  assign \new_[38843]_  = \new_[38842]_  & \new_[38839]_ ;
  assign \new_[38844]_  = \new_[38843]_  & \new_[38836]_ ;
  assign \new_[38848]_  = ~A166 & ~A167;
  assign \new_[38849]_  = ~A169 & \new_[38848]_ ;
  assign \new_[38853]_  = A201 & ~A200;
  assign \new_[38854]_  = A199 & \new_[38853]_ ;
  assign \new_[38855]_  = \new_[38854]_  & \new_[38849]_ ;
  assign \new_[38859]_  = A233 & A232;
  assign \new_[38860]_  = A203 & \new_[38859]_ ;
  assign \new_[38863]_  = A266 & A265;
  assign \new_[38866]_  = A299 & ~A298;
  assign \new_[38867]_  = \new_[38866]_  & \new_[38863]_ ;
  assign \new_[38868]_  = \new_[38867]_  & \new_[38860]_ ;
  assign \new_[38872]_  = ~A166 & ~A167;
  assign \new_[38873]_  = ~A169 & \new_[38872]_ ;
  assign \new_[38877]_  = A201 & ~A200;
  assign \new_[38878]_  = A199 & \new_[38877]_ ;
  assign \new_[38879]_  = \new_[38878]_  & \new_[38873]_ ;
  assign \new_[38883]_  = A233 & A232;
  assign \new_[38884]_  = A203 & \new_[38883]_ ;
  assign \new_[38887]_  = ~A266 & ~A265;
  assign \new_[38890]_  = A299 & ~A298;
  assign \new_[38891]_  = \new_[38890]_  & \new_[38887]_ ;
  assign \new_[38892]_  = \new_[38891]_  & \new_[38884]_ ;
  assign \new_[38896]_  = ~A166 & ~A167;
  assign \new_[38897]_  = ~A169 & \new_[38896]_ ;
  assign \new_[38901]_  = A201 & ~A200;
  assign \new_[38902]_  = A199 & \new_[38901]_ ;
  assign \new_[38903]_  = \new_[38902]_  & \new_[38897]_ ;
  assign \new_[38907]_  = A233 & ~A232;
  assign \new_[38908]_  = A203 & \new_[38907]_ ;
  assign \new_[38911]_  = ~A266 & A265;
  assign \new_[38914]_  = A268 & A267;
  assign \new_[38915]_  = \new_[38914]_  & \new_[38911]_ ;
  assign \new_[38916]_  = \new_[38915]_  & \new_[38908]_ ;
  assign \new_[38920]_  = ~A166 & ~A167;
  assign \new_[38921]_  = ~A169 & \new_[38920]_ ;
  assign \new_[38925]_  = A201 & ~A200;
  assign \new_[38926]_  = A199 & \new_[38925]_ ;
  assign \new_[38927]_  = \new_[38926]_  & \new_[38921]_ ;
  assign \new_[38931]_  = A233 & ~A232;
  assign \new_[38932]_  = A203 & \new_[38931]_ ;
  assign \new_[38935]_  = ~A266 & A265;
  assign \new_[38938]_  = A269 & A267;
  assign \new_[38939]_  = \new_[38938]_  & \new_[38935]_ ;
  assign \new_[38940]_  = \new_[38939]_  & \new_[38932]_ ;
  assign \new_[38944]_  = ~A166 & ~A167;
  assign \new_[38945]_  = ~A169 & \new_[38944]_ ;
  assign \new_[38949]_  = A201 & ~A200;
  assign \new_[38950]_  = A199 & \new_[38949]_ ;
  assign \new_[38951]_  = \new_[38950]_  & \new_[38945]_ ;
  assign \new_[38955]_  = ~A234 & ~A233;
  assign \new_[38956]_  = A203 & \new_[38955]_ ;
  assign \new_[38959]_  = A266 & A265;
  assign \new_[38962]_  = A299 & ~A298;
  assign \new_[38963]_  = \new_[38962]_  & \new_[38959]_ ;
  assign \new_[38964]_  = \new_[38963]_  & \new_[38956]_ ;
  assign \new_[38968]_  = ~A166 & ~A167;
  assign \new_[38969]_  = ~A169 & \new_[38968]_ ;
  assign \new_[38973]_  = A201 & ~A200;
  assign \new_[38974]_  = A199 & \new_[38973]_ ;
  assign \new_[38975]_  = \new_[38974]_  & \new_[38969]_ ;
  assign \new_[38979]_  = ~A234 & ~A233;
  assign \new_[38980]_  = A203 & \new_[38979]_ ;
  assign \new_[38983]_  = ~A267 & ~A266;
  assign \new_[38986]_  = A299 & ~A298;
  assign \new_[38987]_  = \new_[38986]_  & \new_[38983]_ ;
  assign \new_[38988]_  = \new_[38987]_  & \new_[38980]_ ;
  assign \new_[38992]_  = ~A166 & ~A167;
  assign \new_[38993]_  = ~A169 & \new_[38992]_ ;
  assign \new_[38997]_  = A201 & ~A200;
  assign \new_[38998]_  = A199 & \new_[38997]_ ;
  assign \new_[38999]_  = \new_[38998]_  & \new_[38993]_ ;
  assign \new_[39003]_  = ~A234 & ~A233;
  assign \new_[39004]_  = A203 & \new_[39003]_ ;
  assign \new_[39007]_  = ~A266 & ~A265;
  assign \new_[39010]_  = A299 & ~A298;
  assign \new_[39011]_  = \new_[39010]_  & \new_[39007]_ ;
  assign \new_[39012]_  = \new_[39011]_  & \new_[39004]_ ;
  assign \new_[39016]_  = ~A166 & ~A167;
  assign \new_[39017]_  = ~A169 & \new_[39016]_ ;
  assign \new_[39021]_  = A201 & ~A200;
  assign \new_[39022]_  = A199 & \new_[39021]_ ;
  assign \new_[39023]_  = \new_[39022]_  & \new_[39017]_ ;
  assign \new_[39027]_  = ~A233 & A232;
  assign \new_[39028]_  = A203 & \new_[39027]_ ;
  assign \new_[39031]_  = A235 & A234;
  assign \new_[39034]_  = ~A300 & A298;
  assign \new_[39035]_  = \new_[39034]_  & \new_[39031]_ ;
  assign \new_[39036]_  = \new_[39035]_  & \new_[39028]_ ;
  assign \new_[39040]_  = ~A166 & ~A167;
  assign \new_[39041]_  = ~A169 & \new_[39040]_ ;
  assign \new_[39045]_  = A201 & ~A200;
  assign \new_[39046]_  = A199 & \new_[39045]_ ;
  assign \new_[39047]_  = \new_[39046]_  & \new_[39041]_ ;
  assign \new_[39051]_  = ~A233 & A232;
  assign \new_[39052]_  = A203 & \new_[39051]_ ;
  assign \new_[39055]_  = A235 & A234;
  assign \new_[39058]_  = A299 & A298;
  assign \new_[39059]_  = \new_[39058]_  & \new_[39055]_ ;
  assign \new_[39060]_  = \new_[39059]_  & \new_[39052]_ ;
  assign \new_[39064]_  = ~A166 & ~A167;
  assign \new_[39065]_  = ~A169 & \new_[39064]_ ;
  assign \new_[39069]_  = A201 & ~A200;
  assign \new_[39070]_  = A199 & \new_[39069]_ ;
  assign \new_[39071]_  = \new_[39070]_  & \new_[39065]_ ;
  assign \new_[39075]_  = ~A233 & A232;
  assign \new_[39076]_  = A203 & \new_[39075]_ ;
  assign \new_[39079]_  = A235 & A234;
  assign \new_[39082]_  = ~A299 & ~A298;
  assign \new_[39083]_  = \new_[39082]_  & \new_[39079]_ ;
  assign \new_[39084]_  = \new_[39083]_  & \new_[39076]_ ;
  assign \new_[39088]_  = ~A166 & ~A167;
  assign \new_[39089]_  = ~A169 & \new_[39088]_ ;
  assign \new_[39093]_  = A201 & ~A200;
  assign \new_[39094]_  = A199 & \new_[39093]_ ;
  assign \new_[39095]_  = \new_[39094]_  & \new_[39089]_ ;
  assign \new_[39099]_  = ~A233 & A232;
  assign \new_[39100]_  = A203 & \new_[39099]_ ;
  assign \new_[39103]_  = A235 & A234;
  assign \new_[39106]_  = A266 & ~A265;
  assign \new_[39107]_  = \new_[39106]_  & \new_[39103]_ ;
  assign \new_[39108]_  = \new_[39107]_  & \new_[39100]_ ;
  assign \new_[39112]_  = ~A166 & ~A167;
  assign \new_[39113]_  = ~A169 & \new_[39112]_ ;
  assign \new_[39117]_  = A201 & ~A200;
  assign \new_[39118]_  = A199 & \new_[39117]_ ;
  assign \new_[39119]_  = \new_[39118]_  & \new_[39113]_ ;
  assign \new_[39123]_  = ~A233 & A232;
  assign \new_[39124]_  = A203 & \new_[39123]_ ;
  assign \new_[39127]_  = A236 & A234;
  assign \new_[39130]_  = ~A300 & A298;
  assign \new_[39131]_  = \new_[39130]_  & \new_[39127]_ ;
  assign \new_[39132]_  = \new_[39131]_  & \new_[39124]_ ;
  assign \new_[39136]_  = ~A166 & ~A167;
  assign \new_[39137]_  = ~A169 & \new_[39136]_ ;
  assign \new_[39141]_  = A201 & ~A200;
  assign \new_[39142]_  = A199 & \new_[39141]_ ;
  assign \new_[39143]_  = \new_[39142]_  & \new_[39137]_ ;
  assign \new_[39147]_  = ~A233 & A232;
  assign \new_[39148]_  = A203 & \new_[39147]_ ;
  assign \new_[39151]_  = A236 & A234;
  assign \new_[39154]_  = A299 & A298;
  assign \new_[39155]_  = \new_[39154]_  & \new_[39151]_ ;
  assign \new_[39156]_  = \new_[39155]_  & \new_[39148]_ ;
  assign \new_[39160]_  = ~A166 & ~A167;
  assign \new_[39161]_  = ~A169 & \new_[39160]_ ;
  assign \new_[39165]_  = A201 & ~A200;
  assign \new_[39166]_  = A199 & \new_[39165]_ ;
  assign \new_[39167]_  = \new_[39166]_  & \new_[39161]_ ;
  assign \new_[39171]_  = ~A233 & A232;
  assign \new_[39172]_  = A203 & \new_[39171]_ ;
  assign \new_[39175]_  = A236 & A234;
  assign \new_[39178]_  = ~A299 & ~A298;
  assign \new_[39179]_  = \new_[39178]_  & \new_[39175]_ ;
  assign \new_[39180]_  = \new_[39179]_  & \new_[39172]_ ;
  assign \new_[39184]_  = ~A166 & ~A167;
  assign \new_[39185]_  = ~A169 & \new_[39184]_ ;
  assign \new_[39189]_  = A201 & ~A200;
  assign \new_[39190]_  = A199 & \new_[39189]_ ;
  assign \new_[39191]_  = \new_[39190]_  & \new_[39185]_ ;
  assign \new_[39195]_  = ~A233 & A232;
  assign \new_[39196]_  = A203 & \new_[39195]_ ;
  assign \new_[39199]_  = A236 & A234;
  assign \new_[39202]_  = A266 & ~A265;
  assign \new_[39203]_  = \new_[39202]_  & \new_[39199]_ ;
  assign \new_[39204]_  = \new_[39203]_  & \new_[39196]_ ;
  assign \new_[39208]_  = ~A166 & ~A167;
  assign \new_[39209]_  = ~A169 & \new_[39208]_ ;
  assign \new_[39213]_  = A201 & ~A200;
  assign \new_[39214]_  = A199 & \new_[39213]_ ;
  assign \new_[39215]_  = \new_[39214]_  & \new_[39209]_ ;
  assign \new_[39219]_  = ~A233 & ~A232;
  assign \new_[39220]_  = A203 & \new_[39219]_ ;
  assign \new_[39223]_  = A266 & A265;
  assign \new_[39226]_  = A299 & ~A298;
  assign \new_[39227]_  = \new_[39226]_  & \new_[39223]_ ;
  assign \new_[39228]_  = \new_[39227]_  & \new_[39220]_ ;
  assign \new_[39232]_  = ~A166 & ~A167;
  assign \new_[39233]_  = ~A169 & \new_[39232]_ ;
  assign \new_[39237]_  = A201 & ~A200;
  assign \new_[39238]_  = A199 & \new_[39237]_ ;
  assign \new_[39239]_  = \new_[39238]_  & \new_[39233]_ ;
  assign \new_[39243]_  = ~A233 & ~A232;
  assign \new_[39244]_  = A203 & \new_[39243]_ ;
  assign \new_[39247]_  = ~A267 & ~A266;
  assign \new_[39250]_  = A299 & ~A298;
  assign \new_[39251]_  = \new_[39250]_  & \new_[39247]_ ;
  assign \new_[39252]_  = \new_[39251]_  & \new_[39244]_ ;
  assign \new_[39256]_  = ~A166 & ~A167;
  assign \new_[39257]_  = ~A169 & \new_[39256]_ ;
  assign \new_[39261]_  = A201 & ~A200;
  assign \new_[39262]_  = A199 & \new_[39261]_ ;
  assign \new_[39263]_  = \new_[39262]_  & \new_[39257]_ ;
  assign \new_[39267]_  = ~A233 & ~A232;
  assign \new_[39268]_  = A203 & \new_[39267]_ ;
  assign \new_[39271]_  = ~A266 & ~A265;
  assign \new_[39274]_  = A299 & ~A298;
  assign \new_[39275]_  = \new_[39274]_  & \new_[39271]_ ;
  assign \new_[39276]_  = \new_[39275]_  & \new_[39268]_ ;
  assign \new_[39280]_  = A167 & ~A168;
  assign \new_[39281]_  = ~A169 & \new_[39280]_ ;
  assign \new_[39285]_  = A200 & ~A199;
  assign \new_[39286]_  = A166 & \new_[39285]_ ;
  assign \new_[39287]_  = \new_[39286]_  & \new_[39281]_ ;
  assign \new_[39291]_  = A265 & A233;
  assign \new_[39292]_  = A232 & \new_[39291]_ ;
  assign \new_[39295]_  = ~A269 & ~A268;
  assign \new_[39298]_  = A299 & ~A298;
  assign \new_[39299]_  = \new_[39298]_  & \new_[39295]_ ;
  assign \new_[39300]_  = \new_[39299]_  & \new_[39292]_ ;
  assign \new_[39304]_  = A167 & ~A168;
  assign \new_[39305]_  = ~A169 & \new_[39304]_ ;
  assign \new_[39309]_  = A200 & ~A199;
  assign \new_[39310]_  = A166 & \new_[39309]_ ;
  assign \new_[39311]_  = \new_[39310]_  & \new_[39305]_ ;
  assign \new_[39315]_  = ~A236 & ~A235;
  assign \new_[39316]_  = ~A233 & \new_[39315]_ ;
  assign \new_[39319]_  = A266 & A265;
  assign \new_[39322]_  = A299 & ~A298;
  assign \new_[39323]_  = \new_[39322]_  & \new_[39319]_ ;
  assign \new_[39324]_  = \new_[39323]_  & \new_[39316]_ ;
  assign \new_[39328]_  = A167 & ~A168;
  assign \new_[39329]_  = ~A169 & \new_[39328]_ ;
  assign \new_[39333]_  = A200 & ~A199;
  assign \new_[39334]_  = A166 & \new_[39333]_ ;
  assign \new_[39335]_  = \new_[39334]_  & \new_[39329]_ ;
  assign \new_[39339]_  = ~A236 & ~A235;
  assign \new_[39340]_  = ~A233 & \new_[39339]_ ;
  assign \new_[39343]_  = ~A267 & ~A266;
  assign \new_[39346]_  = A299 & ~A298;
  assign \new_[39347]_  = \new_[39346]_  & \new_[39343]_ ;
  assign \new_[39348]_  = \new_[39347]_  & \new_[39340]_ ;
  assign \new_[39352]_  = A167 & ~A168;
  assign \new_[39353]_  = ~A169 & \new_[39352]_ ;
  assign \new_[39357]_  = A200 & ~A199;
  assign \new_[39358]_  = A166 & \new_[39357]_ ;
  assign \new_[39359]_  = \new_[39358]_  & \new_[39353]_ ;
  assign \new_[39363]_  = ~A236 & ~A235;
  assign \new_[39364]_  = ~A233 & \new_[39363]_ ;
  assign \new_[39367]_  = ~A266 & ~A265;
  assign \new_[39370]_  = A299 & ~A298;
  assign \new_[39371]_  = \new_[39370]_  & \new_[39367]_ ;
  assign \new_[39372]_  = \new_[39371]_  & \new_[39364]_ ;
  assign \new_[39376]_  = A167 & ~A168;
  assign \new_[39377]_  = ~A169 & \new_[39376]_ ;
  assign \new_[39381]_  = A200 & ~A199;
  assign \new_[39382]_  = A166 & \new_[39381]_ ;
  assign \new_[39383]_  = \new_[39382]_  & \new_[39377]_ ;
  assign \new_[39387]_  = ~A266 & ~A234;
  assign \new_[39388]_  = ~A233 & \new_[39387]_ ;
  assign \new_[39391]_  = ~A269 & ~A268;
  assign \new_[39394]_  = A299 & ~A298;
  assign \new_[39395]_  = \new_[39394]_  & \new_[39391]_ ;
  assign \new_[39396]_  = \new_[39395]_  & \new_[39388]_ ;
  assign \new_[39400]_  = A167 & ~A168;
  assign \new_[39401]_  = ~A169 & \new_[39400]_ ;
  assign \new_[39405]_  = A200 & ~A199;
  assign \new_[39406]_  = A166 & \new_[39405]_ ;
  assign \new_[39407]_  = \new_[39406]_  & \new_[39401]_ ;
  assign \new_[39411]_  = A234 & ~A233;
  assign \new_[39412]_  = A232 & \new_[39411]_ ;
  assign \new_[39415]_  = A298 & A235;
  assign \new_[39418]_  = ~A302 & ~A301;
  assign \new_[39419]_  = \new_[39418]_  & \new_[39415]_ ;
  assign \new_[39420]_  = \new_[39419]_  & \new_[39412]_ ;
  assign \new_[39424]_  = A167 & ~A168;
  assign \new_[39425]_  = ~A169 & \new_[39424]_ ;
  assign \new_[39429]_  = A200 & ~A199;
  assign \new_[39430]_  = A166 & \new_[39429]_ ;
  assign \new_[39431]_  = \new_[39430]_  & \new_[39425]_ ;
  assign \new_[39435]_  = A234 & ~A233;
  assign \new_[39436]_  = A232 & \new_[39435]_ ;
  assign \new_[39439]_  = A298 & A236;
  assign \new_[39442]_  = ~A302 & ~A301;
  assign \new_[39443]_  = \new_[39442]_  & \new_[39439]_ ;
  assign \new_[39444]_  = \new_[39443]_  & \new_[39436]_ ;
  assign \new_[39448]_  = A167 & ~A168;
  assign \new_[39449]_  = ~A169 & \new_[39448]_ ;
  assign \new_[39453]_  = A200 & ~A199;
  assign \new_[39454]_  = A166 & \new_[39453]_ ;
  assign \new_[39455]_  = \new_[39454]_  & \new_[39449]_ ;
  assign \new_[39459]_  = ~A266 & ~A233;
  assign \new_[39460]_  = ~A232 & \new_[39459]_ ;
  assign \new_[39463]_  = ~A269 & ~A268;
  assign \new_[39466]_  = A299 & ~A298;
  assign \new_[39467]_  = \new_[39466]_  & \new_[39463]_ ;
  assign \new_[39468]_  = \new_[39467]_  & \new_[39460]_ ;
  assign \new_[39472]_  = A167 & ~A168;
  assign \new_[39473]_  = ~A169 & \new_[39472]_ ;
  assign \new_[39477]_  = ~A200 & A199;
  assign \new_[39478]_  = A166 & \new_[39477]_ ;
  assign \new_[39479]_  = \new_[39478]_  & \new_[39473]_ ;
  assign \new_[39483]_  = ~A232 & A202;
  assign \new_[39484]_  = A201 & \new_[39483]_ ;
  assign \new_[39487]_  = ~A299 & A233;
  assign \new_[39490]_  = ~A302 & ~A301;
  assign \new_[39491]_  = \new_[39490]_  & \new_[39487]_ ;
  assign \new_[39492]_  = \new_[39491]_  & \new_[39484]_ ;
  assign \new_[39496]_  = A167 & ~A168;
  assign \new_[39497]_  = ~A169 & \new_[39496]_ ;
  assign \new_[39501]_  = ~A200 & A199;
  assign \new_[39502]_  = A166 & \new_[39501]_ ;
  assign \new_[39503]_  = \new_[39502]_  & \new_[39497]_ ;
  assign \new_[39507]_  = ~A232 & A203;
  assign \new_[39508]_  = A201 & \new_[39507]_ ;
  assign \new_[39511]_  = ~A299 & A233;
  assign \new_[39514]_  = ~A302 & ~A301;
  assign \new_[39515]_  = \new_[39514]_  & \new_[39511]_ ;
  assign \new_[39516]_  = \new_[39515]_  & \new_[39508]_ ;
  assign \new_[39520]_  = A167 & ~A169;
  assign \new_[39521]_  = A170 & \new_[39520]_ ;
  assign \new_[39525]_  = A200 & A199;
  assign \new_[39526]_  = ~A166 & \new_[39525]_ ;
  assign \new_[39527]_  = \new_[39526]_  & \new_[39521]_ ;
  assign \new_[39531]_  = A265 & A233;
  assign \new_[39532]_  = A232 & \new_[39531]_ ;
  assign \new_[39535]_  = ~A269 & ~A268;
  assign \new_[39538]_  = A299 & ~A298;
  assign \new_[39539]_  = \new_[39538]_  & \new_[39535]_ ;
  assign \new_[39540]_  = \new_[39539]_  & \new_[39532]_ ;
  assign \new_[39544]_  = A167 & ~A169;
  assign \new_[39545]_  = A170 & \new_[39544]_ ;
  assign \new_[39549]_  = A200 & A199;
  assign \new_[39550]_  = ~A166 & \new_[39549]_ ;
  assign \new_[39551]_  = \new_[39550]_  & \new_[39545]_ ;
  assign \new_[39555]_  = ~A236 & ~A235;
  assign \new_[39556]_  = ~A233 & \new_[39555]_ ;
  assign \new_[39559]_  = A266 & A265;
  assign \new_[39562]_  = A299 & ~A298;
  assign \new_[39563]_  = \new_[39562]_  & \new_[39559]_ ;
  assign \new_[39564]_  = \new_[39563]_  & \new_[39556]_ ;
  assign \new_[39568]_  = A167 & ~A169;
  assign \new_[39569]_  = A170 & \new_[39568]_ ;
  assign \new_[39573]_  = A200 & A199;
  assign \new_[39574]_  = ~A166 & \new_[39573]_ ;
  assign \new_[39575]_  = \new_[39574]_  & \new_[39569]_ ;
  assign \new_[39579]_  = ~A236 & ~A235;
  assign \new_[39580]_  = ~A233 & \new_[39579]_ ;
  assign \new_[39583]_  = ~A267 & ~A266;
  assign \new_[39586]_  = A299 & ~A298;
  assign \new_[39587]_  = \new_[39586]_  & \new_[39583]_ ;
  assign \new_[39588]_  = \new_[39587]_  & \new_[39580]_ ;
  assign \new_[39592]_  = A167 & ~A169;
  assign \new_[39593]_  = A170 & \new_[39592]_ ;
  assign \new_[39597]_  = A200 & A199;
  assign \new_[39598]_  = ~A166 & \new_[39597]_ ;
  assign \new_[39599]_  = \new_[39598]_  & \new_[39593]_ ;
  assign \new_[39603]_  = ~A236 & ~A235;
  assign \new_[39604]_  = ~A233 & \new_[39603]_ ;
  assign \new_[39607]_  = ~A266 & ~A265;
  assign \new_[39610]_  = A299 & ~A298;
  assign \new_[39611]_  = \new_[39610]_  & \new_[39607]_ ;
  assign \new_[39612]_  = \new_[39611]_  & \new_[39604]_ ;
  assign \new_[39616]_  = A167 & ~A169;
  assign \new_[39617]_  = A170 & \new_[39616]_ ;
  assign \new_[39621]_  = A200 & A199;
  assign \new_[39622]_  = ~A166 & \new_[39621]_ ;
  assign \new_[39623]_  = \new_[39622]_  & \new_[39617]_ ;
  assign \new_[39627]_  = ~A266 & ~A234;
  assign \new_[39628]_  = ~A233 & \new_[39627]_ ;
  assign \new_[39631]_  = ~A269 & ~A268;
  assign \new_[39634]_  = A299 & ~A298;
  assign \new_[39635]_  = \new_[39634]_  & \new_[39631]_ ;
  assign \new_[39636]_  = \new_[39635]_  & \new_[39628]_ ;
  assign \new_[39640]_  = A167 & ~A169;
  assign \new_[39641]_  = A170 & \new_[39640]_ ;
  assign \new_[39645]_  = A200 & A199;
  assign \new_[39646]_  = ~A166 & \new_[39645]_ ;
  assign \new_[39647]_  = \new_[39646]_  & \new_[39641]_ ;
  assign \new_[39651]_  = A234 & ~A233;
  assign \new_[39652]_  = A232 & \new_[39651]_ ;
  assign \new_[39655]_  = A298 & A235;
  assign \new_[39658]_  = ~A302 & ~A301;
  assign \new_[39659]_  = \new_[39658]_  & \new_[39655]_ ;
  assign \new_[39660]_  = \new_[39659]_  & \new_[39652]_ ;
  assign \new_[39664]_  = A167 & ~A169;
  assign \new_[39665]_  = A170 & \new_[39664]_ ;
  assign \new_[39669]_  = A200 & A199;
  assign \new_[39670]_  = ~A166 & \new_[39669]_ ;
  assign \new_[39671]_  = \new_[39670]_  & \new_[39665]_ ;
  assign \new_[39675]_  = A234 & ~A233;
  assign \new_[39676]_  = A232 & \new_[39675]_ ;
  assign \new_[39679]_  = A298 & A236;
  assign \new_[39682]_  = ~A302 & ~A301;
  assign \new_[39683]_  = \new_[39682]_  & \new_[39679]_ ;
  assign \new_[39684]_  = \new_[39683]_  & \new_[39676]_ ;
  assign \new_[39688]_  = A167 & ~A169;
  assign \new_[39689]_  = A170 & \new_[39688]_ ;
  assign \new_[39693]_  = A200 & A199;
  assign \new_[39694]_  = ~A166 & \new_[39693]_ ;
  assign \new_[39695]_  = \new_[39694]_  & \new_[39689]_ ;
  assign \new_[39699]_  = ~A266 & ~A233;
  assign \new_[39700]_  = ~A232 & \new_[39699]_ ;
  assign \new_[39703]_  = ~A269 & ~A268;
  assign \new_[39706]_  = A299 & ~A298;
  assign \new_[39707]_  = \new_[39706]_  & \new_[39703]_ ;
  assign \new_[39708]_  = \new_[39707]_  & \new_[39700]_ ;
  assign \new_[39712]_  = A167 & ~A169;
  assign \new_[39713]_  = A170 & \new_[39712]_ ;
  assign \new_[39717]_  = ~A202 & ~A200;
  assign \new_[39718]_  = ~A166 & \new_[39717]_ ;
  assign \new_[39719]_  = \new_[39718]_  & \new_[39713]_ ;
  assign \new_[39723]_  = A233 & A232;
  assign \new_[39724]_  = ~A203 & \new_[39723]_ ;
  assign \new_[39727]_  = ~A267 & A265;
  assign \new_[39730]_  = A299 & ~A298;
  assign \new_[39731]_  = \new_[39730]_  & \new_[39727]_ ;
  assign \new_[39732]_  = \new_[39731]_  & \new_[39724]_ ;
  assign \new_[39736]_  = A167 & ~A169;
  assign \new_[39737]_  = A170 & \new_[39736]_ ;
  assign \new_[39741]_  = ~A202 & ~A200;
  assign \new_[39742]_  = ~A166 & \new_[39741]_ ;
  assign \new_[39743]_  = \new_[39742]_  & \new_[39737]_ ;
  assign \new_[39747]_  = A233 & A232;
  assign \new_[39748]_  = ~A203 & \new_[39747]_ ;
  assign \new_[39751]_  = A266 & A265;
  assign \new_[39754]_  = A299 & ~A298;
  assign \new_[39755]_  = \new_[39754]_  & \new_[39751]_ ;
  assign \new_[39756]_  = \new_[39755]_  & \new_[39748]_ ;
  assign \new_[39760]_  = A167 & ~A169;
  assign \new_[39761]_  = A170 & \new_[39760]_ ;
  assign \new_[39765]_  = ~A202 & ~A200;
  assign \new_[39766]_  = ~A166 & \new_[39765]_ ;
  assign \new_[39767]_  = \new_[39766]_  & \new_[39761]_ ;
  assign \new_[39771]_  = A233 & A232;
  assign \new_[39772]_  = ~A203 & \new_[39771]_ ;
  assign \new_[39775]_  = ~A266 & ~A265;
  assign \new_[39778]_  = A299 & ~A298;
  assign \new_[39779]_  = \new_[39778]_  & \new_[39775]_ ;
  assign \new_[39780]_  = \new_[39779]_  & \new_[39772]_ ;
  assign \new_[39784]_  = A167 & ~A169;
  assign \new_[39785]_  = A170 & \new_[39784]_ ;
  assign \new_[39789]_  = ~A202 & ~A200;
  assign \new_[39790]_  = ~A166 & \new_[39789]_ ;
  assign \new_[39791]_  = \new_[39790]_  & \new_[39785]_ ;
  assign \new_[39795]_  = A233 & ~A232;
  assign \new_[39796]_  = ~A203 & \new_[39795]_ ;
  assign \new_[39799]_  = ~A266 & A265;
  assign \new_[39802]_  = A268 & A267;
  assign \new_[39803]_  = \new_[39802]_  & \new_[39799]_ ;
  assign \new_[39804]_  = \new_[39803]_  & \new_[39796]_ ;
  assign \new_[39808]_  = A167 & ~A169;
  assign \new_[39809]_  = A170 & \new_[39808]_ ;
  assign \new_[39813]_  = ~A202 & ~A200;
  assign \new_[39814]_  = ~A166 & \new_[39813]_ ;
  assign \new_[39815]_  = \new_[39814]_  & \new_[39809]_ ;
  assign \new_[39819]_  = A233 & ~A232;
  assign \new_[39820]_  = ~A203 & \new_[39819]_ ;
  assign \new_[39823]_  = ~A266 & A265;
  assign \new_[39826]_  = A269 & A267;
  assign \new_[39827]_  = \new_[39826]_  & \new_[39823]_ ;
  assign \new_[39828]_  = \new_[39827]_  & \new_[39820]_ ;
  assign \new_[39832]_  = A167 & ~A169;
  assign \new_[39833]_  = A170 & \new_[39832]_ ;
  assign \new_[39837]_  = ~A202 & ~A200;
  assign \new_[39838]_  = ~A166 & \new_[39837]_ ;
  assign \new_[39839]_  = \new_[39838]_  & \new_[39833]_ ;
  assign \new_[39843]_  = ~A234 & ~A233;
  assign \new_[39844]_  = ~A203 & \new_[39843]_ ;
  assign \new_[39847]_  = A266 & A265;
  assign \new_[39850]_  = A299 & ~A298;
  assign \new_[39851]_  = \new_[39850]_  & \new_[39847]_ ;
  assign \new_[39852]_  = \new_[39851]_  & \new_[39844]_ ;
  assign \new_[39856]_  = A167 & ~A169;
  assign \new_[39857]_  = A170 & \new_[39856]_ ;
  assign \new_[39861]_  = ~A202 & ~A200;
  assign \new_[39862]_  = ~A166 & \new_[39861]_ ;
  assign \new_[39863]_  = \new_[39862]_  & \new_[39857]_ ;
  assign \new_[39867]_  = ~A234 & ~A233;
  assign \new_[39868]_  = ~A203 & \new_[39867]_ ;
  assign \new_[39871]_  = ~A267 & ~A266;
  assign \new_[39874]_  = A299 & ~A298;
  assign \new_[39875]_  = \new_[39874]_  & \new_[39871]_ ;
  assign \new_[39876]_  = \new_[39875]_  & \new_[39868]_ ;
  assign \new_[39880]_  = A167 & ~A169;
  assign \new_[39881]_  = A170 & \new_[39880]_ ;
  assign \new_[39885]_  = ~A202 & ~A200;
  assign \new_[39886]_  = ~A166 & \new_[39885]_ ;
  assign \new_[39887]_  = \new_[39886]_  & \new_[39881]_ ;
  assign \new_[39891]_  = ~A234 & ~A233;
  assign \new_[39892]_  = ~A203 & \new_[39891]_ ;
  assign \new_[39895]_  = ~A266 & ~A265;
  assign \new_[39898]_  = A299 & ~A298;
  assign \new_[39899]_  = \new_[39898]_  & \new_[39895]_ ;
  assign \new_[39900]_  = \new_[39899]_  & \new_[39892]_ ;
  assign \new_[39904]_  = A167 & ~A169;
  assign \new_[39905]_  = A170 & \new_[39904]_ ;
  assign \new_[39909]_  = ~A202 & ~A200;
  assign \new_[39910]_  = ~A166 & \new_[39909]_ ;
  assign \new_[39911]_  = \new_[39910]_  & \new_[39905]_ ;
  assign \new_[39915]_  = ~A233 & A232;
  assign \new_[39916]_  = ~A203 & \new_[39915]_ ;
  assign \new_[39919]_  = A235 & A234;
  assign \new_[39922]_  = ~A300 & A298;
  assign \new_[39923]_  = \new_[39922]_  & \new_[39919]_ ;
  assign \new_[39924]_  = \new_[39923]_  & \new_[39916]_ ;
  assign \new_[39928]_  = A167 & ~A169;
  assign \new_[39929]_  = A170 & \new_[39928]_ ;
  assign \new_[39933]_  = ~A202 & ~A200;
  assign \new_[39934]_  = ~A166 & \new_[39933]_ ;
  assign \new_[39935]_  = \new_[39934]_  & \new_[39929]_ ;
  assign \new_[39939]_  = ~A233 & A232;
  assign \new_[39940]_  = ~A203 & \new_[39939]_ ;
  assign \new_[39943]_  = A235 & A234;
  assign \new_[39946]_  = A299 & A298;
  assign \new_[39947]_  = \new_[39946]_  & \new_[39943]_ ;
  assign \new_[39948]_  = \new_[39947]_  & \new_[39940]_ ;
  assign \new_[39952]_  = A167 & ~A169;
  assign \new_[39953]_  = A170 & \new_[39952]_ ;
  assign \new_[39957]_  = ~A202 & ~A200;
  assign \new_[39958]_  = ~A166 & \new_[39957]_ ;
  assign \new_[39959]_  = \new_[39958]_  & \new_[39953]_ ;
  assign \new_[39963]_  = ~A233 & A232;
  assign \new_[39964]_  = ~A203 & \new_[39963]_ ;
  assign \new_[39967]_  = A235 & A234;
  assign \new_[39970]_  = ~A299 & ~A298;
  assign \new_[39971]_  = \new_[39970]_  & \new_[39967]_ ;
  assign \new_[39972]_  = \new_[39971]_  & \new_[39964]_ ;
  assign \new_[39976]_  = A167 & ~A169;
  assign \new_[39977]_  = A170 & \new_[39976]_ ;
  assign \new_[39981]_  = ~A202 & ~A200;
  assign \new_[39982]_  = ~A166 & \new_[39981]_ ;
  assign \new_[39983]_  = \new_[39982]_  & \new_[39977]_ ;
  assign \new_[39987]_  = ~A233 & A232;
  assign \new_[39988]_  = ~A203 & \new_[39987]_ ;
  assign \new_[39991]_  = A235 & A234;
  assign \new_[39994]_  = A266 & ~A265;
  assign \new_[39995]_  = \new_[39994]_  & \new_[39991]_ ;
  assign \new_[39996]_  = \new_[39995]_  & \new_[39988]_ ;
  assign \new_[40000]_  = A167 & ~A169;
  assign \new_[40001]_  = A170 & \new_[40000]_ ;
  assign \new_[40005]_  = ~A202 & ~A200;
  assign \new_[40006]_  = ~A166 & \new_[40005]_ ;
  assign \new_[40007]_  = \new_[40006]_  & \new_[40001]_ ;
  assign \new_[40011]_  = ~A233 & A232;
  assign \new_[40012]_  = ~A203 & \new_[40011]_ ;
  assign \new_[40015]_  = A236 & A234;
  assign \new_[40018]_  = ~A300 & A298;
  assign \new_[40019]_  = \new_[40018]_  & \new_[40015]_ ;
  assign \new_[40020]_  = \new_[40019]_  & \new_[40012]_ ;
  assign \new_[40024]_  = A167 & ~A169;
  assign \new_[40025]_  = A170 & \new_[40024]_ ;
  assign \new_[40029]_  = ~A202 & ~A200;
  assign \new_[40030]_  = ~A166 & \new_[40029]_ ;
  assign \new_[40031]_  = \new_[40030]_  & \new_[40025]_ ;
  assign \new_[40035]_  = ~A233 & A232;
  assign \new_[40036]_  = ~A203 & \new_[40035]_ ;
  assign \new_[40039]_  = A236 & A234;
  assign \new_[40042]_  = A299 & A298;
  assign \new_[40043]_  = \new_[40042]_  & \new_[40039]_ ;
  assign \new_[40044]_  = \new_[40043]_  & \new_[40036]_ ;
  assign \new_[40048]_  = A167 & ~A169;
  assign \new_[40049]_  = A170 & \new_[40048]_ ;
  assign \new_[40053]_  = ~A202 & ~A200;
  assign \new_[40054]_  = ~A166 & \new_[40053]_ ;
  assign \new_[40055]_  = \new_[40054]_  & \new_[40049]_ ;
  assign \new_[40059]_  = ~A233 & A232;
  assign \new_[40060]_  = ~A203 & \new_[40059]_ ;
  assign \new_[40063]_  = A236 & A234;
  assign \new_[40066]_  = ~A299 & ~A298;
  assign \new_[40067]_  = \new_[40066]_  & \new_[40063]_ ;
  assign \new_[40068]_  = \new_[40067]_  & \new_[40060]_ ;
  assign \new_[40072]_  = A167 & ~A169;
  assign \new_[40073]_  = A170 & \new_[40072]_ ;
  assign \new_[40077]_  = ~A202 & ~A200;
  assign \new_[40078]_  = ~A166 & \new_[40077]_ ;
  assign \new_[40079]_  = \new_[40078]_  & \new_[40073]_ ;
  assign \new_[40083]_  = ~A233 & A232;
  assign \new_[40084]_  = ~A203 & \new_[40083]_ ;
  assign \new_[40087]_  = A236 & A234;
  assign \new_[40090]_  = A266 & ~A265;
  assign \new_[40091]_  = \new_[40090]_  & \new_[40087]_ ;
  assign \new_[40092]_  = \new_[40091]_  & \new_[40084]_ ;
  assign \new_[40096]_  = A167 & ~A169;
  assign \new_[40097]_  = A170 & \new_[40096]_ ;
  assign \new_[40101]_  = ~A202 & ~A200;
  assign \new_[40102]_  = ~A166 & \new_[40101]_ ;
  assign \new_[40103]_  = \new_[40102]_  & \new_[40097]_ ;
  assign \new_[40107]_  = ~A233 & ~A232;
  assign \new_[40108]_  = ~A203 & \new_[40107]_ ;
  assign \new_[40111]_  = A266 & A265;
  assign \new_[40114]_  = A299 & ~A298;
  assign \new_[40115]_  = \new_[40114]_  & \new_[40111]_ ;
  assign \new_[40116]_  = \new_[40115]_  & \new_[40108]_ ;
  assign \new_[40120]_  = A167 & ~A169;
  assign \new_[40121]_  = A170 & \new_[40120]_ ;
  assign \new_[40125]_  = ~A202 & ~A200;
  assign \new_[40126]_  = ~A166 & \new_[40125]_ ;
  assign \new_[40127]_  = \new_[40126]_  & \new_[40121]_ ;
  assign \new_[40131]_  = ~A233 & ~A232;
  assign \new_[40132]_  = ~A203 & \new_[40131]_ ;
  assign \new_[40135]_  = ~A267 & ~A266;
  assign \new_[40138]_  = A299 & ~A298;
  assign \new_[40139]_  = \new_[40138]_  & \new_[40135]_ ;
  assign \new_[40140]_  = \new_[40139]_  & \new_[40132]_ ;
  assign \new_[40144]_  = A167 & ~A169;
  assign \new_[40145]_  = A170 & \new_[40144]_ ;
  assign \new_[40149]_  = ~A202 & ~A200;
  assign \new_[40150]_  = ~A166 & \new_[40149]_ ;
  assign \new_[40151]_  = \new_[40150]_  & \new_[40145]_ ;
  assign \new_[40155]_  = ~A233 & ~A232;
  assign \new_[40156]_  = ~A203 & \new_[40155]_ ;
  assign \new_[40159]_  = ~A266 & ~A265;
  assign \new_[40162]_  = A299 & ~A298;
  assign \new_[40163]_  = \new_[40162]_  & \new_[40159]_ ;
  assign \new_[40164]_  = \new_[40163]_  & \new_[40156]_ ;
  assign \new_[40168]_  = A167 & ~A169;
  assign \new_[40169]_  = A170 & \new_[40168]_ ;
  assign \new_[40173]_  = ~A201 & ~A200;
  assign \new_[40174]_  = ~A166 & \new_[40173]_ ;
  assign \new_[40175]_  = \new_[40174]_  & \new_[40169]_ ;
  assign \new_[40179]_  = A265 & A233;
  assign \new_[40180]_  = A232 & \new_[40179]_ ;
  assign \new_[40183]_  = ~A269 & ~A268;
  assign \new_[40186]_  = A299 & ~A298;
  assign \new_[40187]_  = \new_[40186]_  & \new_[40183]_ ;
  assign \new_[40188]_  = \new_[40187]_  & \new_[40180]_ ;
  assign \new_[40192]_  = A167 & ~A169;
  assign \new_[40193]_  = A170 & \new_[40192]_ ;
  assign \new_[40197]_  = ~A201 & ~A200;
  assign \new_[40198]_  = ~A166 & \new_[40197]_ ;
  assign \new_[40199]_  = \new_[40198]_  & \new_[40193]_ ;
  assign \new_[40203]_  = ~A236 & ~A235;
  assign \new_[40204]_  = ~A233 & \new_[40203]_ ;
  assign \new_[40207]_  = A266 & A265;
  assign \new_[40210]_  = A299 & ~A298;
  assign \new_[40211]_  = \new_[40210]_  & \new_[40207]_ ;
  assign \new_[40212]_  = \new_[40211]_  & \new_[40204]_ ;
  assign \new_[40216]_  = A167 & ~A169;
  assign \new_[40217]_  = A170 & \new_[40216]_ ;
  assign \new_[40221]_  = ~A201 & ~A200;
  assign \new_[40222]_  = ~A166 & \new_[40221]_ ;
  assign \new_[40223]_  = \new_[40222]_  & \new_[40217]_ ;
  assign \new_[40227]_  = ~A236 & ~A235;
  assign \new_[40228]_  = ~A233 & \new_[40227]_ ;
  assign \new_[40231]_  = ~A267 & ~A266;
  assign \new_[40234]_  = A299 & ~A298;
  assign \new_[40235]_  = \new_[40234]_  & \new_[40231]_ ;
  assign \new_[40236]_  = \new_[40235]_  & \new_[40228]_ ;
  assign \new_[40240]_  = A167 & ~A169;
  assign \new_[40241]_  = A170 & \new_[40240]_ ;
  assign \new_[40245]_  = ~A201 & ~A200;
  assign \new_[40246]_  = ~A166 & \new_[40245]_ ;
  assign \new_[40247]_  = \new_[40246]_  & \new_[40241]_ ;
  assign \new_[40251]_  = ~A236 & ~A235;
  assign \new_[40252]_  = ~A233 & \new_[40251]_ ;
  assign \new_[40255]_  = ~A266 & ~A265;
  assign \new_[40258]_  = A299 & ~A298;
  assign \new_[40259]_  = \new_[40258]_  & \new_[40255]_ ;
  assign \new_[40260]_  = \new_[40259]_  & \new_[40252]_ ;
  assign \new_[40264]_  = A167 & ~A169;
  assign \new_[40265]_  = A170 & \new_[40264]_ ;
  assign \new_[40269]_  = ~A201 & ~A200;
  assign \new_[40270]_  = ~A166 & \new_[40269]_ ;
  assign \new_[40271]_  = \new_[40270]_  & \new_[40265]_ ;
  assign \new_[40275]_  = ~A266 & ~A234;
  assign \new_[40276]_  = ~A233 & \new_[40275]_ ;
  assign \new_[40279]_  = ~A269 & ~A268;
  assign \new_[40282]_  = A299 & ~A298;
  assign \new_[40283]_  = \new_[40282]_  & \new_[40279]_ ;
  assign \new_[40284]_  = \new_[40283]_  & \new_[40276]_ ;
  assign \new_[40288]_  = A167 & ~A169;
  assign \new_[40289]_  = A170 & \new_[40288]_ ;
  assign \new_[40293]_  = ~A201 & ~A200;
  assign \new_[40294]_  = ~A166 & \new_[40293]_ ;
  assign \new_[40295]_  = \new_[40294]_  & \new_[40289]_ ;
  assign \new_[40299]_  = A234 & ~A233;
  assign \new_[40300]_  = A232 & \new_[40299]_ ;
  assign \new_[40303]_  = A298 & A235;
  assign \new_[40306]_  = ~A302 & ~A301;
  assign \new_[40307]_  = \new_[40306]_  & \new_[40303]_ ;
  assign \new_[40308]_  = \new_[40307]_  & \new_[40300]_ ;
  assign \new_[40312]_  = A167 & ~A169;
  assign \new_[40313]_  = A170 & \new_[40312]_ ;
  assign \new_[40317]_  = ~A201 & ~A200;
  assign \new_[40318]_  = ~A166 & \new_[40317]_ ;
  assign \new_[40319]_  = \new_[40318]_  & \new_[40313]_ ;
  assign \new_[40323]_  = A234 & ~A233;
  assign \new_[40324]_  = A232 & \new_[40323]_ ;
  assign \new_[40327]_  = A298 & A236;
  assign \new_[40330]_  = ~A302 & ~A301;
  assign \new_[40331]_  = \new_[40330]_  & \new_[40327]_ ;
  assign \new_[40332]_  = \new_[40331]_  & \new_[40324]_ ;
  assign \new_[40336]_  = A167 & ~A169;
  assign \new_[40337]_  = A170 & \new_[40336]_ ;
  assign \new_[40341]_  = ~A201 & ~A200;
  assign \new_[40342]_  = ~A166 & \new_[40341]_ ;
  assign \new_[40343]_  = \new_[40342]_  & \new_[40337]_ ;
  assign \new_[40347]_  = ~A266 & ~A233;
  assign \new_[40348]_  = ~A232 & \new_[40347]_ ;
  assign \new_[40351]_  = ~A269 & ~A268;
  assign \new_[40354]_  = A299 & ~A298;
  assign \new_[40355]_  = \new_[40354]_  & \new_[40351]_ ;
  assign \new_[40356]_  = \new_[40355]_  & \new_[40348]_ ;
  assign \new_[40360]_  = A167 & ~A169;
  assign \new_[40361]_  = A170 & \new_[40360]_ ;
  assign \new_[40365]_  = ~A200 & ~A199;
  assign \new_[40366]_  = ~A166 & \new_[40365]_ ;
  assign \new_[40367]_  = \new_[40366]_  & \new_[40361]_ ;
  assign \new_[40371]_  = A265 & A233;
  assign \new_[40372]_  = A232 & \new_[40371]_ ;
  assign \new_[40375]_  = ~A269 & ~A268;
  assign \new_[40378]_  = A299 & ~A298;
  assign \new_[40379]_  = \new_[40378]_  & \new_[40375]_ ;
  assign \new_[40380]_  = \new_[40379]_  & \new_[40372]_ ;
  assign \new_[40384]_  = A167 & ~A169;
  assign \new_[40385]_  = A170 & \new_[40384]_ ;
  assign \new_[40389]_  = ~A200 & ~A199;
  assign \new_[40390]_  = ~A166 & \new_[40389]_ ;
  assign \new_[40391]_  = \new_[40390]_  & \new_[40385]_ ;
  assign \new_[40395]_  = ~A236 & ~A235;
  assign \new_[40396]_  = ~A233 & \new_[40395]_ ;
  assign \new_[40399]_  = A266 & A265;
  assign \new_[40402]_  = A299 & ~A298;
  assign \new_[40403]_  = \new_[40402]_  & \new_[40399]_ ;
  assign \new_[40404]_  = \new_[40403]_  & \new_[40396]_ ;
  assign \new_[40408]_  = A167 & ~A169;
  assign \new_[40409]_  = A170 & \new_[40408]_ ;
  assign \new_[40413]_  = ~A200 & ~A199;
  assign \new_[40414]_  = ~A166 & \new_[40413]_ ;
  assign \new_[40415]_  = \new_[40414]_  & \new_[40409]_ ;
  assign \new_[40419]_  = ~A236 & ~A235;
  assign \new_[40420]_  = ~A233 & \new_[40419]_ ;
  assign \new_[40423]_  = ~A267 & ~A266;
  assign \new_[40426]_  = A299 & ~A298;
  assign \new_[40427]_  = \new_[40426]_  & \new_[40423]_ ;
  assign \new_[40428]_  = \new_[40427]_  & \new_[40420]_ ;
  assign \new_[40432]_  = A167 & ~A169;
  assign \new_[40433]_  = A170 & \new_[40432]_ ;
  assign \new_[40437]_  = ~A200 & ~A199;
  assign \new_[40438]_  = ~A166 & \new_[40437]_ ;
  assign \new_[40439]_  = \new_[40438]_  & \new_[40433]_ ;
  assign \new_[40443]_  = ~A236 & ~A235;
  assign \new_[40444]_  = ~A233 & \new_[40443]_ ;
  assign \new_[40447]_  = ~A266 & ~A265;
  assign \new_[40450]_  = A299 & ~A298;
  assign \new_[40451]_  = \new_[40450]_  & \new_[40447]_ ;
  assign \new_[40452]_  = \new_[40451]_  & \new_[40444]_ ;
  assign \new_[40456]_  = A167 & ~A169;
  assign \new_[40457]_  = A170 & \new_[40456]_ ;
  assign \new_[40461]_  = ~A200 & ~A199;
  assign \new_[40462]_  = ~A166 & \new_[40461]_ ;
  assign \new_[40463]_  = \new_[40462]_  & \new_[40457]_ ;
  assign \new_[40467]_  = ~A266 & ~A234;
  assign \new_[40468]_  = ~A233 & \new_[40467]_ ;
  assign \new_[40471]_  = ~A269 & ~A268;
  assign \new_[40474]_  = A299 & ~A298;
  assign \new_[40475]_  = \new_[40474]_  & \new_[40471]_ ;
  assign \new_[40476]_  = \new_[40475]_  & \new_[40468]_ ;
  assign \new_[40480]_  = A167 & ~A169;
  assign \new_[40481]_  = A170 & \new_[40480]_ ;
  assign \new_[40485]_  = ~A200 & ~A199;
  assign \new_[40486]_  = ~A166 & \new_[40485]_ ;
  assign \new_[40487]_  = \new_[40486]_  & \new_[40481]_ ;
  assign \new_[40491]_  = A234 & ~A233;
  assign \new_[40492]_  = A232 & \new_[40491]_ ;
  assign \new_[40495]_  = A298 & A235;
  assign \new_[40498]_  = ~A302 & ~A301;
  assign \new_[40499]_  = \new_[40498]_  & \new_[40495]_ ;
  assign \new_[40500]_  = \new_[40499]_  & \new_[40492]_ ;
  assign \new_[40504]_  = A167 & ~A169;
  assign \new_[40505]_  = A170 & \new_[40504]_ ;
  assign \new_[40509]_  = ~A200 & ~A199;
  assign \new_[40510]_  = ~A166 & \new_[40509]_ ;
  assign \new_[40511]_  = \new_[40510]_  & \new_[40505]_ ;
  assign \new_[40515]_  = A234 & ~A233;
  assign \new_[40516]_  = A232 & \new_[40515]_ ;
  assign \new_[40519]_  = A298 & A236;
  assign \new_[40522]_  = ~A302 & ~A301;
  assign \new_[40523]_  = \new_[40522]_  & \new_[40519]_ ;
  assign \new_[40524]_  = \new_[40523]_  & \new_[40516]_ ;
  assign \new_[40528]_  = A167 & ~A169;
  assign \new_[40529]_  = A170 & \new_[40528]_ ;
  assign \new_[40533]_  = ~A200 & ~A199;
  assign \new_[40534]_  = ~A166 & \new_[40533]_ ;
  assign \new_[40535]_  = \new_[40534]_  & \new_[40529]_ ;
  assign \new_[40539]_  = ~A266 & ~A233;
  assign \new_[40540]_  = ~A232 & \new_[40539]_ ;
  assign \new_[40543]_  = ~A269 & ~A268;
  assign \new_[40546]_  = A299 & ~A298;
  assign \new_[40547]_  = \new_[40546]_  & \new_[40543]_ ;
  assign \new_[40548]_  = \new_[40547]_  & \new_[40540]_ ;
  assign \new_[40552]_  = ~A167 & ~A169;
  assign \new_[40553]_  = A170 & \new_[40552]_ ;
  assign \new_[40557]_  = A200 & A199;
  assign \new_[40558]_  = A166 & \new_[40557]_ ;
  assign \new_[40559]_  = \new_[40558]_  & \new_[40553]_ ;
  assign \new_[40563]_  = A265 & A233;
  assign \new_[40564]_  = A232 & \new_[40563]_ ;
  assign \new_[40567]_  = ~A269 & ~A268;
  assign \new_[40570]_  = A299 & ~A298;
  assign \new_[40571]_  = \new_[40570]_  & \new_[40567]_ ;
  assign \new_[40572]_  = \new_[40571]_  & \new_[40564]_ ;
  assign \new_[40576]_  = ~A167 & ~A169;
  assign \new_[40577]_  = A170 & \new_[40576]_ ;
  assign \new_[40581]_  = A200 & A199;
  assign \new_[40582]_  = A166 & \new_[40581]_ ;
  assign \new_[40583]_  = \new_[40582]_  & \new_[40577]_ ;
  assign \new_[40587]_  = ~A236 & ~A235;
  assign \new_[40588]_  = ~A233 & \new_[40587]_ ;
  assign \new_[40591]_  = A266 & A265;
  assign \new_[40594]_  = A299 & ~A298;
  assign \new_[40595]_  = \new_[40594]_  & \new_[40591]_ ;
  assign \new_[40596]_  = \new_[40595]_  & \new_[40588]_ ;
  assign \new_[40600]_  = ~A167 & ~A169;
  assign \new_[40601]_  = A170 & \new_[40600]_ ;
  assign \new_[40605]_  = A200 & A199;
  assign \new_[40606]_  = A166 & \new_[40605]_ ;
  assign \new_[40607]_  = \new_[40606]_  & \new_[40601]_ ;
  assign \new_[40611]_  = ~A236 & ~A235;
  assign \new_[40612]_  = ~A233 & \new_[40611]_ ;
  assign \new_[40615]_  = ~A267 & ~A266;
  assign \new_[40618]_  = A299 & ~A298;
  assign \new_[40619]_  = \new_[40618]_  & \new_[40615]_ ;
  assign \new_[40620]_  = \new_[40619]_  & \new_[40612]_ ;
  assign \new_[40624]_  = ~A167 & ~A169;
  assign \new_[40625]_  = A170 & \new_[40624]_ ;
  assign \new_[40629]_  = A200 & A199;
  assign \new_[40630]_  = A166 & \new_[40629]_ ;
  assign \new_[40631]_  = \new_[40630]_  & \new_[40625]_ ;
  assign \new_[40635]_  = ~A236 & ~A235;
  assign \new_[40636]_  = ~A233 & \new_[40635]_ ;
  assign \new_[40639]_  = ~A266 & ~A265;
  assign \new_[40642]_  = A299 & ~A298;
  assign \new_[40643]_  = \new_[40642]_  & \new_[40639]_ ;
  assign \new_[40644]_  = \new_[40643]_  & \new_[40636]_ ;
  assign \new_[40648]_  = ~A167 & ~A169;
  assign \new_[40649]_  = A170 & \new_[40648]_ ;
  assign \new_[40653]_  = A200 & A199;
  assign \new_[40654]_  = A166 & \new_[40653]_ ;
  assign \new_[40655]_  = \new_[40654]_  & \new_[40649]_ ;
  assign \new_[40659]_  = ~A266 & ~A234;
  assign \new_[40660]_  = ~A233 & \new_[40659]_ ;
  assign \new_[40663]_  = ~A269 & ~A268;
  assign \new_[40666]_  = A299 & ~A298;
  assign \new_[40667]_  = \new_[40666]_  & \new_[40663]_ ;
  assign \new_[40668]_  = \new_[40667]_  & \new_[40660]_ ;
  assign \new_[40672]_  = ~A167 & ~A169;
  assign \new_[40673]_  = A170 & \new_[40672]_ ;
  assign \new_[40677]_  = A200 & A199;
  assign \new_[40678]_  = A166 & \new_[40677]_ ;
  assign \new_[40679]_  = \new_[40678]_  & \new_[40673]_ ;
  assign \new_[40683]_  = A234 & ~A233;
  assign \new_[40684]_  = A232 & \new_[40683]_ ;
  assign \new_[40687]_  = A298 & A235;
  assign \new_[40690]_  = ~A302 & ~A301;
  assign \new_[40691]_  = \new_[40690]_  & \new_[40687]_ ;
  assign \new_[40692]_  = \new_[40691]_  & \new_[40684]_ ;
  assign \new_[40696]_  = ~A167 & ~A169;
  assign \new_[40697]_  = A170 & \new_[40696]_ ;
  assign \new_[40701]_  = A200 & A199;
  assign \new_[40702]_  = A166 & \new_[40701]_ ;
  assign \new_[40703]_  = \new_[40702]_  & \new_[40697]_ ;
  assign \new_[40707]_  = A234 & ~A233;
  assign \new_[40708]_  = A232 & \new_[40707]_ ;
  assign \new_[40711]_  = A298 & A236;
  assign \new_[40714]_  = ~A302 & ~A301;
  assign \new_[40715]_  = \new_[40714]_  & \new_[40711]_ ;
  assign \new_[40716]_  = \new_[40715]_  & \new_[40708]_ ;
  assign \new_[40720]_  = ~A167 & ~A169;
  assign \new_[40721]_  = A170 & \new_[40720]_ ;
  assign \new_[40725]_  = A200 & A199;
  assign \new_[40726]_  = A166 & \new_[40725]_ ;
  assign \new_[40727]_  = \new_[40726]_  & \new_[40721]_ ;
  assign \new_[40731]_  = ~A266 & ~A233;
  assign \new_[40732]_  = ~A232 & \new_[40731]_ ;
  assign \new_[40735]_  = ~A269 & ~A268;
  assign \new_[40738]_  = A299 & ~A298;
  assign \new_[40739]_  = \new_[40738]_  & \new_[40735]_ ;
  assign \new_[40740]_  = \new_[40739]_  & \new_[40732]_ ;
  assign \new_[40744]_  = ~A167 & ~A169;
  assign \new_[40745]_  = A170 & \new_[40744]_ ;
  assign \new_[40749]_  = ~A202 & ~A200;
  assign \new_[40750]_  = A166 & \new_[40749]_ ;
  assign \new_[40751]_  = \new_[40750]_  & \new_[40745]_ ;
  assign \new_[40755]_  = A233 & A232;
  assign \new_[40756]_  = ~A203 & \new_[40755]_ ;
  assign \new_[40759]_  = ~A267 & A265;
  assign \new_[40762]_  = A299 & ~A298;
  assign \new_[40763]_  = \new_[40762]_  & \new_[40759]_ ;
  assign \new_[40764]_  = \new_[40763]_  & \new_[40756]_ ;
  assign \new_[40768]_  = ~A167 & ~A169;
  assign \new_[40769]_  = A170 & \new_[40768]_ ;
  assign \new_[40773]_  = ~A202 & ~A200;
  assign \new_[40774]_  = A166 & \new_[40773]_ ;
  assign \new_[40775]_  = \new_[40774]_  & \new_[40769]_ ;
  assign \new_[40779]_  = A233 & A232;
  assign \new_[40780]_  = ~A203 & \new_[40779]_ ;
  assign \new_[40783]_  = A266 & A265;
  assign \new_[40786]_  = A299 & ~A298;
  assign \new_[40787]_  = \new_[40786]_  & \new_[40783]_ ;
  assign \new_[40788]_  = \new_[40787]_  & \new_[40780]_ ;
  assign \new_[40792]_  = ~A167 & ~A169;
  assign \new_[40793]_  = A170 & \new_[40792]_ ;
  assign \new_[40797]_  = ~A202 & ~A200;
  assign \new_[40798]_  = A166 & \new_[40797]_ ;
  assign \new_[40799]_  = \new_[40798]_  & \new_[40793]_ ;
  assign \new_[40803]_  = A233 & A232;
  assign \new_[40804]_  = ~A203 & \new_[40803]_ ;
  assign \new_[40807]_  = ~A266 & ~A265;
  assign \new_[40810]_  = A299 & ~A298;
  assign \new_[40811]_  = \new_[40810]_  & \new_[40807]_ ;
  assign \new_[40812]_  = \new_[40811]_  & \new_[40804]_ ;
  assign \new_[40816]_  = ~A167 & ~A169;
  assign \new_[40817]_  = A170 & \new_[40816]_ ;
  assign \new_[40821]_  = ~A202 & ~A200;
  assign \new_[40822]_  = A166 & \new_[40821]_ ;
  assign \new_[40823]_  = \new_[40822]_  & \new_[40817]_ ;
  assign \new_[40827]_  = A233 & ~A232;
  assign \new_[40828]_  = ~A203 & \new_[40827]_ ;
  assign \new_[40831]_  = ~A266 & A265;
  assign \new_[40834]_  = A268 & A267;
  assign \new_[40835]_  = \new_[40834]_  & \new_[40831]_ ;
  assign \new_[40836]_  = \new_[40835]_  & \new_[40828]_ ;
  assign \new_[40840]_  = ~A167 & ~A169;
  assign \new_[40841]_  = A170 & \new_[40840]_ ;
  assign \new_[40845]_  = ~A202 & ~A200;
  assign \new_[40846]_  = A166 & \new_[40845]_ ;
  assign \new_[40847]_  = \new_[40846]_  & \new_[40841]_ ;
  assign \new_[40851]_  = A233 & ~A232;
  assign \new_[40852]_  = ~A203 & \new_[40851]_ ;
  assign \new_[40855]_  = ~A266 & A265;
  assign \new_[40858]_  = A269 & A267;
  assign \new_[40859]_  = \new_[40858]_  & \new_[40855]_ ;
  assign \new_[40860]_  = \new_[40859]_  & \new_[40852]_ ;
  assign \new_[40864]_  = ~A167 & ~A169;
  assign \new_[40865]_  = A170 & \new_[40864]_ ;
  assign \new_[40869]_  = ~A202 & ~A200;
  assign \new_[40870]_  = A166 & \new_[40869]_ ;
  assign \new_[40871]_  = \new_[40870]_  & \new_[40865]_ ;
  assign \new_[40875]_  = ~A234 & ~A233;
  assign \new_[40876]_  = ~A203 & \new_[40875]_ ;
  assign \new_[40879]_  = A266 & A265;
  assign \new_[40882]_  = A299 & ~A298;
  assign \new_[40883]_  = \new_[40882]_  & \new_[40879]_ ;
  assign \new_[40884]_  = \new_[40883]_  & \new_[40876]_ ;
  assign \new_[40888]_  = ~A167 & ~A169;
  assign \new_[40889]_  = A170 & \new_[40888]_ ;
  assign \new_[40893]_  = ~A202 & ~A200;
  assign \new_[40894]_  = A166 & \new_[40893]_ ;
  assign \new_[40895]_  = \new_[40894]_  & \new_[40889]_ ;
  assign \new_[40899]_  = ~A234 & ~A233;
  assign \new_[40900]_  = ~A203 & \new_[40899]_ ;
  assign \new_[40903]_  = ~A267 & ~A266;
  assign \new_[40906]_  = A299 & ~A298;
  assign \new_[40907]_  = \new_[40906]_  & \new_[40903]_ ;
  assign \new_[40908]_  = \new_[40907]_  & \new_[40900]_ ;
  assign \new_[40912]_  = ~A167 & ~A169;
  assign \new_[40913]_  = A170 & \new_[40912]_ ;
  assign \new_[40917]_  = ~A202 & ~A200;
  assign \new_[40918]_  = A166 & \new_[40917]_ ;
  assign \new_[40919]_  = \new_[40918]_  & \new_[40913]_ ;
  assign \new_[40923]_  = ~A234 & ~A233;
  assign \new_[40924]_  = ~A203 & \new_[40923]_ ;
  assign \new_[40927]_  = ~A266 & ~A265;
  assign \new_[40930]_  = A299 & ~A298;
  assign \new_[40931]_  = \new_[40930]_  & \new_[40927]_ ;
  assign \new_[40932]_  = \new_[40931]_  & \new_[40924]_ ;
  assign \new_[40936]_  = ~A167 & ~A169;
  assign \new_[40937]_  = A170 & \new_[40936]_ ;
  assign \new_[40941]_  = ~A202 & ~A200;
  assign \new_[40942]_  = A166 & \new_[40941]_ ;
  assign \new_[40943]_  = \new_[40942]_  & \new_[40937]_ ;
  assign \new_[40947]_  = ~A233 & A232;
  assign \new_[40948]_  = ~A203 & \new_[40947]_ ;
  assign \new_[40951]_  = A235 & A234;
  assign \new_[40954]_  = ~A300 & A298;
  assign \new_[40955]_  = \new_[40954]_  & \new_[40951]_ ;
  assign \new_[40956]_  = \new_[40955]_  & \new_[40948]_ ;
  assign \new_[40960]_  = ~A167 & ~A169;
  assign \new_[40961]_  = A170 & \new_[40960]_ ;
  assign \new_[40965]_  = ~A202 & ~A200;
  assign \new_[40966]_  = A166 & \new_[40965]_ ;
  assign \new_[40967]_  = \new_[40966]_  & \new_[40961]_ ;
  assign \new_[40971]_  = ~A233 & A232;
  assign \new_[40972]_  = ~A203 & \new_[40971]_ ;
  assign \new_[40975]_  = A235 & A234;
  assign \new_[40978]_  = A299 & A298;
  assign \new_[40979]_  = \new_[40978]_  & \new_[40975]_ ;
  assign \new_[40980]_  = \new_[40979]_  & \new_[40972]_ ;
  assign \new_[40984]_  = ~A167 & ~A169;
  assign \new_[40985]_  = A170 & \new_[40984]_ ;
  assign \new_[40989]_  = ~A202 & ~A200;
  assign \new_[40990]_  = A166 & \new_[40989]_ ;
  assign \new_[40991]_  = \new_[40990]_  & \new_[40985]_ ;
  assign \new_[40995]_  = ~A233 & A232;
  assign \new_[40996]_  = ~A203 & \new_[40995]_ ;
  assign \new_[40999]_  = A235 & A234;
  assign \new_[41002]_  = ~A299 & ~A298;
  assign \new_[41003]_  = \new_[41002]_  & \new_[40999]_ ;
  assign \new_[41004]_  = \new_[41003]_  & \new_[40996]_ ;
  assign \new_[41008]_  = ~A167 & ~A169;
  assign \new_[41009]_  = A170 & \new_[41008]_ ;
  assign \new_[41013]_  = ~A202 & ~A200;
  assign \new_[41014]_  = A166 & \new_[41013]_ ;
  assign \new_[41015]_  = \new_[41014]_  & \new_[41009]_ ;
  assign \new_[41019]_  = ~A233 & A232;
  assign \new_[41020]_  = ~A203 & \new_[41019]_ ;
  assign \new_[41023]_  = A235 & A234;
  assign \new_[41026]_  = A266 & ~A265;
  assign \new_[41027]_  = \new_[41026]_  & \new_[41023]_ ;
  assign \new_[41028]_  = \new_[41027]_  & \new_[41020]_ ;
  assign \new_[41032]_  = ~A167 & ~A169;
  assign \new_[41033]_  = A170 & \new_[41032]_ ;
  assign \new_[41037]_  = ~A202 & ~A200;
  assign \new_[41038]_  = A166 & \new_[41037]_ ;
  assign \new_[41039]_  = \new_[41038]_  & \new_[41033]_ ;
  assign \new_[41043]_  = ~A233 & A232;
  assign \new_[41044]_  = ~A203 & \new_[41043]_ ;
  assign \new_[41047]_  = A236 & A234;
  assign \new_[41050]_  = ~A300 & A298;
  assign \new_[41051]_  = \new_[41050]_  & \new_[41047]_ ;
  assign \new_[41052]_  = \new_[41051]_  & \new_[41044]_ ;
  assign \new_[41056]_  = ~A167 & ~A169;
  assign \new_[41057]_  = A170 & \new_[41056]_ ;
  assign \new_[41061]_  = ~A202 & ~A200;
  assign \new_[41062]_  = A166 & \new_[41061]_ ;
  assign \new_[41063]_  = \new_[41062]_  & \new_[41057]_ ;
  assign \new_[41067]_  = ~A233 & A232;
  assign \new_[41068]_  = ~A203 & \new_[41067]_ ;
  assign \new_[41071]_  = A236 & A234;
  assign \new_[41074]_  = A299 & A298;
  assign \new_[41075]_  = \new_[41074]_  & \new_[41071]_ ;
  assign \new_[41076]_  = \new_[41075]_  & \new_[41068]_ ;
  assign \new_[41080]_  = ~A167 & ~A169;
  assign \new_[41081]_  = A170 & \new_[41080]_ ;
  assign \new_[41085]_  = ~A202 & ~A200;
  assign \new_[41086]_  = A166 & \new_[41085]_ ;
  assign \new_[41087]_  = \new_[41086]_  & \new_[41081]_ ;
  assign \new_[41091]_  = ~A233 & A232;
  assign \new_[41092]_  = ~A203 & \new_[41091]_ ;
  assign \new_[41095]_  = A236 & A234;
  assign \new_[41098]_  = ~A299 & ~A298;
  assign \new_[41099]_  = \new_[41098]_  & \new_[41095]_ ;
  assign \new_[41100]_  = \new_[41099]_  & \new_[41092]_ ;
  assign \new_[41104]_  = ~A167 & ~A169;
  assign \new_[41105]_  = A170 & \new_[41104]_ ;
  assign \new_[41109]_  = ~A202 & ~A200;
  assign \new_[41110]_  = A166 & \new_[41109]_ ;
  assign \new_[41111]_  = \new_[41110]_  & \new_[41105]_ ;
  assign \new_[41115]_  = ~A233 & A232;
  assign \new_[41116]_  = ~A203 & \new_[41115]_ ;
  assign \new_[41119]_  = A236 & A234;
  assign \new_[41122]_  = A266 & ~A265;
  assign \new_[41123]_  = \new_[41122]_  & \new_[41119]_ ;
  assign \new_[41124]_  = \new_[41123]_  & \new_[41116]_ ;
  assign \new_[41128]_  = ~A167 & ~A169;
  assign \new_[41129]_  = A170 & \new_[41128]_ ;
  assign \new_[41133]_  = ~A202 & ~A200;
  assign \new_[41134]_  = A166 & \new_[41133]_ ;
  assign \new_[41135]_  = \new_[41134]_  & \new_[41129]_ ;
  assign \new_[41139]_  = ~A233 & ~A232;
  assign \new_[41140]_  = ~A203 & \new_[41139]_ ;
  assign \new_[41143]_  = A266 & A265;
  assign \new_[41146]_  = A299 & ~A298;
  assign \new_[41147]_  = \new_[41146]_  & \new_[41143]_ ;
  assign \new_[41148]_  = \new_[41147]_  & \new_[41140]_ ;
  assign \new_[41152]_  = ~A167 & ~A169;
  assign \new_[41153]_  = A170 & \new_[41152]_ ;
  assign \new_[41157]_  = ~A202 & ~A200;
  assign \new_[41158]_  = A166 & \new_[41157]_ ;
  assign \new_[41159]_  = \new_[41158]_  & \new_[41153]_ ;
  assign \new_[41163]_  = ~A233 & ~A232;
  assign \new_[41164]_  = ~A203 & \new_[41163]_ ;
  assign \new_[41167]_  = ~A267 & ~A266;
  assign \new_[41170]_  = A299 & ~A298;
  assign \new_[41171]_  = \new_[41170]_  & \new_[41167]_ ;
  assign \new_[41172]_  = \new_[41171]_  & \new_[41164]_ ;
  assign \new_[41176]_  = ~A167 & ~A169;
  assign \new_[41177]_  = A170 & \new_[41176]_ ;
  assign \new_[41181]_  = ~A202 & ~A200;
  assign \new_[41182]_  = A166 & \new_[41181]_ ;
  assign \new_[41183]_  = \new_[41182]_  & \new_[41177]_ ;
  assign \new_[41187]_  = ~A233 & ~A232;
  assign \new_[41188]_  = ~A203 & \new_[41187]_ ;
  assign \new_[41191]_  = ~A266 & ~A265;
  assign \new_[41194]_  = A299 & ~A298;
  assign \new_[41195]_  = \new_[41194]_  & \new_[41191]_ ;
  assign \new_[41196]_  = \new_[41195]_  & \new_[41188]_ ;
  assign \new_[41200]_  = ~A167 & ~A169;
  assign \new_[41201]_  = A170 & \new_[41200]_ ;
  assign \new_[41205]_  = ~A201 & ~A200;
  assign \new_[41206]_  = A166 & \new_[41205]_ ;
  assign \new_[41207]_  = \new_[41206]_  & \new_[41201]_ ;
  assign \new_[41211]_  = A265 & A233;
  assign \new_[41212]_  = A232 & \new_[41211]_ ;
  assign \new_[41215]_  = ~A269 & ~A268;
  assign \new_[41218]_  = A299 & ~A298;
  assign \new_[41219]_  = \new_[41218]_  & \new_[41215]_ ;
  assign \new_[41220]_  = \new_[41219]_  & \new_[41212]_ ;
  assign \new_[41224]_  = ~A167 & ~A169;
  assign \new_[41225]_  = A170 & \new_[41224]_ ;
  assign \new_[41229]_  = ~A201 & ~A200;
  assign \new_[41230]_  = A166 & \new_[41229]_ ;
  assign \new_[41231]_  = \new_[41230]_  & \new_[41225]_ ;
  assign \new_[41235]_  = ~A236 & ~A235;
  assign \new_[41236]_  = ~A233 & \new_[41235]_ ;
  assign \new_[41239]_  = A266 & A265;
  assign \new_[41242]_  = A299 & ~A298;
  assign \new_[41243]_  = \new_[41242]_  & \new_[41239]_ ;
  assign \new_[41244]_  = \new_[41243]_  & \new_[41236]_ ;
  assign \new_[41248]_  = ~A167 & ~A169;
  assign \new_[41249]_  = A170 & \new_[41248]_ ;
  assign \new_[41253]_  = ~A201 & ~A200;
  assign \new_[41254]_  = A166 & \new_[41253]_ ;
  assign \new_[41255]_  = \new_[41254]_  & \new_[41249]_ ;
  assign \new_[41259]_  = ~A236 & ~A235;
  assign \new_[41260]_  = ~A233 & \new_[41259]_ ;
  assign \new_[41263]_  = ~A267 & ~A266;
  assign \new_[41266]_  = A299 & ~A298;
  assign \new_[41267]_  = \new_[41266]_  & \new_[41263]_ ;
  assign \new_[41268]_  = \new_[41267]_  & \new_[41260]_ ;
  assign \new_[41272]_  = ~A167 & ~A169;
  assign \new_[41273]_  = A170 & \new_[41272]_ ;
  assign \new_[41277]_  = ~A201 & ~A200;
  assign \new_[41278]_  = A166 & \new_[41277]_ ;
  assign \new_[41279]_  = \new_[41278]_  & \new_[41273]_ ;
  assign \new_[41283]_  = ~A236 & ~A235;
  assign \new_[41284]_  = ~A233 & \new_[41283]_ ;
  assign \new_[41287]_  = ~A266 & ~A265;
  assign \new_[41290]_  = A299 & ~A298;
  assign \new_[41291]_  = \new_[41290]_  & \new_[41287]_ ;
  assign \new_[41292]_  = \new_[41291]_  & \new_[41284]_ ;
  assign \new_[41296]_  = ~A167 & ~A169;
  assign \new_[41297]_  = A170 & \new_[41296]_ ;
  assign \new_[41301]_  = ~A201 & ~A200;
  assign \new_[41302]_  = A166 & \new_[41301]_ ;
  assign \new_[41303]_  = \new_[41302]_  & \new_[41297]_ ;
  assign \new_[41307]_  = ~A266 & ~A234;
  assign \new_[41308]_  = ~A233 & \new_[41307]_ ;
  assign \new_[41311]_  = ~A269 & ~A268;
  assign \new_[41314]_  = A299 & ~A298;
  assign \new_[41315]_  = \new_[41314]_  & \new_[41311]_ ;
  assign \new_[41316]_  = \new_[41315]_  & \new_[41308]_ ;
  assign \new_[41320]_  = ~A167 & ~A169;
  assign \new_[41321]_  = A170 & \new_[41320]_ ;
  assign \new_[41325]_  = ~A201 & ~A200;
  assign \new_[41326]_  = A166 & \new_[41325]_ ;
  assign \new_[41327]_  = \new_[41326]_  & \new_[41321]_ ;
  assign \new_[41331]_  = A234 & ~A233;
  assign \new_[41332]_  = A232 & \new_[41331]_ ;
  assign \new_[41335]_  = A298 & A235;
  assign \new_[41338]_  = ~A302 & ~A301;
  assign \new_[41339]_  = \new_[41338]_  & \new_[41335]_ ;
  assign \new_[41340]_  = \new_[41339]_  & \new_[41332]_ ;
  assign \new_[41344]_  = ~A167 & ~A169;
  assign \new_[41345]_  = A170 & \new_[41344]_ ;
  assign \new_[41349]_  = ~A201 & ~A200;
  assign \new_[41350]_  = A166 & \new_[41349]_ ;
  assign \new_[41351]_  = \new_[41350]_  & \new_[41345]_ ;
  assign \new_[41355]_  = A234 & ~A233;
  assign \new_[41356]_  = A232 & \new_[41355]_ ;
  assign \new_[41359]_  = A298 & A236;
  assign \new_[41362]_  = ~A302 & ~A301;
  assign \new_[41363]_  = \new_[41362]_  & \new_[41359]_ ;
  assign \new_[41364]_  = \new_[41363]_  & \new_[41356]_ ;
  assign \new_[41368]_  = ~A167 & ~A169;
  assign \new_[41369]_  = A170 & \new_[41368]_ ;
  assign \new_[41373]_  = ~A201 & ~A200;
  assign \new_[41374]_  = A166 & \new_[41373]_ ;
  assign \new_[41375]_  = \new_[41374]_  & \new_[41369]_ ;
  assign \new_[41379]_  = ~A266 & ~A233;
  assign \new_[41380]_  = ~A232 & \new_[41379]_ ;
  assign \new_[41383]_  = ~A269 & ~A268;
  assign \new_[41386]_  = A299 & ~A298;
  assign \new_[41387]_  = \new_[41386]_  & \new_[41383]_ ;
  assign \new_[41388]_  = \new_[41387]_  & \new_[41380]_ ;
  assign \new_[41392]_  = ~A167 & ~A169;
  assign \new_[41393]_  = A170 & \new_[41392]_ ;
  assign \new_[41397]_  = ~A200 & ~A199;
  assign \new_[41398]_  = A166 & \new_[41397]_ ;
  assign \new_[41399]_  = \new_[41398]_  & \new_[41393]_ ;
  assign \new_[41403]_  = A265 & A233;
  assign \new_[41404]_  = A232 & \new_[41403]_ ;
  assign \new_[41407]_  = ~A269 & ~A268;
  assign \new_[41410]_  = A299 & ~A298;
  assign \new_[41411]_  = \new_[41410]_  & \new_[41407]_ ;
  assign \new_[41412]_  = \new_[41411]_  & \new_[41404]_ ;
  assign \new_[41416]_  = ~A167 & ~A169;
  assign \new_[41417]_  = A170 & \new_[41416]_ ;
  assign \new_[41421]_  = ~A200 & ~A199;
  assign \new_[41422]_  = A166 & \new_[41421]_ ;
  assign \new_[41423]_  = \new_[41422]_  & \new_[41417]_ ;
  assign \new_[41427]_  = ~A236 & ~A235;
  assign \new_[41428]_  = ~A233 & \new_[41427]_ ;
  assign \new_[41431]_  = A266 & A265;
  assign \new_[41434]_  = A299 & ~A298;
  assign \new_[41435]_  = \new_[41434]_  & \new_[41431]_ ;
  assign \new_[41436]_  = \new_[41435]_  & \new_[41428]_ ;
  assign \new_[41440]_  = ~A167 & ~A169;
  assign \new_[41441]_  = A170 & \new_[41440]_ ;
  assign \new_[41445]_  = ~A200 & ~A199;
  assign \new_[41446]_  = A166 & \new_[41445]_ ;
  assign \new_[41447]_  = \new_[41446]_  & \new_[41441]_ ;
  assign \new_[41451]_  = ~A236 & ~A235;
  assign \new_[41452]_  = ~A233 & \new_[41451]_ ;
  assign \new_[41455]_  = ~A267 & ~A266;
  assign \new_[41458]_  = A299 & ~A298;
  assign \new_[41459]_  = \new_[41458]_  & \new_[41455]_ ;
  assign \new_[41460]_  = \new_[41459]_  & \new_[41452]_ ;
  assign \new_[41464]_  = ~A167 & ~A169;
  assign \new_[41465]_  = A170 & \new_[41464]_ ;
  assign \new_[41469]_  = ~A200 & ~A199;
  assign \new_[41470]_  = A166 & \new_[41469]_ ;
  assign \new_[41471]_  = \new_[41470]_  & \new_[41465]_ ;
  assign \new_[41475]_  = ~A236 & ~A235;
  assign \new_[41476]_  = ~A233 & \new_[41475]_ ;
  assign \new_[41479]_  = ~A266 & ~A265;
  assign \new_[41482]_  = A299 & ~A298;
  assign \new_[41483]_  = \new_[41482]_  & \new_[41479]_ ;
  assign \new_[41484]_  = \new_[41483]_  & \new_[41476]_ ;
  assign \new_[41488]_  = ~A167 & ~A169;
  assign \new_[41489]_  = A170 & \new_[41488]_ ;
  assign \new_[41493]_  = ~A200 & ~A199;
  assign \new_[41494]_  = A166 & \new_[41493]_ ;
  assign \new_[41495]_  = \new_[41494]_  & \new_[41489]_ ;
  assign \new_[41499]_  = ~A266 & ~A234;
  assign \new_[41500]_  = ~A233 & \new_[41499]_ ;
  assign \new_[41503]_  = ~A269 & ~A268;
  assign \new_[41506]_  = A299 & ~A298;
  assign \new_[41507]_  = \new_[41506]_  & \new_[41503]_ ;
  assign \new_[41508]_  = \new_[41507]_  & \new_[41500]_ ;
  assign \new_[41512]_  = ~A167 & ~A169;
  assign \new_[41513]_  = A170 & \new_[41512]_ ;
  assign \new_[41517]_  = ~A200 & ~A199;
  assign \new_[41518]_  = A166 & \new_[41517]_ ;
  assign \new_[41519]_  = \new_[41518]_  & \new_[41513]_ ;
  assign \new_[41523]_  = A234 & ~A233;
  assign \new_[41524]_  = A232 & \new_[41523]_ ;
  assign \new_[41527]_  = A298 & A235;
  assign \new_[41530]_  = ~A302 & ~A301;
  assign \new_[41531]_  = \new_[41530]_  & \new_[41527]_ ;
  assign \new_[41532]_  = \new_[41531]_  & \new_[41524]_ ;
  assign \new_[41536]_  = ~A167 & ~A169;
  assign \new_[41537]_  = A170 & \new_[41536]_ ;
  assign \new_[41541]_  = ~A200 & ~A199;
  assign \new_[41542]_  = A166 & \new_[41541]_ ;
  assign \new_[41543]_  = \new_[41542]_  & \new_[41537]_ ;
  assign \new_[41547]_  = A234 & ~A233;
  assign \new_[41548]_  = A232 & \new_[41547]_ ;
  assign \new_[41551]_  = A298 & A236;
  assign \new_[41554]_  = ~A302 & ~A301;
  assign \new_[41555]_  = \new_[41554]_  & \new_[41551]_ ;
  assign \new_[41556]_  = \new_[41555]_  & \new_[41548]_ ;
  assign \new_[41560]_  = ~A167 & ~A169;
  assign \new_[41561]_  = A170 & \new_[41560]_ ;
  assign \new_[41565]_  = ~A200 & ~A199;
  assign \new_[41566]_  = A166 & \new_[41565]_ ;
  assign \new_[41567]_  = \new_[41566]_  & \new_[41561]_ ;
  assign \new_[41571]_  = ~A266 & ~A233;
  assign \new_[41572]_  = ~A232 & \new_[41571]_ ;
  assign \new_[41575]_  = ~A269 & ~A268;
  assign \new_[41578]_  = A299 & ~A298;
  assign \new_[41579]_  = \new_[41578]_  & \new_[41575]_ ;
  assign \new_[41580]_  = \new_[41579]_  & \new_[41572]_ ;
  assign \new_[41584]_  = ~A168 & ~A169;
  assign \new_[41585]_  = ~A170 & \new_[41584]_ ;
  assign \new_[41589]_  = A201 & ~A200;
  assign \new_[41590]_  = A199 & \new_[41589]_ ;
  assign \new_[41591]_  = \new_[41590]_  & \new_[41585]_ ;
  assign \new_[41595]_  = A233 & A232;
  assign \new_[41596]_  = A202 & \new_[41595]_ ;
  assign \new_[41599]_  = ~A267 & A265;
  assign \new_[41602]_  = A299 & ~A298;
  assign \new_[41603]_  = \new_[41602]_  & \new_[41599]_ ;
  assign \new_[41604]_  = \new_[41603]_  & \new_[41596]_ ;
  assign \new_[41608]_  = ~A168 & ~A169;
  assign \new_[41609]_  = ~A170 & \new_[41608]_ ;
  assign \new_[41613]_  = A201 & ~A200;
  assign \new_[41614]_  = A199 & \new_[41613]_ ;
  assign \new_[41615]_  = \new_[41614]_  & \new_[41609]_ ;
  assign \new_[41619]_  = A233 & A232;
  assign \new_[41620]_  = A202 & \new_[41619]_ ;
  assign \new_[41623]_  = A266 & A265;
  assign \new_[41626]_  = A299 & ~A298;
  assign \new_[41627]_  = \new_[41626]_  & \new_[41623]_ ;
  assign \new_[41628]_  = \new_[41627]_  & \new_[41620]_ ;
  assign \new_[41632]_  = ~A168 & ~A169;
  assign \new_[41633]_  = ~A170 & \new_[41632]_ ;
  assign \new_[41637]_  = A201 & ~A200;
  assign \new_[41638]_  = A199 & \new_[41637]_ ;
  assign \new_[41639]_  = \new_[41638]_  & \new_[41633]_ ;
  assign \new_[41643]_  = A233 & A232;
  assign \new_[41644]_  = A202 & \new_[41643]_ ;
  assign \new_[41647]_  = ~A266 & ~A265;
  assign \new_[41650]_  = A299 & ~A298;
  assign \new_[41651]_  = \new_[41650]_  & \new_[41647]_ ;
  assign \new_[41652]_  = \new_[41651]_  & \new_[41644]_ ;
  assign \new_[41656]_  = ~A168 & ~A169;
  assign \new_[41657]_  = ~A170 & \new_[41656]_ ;
  assign \new_[41661]_  = A201 & ~A200;
  assign \new_[41662]_  = A199 & \new_[41661]_ ;
  assign \new_[41663]_  = \new_[41662]_  & \new_[41657]_ ;
  assign \new_[41667]_  = A233 & ~A232;
  assign \new_[41668]_  = A202 & \new_[41667]_ ;
  assign \new_[41671]_  = ~A266 & A265;
  assign \new_[41674]_  = A268 & A267;
  assign \new_[41675]_  = \new_[41674]_  & \new_[41671]_ ;
  assign \new_[41676]_  = \new_[41675]_  & \new_[41668]_ ;
  assign \new_[41680]_  = ~A168 & ~A169;
  assign \new_[41681]_  = ~A170 & \new_[41680]_ ;
  assign \new_[41685]_  = A201 & ~A200;
  assign \new_[41686]_  = A199 & \new_[41685]_ ;
  assign \new_[41687]_  = \new_[41686]_  & \new_[41681]_ ;
  assign \new_[41691]_  = A233 & ~A232;
  assign \new_[41692]_  = A202 & \new_[41691]_ ;
  assign \new_[41695]_  = ~A266 & A265;
  assign \new_[41698]_  = A269 & A267;
  assign \new_[41699]_  = \new_[41698]_  & \new_[41695]_ ;
  assign \new_[41700]_  = \new_[41699]_  & \new_[41692]_ ;
  assign \new_[41704]_  = ~A168 & ~A169;
  assign \new_[41705]_  = ~A170 & \new_[41704]_ ;
  assign \new_[41709]_  = A201 & ~A200;
  assign \new_[41710]_  = A199 & \new_[41709]_ ;
  assign \new_[41711]_  = \new_[41710]_  & \new_[41705]_ ;
  assign \new_[41715]_  = ~A234 & ~A233;
  assign \new_[41716]_  = A202 & \new_[41715]_ ;
  assign \new_[41719]_  = A266 & A265;
  assign \new_[41722]_  = A299 & ~A298;
  assign \new_[41723]_  = \new_[41722]_  & \new_[41719]_ ;
  assign \new_[41724]_  = \new_[41723]_  & \new_[41716]_ ;
  assign \new_[41728]_  = ~A168 & ~A169;
  assign \new_[41729]_  = ~A170 & \new_[41728]_ ;
  assign \new_[41733]_  = A201 & ~A200;
  assign \new_[41734]_  = A199 & \new_[41733]_ ;
  assign \new_[41735]_  = \new_[41734]_  & \new_[41729]_ ;
  assign \new_[41739]_  = ~A234 & ~A233;
  assign \new_[41740]_  = A202 & \new_[41739]_ ;
  assign \new_[41743]_  = ~A267 & ~A266;
  assign \new_[41746]_  = A299 & ~A298;
  assign \new_[41747]_  = \new_[41746]_  & \new_[41743]_ ;
  assign \new_[41748]_  = \new_[41747]_  & \new_[41740]_ ;
  assign \new_[41752]_  = ~A168 & ~A169;
  assign \new_[41753]_  = ~A170 & \new_[41752]_ ;
  assign \new_[41757]_  = A201 & ~A200;
  assign \new_[41758]_  = A199 & \new_[41757]_ ;
  assign \new_[41759]_  = \new_[41758]_  & \new_[41753]_ ;
  assign \new_[41763]_  = ~A234 & ~A233;
  assign \new_[41764]_  = A202 & \new_[41763]_ ;
  assign \new_[41767]_  = ~A266 & ~A265;
  assign \new_[41770]_  = A299 & ~A298;
  assign \new_[41771]_  = \new_[41770]_  & \new_[41767]_ ;
  assign \new_[41772]_  = \new_[41771]_  & \new_[41764]_ ;
  assign \new_[41776]_  = ~A168 & ~A169;
  assign \new_[41777]_  = ~A170 & \new_[41776]_ ;
  assign \new_[41781]_  = A201 & ~A200;
  assign \new_[41782]_  = A199 & \new_[41781]_ ;
  assign \new_[41783]_  = \new_[41782]_  & \new_[41777]_ ;
  assign \new_[41787]_  = ~A233 & A232;
  assign \new_[41788]_  = A202 & \new_[41787]_ ;
  assign \new_[41791]_  = A235 & A234;
  assign \new_[41794]_  = ~A300 & A298;
  assign \new_[41795]_  = \new_[41794]_  & \new_[41791]_ ;
  assign \new_[41796]_  = \new_[41795]_  & \new_[41788]_ ;
  assign \new_[41800]_  = ~A168 & ~A169;
  assign \new_[41801]_  = ~A170 & \new_[41800]_ ;
  assign \new_[41805]_  = A201 & ~A200;
  assign \new_[41806]_  = A199 & \new_[41805]_ ;
  assign \new_[41807]_  = \new_[41806]_  & \new_[41801]_ ;
  assign \new_[41811]_  = ~A233 & A232;
  assign \new_[41812]_  = A202 & \new_[41811]_ ;
  assign \new_[41815]_  = A235 & A234;
  assign \new_[41818]_  = A299 & A298;
  assign \new_[41819]_  = \new_[41818]_  & \new_[41815]_ ;
  assign \new_[41820]_  = \new_[41819]_  & \new_[41812]_ ;
  assign \new_[41824]_  = ~A168 & ~A169;
  assign \new_[41825]_  = ~A170 & \new_[41824]_ ;
  assign \new_[41829]_  = A201 & ~A200;
  assign \new_[41830]_  = A199 & \new_[41829]_ ;
  assign \new_[41831]_  = \new_[41830]_  & \new_[41825]_ ;
  assign \new_[41835]_  = ~A233 & A232;
  assign \new_[41836]_  = A202 & \new_[41835]_ ;
  assign \new_[41839]_  = A235 & A234;
  assign \new_[41842]_  = ~A299 & ~A298;
  assign \new_[41843]_  = \new_[41842]_  & \new_[41839]_ ;
  assign \new_[41844]_  = \new_[41843]_  & \new_[41836]_ ;
  assign \new_[41848]_  = ~A168 & ~A169;
  assign \new_[41849]_  = ~A170 & \new_[41848]_ ;
  assign \new_[41853]_  = A201 & ~A200;
  assign \new_[41854]_  = A199 & \new_[41853]_ ;
  assign \new_[41855]_  = \new_[41854]_  & \new_[41849]_ ;
  assign \new_[41859]_  = ~A233 & A232;
  assign \new_[41860]_  = A202 & \new_[41859]_ ;
  assign \new_[41863]_  = A235 & A234;
  assign \new_[41866]_  = A266 & ~A265;
  assign \new_[41867]_  = \new_[41866]_  & \new_[41863]_ ;
  assign \new_[41868]_  = \new_[41867]_  & \new_[41860]_ ;
  assign \new_[41872]_  = ~A168 & ~A169;
  assign \new_[41873]_  = ~A170 & \new_[41872]_ ;
  assign \new_[41877]_  = A201 & ~A200;
  assign \new_[41878]_  = A199 & \new_[41877]_ ;
  assign \new_[41879]_  = \new_[41878]_  & \new_[41873]_ ;
  assign \new_[41883]_  = ~A233 & A232;
  assign \new_[41884]_  = A202 & \new_[41883]_ ;
  assign \new_[41887]_  = A236 & A234;
  assign \new_[41890]_  = ~A300 & A298;
  assign \new_[41891]_  = \new_[41890]_  & \new_[41887]_ ;
  assign \new_[41892]_  = \new_[41891]_  & \new_[41884]_ ;
  assign \new_[41896]_  = ~A168 & ~A169;
  assign \new_[41897]_  = ~A170 & \new_[41896]_ ;
  assign \new_[41901]_  = A201 & ~A200;
  assign \new_[41902]_  = A199 & \new_[41901]_ ;
  assign \new_[41903]_  = \new_[41902]_  & \new_[41897]_ ;
  assign \new_[41907]_  = ~A233 & A232;
  assign \new_[41908]_  = A202 & \new_[41907]_ ;
  assign \new_[41911]_  = A236 & A234;
  assign \new_[41914]_  = A299 & A298;
  assign \new_[41915]_  = \new_[41914]_  & \new_[41911]_ ;
  assign \new_[41916]_  = \new_[41915]_  & \new_[41908]_ ;
  assign \new_[41920]_  = ~A168 & ~A169;
  assign \new_[41921]_  = ~A170 & \new_[41920]_ ;
  assign \new_[41925]_  = A201 & ~A200;
  assign \new_[41926]_  = A199 & \new_[41925]_ ;
  assign \new_[41927]_  = \new_[41926]_  & \new_[41921]_ ;
  assign \new_[41931]_  = ~A233 & A232;
  assign \new_[41932]_  = A202 & \new_[41931]_ ;
  assign \new_[41935]_  = A236 & A234;
  assign \new_[41938]_  = ~A299 & ~A298;
  assign \new_[41939]_  = \new_[41938]_  & \new_[41935]_ ;
  assign \new_[41940]_  = \new_[41939]_  & \new_[41932]_ ;
  assign \new_[41944]_  = ~A168 & ~A169;
  assign \new_[41945]_  = ~A170 & \new_[41944]_ ;
  assign \new_[41949]_  = A201 & ~A200;
  assign \new_[41950]_  = A199 & \new_[41949]_ ;
  assign \new_[41951]_  = \new_[41950]_  & \new_[41945]_ ;
  assign \new_[41955]_  = ~A233 & A232;
  assign \new_[41956]_  = A202 & \new_[41955]_ ;
  assign \new_[41959]_  = A236 & A234;
  assign \new_[41962]_  = A266 & ~A265;
  assign \new_[41963]_  = \new_[41962]_  & \new_[41959]_ ;
  assign \new_[41964]_  = \new_[41963]_  & \new_[41956]_ ;
  assign \new_[41968]_  = ~A168 & ~A169;
  assign \new_[41969]_  = ~A170 & \new_[41968]_ ;
  assign \new_[41973]_  = A201 & ~A200;
  assign \new_[41974]_  = A199 & \new_[41973]_ ;
  assign \new_[41975]_  = \new_[41974]_  & \new_[41969]_ ;
  assign \new_[41979]_  = ~A233 & ~A232;
  assign \new_[41980]_  = A202 & \new_[41979]_ ;
  assign \new_[41983]_  = A266 & A265;
  assign \new_[41986]_  = A299 & ~A298;
  assign \new_[41987]_  = \new_[41986]_  & \new_[41983]_ ;
  assign \new_[41988]_  = \new_[41987]_  & \new_[41980]_ ;
  assign \new_[41992]_  = ~A168 & ~A169;
  assign \new_[41993]_  = ~A170 & \new_[41992]_ ;
  assign \new_[41997]_  = A201 & ~A200;
  assign \new_[41998]_  = A199 & \new_[41997]_ ;
  assign \new_[41999]_  = \new_[41998]_  & \new_[41993]_ ;
  assign \new_[42003]_  = ~A233 & ~A232;
  assign \new_[42004]_  = A202 & \new_[42003]_ ;
  assign \new_[42007]_  = ~A267 & ~A266;
  assign \new_[42010]_  = A299 & ~A298;
  assign \new_[42011]_  = \new_[42010]_  & \new_[42007]_ ;
  assign \new_[42012]_  = \new_[42011]_  & \new_[42004]_ ;
  assign \new_[42016]_  = ~A168 & ~A169;
  assign \new_[42017]_  = ~A170 & \new_[42016]_ ;
  assign \new_[42021]_  = A201 & ~A200;
  assign \new_[42022]_  = A199 & \new_[42021]_ ;
  assign \new_[42023]_  = \new_[42022]_  & \new_[42017]_ ;
  assign \new_[42027]_  = ~A233 & ~A232;
  assign \new_[42028]_  = A202 & \new_[42027]_ ;
  assign \new_[42031]_  = ~A266 & ~A265;
  assign \new_[42034]_  = A299 & ~A298;
  assign \new_[42035]_  = \new_[42034]_  & \new_[42031]_ ;
  assign \new_[42036]_  = \new_[42035]_  & \new_[42028]_ ;
  assign \new_[42040]_  = ~A168 & ~A169;
  assign \new_[42041]_  = ~A170 & \new_[42040]_ ;
  assign \new_[42045]_  = A201 & ~A200;
  assign \new_[42046]_  = A199 & \new_[42045]_ ;
  assign \new_[42047]_  = \new_[42046]_  & \new_[42041]_ ;
  assign \new_[42051]_  = A233 & A232;
  assign \new_[42052]_  = A203 & \new_[42051]_ ;
  assign \new_[42055]_  = ~A267 & A265;
  assign \new_[42058]_  = A299 & ~A298;
  assign \new_[42059]_  = \new_[42058]_  & \new_[42055]_ ;
  assign \new_[42060]_  = \new_[42059]_  & \new_[42052]_ ;
  assign \new_[42064]_  = ~A168 & ~A169;
  assign \new_[42065]_  = ~A170 & \new_[42064]_ ;
  assign \new_[42069]_  = A201 & ~A200;
  assign \new_[42070]_  = A199 & \new_[42069]_ ;
  assign \new_[42071]_  = \new_[42070]_  & \new_[42065]_ ;
  assign \new_[42075]_  = A233 & A232;
  assign \new_[42076]_  = A203 & \new_[42075]_ ;
  assign \new_[42079]_  = A266 & A265;
  assign \new_[42082]_  = A299 & ~A298;
  assign \new_[42083]_  = \new_[42082]_  & \new_[42079]_ ;
  assign \new_[42084]_  = \new_[42083]_  & \new_[42076]_ ;
  assign \new_[42088]_  = ~A168 & ~A169;
  assign \new_[42089]_  = ~A170 & \new_[42088]_ ;
  assign \new_[42093]_  = A201 & ~A200;
  assign \new_[42094]_  = A199 & \new_[42093]_ ;
  assign \new_[42095]_  = \new_[42094]_  & \new_[42089]_ ;
  assign \new_[42099]_  = A233 & A232;
  assign \new_[42100]_  = A203 & \new_[42099]_ ;
  assign \new_[42103]_  = ~A266 & ~A265;
  assign \new_[42106]_  = A299 & ~A298;
  assign \new_[42107]_  = \new_[42106]_  & \new_[42103]_ ;
  assign \new_[42108]_  = \new_[42107]_  & \new_[42100]_ ;
  assign \new_[42112]_  = ~A168 & ~A169;
  assign \new_[42113]_  = ~A170 & \new_[42112]_ ;
  assign \new_[42117]_  = A201 & ~A200;
  assign \new_[42118]_  = A199 & \new_[42117]_ ;
  assign \new_[42119]_  = \new_[42118]_  & \new_[42113]_ ;
  assign \new_[42123]_  = A233 & ~A232;
  assign \new_[42124]_  = A203 & \new_[42123]_ ;
  assign \new_[42127]_  = ~A266 & A265;
  assign \new_[42130]_  = A268 & A267;
  assign \new_[42131]_  = \new_[42130]_  & \new_[42127]_ ;
  assign \new_[42132]_  = \new_[42131]_  & \new_[42124]_ ;
  assign \new_[42136]_  = ~A168 & ~A169;
  assign \new_[42137]_  = ~A170 & \new_[42136]_ ;
  assign \new_[42141]_  = A201 & ~A200;
  assign \new_[42142]_  = A199 & \new_[42141]_ ;
  assign \new_[42143]_  = \new_[42142]_  & \new_[42137]_ ;
  assign \new_[42147]_  = A233 & ~A232;
  assign \new_[42148]_  = A203 & \new_[42147]_ ;
  assign \new_[42151]_  = ~A266 & A265;
  assign \new_[42154]_  = A269 & A267;
  assign \new_[42155]_  = \new_[42154]_  & \new_[42151]_ ;
  assign \new_[42156]_  = \new_[42155]_  & \new_[42148]_ ;
  assign \new_[42160]_  = ~A168 & ~A169;
  assign \new_[42161]_  = ~A170 & \new_[42160]_ ;
  assign \new_[42165]_  = A201 & ~A200;
  assign \new_[42166]_  = A199 & \new_[42165]_ ;
  assign \new_[42167]_  = \new_[42166]_  & \new_[42161]_ ;
  assign \new_[42171]_  = ~A234 & ~A233;
  assign \new_[42172]_  = A203 & \new_[42171]_ ;
  assign \new_[42175]_  = A266 & A265;
  assign \new_[42178]_  = A299 & ~A298;
  assign \new_[42179]_  = \new_[42178]_  & \new_[42175]_ ;
  assign \new_[42180]_  = \new_[42179]_  & \new_[42172]_ ;
  assign \new_[42184]_  = ~A168 & ~A169;
  assign \new_[42185]_  = ~A170 & \new_[42184]_ ;
  assign \new_[42189]_  = A201 & ~A200;
  assign \new_[42190]_  = A199 & \new_[42189]_ ;
  assign \new_[42191]_  = \new_[42190]_  & \new_[42185]_ ;
  assign \new_[42195]_  = ~A234 & ~A233;
  assign \new_[42196]_  = A203 & \new_[42195]_ ;
  assign \new_[42199]_  = ~A267 & ~A266;
  assign \new_[42202]_  = A299 & ~A298;
  assign \new_[42203]_  = \new_[42202]_  & \new_[42199]_ ;
  assign \new_[42204]_  = \new_[42203]_  & \new_[42196]_ ;
  assign \new_[42208]_  = ~A168 & ~A169;
  assign \new_[42209]_  = ~A170 & \new_[42208]_ ;
  assign \new_[42213]_  = A201 & ~A200;
  assign \new_[42214]_  = A199 & \new_[42213]_ ;
  assign \new_[42215]_  = \new_[42214]_  & \new_[42209]_ ;
  assign \new_[42219]_  = ~A234 & ~A233;
  assign \new_[42220]_  = A203 & \new_[42219]_ ;
  assign \new_[42223]_  = ~A266 & ~A265;
  assign \new_[42226]_  = A299 & ~A298;
  assign \new_[42227]_  = \new_[42226]_  & \new_[42223]_ ;
  assign \new_[42228]_  = \new_[42227]_  & \new_[42220]_ ;
  assign \new_[42232]_  = ~A168 & ~A169;
  assign \new_[42233]_  = ~A170 & \new_[42232]_ ;
  assign \new_[42237]_  = A201 & ~A200;
  assign \new_[42238]_  = A199 & \new_[42237]_ ;
  assign \new_[42239]_  = \new_[42238]_  & \new_[42233]_ ;
  assign \new_[42243]_  = ~A233 & A232;
  assign \new_[42244]_  = A203 & \new_[42243]_ ;
  assign \new_[42247]_  = A235 & A234;
  assign \new_[42250]_  = ~A300 & A298;
  assign \new_[42251]_  = \new_[42250]_  & \new_[42247]_ ;
  assign \new_[42252]_  = \new_[42251]_  & \new_[42244]_ ;
  assign \new_[42256]_  = ~A168 & ~A169;
  assign \new_[42257]_  = ~A170 & \new_[42256]_ ;
  assign \new_[42261]_  = A201 & ~A200;
  assign \new_[42262]_  = A199 & \new_[42261]_ ;
  assign \new_[42263]_  = \new_[42262]_  & \new_[42257]_ ;
  assign \new_[42267]_  = ~A233 & A232;
  assign \new_[42268]_  = A203 & \new_[42267]_ ;
  assign \new_[42271]_  = A235 & A234;
  assign \new_[42274]_  = A299 & A298;
  assign \new_[42275]_  = \new_[42274]_  & \new_[42271]_ ;
  assign \new_[42276]_  = \new_[42275]_  & \new_[42268]_ ;
  assign \new_[42280]_  = ~A168 & ~A169;
  assign \new_[42281]_  = ~A170 & \new_[42280]_ ;
  assign \new_[42285]_  = A201 & ~A200;
  assign \new_[42286]_  = A199 & \new_[42285]_ ;
  assign \new_[42287]_  = \new_[42286]_  & \new_[42281]_ ;
  assign \new_[42291]_  = ~A233 & A232;
  assign \new_[42292]_  = A203 & \new_[42291]_ ;
  assign \new_[42295]_  = A235 & A234;
  assign \new_[42298]_  = ~A299 & ~A298;
  assign \new_[42299]_  = \new_[42298]_  & \new_[42295]_ ;
  assign \new_[42300]_  = \new_[42299]_  & \new_[42292]_ ;
  assign \new_[42304]_  = ~A168 & ~A169;
  assign \new_[42305]_  = ~A170 & \new_[42304]_ ;
  assign \new_[42309]_  = A201 & ~A200;
  assign \new_[42310]_  = A199 & \new_[42309]_ ;
  assign \new_[42311]_  = \new_[42310]_  & \new_[42305]_ ;
  assign \new_[42315]_  = ~A233 & A232;
  assign \new_[42316]_  = A203 & \new_[42315]_ ;
  assign \new_[42319]_  = A235 & A234;
  assign \new_[42322]_  = A266 & ~A265;
  assign \new_[42323]_  = \new_[42322]_  & \new_[42319]_ ;
  assign \new_[42324]_  = \new_[42323]_  & \new_[42316]_ ;
  assign \new_[42328]_  = ~A168 & ~A169;
  assign \new_[42329]_  = ~A170 & \new_[42328]_ ;
  assign \new_[42333]_  = A201 & ~A200;
  assign \new_[42334]_  = A199 & \new_[42333]_ ;
  assign \new_[42335]_  = \new_[42334]_  & \new_[42329]_ ;
  assign \new_[42339]_  = ~A233 & A232;
  assign \new_[42340]_  = A203 & \new_[42339]_ ;
  assign \new_[42343]_  = A236 & A234;
  assign \new_[42346]_  = ~A300 & A298;
  assign \new_[42347]_  = \new_[42346]_  & \new_[42343]_ ;
  assign \new_[42348]_  = \new_[42347]_  & \new_[42340]_ ;
  assign \new_[42352]_  = ~A168 & ~A169;
  assign \new_[42353]_  = ~A170 & \new_[42352]_ ;
  assign \new_[42357]_  = A201 & ~A200;
  assign \new_[42358]_  = A199 & \new_[42357]_ ;
  assign \new_[42359]_  = \new_[42358]_  & \new_[42353]_ ;
  assign \new_[42363]_  = ~A233 & A232;
  assign \new_[42364]_  = A203 & \new_[42363]_ ;
  assign \new_[42367]_  = A236 & A234;
  assign \new_[42370]_  = A299 & A298;
  assign \new_[42371]_  = \new_[42370]_  & \new_[42367]_ ;
  assign \new_[42372]_  = \new_[42371]_  & \new_[42364]_ ;
  assign \new_[42376]_  = ~A168 & ~A169;
  assign \new_[42377]_  = ~A170 & \new_[42376]_ ;
  assign \new_[42381]_  = A201 & ~A200;
  assign \new_[42382]_  = A199 & \new_[42381]_ ;
  assign \new_[42383]_  = \new_[42382]_  & \new_[42377]_ ;
  assign \new_[42387]_  = ~A233 & A232;
  assign \new_[42388]_  = A203 & \new_[42387]_ ;
  assign \new_[42391]_  = A236 & A234;
  assign \new_[42394]_  = ~A299 & ~A298;
  assign \new_[42395]_  = \new_[42394]_  & \new_[42391]_ ;
  assign \new_[42396]_  = \new_[42395]_  & \new_[42388]_ ;
  assign \new_[42400]_  = ~A168 & ~A169;
  assign \new_[42401]_  = ~A170 & \new_[42400]_ ;
  assign \new_[42405]_  = A201 & ~A200;
  assign \new_[42406]_  = A199 & \new_[42405]_ ;
  assign \new_[42407]_  = \new_[42406]_  & \new_[42401]_ ;
  assign \new_[42411]_  = ~A233 & A232;
  assign \new_[42412]_  = A203 & \new_[42411]_ ;
  assign \new_[42415]_  = A236 & A234;
  assign \new_[42418]_  = A266 & ~A265;
  assign \new_[42419]_  = \new_[42418]_  & \new_[42415]_ ;
  assign \new_[42420]_  = \new_[42419]_  & \new_[42412]_ ;
  assign \new_[42424]_  = ~A168 & ~A169;
  assign \new_[42425]_  = ~A170 & \new_[42424]_ ;
  assign \new_[42429]_  = A201 & ~A200;
  assign \new_[42430]_  = A199 & \new_[42429]_ ;
  assign \new_[42431]_  = \new_[42430]_  & \new_[42425]_ ;
  assign \new_[42435]_  = ~A233 & ~A232;
  assign \new_[42436]_  = A203 & \new_[42435]_ ;
  assign \new_[42439]_  = A266 & A265;
  assign \new_[42442]_  = A299 & ~A298;
  assign \new_[42443]_  = \new_[42442]_  & \new_[42439]_ ;
  assign \new_[42444]_  = \new_[42443]_  & \new_[42436]_ ;
  assign \new_[42448]_  = ~A168 & ~A169;
  assign \new_[42449]_  = ~A170 & \new_[42448]_ ;
  assign \new_[42453]_  = A201 & ~A200;
  assign \new_[42454]_  = A199 & \new_[42453]_ ;
  assign \new_[42455]_  = \new_[42454]_  & \new_[42449]_ ;
  assign \new_[42459]_  = ~A233 & ~A232;
  assign \new_[42460]_  = A203 & \new_[42459]_ ;
  assign \new_[42463]_  = ~A267 & ~A266;
  assign \new_[42466]_  = A299 & ~A298;
  assign \new_[42467]_  = \new_[42466]_  & \new_[42463]_ ;
  assign \new_[42468]_  = \new_[42467]_  & \new_[42460]_ ;
  assign \new_[42472]_  = ~A168 & ~A169;
  assign \new_[42473]_  = ~A170 & \new_[42472]_ ;
  assign \new_[42477]_  = A201 & ~A200;
  assign \new_[42478]_  = A199 & \new_[42477]_ ;
  assign \new_[42479]_  = \new_[42478]_  & \new_[42473]_ ;
  assign \new_[42483]_  = ~A233 & ~A232;
  assign \new_[42484]_  = A203 & \new_[42483]_ ;
  assign \new_[42487]_  = ~A266 & ~A265;
  assign \new_[42490]_  = A299 & ~A298;
  assign \new_[42491]_  = \new_[42490]_  & \new_[42487]_ ;
  assign \new_[42492]_  = \new_[42491]_  & \new_[42484]_ ;
  assign \new_[42496]_  = A199 & A166;
  assign \new_[42497]_  = A168 & \new_[42496]_ ;
  assign \new_[42500]_  = ~A233 & A200;
  assign \new_[42503]_  = ~A236 & ~A235;
  assign \new_[42504]_  = \new_[42503]_  & \new_[42500]_ ;
  assign \new_[42505]_  = \new_[42504]_  & \new_[42497]_ ;
  assign \new_[42509]_  = ~A269 & ~A268;
  assign \new_[42510]_  = ~A266 & \new_[42509]_ ;
  assign \new_[42513]_  = ~A299 & A298;
  assign \new_[42516]_  = A301 & A300;
  assign \new_[42517]_  = \new_[42516]_  & \new_[42513]_ ;
  assign \new_[42518]_  = \new_[42517]_  & \new_[42510]_ ;
  assign \new_[42522]_  = A199 & A166;
  assign \new_[42523]_  = A168 & \new_[42522]_ ;
  assign \new_[42526]_  = ~A233 & A200;
  assign \new_[42529]_  = ~A236 & ~A235;
  assign \new_[42530]_  = \new_[42529]_  & \new_[42526]_ ;
  assign \new_[42531]_  = \new_[42530]_  & \new_[42523]_ ;
  assign \new_[42535]_  = ~A269 & ~A268;
  assign \new_[42536]_  = ~A266 & \new_[42535]_ ;
  assign \new_[42539]_  = ~A299 & A298;
  assign \new_[42542]_  = A302 & A300;
  assign \new_[42543]_  = \new_[42542]_  & \new_[42539]_ ;
  assign \new_[42544]_  = \new_[42543]_  & \new_[42536]_ ;
  assign \new_[42548]_  = ~A200 & A166;
  assign \new_[42549]_  = A168 & \new_[42548]_ ;
  assign \new_[42552]_  = ~A203 & ~A202;
  assign \new_[42555]_  = A233 & A232;
  assign \new_[42556]_  = \new_[42555]_  & \new_[42552]_ ;
  assign \new_[42557]_  = \new_[42556]_  & \new_[42549]_ ;
  assign \new_[42561]_  = ~A269 & ~A268;
  assign \new_[42562]_  = A265 & \new_[42561]_ ;
  assign \new_[42565]_  = ~A299 & A298;
  assign \new_[42568]_  = A301 & A300;
  assign \new_[42569]_  = \new_[42568]_  & \new_[42565]_ ;
  assign \new_[42570]_  = \new_[42569]_  & \new_[42562]_ ;
  assign \new_[42574]_  = ~A200 & A166;
  assign \new_[42575]_  = A168 & \new_[42574]_ ;
  assign \new_[42578]_  = ~A203 & ~A202;
  assign \new_[42581]_  = A233 & A232;
  assign \new_[42582]_  = \new_[42581]_  & \new_[42578]_ ;
  assign \new_[42583]_  = \new_[42582]_  & \new_[42575]_ ;
  assign \new_[42587]_  = ~A269 & ~A268;
  assign \new_[42588]_  = A265 & \new_[42587]_ ;
  assign \new_[42591]_  = ~A299 & A298;
  assign \new_[42594]_  = A302 & A300;
  assign \new_[42595]_  = \new_[42594]_  & \new_[42591]_ ;
  assign \new_[42596]_  = \new_[42595]_  & \new_[42588]_ ;
  assign \new_[42600]_  = ~A200 & A166;
  assign \new_[42601]_  = A168 & \new_[42600]_ ;
  assign \new_[42604]_  = ~A203 & ~A202;
  assign \new_[42607]_  = ~A235 & ~A233;
  assign \new_[42608]_  = \new_[42607]_  & \new_[42604]_ ;
  assign \new_[42609]_  = \new_[42608]_  & \new_[42601]_ ;
  assign \new_[42613]_  = A266 & A265;
  assign \new_[42614]_  = ~A236 & \new_[42613]_ ;
  assign \new_[42617]_  = ~A299 & A298;
  assign \new_[42620]_  = A301 & A300;
  assign \new_[42621]_  = \new_[42620]_  & \new_[42617]_ ;
  assign \new_[42622]_  = \new_[42621]_  & \new_[42614]_ ;
  assign \new_[42626]_  = ~A200 & A166;
  assign \new_[42627]_  = A168 & \new_[42626]_ ;
  assign \new_[42630]_  = ~A203 & ~A202;
  assign \new_[42633]_  = ~A235 & ~A233;
  assign \new_[42634]_  = \new_[42633]_  & \new_[42630]_ ;
  assign \new_[42635]_  = \new_[42634]_  & \new_[42627]_ ;
  assign \new_[42639]_  = A266 & A265;
  assign \new_[42640]_  = ~A236 & \new_[42639]_ ;
  assign \new_[42643]_  = ~A299 & A298;
  assign \new_[42646]_  = A302 & A300;
  assign \new_[42647]_  = \new_[42646]_  & \new_[42643]_ ;
  assign \new_[42648]_  = \new_[42647]_  & \new_[42640]_ ;
  assign \new_[42652]_  = ~A200 & A166;
  assign \new_[42653]_  = A168 & \new_[42652]_ ;
  assign \new_[42656]_  = ~A203 & ~A202;
  assign \new_[42659]_  = ~A235 & ~A233;
  assign \new_[42660]_  = \new_[42659]_  & \new_[42656]_ ;
  assign \new_[42661]_  = \new_[42660]_  & \new_[42653]_ ;
  assign \new_[42665]_  = ~A267 & ~A266;
  assign \new_[42666]_  = ~A236 & \new_[42665]_ ;
  assign \new_[42669]_  = ~A299 & A298;
  assign \new_[42672]_  = A301 & A300;
  assign \new_[42673]_  = \new_[42672]_  & \new_[42669]_ ;
  assign \new_[42674]_  = \new_[42673]_  & \new_[42666]_ ;
  assign \new_[42678]_  = ~A200 & A166;
  assign \new_[42679]_  = A168 & \new_[42678]_ ;
  assign \new_[42682]_  = ~A203 & ~A202;
  assign \new_[42685]_  = ~A235 & ~A233;
  assign \new_[42686]_  = \new_[42685]_  & \new_[42682]_ ;
  assign \new_[42687]_  = \new_[42686]_  & \new_[42679]_ ;
  assign \new_[42691]_  = ~A267 & ~A266;
  assign \new_[42692]_  = ~A236 & \new_[42691]_ ;
  assign \new_[42695]_  = ~A299 & A298;
  assign \new_[42698]_  = A302 & A300;
  assign \new_[42699]_  = \new_[42698]_  & \new_[42695]_ ;
  assign \new_[42700]_  = \new_[42699]_  & \new_[42692]_ ;
  assign \new_[42704]_  = ~A200 & A166;
  assign \new_[42705]_  = A168 & \new_[42704]_ ;
  assign \new_[42708]_  = ~A203 & ~A202;
  assign \new_[42711]_  = ~A235 & ~A233;
  assign \new_[42712]_  = \new_[42711]_  & \new_[42708]_ ;
  assign \new_[42713]_  = \new_[42712]_  & \new_[42705]_ ;
  assign \new_[42717]_  = ~A266 & ~A265;
  assign \new_[42718]_  = ~A236 & \new_[42717]_ ;
  assign \new_[42721]_  = ~A299 & A298;
  assign \new_[42724]_  = A301 & A300;
  assign \new_[42725]_  = \new_[42724]_  & \new_[42721]_ ;
  assign \new_[42726]_  = \new_[42725]_  & \new_[42718]_ ;
  assign \new_[42730]_  = ~A200 & A166;
  assign \new_[42731]_  = A168 & \new_[42730]_ ;
  assign \new_[42734]_  = ~A203 & ~A202;
  assign \new_[42737]_  = ~A235 & ~A233;
  assign \new_[42738]_  = \new_[42737]_  & \new_[42734]_ ;
  assign \new_[42739]_  = \new_[42738]_  & \new_[42731]_ ;
  assign \new_[42743]_  = ~A266 & ~A265;
  assign \new_[42744]_  = ~A236 & \new_[42743]_ ;
  assign \new_[42747]_  = ~A299 & A298;
  assign \new_[42750]_  = A302 & A300;
  assign \new_[42751]_  = \new_[42750]_  & \new_[42747]_ ;
  assign \new_[42752]_  = \new_[42751]_  & \new_[42744]_ ;
  assign \new_[42756]_  = ~A200 & A166;
  assign \new_[42757]_  = A168 & \new_[42756]_ ;
  assign \new_[42760]_  = ~A203 & ~A202;
  assign \new_[42763]_  = ~A234 & ~A233;
  assign \new_[42764]_  = \new_[42763]_  & \new_[42760]_ ;
  assign \new_[42765]_  = \new_[42764]_  & \new_[42757]_ ;
  assign \new_[42769]_  = ~A269 & ~A268;
  assign \new_[42770]_  = ~A266 & \new_[42769]_ ;
  assign \new_[42773]_  = ~A299 & A298;
  assign \new_[42776]_  = A301 & A300;
  assign \new_[42777]_  = \new_[42776]_  & \new_[42773]_ ;
  assign \new_[42778]_  = \new_[42777]_  & \new_[42770]_ ;
  assign \new_[42782]_  = ~A200 & A166;
  assign \new_[42783]_  = A168 & \new_[42782]_ ;
  assign \new_[42786]_  = ~A203 & ~A202;
  assign \new_[42789]_  = ~A234 & ~A233;
  assign \new_[42790]_  = \new_[42789]_  & \new_[42786]_ ;
  assign \new_[42791]_  = \new_[42790]_  & \new_[42783]_ ;
  assign \new_[42795]_  = ~A269 & ~A268;
  assign \new_[42796]_  = ~A266 & \new_[42795]_ ;
  assign \new_[42799]_  = ~A299 & A298;
  assign \new_[42802]_  = A302 & A300;
  assign \new_[42803]_  = \new_[42802]_  & \new_[42799]_ ;
  assign \new_[42804]_  = \new_[42803]_  & \new_[42796]_ ;
  assign \new_[42808]_  = ~A200 & A166;
  assign \new_[42809]_  = A168 & \new_[42808]_ ;
  assign \new_[42812]_  = ~A203 & ~A202;
  assign \new_[42815]_  = ~A233 & ~A232;
  assign \new_[42816]_  = \new_[42815]_  & \new_[42812]_ ;
  assign \new_[42817]_  = \new_[42816]_  & \new_[42809]_ ;
  assign \new_[42821]_  = ~A269 & ~A268;
  assign \new_[42822]_  = ~A266 & \new_[42821]_ ;
  assign \new_[42825]_  = ~A299 & A298;
  assign \new_[42828]_  = A301 & A300;
  assign \new_[42829]_  = \new_[42828]_  & \new_[42825]_ ;
  assign \new_[42830]_  = \new_[42829]_  & \new_[42822]_ ;
  assign \new_[42834]_  = ~A200 & A166;
  assign \new_[42835]_  = A168 & \new_[42834]_ ;
  assign \new_[42838]_  = ~A203 & ~A202;
  assign \new_[42841]_  = ~A233 & ~A232;
  assign \new_[42842]_  = \new_[42841]_  & \new_[42838]_ ;
  assign \new_[42843]_  = \new_[42842]_  & \new_[42835]_ ;
  assign \new_[42847]_  = ~A269 & ~A268;
  assign \new_[42848]_  = ~A266 & \new_[42847]_ ;
  assign \new_[42851]_  = ~A299 & A298;
  assign \new_[42854]_  = A302 & A300;
  assign \new_[42855]_  = \new_[42854]_  & \new_[42851]_ ;
  assign \new_[42856]_  = \new_[42855]_  & \new_[42848]_ ;
  assign \new_[42860]_  = ~A200 & A166;
  assign \new_[42861]_  = A168 & \new_[42860]_ ;
  assign \new_[42864]_  = ~A233 & ~A201;
  assign \new_[42867]_  = ~A236 & ~A235;
  assign \new_[42868]_  = \new_[42867]_  & \new_[42864]_ ;
  assign \new_[42869]_  = \new_[42868]_  & \new_[42861]_ ;
  assign \new_[42873]_  = ~A269 & ~A268;
  assign \new_[42874]_  = ~A266 & \new_[42873]_ ;
  assign \new_[42877]_  = ~A299 & A298;
  assign \new_[42880]_  = A301 & A300;
  assign \new_[42881]_  = \new_[42880]_  & \new_[42877]_ ;
  assign \new_[42882]_  = \new_[42881]_  & \new_[42874]_ ;
  assign \new_[42886]_  = ~A200 & A166;
  assign \new_[42887]_  = A168 & \new_[42886]_ ;
  assign \new_[42890]_  = ~A233 & ~A201;
  assign \new_[42893]_  = ~A236 & ~A235;
  assign \new_[42894]_  = \new_[42893]_  & \new_[42890]_ ;
  assign \new_[42895]_  = \new_[42894]_  & \new_[42887]_ ;
  assign \new_[42899]_  = ~A269 & ~A268;
  assign \new_[42900]_  = ~A266 & \new_[42899]_ ;
  assign \new_[42903]_  = ~A299 & A298;
  assign \new_[42906]_  = A302 & A300;
  assign \new_[42907]_  = \new_[42906]_  & \new_[42903]_ ;
  assign \new_[42908]_  = \new_[42907]_  & \new_[42900]_ ;
  assign \new_[42912]_  = ~A199 & A166;
  assign \new_[42913]_  = A168 & \new_[42912]_ ;
  assign \new_[42916]_  = ~A233 & ~A200;
  assign \new_[42919]_  = ~A236 & ~A235;
  assign \new_[42920]_  = \new_[42919]_  & \new_[42916]_ ;
  assign \new_[42921]_  = \new_[42920]_  & \new_[42913]_ ;
  assign \new_[42925]_  = ~A269 & ~A268;
  assign \new_[42926]_  = ~A266 & \new_[42925]_ ;
  assign \new_[42929]_  = ~A299 & A298;
  assign \new_[42932]_  = A301 & A300;
  assign \new_[42933]_  = \new_[42932]_  & \new_[42929]_ ;
  assign \new_[42934]_  = \new_[42933]_  & \new_[42926]_ ;
  assign \new_[42938]_  = ~A199 & A166;
  assign \new_[42939]_  = A168 & \new_[42938]_ ;
  assign \new_[42942]_  = ~A233 & ~A200;
  assign \new_[42945]_  = ~A236 & ~A235;
  assign \new_[42946]_  = \new_[42945]_  & \new_[42942]_ ;
  assign \new_[42947]_  = \new_[42946]_  & \new_[42939]_ ;
  assign \new_[42951]_  = ~A269 & ~A268;
  assign \new_[42952]_  = ~A266 & \new_[42951]_ ;
  assign \new_[42955]_  = ~A299 & A298;
  assign \new_[42958]_  = A302 & A300;
  assign \new_[42959]_  = \new_[42958]_  & \new_[42955]_ ;
  assign \new_[42960]_  = \new_[42959]_  & \new_[42952]_ ;
  assign \new_[42964]_  = A199 & A167;
  assign \new_[42965]_  = A168 & \new_[42964]_ ;
  assign \new_[42968]_  = ~A233 & A200;
  assign \new_[42971]_  = ~A236 & ~A235;
  assign \new_[42972]_  = \new_[42971]_  & \new_[42968]_ ;
  assign \new_[42973]_  = \new_[42972]_  & \new_[42965]_ ;
  assign \new_[42977]_  = ~A269 & ~A268;
  assign \new_[42978]_  = ~A266 & \new_[42977]_ ;
  assign \new_[42981]_  = ~A299 & A298;
  assign \new_[42984]_  = A301 & A300;
  assign \new_[42985]_  = \new_[42984]_  & \new_[42981]_ ;
  assign \new_[42986]_  = \new_[42985]_  & \new_[42978]_ ;
  assign \new_[42990]_  = A199 & A167;
  assign \new_[42991]_  = A168 & \new_[42990]_ ;
  assign \new_[42994]_  = ~A233 & A200;
  assign \new_[42997]_  = ~A236 & ~A235;
  assign \new_[42998]_  = \new_[42997]_  & \new_[42994]_ ;
  assign \new_[42999]_  = \new_[42998]_  & \new_[42991]_ ;
  assign \new_[43003]_  = ~A269 & ~A268;
  assign \new_[43004]_  = ~A266 & \new_[43003]_ ;
  assign \new_[43007]_  = ~A299 & A298;
  assign \new_[43010]_  = A302 & A300;
  assign \new_[43011]_  = \new_[43010]_  & \new_[43007]_ ;
  assign \new_[43012]_  = \new_[43011]_  & \new_[43004]_ ;
  assign \new_[43016]_  = ~A200 & A167;
  assign \new_[43017]_  = A168 & \new_[43016]_ ;
  assign \new_[43020]_  = ~A203 & ~A202;
  assign \new_[43023]_  = A233 & A232;
  assign \new_[43024]_  = \new_[43023]_  & \new_[43020]_ ;
  assign \new_[43025]_  = \new_[43024]_  & \new_[43017]_ ;
  assign \new_[43029]_  = ~A269 & ~A268;
  assign \new_[43030]_  = A265 & \new_[43029]_ ;
  assign \new_[43033]_  = ~A299 & A298;
  assign \new_[43036]_  = A301 & A300;
  assign \new_[43037]_  = \new_[43036]_  & \new_[43033]_ ;
  assign \new_[43038]_  = \new_[43037]_  & \new_[43030]_ ;
  assign \new_[43042]_  = ~A200 & A167;
  assign \new_[43043]_  = A168 & \new_[43042]_ ;
  assign \new_[43046]_  = ~A203 & ~A202;
  assign \new_[43049]_  = A233 & A232;
  assign \new_[43050]_  = \new_[43049]_  & \new_[43046]_ ;
  assign \new_[43051]_  = \new_[43050]_  & \new_[43043]_ ;
  assign \new_[43055]_  = ~A269 & ~A268;
  assign \new_[43056]_  = A265 & \new_[43055]_ ;
  assign \new_[43059]_  = ~A299 & A298;
  assign \new_[43062]_  = A302 & A300;
  assign \new_[43063]_  = \new_[43062]_  & \new_[43059]_ ;
  assign \new_[43064]_  = \new_[43063]_  & \new_[43056]_ ;
  assign \new_[43068]_  = ~A200 & A167;
  assign \new_[43069]_  = A168 & \new_[43068]_ ;
  assign \new_[43072]_  = ~A203 & ~A202;
  assign \new_[43075]_  = ~A235 & ~A233;
  assign \new_[43076]_  = \new_[43075]_  & \new_[43072]_ ;
  assign \new_[43077]_  = \new_[43076]_  & \new_[43069]_ ;
  assign \new_[43081]_  = A266 & A265;
  assign \new_[43082]_  = ~A236 & \new_[43081]_ ;
  assign \new_[43085]_  = ~A299 & A298;
  assign \new_[43088]_  = A301 & A300;
  assign \new_[43089]_  = \new_[43088]_  & \new_[43085]_ ;
  assign \new_[43090]_  = \new_[43089]_  & \new_[43082]_ ;
  assign \new_[43094]_  = ~A200 & A167;
  assign \new_[43095]_  = A168 & \new_[43094]_ ;
  assign \new_[43098]_  = ~A203 & ~A202;
  assign \new_[43101]_  = ~A235 & ~A233;
  assign \new_[43102]_  = \new_[43101]_  & \new_[43098]_ ;
  assign \new_[43103]_  = \new_[43102]_  & \new_[43095]_ ;
  assign \new_[43107]_  = A266 & A265;
  assign \new_[43108]_  = ~A236 & \new_[43107]_ ;
  assign \new_[43111]_  = ~A299 & A298;
  assign \new_[43114]_  = A302 & A300;
  assign \new_[43115]_  = \new_[43114]_  & \new_[43111]_ ;
  assign \new_[43116]_  = \new_[43115]_  & \new_[43108]_ ;
  assign \new_[43120]_  = ~A200 & A167;
  assign \new_[43121]_  = A168 & \new_[43120]_ ;
  assign \new_[43124]_  = ~A203 & ~A202;
  assign \new_[43127]_  = ~A235 & ~A233;
  assign \new_[43128]_  = \new_[43127]_  & \new_[43124]_ ;
  assign \new_[43129]_  = \new_[43128]_  & \new_[43121]_ ;
  assign \new_[43133]_  = ~A267 & ~A266;
  assign \new_[43134]_  = ~A236 & \new_[43133]_ ;
  assign \new_[43137]_  = ~A299 & A298;
  assign \new_[43140]_  = A301 & A300;
  assign \new_[43141]_  = \new_[43140]_  & \new_[43137]_ ;
  assign \new_[43142]_  = \new_[43141]_  & \new_[43134]_ ;
  assign \new_[43146]_  = ~A200 & A167;
  assign \new_[43147]_  = A168 & \new_[43146]_ ;
  assign \new_[43150]_  = ~A203 & ~A202;
  assign \new_[43153]_  = ~A235 & ~A233;
  assign \new_[43154]_  = \new_[43153]_  & \new_[43150]_ ;
  assign \new_[43155]_  = \new_[43154]_  & \new_[43147]_ ;
  assign \new_[43159]_  = ~A267 & ~A266;
  assign \new_[43160]_  = ~A236 & \new_[43159]_ ;
  assign \new_[43163]_  = ~A299 & A298;
  assign \new_[43166]_  = A302 & A300;
  assign \new_[43167]_  = \new_[43166]_  & \new_[43163]_ ;
  assign \new_[43168]_  = \new_[43167]_  & \new_[43160]_ ;
  assign \new_[43172]_  = ~A200 & A167;
  assign \new_[43173]_  = A168 & \new_[43172]_ ;
  assign \new_[43176]_  = ~A203 & ~A202;
  assign \new_[43179]_  = ~A235 & ~A233;
  assign \new_[43180]_  = \new_[43179]_  & \new_[43176]_ ;
  assign \new_[43181]_  = \new_[43180]_  & \new_[43173]_ ;
  assign \new_[43185]_  = ~A266 & ~A265;
  assign \new_[43186]_  = ~A236 & \new_[43185]_ ;
  assign \new_[43189]_  = ~A299 & A298;
  assign \new_[43192]_  = A301 & A300;
  assign \new_[43193]_  = \new_[43192]_  & \new_[43189]_ ;
  assign \new_[43194]_  = \new_[43193]_  & \new_[43186]_ ;
  assign \new_[43198]_  = ~A200 & A167;
  assign \new_[43199]_  = A168 & \new_[43198]_ ;
  assign \new_[43202]_  = ~A203 & ~A202;
  assign \new_[43205]_  = ~A235 & ~A233;
  assign \new_[43206]_  = \new_[43205]_  & \new_[43202]_ ;
  assign \new_[43207]_  = \new_[43206]_  & \new_[43199]_ ;
  assign \new_[43211]_  = ~A266 & ~A265;
  assign \new_[43212]_  = ~A236 & \new_[43211]_ ;
  assign \new_[43215]_  = ~A299 & A298;
  assign \new_[43218]_  = A302 & A300;
  assign \new_[43219]_  = \new_[43218]_  & \new_[43215]_ ;
  assign \new_[43220]_  = \new_[43219]_  & \new_[43212]_ ;
  assign \new_[43224]_  = ~A200 & A167;
  assign \new_[43225]_  = A168 & \new_[43224]_ ;
  assign \new_[43228]_  = ~A203 & ~A202;
  assign \new_[43231]_  = ~A234 & ~A233;
  assign \new_[43232]_  = \new_[43231]_  & \new_[43228]_ ;
  assign \new_[43233]_  = \new_[43232]_  & \new_[43225]_ ;
  assign \new_[43237]_  = ~A269 & ~A268;
  assign \new_[43238]_  = ~A266 & \new_[43237]_ ;
  assign \new_[43241]_  = ~A299 & A298;
  assign \new_[43244]_  = A301 & A300;
  assign \new_[43245]_  = \new_[43244]_  & \new_[43241]_ ;
  assign \new_[43246]_  = \new_[43245]_  & \new_[43238]_ ;
  assign \new_[43250]_  = ~A200 & A167;
  assign \new_[43251]_  = A168 & \new_[43250]_ ;
  assign \new_[43254]_  = ~A203 & ~A202;
  assign \new_[43257]_  = ~A234 & ~A233;
  assign \new_[43258]_  = \new_[43257]_  & \new_[43254]_ ;
  assign \new_[43259]_  = \new_[43258]_  & \new_[43251]_ ;
  assign \new_[43263]_  = ~A269 & ~A268;
  assign \new_[43264]_  = ~A266 & \new_[43263]_ ;
  assign \new_[43267]_  = ~A299 & A298;
  assign \new_[43270]_  = A302 & A300;
  assign \new_[43271]_  = \new_[43270]_  & \new_[43267]_ ;
  assign \new_[43272]_  = \new_[43271]_  & \new_[43264]_ ;
  assign \new_[43276]_  = ~A200 & A167;
  assign \new_[43277]_  = A168 & \new_[43276]_ ;
  assign \new_[43280]_  = ~A203 & ~A202;
  assign \new_[43283]_  = ~A233 & ~A232;
  assign \new_[43284]_  = \new_[43283]_  & \new_[43280]_ ;
  assign \new_[43285]_  = \new_[43284]_  & \new_[43277]_ ;
  assign \new_[43289]_  = ~A269 & ~A268;
  assign \new_[43290]_  = ~A266 & \new_[43289]_ ;
  assign \new_[43293]_  = ~A299 & A298;
  assign \new_[43296]_  = A301 & A300;
  assign \new_[43297]_  = \new_[43296]_  & \new_[43293]_ ;
  assign \new_[43298]_  = \new_[43297]_  & \new_[43290]_ ;
  assign \new_[43302]_  = ~A200 & A167;
  assign \new_[43303]_  = A168 & \new_[43302]_ ;
  assign \new_[43306]_  = ~A203 & ~A202;
  assign \new_[43309]_  = ~A233 & ~A232;
  assign \new_[43310]_  = \new_[43309]_  & \new_[43306]_ ;
  assign \new_[43311]_  = \new_[43310]_  & \new_[43303]_ ;
  assign \new_[43315]_  = ~A269 & ~A268;
  assign \new_[43316]_  = ~A266 & \new_[43315]_ ;
  assign \new_[43319]_  = ~A299 & A298;
  assign \new_[43322]_  = A302 & A300;
  assign \new_[43323]_  = \new_[43322]_  & \new_[43319]_ ;
  assign \new_[43324]_  = \new_[43323]_  & \new_[43316]_ ;
  assign \new_[43328]_  = ~A200 & A167;
  assign \new_[43329]_  = A168 & \new_[43328]_ ;
  assign \new_[43332]_  = ~A233 & ~A201;
  assign \new_[43335]_  = ~A236 & ~A235;
  assign \new_[43336]_  = \new_[43335]_  & \new_[43332]_ ;
  assign \new_[43337]_  = \new_[43336]_  & \new_[43329]_ ;
  assign \new_[43341]_  = ~A269 & ~A268;
  assign \new_[43342]_  = ~A266 & \new_[43341]_ ;
  assign \new_[43345]_  = ~A299 & A298;
  assign \new_[43348]_  = A301 & A300;
  assign \new_[43349]_  = \new_[43348]_  & \new_[43345]_ ;
  assign \new_[43350]_  = \new_[43349]_  & \new_[43342]_ ;
  assign \new_[43354]_  = ~A200 & A167;
  assign \new_[43355]_  = A168 & \new_[43354]_ ;
  assign \new_[43358]_  = ~A233 & ~A201;
  assign \new_[43361]_  = ~A236 & ~A235;
  assign \new_[43362]_  = \new_[43361]_  & \new_[43358]_ ;
  assign \new_[43363]_  = \new_[43362]_  & \new_[43355]_ ;
  assign \new_[43367]_  = ~A269 & ~A268;
  assign \new_[43368]_  = ~A266 & \new_[43367]_ ;
  assign \new_[43371]_  = ~A299 & A298;
  assign \new_[43374]_  = A302 & A300;
  assign \new_[43375]_  = \new_[43374]_  & \new_[43371]_ ;
  assign \new_[43376]_  = \new_[43375]_  & \new_[43368]_ ;
  assign \new_[43380]_  = ~A199 & A167;
  assign \new_[43381]_  = A168 & \new_[43380]_ ;
  assign \new_[43384]_  = ~A233 & ~A200;
  assign \new_[43387]_  = ~A236 & ~A235;
  assign \new_[43388]_  = \new_[43387]_  & \new_[43384]_ ;
  assign \new_[43389]_  = \new_[43388]_  & \new_[43381]_ ;
  assign \new_[43393]_  = ~A269 & ~A268;
  assign \new_[43394]_  = ~A266 & \new_[43393]_ ;
  assign \new_[43397]_  = ~A299 & A298;
  assign \new_[43400]_  = A301 & A300;
  assign \new_[43401]_  = \new_[43400]_  & \new_[43397]_ ;
  assign \new_[43402]_  = \new_[43401]_  & \new_[43394]_ ;
  assign \new_[43406]_  = ~A199 & A167;
  assign \new_[43407]_  = A168 & \new_[43406]_ ;
  assign \new_[43410]_  = ~A233 & ~A200;
  assign \new_[43413]_  = ~A236 & ~A235;
  assign \new_[43414]_  = \new_[43413]_  & \new_[43410]_ ;
  assign \new_[43415]_  = \new_[43414]_  & \new_[43407]_ ;
  assign \new_[43419]_  = ~A269 & ~A268;
  assign \new_[43420]_  = ~A266 & \new_[43419]_ ;
  assign \new_[43423]_  = ~A299 & A298;
  assign \new_[43426]_  = A302 & A300;
  assign \new_[43427]_  = \new_[43426]_  & \new_[43423]_ ;
  assign \new_[43428]_  = \new_[43427]_  & \new_[43420]_ ;
  assign \new_[43432]_  = ~A166 & ~A167;
  assign \new_[43433]_  = A170 & \new_[43432]_ ;
  assign \new_[43436]_  = A200 & ~A199;
  assign \new_[43439]_  = A233 & A232;
  assign \new_[43440]_  = \new_[43439]_  & \new_[43436]_ ;
  assign \new_[43441]_  = \new_[43440]_  & \new_[43433]_ ;
  assign \new_[43445]_  = ~A269 & ~A268;
  assign \new_[43446]_  = A265 & \new_[43445]_ ;
  assign \new_[43449]_  = ~A299 & A298;
  assign \new_[43452]_  = A301 & A300;
  assign \new_[43453]_  = \new_[43452]_  & \new_[43449]_ ;
  assign \new_[43454]_  = \new_[43453]_  & \new_[43446]_ ;
  assign \new_[43458]_  = ~A166 & ~A167;
  assign \new_[43459]_  = A170 & \new_[43458]_ ;
  assign \new_[43462]_  = A200 & ~A199;
  assign \new_[43465]_  = A233 & A232;
  assign \new_[43466]_  = \new_[43465]_  & \new_[43462]_ ;
  assign \new_[43467]_  = \new_[43466]_  & \new_[43459]_ ;
  assign \new_[43471]_  = ~A269 & ~A268;
  assign \new_[43472]_  = A265 & \new_[43471]_ ;
  assign \new_[43475]_  = ~A299 & A298;
  assign \new_[43478]_  = A302 & A300;
  assign \new_[43479]_  = \new_[43478]_  & \new_[43475]_ ;
  assign \new_[43480]_  = \new_[43479]_  & \new_[43472]_ ;
  assign \new_[43484]_  = ~A166 & ~A167;
  assign \new_[43485]_  = A170 & \new_[43484]_ ;
  assign \new_[43488]_  = A200 & ~A199;
  assign \new_[43491]_  = ~A235 & ~A233;
  assign \new_[43492]_  = \new_[43491]_  & \new_[43488]_ ;
  assign \new_[43493]_  = \new_[43492]_  & \new_[43485]_ ;
  assign \new_[43497]_  = A266 & A265;
  assign \new_[43498]_  = ~A236 & \new_[43497]_ ;
  assign \new_[43501]_  = ~A299 & A298;
  assign \new_[43504]_  = A301 & A300;
  assign \new_[43505]_  = \new_[43504]_  & \new_[43501]_ ;
  assign \new_[43506]_  = \new_[43505]_  & \new_[43498]_ ;
  assign \new_[43510]_  = ~A166 & ~A167;
  assign \new_[43511]_  = A170 & \new_[43510]_ ;
  assign \new_[43514]_  = A200 & ~A199;
  assign \new_[43517]_  = ~A235 & ~A233;
  assign \new_[43518]_  = \new_[43517]_  & \new_[43514]_ ;
  assign \new_[43519]_  = \new_[43518]_  & \new_[43511]_ ;
  assign \new_[43523]_  = A266 & A265;
  assign \new_[43524]_  = ~A236 & \new_[43523]_ ;
  assign \new_[43527]_  = ~A299 & A298;
  assign \new_[43530]_  = A302 & A300;
  assign \new_[43531]_  = \new_[43530]_  & \new_[43527]_ ;
  assign \new_[43532]_  = \new_[43531]_  & \new_[43524]_ ;
  assign \new_[43536]_  = ~A166 & ~A167;
  assign \new_[43537]_  = A170 & \new_[43536]_ ;
  assign \new_[43540]_  = A200 & ~A199;
  assign \new_[43543]_  = ~A235 & ~A233;
  assign \new_[43544]_  = \new_[43543]_  & \new_[43540]_ ;
  assign \new_[43545]_  = \new_[43544]_  & \new_[43537]_ ;
  assign \new_[43549]_  = ~A267 & ~A266;
  assign \new_[43550]_  = ~A236 & \new_[43549]_ ;
  assign \new_[43553]_  = ~A299 & A298;
  assign \new_[43556]_  = A301 & A300;
  assign \new_[43557]_  = \new_[43556]_  & \new_[43553]_ ;
  assign \new_[43558]_  = \new_[43557]_  & \new_[43550]_ ;
  assign \new_[43562]_  = ~A166 & ~A167;
  assign \new_[43563]_  = A170 & \new_[43562]_ ;
  assign \new_[43566]_  = A200 & ~A199;
  assign \new_[43569]_  = ~A235 & ~A233;
  assign \new_[43570]_  = \new_[43569]_  & \new_[43566]_ ;
  assign \new_[43571]_  = \new_[43570]_  & \new_[43563]_ ;
  assign \new_[43575]_  = ~A267 & ~A266;
  assign \new_[43576]_  = ~A236 & \new_[43575]_ ;
  assign \new_[43579]_  = ~A299 & A298;
  assign \new_[43582]_  = A302 & A300;
  assign \new_[43583]_  = \new_[43582]_  & \new_[43579]_ ;
  assign \new_[43584]_  = \new_[43583]_  & \new_[43576]_ ;
  assign \new_[43588]_  = ~A166 & ~A167;
  assign \new_[43589]_  = A170 & \new_[43588]_ ;
  assign \new_[43592]_  = A200 & ~A199;
  assign \new_[43595]_  = ~A235 & ~A233;
  assign \new_[43596]_  = \new_[43595]_  & \new_[43592]_ ;
  assign \new_[43597]_  = \new_[43596]_  & \new_[43589]_ ;
  assign \new_[43601]_  = ~A266 & ~A265;
  assign \new_[43602]_  = ~A236 & \new_[43601]_ ;
  assign \new_[43605]_  = ~A299 & A298;
  assign \new_[43608]_  = A301 & A300;
  assign \new_[43609]_  = \new_[43608]_  & \new_[43605]_ ;
  assign \new_[43610]_  = \new_[43609]_  & \new_[43602]_ ;
  assign \new_[43614]_  = ~A166 & ~A167;
  assign \new_[43615]_  = A170 & \new_[43614]_ ;
  assign \new_[43618]_  = A200 & ~A199;
  assign \new_[43621]_  = ~A235 & ~A233;
  assign \new_[43622]_  = \new_[43621]_  & \new_[43618]_ ;
  assign \new_[43623]_  = \new_[43622]_  & \new_[43615]_ ;
  assign \new_[43627]_  = ~A266 & ~A265;
  assign \new_[43628]_  = ~A236 & \new_[43627]_ ;
  assign \new_[43631]_  = ~A299 & A298;
  assign \new_[43634]_  = A302 & A300;
  assign \new_[43635]_  = \new_[43634]_  & \new_[43631]_ ;
  assign \new_[43636]_  = \new_[43635]_  & \new_[43628]_ ;
  assign \new_[43640]_  = ~A166 & ~A167;
  assign \new_[43641]_  = A170 & \new_[43640]_ ;
  assign \new_[43644]_  = A200 & ~A199;
  assign \new_[43647]_  = ~A234 & ~A233;
  assign \new_[43648]_  = \new_[43647]_  & \new_[43644]_ ;
  assign \new_[43649]_  = \new_[43648]_  & \new_[43641]_ ;
  assign \new_[43653]_  = ~A269 & ~A268;
  assign \new_[43654]_  = ~A266 & \new_[43653]_ ;
  assign \new_[43657]_  = ~A299 & A298;
  assign \new_[43660]_  = A301 & A300;
  assign \new_[43661]_  = \new_[43660]_  & \new_[43657]_ ;
  assign \new_[43662]_  = \new_[43661]_  & \new_[43654]_ ;
  assign \new_[43666]_  = ~A166 & ~A167;
  assign \new_[43667]_  = A170 & \new_[43666]_ ;
  assign \new_[43670]_  = A200 & ~A199;
  assign \new_[43673]_  = ~A234 & ~A233;
  assign \new_[43674]_  = \new_[43673]_  & \new_[43670]_ ;
  assign \new_[43675]_  = \new_[43674]_  & \new_[43667]_ ;
  assign \new_[43679]_  = ~A269 & ~A268;
  assign \new_[43680]_  = ~A266 & \new_[43679]_ ;
  assign \new_[43683]_  = ~A299 & A298;
  assign \new_[43686]_  = A302 & A300;
  assign \new_[43687]_  = \new_[43686]_  & \new_[43683]_ ;
  assign \new_[43688]_  = \new_[43687]_  & \new_[43680]_ ;
  assign \new_[43692]_  = ~A166 & ~A167;
  assign \new_[43693]_  = A170 & \new_[43692]_ ;
  assign \new_[43696]_  = A200 & ~A199;
  assign \new_[43699]_  = ~A233 & ~A232;
  assign \new_[43700]_  = \new_[43699]_  & \new_[43696]_ ;
  assign \new_[43701]_  = \new_[43700]_  & \new_[43693]_ ;
  assign \new_[43705]_  = ~A269 & ~A268;
  assign \new_[43706]_  = ~A266 & \new_[43705]_ ;
  assign \new_[43709]_  = ~A299 & A298;
  assign \new_[43712]_  = A301 & A300;
  assign \new_[43713]_  = \new_[43712]_  & \new_[43709]_ ;
  assign \new_[43714]_  = \new_[43713]_  & \new_[43706]_ ;
  assign \new_[43718]_  = ~A166 & ~A167;
  assign \new_[43719]_  = A170 & \new_[43718]_ ;
  assign \new_[43722]_  = A200 & ~A199;
  assign \new_[43725]_  = ~A233 & ~A232;
  assign \new_[43726]_  = \new_[43725]_  & \new_[43722]_ ;
  assign \new_[43727]_  = \new_[43726]_  & \new_[43719]_ ;
  assign \new_[43731]_  = ~A269 & ~A268;
  assign \new_[43732]_  = ~A266 & \new_[43731]_ ;
  assign \new_[43735]_  = ~A299 & A298;
  assign \new_[43738]_  = A302 & A300;
  assign \new_[43739]_  = \new_[43738]_  & \new_[43735]_ ;
  assign \new_[43740]_  = \new_[43739]_  & \new_[43732]_ ;
  assign \new_[43744]_  = ~A166 & ~A167;
  assign \new_[43745]_  = A170 & \new_[43744]_ ;
  assign \new_[43748]_  = ~A200 & A199;
  assign \new_[43751]_  = A202 & A201;
  assign \new_[43752]_  = \new_[43751]_  & \new_[43748]_ ;
  assign \new_[43753]_  = \new_[43752]_  & \new_[43745]_ ;
  assign \new_[43757]_  = A265 & A233;
  assign \new_[43758]_  = A232 & \new_[43757]_ ;
  assign \new_[43761]_  = ~A269 & ~A268;
  assign \new_[43764]_  = A299 & ~A298;
  assign \new_[43765]_  = \new_[43764]_  & \new_[43761]_ ;
  assign \new_[43766]_  = \new_[43765]_  & \new_[43758]_ ;
  assign \new_[43770]_  = ~A166 & ~A167;
  assign \new_[43771]_  = A170 & \new_[43770]_ ;
  assign \new_[43774]_  = ~A200 & A199;
  assign \new_[43777]_  = A202 & A201;
  assign \new_[43778]_  = \new_[43777]_  & \new_[43774]_ ;
  assign \new_[43779]_  = \new_[43778]_  & \new_[43771]_ ;
  assign \new_[43783]_  = ~A236 & ~A235;
  assign \new_[43784]_  = ~A233 & \new_[43783]_ ;
  assign \new_[43787]_  = A266 & A265;
  assign \new_[43790]_  = A299 & ~A298;
  assign \new_[43791]_  = \new_[43790]_  & \new_[43787]_ ;
  assign \new_[43792]_  = \new_[43791]_  & \new_[43784]_ ;
  assign \new_[43796]_  = ~A166 & ~A167;
  assign \new_[43797]_  = A170 & \new_[43796]_ ;
  assign \new_[43800]_  = ~A200 & A199;
  assign \new_[43803]_  = A202 & A201;
  assign \new_[43804]_  = \new_[43803]_  & \new_[43800]_ ;
  assign \new_[43805]_  = \new_[43804]_  & \new_[43797]_ ;
  assign \new_[43809]_  = ~A236 & ~A235;
  assign \new_[43810]_  = ~A233 & \new_[43809]_ ;
  assign \new_[43813]_  = ~A267 & ~A266;
  assign \new_[43816]_  = A299 & ~A298;
  assign \new_[43817]_  = \new_[43816]_  & \new_[43813]_ ;
  assign \new_[43818]_  = \new_[43817]_  & \new_[43810]_ ;
  assign \new_[43822]_  = ~A166 & ~A167;
  assign \new_[43823]_  = A170 & \new_[43822]_ ;
  assign \new_[43826]_  = ~A200 & A199;
  assign \new_[43829]_  = A202 & A201;
  assign \new_[43830]_  = \new_[43829]_  & \new_[43826]_ ;
  assign \new_[43831]_  = \new_[43830]_  & \new_[43823]_ ;
  assign \new_[43835]_  = ~A236 & ~A235;
  assign \new_[43836]_  = ~A233 & \new_[43835]_ ;
  assign \new_[43839]_  = ~A266 & ~A265;
  assign \new_[43842]_  = A299 & ~A298;
  assign \new_[43843]_  = \new_[43842]_  & \new_[43839]_ ;
  assign \new_[43844]_  = \new_[43843]_  & \new_[43836]_ ;
  assign \new_[43848]_  = ~A166 & ~A167;
  assign \new_[43849]_  = A170 & \new_[43848]_ ;
  assign \new_[43852]_  = ~A200 & A199;
  assign \new_[43855]_  = A202 & A201;
  assign \new_[43856]_  = \new_[43855]_  & \new_[43852]_ ;
  assign \new_[43857]_  = \new_[43856]_  & \new_[43849]_ ;
  assign \new_[43861]_  = ~A266 & ~A234;
  assign \new_[43862]_  = ~A233 & \new_[43861]_ ;
  assign \new_[43865]_  = ~A269 & ~A268;
  assign \new_[43868]_  = A299 & ~A298;
  assign \new_[43869]_  = \new_[43868]_  & \new_[43865]_ ;
  assign \new_[43870]_  = \new_[43869]_  & \new_[43862]_ ;
  assign \new_[43874]_  = ~A166 & ~A167;
  assign \new_[43875]_  = A170 & \new_[43874]_ ;
  assign \new_[43878]_  = ~A200 & A199;
  assign \new_[43881]_  = A202 & A201;
  assign \new_[43882]_  = \new_[43881]_  & \new_[43878]_ ;
  assign \new_[43883]_  = \new_[43882]_  & \new_[43875]_ ;
  assign \new_[43887]_  = A234 & ~A233;
  assign \new_[43888]_  = A232 & \new_[43887]_ ;
  assign \new_[43891]_  = A298 & A235;
  assign \new_[43894]_  = ~A302 & ~A301;
  assign \new_[43895]_  = \new_[43894]_  & \new_[43891]_ ;
  assign \new_[43896]_  = \new_[43895]_  & \new_[43888]_ ;
  assign \new_[43900]_  = ~A166 & ~A167;
  assign \new_[43901]_  = A170 & \new_[43900]_ ;
  assign \new_[43904]_  = ~A200 & A199;
  assign \new_[43907]_  = A202 & A201;
  assign \new_[43908]_  = \new_[43907]_  & \new_[43904]_ ;
  assign \new_[43909]_  = \new_[43908]_  & \new_[43901]_ ;
  assign \new_[43913]_  = A234 & ~A233;
  assign \new_[43914]_  = A232 & \new_[43913]_ ;
  assign \new_[43917]_  = A298 & A236;
  assign \new_[43920]_  = ~A302 & ~A301;
  assign \new_[43921]_  = \new_[43920]_  & \new_[43917]_ ;
  assign \new_[43922]_  = \new_[43921]_  & \new_[43914]_ ;
  assign \new_[43926]_  = ~A166 & ~A167;
  assign \new_[43927]_  = A170 & \new_[43926]_ ;
  assign \new_[43930]_  = ~A200 & A199;
  assign \new_[43933]_  = A202 & A201;
  assign \new_[43934]_  = \new_[43933]_  & \new_[43930]_ ;
  assign \new_[43935]_  = \new_[43934]_  & \new_[43927]_ ;
  assign \new_[43939]_  = ~A266 & ~A233;
  assign \new_[43940]_  = ~A232 & \new_[43939]_ ;
  assign \new_[43943]_  = ~A269 & ~A268;
  assign \new_[43946]_  = A299 & ~A298;
  assign \new_[43947]_  = \new_[43946]_  & \new_[43943]_ ;
  assign \new_[43948]_  = \new_[43947]_  & \new_[43940]_ ;
  assign \new_[43952]_  = ~A166 & ~A167;
  assign \new_[43953]_  = A170 & \new_[43952]_ ;
  assign \new_[43956]_  = ~A200 & A199;
  assign \new_[43959]_  = A203 & A201;
  assign \new_[43960]_  = \new_[43959]_  & \new_[43956]_ ;
  assign \new_[43961]_  = \new_[43960]_  & \new_[43953]_ ;
  assign \new_[43965]_  = A265 & A233;
  assign \new_[43966]_  = A232 & \new_[43965]_ ;
  assign \new_[43969]_  = ~A269 & ~A268;
  assign \new_[43972]_  = A299 & ~A298;
  assign \new_[43973]_  = \new_[43972]_  & \new_[43969]_ ;
  assign \new_[43974]_  = \new_[43973]_  & \new_[43966]_ ;
  assign \new_[43978]_  = ~A166 & ~A167;
  assign \new_[43979]_  = A170 & \new_[43978]_ ;
  assign \new_[43982]_  = ~A200 & A199;
  assign \new_[43985]_  = A203 & A201;
  assign \new_[43986]_  = \new_[43985]_  & \new_[43982]_ ;
  assign \new_[43987]_  = \new_[43986]_  & \new_[43979]_ ;
  assign \new_[43991]_  = ~A236 & ~A235;
  assign \new_[43992]_  = ~A233 & \new_[43991]_ ;
  assign \new_[43995]_  = A266 & A265;
  assign \new_[43998]_  = A299 & ~A298;
  assign \new_[43999]_  = \new_[43998]_  & \new_[43995]_ ;
  assign \new_[44000]_  = \new_[43999]_  & \new_[43992]_ ;
  assign \new_[44004]_  = ~A166 & ~A167;
  assign \new_[44005]_  = A170 & \new_[44004]_ ;
  assign \new_[44008]_  = ~A200 & A199;
  assign \new_[44011]_  = A203 & A201;
  assign \new_[44012]_  = \new_[44011]_  & \new_[44008]_ ;
  assign \new_[44013]_  = \new_[44012]_  & \new_[44005]_ ;
  assign \new_[44017]_  = ~A236 & ~A235;
  assign \new_[44018]_  = ~A233 & \new_[44017]_ ;
  assign \new_[44021]_  = ~A267 & ~A266;
  assign \new_[44024]_  = A299 & ~A298;
  assign \new_[44025]_  = \new_[44024]_  & \new_[44021]_ ;
  assign \new_[44026]_  = \new_[44025]_  & \new_[44018]_ ;
  assign \new_[44030]_  = ~A166 & ~A167;
  assign \new_[44031]_  = A170 & \new_[44030]_ ;
  assign \new_[44034]_  = ~A200 & A199;
  assign \new_[44037]_  = A203 & A201;
  assign \new_[44038]_  = \new_[44037]_  & \new_[44034]_ ;
  assign \new_[44039]_  = \new_[44038]_  & \new_[44031]_ ;
  assign \new_[44043]_  = ~A236 & ~A235;
  assign \new_[44044]_  = ~A233 & \new_[44043]_ ;
  assign \new_[44047]_  = ~A266 & ~A265;
  assign \new_[44050]_  = A299 & ~A298;
  assign \new_[44051]_  = \new_[44050]_  & \new_[44047]_ ;
  assign \new_[44052]_  = \new_[44051]_  & \new_[44044]_ ;
  assign \new_[44056]_  = ~A166 & ~A167;
  assign \new_[44057]_  = A170 & \new_[44056]_ ;
  assign \new_[44060]_  = ~A200 & A199;
  assign \new_[44063]_  = A203 & A201;
  assign \new_[44064]_  = \new_[44063]_  & \new_[44060]_ ;
  assign \new_[44065]_  = \new_[44064]_  & \new_[44057]_ ;
  assign \new_[44069]_  = ~A266 & ~A234;
  assign \new_[44070]_  = ~A233 & \new_[44069]_ ;
  assign \new_[44073]_  = ~A269 & ~A268;
  assign \new_[44076]_  = A299 & ~A298;
  assign \new_[44077]_  = \new_[44076]_  & \new_[44073]_ ;
  assign \new_[44078]_  = \new_[44077]_  & \new_[44070]_ ;
  assign \new_[44082]_  = ~A166 & ~A167;
  assign \new_[44083]_  = A170 & \new_[44082]_ ;
  assign \new_[44086]_  = ~A200 & A199;
  assign \new_[44089]_  = A203 & A201;
  assign \new_[44090]_  = \new_[44089]_  & \new_[44086]_ ;
  assign \new_[44091]_  = \new_[44090]_  & \new_[44083]_ ;
  assign \new_[44095]_  = A234 & ~A233;
  assign \new_[44096]_  = A232 & \new_[44095]_ ;
  assign \new_[44099]_  = A298 & A235;
  assign \new_[44102]_  = ~A302 & ~A301;
  assign \new_[44103]_  = \new_[44102]_  & \new_[44099]_ ;
  assign \new_[44104]_  = \new_[44103]_  & \new_[44096]_ ;
  assign \new_[44108]_  = ~A166 & ~A167;
  assign \new_[44109]_  = A170 & \new_[44108]_ ;
  assign \new_[44112]_  = ~A200 & A199;
  assign \new_[44115]_  = A203 & A201;
  assign \new_[44116]_  = \new_[44115]_  & \new_[44112]_ ;
  assign \new_[44117]_  = \new_[44116]_  & \new_[44109]_ ;
  assign \new_[44121]_  = A234 & ~A233;
  assign \new_[44122]_  = A232 & \new_[44121]_ ;
  assign \new_[44125]_  = A298 & A236;
  assign \new_[44128]_  = ~A302 & ~A301;
  assign \new_[44129]_  = \new_[44128]_  & \new_[44125]_ ;
  assign \new_[44130]_  = \new_[44129]_  & \new_[44122]_ ;
  assign \new_[44134]_  = ~A166 & ~A167;
  assign \new_[44135]_  = A170 & \new_[44134]_ ;
  assign \new_[44138]_  = ~A200 & A199;
  assign \new_[44141]_  = A203 & A201;
  assign \new_[44142]_  = \new_[44141]_  & \new_[44138]_ ;
  assign \new_[44143]_  = \new_[44142]_  & \new_[44135]_ ;
  assign \new_[44147]_  = ~A266 & ~A233;
  assign \new_[44148]_  = ~A232 & \new_[44147]_ ;
  assign \new_[44151]_  = ~A269 & ~A268;
  assign \new_[44154]_  = A299 & ~A298;
  assign \new_[44155]_  = \new_[44154]_  & \new_[44151]_ ;
  assign \new_[44156]_  = \new_[44155]_  & \new_[44148]_ ;
  assign \new_[44160]_  = A167 & ~A168;
  assign \new_[44161]_  = A170 & \new_[44160]_ ;
  assign \new_[44164]_  = ~A199 & A166;
  assign \new_[44167]_  = A232 & A200;
  assign \new_[44168]_  = \new_[44167]_  & \new_[44164]_ ;
  assign \new_[44169]_  = \new_[44168]_  & \new_[44161]_ ;
  assign \new_[44173]_  = ~A267 & A265;
  assign \new_[44174]_  = A233 & \new_[44173]_ ;
  assign \new_[44177]_  = ~A299 & A298;
  assign \new_[44180]_  = A301 & A300;
  assign \new_[44181]_  = \new_[44180]_  & \new_[44177]_ ;
  assign \new_[44182]_  = \new_[44181]_  & \new_[44174]_ ;
  assign \new_[44186]_  = A167 & ~A168;
  assign \new_[44187]_  = A170 & \new_[44186]_ ;
  assign \new_[44190]_  = ~A199 & A166;
  assign \new_[44193]_  = A232 & A200;
  assign \new_[44194]_  = \new_[44193]_  & \new_[44190]_ ;
  assign \new_[44195]_  = \new_[44194]_  & \new_[44187]_ ;
  assign \new_[44199]_  = ~A267 & A265;
  assign \new_[44200]_  = A233 & \new_[44199]_ ;
  assign \new_[44203]_  = ~A299 & A298;
  assign \new_[44206]_  = A302 & A300;
  assign \new_[44207]_  = \new_[44206]_  & \new_[44203]_ ;
  assign \new_[44208]_  = \new_[44207]_  & \new_[44200]_ ;
  assign \new_[44212]_  = A167 & ~A168;
  assign \new_[44213]_  = A170 & \new_[44212]_ ;
  assign \new_[44216]_  = ~A199 & A166;
  assign \new_[44219]_  = A232 & A200;
  assign \new_[44220]_  = \new_[44219]_  & \new_[44216]_ ;
  assign \new_[44221]_  = \new_[44220]_  & \new_[44213]_ ;
  assign \new_[44225]_  = A266 & A265;
  assign \new_[44226]_  = A233 & \new_[44225]_ ;
  assign \new_[44229]_  = ~A299 & A298;
  assign \new_[44232]_  = A301 & A300;
  assign \new_[44233]_  = \new_[44232]_  & \new_[44229]_ ;
  assign \new_[44234]_  = \new_[44233]_  & \new_[44226]_ ;
  assign \new_[44238]_  = A167 & ~A168;
  assign \new_[44239]_  = A170 & \new_[44238]_ ;
  assign \new_[44242]_  = ~A199 & A166;
  assign \new_[44245]_  = A232 & A200;
  assign \new_[44246]_  = \new_[44245]_  & \new_[44242]_ ;
  assign \new_[44247]_  = \new_[44246]_  & \new_[44239]_ ;
  assign \new_[44251]_  = A266 & A265;
  assign \new_[44252]_  = A233 & \new_[44251]_ ;
  assign \new_[44255]_  = ~A299 & A298;
  assign \new_[44258]_  = A302 & A300;
  assign \new_[44259]_  = \new_[44258]_  & \new_[44255]_ ;
  assign \new_[44260]_  = \new_[44259]_  & \new_[44252]_ ;
  assign \new_[44264]_  = A167 & ~A168;
  assign \new_[44265]_  = A170 & \new_[44264]_ ;
  assign \new_[44268]_  = ~A199 & A166;
  assign \new_[44271]_  = A232 & A200;
  assign \new_[44272]_  = \new_[44271]_  & \new_[44268]_ ;
  assign \new_[44273]_  = \new_[44272]_  & \new_[44265]_ ;
  assign \new_[44277]_  = ~A266 & ~A265;
  assign \new_[44278]_  = A233 & \new_[44277]_ ;
  assign \new_[44281]_  = ~A299 & A298;
  assign \new_[44284]_  = A301 & A300;
  assign \new_[44285]_  = \new_[44284]_  & \new_[44281]_ ;
  assign \new_[44286]_  = \new_[44285]_  & \new_[44278]_ ;
  assign \new_[44290]_  = A167 & ~A168;
  assign \new_[44291]_  = A170 & \new_[44290]_ ;
  assign \new_[44294]_  = ~A199 & A166;
  assign \new_[44297]_  = A232 & A200;
  assign \new_[44298]_  = \new_[44297]_  & \new_[44294]_ ;
  assign \new_[44299]_  = \new_[44298]_  & \new_[44291]_ ;
  assign \new_[44303]_  = ~A266 & ~A265;
  assign \new_[44304]_  = A233 & \new_[44303]_ ;
  assign \new_[44307]_  = ~A299 & A298;
  assign \new_[44310]_  = A302 & A300;
  assign \new_[44311]_  = \new_[44310]_  & \new_[44307]_ ;
  assign \new_[44312]_  = \new_[44311]_  & \new_[44304]_ ;
  assign \new_[44316]_  = A167 & ~A168;
  assign \new_[44317]_  = A170 & \new_[44316]_ ;
  assign \new_[44320]_  = ~A199 & A166;
  assign \new_[44323]_  = ~A233 & A200;
  assign \new_[44324]_  = \new_[44323]_  & \new_[44320]_ ;
  assign \new_[44325]_  = \new_[44324]_  & \new_[44317]_ ;
  assign \new_[44329]_  = ~A266 & ~A236;
  assign \new_[44330]_  = ~A235 & \new_[44329]_ ;
  assign \new_[44333]_  = ~A269 & ~A268;
  assign \new_[44336]_  = A299 & ~A298;
  assign \new_[44337]_  = \new_[44336]_  & \new_[44333]_ ;
  assign \new_[44338]_  = \new_[44337]_  & \new_[44330]_ ;
  assign \new_[44342]_  = A167 & ~A168;
  assign \new_[44343]_  = A170 & \new_[44342]_ ;
  assign \new_[44346]_  = ~A199 & A166;
  assign \new_[44349]_  = ~A233 & A200;
  assign \new_[44350]_  = \new_[44349]_  & \new_[44346]_ ;
  assign \new_[44351]_  = \new_[44350]_  & \new_[44343]_ ;
  assign \new_[44355]_  = A266 & A265;
  assign \new_[44356]_  = ~A234 & \new_[44355]_ ;
  assign \new_[44359]_  = ~A299 & A298;
  assign \new_[44362]_  = A301 & A300;
  assign \new_[44363]_  = \new_[44362]_  & \new_[44359]_ ;
  assign \new_[44364]_  = \new_[44363]_  & \new_[44356]_ ;
  assign \new_[44368]_  = A167 & ~A168;
  assign \new_[44369]_  = A170 & \new_[44368]_ ;
  assign \new_[44372]_  = ~A199 & A166;
  assign \new_[44375]_  = ~A233 & A200;
  assign \new_[44376]_  = \new_[44375]_  & \new_[44372]_ ;
  assign \new_[44377]_  = \new_[44376]_  & \new_[44369]_ ;
  assign \new_[44381]_  = A266 & A265;
  assign \new_[44382]_  = ~A234 & \new_[44381]_ ;
  assign \new_[44385]_  = ~A299 & A298;
  assign \new_[44388]_  = A302 & A300;
  assign \new_[44389]_  = \new_[44388]_  & \new_[44385]_ ;
  assign \new_[44390]_  = \new_[44389]_  & \new_[44382]_ ;
  assign \new_[44394]_  = A167 & ~A168;
  assign \new_[44395]_  = A170 & \new_[44394]_ ;
  assign \new_[44398]_  = ~A199 & A166;
  assign \new_[44401]_  = ~A233 & A200;
  assign \new_[44402]_  = \new_[44401]_  & \new_[44398]_ ;
  assign \new_[44403]_  = \new_[44402]_  & \new_[44395]_ ;
  assign \new_[44407]_  = ~A267 & ~A266;
  assign \new_[44408]_  = ~A234 & \new_[44407]_ ;
  assign \new_[44411]_  = ~A299 & A298;
  assign \new_[44414]_  = A301 & A300;
  assign \new_[44415]_  = \new_[44414]_  & \new_[44411]_ ;
  assign \new_[44416]_  = \new_[44415]_  & \new_[44408]_ ;
  assign \new_[44420]_  = A167 & ~A168;
  assign \new_[44421]_  = A170 & \new_[44420]_ ;
  assign \new_[44424]_  = ~A199 & A166;
  assign \new_[44427]_  = ~A233 & A200;
  assign \new_[44428]_  = \new_[44427]_  & \new_[44424]_ ;
  assign \new_[44429]_  = \new_[44428]_  & \new_[44421]_ ;
  assign \new_[44433]_  = ~A267 & ~A266;
  assign \new_[44434]_  = ~A234 & \new_[44433]_ ;
  assign \new_[44437]_  = ~A299 & A298;
  assign \new_[44440]_  = A302 & A300;
  assign \new_[44441]_  = \new_[44440]_  & \new_[44437]_ ;
  assign \new_[44442]_  = \new_[44441]_  & \new_[44434]_ ;
  assign \new_[44446]_  = A167 & ~A168;
  assign \new_[44447]_  = A170 & \new_[44446]_ ;
  assign \new_[44450]_  = ~A199 & A166;
  assign \new_[44453]_  = ~A233 & A200;
  assign \new_[44454]_  = \new_[44453]_  & \new_[44450]_ ;
  assign \new_[44455]_  = \new_[44454]_  & \new_[44447]_ ;
  assign \new_[44459]_  = ~A266 & ~A265;
  assign \new_[44460]_  = ~A234 & \new_[44459]_ ;
  assign \new_[44463]_  = ~A299 & A298;
  assign \new_[44466]_  = A301 & A300;
  assign \new_[44467]_  = \new_[44466]_  & \new_[44463]_ ;
  assign \new_[44468]_  = \new_[44467]_  & \new_[44460]_ ;
  assign \new_[44472]_  = A167 & ~A168;
  assign \new_[44473]_  = A170 & \new_[44472]_ ;
  assign \new_[44476]_  = ~A199 & A166;
  assign \new_[44479]_  = ~A233 & A200;
  assign \new_[44480]_  = \new_[44479]_  & \new_[44476]_ ;
  assign \new_[44481]_  = \new_[44480]_  & \new_[44473]_ ;
  assign \new_[44485]_  = ~A266 & ~A265;
  assign \new_[44486]_  = ~A234 & \new_[44485]_ ;
  assign \new_[44489]_  = ~A299 & A298;
  assign \new_[44492]_  = A302 & A300;
  assign \new_[44493]_  = \new_[44492]_  & \new_[44489]_ ;
  assign \new_[44494]_  = \new_[44493]_  & \new_[44486]_ ;
  assign \new_[44498]_  = A167 & ~A168;
  assign \new_[44499]_  = A170 & \new_[44498]_ ;
  assign \new_[44502]_  = ~A199 & A166;
  assign \new_[44505]_  = A232 & A200;
  assign \new_[44506]_  = \new_[44505]_  & \new_[44502]_ ;
  assign \new_[44507]_  = \new_[44506]_  & \new_[44499]_ ;
  assign \new_[44511]_  = A235 & A234;
  assign \new_[44512]_  = ~A233 & \new_[44511]_ ;
  assign \new_[44515]_  = ~A266 & A265;
  assign \new_[44518]_  = A268 & A267;
  assign \new_[44519]_  = \new_[44518]_  & \new_[44515]_ ;
  assign \new_[44520]_  = \new_[44519]_  & \new_[44512]_ ;
  assign \new_[44524]_  = A167 & ~A168;
  assign \new_[44525]_  = A170 & \new_[44524]_ ;
  assign \new_[44528]_  = ~A199 & A166;
  assign \new_[44531]_  = A232 & A200;
  assign \new_[44532]_  = \new_[44531]_  & \new_[44528]_ ;
  assign \new_[44533]_  = \new_[44532]_  & \new_[44525]_ ;
  assign \new_[44537]_  = A235 & A234;
  assign \new_[44538]_  = ~A233 & \new_[44537]_ ;
  assign \new_[44541]_  = ~A266 & A265;
  assign \new_[44544]_  = A269 & A267;
  assign \new_[44545]_  = \new_[44544]_  & \new_[44541]_ ;
  assign \new_[44546]_  = \new_[44545]_  & \new_[44538]_ ;
  assign \new_[44550]_  = A167 & ~A168;
  assign \new_[44551]_  = A170 & \new_[44550]_ ;
  assign \new_[44554]_  = ~A199 & A166;
  assign \new_[44557]_  = A232 & A200;
  assign \new_[44558]_  = \new_[44557]_  & \new_[44554]_ ;
  assign \new_[44559]_  = \new_[44558]_  & \new_[44551]_ ;
  assign \new_[44563]_  = A236 & A234;
  assign \new_[44564]_  = ~A233 & \new_[44563]_ ;
  assign \new_[44567]_  = ~A266 & A265;
  assign \new_[44570]_  = A268 & A267;
  assign \new_[44571]_  = \new_[44570]_  & \new_[44567]_ ;
  assign \new_[44572]_  = \new_[44571]_  & \new_[44564]_ ;
  assign \new_[44576]_  = A167 & ~A168;
  assign \new_[44577]_  = A170 & \new_[44576]_ ;
  assign \new_[44580]_  = ~A199 & A166;
  assign \new_[44583]_  = A232 & A200;
  assign \new_[44584]_  = \new_[44583]_  & \new_[44580]_ ;
  assign \new_[44585]_  = \new_[44584]_  & \new_[44577]_ ;
  assign \new_[44589]_  = A236 & A234;
  assign \new_[44590]_  = ~A233 & \new_[44589]_ ;
  assign \new_[44593]_  = ~A266 & A265;
  assign \new_[44596]_  = A269 & A267;
  assign \new_[44597]_  = \new_[44596]_  & \new_[44593]_ ;
  assign \new_[44598]_  = \new_[44597]_  & \new_[44590]_ ;
  assign \new_[44602]_  = A167 & ~A168;
  assign \new_[44603]_  = A170 & \new_[44602]_ ;
  assign \new_[44606]_  = ~A199 & A166;
  assign \new_[44609]_  = ~A232 & A200;
  assign \new_[44610]_  = \new_[44609]_  & \new_[44606]_ ;
  assign \new_[44611]_  = \new_[44610]_  & \new_[44603]_ ;
  assign \new_[44615]_  = A266 & A265;
  assign \new_[44616]_  = ~A233 & \new_[44615]_ ;
  assign \new_[44619]_  = ~A299 & A298;
  assign \new_[44622]_  = A301 & A300;
  assign \new_[44623]_  = \new_[44622]_  & \new_[44619]_ ;
  assign \new_[44624]_  = \new_[44623]_  & \new_[44616]_ ;
  assign \new_[44628]_  = A167 & ~A168;
  assign \new_[44629]_  = A170 & \new_[44628]_ ;
  assign \new_[44632]_  = ~A199 & A166;
  assign \new_[44635]_  = ~A232 & A200;
  assign \new_[44636]_  = \new_[44635]_  & \new_[44632]_ ;
  assign \new_[44637]_  = \new_[44636]_  & \new_[44629]_ ;
  assign \new_[44641]_  = A266 & A265;
  assign \new_[44642]_  = ~A233 & \new_[44641]_ ;
  assign \new_[44645]_  = ~A299 & A298;
  assign \new_[44648]_  = A302 & A300;
  assign \new_[44649]_  = \new_[44648]_  & \new_[44645]_ ;
  assign \new_[44650]_  = \new_[44649]_  & \new_[44642]_ ;
  assign \new_[44654]_  = A167 & ~A168;
  assign \new_[44655]_  = A170 & \new_[44654]_ ;
  assign \new_[44658]_  = ~A199 & A166;
  assign \new_[44661]_  = ~A232 & A200;
  assign \new_[44662]_  = \new_[44661]_  & \new_[44658]_ ;
  assign \new_[44663]_  = \new_[44662]_  & \new_[44655]_ ;
  assign \new_[44667]_  = ~A267 & ~A266;
  assign \new_[44668]_  = ~A233 & \new_[44667]_ ;
  assign \new_[44671]_  = ~A299 & A298;
  assign \new_[44674]_  = A301 & A300;
  assign \new_[44675]_  = \new_[44674]_  & \new_[44671]_ ;
  assign \new_[44676]_  = \new_[44675]_  & \new_[44668]_ ;
  assign \new_[44680]_  = A167 & ~A168;
  assign \new_[44681]_  = A170 & \new_[44680]_ ;
  assign \new_[44684]_  = ~A199 & A166;
  assign \new_[44687]_  = ~A232 & A200;
  assign \new_[44688]_  = \new_[44687]_  & \new_[44684]_ ;
  assign \new_[44689]_  = \new_[44688]_  & \new_[44681]_ ;
  assign \new_[44693]_  = ~A267 & ~A266;
  assign \new_[44694]_  = ~A233 & \new_[44693]_ ;
  assign \new_[44697]_  = ~A299 & A298;
  assign \new_[44700]_  = A302 & A300;
  assign \new_[44701]_  = \new_[44700]_  & \new_[44697]_ ;
  assign \new_[44702]_  = \new_[44701]_  & \new_[44694]_ ;
  assign \new_[44706]_  = A167 & ~A168;
  assign \new_[44707]_  = A170 & \new_[44706]_ ;
  assign \new_[44710]_  = ~A199 & A166;
  assign \new_[44713]_  = ~A232 & A200;
  assign \new_[44714]_  = \new_[44713]_  & \new_[44710]_ ;
  assign \new_[44715]_  = \new_[44714]_  & \new_[44707]_ ;
  assign \new_[44719]_  = ~A266 & ~A265;
  assign \new_[44720]_  = ~A233 & \new_[44719]_ ;
  assign \new_[44723]_  = ~A299 & A298;
  assign \new_[44726]_  = A301 & A300;
  assign \new_[44727]_  = \new_[44726]_  & \new_[44723]_ ;
  assign \new_[44728]_  = \new_[44727]_  & \new_[44720]_ ;
  assign \new_[44732]_  = A167 & ~A168;
  assign \new_[44733]_  = A170 & \new_[44732]_ ;
  assign \new_[44736]_  = ~A199 & A166;
  assign \new_[44739]_  = ~A232 & A200;
  assign \new_[44740]_  = \new_[44739]_  & \new_[44736]_ ;
  assign \new_[44741]_  = \new_[44740]_  & \new_[44733]_ ;
  assign \new_[44745]_  = ~A266 & ~A265;
  assign \new_[44746]_  = ~A233 & \new_[44745]_ ;
  assign \new_[44749]_  = ~A299 & A298;
  assign \new_[44752]_  = A302 & A300;
  assign \new_[44753]_  = \new_[44752]_  & \new_[44749]_ ;
  assign \new_[44754]_  = \new_[44753]_  & \new_[44746]_ ;
  assign \new_[44758]_  = A167 & ~A168;
  assign \new_[44759]_  = ~A170 & \new_[44758]_ ;
  assign \new_[44762]_  = ~A199 & ~A166;
  assign \new_[44765]_  = A232 & A200;
  assign \new_[44766]_  = \new_[44765]_  & \new_[44762]_ ;
  assign \new_[44767]_  = \new_[44766]_  & \new_[44759]_ ;
  assign \new_[44771]_  = ~A267 & A265;
  assign \new_[44772]_  = A233 & \new_[44771]_ ;
  assign \new_[44775]_  = ~A299 & A298;
  assign \new_[44778]_  = A301 & A300;
  assign \new_[44779]_  = \new_[44778]_  & \new_[44775]_ ;
  assign \new_[44780]_  = \new_[44779]_  & \new_[44772]_ ;
  assign \new_[44784]_  = A167 & ~A168;
  assign \new_[44785]_  = ~A170 & \new_[44784]_ ;
  assign \new_[44788]_  = ~A199 & ~A166;
  assign \new_[44791]_  = A232 & A200;
  assign \new_[44792]_  = \new_[44791]_  & \new_[44788]_ ;
  assign \new_[44793]_  = \new_[44792]_  & \new_[44785]_ ;
  assign \new_[44797]_  = ~A267 & A265;
  assign \new_[44798]_  = A233 & \new_[44797]_ ;
  assign \new_[44801]_  = ~A299 & A298;
  assign \new_[44804]_  = A302 & A300;
  assign \new_[44805]_  = \new_[44804]_  & \new_[44801]_ ;
  assign \new_[44806]_  = \new_[44805]_  & \new_[44798]_ ;
  assign \new_[44810]_  = A167 & ~A168;
  assign \new_[44811]_  = ~A170 & \new_[44810]_ ;
  assign \new_[44814]_  = ~A199 & ~A166;
  assign \new_[44817]_  = A232 & A200;
  assign \new_[44818]_  = \new_[44817]_  & \new_[44814]_ ;
  assign \new_[44819]_  = \new_[44818]_  & \new_[44811]_ ;
  assign \new_[44823]_  = A266 & A265;
  assign \new_[44824]_  = A233 & \new_[44823]_ ;
  assign \new_[44827]_  = ~A299 & A298;
  assign \new_[44830]_  = A301 & A300;
  assign \new_[44831]_  = \new_[44830]_  & \new_[44827]_ ;
  assign \new_[44832]_  = \new_[44831]_  & \new_[44824]_ ;
  assign \new_[44836]_  = A167 & ~A168;
  assign \new_[44837]_  = ~A170 & \new_[44836]_ ;
  assign \new_[44840]_  = ~A199 & ~A166;
  assign \new_[44843]_  = A232 & A200;
  assign \new_[44844]_  = \new_[44843]_  & \new_[44840]_ ;
  assign \new_[44845]_  = \new_[44844]_  & \new_[44837]_ ;
  assign \new_[44849]_  = A266 & A265;
  assign \new_[44850]_  = A233 & \new_[44849]_ ;
  assign \new_[44853]_  = ~A299 & A298;
  assign \new_[44856]_  = A302 & A300;
  assign \new_[44857]_  = \new_[44856]_  & \new_[44853]_ ;
  assign \new_[44858]_  = \new_[44857]_  & \new_[44850]_ ;
  assign \new_[44862]_  = A167 & ~A168;
  assign \new_[44863]_  = ~A170 & \new_[44862]_ ;
  assign \new_[44866]_  = ~A199 & ~A166;
  assign \new_[44869]_  = A232 & A200;
  assign \new_[44870]_  = \new_[44869]_  & \new_[44866]_ ;
  assign \new_[44871]_  = \new_[44870]_  & \new_[44863]_ ;
  assign \new_[44875]_  = ~A266 & ~A265;
  assign \new_[44876]_  = A233 & \new_[44875]_ ;
  assign \new_[44879]_  = ~A299 & A298;
  assign \new_[44882]_  = A301 & A300;
  assign \new_[44883]_  = \new_[44882]_  & \new_[44879]_ ;
  assign \new_[44884]_  = \new_[44883]_  & \new_[44876]_ ;
  assign \new_[44888]_  = A167 & ~A168;
  assign \new_[44889]_  = ~A170 & \new_[44888]_ ;
  assign \new_[44892]_  = ~A199 & ~A166;
  assign \new_[44895]_  = A232 & A200;
  assign \new_[44896]_  = \new_[44895]_  & \new_[44892]_ ;
  assign \new_[44897]_  = \new_[44896]_  & \new_[44889]_ ;
  assign \new_[44901]_  = ~A266 & ~A265;
  assign \new_[44902]_  = A233 & \new_[44901]_ ;
  assign \new_[44905]_  = ~A299 & A298;
  assign \new_[44908]_  = A302 & A300;
  assign \new_[44909]_  = \new_[44908]_  & \new_[44905]_ ;
  assign \new_[44910]_  = \new_[44909]_  & \new_[44902]_ ;
  assign \new_[44914]_  = A167 & ~A168;
  assign \new_[44915]_  = ~A170 & \new_[44914]_ ;
  assign \new_[44918]_  = ~A199 & ~A166;
  assign \new_[44921]_  = ~A233 & A200;
  assign \new_[44922]_  = \new_[44921]_  & \new_[44918]_ ;
  assign \new_[44923]_  = \new_[44922]_  & \new_[44915]_ ;
  assign \new_[44927]_  = ~A266 & ~A236;
  assign \new_[44928]_  = ~A235 & \new_[44927]_ ;
  assign \new_[44931]_  = ~A269 & ~A268;
  assign \new_[44934]_  = A299 & ~A298;
  assign \new_[44935]_  = \new_[44934]_  & \new_[44931]_ ;
  assign \new_[44936]_  = \new_[44935]_  & \new_[44928]_ ;
  assign \new_[44940]_  = A167 & ~A168;
  assign \new_[44941]_  = ~A170 & \new_[44940]_ ;
  assign \new_[44944]_  = ~A199 & ~A166;
  assign \new_[44947]_  = ~A233 & A200;
  assign \new_[44948]_  = \new_[44947]_  & \new_[44944]_ ;
  assign \new_[44949]_  = \new_[44948]_  & \new_[44941]_ ;
  assign \new_[44953]_  = A266 & A265;
  assign \new_[44954]_  = ~A234 & \new_[44953]_ ;
  assign \new_[44957]_  = ~A299 & A298;
  assign \new_[44960]_  = A301 & A300;
  assign \new_[44961]_  = \new_[44960]_  & \new_[44957]_ ;
  assign \new_[44962]_  = \new_[44961]_  & \new_[44954]_ ;
  assign \new_[44966]_  = A167 & ~A168;
  assign \new_[44967]_  = ~A170 & \new_[44966]_ ;
  assign \new_[44970]_  = ~A199 & ~A166;
  assign \new_[44973]_  = ~A233 & A200;
  assign \new_[44974]_  = \new_[44973]_  & \new_[44970]_ ;
  assign \new_[44975]_  = \new_[44974]_  & \new_[44967]_ ;
  assign \new_[44979]_  = A266 & A265;
  assign \new_[44980]_  = ~A234 & \new_[44979]_ ;
  assign \new_[44983]_  = ~A299 & A298;
  assign \new_[44986]_  = A302 & A300;
  assign \new_[44987]_  = \new_[44986]_  & \new_[44983]_ ;
  assign \new_[44988]_  = \new_[44987]_  & \new_[44980]_ ;
  assign \new_[44992]_  = A167 & ~A168;
  assign \new_[44993]_  = ~A170 & \new_[44992]_ ;
  assign \new_[44996]_  = ~A199 & ~A166;
  assign \new_[44999]_  = ~A233 & A200;
  assign \new_[45000]_  = \new_[44999]_  & \new_[44996]_ ;
  assign \new_[45001]_  = \new_[45000]_  & \new_[44993]_ ;
  assign \new_[45005]_  = ~A267 & ~A266;
  assign \new_[45006]_  = ~A234 & \new_[45005]_ ;
  assign \new_[45009]_  = ~A299 & A298;
  assign \new_[45012]_  = A301 & A300;
  assign \new_[45013]_  = \new_[45012]_  & \new_[45009]_ ;
  assign \new_[45014]_  = \new_[45013]_  & \new_[45006]_ ;
  assign \new_[45018]_  = A167 & ~A168;
  assign \new_[45019]_  = ~A170 & \new_[45018]_ ;
  assign \new_[45022]_  = ~A199 & ~A166;
  assign \new_[45025]_  = ~A233 & A200;
  assign \new_[45026]_  = \new_[45025]_  & \new_[45022]_ ;
  assign \new_[45027]_  = \new_[45026]_  & \new_[45019]_ ;
  assign \new_[45031]_  = ~A267 & ~A266;
  assign \new_[45032]_  = ~A234 & \new_[45031]_ ;
  assign \new_[45035]_  = ~A299 & A298;
  assign \new_[45038]_  = A302 & A300;
  assign \new_[45039]_  = \new_[45038]_  & \new_[45035]_ ;
  assign \new_[45040]_  = \new_[45039]_  & \new_[45032]_ ;
  assign \new_[45044]_  = A167 & ~A168;
  assign \new_[45045]_  = ~A170 & \new_[45044]_ ;
  assign \new_[45048]_  = ~A199 & ~A166;
  assign \new_[45051]_  = ~A233 & A200;
  assign \new_[45052]_  = \new_[45051]_  & \new_[45048]_ ;
  assign \new_[45053]_  = \new_[45052]_  & \new_[45045]_ ;
  assign \new_[45057]_  = ~A266 & ~A265;
  assign \new_[45058]_  = ~A234 & \new_[45057]_ ;
  assign \new_[45061]_  = ~A299 & A298;
  assign \new_[45064]_  = A301 & A300;
  assign \new_[45065]_  = \new_[45064]_  & \new_[45061]_ ;
  assign \new_[45066]_  = \new_[45065]_  & \new_[45058]_ ;
  assign \new_[45070]_  = A167 & ~A168;
  assign \new_[45071]_  = ~A170 & \new_[45070]_ ;
  assign \new_[45074]_  = ~A199 & ~A166;
  assign \new_[45077]_  = ~A233 & A200;
  assign \new_[45078]_  = \new_[45077]_  & \new_[45074]_ ;
  assign \new_[45079]_  = \new_[45078]_  & \new_[45071]_ ;
  assign \new_[45083]_  = ~A266 & ~A265;
  assign \new_[45084]_  = ~A234 & \new_[45083]_ ;
  assign \new_[45087]_  = ~A299 & A298;
  assign \new_[45090]_  = A302 & A300;
  assign \new_[45091]_  = \new_[45090]_  & \new_[45087]_ ;
  assign \new_[45092]_  = \new_[45091]_  & \new_[45084]_ ;
  assign \new_[45096]_  = A167 & ~A168;
  assign \new_[45097]_  = ~A170 & \new_[45096]_ ;
  assign \new_[45100]_  = ~A199 & ~A166;
  assign \new_[45103]_  = A232 & A200;
  assign \new_[45104]_  = \new_[45103]_  & \new_[45100]_ ;
  assign \new_[45105]_  = \new_[45104]_  & \new_[45097]_ ;
  assign \new_[45109]_  = A235 & A234;
  assign \new_[45110]_  = ~A233 & \new_[45109]_ ;
  assign \new_[45113]_  = ~A266 & A265;
  assign \new_[45116]_  = A268 & A267;
  assign \new_[45117]_  = \new_[45116]_  & \new_[45113]_ ;
  assign \new_[45118]_  = \new_[45117]_  & \new_[45110]_ ;
  assign \new_[45122]_  = A167 & ~A168;
  assign \new_[45123]_  = ~A170 & \new_[45122]_ ;
  assign \new_[45126]_  = ~A199 & ~A166;
  assign \new_[45129]_  = A232 & A200;
  assign \new_[45130]_  = \new_[45129]_  & \new_[45126]_ ;
  assign \new_[45131]_  = \new_[45130]_  & \new_[45123]_ ;
  assign \new_[45135]_  = A235 & A234;
  assign \new_[45136]_  = ~A233 & \new_[45135]_ ;
  assign \new_[45139]_  = ~A266 & A265;
  assign \new_[45142]_  = A269 & A267;
  assign \new_[45143]_  = \new_[45142]_  & \new_[45139]_ ;
  assign \new_[45144]_  = \new_[45143]_  & \new_[45136]_ ;
  assign \new_[45148]_  = A167 & ~A168;
  assign \new_[45149]_  = ~A170 & \new_[45148]_ ;
  assign \new_[45152]_  = ~A199 & ~A166;
  assign \new_[45155]_  = A232 & A200;
  assign \new_[45156]_  = \new_[45155]_  & \new_[45152]_ ;
  assign \new_[45157]_  = \new_[45156]_  & \new_[45149]_ ;
  assign \new_[45161]_  = A236 & A234;
  assign \new_[45162]_  = ~A233 & \new_[45161]_ ;
  assign \new_[45165]_  = ~A266 & A265;
  assign \new_[45168]_  = A268 & A267;
  assign \new_[45169]_  = \new_[45168]_  & \new_[45165]_ ;
  assign \new_[45170]_  = \new_[45169]_  & \new_[45162]_ ;
  assign \new_[45174]_  = A167 & ~A168;
  assign \new_[45175]_  = ~A170 & \new_[45174]_ ;
  assign \new_[45178]_  = ~A199 & ~A166;
  assign \new_[45181]_  = A232 & A200;
  assign \new_[45182]_  = \new_[45181]_  & \new_[45178]_ ;
  assign \new_[45183]_  = \new_[45182]_  & \new_[45175]_ ;
  assign \new_[45187]_  = A236 & A234;
  assign \new_[45188]_  = ~A233 & \new_[45187]_ ;
  assign \new_[45191]_  = ~A266 & A265;
  assign \new_[45194]_  = A269 & A267;
  assign \new_[45195]_  = \new_[45194]_  & \new_[45191]_ ;
  assign \new_[45196]_  = \new_[45195]_  & \new_[45188]_ ;
  assign \new_[45200]_  = A167 & ~A168;
  assign \new_[45201]_  = ~A170 & \new_[45200]_ ;
  assign \new_[45204]_  = ~A199 & ~A166;
  assign \new_[45207]_  = ~A232 & A200;
  assign \new_[45208]_  = \new_[45207]_  & \new_[45204]_ ;
  assign \new_[45209]_  = \new_[45208]_  & \new_[45201]_ ;
  assign \new_[45213]_  = A266 & A265;
  assign \new_[45214]_  = ~A233 & \new_[45213]_ ;
  assign \new_[45217]_  = ~A299 & A298;
  assign \new_[45220]_  = A301 & A300;
  assign \new_[45221]_  = \new_[45220]_  & \new_[45217]_ ;
  assign \new_[45222]_  = \new_[45221]_  & \new_[45214]_ ;
  assign \new_[45226]_  = A167 & ~A168;
  assign \new_[45227]_  = ~A170 & \new_[45226]_ ;
  assign \new_[45230]_  = ~A199 & ~A166;
  assign \new_[45233]_  = ~A232 & A200;
  assign \new_[45234]_  = \new_[45233]_  & \new_[45230]_ ;
  assign \new_[45235]_  = \new_[45234]_  & \new_[45227]_ ;
  assign \new_[45239]_  = A266 & A265;
  assign \new_[45240]_  = ~A233 & \new_[45239]_ ;
  assign \new_[45243]_  = ~A299 & A298;
  assign \new_[45246]_  = A302 & A300;
  assign \new_[45247]_  = \new_[45246]_  & \new_[45243]_ ;
  assign \new_[45248]_  = \new_[45247]_  & \new_[45240]_ ;
  assign \new_[45252]_  = A167 & ~A168;
  assign \new_[45253]_  = ~A170 & \new_[45252]_ ;
  assign \new_[45256]_  = ~A199 & ~A166;
  assign \new_[45259]_  = ~A232 & A200;
  assign \new_[45260]_  = \new_[45259]_  & \new_[45256]_ ;
  assign \new_[45261]_  = \new_[45260]_  & \new_[45253]_ ;
  assign \new_[45265]_  = ~A267 & ~A266;
  assign \new_[45266]_  = ~A233 & \new_[45265]_ ;
  assign \new_[45269]_  = ~A299 & A298;
  assign \new_[45272]_  = A301 & A300;
  assign \new_[45273]_  = \new_[45272]_  & \new_[45269]_ ;
  assign \new_[45274]_  = \new_[45273]_  & \new_[45266]_ ;
  assign \new_[45278]_  = A167 & ~A168;
  assign \new_[45279]_  = ~A170 & \new_[45278]_ ;
  assign \new_[45282]_  = ~A199 & ~A166;
  assign \new_[45285]_  = ~A232 & A200;
  assign \new_[45286]_  = \new_[45285]_  & \new_[45282]_ ;
  assign \new_[45287]_  = \new_[45286]_  & \new_[45279]_ ;
  assign \new_[45291]_  = ~A267 & ~A266;
  assign \new_[45292]_  = ~A233 & \new_[45291]_ ;
  assign \new_[45295]_  = ~A299 & A298;
  assign \new_[45298]_  = A302 & A300;
  assign \new_[45299]_  = \new_[45298]_  & \new_[45295]_ ;
  assign \new_[45300]_  = \new_[45299]_  & \new_[45292]_ ;
  assign \new_[45304]_  = A167 & ~A168;
  assign \new_[45305]_  = ~A170 & \new_[45304]_ ;
  assign \new_[45308]_  = ~A199 & ~A166;
  assign \new_[45311]_  = ~A232 & A200;
  assign \new_[45312]_  = \new_[45311]_  & \new_[45308]_ ;
  assign \new_[45313]_  = \new_[45312]_  & \new_[45305]_ ;
  assign \new_[45317]_  = ~A266 & ~A265;
  assign \new_[45318]_  = ~A233 & \new_[45317]_ ;
  assign \new_[45321]_  = ~A299 & A298;
  assign \new_[45324]_  = A301 & A300;
  assign \new_[45325]_  = \new_[45324]_  & \new_[45321]_ ;
  assign \new_[45326]_  = \new_[45325]_  & \new_[45318]_ ;
  assign \new_[45330]_  = A167 & ~A168;
  assign \new_[45331]_  = ~A170 & \new_[45330]_ ;
  assign \new_[45334]_  = ~A199 & ~A166;
  assign \new_[45337]_  = ~A232 & A200;
  assign \new_[45338]_  = \new_[45337]_  & \new_[45334]_ ;
  assign \new_[45339]_  = \new_[45338]_  & \new_[45331]_ ;
  assign \new_[45343]_  = ~A266 & ~A265;
  assign \new_[45344]_  = ~A233 & \new_[45343]_ ;
  assign \new_[45347]_  = ~A299 & A298;
  assign \new_[45350]_  = A302 & A300;
  assign \new_[45351]_  = \new_[45350]_  & \new_[45347]_ ;
  assign \new_[45352]_  = \new_[45351]_  & \new_[45344]_ ;
  assign \new_[45356]_  = ~A167 & ~A168;
  assign \new_[45357]_  = ~A170 & \new_[45356]_ ;
  assign \new_[45360]_  = ~A199 & A166;
  assign \new_[45363]_  = A232 & A200;
  assign \new_[45364]_  = \new_[45363]_  & \new_[45360]_ ;
  assign \new_[45365]_  = \new_[45364]_  & \new_[45357]_ ;
  assign \new_[45369]_  = ~A267 & A265;
  assign \new_[45370]_  = A233 & \new_[45369]_ ;
  assign \new_[45373]_  = ~A299 & A298;
  assign \new_[45376]_  = A301 & A300;
  assign \new_[45377]_  = \new_[45376]_  & \new_[45373]_ ;
  assign \new_[45378]_  = \new_[45377]_  & \new_[45370]_ ;
  assign \new_[45382]_  = ~A167 & ~A168;
  assign \new_[45383]_  = ~A170 & \new_[45382]_ ;
  assign \new_[45386]_  = ~A199 & A166;
  assign \new_[45389]_  = A232 & A200;
  assign \new_[45390]_  = \new_[45389]_  & \new_[45386]_ ;
  assign \new_[45391]_  = \new_[45390]_  & \new_[45383]_ ;
  assign \new_[45395]_  = ~A267 & A265;
  assign \new_[45396]_  = A233 & \new_[45395]_ ;
  assign \new_[45399]_  = ~A299 & A298;
  assign \new_[45402]_  = A302 & A300;
  assign \new_[45403]_  = \new_[45402]_  & \new_[45399]_ ;
  assign \new_[45404]_  = \new_[45403]_  & \new_[45396]_ ;
  assign \new_[45408]_  = ~A167 & ~A168;
  assign \new_[45409]_  = ~A170 & \new_[45408]_ ;
  assign \new_[45412]_  = ~A199 & A166;
  assign \new_[45415]_  = A232 & A200;
  assign \new_[45416]_  = \new_[45415]_  & \new_[45412]_ ;
  assign \new_[45417]_  = \new_[45416]_  & \new_[45409]_ ;
  assign \new_[45421]_  = A266 & A265;
  assign \new_[45422]_  = A233 & \new_[45421]_ ;
  assign \new_[45425]_  = ~A299 & A298;
  assign \new_[45428]_  = A301 & A300;
  assign \new_[45429]_  = \new_[45428]_  & \new_[45425]_ ;
  assign \new_[45430]_  = \new_[45429]_  & \new_[45422]_ ;
  assign \new_[45434]_  = ~A167 & ~A168;
  assign \new_[45435]_  = ~A170 & \new_[45434]_ ;
  assign \new_[45438]_  = ~A199 & A166;
  assign \new_[45441]_  = A232 & A200;
  assign \new_[45442]_  = \new_[45441]_  & \new_[45438]_ ;
  assign \new_[45443]_  = \new_[45442]_  & \new_[45435]_ ;
  assign \new_[45447]_  = A266 & A265;
  assign \new_[45448]_  = A233 & \new_[45447]_ ;
  assign \new_[45451]_  = ~A299 & A298;
  assign \new_[45454]_  = A302 & A300;
  assign \new_[45455]_  = \new_[45454]_  & \new_[45451]_ ;
  assign \new_[45456]_  = \new_[45455]_  & \new_[45448]_ ;
  assign \new_[45460]_  = ~A167 & ~A168;
  assign \new_[45461]_  = ~A170 & \new_[45460]_ ;
  assign \new_[45464]_  = ~A199 & A166;
  assign \new_[45467]_  = A232 & A200;
  assign \new_[45468]_  = \new_[45467]_  & \new_[45464]_ ;
  assign \new_[45469]_  = \new_[45468]_  & \new_[45461]_ ;
  assign \new_[45473]_  = ~A266 & ~A265;
  assign \new_[45474]_  = A233 & \new_[45473]_ ;
  assign \new_[45477]_  = ~A299 & A298;
  assign \new_[45480]_  = A301 & A300;
  assign \new_[45481]_  = \new_[45480]_  & \new_[45477]_ ;
  assign \new_[45482]_  = \new_[45481]_  & \new_[45474]_ ;
  assign \new_[45486]_  = ~A167 & ~A168;
  assign \new_[45487]_  = ~A170 & \new_[45486]_ ;
  assign \new_[45490]_  = ~A199 & A166;
  assign \new_[45493]_  = A232 & A200;
  assign \new_[45494]_  = \new_[45493]_  & \new_[45490]_ ;
  assign \new_[45495]_  = \new_[45494]_  & \new_[45487]_ ;
  assign \new_[45499]_  = ~A266 & ~A265;
  assign \new_[45500]_  = A233 & \new_[45499]_ ;
  assign \new_[45503]_  = ~A299 & A298;
  assign \new_[45506]_  = A302 & A300;
  assign \new_[45507]_  = \new_[45506]_  & \new_[45503]_ ;
  assign \new_[45508]_  = \new_[45507]_  & \new_[45500]_ ;
  assign \new_[45512]_  = ~A167 & ~A168;
  assign \new_[45513]_  = ~A170 & \new_[45512]_ ;
  assign \new_[45516]_  = ~A199 & A166;
  assign \new_[45519]_  = ~A233 & A200;
  assign \new_[45520]_  = \new_[45519]_  & \new_[45516]_ ;
  assign \new_[45521]_  = \new_[45520]_  & \new_[45513]_ ;
  assign \new_[45525]_  = ~A266 & ~A236;
  assign \new_[45526]_  = ~A235 & \new_[45525]_ ;
  assign \new_[45529]_  = ~A269 & ~A268;
  assign \new_[45532]_  = A299 & ~A298;
  assign \new_[45533]_  = \new_[45532]_  & \new_[45529]_ ;
  assign \new_[45534]_  = \new_[45533]_  & \new_[45526]_ ;
  assign \new_[45538]_  = ~A167 & ~A168;
  assign \new_[45539]_  = ~A170 & \new_[45538]_ ;
  assign \new_[45542]_  = ~A199 & A166;
  assign \new_[45545]_  = ~A233 & A200;
  assign \new_[45546]_  = \new_[45545]_  & \new_[45542]_ ;
  assign \new_[45547]_  = \new_[45546]_  & \new_[45539]_ ;
  assign \new_[45551]_  = A266 & A265;
  assign \new_[45552]_  = ~A234 & \new_[45551]_ ;
  assign \new_[45555]_  = ~A299 & A298;
  assign \new_[45558]_  = A301 & A300;
  assign \new_[45559]_  = \new_[45558]_  & \new_[45555]_ ;
  assign \new_[45560]_  = \new_[45559]_  & \new_[45552]_ ;
  assign \new_[45564]_  = ~A167 & ~A168;
  assign \new_[45565]_  = ~A170 & \new_[45564]_ ;
  assign \new_[45568]_  = ~A199 & A166;
  assign \new_[45571]_  = ~A233 & A200;
  assign \new_[45572]_  = \new_[45571]_  & \new_[45568]_ ;
  assign \new_[45573]_  = \new_[45572]_  & \new_[45565]_ ;
  assign \new_[45577]_  = A266 & A265;
  assign \new_[45578]_  = ~A234 & \new_[45577]_ ;
  assign \new_[45581]_  = ~A299 & A298;
  assign \new_[45584]_  = A302 & A300;
  assign \new_[45585]_  = \new_[45584]_  & \new_[45581]_ ;
  assign \new_[45586]_  = \new_[45585]_  & \new_[45578]_ ;
  assign \new_[45590]_  = ~A167 & ~A168;
  assign \new_[45591]_  = ~A170 & \new_[45590]_ ;
  assign \new_[45594]_  = ~A199 & A166;
  assign \new_[45597]_  = ~A233 & A200;
  assign \new_[45598]_  = \new_[45597]_  & \new_[45594]_ ;
  assign \new_[45599]_  = \new_[45598]_  & \new_[45591]_ ;
  assign \new_[45603]_  = ~A267 & ~A266;
  assign \new_[45604]_  = ~A234 & \new_[45603]_ ;
  assign \new_[45607]_  = ~A299 & A298;
  assign \new_[45610]_  = A301 & A300;
  assign \new_[45611]_  = \new_[45610]_  & \new_[45607]_ ;
  assign \new_[45612]_  = \new_[45611]_  & \new_[45604]_ ;
  assign \new_[45616]_  = ~A167 & ~A168;
  assign \new_[45617]_  = ~A170 & \new_[45616]_ ;
  assign \new_[45620]_  = ~A199 & A166;
  assign \new_[45623]_  = ~A233 & A200;
  assign \new_[45624]_  = \new_[45623]_  & \new_[45620]_ ;
  assign \new_[45625]_  = \new_[45624]_  & \new_[45617]_ ;
  assign \new_[45629]_  = ~A267 & ~A266;
  assign \new_[45630]_  = ~A234 & \new_[45629]_ ;
  assign \new_[45633]_  = ~A299 & A298;
  assign \new_[45636]_  = A302 & A300;
  assign \new_[45637]_  = \new_[45636]_  & \new_[45633]_ ;
  assign \new_[45638]_  = \new_[45637]_  & \new_[45630]_ ;
  assign \new_[45642]_  = ~A167 & ~A168;
  assign \new_[45643]_  = ~A170 & \new_[45642]_ ;
  assign \new_[45646]_  = ~A199 & A166;
  assign \new_[45649]_  = ~A233 & A200;
  assign \new_[45650]_  = \new_[45649]_  & \new_[45646]_ ;
  assign \new_[45651]_  = \new_[45650]_  & \new_[45643]_ ;
  assign \new_[45655]_  = ~A266 & ~A265;
  assign \new_[45656]_  = ~A234 & \new_[45655]_ ;
  assign \new_[45659]_  = ~A299 & A298;
  assign \new_[45662]_  = A301 & A300;
  assign \new_[45663]_  = \new_[45662]_  & \new_[45659]_ ;
  assign \new_[45664]_  = \new_[45663]_  & \new_[45656]_ ;
  assign \new_[45668]_  = ~A167 & ~A168;
  assign \new_[45669]_  = ~A170 & \new_[45668]_ ;
  assign \new_[45672]_  = ~A199 & A166;
  assign \new_[45675]_  = ~A233 & A200;
  assign \new_[45676]_  = \new_[45675]_  & \new_[45672]_ ;
  assign \new_[45677]_  = \new_[45676]_  & \new_[45669]_ ;
  assign \new_[45681]_  = ~A266 & ~A265;
  assign \new_[45682]_  = ~A234 & \new_[45681]_ ;
  assign \new_[45685]_  = ~A299 & A298;
  assign \new_[45688]_  = A302 & A300;
  assign \new_[45689]_  = \new_[45688]_  & \new_[45685]_ ;
  assign \new_[45690]_  = \new_[45689]_  & \new_[45682]_ ;
  assign \new_[45694]_  = ~A167 & ~A168;
  assign \new_[45695]_  = ~A170 & \new_[45694]_ ;
  assign \new_[45698]_  = ~A199 & A166;
  assign \new_[45701]_  = A232 & A200;
  assign \new_[45702]_  = \new_[45701]_  & \new_[45698]_ ;
  assign \new_[45703]_  = \new_[45702]_  & \new_[45695]_ ;
  assign \new_[45707]_  = A235 & A234;
  assign \new_[45708]_  = ~A233 & \new_[45707]_ ;
  assign \new_[45711]_  = ~A266 & A265;
  assign \new_[45714]_  = A268 & A267;
  assign \new_[45715]_  = \new_[45714]_  & \new_[45711]_ ;
  assign \new_[45716]_  = \new_[45715]_  & \new_[45708]_ ;
  assign \new_[45720]_  = ~A167 & ~A168;
  assign \new_[45721]_  = ~A170 & \new_[45720]_ ;
  assign \new_[45724]_  = ~A199 & A166;
  assign \new_[45727]_  = A232 & A200;
  assign \new_[45728]_  = \new_[45727]_  & \new_[45724]_ ;
  assign \new_[45729]_  = \new_[45728]_  & \new_[45721]_ ;
  assign \new_[45733]_  = A235 & A234;
  assign \new_[45734]_  = ~A233 & \new_[45733]_ ;
  assign \new_[45737]_  = ~A266 & A265;
  assign \new_[45740]_  = A269 & A267;
  assign \new_[45741]_  = \new_[45740]_  & \new_[45737]_ ;
  assign \new_[45742]_  = \new_[45741]_  & \new_[45734]_ ;
  assign \new_[45746]_  = ~A167 & ~A168;
  assign \new_[45747]_  = ~A170 & \new_[45746]_ ;
  assign \new_[45750]_  = ~A199 & A166;
  assign \new_[45753]_  = A232 & A200;
  assign \new_[45754]_  = \new_[45753]_  & \new_[45750]_ ;
  assign \new_[45755]_  = \new_[45754]_  & \new_[45747]_ ;
  assign \new_[45759]_  = A236 & A234;
  assign \new_[45760]_  = ~A233 & \new_[45759]_ ;
  assign \new_[45763]_  = ~A266 & A265;
  assign \new_[45766]_  = A268 & A267;
  assign \new_[45767]_  = \new_[45766]_  & \new_[45763]_ ;
  assign \new_[45768]_  = \new_[45767]_  & \new_[45760]_ ;
  assign \new_[45772]_  = ~A167 & ~A168;
  assign \new_[45773]_  = ~A170 & \new_[45772]_ ;
  assign \new_[45776]_  = ~A199 & A166;
  assign \new_[45779]_  = A232 & A200;
  assign \new_[45780]_  = \new_[45779]_  & \new_[45776]_ ;
  assign \new_[45781]_  = \new_[45780]_  & \new_[45773]_ ;
  assign \new_[45785]_  = A236 & A234;
  assign \new_[45786]_  = ~A233 & \new_[45785]_ ;
  assign \new_[45789]_  = ~A266 & A265;
  assign \new_[45792]_  = A269 & A267;
  assign \new_[45793]_  = \new_[45792]_  & \new_[45789]_ ;
  assign \new_[45794]_  = \new_[45793]_  & \new_[45786]_ ;
  assign \new_[45798]_  = ~A167 & ~A168;
  assign \new_[45799]_  = ~A170 & \new_[45798]_ ;
  assign \new_[45802]_  = ~A199 & A166;
  assign \new_[45805]_  = ~A232 & A200;
  assign \new_[45806]_  = \new_[45805]_  & \new_[45802]_ ;
  assign \new_[45807]_  = \new_[45806]_  & \new_[45799]_ ;
  assign \new_[45811]_  = A266 & A265;
  assign \new_[45812]_  = ~A233 & \new_[45811]_ ;
  assign \new_[45815]_  = ~A299 & A298;
  assign \new_[45818]_  = A301 & A300;
  assign \new_[45819]_  = \new_[45818]_  & \new_[45815]_ ;
  assign \new_[45820]_  = \new_[45819]_  & \new_[45812]_ ;
  assign \new_[45824]_  = ~A167 & ~A168;
  assign \new_[45825]_  = ~A170 & \new_[45824]_ ;
  assign \new_[45828]_  = ~A199 & A166;
  assign \new_[45831]_  = ~A232 & A200;
  assign \new_[45832]_  = \new_[45831]_  & \new_[45828]_ ;
  assign \new_[45833]_  = \new_[45832]_  & \new_[45825]_ ;
  assign \new_[45837]_  = A266 & A265;
  assign \new_[45838]_  = ~A233 & \new_[45837]_ ;
  assign \new_[45841]_  = ~A299 & A298;
  assign \new_[45844]_  = A302 & A300;
  assign \new_[45845]_  = \new_[45844]_  & \new_[45841]_ ;
  assign \new_[45846]_  = \new_[45845]_  & \new_[45838]_ ;
  assign \new_[45850]_  = ~A167 & ~A168;
  assign \new_[45851]_  = ~A170 & \new_[45850]_ ;
  assign \new_[45854]_  = ~A199 & A166;
  assign \new_[45857]_  = ~A232 & A200;
  assign \new_[45858]_  = \new_[45857]_  & \new_[45854]_ ;
  assign \new_[45859]_  = \new_[45858]_  & \new_[45851]_ ;
  assign \new_[45863]_  = ~A267 & ~A266;
  assign \new_[45864]_  = ~A233 & \new_[45863]_ ;
  assign \new_[45867]_  = ~A299 & A298;
  assign \new_[45870]_  = A301 & A300;
  assign \new_[45871]_  = \new_[45870]_  & \new_[45867]_ ;
  assign \new_[45872]_  = \new_[45871]_  & \new_[45864]_ ;
  assign \new_[45876]_  = ~A167 & ~A168;
  assign \new_[45877]_  = ~A170 & \new_[45876]_ ;
  assign \new_[45880]_  = ~A199 & A166;
  assign \new_[45883]_  = ~A232 & A200;
  assign \new_[45884]_  = \new_[45883]_  & \new_[45880]_ ;
  assign \new_[45885]_  = \new_[45884]_  & \new_[45877]_ ;
  assign \new_[45889]_  = ~A267 & ~A266;
  assign \new_[45890]_  = ~A233 & \new_[45889]_ ;
  assign \new_[45893]_  = ~A299 & A298;
  assign \new_[45896]_  = A302 & A300;
  assign \new_[45897]_  = \new_[45896]_  & \new_[45893]_ ;
  assign \new_[45898]_  = \new_[45897]_  & \new_[45890]_ ;
  assign \new_[45902]_  = ~A167 & ~A168;
  assign \new_[45903]_  = ~A170 & \new_[45902]_ ;
  assign \new_[45906]_  = ~A199 & A166;
  assign \new_[45909]_  = ~A232 & A200;
  assign \new_[45910]_  = \new_[45909]_  & \new_[45906]_ ;
  assign \new_[45911]_  = \new_[45910]_  & \new_[45903]_ ;
  assign \new_[45915]_  = ~A266 & ~A265;
  assign \new_[45916]_  = ~A233 & \new_[45915]_ ;
  assign \new_[45919]_  = ~A299 & A298;
  assign \new_[45922]_  = A301 & A300;
  assign \new_[45923]_  = \new_[45922]_  & \new_[45919]_ ;
  assign \new_[45924]_  = \new_[45923]_  & \new_[45916]_ ;
  assign \new_[45928]_  = ~A167 & ~A168;
  assign \new_[45929]_  = ~A170 & \new_[45928]_ ;
  assign \new_[45932]_  = ~A199 & A166;
  assign \new_[45935]_  = ~A232 & A200;
  assign \new_[45936]_  = \new_[45935]_  & \new_[45932]_ ;
  assign \new_[45937]_  = \new_[45936]_  & \new_[45929]_ ;
  assign \new_[45941]_  = ~A266 & ~A265;
  assign \new_[45942]_  = ~A233 & \new_[45941]_ ;
  assign \new_[45945]_  = ~A299 & A298;
  assign \new_[45948]_  = A302 & A300;
  assign \new_[45949]_  = \new_[45948]_  & \new_[45945]_ ;
  assign \new_[45950]_  = \new_[45949]_  & \new_[45942]_ ;
  assign \new_[45954]_  = A167 & ~A168;
  assign \new_[45955]_  = A169 & \new_[45954]_ ;
  assign \new_[45958]_  = ~A199 & ~A166;
  assign \new_[45961]_  = A232 & A200;
  assign \new_[45962]_  = \new_[45961]_  & \new_[45958]_ ;
  assign \new_[45963]_  = \new_[45962]_  & \new_[45955]_ ;
  assign \new_[45967]_  = ~A267 & A265;
  assign \new_[45968]_  = A233 & \new_[45967]_ ;
  assign \new_[45971]_  = ~A299 & A298;
  assign \new_[45974]_  = A301 & A300;
  assign \new_[45975]_  = \new_[45974]_  & \new_[45971]_ ;
  assign \new_[45976]_  = \new_[45975]_  & \new_[45968]_ ;
  assign \new_[45980]_  = A167 & ~A168;
  assign \new_[45981]_  = A169 & \new_[45980]_ ;
  assign \new_[45984]_  = ~A199 & ~A166;
  assign \new_[45987]_  = A232 & A200;
  assign \new_[45988]_  = \new_[45987]_  & \new_[45984]_ ;
  assign \new_[45989]_  = \new_[45988]_  & \new_[45981]_ ;
  assign \new_[45993]_  = ~A267 & A265;
  assign \new_[45994]_  = A233 & \new_[45993]_ ;
  assign \new_[45997]_  = ~A299 & A298;
  assign \new_[46000]_  = A302 & A300;
  assign \new_[46001]_  = \new_[46000]_  & \new_[45997]_ ;
  assign \new_[46002]_  = \new_[46001]_  & \new_[45994]_ ;
  assign \new_[46006]_  = A167 & ~A168;
  assign \new_[46007]_  = A169 & \new_[46006]_ ;
  assign \new_[46010]_  = ~A199 & ~A166;
  assign \new_[46013]_  = A232 & A200;
  assign \new_[46014]_  = \new_[46013]_  & \new_[46010]_ ;
  assign \new_[46015]_  = \new_[46014]_  & \new_[46007]_ ;
  assign \new_[46019]_  = A266 & A265;
  assign \new_[46020]_  = A233 & \new_[46019]_ ;
  assign \new_[46023]_  = ~A299 & A298;
  assign \new_[46026]_  = A301 & A300;
  assign \new_[46027]_  = \new_[46026]_  & \new_[46023]_ ;
  assign \new_[46028]_  = \new_[46027]_  & \new_[46020]_ ;
  assign \new_[46032]_  = A167 & ~A168;
  assign \new_[46033]_  = A169 & \new_[46032]_ ;
  assign \new_[46036]_  = ~A199 & ~A166;
  assign \new_[46039]_  = A232 & A200;
  assign \new_[46040]_  = \new_[46039]_  & \new_[46036]_ ;
  assign \new_[46041]_  = \new_[46040]_  & \new_[46033]_ ;
  assign \new_[46045]_  = A266 & A265;
  assign \new_[46046]_  = A233 & \new_[46045]_ ;
  assign \new_[46049]_  = ~A299 & A298;
  assign \new_[46052]_  = A302 & A300;
  assign \new_[46053]_  = \new_[46052]_  & \new_[46049]_ ;
  assign \new_[46054]_  = \new_[46053]_  & \new_[46046]_ ;
  assign \new_[46058]_  = A167 & ~A168;
  assign \new_[46059]_  = A169 & \new_[46058]_ ;
  assign \new_[46062]_  = ~A199 & ~A166;
  assign \new_[46065]_  = A232 & A200;
  assign \new_[46066]_  = \new_[46065]_  & \new_[46062]_ ;
  assign \new_[46067]_  = \new_[46066]_  & \new_[46059]_ ;
  assign \new_[46071]_  = ~A266 & ~A265;
  assign \new_[46072]_  = A233 & \new_[46071]_ ;
  assign \new_[46075]_  = ~A299 & A298;
  assign \new_[46078]_  = A301 & A300;
  assign \new_[46079]_  = \new_[46078]_  & \new_[46075]_ ;
  assign \new_[46080]_  = \new_[46079]_  & \new_[46072]_ ;
  assign \new_[46084]_  = A167 & ~A168;
  assign \new_[46085]_  = A169 & \new_[46084]_ ;
  assign \new_[46088]_  = ~A199 & ~A166;
  assign \new_[46091]_  = A232 & A200;
  assign \new_[46092]_  = \new_[46091]_  & \new_[46088]_ ;
  assign \new_[46093]_  = \new_[46092]_  & \new_[46085]_ ;
  assign \new_[46097]_  = ~A266 & ~A265;
  assign \new_[46098]_  = A233 & \new_[46097]_ ;
  assign \new_[46101]_  = ~A299 & A298;
  assign \new_[46104]_  = A302 & A300;
  assign \new_[46105]_  = \new_[46104]_  & \new_[46101]_ ;
  assign \new_[46106]_  = \new_[46105]_  & \new_[46098]_ ;
  assign \new_[46110]_  = A167 & ~A168;
  assign \new_[46111]_  = A169 & \new_[46110]_ ;
  assign \new_[46114]_  = ~A199 & ~A166;
  assign \new_[46117]_  = ~A233 & A200;
  assign \new_[46118]_  = \new_[46117]_  & \new_[46114]_ ;
  assign \new_[46119]_  = \new_[46118]_  & \new_[46111]_ ;
  assign \new_[46123]_  = ~A266 & ~A236;
  assign \new_[46124]_  = ~A235 & \new_[46123]_ ;
  assign \new_[46127]_  = ~A269 & ~A268;
  assign \new_[46130]_  = A299 & ~A298;
  assign \new_[46131]_  = \new_[46130]_  & \new_[46127]_ ;
  assign \new_[46132]_  = \new_[46131]_  & \new_[46124]_ ;
  assign \new_[46136]_  = A167 & ~A168;
  assign \new_[46137]_  = A169 & \new_[46136]_ ;
  assign \new_[46140]_  = ~A199 & ~A166;
  assign \new_[46143]_  = ~A233 & A200;
  assign \new_[46144]_  = \new_[46143]_  & \new_[46140]_ ;
  assign \new_[46145]_  = \new_[46144]_  & \new_[46137]_ ;
  assign \new_[46149]_  = A266 & A265;
  assign \new_[46150]_  = ~A234 & \new_[46149]_ ;
  assign \new_[46153]_  = ~A299 & A298;
  assign \new_[46156]_  = A301 & A300;
  assign \new_[46157]_  = \new_[46156]_  & \new_[46153]_ ;
  assign \new_[46158]_  = \new_[46157]_  & \new_[46150]_ ;
  assign \new_[46162]_  = A167 & ~A168;
  assign \new_[46163]_  = A169 & \new_[46162]_ ;
  assign \new_[46166]_  = ~A199 & ~A166;
  assign \new_[46169]_  = ~A233 & A200;
  assign \new_[46170]_  = \new_[46169]_  & \new_[46166]_ ;
  assign \new_[46171]_  = \new_[46170]_  & \new_[46163]_ ;
  assign \new_[46175]_  = A266 & A265;
  assign \new_[46176]_  = ~A234 & \new_[46175]_ ;
  assign \new_[46179]_  = ~A299 & A298;
  assign \new_[46182]_  = A302 & A300;
  assign \new_[46183]_  = \new_[46182]_  & \new_[46179]_ ;
  assign \new_[46184]_  = \new_[46183]_  & \new_[46176]_ ;
  assign \new_[46188]_  = A167 & ~A168;
  assign \new_[46189]_  = A169 & \new_[46188]_ ;
  assign \new_[46192]_  = ~A199 & ~A166;
  assign \new_[46195]_  = ~A233 & A200;
  assign \new_[46196]_  = \new_[46195]_  & \new_[46192]_ ;
  assign \new_[46197]_  = \new_[46196]_  & \new_[46189]_ ;
  assign \new_[46201]_  = ~A267 & ~A266;
  assign \new_[46202]_  = ~A234 & \new_[46201]_ ;
  assign \new_[46205]_  = ~A299 & A298;
  assign \new_[46208]_  = A301 & A300;
  assign \new_[46209]_  = \new_[46208]_  & \new_[46205]_ ;
  assign \new_[46210]_  = \new_[46209]_  & \new_[46202]_ ;
  assign \new_[46214]_  = A167 & ~A168;
  assign \new_[46215]_  = A169 & \new_[46214]_ ;
  assign \new_[46218]_  = ~A199 & ~A166;
  assign \new_[46221]_  = ~A233 & A200;
  assign \new_[46222]_  = \new_[46221]_  & \new_[46218]_ ;
  assign \new_[46223]_  = \new_[46222]_  & \new_[46215]_ ;
  assign \new_[46227]_  = ~A267 & ~A266;
  assign \new_[46228]_  = ~A234 & \new_[46227]_ ;
  assign \new_[46231]_  = ~A299 & A298;
  assign \new_[46234]_  = A302 & A300;
  assign \new_[46235]_  = \new_[46234]_  & \new_[46231]_ ;
  assign \new_[46236]_  = \new_[46235]_  & \new_[46228]_ ;
  assign \new_[46240]_  = A167 & ~A168;
  assign \new_[46241]_  = A169 & \new_[46240]_ ;
  assign \new_[46244]_  = ~A199 & ~A166;
  assign \new_[46247]_  = ~A233 & A200;
  assign \new_[46248]_  = \new_[46247]_  & \new_[46244]_ ;
  assign \new_[46249]_  = \new_[46248]_  & \new_[46241]_ ;
  assign \new_[46253]_  = ~A266 & ~A265;
  assign \new_[46254]_  = ~A234 & \new_[46253]_ ;
  assign \new_[46257]_  = ~A299 & A298;
  assign \new_[46260]_  = A301 & A300;
  assign \new_[46261]_  = \new_[46260]_  & \new_[46257]_ ;
  assign \new_[46262]_  = \new_[46261]_  & \new_[46254]_ ;
  assign \new_[46266]_  = A167 & ~A168;
  assign \new_[46267]_  = A169 & \new_[46266]_ ;
  assign \new_[46270]_  = ~A199 & ~A166;
  assign \new_[46273]_  = ~A233 & A200;
  assign \new_[46274]_  = \new_[46273]_  & \new_[46270]_ ;
  assign \new_[46275]_  = \new_[46274]_  & \new_[46267]_ ;
  assign \new_[46279]_  = ~A266 & ~A265;
  assign \new_[46280]_  = ~A234 & \new_[46279]_ ;
  assign \new_[46283]_  = ~A299 & A298;
  assign \new_[46286]_  = A302 & A300;
  assign \new_[46287]_  = \new_[46286]_  & \new_[46283]_ ;
  assign \new_[46288]_  = \new_[46287]_  & \new_[46280]_ ;
  assign \new_[46292]_  = A167 & ~A168;
  assign \new_[46293]_  = A169 & \new_[46292]_ ;
  assign \new_[46296]_  = ~A199 & ~A166;
  assign \new_[46299]_  = A232 & A200;
  assign \new_[46300]_  = \new_[46299]_  & \new_[46296]_ ;
  assign \new_[46301]_  = \new_[46300]_  & \new_[46293]_ ;
  assign \new_[46305]_  = A235 & A234;
  assign \new_[46306]_  = ~A233 & \new_[46305]_ ;
  assign \new_[46309]_  = ~A266 & A265;
  assign \new_[46312]_  = A268 & A267;
  assign \new_[46313]_  = \new_[46312]_  & \new_[46309]_ ;
  assign \new_[46314]_  = \new_[46313]_  & \new_[46306]_ ;
  assign \new_[46318]_  = A167 & ~A168;
  assign \new_[46319]_  = A169 & \new_[46318]_ ;
  assign \new_[46322]_  = ~A199 & ~A166;
  assign \new_[46325]_  = A232 & A200;
  assign \new_[46326]_  = \new_[46325]_  & \new_[46322]_ ;
  assign \new_[46327]_  = \new_[46326]_  & \new_[46319]_ ;
  assign \new_[46331]_  = A235 & A234;
  assign \new_[46332]_  = ~A233 & \new_[46331]_ ;
  assign \new_[46335]_  = ~A266 & A265;
  assign \new_[46338]_  = A269 & A267;
  assign \new_[46339]_  = \new_[46338]_  & \new_[46335]_ ;
  assign \new_[46340]_  = \new_[46339]_  & \new_[46332]_ ;
  assign \new_[46344]_  = A167 & ~A168;
  assign \new_[46345]_  = A169 & \new_[46344]_ ;
  assign \new_[46348]_  = ~A199 & ~A166;
  assign \new_[46351]_  = A232 & A200;
  assign \new_[46352]_  = \new_[46351]_  & \new_[46348]_ ;
  assign \new_[46353]_  = \new_[46352]_  & \new_[46345]_ ;
  assign \new_[46357]_  = A236 & A234;
  assign \new_[46358]_  = ~A233 & \new_[46357]_ ;
  assign \new_[46361]_  = ~A266 & A265;
  assign \new_[46364]_  = A268 & A267;
  assign \new_[46365]_  = \new_[46364]_  & \new_[46361]_ ;
  assign \new_[46366]_  = \new_[46365]_  & \new_[46358]_ ;
  assign \new_[46370]_  = A167 & ~A168;
  assign \new_[46371]_  = A169 & \new_[46370]_ ;
  assign \new_[46374]_  = ~A199 & ~A166;
  assign \new_[46377]_  = A232 & A200;
  assign \new_[46378]_  = \new_[46377]_  & \new_[46374]_ ;
  assign \new_[46379]_  = \new_[46378]_  & \new_[46371]_ ;
  assign \new_[46383]_  = A236 & A234;
  assign \new_[46384]_  = ~A233 & \new_[46383]_ ;
  assign \new_[46387]_  = ~A266 & A265;
  assign \new_[46390]_  = A269 & A267;
  assign \new_[46391]_  = \new_[46390]_  & \new_[46387]_ ;
  assign \new_[46392]_  = \new_[46391]_  & \new_[46384]_ ;
  assign \new_[46396]_  = A167 & ~A168;
  assign \new_[46397]_  = A169 & \new_[46396]_ ;
  assign \new_[46400]_  = ~A199 & ~A166;
  assign \new_[46403]_  = ~A232 & A200;
  assign \new_[46404]_  = \new_[46403]_  & \new_[46400]_ ;
  assign \new_[46405]_  = \new_[46404]_  & \new_[46397]_ ;
  assign \new_[46409]_  = A266 & A265;
  assign \new_[46410]_  = ~A233 & \new_[46409]_ ;
  assign \new_[46413]_  = ~A299 & A298;
  assign \new_[46416]_  = A301 & A300;
  assign \new_[46417]_  = \new_[46416]_  & \new_[46413]_ ;
  assign \new_[46418]_  = \new_[46417]_  & \new_[46410]_ ;
  assign \new_[46422]_  = A167 & ~A168;
  assign \new_[46423]_  = A169 & \new_[46422]_ ;
  assign \new_[46426]_  = ~A199 & ~A166;
  assign \new_[46429]_  = ~A232 & A200;
  assign \new_[46430]_  = \new_[46429]_  & \new_[46426]_ ;
  assign \new_[46431]_  = \new_[46430]_  & \new_[46423]_ ;
  assign \new_[46435]_  = A266 & A265;
  assign \new_[46436]_  = ~A233 & \new_[46435]_ ;
  assign \new_[46439]_  = ~A299 & A298;
  assign \new_[46442]_  = A302 & A300;
  assign \new_[46443]_  = \new_[46442]_  & \new_[46439]_ ;
  assign \new_[46444]_  = \new_[46443]_  & \new_[46436]_ ;
  assign \new_[46448]_  = A167 & ~A168;
  assign \new_[46449]_  = A169 & \new_[46448]_ ;
  assign \new_[46452]_  = ~A199 & ~A166;
  assign \new_[46455]_  = ~A232 & A200;
  assign \new_[46456]_  = \new_[46455]_  & \new_[46452]_ ;
  assign \new_[46457]_  = \new_[46456]_  & \new_[46449]_ ;
  assign \new_[46461]_  = ~A267 & ~A266;
  assign \new_[46462]_  = ~A233 & \new_[46461]_ ;
  assign \new_[46465]_  = ~A299 & A298;
  assign \new_[46468]_  = A301 & A300;
  assign \new_[46469]_  = \new_[46468]_  & \new_[46465]_ ;
  assign \new_[46470]_  = \new_[46469]_  & \new_[46462]_ ;
  assign \new_[46474]_  = A167 & ~A168;
  assign \new_[46475]_  = A169 & \new_[46474]_ ;
  assign \new_[46478]_  = ~A199 & ~A166;
  assign \new_[46481]_  = ~A232 & A200;
  assign \new_[46482]_  = \new_[46481]_  & \new_[46478]_ ;
  assign \new_[46483]_  = \new_[46482]_  & \new_[46475]_ ;
  assign \new_[46487]_  = ~A267 & ~A266;
  assign \new_[46488]_  = ~A233 & \new_[46487]_ ;
  assign \new_[46491]_  = ~A299 & A298;
  assign \new_[46494]_  = A302 & A300;
  assign \new_[46495]_  = \new_[46494]_  & \new_[46491]_ ;
  assign \new_[46496]_  = \new_[46495]_  & \new_[46488]_ ;
  assign \new_[46500]_  = A167 & ~A168;
  assign \new_[46501]_  = A169 & \new_[46500]_ ;
  assign \new_[46504]_  = ~A199 & ~A166;
  assign \new_[46507]_  = ~A232 & A200;
  assign \new_[46508]_  = \new_[46507]_  & \new_[46504]_ ;
  assign \new_[46509]_  = \new_[46508]_  & \new_[46501]_ ;
  assign \new_[46513]_  = ~A266 & ~A265;
  assign \new_[46514]_  = ~A233 & \new_[46513]_ ;
  assign \new_[46517]_  = ~A299 & A298;
  assign \new_[46520]_  = A301 & A300;
  assign \new_[46521]_  = \new_[46520]_  & \new_[46517]_ ;
  assign \new_[46522]_  = \new_[46521]_  & \new_[46514]_ ;
  assign \new_[46526]_  = A167 & ~A168;
  assign \new_[46527]_  = A169 & \new_[46526]_ ;
  assign \new_[46530]_  = ~A199 & ~A166;
  assign \new_[46533]_  = ~A232 & A200;
  assign \new_[46534]_  = \new_[46533]_  & \new_[46530]_ ;
  assign \new_[46535]_  = \new_[46534]_  & \new_[46527]_ ;
  assign \new_[46539]_  = ~A266 & ~A265;
  assign \new_[46540]_  = ~A233 & \new_[46539]_ ;
  assign \new_[46543]_  = ~A299 & A298;
  assign \new_[46546]_  = A302 & A300;
  assign \new_[46547]_  = \new_[46546]_  & \new_[46543]_ ;
  assign \new_[46548]_  = \new_[46547]_  & \new_[46540]_ ;
  assign \new_[46552]_  = A167 & ~A168;
  assign \new_[46553]_  = A169 & \new_[46552]_ ;
  assign \new_[46556]_  = A199 & ~A166;
  assign \new_[46559]_  = A201 & ~A200;
  assign \new_[46560]_  = \new_[46559]_  & \new_[46556]_ ;
  assign \new_[46561]_  = \new_[46560]_  & \new_[46553]_ ;
  assign \new_[46565]_  = A233 & A232;
  assign \new_[46566]_  = A202 & \new_[46565]_ ;
  assign \new_[46569]_  = ~A267 & A265;
  assign \new_[46572]_  = A299 & ~A298;
  assign \new_[46573]_  = \new_[46572]_  & \new_[46569]_ ;
  assign \new_[46574]_  = \new_[46573]_  & \new_[46566]_ ;
  assign \new_[46578]_  = A167 & ~A168;
  assign \new_[46579]_  = A169 & \new_[46578]_ ;
  assign \new_[46582]_  = A199 & ~A166;
  assign \new_[46585]_  = A201 & ~A200;
  assign \new_[46586]_  = \new_[46585]_  & \new_[46582]_ ;
  assign \new_[46587]_  = \new_[46586]_  & \new_[46579]_ ;
  assign \new_[46591]_  = A233 & A232;
  assign \new_[46592]_  = A202 & \new_[46591]_ ;
  assign \new_[46595]_  = A266 & A265;
  assign \new_[46598]_  = A299 & ~A298;
  assign \new_[46599]_  = \new_[46598]_  & \new_[46595]_ ;
  assign \new_[46600]_  = \new_[46599]_  & \new_[46592]_ ;
  assign \new_[46604]_  = A167 & ~A168;
  assign \new_[46605]_  = A169 & \new_[46604]_ ;
  assign \new_[46608]_  = A199 & ~A166;
  assign \new_[46611]_  = A201 & ~A200;
  assign \new_[46612]_  = \new_[46611]_  & \new_[46608]_ ;
  assign \new_[46613]_  = \new_[46612]_  & \new_[46605]_ ;
  assign \new_[46617]_  = A233 & A232;
  assign \new_[46618]_  = A202 & \new_[46617]_ ;
  assign \new_[46621]_  = ~A266 & ~A265;
  assign \new_[46624]_  = A299 & ~A298;
  assign \new_[46625]_  = \new_[46624]_  & \new_[46621]_ ;
  assign \new_[46626]_  = \new_[46625]_  & \new_[46618]_ ;
  assign \new_[46630]_  = A167 & ~A168;
  assign \new_[46631]_  = A169 & \new_[46630]_ ;
  assign \new_[46634]_  = A199 & ~A166;
  assign \new_[46637]_  = A201 & ~A200;
  assign \new_[46638]_  = \new_[46637]_  & \new_[46634]_ ;
  assign \new_[46639]_  = \new_[46638]_  & \new_[46631]_ ;
  assign \new_[46643]_  = A233 & ~A232;
  assign \new_[46644]_  = A202 & \new_[46643]_ ;
  assign \new_[46647]_  = ~A266 & A265;
  assign \new_[46650]_  = A268 & A267;
  assign \new_[46651]_  = \new_[46650]_  & \new_[46647]_ ;
  assign \new_[46652]_  = \new_[46651]_  & \new_[46644]_ ;
  assign \new_[46656]_  = A167 & ~A168;
  assign \new_[46657]_  = A169 & \new_[46656]_ ;
  assign \new_[46660]_  = A199 & ~A166;
  assign \new_[46663]_  = A201 & ~A200;
  assign \new_[46664]_  = \new_[46663]_  & \new_[46660]_ ;
  assign \new_[46665]_  = \new_[46664]_  & \new_[46657]_ ;
  assign \new_[46669]_  = A233 & ~A232;
  assign \new_[46670]_  = A202 & \new_[46669]_ ;
  assign \new_[46673]_  = ~A266 & A265;
  assign \new_[46676]_  = A269 & A267;
  assign \new_[46677]_  = \new_[46676]_  & \new_[46673]_ ;
  assign \new_[46678]_  = \new_[46677]_  & \new_[46670]_ ;
  assign \new_[46682]_  = A167 & ~A168;
  assign \new_[46683]_  = A169 & \new_[46682]_ ;
  assign \new_[46686]_  = A199 & ~A166;
  assign \new_[46689]_  = A201 & ~A200;
  assign \new_[46690]_  = \new_[46689]_  & \new_[46686]_ ;
  assign \new_[46691]_  = \new_[46690]_  & \new_[46683]_ ;
  assign \new_[46695]_  = ~A234 & ~A233;
  assign \new_[46696]_  = A202 & \new_[46695]_ ;
  assign \new_[46699]_  = A266 & A265;
  assign \new_[46702]_  = A299 & ~A298;
  assign \new_[46703]_  = \new_[46702]_  & \new_[46699]_ ;
  assign \new_[46704]_  = \new_[46703]_  & \new_[46696]_ ;
  assign \new_[46708]_  = A167 & ~A168;
  assign \new_[46709]_  = A169 & \new_[46708]_ ;
  assign \new_[46712]_  = A199 & ~A166;
  assign \new_[46715]_  = A201 & ~A200;
  assign \new_[46716]_  = \new_[46715]_  & \new_[46712]_ ;
  assign \new_[46717]_  = \new_[46716]_  & \new_[46709]_ ;
  assign \new_[46721]_  = ~A234 & ~A233;
  assign \new_[46722]_  = A202 & \new_[46721]_ ;
  assign \new_[46725]_  = ~A267 & ~A266;
  assign \new_[46728]_  = A299 & ~A298;
  assign \new_[46729]_  = \new_[46728]_  & \new_[46725]_ ;
  assign \new_[46730]_  = \new_[46729]_  & \new_[46722]_ ;
  assign \new_[46734]_  = A167 & ~A168;
  assign \new_[46735]_  = A169 & \new_[46734]_ ;
  assign \new_[46738]_  = A199 & ~A166;
  assign \new_[46741]_  = A201 & ~A200;
  assign \new_[46742]_  = \new_[46741]_  & \new_[46738]_ ;
  assign \new_[46743]_  = \new_[46742]_  & \new_[46735]_ ;
  assign \new_[46747]_  = ~A234 & ~A233;
  assign \new_[46748]_  = A202 & \new_[46747]_ ;
  assign \new_[46751]_  = ~A266 & ~A265;
  assign \new_[46754]_  = A299 & ~A298;
  assign \new_[46755]_  = \new_[46754]_  & \new_[46751]_ ;
  assign \new_[46756]_  = \new_[46755]_  & \new_[46748]_ ;
  assign \new_[46760]_  = A167 & ~A168;
  assign \new_[46761]_  = A169 & \new_[46760]_ ;
  assign \new_[46764]_  = A199 & ~A166;
  assign \new_[46767]_  = A201 & ~A200;
  assign \new_[46768]_  = \new_[46767]_  & \new_[46764]_ ;
  assign \new_[46769]_  = \new_[46768]_  & \new_[46761]_ ;
  assign \new_[46773]_  = ~A233 & A232;
  assign \new_[46774]_  = A202 & \new_[46773]_ ;
  assign \new_[46777]_  = A235 & A234;
  assign \new_[46780]_  = ~A300 & A298;
  assign \new_[46781]_  = \new_[46780]_  & \new_[46777]_ ;
  assign \new_[46782]_  = \new_[46781]_  & \new_[46774]_ ;
  assign \new_[46786]_  = A167 & ~A168;
  assign \new_[46787]_  = A169 & \new_[46786]_ ;
  assign \new_[46790]_  = A199 & ~A166;
  assign \new_[46793]_  = A201 & ~A200;
  assign \new_[46794]_  = \new_[46793]_  & \new_[46790]_ ;
  assign \new_[46795]_  = \new_[46794]_  & \new_[46787]_ ;
  assign \new_[46799]_  = ~A233 & A232;
  assign \new_[46800]_  = A202 & \new_[46799]_ ;
  assign \new_[46803]_  = A235 & A234;
  assign \new_[46806]_  = A299 & A298;
  assign \new_[46807]_  = \new_[46806]_  & \new_[46803]_ ;
  assign \new_[46808]_  = \new_[46807]_  & \new_[46800]_ ;
  assign \new_[46812]_  = A167 & ~A168;
  assign \new_[46813]_  = A169 & \new_[46812]_ ;
  assign \new_[46816]_  = A199 & ~A166;
  assign \new_[46819]_  = A201 & ~A200;
  assign \new_[46820]_  = \new_[46819]_  & \new_[46816]_ ;
  assign \new_[46821]_  = \new_[46820]_  & \new_[46813]_ ;
  assign \new_[46825]_  = ~A233 & A232;
  assign \new_[46826]_  = A202 & \new_[46825]_ ;
  assign \new_[46829]_  = A235 & A234;
  assign \new_[46832]_  = ~A299 & ~A298;
  assign \new_[46833]_  = \new_[46832]_  & \new_[46829]_ ;
  assign \new_[46834]_  = \new_[46833]_  & \new_[46826]_ ;
  assign \new_[46838]_  = A167 & ~A168;
  assign \new_[46839]_  = A169 & \new_[46838]_ ;
  assign \new_[46842]_  = A199 & ~A166;
  assign \new_[46845]_  = A201 & ~A200;
  assign \new_[46846]_  = \new_[46845]_  & \new_[46842]_ ;
  assign \new_[46847]_  = \new_[46846]_  & \new_[46839]_ ;
  assign \new_[46851]_  = ~A233 & A232;
  assign \new_[46852]_  = A202 & \new_[46851]_ ;
  assign \new_[46855]_  = A235 & A234;
  assign \new_[46858]_  = A266 & ~A265;
  assign \new_[46859]_  = \new_[46858]_  & \new_[46855]_ ;
  assign \new_[46860]_  = \new_[46859]_  & \new_[46852]_ ;
  assign \new_[46864]_  = A167 & ~A168;
  assign \new_[46865]_  = A169 & \new_[46864]_ ;
  assign \new_[46868]_  = A199 & ~A166;
  assign \new_[46871]_  = A201 & ~A200;
  assign \new_[46872]_  = \new_[46871]_  & \new_[46868]_ ;
  assign \new_[46873]_  = \new_[46872]_  & \new_[46865]_ ;
  assign \new_[46877]_  = ~A233 & A232;
  assign \new_[46878]_  = A202 & \new_[46877]_ ;
  assign \new_[46881]_  = A236 & A234;
  assign \new_[46884]_  = ~A300 & A298;
  assign \new_[46885]_  = \new_[46884]_  & \new_[46881]_ ;
  assign \new_[46886]_  = \new_[46885]_  & \new_[46878]_ ;
  assign \new_[46890]_  = A167 & ~A168;
  assign \new_[46891]_  = A169 & \new_[46890]_ ;
  assign \new_[46894]_  = A199 & ~A166;
  assign \new_[46897]_  = A201 & ~A200;
  assign \new_[46898]_  = \new_[46897]_  & \new_[46894]_ ;
  assign \new_[46899]_  = \new_[46898]_  & \new_[46891]_ ;
  assign \new_[46903]_  = ~A233 & A232;
  assign \new_[46904]_  = A202 & \new_[46903]_ ;
  assign \new_[46907]_  = A236 & A234;
  assign \new_[46910]_  = A299 & A298;
  assign \new_[46911]_  = \new_[46910]_  & \new_[46907]_ ;
  assign \new_[46912]_  = \new_[46911]_  & \new_[46904]_ ;
  assign \new_[46916]_  = A167 & ~A168;
  assign \new_[46917]_  = A169 & \new_[46916]_ ;
  assign \new_[46920]_  = A199 & ~A166;
  assign \new_[46923]_  = A201 & ~A200;
  assign \new_[46924]_  = \new_[46923]_  & \new_[46920]_ ;
  assign \new_[46925]_  = \new_[46924]_  & \new_[46917]_ ;
  assign \new_[46929]_  = ~A233 & A232;
  assign \new_[46930]_  = A202 & \new_[46929]_ ;
  assign \new_[46933]_  = A236 & A234;
  assign \new_[46936]_  = ~A299 & ~A298;
  assign \new_[46937]_  = \new_[46936]_  & \new_[46933]_ ;
  assign \new_[46938]_  = \new_[46937]_  & \new_[46930]_ ;
  assign \new_[46942]_  = A167 & ~A168;
  assign \new_[46943]_  = A169 & \new_[46942]_ ;
  assign \new_[46946]_  = A199 & ~A166;
  assign \new_[46949]_  = A201 & ~A200;
  assign \new_[46950]_  = \new_[46949]_  & \new_[46946]_ ;
  assign \new_[46951]_  = \new_[46950]_  & \new_[46943]_ ;
  assign \new_[46955]_  = ~A233 & A232;
  assign \new_[46956]_  = A202 & \new_[46955]_ ;
  assign \new_[46959]_  = A236 & A234;
  assign \new_[46962]_  = A266 & ~A265;
  assign \new_[46963]_  = \new_[46962]_  & \new_[46959]_ ;
  assign \new_[46964]_  = \new_[46963]_  & \new_[46956]_ ;
  assign \new_[46968]_  = A167 & ~A168;
  assign \new_[46969]_  = A169 & \new_[46968]_ ;
  assign \new_[46972]_  = A199 & ~A166;
  assign \new_[46975]_  = A201 & ~A200;
  assign \new_[46976]_  = \new_[46975]_  & \new_[46972]_ ;
  assign \new_[46977]_  = \new_[46976]_  & \new_[46969]_ ;
  assign \new_[46981]_  = ~A233 & ~A232;
  assign \new_[46982]_  = A202 & \new_[46981]_ ;
  assign \new_[46985]_  = A266 & A265;
  assign \new_[46988]_  = A299 & ~A298;
  assign \new_[46989]_  = \new_[46988]_  & \new_[46985]_ ;
  assign \new_[46990]_  = \new_[46989]_  & \new_[46982]_ ;
  assign \new_[46994]_  = A167 & ~A168;
  assign \new_[46995]_  = A169 & \new_[46994]_ ;
  assign \new_[46998]_  = A199 & ~A166;
  assign \new_[47001]_  = A201 & ~A200;
  assign \new_[47002]_  = \new_[47001]_  & \new_[46998]_ ;
  assign \new_[47003]_  = \new_[47002]_  & \new_[46995]_ ;
  assign \new_[47007]_  = ~A233 & ~A232;
  assign \new_[47008]_  = A202 & \new_[47007]_ ;
  assign \new_[47011]_  = ~A267 & ~A266;
  assign \new_[47014]_  = A299 & ~A298;
  assign \new_[47015]_  = \new_[47014]_  & \new_[47011]_ ;
  assign \new_[47016]_  = \new_[47015]_  & \new_[47008]_ ;
  assign \new_[47020]_  = A167 & ~A168;
  assign \new_[47021]_  = A169 & \new_[47020]_ ;
  assign \new_[47024]_  = A199 & ~A166;
  assign \new_[47027]_  = A201 & ~A200;
  assign \new_[47028]_  = \new_[47027]_  & \new_[47024]_ ;
  assign \new_[47029]_  = \new_[47028]_  & \new_[47021]_ ;
  assign \new_[47033]_  = ~A233 & ~A232;
  assign \new_[47034]_  = A202 & \new_[47033]_ ;
  assign \new_[47037]_  = ~A266 & ~A265;
  assign \new_[47040]_  = A299 & ~A298;
  assign \new_[47041]_  = \new_[47040]_  & \new_[47037]_ ;
  assign \new_[47042]_  = \new_[47041]_  & \new_[47034]_ ;
  assign \new_[47046]_  = A167 & ~A168;
  assign \new_[47047]_  = A169 & \new_[47046]_ ;
  assign \new_[47050]_  = A199 & ~A166;
  assign \new_[47053]_  = A201 & ~A200;
  assign \new_[47054]_  = \new_[47053]_  & \new_[47050]_ ;
  assign \new_[47055]_  = \new_[47054]_  & \new_[47047]_ ;
  assign \new_[47059]_  = A233 & A232;
  assign \new_[47060]_  = A203 & \new_[47059]_ ;
  assign \new_[47063]_  = ~A267 & A265;
  assign \new_[47066]_  = A299 & ~A298;
  assign \new_[47067]_  = \new_[47066]_  & \new_[47063]_ ;
  assign \new_[47068]_  = \new_[47067]_  & \new_[47060]_ ;
  assign \new_[47072]_  = A167 & ~A168;
  assign \new_[47073]_  = A169 & \new_[47072]_ ;
  assign \new_[47076]_  = A199 & ~A166;
  assign \new_[47079]_  = A201 & ~A200;
  assign \new_[47080]_  = \new_[47079]_  & \new_[47076]_ ;
  assign \new_[47081]_  = \new_[47080]_  & \new_[47073]_ ;
  assign \new_[47085]_  = A233 & A232;
  assign \new_[47086]_  = A203 & \new_[47085]_ ;
  assign \new_[47089]_  = A266 & A265;
  assign \new_[47092]_  = A299 & ~A298;
  assign \new_[47093]_  = \new_[47092]_  & \new_[47089]_ ;
  assign \new_[47094]_  = \new_[47093]_  & \new_[47086]_ ;
  assign \new_[47098]_  = A167 & ~A168;
  assign \new_[47099]_  = A169 & \new_[47098]_ ;
  assign \new_[47102]_  = A199 & ~A166;
  assign \new_[47105]_  = A201 & ~A200;
  assign \new_[47106]_  = \new_[47105]_  & \new_[47102]_ ;
  assign \new_[47107]_  = \new_[47106]_  & \new_[47099]_ ;
  assign \new_[47111]_  = A233 & A232;
  assign \new_[47112]_  = A203 & \new_[47111]_ ;
  assign \new_[47115]_  = ~A266 & ~A265;
  assign \new_[47118]_  = A299 & ~A298;
  assign \new_[47119]_  = \new_[47118]_  & \new_[47115]_ ;
  assign \new_[47120]_  = \new_[47119]_  & \new_[47112]_ ;
  assign \new_[47124]_  = A167 & ~A168;
  assign \new_[47125]_  = A169 & \new_[47124]_ ;
  assign \new_[47128]_  = A199 & ~A166;
  assign \new_[47131]_  = A201 & ~A200;
  assign \new_[47132]_  = \new_[47131]_  & \new_[47128]_ ;
  assign \new_[47133]_  = \new_[47132]_  & \new_[47125]_ ;
  assign \new_[47137]_  = A233 & ~A232;
  assign \new_[47138]_  = A203 & \new_[47137]_ ;
  assign \new_[47141]_  = ~A266 & A265;
  assign \new_[47144]_  = A268 & A267;
  assign \new_[47145]_  = \new_[47144]_  & \new_[47141]_ ;
  assign \new_[47146]_  = \new_[47145]_  & \new_[47138]_ ;
  assign \new_[47150]_  = A167 & ~A168;
  assign \new_[47151]_  = A169 & \new_[47150]_ ;
  assign \new_[47154]_  = A199 & ~A166;
  assign \new_[47157]_  = A201 & ~A200;
  assign \new_[47158]_  = \new_[47157]_  & \new_[47154]_ ;
  assign \new_[47159]_  = \new_[47158]_  & \new_[47151]_ ;
  assign \new_[47163]_  = A233 & ~A232;
  assign \new_[47164]_  = A203 & \new_[47163]_ ;
  assign \new_[47167]_  = ~A266 & A265;
  assign \new_[47170]_  = A269 & A267;
  assign \new_[47171]_  = \new_[47170]_  & \new_[47167]_ ;
  assign \new_[47172]_  = \new_[47171]_  & \new_[47164]_ ;
  assign \new_[47176]_  = A167 & ~A168;
  assign \new_[47177]_  = A169 & \new_[47176]_ ;
  assign \new_[47180]_  = A199 & ~A166;
  assign \new_[47183]_  = A201 & ~A200;
  assign \new_[47184]_  = \new_[47183]_  & \new_[47180]_ ;
  assign \new_[47185]_  = \new_[47184]_  & \new_[47177]_ ;
  assign \new_[47189]_  = ~A234 & ~A233;
  assign \new_[47190]_  = A203 & \new_[47189]_ ;
  assign \new_[47193]_  = A266 & A265;
  assign \new_[47196]_  = A299 & ~A298;
  assign \new_[47197]_  = \new_[47196]_  & \new_[47193]_ ;
  assign \new_[47198]_  = \new_[47197]_  & \new_[47190]_ ;
  assign \new_[47202]_  = A167 & ~A168;
  assign \new_[47203]_  = A169 & \new_[47202]_ ;
  assign \new_[47206]_  = A199 & ~A166;
  assign \new_[47209]_  = A201 & ~A200;
  assign \new_[47210]_  = \new_[47209]_  & \new_[47206]_ ;
  assign \new_[47211]_  = \new_[47210]_  & \new_[47203]_ ;
  assign \new_[47215]_  = ~A234 & ~A233;
  assign \new_[47216]_  = A203 & \new_[47215]_ ;
  assign \new_[47219]_  = ~A267 & ~A266;
  assign \new_[47222]_  = A299 & ~A298;
  assign \new_[47223]_  = \new_[47222]_  & \new_[47219]_ ;
  assign \new_[47224]_  = \new_[47223]_  & \new_[47216]_ ;
  assign \new_[47228]_  = A167 & ~A168;
  assign \new_[47229]_  = A169 & \new_[47228]_ ;
  assign \new_[47232]_  = A199 & ~A166;
  assign \new_[47235]_  = A201 & ~A200;
  assign \new_[47236]_  = \new_[47235]_  & \new_[47232]_ ;
  assign \new_[47237]_  = \new_[47236]_  & \new_[47229]_ ;
  assign \new_[47241]_  = ~A234 & ~A233;
  assign \new_[47242]_  = A203 & \new_[47241]_ ;
  assign \new_[47245]_  = ~A266 & ~A265;
  assign \new_[47248]_  = A299 & ~A298;
  assign \new_[47249]_  = \new_[47248]_  & \new_[47245]_ ;
  assign \new_[47250]_  = \new_[47249]_  & \new_[47242]_ ;
  assign \new_[47254]_  = A167 & ~A168;
  assign \new_[47255]_  = A169 & \new_[47254]_ ;
  assign \new_[47258]_  = A199 & ~A166;
  assign \new_[47261]_  = A201 & ~A200;
  assign \new_[47262]_  = \new_[47261]_  & \new_[47258]_ ;
  assign \new_[47263]_  = \new_[47262]_  & \new_[47255]_ ;
  assign \new_[47267]_  = ~A233 & A232;
  assign \new_[47268]_  = A203 & \new_[47267]_ ;
  assign \new_[47271]_  = A235 & A234;
  assign \new_[47274]_  = ~A300 & A298;
  assign \new_[47275]_  = \new_[47274]_  & \new_[47271]_ ;
  assign \new_[47276]_  = \new_[47275]_  & \new_[47268]_ ;
  assign \new_[47280]_  = A167 & ~A168;
  assign \new_[47281]_  = A169 & \new_[47280]_ ;
  assign \new_[47284]_  = A199 & ~A166;
  assign \new_[47287]_  = A201 & ~A200;
  assign \new_[47288]_  = \new_[47287]_  & \new_[47284]_ ;
  assign \new_[47289]_  = \new_[47288]_  & \new_[47281]_ ;
  assign \new_[47293]_  = ~A233 & A232;
  assign \new_[47294]_  = A203 & \new_[47293]_ ;
  assign \new_[47297]_  = A235 & A234;
  assign \new_[47300]_  = A299 & A298;
  assign \new_[47301]_  = \new_[47300]_  & \new_[47297]_ ;
  assign \new_[47302]_  = \new_[47301]_  & \new_[47294]_ ;
  assign \new_[47306]_  = A167 & ~A168;
  assign \new_[47307]_  = A169 & \new_[47306]_ ;
  assign \new_[47310]_  = A199 & ~A166;
  assign \new_[47313]_  = A201 & ~A200;
  assign \new_[47314]_  = \new_[47313]_  & \new_[47310]_ ;
  assign \new_[47315]_  = \new_[47314]_  & \new_[47307]_ ;
  assign \new_[47319]_  = ~A233 & A232;
  assign \new_[47320]_  = A203 & \new_[47319]_ ;
  assign \new_[47323]_  = A235 & A234;
  assign \new_[47326]_  = ~A299 & ~A298;
  assign \new_[47327]_  = \new_[47326]_  & \new_[47323]_ ;
  assign \new_[47328]_  = \new_[47327]_  & \new_[47320]_ ;
  assign \new_[47332]_  = A167 & ~A168;
  assign \new_[47333]_  = A169 & \new_[47332]_ ;
  assign \new_[47336]_  = A199 & ~A166;
  assign \new_[47339]_  = A201 & ~A200;
  assign \new_[47340]_  = \new_[47339]_  & \new_[47336]_ ;
  assign \new_[47341]_  = \new_[47340]_  & \new_[47333]_ ;
  assign \new_[47345]_  = ~A233 & A232;
  assign \new_[47346]_  = A203 & \new_[47345]_ ;
  assign \new_[47349]_  = A235 & A234;
  assign \new_[47352]_  = A266 & ~A265;
  assign \new_[47353]_  = \new_[47352]_  & \new_[47349]_ ;
  assign \new_[47354]_  = \new_[47353]_  & \new_[47346]_ ;
  assign \new_[47358]_  = A167 & ~A168;
  assign \new_[47359]_  = A169 & \new_[47358]_ ;
  assign \new_[47362]_  = A199 & ~A166;
  assign \new_[47365]_  = A201 & ~A200;
  assign \new_[47366]_  = \new_[47365]_  & \new_[47362]_ ;
  assign \new_[47367]_  = \new_[47366]_  & \new_[47359]_ ;
  assign \new_[47371]_  = ~A233 & A232;
  assign \new_[47372]_  = A203 & \new_[47371]_ ;
  assign \new_[47375]_  = A236 & A234;
  assign \new_[47378]_  = ~A300 & A298;
  assign \new_[47379]_  = \new_[47378]_  & \new_[47375]_ ;
  assign \new_[47380]_  = \new_[47379]_  & \new_[47372]_ ;
  assign \new_[47384]_  = A167 & ~A168;
  assign \new_[47385]_  = A169 & \new_[47384]_ ;
  assign \new_[47388]_  = A199 & ~A166;
  assign \new_[47391]_  = A201 & ~A200;
  assign \new_[47392]_  = \new_[47391]_  & \new_[47388]_ ;
  assign \new_[47393]_  = \new_[47392]_  & \new_[47385]_ ;
  assign \new_[47397]_  = ~A233 & A232;
  assign \new_[47398]_  = A203 & \new_[47397]_ ;
  assign \new_[47401]_  = A236 & A234;
  assign \new_[47404]_  = A299 & A298;
  assign \new_[47405]_  = \new_[47404]_  & \new_[47401]_ ;
  assign \new_[47406]_  = \new_[47405]_  & \new_[47398]_ ;
  assign \new_[47410]_  = A167 & ~A168;
  assign \new_[47411]_  = A169 & \new_[47410]_ ;
  assign \new_[47414]_  = A199 & ~A166;
  assign \new_[47417]_  = A201 & ~A200;
  assign \new_[47418]_  = \new_[47417]_  & \new_[47414]_ ;
  assign \new_[47419]_  = \new_[47418]_  & \new_[47411]_ ;
  assign \new_[47423]_  = ~A233 & A232;
  assign \new_[47424]_  = A203 & \new_[47423]_ ;
  assign \new_[47427]_  = A236 & A234;
  assign \new_[47430]_  = ~A299 & ~A298;
  assign \new_[47431]_  = \new_[47430]_  & \new_[47427]_ ;
  assign \new_[47432]_  = \new_[47431]_  & \new_[47424]_ ;
  assign \new_[47436]_  = A167 & ~A168;
  assign \new_[47437]_  = A169 & \new_[47436]_ ;
  assign \new_[47440]_  = A199 & ~A166;
  assign \new_[47443]_  = A201 & ~A200;
  assign \new_[47444]_  = \new_[47443]_  & \new_[47440]_ ;
  assign \new_[47445]_  = \new_[47444]_  & \new_[47437]_ ;
  assign \new_[47449]_  = ~A233 & A232;
  assign \new_[47450]_  = A203 & \new_[47449]_ ;
  assign \new_[47453]_  = A236 & A234;
  assign \new_[47456]_  = A266 & ~A265;
  assign \new_[47457]_  = \new_[47456]_  & \new_[47453]_ ;
  assign \new_[47458]_  = \new_[47457]_  & \new_[47450]_ ;
  assign \new_[47462]_  = A167 & ~A168;
  assign \new_[47463]_  = A169 & \new_[47462]_ ;
  assign \new_[47466]_  = A199 & ~A166;
  assign \new_[47469]_  = A201 & ~A200;
  assign \new_[47470]_  = \new_[47469]_  & \new_[47466]_ ;
  assign \new_[47471]_  = \new_[47470]_  & \new_[47463]_ ;
  assign \new_[47475]_  = ~A233 & ~A232;
  assign \new_[47476]_  = A203 & \new_[47475]_ ;
  assign \new_[47479]_  = A266 & A265;
  assign \new_[47482]_  = A299 & ~A298;
  assign \new_[47483]_  = \new_[47482]_  & \new_[47479]_ ;
  assign \new_[47484]_  = \new_[47483]_  & \new_[47476]_ ;
  assign \new_[47488]_  = A167 & ~A168;
  assign \new_[47489]_  = A169 & \new_[47488]_ ;
  assign \new_[47492]_  = A199 & ~A166;
  assign \new_[47495]_  = A201 & ~A200;
  assign \new_[47496]_  = \new_[47495]_  & \new_[47492]_ ;
  assign \new_[47497]_  = \new_[47496]_  & \new_[47489]_ ;
  assign \new_[47501]_  = ~A233 & ~A232;
  assign \new_[47502]_  = A203 & \new_[47501]_ ;
  assign \new_[47505]_  = ~A267 & ~A266;
  assign \new_[47508]_  = A299 & ~A298;
  assign \new_[47509]_  = \new_[47508]_  & \new_[47505]_ ;
  assign \new_[47510]_  = \new_[47509]_  & \new_[47502]_ ;
  assign \new_[47514]_  = A167 & ~A168;
  assign \new_[47515]_  = A169 & \new_[47514]_ ;
  assign \new_[47518]_  = A199 & ~A166;
  assign \new_[47521]_  = A201 & ~A200;
  assign \new_[47522]_  = \new_[47521]_  & \new_[47518]_ ;
  assign \new_[47523]_  = \new_[47522]_  & \new_[47515]_ ;
  assign \new_[47527]_  = ~A233 & ~A232;
  assign \new_[47528]_  = A203 & \new_[47527]_ ;
  assign \new_[47531]_  = ~A266 & ~A265;
  assign \new_[47534]_  = A299 & ~A298;
  assign \new_[47535]_  = \new_[47534]_  & \new_[47531]_ ;
  assign \new_[47536]_  = \new_[47535]_  & \new_[47528]_ ;
  assign \new_[47540]_  = ~A167 & ~A168;
  assign \new_[47541]_  = A169 & \new_[47540]_ ;
  assign \new_[47544]_  = ~A199 & A166;
  assign \new_[47547]_  = A232 & A200;
  assign \new_[47548]_  = \new_[47547]_  & \new_[47544]_ ;
  assign \new_[47549]_  = \new_[47548]_  & \new_[47541]_ ;
  assign \new_[47553]_  = ~A267 & A265;
  assign \new_[47554]_  = A233 & \new_[47553]_ ;
  assign \new_[47557]_  = ~A299 & A298;
  assign \new_[47560]_  = A301 & A300;
  assign \new_[47561]_  = \new_[47560]_  & \new_[47557]_ ;
  assign \new_[47562]_  = \new_[47561]_  & \new_[47554]_ ;
  assign \new_[47566]_  = ~A167 & ~A168;
  assign \new_[47567]_  = A169 & \new_[47566]_ ;
  assign \new_[47570]_  = ~A199 & A166;
  assign \new_[47573]_  = A232 & A200;
  assign \new_[47574]_  = \new_[47573]_  & \new_[47570]_ ;
  assign \new_[47575]_  = \new_[47574]_  & \new_[47567]_ ;
  assign \new_[47579]_  = ~A267 & A265;
  assign \new_[47580]_  = A233 & \new_[47579]_ ;
  assign \new_[47583]_  = ~A299 & A298;
  assign \new_[47586]_  = A302 & A300;
  assign \new_[47587]_  = \new_[47586]_  & \new_[47583]_ ;
  assign \new_[47588]_  = \new_[47587]_  & \new_[47580]_ ;
  assign \new_[47592]_  = ~A167 & ~A168;
  assign \new_[47593]_  = A169 & \new_[47592]_ ;
  assign \new_[47596]_  = ~A199 & A166;
  assign \new_[47599]_  = A232 & A200;
  assign \new_[47600]_  = \new_[47599]_  & \new_[47596]_ ;
  assign \new_[47601]_  = \new_[47600]_  & \new_[47593]_ ;
  assign \new_[47605]_  = A266 & A265;
  assign \new_[47606]_  = A233 & \new_[47605]_ ;
  assign \new_[47609]_  = ~A299 & A298;
  assign \new_[47612]_  = A301 & A300;
  assign \new_[47613]_  = \new_[47612]_  & \new_[47609]_ ;
  assign \new_[47614]_  = \new_[47613]_  & \new_[47606]_ ;
  assign \new_[47618]_  = ~A167 & ~A168;
  assign \new_[47619]_  = A169 & \new_[47618]_ ;
  assign \new_[47622]_  = ~A199 & A166;
  assign \new_[47625]_  = A232 & A200;
  assign \new_[47626]_  = \new_[47625]_  & \new_[47622]_ ;
  assign \new_[47627]_  = \new_[47626]_  & \new_[47619]_ ;
  assign \new_[47631]_  = A266 & A265;
  assign \new_[47632]_  = A233 & \new_[47631]_ ;
  assign \new_[47635]_  = ~A299 & A298;
  assign \new_[47638]_  = A302 & A300;
  assign \new_[47639]_  = \new_[47638]_  & \new_[47635]_ ;
  assign \new_[47640]_  = \new_[47639]_  & \new_[47632]_ ;
  assign \new_[47644]_  = ~A167 & ~A168;
  assign \new_[47645]_  = A169 & \new_[47644]_ ;
  assign \new_[47648]_  = ~A199 & A166;
  assign \new_[47651]_  = A232 & A200;
  assign \new_[47652]_  = \new_[47651]_  & \new_[47648]_ ;
  assign \new_[47653]_  = \new_[47652]_  & \new_[47645]_ ;
  assign \new_[47657]_  = ~A266 & ~A265;
  assign \new_[47658]_  = A233 & \new_[47657]_ ;
  assign \new_[47661]_  = ~A299 & A298;
  assign \new_[47664]_  = A301 & A300;
  assign \new_[47665]_  = \new_[47664]_  & \new_[47661]_ ;
  assign \new_[47666]_  = \new_[47665]_  & \new_[47658]_ ;
  assign \new_[47670]_  = ~A167 & ~A168;
  assign \new_[47671]_  = A169 & \new_[47670]_ ;
  assign \new_[47674]_  = ~A199 & A166;
  assign \new_[47677]_  = A232 & A200;
  assign \new_[47678]_  = \new_[47677]_  & \new_[47674]_ ;
  assign \new_[47679]_  = \new_[47678]_  & \new_[47671]_ ;
  assign \new_[47683]_  = ~A266 & ~A265;
  assign \new_[47684]_  = A233 & \new_[47683]_ ;
  assign \new_[47687]_  = ~A299 & A298;
  assign \new_[47690]_  = A302 & A300;
  assign \new_[47691]_  = \new_[47690]_  & \new_[47687]_ ;
  assign \new_[47692]_  = \new_[47691]_  & \new_[47684]_ ;
  assign \new_[47696]_  = ~A167 & ~A168;
  assign \new_[47697]_  = A169 & \new_[47696]_ ;
  assign \new_[47700]_  = ~A199 & A166;
  assign \new_[47703]_  = ~A233 & A200;
  assign \new_[47704]_  = \new_[47703]_  & \new_[47700]_ ;
  assign \new_[47705]_  = \new_[47704]_  & \new_[47697]_ ;
  assign \new_[47709]_  = ~A266 & ~A236;
  assign \new_[47710]_  = ~A235 & \new_[47709]_ ;
  assign \new_[47713]_  = ~A269 & ~A268;
  assign \new_[47716]_  = A299 & ~A298;
  assign \new_[47717]_  = \new_[47716]_  & \new_[47713]_ ;
  assign \new_[47718]_  = \new_[47717]_  & \new_[47710]_ ;
  assign \new_[47722]_  = ~A167 & ~A168;
  assign \new_[47723]_  = A169 & \new_[47722]_ ;
  assign \new_[47726]_  = ~A199 & A166;
  assign \new_[47729]_  = ~A233 & A200;
  assign \new_[47730]_  = \new_[47729]_  & \new_[47726]_ ;
  assign \new_[47731]_  = \new_[47730]_  & \new_[47723]_ ;
  assign \new_[47735]_  = A266 & A265;
  assign \new_[47736]_  = ~A234 & \new_[47735]_ ;
  assign \new_[47739]_  = ~A299 & A298;
  assign \new_[47742]_  = A301 & A300;
  assign \new_[47743]_  = \new_[47742]_  & \new_[47739]_ ;
  assign \new_[47744]_  = \new_[47743]_  & \new_[47736]_ ;
  assign \new_[47748]_  = ~A167 & ~A168;
  assign \new_[47749]_  = A169 & \new_[47748]_ ;
  assign \new_[47752]_  = ~A199 & A166;
  assign \new_[47755]_  = ~A233 & A200;
  assign \new_[47756]_  = \new_[47755]_  & \new_[47752]_ ;
  assign \new_[47757]_  = \new_[47756]_  & \new_[47749]_ ;
  assign \new_[47761]_  = A266 & A265;
  assign \new_[47762]_  = ~A234 & \new_[47761]_ ;
  assign \new_[47765]_  = ~A299 & A298;
  assign \new_[47768]_  = A302 & A300;
  assign \new_[47769]_  = \new_[47768]_  & \new_[47765]_ ;
  assign \new_[47770]_  = \new_[47769]_  & \new_[47762]_ ;
  assign \new_[47774]_  = ~A167 & ~A168;
  assign \new_[47775]_  = A169 & \new_[47774]_ ;
  assign \new_[47778]_  = ~A199 & A166;
  assign \new_[47781]_  = ~A233 & A200;
  assign \new_[47782]_  = \new_[47781]_  & \new_[47778]_ ;
  assign \new_[47783]_  = \new_[47782]_  & \new_[47775]_ ;
  assign \new_[47787]_  = ~A267 & ~A266;
  assign \new_[47788]_  = ~A234 & \new_[47787]_ ;
  assign \new_[47791]_  = ~A299 & A298;
  assign \new_[47794]_  = A301 & A300;
  assign \new_[47795]_  = \new_[47794]_  & \new_[47791]_ ;
  assign \new_[47796]_  = \new_[47795]_  & \new_[47788]_ ;
  assign \new_[47800]_  = ~A167 & ~A168;
  assign \new_[47801]_  = A169 & \new_[47800]_ ;
  assign \new_[47804]_  = ~A199 & A166;
  assign \new_[47807]_  = ~A233 & A200;
  assign \new_[47808]_  = \new_[47807]_  & \new_[47804]_ ;
  assign \new_[47809]_  = \new_[47808]_  & \new_[47801]_ ;
  assign \new_[47813]_  = ~A267 & ~A266;
  assign \new_[47814]_  = ~A234 & \new_[47813]_ ;
  assign \new_[47817]_  = ~A299 & A298;
  assign \new_[47820]_  = A302 & A300;
  assign \new_[47821]_  = \new_[47820]_  & \new_[47817]_ ;
  assign \new_[47822]_  = \new_[47821]_  & \new_[47814]_ ;
  assign \new_[47826]_  = ~A167 & ~A168;
  assign \new_[47827]_  = A169 & \new_[47826]_ ;
  assign \new_[47830]_  = ~A199 & A166;
  assign \new_[47833]_  = ~A233 & A200;
  assign \new_[47834]_  = \new_[47833]_  & \new_[47830]_ ;
  assign \new_[47835]_  = \new_[47834]_  & \new_[47827]_ ;
  assign \new_[47839]_  = ~A266 & ~A265;
  assign \new_[47840]_  = ~A234 & \new_[47839]_ ;
  assign \new_[47843]_  = ~A299 & A298;
  assign \new_[47846]_  = A301 & A300;
  assign \new_[47847]_  = \new_[47846]_  & \new_[47843]_ ;
  assign \new_[47848]_  = \new_[47847]_  & \new_[47840]_ ;
  assign \new_[47852]_  = ~A167 & ~A168;
  assign \new_[47853]_  = A169 & \new_[47852]_ ;
  assign \new_[47856]_  = ~A199 & A166;
  assign \new_[47859]_  = ~A233 & A200;
  assign \new_[47860]_  = \new_[47859]_  & \new_[47856]_ ;
  assign \new_[47861]_  = \new_[47860]_  & \new_[47853]_ ;
  assign \new_[47865]_  = ~A266 & ~A265;
  assign \new_[47866]_  = ~A234 & \new_[47865]_ ;
  assign \new_[47869]_  = ~A299 & A298;
  assign \new_[47872]_  = A302 & A300;
  assign \new_[47873]_  = \new_[47872]_  & \new_[47869]_ ;
  assign \new_[47874]_  = \new_[47873]_  & \new_[47866]_ ;
  assign \new_[47878]_  = ~A167 & ~A168;
  assign \new_[47879]_  = A169 & \new_[47878]_ ;
  assign \new_[47882]_  = ~A199 & A166;
  assign \new_[47885]_  = A232 & A200;
  assign \new_[47886]_  = \new_[47885]_  & \new_[47882]_ ;
  assign \new_[47887]_  = \new_[47886]_  & \new_[47879]_ ;
  assign \new_[47891]_  = A235 & A234;
  assign \new_[47892]_  = ~A233 & \new_[47891]_ ;
  assign \new_[47895]_  = ~A266 & A265;
  assign \new_[47898]_  = A268 & A267;
  assign \new_[47899]_  = \new_[47898]_  & \new_[47895]_ ;
  assign \new_[47900]_  = \new_[47899]_  & \new_[47892]_ ;
  assign \new_[47904]_  = ~A167 & ~A168;
  assign \new_[47905]_  = A169 & \new_[47904]_ ;
  assign \new_[47908]_  = ~A199 & A166;
  assign \new_[47911]_  = A232 & A200;
  assign \new_[47912]_  = \new_[47911]_  & \new_[47908]_ ;
  assign \new_[47913]_  = \new_[47912]_  & \new_[47905]_ ;
  assign \new_[47917]_  = A235 & A234;
  assign \new_[47918]_  = ~A233 & \new_[47917]_ ;
  assign \new_[47921]_  = ~A266 & A265;
  assign \new_[47924]_  = A269 & A267;
  assign \new_[47925]_  = \new_[47924]_  & \new_[47921]_ ;
  assign \new_[47926]_  = \new_[47925]_  & \new_[47918]_ ;
  assign \new_[47930]_  = ~A167 & ~A168;
  assign \new_[47931]_  = A169 & \new_[47930]_ ;
  assign \new_[47934]_  = ~A199 & A166;
  assign \new_[47937]_  = A232 & A200;
  assign \new_[47938]_  = \new_[47937]_  & \new_[47934]_ ;
  assign \new_[47939]_  = \new_[47938]_  & \new_[47931]_ ;
  assign \new_[47943]_  = A236 & A234;
  assign \new_[47944]_  = ~A233 & \new_[47943]_ ;
  assign \new_[47947]_  = ~A266 & A265;
  assign \new_[47950]_  = A268 & A267;
  assign \new_[47951]_  = \new_[47950]_  & \new_[47947]_ ;
  assign \new_[47952]_  = \new_[47951]_  & \new_[47944]_ ;
  assign \new_[47956]_  = ~A167 & ~A168;
  assign \new_[47957]_  = A169 & \new_[47956]_ ;
  assign \new_[47960]_  = ~A199 & A166;
  assign \new_[47963]_  = A232 & A200;
  assign \new_[47964]_  = \new_[47963]_  & \new_[47960]_ ;
  assign \new_[47965]_  = \new_[47964]_  & \new_[47957]_ ;
  assign \new_[47969]_  = A236 & A234;
  assign \new_[47970]_  = ~A233 & \new_[47969]_ ;
  assign \new_[47973]_  = ~A266 & A265;
  assign \new_[47976]_  = A269 & A267;
  assign \new_[47977]_  = \new_[47976]_  & \new_[47973]_ ;
  assign \new_[47978]_  = \new_[47977]_  & \new_[47970]_ ;
  assign \new_[47982]_  = ~A167 & ~A168;
  assign \new_[47983]_  = A169 & \new_[47982]_ ;
  assign \new_[47986]_  = ~A199 & A166;
  assign \new_[47989]_  = ~A232 & A200;
  assign \new_[47990]_  = \new_[47989]_  & \new_[47986]_ ;
  assign \new_[47991]_  = \new_[47990]_  & \new_[47983]_ ;
  assign \new_[47995]_  = A266 & A265;
  assign \new_[47996]_  = ~A233 & \new_[47995]_ ;
  assign \new_[47999]_  = ~A299 & A298;
  assign \new_[48002]_  = A301 & A300;
  assign \new_[48003]_  = \new_[48002]_  & \new_[47999]_ ;
  assign \new_[48004]_  = \new_[48003]_  & \new_[47996]_ ;
  assign \new_[48008]_  = ~A167 & ~A168;
  assign \new_[48009]_  = A169 & \new_[48008]_ ;
  assign \new_[48012]_  = ~A199 & A166;
  assign \new_[48015]_  = ~A232 & A200;
  assign \new_[48016]_  = \new_[48015]_  & \new_[48012]_ ;
  assign \new_[48017]_  = \new_[48016]_  & \new_[48009]_ ;
  assign \new_[48021]_  = A266 & A265;
  assign \new_[48022]_  = ~A233 & \new_[48021]_ ;
  assign \new_[48025]_  = ~A299 & A298;
  assign \new_[48028]_  = A302 & A300;
  assign \new_[48029]_  = \new_[48028]_  & \new_[48025]_ ;
  assign \new_[48030]_  = \new_[48029]_  & \new_[48022]_ ;
  assign \new_[48034]_  = ~A167 & ~A168;
  assign \new_[48035]_  = A169 & \new_[48034]_ ;
  assign \new_[48038]_  = ~A199 & A166;
  assign \new_[48041]_  = ~A232 & A200;
  assign \new_[48042]_  = \new_[48041]_  & \new_[48038]_ ;
  assign \new_[48043]_  = \new_[48042]_  & \new_[48035]_ ;
  assign \new_[48047]_  = ~A267 & ~A266;
  assign \new_[48048]_  = ~A233 & \new_[48047]_ ;
  assign \new_[48051]_  = ~A299 & A298;
  assign \new_[48054]_  = A301 & A300;
  assign \new_[48055]_  = \new_[48054]_  & \new_[48051]_ ;
  assign \new_[48056]_  = \new_[48055]_  & \new_[48048]_ ;
  assign \new_[48060]_  = ~A167 & ~A168;
  assign \new_[48061]_  = A169 & \new_[48060]_ ;
  assign \new_[48064]_  = ~A199 & A166;
  assign \new_[48067]_  = ~A232 & A200;
  assign \new_[48068]_  = \new_[48067]_  & \new_[48064]_ ;
  assign \new_[48069]_  = \new_[48068]_  & \new_[48061]_ ;
  assign \new_[48073]_  = ~A267 & ~A266;
  assign \new_[48074]_  = ~A233 & \new_[48073]_ ;
  assign \new_[48077]_  = ~A299 & A298;
  assign \new_[48080]_  = A302 & A300;
  assign \new_[48081]_  = \new_[48080]_  & \new_[48077]_ ;
  assign \new_[48082]_  = \new_[48081]_  & \new_[48074]_ ;
  assign \new_[48086]_  = ~A167 & ~A168;
  assign \new_[48087]_  = A169 & \new_[48086]_ ;
  assign \new_[48090]_  = ~A199 & A166;
  assign \new_[48093]_  = ~A232 & A200;
  assign \new_[48094]_  = \new_[48093]_  & \new_[48090]_ ;
  assign \new_[48095]_  = \new_[48094]_  & \new_[48087]_ ;
  assign \new_[48099]_  = ~A266 & ~A265;
  assign \new_[48100]_  = ~A233 & \new_[48099]_ ;
  assign \new_[48103]_  = ~A299 & A298;
  assign \new_[48106]_  = A301 & A300;
  assign \new_[48107]_  = \new_[48106]_  & \new_[48103]_ ;
  assign \new_[48108]_  = \new_[48107]_  & \new_[48100]_ ;
  assign \new_[48112]_  = ~A167 & ~A168;
  assign \new_[48113]_  = A169 & \new_[48112]_ ;
  assign \new_[48116]_  = ~A199 & A166;
  assign \new_[48119]_  = ~A232 & A200;
  assign \new_[48120]_  = \new_[48119]_  & \new_[48116]_ ;
  assign \new_[48121]_  = \new_[48120]_  & \new_[48113]_ ;
  assign \new_[48125]_  = ~A266 & ~A265;
  assign \new_[48126]_  = ~A233 & \new_[48125]_ ;
  assign \new_[48129]_  = ~A299 & A298;
  assign \new_[48132]_  = A302 & A300;
  assign \new_[48133]_  = \new_[48132]_  & \new_[48129]_ ;
  assign \new_[48134]_  = \new_[48133]_  & \new_[48126]_ ;
  assign \new_[48138]_  = ~A167 & ~A168;
  assign \new_[48139]_  = A169 & \new_[48138]_ ;
  assign \new_[48142]_  = A199 & A166;
  assign \new_[48145]_  = A201 & ~A200;
  assign \new_[48146]_  = \new_[48145]_  & \new_[48142]_ ;
  assign \new_[48147]_  = \new_[48146]_  & \new_[48139]_ ;
  assign \new_[48151]_  = A233 & A232;
  assign \new_[48152]_  = A202 & \new_[48151]_ ;
  assign \new_[48155]_  = ~A267 & A265;
  assign \new_[48158]_  = A299 & ~A298;
  assign \new_[48159]_  = \new_[48158]_  & \new_[48155]_ ;
  assign \new_[48160]_  = \new_[48159]_  & \new_[48152]_ ;
  assign \new_[48164]_  = ~A167 & ~A168;
  assign \new_[48165]_  = A169 & \new_[48164]_ ;
  assign \new_[48168]_  = A199 & A166;
  assign \new_[48171]_  = A201 & ~A200;
  assign \new_[48172]_  = \new_[48171]_  & \new_[48168]_ ;
  assign \new_[48173]_  = \new_[48172]_  & \new_[48165]_ ;
  assign \new_[48177]_  = A233 & A232;
  assign \new_[48178]_  = A202 & \new_[48177]_ ;
  assign \new_[48181]_  = A266 & A265;
  assign \new_[48184]_  = A299 & ~A298;
  assign \new_[48185]_  = \new_[48184]_  & \new_[48181]_ ;
  assign \new_[48186]_  = \new_[48185]_  & \new_[48178]_ ;
  assign \new_[48190]_  = ~A167 & ~A168;
  assign \new_[48191]_  = A169 & \new_[48190]_ ;
  assign \new_[48194]_  = A199 & A166;
  assign \new_[48197]_  = A201 & ~A200;
  assign \new_[48198]_  = \new_[48197]_  & \new_[48194]_ ;
  assign \new_[48199]_  = \new_[48198]_  & \new_[48191]_ ;
  assign \new_[48203]_  = A233 & A232;
  assign \new_[48204]_  = A202 & \new_[48203]_ ;
  assign \new_[48207]_  = ~A266 & ~A265;
  assign \new_[48210]_  = A299 & ~A298;
  assign \new_[48211]_  = \new_[48210]_  & \new_[48207]_ ;
  assign \new_[48212]_  = \new_[48211]_  & \new_[48204]_ ;
  assign \new_[48216]_  = ~A167 & ~A168;
  assign \new_[48217]_  = A169 & \new_[48216]_ ;
  assign \new_[48220]_  = A199 & A166;
  assign \new_[48223]_  = A201 & ~A200;
  assign \new_[48224]_  = \new_[48223]_  & \new_[48220]_ ;
  assign \new_[48225]_  = \new_[48224]_  & \new_[48217]_ ;
  assign \new_[48229]_  = A233 & ~A232;
  assign \new_[48230]_  = A202 & \new_[48229]_ ;
  assign \new_[48233]_  = ~A266 & A265;
  assign \new_[48236]_  = A268 & A267;
  assign \new_[48237]_  = \new_[48236]_  & \new_[48233]_ ;
  assign \new_[48238]_  = \new_[48237]_  & \new_[48230]_ ;
  assign \new_[48242]_  = ~A167 & ~A168;
  assign \new_[48243]_  = A169 & \new_[48242]_ ;
  assign \new_[48246]_  = A199 & A166;
  assign \new_[48249]_  = A201 & ~A200;
  assign \new_[48250]_  = \new_[48249]_  & \new_[48246]_ ;
  assign \new_[48251]_  = \new_[48250]_  & \new_[48243]_ ;
  assign \new_[48255]_  = A233 & ~A232;
  assign \new_[48256]_  = A202 & \new_[48255]_ ;
  assign \new_[48259]_  = ~A266 & A265;
  assign \new_[48262]_  = A269 & A267;
  assign \new_[48263]_  = \new_[48262]_  & \new_[48259]_ ;
  assign \new_[48264]_  = \new_[48263]_  & \new_[48256]_ ;
  assign \new_[48268]_  = ~A167 & ~A168;
  assign \new_[48269]_  = A169 & \new_[48268]_ ;
  assign \new_[48272]_  = A199 & A166;
  assign \new_[48275]_  = A201 & ~A200;
  assign \new_[48276]_  = \new_[48275]_  & \new_[48272]_ ;
  assign \new_[48277]_  = \new_[48276]_  & \new_[48269]_ ;
  assign \new_[48281]_  = ~A234 & ~A233;
  assign \new_[48282]_  = A202 & \new_[48281]_ ;
  assign \new_[48285]_  = A266 & A265;
  assign \new_[48288]_  = A299 & ~A298;
  assign \new_[48289]_  = \new_[48288]_  & \new_[48285]_ ;
  assign \new_[48290]_  = \new_[48289]_  & \new_[48282]_ ;
  assign \new_[48294]_  = ~A167 & ~A168;
  assign \new_[48295]_  = A169 & \new_[48294]_ ;
  assign \new_[48298]_  = A199 & A166;
  assign \new_[48301]_  = A201 & ~A200;
  assign \new_[48302]_  = \new_[48301]_  & \new_[48298]_ ;
  assign \new_[48303]_  = \new_[48302]_  & \new_[48295]_ ;
  assign \new_[48307]_  = ~A234 & ~A233;
  assign \new_[48308]_  = A202 & \new_[48307]_ ;
  assign \new_[48311]_  = ~A267 & ~A266;
  assign \new_[48314]_  = A299 & ~A298;
  assign \new_[48315]_  = \new_[48314]_  & \new_[48311]_ ;
  assign \new_[48316]_  = \new_[48315]_  & \new_[48308]_ ;
  assign \new_[48320]_  = ~A167 & ~A168;
  assign \new_[48321]_  = A169 & \new_[48320]_ ;
  assign \new_[48324]_  = A199 & A166;
  assign \new_[48327]_  = A201 & ~A200;
  assign \new_[48328]_  = \new_[48327]_  & \new_[48324]_ ;
  assign \new_[48329]_  = \new_[48328]_  & \new_[48321]_ ;
  assign \new_[48333]_  = ~A234 & ~A233;
  assign \new_[48334]_  = A202 & \new_[48333]_ ;
  assign \new_[48337]_  = ~A266 & ~A265;
  assign \new_[48340]_  = A299 & ~A298;
  assign \new_[48341]_  = \new_[48340]_  & \new_[48337]_ ;
  assign \new_[48342]_  = \new_[48341]_  & \new_[48334]_ ;
  assign \new_[48346]_  = ~A167 & ~A168;
  assign \new_[48347]_  = A169 & \new_[48346]_ ;
  assign \new_[48350]_  = A199 & A166;
  assign \new_[48353]_  = A201 & ~A200;
  assign \new_[48354]_  = \new_[48353]_  & \new_[48350]_ ;
  assign \new_[48355]_  = \new_[48354]_  & \new_[48347]_ ;
  assign \new_[48359]_  = ~A233 & A232;
  assign \new_[48360]_  = A202 & \new_[48359]_ ;
  assign \new_[48363]_  = A235 & A234;
  assign \new_[48366]_  = ~A300 & A298;
  assign \new_[48367]_  = \new_[48366]_  & \new_[48363]_ ;
  assign \new_[48368]_  = \new_[48367]_  & \new_[48360]_ ;
  assign \new_[48372]_  = ~A167 & ~A168;
  assign \new_[48373]_  = A169 & \new_[48372]_ ;
  assign \new_[48376]_  = A199 & A166;
  assign \new_[48379]_  = A201 & ~A200;
  assign \new_[48380]_  = \new_[48379]_  & \new_[48376]_ ;
  assign \new_[48381]_  = \new_[48380]_  & \new_[48373]_ ;
  assign \new_[48385]_  = ~A233 & A232;
  assign \new_[48386]_  = A202 & \new_[48385]_ ;
  assign \new_[48389]_  = A235 & A234;
  assign \new_[48392]_  = A299 & A298;
  assign \new_[48393]_  = \new_[48392]_  & \new_[48389]_ ;
  assign \new_[48394]_  = \new_[48393]_  & \new_[48386]_ ;
  assign \new_[48398]_  = ~A167 & ~A168;
  assign \new_[48399]_  = A169 & \new_[48398]_ ;
  assign \new_[48402]_  = A199 & A166;
  assign \new_[48405]_  = A201 & ~A200;
  assign \new_[48406]_  = \new_[48405]_  & \new_[48402]_ ;
  assign \new_[48407]_  = \new_[48406]_  & \new_[48399]_ ;
  assign \new_[48411]_  = ~A233 & A232;
  assign \new_[48412]_  = A202 & \new_[48411]_ ;
  assign \new_[48415]_  = A235 & A234;
  assign \new_[48418]_  = ~A299 & ~A298;
  assign \new_[48419]_  = \new_[48418]_  & \new_[48415]_ ;
  assign \new_[48420]_  = \new_[48419]_  & \new_[48412]_ ;
  assign \new_[48424]_  = ~A167 & ~A168;
  assign \new_[48425]_  = A169 & \new_[48424]_ ;
  assign \new_[48428]_  = A199 & A166;
  assign \new_[48431]_  = A201 & ~A200;
  assign \new_[48432]_  = \new_[48431]_  & \new_[48428]_ ;
  assign \new_[48433]_  = \new_[48432]_  & \new_[48425]_ ;
  assign \new_[48437]_  = ~A233 & A232;
  assign \new_[48438]_  = A202 & \new_[48437]_ ;
  assign \new_[48441]_  = A235 & A234;
  assign \new_[48444]_  = A266 & ~A265;
  assign \new_[48445]_  = \new_[48444]_  & \new_[48441]_ ;
  assign \new_[48446]_  = \new_[48445]_  & \new_[48438]_ ;
  assign \new_[48450]_  = ~A167 & ~A168;
  assign \new_[48451]_  = A169 & \new_[48450]_ ;
  assign \new_[48454]_  = A199 & A166;
  assign \new_[48457]_  = A201 & ~A200;
  assign \new_[48458]_  = \new_[48457]_  & \new_[48454]_ ;
  assign \new_[48459]_  = \new_[48458]_  & \new_[48451]_ ;
  assign \new_[48463]_  = ~A233 & A232;
  assign \new_[48464]_  = A202 & \new_[48463]_ ;
  assign \new_[48467]_  = A236 & A234;
  assign \new_[48470]_  = ~A300 & A298;
  assign \new_[48471]_  = \new_[48470]_  & \new_[48467]_ ;
  assign \new_[48472]_  = \new_[48471]_  & \new_[48464]_ ;
  assign \new_[48476]_  = ~A167 & ~A168;
  assign \new_[48477]_  = A169 & \new_[48476]_ ;
  assign \new_[48480]_  = A199 & A166;
  assign \new_[48483]_  = A201 & ~A200;
  assign \new_[48484]_  = \new_[48483]_  & \new_[48480]_ ;
  assign \new_[48485]_  = \new_[48484]_  & \new_[48477]_ ;
  assign \new_[48489]_  = ~A233 & A232;
  assign \new_[48490]_  = A202 & \new_[48489]_ ;
  assign \new_[48493]_  = A236 & A234;
  assign \new_[48496]_  = A299 & A298;
  assign \new_[48497]_  = \new_[48496]_  & \new_[48493]_ ;
  assign \new_[48498]_  = \new_[48497]_  & \new_[48490]_ ;
  assign \new_[48502]_  = ~A167 & ~A168;
  assign \new_[48503]_  = A169 & \new_[48502]_ ;
  assign \new_[48506]_  = A199 & A166;
  assign \new_[48509]_  = A201 & ~A200;
  assign \new_[48510]_  = \new_[48509]_  & \new_[48506]_ ;
  assign \new_[48511]_  = \new_[48510]_  & \new_[48503]_ ;
  assign \new_[48515]_  = ~A233 & A232;
  assign \new_[48516]_  = A202 & \new_[48515]_ ;
  assign \new_[48519]_  = A236 & A234;
  assign \new_[48522]_  = ~A299 & ~A298;
  assign \new_[48523]_  = \new_[48522]_  & \new_[48519]_ ;
  assign \new_[48524]_  = \new_[48523]_  & \new_[48516]_ ;
  assign \new_[48528]_  = ~A167 & ~A168;
  assign \new_[48529]_  = A169 & \new_[48528]_ ;
  assign \new_[48532]_  = A199 & A166;
  assign \new_[48535]_  = A201 & ~A200;
  assign \new_[48536]_  = \new_[48535]_  & \new_[48532]_ ;
  assign \new_[48537]_  = \new_[48536]_  & \new_[48529]_ ;
  assign \new_[48541]_  = ~A233 & A232;
  assign \new_[48542]_  = A202 & \new_[48541]_ ;
  assign \new_[48545]_  = A236 & A234;
  assign \new_[48548]_  = A266 & ~A265;
  assign \new_[48549]_  = \new_[48548]_  & \new_[48545]_ ;
  assign \new_[48550]_  = \new_[48549]_  & \new_[48542]_ ;
  assign \new_[48554]_  = ~A167 & ~A168;
  assign \new_[48555]_  = A169 & \new_[48554]_ ;
  assign \new_[48558]_  = A199 & A166;
  assign \new_[48561]_  = A201 & ~A200;
  assign \new_[48562]_  = \new_[48561]_  & \new_[48558]_ ;
  assign \new_[48563]_  = \new_[48562]_  & \new_[48555]_ ;
  assign \new_[48567]_  = ~A233 & ~A232;
  assign \new_[48568]_  = A202 & \new_[48567]_ ;
  assign \new_[48571]_  = A266 & A265;
  assign \new_[48574]_  = A299 & ~A298;
  assign \new_[48575]_  = \new_[48574]_  & \new_[48571]_ ;
  assign \new_[48576]_  = \new_[48575]_  & \new_[48568]_ ;
  assign \new_[48580]_  = ~A167 & ~A168;
  assign \new_[48581]_  = A169 & \new_[48580]_ ;
  assign \new_[48584]_  = A199 & A166;
  assign \new_[48587]_  = A201 & ~A200;
  assign \new_[48588]_  = \new_[48587]_  & \new_[48584]_ ;
  assign \new_[48589]_  = \new_[48588]_  & \new_[48581]_ ;
  assign \new_[48593]_  = ~A233 & ~A232;
  assign \new_[48594]_  = A202 & \new_[48593]_ ;
  assign \new_[48597]_  = ~A267 & ~A266;
  assign \new_[48600]_  = A299 & ~A298;
  assign \new_[48601]_  = \new_[48600]_  & \new_[48597]_ ;
  assign \new_[48602]_  = \new_[48601]_  & \new_[48594]_ ;
  assign \new_[48606]_  = ~A167 & ~A168;
  assign \new_[48607]_  = A169 & \new_[48606]_ ;
  assign \new_[48610]_  = A199 & A166;
  assign \new_[48613]_  = A201 & ~A200;
  assign \new_[48614]_  = \new_[48613]_  & \new_[48610]_ ;
  assign \new_[48615]_  = \new_[48614]_  & \new_[48607]_ ;
  assign \new_[48619]_  = ~A233 & ~A232;
  assign \new_[48620]_  = A202 & \new_[48619]_ ;
  assign \new_[48623]_  = ~A266 & ~A265;
  assign \new_[48626]_  = A299 & ~A298;
  assign \new_[48627]_  = \new_[48626]_  & \new_[48623]_ ;
  assign \new_[48628]_  = \new_[48627]_  & \new_[48620]_ ;
  assign \new_[48632]_  = ~A167 & ~A168;
  assign \new_[48633]_  = A169 & \new_[48632]_ ;
  assign \new_[48636]_  = A199 & A166;
  assign \new_[48639]_  = A201 & ~A200;
  assign \new_[48640]_  = \new_[48639]_  & \new_[48636]_ ;
  assign \new_[48641]_  = \new_[48640]_  & \new_[48633]_ ;
  assign \new_[48645]_  = A233 & A232;
  assign \new_[48646]_  = A203 & \new_[48645]_ ;
  assign \new_[48649]_  = ~A267 & A265;
  assign \new_[48652]_  = A299 & ~A298;
  assign \new_[48653]_  = \new_[48652]_  & \new_[48649]_ ;
  assign \new_[48654]_  = \new_[48653]_  & \new_[48646]_ ;
  assign \new_[48658]_  = ~A167 & ~A168;
  assign \new_[48659]_  = A169 & \new_[48658]_ ;
  assign \new_[48662]_  = A199 & A166;
  assign \new_[48665]_  = A201 & ~A200;
  assign \new_[48666]_  = \new_[48665]_  & \new_[48662]_ ;
  assign \new_[48667]_  = \new_[48666]_  & \new_[48659]_ ;
  assign \new_[48671]_  = A233 & A232;
  assign \new_[48672]_  = A203 & \new_[48671]_ ;
  assign \new_[48675]_  = A266 & A265;
  assign \new_[48678]_  = A299 & ~A298;
  assign \new_[48679]_  = \new_[48678]_  & \new_[48675]_ ;
  assign \new_[48680]_  = \new_[48679]_  & \new_[48672]_ ;
  assign \new_[48684]_  = ~A167 & ~A168;
  assign \new_[48685]_  = A169 & \new_[48684]_ ;
  assign \new_[48688]_  = A199 & A166;
  assign \new_[48691]_  = A201 & ~A200;
  assign \new_[48692]_  = \new_[48691]_  & \new_[48688]_ ;
  assign \new_[48693]_  = \new_[48692]_  & \new_[48685]_ ;
  assign \new_[48697]_  = A233 & A232;
  assign \new_[48698]_  = A203 & \new_[48697]_ ;
  assign \new_[48701]_  = ~A266 & ~A265;
  assign \new_[48704]_  = A299 & ~A298;
  assign \new_[48705]_  = \new_[48704]_  & \new_[48701]_ ;
  assign \new_[48706]_  = \new_[48705]_  & \new_[48698]_ ;
  assign \new_[48710]_  = ~A167 & ~A168;
  assign \new_[48711]_  = A169 & \new_[48710]_ ;
  assign \new_[48714]_  = A199 & A166;
  assign \new_[48717]_  = A201 & ~A200;
  assign \new_[48718]_  = \new_[48717]_  & \new_[48714]_ ;
  assign \new_[48719]_  = \new_[48718]_  & \new_[48711]_ ;
  assign \new_[48723]_  = A233 & ~A232;
  assign \new_[48724]_  = A203 & \new_[48723]_ ;
  assign \new_[48727]_  = ~A266 & A265;
  assign \new_[48730]_  = A268 & A267;
  assign \new_[48731]_  = \new_[48730]_  & \new_[48727]_ ;
  assign \new_[48732]_  = \new_[48731]_  & \new_[48724]_ ;
  assign \new_[48736]_  = ~A167 & ~A168;
  assign \new_[48737]_  = A169 & \new_[48736]_ ;
  assign \new_[48740]_  = A199 & A166;
  assign \new_[48743]_  = A201 & ~A200;
  assign \new_[48744]_  = \new_[48743]_  & \new_[48740]_ ;
  assign \new_[48745]_  = \new_[48744]_  & \new_[48737]_ ;
  assign \new_[48749]_  = A233 & ~A232;
  assign \new_[48750]_  = A203 & \new_[48749]_ ;
  assign \new_[48753]_  = ~A266 & A265;
  assign \new_[48756]_  = A269 & A267;
  assign \new_[48757]_  = \new_[48756]_  & \new_[48753]_ ;
  assign \new_[48758]_  = \new_[48757]_  & \new_[48750]_ ;
  assign \new_[48762]_  = ~A167 & ~A168;
  assign \new_[48763]_  = A169 & \new_[48762]_ ;
  assign \new_[48766]_  = A199 & A166;
  assign \new_[48769]_  = A201 & ~A200;
  assign \new_[48770]_  = \new_[48769]_  & \new_[48766]_ ;
  assign \new_[48771]_  = \new_[48770]_  & \new_[48763]_ ;
  assign \new_[48775]_  = ~A234 & ~A233;
  assign \new_[48776]_  = A203 & \new_[48775]_ ;
  assign \new_[48779]_  = A266 & A265;
  assign \new_[48782]_  = A299 & ~A298;
  assign \new_[48783]_  = \new_[48782]_  & \new_[48779]_ ;
  assign \new_[48784]_  = \new_[48783]_  & \new_[48776]_ ;
  assign \new_[48788]_  = ~A167 & ~A168;
  assign \new_[48789]_  = A169 & \new_[48788]_ ;
  assign \new_[48792]_  = A199 & A166;
  assign \new_[48795]_  = A201 & ~A200;
  assign \new_[48796]_  = \new_[48795]_  & \new_[48792]_ ;
  assign \new_[48797]_  = \new_[48796]_  & \new_[48789]_ ;
  assign \new_[48801]_  = ~A234 & ~A233;
  assign \new_[48802]_  = A203 & \new_[48801]_ ;
  assign \new_[48805]_  = ~A267 & ~A266;
  assign \new_[48808]_  = A299 & ~A298;
  assign \new_[48809]_  = \new_[48808]_  & \new_[48805]_ ;
  assign \new_[48810]_  = \new_[48809]_  & \new_[48802]_ ;
  assign \new_[48814]_  = ~A167 & ~A168;
  assign \new_[48815]_  = A169 & \new_[48814]_ ;
  assign \new_[48818]_  = A199 & A166;
  assign \new_[48821]_  = A201 & ~A200;
  assign \new_[48822]_  = \new_[48821]_  & \new_[48818]_ ;
  assign \new_[48823]_  = \new_[48822]_  & \new_[48815]_ ;
  assign \new_[48827]_  = ~A234 & ~A233;
  assign \new_[48828]_  = A203 & \new_[48827]_ ;
  assign \new_[48831]_  = ~A266 & ~A265;
  assign \new_[48834]_  = A299 & ~A298;
  assign \new_[48835]_  = \new_[48834]_  & \new_[48831]_ ;
  assign \new_[48836]_  = \new_[48835]_  & \new_[48828]_ ;
  assign \new_[48840]_  = ~A167 & ~A168;
  assign \new_[48841]_  = A169 & \new_[48840]_ ;
  assign \new_[48844]_  = A199 & A166;
  assign \new_[48847]_  = A201 & ~A200;
  assign \new_[48848]_  = \new_[48847]_  & \new_[48844]_ ;
  assign \new_[48849]_  = \new_[48848]_  & \new_[48841]_ ;
  assign \new_[48853]_  = ~A233 & A232;
  assign \new_[48854]_  = A203 & \new_[48853]_ ;
  assign \new_[48857]_  = A235 & A234;
  assign \new_[48860]_  = ~A300 & A298;
  assign \new_[48861]_  = \new_[48860]_  & \new_[48857]_ ;
  assign \new_[48862]_  = \new_[48861]_  & \new_[48854]_ ;
  assign \new_[48866]_  = ~A167 & ~A168;
  assign \new_[48867]_  = A169 & \new_[48866]_ ;
  assign \new_[48870]_  = A199 & A166;
  assign \new_[48873]_  = A201 & ~A200;
  assign \new_[48874]_  = \new_[48873]_  & \new_[48870]_ ;
  assign \new_[48875]_  = \new_[48874]_  & \new_[48867]_ ;
  assign \new_[48879]_  = ~A233 & A232;
  assign \new_[48880]_  = A203 & \new_[48879]_ ;
  assign \new_[48883]_  = A235 & A234;
  assign \new_[48886]_  = A299 & A298;
  assign \new_[48887]_  = \new_[48886]_  & \new_[48883]_ ;
  assign \new_[48888]_  = \new_[48887]_  & \new_[48880]_ ;
  assign \new_[48892]_  = ~A167 & ~A168;
  assign \new_[48893]_  = A169 & \new_[48892]_ ;
  assign \new_[48896]_  = A199 & A166;
  assign \new_[48899]_  = A201 & ~A200;
  assign \new_[48900]_  = \new_[48899]_  & \new_[48896]_ ;
  assign \new_[48901]_  = \new_[48900]_  & \new_[48893]_ ;
  assign \new_[48905]_  = ~A233 & A232;
  assign \new_[48906]_  = A203 & \new_[48905]_ ;
  assign \new_[48909]_  = A235 & A234;
  assign \new_[48912]_  = ~A299 & ~A298;
  assign \new_[48913]_  = \new_[48912]_  & \new_[48909]_ ;
  assign \new_[48914]_  = \new_[48913]_  & \new_[48906]_ ;
  assign \new_[48918]_  = ~A167 & ~A168;
  assign \new_[48919]_  = A169 & \new_[48918]_ ;
  assign \new_[48922]_  = A199 & A166;
  assign \new_[48925]_  = A201 & ~A200;
  assign \new_[48926]_  = \new_[48925]_  & \new_[48922]_ ;
  assign \new_[48927]_  = \new_[48926]_  & \new_[48919]_ ;
  assign \new_[48931]_  = ~A233 & A232;
  assign \new_[48932]_  = A203 & \new_[48931]_ ;
  assign \new_[48935]_  = A235 & A234;
  assign \new_[48938]_  = A266 & ~A265;
  assign \new_[48939]_  = \new_[48938]_  & \new_[48935]_ ;
  assign \new_[48940]_  = \new_[48939]_  & \new_[48932]_ ;
  assign \new_[48944]_  = ~A167 & ~A168;
  assign \new_[48945]_  = A169 & \new_[48944]_ ;
  assign \new_[48948]_  = A199 & A166;
  assign \new_[48951]_  = A201 & ~A200;
  assign \new_[48952]_  = \new_[48951]_  & \new_[48948]_ ;
  assign \new_[48953]_  = \new_[48952]_  & \new_[48945]_ ;
  assign \new_[48957]_  = ~A233 & A232;
  assign \new_[48958]_  = A203 & \new_[48957]_ ;
  assign \new_[48961]_  = A236 & A234;
  assign \new_[48964]_  = ~A300 & A298;
  assign \new_[48965]_  = \new_[48964]_  & \new_[48961]_ ;
  assign \new_[48966]_  = \new_[48965]_  & \new_[48958]_ ;
  assign \new_[48970]_  = ~A167 & ~A168;
  assign \new_[48971]_  = A169 & \new_[48970]_ ;
  assign \new_[48974]_  = A199 & A166;
  assign \new_[48977]_  = A201 & ~A200;
  assign \new_[48978]_  = \new_[48977]_  & \new_[48974]_ ;
  assign \new_[48979]_  = \new_[48978]_  & \new_[48971]_ ;
  assign \new_[48983]_  = ~A233 & A232;
  assign \new_[48984]_  = A203 & \new_[48983]_ ;
  assign \new_[48987]_  = A236 & A234;
  assign \new_[48990]_  = A299 & A298;
  assign \new_[48991]_  = \new_[48990]_  & \new_[48987]_ ;
  assign \new_[48992]_  = \new_[48991]_  & \new_[48984]_ ;
  assign \new_[48996]_  = ~A167 & ~A168;
  assign \new_[48997]_  = A169 & \new_[48996]_ ;
  assign \new_[49000]_  = A199 & A166;
  assign \new_[49003]_  = A201 & ~A200;
  assign \new_[49004]_  = \new_[49003]_  & \new_[49000]_ ;
  assign \new_[49005]_  = \new_[49004]_  & \new_[48997]_ ;
  assign \new_[49009]_  = ~A233 & A232;
  assign \new_[49010]_  = A203 & \new_[49009]_ ;
  assign \new_[49013]_  = A236 & A234;
  assign \new_[49016]_  = ~A299 & ~A298;
  assign \new_[49017]_  = \new_[49016]_  & \new_[49013]_ ;
  assign \new_[49018]_  = \new_[49017]_  & \new_[49010]_ ;
  assign \new_[49022]_  = ~A167 & ~A168;
  assign \new_[49023]_  = A169 & \new_[49022]_ ;
  assign \new_[49026]_  = A199 & A166;
  assign \new_[49029]_  = A201 & ~A200;
  assign \new_[49030]_  = \new_[49029]_  & \new_[49026]_ ;
  assign \new_[49031]_  = \new_[49030]_  & \new_[49023]_ ;
  assign \new_[49035]_  = ~A233 & A232;
  assign \new_[49036]_  = A203 & \new_[49035]_ ;
  assign \new_[49039]_  = A236 & A234;
  assign \new_[49042]_  = A266 & ~A265;
  assign \new_[49043]_  = \new_[49042]_  & \new_[49039]_ ;
  assign \new_[49044]_  = \new_[49043]_  & \new_[49036]_ ;
  assign \new_[49048]_  = ~A167 & ~A168;
  assign \new_[49049]_  = A169 & \new_[49048]_ ;
  assign \new_[49052]_  = A199 & A166;
  assign \new_[49055]_  = A201 & ~A200;
  assign \new_[49056]_  = \new_[49055]_  & \new_[49052]_ ;
  assign \new_[49057]_  = \new_[49056]_  & \new_[49049]_ ;
  assign \new_[49061]_  = ~A233 & ~A232;
  assign \new_[49062]_  = A203 & \new_[49061]_ ;
  assign \new_[49065]_  = A266 & A265;
  assign \new_[49068]_  = A299 & ~A298;
  assign \new_[49069]_  = \new_[49068]_  & \new_[49065]_ ;
  assign \new_[49070]_  = \new_[49069]_  & \new_[49062]_ ;
  assign \new_[49074]_  = ~A167 & ~A168;
  assign \new_[49075]_  = A169 & \new_[49074]_ ;
  assign \new_[49078]_  = A199 & A166;
  assign \new_[49081]_  = A201 & ~A200;
  assign \new_[49082]_  = \new_[49081]_  & \new_[49078]_ ;
  assign \new_[49083]_  = \new_[49082]_  & \new_[49075]_ ;
  assign \new_[49087]_  = ~A233 & ~A232;
  assign \new_[49088]_  = A203 & \new_[49087]_ ;
  assign \new_[49091]_  = ~A267 & ~A266;
  assign \new_[49094]_  = A299 & ~A298;
  assign \new_[49095]_  = \new_[49094]_  & \new_[49091]_ ;
  assign \new_[49096]_  = \new_[49095]_  & \new_[49088]_ ;
  assign \new_[49100]_  = ~A167 & ~A168;
  assign \new_[49101]_  = A169 & \new_[49100]_ ;
  assign \new_[49104]_  = A199 & A166;
  assign \new_[49107]_  = A201 & ~A200;
  assign \new_[49108]_  = \new_[49107]_  & \new_[49104]_ ;
  assign \new_[49109]_  = \new_[49108]_  & \new_[49101]_ ;
  assign \new_[49113]_  = ~A233 & ~A232;
  assign \new_[49114]_  = A203 & \new_[49113]_ ;
  assign \new_[49117]_  = ~A266 & ~A265;
  assign \new_[49120]_  = A299 & ~A298;
  assign \new_[49121]_  = \new_[49120]_  & \new_[49117]_ ;
  assign \new_[49122]_  = \new_[49121]_  & \new_[49114]_ ;
  assign \new_[49126]_  = ~A168 & A169;
  assign \new_[49127]_  = A170 & \new_[49126]_ ;
  assign \new_[49130]_  = ~A200 & A199;
  assign \new_[49133]_  = A202 & A201;
  assign \new_[49134]_  = \new_[49133]_  & \new_[49130]_ ;
  assign \new_[49135]_  = \new_[49134]_  & \new_[49127]_ ;
  assign \new_[49139]_  = A265 & A233;
  assign \new_[49140]_  = A232 & \new_[49139]_ ;
  assign \new_[49143]_  = ~A269 & ~A268;
  assign \new_[49146]_  = A299 & ~A298;
  assign \new_[49147]_  = \new_[49146]_  & \new_[49143]_ ;
  assign \new_[49148]_  = \new_[49147]_  & \new_[49140]_ ;
  assign \new_[49152]_  = ~A168 & A169;
  assign \new_[49153]_  = A170 & \new_[49152]_ ;
  assign \new_[49156]_  = ~A200 & A199;
  assign \new_[49159]_  = A202 & A201;
  assign \new_[49160]_  = \new_[49159]_  & \new_[49156]_ ;
  assign \new_[49161]_  = \new_[49160]_  & \new_[49153]_ ;
  assign \new_[49165]_  = ~A236 & ~A235;
  assign \new_[49166]_  = ~A233 & \new_[49165]_ ;
  assign \new_[49169]_  = A266 & A265;
  assign \new_[49172]_  = A299 & ~A298;
  assign \new_[49173]_  = \new_[49172]_  & \new_[49169]_ ;
  assign \new_[49174]_  = \new_[49173]_  & \new_[49166]_ ;
  assign \new_[49178]_  = ~A168 & A169;
  assign \new_[49179]_  = A170 & \new_[49178]_ ;
  assign \new_[49182]_  = ~A200 & A199;
  assign \new_[49185]_  = A202 & A201;
  assign \new_[49186]_  = \new_[49185]_  & \new_[49182]_ ;
  assign \new_[49187]_  = \new_[49186]_  & \new_[49179]_ ;
  assign \new_[49191]_  = ~A236 & ~A235;
  assign \new_[49192]_  = ~A233 & \new_[49191]_ ;
  assign \new_[49195]_  = ~A267 & ~A266;
  assign \new_[49198]_  = A299 & ~A298;
  assign \new_[49199]_  = \new_[49198]_  & \new_[49195]_ ;
  assign \new_[49200]_  = \new_[49199]_  & \new_[49192]_ ;
  assign \new_[49204]_  = ~A168 & A169;
  assign \new_[49205]_  = A170 & \new_[49204]_ ;
  assign \new_[49208]_  = ~A200 & A199;
  assign \new_[49211]_  = A202 & A201;
  assign \new_[49212]_  = \new_[49211]_  & \new_[49208]_ ;
  assign \new_[49213]_  = \new_[49212]_  & \new_[49205]_ ;
  assign \new_[49217]_  = ~A236 & ~A235;
  assign \new_[49218]_  = ~A233 & \new_[49217]_ ;
  assign \new_[49221]_  = ~A266 & ~A265;
  assign \new_[49224]_  = A299 & ~A298;
  assign \new_[49225]_  = \new_[49224]_  & \new_[49221]_ ;
  assign \new_[49226]_  = \new_[49225]_  & \new_[49218]_ ;
  assign \new_[49230]_  = ~A168 & A169;
  assign \new_[49231]_  = A170 & \new_[49230]_ ;
  assign \new_[49234]_  = ~A200 & A199;
  assign \new_[49237]_  = A202 & A201;
  assign \new_[49238]_  = \new_[49237]_  & \new_[49234]_ ;
  assign \new_[49239]_  = \new_[49238]_  & \new_[49231]_ ;
  assign \new_[49243]_  = ~A266 & ~A234;
  assign \new_[49244]_  = ~A233 & \new_[49243]_ ;
  assign \new_[49247]_  = ~A269 & ~A268;
  assign \new_[49250]_  = A299 & ~A298;
  assign \new_[49251]_  = \new_[49250]_  & \new_[49247]_ ;
  assign \new_[49252]_  = \new_[49251]_  & \new_[49244]_ ;
  assign \new_[49256]_  = ~A168 & A169;
  assign \new_[49257]_  = A170 & \new_[49256]_ ;
  assign \new_[49260]_  = ~A200 & A199;
  assign \new_[49263]_  = A202 & A201;
  assign \new_[49264]_  = \new_[49263]_  & \new_[49260]_ ;
  assign \new_[49265]_  = \new_[49264]_  & \new_[49257]_ ;
  assign \new_[49269]_  = A234 & ~A233;
  assign \new_[49270]_  = A232 & \new_[49269]_ ;
  assign \new_[49273]_  = A298 & A235;
  assign \new_[49276]_  = ~A302 & ~A301;
  assign \new_[49277]_  = \new_[49276]_  & \new_[49273]_ ;
  assign \new_[49278]_  = \new_[49277]_  & \new_[49270]_ ;
  assign \new_[49282]_  = ~A168 & A169;
  assign \new_[49283]_  = A170 & \new_[49282]_ ;
  assign \new_[49286]_  = ~A200 & A199;
  assign \new_[49289]_  = A202 & A201;
  assign \new_[49290]_  = \new_[49289]_  & \new_[49286]_ ;
  assign \new_[49291]_  = \new_[49290]_  & \new_[49283]_ ;
  assign \new_[49295]_  = A234 & ~A233;
  assign \new_[49296]_  = A232 & \new_[49295]_ ;
  assign \new_[49299]_  = A298 & A236;
  assign \new_[49302]_  = ~A302 & ~A301;
  assign \new_[49303]_  = \new_[49302]_  & \new_[49299]_ ;
  assign \new_[49304]_  = \new_[49303]_  & \new_[49296]_ ;
  assign \new_[49308]_  = ~A168 & A169;
  assign \new_[49309]_  = A170 & \new_[49308]_ ;
  assign \new_[49312]_  = ~A200 & A199;
  assign \new_[49315]_  = A202 & A201;
  assign \new_[49316]_  = \new_[49315]_  & \new_[49312]_ ;
  assign \new_[49317]_  = \new_[49316]_  & \new_[49309]_ ;
  assign \new_[49321]_  = ~A266 & ~A233;
  assign \new_[49322]_  = ~A232 & \new_[49321]_ ;
  assign \new_[49325]_  = ~A269 & ~A268;
  assign \new_[49328]_  = A299 & ~A298;
  assign \new_[49329]_  = \new_[49328]_  & \new_[49325]_ ;
  assign \new_[49330]_  = \new_[49329]_  & \new_[49322]_ ;
  assign \new_[49334]_  = ~A168 & A169;
  assign \new_[49335]_  = A170 & \new_[49334]_ ;
  assign \new_[49338]_  = ~A200 & A199;
  assign \new_[49341]_  = A203 & A201;
  assign \new_[49342]_  = \new_[49341]_  & \new_[49338]_ ;
  assign \new_[49343]_  = \new_[49342]_  & \new_[49335]_ ;
  assign \new_[49347]_  = A265 & A233;
  assign \new_[49348]_  = A232 & \new_[49347]_ ;
  assign \new_[49351]_  = ~A269 & ~A268;
  assign \new_[49354]_  = A299 & ~A298;
  assign \new_[49355]_  = \new_[49354]_  & \new_[49351]_ ;
  assign \new_[49356]_  = \new_[49355]_  & \new_[49348]_ ;
  assign \new_[49360]_  = ~A168 & A169;
  assign \new_[49361]_  = A170 & \new_[49360]_ ;
  assign \new_[49364]_  = ~A200 & A199;
  assign \new_[49367]_  = A203 & A201;
  assign \new_[49368]_  = \new_[49367]_  & \new_[49364]_ ;
  assign \new_[49369]_  = \new_[49368]_  & \new_[49361]_ ;
  assign \new_[49373]_  = ~A236 & ~A235;
  assign \new_[49374]_  = ~A233 & \new_[49373]_ ;
  assign \new_[49377]_  = A266 & A265;
  assign \new_[49380]_  = A299 & ~A298;
  assign \new_[49381]_  = \new_[49380]_  & \new_[49377]_ ;
  assign \new_[49382]_  = \new_[49381]_  & \new_[49374]_ ;
  assign \new_[49386]_  = ~A168 & A169;
  assign \new_[49387]_  = A170 & \new_[49386]_ ;
  assign \new_[49390]_  = ~A200 & A199;
  assign \new_[49393]_  = A203 & A201;
  assign \new_[49394]_  = \new_[49393]_  & \new_[49390]_ ;
  assign \new_[49395]_  = \new_[49394]_  & \new_[49387]_ ;
  assign \new_[49399]_  = ~A236 & ~A235;
  assign \new_[49400]_  = ~A233 & \new_[49399]_ ;
  assign \new_[49403]_  = ~A267 & ~A266;
  assign \new_[49406]_  = A299 & ~A298;
  assign \new_[49407]_  = \new_[49406]_  & \new_[49403]_ ;
  assign \new_[49408]_  = \new_[49407]_  & \new_[49400]_ ;
  assign \new_[49412]_  = ~A168 & A169;
  assign \new_[49413]_  = A170 & \new_[49412]_ ;
  assign \new_[49416]_  = ~A200 & A199;
  assign \new_[49419]_  = A203 & A201;
  assign \new_[49420]_  = \new_[49419]_  & \new_[49416]_ ;
  assign \new_[49421]_  = \new_[49420]_  & \new_[49413]_ ;
  assign \new_[49425]_  = ~A236 & ~A235;
  assign \new_[49426]_  = ~A233 & \new_[49425]_ ;
  assign \new_[49429]_  = ~A266 & ~A265;
  assign \new_[49432]_  = A299 & ~A298;
  assign \new_[49433]_  = \new_[49432]_  & \new_[49429]_ ;
  assign \new_[49434]_  = \new_[49433]_  & \new_[49426]_ ;
  assign \new_[49438]_  = ~A168 & A169;
  assign \new_[49439]_  = A170 & \new_[49438]_ ;
  assign \new_[49442]_  = ~A200 & A199;
  assign \new_[49445]_  = A203 & A201;
  assign \new_[49446]_  = \new_[49445]_  & \new_[49442]_ ;
  assign \new_[49447]_  = \new_[49446]_  & \new_[49439]_ ;
  assign \new_[49451]_  = ~A266 & ~A234;
  assign \new_[49452]_  = ~A233 & \new_[49451]_ ;
  assign \new_[49455]_  = ~A269 & ~A268;
  assign \new_[49458]_  = A299 & ~A298;
  assign \new_[49459]_  = \new_[49458]_  & \new_[49455]_ ;
  assign \new_[49460]_  = \new_[49459]_  & \new_[49452]_ ;
  assign \new_[49464]_  = ~A168 & A169;
  assign \new_[49465]_  = A170 & \new_[49464]_ ;
  assign \new_[49468]_  = ~A200 & A199;
  assign \new_[49471]_  = A203 & A201;
  assign \new_[49472]_  = \new_[49471]_  & \new_[49468]_ ;
  assign \new_[49473]_  = \new_[49472]_  & \new_[49465]_ ;
  assign \new_[49477]_  = A234 & ~A233;
  assign \new_[49478]_  = A232 & \new_[49477]_ ;
  assign \new_[49481]_  = A298 & A235;
  assign \new_[49484]_  = ~A302 & ~A301;
  assign \new_[49485]_  = \new_[49484]_  & \new_[49481]_ ;
  assign \new_[49486]_  = \new_[49485]_  & \new_[49478]_ ;
  assign \new_[49490]_  = ~A168 & A169;
  assign \new_[49491]_  = A170 & \new_[49490]_ ;
  assign \new_[49494]_  = ~A200 & A199;
  assign \new_[49497]_  = A203 & A201;
  assign \new_[49498]_  = \new_[49497]_  & \new_[49494]_ ;
  assign \new_[49499]_  = \new_[49498]_  & \new_[49491]_ ;
  assign \new_[49503]_  = A234 & ~A233;
  assign \new_[49504]_  = A232 & \new_[49503]_ ;
  assign \new_[49507]_  = A298 & A236;
  assign \new_[49510]_  = ~A302 & ~A301;
  assign \new_[49511]_  = \new_[49510]_  & \new_[49507]_ ;
  assign \new_[49512]_  = \new_[49511]_  & \new_[49504]_ ;
  assign \new_[49516]_  = ~A168 & A169;
  assign \new_[49517]_  = A170 & \new_[49516]_ ;
  assign \new_[49520]_  = ~A200 & A199;
  assign \new_[49523]_  = A203 & A201;
  assign \new_[49524]_  = \new_[49523]_  & \new_[49520]_ ;
  assign \new_[49525]_  = \new_[49524]_  & \new_[49517]_ ;
  assign \new_[49529]_  = ~A266 & ~A233;
  assign \new_[49530]_  = ~A232 & \new_[49529]_ ;
  assign \new_[49533]_  = ~A269 & ~A268;
  assign \new_[49536]_  = A299 & ~A298;
  assign \new_[49537]_  = \new_[49536]_  & \new_[49533]_ ;
  assign \new_[49538]_  = \new_[49537]_  & \new_[49530]_ ;
  assign \new_[49542]_  = A167 & A169;
  assign \new_[49543]_  = ~A170 & \new_[49542]_ ;
  assign \new_[49546]_  = A199 & A166;
  assign \new_[49549]_  = A232 & A200;
  assign \new_[49550]_  = \new_[49549]_  & \new_[49546]_ ;
  assign \new_[49551]_  = \new_[49550]_  & \new_[49543]_ ;
  assign \new_[49555]_  = ~A267 & A265;
  assign \new_[49556]_  = A233 & \new_[49555]_ ;
  assign \new_[49559]_  = ~A299 & A298;
  assign \new_[49562]_  = A301 & A300;
  assign \new_[49563]_  = \new_[49562]_  & \new_[49559]_ ;
  assign \new_[49564]_  = \new_[49563]_  & \new_[49556]_ ;
  assign \new_[49568]_  = A167 & A169;
  assign \new_[49569]_  = ~A170 & \new_[49568]_ ;
  assign \new_[49572]_  = A199 & A166;
  assign \new_[49575]_  = A232 & A200;
  assign \new_[49576]_  = \new_[49575]_  & \new_[49572]_ ;
  assign \new_[49577]_  = \new_[49576]_  & \new_[49569]_ ;
  assign \new_[49581]_  = ~A267 & A265;
  assign \new_[49582]_  = A233 & \new_[49581]_ ;
  assign \new_[49585]_  = ~A299 & A298;
  assign \new_[49588]_  = A302 & A300;
  assign \new_[49589]_  = \new_[49588]_  & \new_[49585]_ ;
  assign \new_[49590]_  = \new_[49589]_  & \new_[49582]_ ;
  assign \new_[49594]_  = A167 & A169;
  assign \new_[49595]_  = ~A170 & \new_[49594]_ ;
  assign \new_[49598]_  = A199 & A166;
  assign \new_[49601]_  = A232 & A200;
  assign \new_[49602]_  = \new_[49601]_  & \new_[49598]_ ;
  assign \new_[49603]_  = \new_[49602]_  & \new_[49595]_ ;
  assign \new_[49607]_  = A266 & A265;
  assign \new_[49608]_  = A233 & \new_[49607]_ ;
  assign \new_[49611]_  = ~A299 & A298;
  assign \new_[49614]_  = A301 & A300;
  assign \new_[49615]_  = \new_[49614]_  & \new_[49611]_ ;
  assign \new_[49616]_  = \new_[49615]_  & \new_[49608]_ ;
  assign \new_[49620]_  = A167 & A169;
  assign \new_[49621]_  = ~A170 & \new_[49620]_ ;
  assign \new_[49624]_  = A199 & A166;
  assign \new_[49627]_  = A232 & A200;
  assign \new_[49628]_  = \new_[49627]_  & \new_[49624]_ ;
  assign \new_[49629]_  = \new_[49628]_  & \new_[49621]_ ;
  assign \new_[49633]_  = A266 & A265;
  assign \new_[49634]_  = A233 & \new_[49633]_ ;
  assign \new_[49637]_  = ~A299 & A298;
  assign \new_[49640]_  = A302 & A300;
  assign \new_[49641]_  = \new_[49640]_  & \new_[49637]_ ;
  assign \new_[49642]_  = \new_[49641]_  & \new_[49634]_ ;
  assign \new_[49646]_  = A167 & A169;
  assign \new_[49647]_  = ~A170 & \new_[49646]_ ;
  assign \new_[49650]_  = A199 & A166;
  assign \new_[49653]_  = A232 & A200;
  assign \new_[49654]_  = \new_[49653]_  & \new_[49650]_ ;
  assign \new_[49655]_  = \new_[49654]_  & \new_[49647]_ ;
  assign \new_[49659]_  = ~A266 & ~A265;
  assign \new_[49660]_  = A233 & \new_[49659]_ ;
  assign \new_[49663]_  = ~A299 & A298;
  assign \new_[49666]_  = A301 & A300;
  assign \new_[49667]_  = \new_[49666]_  & \new_[49663]_ ;
  assign \new_[49668]_  = \new_[49667]_  & \new_[49660]_ ;
  assign \new_[49672]_  = A167 & A169;
  assign \new_[49673]_  = ~A170 & \new_[49672]_ ;
  assign \new_[49676]_  = A199 & A166;
  assign \new_[49679]_  = A232 & A200;
  assign \new_[49680]_  = \new_[49679]_  & \new_[49676]_ ;
  assign \new_[49681]_  = \new_[49680]_  & \new_[49673]_ ;
  assign \new_[49685]_  = ~A266 & ~A265;
  assign \new_[49686]_  = A233 & \new_[49685]_ ;
  assign \new_[49689]_  = ~A299 & A298;
  assign \new_[49692]_  = A302 & A300;
  assign \new_[49693]_  = \new_[49692]_  & \new_[49689]_ ;
  assign \new_[49694]_  = \new_[49693]_  & \new_[49686]_ ;
  assign \new_[49698]_  = A167 & A169;
  assign \new_[49699]_  = ~A170 & \new_[49698]_ ;
  assign \new_[49702]_  = A199 & A166;
  assign \new_[49705]_  = ~A233 & A200;
  assign \new_[49706]_  = \new_[49705]_  & \new_[49702]_ ;
  assign \new_[49707]_  = \new_[49706]_  & \new_[49699]_ ;
  assign \new_[49711]_  = ~A266 & ~A236;
  assign \new_[49712]_  = ~A235 & \new_[49711]_ ;
  assign \new_[49715]_  = ~A269 & ~A268;
  assign \new_[49718]_  = A299 & ~A298;
  assign \new_[49719]_  = \new_[49718]_  & \new_[49715]_ ;
  assign \new_[49720]_  = \new_[49719]_  & \new_[49712]_ ;
  assign \new_[49724]_  = A167 & A169;
  assign \new_[49725]_  = ~A170 & \new_[49724]_ ;
  assign \new_[49728]_  = A199 & A166;
  assign \new_[49731]_  = ~A233 & A200;
  assign \new_[49732]_  = \new_[49731]_  & \new_[49728]_ ;
  assign \new_[49733]_  = \new_[49732]_  & \new_[49725]_ ;
  assign \new_[49737]_  = A266 & A265;
  assign \new_[49738]_  = ~A234 & \new_[49737]_ ;
  assign \new_[49741]_  = ~A299 & A298;
  assign \new_[49744]_  = A301 & A300;
  assign \new_[49745]_  = \new_[49744]_  & \new_[49741]_ ;
  assign \new_[49746]_  = \new_[49745]_  & \new_[49738]_ ;
  assign \new_[49750]_  = A167 & A169;
  assign \new_[49751]_  = ~A170 & \new_[49750]_ ;
  assign \new_[49754]_  = A199 & A166;
  assign \new_[49757]_  = ~A233 & A200;
  assign \new_[49758]_  = \new_[49757]_  & \new_[49754]_ ;
  assign \new_[49759]_  = \new_[49758]_  & \new_[49751]_ ;
  assign \new_[49763]_  = A266 & A265;
  assign \new_[49764]_  = ~A234 & \new_[49763]_ ;
  assign \new_[49767]_  = ~A299 & A298;
  assign \new_[49770]_  = A302 & A300;
  assign \new_[49771]_  = \new_[49770]_  & \new_[49767]_ ;
  assign \new_[49772]_  = \new_[49771]_  & \new_[49764]_ ;
  assign \new_[49776]_  = A167 & A169;
  assign \new_[49777]_  = ~A170 & \new_[49776]_ ;
  assign \new_[49780]_  = A199 & A166;
  assign \new_[49783]_  = ~A233 & A200;
  assign \new_[49784]_  = \new_[49783]_  & \new_[49780]_ ;
  assign \new_[49785]_  = \new_[49784]_  & \new_[49777]_ ;
  assign \new_[49789]_  = ~A267 & ~A266;
  assign \new_[49790]_  = ~A234 & \new_[49789]_ ;
  assign \new_[49793]_  = ~A299 & A298;
  assign \new_[49796]_  = A301 & A300;
  assign \new_[49797]_  = \new_[49796]_  & \new_[49793]_ ;
  assign \new_[49798]_  = \new_[49797]_  & \new_[49790]_ ;
  assign \new_[49802]_  = A167 & A169;
  assign \new_[49803]_  = ~A170 & \new_[49802]_ ;
  assign \new_[49806]_  = A199 & A166;
  assign \new_[49809]_  = ~A233 & A200;
  assign \new_[49810]_  = \new_[49809]_  & \new_[49806]_ ;
  assign \new_[49811]_  = \new_[49810]_  & \new_[49803]_ ;
  assign \new_[49815]_  = ~A267 & ~A266;
  assign \new_[49816]_  = ~A234 & \new_[49815]_ ;
  assign \new_[49819]_  = ~A299 & A298;
  assign \new_[49822]_  = A302 & A300;
  assign \new_[49823]_  = \new_[49822]_  & \new_[49819]_ ;
  assign \new_[49824]_  = \new_[49823]_  & \new_[49816]_ ;
  assign \new_[49828]_  = A167 & A169;
  assign \new_[49829]_  = ~A170 & \new_[49828]_ ;
  assign \new_[49832]_  = A199 & A166;
  assign \new_[49835]_  = ~A233 & A200;
  assign \new_[49836]_  = \new_[49835]_  & \new_[49832]_ ;
  assign \new_[49837]_  = \new_[49836]_  & \new_[49829]_ ;
  assign \new_[49841]_  = ~A266 & ~A265;
  assign \new_[49842]_  = ~A234 & \new_[49841]_ ;
  assign \new_[49845]_  = ~A299 & A298;
  assign \new_[49848]_  = A301 & A300;
  assign \new_[49849]_  = \new_[49848]_  & \new_[49845]_ ;
  assign \new_[49850]_  = \new_[49849]_  & \new_[49842]_ ;
  assign \new_[49854]_  = A167 & A169;
  assign \new_[49855]_  = ~A170 & \new_[49854]_ ;
  assign \new_[49858]_  = A199 & A166;
  assign \new_[49861]_  = ~A233 & A200;
  assign \new_[49862]_  = \new_[49861]_  & \new_[49858]_ ;
  assign \new_[49863]_  = \new_[49862]_  & \new_[49855]_ ;
  assign \new_[49867]_  = ~A266 & ~A265;
  assign \new_[49868]_  = ~A234 & \new_[49867]_ ;
  assign \new_[49871]_  = ~A299 & A298;
  assign \new_[49874]_  = A302 & A300;
  assign \new_[49875]_  = \new_[49874]_  & \new_[49871]_ ;
  assign \new_[49876]_  = \new_[49875]_  & \new_[49868]_ ;
  assign \new_[49880]_  = A167 & A169;
  assign \new_[49881]_  = ~A170 & \new_[49880]_ ;
  assign \new_[49884]_  = A199 & A166;
  assign \new_[49887]_  = A232 & A200;
  assign \new_[49888]_  = \new_[49887]_  & \new_[49884]_ ;
  assign \new_[49889]_  = \new_[49888]_  & \new_[49881]_ ;
  assign \new_[49893]_  = A235 & A234;
  assign \new_[49894]_  = ~A233 & \new_[49893]_ ;
  assign \new_[49897]_  = ~A266 & A265;
  assign \new_[49900]_  = A268 & A267;
  assign \new_[49901]_  = \new_[49900]_  & \new_[49897]_ ;
  assign \new_[49902]_  = \new_[49901]_  & \new_[49894]_ ;
  assign \new_[49906]_  = A167 & A169;
  assign \new_[49907]_  = ~A170 & \new_[49906]_ ;
  assign \new_[49910]_  = A199 & A166;
  assign \new_[49913]_  = A232 & A200;
  assign \new_[49914]_  = \new_[49913]_  & \new_[49910]_ ;
  assign \new_[49915]_  = \new_[49914]_  & \new_[49907]_ ;
  assign \new_[49919]_  = A235 & A234;
  assign \new_[49920]_  = ~A233 & \new_[49919]_ ;
  assign \new_[49923]_  = ~A266 & A265;
  assign \new_[49926]_  = A269 & A267;
  assign \new_[49927]_  = \new_[49926]_  & \new_[49923]_ ;
  assign \new_[49928]_  = \new_[49927]_  & \new_[49920]_ ;
  assign \new_[49932]_  = A167 & A169;
  assign \new_[49933]_  = ~A170 & \new_[49932]_ ;
  assign \new_[49936]_  = A199 & A166;
  assign \new_[49939]_  = A232 & A200;
  assign \new_[49940]_  = \new_[49939]_  & \new_[49936]_ ;
  assign \new_[49941]_  = \new_[49940]_  & \new_[49933]_ ;
  assign \new_[49945]_  = A236 & A234;
  assign \new_[49946]_  = ~A233 & \new_[49945]_ ;
  assign \new_[49949]_  = ~A266 & A265;
  assign \new_[49952]_  = A268 & A267;
  assign \new_[49953]_  = \new_[49952]_  & \new_[49949]_ ;
  assign \new_[49954]_  = \new_[49953]_  & \new_[49946]_ ;
  assign \new_[49958]_  = A167 & A169;
  assign \new_[49959]_  = ~A170 & \new_[49958]_ ;
  assign \new_[49962]_  = A199 & A166;
  assign \new_[49965]_  = A232 & A200;
  assign \new_[49966]_  = \new_[49965]_  & \new_[49962]_ ;
  assign \new_[49967]_  = \new_[49966]_  & \new_[49959]_ ;
  assign \new_[49971]_  = A236 & A234;
  assign \new_[49972]_  = ~A233 & \new_[49971]_ ;
  assign \new_[49975]_  = ~A266 & A265;
  assign \new_[49978]_  = A269 & A267;
  assign \new_[49979]_  = \new_[49978]_  & \new_[49975]_ ;
  assign \new_[49980]_  = \new_[49979]_  & \new_[49972]_ ;
  assign \new_[49984]_  = A167 & A169;
  assign \new_[49985]_  = ~A170 & \new_[49984]_ ;
  assign \new_[49988]_  = A199 & A166;
  assign \new_[49991]_  = ~A232 & A200;
  assign \new_[49992]_  = \new_[49991]_  & \new_[49988]_ ;
  assign \new_[49993]_  = \new_[49992]_  & \new_[49985]_ ;
  assign \new_[49997]_  = A266 & A265;
  assign \new_[49998]_  = ~A233 & \new_[49997]_ ;
  assign \new_[50001]_  = ~A299 & A298;
  assign \new_[50004]_  = A301 & A300;
  assign \new_[50005]_  = \new_[50004]_  & \new_[50001]_ ;
  assign \new_[50006]_  = \new_[50005]_  & \new_[49998]_ ;
  assign \new_[50010]_  = A167 & A169;
  assign \new_[50011]_  = ~A170 & \new_[50010]_ ;
  assign \new_[50014]_  = A199 & A166;
  assign \new_[50017]_  = ~A232 & A200;
  assign \new_[50018]_  = \new_[50017]_  & \new_[50014]_ ;
  assign \new_[50019]_  = \new_[50018]_  & \new_[50011]_ ;
  assign \new_[50023]_  = A266 & A265;
  assign \new_[50024]_  = ~A233 & \new_[50023]_ ;
  assign \new_[50027]_  = ~A299 & A298;
  assign \new_[50030]_  = A302 & A300;
  assign \new_[50031]_  = \new_[50030]_  & \new_[50027]_ ;
  assign \new_[50032]_  = \new_[50031]_  & \new_[50024]_ ;
  assign \new_[50036]_  = A167 & A169;
  assign \new_[50037]_  = ~A170 & \new_[50036]_ ;
  assign \new_[50040]_  = A199 & A166;
  assign \new_[50043]_  = ~A232 & A200;
  assign \new_[50044]_  = \new_[50043]_  & \new_[50040]_ ;
  assign \new_[50045]_  = \new_[50044]_  & \new_[50037]_ ;
  assign \new_[50049]_  = ~A267 & ~A266;
  assign \new_[50050]_  = ~A233 & \new_[50049]_ ;
  assign \new_[50053]_  = ~A299 & A298;
  assign \new_[50056]_  = A301 & A300;
  assign \new_[50057]_  = \new_[50056]_  & \new_[50053]_ ;
  assign \new_[50058]_  = \new_[50057]_  & \new_[50050]_ ;
  assign \new_[50062]_  = A167 & A169;
  assign \new_[50063]_  = ~A170 & \new_[50062]_ ;
  assign \new_[50066]_  = A199 & A166;
  assign \new_[50069]_  = ~A232 & A200;
  assign \new_[50070]_  = \new_[50069]_  & \new_[50066]_ ;
  assign \new_[50071]_  = \new_[50070]_  & \new_[50063]_ ;
  assign \new_[50075]_  = ~A267 & ~A266;
  assign \new_[50076]_  = ~A233 & \new_[50075]_ ;
  assign \new_[50079]_  = ~A299 & A298;
  assign \new_[50082]_  = A302 & A300;
  assign \new_[50083]_  = \new_[50082]_  & \new_[50079]_ ;
  assign \new_[50084]_  = \new_[50083]_  & \new_[50076]_ ;
  assign \new_[50088]_  = A167 & A169;
  assign \new_[50089]_  = ~A170 & \new_[50088]_ ;
  assign \new_[50092]_  = A199 & A166;
  assign \new_[50095]_  = ~A232 & A200;
  assign \new_[50096]_  = \new_[50095]_  & \new_[50092]_ ;
  assign \new_[50097]_  = \new_[50096]_  & \new_[50089]_ ;
  assign \new_[50101]_  = ~A266 & ~A265;
  assign \new_[50102]_  = ~A233 & \new_[50101]_ ;
  assign \new_[50105]_  = ~A299 & A298;
  assign \new_[50108]_  = A301 & A300;
  assign \new_[50109]_  = \new_[50108]_  & \new_[50105]_ ;
  assign \new_[50110]_  = \new_[50109]_  & \new_[50102]_ ;
  assign \new_[50114]_  = A167 & A169;
  assign \new_[50115]_  = ~A170 & \new_[50114]_ ;
  assign \new_[50118]_  = A199 & A166;
  assign \new_[50121]_  = ~A232 & A200;
  assign \new_[50122]_  = \new_[50121]_  & \new_[50118]_ ;
  assign \new_[50123]_  = \new_[50122]_  & \new_[50115]_ ;
  assign \new_[50127]_  = ~A266 & ~A265;
  assign \new_[50128]_  = ~A233 & \new_[50127]_ ;
  assign \new_[50131]_  = ~A299 & A298;
  assign \new_[50134]_  = A302 & A300;
  assign \new_[50135]_  = \new_[50134]_  & \new_[50131]_ ;
  assign \new_[50136]_  = \new_[50135]_  & \new_[50128]_ ;
  assign \new_[50140]_  = A167 & A169;
  assign \new_[50141]_  = ~A170 & \new_[50140]_ ;
  assign \new_[50144]_  = ~A200 & A166;
  assign \new_[50147]_  = ~A203 & ~A202;
  assign \new_[50148]_  = \new_[50147]_  & \new_[50144]_ ;
  assign \new_[50149]_  = \new_[50148]_  & \new_[50141]_ ;
  assign \new_[50153]_  = A265 & A233;
  assign \new_[50154]_  = A232 & \new_[50153]_ ;
  assign \new_[50157]_  = ~A269 & ~A268;
  assign \new_[50160]_  = A299 & ~A298;
  assign \new_[50161]_  = \new_[50160]_  & \new_[50157]_ ;
  assign \new_[50162]_  = \new_[50161]_  & \new_[50154]_ ;
  assign \new_[50166]_  = A167 & A169;
  assign \new_[50167]_  = ~A170 & \new_[50166]_ ;
  assign \new_[50170]_  = ~A200 & A166;
  assign \new_[50173]_  = ~A203 & ~A202;
  assign \new_[50174]_  = \new_[50173]_  & \new_[50170]_ ;
  assign \new_[50175]_  = \new_[50174]_  & \new_[50167]_ ;
  assign \new_[50179]_  = ~A236 & ~A235;
  assign \new_[50180]_  = ~A233 & \new_[50179]_ ;
  assign \new_[50183]_  = A266 & A265;
  assign \new_[50186]_  = A299 & ~A298;
  assign \new_[50187]_  = \new_[50186]_  & \new_[50183]_ ;
  assign \new_[50188]_  = \new_[50187]_  & \new_[50180]_ ;
  assign \new_[50192]_  = A167 & A169;
  assign \new_[50193]_  = ~A170 & \new_[50192]_ ;
  assign \new_[50196]_  = ~A200 & A166;
  assign \new_[50199]_  = ~A203 & ~A202;
  assign \new_[50200]_  = \new_[50199]_  & \new_[50196]_ ;
  assign \new_[50201]_  = \new_[50200]_  & \new_[50193]_ ;
  assign \new_[50205]_  = ~A236 & ~A235;
  assign \new_[50206]_  = ~A233 & \new_[50205]_ ;
  assign \new_[50209]_  = ~A267 & ~A266;
  assign \new_[50212]_  = A299 & ~A298;
  assign \new_[50213]_  = \new_[50212]_  & \new_[50209]_ ;
  assign \new_[50214]_  = \new_[50213]_  & \new_[50206]_ ;
  assign \new_[50218]_  = A167 & A169;
  assign \new_[50219]_  = ~A170 & \new_[50218]_ ;
  assign \new_[50222]_  = ~A200 & A166;
  assign \new_[50225]_  = ~A203 & ~A202;
  assign \new_[50226]_  = \new_[50225]_  & \new_[50222]_ ;
  assign \new_[50227]_  = \new_[50226]_  & \new_[50219]_ ;
  assign \new_[50231]_  = ~A236 & ~A235;
  assign \new_[50232]_  = ~A233 & \new_[50231]_ ;
  assign \new_[50235]_  = ~A266 & ~A265;
  assign \new_[50238]_  = A299 & ~A298;
  assign \new_[50239]_  = \new_[50238]_  & \new_[50235]_ ;
  assign \new_[50240]_  = \new_[50239]_  & \new_[50232]_ ;
  assign \new_[50244]_  = A167 & A169;
  assign \new_[50245]_  = ~A170 & \new_[50244]_ ;
  assign \new_[50248]_  = ~A200 & A166;
  assign \new_[50251]_  = ~A203 & ~A202;
  assign \new_[50252]_  = \new_[50251]_  & \new_[50248]_ ;
  assign \new_[50253]_  = \new_[50252]_  & \new_[50245]_ ;
  assign \new_[50257]_  = ~A266 & ~A234;
  assign \new_[50258]_  = ~A233 & \new_[50257]_ ;
  assign \new_[50261]_  = ~A269 & ~A268;
  assign \new_[50264]_  = A299 & ~A298;
  assign \new_[50265]_  = \new_[50264]_  & \new_[50261]_ ;
  assign \new_[50266]_  = \new_[50265]_  & \new_[50258]_ ;
  assign \new_[50270]_  = A167 & A169;
  assign \new_[50271]_  = ~A170 & \new_[50270]_ ;
  assign \new_[50274]_  = ~A200 & A166;
  assign \new_[50277]_  = ~A203 & ~A202;
  assign \new_[50278]_  = \new_[50277]_  & \new_[50274]_ ;
  assign \new_[50279]_  = \new_[50278]_  & \new_[50271]_ ;
  assign \new_[50283]_  = A234 & ~A233;
  assign \new_[50284]_  = A232 & \new_[50283]_ ;
  assign \new_[50287]_  = A298 & A235;
  assign \new_[50290]_  = ~A302 & ~A301;
  assign \new_[50291]_  = \new_[50290]_  & \new_[50287]_ ;
  assign \new_[50292]_  = \new_[50291]_  & \new_[50284]_ ;
  assign \new_[50296]_  = A167 & A169;
  assign \new_[50297]_  = ~A170 & \new_[50296]_ ;
  assign \new_[50300]_  = ~A200 & A166;
  assign \new_[50303]_  = ~A203 & ~A202;
  assign \new_[50304]_  = \new_[50303]_  & \new_[50300]_ ;
  assign \new_[50305]_  = \new_[50304]_  & \new_[50297]_ ;
  assign \new_[50309]_  = A234 & ~A233;
  assign \new_[50310]_  = A232 & \new_[50309]_ ;
  assign \new_[50313]_  = A298 & A236;
  assign \new_[50316]_  = ~A302 & ~A301;
  assign \new_[50317]_  = \new_[50316]_  & \new_[50313]_ ;
  assign \new_[50318]_  = \new_[50317]_  & \new_[50310]_ ;
  assign \new_[50322]_  = A167 & A169;
  assign \new_[50323]_  = ~A170 & \new_[50322]_ ;
  assign \new_[50326]_  = ~A200 & A166;
  assign \new_[50329]_  = ~A203 & ~A202;
  assign \new_[50330]_  = \new_[50329]_  & \new_[50326]_ ;
  assign \new_[50331]_  = \new_[50330]_  & \new_[50323]_ ;
  assign \new_[50335]_  = ~A266 & ~A233;
  assign \new_[50336]_  = ~A232 & \new_[50335]_ ;
  assign \new_[50339]_  = ~A269 & ~A268;
  assign \new_[50342]_  = A299 & ~A298;
  assign \new_[50343]_  = \new_[50342]_  & \new_[50339]_ ;
  assign \new_[50344]_  = \new_[50343]_  & \new_[50336]_ ;
  assign \new_[50348]_  = A167 & A169;
  assign \new_[50349]_  = ~A170 & \new_[50348]_ ;
  assign \new_[50352]_  = ~A200 & A166;
  assign \new_[50355]_  = A232 & ~A201;
  assign \new_[50356]_  = \new_[50355]_  & \new_[50352]_ ;
  assign \new_[50357]_  = \new_[50356]_  & \new_[50349]_ ;
  assign \new_[50361]_  = ~A267 & A265;
  assign \new_[50362]_  = A233 & \new_[50361]_ ;
  assign \new_[50365]_  = ~A299 & A298;
  assign \new_[50368]_  = A301 & A300;
  assign \new_[50369]_  = \new_[50368]_  & \new_[50365]_ ;
  assign \new_[50370]_  = \new_[50369]_  & \new_[50362]_ ;
  assign \new_[50374]_  = A167 & A169;
  assign \new_[50375]_  = ~A170 & \new_[50374]_ ;
  assign \new_[50378]_  = ~A200 & A166;
  assign \new_[50381]_  = A232 & ~A201;
  assign \new_[50382]_  = \new_[50381]_  & \new_[50378]_ ;
  assign \new_[50383]_  = \new_[50382]_  & \new_[50375]_ ;
  assign \new_[50387]_  = ~A267 & A265;
  assign \new_[50388]_  = A233 & \new_[50387]_ ;
  assign \new_[50391]_  = ~A299 & A298;
  assign \new_[50394]_  = A302 & A300;
  assign \new_[50395]_  = \new_[50394]_  & \new_[50391]_ ;
  assign \new_[50396]_  = \new_[50395]_  & \new_[50388]_ ;
  assign \new_[50400]_  = A167 & A169;
  assign \new_[50401]_  = ~A170 & \new_[50400]_ ;
  assign \new_[50404]_  = ~A200 & A166;
  assign \new_[50407]_  = A232 & ~A201;
  assign \new_[50408]_  = \new_[50407]_  & \new_[50404]_ ;
  assign \new_[50409]_  = \new_[50408]_  & \new_[50401]_ ;
  assign \new_[50413]_  = A266 & A265;
  assign \new_[50414]_  = A233 & \new_[50413]_ ;
  assign \new_[50417]_  = ~A299 & A298;
  assign \new_[50420]_  = A301 & A300;
  assign \new_[50421]_  = \new_[50420]_  & \new_[50417]_ ;
  assign \new_[50422]_  = \new_[50421]_  & \new_[50414]_ ;
  assign \new_[50426]_  = A167 & A169;
  assign \new_[50427]_  = ~A170 & \new_[50426]_ ;
  assign \new_[50430]_  = ~A200 & A166;
  assign \new_[50433]_  = A232 & ~A201;
  assign \new_[50434]_  = \new_[50433]_  & \new_[50430]_ ;
  assign \new_[50435]_  = \new_[50434]_  & \new_[50427]_ ;
  assign \new_[50439]_  = A266 & A265;
  assign \new_[50440]_  = A233 & \new_[50439]_ ;
  assign \new_[50443]_  = ~A299 & A298;
  assign \new_[50446]_  = A302 & A300;
  assign \new_[50447]_  = \new_[50446]_  & \new_[50443]_ ;
  assign \new_[50448]_  = \new_[50447]_  & \new_[50440]_ ;
  assign \new_[50452]_  = A167 & A169;
  assign \new_[50453]_  = ~A170 & \new_[50452]_ ;
  assign \new_[50456]_  = ~A200 & A166;
  assign \new_[50459]_  = A232 & ~A201;
  assign \new_[50460]_  = \new_[50459]_  & \new_[50456]_ ;
  assign \new_[50461]_  = \new_[50460]_  & \new_[50453]_ ;
  assign \new_[50465]_  = ~A266 & ~A265;
  assign \new_[50466]_  = A233 & \new_[50465]_ ;
  assign \new_[50469]_  = ~A299 & A298;
  assign \new_[50472]_  = A301 & A300;
  assign \new_[50473]_  = \new_[50472]_  & \new_[50469]_ ;
  assign \new_[50474]_  = \new_[50473]_  & \new_[50466]_ ;
  assign \new_[50478]_  = A167 & A169;
  assign \new_[50479]_  = ~A170 & \new_[50478]_ ;
  assign \new_[50482]_  = ~A200 & A166;
  assign \new_[50485]_  = A232 & ~A201;
  assign \new_[50486]_  = \new_[50485]_  & \new_[50482]_ ;
  assign \new_[50487]_  = \new_[50486]_  & \new_[50479]_ ;
  assign \new_[50491]_  = ~A266 & ~A265;
  assign \new_[50492]_  = A233 & \new_[50491]_ ;
  assign \new_[50495]_  = ~A299 & A298;
  assign \new_[50498]_  = A302 & A300;
  assign \new_[50499]_  = \new_[50498]_  & \new_[50495]_ ;
  assign \new_[50500]_  = \new_[50499]_  & \new_[50492]_ ;
  assign \new_[50504]_  = A167 & A169;
  assign \new_[50505]_  = ~A170 & \new_[50504]_ ;
  assign \new_[50508]_  = ~A200 & A166;
  assign \new_[50511]_  = ~A233 & ~A201;
  assign \new_[50512]_  = \new_[50511]_  & \new_[50508]_ ;
  assign \new_[50513]_  = \new_[50512]_  & \new_[50505]_ ;
  assign \new_[50517]_  = ~A266 & ~A236;
  assign \new_[50518]_  = ~A235 & \new_[50517]_ ;
  assign \new_[50521]_  = ~A269 & ~A268;
  assign \new_[50524]_  = A299 & ~A298;
  assign \new_[50525]_  = \new_[50524]_  & \new_[50521]_ ;
  assign \new_[50526]_  = \new_[50525]_  & \new_[50518]_ ;
  assign \new_[50530]_  = A167 & A169;
  assign \new_[50531]_  = ~A170 & \new_[50530]_ ;
  assign \new_[50534]_  = ~A200 & A166;
  assign \new_[50537]_  = ~A233 & ~A201;
  assign \new_[50538]_  = \new_[50537]_  & \new_[50534]_ ;
  assign \new_[50539]_  = \new_[50538]_  & \new_[50531]_ ;
  assign \new_[50543]_  = A266 & A265;
  assign \new_[50544]_  = ~A234 & \new_[50543]_ ;
  assign \new_[50547]_  = ~A299 & A298;
  assign \new_[50550]_  = A301 & A300;
  assign \new_[50551]_  = \new_[50550]_  & \new_[50547]_ ;
  assign \new_[50552]_  = \new_[50551]_  & \new_[50544]_ ;
  assign \new_[50556]_  = A167 & A169;
  assign \new_[50557]_  = ~A170 & \new_[50556]_ ;
  assign \new_[50560]_  = ~A200 & A166;
  assign \new_[50563]_  = ~A233 & ~A201;
  assign \new_[50564]_  = \new_[50563]_  & \new_[50560]_ ;
  assign \new_[50565]_  = \new_[50564]_  & \new_[50557]_ ;
  assign \new_[50569]_  = A266 & A265;
  assign \new_[50570]_  = ~A234 & \new_[50569]_ ;
  assign \new_[50573]_  = ~A299 & A298;
  assign \new_[50576]_  = A302 & A300;
  assign \new_[50577]_  = \new_[50576]_  & \new_[50573]_ ;
  assign \new_[50578]_  = \new_[50577]_  & \new_[50570]_ ;
  assign \new_[50582]_  = A167 & A169;
  assign \new_[50583]_  = ~A170 & \new_[50582]_ ;
  assign \new_[50586]_  = ~A200 & A166;
  assign \new_[50589]_  = ~A233 & ~A201;
  assign \new_[50590]_  = \new_[50589]_  & \new_[50586]_ ;
  assign \new_[50591]_  = \new_[50590]_  & \new_[50583]_ ;
  assign \new_[50595]_  = ~A267 & ~A266;
  assign \new_[50596]_  = ~A234 & \new_[50595]_ ;
  assign \new_[50599]_  = ~A299 & A298;
  assign \new_[50602]_  = A301 & A300;
  assign \new_[50603]_  = \new_[50602]_  & \new_[50599]_ ;
  assign \new_[50604]_  = \new_[50603]_  & \new_[50596]_ ;
  assign \new_[50608]_  = A167 & A169;
  assign \new_[50609]_  = ~A170 & \new_[50608]_ ;
  assign \new_[50612]_  = ~A200 & A166;
  assign \new_[50615]_  = ~A233 & ~A201;
  assign \new_[50616]_  = \new_[50615]_  & \new_[50612]_ ;
  assign \new_[50617]_  = \new_[50616]_  & \new_[50609]_ ;
  assign \new_[50621]_  = ~A267 & ~A266;
  assign \new_[50622]_  = ~A234 & \new_[50621]_ ;
  assign \new_[50625]_  = ~A299 & A298;
  assign \new_[50628]_  = A302 & A300;
  assign \new_[50629]_  = \new_[50628]_  & \new_[50625]_ ;
  assign \new_[50630]_  = \new_[50629]_  & \new_[50622]_ ;
  assign \new_[50634]_  = A167 & A169;
  assign \new_[50635]_  = ~A170 & \new_[50634]_ ;
  assign \new_[50638]_  = ~A200 & A166;
  assign \new_[50641]_  = ~A233 & ~A201;
  assign \new_[50642]_  = \new_[50641]_  & \new_[50638]_ ;
  assign \new_[50643]_  = \new_[50642]_  & \new_[50635]_ ;
  assign \new_[50647]_  = ~A266 & ~A265;
  assign \new_[50648]_  = ~A234 & \new_[50647]_ ;
  assign \new_[50651]_  = ~A299 & A298;
  assign \new_[50654]_  = A301 & A300;
  assign \new_[50655]_  = \new_[50654]_  & \new_[50651]_ ;
  assign \new_[50656]_  = \new_[50655]_  & \new_[50648]_ ;
  assign \new_[50660]_  = A167 & A169;
  assign \new_[50661]_  = ~A170 & \new_[50660]_ ;
  assign \new_[50664]_  = ~A200 & A166;
  assign \new_[50667]_  = ~A233 & ~A201;
  assign \new_[50668]_  = \new_[50667]_  & \new_[50664]_ ;
  assign \new_[50669]_  = \new_[50668]_  & \new_[50661]_ ;
  assign \new_[50673]_  = ~A266 & ~A265;
  assign \new_[50674]_  = ~A234 & \new_[50673]_ ;
  assign \new_[50677]_  = ~A299 & A298;
  assign \new_[50680]_  = A302 & A300;
  assign \new_[50681]_  = \new_[50680]_  & \new_[50677]_ ;
  assign \new_[50682]_  = \new_[50681]_  & \new_[50674]_ ;
  assign \new_[50686]_  = A167 & A169;
  assign \new_[50687]_  = ~A170 & \new_[50686]_ ;
  assign \new_[50690]_  = ~A200 & A166;
  assign \new_[50693]_  = A232 & ~A201;
  assign \new_[50694]_  = \new_[50693]_  & \new_[50690]_ ;
  assign \new_[50695]_  = \new_[50694]_  & \new_[50687]_ ;
  assign \new_[50699]_  = A235 & A234;
  assign \new_[50700]_  = ~A233 & \new_[50699]_ ;
  assign \new_[50703]_  = ~A266 & A265;
  assign \new_[50706]_  = A268 & A267;
  assign \new_[50707]_  = \new_[50706]_  & \new_[50703]_ ;
  assign \new_[50708]_  = \new_[50707]_  & \new_[50700]_ ;
  assign \new_[50712]_  = A167 & A169;
  assign \new_[50713]_  = ~A170 & \new_[50712]_ ;
  assign \new_[50716]_  = ~A200 & A166;
  assign \new_[50719]_  = A232 & ~A201;
  assign \new_[50720]_  = \new_[50719]_  & \new_[50716]_ ;
  assign \new_[50721]_  = \new_[50720]_  & \new_[50713]_ ;
  assign \new_[50725]_  = A235 & A234;
  assign \new_[50726]_  = ~A233 & \new_[50725]_ ;
  assign \new_[50729]_  = ~A266 & A265;
  assign \new_[50732]_  = A269 & A267;
  assign \new_[50733]_  = \new_[50732]_  & \new_[50729]_ ;
  assign \new_[50734]_  = \new_[50733]_  & \new_[50726]_ ;
  assign \new_[50738]_  = A167 & A169;
  assign \new_[50739]_  = ~A170 & \new_[50738]_ ;
  assign \new_[50742]_  = ~A200 & A166;
  assign \new_[50745]_  = A232 & ~A201;
  assign \new_[50746]_  = \new_[50745]_  & \new_[50742]_ ;
  assign \new_[50747]_  = \new_[50746]_  & \new_[50739]_ ;
  assign \new_[50751]_  = A236 & A234;
  assign \new_[50752]_  = ~A233 & \new_[50751]_ ;
  assign \new_[50755]_  = ~A266 & A265;
  assign \new_[50758]_  = A268 & A267;
  assign \new_[50759]_  = \new_[50758]_  & \new_[50755]_ ;
  assign \new_[50760]_  = \new_[50759]_  & \new_[50752]_ ;
  assign \new_[50764]_  = A167 & A169;
  assign \new_[50765]_  = ~A170 & \new_[50764]_ ;
  assign \new_[50768]_  = ~A200 & A166;
  assign \new_[50771]_  = A232 & ~A201;
  assign \new_[50772]_  = \new_[50771]_  & \new_[50768]_ ;
  assign \new_[50773]_  = \new_[50772]_  & \new_[50765]_ ;
  assign \new_[50777]_  = A236 & A234;
  assign \new_[50778]_  = ~A233 & \new_[50777]_ ;
  assign \new_[50781]_  = ~A266 & A265;
  assign \new_[50784]_  = A269 & A267;
  assign \new_[50785]_  = \new_[50784]_  & \new_[50781]_ ;
  assign \new_[50786]_  = \new_[50785]_  & \new_[50778]_ ;
  assign \new_[50790]_  = A167 & A169;
  assign \new_[50791]_  = ~A170 & \new_[50790]_ ;
  assign \new_[50794]_  = ~A200 & A166;
  assign \new_[50797]_  = ~A232 & ~A201;
  assign \new_[50798]_  = \new_[50797]_  & \new_[50794]_ ;
  assign \new_[50799]_  = \new_[50798]_  & \new_[50791]_ ;
  assign \new_[50803]_  = A266 & A265;
  assign \new_[50804]_  = ~A233 & \new_[50803]_ ;
  assign \new_[50807]_  = ~A299 & A298;
  assign \new_[50810]_  = A301 & A300;
  assign \new_[50811]_  = \new_[50810]_  & \new_[50807]_ ;
  assign \new_[50812]_  = \new_[50811]_  & \new_[50804]_ ;
  assign \new_[50816]_  = A167 & A169;
  assign \new_[50817]_  = ~A170 & \new_[50816]_ ;
  assign \new_[50820]_  = ~A200 & A166;
  assign \new_[50823]_  = ~A232 & ~A201;
  assign \new_[50824]_  = \new_[50823]_  & \new_[50820]_ ;
  assign \new_[50825]_  = \new_[50824]_  & \new_[50817]_ ;
  assign \new_[50829]_  = A266 & A265;
  assign \new_[50830]_  = ~A233 & \new_[50829]_ ;
  assign \new_[50833]_  = ~A299 & A298;
  assign \new_[50836]_  = A302 & A300;
  assign \new_[50837]_  = \new_[50836]_  & \new_[50833]_ ;
  assign \new_[50838]_  = \new_[50837]_  & \new_[50830]_ ;
  assign \new_[50842]_  = A167 & A169;
  assign \new_[50843]_  = ~A170 & \new_[50842]_ ;
  assign \new_[50846]_  = ~A200 & A166;
  assign \new_[50849]_  = ~A232 & ~A201;
  assign \new_[50850]_  = \new_[50849]_  & \new_[50846]_ ;
  assign \new_[50851]_  = \new_[50850]_  & \new_[50843]_ ;
  assign \new_[50855]_  = ~A267 & ~A266;
  assign \new_[50856]_  = ~A233 & \new_[50855]_ ;
  assign \new_[50859]_  = ~A299 & A298;
  assign \new_[50862]_  = A301 & A300;
  assign \new_[50863]_  = \new_[50862]_  & \new_[50859]_ ;
  assign \new_[50864]_  = \new_[50863]_  & \new_[50856]_ ;
  assign \new_[50868]_  = A167 & A169;
  assign \new_[50869]_  = ~A170 & \new_[50868]_ ;
  assign \new_[50872]_  = ~A200 & A166;
  assign \new_[50875]_  = ~A232 & ~A201;
  assign \new_[50876]_  = \new_[50875]_  & \new_[50872]_ ;
  assign \new_[50877]_  = \new_[50876]_  & \new_[50869]_ ;
  assign \new_[50881]_  = ~A267 & ~A266;
  assign \new_[50882]_  = ~A233 & \new_[50881]_ ;
  assign \new_[50885]_  = ~A299 & A298;
  assign \new_[50888]_  = A302 & A300;
  assign \new_[50889]_  = \new_[50888]_  & \new_[50885]_ ;
  assign \new_[50890]_  = \new_[50889]_  & \new_[50882]_ ;
  assign \new_[50894]_  = A167 & A169;
  assign \new_[50895]_  = ~A170 & \new_[50894]_ ;
  assign \new_[50898]_  = ~A200 & A166;
  assign \new_[50901]_  = ~A232 & ~A201;
  assign \new_[50902]_  = \new_[50901]_  & \new_[50898]_ ;
  assign \new_[50903]_  = \new_[50902]_  & \new_[50895]_ ;
  assign \new_[50907]_  = ~A266 & ~A265;
  assign \new_[50908]_  = ~A233 & \new_[50907]_ ;
  assign \new_[50911]_  = ~A299 & A298;
  assign \new_[50914]_  = A301 & A300;
  assign \new_[50915]_  = \new_[50914]_  & \new_[50911]_ ;
  assign \new_[50916]_  = \new_[50915]_  & \new_[50908]_ ;
  assign \new_[50920]_  = A167 & A169;
  assign \new_[50921]_  = ~A170 & \new_[50920]_ ;
  assign \new_[50924]_  = ~A200 & A166;
  assign \new_[50927]_  = ~A232 & ~A201;
  assign \new_[50928]_  = \new_[50927]_  & \new_[50924]_ ;
  assign \new_[50929]_  = \new_[50928]_  & \new_[50921]_ ;
  assign \new_[50933]_  = ~A266 & ~A265;
  assign \new_[50934]_  = ~A233 & \new_[50933]_ ;
  assign \new_[50937]_  = ~A299 & A298;
  assign \new_[50940]_  = A302 & A300;
  assign \new_[50941]_  = \new_[50940]_  & \new_[50937]_ ;
  assign \new_[50942]_  = \new_[50941]_  & \new_[50934]_ ;
  assign \new_[50946]_  = A167 & A169;
  assign \new_[50947]_  = ~A170 & \new_[50946]_ ;
  assign \new_[50950]_  = ~A199 & A166;
  assign \new_[50953]_  = A232 & ~A200;
  assign \new_[50954]_  = \new_[50953]_  & \new_[50950]_ ;
  assign \new_[50955]_  = \new_[50954]_  & \new_[50947]_ ;
  assign \new_[50959]_  = ~A267 & A265;
  assign \new_[50960]_  = A233 & \new_[50959]_ ;
  assign \new_[50963]_  = ~A299 & A298;
  assign \new_[50966]_  = A301 & A300;
  assign \new_[50967]_  = \new_[50966]_  & \new_[50963]_ ;
  assign \new_[50968]_  = \new_[50967]_  & \new_[50960]_ ;
  assign \new_[50972]_  = A167 & A169;
  assign \new_[50973]_  = ~A170 & \new_[50972]_ ;
  assign \new_[50976]_  = ~A199 & A166;
  assign \new_[50979]_  = A232 & ~A200;
  assign \new_[50980]_  = \new_[50979]_  & \new_[50976]_ ;
  assign \new_[50981]_  = \new_[50980]_  & \new_[50973]_ ;
  assign \new_[50985]_  = ~A267 & A265;
  assign \new_[50986]_  = A233 & \new_[50985]_ ;
  assign \new_[50989]_  = ~A299 & A298;
  assign \new_[50992]_  = A302 & A300;
  assign \new_[50993]_  = \new_[50992]_  & \new_[50989]_ ;
  assign \new_[50994]_  = \new_[50993]_  & \new_[50986]_ ;
  assign \new_[50998]_  = A167 & A169;
  assign \new_[50999]_  = ~A170 & \new_[50998]_ ;
  assign \new_[51002]_  = ~A199 & A166;
  assign \new_[51005]_  = A232 & ~A200;
  assign \new_[51006]_  = \new_[51005]_  & \new_[51002]_ ;
  assign \new_[51007]_  = \new_[51006]_  & \new_[50999]_ ;
  assign \new_[51011]_  = A266 & A265;
  assign \new_[51012]_  = A233 & \new_[51011]_ ;
  assign \new_[51015]_  = ~A299 & A298;
  assign \new_[51018]_  = A301 & A300;
  assign \new_[51019]_  = \new_[51018]_  & \new_[51015]_ ;
  assign \new_[51020]_  = \new_[51019]_  & \new_[51012]_ ;
  assign \new_[51024]_  = A167 & A169;
  assign \new_[51025]_  = ~A170 & \new_[51024]_ ;
  assign \new_[51028]_  = ~A199 & A166;
  assign \new_[51031]_  = A232 & ~A200;
  assign \new_[51032]_  = \new_[51031]_  & \new_[51028]_ ;
  assign \new_[51033]_  = \new_[51032]_  & \new_[51025]_ ;
  assign \new_[51037]_  = A266 & A265;
  assign \new_[51038]_  = A233 & \new_[51037]_ ;
  assign \new_[51041]_  = ~A299 & A298;
  assign \new_[51044]_  = A302 & A300;
  assign \new_[51045]_  = \new_[51044]_  & \new_[51041]_ ;
  assign \new_[51046]_  = \new_[51045]_  & \new_[51038]_ ;
  assign \new_[51050]_  = A167 & A169;
  assign \new_[51051]_  = ~A170 & \new_[51050]_ ;
  assign \new_[51054]_  = ~A199 & A166;
  assign \new_[51057]_  = A232 & ~A200;
  assign \new_[51058]_  = \new_[51057]_  & \new_[51054]_ ;
  assign \new_[51059]_  = \new_[51058]_  & \new_[51051]_ ;
  assign \new_[51063]_  = ~A266 & ~A265;
  assign \new_[51064]_  = A233 & \new_[51063]_ ;
  assign \new_[51067]_  = ~A299 & A298;
  assign \new_[51070]_  = A301 & A300;
  assign \new_[51071]_  = \new_[51070]_  & \new_[51067]_ ;
  assign \new_[51072]_  = \new_[51071]_  & \new_[51064]_ ;
  assign \new_[51076]_  = A167 & A169;
  assign \new_[51077]_  = ~A170 & \new_[51076]_ ;
  assign \new_[51080]_  = ~A199 & A166;
  assign \new_[51083]_  = A232 & ~A200;
  assign \new_[51084]_  = \new_[51083]_  & \new_[51080]_ ;
  assign \new_[51085]_  = \new_[51084]_  & \new_[51077]_ ;
  assign \new_[51089]_  = ~A266 & ~A265;
  assign \new_[51090]_  = A233 & \new_[51089]_ ;
  assign \new_[51093]_  = ~A299 & A298;
  assign \new_[51096]_  = A302 & A300;
  assign \new_[51097]_  = \new_[51096]_  & \new_[51093]_ ;
  assign \new_[51098]_  = \new_[51097]_  & \new_[51090]_ ;
  assign \new_[51102]_  = A167 & A169;
  assign \new_[51103]_  = ~A170 & \new_[51102]_ ;
  assign \new_[51106]_  = ~A199 & A166;
  assign \new_[51109]_  = ~A233 & ~A200;
  assign \new_[51110]_  = \new_[51109]_  & \new_[51106]_ ;
  assign \new_[51111]_  = \new_[51110]_  & \new_[51103]_ ;
  assign \new_[51115]_  = ~A266 & ~A236;
  assign \new_[51116]_  = ~A235 & \new_[51115]_ ;
  assign \new_[51119]_  = ~A269 & ~A268;
  assign \new_[51122]_  = A299 & ~A298;
  assign \new_[51123]_  = \new_[51122]_  & \new_[51119]_ ;
  assign \new_[51124]_  = \new_[51123]_  & \new_[51116]_ ;
  assign \new_[51128]_  = A167 & A169;
  assign \new_[51129]_  = ~A170 & \new_[51128]_ ;
  assign \new_[51132]_  = ~A199 & A166;
  assign \new_[51135]_  = ~A233 & ~A200;
  assign \new_[51136]_  = \new_[51135]_  & \new_[51132]_ ;
  assign \new_[51137]_  = \new_[51136]_  & \new_[51129]_ ;
  assign \new_[51141]_  = A266 & A265;
  assign \new_[51142]_  = ~A234 & \new_[51141]_ ;
  assign \new_[51145]_  = ~A299 & A298;
  assign \new_[51148]_  = A301 & A300;
  assign \new_[51149]_  = \new_[51148]_  & \new_[51145]_ ;
  assign \new_[51150]_  = \new_[51149]_  & \new_[51142]_ ;
  assign \new_[51154]_  = A167 & A169;
  assign \new_[51155]_  = ~A170 & \new_[51154]_ ;
  assign \new_[51158]_  = ~A199 & A166;
  assign \new_[51161]_  = ~A233 & ~A200;
  assign \new_[51162]_  = \new_[51161]_  & \new_[51158]_ ;
  assign \new_[51163]_  = \new_[51162]_  & \new_[51155]_ ;
  assign \new_[51167]_  = A266 & A265;
  assign \new_[51168]_  = ~A234 & \new_[51167]_ ;
  assign \new_[51171]_  = ~A299 & A298;
  assign \new_[51174]_  = A302 & A300;
  assign \new_[51175]_  = \new_[51174]_  & \new_[51171]_ ;
  assign \new_[51176]_  = \new_[51175]_  & \new_[51168]_ ;
  assign \new_[51180]_  = A167 & A169;
  assign \new_[51181]_  = ~A170 & \new_[51180]_ ;
  assign \new_[51184]_  = ~A199 & A166;
  assign \new_[51187]_  = ~A233 & ~A200;
  assign \new_[51188]_  = \new_[51187]_  & \new_[51184]_ ;
  assign \new_[51189]_  = \new_[51188]_  & \new_[51181]_ ;
  assign \new_[51193]_  = ~A267 & ~A266;
  assign \new_[51194]_  = ~A234 & \new_[51193]_ ;
  assign \new_[51197]_  = ~A299 & A298;
  assign \new_[51200]_  = A301 & A300;
  assign \new_[51201]_  = \new_[51200]_  & \new_[51197]_ ;
  assign \new_[51202]_  = \new_[51201]_  & \new_[51194]_ ;
  assign \new_[51206]_  = A167 & A169;
  assign \new_[51207]_  = ~A170 & \new_[51206]_ ;
  assign \new_[51210]_  = ~A199 & A166;
  assign \new_[51213]_  = ~A233 & ~A200;
  assign \new_[51214]_  = \new_[51213]_  & \new_[51210]_ ;
  assign \new_[51215]_  = \new_[51214]_  & \new_[51207]_ ;
  assign \new_[51219]_  = ~A267 & ~A266;
  assign \new_[51220]_  = ~A234 & \new_[51219]_ ;
  assign \new_[51223]_  = ~A299 & A298;
  assign \new_[51226]_  = A302 & A300;
  assign \new_[51227]_  = \new_[51226]_  & \new_[51223]_ ;
  assign \new_[51228]_  = \new_[51227]_  & \new_[51220]_ ;
  assign \new_[51232]_  = A167 & A169;
  assign \new_[51233]_  = ~A170 & \new_[51232]_ ;
  assign \new_[51236]_  = ~A199 & A166;
  assign \new_[51239]_  = ~A233 & ~A200;
  assign \new_[51240]_  = \new_[51239]_  & \new_[51236]_ ;
  assign \new_[51241]_  = \new_[51240]_  & \new_[51233]_ ;
  assign \new_[51245]_  = ~A266 & ~A265;
  assign \new_[51246]_  = ~A234 & \new_[51245]_ ;
  assign \new_[51249]_  = ~A299 & A298;
  assign \new_[51252]_  = A301 & A300;
  assign \new_[51253]_  = \new_[51252]_  & \new_[51249]_ ;
  assign \new_[51254]_  = \new_[51253]_  & \new_[51246]_ ;
  assign \new_[51258]_  = A167 & A169;
  assign \new_[51259]_  = ~A170 & \new_[51258]_ ;
  assign \new_[51262]_  = ~A199 & A166;
  assign \new_[51265]_  = ~A233 & ~A200;
  assign \new_[51266]_  = \new_[51265]_  & \new_[51262]_ ;
  assign \new_[51267]_  = \new_[51266]_  & \new_[51259]_ ;
  assign \new_[51271]_  = ~A266 & ~A265;
  assign \new_[51272]_  = ~A234 & \new_[51271]_ ;
  assign \new_[51275]_  = ~A299 & A298;
  assign \new_[51278]_  = A302 & A300;
  assign \new_[51279]_  = \new_[51278]_  & \new_[51275]_ ;
  assign \new_[51280]_  = \new_[51279]_  & \new_[51272]_ ;
  assign \new_[51284]_  = A167 & A169;
  assign \new_[51285]_  = ~A170 & \new_[51284]_ ;
  assign \new_[51288]_  = ~A199 & A166;
  assign \new_[51291]_  = A232 & ~A200;
  assign \new_[51292]_  = \new_[51291]_  & \new_[51288]_ ;
  assign \new_[51293]_  = \new_[51292]_  & \new_[51285]_ ;
  assign \new_[51297]_  = A235 & A234;
  assign \new_[51298]_  = ~A233 & \new_[51297]_ ;
  assign \new_[51301]_  = ~A266 & A265;
  assign \new_[51304]_  = A268 & A267;
  assign \new_[51305]_  = \new_[51304]_  & \new_[51301]_ ;
  assign \new_[51306]_  = \new_[51305]_  & \new_[51298]_ ;
  assign \new_[51310]_  = A167 & A169;
  assign \new_[51311]_  = ~A170 & \new_[51310]_ ;
  assign \new_[51314]_  = ~A199 & A166;
  assign \new_[51317]_  = A232 & ~A200;
  assign \new_[51318]_  = \new_[51317]_  & \new_[51314]_ ;
  assign \new_[51319]_  = \new_[51318]_  & \new_[51311]_ ;
  assign \new_[51323]_  = A235 & A234;
  assign \new_[51324]_  = ~A233 & \new_[51323]_ ;
  assign \new_[51327]_  = ~A266 & A265;
  assign \new_[51330]_  = A269 & A267;
  assign \new_[51331]_  = \new_[51330]_  & \new_[51327]_ ;
  assign \new_[51332]_  = \new_[51331]_  & \new_[51324]_ ;
  assign \new_[51336]_  = A167 & A169;
  assign \new_[51337]_  = ~A170 & \new_[51336]_ ;
  assign \new_[51340]_  = ~A199 & A166;
  assign \new_[51343]_  = A232 & ~A200;
  assign \new_[51344]_  = \new_[51343]_  & \new_[51340]_ ;
  assign \new_[51345]_  = \new_[51344]_  & \new_[51337]_ ;
  assign \new_[51349]_  = A236 & A234;
  assign \new_[51350]_  = ~A233 & \new_[51349]_ ;
  assign \new_[51353]_  = ~A266 & A265;
  assign \new_[51356]_  = A268 & A267;
  assign \new_[51357]_  = \new_[51356]_  & \new_[51353]_ ;
  assign \new_[51358]_  = \new_[51357]_  & \new_[51350]_ ;
  assign \new_[51362]_  = A167 & A169;
  assign \new_[51363]_  = ~A170 & \new_[51362]_ ;
  assign \new_[51366]_  = ~A199 & A166;
  assign \new_[51369]_  = A232 & ~A200;
  assign \new_[51370]_  = \new_[51369]_  & \new_[51366]_ ;
  assign \new_[51371]_  = \new_[51370]_  & \new_[51363]_ ;
  assign \new_[51375]_  = A236 & A234;
  assign \new_[51376]_  = ~A233 & \new_[51375]_ ;
  assign \new_[51379]_  = ~A266 & A265;
  assign \new_[51382]_  = A269 & A267;
  assign \new_[51383]_  = \new_[51382]_  & \new_[51379]_ ;
  assign \new_[51384]_  = \new_[51383]_  & \new_[51376]_ ;
  assign \new_[51388]_  = A167 & A169;
  assign \new_[51389]_  = ~A170 & \new_[51388]_ ;
  assign \new_[51392]_  = ~A199 & A166;
  assign \new_[51395]_  = ~A232 & ~A200;
  assign \new_[51396]_  = \new_[51395]_  & \new_[51392]_ ;
  assign \new_[51397]_  = \new_[51396]_  & \new_[51389]_ ;
  assign \new_[51401]_  = A266 & A265;
  assign \new_[51402]_  = ~A233 & \new_[51401]_ ;
  assign \new_[51405]_  = ~A299 & A298;
  assign \new_[51408]_  = A301 & A300;
  assign \new_[51409]_  = \new_[51408]_  & \new_[51405]_ ;
  assign \new_[51410]_  = \new_[51409]_  & \new_[51402]_ ;
  assign \new_[51414]_  = A167 & A169;
  assign \new_[51415]_  = ~A170 & \new_[51414]_ ;
  assign \new_[51418]_  = ~A199 & A166;
  assign \new_[51421]_  = ~A232 & ~A200;
  assign \new_[51422]_  = \new_[51421]_  & \new_[51418]_ ;
  assign \new_[51423]_  = \new_[51422]_  & \new_[51415]_ ;
  assign \new_[51427]_  = A266 & A265;
  assign \new_[51428]_  = ~A233 & \new_[51427]_ ;
  assign \new_[51431]_  = ~A299 & A298;
  assign \new_[51434]_  = A302 & A300;
  assign \new_[51435]_  = \new_[51434]_  & \new_[51431]_ ;
  assign \new_[51436]_  = \new_[51435]_  & \new_[51428]_ ;
  assign \new_[51440]_  = A167 & A169;
  assign \new_[51441]_  = ~A170 & \new_[51440]_ ;
  assign \new_[51444]_  = ~A199 & A166;
  assign \new_[51447]_  = ~A232 & ~A200;
  assign \new_[51448]_  = \new_[51447]_  & \new_[51444]_ ;
  assign \new_[51449]_  = \new_[51448]_  & \new_[51441]_ ;
  assign \new_[51453]_  = ~A267 & ~A266;
  assign \new_[51454]_  = ~A233 & \new_[51453]_ ;
  assign \new_[51457]_  = ~A299 & A298;
  assign \new_[51460]_  = A301 & A300;
  assign \new_[51461]_  = \new_[51460]_  & \new_[51457]_ ;
  assign \new_[51462]_  = \new_[51461]_  & \new_[51454]_ ;
  assign \new_[51466]_  = A167 & A169;
  assign \new_[51467]_  = ~A170 & \new_[51466]_ ;
  assign \new_[51470]_  = ~A199 & A166;
  assign \new_[51473]_  = ~A232 & ~A200;
  assign \new_[51474]_  = \new_[51473]_  & \new_[51470]_ ;
  assign \new_[51475]_  = \new_[51474]_  & \new_[51467]_ ;
  assign \new_[51479]_  = ~A267 & ~A266;
  assign \new_[51480]_  = ~A233 & \new_[51479]_ ;
  assign \new_[51483]_  = ~A299 & A298;
  assign \new_[51486]_  = A302 & A300;
  assign \new_[51487]_  = \new_[51486]_  & \new_[51483]_ ;
  assign \new_[51488]_  = \new_[51487]_  & \new_[51480]_ ;
  assign \new_[51492]_  = A167 & A169;
  assign \new_[51493]_  = ~A170 & \new_[51492]_ ;
  assign \new_[51496]_  = ~A199 & A166;
  assign \new_[51499]_  = ~A232 & ~A200;
  assign \new_[51500]_  = \new_[51499]_  & \new_[51496]_ ;
  assign \new_[51501]_  = \new_[51500]_  & \new_[51493]_ ;
  assign \new_[51505]_  = ~A266 & ~A265;
  assign \new_[51506]_  = ~A233 & \new_[51505]_ ;
  assign \new_[51509]_  = ~A299 & A298;
  assign \new_[51512]_  = A301 & A300;
  assign \new_[51513]_  = \new_[51512]_  & \new_[51509]_ ;
  assign \new_[51514]_  = \new_[51513]_  & \new_[51506]_ ;
  assign \new_[51518]_  = A167 & A169;
  assign \new_[51519]_  = ~A170 & \new_[51518]_ ;
  assign \new_[51522]_  = ~A199 & A166;
  assign \new_[51525]_  = ~A232 & ~A200;
  assign \new_[51526]_  = \new_[51525]_  & \new_[51522]_ ;
  assign \new_[51527]_  = \new_[51526]_  & \new_[51519]_ ;
  assign \new_[51531]_  = ~A266 & ~A265;
  assign \new_[51532]_  = ~A233 & \new_[51531]_ ;
  assign \new_[51535]_  = ~A299 & A298;
  assign \new_[51538]_  = A302 & A300;
  assign \new_[51539]_  = \new_[51538]_  & \new_[51535]_ ;
  assign \new_[51540]_  = \new_[51539]_  & \new_[51532]_ ;
  assign \new_[51544]_  = ~A167 & A169;
  assign \new_[51545]_  = ~A170 & \new_[51544]_ ;
  assign \new_[51548]_  = A199 & ~A166;
  assign \new_[51551]_  = A232 & A200;
  assign \new_[51552]_  = \new_[51551]_  & \new_[51548]_ ;
  assign \new_[51553]_  = \new_[51552]_  & \new_[51545]_ ;
  assign \new_[51557]_  = ~A267 & A265;
  assign \new_[51558]_  = A233 & \new_[51557]_ ;
  assign \new_[51561]_  = ~A299 & A298;
  assign \new_[51564]_  = A301 & A300;
  assign \new_[51565]_  = \new_[51564]_  & \new_[51561]_ ;
  assign \new_[51566]_  = \new_[51565]_  & \new_[51558]_ ;
  assign \new_[51570]_  = ~A167 & A169;
  assign \new_[51571]_  = ~A170 & \new_[51570]_ ;
  assign \new_[51574]_  = A199 & ~A166;
  assign \new_[51577]_  = A232 & A200;
  assign \new_[51578]_  = \new_[51577]_  & \new_[51574]_ ;
  assign \new_[51579]_  = \new_[51578]_  & \new_[51571]_ ;
  assign \new_[51583]_  = ~A267 & A265;
  assign \new_[51584]_  = A233 & \new_[51583]_ ;
  assign \new_[51587]_  = ~A299 & A298;
  assign \new_[51590]_  = A302 & A300;
  assign \new_[51591]_  = \new_[51590]_  & \new_[51587]_ ;
  assign \new_[51592]_  = \new_[51591]_  & \new_[51584]_ ;
  assign \new_[51596]_  = ~A167 & A169;
  assign \new_[51597]_  = ~A170 & \new_[51596]_ ;
  assign \new_[51600]_  = A199 & ~A166;
  assign \new_[51603]_  = A232 & A200;
  assign \new_[51604]_  = \new_[51603]_  & \new_[51600]_ ;
  assign \new_[51605]_  = \new_[51604]_  & \new_[51597]_ ;
  assign \new_[51609]_  = A266 & A265;
  assign \new_[51610]_  = A233 & \new_[51609]_ ;
  assign \new_[51613]_  = ~A299 & A298;
  assign \new_[51616]_  = A301 & A300;
  assign \new_[51617]_  = \new_[51616]_  & \new_[51613]_ ;
  assign \new_[51618]_  = \new_[51617]_  & \new_[51610]_ ;
  assign \new_[51622]_  = ~A167 & A169;
  assign \new_[51623]_  = ~A170 & \new_[51622]_ ;
  assign \new_[51626]_  = A199 & ~A166;
  assign \new_[51629]_  = A232 & A200;
  assign \new_[51630]_  = \new_[51629]_  & \new_[51626]_ ;
  assign \new_[51631]_  = \new_[51630]_  & \new_[51623]_ ;
  assign \new_[51635]_  = A266 & A265;
  assign \new_[51636]_  = A233 & \new_[51635]_ ;
  assign \new_[51639]_  = ~A299 & A298;
  assign \new_[51642]_  = A302 & A300;
  assign \new_[51643]_  = \new_[51642]_  & \new_[51639]_ ;
  assign \new_[51644]_  = \new_[51643]_  & \new_[51636]_ ;
  assign \new_[51648]_  = ~A167 & A169;
  assign \new_[51649]_  = ~A170 & \new_[51648]_ ;
  assign \new_[51652]_  = A199 & ~A166;
  assign \new_[51655]_  = A232 & A200;
  assign \new_[51656]_  = \new_[51655]_  & \new_[51652]_ ;
  assign \new_[51657]_  = \new_[51656]_  & \new_[51649]_ ;
  assign \new_[51661]_  = ~A266 & ~A265;
  assign \new_[51662]_  = A233 & \new_[51661]_ ;
  assign \new_[51665]_  = ~A299 & A298;
  assign \new_[51668]_  = A301 & A300;
  assign \new_[51669]_  = \new_[51668]_  & \new_[51665]_ ;
  assign \new_[51670]_  = \new_[51669]_  & \new_[51662]_ ;
  assign \new_[51674]_  = ~A167 & A169;
  assign \new_[51675]_  = ~A170 & \new_[51674]_ ;
  assign \new_[51678]_  = A199 & ~A166;
  assign \new_[51681]_  = A232 & A200;
  assign \new_[51682]_  = \new_[51681]_  & \new_[51678]_ ;
  assign \new_[51683]_  = \new_[51682]_  & \new_[51675]_ ;
  assign \new_[51687]_  = ~A266 & ~A265;
  assign \new_[51688]_  = A233 & \new_[51687]_ ;
  assign \new_[51691]_  = ~A299 & A298;
  assign \new_[51694]_  = A302 & A300;
  assign \new_[51695]_  = \new_[51694]_  & \new_[51691]_ ;
  assign \new_[51696]_  = \new_[51695]_  & \new_[51688]_ ;
  assign \new_[51700]_  = ~A167 & A169;
  assign \new_[51701]_  = ~A170 & \new_[51700]_ ;
  assign \new_[51704]_  = A199 & ~A166;
  assign \new_[51707]_  = ~A233 & A200;
  assign \new_[51708]_  = \new_[51707]_  & \new_[51704]_ ;
  assign \new_[51709]_  = \new_[51708]_  & \new_[51701]_ ;
  assign \new_[51713]_  = ~A266 & ~A236;
  assign \new_[51714]_  = ~A235 & \new_[51713]_ ;
  assign \new_[51717]_  = ~A269 & ~A268;
  assign \new_[51720]_  = A299 & ~A298;
  assign \new_[51721]_  = \new_[51720]_  & \new_[51717]_ ;
  assign \new_[51722]_  = \new_[51721]_  & \new_[51714]_ ;
  assign \new_[51726]_  = ~A167 & A169;
  assign \new_[51727]_  = ~A170 & \new_[51726]_ ;
  assign \new_[51730]_  = A199 & ~A166;
  assign \new_[51733]_  = ~A233 & A200;
  assign \new_[51734]_  = \new_[51733]_  & \new_[51730]_ ;
  assign \new_[51735]_  = \new_[51734]_  & \new_[51727]_ ;
  assign \new_[51739]_  = A266 & A265;
  assign \new_[51740]_  = ~A234 & \new_[51739]_ ;
  assign \new_[51743]_  = ~A299 & A298;
  assign \new_[51746]_  = A301 & A300;
  assign \new_[51747]_  = \new_[51746]_  & \new_[51743]_ ;
  assign \new_[51748]_  = \new_[51747]_  & \new_[51740]_ ;
  assign \new_[51752]_  = ~A167 & A169;
  assign \new_[51753]_  = ~A170 & \new_[51752]_ ;
  assign \new_[51756]_  = A199 & ~A166;
  assign \new_[51759]_  = ~A233 & A200;
  assign \new_[51760]_  = \new_[51759]_  & \new_[51756]_ ;
  assign \new_[51761]_  = \new_[51760]_  & \new_[51753]_ ;
  assign \new_[51765]_  = A266 & A265;
  assign \new_[51766]_  = ~A234 & \new_[51765]_ ;
  assign \new_[51769]_  = ~A299 & A298;
  assign \new_[51772]_  = A302 & A300;
  assign \new_[51773]_  = \new_[51772]_  & \new_[51769]_ ;
  assign \new_[51774]_  = \new_[51773]_  & \new_[51766]_ ;
  assign \new_[51778]_  = ~A167 & A169;
  assign \new_[51779]_  = ~A170 & \new_[51778]_ ;
  assign \new_[51782]_  = A199 & ~A166;
  assign \new_[51785]_  = ~A233 & A200;
  assign \new_[51786]_  = \new_[51785]_  & \new_[51782]_ ;
  assign \new_[51787]_  = \new_[51786]_  & \new_[51779]_ ;
  assign \new_[51791]_  = ~A267 & ~A266;
  assign \new_[51792]_  = ~A234 & \new_[51791]_ ;
  assign \new_[51795]_  = ~A299 & A298;
  assign \new_[51798]_  = A301 & A300;
  assign \new_[51799]_  = \new_[51798]_  & \new_[51795]_ ;
  assign \new_[51800]_  = \new_[51799]_  & \new_[51792]_ ;
  assign \new_[51804]_  = ~A167 & A169;
  assign \new_[51805]_  = ~A170 & \new_[51804]_ ;
  assign \new_[51808]_  = A199 & ~A166;
  assign \new_[51811]_  = ~A233 & A200;
  assign \new_[51812]_  = \new_[51811]_  & \new_[51808]_ ;
  assign \new_[51813]_  = \new_[51812]_  & \new_[51805]_ ;
  assign \new_[51817]_  = ~A267 & ~A266;
  assign \new_[51818]_  = ~A234 & \new_[51817]_ ;
  assign \new_[51821]_  = ~A299 & A298;
  assign \new_[51824]_  = A302 & A300;
  assign \new_[51825]_  = \new_[51824]_  & \new_[51821]_ ;
  assign \new_[51826]_  = \new_[51825]_  & \new_[51818]_ ;
  assign \new_[51830]_  = ~A167 & A169;
  assign \new_[51831]_  = ~A170 & \new_[51830]_ ;
  assign \new_[51834]_  = A199 & ~A166;
  assign \new_[51837]_  = ~A233 & A200;
  assign \new_[51838]_  = \new_[51837]_  & \new_[51834]_ ;
  assign \new_[51839]_  = \new_[51838]_  & \new_[51831]_ ;
  assign \new_[51843]_  = ~A266 & ~A265;
  assign \new_[51844]_  = ~A234 & \new_[51843]_ ;
  assign \new_[51847]_  = ~A299 & A298;
  assign \new_[51850]_  = A301 & A300;
  assign \new_[51851]_  = \new_[51850]_  & \new_[51847]_ ;
  assign \new_[51852]_  = \new_[51851]_  & \new_[51844]_ ;
  assign \new_[51856]_  = ~A167 & A169;
  assign \new_[51857]_  = ~A170 & \new_[51856]_ ;
  assign \new_[51860]_  = A199 & ~A166;
  assign \new_[51863]_  = ~A233 & A200;
  assign \new_[51864]_  = \new_[51863]_  & \new_[51860]_ ;
  assign \new_[51865]_  = \new_[51864]_  & \new_[51857]_ ;
  assign \new_[51869]_  = ~A266 & ~A265;
  assign \new_[51870]_  = ~A234 & \new_[51869]_ ;
  assign \new_[51873]_  = ~A299 & A298;
  assign \new_[51876]_  = A302 & A300;
  assign \new_[51877]_  = \new_[51876]_  & \new_[51873]_ ;
  assign \new_[51878]_  = \new_[51877]_  & \new_[51870]_ ;
  assign \new_[51882]_  = ~A167 & A169;
  assign \new_[51883]_  = ~A170 & \new_[51882]_ ;
  assign \new_[51886]_  = A199 & ~A166;
  assign \new_[51889]_  = A232 & A200;
  assign \new_[51890]_  = \new_[51889]_  & \new_[51886]_ ;
  assign \new_[51891]_  = \new_[51890]_  & \new_[51883]_ ;
  assign \new_[51895]_  = A235 & A234;
  assign \new_[51896]_  = ~A233 & \new_[51895]_ ;
  assign \new_[51899]_  = ~A266 & A265;
  assign \new_[51902]_  = A268 & A267;
  assign \new_[51903]_  = \new_[51902]_  & \new_[51899]_ ;
  assign \new_[51904]_  = \new_[51903]_  & \new_[51896]_ ;
  assign \new_[51908]_  = ~A167 & A169;
  assign \new_[51909]_  = ~A170 & \new_[51908]_ ;
  assign \new_[51912]_  = A199 & ~A166;
  assign \new_[51915]_  = A232 & A200;
  assign \new_[51916]_  = \new_[51915]_  & \new_[51912]_ ;
  assign \new_[51917]_  = \new_[51916]_  & \new_[51909]_ ;
  assign \new_[51921]_  = A235 & A234;
  assign \new_[51922]_  = ~A233 & \new_[51921]_ ;
  assign \new_[51925]_  = ~A266 & A265;
  assign \new_[51928]_  = A269 & A267;
  assign \new_[51929]_  = \new_[51928]_  & \new_[51925]_ ;
  assign \new_[51930]_  = \new_[51929]_  & \new_[51922]_ ;
  assign \new_[51934]_  = ~A167 & A169;
  assign \new_[51935]_  = ~A170 & \new_[51934]_ ;
  assign \new_[51938]_  = A199 & ~A166;
  assign \new_[51941]_  = A232 & A200;
  assign \new_[51942]_  = \new_[51941]_  & \new_[51938]_ ;
  assign \new_[51943]_  = \new_[51942]_  & \new_[51935]_ ;
  assign \new_[51947]_  = A236 & A234;
  assign \new_[51948]_  = ~A233 & \new_[51947]_ ;
  assign \new_[51951]_  = ~A266 & A265;
  assign \new_[51954]_  = A268 & A267;
  assign \new_[51955]_  = \new_[51954]_  & \new_[51951]_ ;
  assign \new_[51956]_  = \new_[51955]_  & \new_[51948]_ ;
  assign \new_[51960]_  = ~A167 & A169;
  assign \new_[51961]_  = ~A170 & \new_[51960]_ ;
  assign \new_[51964]_  = A199 & ~A166;
  assign \new_[51967]_  = A232 & A200;
  assign \new_[51968]_  = \new_[51967]_  & \new_[51964]_ ;
  assign \new_[51969]_  = \new_[51968]_  & \new_[51961]_ ;
  assign \new_[51973]_  = A236 & A234;
  assign \new_[51974]_  = ~A233 & \new_[51973]_ ;
  assign \new_[51977]_  = ~A266 & A265;
  assign \new_[51980]_  = A269 & A267;
  assign \new_[51981]_  = \new_[51980]_  & \new_[51977]_ ;
  assign \new_[51982]_  = \new_[51981]_  & \new_[51974]_ ;
  assign \new_[51986]_  = ~A167 & A169;
  assign \new_[51987]_  = ~A170 & \new_[51986]_ ;
  assign \new_[51990]_  = A199 & ~A166;
  assign \new_[51993]_  = ~A232 & A200;
  assign \new_[51994]_  = \new_[51993]_  & \new_[51990]_ ;
  assign \new_[51995]_  = \new_[51994]_  & \new_[51987]_ ;
  assign \new_[51999]_  = A266 & A265;
  assign \new_[52000]_  = ~A233 & \new_[51999]_ ;
  assign \new_[52003]_  = ~A299 & A298;
  assign \new_[52006]_  = A301 & A300;
  assign \new_[52007]_  = \new_[52006]_  & \new_[52003]_ ;
  assign \new_[52008]_  = \new_[52007]_  & \new_[52000]_ ;
  assign \new_[52012]_  = ~A167 & A169;
  assign \new_[52013]_  = ~A170 & \new_[52012]_ ;
  assign \new_[52016]_  = A199 & ~A166;
  assign \new_[52019]_  = ~A232 & A200;
  assign \new_[52020]_  = \new_[52019]_  & \new_[52016]_ ;
  assign \new_[52021]_  = \new_[52020]_  & \new_[52013]_ ;
  assign \new_[52025]_  = A266 & A265;
  assign \new_[52026]_  = ~A233 & \new_[52025]_ ;
  assign \new_[52029]_  = ~A299 & A298;
  assign \new_[52032]_  = A302 & A300;
  assign \new_[52033]_  = \new_[52032]_  & \new_[52029]_ ;
  assign \new_[52034]_  = \new_[52033]_  & \new_[52026]_ ;
  assign \new_[52038]_  = ~A167 & A169;
  assign \new_[52039]_  = ~A170 & \new_[52038]_ ;
  assign \new_[52042]_  = A199 & ~A166;
  assign \new_[52045]_  = ~A232 & A200;
  assign \new_[52046]_  = \new_[52045]_  & \new_[52042]_ ;
  assign \new_[52047]_  = \new_[52046]_  & \new_[52039]_ ;
  assign \new_[52051]_  = ~A267 & ~A266;
  assign \new_[52052]_  = ~A233 & \new_[52051]_ ;
  assign \new_[52055]_  = ~A299 & A298;
  assign \new_[52058]_  = A301 & A300;
  assign \new_[52059]_  = \new_[52058]_  & \new_[52055]_ ;
  assign \new_[52060]_  = \new_[52059]_  & \new_[52052]_ ;
  assign \new_[52064]_  = ~A167 & A169;
  assign \new_[52065]_  = ~A170 & \new_[52064]_ ;
  assign \new_[52068]_  = A199 & ~A166;
  assign \new_[52071]_  = ~A232 & A200;
  assign \new_[52072]_  = \new_[52071]_  & \new_[52068]_ ;
  assign \new_[52073]_  = \new_[52072]_  & \new_[52065]_ ;
  assign \new_[52077]_  = ~A267 & ~A266;
  assign \new_[52078]_  = ~A233 & \new_[52077]_ ;
  assign \new_[52081]_  = ~A299 & A298;
  assign \new_[52084]_  = A302 & A300;
  assign \new_[52085]_  = \new_[52084]_  & \new_[52081]_ ;
  assign \new_[52086]_  = \new_[52085]_  & \new_[52078]_ ;
  assign \new_[52090]_  = ~A167 & A169;
  assign \new_[52091]_  = ~A170 & \new_[52090]_ ;
  assign \new_[52094]_  = A199 & ~A166;
  assign \new_[52097]_  = ~A232 & A200;
  assign \new_[52098]_  = \new_[52097]_  & \new_[52094]_ ;
  assign \new_[52099]_  = \new_[52098]_  & \new_[52091]_ ;
  assign \new_[52103]_  = ~A266 & ~A265;
  assign \new_[52104]_  = ~A233 & \new_[52103]_ ;
  assign \new_[52107]_  = ~A299 & A298;
  assign \new_[52110]_  = A301 & A300;
  assign \new_[52111]_  = \new_[52110]_  & \new_[52107]_ ;
  assign \new_[52112]_  = \new_[52111]_  & \new_[52104]_ ;
  assign \new_[52116]_  = ~A167 & A169;
  assign \new_[52117]_  = ~A170 & \new_[52116]_ ;
  assign \new_[52120]_  = A199 & ~A166;
  assign \new_[52123]_  = ~A232 & A200;
  assign \new_[52124]_  = \new_[52123]_  & \new_[52120]_ ;
  assign \new_[52125]_  = \new_[52124]_  & \new_[52117]_ ;
  assign \new_[52129]_  = ~A266 & ~A265;
  assign \new_[52130]_  = ~A233 & \new_[52129]_ ;
  assign \new_[52133]_  = ~A299 & A298;
  assign \new_[52136]_  = A302 & A300;
  assign \new_[52137]_  = \new_[52136]_  & \new_[52133]_ ;
  assign \new_[52138]_  = \new_[52137]_  & \new_[52130]_ ;
  assign \new_[52142]_  = ~A167 & A169;
  assign \new_[52143]_  = ~A170 & \new_[52142]_ ;
  assign \new_[52146]_  = ~A200 & ~A166;
  assign \new_[52149]_  = ~A203 & ~A202;
  assign \new_[52150]_  = \new_[52149]_  & \new_[52146]_ ;
  assign \new_[52151]_  = \new_[52150]_  & \new_[52143]_ ;
  assign \new_[52155]_  = A265 & A233;
  assign \new_[52156]_  = A232 & \new_[52155]_ ;
  assign \new_[52159]_  = ~A269 & ~A268;
  assign \new_[52162]_  = A299 & ~A298;
  assign \new_[52163]_  = \new_[52162]_  & \new_[52159]_ ;
  assign \new_[52164]_  = \new_[52163]_  & \new_[52156]_ ;
  assign \new_[52168]_  = ~A167 & A169;
  assign \new_[52169]_  = ~A170 & \new_[52168]_ ;
  assign \new_[52172]_  = ~A200 & ~A166;
  assign \new_[52175]_  = ~A203 & ~A202;
  assign \new_[52176]_  = \new_[52175]_  & \new_[52172]_ ;
  assign \new_[52177]_  = \new_[52176]_  & \new_[52169]_ ;
  assign \new_[52181]_  = ~A236 & ~A235;
  assign \new_[52182]_  = ~A233 & \new_[52181]_ ;
  assign \new_[52185]_  = A266 & A265;
  assign \new_[52188]_  = A299 & ~A298;
  assign \new_[52189]_  = \new_[52188]_  & \new_[52185]_ ;
  assign \new_[52190]_  = \new_[52189]_  & \new_[52182]_ ;
  assign \new_[52194]_  = ~A167 & A169;
  assign \new_[52195]_  = ~A170 & \new_[52194]_ ;
  assign \new_[52198]_  = ~A200 & ~A166;
  assign \new_[52201]_  = ~A203 & ~A202;
  assign \new_[52202]_  = \new_[52201]_  & \new_[52198]_ ;
  assign \new_[52203]_  = \new_[52202]_  & \new_[52195]_ ;
  assign \new_[52207]_  = ~A236 & ~A235;
  assign \new_[52208]_  = ~A233 & \new_[52207]_ ;
  assign \new_[52211]_  = ~A267 & ~A266;
  assign \new_[52214]_  = A299 & ~A298;
  assign \new_[52215]_  = \new_[52214]_  & \new_[52211]_ ;
  assign \new_[52216]_  = \new_[52215]_  & \new_[52208]_ ;
  assign \new_[52220]_  = ~A167 & A169;
  assign \new_[52221]_  = ~A170 & \new_[52220]_ ;
  assign \new_[52224]_  = ~A200 & ~A166;
  assign \new_[52227]_  = ~A203 & ~A202;
  assign \new_[52228]_  = \new_[52227]_  & \new_[52224]_ ;
  assign \new_[52229]_  = \new_[52228]_  & \new_[52221]_ ;
  assign \new_[52233]_  = ~A236 & ~A235;
  assign \new_[52234]_  = ~A233 & \new_[52233]_ ;
  assign \new_[52237]_  = ~A266 & ~A265;
  assign \new_[52240]_  = A299 & ~A298;
  assign \new_[52241]_  = \new_[52240]_  & \new_[52237]_ ;
  assign \new_[52242]_  = \new_[52241]_  & \new_[52234]_ ;
  assign \new_[52246]_  = ~A167 & A169;
  assign \new_[52247]_  = ~A170 & \new_[52246]_ ;
  assign \new_[52250]_  = ~A200 & ~A166;
  assign \new_[52253]_  = ~A203 & ~A202;
  assign \new_[52254]_  = \new_[52253]_  & \new_[52250]_ ;
  assign \new_[52255]_  = \new_[52254]_  & \new_[52247]_ ;
  assign \new_[52259]_  = ~A266 & ~A234;
  assign \new_[52260]_  = ~A233 & \new_[52259]_ ;
  assign \new_[52263]_  = ~A269 & ~A268;
  assign \new_[52266]_  = A299 & ~A298;
  assign \new_[52267]_  = \new_[52266]_  & \new_[52263]_ ;
  assign \new_[52268]_  = \new_[52267]_  & \new_[52260]_ ;
  assign \new_[52272]_  = ~A167 & A169;
  assign \new_[52273]_  = ~A170 & \new_[52272]_ ;
  assign \new_[52276]_  = ~A200 & ~A166;
  assign \new_[52279]_  = ~A203 & ~A202;
  assign \new_[52280]_  = \new_[52279]_  & \new_[52276]_ ;
  assign \new_[52281]_  = \new_[52280]_  & \new_[52273]_ ;
  assign \new_[52285]_  = A234 & ~A233;
  assign \new_[52286]_  = A232 & \new_[52285]_ ;
  assign \new_[52289]_  = A298 & A235;
  assign \new_[52292]_  = ~A302 & ~A301;
  assign \new_[52293]_  = \new_[52292]_  & \new_[52289]_ ;
  assign \new_[52294]_  = \new_[52293]_  & \new_[52286]_ ;
  assign \new_[52298]_  = ~A167 & A169;
  assign \new_[52299]_  = ~A170 & \new_[52298]_ ;
  assign \new_[52302]_  = ~A200 & ~A166;
  assign \new_[52305]_  = ~A203 & ~A202;
  assign \new_[52306]_  = \new_[52305]_  & \new_[52302]_ ;
  assign \new_[52307]_  = \new_[52306]_  & \new_[52299]_ ;
  assign \new_[52311]_  = A234 & ~A233;
  assign \new_[52312]_  = A232 & \new_[52311]_ ;
  assign \new_[52315]_  = A298 & A236;
  assign \new_[52318]_  = ~A302 & ~A301;
  assign \new_[52319]_  = \new_[52318]_  & \new_[52315]_ ;
  assign \new_[52320]_  = \new_[52319]_  & \new_[52312]_ ;
  assign \new_[52324]_  = ~A167 & A169;
  assign \new_[52325]_  = ~A170 & \new_[52324]_ ;
  assign \new_[52328]_  = ~A200 & ~A166;
  assign \new_[52331]_  = ~A203 & ~A202;
  assign \new_[52332]_  = \new_[52331]_  & \new_[52328]_ ;
  assign \new_[52333]_  = \new_[52332]_  & \new_[52325]_ ;
  assign \new_[52337]_  = ~A266 & ~A233;
  assign \new_[52338]_  = ~A232 & \new_[52337]_ ;
  assign \new_[52341]_  = ~A269 & ~A268;
  assign \new_[52344]_  = A299 & ~A298;
  assign \new_[52345]_  = \new_[52344]_  & \new_[52341]_ ;
  assign \new_[52346]_  = \new_[52345]_  & \new_[52338]_ ;
  assign \new_[52350]_  = ~A167 & A169;
  assign \new_[52351]_  = ~A170 & \new_[52350]_ ;
  assign \new_[52354]_  = ~A200 & ~A166;
  assign \new_[52357]_  = A232 & ~A201;
  assign \new_[52358]_  = \new_[52357]_  & \new_[52354]_ ;
  assign \new_[52359]_  = \new_[52358]_  & \new_[52351]_ ;
  assign \new_[52363]_  = ~A267 & A265;
  assign \new_[52364]_  = A233 & \new_[52363]_ ;
  assign \new_[52367]_  = ~A299 & A298;
  assign \new_[52370]_  = A301 & A300;
  assign \new_[52371]_  = \new_[52370]_  & \new_[52367]_ ;
  assign \new_[52372]_  = \new_[52371]_  & \new_[52364]_ ;
  assign \new_[52376]_  = ~A167 & A169;
  assign \new_[52377]_  = ~A170 & \new_[52376]_ ;
  assign \new_[52380]_  = ~A200 & ~A166;
  assign \new_[52383]_  = A232 & ~A201;
  assign \new_[52384]_  = \new_[52383]_  & \new_[52380]_ ;
  assign \new_[52385]_  = \new_[52384]_  & \new_[52377]_ ;
  assign \new_[52389]_  = ~A267 & A265;
  assign \new_[52390]_  = A233 & \new_[52389]_ ;
  assign \new_[52393]_  = ~A299 & A298;
  assign \new_[52396]_  = A302 & A300;
  assign \new_[52397]_  = \new_[52396]_  & \new_[52393]_ ;
  assign \new_[52398]_  = \new_[52397]_  & \new_[52390]_ ;
  assign \new_[52402]_  = ~A167 & A169;
  assign \new_[52403]_  = ~A170 & \new_[52402]_ ;
  assign \new_[52406]_  = ~A200 & ~A166;
  assign \new_[52409]_  = A232 & ~A201;
  assign \new_[52410]_  = \new_[52409]_  & \new_[52406]_ ;
  assign \new_[52411]_  = \new_[52410]_  & \new_[52403]_ ;
  assign \new_[52415]_  = A266 & A265;
  assign \new_[52416]_  = A233 & \new_[52415]_ ;
  assign \new_[52419]_  = ~A299 & A298;
  assign \new_[52422]_  = A301 & A300;
  assign \new_[52423]_  = \new_[52422]_  & \new_[52419]_ ;
  assign \new_[52424]_  = \new_[52423]_  & \new_[52416]_ ;
  assign \new_[52428]_  = ~A167 & A169;
  assign \new_[52429]_  = ~A170 & \new_[52428]_ ;
  assign \new_[52432]_  = ~A200 & ~A166;
  assign \new_[52435]_  = A232 & ~A201;
  assign \new_[52436]_  = \new_[52435]_  & \new_[52432]_ ;
  assign \new_[52437]_  = \new_[52436]_  & \new_[52429]_ ;
  assign \new_[52441]_  = A266 & A265;
  assign \new_[52442]_  = A233 & \new_[52441]_ ;
  assign \new_[52445]_  = ~A299 & A298;
  assign \new_[52448]_  = A302 & A300;
  assign \new_[52449]_  = \new_[52448]_  & \new_[52445]_ ;
  assign \new_[52450]_  = \new_[52449]_  & \new_[52442]_ ;
  assign \new_[52454]_  = ~A167 & A169;
  assign \new_[52455]_  = ~A170 & \new_[52454]_ ;
  assign \new_[52458]_  = ~A200 & ~A166;
  assign \new_[52461]_  = A232 & ~A201;
  assign \new_[52462]_  = \new_[52461]_  & \new_[52458]_ ;
  assign \new_[52463]_  = \new_[52462]_  & \new_[52455]_ ;
  assign \new_[52467]_  = ~A266 & ~A265;
  assign \new_[52468]_  = A233 & \new_[52467]_ ;
  assign \new_[52471]_  = ~A299 & A298;
  assign \new_[52474]_  = A301 & A300;
  assign \new_[52475]_  = \new_[52474]_  & \new_[52471]_ ;
  assign \new_[52476]_  = \new_[52475]_  & \new_[52468]_ ;
  assign \new_[52480]_  = ~A167 & A169;
  assign \new_[52481]_  = ~A170 & \new_[52480]_ ;
  assign \new_[52484]_  = ~A200 & ~A166;
  assign \new_[52487]_  = A232 & ~A201;
  assign \new_[52488]_  = \new_[52487]_  & \new_[52484]_ ;
  assign \new_[52489]_  = \new_[52488]_  & \new_[52481]_ ;
  assign \new_[52493]_  = ~A266 & ~A265;
  assign \new_[52494]_  = A233 & \new_[52493]_ ;
  assign \new_[52497]_  = ~A299 & A298;
  assign \new_[52500]_  = A302 & A300;
  assign \new_[52501]_  = \new_[52500]_  & \new_[52497]_ ;
  assign \new_[52502]_  = \new_[52501]_  & \new_[52494]_ ;
  assign \new_[52506]_  = ~A167 & A169;
  assign \new_[52507]_  = ~A170 & \new_[52506]_ ;
  assign \new_[52510]_  = ~A200 & ~A166;
  assign \new_[52513]_  = ~A233 & ~A201;
  assign \new_[52514]_  = \new_[52513]_  & \new_[52510]_ ;
  assign \new_[52515]_  = \new_[52514]_  & \new_[52507]_ ;
  assign \new_[52519]_  = ~A266 & ~A236;
  assign \new_[52520]_  = ~A235 & \new_[52519]_ ;
  assign \new_[52523]_  = ~A269 & ~A268;
  assign \new_[52526]_  = A299 & ~A298;
  assign \new_[52527]_  = \new_[52526]_  & \new_[52523]_ ;
  assign \new_[52528]_  = \new_[52527]_  & \new_[52520]_ ;
  assign \new_[52532]_  = ~A167 & A169;
  assign \new_[52533]_  = ~A170 & \new_[52532]_ ;
  assign \new_[52536]_  = ~A200 & ~A166;
  assign \new_[52539]_  = ~A233 & ~A201;
  assign \new_[52540]_  = \new_[52539]_  & \new_[52536]_ ;
  assign \new_[52541]_  = \new_[52540]_  & \new_[52533]_ ;
  assign \new_[52545]_  = A266 & A265;
  assign \new_[52546]_  = ~A234 & \new_[52545]_ ;
  assign \new_[52549]_  = ~A299 & A298;
  assign \new_[52552]_  = A301 & A300;
  assign \new_[52553]_  = \new_[52552]_  & \new_[52549]_ ;
  assign \new_[52554]_  = \new_[52553]_  & \new_[52546]_ ;
  assign \new_[52558]_  = ~A167 & A169;
  assign \new_[52559]_  = ~A170 & \new_[52558]_ ;
  assign \new_[52562]_  = ~A200 & ~A166;
  assign \new_[52565]_  = ~A233 & ~A201;
  assign \new_[52566]_  = \new_[52565]_  & \new_[52562]_ ;
  assign \new_[52567]_  = \new_[52566]_  & \new_[52559]_ ;
  assign \new_[52571]_  = A266 & A265;
  assign \new_[52572]_  = ~A234 & \new_[52571]_ ;
  assign \new_[52575]_  = ~A299 & A298;
  assign \new_[52578]_  = A302 & A300;
  assign \new_[52579]_  = \new_[52578]_  & \new_[52575]_ ;
  assign \new_[52580]_  = \new_[52579]_  & \new_[52572]_ ;
  assign \new_[52584]_  = ~A167 & A169;
  assign \new_[52585]_  = ~A170 & \new_[52584]_ ;
  assign \new_[52588]_  = ~A200 & ~A166;
  assign \new_[52591]_  = ~A233 & ~A201;
  assign \new_[52592]_  = \new_[52591]_  & \new_[52588]_ ;
  assign \new_[52593]_  = \new_[52592]_  & \new_[52585]_ ;
  assign \new_[52597]_  = ~A267 & ~A266;
  assign \new_[52598]_  = ~A234 & \new_[52597]_ ;
  assign \new_[52601]_  = ~A299 & A298;
  assign \new_[52604]_  = A301 & A300;
  assign \new_[52605]_  = \new_[52604]_  & \new_[52601]_ ;
  assign \new_[52606]_  = \new_[52605]_  & \new_[52598]_ ;
  assign \new_[52610]_  = ~A167 & A169;
  assign \new_[52611]_  = ~A170 & \new_[52610]_ ;
  assign \new_[52614]_  = ~A200 & ~A166;
  assign \new_[52617]_  = ~A233 & ~A201;
  assign \new_[52618]_  = \new_[52617]_  & \new_[52614]_ ;
  assign \new_[52619]_  = \new_[52618]_  & \new_[52611]_ ;
  assign \new_[52623]_  = ~A267 & ~A266;
  assign \new_[52624]_  = ~A234 & \new_[52623]_ ;
  assign \new_[52627]_  = ~A299 & A298;
  assign \new_[52630]_  = A302 & A300;
  assign \new_[52631]_  = \new_[52630]_  & \new_[52627]_ ;
  assign \new_[52632]_  = \new_[52631]_  & \new_[52624]_ ;
  assign \new_[52636]_  = ~A167 & A169;
  assign \new_[52637]_  = ~A170 & \new_[52636]_ ;
  assign \new_[52640]_  = ~A200 & ~A166;
  assign \new_[52643]_  = ~A233 & ~A201;
  assign \new_[52644]_  = \new_[52643]_  & \new_[52640]_ ;
  assign \new_[52645]_  = \new_[52644]_  & \new_[52637]_ ;
  assign \new_[52649]_  = ~A266 & ~A265;
  assign \new_[52650]_  = ~A234 & \new_[52649]_ ;
  assign \new_[52653]_  = ~A299 & A298;
  assign \new_[52656]_  = A301 & A300;
  assign \new_[52657]_  = \new_[52656]_  & \new_[52653]_ ;
  assign \new_[52658]_  = \new_[52657]_  & \new_[52650]_ ;
  assign \new_[52662]_  = ~A167 & A169;
  assign \new_[52663]_  = ~A170 & \new_[52662]_ ;
  assign \new_[52666]_  = ~A200 & ~A166;
  assign \new_[52669]_  = ~A233 & ~A201;
  assign \new_[52670]_  = \new_[52669]_  & \new_[52666]_ ;
  assign \new_[52671]_  = \new_[52670]_  & \new_[52663]_ ;
  assign \new_[52675]_  = ~A266 & ~A265;
  assign \new_[52676]_  = ~A234 & \new_[52675]_ ;
  assign \new_[52679]_  = ~A299 & A298;
  assign \new_[52682]_  = A302 & A300;
  assign \new_[52683]_  = \new_[52682]_  & \new_[52679]_ ;
  assign \new_[52684]_  = \new_[52683]_  & \new_[52676]_ ;
  assign \new_[52688]_  = ~A167 & A169;
  assign \new_[52689]_  = ~A170 & \new_[52688]_ ;
  assign \new_[52692]_  = ~A200 & ~A166;
  assign \new_[52695]_  = A232 & ~A201;
  assign \new_[52696]_  = \new_[52695]_  & \new_[52692]_ ;
  assign \new_[52697]_  = \new_[52696]_  & \new_[52689]_ ;
  assign \new_[52701]_  = A235 & A234;
  assign \new_[52702]_  = ~A233 & \new_[52701]_ ;
  assign \new_[52705]_  = ~A266 & A265;
  assign \new_[52708]_  = A268 & A267;
  assign \new_[52709]_  = \new_[52708]_  & \new_[52705]_ ;
  assign \new_[52710]_  = \new_[52709]_  & \new_[52702]_ ;
  assign \new_[52714]_  = ~A167 & A169;
  assign \new_[52715]_  = ~A170 & \new_[52714]_ ;
  assign \new_[52718]_  = ~A200 & ~A166;
  assign \new_[52721]_  = A232 & ~A201;
  assign \new_[52722]_  = \new_[52721]_  & \new_[52718]_ ;
  assign \new_[52723]_  = \new_[52722]_  & \new_[52715]_ ;
  assign \new_[52727]_  = A235 & A234;
  assign \new_[52728]_  = ~A233 & \new_[52727]_ ;
  assign \new_[52731]_  = ~A266 & A265;
  assign \new_[52734]_  = A269 & A267;
  assign \new_[52735]_  = \new_[52734]_  & \new_[52731]_ ;
  assign \new_[52736]_  = \new_[52735]_  & \new_[52728]_ ;
  assign \new_[52740]_  = ~A167 & A169;
  assign \new_[52741]_  = ~A170 & \new_[52740]_ ;
  assign \new_[52744]_  = ~A200 & ~A166;
  assign \new_[52747]_  = A232 & ~A201;
  assign \new_[52748]_  = \new_[52747]_  & \new_[52744]_ ;
  assign \new_[52749]_  = \new_[52748]_  & \new_[52741]_ ;
  assign \new_[52753]_  = A236 & A234;
  assign \new_[52754]_  = ~A233 & \new_[52753]_ ;
  assign \new_[52757]_  = ~A266 & A265;
  assign \new_[52760]_  = A268 & A267;
  assign \new_[52761]_  = \new_[52760]_  & \new_[52757]_ ;
  assign \new_[52762]_  = \new_[52761]_  & \new_[52754]_ ;
  assign \new_[52766]_  = ~A167 & A169;
  assign \new_[52767]_  = ~A170 & \new_[52766]_ ;
  assign \new_[52770]_  = ~A200 & ~A166;
  assign \new_[52773]_  = A232 & ~A201;
  assign \new_[52774]_  = \new_[52773]_  & \new_[52770]_ ;
  assign \new_[52775]_  = \new_[52774]_  & \new_[52767]_ ;
  assign \new_[52779]_  = A236 & A234;
  assign \new_[52780]_  = ~A233 & \new_[52779]_ ;
  assign \new_[52783]_  = ~A266 & A265;
  assign \new_[52786]_  = A269 & A267;
  assign \new_[52787]_  = \new_[52786]_  & \new_[52783]_ ;
  assign \new_[52788]_  = \new_[52787]_  & \new_[52780]_ ;
  assign \new_[52792]_  = ~A167 & A169;
  assign \new_[52793]_  = ~A170 & \new_[52792]_ ;
  assign \new_[52796]_  = ~A200 & ~A166;
  assign \new_[52799]_  = ~A232 & ~A201;
  assign \new_[52800]_  = \new_[52799]_  & \new_[52796]_ ;
  assign \new_[52801]_  = \new_[52800]_  & \new_[52793]_ ;
  assign \new_[52805]_  = A266 & A265;
  assign \new_[52806]_  = ~A233 & \new_[52805]_ ;
  assign \new_[52809]_  = ~A299 & A298;
  assign \new_[52812]_  = A301 & A300;
  assign \new_[52813]_  = \new_[52812]_  & \new_[52809]_ ;
  assign \new_[52814]_  = \new_[52813]_  & \new_[52806]_ ;
  assign \new_[52818]_  = ~A167 & A169;
  assign \new_[52819]_  = ~A170 & \new_[52818]_ ;
  assign \new_[52822]_  = ~A200 & ~A166;
  assign \new_[52825]_  = ~A232 & ~A201;
  assign \new_[52826]_  = \new_[52825]_  & \new_[52822]_ ;
  assign \new_[52827]_  = \new_[52826]_  & \new_[52819]_ ;
  assign \new_[52831]_  = A266 & A265;
  assign \new_[52832]_  = ~A233 & \new_[52831]_ ;
  assign \new_[52835]_  = ~A299 & A298;
  assign \new_[52838]_  = A302 & A300;
  assign \new_[52839]_  = \new_[52838]_  & \new_[52835]_ ;
  assign \new_[52840]_  = \new_[52839]_  & \new_[52832]_ ;
  assign \new_[52844]_  = ~A167 & A169;
  assign \new_[52845]_  = ~A170 & \new_[52844]_ ;
  assign \new_[52848]_  = ~A200 & ~A166;
  assign \new_[52851]_  = ~A232 & ~A201;
  assign \new_[52852]_  = \new_[52851]_  & \new_[52848]_ ;
  assign \new_[52853]_  = \new_[52852]_  & \new_[52845]_ ;
  assign \new_[52857]_  = ~A267 & ~A266;
  assign \new_[52858]_  = ~A233 & \new_[52857]_ ;
  assign \new_[52861]_  = ~A299 & A298;
  assign \new_[52864]_  = A301 & A300;
  assign \new_[52865]_  = \new_[52864]_  & \new_[52861]_ ;
  assign \new_[52866]_  = \new_[52865]_  & \new_[52858]_ ;
  assign \new_[52870]_  = ~A167 & A169;
  assign \new_[52871]_  = ~A170 & \new_[52870]_ ;
  assign \new_[52874]_  = ~A200 & ~A166;
  assign \new_[52877]_  = ~A232 & ~A201;
  assign \new_[52878]_  = \new_[52877]_  & \new_[52874]_ ;
  assign \new_[52879]_  = \new_[52878]_  & \new_[52871]_ ;
  assign \new_[52883]_  = ~A267 & ~A266;
  assign \new_[52884]_  = ~A233 & \new_[52883]_ ;
  assign \new_[52887]_  = ~A299 & A298;
  assign \new_[52890]_  = A302 & A300;
  assign \new_[52891]_  = \new_[52890]_  & \new_[52887]_ ;
  assign \new_[52892]_  = \new_[52891]_  & \new_[52884]_ ;
  assign \new_[52896]_  = ~A167 & A169;
  assign \new_[52897]_  = ~A170 & \new_[52896]_ ;
  assign \new_[52900]_  = ~A200 & ~A166;
  assign \new_[52903]_  = ~A232 & ~A201;
  assign \new_[52904]_  = \new_[52903]_  & \new_[52900]_ ;
  assign \new_[52905]_  = \new_[52904]_  & \new_[52897]_ ;
  assign \new_[52909]_  = ~A266 & ~A265;
  assign \new_[52910]_  = ~A233 & \new_[52909]_ ;
  assign \new_[52913]_  = ~A299 & A298;
  assign \new_[52916]_  = A301 & A300;
  assign \new_[52917]_  = \new_[52916]_  & \new_[52913]_ ;
  assign \new_[52918]_  = \new_[52917]_  & \new_[52910]_ ;
  assign \new_[52922]_  = ~A167 & A169;
  assign \new_[52923]_  = ~A170 & \new_[52922]_ ;
  assign \new_[52926]_  = ~A200 & ~A166;
  assign \new_[52929]_  = ~A232 & ~A201;
  assign \new_[52930]_  = \new_[52929]_  & \new_[52926]_ ;
  assign \new_[52931]_  = \new_[52930]_  & \new_[52923]_ ;
  assign \new_[52935]_  = ~A266 & ~A265;
  assign \new_[52936]_  = ~A233 & \new_[52935]_ ;
  assign \new_[52939]_  = ~A299 & A298;
  assign \new_[52942]_  = A302 & A300;
  assign \new_[52943]_  = \new_[52942]_  & \new_[52939]_ ;
  assign \new_[52944]_  = \new_[52943]_  & \new_[52936]_ ;
  assign \new_[52948]_  = ~A167 & A169;
  assign \new_[52949]_  = ~A170 & \new_[52948]_ ;
  assign \new_[52952]_  = ~A199 & ~A166;
  assign \new_[52955]_  = A232 & ~A200;
  assign \new_[52956]_  = \new_[52955]_  & \new_[52952]_ ;
  assign \new_[52957]_  = \new_[52956]_  & \new_[52949]_ ;
  assign \new_[52961]_  = ~A267 & A265;
  assign \new_[52962]_  = A233 & \new_[52961]_ ;
  assign \new_[52965]_  = ~A299 & A298;
  assign \new_[52968]_  = A301 & A300;
  assign \new_[52969]_  = \new_[52968]_  & \new_[52965]_ ;
  assign \new_[52970]_  = \new_[52969]_  & \new_[52962]_ ;
  assign \new_[52974]_  = ~A167 & A169;
  assign \new_[52975]_  = ~A170 & \new_[52974]_ ;
  assign \new_[52978]_  = ~A199 & ~A166;
  assign \new_[52981]_  = A232 & ~A200;
  assign \new_[52982]_  = \new_[52981]_  & \new_[52978]_ ;
  assign \new_[52983]_  = \new_[52982]_  & \new_[52975]_ ;
  assign \new_[52987]_  = ~A267 & A265;
  assign \new_[52988]_  = A233 & \new_[52987]_ ;
  assign \new_[52991]_  = ~A299 & A298;
  assign \new_[52994]_  = A302 & A300;
  assign \new_[52995]_  = \new_[52994]_  & \new_[52991]_ ;
  assign \new_[52996]_  = \new_[52995]_  & \new_[52988]_ ;
  assign \new_[53000]_  = ~A167 & A169;
  assign \new_[53001]_  = ~A170 & \new_[53000]_ ;
  assign \new_[53004]_  = ~A199 & ~A166;
  assign \new_[53007]_  = A232 & ~A200;
  assign \new_[53008]_  = \new_[53007]_  & \new_[53004]_ ;
  assign \new_[53009]_  = \new_[53008]_  & \new_[53001]_ ;
  assign \new_[53013]_  = A266 & A265;
  assign \new_[53014]_  = A233 & \new_[53013]_ ;
  assign \new_[53017]_  = ~A299 & A298;
  assign \new_[53020]_  = A301 & A300;
  assign \new_[53021]_  = \new_[53020]_  & \new_[53017]_ ;
  assign \new_[53022]_  = \new_[53021]_  & \new_[53014]_ ;
  assign \new_[53026]_  = ~A167 & A169;
  assign \new_[53027]_  = ~A170 & \new_[53026]_ ;
  assign \new_[53030]_  = ~A199 & ~A166;
  assign \new_[53033]_  = A232 & ~A200;
  assign \new_[53034]_  = \new_[53033]_  & \new_[53030]_ ;
  assign \new_[53035]_  = \new_[53034]_  & \new_[53027]_ ;
  assign \new_[53039]_  = A266 & A265;
  assign \new_[53040]_  = A233 & \new_[53039]_ ;
  assign \new_[53043]_  = ~A299 & A298;
  assign \new_[53046]_  = A302 & A300;
  assign \new_[53047]_  = \new_[53046]_  & \new_[53043]_ ;
  assign \new_[53048]_  = \new_[53047]_  & \new_[53040]_ ;
  assign \new_[53052]_  = ~A167 & A169;
  assign \new_[53053]_  = ~A170 & \new_[53052]_ ;
  assign \new_[53056]_  = ~A199 & ~A166;
  assign \new_[53059]_  = A232 & ~A200;
  assign \new_[53060]_  = \new_[53059]_  & \new_[53056]_ ;
  assign \new_[53061]_  = \new_[53060]_  & \new_[53053]_ ;
  assign \new_[53065]_  = ~A266 & ~A265;
  assign \new_[53066]_  = A233 & \new_[53065]_ ;
  assign \new_[53069]_  = ~A299 & A298;
  assign \new_[53072]_  = A301 & A300;
  assign \new_[53073]_  = \new_[53072]_  & \new_[53069]_ ;
  assign \new_[53074]_  = \new_[53073]_  & \new_[53066]_ ;
  assign \new_[53078]_  = ~A167 & A169;
  assign \new_[53079]_  = ~A170 & \new_[53078]_ ;
  assign \new_[53082]_  = ~A199 & ~A166;
  assign \new_[53085]_  = A232 & ~A200;
  assign \new_[53086]_  = \new_[53085]_  & \new_[53082]_ ;
  assign \new_[53087]_  = \new_[53086]_  & \new_[53079]_ ;
  assign \new_[53091]_  = ~A266 & ~A265;
  assign \new_[53092]_  = A233 & \new_[53091]_ ;
  assign \new_[53095]_  = ~A299 & A298;
  assign \new_[53098]_  = A302 & A300;
  assign \new_[53099]_  = \new_[53098]_  & \new_[53095]_ ;
  assign \new_[53100]_  = \new_[53099]_  & \new_[53092]_ ;
  assign \new_[53104]_  = ~A167 & A169;
  assign \new_[53105]_  = ~A170 & \new_[53104]_ ;
  assign \new_[53108]_  = ~A199 & ~A166;
  assign \new_[53111]_  = ~A233 & ~A200;
  assign \new_[53112]_  = \new_[53111]_  & \new_[53108]_ ;
  assign \new_[53113]_  = \new_[53112]_  & \new_[53105]_ ;
  assign \new_[53117]_  = ~A266 & ~A236;
  assign \new_[53118]_  = ~A235 & \new_[53117]_ ;
  assign \new_[53121]_  = ~A269 & ~A268;
  assign \new_[53124]_  = A299 & ~A298;
  assign \new_[53125]_  = \new_[53124]_  & \new_[53121]_ ;
  assign \new_[53126]_  = \new_[53125]_  & \new_[53118]_ ;
  assign \new_[53130]_  = ~A167 & A169;
  assign \new_[53131]_  = ~A170 & \new_[53130]_ ;
  assign \new_[53134]_  = ~A199 & ~A166;
  assign \new_[53137]_  = ~A233 & ~A200;
  assign \new_[53138]_  = \new_[53137]_  & \new_[53134]_ ;
  assign \new_[53139]_  = \new_[53138]_  & \new_[53131]_ ;
  assign \new_[53143]_  = A266 & A265;
  assign \new_[53144]_  = ~A234 & \new_[53143]_ ;
  assign \new_[53147]_  = ~A299 & A298;
  assign \new_[53150]_  = A301 & A300;
  assign \new_[53151]_  = \new_[53150]_  & \new_[53147]_ ;
  assign \new_[53152]_  = \new_[53151]_  & \new_[53144]_ ;
  assign \new_[53156]_  = ~A167 & A169;
  assign \new_[53157]_  = ~A170 & \new_[53156]_ ;
  assign \new_[53160]_  = ~A199 & ~A166;
  assign \new_[53163]_  = ~A233 & ~A200;
  assign \new_[53164]_  = \new_[53163]_  & \new_[53160]_ ;
  assign \new_[53165]_  = \new_[53164]_  & \new_[53157]_ ;
  assign \new_[53169]_  = A266 & A265;
  assign \new_[53170]_  = ~A234 & \new_[53169]_ ;
  assign \new_[53173]_  = ~A299 & A298;
  assign \new_[53176]_  = A302 & A300;
  assign \new_[53177]_  = \new_[53176]_  & \new_[53173]_ ;
  assign \new_[53178]_  = \new_[53177]_  & \new_[53170]_ ;
  assign \new_[53182]_  = ~A167 & A169;
  assign \new_[53183]_  = ~A170 & \new_[53182]_ ;
  assign \new_[53186]_  = ~A199 & ~A166;
  assign \new_[53189]_  = ~A233 & ~A200;
  assign \new_[53190]_  = \new_[53189]_  & \new_[53186]_ ;
  assign \new_[53191]_  = \new_[53190]_  & \new_[53183]_ ;
  assign \new_[53195]_  = ~A267 & ~A266;
  assign \new_[53196]_  = ~A234 & \new_[53195]_ ;
  assign \new_[53199]_  = ~A299 & A298;
  assign \new_[53202]_  = A301 & A300;
  assign \new_[53203]_  = \new_[53202]_  & \new_[53199]_ ;
  assign \new_[53204]_  = \new_[53203]_  & \new_[53196]_ ;
  assign \new_[53208]_  = ~A167 & A169;
  assign \new_[53209]_  = ~A170 & \new_[53208]_ ;
  assign \new_[53212]_  = ~A199 & ~A166;
  assign \new_[53215]_  = ~A233 & ~A200;
  assign \new_[53216]_  = \new_[53215]_  & \new_[53212]_ ;
  assign \new_[53217]_  = \new_[53216]_  & \new_[53209]_ ;
  assign \new_[53221]_  = ~A267 & ~A266;
  assign \new_[53222]_  = ~A234 & \new_[53221]_ ;
  assign \new_[53225]_  = ~A299 & A298;
  assign \new_[53228]_  = A302 & A300;
  assign \new_[53229]_  = \new_[53228]_  & \new_[53225]_ ;
  assign \new_[53230]_  = \new_[53229]_  & \new_[53222]_ ;
  assign \new_[53234]_  = ~A167 & A169;
  assign \new_[53235]_  = ~A170 & \new_[53234]_ ;
  assign \new_[53238]_  = ~A199 & ~A166;
  assign \new_[53241]_  = ~A233 & ~A200;
  assign \new_[53242]_  = \new_[53241]_  & \new_[53238]_ ;
  assign \new_[53243]_  = \new_[53242]_  & \new_[53235]_ ;
  assign \new_[53247]_  = ~A266 & ~A265;
  assign \new_[53248]_  = ~A234 & \new_[53247]_ ;
  assign \new_[53251]_  = ~A299 & A298;
  assign \new_[53254]_  = A301 & A300;
  assign \new_[53255]_  = \new_[53254]_  & \new_[53251]_ ;
  assign \new_[53256]_  = \new_[53255]_  & \new_[53248]_ ;
  assign \new_[53260]_  = ~A167 & A169;
  assign \new_[53261]_  = ~A170 & \new_[53260]_ ;
  assign \new_[53264]_  = ~A199 & ~A166;
  assign \new_[53267]_  = ~A233 & ~A200;
  assign \new_[53268]_  = \new_[53267]_  & \new_[53264]_ ;
  assign \new_[53269]_  = \new_[53268]_  & \new_[53261]_ ;
  assign \new_[53273]_  = ~A266 & ~A265;
  assign \new_[53274]_  = ~A234 & \new_[53273]_ ;
  assign \new_[53277]_  = ~A299 & A298;
  assign \new_[53280]_  = A302 & A300;
  assign \new_[53281]_  = \new_[53280]_  & \new_[53277]_ ;
  assign \new_[53282]_  = \new_[53281]_  & \new_[53274]_ ;
  assign \new_[53286]_  = ~A167 & A169;
  assign \new_[53287]_  = ~A170 & \new_[53286]_ ;
  assign \new_[53290]_  = ~A199 & ~A166;
  assign \new_[53293]_  = A232 & ~A200;
  assign \new_[53294]_  = \new_[53293]_  & \new_[53290]_ ;
  assign \new_[53295]_  = \new_[53294]_  & \new_[53287]_ ;
  assign \new_[53299]_  = A235 & A234;
  assign \new_[53300]_  = ~A233 & \new_[53299]_ ;
  assign \new_[53303]_  = ~A266 & A265;
  assign \new_[53306]_  = A268 & A267;
  assign \new_[53307]_  = \new_[53306]_  & \new_[53303]_ ;
  assign \new_[53308]_  = \new_[53307]_  & \new_[53300]_ ;
  assign \new_[53312]_  = ~A167 & A169;
  assign \new_[53313]_  = ~A170 & \new_[53312]_ ;
  assign \new_[53316]_  = ~A199 & ~A166;
  assign \new_[53319]_  = A232 & ~A200;
  assign \new_[53320]_  = \new_[53319]_  & \new_[53316]_ ;
  assign \new_[53321]_  = \new_[53320]_  & \new_[53313]_ ;
  assign \new_[53325]_  = A235 & A234;
  assign \new_[53326]_  = ~A233 & \new_[53325]_ ;
  assign \new_[53329]_  = ~A266 & A265;
  assign \new_[53332]_  = A269 & A267;
  assign \new_[53333]_  = \new_[53332]_  & \new_[53329]_ ;
  assign \new_[53334]_  = \new_[53333]_  & \new_[53326]_ ;
  assign \new_[53338]_  = ~A167 & A169;
  assign \new_[53339]_  = ~A170 & \new_[53338]_ ;
  assign \new_[53342]_  = ~A199 & ~A166;
  assign \new_[53345]_  = A232 & ~A200;
  assign \new_[53346]_  = \new_[53345]_  & \new_[53342]_ ;
  assign \new_[53347]_  = \new_[53346]_  & \new_[53339]_ ;
  assign \new_[53351]_  = A236 & A234;
  assign \new_[53352]_  = ~A233 & \new_[53351]_ ;
  assign \new_[53355]_  = ~A266 & A265;
  assign \new_[53358]_  = A268 & A267;
  assign \new_[53359]_  = \new_[53358]_  & \new_[53355]_ ;
  assign \new_[53360]_  = \new_[53359]_  & \new_[53352]_ ;
  assign \new_[53364]_  = ~A167 & A169;
  assign \new_[53365]_  = ~A170 & \new_[53364]_ ;
  assign \new_[53368]_  = ~A199 & ~A166;
  assign \new_[53371]_  = A232 & ~A200;
  assign \new_[53372]_  = \new_[53371]_  & \new_[53368]_ ;
  assign \new_[53373]_  = \new_[53372]_  & \new_[53365]_ ;
  assign \new_[53377]_  = A236 & A234;
  assign \new_[53378]_  = ~A233 & \new_[53377]_ ;
  assign \new_[53381]_  = ~A266 & A265;
  assign \new_[53384]_  = A269 & A267;
  assign \new_[53385]_  = \new_[53384]_  & \new_[53381]_ ;
  assign \new_[53386]_  = \new_[53385]_  & \new_[53378]_ ;
  assign \new_[53390]_  = ~A167 & A169;
  assign \new_[53391]_  = ~A170 & \new_[53390]_ ;
  assign \new_[53394]_  = ~A199 & ~A166;
  assign \new_[53397]_  = ~A232 & ~A200;
  assign \new_[53398]_  = \new_[53397]_  & \new_[53394]_ ;
  assign \new_[53399]_  = \new_[53398]_  & \new_[53391]_ ;
  assign \new_[53403]_  = A266 & A265;
  assign \new_[53404]_  = ~A233 & \new_[53403]_ ;
  assign \new_[53407]_  = ~A299 & A298;
  assign \new_[53410]_  = A301 & A300;
  assign \new_[53411]_  = \new_[53410]_  & \new_[53407]_ ;
  assign \new_[53412]_  = \new_[53411]_  & \new_[53404]_ ;
  assign \new_[53416]_  = ~A167 & A169;
  assign \new_[53417]_  = ~A170 & \new_[53416]_ ;
  assign \new_[53420]_  = ~A199 & ~A166;
  assign \new_[53423]_  = ~A232 & ~A200;
  assign \new_[53424]_  = \new_[53423]_  & \new_[53420]_ ;
  assign \new_[53425]_  = \new_[53424]_  & \new_[53417]_ ;
  assign \new_[53429]_  = A266 & A265;
  assign \new_[53430]_  = ~A233 & \new_[53429]_ ;
  assign \new_[53433]_  = ~A299 & A298;
  assign \new_[53436]_  = A302 & A300;
  assign \new_[53437]_  = \new_[53436]_  & \new_[53433]_ ;
  assign \new_[53438]_  = \new_[53437]_  & \new_[53430]_ ;
  assign \new_[53442]_  = ~A167 & A169;
  assign \new_[53443]_  = ~A170 & \new_[53442]_ ;
  assign \new_[53446]_  = ~A199 & ~A166;
  assign \new_[53449]_  = ~A232 & ~A200;
  assign \new_[53450]_  = \new_[53449]_  & \new_[53446]_ ;
  assign \new_[53451]_  = \new_[53450]_  & \new_[53443]_ ;
  assign \new_[53455]_  = ~A267 & ~A266;
  assign \new_[53456]_  = ~A233 & \new_[53455]_ ;
  assign \new_[53459]_  = ~A299 & A298;
  assign \new_[53462]_  = A301 & A300;
  assign \new_[53463]_  = \new_[53462]_  & \new_[53459]_ ;
  assign \new_[53464]_  = \new_[53463]_  & \new_[53456]_ ;
  assign \new_[53468]_  = ~A167 & A169;
  assign \new_[53469]_  = ~A170 & \new_[53468]_ ;
  assign \new_[53472]_  = ~A199 & ~A166;
  assign \new_[53475]_  = ~A232 & ~A200;
  assign \new_[53476]_  = \new_[53475]_  & \new_[53472]_ ;
  assign \new_[53477]_  = \new_[53476]_  & \new_[53469]_ ;
  assign \new_[53481]_  = ~A267 & ~A266;
  assign \new_[53482]_  = ~A233 & \new_[53481]_ ;
  assign \new_[53485]_  = ~A299 & A298;
  assign \new_[53488]_  = A302 & A300;
  assign \new_[53489]_  = \new_[53488]_  & \new_[53485]_ ;
  assign \new_[53490]_  = \new_[53489]_  & \new_[53482]_ ;
  assign \new_[53494]_  = ~A167 & A169;
  assign \new_[53495]_  = ~A170 & \new_[53494]_ ;
  assign \new_[53498]_  = ~A199 & ~A166;
  assign \new_[53501]_  = ~A232 & ~A200;
  assign \new_[53502]_  = \new_[53501]_  & \new_[53498]_ ;
  assign \new_[53503]_  = \new_[53502]_  & \new_[53495]_ ;
  assign \new_[53507]_  = ~A266 & ~A265;
  assign \new_[53508]_  = ~A233 & \new_[53507]_ ;
  assign \new_[53511]_  = ~A299 & A298;
  assign \new_[53514]_  = A301 & A300;
  assign \new_[53515]_  = \new_[53514]_  & \new_[53511]_ ;
  assign \new_[53516]_  = \new_[53515]_  & \new_[53508]_ ;
  assign \new_[53520]_  = ~A167 & A169;
  assign \new_[53521]_  = ~A170 & \new_[53520]_ ;
  assign \new_[53524]_  = ~A199 & ~A166;
  assign \new_[53527]_  = ~A232 & ~A200;
  assign \new_[53528]_  = \new_[53527]_  & \new_[53524]_ ;
  assign \new_[53529]_  = \new_[53528]_  & \new_[53521]_ ;
  assign \new_[53533]_  = ~A266 & ~A265;
  assign \new_[53534]_  = ~A233 & \new_[53533]_ ;
  assign \new_[53537]_  = ~A299 & A298;
  assign \new_[53540]_  = A302 & A300;
  assign \new_[53541]_  = \new_[53540]_  & \new_[53537]_ ;
  assign \new_[53542]_  = \new_[53541]_  & \new_[53534]_ ;
  assign \new_[53546]_  = ~A166 & ~A167;
  assign \new_[53547]_  = ~A169 & \new_[53546]_ ;
  assign \new_[53550]_  = A200 & ~A199;
  assign \new_[53553]_  = A233 & A232;
  assign \new_[53554]_  = \new_[53553]_  & \new_[53550]_ ;
  assign \new_[53555]_  = \new_[53554]_  & \new_[53547]_ ;
  assign \new_[53559]_  = ~A269 & ~A268;
  assign \new_[53560]_  = A265 & \new_[53559]_ ;
  assign \new_[53563]_  = ~A299 & A298;
  assign \new_[53566]_  = A301 & A300;
  assign \new_[53567]_  = \new_[53566]_  & \new_[53563]_ ;
  assign \new_[53568]_  = \new_[53567]_  & \new_[53560]_ ;
  assign \new_[53572]_  = ~A166 & ~A167;
  assign \new_[53573]_  = ~A169 & \new_[53572]_ ;
  assign \new_[53576]_  = A200 & ~A199;
  assign \new_[53579]_  = A233 & A232;
  assign \new_[53580]_  = \new_[53579]_  & \new_[53576]_ ;
  assign \new_[53581]_  = \new_[53580]_  & \new_[53573]_ ;
  assign \new_[53585]_  = ~A269 & ~A268;
  assign \new_[53586]_  = A265 & \new_[53585]_ ;
  assign \new_[53589]_  = ~A299 & A298;
  assign \new_[53592]_  = A302 & A300;
  assign \new_[53593]_  = \new_[53592]_  & \new_[53589]_ ;
  assign \new_[53594]_  = \new_[53593]_  & \new_[53586]_ ;
  assign \new_[53598]_  = ~A166 & ~A167;
  assign \new_[53599]_  = ~A169 & \new_[53598]_ ;
  assign \new_[53602]_  = A200 & ~A199;
  assign \new_[53605]_  = ~A235 & ~A233;
  assign \new_[53606]_  = \new_[53605]_  & \new_[53602]_ ;
  assign \new_[53607]_  = \new_[53606]_  & \new_[53599]_ ;
  assign \new_[53611]_  = A266 & A265;
  assign \new_[53612]_  = ~A236 & \new_[53611]_ ;
  assign \new_[53615]_  = ~A299 & A298;
  assign \new_[53618]_  = A301 & A300;
  assign \new_[53619]_  = \new_[53618]_  & \new_[53615]_ ;
  assign \new_[53620]_  = \new_[53619]_  & \new_[53612]_ ;
  assign \new_[53624]_  = ~A166 & ~A167;
  assign \new_[53625]_  = ~A169 & \new_[53624]_ ;
  assign \new_[53628]_  = A200 & ~A199;
  assign \new_[53631]_  = ~A235 & ~A233;
  assign \new_[53632]_  = \new_[53631]_  & \new_[53628]_ ;
  assign \new_[53633]_  = \new_[53632]_  & \new_[53625]_ ;
  assign \new_[53637]_  = A266 & A265;
  assign \new_[53638]_  = ~A236 & \new_[53637]_ ;
  assign \new_[53641]_  = ~A299 & A298;
  assign \new_[53644]_  = A302 & A300;
  assign \new_[53645]_  = \new_[53644]_  & \new_[53641]_ ;
  assign \new_[53646]_  = \new_[53645]_  & \new_[53638]_ ;
  assign \new_[53650]_  = ~A166 & ~A167;
  assign \new_[53651]_  = ~A169 & \new_[53650]_ ;
  assign \new_[53654]_  = A200 & ~A199;
  assign \new_[53657]_  = ~A235 & ~A233;
  assign \new_[53658]_  = \new_[53657]_  & \new_[53654]_ ;
  assign \new_[53659]_  = \new_[53658]_  & \new_[53651]_ ;
  assign \new_[53663]_  = ~A267 & ~A266;
  assign \new_[53664]_  = ~A236 & \new_[53663]_ ;
  assign \new_[53667]_  = ~A299 & A298;
  assign \new_[53670]_  = A301 & A300;
  assign \new_[53671]_  = \new_[53670]_  & \new_[53667]_ ;
  assign \new_[53672]_  = \new_[53671]_  & \new_[53664]_ ;
  assign \new_[53676]_  = ~A166 & ~A167;
  assign \new_[53677]_  = ~A169 & \new_[53676]_ ;
  assign \new_[53680]_  = A200 & ~A199;
  assign \new_[53683]_  = ~A235 & ~A233;
  assign \new_[53684]_  = \new_[53683]_  & \new_[53680]_ ;
  assign \new_[53685]_  = \new_[53684]_  & \new_[53677]_ ;
  assign \new_[53689]_  = ~A267 & ~A266;
  assign \new_[53690]_  = ~A236 & \new_[53689]_ ;
  assign \new_[53693]_  = ~A299 & A298;
  assign \new_[53696]_  = A302 & A300;
  assign \new_[53697]_  = \new_[53696]_  & \new_[53693]_ ;
  assign \new_[53698]_  = \new_[53697]_  & \new_[53690]_ ;
  assign \new_[53702]_  = ~A166 & ~A167;
  assign \new_[53703]_  = ~A169 & \new_[53702]_ ;
  assign \new_[53706]_  = A200 & ~A199;
  assign \new_[53709]_  = ~A235 & ~A233;
  assign \new_[53710]_  = \new_[53709]_  & \new_[53706]_ ;
  assign \new_[53711]_  = \new_[53710]_  & \new_[53703]_ ;
  assign \new_[53715]_  = ~A266 & ~A265;
  assign \new_[53716]_  = ~A236 & \new_[53715]_ ;
  assign \new_[53719]_  = ~A299 & A298;
  assign \new_[53722]_  = A301 & A300;
  assign \new_[53723]_  = \new_[53722]_  & \new_[53719]_ ;
  assign \new_[53724]_  = \new_[53723]_  & \new_[53716]_ ;
  assign \new_[53728]_  = ~A166 & ~A167;
  assign \new_[53729]_  = ~A169 & \new_[53728]_ ;
  assign \new_[53732]_  = A200 & ~A199;
  assign \new_[53735]_  = ~A235 & ~A233;
  assign \new_[53736]_  = \new_[53735]_  & \new_[53732]_ ;
  assign \new_[53737]_  = \new_[53736]_  & \new_[53729]_ ;
  assign \new_[53741]_  = ~A266 & ~A265;
  assign \new_[53742]_  = ~A236 & \new_[53741]_ ;
  assign \new_[53745]_  = ~A299 & A298;
  assign \new_[53748]_  = A302 & A300;
  assign \new_[53749]_  = \new_[53748]_  & \new_[53745]_ ;
  assign \new_[53750]_  = \new_[53749]_  & \new_[53742]_ ;
  assign \new_[53754]_  = ~A166 & ~A167;
  assign \new_[53755]_  = ~A169 & \new_[53754]_ ;
  assign \new_[53758]_  = A200 & ~A199;
  assign \new_[53761]_  = ~A234 & ~A233;
  assign \new_[53762]_  = \new_[53761]_  & \new_[53758]_ ;
  assign \new_[53763]_  = \new_[53762]_  & \new_[53755]_ ;
  assign \new_[53767]_  = ~A269 & ~A268;
  assign \new_[53768]_  = ~A266 & \new_[53767]_ ;
  assign \new_[53771]_  = ~A299 & A298;
  assign \new_[53774]_  = A301 & A300;
  assign \new_[53775]_  = \new_[53774]_  & \new_[53771]_ ;
  assign \new_[53776]_  = \new_[53775]_  & \new_[53768]_ ;
  assign \new_[53780]_  = ~A166 & ~A167;
  assign \new_[53781]_  = ~A169 & \new_[53780]_ ;
  assign \new_[53784]_  = A200 & ~A199;
  assign \new_[53787]_  = ~A234 & ~A233;
  assign \new_[53788]_  = \new_[53787]_  & \new_[53784]_ ;
  assign \new_[53789]_  = \new_[53788]_  & \new_[53781]_ ;
  assign \new_[53793]_  = ~A269 & ~A268;
  assign \new_[53794]_  = ~A266 & \new_[53793]_ ;
  assign \new_[53797]_  = ~A299 & A298;
  assign \new_[53800]_  = A302 & A300;
  assign \new_[53801]_  = \new_[53800]_  & \new_[53797]_ ;
  assign \new_[53802]_  = \new_[53801]_  & \new_[53794]_ ;
  assign \new_[53806]_  = ~A166 & ~A167;
  assign \new_[53807]_  = ~A169 & \new_[53806]_ ;
  assign \new_[53810]_  = A200 & ~A199;
  assign \new_[53813]_  = ~A233 & ~A232;
  assign \new_[53814]_  = \new_[53813]_  & \new_[53810]_ ;
  assign \new_[53815]_  = \new_[53814]_  & \new_[53807]_ ;
  assign \new_[53819]_  = ~A269 & ~A268;
  assign \new_[53820]_  = ~A266 & \new_[53819]_ ;
  assign \new_[53823]_  = ~A299 & A298;
  assign \new_[53826]_  = A301 & A300;
  assign \new_[53827]_  = \new_[53826]_  & \new_[53823]_ ;
  assign \new_[53828]_  = \new_[53827]_  & \new_[53820]_ ;
  assign \new_[53832]_  = ~A166 & ~A167;
  assign \new_[53833]_  = ~A169 & \new_[53832]_ ;
  assign \new_[53836]_  = A200 & ~A199;
  assign \new_[53839]_  = ~A233 & ~A232;
  assign \new_[53840]_  = \new_[53839]_  & \new_[53836]_ ;
  assign \new_[53841]_  = \new_[53840]_  & \new_[53833]_ ;
  assign \new_[53845]_  = ~A269 & ~A268;
  assign \new_[53846]_  = ~A266 & \new_[53845]_ ;
  assign \new_[53849]_  = ~A299 & A298;
  assign \new_[53852]_  = A302 & A300;
  assign \new_[53853]_  = \new_[53852]_  & \new_[53849]_ ;
  assign \new_[53854]_  = \new_[53853]_  & \new_[53846]_ ;
  assign \new_[53858]_  = ~A166 & ~A167;
  assign \new_[53859]_  = ~A169 & \new_[53858]_ ;
  assign \new_[53862]_  = ~A200 & A199;
  assign \new_[53865]_  = A202 & A201;
  assign \new_[53866]_  = \new_[53865]_  & \new_[53862]_ ;
  assign \new_[53867]_  = \new_[53866]_  & \new_[53859]_ ;
  assign \new_[53871]_  = A265 & A233;
  assign \new_[53872]_  = A232 & \new_[53871]_ ;
  assign \new_[53875]_  = ~A269 & ~A268;
  assign \new_[53878]_  = A299 & ~A298;
  assign \new_[53879]_  = \new_[53878]_  & \new_[53875]_ ;
  assign \new_[53880]_  = \new_[53879]_  & \new_[53872]_ ;
  assign \new_[53884]_  = ~A166 & ~A167;
  assign \new_[53885]_  = ~A169 & \new_[53884]_ ;
  assign \new_[53888]_  = ~A200 & A199;
  assign \new_[53891]_  = A202 & A201;
  assign \new_[53892]_  = \new_[53891]_  & \new_[53888]_ ;
  assign \new_[53893]_  = \new_[53892]_  & \new_[53885]_ ;
  assign \new_[53897]_  = ~A236 & ~A235;
  assign \new_[53898]_  = ~A233 & \new_[53897]_ ;
  assign \new_[53901]_  = A266 & A265;
  assign \new_[53904]_  = A299 & ~A298;
  assign \new_[53905]_  = \new_[53904]_  & \new_[53901]_ ;
  assign \new_[53906]_  = \new_[53905]_  & \new_[53898]_ ;
  assign \new_[53910]_  = ~A166 & ~A167;
  assign \new_[53911]_  = ~A169 & \new_[53910]_ ;
  assign \new_[53914]_  = ~A200 & A199;
  assign \new_[53917]_  = A202 & A201;
  assign \new_[53918]_  = \new_[53917]_  & \new_[53914]_ ;
  assign \new_[53919]_  = \new_[53918]_  & \new_[53911]_ ;
  assign \new_[53923]_  = ~A236 & ~A235;
  assign \new_[53924]_  = ~A233 & \new_[53923]_ ;
  assign \new_[53927]_  = ~A267 & ~A266;
  assign \new_[53930]_  = A299 & ~A298;
  assign \new_[53931]_  = \new_[53930]_  & \new_[53927]_ ;
  assign \new_[53932]_  = \new_[53931]_  & \new_[53924]_ ;
  assign \new_[53936]_  = ~A166 & ~A167;
  assign \new_[53937]_  = ~A169 & \new_[53936]_ ;
  assign \new_[53940]_  = ~A200 & A199;
  assign \new_[53943]_  = A202 & A201;
  assign \new_[53944]_  = \new_[53943]_  & \new_[53940]_ ;
  assign \new_[53945]_  = \new_[53944]_  & \new_[53937]_ ;
  assign \new_[53949]_  = ~A236 & ~A235;
  assign \new_[53950]_  = ~A233 & \new_[53949]_ ;
  assign \new_[53953]_  = ~A266 & ~A265;
  assign \new_[53956]_  = A299 & ~A298;
  assign \new_[53957]_  = \new_[53956]_  & \new_[53953]_ ;
  assign \new_[53958]_  = \new_[53957]_  & \new_[53950]_ ;
  assign \new_[53962]_  = ~A166 & ~A167;
  assign \new_[53963]_  = ~A169 & \new_[53962]_ ;
  assign \new_[53966]_  = ~A200 & A199;
  assign \new_[53969]_  = A202 & A201;
  assign \new_[53970]_  = \new_[53969]_  & \new_[53966]_ ;
  assign \new_[53971]_  = \new_[53970]_  & \new_[53963]_ ;
  assign \new_[53975]_  = ~A266 & ~A234;
  assign \new_[53976]_  = ~A233 & \new_[53975]_ ;
  assign \new_[53979]_  = ~A269 & ~A268;
  assign \new_[53982]_  = A299 & ~A298;
  assign \new_[53983]_  = \new_[53982]_  & \new_[53979]_ ;
  assign \new_[53984]_  = \new_[53983]_  & \new_[53976]_ ;
  assign \new_[53988]_  = ~A166 & ~A167;
  assign \new_[53989]_  = ~A169 & \new_[53988]_ ;
  assign \new_[53992]_  = ~A200 & A199;
  assign \new_[53995]_  = A202 & A201;
  assign \new_[53996]_  = \new_[53995]_  & \new_[53992]_ ;
  assign \new_[53997]_  = \new_[53996]_  & \new_[53989]_ ;
  assign \new_[54001]_  = A234 & ~A233;
  assign \new_[54002]_  = A232 & \new_[54001]_ ;
  assign \new_[54005]_  = A298 & A235;
  assign \new_[54008]_  = ~A302 & ~A301;
  assign \new_[54009]_  = \new_[54008]_  & \new_[54005]_ ;
  assign \new_[54010]_  = \new_[54009]_  & \new_[54002]_ ;
  assign \new_[54014]_  = ~A166 & ~A167;
  assign \new_[54015]_  = ~A169 & \new_[54014]_ ;
  assign \new_[54018]_  = ~A200 & A199;
  assign \new_[54021]_  = A202 & A201;
  assign \new_[54022]_  = \new_[54021]_  & \new_[54018]_ ;
  assign \new_[54023]_  = \new_[54022]_  & \new_[54015]_ ;
  assign \new_[54027]_  = A234 & ~A233;
  assign \new_[54028]_  = A232 & \new_[54027]_ ;
  assign \new_[54031]_  = A298 & A236;
  assign \new_[54034]_  = ~A302 & ~A301;
  assign \new_[54035]_  = \new_[54034]_  & \new_[54031]_ ;
  assign \new_[54036]_  = \new_[54035]_  & \new_[54028]_ ;
  assign \new_[54040]_  = ~A166 & ~A167;
  assign \new_[54041]_  = ~A169 & \new_[54040]_ ;
  assign \new_[54044]_  = ~A200 & A199;
  assign \new_[54047]_  = A202 & A201;
  assign \new_[54048]_  = \new_[54047]_  & \new_[54044]_ ;
  assign \new_[54049]_  = \new_[54048]_  & \new_[54041]_ ;
  assign \new_[54053]_  = ~A266 & ~A233;
  assign \new_[54054]_  = ~A232 & \new_[54053]_ ;
  assign \new_[54057]_  = ~A269 & ~A268;
  assign \new_[54060]_  = A299 & ~A298;
  assign \new_[54061]_  = \new_[54060]_  & \new_[54057]_ ;
  assign \new_[54062]_  = \new_[54061]_  & \new_[54054]_ ;
  assign \new_[54066]_  = ~A166 & ~A167;
  assign \new_[54067]_  = ~A169 & \new_[54066]_ ;
  assign \new_[54070]_  = ~A200 & A199;
  assign \new_[54073]_  = A203 & A201;
  assign \new_[54074]_  = \new_[54073]_  & \new_[54070]_ ;
  assign \new_[54075]_  = \new_[54074]_  & \new_[54067]_ ;
  assign \new_[54079]_  = A265 & A233;
  assign \new_[54080]_  = A232 & \new_[54079]_ ;
  assign \new_[54083]_  = ~A269 & ~A268;
  assign \new_[54086]_  = A299 & ~A298;
  assign \new_[54087]_  = \new_[54086]_  & \new_[54083]_ ;
  assign \new_[54088]_  = \new_[54087]_  & \new_[54080]_ ;
  assign \new_[54092]_  = ~A166 & ~A167;
  assign \new_[54093]_  = ~A169 & \new_[54092]_ ;
  assign \new_[54096]_  = ~A200 & A199;
  assign \new_[54099]_  = A203 & A201;
  assign \new_[54100]_  = \new_[54099]_  & \new_[54096]_ ;
  assign \new_[54101]_  = \new_[54100]_  & \new_[54093]_ ;
  assign \new_[54105]_  = ~A236 & ~A235;
  assign \new_[54106]_  = ~A233 & \new_[54105]_ ;
  assign \new_[54109]_  = A266 & A265;
  assign \new_[54112]_  = A299 & ~A298;
  assign \new_[54113]_  = \new_[54112]_  & \new_[54109]_ ;
  assign \new_[54114]_  = \new_[54113]_  & \new_[54106]_ ;
  assign \new_[54118]_  = ~A166 & ~A167;
  assign \new_[54119]_  = ~A169 & \new_[54118]_ ;
  assign \new_[54122]_  = ~A200 & A199;
  assign \new_[54125]_  = A203 & A201;
  assign \new_[54126]_  = \new_[54125]_  & \new_[54122]_ ;
  assign \new_[54127]_  = \new_[54126]_  & \new_[54119]_ ;
  assign \new_[54131]_  = ~A236 & ~A235;
  assign \new_[54132]_  = ~A233 & \new_[54131]_ ;
  assign \new_[54135]_  = ~A267 & ~A266;
  assign \new_[54138]_  = A299 & ~A298;
  assign \new_[54139]_  = \new_[54138]_  & \new_[54135]_ ;
  assign \new_[54140]_  = \new_[54139]_  & \new_[54132]_ ;
  assign \new_[54144]_  = ~A166 & ~A167;
  assign \new_[54145]_  = ~A169 & \new_[54144]_ ;
  assign \new_[54148]_  = ~A200 & A199;
  assign \new_[54151]_  = A203 & A201;
  assign \new_[54152]_  = \new_[54151]_  & \new_[54148]_ ;
  assign \new_[54153]_  = \new_[54152]_  & \new_[54145]_ ;
  assign \new_[54157]_  = ~A236 & ~A235;
  assign \new_[54158]_  = ~A233 & \new_[54157]_ ;
  assign \new_[54161]_  = ~A266 & ~A265;
  assign \new_[54164]_  = A299 & ~A298;
  assign \new_[54165]_  = \new_[54164]_  & \new_[54161]_ ;
  assign \new_[54166]_  = \new_[54165]_  & \new_[54158]_ ;
  assign \new_[54170]_  = ~A166 & ~A167;
  assign \new_[54171]_  = ~A169 & \new_[54170]_ ;
  assign \new_[54174]_  = ~A200 & A199;
  assign \new_[54177]_  = A203 & A201;
  assign \new_[54178]_  = \new_[54177]_  & \new_[54174]_ ;
  assign \new_[54179]_  = \new_[54178]_  & \new_[54171]_ ;
  assign \new_[54183]_  = ~A266 & ~A234;
  assign \new_[54184]_  = ~A233 & \new_[54183]_ ;
  assign \new_[54187]_  = ~A269 & ~A268;
  assign \new_[54190]_  = A299 & ~A298;
  assign \new_[54191]_  = \new_[54190]_  & \new_[54187]_ ;
  assign \new_[54192]_  = \new_[54191]_  & \new_[54184]_ ;
  assign \new_[54196]_  = ~A166 & ~A167;
  assign \new_[54197]_  = ~A169 & \new_[54196]_ ;
  assign \new_[54200]_  = ~A200 & A199;
  assign \new_[54203]_  = A203 & A201;
  assign \new_[54204]_  = \new_[54203]_  & \new_[54200]_ ;
  assign \new_[54205]_  = \new_[54204]_  & \new_[54197]_ ;
  assign \new_[54209]_  = A234 & ~A233;
  assign \new_[54210]_  = A232 & \new_[54209]_ ;
  assign \new_[54213]_  = A298 & A235;
  assign \new_[54216]_  = ~A302 & ~A301;
  assign \new_[54217]_  = \new_[54216]_  & \new_[54213]_ ;
  assign \new_[54218]_  = \new_[54217]_  & \new_[54210]_ ;
  assign \new_[54222]_  = ~A166 & ~A167;
  assign \new_[54223]_  = ~A169 & \new_[54222]_ ;
  assign \new_[54226]_  = ~A200 & A199;
  assign \new_[54229]_  = A203 & A201;
  assign \new_[54230]_  = \new_[54229]_  & \new_[54226]_ ;
  assign \new_[54231]_  = \new_[54230]_  & \new_[54223]_ ;
  assign \new_[54235]_  = A234 & ~A233;
  assign \new_[54236]_  = A232 & \new_[54235]_ ;
  assign \new_[54239]_  = A298 & A236;
  assign \new_[54242]_  = ~A302 & ~A301;
  assign \new_[54243]_  = \new_[54242]_  & \new_[54239]_ ;
  assign \new_[54244]_  = \new_[54243]_  & \new_[54236]_ ;
  assign \new_[54248]_  = ~A166 & ~A167;
  assign \new_[54249]_  = ~A169 & \new_[54248]_ ;
  assign \new_[54252]_  = ~A200 & A199;
  assign \new_[54255]_  = A203 & A201;
  assign \new_[54256]_  = \new_[54255]_  & \new_[54252]_ ;
  assign \new_[54257]_  = \new_[54256]_  & \new_[54249]_ ;
  assign \new_[54261]_  = ~A266 & ~A233;
  assign \new_[54262]_  = ~A232 & \new_[54261]_ ;
  assign \new_[54265]_  = ~A269 & ~A268;
  assign \new_[54268]_  = A299 & ~A298;
  assign \new_[54269]_  = \new_[54268]_  & \new_[54265]_ ;
  assign \new_[54270]_  = \new_[54269]_  & \new_[54262]_ ;
  assign \new_[54274]_  = A167 & ~A168;
  assign \new_[54275]_  = ~A169 & \new_[54274]_ ;
  assign \new_[54278]_  = ~A199 & A166;
  assign \new_[54281]_  = A232 & A200;
  assign \new_[54282]_  = \new_[54281]_  & \new_[54278]_ ;
  assign \new_[54283]_  = \new_[54282]_  & \new_[54275]_ ;
  assign \new_[54287]_  = ~A267 & A265;
  assign \new_[54288]_  = A233 & \new_[54287]_ ;
  assign \new_[54291]_  = ~A299 & A298;
  assign \new_[54294]_  = A301 & A300;
  assign \new_[54295]_  = \new_[54294]_  & \new_[54291]_ ;
  assign \new_[54296]_  = \new_[54295]_  & \new_[54288]_ ;
  assign \new_[54300]_  = A167 & ~A168;
  assign \new_[54301]_  = ~A169 & \new_[54300]_ ;
  assign \new_[54304]_  = ~A199 & A166;
  assign \new_[54307]_  = A232 & A200;
  assign \new_[54308]_  = \new_[54307]_  & \new_[54304]_ ;
  assign \new_[54309]_  = \new_[54308]_  & \new_[54301]_ ;
  assign \new_[54313]_  = ~A267 & A265;
  assign \new_[54314]_  = A233 & \new_[54313]_ ;
  assign \new_[54317]_  = ~A299 & A298;
  assign \new_[54320]_  = A302 & A300;
  assign \new_[54321]_  = \new_[54320]_  & \new_[54317]_ ;
  assign \new_[54322]_  = \new_[54321]_  & \new_[54314]_ ;
  assign \new_[54326]_  = A167 & ~A168;
  assign \new_[54327]_  = ~A169 & \new_[54326]_ ;
  assign \new_[54330]_  = ~A199 & A166;
  assign \new_[54333]_  = A232 & A200;
  assign \new_[54334]_  = \new_[54333]_  & \new_[54330]_ ;
  assign \new_[54335]_  = \new_[54334]_  & \new_[54327]_ ;
  assign \new_[54339]_  = A266 & A265;
  assign \new_[54340]_  = A233 & \new_[54339]_ ;
  assign \new_[54343]_  = ~A299 & A298;
  assign \new_[54346]_  = A301 & A300;
  assign \new_[54347]_  = \new_[54346]_  & \new_[54343]_ ;
  assign \new_[54348]_  = \new_[54347]_  & \new_[54340]_ ;
  assign \new_[54352]_  = A167 & ~A168;
  assign \new_[54353]_  = ~A169 & \new_[54352]_ ;
  assign \new_[54356]_  = ~A199 & A166;
  assign \new_[54359]_  = A232 & A200;
  assign \new_[54360]_  = \new_[54359]_  & \new_[54356]_ ;
  assign \new_[54361]_  = \new_[54360]_  & \new_[54353]_ ;
  assign \new_[54365]_  = A266 & A265;
  assign \new_[54366]_  = A233 & \new_[54365]_ ;
  assign \new_[54369]_  = ~A299 & A298;
  assign \new_[54372]_  = A302 & A300;
  assign \new_[54373]_  = \new_[54372]_  & \new_[54369]_ ;
  assign \new_[54374]_  = \new_[54373]_  & \new_[54366]_ ;
  assign \new_[54378]_  = A167 & ~A168;
  assign \new_[54379]_  = ~A169 & \new_[54378]_ ;
  assign \new_[54382]_  = ~A199 & A166;
  assign \new_[54385]_  = A232 & A200;
  assign \new_[54386]_  = \new_[54385]_  & \new_[54382]_ ;
  assign \new_[54387]_  = \new_[54386]_  & \new_[54379]_ ;
  assign \new_[54391]_  = ~A266 & ~A265;
  assign \new_[54392]_  = A233 & \new_[54391]_ ;
  assign \new_[54395]_  = ~A299 & A298;
  assign \new_[54398]_  = A301 & A300;
  assign \new_[54399]_  = \new_[54398]_  & \new_[54395]_ ;
  assign \new_[54400]_  = \new_[54399]_  & \new_[54392]_ ;
  assign \new_[54404]_  = A167 & ~A168;
  assign \new_[54405]_  = ~A169 & \new_[54404]_ ;
  assign \new_[54408]_  = ~A199 & A166;
  assign \new_[54411]_  = A232 & A200;
  assign \new_[54412]_  = \new_[54411]_  & \new_[54408]_ ;
  assign \new_[54413]_  = \new_[54412]_  & \new_[54405]_ ;
  assign \new_[54417]_  = ~A266 & ~A265;
  assign \new_[54418]_  = A233 & \new_[54417]_ ;
  assign \new_[54421]_  = ~A299 & A298;
  assign \new_[54424]_  = A302 & A300;
  assign \new_[54425]_  = \new_[54424]_  & \new_[54421]_ ;
  assign \new_[54426]_  = \new_[54425]_  & \new_[54418]_ ;
  assign \new_[54430]_  = A167 & ~A168;
  assign \new_[54431]_  = ~A169 & \new_[54430]_ ;
  assign \new_[54434]_  = ~A199 & A166;
  assign \new_[54437]_  = ~A233 & A200;
  assign \new_[54438]_  = \new_[54437]_  & \new_[54434]_ ;
  assign \new_[54439]_  = \new_[54438]_  & \new_[54431]_ ;
  assign \new_[54443]_  = ~A266 & ~A236;
  assign \new_[54444]_  = ~A235 & \new_[54443]_ ;
  assign \new_[54447]_  = ~A269 & ~A268;
  assign \new_[54450]_  = A299 & ~A298;
  assign \new_[54451]_  = \new_[54450]_  & \new_[54447]_ ;
  assign \new_[54452]_  = \new_[54451]_  & \new_[54444]_ ;
  assign \new_[54456]_  = A167 & ~A168;
  assign \new_[54457]_  = ~A169 & \new_[54456]_ ;
  assign \new_[54460]_  = ~A199 & A166;
  assign \new_[54463]_  = ~A233 & A200;
  assign \new_[54464]_  = \new_[54463]_  & \new_[54460]_ ;
  assign \new_[54465]_  = \new_[54464]_  & \new_[54457]_ ;
  assign \new_[54469]_  = A266 & A265;
  assign \new_[54470]_  = ~A234 & \new_[54469]_ ;
  assign \new_[54473]_  = ~A299 & A298;
  assign \new_[54476]_  = A301 & A300;
  assign \new_[54477]_  = \new_[54476]_  & \new_[54473]_ ;
  assign \new_[54478]_  = \new_[54477]_  & \new_[54470]_ ;
  assign \new_[54482]_  = A167 & ~A168;
  assign \new_[54483]_  = ~A169 & \new_[54482]_ ;
  assign \new_[54486]_  = ~A199 & A166;
  assign \new_[54489]_  = ~A233 & A200;
  assign \new_[54490]_  = \new_[54489]_  & \new_[54486]_ ;
  assign \new_[54491]_  = \new_[54490]_  & \new_[54483]_ ;
  assign \new_[54495]_  = A266 & A265;
  assign \new_[54496]_  = ~A234 & \new_[54495]_ ;
  assign \new_[54499]_  = ~A299 & A298;
  assign \new_[54502]_  = A302 & A300;
  assign \new_[54503]_  = \new_[54502]_  & \new_[54499]_ ;
  assign \new_[54504]_  = \new_[54503]_  & \new_[54496]_ ;
  assign \new_[54508]_  = A167 & ~A168;
  assign \new_[54509]_  = ~A169 & \new_[54508]_ ;
  assign \new_[54512]_  = ~A199 & A166;
  assign \new_[54515]_  = ~A233 & A200;
  assign \new_[54516]_  = \new_[54515]_  & \new_[54512]_ ;
  assign \new_[54517]_  = \new_[54516]_  & \new_[54509]_ ;
  assign \new_[54521]_  = ~A267 & ~A266;
  assign \new_[54522]_  = ~A234 & \new_[54521]_ ;
  assign \new_[54525]_  = ~A299 & A298;
  assign \new_[54528]_  = A301 & A300;
  assign \new_[54529]_  = \new_[54528]_  & \new_[54525]_ ;
  assign \new_[54530]_  = \new_[54529]_  & \new_[54522]_ ;
  assign \new_[54534]_  = A167 & ~A168;
  assign \new_[54535]_  = ~A169 & \new_[54534]_ ;
  assign \new_[54538]_  = ~A199 & A166;
  assign \new_[54541]_  = ~A233 & A200;
  assign \new_[54542]_  = \new_[54541]_  & \new_[54538]_ ;
  assign \new_[54543]_  = \new_[54542]_  & \new_[54535]_ ;
  assign \new_[54547]_  = ~A267 & ~A266;
  assign \new_[54548]_  = ~A234 & \new_[54547]_ ;
  assign \new_[54551]_  = ~A299 & A298;
  assign \new_[54554]_  = A302 & A300;
  assign \new_[54555]_  = \new_[54554]_  & \new_[54551]_ ;
  assign \new_[54556]_  = \new_[54555]_  & \new_[54548]_ ;
  assign \new_[54560]_  = A167 & ~A168;
  assign \new_[54561]_  = ~A169 & \new_[54560]_ ;
  assign \new_[54564]_  = ~A199 & A166;
  assign \new_[54567]_  = ~A233 & A200;
  assign \new_[54568]_  = \new_[54567]_  & \new_[54564]_ ;
  assign \new_[54569]_  = \new_[54568]_  & \new_[54561]_ ;
  assign \new_[54573]_  = ~A266 & ~A265;
  assign \new_[54574]_  = ~A234 & \new_[54573]_ ;
  assign \new_[54577]_  = ~A299 & A298;
  assign \new_[54580]_  = A301 & A300;
  assign \new_[54581]_  = \new_[54580]_  & \new_[54577]_ ;
  assign \new_[54582]_  = \new_[54581]_  & \new_[54574]_ ;
  assign \new_[54586]_  = A167 & ~A168;
  assign \new_[54587]_  = ~A169 & \new_[54586]_ ;
  assign \new_[54590]_  = ~A199 & A166;
  assign \new_[54593]_  = ~A233 & A200;
  assign \new_[54594]_  = \new_[54593]_  & \new_[54590]_ ;
  assign \new_[54595]_  = \new_[54594]_  & \new_[54587]_ ;
  assign \new_[54599]_  = ~A266 & ~A265;
  assign \new_[54600]_  = ~A234 & \new_[54599]_ ;
  assign \new_[54603]_  = ~A299 & A298;
  assign \new_[54606]_  = A302 & A300;
  assign \new_[54607]_  = \new_[54606]_  & \new_[54603]_ ;
  assign \new_[54608]_  = \new_[54607]_  & \new_[54600]_ ;
  assign \new_[54612]_  = A167 & ~A168;
  assign \new_[54613]_  = ~A169 & \new_[54612]_ ;
  assign \new_[54616]_  = ~A199 & A166;
  assign \new_[54619]_  = A232 & A200;
  assign \new_[54620]_  = \new_[54619]_  & \new_[54616]_ ;
  assign \new_[54621]_  = \new_[54620]_  & \new_[54613]_ ;
  assign \new_[54625]_  = A235 & A234;
  assign \new_[54626]_  = ~A233 & \new_[54625]_ ;
  assign \new_[54629]_  = ~A266 & A265;
  assign \new_[54632]_  = A268 & A267;
  assign \new_[54633]_  = \new_[54632]_  & \new_[54629]_ ;
  assign \new_[54634]_  = \new_[54633]_  & \new_[54626]_ ;
  assign \new_[54638]_  = A167 & ~A168;
  assign \new_[54639]_  = ~A169 & \new_[54638]_ ;
  assign \new_[54642]_  = ~A199 & A166;
  assign \new_[54645]_  = A232 & A200;
  assign \new_[54646]_  = \new_[54645]_  & \new_[54642]_ ;
  assign \new_[54647]_  = \new_[54646]_  & \new_[54639]_ ;
  assign \new_[54651]_  = A235 & A234;
  assign \new_[54652]_  = ~A233 & \new_[54651]_ ;
  assign \new_[54655]_  = ~A266 & A265;
  assign \new_[54658]_  = A269 & A267;
  assign \new_[54659]_  = \new_[54658]_  & \new_[54655]_ ;
  assign \new_[54660]_  = \new_[54659]_  & \new_[54652]_ ;
  assign \new_[54664]_  = A167 & ~A168;
  assign \new_[54665]_  = ~A169 & \new_[54664]_ ;
  assign \new_[54668]_  = ~A199 & A166;
  assign \new_[54671]_  = A232 & A200;
  assign \new_[54672]_  = \new_[54671]_  & \new_[54668]_ ;
  assign \new_[54673]_  = \new_[54672]_  & \new_[54665]_ ;
  assign \new_[54677]_  = A236 & A234;
  assign \new_[54678]_  = ~A233 & \new_[54677]_ ;
  assign \new_[54681]_  = ~A266 & A265;
  assign \new_[54684]_  = A268 & A267;
  assign \new_[54685]_  = \new_[54684]_  & \new_[54681]_ ;
  assign \new_[54686]_  = \new_[54685]_  & \new_[54678]_ ;
  assign \new_[54690]_  = A167 & ~A168;
  assign \new_[54691]_  = ~A169 & \new_[54690]_ ;
  assign \new_[54694]_  = ~A199 & A166;
  assign \new_[54697]_  = A232 & A200;
  assign \new_[54698]_  = \new_[54697]_  & \new_[54694]_ ;
  assign \new_[54699]_  = \new_[54698]_  & \new_[54691]_ ;
  assign \new_[54703]_  = A236 & A234;
  assign \new_[54704]_  = ~A233 & \new_[54703]_ ;
  assign \new_[54707]_  = ~A266 & A265;
  assign \new_[54710]_  = A269 & A267;
  assign \new_[54711]_  = \new_[54710]_  & \new_[54707]_ ;
  assign \new_[54712]_  = \new_[54711]_  & \new_[54704]_ ;
  assign \new_[54716]_  = A167 & ~A168;
  assign \new_[54717]_  = ~A169 & \new_[54716]_ ;
  assign \new_[54720]_  = ~A199 & A166;
  assign \new_[54723]_  = ~A232 & A200;
  assign \new_[54724]_  = \new_[54723]_  & \new_[54720]_ ;
  assign \new_[54725]_  = \new_[54724]_  & \new_[54717]_ ;
  assign \new_[54729]_  = A266 & A265;
  assign \new_[54730]_  = ~A233 & \new_[54729]_ ;
  assign \new_[54733]_  = ~A299 & A298;
  assign \new_[54736]_  = A301 & A300;
  assign \new_[54737]_  = \new_[54736]_  & \new_[54733]_ ;
  assign \new_[54738]_  = \new_[54737]_  & \new_[54730]_ ;
  assign \new_[54742]_  = A167 & ~A168;
  assign \new_[54743]_  = ~A169 & \new_[54742]_ ;
  assign \new_[54746]_  = ~A199 & A166;
  assign \new_[54749]_  = ~A232 & A200;
  assign \new_[54750]_  = \new_[54749]_  & \new_[54746]_ ;
  assign \new_[54751]_  = \new_[54750]_  & \new_[54743]_ ;
  assign \new_[54755]_  = A266 & A265;
  assign \new_[54756]_  = ~A233 & \new_[54755]_ ;
  assign \new_[54759]_  = ~A299 & A298;
  assign \new_[54762]_  = A302 & A300;
  assign \new_[54763]_  = \new_[54762]_  & \new_[54759]_ ;
  assign \new_[54764]_  = \new_[54763]_  & \new_[54756]_ ;
  assign \new_[54768]_  = A167 & ~A168;
  assign \new_[54769]_  = ~A169 & \new_[54768]_ ;
  assign \new_[54772]_  = ~A199 & A166;
  assign \new_[54775]_  = ~A232 & A200;
  assign \new_[54776]_  = \new_[54775]_  & \new_[54772]_ ;
  assign \new_[54777]_  = \new_[54776]_  & \new_[54769]_ ;
  assign \new_[54781]_  = ~A267 & ~A266;
  assign \new_[54782]_  = ~A233 & \new_[54781]_ ;
  assign \new_[54785]_  = ~A299 & A298;
  assign \new_[54788]_  = A301 & A300;
  assign \new_[54789]_  = \new_[54788]_  & \new_[54785]_ ;
  assign \new_[54790]_  = \new_[54789]_  & \new_[54782]_ ;
  assign \new_[54794]_  = A167 & ~A168;
  assign \new_[54795]_  = ~A169 & \new_[54794]_ ;
  assign \new_[54798]_  = ~A199 & A166;
  assign \new_[54801]_  = ~A232 & A200;
  assign \new_[54802]_  = \new_[54801]_  & \new_[54798]_ ;
  assign \new_[54803]_  = \new_[54802]_  & \new_[54795]_ ;
  assign \new_[54807]_  = ~A267 & ~A266;
  assign \new_[54808]_  = ~A233 & \new_[54807]_ ;
  assign \new_[54811]_  = ~A299 & A298;
  assign \new_[54814]_  = A302 & A300;
  assign \new_[54815]_  = \new_[54814]_  & \new_[54811]_ ;
  assign \new_[54816]_  = \new_[54815]_  & \new_[54808]_ ;
  assign \new_[54820]_  = A167 & ~A168;
  assign \new_[54821]_  = ~A169 & \new_[54820]_ ;
  assign \new_[54824]_  = ~A199 & A166;
  assign \new_[54827]_  = ~A232 & A200;
  assign \new_[54828]_  = \new_[54827]_  & \new_[54824]_ ;
  assign \new_[54829]_  = \new_[54828]_  & \new_[54821]_ ;
  assign \new_[54833]_  = ~A266 & ~A265;
  assign \new_[54834]_  = ~A233 & \new_[54833]_ ;
  assign \new_[54837]_  = ~A299 & A298;
  assign \new_[54840]_  = A301 & A300;
  assign \new_[54841]_  = \new_[54840]_  & \new_[54837]_ ;
  assign \new_[54842]_  = \new_[54841]_  & \new_[54834]_ ;
  assign \new_[54846]_  = A167 & ~A168;
  assign \new_[54847]_  = ~A169 & \new_[54846]_ ;
  assign \new_[54850]_  = ~A199 & A166;
  assign \new_[54853]_  = ~A232 & A200;
  assign \new_[54854]_  = \new_[54853]_  & \new_[54850]_ ;
  assign \new_[54855]_  = \new_[54854]_  & \new_[54847]_ ;
  assign \new_[54859]_  = ~A266 & ~A265;
  assign \new_[54860]_  = ~A233 & \new_[54859]_ ;
  assign \new_[54863]_  = ~A299 & A298;
  assign \new_[54866]_  = A302 & A300;
  assign \new_[54867]_  = \new_[54866]_  & \new_[54863]_ ;
  assign \new_[54868]_  = \new_[54867]_  & \new_[54860]_ ;
  assign \new_[54872]_  = A167 & ~A168;
  assign \new_[54873]_  = ~A169 & \new_[54872]_ ;
  assign \new_[54876]_  = A199 & A166;
  assign \new_[54879]_  = A201 & ~A200;
  assign \new_[54880]_  = \new_[54879]_  & \new_[54876]_ ;
  assign \new_[54881]_  = \new_[54880]_  & \new_[54873]_ ;
  assign \new_[54885]_  = A233 & A232;
  assign \new_[54886]_  = A202 & \new_[54885]_ ;
  assign \new_[54889]_  = ~A267 & A265;
  assign \new_[54892]_  = A299 & ~A298;
  assign \new_[54893]_  = \new_[54892]_  & \new_[54889]_ ;
  assign \new_[54894]_  = \new_[54893]_  & \new_[54886]_ ;
  assign \new_[54898]_  = A167 & ~A168;
  assign \new_[54899]_  = ~A169 & \new_[54898]_ ;
  assign \new_[54902]_  = A199 & A166;
  assign \new_[54905]_  = A201 & ~A200;
  assign \new_[54906]_  = \new_[54905]_  & \new_[54902]_ ;
  assign \new_[54907]_  = \new_[54906]_  & \new_[54899]_ ;
  assign \new_[54911]_  = A233 & A232;
  assign \new_[54912]_  = A202 & \new_[54911]_ ;
  assign \new_[54915]_  = A266 & A265;
  assign \new_[54918]_  = A299 & ~A298;
  assign \new_[54919]_  = \new_[54918]_  & \new_[54915]_ ;
  assign \new_[54920]_  = \new_[54919]_  & \new_[54912]_ ;
  assign \new_[54924]_  = A167 & ~A168;
  assign \new_[54925]_  = ~A169 & \new_[54924]_ ;
  assign \new_[54928]_  = A199 & A166;
  assign \new_[54931]_  = A201 & ~A200;
  assign \new_[54932]_  = \new_[54931]_  & \new_[54928]_ ;
  assign \new_[54933]_  = \new_[54932]_  & \new_[54925]_ ;
  assign \new_[54937]_  = A233 & A232;
  assign \new_[54938]_  = A202 & \new_[54937]_ ;
  assign \new_[54941]_  = ~A266 & ~A265;
  assign \new_[54944]_  = A299 & ~A298;
  assign \new_[54945]_  = \new_[54944]_  & \new_[54941]_ ;
  assign \new_[54946]_  = \new_[54945]_  & \new_[54938]_ ;
  assign \new_[54950]_  = A167 & ~A168;
  assign \new_[54951]_  = ~A169 & \new_[54950]_ ;
  assign \new_[54954]_  = A199 & A166;
  assign \new_[54957]_  = A201 & ~A200;
  assign \new_[54958]_  = \new_[54957]_  & \new_[54954]_ ;
  assign \new_[54959]_  = \new_[54958]_  & \new_[54951]_ ;
  assign \new_[54963]_  = A233 & ~A232;
  assign \new_[54964]_  = A202 & \new_[54963]_ ;
  assign \new_[54967]_  = ~A266 & A265;
  assign \new_[54970]_  = A268 & A267;
  assign \new_[54971]_  = \new_[54970]_  & \new_[54967]_ ;
  assign \new_[54972]_  = \new_[54971]_  & \new_[54964]_ ;
  assign \new_[54976]_  = A167 & ~A168;
  assign \new_[54977]_  = ~A169 & \new_[54976]_ ;
  assign \new_[54980]_  = A199 & A166;
  assign \new_[54983]_  = A201 & ~A200;
  assign \new_[54984]_  = \new_[54983]_  & \new_[54980]_ ;
  assign \new_[54985]_  = \new_[54984]_  & \new_[54977]_ ;
  assign \new_[54989]_  = A233 & ~A232;
  assign \new_[54990]_  = A202 & \new_[54989]_ ;
  assign \new_[54993]_  = ~A266 & A265;
  assign \new_[54996]_  = A269 & A267;
  assign \new_[54997]_  = \new_[54996]_  & \new_[54993]_ ;
  assign \new_[54998]_  = \new_[54997]_  & \new_[54990]_ ;
  assign \new_[55002]_  = A167 & ~A168;
  assign \new_[55003]_  = ~A169 & \new_[55002]_ ;
  assign \new_[55006]_  = A199 & A166;
  assign \new_[55009]_  = A201 & ~A200;
  assign \new_[55010]_  = \new_[55009]_  & \new_[55006]_ ;
  assign \new_[55011]_  = \new_[55010]_  & \new_[55003]_ ;
  assign \new_[55015]_  = ~A234 & ~A233;
  assign \new_[55016]_  = A202 & \new_[55015]_ ;
  assign \new_[55019]_  = A266 & A265;
  assign \new_[55022]_  = A299 & ~A298;
  assign \new_[55023]_  = \new_[55022]_  & \new_[55019]_ ;
  assign \new_[55024]_  = \new_[55023]_  & \new_[55016]_ ;
  assign \new_[55028]_  = A167 & ~A168;
  assign \new_[55029]_  = ~A169 & \new_[55028]_ ;
  assign \new_[55032]_  = A199 & A166;
  assign \new_[55035]_  = A201 & ~A200;
  assign \new_[55036]_  = \new_[55035]_  & \new_[55032]_ ;
  assign \new_[55037]_  = \new_[55036]_  & \new_[55029]_ ;
  assign \new_[55041]_  = ~A234 & ~A233;
  assign \new_[55042]_  = A202 & \new_[55041]_ ;
  assign \new_[55045]_  = ~A267 & ~A266;
  assign \new_[55048]_  = A299 & ~A298;
  assign \new_[55049]_  = \new_[55048]_  & \new_[55045]_ ;
  assign \new_[55050]_  = \new_[55049]_  & \new_[55042]_ ;
  assign \new_[55054]_  = A167 & ~A168;
  assign \new_[55055]_  = ~A169 & \new_[55054]_ ;
  assign \new_[55058]_  = A199 & A166;
  assign \new_[55061]_  = A201 & ~A200;
  assign \new_[55062]_  = \new_[55061]_  & \new_[55058]_ ;
  assign \new_[55063]_  = \new_[55062]_  & \new_[55055]_ ;
  assign \new_[55067]_  = ~A234 & ~A233;
  assign \new_[55068]_  = A202 & \new_[55067]_ ;
  assign \new_[55071]_  = ~A266 & ~A265;
  assign \new_[55074]_  = A299 & ~A298;
  assign \new_[55075]_  = \new_[55074]_  & \new_[55071]_ ;
  assign \new_[55076]_  = \new_[55075]_  & \new_[55068]_ ;
  assign \new_[55080]_  = A167 & ~A168;
  assign \new_[55081]_  = ~A169 & \new_[55080]_ ;
  assign \new_[55084]_  = A199 & A166;
  assign \new_[55087]_  = A201 & ~A200;
  assign \new_[55088]_  = \new_[55087]_  & \new_[55084]_ ;
  assign \new_[55089]_  = \new_[55088]_  & \new_[55081]_ ;
  assign \new_[55093]_  = ~A233 & A232;
  assign \new_[55094]_  = A202 & \new_[55093]_ ;
  assign \new_[55097]_  = A235 & A234;
  assign \new_[55100]_  = ~A300 & A298;
  assign \new_[55101]_  = \new_[55100]_  & \new_[55097]_ ;
  assign \new_[55102]_  = \new_[55101]_  & \new_[55094]_ ;
  assign \new_[55106]_  = A167 & ~A168;
  assign \new_[55107]_  = ~A169 & \new_[55106]_ ;
  assign \new_[55110]_  = A199 & A166;
  assign \new_[55113]_  = A201 & ~A200;
  assign \new_[55114]_  = \new_[55113]_  & \new_[55110]_ ;
  assign \new_[55115]_  = \new_[55114]_  & \new_[55107]_ ;
  assign \new_[55119]_  = ~A233 & A232;
  assign \new_[55120]_  = A202 & \new_[55119]_ ;
  assign \new_[55123]_  = A235 & A234;
  assign \new_[55126]_  = A299 & A298;
  assign \new_[55127]_  = \new_[55126]_  & \new_[55123]_ ;
  assign \new_[55128]_  = \new_[55127]_  & \new_[55120]_ ;
  assign \new_[55132]_  = A167 & ~A168;
  assign \new_[55133]_  = ~A169 & \new_[55132]_ ;
  assign \new_[55136]_  = A199 & A166;
  assign \new_[55139]_  = A201 & ~A200;
  assign \new_[55140]_  = \new_[55139]_  & \new_[55136]_ ;
  assign \new_[55141]_  = \new_[55140]_  & \new_[55133]_ ;
  assign \new_[55145]_  = ~A233 & A232;
  assign \new_[55146]_  = A202 & \new_[55145]_ ;
  assign \new_[55149]_  = A235 & A234;
  assign \new_[55152]_  = ~A299 & ~A298;
  assign \new_[55153]_  = \new_[55152]_  & \new_[55149]_ ;
  assign \new_[55154]_  = \new_[55153]_  & \new_[55146]_ ;
  assign \new_[55158]_  = A167 & ~A168;
  assign \new_[55159]_  = ~A169 & \new_[55158]_ ;
  assign \new_[55162]_  = A199 & A166;
  assign \new_[55165]_  = A201 & ~A200;
  assign \new_[55166]_  = \new_[55165]_  & \new_[55162]_ ;
  assign \new_[55167]_  = \new_[55166]_  & \new_[55159]_ ;
  assign \new_[55171]_  = ~A233 & A232;
  assign \new_[55172]_  = A202 & \new_[55171]_ ;
  assign \new_[55175]_  = A235 & A234;
  assign \new_[55178]_  = A266 & ~A265;
  assign \new_[55179]_  = \new_[55178]_  & \new_[55175]_ ;
  assign \new_[55180]_  = \new_[55179]_  & \new_[55172]_ ;
  assign \new_[55184]_  = A167 & ~A168;
  assign \new_[55185]_  = ~A169 & \new_[55184]_ ;
  assign \new_[55188]_  = A199 & A166;
  assign \new_[55191]_  = A201 & ~A200;
  assign \new_[55192]_  = \new_[55191]_  & \new_[55188]_ ;
  assign \new_[55193]_  = \new_[55192]_  & \new_[55185]_ ;
  assign \new_[55197]_  = ~A233 & A232;
  assign \new_[55198]_  = A202 & \new_[55197]_ ;
  assign \new_[55201]_  = A236 & A234;
  assign \new_[55204]_  = ~A300 & A298;
  assign \new_[55205]_  = \new_[55204]_  & \new_[55201]_ ;
  assign \new_[55206]_  = \new_[55205]_  & \new_[55198]_ ;
  assign \new_[55210]_  = A167 & ~A168;
  assign \new_[55211]_  = ~A169 & \new_[55210]_ ;
  assign \new_[55214]_  = A199 & A166;
  assign \new_[55217]_  = A201 & ~A200;
  assign \new_[55218]_  = \new_[55217]_  & \new_[55214]_ ;
  assign \new_[55219]_  = \new_[55218]_  & \new_[55211]_ ;
  assign \new_[55223]_  = ~A233 & A232;
  assign \new_[55224]_  = A202 & \new_[55223]_ ;
  assign \new_[55227]_  = A236 & A234;
  assign \new_[55230]_  = A299 & A298;
  assign \new_[55231]_  = \new_[55230]_  & \new_[55227]_ ;
  assign \new_[55232]_  = \new_[55231]_  & \new_[55224]_ ;
  assign \new_[55236]_  = A167 & ~A168;
  assign \new_[55237]_  = ~A169 & \new_[55236]_ ;
  assign \new_[55240]_  = A199 & A166;
  assign \new_[55243]_  = A201 & ~A200;
  assign \new_[55244]_  = \new_[55243]_  & \new_[55240]_ ;
  assign \new_[55245]_  = \new_[55244]_  & \new_[55237]_ ;
  assign \new_[55249]_  = ~A233 & A232;
  assign \new_[55250]_  = A202 & \new_[55249]_ ;
  assign \new_[55253]_  = A236 & A234;
  assign \new_[55256]_  = ~A299 & ~A298;
  assign \new_[55257]_  = \new_[55256]_  & \new_[55253]_ ;
  assign \new_[55258]_  = \new_[55257]_  & \new_[55250]_ ;
  assign \new_[55262]_  = A167 & ~A168;
  assign \new_[55263]_  = ~A169 & \new_[55262]_ ;
  assign \new_[55266]_  = A199 & A166;
  assign \new_[55269]_  = A201 & ~A200;
  assign \new_[55270]_  = \new_[55269]_  & \new_[55266]_ ;
  assign \new_[55271]_  = \new_[55270]_  & \new_[55263]_ ;
  assign \new_[55275]_  = ~A233 & A232;
  assign \new_[55276]_  = A202 & \new_[55275]_ ;
  assign \new_[55279]_  = A236 & A234;
  assign \new_[55282]_  = A266 & ~A265;
  assign \new_[55283]_  = \new_[55282]_  & \new_[55279]_ ;
  assign \new_[55284]_  = \new_[55283]_  & \new_[55276]_ ;
  assign \new_[55288]_  = A167 & ~A168;
  assign \new_[55289]_  = ~A169 & \new_[55288]_ ;
  assign \new_[55292]_  = A199 & A166;
  assign \new_[55295]_  = A201 & ~A200;
  assign \new_[55296]_  = \new_[55295]_  & \new_[55292]_ ;
  assign \new_[55297]_  = \new_[55296]_  & \new_[55289]_ ;
  assign \new_[55301]_  = ~A233 & ~A232;
  assign \new_[55302]_  = A202 & \new_[55301]_ ;
  assign \new_[55305]_  = A266 & A265;
  assign \new_[55308]_  = A299 & ~A298;
  assign \new_[55309]_  = \new_[55308]_  & \new_[55305]_ ;
  assign \new_[55310]_  = \new_[55309]_  & \new_[55302]_ ;
  assign \new_[55314]_  = A167 & ~A168;
  assign \new_[55315]_  = ~A169 & \new_[55314]_ ;
  assign \new_[55318]_  = A199 & A166;
  assign \new_[55321]_  = A201 & ~A200;
  assign \new_[55322]_  = \new_[55321]_  & \new_[55318]_ ;
  assign \new_[55323]_  = \new_[55322]_  & \new_[55315]_ ;
  assign \new_[55327]_  = ~A233 & ~A232;
  assign \new_[55328]_  = A202 & \new_[55327]_ ;
  assign \new_[55331]_  = ~A267 & ~A266;
  assign \new_[55334]_  = A299 & ~A298;
  assign \new_[55335]_  = \new_[55334]_  & \new_[55331]_ ;
  assign \new_[55336]_  = \new_[55335]_  & \new_[55328]_ ;
  assign \new_[55340]_  = A167 & ~A168;
  assign \new_[55341]_  = ~A169 & \new_[55340]_ ;
  assign \new_[55344]_  = A199 & A166;
  assign \new_[55347]_  = A201 & ~A200;
  assign \new_[55348]_  = \new_[55347]_  & \new_[55344]_ ;
  assign \new_[55349]_  = \new_[55348]_  & \new_[55341]_ ;
  assign \new_[55353]_  = ~A233 & ~A232;
  assign \new_[55354]_  = A202 & \new_[55353]_ ;
  assign \new_[55357]_  = ~A266 & ~A265;
  assign \new_[55360]_  = A299 & ~A298;
  assign \new_[55361]_  = \new_[55360]_  & \new_[55357]_ ;
  assign \new_[55362]_  = \new_[55361]_  & \new_[55354]_ ;
  assign \new_[55366]_  = A167 & ~A168;
  assign \new_[55367]_  = ~A169 & \new_[55366]_ ;
  assign \new_[55370]_  = A199 & A166;
  assign \new_[55373]_  = A201 & ~A200;
  assign \new_[55374]_  = \new_[55373]_  & \new_[55370]_ ;
  assign \new_[55375]_  = \new_[55374]_  & \new_[55367]_ ;
  assign \new_[55379]_  = A233 & A232;
  assign \new_[55380]_  = A203 & \new_[55379]_ ;
  assign \new_[55383]_  = ~A267 & A265;
  assign \new_[55386]_  = A299 & ~A298;
  assign \new_[55387]_  = \new_[55386]_  & \new_[55383]_ ;
  assign \new_[55388]_  = \new_[55387]_  & \new_[55380]_ ;
  assign \new_[55392]_  = A167 & ~A168;
  assign \new_[55393]_  = ~A169 & \new_[55392]_ ;
  assign \new_[55396]_  = A199 & A166;
  assign \new_[55399]_  = A201 & ~A200;
  assign \new_[55400]_  = \new_[55399]_  & \new_[55396]_ ;
  assign \new_[55401]_  = \new_[55400]_  & \new_[55393]_ ;
  assign \new_[55405]_  = A233 & A232;
  assign \new_[55406]_  = A203 & \new_[55405]_ ;
  assign \new_[55409]_  = A266 & A265;
  assign \new_[55412]_  = A299 & ~A298;
  assign \new_[55413]_  = \new_[55412]_  & \new_[55409]_ ;
  assign \new_[55414]_  = \new_[55413]_  & \new_[55406]_ ;
  assign \new_[55418]_  = A167 & ~A168;
  assign \new_[55419]_  = ~A169 & \new_[55418]_ ;
  assign \new_[55422]_  = A199 & A166;
  assign \new_[55425]_  = A201 & ~A200;
  assign \new_[55426]_  = \new_[55425]_  & \new_[55422]_ ;
  assign \new_[55427]_  = \new_[55426]_  & \new_[55419]_ ;
  assign \new_[55431]_  = A233 & A232;
  assign \new_[55432]_  = A203 & \new_[55431]_ ;
  assign \new_[55435]_  = ~A266 & ~A265;
  assign \new_[55438]_  = A299 & ~A298;
  assign \new_[55439]_  = \new_[55438]_  & \new_[55435]_ ;
  assign \new_[55440]_  = \new_[55439]_  & \new_[55432]_ ;
  assign \new_[55444]_  = A167 & ~A168;
  assign \new_[55445]_  = ~A169 & \new_[55444]_ ;
  assign \new_[55448]_  = A199 & A166;
  assign \new_[55451]_  = A201 & ~A200;
  assign \new_[55452]_  = \new_[55451]_  & \new_[55448]_ ;
  assign \new_[55453]_  = \new_[55452]_  & \new_[55445]_ ;
  assign \new_[55457]_  = A233 & ~A232;
  assign \new_[55458]_  = A203 & \new_[55457]_ ;
  assign \new_[55461]_  = ~A266 & A265;
  assign \new_[55464]_  = A268 & A267;
  assign \new_[55465]_  = \new_[55464]_  & \new_[55461]_ ;
  assign \new_[55466]_  = \new_[55465]_  & \new_[55458]_ ;
  assign \new_[55470]_  = A167 & ~A168;
  assign \new_[55471]_  = ~A169 & \new_[55470]_ ;
  assign \new_[55474]_  = A199 & A166;
  assign \new_[55477]_  = A201 & ~A200;
  assign \new_[55478]_  = \new_[55477]_  & \new_[55474]_ ;
  assign \new_[55479]_  = \new_[55478]_  & \new_[55471]_ ;
  assign \new_[55483]_  = A233 & ~A232;
  assign \new_[55484]_  = A203 & \new_[55483]_ ;
  assign \new_[55487]_  = ~A266 & A265;
  assign \new_[55490]_  = A269 & A267;
  assign \new_[55491]_  = \new_[55490]_  & \new_[55487]_ ;
  assign \new_[55492]_  = \new_[55491]_  & \new_[55484]_ ;
  assign \new_[55496]_  = A167 & ~A168;
  assign \new_[55497]_  = ~A169 & \new_[55496]_ ;
  assign \new_[55500]_  = A199 & A166;
  assign \new_[55503]_  = A201 & ~A200;
  assign \new_[55504]_  = \new_[55503]_  & \new_[55500]_ ;
  assign \new_[55505]_  = \new_[55504]_  & \new_[55497]_ ;
  assign \new_[55509]_  = ~A234 & ~A233;
  assign \new_[55510]_  = A203 & \new_[55509]_ ;
  assign \new_[55513]_  = A266 & A265;
  assign \new_[55516]_  = A299 & ~A298;
  assign \new_[55517]_  = \new_[55516]_  & \new_[55513]_ ;
  assign \new_[55518]_  = \new_[55517]_  & \new_[55510]_ ;
  assign \new_[55522]_  = A167 & ~A168;
  assign \new_[55523]_  = ~A169 & \new_[55522]_ ;
  assign \new_[55526]_  = A199 & A166;
  assign \new_[55529]_  = A201 & ~A200;
  assign \new_[55530]_  = \new_[55529]_  & \new_[55526]_ ;
  assign \new_[55531]_  = \new_[55530]_  & \new_[55523]_ ;
  assign \new_[55535]_  = ~A234 & ~A233;
  assign \new_[55536]_  = A203 & \new_[55535]_ ;
  assign \new_[55539]_  = ~A267 & ~A266;
  assign \new_[55542]_  = A299 & ~A298;
  assign \new_[55543]_  = \new_[55542]_  & \new_[55539]_ ;
  assign \new_[55544]_  = \new_[55543]_  & \new_[55536]_ ;
  assign \new_[55548]_  = A167 & ~A168;
  assign \new_[55549]_  = ~A169 & \new_[55548]_ ;
  assign \new_[55552]_  = A199 & A166;
  assign \new_[55555]_  = A201 & ~A200;
  assign \new_[55556]_  = \new_[55555]_  & \new_[55552]_ ;
  assign \new_[55557]_  = \new_[55556]_  & \new_[55549]_ ;
  assign \new_[55561]_  = ~A234 & ~A233;
  assign \new_[55562]_  = A203 & \new_[55561]_ ;
  assign \new_[55565]_  = ~A266 & ~A265;
  assign \new_[55568]_  = A299 & ~A298;
  assign \new_[55569]_  = \new_[55568]_  & \new_[55565]_ ;
  assign \new_[55570]_  = \new_[55569]_  & \new_[55562]_ ;
  assign \new_[55574]_  = A167 & ~A168;
  assign \new_[55575]_  = ~A169 & \new_[55574]_ ;
  assign \new_[55578]_  = A199 & A166;
  assign \new_[55581]_  = A201 & ~A200;
  assign \new_[55582]_  = \new_[55581]_  & \new_[55578]_ ;
  assign \new_[55583]_  = \new_[55582]_  & \new_[55575]_ ;
  assign \new_[55587]_  = ~A233 & A232;
  assign \new_[55588]_  = A203 & \new_[55587]_ ;
  assign \new_[55591]_  = A235 & A234;
  assign \new_[55594]_  = ~A300 & A298;
  assign \new_[55595]_  = \new_[55594]_  & \new_[55591]_ ;
  assign \new_[55596]_  = \new_[55595]_  & \new_[55588]_ ;
  assign \new_[55600]_  = A167 & ~A168;
  assign \new_[55601]_  = ~A169 & \new_[55600]_ ;
  assign \new_[55604]_  = A199 & A166;
  assign \new_[55607]_  = A201 & ~A200;
  assign \new_[55608]_  = \new_[55607]_  & \new_[55604]_ ;
  assign \new_[55609]_  = \new_[55608]_  & \new_[55601]_ ;
  assign \new_[55613]_  = ~A233 & A232;
  assign \new_[55614]_  = A203 & \new_[55613]_ ;
  assign \new_[55617]_  = A235 & A234;
  assign \new_[55620]_  = A299 & A298;
  assign \new_[55621]_  = \new_[55620]_  & \new_[55617]_ ;
  assign \new_[55622]_  = \new_[55621]_  & \new_[55614]_ ;
  assign \new_[55626]_  = A167 & ~A168;
  assign \new_[55627]_  = ~A169 & \new_[55626]_ ;
  assign \new_[55630]_  = A199 & A166;
  assign \new_[55633]_  = A201 & ~A200;
  assign \new_[55634]_  = \new_[55633]_  & \new_[55630]_ ;
  assign \new_[55635]_  = \new_[55634]_  & \new_[55627]_ ;
  assign \new_[55639]_  = ~A233 & A232;
  assign \new_[55640]_  = A203 & \new_[55639]_ ;
  assign \new_[55643]_  = A235 & A234;
  assign \new_[55646]_  = ~A299 & ~A298;
  assign \new_[55647]_  = \new_[55646]_  & \new_[55643]_ ;
  assign \new_[55648]_  = \new_[55647]_  & \new_[55640]_ ;
  assign \new_[55652]_  = A167 & ~A168;
  assign \new_[55653]_  = ~A169 & \new_[55652]_ ;
  assign \new_[55656]_  = A199 & A166;
  assign \new_[55659]_  = A201 & ~A200;
  assign \new_[55660]_  = \new_[55659]_  & \new_[55656]_ ;
  assign \new_[55661]_  = \new_[55660]_  & \new_[55653]_ ;
  assign \new_[55665]_  = ~A233 & A232;
  assign \new_[55666]_  = A203 & \new_[55665]_ ;
  assign \new_[55669]_  = A235 & A234;
  assign \new_[55672]_  = A266 & ~A265;
  assign \new_[55673]_  = \new_[55672]_  & \new_[55669]_ ;
  assign \new_[55674]_  = \new_[55673]_  & \new_[55666]_ ;
  assign \new_[55678]_  = A167 & ~A168;
  assign \new_[55679]_  = ~A169 & \new_[55678]_ ;
  assign \new_[55682]_  = A199 & A166;
  assign \new_[55685]_  = A201 & ~A200;
  assign \new_[55686]_  = \new_[55685]_  & \new_[55682]_ ;
  assign \new_[55687]_  = \new_[55686]_  & \new_[55679]_ ;
  assign \new_[55691]_  = ~A233 & A232;
  assign \new_[55692]_  = A203 & \new_[55691]_ ;
  assign \new_[55695]_  = A236 & A234;
  assign \new_[55698]_  = ~A300 & A298;
  assign \new_[55699]_  = \new_[55698]_  & \new_[55695]_ ;
  assign \new_[55700]_  = \new_[55699]_  & \new_[55692]_ ;
  assign \new_[55704]_  = A167 & ~A168;
  assign \new_[55705]_  = ~A169 & \new_[55704]_ ;
  assign \new_[55708]_  = A199 & A166;
  assign \new_[55711]_  = A201 & ~A200;
  assign \new_[55712]_  = \new_[55711]_  & \new_[55708]_ ;
  assign \new_[55713]_  = \new_[55712]_  & \new_[55705]_ ;
  assign \new_[55717]_  = ~A233 & A232;
  assign \new_[55718]_  = A203 & \new_[55717]_ ;
  assign \new_[55721]_  = A236 & A234;
  assign \new_[55724]_  = A299 & A298;
  assign \new_[55725]_  = \new_[55724]_  & \new_[55721]_ ;
  assign \new_[55726]_  = \new_[55725]_  & \new_[55718]_ ;
  assign \new_[55730]_  = A167 & ~A168;
  assign \new_[55731]_  = ~A169 & \new_[55730]_ ;
  assign \new_[55734]_  = A199 & A166;
  assign \new_[55737]_  = A201 & ~A200;
  assign \new_[55738]_  = \new_[55737]_  & \new_[55734]_ ;
  assign \new_[55739]_  = \new_[55738]_  & \new_[55731]_ ;
  assign \new_[55743]_  = ~A233 & A232;
  assign \new_[55744]_  = A203 & \new_[55743]_ ;
  assign \new_[55747]_  = A236 & A234;
  assign \new_[55750]_  = ~A299 & ~A298;
  assign \new_[55751]_  = \new_[55750]_  & \new_[55747]_ ;
  assign \new_[55752]_  = \new_[55751]_  & \new_[55744]_ ;
  assign \new_[55756]_  = A167 & ~A168;
  assign \new_[55757]_  = ~A169 & \new_[55756]_ ;
  assign \new_[55760]_  = A199 & A166;
  assign \new_[55763]_  = A201 & ~A200;
  assign \new_[55764]_  = \new_[55763]_  & \new_[55760]_ ;
  assign \new_[55765]_  = \new_[55764]_  & \new_[55757]_ ;
  assign \new_[55769]_  = ~A233 & A232;
  assign \new_[55770]_  = A203 & \new_[55769]_ ;
  assign \new_[55773]_  = A236 & A234;
  assign \new_[55776]_  = A266 & ~A265;
  assign \new_[55777]_  = \new_[55776]_  & \new_[55773]_ ;
  assign \new_[55778]_  = \new_[55777]_  & \new_[55770]_ ;
  assign \new_[55782]_  = A167 & ~A168;
  assign \new_[55783]_  = ~A169 & \new_[55782]_ ;
  assign \new_[55786]_  = A199 & A166;
  assign \new_[55789]_  = A201 & ~A200;
  assign \new_[55790]_  = \new_[55789]_  & \new_[55786]_ ;
  assign \new_[55791]_  = \new_[55790]_  & \new_[55783]_ ;
  assign \new_[55795]_  = ~A233 & ~A232;
  assign \new_[55796]_  = A203 & \new_[55795]_ ;
  assign \new_[55799]_  = A266 & A265;
  assign \new_[55802]_  = A299 & ~A298;
  assign \new_[55803]_  = \new_[55802]_  & \new_[55799]_ ;
  assign \new_[55804]_  = \new_[55803]_  & \new_[55796]_ ;
  assign \new_[55808]_  = A167 & ~A168;
  assign \new_[55809]_  = ~A169 & \new_[55808]_ ;
  assign \new_[55812]_  = A199 & A166;
  assign \new_[55815]_  = A201 & ~A200;
  assign \new_[55816]_  = \new_[55815]_  & \new_[55812]_ ;
  assign \new_[55817]_  = \new_[55816]_  & \new_[55809]_ ;
  assign \new_[55821]_  = ~A233 & ~A232;
  assign \new_[55822]_  = A203 & \new_[55821]_ ;
  assign \new_[55825]_  = ~A267 & ~A266;
  assign \new_[55828]_  = A299 & ~A298;
  assign \new_[55829]_  = \new_[55828]_  & \new_[55825]_ ;
  assign \new_[55830]_  = \new_[55829]_  & \new_[55822]_ ;
  assign \new_[55834]_  = A167 & ~A168;
  assign \new_[55835]_  = ~A169 & \new_[55834]_ ;
  assign \new_[55838]_  = A199 & A166;
  assign \new_[55841]_  = A201 & ~A200;
  assign \new_[55842]_  = \new_[55841]_  & \new_[55838]_ ;
  assign \new_[55843]_  = \new_[55842]_  & \new_[55835]_ ;
  assign \new_[55847]_  = ~A233 & ~A232;
  assign \new_[55848]_  = A203 & \new_[55847]_ ;
  assign \new_[55851]_  = ~A266 & ~A265;
  assign \new_[55854]_  = A299 & ~A298;
  assign \new_[55855]_  = \new_[55854]_  & \new_[55851]_ ;
  assign \new_[55856]_  = \new_[55855]_  & \new_[55848]_ ;
  assign \new_[55860]_  = A167 & ~A169;
  assign \new_[55861]_  = A170 & \new_[55860]_ ;
  assign \new_[55864]_  = A199 & ~A166;
  assign \new_[55867]_  = A232 & A200;
  assign \new_[55868]_  = \new_[55867]_  & \new_[55864]_ ;
  assign \new_[55869]_  = \new_[55868]_  & \new_[55861]_ ;
  assign \new_[55873]_  = ~A267 & A265;
  assign \new_[55874]_  = A233 & \new_[55873]_ ;
  assign \new_[55877]_  = ~A299 & A298;
  assign \new_[55880]_  = A301 & A300;
  assign \new_[55881]_  = \new_[55880]_  & \new_[55877]_ ;
  assign \new_[55882]_  = \new_[55881]_  & \new_[55874]_ ;
  assign \new_[55886]_  = A167 & ~A169;
  assign \new_[55887]_  = A170 & \new_[55886]_ ;
  assign \new_[55890]_  = A199 & ~A166;
  assign \new_[55893]_  = A232 & A200;
  assign \new_[55894]_  = \new_[55893]_  & \new_[55890]_ ;
  assign \new_[55895]_  = \new_[55894]_  & \new_[55887]_ ;
  assign \new_[55899]_  = ~A267 & A265;
  assign \new_[55900]_  = A233 & \new_[55899]_ ;
  assign \new_[55903]_  = ~A299 & A298;
  assign \new_[55906]_  = A302 & A300;
  assign \new_[55907]_  = \new_[55906]_  & \new_[55903]_ ;
  assign \new_[55908]_  = \new_[55907]_  & \new_[55900]_ ;
  assign \new_[55912]_  = A167 & ~A169;
  assign \new_[55913]_  = A170 & \new_[55912]_ ;
  assign \new_[55916]_  = A199 & ~A166;
  assign \new_[55919]_  = A232 & A200;
  assign \new_[55920]_  = \new_[55919]_  & \new_[55916]_ ;
  assign \new_[55921]_  = \new_[55920]_  & \new_[55913]_ ;
  assign \new_[55925]_  = A266 & A265;
  assign \new_[55926]_  = A233 & \new_[55925]_ ;
  assign \new_[55929]_  = ~A299 & A298;
  assign \new_[55932]_  = A301 & A300;
  assign \new_[55933]_  = \new_[55932]_  & \new_[55929]_ ;
  assign \new_[55934]_  = \new_[55933]_  & \new_[55926]_ ;
  assign \new_[55938]_  = A167 & ~A169;
  assign \new_[55939]_  = A170 & \new_[55938]_ ;
  assign \new_[55942]_  = A199 & ~A166;
  assign \new_[55945]_  = A232 & A200;
  assign \new_[55946]_  = \new_[55945]_  & \new_[55942]_ ;
  assign \new_[55947]_  = \new_[55946]_  & \new_[55939]_ ;
  assign \new_[55951]_  = A266 & A265;
  assign \new_[55952]_  = A233 & \new_[55951]_ ;
  assign \new_[55955]_  = ~A299 & A298;
  assign \new_[55958]_  = A302 & A300;
  assign \new_[55959]_  = \new_[55958]_  & \new_[55955]_ ;
  assign \new_[55960]_  = \new_[55959]_  & \new_[55952]_ ;
  assign \new_[55964]_  = A167 & ~A169;
  assign \new_[55965]_  = A170 & \new_[55964]_ ;
  assign \new_[55968]_  = A199 & ~A166;
  assign \new_[55971]_  = A232 & A200;
  assign \new_[55972]_  = \new_[55971]_  & \new_[55968]_ ;
  assign \new_[55973]_  = \new_[55972]_  & \new_[55965]_ ;
  assign \new_[55977]_  = ~A266 & ~A265;
  assign \new_[55978]_  = A233 & \new_[55977]_ ;
  assign \new_[55981]_  = ~A299 & A298;
  assign \new_[55984]_  = A301 & A300;
  assign \new_[55985]_  = \new_[55984]_  & \new_[55981]_ ;
  assign \new_[55986]_  = \new_[55985]_  & \new_[55978]_ ;
  assign \new_[55990]_  = A167 & ~A169;
  assign \new_[55991]_  = A170 & \new_[55990]_ ;
  assign \new_[55994]_  = A199 & ~A166;
  assign \new_[55997]_  = A232 & A200;
  assign \new_[55998]_  = \new_[55997]_  & \new_[55994]_ ;
  assign \new_[55999]_  = \new_[55998]_  & \new_[55991]_ ;
  assign \new_[56003]_  = ~A266 & ~A265;
  assign \new_[56004]_  = A233 & \new_[56003]_ ;
  assign \new_[56007]_  = ~A299 & A298;
  assign \new_[56010]_  = A302 & A300;
  assign \new_[56011]_  = \new_[56010]_  & \new_[56007]_ ;
  assign \new_[56012]_  = \new_[56011]_  & \new_[56004]_ ;
  assign \new_[56016]_  = A167 & ~A169;
  assign \new_[56017]_  = A170 & \new_[56016]_ ;
  assign \new_[56020]_  = A199 & ~A166;
  assign \new_[56023]_  = ~A233 & A200;
  assign \new_[56024]_  = \new_[56023]_  & \new_[56020]_ ;
  assign \new_[56025]_  = \new_[56024]_  & \new_[56017]_ ;
  assign \new_[56029]_  = ~A266 & ~A236;
  assign \new_[56030]_  = ~A235 & \new_[56029]_ ;
  assign \new_[56033]_  = ~A269 & ~A268;
  assign \new_[56036]_  = A299 & ~A298;
  assign \new_[56037]_  = \new_[56036]_  & \new_[56033]_ ;
  assign \new_[56038]_  = \new_[56037]_  & \new_[56030]_ ;
  assign \new_[56042]_  = A167 & ~A169;
  assign \new_[56043]_  = A170 & \new_[56042]_ ;
  assign \new_[56046]_  = A199 & ~A166;
  assign \new_[56049]_  = ~A233 & A200;
  assign \new_[56050]_  = \new_[56049]_  & \new_[56046]_ ;
  assign \new_[56051]_  = \new_[56050]_  & \new_[56043]_ ;
  assign \new_[56055]_  = A266 & A265;
  assign \new_[56056]_  = ~A234 & \new_[56055]_ ;
  assign \new_[56059]_  = ~A299 & A298;
  assign \new_[56062]_  = A301 & A300;
  assign \new_[56063]_  = \new_[56062]_  & \new_[56059]_ ;
  assign \new_[56064]_  = \new_[56063]_  & \new_[56056]_ ;
  assign \new_[56068]_  = A167 & ~A169;
  assign \new_[56069]_  = A170 & \new_[56068]_ ;
  assign \new_[56072]_  = A199 & ~A166;
  assign \new_[56075]_  = ~A233 & A200;
  assign \new_[56076]_  = \new_[56075]_  & \new_[56072]_ ;
  assign \new_[56077]_  = \new_[56076]_  & \new_[56069]_ ;
  assign \new_[56081]_  = A266 & A265;
  assign \new_[56082]_  = ~A234 & \new_[56081]_ ;
  assign \new_[56085]_  = ~A299 & A298;
  assign \new_[56088]_  = A302 & A300;
  assign \new_[56089]_  = \new_[56088]_  & \new_[56085]_ ;
  assign \new_[56090]_  = \new_[56089]_  & \new_[56082]_ ;
  assign \new_[56094]_  = A167 & ~A169;
  assign \new_[56095]_  = A170 & \new_[56094]_ ;
  assign \new_[56098]_  = A199 & ~A166;
  assign \new_[56101]_  = ~A233 & A200;
  assign \new_[56102]_  = \new_[56101]_  & \new_[56098]_ ;
  assign \new_[56103]_  = \new_[56102]_  & \new_[56095]_ ;
  assign \new_[56107]_  = ~A267 & ~A266;
  assign \new_[56108]_  = ~A234 & \new_[56107]_ ;
  assign \new_[56111]_  = ~A299 & A298;
  assign \new_[56114]_  = A301 & A300;
  assign \new_[56115]_  = \new_[56114]_  & \new_[56111]_ ;
  assign \new_[56116]_  = \new_[56115]_  & \new_[56108]_ ;
  assign \new_[56120]_  = A167 & ~A169;
  assign \new_[56121]_  = A170 & \new_[56120]_ ;
  assign \new_[56124]_  = A199 & ~A166;
  assign \new_[56127]_  = ~A233 & A200;
  assign \new_[56128]_  = \new_[56127]_  & \new_[56124]_ ;
  assign \new_[56129]_  = \new_[56128]_  & \new_[56121]_ ;
  assign \new_[56133]_  = ~A267 & ~A266;
  assign \new_[56134]_  = ~A234 & \new_[56133]_ ;
  assign \new_[56137]_  = ~A299 & A298;
  assign \new_[56140]_  = A302 & A300;
  assign \new_[56141]_  = \new_[56140]_  & \new_[56137]_ ;
  assign \new_[56142]_  = \new_[56141]_  & \new_[56134]_ ;
  assign \new_[56146]_  = A167 & ~A169;
  assign \new_[56147]_  = A170 & \new_[56146]_ ;
  assign \new_[56150]_  = A199 & ~A166;
  assign \new_[56153]_  = ~A233 & A200;
  assign \new_[56154]_  = \new_[56153]_  & \new_[56150]_ ;
  assign \new_[56155]_  = \new_[56154]_  & \new_[56147]_ ;
  assign \new_[56159]_  = ~A266 & ~A265;
  assign \new_[56160]_  = ~A234 & \new_[56159]_ ;
  assign \new_[56163]_  = ~A299 & A298;
  assign \new_[56166]_  = A301 & A300;
  assign \new_[56167]_  = \new_[56166]_  & \new_[56163]_ ;
  assign \new_[56168]_  = \new_[56167]_  & \new_[56160]_ ;
  assign \new_[56172]_  = A167 & ~A169;
  assign \new_[56173]_  = A170 & \new_[56172]_ ;
  assign \new_[56176]_  = A199 & ~A166;
  assign \new_[56179]_  = ~A233 & A200;
  assign \new_[56180]_  = \new_[56179]_  & \new_[56176]_ ;
  assign \new_[56181]_  = \new_[56180]_  & \new_[56173]_ ;
  assign \new_[56185]_  = ~A266 & ~A265;
  assign \new_[56186]_  = ~A234 & \new_[56185]_ ;
  assign \new_[56189]_  = ~A299 & A298;
  assign \new_[56192]_  = A302 & A300;
  assign \new_[56193]_  = \new_[56192]_  & \new_[56189]_ ;
  assign \new_[56194]_  = \new_[56193]_  & \new_[56186]_ ;
  assign \new_[56198]_  = A167 & ~A169;
  assign \new_[56199]_  = A170 & \new_[56198]_ ;
  assign \new_[56202]_  = A199 & ~A166;
  assign \new_[56205]_  = A232 & A200;
  assign \new_[56206]_  = \new_[56205]_  & \new_[56202]_ ;
  assign \new_[56207]_  = \new_[56206]_  & \new_[56199]_ ;
  assign \new_[56211]_  = A235 & A234;
  assign \new_[56212]_  = ~A233 & \new_[56211]_ ;
  assign \new_[56215]_  = ~A266 & A265;
  assign \new_[56218]_  = A268 & A267;
  assign \new_[56219]_  = \new_[56218]_  & \new_[56215]_ ;
  assign \new_[56220]_  = \new_[56219]_  & \new_[56212]_ ;
  assign \new_[56224]_  = A167 & ~A169;
  assign \new_[56225]_  = A170 & \new_[56224]_ ;
  assign \new_[56228]_  = A199 & ~A166;
  assign \new_[56231]_  = A232 & A200;
  assign \new_[56232]_  = \new_[56231]_  & \new_[56228]_ ;
  assign \new_[56233]_  = \new_[56232]_  & \new_[56225]_ ;
  assign \new_[56237]_  = A235 & A234;
  assign \new_[56238]_  = ~A233 & \new_[56237]_ ;
  assign \new_[56241]_  = ~A266 & A265;
  assign \new_[56244]_  = A269 & A267;
  assign \new_[56245]_  = \new_[56244]_  & \new_[56241]_ ;
  assign \new_[56246]_  = \new_[56245]_  & \new_[56238]_ ;
  assign \new_[56250]_  = A167 & ~A169;
  assign \new_[56251]_  = A170 & \new_[56250]_ ;
  assign \new_[56254]_  = A199 & ~A166;
  assign \new_[56257]_  = A232 & A200;
  assign \new_[56258]_  = \new_[56257]_  & \new_[56254]_ ;
  assign \new_[56259]_  = \new_[56258]_  & \new_[56251]_ ;
  assign \new_[56263]_  = A236 & A234;
  assign \new_[56264]_  = ~A233 & \new_[56263]_ ;
  assign \new_[56267]_  = ~A266 & A265;
  assign \new_[56270]_  = A268 & A267;
  assign \new_[56271]_  = \new_[56270]_  & \new_[56267]_ ;
  assign \new_[56272]_  = \new_[56271]_  & \new_[56264]_ ;
  assign \new_[56276]_  = A167 & ~A169;
  assign \new_[56277]_  = A170 & \new_[56276]_ ;
  assign \new_[56280]_  = A199 & ~A166;
  assign \new_[56283]_  = A232 & A200;
  assign \new_[56284]_  = \new_[56283]_  & \new_[56280]_ ;
  assign \new_[56285]_  = \new_[56284]_  & \new_[56277]_ ;
  assign \new_[56289]_  = A236 & A234;
  assign \new_[56290]_  = ~A233 & \new_[56289]_ ;
  assign \new_[56293]_  = ~A266 & A265;
  assign \new_[56296]_  = A269 & A267;
  assign \new_[56297]_  = \new_[56296]_  & \new_[56293]_ ;
  assign \new_[56298]_  = \new_[56297]_  & \new_[56290]_ ;
  assign \new_[56302]_  = A167 & ~A169;
  assign \new_[56303]_  = A170 & \new_[56302]_ ;
  assign \new_[56306]_  = A199 & ~A166;
  assign \new_[56309]_  = ~A232 & A200;
  assign \new_[56310]_  = \new_[56309]_  & \new_[56306]_ ;
  assign \new_[56311]_  = \new_[56310]_  & \new_[56303]_ ;
  assign \new_[56315]_  = A266 & A265;
  assign \new_[56316]_  = ~A233 & \new_[56315]_ ;
  assign \new_[56319]_  = ~A299 & A298;
  assign \new_[56322]_  = A301 & A300;
  assign \new_[56323]_  = \new_[56322]_  & \new_[56319]_ ;
  assign \new_[56324]_  = \new_[56323]_  & \new_[56316]_ ;
  assign \new_[56328]_  = A167 & ~A169;
  assign \new_[56329]_  = A170 & \new_[56328]_ ;
  assign \new_[56332]_  = A199 & ~A166;
  assign \new_[56335]_  = ~A232 & A200;
  assign \new_[56336]_  = \new_[56335]_  & \new_[56332]_ ;
  assign \new_[56337]_  = \new_[56336]_  & \new_[56329]_ ;
  assign \new_[56341]_  = A266 & A265;
  assign \new_[56342]_  = ~A233 & \new_[56341]_ ;
  assign \new_[56345]_  = ~A299 & A298;
  assign \new_[56348]_  = A302 & A300;
  assign \new_[56349]_  = \new_[56348]_  & \new_[56345]_ ;
  assign \new_[56350]_  = \new_[56349]_  & \new_[56342]_ ;
  assign \new_[56354]_  = A167 & ~A169;
  assign \new_[56355]_  = A170 & \new_[56354]_ ;
  assign \new_[56358]_  = A199 & ~A166;
  assign \new_[56361]_  = ~A232 & A200;
  assign \new_[56362]_  = \new_[56361]_  & \new_[56358]_ ;
  assign \new_[56363]_  = \new_[56362]_  & \new_[56355]_ ;
  assign \new_[56367]_  = ~A267 & ~A266;
  assign \new_[56368]_  = ~A233 & \new_[56367]_ ;
  assign \new_[56371]_  = ~A299 & A298;
  assign \new_[56374]_  = A301 & A300;
  assign \new_[56375]_  = \new_[56374]_  & \new_[56371]_ ;
  assign \new_[56376]_  = \new_[56375]_  & \new_[56368]_ ;
  assign \new_[56380]_  = A167 & ~A169;
  assign \new_[56381]_  = A170 & \new_[56380]_ ;
  assign \new_[56384]_  = A199 & ~A166;
  assign \new_[56387]_  = ~A232 & A200;
  assign \new_[56388]_  = \new_[56387]_  & \new_[56384]_ ;
  assign \new_[56389]_  = \new_[56388]_  & \new_[56381]_ ;
  assign \new_[56393]_  = ~A267 & ~A266;
  assign \new_[56394]_  = ~A233 & \new_[56393]_ ;
  assign \new_[56397]_  = ~A299 & A298;
  assign \new_[56400]_  = A302 & A300;
  assign \new_[56401]_  = \new_[56400]_  & \new_[56397]_ ;
  assign \new_[56402]_  = \new_[56401]_  & \new_[56394]_ ;
  assign \new_[56406]_  = A167 & ~A169;
  assign \new_[56407]_  = A170 & \new_[56406]_ ;
  assign \new_[56410]_  = A199 & ~A166;
  assign \new_[56413]_  = ~A232 & A200;
  assign \new_[56414]_  = \new_[56413]_  & \new_[56410]_ ;
  assign \new_[56415]_  = \new_[56414]_  & \new_[56407]_ ;
  assign \new_[56419]_  = ~A266 & ~A265;
  assign \new_[56420]_  = ~A233 & \new_[56419]_ ;
  assign \new_[56423]_  = ~A299 & A298;
  assign \new_[56426]_  = A301 & A300;
  assign \new_[56427]_  = \new_[56426]_  & \new_[56423]_ ;
  assign \new_[56428]_  = \new_[56427]_  & \new_[56420]_ ;
  assign \new_[56432]_  = A167 & ~A169;
  assign \new_[56433]_  = A170 & \new_[56432]_ ;
  assign \new_[56436]_  = A199 & ~A166;
  assign \new_[56439]_  = ~A232 & A200;
  assign \new_[56440]_  = \new_[56439]_  & \new_[56436]_ ;
  assign \new_[56441]_  = \new_[56440]_  & \new_[56433]_ ;
  assign \new_[56445]_  = ~A266 & ~A265;
  assign \new_[56446]_  = ~A233 & \new_[56445]_ ;
  assign \new_[56449]_  = ~A299 & A298;
  assign \new_[56452]_  = A302 & A300;
  assign \new_[56453]_  = \new_[56452]_  & \new_[56449]_ ;
  assign \new_[56454]_  = \new_[56453]_  & \new_[56446]_ ;
  assign \new_[56458]_  = A167 & ~A169;
  assign \new_[56459]_  = A170 & \new_[56458]_ ;
  assign \new_[56462]_  = ~A200 & ~A166;
  assign \new_[56465]_  = ~A203 & ~A202;
  assign \new_[56466]_  = \new_[56465]_  & \new_[56462]_ ;
  assign \new_[56467]_  = \new_[56466]_  & \new_[56459]_ ;
  assign \new_[56471]_  = A265 & A233;
  assign \new_[56472]_  = A232 & \new_[56471]_ ;
  assign \new_[56475]_  = ~A269 & ~A268;
  assign \new_[56478]_  = A299 & ~A298;
  assign \new_[56479]_  = \new_[56478]_  & \new_[56475]_ ;
  assign \new_[56480]_  = \new_[56479]_  & \new_[56472]_ ;
  assign \new_[56484]_  = A167 & ~A169;
  assign \new_[56485]_  = A170 & \new_[56484]_ ;
  assign \new_[56488]_  = ~A200 & ~A166;
  assign \new_[56491]_  = ~A203 & ~A202;
  assign \new_[56492]_  = \new_[56491]_  & \new_[56488]_ ;
  assign \new_[56493]_  = \new_[56492]_  & \new_[56485]_ ;
  assign \new_[56497]_  = ~A236 & ~A235;
  assign \new_[56498]_  = ~A233 & \new_[56497]_ ;
  assign \new_[56501]_  = A266 & A265;
  assign \new_[56504]_  = A299 & ~A298;
  assign \new_[56505]_  = \new_[56504]_  & \new_[56501]_ ;
  assign \new_[56506]_  = \new_[56505]_  & \new_[56498]_ ;
  assign \new_[56510]_  = A167 & ~A169;
  assign \new_[56511]_  = A170 & \new_[56510]_ ;
  assign \new_[56514]_  = ~A200 & ~A166;
  assign \new_[56517]_  = ~A203 & ~A202;
  assign \new_[56518]_  = \new_[56517]_  & \new_[56514]_ ;
  assign \new_[56519]_  = \new_[56518]_  & \new_[56511]_ ;
  assign \new_[56523]_  = ~A236 & ~A235;
  assign \new_[56524]_  = ~A233 & \new_[56523]_ ;
  assign \new_[56527]_  = ~A267 & ~A266;
  assign \new_[56530]_  = A299 & ~A298;
  assign \new_[56531]_  = \new_[56530]_  & \new_[56527]_ ;
  assign \new_[56532]_  = \new_[56531]_  & \new_[56524]_ ;
  assign \new_[56536]_  = A167 & ~A169;
  assign \new_[56537]_  = A170 & \new_[56536]_ ;
  assign \new_[56540]_  = ~A200 & ~A166;
  assign \new_[56543]_  = ~A203 & ~A202;
  assign \new_[56544]_  = \new_[56543]_  & \new_[56540]_ ;
  assign \new_[56545]_  = \new_[56544]_  & \new_[56537]_ ;
  assign \new_[56549]_  = ~A236 & ~A235;
  assign \new_[56550]_  = ~A233 & \new_[56549]_ ;
  assign \new_[56553]_  = ~A266 & ~A265;
  assign \new_[56556]_  = A299 & ~A298;
  assign \new_[56557]_  = \new_[56556]_  & \new_[56553]_ ;
  assign \new_[56558]_  = \new_[56557]_  & \new_[56550]_ ;
  assign \new_[56562]_  = A167 & ~A169;
  assign \new_[56563]_  = A170 & \new_[56562]_ ;
  assign \new_[56566]_  = ~A200 & ~A166;
  assign \new_[56569]_  = ~A203 & ~A202;
  assign \new_[56570]_  = \new_[56569]_  & \new_[56566]_ ;
  assign \new_[56571]_  = \new_[56570]_  & \new_[56563]_ ;
  assign \new_[56575]_  = ~A266 & ~A234;
  assign \new_[56576]_  = ~A233 & \new_[56575]_ ;
  assign \new_[56579]_  = ~A269 & ~A268;
  assign \new_[56582]_  = A299 & ~A298;
  assign \new_[56583]_  = \new_[56582]_  & \new_[56579]_ ;
  assign \new_[56584]_  = \new_[56583]_  & \new_[56576]_ ;
  assign \new_[56588]_  = A167 & ~A169;
  assign \new_[56589]_  = A170 & \new_[56588]_ ;
  assign \new_[56592]_  = ~A200 & ~A166;
  assign \new_[56595]_  = ~A203 & ~A202;
  assign \new_[56596]_  = \new_[56595]_  & \new_[56592]_ ;
  assign \new_[56597]_  = \new_[56596]_  & \new_[56589]_ ;
  assign \new_[56601]_  = A234 & ~A233;
  assign \new_[56602]_  = A232 & \new_[56601]_ ;
  assign \new_[56605]_  = A298 & A235;
  assign \new_[56608]_  = ~A302 & ~A301;
  assign \new_[56609]_  = \new_[56608]_  & \new_[56605]_ ;
  assign \new_[56610]_  = \new_[56609]_  & \new_[56602]_ ;
  assign \new_[56614]_  = A167 & ~A169;
  assign \new_[56615]_  = A170 & \new_[56614]_ ;
  assign \new_[56618]_  = ~A200 & ~A166;
  assign \new_[56621]_  = ~A203 & ~A202;
  assign \new_[56622]_  = \new_[56621]_  & \new_[56618]_ ;
  assign \new_[56623]_  = \new_[56622]_  & \new_[56615]_ ;
  assign \new_[56627]_  = A234 & ~A233;
  assign \new_[56628]_  = A232 & \new_[56627]_ ;
  assign \new_[56631]_  = A298 & A236;
  assign \new_[56634]_  = ~A302 & ~A301;
  assign \new_[56635]_  = \new_[56634]_  & \new_[56631]_ ;
  assign \new_[56636]_  = \new_[56635]_  & \new_[56628]_ ;
  assign \new_[56640]_  = A167 & ~A169;
  assign \new_[56641]_  = A170 & \new_[56640]_ ;
  assign \new_[56644]_  = ~A200 & ~A166;
  assign \new_[56647]_  = ~A203 & ~A202;
  assign \new_[56648]_  = \new_[56647]_  & \new_[56644]_ ;
  assign \new_[56649]_  = \new_[56648]_  & \new_[56641]_ ;
  assign \new_[56653]_  = ~A266 & ~A233;
  assign \new_[56654]_  = ~A232 & \new_[56653]_ ;
  assign \new_[56657]_  = ~A269 & ~A268;
  assign \new_[56660]_  = A299 & ~A298;
  assign \new_[56661]_  = \new_[56660]_  & \new_[56657]_ ;
  assign \new_[56662]_  = \new_[56661]_  & \new_[56654]_ ;
  assign \new_[56666]_  = A167 & ~A169;
  assign \new_[56667]_  = A170 & \new_[56666]_ ;
  assign \new_[56670]_  = ~A200 & ~A166;
  assign \new_[56673]_  = A232 & ~A201;
  assign \new_[56674]_  = \new_[56673]_  & \new_[56670]_ ;
  assign \new_[56675]_  = \new_[56674]_  & \new_[56667]_ ;
  assign \new_[56679]_  = ~A267 & A265;
  assign \new_[56680]_  = A233 & \new_[56679]_ ;
  assign \new_[56683]_  = ~A299 & A298;
  assign \new_[56686]_  = A301 & A300;
  assign \new_[56687]_  = \new_[56686]_  & \new_[56683]_ ;
  assign \new_[56688]_  = \new_[56687]_  & \new_[56680]_ ;
  assign \new_[56692]_  = A167 & ~A169;
  assign \new_[56693]_  = A170 & \new_[56692]_ ;
  assign \new_[56696]_  = ~A200 & ~A166;
  assign \new_[56699]_  = A232 & ~A201;
  assign \new_[56700]_  = \new_[56699]_  & \new_[56696]_ ;
  assign \new_[56701]_  = \new_[56700]_  & \new_[56693]_ ;
  assign \new_[56705]_  = ~A267 & A265;
  assign \new_[56706]_  = A233 & \new_[56705]_ ;
  assign \new_[56709]_  = ~A299 & A298;
  assign \new_[56712]_  = A302 & A300;
  assign \new_[56713]_  = \new_[56712]_  & \new_[56709]_ ;
  assign \new_[56714]_  = \new_[56713]_  & \new_[56706]_ ;
  assign \new_[56718]_  = A167 & ~A169;
  assign \new_[56719]_  = A170 & \new_[56718]_ ;
  assign \new_[56722]_  = ~A200 & ~A166;
  assign \new_[56725]_  = A232 & ~A201;
  assign \new_[56726]_  = \new_[56725]_  & \new_[56722]_ ;
  assign \new_[56727]_  = \new_[56726]_  & \new_[56719]_ ;
  assign \new_[56731]_  = A266 & A265;
  assign \new_[56732]_  = A233 & \new_[56731]_ ;
  assign \new_[56735]_  = ~A299 & A298;
  assign \new_[56738]_  = A301 & A300;
  assign \new_[56739]_  = \new_[56738]_  & \new_[56735]_ ;
  assign \new_[56740]_  = \new_[56739]_  & \new_[56732]_ ;
  assign \new_[56744]_  = A167 & ~A169;
  assign \new_[56745]_  = A170 & \new_[56744]_ ;
  assign \new_[56748]_  = ~A200 & ~A166;
  assign \new_[56751]_  = A232 & ~A201;
  assign \new_[56752]_  = \new_[56751]_  & \new_[56748]_ ;
  assign \new_[56753]_  = \new_[56752]_  & \new_[56745]_ ;
  assign \new_[56757]_  = A266 & A265;
  assign \new_[56758]_  = A233 & \new_[56757]_ ;
  assign \new_[56761]_  = ~A299 & A298;
  assign \new_[56764]_  = A302 & A300;
  assign \new_[56765]_  = \new_[56764]_  & \new_[56761]_ ;
  assign \new_[56766]_  = \new_[56765]_  & \new_[56758]_ ;
  assign \new_[56770]_  = A167 & ~A169;
  assign \new_[56771]_  = A170 & \new_[56770]_ ;
  assign \new_[56774]_  = ~A200 & ~A166;
  assign \new_[56777]_  = A232 & ~A201;
  assign \new_[56778]_  = \new_[56777]_  & \new_[56774]_ ;
  assign \new_[56779]_  = \new_[56778]_  & \new_[56771]_ ;
  assign \new_[56783]_  = ~A266 & ~A265;
  assign \new_[56784]_  = A233 & \new_[56783]_ ;
  assign \new_[56787]_  = ~A299 & A298;
  assign \new_[56790]_  = A301 & A300;
  assign \new_[56791]_  = \new_[56790]_  & \new_[56787]_ ;
  assign \new_[56792]_  = \new_[56791]_  & \new_[56784]_ ;
  assign \new_[56796]_  = A167 & ~A169;
  assign \new_[56797]_  = A170 & \new_[56796]_ ;
  assign \new_[56800]_  = ~A200 & ~A166;
  assign \new_[56803]_  = A232 & ~A201;
  assign \new_[56804]_  = \new_[56803]_  & \new_[56800]_ ;
  assign \new_[56805]_  = \new_[56804]_  & \new_[56797]_ ;
  assign \new_[56809]_  = ~A266 & ~A265;
  assign \new_[56810]_  = A233 & \new_[56809]_ ;
  assign \new_[56813]_  = ~A299 & A298;
  assign \new_[56816]_  = A302 & A300;
  assign \new_[56817]_  = \new_[56816]_  & \new_[56813]_ ;
  assign \new_[56818]_  = \new_[56817]_  & \new_[56810]_ ;
  assign \new_[56822]_  = A167 & ~A169;
  assign \new_[56823]_  = A170 & \new_[56822]_ ;
  assign \new_[56826]_  = ~A200 & ~A166;
  assign \new_[56829]_  = ~A233 & ~A201;
  assign \new_[56830]_  = \new_[56829]_  & \new_[56826]_ ;
  assign \new_[56831]_  = \new_[56830]_  & \new_[56823]_ ;
  assign \new_[56835]_  = ~A266 & ~A236;
  assign \new_[56836]_  = ~A235 & \new_[56835]_ ;
  assign \new_[56839]_  = ~A269 & ~A268;
  assign \new_[56842]_  = A299 & ~A298;
  assign \new_[56843]_  = \new_[56842]_  & \new_[56839]_ ;
  assign \new_[56844]_  = \new_[56843]_  & \new_[56836]_ ;
  assign \new_[56848]_  = A167 & ~A169;
  assign \new_[56849]_  = A170 & \new_[56848]_ ;
  assign \new_[56852]_  = ~A200 & ~A166;
  assign \new_[56855]_  = ~A233 & ~A201;
  assign \new_[56856]_  = \new_[56855]_  & \new_[56852]_ ;
  assign \new_[56857]_  = \new_[56856]_  & \new_[56849]_ ;
  assign \new_[56861]_  = A266 & A265;
  assign \new_[56862]_  = ~A234 & \new_[56861]_ ;
  assign \new_[56865]_  = ~A299 & A298;
  assign \new_[56868]_  = A301 & A300;
  assign \new_[56869]_  = \new_[56868]_  & \new_[56865]_ ;
  assign \new_[56870]_  = \new_[56869]_  & \new_[56862]_ ;
  assign \new_[56874]_  = A167 & ~A169;
  assign \new_[56875]_  = A170 & \new_[56874]_ ;
  assign \new_[56878]_  = ~A200 & ~A166;
  assign \new_[56881]_  = ~A233 & ~A201;
  assign \new_[56882]_  = \new_[56881]_  & \new_[56878]_ ;
  assign \new_[56883]_  = \new_[56882]_  & \new_[56875]_ ;
  assign \new_[56887]_  = A266 & A265;
  assign \new_[56888]_  = ~A234 & \new_[56887]_ ;
  assign \new_[56891]_  = ~A299 & A298;
  assign \new_[56894]_  = A302 & A300;
  assign \new_[56895]_  = \new_[56894]_  & \new_[56891]_ ;
  assign \new_[56896]_  = \new_[56895]_  & \new_[56888]_ ;
  assign \new_[56900]_  = A167 & ~A169;
  assign \new_[56901]_  = A170 & \new_[56900]_ ;
  assign \new_[56904]_  = ~A200 & ~A166;
  assign \new_[56907]_  = ~A233 & ~A201;
  assign \new_[56908]_  = \new_[56907]_  & \new_[56904]_ ;
  assign \new_[56909]_  = \new_[56908]_  & \new_[56901]_ ;
  assign \new_[56913]_  = ~A267 & ~A266;
  assign \new_[56914]_  = ~A234 & \new_[56913]_ ;
  assign \new_[56917]_  = ~A299 & A298;
  assign \new_[56920]_  = A301 & A300;
  assign \new_[56921]_  = \new_[56920]_  & \new_[56917]_ ;
  assign \new_[56922]_  = \new_[56921]_  & \new_[56914]_ ;
  assign \new_[56926]_  = A167 & ~A169;
  assign \new_[56927]_  = A170 & \new_[56926]_ ;
  assign \new_[56930]_  = ~A200 & ~A166;
  assign \new_[56933]_  = ~A233 & ~A201;
  assign \new_[56934]_  = \new_[56933]_  & \new_[56930]_ ;
  assign \new_[56935]_  = \new_[56934]_  & \new_[56927]_ ;
  assign \new_[56939]_  = ~A267 & ~A266;
  assign \new_[56940]_  = ~A234 & \new_[56939]_ ;
  assign \new_[56943]_  = ~A299 & A298;
  assign \new_[56946]_  = A302 & A300;
  assign \new_[56947]_  = \new_[56946]_  & \new_[56943]_ ;
  assign \new_[56948]_  = \new_[56947]_  & \new_[56940]_ ;
  assign \new_[56952]_  = A167 & ~A169;
  assign \new_[56953]_  = A170 & \new_[56952]_ ;
  assign \new_[56956]_  = ~A200 & ~A166;
  assign \new_[56959]_  = ~A233 & ~A201;
  assign \new_[56960]_  = \new_[56959]_  & \new_[56956]_ ;
  assign \new_[56961]_  = \new_[56960]_  & \new_[56953]_ ;
  assign \new_[56965]_  = ~A266 & ~A265;
  assign \new_[56966]_  = ~A234 & \new_[56965]_ ;
  assign \new_[56969]_  = ~A299 & A298;
  assign \new_[56972]_  = A301 & A300;
  assign \new_[56973]_  = \new_[56972]_  & \new_[56969]_ ;
  assign \new_[56974]_  = \new_[56973]_  & \new_[56966]_ ;
  assign \new_[56978]_  = A167 & ~A169;
  assign \new_[56979]_  = A170 & \new_[56978]_ ;
  assign \new_[56982]_  = ~A200 & ~A166;
  assign \new_[56985]_  = ~A233 & ~A201;
  assign \new_[56986]_  = \new_[56985]_  & \new_[56982]_ ;
  assign \new_[56987]_  = \new_[56986]_  & \new_[56979]_ ;
  assign \new_[56991]_  = ~A266 & ~A265;
  assign \new_[56992]_  = ~A234 & \new_[56991]_ ;
  assign \new_[56995]_  = ~A299 & A298;
  assign \new_[56998]_  = A302 & A300;
  assign \new_[56999]_  = \new_[56998]_  & \new_[56995]_ ;
  assign \new_[57000]_  = \new_[56999]_  & \new_[56992]_ ;
  assign \new_[57004]_  = A167 & ~A169;
  assign \new_[57005]_  = A170 & \new_[57004]_ ;
  assign \new_[57008]_  = ~A200 & ~A166;
  assign \new_[57011]_  = A232 & ~A201;
  assign \new_[57012]_  = \new_[57011]_  & \new_[57008]_ ;
  assign \new_[57013]_  = \new_[57012]_  & \new_[57005]_ ;
  assign \new_[57017]_  = A235 & A234;
  assign \new_[57018]_  = ~A233 & \new_[57017]_ ;
  assign \new_[57021]_  = ~A266 & A265;
  assign \new_[57024]_  = A268 & A267;
  assign \new_[57025]_  = \new_[57024]_  & \new_[57021]_ ;
  assign \new_[57026]_  = \new_[57025]_  & \new_[57018]_ ;
  assign \new_[57030]_  = A167 & ~A169;
  assign \new_[57031]_  = A170 & \new_[57030]_ ;
  assign \new_[57034]_  = ~A200 & ~A166;
  assign \new_[57037]_  = A232 & ~A201;
  assign \new_[57038]_  = \new_[57037]_  & \new_[57034]_ ;
  assign \new_[57039]_  = \new_[57038]_  & \new_[57031]_ ;
  assign \new_[57043]_  = A235 & A234;
  assign \new_[57044]_  = ~A233 & \new_[57043]_ ;
  assign \new_[57047]_  = ~A266 & A265;
  assign \new_[57050]_  = A269 & A267;
  assign \new_[57051]_  = \new_[57050]_  & \new_[57047]_ ;
  assign \new_[57052]_  = \new_[57051]_  & \new_[57044]_ ;
  assign \new_[57056]_  = A167 & ~A169;
  assign \new_[57057]_  = A170 & \new_[57056]_ ;
  assign \new_[57060]_  = ~A200 & ~A166;
  assign \new_[57063]_  = A232 & ~A201;
  assign \new_[57064]_  = \new_[57063]_  & \new_[57060]_ ;
  assign \new_[57065]_  = \new_[57064]_  & \new_[57057]_ ;
  assign \new_[57069]_  = A236 & A234;
  assign \new_[57070]_  = ~A233 & \new_[57069]_ ;
  assign \new_[57073]_  = ~A266 & A265;
  assign \new_[57076]_  = A268 & A267;
  assign \new_[57077]_  = \new_[57076]_  & \new_[57073]_ ;
  assign \new_[57078]_  = \new_[57077]_  & \new_[57070]_ ;
  assign \new_[57082]_  = A167 & ~A169;
  assign \new_[57083]_  = A170 & \new_[57082]_ ;
  assign \new_[57086]_  = ~A200 & ~A166;
  assign \new_[57089]_  = A232 & ~A201;
  assign \new_[57090]_  = \new_[57089]_  & \new_[57086]_ ;
  assign \new_[57091]_  = \new_[57090]_  & \new_[57083]_ ;
  assign \new_[57095]_  = A236 & A234;
  assign \new_[57096]_  = ~A233 & \new_[57095]_ ;
  assign \new_[57099]_  = ~A266 & A265;
  assign \new_[57102]_  = A269 & A267;
  assign \new_[57103]_  = \new_[57102]_  & \new_[57099]_ ;
  assign \new_[57104]_  = \new_[57103]_  & \new_[57096]_ ;
  assign \new_[57108]_  = A167 & ~A169;
  assign \new_[57109]_  = A170 & \new_[57108]_ ;
  assign \new_[57112]_  = ~A200 & ~A166;
  assign \new_[57115]_  = ~A232 & ~A201;
  assign \new_[57116]_  = \new_[57115]_  & \new_[57112]_ ;
  assign \new_[57117]_  = \new_[57116]_  & \new_[57109]_ ;
  assign \new_[57121]_  = A266 & A265;
  assign \new_[57122]_  = ~A233 & \new_[57121]_ ;
  assign \new_[57125]_  = ~A299 & A298;
  assign \new_[57128]_  = A301 & A300;
  assign \new_[57129]_  = \new_[57128]_  & \new_[57125]_ ;
  assign \new_[57130]_  = \new_[57129]_  & \new_[57122]_ ;
  assign \new_[57134]_  = A167 & ~A169;
  assign \new_[57135]_  = A170 & \new_[57134]_ ;
  assign \new_[57138]_  = ~A200 & ~A166;
  assign \new_[57141]_  = ~A232 & ~A201;
  assign \new_[57142]_  = \new_[57141]_  & \new_[57138]_ ;
  assign \new_[57143]_  = \new_[57142]_  & \new_[57135]_ ;
  assign \new_[57147]_  = A266 & A265;
  assign \new_[57148]_  = ~A233 & \new_[57147]_ ;
  assign \new_[57151]_  = ~A299 & A298;
  assign \new_[57154]_  = A302 & A300;
  assign \new_[57155]_  = \new_[57154]_  & \new_[57151]_ ;
  assign \new_[57156]_  = \new_[57155]_  & \new_[57148]_ ;
  assign \new_[57160]_  = A167 & ~A169;
  assign \new_[57161]_  = A170 & \new_[57160]_ ;
  assign \new_[57164]_  = ~A200 & ~A166;
  assign \new_[57167]_  = ~A232 & ~A201;
  assign \new_[57168]_  = \new_[57167]_  & \new_[57164]_ ;
  assign \new_[57169]_  = \new_[57168]_  & \new_[57161]_ ;
  assign \new_[57173]_  = ~A267 & ~A266;
  assign \new_[57174]_  = ~A233 & \new_[57173]_ ;
  assign \new_[57177]_  = ~A299 & A298;
  assign \new_[57180]_  = A301 & A300;
  assign \new_[57181]_  = \new_[57180]_  & \new_[57177]_ ;
  assign \new_[57182]_  = \new_[57181]_  & \new_[57174]_ ;
  assign \new_[57186]_  = A167 & ~A169;
  assign \new_[57187]_  = A170 & \new_[57186]_ ;
  assign \new_[57190]_  = ~A200 & ~A166;
  assign \new_[57193]_  = ~A232 & ~A201;
  assign \new_[57194]_  = \new_[57193]_  & \new_[57190]_ ;
  assign \new_[57195]_  = \new_[57194]_  & \new_[57187]_ ;
  assign \new_[57199]_  = ~A267 & ~A266;
  assign \new_[57200]_  = ~A233 & \new_[57199]_ ;
  assign \new_[57203]_  = ~A299 & A298;
  assign \new_[57206]_  = A302 & A300;
  assign \new_[57207]_  = \new_[57206]_  & \new_[57203]_ ;
  assign \new_[57208]_  = \new_[57207]_  & \new_[57200]_ ;
  assign \new_[57212]_  = A167 & ~A169;
  assign \new_[57213]_  = A170 & \new_[57212]_ ;
  assign \new_[57216]_  = ~A200 & ~A166;
  assign \new_[57219]_  = ~A232 & ~A201;
  assign \new_[57220]_  = \new_[57219]_  & \new_[57216]_ ;
  assign \new_[57221]_  = \new_[57220]_  & \new_[57213]_ ;
  assign \new_[57225]_  = ~A266 & ~A265;
  assign \new_[57226]_  = ~A233 & \new_[57225]_ ;
  assign \new_[57229]_  = ~A299 & A298;
  assign \new_[57232]_  = A301 & A300;
  assign \new_[57233]_  = \new_[57232]_  & \new_[57229]_ ;
  assign \new_[57234]_  = \new_[57233]_  & \new_[57226]_ ;
  assign \new_[57238]_  = A167 & ~A169;
  assign \new_[57239]_  = A170 & \new_[57238]_ ;
  assign \new_[57242]_  = ~A200 & ~A166;
  assign \new_[57245]_  = ~A232 & ~A201;
  assign \new_[57246]_  = \new_[57245]_  & \new_[57242]_ ;
  assign \new_[57247]_  = \new_[57246]_  & \new_[57239]_ ;
  assign \new_[57251]_  = ~A266 & ~A265;
  assign \new_[57252]_  = ~A233 & \new_[57251]_ ;
  assign \new_[57255]_  = ~A299 & A298;
  assign \new_[57258]_  = A302 & A300;
  assign \new_[57259]_  = \new_[57258]_  & \new_[57255]_ ;
  assign \new_[57260]_  = \new_[57259]_  & \new_[57252]_ ;
  assign \new_[57264]_  = A167 & ~A169;
  assign \new_[57265]_  = A170 & \new_[57264]_ ;
  assign \new_[57268]_  = ~A199 & ~A166;
  assign \new_[57271]_  = A232 & ~A200;
  assign \new_[57272]_  = \new_[57271]_  & \new_[57268]_ ;
  assign \new_[57273]_  = \new_[57272]_  & \new_[57265]_ ;
  assign \new_[57277]_  = ~A267 & A265;
  assign \new_[57278]_  = A233 & \new_[57277]_ ;
  assign \new_[57281]_  = ~A299 & A298;
  assign \new_[57284]_  = A301 & A300;
  assign \new_[57285]_  = \new_[57284]_  & \new_[57281]_ ;
  assign \new_[57286]_  = \new_[57285]_  & \new_[57278]_ ;
  assign \new_[57290]_  = A167 & ~A169;
  assign \new_[57291]_  = A170 & \new_[57290]_ ;
  assign \new_[57294]_  = ~A199 & ~A166;
  assign \new_[57297]_  = A232 & ~A200;
  assign \new_[57298]_  = \new_[57297]_  & \new_[57294]_ ;
  assign \new_[57299]_  = \new_[57298]_  & \new_[57291]_ ;
  assign \new_[57303]_  = ~A267 & A265;
  assign \new_[57304]_  = A233 & \new_[57303]_ ;
  assign \new_[57307]_  = ~A299 & A298;
  assign \new_[57310]_  = A302 & A300;
  assign \new_[57311]_  = \new_[57310]_  & \new_[57307]_ ;
  assign \new_[57312]_  = \new_[57311]_  & \new_[57304]_ ;
  assign \new_[57316]_  = A167 & ~A169;
  assign \new_[57317]_  = A170 & \new_[57316]_ ;
  assign \new_[57320]_  = ~A199 & ~A166;
  assign \new_[57323]_  = A232 & ~A200;
  assign \new_[57324]_  = \new_[57323]_  & \new_[57320]_ ;
  assign \new_[57325]_  = \new_[57324]_  & \new_[57317]_ ;
  assign \new_[57329]_  = A266 & A265;
  assign \new_[57330]_  = A233 & \new_[57329]_ ;
  assign \new_[57333]_  = ~A299 & A298;
  assign \new_[57336]_  = A301 & A300;
  assign \new_[57337]_  = \new_[57336]_  & \new_[57333]_ ;
  assign \new_[57338]_  = \new_[57337]_  & \new_[57330]_ ;
  assign \new_[57342]_  = A167 & ~A169;
  assign \new_[57343]_  = A170 & \new_[57342]_ ;
  assign \new_[57346]_  = ~A199 & ~A166;
  assign \new_[57349]_  = A232 & ~A200;
  assign \new_[57350]_  = \new_[57349]_  & \new_[57346]_ ;
  assign \new_[57351]_  = \new_[57350]_  & \new_[57343]_ ;
  assign \new_[57355]_  = A266 & A265;
  assign \new_[57356]_  = A233 & \new_[57355]_ ;
  assign \new_[57359]_  = ~A299 & A298;
  assign \new_[57362]_  = A302 & A300;
  assign \new_[57363]_  = \new_[57362]_  & \new_[57359]_ ;
  assign \new_[57364]_  = \new_[57363]_  & \new_[57356]_ ;
  assign \new_[57368]_  = A167 & ~A169;
  assign \new_[57369]_  = A170 & \new_[57368]_ ;
  assign \new_[57372]_  = ~A199 & ~A166;
  assign \new_[57375]_  = A232 & ~A200;
  assign \new_[57376]_  = \new_[57375]_  & \new_[57372]_ ;
  assign \new_[57377]_  = \new_[57376]_  & \new_[57369]_ ;
  assign \new_[57381]_  = ~A266 & ~A265;
  assign \new_[57382]_  = A233 & \new_[57381]_ ;
  assign \new_[57385]_  = ~A299 & A298;
  assign \new_[57388]_  = A301 & A300;
  assign \new_[57389]_  = \new_[57388]_  & \new_[57385]_ ;
  assign \new_[57390]_  = \new_[57389]_  & \new_[57382]_ ;
  assign \new_[57394]_  = A167 & ~A169;
  assign \new_[57395]_  = A170 & \new_[57394]_ ;
  assign \new_[57398]_  = ~A199 & ~A166;
  assign \new_[57401]_  = A232 & ~A200;
  assign \new_[57402]_  = \new_[57401]_  & \new_[57398]_ ;
  assign \new_[57403]_  = \new_[57402]_  & \new_[57395]_ ;
  assign \new_[57407]_  = ~A266 & ~A265;
  assign \new_[57408]_  = A233 & \new_[57407]_ ;
  assign \new_[57411]_  = ~A299 & A298;
  assign \new_[57414]_  = A302 & A300;
  assign \new_[57415]_  = \new_[57414]_  & \new_[57411]_ ;
  assign \new_[57416]_  = \new_[57415]_  & \new_[57408]_ ;
  assign \new_[57420]_  = A167 & ~A169;
  assign \new_[57421]_  = A170 & \new_[57420]_ ;
  assign \new_[57424]_  = ~A199 & ~A166;
  assign \new_[57427]_  = ~A233 & ~A200;
  assign \new_[57428]_  = \new_[57427]_  & \new_[57424]_ ;
  assign \new_[57429]_  = \new_[57428]_  & \new_[57421]_ ;
  assign \new_[57433]_  = ~A266 & ~A236;
  assign \new_[57434]_  = ~A235 & \new_[57433]_ ;
  assign \new_[57437]_  = ~A269 & ~A268;
  assign \new_[57440]_  = A299 & ~A298;
  assign \new_[57441]_  = \new_[57440]_  & \new_[57437]_ ;
  assign \new_[57442]_  = \new_[57441]_  & \new_[57434]_ ;
  assign \new_[57446]_  = A167 & ~A169;
  assign \new_[57447]_  = A170 & \new_[57446]_ ;
  assign \new_[57450]_  = ~A199 & ~A166;
  assign \new_[57453]_  = ~A233 & ~A200;
  assign \new_[57454]_  = \new_[57453]_  & \new_[57450]_ ;
  assign \new_[57455]_  = \new_[57454]_  & \new_[57447]_ ;
  assign \new_[57459]_  = A266 & A265;
  assign \new_[57460]_  = ~A234 & \new_[57459]_ ;
  assign \new_[57463]_  = ~A299 & A298;
  assign \new_[57466]_  = A301 & A300;
  assign \new_[57467]_  = \new_[57466]_  & \new_[57463]_ ;
  assign \new_[57468]_  = \new_[57467]_  & \new_[57460]_ ;
  assign \new_[57472]_  = A167 & ~A169;
  assign \new_[57473]_  = A170 & \new_[57472]_ ;
  assign \new_[57476]_  = ~A199 & ~A166;
  assign \new_[57479]_  = ~A233 & ~A200;
  assign \new_[57480]_  = \new_[57479]_  & \new_[57476]_ ;
  assign \new_[57481]_  = \new_[57480]_  & \new_[57473]_ ;
  assign \new_[57485]_  = A266 & A265;
  assign \new_[57486]_  = ~A234 & \new_[57485]_ ;
  assign \new_[57489]_  = ~A299 & A298;
  assign \new_[57492]_  = A302 & A300;
  assign \new_[57493]_  = \new_[57492]_  & \new_[57489]_ ;
  assign \new_[57494]_  = \new_[57493]_  & \new_[57486]_ ;
  assign \new_[57498]_  = A167 & ~A169;
  assign \new_[57499]_  = A170 & \new_[57498]_ ;
  assign \new_[57502]_  = ~A199 & ~A166;
  assign \new_[57505]_  = ~A233 & ~A200;
  assign \new_[57506]_  = \new_[57505]_  & \new_[57502]_ ;
  assign \new_[57507]_  = \new_[57506]_  & \new_[57499]_ ;
  assign \new_[57511]_  = ~A267 & ~A266;
  assign \new_[57512]_  = ~A234 & \new_[57511]_ ;
  assign \new_[57515]_  = ~A299 & A298;
  assign \new_[57518]_  = A301 & A300;
  assign \new_[57519]_  = \new_[57518]_  & \new_[57515]_ ;
  assign \new_[57520]_  = \new_[57519]_  & \new_[57512]_ ;
  assign \new_[57524]_  = A167 & ~A169;
  assign \new_[57525]_  = A170 & \new_[57524]_ ;
  assign \new_[57528]_  = ~A199 & ~A166;
  assign \new_[57531]_  = ~A233 & ~A200;
  assign \new_[57532]_  = \new_[57531]_  & \new_[57528]_ ;
  assign \new_[57533]_  = \new_[57532]_  & \new_[57525]_ ;
  assign \new_[57537]_  = ~A267 & ~A266;
  assign \new_[57538]_  = ~A234 & \new_[57537]_ ;
  assign \new_[57541]_  = ~A299 & A298;
  assign \new_[57544]_  = A302 & A300;
  assign \new_[57545]_  = \new_[57544]_  & \new_[57541]_ ;
  assign \new_[57546]_  = \new_[57545]_  & \new_[57538]_ ;
  assign \new_[57550]_  = A167 & ~A169;
  assign \new_[57551]_  = A170 & \new_[57550]_ ;
  assign \new_[57554]_  = ~A199 & ~A166;
  assign \new_[57557]_  = ~A233 & ~A200;
  assign \new_[57558]_  = \new_[57557]_  & \new_[57554]_ ;
  assign \new_[57559]_  = \new_[57558]_  & \new_[57551]_ ;
  assign \new_[57563]_  = ~A266 & ~A265;
  assign \new_[57564]_  = ~A234 & \new_[57563]_ ;
  assign \new_[57567]_  = ~A299 & A298;
  assign \new_[57570]_  = A301 & A300;
  assign \new_[57571]_  = \new_[57570]_  & \new_[57567]_ ;
  assign \new_[57572]_  = \new_[57571]_  & \new_[57564]_ ;
  assign \new_[57576]_  = A167 & ~A169;
  assign \new_[57577]_  = A170 & \new_[57576]_ ;
  assign \new_[57580]_  = ~A199 & ~A166;
  assign \new_[57583]_  = ~A233 & ~A200;
  assign \new_[57584]_  = \new_[57583]_  & \new_[57580]_ ;
  assign \new_[57585]_  = \new_[57584]_  & \new_[57577]_ ;
  assign \new_[57589]_  = ~A266 & ~A265;
  assign \new_[57590]_  = ~A234 & \new_[57589]_ ;
  assign \new_[57593]_  = ~A299 & A298;
  assign \new_[57596]_  = A302 & A300;
  assign \new_[57597]_  = \new_[57596]_  & \new_[57593]_ ;
  assign \new_[57598]_  = \new_[57597]_  & \new_[57590]_ ;
  assign \new_[57602]_  = A167 & ~A169;
  assign \new_[57603]_  = A170 & \new_[57602]_ ;
  assign \new_[57606]_  = ~A199 & ~A166;
  assign \new_[57609]_  = A232 & ~A200;
  assign \new_[57610]_  = \new_[57609]_  & \new_[57606]_ ;
  assign \new_[57611]_  = \new_[57610]_  & \new_[57603]_ ;
  assign \new_[57615]_  = A235 & A234;
  assign \new_[57616]_  = ~A233 & \new_[57615]_ ;
  assign \new_[57619]_  = ~A266 & A265;
  assign \new_[57622]_  = A268 & A267;
  assign \new_[57623]_  = \new_[57622]_  & \new_[57619]_ ;
  assign \new_[57624]_  = \new_[57623]_  & \new_[57616]_ ;
  assign \new_[57628]_  = A167 & ~A169;
  assign \new_[57629]_  = A170 & \new_[57628]_ ;
  assign \new_[57632]_  = ~A199 & ~A166;
  assign \new_[57635]_  = A232 & ~A200;
  assign \new_[57636]_  = \new_[57635]_  & \new_[57632]_ ;
  assign \new_[57637]_  = \new_[57636]_  & \new_[57629]_ ;
  assign \new_[57641]_  = A235 & A234;
  assign \new_[57642]_  = ~A233 & \new_[57641]_ ;
  assign \new_[57645]_  = ~A266 & A265;
  assign \new_[57648]_  = A269 & A267;
  assign \new_[57649]_  = \new_[57648]_  & \new_[57645]_ ;
  assign \new_[57650]_  = \new_[57649]_  & \new_[57642]_ ;
  assign \new_[57654]_  = A167 & ~A169;
  assign \new_[57655]_  = A170 & \new_[57654]_ ;
  assign \new_[57658]_  = ~A199 & ~A166;
  assign \new_[57661]_  = A232 & ~A200;
  assign \new_[57662]_  = \new_[57661]_  & \new_[57658]_ ;
  assign \new_[57663]_  = \new_[57662]_  & \new_[57655]_ ;
  assign \new_[57667]_  = A236 & A234;
  assign \new_[57668]_  = ~A233 & \new_[57667]_ ;
  assign \new_[57671]_  = ~A266 & A265;
  assign \new_[57674]_  = A268 & A267;
  assign \new_[57675]_  = \new_[57674]_  & \new_[57671]_ ;
  assign \new_[57676]_  = \new_[57675]_  & \new_[57668]_ ;
  assign \new_[57680]_  = A167 & ~A169;
  assign \new_[57681]_  = A170 & \new_[57680]_ ;
  assign \new_[57684]_  = ~A199 & ~A166;
  assign \new_[57687]_  = A232 & ~A200;
  assign \new_[57688]_  = \new_[57687]_  & \new_[57684]_ ;
  assign \new_[57689]_  = \new_[57688]_  & \new_[57681]_ ;
  assign \new_[57693]_  = A236 & A234;
  assign \new_[57694]_  = ~A233 & \new_[57693]_ ;
  assign \new_[57697]_  = ~A266 & A265;
  assign \new_[57700]_  = A269 & A267;
  assign \new_[57701]_  = \new_[57700]_  & \new_[57697]_ ;
  assign \new_[57702]_  = \new_[57701]_  & \new_[57694]_ ;
  assign \new_[57706]_  = A167 & ~A169;
  assign \new_[57707]_  = A170 & \new_[57706]_ ;
  assign \new_[57710]_  = ~A199 & ~A166;
  assign \new_[57713]_  = ~A232 & ~A200;
  assign \new_[57714]_  = \new_[57713]_  & \new_[57710]_ ;
  assign \new_[57715]_  = \new_[57714]_  & \new_[57707]_ ;
  assign \new_[57719]_  = A266 & A265;
  assign \new_[57720]_  = ~A233 & \new_[57719]_ ;
  assign \new_[57723]_  = ~A299 & A298;
  assign \new_[57726]_  = A301 & A300;
  assign \new_[57727]_  = \new_[57726]_  & \new_[57723]_ ;
  assign \new_[57728]_  = \new_[57727]_  & \new_[57720]_ ;
  assign \new_[57732]_  = A167 & ~A169;
  assign \new_[57733]_  = A170 & \new_[57732]_ ;
  assign \new_[57736]_  = ~A199 & ~A166;
  assign \new_[57739]_  = ~A232 & ~A200;
  assign \new_[57740]_  = \new_[57739]_  & \new_[57736]_ ;
  assign \new_[57741]_  = \new_[57740]_  & \new_[57733]_ ;
  assign \new_[57745]_  = A266 & A265;
  assign \new_[57746]_  = ~A233 & \new_[57745]_ ;
  assign \new_[57749]_  = ~A299 & A298;
  assign \new_[57752]_  = A302 & A300;
  assign \new_[57753]_  = \new_[57752]_  & \new_[57749]_ ;
  assign \new_[57754]_  = \new_[57753]_  & \new_[57746]_ ;
  assign \new_[57758]_  = A167 & ~A169;
  assign \new_[57759]_  = A170 & \new_[57758]_ ;
  assign \new_[57762]_  = ~A199 & ~A166;
  assign \new_[57765]_  = ~A232 & ~A200;
  assign \new_[57766]_  = \new_[57765]_  & \new_[57762]_ ;
  assign \new_[57767]_  = \new_[57766]_  & \new_[57759]_ ;
  assign \new_[57771]_  = ~A267 & ~A266;
  assign \new_[57772]_  = ~A233 & \new_[57771]_ ;
  assign \new_[57775]_  = ~A299 & A298;
  assign \new_[57778]_  = A301 & A300;
  assign \new_[57779]_  = \new_[57778]_  & \new_[57775]_ ;
  assign \new_[57780]_  = \new_[57779]_  & \new_[57772]_ ;
  assign \new_[57784]_  = A167 & ~A169;
  assign \new_[57785]_  = A170 & \new_[57784]_ ;
  assign \new_[57788]_  = ~A199 & ~A166;
  assign \new_[57791]_  = ~A232 & ~A200;
  assign \new_[57792]_  = \new_[57791]_  & \new_[57788]_ ;
  assign \new_[57793]_  = \new_[57792]_  & \new_[57785]_ ;
  assign \new_[57797]_  = ~A267 & ~A266;
  assign \new_[57798]_  = ~A233 & \new_[57797]_ ;
  assign \new_[57801]_  = ~A299 & A298;
  assign \new_[57804]_  = A302 & A300;
  assign \new_[57805]_  = \new_[57804]_  & \new_[57801]_ ;
  assign \new_[57806]_  = \new_[57805]_  & \new_[57798]_ ;
  assign \new_[57810]_  = A167 & ~A169;
  assign \new_[57811]_  = A170 & \new_[57810]_ ;
  assign \new_[57814]_  = ~A199 & ~A166;
  assign \new_[57817]_  = ~A232 & ~A200;
  assign \new_[57818]_  = \new_[57817]_  & \new_[57814]_ ;
  assign \new_[57819]_  = \new_[57818]_  & \new_[57811]_ ;
  assign \new_[57823]_  = ~A266 & ~A265;
  assign \new_[57824]_  = ~A233 & \new_[57823]_ ;
  assign \new_[57827]_  = ~A299 & A298;
  assign \new_[57830]_  = A301 & A300;
  assign \new_[57831]_  = \new_[57830]_  & \new_[57827]_ ;
  assign \new_[57832]_  = \new_[57831]_  & \new_[57824]_ ;
  assign \new_[57836]_  = A167 & ~A169;
  assign \new_[57837]_  = A170 & \new_[57836]_ ;
  assign \new_[57840]_  = ~A199 & ~A166;
  assign \new_[57843]_  = ~A232 & ~A200;
  assign \new_[57844]_  = \new_[57843]_  & \new_[57840]_ ;
  assign \new_[57845]_  = \new_[57844]_  & \new_[57837]_ ;
  assign \new_[57849]_  = ~A266 & ~A265;
  assign \new_[57850]_  = ~A233 & \new_[57849]_ ;
  assign \new_[57853]_  = ~A299 & A298;
  assign \new_[57856]_  = A302 & A300;
  assign \new_[57857]_  = \new_[57856]_  & \new_[57853]_ ;
  assign \new_[57858]_  = \new_[57857]_  & \new_[57850]_ ;
  assign \new_[57862]_  = ~A167 & ~A169;
  assign \new_[57863]_  = A170 & \new_[57862]_ ;
  assign \new_[57866]_  = A199 & A166;
  assign \new_[57869]_  = A232 & A200;
  assign \new_[57870]_  = \new_[57869]_  & \new_[57866]_ ;
  assign \new_[57871]_  = \new_[57870]_  & \new_[57863]_ ;
  assign \new_[57875]_  = ~A267 & A265;
  assign \new_[57876]_  = A233 & \new_[57875]_ ;
  assign \new_[57879]_  = ~A299 & A298;
  assign \new_[57882]_  = A301 & A300;
  assign \new_[57883]_  = \new_[57882]_  & \new_[57879]_ ;
  assign \new_[57884]_  = \new_[57883]_  & \new_[57876]_ ;
  assign \new_[57888]_  = ~A167 & ~A169;
  assign \new_[57889]_  = A170 & \new_[57888]_ ;
  assign \new_[57892]_  = A199 & A166;
  assign \new_[57895]_  = A232 & A200;
  assign \new_[57896]_  = \new_[57895]_  & \new_[57892]_ ;
  assign \new_[57897]_  = \new_[57896]_  & \new_[57889]_ ;
  assign \new_[57901]_  = ~A267 & A265;
  assign \new_[57902]_  = A233 & \new_[57901]_ ;
  assign \new_[57905]_  = ~A299 & A298;
  assign \new_[57908]_  = A302 & A300;
  assign \new_[57909]_  = \new_[57908]_  & \new_[57905]_ ;
  assign \new_[57910]_  = \new_[57909]_  & \new_[57902]_ ;
  assign \new_[57914]_  = ~A167 & ~A169;
  assign \new_[57915]_  = A170 & \new_[57914]_ ;
  assign \new_[57918]_  = A199 & A166;
  assign \new_[57921]_  = A232 & A200;
  assign \new_[57922]_  = \new_[57921]_  & \new_[57918]_ ;
  assign \new_[57923]_  = \new_[57922]_  & \new_[57915]_ ;
  assign \new_[57927]_  = A266 & A265;
  assign \new_[57928]_  = A233 & \new_[57927]_ ;
  assign \new_[57931]_  = ~A299 & A298;
  assign \new_[57934]_  = A301 & A300;
  assign \new_[57935]_  = \new_[57934]_  & \new_[57931]_ ;
  assign \new_[57936]_  = \new_[57935]_  & \new_[57928]_ ;
  assign \new_[57940]_  = ~A167 & ~A169;
  assign \new_[57941]_  = A170 & \new_[57940]_ ;
  assign \new_[57944]_  = A199 & A166;
  assign \new_[57947]_  = A232 & A200;
  assign \new_[57948]_  = \new_[57947]_  & \new_[57944]_ ;
  assign \new_[57949]_  = \new_[57948]_  & \new_[57941]_ ;
  assign \new_[57953]_  = A266 & A265;
  assign \new_[57954]_  = A233 & \new_[57953]_ ;
  assign \new_[57957]_  = ~A299 & A298;
  assign \new_[57960]_  = A302 & A300;
  assign \new_[57961]_  = \new_[57960]_  & \new_[57957]_ ;
  assign \new_[57962]_  = \new_[57961]_  & \new_[57954]_ ;
  assign \new_[57966]_  = ~A167 & ~A169;
  assign \new_[57967]_  = A170 & \new_[57966]_ ;
  assign \new_[57970]_  = A199 & A166;
  assign \new_[57973]_  = A232 & A200;
  assign \new_[57974]_  = \new_[57973]_  & \new_[57970]_ ;
  assign \new_[57975]_  = \new_[57974]_  & \new_[57967]_ ;
  assign \new_[57979]_  = ~A266 & ~A265;
  assign \new_[57980]_  = A233 & \new_[57979]_ ;
  assign \new_[57983]_  = ~A299 & A298;
  assign \new_[57986]_  = A301 & A300;
  assign \new_[57987]_  = \new_[57986]_  & \new_[57983]_ ;
  assign \new_[57988]_  = \new_[57987]_  & \new_[57980]_ ;
  assign \new_[57992]_  = ~A167 & ~A169;
  assign \new_[57993]_  = A170 & \new_[57992]_ ;
  assign \new_[57996]_  = A199 & A166;
  assign \new_[57999]_  = A232 & A200;
  assign \new_[58000]_  = \new_[57999]_  & \new_[57996]_ ;
  assign \new_[58001]_  = \new_[58000]_  & \new_[57993]_ ;
  assign \new_[58005]_  = ~A266 & ~A265;
  assign \new_[58006]_  = A233 & \new_[58005]_ ;
  assign \new_[58009]_  = ~A299 & A298;
  assign \new_[58012]_  = A302 & A300;
  assign \new_[58013]_  = \new_[58012]_  & \new_[58009]_ ;
  assign \new_[58014]_  = \new_[58013]_  & \new_[58006]_ ;
  assign \new_[58018]_  = ~A167 & ~A169;
  assign \new_[58019]_  = A170 & \new_[58018]_ ;
  assign \new_[58022]_  = A199 & A166;
  assign \new_[58025]_  = ~A233 & A200;
  assign \new_[58026]_  = \new_[58025]_  & \new_[58022]_ ;
  assign \new_[58027]_  = \new_[58026]_  & \new_[58019]_ ;
  assign \new_[58031]_  = ~A266 & ~A236;
  assign \new_[58032]_  = ~A235 & \new_[58031]_ ;
  assign \new_[58035]_  = ~A269 & ~A268;
  assign \new_[58038]_  = A299 & ~A298;
  assign \new_[58039]_  = \new_[58038]_  & \new_[58035]_ ;
  assign \new_[58040]_  = \new_[58039]_  & \new_[58032]_ ;
  assign \new_[58044]_  = ~A167 & ~A169;
  assign \new_[58045]_  = A170 & \new_[58044]_ ;
  assign \new_[58048]_  = A199 & A166;
  assign \new_[58051]_  = ~A233 & A200;
  assign \new_[58052]_  = \new_[58051]_  & \new_[58048]_ ;
  assign \new_[58053]_  = \new_[58052]_  & \new_[58045]_ ;
  assign \new_[58057]_  = A266 & A265;
  assign \new_[58058]_  = ~A234 & \new_[58057]_ ;
  assign \new_[58061]_  = ~A299 & A298;
  assign \new_[58064]_  = A301 & A300;
  assign \new_[58065]_  = \new_[58064]_  & \new_[58061]_ ;
  assign \new_[58066]_  = \new_[58065]_  & \new_[58058]_ ;
  assign \new_[58070]_  = ~A167 & ~A169;
  assign \new_[58071]_  = A170 & \new_[58070]_ ;
  assign \new_[58074]_  = A199 & A166;
  assign \new_[58077]_  = ~A233 & A200;
  assign \new_[58078]_  = \new_[58077]_  & \new_[58074]_ ;
  assign \new_[58079]_  = \new_[58078]_  & \new_[58071]_ ;
  assign \new_[58083]_  = A266 & A265;
  assign \new_[58084]_  = ~A234 & \new_[58083]_ ;
  assign \new_[58087]_  = ~A299 & A298;
  assign \new_[58090]_  = A302 & A300;
  assign \new_[58091]_  = \new_[58090]_  & \new_[58087]_ ;
  assign \new_[58092]_  = \new_[58091]_  & \new_[58084]_ ;
  assign \new_[58096]_  = ~A167 & ~A169;
  assign \new_[58097]_  = A170 & \new_[58096]_ ;
  assign \new_[58100]_  = A199 & A166;
  assign \new_[58103]_  = ~A233 & A200;
  assign \new_[58104]_  = \new_[58103]_  & \new_[58100]_ ;
  assign \new_[58105]_  = \new_[58104]_  & \new_[58097]_ ;
  assign \new_[58109]_  = ~A267 & ~A266;
  assign \new_[58110]_  = ~A234 & \new_[58109]_ ;
  assign \new_[58113]_  = ~A299 & A298;
  assign \new_[58116]_  = A301 & A300;
  assign \new_[58117]_  = \new_[58116]_  & \new_[58113]_ ;
  assign \new_[58118]_  = \new_[58117]_  & \new_[58110]_ ;
  assign \new_[58122]_  = ~A167 & ~A169;
  assign \new_[58123]_  = A170 & \new_[58122]_ ;
  assign \new_[58126]_  = A199 & A166;
  assign \new_[58129]_  = ~A233 & A200;
  assign \new_[58130]_  = \new_[58129]_  & \new_[58126]_ ;
  assign \new_[58131]_  = \new_[58130]_  & \new_[58123]_ ;
  assign \new_[58135]_  = ~A267 & ~A266;
  assign \new_[58136]_  = ~A234 & \new_[58135]_ ;
  assign \new_[58139]_  = ~A299 & A298;
  assign \new_[58142]_  = A302 & A300;
  assign \new_[58143]_  = \new_[58142]_  & \new_[58139]_ ;
  assign \new_[58144]_  = \new_[58143]_  & \new_[58136]_ ;
  assign \new_[58148]_  = ~A167 & ~A169;
  assign \new_[58149]_  = A170 & \new_[58148]_ ;
  assign \new_[58152]_  = A199 & A166;
  assign \new_[58155]_  = ~A233 & A200;
  assign \new_[58156]_  = \new_[58155]_  & \new_[58152]_ ;
  assign \new_[58157]_  = \new_[58156]_  & \new_[58149]_ ;
  assign \new_[58161]_  = ~A266 & ~A265;
  assign \new_[58162]_  = ~A234 & \new_[58161]_ ;
  assign \new_[58165]_  = ~A299 & A298;
  assign \new_[58168]_  = A301 & A300;
  assign \new_[58169]_  = \new_[58168]_  & \new_[58165]_ ;
  assign \new_[58170]_  = \new_[58169]_  & \new_[58162]_ ;
  assign \new_[58174]_  = ~A167 & ~A169;
  assign \new_[58175]_  = A170 & \new_[58174]_ ;
  assign \new_[58178]_  = A199 & A166;
  assign \new_[58181]_  = ~A233 & A200;
  assign \new_[58182]_  = \new_[58181]_  & \new_[58178]_ ;
  assign \new_[58183]_  = \new_[58182]_  & \new_[58175]_ ;
  assign \new_[58187]_  = ~A266 & ~A265;
  assign \new_[58188]_  = ~A234 & \new_[58187]_ ;
  assign \new_[58191]_  = ~A299 & A298;
  assign \new_[58194]_  = A302 & A300;
  assign \new_[58195]_  = \new_[58194]_  & \new_[58191]_ ;
  assign \new_[58196]_  = \new_[58195]_  & \new_[58188]_ ;
  assign \new_[58200]_  = ~A167 & ~A169;
  assign \new_[58201]_  = A170 & \new_[58200]_ ;
  assign \new_[58204]_  = A199 & A166;
  assign \new_[58207]_  = A232 & A200;
  assign \new_[58208]_  = \new_[58207]_  & \new_[58204]_ ;
  assign \new_[58209]_  = \new_[58208]_  & \new_[58201]_ ;
  assign \new_[58213]_  = A235 & A234;
  assign \new_[58214]_  = ~A233 & \new_[58213]_ ;
  assign \new_[58217]_  = ~A266 & A265;
  assign \new_[58220]_  = A268 & A267;
  assign \new_[58221]_  = \new_[58220]_  & \new_[58217]_ ;
  assign \new_[58222]_  = \new_[58221]_  & \new_[58214]_ ;
  assign \new_[58226]_  = ~A167 & ~A169;
  assign \new_[58227]_  = A170 & \new_[58226]_ ;
  assign \new_[58230]_  = A199 & A166;
  assign \new_[58233]_  = A232 & A200;
  assign \new_[58234]_  = \new_[58233]_  & \new_[58230]_ ;
  assign \new_[58235]_  = \new_[58234]_  & \new_[58227]_ ;
  assign \new_[58239]_  = A235 & A234;
  assign \new_[58240]_  = ~A233 & \new_[58239]_ ;
  assign \new_[58243]_  = ~A266 & A265;
  assign \new_[58246]_  = A269 & A267;
  assign \new_[58247]_  = \new_[58246]_  & \new_[58243]_ ;
  assign \new_[58248]_  = \new_[58247]_  & \new_[58240]_ ;
  assign \new_[58252]_  = ~A167 & ~A169;
  assign \new_[58253]_  = A170 & \new_[58252]_ ;
  assign \new_[58256]_  = A199 & A166;
  assign \new_[58259]_  = A232 & A200;
  assign \new_[58260]_  = \new_[58259]_  & \new_[58256]_ ;
  assign \new_[58261]_  = \new_[58260]_  & \new_[58253]_ ;
  assign \new_[58265]_  = A236 & A234;
  assign \new_[58266]_  = ~A233 & \new_[58265]_ ;
  assign \new_[58269]_  = ~A266 & A265;
  assign \new_[58272]_  = A268 & A267;
  assign \new_[58273]_  = \new_[58272]_  & \new_[58269]_ ;
  assign \new_[58274]_  = \new_[58273]_  & \new_[58266]_ ;
  assign \new_[58278]_  = ~A167 & ~A169;
  assign \new_[58279]_  = A170 & \new_[58278]_ ;
  assign \new_[58282]_  = A199 & A166;
  assign \new_[58285]_  = A232 & A200;
  assign \new_[58286]_  = \new_[58285]_  & \new_[58282]_ ;
  assign \new_[58287]_  = \new_[58286]_  & \new_[58279]_ ;
  assign \new_[58291]_  = A236 & A234;
  assign \new_[58292]_  = ~A233 & \new_[58291]_ ;
  assign \new_[58295]_  = ~A266 & A265;
  assign \new_[58298]_  = A269 & A267;
  assign \new_[58299]_  = \new_[58298]_  & \new_[58295]_ ;
  assign \new_[58300]_  = \new_[58299]_  & \new_[58292]_ ;
  assign \new_[58304]_  = ~A167 & ~A169;
  assign \new_[58305]_  = A170 & \new_[58304]_ ;
  assign \new_[58308]_  = A199 & A166;
  assign \new_[58311]_  = ~A232 & A200;
  assign \new_[58312]_  = \new_[58311]_  & \new_[58308]_ ;
  assign \new_[58313]_  = \new_[58312]_  & \new_[58305]_ ;
  assign \new_[58317]_  = A266 & A265;
  assign \new_[58318]_  = ~A233 & \new_[58317]_ ;
  assign \new_[58321]_  = ~A299 & A298;
  assign \new_[58324]_  = A301 & A300;
  assign \new_[58325]_  = \new_[58324]_  & \new_[58321]_ ;
  assign \new_[58326]_  = \new_[58325]_  & \new_[58318]_ ;
  assign \new_[58330]_  = ~A167 & ~A169;
  assign \new_[58331]_  = A170 & \new_[58330]_ ;
  assign \new_[58334]_  = A199 & A166;
  assign \new_[58337]_  = ~A232 & A200;
  assign \new_[58338]_  = \new_[58337]_  & \new_[58334]_ ;
  assign \new_[58339]_  = \new_[58338]_  & \new_[58331]_ ;
  assign \new_[58343]_  = A266 & A265;
  assign \new_[58344]_  = ~A233 & \new_[58343]_ ;
  assign \new_[58347]_  = ~A299 & A298;
  assign \new_[58350]_  = A302 & A300;
  assign \new_[58351]_  = \new_[58350]_  & \new_[58347]_ ;
  assign \new_[58352]_  = \new_[58351]_  & \new_[58344]_ ;
  assign \new_[58356]_  = ~A167 & ~A169;
  assign \new_[58357]_  = A170 & \new_[58356]_ ;
  assign \new_[58360]_  = A199 & A166;
  assign \new_[58363]_  = ~A232 & A200;
  assign \new_[58364]_  = \new_[58363]_  & \new_[58360]_ ;
  assign \new_[58365]_  = \new_[58364]_  & \new_[58357]_ ;
  assign \new_[58369]_  = ~A267 & ~A266;
  assign \new_[58370]_  = ~A233 & \new_[58369]_ ;
  assign \new_[58373]_  = ~A299 & A298;
  assign \new_[58376]_  = A301 & A300;
  assign \new_[58377]_  = \new_[58376]_  & \new_[58373]_ ;
  assign \new_[58378]_  = \new_[58377]_  & \new_[58370]_ ;
  assign \new_[58382]_  = ~A167 & ~A169;
  assign \new_[58383]_  = A170 & \new_[58382]_ ;
  assign \new_[58386]_  = A199 & A166;
  assign \new_[58389]_  = ~A232 & A200;
  assign \new_[58390]_  = \new_[58389]_  & \new_[58386]_ ;
  assign \new_[58391]_  = \new_[58390]_  & \new_[58383]_ ;
  assign \new_[58395]_  = ~A267 & ~A266;
  assign \new_[58396]_  = ~A233 & \new_[58395]_ ;
  assign \new_[58399]_  = ~A299 & A298;
  assign \new_[58402]_  = A302 & A300;
  assign \new_[58403]_  = \new_[58402]_  & \new_[58399]_ ;
  assign \new_[58404]_  = \new_[58403]_  & \new_[58396]_ ;
  assign \new_[58408]_  = ~A167 & ~A169;
  assign \new_[58409]_  = A170 & \new_[58408]_ ;
  assign \new_[58412]_  = A199 & A166;
  assign \new_[58415]_  = ~A232 & A200;
  assign \new_[58416]_  = \new_[58415]_  & \new_[58412]_ ;
  assign \new_[58417]_  = \new_[58416]_  & \new_[58409]_ ;
  assign \new_[58421]_  = ~A266 & ~A265;
  assign \new_[58422]_  = ~A233 & \new_[58421]_ ;
  assign \new_[58425]_  = ~A299 & A298;
  assign \new_[58428]_  = A301 & A300;
  assign \new_[58429]_  = \new_[58428]_  & \new_[58425]_ ;
  assign \new_[58430]_  = \new_[58429]_  & \new_[58422]_ ;
  assign \new_[58434]_  = ~A167 & ~A169;
  assign \new_[58435]_  = A170 & \new_[58434]_ ;
  assign \new_[58438]_  = A199 & A166;
  assign \new_[58441]_  = ~A232 & A200;
  assign \new_[58442]_  = \new_[58441]_  & \new_[58438]_ ;
  assign \new_[58443]_  = \new_[58442]_  & \new_[58435]_ ;
  assign \new_[58447]_  = ~A266 & ~A265;
  assign \new_[58448]_  = ~A233 & \new_[58447]_ ;
  assign \new_[58451]_  = ~A299 & A298;
  assign \new_[58454]_  = A302 & A300;
  assign \new_[58455]_  = \new_[58454]_  & \new_[58451]_ ;
  assign \new_[58456]_  = \new_[58455]_  & \new_[58448]_ ;
  assign \new_[58460]_  = ~A167 & ~A169;
  assign \new_[58461]_  = A170 & \new_[58460]_ ;
  assign \new_[58464]_  = ~A200 & A166;
  assign \new_[58467]_  = ~A203 & ~A202;
  assign \new_[58468]_  = \new_[58467]_  & \new_[58464]_ ;
  assign \new_[58469]_  = \new_[58468]_  & \new_[58461]_ ;
  assign \new_[58473]_  = A265 & A233;
  assign \new_[58474]_  = A232 & \new_[58473]_ ;
  assign \new_[58477]_  = ~A269 & ~A268;
  assign \new_[58480]_  = A299 & ~A298;
  assign \new_[58481]_  = \new_[58480]_  & \new_[58477]_ ;
  assign \new_[58482]_  = \new_[58481]_  & \new_[58474]_ ;
  assign \new_[58486]_  = ~A167 & ~A169;
  assign \new_[58487]_  = A170 & \new_[58486]_ ;
  assign \new_[58490]_  = ~A200 & A166;
  assign \new_[58493]_  = ~A203 & ~A202;
  assign \new_[58494]_  = \new_[58493]_  & \new_[58490]_ ;
  assign \new_[58495]_  = \new_[58494]_  & \new_[58487]_ ;
  assign \new_[58499]_  = ~A236 & ~A235;
  assign \new_[58500]_  = ~A233 & \new_[58499]_ ;
  assign \new_[58503]_  = A266 & A265;
  assign \new_[58506]_  = A299 & ~A298;
  assign \new_[58507]_  = \new_[58506]_  & \new_[58503]_ ;
  assign \new_[58508]_  = \new_[58507]_  & \new_[58500]_ ;
  assign \new_[58512]_  = ~A167 & ~A169;
  assign \new_[58513]_  = A170 & \new_[58512]_ ;
  assign \new_[58516]_  = ~A200 & A166;
  assign \new_[58519]_  = ~A203 & ~A202;
  assign \new_[58520]_  = \new_[58519]_  & \new_[58516]_ ;
  assign \new_[58521]_  = \new_[58520]_  & \new_[58513]_ ;
  assign \new_[58525]_  = ~A236 & ~A235;
  assign \new_[58526]_  = ~A233 & \new_[58525]_ ;
  assign \new_[58529]_  = ~A267 & ~A266;
  assign \new_[58532]_  = A299 & ~A298;
  assign \new_[58533]_  = \new_[58532]_  & \new_[58529]_ ;
  assign \new_[58534]_  = \new_[58533]_  & \new_[58526]_ ;
  assign \new_[58538]_  = ~A167 & ~A169;
  assign \new_[58539]_  = A170 & \new_[58538]_ ;
  assign \new_[58542]_  = ~A200 & A166;
  assign \new_[58545]_  = ~A203 & ~A202;
  assign \new_[58546]_  = \new_[58545]_  & \new_[58542]_ ;
  assign \new_[58547]_  = \new_[58546]_  & \new_[58539]_ ;
  assign \new_[58551]_  = ~A236 & ~A235;
  assign \new_[58552]_  = ~A233 & \new_[58551]_ ;
  assign \new_[58555]_  = ~A266 & ~A265;
  assign \new_[58558]_  = A299 & ~A298;
  assign \new_[58559]_  = \new_[58558]_  & \new_[58555]_ ;
  assign \new_[58560]_  = \new_[58559]_  & \new_[58552]_ ;
  assign \new_[58564]_  = ~A167 & ~A169;
  assign \new_[58565]_  = A170 & \new_[58564]_ ;
  assign \new_[58568]_  = ~A200 & A166;
  assign \new_[58571]_  = ~A203 & ~A202;
  assign \new_[58572]_  = \new_[58571]_  & \new_[58568]_ ;
  assign \new_[58573]_  = \new_[58572]_  & \new_[58565]_ ;
  assign \new_[58577]_  = ~A266 & ~A234;
  assign \new_[58578]_  = ~A233 & \new_[58577]_ ;
  assign \new_[58581]_  = ~A269 & ~A268;
  assign \new_[58584]_  = A299 & ~A298;
  assign \new_[58585]_  = \new_[58584]_  & \new_[58581]_ ;
  assign \new_[58586]_  = \new_[58585]_  & \new_[58578]_ ;
  assign \new_[58590]_  = ~A167 & ~A169;
  assign \new_[58591]_  = A170 & \new_[58590]_ ;
  assign \new_[58594]_  = ~A200 & A166;
  assign \new_[58597]_  = ~A203 & ~A202;
  assign \new_[58598]_  = \new_[58597]_  & \new_[58594]_ ;
  assign \new_[58599]_  = \new_[58598]_  & \new_[58591]_ ;
  assign \new_[58603]_  = A234 & ~A233;
  assign \new_[58604]_  = A232 & \new_[58603]_ ;
  assign \new_[58607]_  = A298 & A235;
  assign \new_[58610]_  = ~A302 & ~A301;
  assign \new_[58611]_  = \new_[58610]_  & \new_[58607]_ ;
  assign \new_[58612]_  = \new_[58611]_  & \new_[58604]_ ;
  assign \new_[58616]_  = ~A167 & ~A169;
  assign \new_[58617]_  = A170 & \new_[58616]_ ;
  assign \new_[58620]_  = ~A200 & A166;
  assign \new_[58623]_  = ~A203 & ~A202;
  assign \new_[58624]_  = \new_[58623]_  & \new_[58620]_ ;
  assign \new_[58625]_  = \new_[58624]_  & \new_[58617]_ ;
  assign \new_[58629]_  = A234 & ~A233;
  assign \new_[58630]_  = A232 & \new_[58629]_ ;
  assign \new_[58633]_  = A298 & A236;
  assign \new_[58636]_  = ~A302 & ~A301;
  assign \new_[58637]_  = \new_[58636]_  & \new_[58633]_ ;
  assign \new_[58638]_  = \new_[58637]_  & \new_[58630]_ ;
  assign \new_[58642]_  = ~A167 & ~A169;
  assign \new_[58643]_  = A170 & \new_[58642]_ ;
  assign \new_[58646]_  = ~A200 & A166;
  assign \new_[58649]_  = ~A203 & ~A202;
  assign \new_[58650]_  = \new_[58649]_  & \new_[58646]_ ;
  assign \new_[58651]_  = \new_[58650]_  & \new_[58643]_ ;
  assign \new_[58655]_  = ~A266 & ~A233;
  assign \new_[58656]_  = ~A232 & \new_[58655]_ ;
  assign \new_[58659]_  = ~A269 & ~A268;
  assign \new_[58662]_  = A299 & ~A298;
  assign \new_[58663]_  = \new_[58662]_  & \new_[58659]_ ;
  assign \new_[58664]_  = \new_[58663]_  & \new_[58656]_ ;
  assign \new_[58668]_  = ~A167 & ~A169;
  assign \new_[58669]_  = A170 & \new_[58668]_ ;
  assign \new_[58672]_  = ~A200 & A166;
  assign \new_[58675]_  = A232 & ~A201;
  assign \new_[58676]_  = \new_[58675]_  & \new_[58672]_ ;
  assign \new_[58677]_  = \new_[58676]_  & \new_[58669]_ ;
  assign \new_[58681]_  = ~A267 & A265;
  assign \new_[58682]_  = A233 & \new_[58681]_ ;
  assign \new_[58685]_  = ~A299 & A298;
  assign \new_[58688]_  = A301 & A300;
  assign \new_[58689]_  = \new_[58688]_  & \new_[58685]_ ;
  assign \new_[58690]_  = \new_[58689]_  & \new_[58682]_ ;
  assign \new_[58694]_  = ~A167 & ~A169;
  assign \new_[58695]_  = A170 & \new_[58694]_ ;
  assign \new_[58698]_  = ~A200 & A166;
  assign \new_[58701]_  = A232 & ~A201;
  assign \new_[58702]_  = \new_[58701]_  & \new_[58698]_ ;
  assign \new_[58703]_  = \new_[58702]_  & \new_[58695]_ ;
  assign \new_[58707]_  = ~A267 & A265;
  assign \new_[58708]_  = A233 & \new_[58707]_ ;
  assign \new_[58711]_  = ~A299 & A298;
  assign \new_[58714]_  = A302 & A300;
  assign \new_[58715]_  = \new_[58714]_  & \new_[58711]_ ;
  assign \new_[58716]_  = \new_[58715]_  & \new_[58708]_ ;
  assign \new_[58720]_  = ~A167 & ~A169;
  assign \new_[58721]_  = A170 & \new_[58720]_ ;
  assign \new_[58724]_  = ~A200 & A166;
  assign \new_[58727]_  = A232 & ~A201;
  assign \new_[58728]_  = \new_[58727]_  & \new_[58724]_ ;
  assign \new_[58729]_  = \new_[58728]_  & \new_[58721]_ ;
  assign \new_[58733]_  = A266 & A265;
  assign \new_[58734]_  = A233 & \new_[58733]_ ;
  assign \new_[58737]_  = ~A299 & A298;
  assign \new_[58740]_  = A301 & A300;
  assign \new_[58741]_  = \new_[58740]_  & \new_[58737]_ ;
  assign \new_[58742]_  = \new_[58741]_  & \new_[58734]_ ;
  assign \new_[58746]_  = ~A167 & ~A169;
  assign \new_[58747]_  = A170 & \new_[58746]_ ;
  assign \new_[58750]_  = ~A200 & A166;
  assign \new_[58753]_  = A232 & ~A201;
  assign \new_[58754]_  = \new_[58753]_  & \new_[58750]_ ;
  assign \new_[58755]_  = \new_[58754]_  & \new_[58747]_ ;
  assign \new_[58759]_  = A266 & A265;
  assign \new_[58760]_  = A233 & \new_[58759]_ ;
  assign \new_[58763]_  = ~A299 & A298;
  assign \new_[58766]_  = A302 & A300;
  assign \new_[58767]_  = \new_[58766]_  & \new_[58763]_ ;
  assign \new_[58768]_  = \new_[58767]_  & \new_[58760]_ ;
  assign \new_[58772]_  = ~A167 & ~A169;
  assign \new_[58773]_  = A170 & \new_[58772]_ ;
  assign \new_[58776]_  = ~A200 & A166;
  assign \new_[58779]_  = A232 & ~A201;
  assign \new_[58780]_  = \new_[58779]_  & \new_[58776]_ ;
  assign \new_[58781]_  = \new_[58780]_  & \new_[58773]_ ;
  assign \new_[58785]_  = ~A266 & ~A265;
  assign \new_[58786]_  = A233 & \new_[58785]_ ;
  assign \new_[58789]_  = ~A299 & A298;
  assign \new_[58792]_  = A301 & A300;
  assign \new_[58793]_  = \new_[58792]_  & \new_[58789]_ ;
  assign \new_[58794]_  = \new_[58793]_  & \new_[58786]_ ;
  assign \new_[58798]_  = ~A167 & ~A169;
  assign \new_[58799]_  = A170 & \new_[58798]_ ;
  assign \new_[58802]_  = ~A200 & A166;
  assign \new_[58805]_  = A232 & ~A201;
  assign \new_[58806]_  = \new_[58805]_  & \new_[58802]_ ;
  assign \new_[58807]_  = \new_[58806]_  & \new_[58799]_ ;
  assign \new_[58811]_  = ~A266 & ~A265;
  assign \new_[58812]_  = A233 & \new_[58811]_ ;
  assign \new_[58815]_  = ~A299 & A298;
  assign \new_[58818]_  = A302 & A300;
  assign \new_[58819]_  = \new_[58818]_  & \new_[58815]_ ;
  assign \new_[58820]_  = \new_[58819]_  & \new_[58812]_ ;
  assign \new_[58824]_  = ~A167 & ~A169;
  assign \new_[58825]_  = A170 & \new_[58824]_ ;
  assign \new_[58828]_  = ~A200 & A166;
  assign \new_[58831]_  = ~A233 & ~A201;
  assign \new_[58832]_  = \new_[58831]_  & \new_[58828]_ ;
  assign \new_[58833]_  = \new_[58832]_  & \new_[58825]_ ;
  assign \new_[58837]_  = ~A266 & ~A236;
  assign \new_[58838]_  = ~A235 & \new_[58837]_ ;
  assign \new_[58841]_  = ~A269 & ~A268;
  assign \new_[58844]_  = A299 & ~A298;
  assign \new_[58845]_  = \new_[58844]_  & \new_[58841]_ ;
  assign \new_[58846]_  = \new_[58845]_  & \new_[58838]_ ;
  assign \new_[58850]_  = ~A167 & ~A169;
  assign \new_[58851]_  = A170 & \new_[58850]_ ;
  assign \new_[58854]_  = ~A200 & A166;
  assign \new_[58857]_  = ~A233 & ~A201;
  assign \new_[58858]_  = \new_[58857]_  & \new_[58854]_ ;
  assign \new_[58859]_  = \new_[58858]_  & \new_[58851]_ ;
  assign \new_[58863]_  = A266 & A265;
  assign \new_[58864]_  = ~A234 & \new_[58863]_ ;
  assign \new_[58867]_  = ~A299 & A298;
  assign \new_[58870]_  = A301 & A300;
  assign \new_[58871]_  = \new_[58870]_  & \new_[58867]_ ;
  assign \new_[58872]_  = \new_[58871]_  & \new_[58864]_ ;
  assign \new_[58876]_  = ~A167 & ~A169;
  assign \new_[58877]_  = A170 & \new_[58876]_ ;
  assign \new_[58880]_  = ~A200 & A166;
  assign \new_[58883]_  = ~A233 & ~A201;
  assign \new_[58884]_  = \new_[58883]_  & \new_[58880]_ ;
  assign \new_[58885]_  = \new_[58884]_  & \new_[58877]_ ;
  assign \new_[58889]_  = A266 & A265;
  assign \new_[58890]_  = ~A234 & \new_[58889]_ ;
  assign \new_[58893]_  = ~A299 & A298;
  assign \new_[58896]_  = A302 & A300;
  assign \new_[58897]_  = \new_[58896]_  & \new_[58893]_ ;
  assign \new_[58898]_  = \new_[58897]_  & \new_[58890]_ ;
  assign \new_[58902]_  = ~A167 & ~A169;
  assign \new_[58903]_  = A170 & \new_[58902]_ ;
  assign \new_[58906]_  = ~A200 & A166;
  assign \new_[58909]_  = ~A233 & ~A201;
  assign \new_[58910]_  = \new_[58909]_  & \new_[58906]_ ;
  assign \new_[58911]_  = \new_[58910]_  & \new_[58903]_ ;
  assign \new_[58915]_  = ~A267 & ~A266;
  assign \new_[58916]_  = ~A234 & \new_[58915]_ ;
  assign \new_[58919]_  = ~A299 & A298;
  assign \new_[58922]_  = A301 & A300;
  assign \new_[58923]_  = \new_[58922]_  & \new_[58919]_ ;
  assign \new_[58924]_  = \new_[58923]_  & \new_[58916]_ ;
  assign \new_[58928]_  = ~A167 & ~A169;
  assign \new_[58929]_  = A170 & \new_[58928]_ ;
  assign \new_[58932]_  = ~A200 & A166;
  assign \new_[58935]_  = ~A233 & ~A201;
  assign \new_[58936]_  = \new_[58935]_  & \new_[58932]_ ;
  assign \new_[58937]_  = \new_[58936]_  & \new_[58929]_ ;
  assign \new_[58941]_  = ~A267 & ~A266;
  assign \new_[58942]_  = ~A234 & \new_[58941]_ ;
  assign \new_[58945]_  = ~A299 & A298;
  assign \new_[58948]_  = A302 & A300;
  assign \new_[58949]_  = \new_[58948]_  & \new_[58945]_ ;
  assign \new_[58950]_  = \new_[58949]_  & \new_[58942]_ ;
  assign \new_[58954]_  = ~A167 & ~A169;
  assign \new_[58955]_  = A170 & \new_[58954]_ ;
  assign \new_[58958]_  = ~A200 & A166;
  assign \new_[58961]_  = ~A233 & ~A201;
  assign \new_[58962]_  = \new_[58961]_  & \new_[58958]_ ;
  assign \new_[58963]_  = \new_[58962]_  & \new_[58955]_ ;
  assign \new_[58967]_  = ~A266 & ~A265;
  assign \new_[58968]_  = ~A234 & \new_[58967]_ ;
  assign \new_[58971]_  = ~A299 & A298;
  assign \new_[58974]_  = A301 & A300;
  assign \new_[58975]_  = \new_[58974]_  & \new_[58971]_ ;
  assign \new_[58976]_  = \new_[58975]_  & \new_[58968]_ ;
  assign \new_[58980]_  = ~A167 & ~A169;
  assign \new_[58981]_  = A170 & \new_[58980]_ ;
  assign \new_[58984]_  = ~A200 & A166;
  assign \new_[58987]_  = ~A233 & ~A201;
  assign \new_[58988]_  = \new_[58987]_  & \new_[58984]_ ;
  assign \new_[58989]_  = \new_[58988]_  & \new_[58981]_ ;
  assign \new_[58993]_  = ~A266 & ~A265;
  assign \new_[58994]_  = ~A234 & \new_[58993]_ ;
  assign \new_[58997]_  = ~A299 & A298;
  assign \new_[59000]_  = A302 & A300;
  assign \new_[59001]_  = \new_[59000]_  & \new_[58997]_ ;
  assign \new_[59002]_  = \new_[59001]_  & \new_[58994]_ ;
  assign \new_[59006]_  = ~A167 & ~A169;
  assign \new_[59007]_  = A170 & \new_[59006]_ ;
  assign \new_[59010]_  = ~A200 & A166;
  assign \new_[59013]_  = A232 & ~A201;
  assign \new_[59014]_  = \new_[59013]_  & \new_[59010]_ ;
  assign \new_[59015]_  = \new_[59014]_  & \new_[59007]_ ;
  assign \new_[59019]_  = A235 & A234;
  assign \new_[59020]_  = ~A233 & \new_[59019]_ ;
  assign \new_[59023]_  = ~A266 & A265;
  assign \new_[59026]_  = A268 & A267;
  assign \new_[59027]_  = \new_[59026]_  & \new_[59023]_ ;
  assign \new_[59028]_  = \new_[59027]_  & \new_[59020]_ ;
  assign \new_[59032]_  = ~A167 & ~A169;
  assign \new_[59033]_  = A170 & \new_[59032]_ ;
  assign \new_[59036]_  = ~A200 & A166;
  assign \new_[59039]_  = A232 & ~A201;
  assign \new_[59040]_  = \new_[59039]_  & \new_[59036]_ ;
  assign \new_[59041]_  = \new_[59040]_  & \new_[59033]_ ;
  assign \new_[59045]_  = A235 & A234;
  assign \new_[59046]_  = ~A233 & \new_[59045]_ ;
  assign \new_[59049]_  = ~A266 & A265;
  assign \new_[59052]_  = A269 & A267;
  assign \new_[59053]_  = \new_[59052]_  & \new_[59049]_ ;
  assign \new_[59054]_  = \new_[59053]_  & \new_[59046]_ ;
  assign \new_[59058]_  = ~A167 & ~A169;
  assign \new_[59059]_  = A170 & \new_[59058]_ ;
  assign \new_[59062]_  = ~A200 & A166;
  assign \new_[59065]_  = A232 & ~A201;
  assign \new_[59066]_  = \new_[59065]_  & \new_[59062]_ ;
  assign \new_[59067]_  = \new_[59066]_  & \new_[59059]_ ;
  assign \new_[59071]_  = A236 & A234;
  assign \new_[59072]_  = ~A233 & \new_[59071]_ ;
  assign \new_[59075]_  = ~A266 & A265;
  assign \new_[59078]_  = A268 & A267;
  assign \new_[59079]_  = \new_[59078]_  & \new_[59075]_ ;
  assign \new_[59080]_  = \new_[59079]_  & \new_[59072]_ ;
  assign \new_[59084]_  = ~A167 & ~A169;
  assign \new_[59085]_  = A170 & \new_[59084]_ ;
  assign \new_[59088]_  = ~A200 & A166;
  assign \new_[59091]_  = A232 & ~A201;
  assign \new_[59092]_  = \new_[59091]_  & \new_[59088]_ ;
  assign \new_[59093]_  = \new_[59092]_  & \new_[59085]_ ;
  assign \new_[59097]_  = A236 & A234;
  assign \new_[59098]_  = ~A233 & \new_[59097]_ ;
  assign \new_[59101]_  = ~A266 & A265;
  assign \new_[59104]_  = A269 & A267;
  assign \new_[59105]_  = \new_[59104]_  & \new_[59101]_ ;
  assign \new_[59106]_  = \new_[59105]_  & \new_[59098]_ ;
  assign \new_[59110]_  = ~A167 & ~A169;
  assign \new_[59111]_  = A170 & \new_[59110]_ ;
  assign \new_[59114]_  = ~A200 & A166;
  assign \new_[59117]_  = ~A232 & ~A201;
  assign \new_[59118]_  = \new_[59117]_  & \new_[59114]_ ;
  assign \new_[59119]_  = \new_[59118]_  & \new_[59111]_ ;
  assign \new_[59123]_  = A266 & A265;
  assign \new_[59124]_  = ~A233 & \new_[59123]_ ;
  assign \new_[59127]_  = ~A299 & A298;
  assign \new_[59130]_  = A301 & A300;
  assign \new_[59131]_  = \new_[59130]_  & \new_[59127]_ ;
  assign \new_[59132]_  = \new_[59131]_  & \new_[59124]_ ;
  assign \new_[59136]_  = ~A167 & ~A169;
  assign \new_[59137]_  = A170 & \new_[59136]_ ;
  assign \new_[59140]_  = ~A200 & A166;
  assign \new_[59143]_  = ~A232 & ~A201;
  assign \new_[59144]_  = \new_[59143]_  & \new_[59140]_ ;
  assign \new_[59145]_  = \new_[59144]_  & \new_[59137]_ ;
  assign \new_[59149]_  = A266 & A265;
  assign \new_[59150]_  = ~A233 & \new_[59149]_ ;
  assign \new_[59153]_  = ~A299 & A298;
  assign \new_[59156]_  = A302 & A300;
  assign \new_[59157]_  = \new_[59156]_  & \new_[59153]_ ;
  assign \new_[59158]_  = \new_[59157]_  & \new_[59150]_ ;
  assign \new_[59162]_  = ~A167 & ~A169;
  assign \new_[59163]_  = A170 & \new_[59162]_ ;
  assign \new_[59166]_  = ~A200 & A166;
  assign \new_[59169]_  = ~A232 & ~A201;
  assign \new_[59170]_  = \new_[59169]_  & \new_[59166]_ ;
  assign \new_[59171]_  = \new_[59170]_  & \new_[59163]_ ;
  assign \new_[59175]_  = ~A267 & ~A266;
  assign \new_[59176]_  = ~A233 & \new_[59175]_ ;
  assign \new_[59179]_  = ~A299 & A298;
  assign \new_[59182]_  = A301 & A300;
  assign \new_[59183]_  = \new_[59182]_  & \new_[59179]_ ;
  assign \new_[59184]_  = \new_[59183]_  & \new_[59176]_ ;
  assign \new_[59188]_  = ~A167 & ~A169;
  assign \new_[59189]_  = A170 & \new_[59188]_ ;
  assign \new_[59192]_  = ~A200 & A166;
  assign \new_[59195]_  = ~A232 & ~A201;
  assign \new_[59196]_  = \new_[59195]_  & \new_[59192]_ ;
  assign \new_[59197]_  = \new_[59196]_  & \new_[59189]_ ;
  assign \new_[59201]_  = ~A267 & ~A266;
  assign \new_[59202]_  = ~A233 & \new_[59201]_ ;
  assign \new_[59205]_  = ~A299 & A298;
  assign \new_[59208]_  = A302 & A300;
  assign \new_[59209]_  = \new_[59208]_  & \new_[59205]_ ;
  assign \new_[59210]_  = \new_[59209]_  & \new_[59202]_ ;
  assign \new_[59214]_  = ~A167 & ~A169;
  assign \new_[59215]_  = A170 & \new_[59214]_ ;
  assign \new_[59218]_  = ~A200 & A166;
  assign \new_[59221]_  = ~A232 & ~A201;
  assign \new_[59222]_  = \new_[59221]_  & \new_[59218]_ ;
  assign \new_[59223]_  = \new_[59222]_  & \new_[59215]_ ;
  assign \new_[59227]_  = ~A266 & ~A265;
  assign \new_[59228]_  = ~A233 & \new_[59227]_ ;
  assign \new_[59231]_  = ~A299 & A298;
  assign \new_[59234]_  = A301 & A300;
  assign \new_[59235]_  = \new_[59234]_  & \new_[59231]_ ;
  assign \new_[59236]_  = \new_[59235]_  & \new_[59228]_ ;
  assign \new_[59240]_  = ~A167 & ~A169;
  assign \new_[59241]_  = A170 & \new_[59240]_ ;
  assign \new_[59244]_  = ~A200 & A166;
  assign \new_[59247]_  = ~A232 & ~A201;
  assign \new_[59248]_  = \new_[59247]_  & \new_[59244]_ ;
  assign \new_[59249]_  = \new_[59248]_  & \new_[59241]_ ;
  assign \new_[59253]_  = ~A266 & ~A265;
  assign \new_[59254]_  = ~A233 & \new_[59253]_ ;
  assign \new_[59257]_  = ~A299 & A298;
  assign \new_[59260]_  = A302 & A300;
  assign \new_[59261]_  = \new_[59260]_  & \new_[59257]_ ;
  assign \new_[59262]_  = \new_[59261]_  & \new_[59254]_ ;
  assign \new_[59266]_  = ~A167 & ~A169;
  assign \new_[59267]_  = A170 & \new_[59266]_ ;
  assign \new_[59270]_  = ~A199 & A166;
  assign \new_[59273]_  = A232 & ~A200;
  assign \new_[59274]_  = \new_[59273]_  & \new_[59270]_ ;
  assign \new_[59275]_  = \new_[59274]_  & \new_[59267]_ ;
  assign \new_[59279]_  = ~A267 & A265;
  assign \new_[59280]_  = A233 & \new_[59279]_ ;
  assign \new_[59283]_  = ~A299 & A298;
  assign \new_[59286]_  = A301 & A300;
  assign \new_[59287]_  = \new_[59286]_  & \new_[59283]_ ;
  assign \new_[59288]_  = \new_[59287]_  & \new_[59280]_ ;
  assign \new_[59292]_  = ~A167 & ~A169;
  assign \new_[59293]_  = A170 & \new_[59292]_ ;
  assign \new_[59296]_  = ~A199 & A166;
  assign \new_[59299]_  = A232 & ~A200;
  assign \new_[59300]_  = \new_[59299]_  & \new_[59296]_ ;
  assign \new_[59301]_  = \new_[59300]_  & \new_[59293]_ ;
  assign \new_[59305]_  = ~A267 & A265;
  assign \new_[59306]_  = A233 & \new_[59305]_ ;
  assign \new_[59309]_  = ~A299 & A298;
  assign \new_[59312]_  = A302 & A300;
  assign \new_[59313]_  = \new_[59312]_  & \new_[59309]_ ;
  assign \new_[59314]_  = \new_[59313]_  & \new_[59306]_ ;
  assign \new_[59318]_  = ~A167 & ~A169;
  assign \new_[59319]_  = A170 & \new_[59318]_ ;
  assign \new_[59322]_  = ~A199 & A166;
  assign \new_[59325]_  = A232 & ~A200;
  assign \new_[59326]_  = \new_[59325]_  & \new_[59322]_ ;
  assign \new_[59327]_  = \new_[59326]_  & \new_[59319]_ ;
  assign \new_[59331]_  = A266 & A265;
  assign \new_[59332]_  = A233 & \new_[59331]_ ;
  assign \new_[59335]_  = ~A299 & A298;
  assign \new_[59338]_  = A301 & A300;
  assign \new_[59339]_  = \new_[59338]_  & \new_[59335]_ ;
  assign \new_[59340]_  = \new_[59339]_  & \new_[59332]_ ;
  assign \new_[59344]_  = ~A167 & ~A169;
  assign \new_[59345]_  = A170 & \new_[59344]_ ;
  assign \new_[59348]_  = ~A199 & A166;
  assign \new_[59351]_  = A232 & ~A200;
  assign \new_[59352]_  = \new_[59351]_  & \new_[59348]_ ;
  assign \new_[59353]_  = \new_[59352]_  & \new_[59345]_ ;
  assign \new_[59357]_  = A266 & A265;
  assign \new_[59358]_  = A233 & \new_[59357]_ ;
  assign \new_[59361]_  = ~A299 & A298;
  assign \new_[59364]_  = A302 & A300;
  assign \new_[59365]_  = \new_[59364]_  & \new_[59361]_ ;
  assign \new_[59366]_  = \new_[59365]_  & \new_[59358]_ ;
  assign \new_[59370]_  = ~A167 & ~A169;
  assign \new_[59371]_  = A170 & \new_[59370]_ ;
  assign \new_[59374]_  = ~A199 & A166;
  assign \new_[59377]_  = A232 & ~A200;
  assign \new_[59378]_  = \new_[59377]_  & \new_[59374]_ ;
  assign \new_[59379]_  = \new_[59378]_  & \new_[59371]_ ;
  assign \new_[59383]_  = ~A266 & ~A265;
  assign \new_[59384]_  = A233 & \new_[59383]_ ;
  assign \new_[59387]_  = ~A299 & A298;
  assign \new_[59390]_  = A301 & A300;
  assign \new_[59391]_  = \new_[59390]_  & \new_[59387]_ ;
  assign \new_[59392]_  = \new_[59391]_  & \new_[59384]_ ;
  assign \new_[59396]_  = ~A167 & ~A169;
  assign \new_[59397]_  = A170 & \new_[59396]_ ;
  assign \new_[59400]_  = ~A199 & A166;
  assign \new_[59403]_  = A232 & ~A200;
  assign \new_[59404]_  = \new_[59403]_  & \new_[59400]_ ;
  assign \new_[59405]_  = \new_[59404]_  & \new_[59397]_ ;
  assign \new_[59409]_  = ~A266 & ~A265;
  assign \new_[59410]_  = A233 & \new_[59409]_ ;
  assign \new_[59413]_  = ~A299 & A298;
  assign \new_[59416]_  = A302 & A300;
  assign \new_[59417]_  = \new_[59416]_  & \new_[59413]_ ;
  assign \new_[59418]_  = \new_[59417]_  & \new_[59410]_ ;
  assign \new_[59422]_  = ~A167 & ~A169;
  assign \new_[59423]_  = A170 & \new_[59422]_ ;
  assign \new_[59426]_  = ~A199 & A166;
  assign \new_[59429]_  = ~A233 & ~A200;
  assign \new_[59430]_  = \new_[59429]_  & \new_[59426]_ ;
  assign \new_[59431]_  = \new_[59430]_  & \new_[59423]_ ;
  assign \new_[59435]_  = ~A266 & ~A236;
  assign \new_[59436]_  = ~A235 & \new_[59435]_ ;
  assign \new_[59439]_  = ~A269 & ~A268;
  assign \new_[59442]_  = A299 & ~A298;
  assign \new_[59443]_  = \new_[59442]_  & \new_[59439]_ ;
  assign \new_[59444]_  = \new_[59443]_  & \new_[59436]_ ;
  assign \new_[59448]_  = ~A167 & ~A169;
  assign \new_[59449]_  = A170 & \new_[59448]_ ;
  assign \new_[59452]_  = ~A199 & A166;
  assign \new_[59455]_  = ~A233 & ~A200;
  assign \new_[59456]_  = \new_[59455]_  & \new_[59452]_ ;
  assign \new_[59457]_  = \new_[59456]_  & \new_[59449]_ ;
  assign \new_[59461]_  = A266 & A265;
  assign \new_[59462]_  = ~A234 & \new_[59461]_ ;
  assign \new_[59465]_  = ~A299 & A298;
  assign \new_[59468]_  = A301 & A300;
  assign \new_[59469]_  = \new_[59468]_  & \new_[59465]_ ;
  assign \new_[59470]_  = \new_[59469]_  & \new_[59462]_ ;
  assign \new_[59474]_  = ~A167 & ~A169;
  assign \new_[59475]_  = A170 & \new_[59474]_ ;
  assign \new_[59478]_  = ~A199 & A166;
  assign \new_[59481]_  = ~A233 & ~A200;
  assign \new_[59482]_  = \new_[59481]_  & \new_[59478]_ ;
  assign \new_[59483]_  = \new_[59482]_  & \new_[59475]_ ;
  assign \new_[59487]_  = A266 & A265;
  assign \new_[59488]_  = ~A234 & \new_[59487]_ ;
  assign \new_[59491]_  = ~A299 & A298;
  assign \new_[59494]_  = A302 & A300;
  assign \new_[59495]_  = \new_[59494]_  & \new_[59491]_ ;
  assign \new_[59496]_  = \new_[59495]_  & \new_[59488]_ ;
  assign \new_[59500]_  = ~A167 & ~A169;
  assign \new_[59501]_  = A170 & \new_[59500]_ ;
  assign \new_[59504]_  = ~A199 & A166;
  assign \new_[59507]_  = ~A233 & ~A200;
  assign \new_[59508]_  = \new_[59507]_  & \new_[59504]_ ;
  assign \new_[59509]_  = \new_[59508]_  & \new_[59501]_ ;
  assign \new_[59513]_  = ~A267 & ~A266;
  assign \new_[59514]_  = ~A234 & \new_[59513]_ ;
  assign \new_[59517]_  = ~A299 & A298;
  assign \new_[59520]_  = A301 & A300;
  assign \new_[59521]_  = \new_[59520]_  & \new_[59517]_ ;
  assign \new_[59522]_  = \new_[59521]_  & \new_[59514]_ ;
  assign \new_[59526]_  = ~A167 & ~A169;
  assign \new_[59527]_  = A170 & \new_[59526]_ ;
  assign \new_[59530]_  = ~A199 & A166;
  assign \new_[59533]_  = ~A233 & ~A200;
  assign \new_[59534]_  = \new_[59533]_  & \new_[59530]_ ;
  assign \new_[59535]_  = \new_[59534]_  & \new_[59527]_ ;
  assign \new_[59539]_  = ~A267 & ~A266;
  assign \new_[59540]_  = ~A234 & \new_[59539]_ ;
  assign \new_[59543]_  = ~A299 & A298;
  assign \new_[59546]_  = A302 & A300;
  assign \new_[59547]_  = \new_[59546]_  & \new_[59543]_ ;
  assign \new_[59548]_  = \new_[59547]_  & \new_[59540]_ ;
  assign \new_[59552]_  = ~A167 & ~A169;
  assign \new_[59553]_  = A170 & \new_[59552]_ ;
  assign \new_[59556]_  = ~A199 & A166;
  assign \new_[59559]_  = ~A233 & ~A200;
  assign \new_[59560]_  = \new_[59559]_  & \new_[59556]_ ;
  assign \new_[59561]_  = \new_[59560]_  & \new_[59553]_ ;
  assign \new_[59565]_  = ~A266 & ~A265;
  assign \new_[59566]_  = ~A234 & \new_[59565]_ ;
  assign \new_[59569]_  = ~A299 & A298;
  assign \new_[59572]_  = A301 & A300;
  assign \new_[59573]_  = \new_[59572]_  & \new_[59569]_ ;
  assign \new_[59574]_  = \new_[59573]_  & \new_[59566]_ ;
  assign \new_[59578]_  = ~A167 & ~A169;
  assign \new_[59579]_  = A170 & \new_[59578]_ ;
  assign \new_[59582]_  = ~A199 & A166;
  assign \new_[59585]_  = ~A233 & ~A200;
  assign \new_[59586]_  = \new_[59585]_  & \new_[59582]_ ;
  assign \new_[59587]_  = \new_[59586]_  & \new_[59579]_ ;
  assign \new_[59591]_  = ~A266 & ~A265;
  assign \new_[59592]_  = ~A234 & \new_[59591]_ ;
  assign \new_[59595]_  = ~A299 & A298;
  assign \new_[59598]_  = A302 & A300;
  assign \new_[59599]_  = \new_[59598]_  & \new_[59595]_ ;
  assign \new_[59600]_  = \new_[59599]_  & \new_[59592]_ ;
  assign \new_[59604]_  = ~A167 & ~A169;
  assign \new_[59605]_  = A170 & \new_[59604]_ ;
  assign \new_[59608]_  = ~A199 & A166;
  assign \new_[59611]_  = A232 & ~A200;
  assign \new_[59612]_  = \new_[59611]_  & \new_[59608]_ ;
  assign \new_[59613]_  = \new_[59612]_  & \new_[59605]_ ;
  assign \new_[59617]_  = A235 & A234;
  assign \new_[59618]_  = ~A233 & \new_[59617]_ ;
  assign \new_[59621]_  = ~A266 & A265;
  assign \new_[59624]_  = A268 & A267;
  assign \new_[59625]_  = \new_[59624]_  & \new_[59621]_ ;
  assign \new_[59626]_  = \new_[59625]_  & \new_[59618]_ ;
  assign \new_[59630]_  = ~A167 & ~A169;
  assign \new_[59631]_  = A170 & \new_[59630]_ ;
  assign \new_[59634]_  = ~A199 & A166;
  assign \new_[59637]_  = A232 & ~A200;
  assign \new_[59638]_  = \new_[59637]_  & \new_[59634]_ ;
  assign \new_[59639]_  = \new_[59638]_  & \new_[59631]_ ;
  assign \new_[59643]_  = A235 & A234;
  assign \new_[59644]_  = ~A233 & \new_[59643]_ ;
  assign \new_[59647]_  = ~A266 & A265;
  assign \new_[59650]_  = A269 & A267;
  assign \new_[59651]_  = \new_[59650]_  & \new_[59647]_ ;
  assign \new_[59652]_  = \new_[59651]_  & \new_[59644]_ ;
  assign \new_[59656]_  = ~A167 & ~A169;
  assign \new_[59657]_  = A170 & \new_[59656]_ ;
  assign \new_[59660]_  = ~A199 & A166;
  assign \new_[59663]_  = A232 & ~A200;
  assign \new_[59664]_  = \new_[59663]_  & \new_[59660]_ ;
  assign \new_[59665]_  = \new_[59664]_  & \new_[59657]_ ;
  assign \new_[59669]_  = A236 & A234;
  assign \new_[59670]_  = ~A233 & \new_[59669]_ ;
  assign \new_[59673]_  = ~A266 & A265;
  assign \new_[59676]_  = A268 & A267;
  assign \new_[59677]_  = \new_[59676]_  & \new_[59673]_ ;
  assign \new_[59678]_  = \new_[59677]_  & \new_[59670]_ ;
  assign \new_[59682]_  = ~A167 & ~A169;
  assign \new_[59683]_  = A170 & \new_[59682]_ ;
  assign \new_[59686]_  = ~A199 & A166;
  assign \new_[59689]_  = A232 & ~A200;
  assign \new_[59690]_  = \new_[59689]_  & \new_[59686]_ ;
  assign \new_[59691]_  = \new_[59690]_  & \new_[59683]_ ;
  assign \new_[59695]_  = A236 & A234;
  assign \new_[59696]_  = ~A233 & \new_[59695]_ ;
  assign \new_[59699]_  = ~A266 & A265;
  assign \new_[59702]_  = A269 & A267;
  assign \new_[59703]_  = \new_[59702]_  & \new_[59699]_ ;
  assign \new_[59704]_  = \new_[59703]_  & \new_[59696]_ ;
  assign \new_[59708]_  = ~A167 & ~A169;
  assign \new_[59709]_  = A170 & \new_[59708]_ ;
  assign \new_[59712]_  = ~A199 & A166;
  assign \new_[59715]_  = ~A232 & ~A200;
  assign \new_[59716]_  = \new_[59715]_  & \new_[59712]_ ;
  assign \new_[59717]_  = \new_[59716]_  & \new_[59709]_ ;
  assign \new_[59721]_  = A266 & A265;
  assign \new_[59722]_  = ~A233 & \new_[59721]_ ;
  assign \new_[59725]_  = ~A299 & A298;
  assign \new_[59728]_  = A301 & A300;
  assign \new_[59729]_  = \new_[59728]_  & \new_[59725]_ ;
  assign \new_[59730]_  = \new_[59729]_  & \new_[59722]_ ;
  assign \new_[59734]_  = ~A167 & ~A169;
  assign \new_[59735]_  = A170 & \new_[59734]_ ;
  assign \new_[59738]_  = ~A199 & A166;
  assign \new_[59741]_  = ~A232 & ~A200;
  assign \new_[59742]_  = \new_[59741]_  & \new_[59738]_ ;
  assign \new_[59743]_  = \new_[59742]_  & \new_[59735]_ ;
  assign \new_[59747]_  = A266 & A265;
  assign \new_[59748]_  = ~A233 & \new_[59747]_ ;
  assign \new_[59751]_  = ~A299 & A298;
  assign \new_[59754]_  = A302 & A300;
  assign \new_[59755]_  = \new_[59754]_  & \new_[59751]_ ;
  assign \new_[59756]_  = \new_[59755]_  & \new_[59748]_ ;
  assign \new_[59760]_  = ~A167 & ~A169;
  assign \new_[59761]_  = A170 & \new_[59760]_ ;
  assign \new_[59764]_  = ~A199 & A166;
  assign \new_[59767]_  = ~A232 & ~A200;
  assign \new_[59768]_  = \new_[59767]_  & \new_[59764]_ ;
  assign \new_[59769]_  = \new_[59768]_  & \new_[59761]_ ;
  assign \new_[59773]_  = ~A267 & ~A266;
  assign \new_[59774]_  = ~A233 & \new_[59773]_ ;
  assign \new_[59777]_  = ~A299 & A298;
  assign \new_[59780]_  = A301 & A300;
  assign \new_[59781]_  = \new_[59780]_  & \new_[59777]_ ;
  assign \new_[59782]_  = \new_[59781]_  & \new_[59774]_ ;
  assign \new_[59786]_  = ~A167 & ~A169;
  assign \new_[59787]_  = A170 & \new_[59786]_ ;
  assign \new_[59790]_  = ~A199 & A166;
  assign \new_[59793]_  = ~A232 & ~A200;
  assign \new_[59794]_  = \new_[59793]_  & \new_[59790]_ ;
  assign \new_[59795]_  = \new_[59794]_  & \new_[59787]_ ;
  assign \new_[59799]_  = ~A267 & ~A266;
  assign \new_[59800]_  = ~A233 & \new_[59799]_ ;
  assign \new_[59803]_  = ~A299 & A298;
  assign \new_[59806]_  = A302 & A300;
  assign \new_[59807]_  = \new_[59806]_  & \new_[59803]_ ;
  assign \new_[59808]_  = \new_[59807]_  & \new_[59800]_ ;
  assign \new_[59812]_  = ~A167 & ~A169;
  assign \new_[59813]_  = A170 & \new_[59812]_ ;
  assign \new_[59816]_  = ~A199 & A166;
  assign \new_[59819]_  = ~A232 & ~A200;
  assign \new_[59820]_  = \new_[59819]_  & \new_[59816]_ ;
  assign \new_[59821]_  = \new_[59820]_  & \new_[59813]_ ;
  assign \new_[59825]_  = ~A266 & ~A265;
  assign \new_[59826]_  = ~A233 & \new_[59825]_ ;
  assign \new_[59829]_  = ~A299 & A298;
  assign \new_[59832]_  = A301 & A300;
  assign \new_[59833]_  = \new_[59832]_  & \new_[59829]_ ;
  assign \new_[59834]_  = \new_[59833]_  & \new_[59826]_ ;
  assign \new_[59838]_  = ~A167 & ~A169;
  assign \new_[59839]_  = A170 & \new_[59838]_ ;
  assign \new_[59842]_  = ~A199 & A166;
  assign \new_[59845]_  = ~A232 & ~A200;
  assign \new_[59846]_  = \new_[59845]_  & \new_[59842]_ ;
  assign \new_[59847]_  = \new_[59846]_  & \new_[59839]_ ;
  assign \new_[59851]_  = ~A266 & ~A265;
  assign \new_[59852]_  = ~A233 & \new_[59851]_ ;
  assign \new_[59855]_  = ~A299 & A298;
  assign \new_[59858]_  = A302 & A300;
  assign \new_[59859]_  = \new_[59858]_  & \new_[59855]_ ;
  assign \new_[59860]_  = \new_[59859]_  & \new_[59852]_ ;
  assign \new_[59864]_  = ~A168 & ~A169;
  assign \new_[59865]_  = ~A170 & \new_[59864]_ ;
  assign \new_[59868]_  = ~A200 & A199;
  assign \new_[59871]_  = A202 & A201;
  assign \new_[59872]_  = \new_[59871]_  & \new_[59868]_ ;
  assign \new_[59873]_  = \new_[59872]_  & \new_[59865]_ ;
  assign \new_[59877]_  = A265 & A233;
  assign \new_[59878]_  = A232 & \new_[59877]_ ;
  assign \new_[59881]_  = ~A269 & ~A268;
  assign \new_[59884]_  = A299 & ~A298;
  assign \new_[59885]_  = \new_[59884]_  & \new_[59881]_ ;
  assign \new_[59886]_  = \new_[59885]_  & \new_[59878]_ ;
  assign \new_[59890]_  = ~A168 & ~A169;
  assign \new_[59891]_  = ~A170 & \new_[59890]_ ;
  assign \new_[59894]_  = ~A200 & A199;
  assign \new_[59897]_  = A202 & A201;
  assign \new_[59898]_  = \new_[59897]_  & \new_[59894]_ ;
  assign \new_[59899]_  = \new_[59898]_  & \new_[59891]_ ;
  assign \new_[59903]_  = ~A236 & ~A235;
  assign \new_[59904]_  = ~A233 & \new_[59903]_ ;
  assign \new_[59907]_  = A266 & A265;
  assign \new_[59910]_  = A299 & ~A298;
  assign \new_[59911]_  = \new_[59910]_  & \new_[59907]_ ;
  assign \new_[59912]_  = \new_[59911]_  & \new_[59904]_ ;
  assign \new_[59916]_  = ~A168 & ~A169;
  assign \new_[59917]_  = ~A170 & \new_[59916]_ ;
  assign \new_[59920]_  = ~A200 & A199;
  assign \new_[59923]_  = A202 & A201;
  assign \new_[59924]_  = \new_[59923]_  & \new_[59920]_ ;
  assign \new_[59925]_  = \new_[59924]_  & \new_[59917]_ ;
  assign \new_[59929]_  = ~A236 & ~A235;
  assign \new_[59930]_  = ~A233 & \new_[59929]_ ;
  assign \new_[59933]_  = ~A267 & ~A266;
  assign \new_[59936]_  = A299 & ~A298;
  assign \new_[59937]_  = \new_[59936]_  & \new_[59933]_ ;
  assign \new_[59938]_  = \new_[59937]_  & \new_[59930]_ ;
  assign \new_[59942]_  = ~A168 & ~A169;
  assign \new_[59943]_  = ~A170 & \new_[59942]_ ;
  assign \new_[59946]_  = ~A200 & A199;
  assign \new_[59949]_  = A202 & A201;
  assign \new_[59950]_  = \new_[59949]_  & \new_[59946]_ ;
  assign \new_[59951]_  = \new_[59950]_  & \new_[59943]_ ;
  assign \new_[59955]_  = ~A236 & ~A235;
  assign \new_[59956]_  = ~A233 & \new_[59955]_ ;
  assign \new_[59959]_  = ~A266 & ~A265;
  assign \new_[59962]_  = A299 & ~A298;
  assign \new_[59963]_  = \new_[59962]_  & \new_[59959]_ ;
  assign \new_[59964]_  = \new_[59963]_  & \new_[59956]_ ;
  assign \new_[59968]_  = ~A168 & ~A169;
  assign \new_[59969]_  = ~A170 & \new_[59968]_ ;
  assign \new_[59972]_  = ~A200 & A199;
  assign \new_[59975]_  = A202 & A201;
  assign \new_[59976]_  = \new_[59975]_  & \new_[59972]_ ;
  assign \new_[59977]_  = \new_[59976]_  & \new_[59969]_ ;
  assign \new_[59981]_  = ~A266 & ~A234;
  assign \new_[59982]_  = ~A233 & \new_[59981]_ ;
  assign \new_[59985]_  = ~A269 & ~A268;
  assign \new_[59988]_  = A299 & ~A298;
  assign \new_[59989]_  = \new_[59988]_  & \new_[59985]_ ;
  assign \new_[59990]_  = \new_[59989]_  & \new_[59982]_ ;
  assign \new_[59994]_  = ~A168 & ~A169;
  assign \new_[59995]_  = ~A170 & \new_[59994]_ ;
  assign \new_[59998]_  = ~A200 & A199;
  assign \new_[60001]_  = A202 & A201;
  assign \new_[60002]_  = \new_[60001]_  & \new_[59998]_ ;
  assign \new_[60003]_  = \new_[60002]_  & \new_[59995]_ ;
  assign \new_[60007]_  = A234 & ~A233;
  assign \new_[60008]_  = A232 & \new_[60007]_ ;
  assign \new_[60011]_  = A298 & A235;
  assign \new_[60014]_  = ~A302 & ~A301;
  assign \new_[60015]_  = \new_[60014]_  & \new_[60011]_ ;
  assign \new_[60016]_  = \new_[60015]_  & \new_[60008]_ ;
  assign \new_[60020]_  = ~A168 & ~A169;
  assign \new_[60021]_  = ~A170 & \new_[60020]_ ;
  assign \new_[60024]_  = ~A200 & A199;
  assign \new_[60027]_  = A202 & A201;
  assign \new_[60028]_  = \new_[60027]_  & \new_[60024]_ ;
  assign \new_[60029]_  = \new_[60028]_  & \new_[60021]_ ;
  assign \new_[60033]_  = A234 & ~A233;
  assign \new_[60034]_  = A232 & \new_[60033]_ ;
  assign \new_[60037]_  = A298 & A236;
  assign \new_[60040]_  = ~A302 & ~A301;
  assign \new_[60041]_  = \new_[60040]_  & \new_[60037]_ ;
  assign \new_[60042]_  = \new_[60041]_  & \new_[60034]_ ;
  assign \new_[60046]_  = ~A168 & ~A169;
  assign \new_[60047]_  = ~A170 & \new_[60046]_ ;
  assign \new_[60050]_  = ~A200 & A199;
  assign \new_[60053]_  = A202 & A201;
  assign \new_[60054]_  = \new_[60053]_  & \new_[60050]_ ;
  assign \new_[60055]_  = \new_[60054]_  & \new_[60047]_ ;
  assign \new_[60059]_  = ~A266 & ~A233;
  assign \new_[60060]_  = ~A232 & \new_[60059]_ ;
  assign \new_[60063]_  = ~A269 & ~A268;
  assign \new_[60066]_  = A299 & ~A298;
  assign \new_[60067]_  = \new_[60066]_  & \new_[60063]_ ;
  assign \new_[60068]_  = \new_[60067]_  & \new_[60060]_ ;
  assign \new_[60072]_  = ~A168 & ~A169;
  assign \new_[60073]_  = ~A170 & \new_[60072]_ ;
  assign \new_[60076]_  = ~A200 & A199;
  assign \new_[60079]_  = A203 & A201;
  assign \new_[60080]_  = \new_[60079]_  & \new_[60076]_ ;
  assign \new_[60081]_  = \new_[60080]_  & \new_[60073]_ ;
  assign \new_[60085]_  = A265 & A233;
  assign \new_[60086]_  = A232 & \new_[60085]_ ;
  assign \new_[60089]_  = ~A269 & ~A268;
  assign \new_[60092]_  = A299 & ~A298;
  assign \new_[60093]_  = \new_[60092]_  & \new_[60089]_ ;
  assign \new_[60094]_  = \new_[60093]_  & \new_[60086]_ ;
  assign \new_[60098]_  = ~A168 & ~A169;
  assign \new_[60099]_  = ~A170 & \new_[60098]_ ;
  assign \new_[60102]_  = ~A200 & A199;
  assign \new_[60105]_  = A203 & A201;
  assign \new_[60106]_  = \new_[60105]_  & \new_[60102]_ ;
  assign \new_[60107]_  = \new_[60106]_  & \new_[60099]_ ;
  assign \new_[60111]_  = ~A236 & ~A235;
  assign \new_[60112]_  = ~A233 & \new_[60111]_ ;
  assign \new_[60115]_  = A266 & A265;
  assign \new_[60118]_  = A299 & ~A298;
  assign \new_[60119]_  = \new_[60118]_  & \new_[60115]_ ;
  assign \new_[60120]_  = \new_[60119]_  & \new_[60112]_ ;
  assign \new_[60124]_  = ~A168 & ~A169;
  assign \new_[60125]_  = ~A170 & \new_[60124]_ ;
  assign \new_[60128]_  = ~A200 & A199;
  assign \new_[60131]_  = A203 & A201;
  assign \new_[60132]_  = \new_[60131]_  & \new_[60128]_ ;
  assign \new_[60133]_  = \new_[60132]_  & \new_[60125]_ ;
  assign \new_[60137]_  = ~A236 & ~A235;
  assign \new_[60138]_  = ~A233 & \new_[60137]_ ;
  assign \new_[60141]_  = ~A267 & ~A266;
  assign \new_[60144]_  = A299 & ~A298;
  assign \new_[60145]_  = \new_[60144]_  & \new_[60141]_ ;
  assign \new_[60146]_  = \new_[60145]_  & \new_[60138]_ ;
  assign \new_[60150]_  = ~A168 & ~A169;
  assign \new_[60151]_  = ~A170 & \new_[60150]_ ;
  assign \new_[60154]_  = ~A200 & A199;
  assign \new_[60157]_  = A203 & A201;
  assign \new_[60158]_  = \new_[60157]_  & \new_[60154]_ ;
  assign \new_[60159]_  = \new_[60158]_  & \new_[60151]_ ;
  assign \new_[60163]_  = ~A236 & ~A235;
  assign \new_[60164]_  = ~A233 & \new_[60163]_ ;
  assign \new_[60167]_  = ~A266 & ~A265;
  assign \new_[60170]_  = A299 & ~A298;
  assign \new_[60171]_  = \new_[60170]_  & \new_[60167]_ ;
  assign \new_[60172]_  = \new_[60171]_  & \new_[60164]_ ;
  assign \new_[60176]_  = ~A168 & ~A169;
  assign \new_[60177]_  = ~A170 & \new_[60176]_ ;
  assign \new_[60180]_  = ~A200 & A199;
  assign \new_[60183]_  = A203 & A201;
  assign \new_[60184]_  = \new_[60183]_  & \new_[60180]_ ;
  assign \new_[60185]_  = \new_[60184]_  & \new_[60177]_ ;
  assign \new_[60189]_  = ~A266 & ~A234;
  assign \new_[60190]_  = ~A233 & \new_[60189]_ ;
  assign \new_[60193]_  = ~A269 & ~A268;
  assign \new_[60196]_  = A299 & ~A298;
  assign \new_[60197]_  = \new_[60196]_  & \new_[60193]_ ;
  assign \new_[60198]_  = \new_[60197]_  & \new_[60190]_ ;
  assign \new_[60202]_  = ~A168 & ~A169;
  assign \new_[60203]_  = ~A170 & \new_[60202]_ ;
  assign \new_[60206]_  = ~A200 & A199;
  assign \new_[60209]_  = A203 & A201;
  assign \new_[60210]_  = \new_[60209]_  & \new_[60206]_ ;
  assign \new_[60211]_  = \new_[60210]_  & \new_[60203]_ ;
  assign \new_[60215]_  = A234 & ~A233;
  assign \new_[60216]_  = A232 & \new_[60215]_ ;
  assign \new_[60219]_  = A298 & A235;
  assign \new_[60222]_  = ~A302 & ~A301;
  assign \new_[60223]_  = \new_[60222]_  & \new_[60219]_ ;
  assign \new_[60224]_  = \new_[60223]_  & \new_[60216]_ ;
  assign \new_[60228]_  = ~A168 & ~A169;
  assign \new_[60229]_  = ~A170 & \new_[60228]_ ;
  assign \new_[60232]_  = ~A200 & A199;
  assign \new_[60235]_  = A203 & A201;
  assign \new_[60236]_  = \new_[60235]_  & \new_[60232]_ ;
  assign \new_[60237]_  = \new_[60236]_  & \new_[60229]_ ;
  assign \new_[60241]_  = A234 & ~A233;
  assign \new_[60242]_  = A232 & \new_[60241]_ ;
  assign \new_[60245]_  = A298 & A236;
  assign \new_[60248]_  = ~A302 & ~A301;
  assign \new_[60249]_  = \new_[60248]_  & \new_[60245]_ ;
  assign \new_[60250]_  = \new_[60249]_  & \new_[60242]_ ;
  assign \new_[60254]_  = ~A168 & ~A169;
  assign \new_[60255]_  = ~A170 & \new_[60254]_ ;
  assign \new_[60258]_  = ~A200 & A199;
  assign \new_[60261]_  = A203 & A201;
  assign \new_[60262]_  = \new_[60261]_  & \new_[60258]_ ;
  assign \new_[60263]_  = \new_[60262]_  & \new_[60255]_ ;
  assign \new_[60267]_  = ~A266 & ~A233;
  assign \new_[60268]_  = ~A232 & \new_[60267]_ ;
  assign \new_[60271]_  = ~A269 & ~A268;
  assign \new_[60274]_  = A299 & ~A298;
  assign \new_[60275]_  = \new_[60274]_  & \new_[60271]_ ;
  assign \new_[60276]_  = \new_[60275]_  & \new_[60268]_ ;
  assign \new_[60280]_  = ~A200 & A166;
  assign \new_[60281]_  = A168 & \new_[60280]_ ;
  assign \new_[60284]_  = ~A203 & ~A202;
  assign \new_[60287]_  = ~A235 & ~A233;
  assign \new_[60288]_  = \new_[60287]_  & \new_[60284]_ ;
  assign \new_[60289]_  = \new_[60288]_  & \new_[60281]_ ;
  assign \new_[60292]_  = ~A266 & ~A236;
  assign \new_[60295]_  = ~A269 & ~A268;
  assign \new_[60296]_  = \new_[60295]_  & \new_[60292]_ ;
  assign \new_[60299]_  = ~A299 & A298;
  assign \new_[60302]_  = A301 & A300;
  assign \new_[60303]_  = \new_[60302]_  & \new_[60299]_ ;
  assign \new_[60304]_  = \new_[60303]_  & \new_[60296]_ ;
  assign \new_[60308]_  = ~A200 & A166;
  assign \new_[60309]_  = A168 & \new_[60308]_ ;
  assign \new_[60312]_  = ~A203 & ~A202;
  assign \new_[60315]_  = ~A235 & ~A233;
  assign \new_[60316]_  = \new_[60315]_  & \new_[60312]_ ;
  assign \new_[60317]_  = \new_[60316]_  & \new_[60309]_ ;
  assign \new_[60320]_  = ~A266 & ~A236;
  assign \new_[60323]_  = ~A269 & ~A268;
  assign \new_[60324]_  = \new_[60323]_  & \new_[60320]_ ;
  assign \new_[60327]_  = ~A299 & A298;
  assign \new_[60330]_  = A302 & A300;
  assign \new_[60331]_  = \new_[60330]_  & \new_[60327]_ ;
  assign \new_[60332]_  = \new_[60331]_  & \new_[60324]_ ;
  assign \new_[60336]_  = ~A200 & A167;
  assign \new_[60337]_  = A168 & \new_[60336]_ ;
  assign \new_[60340]_  = ~A203 & ~A202;
  assign \new_[60343]_  = ~A235 & ~A233;
  assign \new_[60344]_  = \new_[60343]_  & \new_[60340]_ ;
  assign \new_[60345]_  = \new_[60344]_  & \new_[60337]_ ;
  assign \new_[60348]_  = ~A266 & ~A236;
  assign \new_[60351]_  = ~A269 & ~A268;
  assign \new_[60352]_  = \new_[60351]_  & \new_[60348]_ ;
  assign \new_[60355]_  = ~A299 & A298;
  assign \new_[60358]_  = A301 & A300;
  assign \new_[60359]_  = \new_[60358]_  & \new_[60355]_ ;
  assign \new_[60360]_  = \new_[60359]_  & \new_[60352]_ ;
  assign \new_[60364]_  = ~A200 & A167;
  assign \new_[60365]_  = A168 & \new_[60364]_ ;
  assign \new_[60368]_  = ~A203 & ~A202;
  assign \new_[60371]_  = ~A235 & ~A233;
  assign \new_[60372]_  = \new_[60371]_  & \new_[60368]_ ;
  assign \new_[60373]_  = \new_[60372]_  & \new_[60365]_ ;
  assign \new_[60376]_  = ~A266 & ~A236;
  assign \new_[60379]_  = ~A269 & ~A268;
  assign \new_[60380]_  = \new_[60379]_  & \new_[60376]_ ;
  assign \new_[60383]_  = ~A299 & A298;
  assign \new_[60386]_  = A302 & A300;
  assign \new_[60387]_  = \new_[60386]_  & \new_[60383]_ ;
  assign \new_[60388]_  = \new_[60387]_  & \new_[60380]_ ;
  assign \new_[60392]_  = ~A166 & ~A167;
  assign \new_[60393]_  = A170 & \new_[60392]_ ;
  assign \new_[60396]_  = A200 & ~A199;
  assign \new_[60399]_  = ~A235 & ~A233;
  assign \new_[60400]_  = \new_[60399]_  & \new_[60396]_ ;
  assign \new_[60401]_  = \new_[60400]_  & \new_[60393]_ ;
  assign \new_[60404]_  = ~A266 & ~A236;
  assign \new_[60407]_  = ~A269 & ~A268;
  assign \new_[60408]_  = \new_[60407]_  & \new_[60404]_ ;
  assign \new_[60411]_  = ~A299 & A298;
  assign \new_[60414]_  = A301 & A300;
  assign \new_[60415]_  = \new_[60414]_  & \new_[60411]_ ;
  assign \new_[60416]_  = \new_[60415]_  & \new_[60408]_ ;
  assign \new_[60420]_  = ~A166 & ~A167;
  assign \new_[60421]_  = A170 & \new_[60420]_ ;
  assign \new_[60424]_  = A200 & ~A199;
  assign \new_[60427]_  = ~A235 & ~A233;
  assign \new_[60428]_  = \new_[60427]_  & \new_[60424]_ ;
  assign \new_[60429]_  = \new_[60428]_  & \new_[60421]_ ;
  assign \new_[60432]_  = ~A266 & ~A236;
  assign \new_[60435]_  = ~A269 & ~A268;
  assign \new_[60436]_  = \new_[60435]_  & \new_[60432]_ ;
  assign \new_[60439]_  = ~A299 & A298;
  assign \new_[60442]_  = A302 & A300;
  assign \new_[60443]_  = \new_[60442]_  & \new_[60439]_ ;
  assign \new_[60444]_  = \new_[60443]_  & \new_[60436]_ ;
  assign \new_[60448]_  = ~A166 & ~A167;
  assign \new_[60449]_  = A170 & \new_[60448]_ ;
  assign \new_[60452]_  = ~A200 & A199;
  assign \new_[60455]_  = A202 & A201;
  assign \new_[60456]_  = \new_[60455]_  & \new_[60452]_ ;
  assign \new_[60457]_  = \new_[60456]_  & \new_[60449]_ ;
  assign \new_[60460]_  = A233 & A232;
  assign \new_[60463]_  = ~A267 & A265;
  assign \new_[60464]_  = \new_[60463]_  & \new_[60460]_ ;
  assign \new_[60467]_  = ~A299 & A298;
  assign \new_[60470]_  = A301 & A300;
  assign \new_[60471]_  = \new_[60470]_  & \new_[60467]_ ;
  assign \new_[60472]_  = \new_[60471]_  & \new_[60464]_ ;
  assign \new_[60476]_  = ~A166 & ~A167;
  assign \new_[60477]_  = A170 & \new_[60476]_ ;
  assign \new_[60480]_  = ~A200 & A199;
  assign \new_[60483]_  = A202 & A201;
  assign \new_[60484]_  = \new_[60483]_  & \new_[60480]_ ;
  assign \new_[60485]_  = \new_[60484]_  & \new_[60477]_ ;
  assign \new_[60488]_  = A233 & A232;
  assign \new_[60491]_  = ~A267 & A265;
  assign \new_[60492]_  = \new_[60491]_  & \new_[60488]_ ;
  assign \new_[60495]_  = ~A299 & A298;
  assign \new_[60498]_  = A302 & A300;
  assign \new_[60499]_  = \new_[60498]_  & \new_[60495]_ ;
  assign \new_[60500]_  = \new_[60499]_  & \new_[60492]_ ;
  assign \new_[60504]_  = ~A166 & ~A167;
  assign \new_[60505]_  = A170 & \new_[60504]_ ;
  assign \new_[60508]_  = ~A200 & A199;
  assign \new_[60511]_  = A202 & A201;
  assign \new_[60512]_  = \new_[60511]_  & \new_[60508]_ ;
  assign \new_[60513]_  = \new_[60512]_  & \new_[60505]_ ;
  assign \new_[60516]_  = A233 & A232;
  assign \new_[60519]_  = A266 & A265;
  assign \new_[60520]_  = \new_[60519]_  & \new_[60516]_ ;
  assign \new_[60523]_  = ~A299 & A298;
  assign \new_[60526]_  = A301 & A300;
  assign \new_[60527]_  = \new_[60526]_  & \new_[60523]_ ;
  assign \new_[60528]_  = \new_[60527]_  & \new_[60520]_ ;
  assign \new_[60532]_  = ~A166 & ~A167;
  assign \new_[60533]_  = A170 & \new_[60532]_ ;
  assign \new_[60536]_  = ~A200 & A199;
  assign \new_[60539]_  = A202 & A201;
  assign \new_[60540]_  = \new_[60539]_  & \new_[60536]_ ;
  assign \new_[60541]_  = \new_[60540]_  & \new_[60533]_ ;
  assign \new_[60544]_  = A233 & A232;
  assign \new_[60547]_  = A266 & A265;
  assign \new_[60548]_  = \new_[60547]_  & \new_[60544]_ ;
  assign \new_[60551]_  = ~A299 & A298;
  assign \new_[60554]_  = A302 & A300;
  assign \new_[60555]_  = \new_[60554]_  & \new_[60551]_ ;
  assign \new_[60556]_  = \new_[60555]_  & \new_[60548]_ ;
  assign \new_[60560]_  = ~A166 & ~A167;
  assign \new_[60561]_  = A170 & \new_[60560]_ ;
  assign \new_[60564]_  = ~A200 & A199;
  assign \new_[60567]_  = A202 & A201;
  assign \new_[60568]_  = \new_[60567]_  & \new_[60564]_ ;
  assign \new_[60569]_  = \new_[60568]_  & \new_[60561]_ ;
  assign \new_[60572]_  = A233 & A232;
  assign \new_[60575]_  = ~A266 & ~A265;
  assign \new_[60576]_  = \new_[60575]_  & \new_[60572]_ ;
  assign \new_[60579]_  = ~A299 & A298;
  assign \new_[60582]_  = A301 & A300;
  assign \new_[60583]_  = \new_[60582]_  & \new_[60579]_ ;
  assign \new_[60584]_  = \new_[60583]_  & \new_[60576]_ ;
  assign \new_[60588]_  = ~A166 & ~A167;
  assign \new_[60589]_  = A170 & \new_[60588]_ ;
  assign \new_[60592]_  = ~A200 & A199;
  assign \new_[60595]_  = A202 & A201;
  assign \new_[60596]_  = \new_[60595]_  & \new_[60592]_ ;
  assign \new_[60597]_  = \new_[60596]_  & \new_[60589]_ ;
  assign \new_[60600]_  = A233 & A232;
  assign \new_[60603]_  = ~A266 & ~A265;
  assign \new_[60604]_  = \new_[60603]_  & \new_[60600]_ ;
  assign \new_[60607]_  = ~A299 & A298;
  assign \new_[60610]_  = A302 & A300;
  assign \new_[60611]_  = \new_[60610]_  & \new_[60607]_ ;
  assign \new_[60612]_  = \new_[60611]_  & \new_[60604]_ ;
  assign \new_[60616]_  = ~A166 & ~A167;
  assign \new_[60617]_  = A170 & \new_[60616]_ ;
  assign \new_[60620]_  = ~A200 & A199;
  assign \new_[60623]_  = A202 & A201;
  assign \new_[60624]_  = \new_[60623]_  & \new_[60620]_ ;
  assign \new_[60625]_  = \new_[60624]_  & \new_[60617]_ ;
  assign \new_[60628]_  = ~A235 & ~A233;
  assign \new_[60631]_  = ~A266 & ~A236;
  assign \new_[60632]_  = \new_[60631]_  & \new_[60628]_ ;
  assign \new_[60635]_  = ~A269 & ~A268;
  assign \new_[60638]_  = A299 & ~A298;
  assign \new_[60639]_  = \new_[60638]_  & \new_[60635]_ ;
  assign \new_[60640]_  = \new_[60639]_  & \new_[60632]_ ;
  assign \new_[60644]_  = ~A166 & ~A167;
  assign \new_[60645]_  = A170 & \new_[60644]_ ;
  assign \new_[60648]_  = ~A200 & A199;
  assign \new_[60651]_  = A202 & A201;
  assign \new_[60652]_  = \new_[60651]_  & \new_[60648]_ ;
  assign \new_[60653]_  = \new_[60652]_  & \new_[60645]_ ;
  assign \new_[60656]_  = ~A234 & ~A233;
  assign \new_[60659]_  = A266 & A265;
  assign \new_[60660]_  = \new_[60659]_  & \new_[60656]_ ;
  assign \new_[60663]_  = ~A299 & A298;
  assign \new_[60666]_  = A301 & A300;
  assign \new_[60667]_  = \new_[60666]_  & \new_[60663]_ ;
  assign \new_[60668]_  = \new_[60667]_  & \new_[60660]_ ;
  assign \new_[60672]_  = ~A166 & ~A167;
  assign \new_[60673]_  = A170 & \new_[60672]_ ;
  assign \new_[60676]_  = ~A200 & A199;
  assign \new_[60679]_  = A202 & A201;
  assign \new_[60680]_  = \new_[60679]_  & \new_[60676]_ ;
  assign \new_[60681]_  = \new_[60680]_  & \new_[60673]_ ;
  assign \new_[60684]_  = ~A234 & ~A233;
  assign \new_[60687]_  = A266 & A265;
  assign \new_[60688]_  = \new_[60687]_  & \new_[60684]_ ;
  assign \new_[60691]_  = ~A299 & A298;
  assign \new_[60694]_  = A302 & A300;
  assign \new_[60695]_  = \new_[60694]_  & \new_[60691]_ ;
  assign \new_[60696]_  = \new_[60695]_  & \new_[60688]_ ;
  assign \new_[60700]_  = ~A166 & ~A167;
  assign \new_[60701]_  = A170 & \new_[60700]_ ;
  assign \new_[60704]_  = ~A200 & A199;
  assign \new_[60707]_  = A202 & A201;
  assign \new_[60708]_  = \new_[60707]_  & \new_[60704]_ ;
  assign \new_[60709]_  = \new_[60708]_  & \new_[60701]_ ;
  assign \new_[60712]_  = ~A234 & ~A233;
  assign \new_[60715]_  = ~A267 & ~A266;
  assign \new_[60716]_  = \new_[60715]_  & \new_[60712]_ ;
  assign \new_[60719]_  = ~A299 & A298;
  assign \new_[60722]_  = A301 & A300;
  assign \new_[60723]_  = \new_[60722]_  & \new_[60719]_ ;
  assign \new_[60724]_  = \new_[60723]_  & \new_[60716]_ ;
  assign \new_[60728]_  = ~A166 & ~A167;
  assign \new_[60729]_  = A170 & \new_[60728]_ ;
  assign \new_[60732]_  = ~A200 & A199;
  assign \new_[60735]_  = A202 & A201;
  assign \new_[60736]_  = \new_[60735]_  & \new_[60732]_ ;
  assign \new_[60737]_  = \new_[60736]_  & \new_[60729]_ ;
  assign \new_[60740]_  = ~A234 & ~A233;
  assign \new_[60743]_  = ~A267 & ~A266;
  assign \new_[60744]_  = \new_[60743]_  & \new_[60740]_ ;
  assign \new_[60747]_  = ~A299 & A298;
  assign \new_[60750]_  = A302 & A300;
  assign \new_[60751]_  = \new_[60750]_  & \new_[60747]_ ;
  assign \new_[60752]_  = \new_[60751]_  & \new_[60744]_ ;
  assign \new_[60756]_  = ~A166 & ~A167;
  assign \new_[60757]_  = A170 & \new_[60756]_ ;
  assign \new_[60760]_  = ~A200 & A199;
  assign \new_[60763]_  = A202 & A201;
  assign \new_[60764]_  = \new_[60763]_  & \new_[60760]_ ;
  assign \new_[60765]_  = \new_[60764]_  & \new_[60757]_ ;
  assign \new_[60768]_  = ~A234 & ~A233;
  assign \new_[60771]_  = ~A266 & ~A265;
  assign \new_[60772]_  = \new_[60771]_  & \new_[60768]_ ;
  assign \new_[60775]_  = ~A299 & A298;
  assign \new_[60778]_  = A301 & A300;
  assign \new_[60779]_  = \new_[60778]_  & \new_[60775]_ ;
  assign \new_[60780]_  = \new_[60779]_  & \new_[60772]_ ;
  assign \new_[60784]_  = ~A166 & ~A167;
  assign \new_[60785]_  = A170 & \new_[60784]_ ;
  assign \new_[60788]_  = ~A200 & A199;
  assign \new_[60791]_  = A202 & A201;
  assign \new_[60792]_  = \new_[60791]_  & \new_[60788]_ ;
  assign \new_[60793]_  = \new_[60792]_  & \new_[60785]_ ;
  assign \new_[60796]_  = ~A234 & ~A233;
  assign \new_[60799]_  = ~A266 & ~A265;
  assign \new_[60800]_  = \new_[60799]_  & \new_[60796]_ ;
  assign \new_[60803]_  = ~A299 & A298;
  assign \new_[60806]_  = A302 & A300;
  assign \new_[60807]_  = \new_[60806]_  & \new_[60803]_ ;
  assign \new_[60808]_  = \new_[60807]_  & \new_[60800]_ ;
  assign \new_[60812]_  = ~A166 & ~A167;
  assign \new_[60813]_  = A170 & \new_[60812]_ ;
  assign \new_[60816]_  = ~A200 & A199;
  assign \new_[60819]_  = A202 & A201;
  assign \new_[60820]_  = \new_[60819]_  & \new_[60816]_ ;
  assign \new_[60821]_  = \new_[60820]_  & \new_[60813]_ ;
  assign \new_[60824]_  = ~A233 & A232;
  assign \new_[60827]_  = A235 & A234;
  assign \new_[60828]_  = \new_[60827]_  & \new_[60824]_ ;
  assign \new_[60831]_  = ~A266 & A265;
  assign \new_[60834]_  = A268 & A267;
  assign \new_[60835]_  = \new_[60834]_  & \new_[60831]_ ;
  assign \new_[60836]_  = \new_[60835]_  & \new_[60828]_ ;
  assign \new_[60840]_  = ~A166 & ~A167;
  assign \new_[60841]_  = A170 & \new_[60840]_ ;
  assign \new_[60844]_  = ~A200 & A199;
  assign \new_[60847]_  = A202 & A201;
  assign \new_[60848]_  = \new_[60847]_  & \new_[60844]_ ;
  assign \new_[60849]_  = \new_[60848]_  & \new_[60841]_ ;
  assign \new_[60852]_  = ~A233 & A232;
  assign \new_[60855]_  = A235 & A234;
  assign \new_[60856]_  = \new_[60855]_  & \new_[60852]_ ;
  assign \new_[60859]_  = ~A266 & A265;
  assign \new_[60862]_  = A269 & A267;
  assign \new_[60863]_  = \new_[60862]_  & \new_[60859]_ ;
  assign \new_[60864]_  = \new_[60863]_  & \new_[60856]_ ;
  assign \new_[60868]_  = ~A166 & ~A167;
  assign \new_[60869]_  = A170 & \new_[60868]_ ;
  assign \new_[60872]_  = ~A200 & A199;
  assign \new_[60875]_  = A202 & A201;
  assign \new_[60876]_  = \new_[60875]_  & \new_[60872]_ ;
  assign \new_[60877]_  = \new_[60876]_  & \new_[60869]_ ;
  assign \new_[60880]_  = ~A233 & A232;
  assign \new_[60883]_  = A236 & A234;
  assign \new_[60884]_  = \new_[60883]_  & \new_[60880]_ ;
  assign \new_[60887]_  = ~A266 & A265;
  assign \new_[60890]_  = A268 & A267;
  assign \new_[60891]_  = \new_[60890]_  & \new_[60887]_ ;
  assign \new_[60892]_  = \new_[60891]_  & \new_[60884]_ ;
  assign \new_[60896]_  = ~A166 & ~A167;
  assign \new_[60897]_  = A170 & \new_[60896]_ ;
  assign \new_[60900]_  = ~A200 & A199;
  assign \new_[60903]_  = A202 & A201;
  assign \new_[60904]_  = \new_[60903]_  & \new_[60900]_ ;
  assign \new_[60905]_  = \new_[60904]_  & \new_[60897]_ ;
  assign \new_[60908]_  = ~A233 & A232;
  assign \new_[60911]_  = A236 & A234;
  assign \new_[60912]_  = \new_[60911]_  & \new_[60908]_ ;
  assign \new_[60915]_  = ~A266 & A265;
  assign \new_[60918]_  = A269 & A267;
  assign \new_[60919]_  = \new_[60918]_  & \new_[60915]_ ;
  assign \new_[60920]_  = \new_[60919]_  & \new_[60912]_ ;
  assign \new_[60924]_  = ~A166 & ~A167;
  assign \new_[60925]_  = A170 & \new_[60924]_ ;
  assign \new_[60928]_  = ~A200 & A199;
  assign \new_[60931]_  = A202 & A201;
  assign \new_[60932]_  = \new_[60931]_  & \new_[60928]_ ;
  assign \new_[60933]_  = \new_[60932]_  & \new_[60925]_ ;
  assign \new_[60936]_  = ~A233 & ~A232;
  assign \new_[60939]_  = A266 & A265;
  assign \new_[60940]_  = \new_[60939]_  & \new_[60936]_ ;
  assign \new_[60943]_  = ~A299 & A298;
  assign \new_[60946]_  = A301 & A300;
  assign \new_[60947]_  = \new_[60946]_  & \new_[60943]_ ;
  assign \new_[60948]_  = \new_[60947]_  & \new_[60940]_ ;
  assign \new_[60952]_  = ~A166 & ~A167;
  assign \new_[60953]_  = A170 & \new_[60952]_ ;
  assign \new_[60956]_  = ~A200 & A199;
  assign \new_[60959]_  = A202 & A201;
  assign \new_[60960]_  = \new_[60959]_  & \new_[60956]_ ;
  assign \new_[60961]_  = \new_[60960]_  & \new_[60953]_ ;
  assign \new_[60964]_  = ~A233 & ~A232;
  assign \new_[60967]_  = A266 & A265;
  assign \new_[60968]_  = \new_[60967]_  & \new_[60964]_ ;
  assign \new_[60971]_  = ~A299 & A298;
  assign \new_[60974]_  = A302 & A300;
  assign \new_[60975]_  = \new_[60974]_  & \new_[60971]_ ;
  assign \new_[60976]_  = \new_[60975]_  & \new_[60968]_ ;
  assign \new_[60980]_  = ~A166 & ~A167;
  assign \new_[60981]_  = A170 & \new_[60980]_ ;
  assign \new_[60984]_  = ~A200 & A199;
  assign \new_[60987]_  = A202 & A201;
  assign \new_[60988]_  = \new_[60987]_  & \new_[60984]_ ;
  assign \new_[60989]_  = \new_[60988]_  & \new_[60981]_ ;
  assign \new_[60992]_  = ~A233 & ~A232;
  assign \new_[60995]_  = ~A267 & ~A266;
  assign \new_[60996]_  = \new_[60995]_  & \new_[60992]_ ;
  assign \new_[60999]_  = ~A299 & A298;
  assign \new_[61002]_  = A301 & A300;
  assign \new_[61003]_  = \new_[61002]_  & \new_[60999]_ ;
  assign \new_[61004]_  = \new_[61003]_  & \new_[60996]_ ;
  assign \new_[61008]_  = ~A166 & ~A167;
  assign \new_[61009]_  = A170 & \new_[61008]_ ;
  assign \new_[61012]_  = ~A200 & A199;
  assign \new_[61015]_  = A202 & A201;
  assign \new_[61016]_  = \new_[61015]_  & \new_[61012]_ ;
  assign \new_[61017]_  = \new_[61016]_  & \new_[61009]_ ;
  assign \new_[61020]_  = ~A233 & ~A232;
  assign \new_[61023]_  = ~A267 & ~A266;
  assign \new_[61024]_  = \new_[61023]_  & \new_[61020]_ ;
  assign \new_[61027]_  = ~A299 & A298;
  assign \new_[61030]_  = A302 & A300;
  assign \new_[61031]_  = \new_[61030]_  & \new_[61027]_ ;
  assign \new_[61032]_  = \new_[61031]_  & \new_[61024]_ ;
  assign \new_[61036]_  = ~A166 & ~A167;
  assign \new_[61037]_  = A170 & \new_[61036]_ ;
  assign \new_[61040]_  = ~A200 & A199;
  assign \new_[61043]_  = A202 & A201;
  assign \new_[61044]_  = \new_[61043]_  & \new_[61040]_ ;
  assign \new_[61045]_  = \new_[61044]_  & \new_[61037]_ ;
  assign \new_[61048]_  = ~A233 & ~A232;
  assign \new_[61051]_  = ~A266 & ~A265;
  assign \new_[61052]_  = \new_[61051]_  & \new_[61048]_ ;
  assign \new_[61055]_  = ~A299 & A298;
  assign \new_[61058]_  = A301 & A300;
  assign \new_[61059]_  = \new_[61058]_  & \new_[61055]_ ;
  assign \new_[61060]_  = \new_[61059]_  & \new_[61052]_ ;
  assign \new_[61064]_  = ~A166 & ~A167;
  assign \new_[61065]_  = A170 & \new_[61064]_ ;
  assign \new_[61068]_  = ~A200 & A199;
  assign \new_[61071]_  = A202 & A201;
  assign \new_[61072]_  = \new_[61071]_  & \new_[61068]_ ;
  assign \new_[61073]_  = \new_[61072]_  & \new_[61065]_ ;
  assign \new_[61076]_  = ~A233 & ~A232;
  assign \new_[61079]_  = ~A266 & ~A265;
  assign \new_[61080]_  = \new_[61079]_  & \new_[61076]_ ;
  assign \new_[61083]_  = ~A299 & A298;
  assign \new_[61086]_  = A302 & A300;
  assign \new_[61087]_  = \new_[61086]_  & \new_[61083]_ ;
  assign \new_[61088]_  = \new_[61087]_  & \new_[61080]_ ;
  assign \new_[61092]_  = ~A166 & ~A167;
  assign \new_[61093]_  = A170 & \new_[61092]_ ;
  assign \new_[61096]_  = ~A200 & A199;
  assign \new_[61099]_  = A203 & A201;
  assign \new_[61100]_  = \new_[61099]_  & \new_[61096]_ ;
  assign \new_[61101]_  = \new_[61100]_  & \new_[61093]_ ;
  assign \new_[61104]_  = A233 & A232;
  assign \new_[61107]_  = ~A267 & A265;
  assign \new_[61108]_  = \new_[61107]_  & \new_[61104]_ ;
  assign \new_[61111]_  = ~A299 & A298;
  assign \new_[61114]_  = A301 & A300;
  assign \new_[61115]_  = \new_[61114]_  & \new_[61111]_ ;
  assign \new_[61116]_  = \new_[61115]_  & \new_[61108]_ ;
  assign \new_[61120]_  = ~A166 & ~A167;
  assign \new_[61121]_  = A170 & \new_[61120]_ ;
  assign \new_[61124]_  = ~A200 & A199;
  assign \new_[61127]_  = A203 & A201;
  assign \new_[61128]_  = \new_[61127]_  & \new_[61124]_ ;
  assign \new_[61129]_  = \new_[61128]_  & \new_[61121]_ ;
  assign \new_[61132]_  = A233 & A232;
  assign \new_[61135]_  = ~A267 & A265;
  assign \new_[61136]_  = \new_[61135]_  & \new_[61132]_ ;
  assign \new_[61139]_  = ~A299 & A298;
  assign \new_[61142]_  = A302 & A300;
  assign \new_[61143]_  = \new_[61142]_  & \new_[61139]_ ;
  assign \new_[61144]_  = \new_[61143]_  & \new_[61136]_ ;
  assign \new_[61148]_  = ~A166 & ~A167;
  assign \new_[61149]_  = A170 & \new_[61148]_ ;
  assign \new_[61152]_  = ~A200 & A199;
  assign \new_[61155]_  = A203 & A201;
  assign \new_[61156]_  = \new_[61155]_  & \new_[61152]_ ;
  assign \new_[61157]_  = \new_[61156]_  & \new_[61149]_ ;
  assign \new_[61160]_  = A233 & A232;
  assign \new_[61163]_  = A266 & A265;
  assign \new_[61164]_  = \new_[61163]_  & \new_[61160]_ ;
  assign \new_[61167]_  = ~A299 & A298;
  assign \new_[61170]_  = A301 & A300;
  assign \new_[61171]_  = \new_[61170]_  & \new_[61167]_ ;
  assign \new_[61172]_  = \new_[61171]_  & \new_[61164]_ ;
  assign \new_[61176]_  = ~A166 & ~A167;
  assign \new_[61177]_  = A170 & \new_[61176]_ ;
  assign \new_[61180]_  = ~A200 & A199;
  assign \new_[61183]_  = A203 & A201;
  assign \new_[61184]_  = \new_[61183]_  & \new_[61180]_ ;
  assign \new_[61185]_  = \new_[61184]_  & \new_[61177]_ ;
  assign \new_[61188]_  = A233 & A232;
  assign \new_[61191]_  = A266 & A265;
  assign \new_[61192]_  = \new_[61191]_  & \new_[61188]_ ;
  assign \new_[61195]_  = ~A299 & A298;
  assign \new_[61198]_  = A302 & A300;
  assign \new_[61199]_  = \new_[61198]_  & \new_[61195]_ ;
  assign \new_[61200]_  = \new_[61199]_  & \new_[61192]_ ;
  assign \new_[61204]_  = ~A166 & ~A167;
  assign \new_[61205]_  = A170 & \new_[61204]_ ;
  assign \new_[61208]_  = ~A200 & A199;
  assign \new_[61211]_  = A203 & A201;
  assign \new_[61212]_  = \new_[61211]_  & \new_[61208]_ ;
  assign \new_[61213]_  = \new_[61212]_  & \new_[61205]_ ;
  assign \new_[61216]_  = A233 & A232;
  assign \new_[61219]_  = ~A266 & ~A265;
  assign \new_[61220]_  = \new_[61219]_  & \new_[61216]_ ;
  assign \new_[61223]_  = ~A299 & A298;
  assign \new_[61226]_  = A301 & A300;
  assign \new_[61227]_  = \new_[61226]_  & \new_[61223]_ ;
  assign \new_[61228]_  = \new_[61227]_  & \new_[61220]_ ;
  assign \new_[61232]_  = ~A166 & ~A167;
  assign \new_[61233]_  = A170 & \new_[61232]_ ;
  assign \new_[61236]_  = ~A200 & A199;
  assign \new_[61239]_  = A203 & A201;
  assign \new_[61240]_  = \new_[61239]_  & \new_[61236]_ ;
  assign \new_[61241]_  = \new_[61240]_  & \new_[61233]_ ;
  assign \new_[61244]_  = A233 & A232;
  assign \new_[61247]_  = ~A266 & ~A265;
  assign \new_[61248]_  = \new_[61247]_  & \new_[61244]_ ;
  assign \new_[61251]_  = ~A299 & A298;
  assign \new_[61254]_  = A302 & A300;
  assign \new_[61255]_  = \new_[61254]_  & \new_[61251]_ ;
  assign \new_[61256]_  = \new_[61255]_  & \new_[61248]_ ;
  assign \new_[61260]_  = ~A166 & ~A167;
  assign \new_[61261]_  = A170 & \new_[61260]_ ;
  assign \new_[61264]_  = ~A200 & A199;
  assign \new_[61267]_  = A203 & A201;
  assign \new_[61268]_  = \new_[61267]_  & \new_[61264]_ ;
  assign \new_[61269]_  = \new_[61268]_  & \new_[61261]_ ;
  assign \new_[61272]_  = ~A235 & ~A233;
  assign \new_[61275]_  = ~A266 & ~A236;
  assign \new_[61276]_  = \new_[61275]_  & \new_[61272]_ ;
  assign \new_[61279]_  = ~A269 & ~A268;
  assign \new_[61282]_  = A299 & ~A298;
  assign \new_[61283]_  = \new_[61282]_  & \new_[61279]_ ;
  assign \new_[61284]_  = \new_[61283]_  & \new_[61276]_ ;
  assign \new_[61288]_  = ~A166 & ~A167;
  assign \new_[61289]_  = A170 & \new_[61288]_ ;
  assign \new_[61292]_  = ~A200 & A199;
  assign \new_[61295]_  = A203 & A201;
  assign \new_[61296]_  = \new_[61295]_  & \new_[61292]_ ;
  assign \new_[61297]_  = \new_[61296]_  & \new_[61289]_ ;
  assign \new_[61300]_  = ~A234 & ~A233;
  assign \new_[61303]_  = A266 & A265;
  assign \new_[61304]_  = \new_[61303]_  & \new_[61300]_ ;
  assign \new_[61307]_  = ~A299 & A298;
  assign \new_[61310]_  = A301 & A300;
  assign \new_[61311]_  = \new_[61310]_  & \new_[61307]_ ;
  assign \new_[61312]_  = \new_[61311]_  & \new_[61304]_ ;
  assign \new_[61316]_  = ~A166 & ~A167;
  assign \new_[61317]_  = A170 & \new_[61316]_ ;
  assign \new_[61320]_  = ~A200 & A199;
  assign \new_[61323]_  = A203 & A201;
  assign \new_[61324]_  = \new_[61323]_  & \new_[61320]_ ;
  assign \new_[61325]_  = \new_[61324]_  & \new_[61317]_ ;
  assign \new_[61328]_  = ~A234 & ~A233;
  assign \new_[61331]_  = A266 & A265;
  assign \new_[61332]_  = \new_[61331]_  & \new_[61328]_ ;
  assign \new_[61335]_  = ~A299 & A298;
  assign \new_[61338]_  = A302 & A300;
  assign \new_[61339]_  = \new_[61338]_  & \new_[61335]_ ;
  assign \new_[61340]_  = \new_[61339]_  & \new_[61332]_ ;
  assign \new_[61344]_  = ~A166 & ~A167;
  assign \new_[61345]_  = A170 & \new_[61344]_ ;
  assign \new_[61348]_  = ~A200 & A199;
  assign \new_[61351]_  = A203 & A201;
  assign \new_[61352]_  = \new_[61351]_  & \new_[61348]_ ;
  assign \new_[61353]_  = \new_[61352]_  & \new_[61345]_ ;
  assign \new_[61356]_  = ~A234 & ~A233;
  assign \new_[61359]_  = ~A267 & ~A266;
  assign \new_[61360]_  = \new_[61359]_  & \new_[61356]_ ;
  assign \new_[61363]_  = ~A299 & A298;
  assign \new_[61366]_  = A301 & A300;
  assign \new_[61367]_  = \new_[61366]_  & \new_[61363]_ ;
  assign \new_[61368]_  = \new_[61367]_  & \new_[61360]_ ;
  assign \new_[61372]_  = ~A166 & ~A167;
  assign \new_[61373]_  = A170 & \new_[61372]_ ;
  assign \new_[61376]_  = ~A200 & A199;
  assign \new_[61379]_  = A203 & A201;
  assign \new_[61380]_  = \new_[61379]_  & \new_[61376]_ ;
  assign \new_[61381]_  = \new_[61380]_  & \new_[61373]_ ;
  assign \new_[61384]_  = ~A234 & ~A233;
  assign \new_[61387]_  = ~A267 & ~A266;
  assign \new_[61388]_  = \new_[61387]_  & \new_[61384]_ ;
  assign \new_[61391]_  = ~A299 & A298;
  assign \new_[61394]_  = A302 & A300;
  assign \new_[61395]_  = \new_[61394]_  & \new_[61391]_ ;
  assign \new_[61396]_  = \new_[61395]_  & \new_[61388]_ ;
  assign \new_[61400]_  = ~A166 & ~A167;
  assign \new_[61401]_  = A170 & \new_[61400]_ ;
  assign \new_[61404]_  = ~A200 & A199;
  assign \new_[61407]_  = A203 & A201;
  assign \new_[61408]_  = \new_[61407]_  & \new_[61404]_ ;
  assign \new_[61409]_  = \new_[61408]_  & \new_[61401]_ ;
  assign \new_[61412]_  = ~A234 & ~A233;
  assign \new_[61415]_  = ~A266 & ~A265;
  assign \new_[61416]_  = \new_[61415]_  & \new_[61412]_ ;
  assign \new_[61419]_  = ~A299 & A298;
  assign \new_[61422]_  = A301 & A300;
  assign \new_[61423]_  = \new_[61422]_  & \new_[61419]_ ;
  assign \new_[61424]_  = \new_[61423]_  & \new_[61416]_ ;
  assign \new_[61428]_  = ~A166 & ~A167;
  assign \new_[61429]_  = A170 & \new_[61428]_ ;
  assign \new_[61432]_  = ~A200 & A199;
  assign \new_[61435]_  = A203 & A201;
  assign \new_[61436]_  = \new_[61435]_  & \new_[61432]_ ;
  assign \new_[61437]_  = \new_[61436]_  & \new_[61429]_ ;
  assign \new_[61440]_  = ~A234 & ~A233;
  assign \new_[61443]_  = ~A266 & ~A265;
  assign \new_[61444]_  = \new_[61443]_  & \new_[61440]_ ;
  assign \new_[61447]_  = ~A299 & A298;
  assign \new_[61450]_  = A302 & A300;
  assign \new_[61451]_  = \new_[61450]_  & \new_[61447]_ ;
  assign \new_[61452]_  = \new_[61451]_  & \new_[61444]_ ;
  assign \new_[61456]_  = ~A166 & ~A167;
  assign \new_[61457]_  = A170 & \new_[61456]_ ;
  assign \new_[61460]_  = ~A200 & A199;
  assign \new_[61463]_  = A203 & A201;
  assign \new_[61464]_  = \new_[61463]_  & \new_[61460]_ ;
  assign \new_[61465]_  = \new_[61464]_  & \new_[61457]_ ;
  assign \new_[61468]_  = ~A233 & A232;
  assign \new_[61471]_  = A235 & A234;
  assign \new_[61472]_  = \new_[61471]_  & \new_[61468]_ ;
  assign \new_[61475]_  = ~A266 & A265;
  assign \new_[61478]_  = A268 & A267;
  assign \new_[61479]_  = \new_[61478]_  & \new_[61475]_ ;
  assign \new_[61480]_  = \new_[61479]_  & \new_[61472]_ ;
  assign \new_[61484]_  = ~A166 & ~A167;
  assign \new_[61485]_  = A170 & \new_[61484]_ ;
  assign \new_[61488]_  = ~A200 & A199;
  assign \new_[61491]_  = A203 & A201;
  assign \new_[61492]_  = \new_[61491]_  & \new_[61488]_ ;
  assign \new_[61493]_  = \new_[61492]_  & \new_[61485]_ ;
  assign \new_[61496]_  = ~A233 & A232;
  assign \new_[61499]_  = A235 & A234;
  assign \new_[61500]_  = \new_[61499]_  & \new_[61496]_ ;
  assign \new_[61503]_  = ~A266 & A265;
  assign \new_[61506]_  = A269 & A267;
  assign \new_[61507]_  = \new_[61506]_  & \new_[61503]_ ;
  assign \new_[61508]_  = \new_[61507]_  & \new_[61500]_ ;
  assign \new_[61512]_  = ~A166 & ~A167;
  assign \new_[61513]_  = A170 & \new_[61512]_ ;
  assign \new_[61516]_  = ~A200 & A199;
  assign \new_[61519]_  = A203 & A201;
  assign \new_[61520]_  = \new_[61519]_  & \new_[61516]_ ;
  assign \new_[61521]_  = \new_[61520]_  & \new_[61513]_ ;
  assign \new_[61524]_  = ~A233 & A232;
  assign \new_[61527]_  = A236 & A234;
  assign \new_[61528]_  = \new_[61527]_  & \new_[61524]_ ;
  assign \new_[61531]_  = ~A266 & A265;
  assign \new_[61534]_  = A268 & A267;
  assign \new_[61535]_  = \new_[61534]_  & \new_[61531]_ ;
  assign \new_[61536]_  = \new_[61535]_  & \new_[61528]_ ;
  assign \new_[61540]_  = ~A166 & ~A167;
  assign \new_[61541]_  = A170 & \new_[61540]_ ;
  assign \new_[61544]_  = ~A200 & A199;
  assign \new_[61547]_  = A203 & A201;
  assign \new_[61548]_  = \new_[61547]_  & \new_[61544]_ ;
  assign \new_[61549]_  = \new_[61548]_  & \new_[61541]_ ;
  assign \new_[61552]_  = ~A233 & A232;
  assign \new_[61555]_  = A236 & A234;
  assign \new_[61556]_  = \new_[61555]_  & \new_[61552]_ ;
  assign \new_[61559]_  = ~A266 & A265;
  assign \new_[61562]_  = A269 & A267;
  assign \new_[61563]_  = \new_[61562]_  & \new_[61559]_ ;
  assign \new_[61564]_  = \new_[61563]_  & \new_[61556]_ ;
  assign \new_[61568]_  = ~A166 & ~A167;
  assign \new_[61569]_  = A170 & \new_[61568]_ ;
  assign \new_[61572]_  = ~A200 & A199;
  assign \new_[61575]_  = A203 & A201;
  assign \new_[61576]_  = \new_[61575]_  & \new_[61572]_ ;
  assign \new_[61577]_  = \new_[61576]_  & \new_[61569]_ ;
  assign \new_[61580]_  = ~A233 & ~A232;
  assign \new_[61583]_  = A266 & A265;
  assign \new_[61584]_  = \new_[61583]_  & \new_[61580]_ ;
  assign \new_[61587]_  = ~A299 & A298;
  assign \new_[61590]_  = A301 & A300;
  assign \new_[61591]_  = \new_[61590]_  & \new_[61587]_ ;
  assign \new_[61592]_  = \new_[61591]_  & \new_[61584]_ ;
  assign \new_[61596]_  = ~A166 & ~A167;
  assign \new_[61597]_  = A170 & \new_[61596]_ ;
  assign \new_[61600]_  = ~A200 & A199;
  assign \new_[61603]_  = A203 & A201;
  assign \new_[61604]_  = \new_[61603]_  & \new_[61600]_ ;
  assign \new_[61605]_  = \new_[61604]_  & \new_[61597]_ ;
  assign \new_[61608]_  = ~A233 & ~A232;
  assign \new_[61611]_  = A266 & A265;
  assign \new_[61612]_  = \new_[61611]_  & \new_[61608]_ ;
  assign \new_[61615]_  = ~A299 & A298;
  assign \new_[61618]_  = A302 & A300;
  assign \new_[61619]_  = \new_[61618]_  & \new_[61615]_ ;
  assign \new_[61620]_  = \new_[61619]_  & \new_[61612]_ ;
  assign \new_[61624]_  = ~A166 & ~A167;
  assign \new_[61625]_  = A170 & \new_[61624]_ ;
  assign \new_[61628]_  = ~A200 & A199;
  assign \new_[61631]_  = A203 & A201;
  assign \new_[61632]_  = \new_[61631]_  & \new_[61628]_ ;
  assign \new_[61633]_  = \new_[61632]_  & \new_[61625]_ ;
  assign \new_[61636]_  = ~A233 & ~A232;
  assign \new_[61639]_  = ~A267 & ~A266;
  assign \new_[61640]_  = \new_[61639]_  & \new_[61636]_ ;
  assign \new_[61643]_  = ~A299 & A298;
  assign \new_[61646]_  = A301 & A300;
  assign \new_[61647]_  = \new_[61646]_  & \new_[61643]_ ;
  assign \new_[61648]_  = \new_[61647]_  & \new_[61640]_ ;
  assign \new_[61652]_  = ~A166 & ~A167;
  assign \new_[61653]_  = A170 & \new_[61652]_ ;
  assign \new_[61656]_  = ~A200 & A199;
  assign \new_[61659]_  = A203 & A201;
  assign \new_[61660]_  = \new_[61659]_  & \new_[61656]_ ;
  assign \new_[61661]_  = \new_[61660]_  & \new_[61653]_ ;
  assign \new_[61664]_  = ~A233 & ~A232;
  assign \new_[61667]_  = ~A267 & ~A266;
  assign \new_[61668]_  = \new_[61667]_  & \new_[61664]_ ;
  assign \new_[61671]_  = ~A299 & A298;
  assign \new_[61674]_  = A302 & A300;
  assign \new_[61675]_  = \new_[61674]_  & \new_[61671]_ ;
  assign \new_[61676]_  = \new_[61675]_  & \new_[61668]_ ;
  assign \new_[61680]_  = ~A166 & ~A167;
  assign \new_[61681]_  = A170 & \new_[61680]_ ;
  assign \new_[61684]_  = ~A200 & A199;
  assign \new_[61687]_  = A203 & A201;
  assign \new_[61688]_  = \new_[61687]_  & \new_[61684]_ ;
  assign \new_[61689]_  = \new_[61688]_  & \new_[61681]_ ;
  assign \new_[61692]_  = ~A233 & ~A232;
  assign \new_[61695]_  = ~A266 & ~A265;
  assign \new_[61696]_  = \new_[61695]_  & \new_[61692]_ ;
  assign \new_[61699]_  = ~A299 & A298;
  assign \new_[61702]_  = A301 & A300;
  assign \new_[61703]_  = \new_[61702]_  & \new_[61699]_ ;
  assign \new_[61704]_  = \new_[61703]_  & \new_[61696]_ ;
  assign \new_[61708]_  = ~A166 & ~A167;
  assign \new_[61709]_  = A170 & \new_[61708]_ ;
  assign \new_[61712]_  = ~A200 & A199;
  assign \new_[61715]_  = A203 & A201;
  assign \new_[61716]_  = \new_[61715]_  & \new_[61712]_ ;
  assign \new_[61717]_  = \new_[61716]_  & \new_[61709]_ ;
  assign \new_[61720]_  = ~A233 & ~A232;
  assign \new_[61723]_  = ~A266 & ~A265;
  assign \new_[61724]_  = \new_[61723]_  & \new_[61720]_ ;
  assign \new_[61727]_  = ~A299 & A298;
  assign \new_[61730]_  = A302 & A300;
  assign \new_[61731]_  = \new_[61730]_  & \new_[61727]_ ;
  assign \new_[61732]_  = \new_[61731]_  & \new_[61724]_ ;
  assign \new_[61736]_  = A167 & ~A168;
  assign \new_[61737]_  = A170 & \new_[61736]_ ;
  assign \new_[61740]_  = ~A199 & A166;
  assign \new_[61743]_  = A232 & A200;
  assign \new_[61744]_  = \new_[61743]_  & \new_[61740]_ ;
  assign \new_[61745]_  = \new_[61744]_  & \new_[61737]_ ;
  assign \new_[61748]_  = A265 & A233;
  assign \new_[61751]_  = ~A269 & ~A268;
  assign \new_[61752]_  = \new_[61751]_  & \new_[61748]_ ;
  assign \new_[61755]_  = ~A299 & A298;
  assign \new_[61758]_  = A301 & A300;
  assign \new_[61759]_  = \new_[61758]_  & \new_[61755]_ ;
  assign \new_[61760]_  = \new_[61759]_  & \new_[61752]_ ;
  assign \new_[61764]_  = A167 & ~A168;
  assign \new_[61765]_  = A170 & \new_[61764]_ ;
  assign \new_[61768]_  = ~A199 & A166;
  assign \new_[61771]_  = A232 & A200;
  assign \new_[61772]_  = \new_[61771]_  & \new_[61768]_ ;
  assign \new_[61773]_  = \new_[61772]_  & \new_[61765]_ ;
  assign \new_[61776]_  = A265 & A233;
  assign \new_[61779]_  = ~A269 & ~A268;
  assign \new_[61780]_  = \new_[61779]_  & \new_[61776]_ ;
  assign \new_[61783]_  = ~A299 & A298;
  assign \new_[61786]_  = A302 & A300;
  assign \new_[61787]_  = \new_[61786]_  & \new_[61783]_ ;
  assign \new_[61788]_  = \new_[61787]_  & \new_[61780]_ ;
  assign \new_[61792]_  = A167 & ~A168;
  assign \new_[61793]_  = A170 & \new_[61792]_ ;
  assign \new_[61796]_  = ~A199 & A166;
  assign \new_[61799]_  = ~A233 & A200;
  assign \new_[61800]_  = \new_[61799]_  & \new_[61796]_ ;
  assign \new_[61801]_  = \new_[61800]_  & \new_[61793]_ ;
  assign \new_[61804]_  = ~A236 & ~A235;
  assign \new_[61807]_  = A266 & A265;
  assign \new_[61808]_  = \new_[61807]_  & \new_[61804]_ ;
  assign \new_[61811]_  = ~A299 & A298;
  assign \new_[61814]_  = A301 & A300;
  assign \new_[61815]_  = \new_[61814]_  & \new_[61811]_ ;
  assign \new_[61816]_  = \new_[61815]_  & \new_[61808]_ ;
  assign \new_[61820]_  = A167 & ~A168;
  assign \new_[61821]_  = A170 & \new_[61820]_ ;
  assign \new_[61824]_  = ~A199 & A166;
  assign \new_[61827]_  = ~A233 & A200;
  assign \new_[61828]_  = \new_[61827]_  & \new_[61824]_ ;
  assign \new_[61829]_  = \new_[61828]_  & \new_[61821]_ ;
  assign \new_[61832]_  = ~A236 & ~A235;
  assign \new_[61835]_  = A266 & A265;
  assign \new_[61836]_  = \new_[61835]_  & \new_[61832]_ ;
  assign \new_[61839]_  = ~A299 & A298;
  assign \new_[61842]_  = A302 & A300;
  assign \new_[61843]_  = \new_[61842]_  & \new_[61839]_ ;
  assign \new_[61844]_  = \new_[61843]_  & \new_[61836]_ ;
  assign \new_[61848]_  = A167 & ~A168;
  assign \new_[61849]_  = A170 & \new_[61848]_ ;
  assign \new_[61852]_  = ~A199 & A166;
  assign \new_[61855]_  = ~A233 & A200;
  assign \new_[61856]_  = \new_[61855]_  & \new_[61852]_ ;
  assign \new_[61857]_  = \new_[61856]_  & \new_[61849]_ ;
  assign \new_[61860]_  = ~A236 & ~A235;
  assign \new_[61863]_  = ~A267 & ~A266;
  assign \new_[61864]_  = \new_[61863]_  & \new_[61860]_ ;
  assign \new_[61867]_  = ~A299 & A298;
  assign \new_[61870]_  = A301 & A300;
  assign \new_[61871]_  = \new_[61870]_  & \new_[61867]_ ;
  assign \new_[61872]_  = \new_[61871]_  & \new_[61864]_ ;
  assign \new_[61876]_  = A167 & ~A168;
  assign \new_[61877]_  = A170 & \new_[61876]_ ;
  assign \new_[61880]_  = ~A199 & A166;
  assign \new_[61883]_  = ~A233 & A200;
  assign \new_[61884]_  = \new_[61883]_  & \new_[61880]_ ;
  assign \new_[61885]_  = \new_[61884]_  & \new_[61877]_ ;
  assign \new_[61888]_  = ~A236 & ~A235;
  assign \new_[61891]_  = ~A267 & ~A266;
  assign \new_[61892]_  = \new_[61891]_  & \new_[61888]_ ;
  assign \new_[61895]_  = ~A299 & A298;
  assign \new_[61898]_  = A302 & A300;
  assign \new_[61899]_  = \new_[61898]_  & \new_[61895]_ ;
  assign \new_[61900]_  = \new_[61899]_  & \new_[61892]_ ;
  assign \new_[61904]_  = A167 & ~A168;
  assign \new_[61905]_  = A170 & \new_[61904]_ ;
  assign \new_[61908]_  = ~A199 & A166;
  assign \new_[61911]_  = ~A233 & A200;
  assign \new_[61912]_  = \new_[61911]_  & \new_[61908]_ ;
  assign \new_[61913]_  = \new_[61912]_  & \new_[61905]_ ;
  assign \new_[61916]_  = ~A236 & ~A235;
  assign \new_[61919]_  = ~A266 & ~A265;
  assign \new_[61920]_  = \new_[61919]_  & \new_[61916]_ ;
  assign \new_[61923]_  = ~A299 & A298;
  assign \new_[61926]_  = A301 & A300;
  assign \new_[61927]_  = \new_[61926]_  & \new_[61923]_ ;
  assign \new_[61928]_  = \new_[61927]_  & \new_[61920]_ ;
  assign \new_[61932]_  = A167 & ~A168;
  assign \new_[61933]_  = A170 & \new_[61932]_ ;
  assign \new_[61936]_  = ~A199 & A166;
  assign \new_[61939]_  = ~A233 & A200;
  assign \new_[61940]_  = \new_[61939]_  & \new_[61936]_ ;
  assign \new_[61941]_  = \new_[61940]_  & \new_[61933]_ ;
  assign \new_[61944]_  = ~A236 & ~A235;
  assign \new_[61947]_  = ~A266 & ~A265;
  assign \new_[61948]_  = \new_[61947]_  & \new_[61944]_ ;
  assign \new_[61951]_  = ~A299 & A298;
  assign \new_[61954]_  = A302 & A300;
  assign \new_[61955]_  = \new_[61954]_  & \new_[61951]_ ;
  assign \new_[61956]_  = \new_[61955]_  & \new_[61948]_ ;
  assign \new_[61960]_  = A167 & ~A168;
  assign \new_[61961]_  = A170 & \new_[61960]_ ;
  assign \new_[61964]_  = ~A199 & A166;
  assign \new_[61967]_  = ~A233 & A200;
  assign \new_[61968]_  = \new_[61967]_  & \new_[61964]_ ;
  assign \new_[61969]_  = \new_[61968]_  & \new_[61961]_ ;
  assign \new_[61972]_  = ~A266 & ~A234;
  assign \new_[61975]_  = ~A269 & ~A268;
  assign \new_[61976]_  = \new_[61975]_  & \new_[61972]_ ;
  assign \new_[61979]_  = ~A299 & A298;
  assign \new_[61982]_  = A301 & A300;
  assign \new_[61983]_  = \new_[61982]_  & \new_[61979]_ ;
  assign \new_[61984]_  = \new_[61983]_  & \new_[61976]_ ;
  assign \new_[61988]_  = A167 & ~A168;
  assign \new_[61989]_  = A170 & \new_[61988]_ ;
  assign \new_[61992]_  = ~A199 & A166;
  assign \new_[61995]_  = ~A233 & A200;
  assign \new_[61996]_  = \new_[61995]_  & \new_[61992]_ ;
  assign \new_[61997]_  = \new_[61996]_  & \new_[61989]_ ;
  assign \new_[62000]_  = ~A266 & ~A234;
  assign \new_[62003]_  = ~A269 & ~A268;
  assign \new_[62004]_  = \new_[62003]_  & \new_[62000]_ ;
  assign \new_[62007]_  = ~A299 & A298;
  assign \new_[62010]_  = A302 & A300;
  assign \new_[62011]_  = \new_[62010]_  & \new_[62007]_ ;
  assign \new_[62012]_  = \new_[62011]_  & \new_[62004]_ ;
  assign \new_[62016]_  = A167 & ~A168;
  assign \new_[62017]_  = A170 & \new_[62016]_ ;
  assign \new_[62020]_  = ~A199 & A166;
  assign \new_[62023]_  = ~A232 & A200;
  assign \new_[62024]_  = \new_[62023]_  & \new_[62020]_ ;
  assign \new_[62025]_  = \new_[62024]_  & \new_[62017]_ ;
  assign \new_[62028]_  = ~A266 & ~A233;
  assign \new_[62031]_  = ~A269 & ~A268;
  assign \new_[62032]_  = \new_[62031]_  & \new_[62028]_ ;
  assign \new_[62035]_  = ~A299 & A298;
  assign \new_[62038]_  = A301 & A300;
  assign \new_[62039]_  = \new_[62038]_  & \new_[62035]_ ;
  assign \new_[62040]_  = \new_[62039]_  & \new_[62032]_ ;
  assign \new_[62044]_  = A167 & ~A168;
  assign \new_[62045]_  = A170 & \new_[62044]_ ;
  assign \new_[62048]_  = ~A199 & A166;
  assign \new_[62051]_  = ~A232 & A200;
  assign \new_[62052]_  = \new_[62051]_  & \new_[62048]_ ;
  assign \new_[62053]_  = \new_[62052]_  & \new_[62045]_ ;
  assign \new_[62056]_  = ~A266 & ~A233;
  assign \new_[62059]_  = ~A269 & ~A268;
  assign \new_[62060]_  = \new_[62059]_  & \new_[62056]_ ;
  assign \new_[62063]_  = ~A299 & A298;
  assign \new_[62066]_  = A302 & A300;
  assign \new_[62067]_  = \new_[62066]_  & \new_[62063]_ ;
  assign \new_[62068]_  = \new_[62067]_  & \new_[62060]_ ;
  assign \new_[62072]_  = A167 & ~A168;
  assign \new_[62073]_  = ~A170 & \new_[62072]_ ;
  assign \new_[62076]_  = ~A199 & ~A166;
  assign \new_[62079]_  = A232 & A200;
  assign \new_[62080]_  = \new_[62079]_  & \new_[62076]_ ;
  assign \new_[62081]_  = \new_[62080]_  & \new_[62073]_ ;
  assign \new_[62084]_  = A265 & A233;
  assign \new_[62087]_  = ~A269 & ~A268;
  assign \new_[62088]_  = \new_[62087]_  & \new_[62084]_ ;
  assign \new_[62091]_  = ~A299 & A298;
  assign \new_[62094]_  = A301 & A300;
  assign \new_[62095]_  = \new_[62094]_  & \new_[62091]_ ;
  assign \new_[62096]_  = \new_[62095]_  & \new_[62088]_ ;
  assign \new_[62100]_  = A167 & ~A168;
  assign \new_[62101]_  = ~A170 & \new_[62100]_ ;
  assign \new_[62104]_  = ~A199 & ~A166;
  assign \new_[62107]_  = A232 & A200;
  assign \new_[62108]_  = \new_[62107]_  & \new_[62104]_ ;
  assign \new_[62109]_  = \new_[62108]_  & \new_[62101]_ ;
  assign \new_[62112]_  = A265 & A233;
  assign \new_[62115]_  = ~A269 & ~A268;
  assign \new_[62116]_  = \new_[62115]_  & \new_[62112]_ ;
  assign \new_[62119]_  = ~A299 & A298;
  assign \new_[62122]_  = A302 & A300;
  assign \new_[62123]_  = \new_[62122]_  & \new_[62119]_ ;
  assign \new_[62124]_  = \new_[62123]_  & \new_[62116]_ ;
  assign \new_[62128]_  = A167 & ~A168;
  assign \new_[62129]_  = ~A170 & \new_[62128]_ ;
  assign \new_[62132]_  = ~A199 & ~A166;
  assign \new_[62135]_  = ~A233 & A200;
  assign \new_[62136]_  = \new_[62135]_  & \new_[62132]_ ;
  assign \new_[62137]_  = \new_[62136]_  & \new_[62129]_ ;
  assign \new_[62140]_  = ~A236 & ~A235;
  assign \new_[62143]_  = A266 & A265;
  assign \new_[62144]_  = \new_[62143]_  & \new_[62140]_ ;
  assign \new_[62147]_  = ~A299 & A298;
  assign \new_[62150]_  = A301 & A300;
  assign \new_[62151]_  = \new_[62150]_  & \new_[62147]_ ;
  assign \new_[62152]_  = \new_[62151]_  & \new_[62144]_ ;
  assign \new_[62156]_  = A167 & ~A168;
  assign \new_[62157]_  = ~A170 & \new_[62156]_ ;
  assign \new_[62160]_  = ~A199 & ~A166;
  assign \new_[62163]_  = ~A233 & A200;
  assign \new_[62164]_  = \new_[62163]_  & \new_[62160]_ ;
  assign \new_[62165]_  = \new_[62164]_  & \new_[62157]_ ;
  assign \new_[62168]_  = ~A236 & ~A235;
  assign \new_[62171]_  = A266 & A265;
  assign \new_[62172]_  = \new_[62171]_  & \new_[62168]_ ;
  assign \new_[62175]_  = ~A299 & A298;
  assign \new_[62178]_  = A302 & A300;
  assign \new_[62179]_  = \new_[62178]_  & \new_[62175]_ ;
  assign \new_[62180]_  = \new_[62179]_  & \new_[62172]_ ;
  assign \new_[62184]_  = A167 & ~A168;
  assign \new_[62185]_  = ~A170 & \new_[62184]_ ;
  assign \new_[62188]_  = ~A199 & ~A166;
  assign \new_[62191]_  = ~A233 & A200;
  assign \new_[62192]_  = \new_[62191]_  & \new_[62188]_ ;
  assign \new_[62193]_  = \new_[62192]_  & \new_[62185]_ ;
  assign \new_[62196]_  = ~A236 & ~A235;
  assign \new_[62199]_  = ~A267 & ~A266;
  assign \new_[62200]_  = \new_[62199]_  & \new_[62196]_ ;
  assign \new_[62203]_  = ~A299 & A298;
  assign \new_[62206]_  = A301 & A300;
  assign \new_[62207]_  = \new_[62206]_  & \new_[62203]_ ;
  assign \new_[62208]_  = \new_[62207]_  & \new_[62200]_ ;
  assign \new_[62212]_  = A167 & ~A168;
  assign \new_[62213]_  = ~A170 & \new_[62212]_ ;
  assign \new_[62216]_  = ~A199 & ~A166;
  assign \new_[62219]_  = ~A233 & A200;
  assign \new_[62220]_  = \new_[62219]_  & \new_[62216]_ ;
  assign \new_[62221]_  = \new_[62220]_  & \new_[62213]_ ;
  assign \new_[62224]_  = ~A236 & ~A235;
  assign \new_[62227]_  = ~A267 & ~A266;
  assign \new_[62228]_  = \new_[62227]_  & \new_[62224]_ ;
  assign \new_[62231]_  = ~A299 & A298;
  assign \new_[62234]_  = A302 & A300;
  assign \new_[62235]_  = \new_[62234]_  & \new_[62231]_ ;
  assign \new_[62236]_  = \new_[62235]_  & \new_[62228]_ ;
  assign \new_[62240]_  = A167 & ~A168;
  assign \new_[62241]_  = ~A170 & \new_[62240]_ ;
  assign \new_[62244]_  = ~A199 & ~A166;
  assign \new_[62247]_  = ~A233 & A200;
  assign \new_[62248]_  = \new_[62247]_  & \new_[62244]_ ;
  assign \new_[62249]_  = \new_[62248]_  & \new_[62241]_ ;
  assign \new_[62252]_  = ~A236 & ~A235;
  assign \new_[62255]_  = ~A266 & ~A265;
  assign \new_[62256]_  = \new_[62255]_  & \new_[62252]_ ;
  assign \new_[62259]_  = ~A299 & A298;
  assign \new_[62262]_  = A301 & A300;
  assign \new_[62263]_  = \new_[62262]_  & \new_[62259]_ ;
  assign \new_[62264]_  = \new_[62263]_  & \new_[62256]_ ;
  assign \new_[62268]_  = A167 & ~A168;
  assign \new_[62269]_  = ~A170 & \new_[62268]_ ;
  assign \new_[62272]_  = ~A199 & ~A166;
  assign \new_[62275]_  = ~A233 & A200;
  assign \new_[62276]_  = \new_[62275]_  & \new_[62272]_ ;
  assign \new_[62277]_  = \new_[62276]_  & \new_[62269]_ ;
  assign \new_[62280]_  = ~A236 & ~A235;
  assign \new_[62283]_  = ~A266 & ~A265;
  assign \new_[62284]_  = \new_[62283]_  & \new_[62280]_ ;
  assign \new_[62287]_  = ~A299 & A298;
  assign \new_[62290]_  = A302 & A300;
  assign \new_[62291]_  = \new_[62290]_  & \new_[62287]_ ;
  assign \new_[62292]_  = \new_[62291]_  & \new_[62284]_ ;
  assign \new_[62296]_  = A167 & ~A168;
  assign \new_[62297]_  = ~A170 & \new_[62296]_ ;
  assign \new_[62300]_  = ~A199 & ~A166;
  assign \new_[62303]_  = ~A233 & A200;
  assign \new_[62304]_  = \new_[62303]_  & \new_[62300]_ ;
  assign \new_[62305]_  = \new_[62304]_  & \new_[62297]_ ;
  assign \new_[62308]_  = ~A266 & ~A234;
  assign \new_[62311]_  = ~A269 & ~A268;
  assign \new_[62312]_  = \new_[62311]_  & \new_[62308]_ ;
  assign \new_[62315]_  = ~A299 & A298;
  assign \new_[62318]_  = A301 & A300;
  assign \new_[62319]_  = \new_[62318]_  & \new_[62315]_ ;
  assign \new_[62320]_  = \new_[62319]_  & \new_[62312]_ ;
  assign \new_[62324]_  = A167 & ~A168;
  assign \new_[62325]_  = ~A170 & \new_[62324]_ ;
  assign \new_[62328]_  = ~A199 & ~A166;
  assign \new_[62331]_  = ~A233 & A200;
  assign \new_[62332]_  = \new_[62331]_  & \new_[62328]_ ;
  assign \new_[62333]_  = \new_[62332]_  & \new_[62325]_ ;
  assign \new_[62336]_  = ~A266 & ~A234;
  assign \new_[62339]_  = ~A269 & ~A268;
  assign \new_[62340]_  = \new_[62339]_  & \new_[62336]_ ;
  assign \new_[62343]_  = ~A299 & A298;
  assign \new_[62346]_  = A302 & A300;
  assign \new_[62347]_  = \new_[62346]_  & \new_[62343]_ ;
  assign \new_[62348]_  = \new_[62347]_  & \new_[62340]_ ;
  assign \new_[62352]_  = A167 & ~A168;
  assign \new_[62353]_  = ~A170 & \new_[62352]_ ;
  assign \new_[62356]_  = ~A199 & ~A166;
  assign \new_[62359]_  = ~A232 & A200;
  assign \new_[62360]_  = \new_[62359]_  & \new_[62356]_ ;
  assign \new_[62361]_  = \new_[62360]_  & \new_[62353]_ ;
  assign \new_[62364]_  = ~A266 & ~A233;
  assign \new_[62367]_  = ~A269 & ~A268;
  assign \new_[62368]_  = \new_[62367]_  & \new_[62364]_ ;
  assign \new_[62371]_  = ~A299 & A298;
  assign \new_[62374]_  = A301 & A300;
  assign \new_[62375]_  = \new_[62374]_  & \new_[62371]_ ;
  assign \new_[62376]_  = \new_[62375]_  & \new_[62368]_ ;
  assign \new_[62380]_  = A167 & ~A168;
  assign \new_[62381]_  = ~A170 & \new_[62380]_ ;
  assign \new_[62384]_  = ~A199 & ~A166;
  assign \new_[62387]_  = ~A232 & A200;
  assign \new_[62388]_  = \new_[62387]_  & \new_[62384]_ ;
  assign \new_[62389]_  = \new_[62388]_  & \new_[62381]_ ;
  assign \new_[62392]_  = ~A266 & ~A233;
  assign \new_[62395]_  = ~A269 & ~A268;
  assign \new_[62396]_  = \new_[62395]_  & \new_[62392]_ ;
  assign \new_[62399]_  = ~A299 & A298;
  assign \new_[62402]_  = A302 & A300;
  assign \new_[62403]_  = \new_[62402]_  & \new_[62399]_ ;
  assign \new_[62404]_  = \new_[62403]_  & \new_[62396]_ ;
  assign \new_[62408]_  = ~A167 & ~A168;
  assign \new_[62409]_  = ~A170 & \new_[62408]_ ;
  assign \new_[62412]_  = ~A199 & A166;
  assign \new_[62415]_  = A232 & A200;
  assign \new_[62416]_  = \new_[62415]_  & \new_[62412]_ ;
  assign \new_[62417]_  = \new_[62416]_  & \new_[62409]_ ;
  assign \new_[62420]_  = A265 & A233;
  assign \new_[62423]_  = ~A269 & ~A268;
  assign \new_[62424]_  = \new_[62423]_  & \new_[62420]_ ;
  assign \new_[62427]_  = ~A299 & A298;
  assign \new_[62430]_  = A301 & A300;
  assign \new_[62431]_  = \new_[62430]_  & \new_[62427]_ ;
  assign \new_[62432]_  = \new_[62431]_  & \new_[62424]_ ;
  assign \new_[62436]_  = ~A167 & ~A168;
  assign \new_[62437]_  = ~A170 & \new_[62436]_ ;
  assign \new_[62440]_  = ~A199 & A166;
  assign \new_[62443]_  = A232 & A200;
  assign \new_[62444]_  = \new_[62443]_  & \new_[62440]_ ;
  assign \new_[62445]_  = \new_[62444]_  & \new_[62437]_ ;
  assign \new_[62448]_  = A265 & A233;
  assign \new_[62451]_  = ~A269 & ~A268;
  assign \new_[62452]_  = \new_[62451]_  & \new_[62448]_ ;
  assign \new_[62455]_  = ~A299 & A298;
  assign \new_[62458]_  = A302 & A300;
  assign \new_[62459]_  = \new_[62458]_  & \new_[62455]_ ;
  assign \new_[62460]_  = \new_[62459]_  & \new_[62452]_ ;
  assign \new_[62464]_  = ~A167 & ~A168;
  assign \new_[62465]_  = ~A170 & \new_[62464]_ ;
  assign \new_[62468]_  = ~A199 & A166;
  assign \new_[62471]_  = ~A233 & A200;
  assign \new_[62472]_  = \new_[62471]_  & \new_[62468]_ ;
  assign \new_[62473]_  = \new_[62472]_  & \new_[62465]_ ;
  assign \new_[62476]_  = ~A236 & ~A235;
  assign \new_[62479]_  = A266 & A265;
  assign \new_[62480]_  = \new_[62479]_  & \new_[62476]_ ;
  assign \new_[62483]_  = ~A299 & A298;
  assign \new_[62486]_  = A301 & A300;
  assign \new_[62487]_  = \new_[62486]_  & \new_[62483]_ ;
  assign \new_[62488]_  = \new_[62487]_  & \new_[62480]_ ;
  assign \new_[62492]_  = ~A167 & ~A168;
  assign \new_[62493]_  = ~A170 & \new_[62492]_ ;
  assign \new_[62496]_  = ~A199 & A166;
  assign \new_[62499]_  = ~A233 & A200;
  assign \new_[62500]_  = \new_[62499]_  & \new_[62496]_ ;
  assign \new_[62501]_  = \new_[62500]_  & \new_[62493]_ ;
  assign \new_[62504]_  = ~A236 & ~A235;
  assign \new_[62507]_  = A266 & A265;
  assign \new_[62508]_  = \new_[62507]_  & \new_[62504]_ ;
  assign \new_[62511]_  = ~A299 & A298;
  assign \new_[62514]_  = A302 & A300;
  assign \new_[62515]_  = \new_[62514]_  & \new_[62511]_ ;
  assign \new_[62516]_  = \new_[62515]_  & \new_[62508]_ ;
  assign \new_[62520]_  = ~A167 & ~A168;
  assign \new_[62521]_  = ~A170 & \new_[62520]_ ;
  assign \new_[62524]_  = ~A199 & A166;
  assign \new_[62527]_  = ~A233 & A200;
  assign \new_[62528]_  = \new_[62527]_  & \new_[62524]_ ;
  assign \new_[62529]_  = \new_[62528]_  & \new_[62521]_ ;
  assign \new_[62532]_  = ~A236 & ~A235;
  assign \new_[62535]_  = ~A267 & ~A266;
  assign \new_[62536]_  = \new_[62535]_  & \new_[62532]_ ;
  assign \new_[62539]_  = ~A299 & A298;
  assign \new_[62542]_  = A301 & A300;
  assign \new_[62543]_  = \new_[62542]_  & \new_[62539]_ ;
  assign \new_[62544]_  = \new_[62543]_  & \new_[62536]_ ;
  assign \new_[62548]_  = ~A167 & ~A168;
  assign \new_[62549]_  = ~A170 & \new_[62548]_ ;
  assign \new_[62552]_  = ~A199 & A166;
  assign \new_[62555]_  = ~A233 & A200;
  assign \new_[62556]_  = \new_[62555]_  & \new_[62552]_ ;
  assign \new_[62557]_  = \new_[62556]_  & \new_[62549]_ ;
  assign \new_[62560]_  = ~A236 & ~A235;
  assign \new_[62563]_  = ~A267 & ~A266;
  assign \new_[62564]_  = \new_[62563]_  & \new_[62560]_ ;
  assign \new_[62567]_  = ~A299 & A298;
  assign \new_[62570]_  = A302 & A300;
  assign \new_[62571]_  = \new_[62570]_  & \new_[62567]_ ;
  assign \new_[62572]_  = \new_[62571]_  & \new_[62564]_ ;
  assign \new_[62576]_  = ~A167 & ~A168;
  assign \new_[62577]_  = ~A170 & \new_[62576]_ ;
  assign \new_[62580]_  = ~A199 & A166;
  assign \new_[62583]_  = ~A233 & A200;
  assign \new_[62584]_  = \new_[62583]_  & \new_[62580]_ ;
  assign \new_[62585]_  = \new_[62584]_  & \new_[62577]_ ;
  assign \new_[62588]_  = ~A236 & ~A235;
  assign \new_[62591]_  = ~A266 & ~A265;
  assign \new_[62592]_  = \new_[62591]_  & \new_[62588]_ ;
  assign \new_[62595]_  = ~A299 & A298;
  assign \new_[62598]_  = A301 & A300;
  assign \new_[62599]_  = \new_[62598]_  & \new_[62595]_ ;
  assign \new_[62600]_  = \new_[62599]_  & \new_[62592]_ ;
  assign \new_[62604]_  = ~A167 & ~A168;
  assign \new_[62605]_  = ~A170 & \new_[62604]_ ;
  assign \new_[62608]_  = ~A199 & A166;
  assign \new_[62611]_  = ~A233 & A200;
  assign \new_[62612]_  = \new_[62611]_  & \new_[62608]_ ;
  assign \new_[62613]_  = \new_[62612]_  & \new_[62605]_ ;
  assign \new_[62616]_  = ~A236 & ~A235;
  assign \new_[62619]_  = ~A266 & ~A265;
  assign \new_[62620]_  = \new_[62619]_  & \new_[62616]_ ;
  assign \new_[62623]_  = ~A299 & A298;
  assign \new_[62626]_  = A302 & A300;
  assign \new_[62627]_  = \new_[62626]_  & \new_[62623]_ ;
  assign \new_[62628]_  = \new_[62627]_  & \new_[62620]_ ;
  assign \new_[62632]_  = ~A167 & ~A168;
  assign \new_[62633]_  = ~A170 & \new_[62632]_ ;
  assign \new_[62636]_  = ~A199 & A166;
  assign \new_[62639]_  = ~A233 & A200;
  assign \new_[62640]_  = \new_[62639]_  & \new_[62636]_ ;
  assign \new_[62641]_  = \new_[62640]_  & \new_[62633]_ ;
  assign \new_[62644]_  = ~A266 & ~A234;
  assign \new_[62647]_  = ~A269 & ~A268;
  assign \new_[62648]_  = \new_[62647]_  & \new_[62644]_ ;
  assign \new_[62651]_  = ~A299 & A298;
  assign \new_[62654]_  = A301 & A300;
  assign \new_[62655]_  = \new_[62654]_  & \new_[62651]_ ;
  assign \new_[62656]_  = \new_[62655]_  & \new_[62648]_ ;
  assign \new_[62660]_  = ~A167 & ~A168;
  assign \new_[62661]_  = ~A170 & \new_[62660]_ ;
  assign \new_[62664]_  = ~A199 & A166;
  assign \new_[62667]_  = ~A233 & A200;
  assign \new_[62668]_  = \new_[62667]_  & \new_[62664]_ ;
  assign \new_[62669]_  = \new_[62668]_  & \new_[62661]_ ;
  assign \new_[62672]_  = ~A266 & ~A234;
  assign \new_[62675]_  = ~A269 & ~A268;
  assign \new_[62676]_  = \new_[62675]_  & \new_[62672]_ ;
  assign \new_[62679]_  = ~A299 & A298;
  assign \new_[62682]_  = A302 & A300;
  assign \new_[62683]_  = \new_[62682]_  & \new_[62679]_ ;
  assign \new_[62684]_  = \new_[62683]_  & \new_[62676]_ ;
  assign \new_[62688]_  = ~A167 & ~A168;
  assign \new_[62689]_  = ~A170 & \new_[62688]_ ;
  assign \new_[62692]_  = ~A199 & A166;
  assign \new_[62695]_  = ~A232 & A200;
  assign \new_[62696]_  = \new_[62695]_  & \new_[62692]_ ;
  assign \new_[62697]_  = \new_[62696]_  & \new_[62689]_ ;
  assign \new_[62700]_  = ~A266 & ~A233;
  assign \new_[62703]_  = ~A269 & ~A268;
  assign \new_[62704]_  = \new_[62703]_  & \new_[62700]_ ;
  assign \new_[62707]_  = ~A299 & A298;
  assign \new_[62710]_  = A301 & A300;
  assign \new_[62711]_  = \new_[62710]_  & \new_[62707]_ ;
  assign \new_[62712]_  = \new_[62711]_  & \new_[62704]_ ;
  assign \new_[62716]_  = ~A167 & ~A168;
  assign \new_[62717]_  = ~A170 & \new_[62716]_ ;
  assign \new_[62720]_  = ~A199 & A166;
  assign \new_[62723]_  = ~A232 & A200;
  assign \new_[62724]_  = \new_[62723]_  & \new_[62720]_ ;
  assign \new_[62725]_  = \new_[62724]_  & \new_[62717]_ ;
  assign \new_[62728]_  = ~A266 & ~A233;
  assign \new_[62731]_  = ~A269 & ~A268;
  assign \new_[62732]_  = \new_[62731]_  & \new_[62728]_ ;
  assign \new_[62735]_  = ~A299 & A298;
  assign \new_[62738]_  = A302 & A300;
  assign \new_[62739]_  = \new_[62738]_  & \new_[62735]_ ;
  assign \new_[62740]_  = \new_[62739]_  & \new_[62732]_ ;
  assign \new_[62744]_  = A167 & ~A168;
  assign \new_[62745]_  = A169 & \new_[62744]_ ;
  assign \new_[62748]_  = ~A199 & ~A166;
  assign \new_[62751]_  = A232 & A200;
  assign \new_[62752]_  = \new_[62751]_  & \new_[62748]_ ;
  assign \new_[62753]_  = \new_[62752]_  & \new_[62745]_ ;
  assign \new_[62756]_  = A265 & A233;
  assign \new_[62759]_  = ~A269 & ~A268;
  assign \new_[62760]_  = \new_[62759]_  & \new_[62756]_ ;
  assign \new_[62763]_  = ~A299 & A298;
  assign \new_[62766]_  = A301 & A300;
  assign \new_[62767]_  = \new_[62766]_  & \new_[62763]_ ;
  assign \new_[62768]_  = \new_[62767]_  & \new_[62760]_ ;
  assign \new_[62772]_  = A167 & ~A168;
  assign \new_[62773]_  = A169 & \new_[62772]_ ;
  assign \new_[62776]_  = ~A199 & ~A166;
  assign \new_[62779]_  = A232 & A200;
  assign \new_[62780]_  = \new_[62779]_  & \new_[62776]_ ;
  assign \new_[62781]_  = \new_[62780]_  & \new_[62773]_ ;
  assign \new_[62784]_  = A265 & A233;
  assign \new_[62787]_  = ~A269 & ~A268;
  assign \new_[62788]_  = \new_[62787]_  & \new_[62784]_ ;
  assign \new_[62791]_  = ~A299 & A298;
  assign \new_[62794]_  = A302 & A300;
  assign \new_[62795]_  = \new_[62794]_  & \new_[62791]_ ;
  assign \new_[62796]_  = \new_[62795]_  & \new_[62788]_ ;
  assign \new_[62800]_  = A167 & ~A168;
  assign \new_[62801]_  = A169 & \new_[62800]_ ;
  assign \new_[62804]_  = ~A199 & ~A166;
  assign \new_[62807]_  = ~A233 & A200;
  assign \new_[62808]_  = \new_[62807]_  & \new_[62804]_ ;
  assign \new_[62809]_  = \new_[62808]_  & \new_[62801]_ ;
  assign \new_[62812]_  = ~A236 & ~A235;
  assign \new_[62815]_  = A266 & A265;
  assign \new_[62816]_  = \new_[62815]_  & \new_[62812]_ ;
  assign \new_[62819]_  = ~A299 & A298;
  assign \new_[62822]_  = A301 & A300;
  assign \new_[62823]_  = \new_[62822]_  & \new_[62819]_ ;
  assign \new_[62824]_  = \new_[62823]_  & \new_[62816]_ ;
  assign \new_[62828]_  = A167 & ~A168;
  assign \new_[62829]_  = A169 & \new_[62828]_ ;
  assign \new_[62832]_  = ~A199 & ~A166;
  assign \new_[62835]_  = ~A233 & A200;
  assign \new_[62836]_  = \new_[62835]_  & \new_[62832]_ ;
  assign \new_[62837]_  = \new_[62836]_  & \new_[62829]_ ;
  assign \new_[62840]_  = ~A236 & ~A235;
  assign \new_[62843]_  = A266 & A265;
  assign \new_[62844]_  = \new_[62843]_  & \new_[62840]_ ;
  assign \new_[62847]_  = ~A299 & A298;
  assign \new_[62850]_  = A302 & A300;
  assign \new_[62851]_  = \new_[62850]_  & \new_[62847]_ ;
  assign \new_[62852]_  = \new_[62851]_  & \new_[62844]_ ;
  assign \new_[62856]_  = A167 & ~A168;
  assign \new_[62857]_  = A169 & \new_[62856]_ ;
  assign \new_[62860]_  = ~A199 & ~A166;
  assign \new_[62863]_  = ~A233 & A200;
  assign \new_[62864]_  = \new_[62863]_  & \new_[62860]_ ;
  assign \new_[62865]_  = \new_[62864]_  & \new_[62857]_ ;
  assign \new_[62868]_  = ~A236 & ~A235;
  assign \new_[62871]_  = ~A267 & ~A266;
  assign \new_[62872]_  = \new_[62871]_  & \new_[62868]_ ;
  assign \new_[62875]_  = ~A299 & A298;
  assign \new_[62878]_  = A301 & A300;
  assign \new_[62879]_  = \new_[62878]_  & \new_[62875]_ ;
  assign \new_[62880]_  = \new_[62879]_  & \new_[62872]_ ;
  assign \new_[62884]_  = A167 & ~A168;
  assign \new_[62885]_  = A169 & \new_[62884]_ ;
  assign \new_[62888]_  = ~A199 & ~A166;
  assign \new_[62891]_  = ~A233 & A200;
  assign \new_[62892]_  = \new_[62891]_  & \new_[62888]_ ;
  assign \new_[62893]_  = \new_[62892]_  & \new_[62885]_ ;
  assign \new_[62896]_  = ~A236 & ~A235;
  assign \new_[62899]_  = ~A267 & ~A266;
  assign \new_[62900]_  = \new_[62899]_  & \new_[62896]_ ;
  assign \new_[62903]_  = ~A299 & A298;
  assign \new_[62906]_  = A302 & A300;
  assign \new_[62907]_  = \new_[62906]_  & \new_[62903]_ ;
  assign \new_[62908]_  = \new_[62907]_  & \new_[62900]_ ;
  assign \new_[62912]_  = A167 & ~A168;
  assign \new_[62913]_  = A169 & \new_[62912]_ ;
  assign \new_[62916]_  = ~A199 & ~A166;
  assign \new_[62919]_  = ~A233 & A200;
  assign \new_[62920]_  = \new_[62919]_  & \new_[62916]_ ;
  assign \new_[62921]_  = \new_[62920]_  & \new_[62913]_ ;
  assign \new_[62924]_  = ~A236 & ~A235;
  assign \new_[62927]_  = ~A266 & ~A265;
  assign \new_[62928]_  = \new_[62927]_  & \new_[62924]_ ;
  assign \new_[62931]_  = ~A299 & A298;
  assign \new_[62934]_  = A301 & A300;
  assign \new_[62935]_  = \new_[62934]_  & \new_[62931]_ ;
  assign \new_[62936]_  = \new_[62935]_  & \new_[62928]_ ;
  assign \new_[62940]_  = A167 & ~A168;
  assign \new_[62941]_  = A169 & \new_[62940]_ ;
  assign \new_[62944]_  = ~A199 & ~A166;
  assign \new_[62947]_  = ~A233 & A200;
  assign \new_[62948]_  = \new_[62947]_  & \new_[62944]_ ;
  assign \new_[62949]_  = \new_[62948]_  & \new_[62941]_ ;
  assign \new_[62952]_  = ~A236 & ~A235;
  assign \new_[62955]_  = ~A266 & ~A265;
  assign \new_[62956]_  = \new_[62955]_  & \new_[62952]_ ;
  assign \new_[62959]_  = ~A299 & A298;
  assign \new_[62962]_  = A302 & A300;
  assign \new_[62963]_  = \new_[62962]_  & \new_[62959]_ ;
  assign \new_[62964]_  = \new_[62963]_  & \new_[62956]_ ;
  assign \new_[62968]_  = A167 & ~A168;
  assign \new_[62969]_  = A169 & \new_[62968]_ ;
  assign \new_[62972]_  = ~A199 & ~A166;
  assign \new_[62975]_  = ~A233 & A200;
  assign \new_[62976]_  = \new_[62975]_  & \new_[62972]_ ;
  assign \new_[62977]_  = \new_[62976]_  & \new_[62969]_ ;
  assign \new_[62980]_  = ~A266 & ~A234;
  assign \new_[62983]_  = ~A269 & ~A268;
  assign \new_[62984]_  = \new_[62983]_  & \new_[62980]_ ;
  assign \new_[62987]_  = ~A299 & A298;
  assign \new_[62990]_  = A301 & A300;
  assign \new_[62991]_  = \new_[62990]_  & \new_[62987]_ ;
  assign \new_[62992]_  = \new_[62991]_  & \new_[62984]_ ;
  assign \new_[62996]_  = A167 & ~A168;
  assign \new_[62997]_  = A169 & \new_[62996]_ ;
  assign \new_[63000]_  = ~A199 & ~A166;
  assign \new_[63003]_  = ~A233 & A200;
  assign \new_[63004]_  = \new_[63003]_  & \new_[63000]_ ;
  assign \new_[63005]_  = \new_[63004]_  & \new_[62997]_ ;
  assign \new_[63008]_  = ~A266 & ~A234;
  assign \new_[63011]_  = ~A269 & ~A268;
  assign \new_[63012]_  = \new_[63011]_  & \new_[63008]_ ;
  assign \new_[63015]_  = ~A299 & A298;
  assign \new_[63018]_  = A302 & A300;
  assign \new_[63019]_  = \new_[63018]_  & \new_[63015]_ ;
  assign \new_[63020]_  = \new_[63019]_  & \new_[63012]_ ;
  assign \new_[63024]_  = A167 & ~A168;
  assign \new_[63025]_  = A169 & \new_[63024]_ ;
  assign \new_[63028]_  = ~A199 & ~A166;
  assign \new_[63031]_  = ~A232 & A200;
  assign \new_[63032]_  = \new_[63031]_  & \new_[63028]_ ;
  assign \new_[63033]_  = \new_[63032]_  & \new_[63025]_ ;
  assign \new_[63036]_  = ~A266 & ~A233;
  assign \new_[63039]_  = ~A269 & ~A268;
  assign \new_[63040]_  = \new_[63039]_  & \new_[63036]_ ;
  assign \new_[63043]_  = ~A299 & A298;
  assign \new_[63046]_  = A301 & A300;
  assign \new_[63047]_  = \new_[63046]_  & \new_[63043]_ ;
  assign \new_[63048]_  = \new_[63047]_  & \new_[63040]_ ;
  assign \new_[63052]_  = A167 & ~A168;
  assign \new_[63053]_  = A169 & \new_[63052]_ ;
  assign \new_[63056]_  = ~A199 & ~A166;
  assign \new_[63059]_  = ~A232 & A200;
  assign \new_[63060]_  = \new_[63059]_  & \new_[63056]_ ;
  assign \new_[63061]_  = \new_[63060]_  & \new_[63053]_ ;
  assign \new_[63064]_  = ~A266 & ~A233;
  assign \new_[63067]_  = ~A269 & ~A268;
  assign \new_[63068]_  = \new_[63067]_  & \new_[63064]_ ;
  assign \new_[63071]_  = ~A299 & A298;
  assign \new_[63074]_  = A302 & A300;
  assign \new_[63075]_  = \new_[63074]_  & \new_[63071]_ ;
  assign \new_[63076]_  = \new_[63075]_  & \new_[63068]_ ;
  assign \new_[63080]_  = A167 & ~A168;
  assign \new_[63081]_  = A169 & \new_[63080]_ ;
  assign \new_[63084]_  = A199 & ~A166;
  assign \new_[63087]_  = A201 & ~A200;
  assign \new_[63088]_  = \new_[63087]_  & \new_[63084]_ ;
  assign \new_[63089]_  = \new_[63088]_  & \new_[63081]_ ;
  assign \new_[63092]_  = A232 & A202;
  assign \new_[63095]_  = A265 & A233;
  assign \new_[63096]_  = \new_[63095]_  & \new_[63092]_ ;
  assign \new_[63099]_  = ~A269 & ~A268;
  assign \new_[63102]_  = A299 & ~A298;
  assign \new_[63103]_  = \new_[63102]_  & \new_[63099]_ ;
  assign \new_[63104]_  = \new_[63103]_  & \new_[63096]_ ;
  assign \new_[63108]_  = A167 & ~A168;
  assign \new_[63109]_  = A169 & \new_[63108]_ ;
  assign \new_[63112]_  = A199 & ~A166;
  assign \new_[63115]_  = A201 & ~A200;
  assign \new_[63116]_  = \new_[63115]_  & \new_[63112]_ ;
  assign \new_[63117]_  = \new_[63116]_  & \new_[63109]_ ;
  assign \new_[63120]_  = ~A233 & A202;
  assign \new_[63123]_  = ~A236 & ~A235;
  assign \new_[63124]_  = \new_[63123]_  & \new_[63120]_ ;
  assign \new_[63127]_  = A266 & A265;
  assign \new_[63130]_  = A299 & ~A298;
  assign \new_[63131]_  = \new_[63130]_  & \new_[63127]_ ;
  assign \new_[63132]_  = \new_[63131]_  & \new_[63124]_ ;
  assign \new_[63136]_  = A167 & ~A168;
  assign \new_[63137]_  = A169 & \new_[63136]_ ;
  assign \new_[63140]_  = A199 & ~A166;
  assign \new_[63143]_  = A201 & ~A200;
  assign \new_[63144]_  = \new_[63143]_  & \new_[63140]_ ;
  assign \new_[63145]_  = \new_[63144]_  & \new_[63137]_ ;
  assign \new_[63148]_  = ~A233 & A202;
  assign \new_[63151]_  = ~A236 & ~A235;
  assign \new_[63152]_  = \new_[63151]_  & \new_[63148]_ ;
  assign \new_[63155]_  = ~A267 & ~A266;
  assign \new_[63158]_  = A299 & ~A298;
  assign \new_[63159]_  = \new_[63158]_  & \new_[63155]_ ;
  assign \new_[63160]_  = \new_[63159]_  & \new_[63152]_ ;
  assign \new_[63164]_  = A167 & ~A168;
  assign \new_[63165]_  = A169 & \new_[63164]_ ;
  assign \new_[63168]_  = A199 & ~A166;
  assign \new_[63171]_  = A201 & ~A200;
  assign \new_[63172]_  = \new_[63171]_  & \new_[63168]_ ;
  assign \new_[63173]_  = \new_[63172]_  & \new_[63165]_ ;
  assign \new_[63176]_  = ~A233 & A202;
  assign \new_[63179]_  = ~A236 & ~A235;
  assign \new_[63180]_  = \new_[63179]_  & \new_[63176]_ ;
  assign \new_[63183]_  = ~A266 & ~A265;
  assign \new_[63186]_  = A299 & ~A298;
  assign \new_[63187]_  = \new_[63186]_  & \new_[63183]_ ;
  assign \new_[63188]_  = \new_[63187]_  & \new_[63180]_ ;
  assign \new_[63192]_  = A167 & ~A168;
  assign \new_[63193]_  = A169 & \new_[63192]_ ;
  assign \new_[63196]_  = A199 & ~A166;
  assign \new_[63199]_  = A201 & ~A200;
  assign \new_[63200]_  = \new_[63199]_  & \new_[63196]_ ;
  assign \new_[63201]_  = \new_[63200]_  & \new_[63193]_ ;
  assign \new_[63204]_  = ~A233 & A202;
  assign \new_[63207]_  = ~A266 & ~A234;
  assign \new_[63208]_  = \new_[63207]_  & \new_[63204]_ ;
  assign \new_[63211]_  = ~A269 & ~A268;
  assign \new_[63214]_  = A299 & ~A298;
  assign \new_[63215]_  = \new_[63214]_  & \new_[63211]_ ;
  assign \new_[63216]_  = \new_[63215]_  & \new_[63208]_ ;
  assign \new_[63220]_  = A167 & ~A168;
  assign \new_[63221]_  = A169 & \new_[63220]_ ;
  assign \new_[63224]_  = A199 & ~A166;
  assign \new_[63227]_  = A201 & ~A200;
  assign \new_[63228]_  = \new_[63227]_  & \new_[63224]_ ;
  assign \new_[63229]_  = \new_[63228]_  & \new_[63221]_ ;
  assign \new_[63232]_  = A232 & A202;
  assign \new_[63235]_  = A234 & ~A233;
  assign \new_[63236]_  = \new_[63235]_  & \new_[63232]_ ;
  assign \new_[63239]_  = A298 & A235;
  assign \new_[63242]_  = ~A302 & ~A301;
  assign \new_[63243]_  = \new_[63242]_  & \new_[63239]_ ;
  assign \new_[63244]_  = \new_[63243]_  & \new_[63236]_ ;
  assign \new_[63248]_  = A167 & ~A168;
  assign \new_[63249]_  = A169 & \new_[63248]_ ;
  assign \new_[63252]_  = A199 & ~A166;
  assign \new_[63255]_  = A201 & ~A200;
  assign \new_[63256]_  = \new_[63255]_  & \new_[63252]_ ;
  assign \new_[63257]_  = \new_[63256]_  & \new_[63249]_ ;
  assign \new_[63260]_  = A232 & A202;
  assign \new_[63263]_  = A234 & ~A233;
  assign \new_[63264]_  = \new_[63263]_  & \new_[63260]_ ;
  assign \new_[63267]_  = A298 & A236;
  assign \new_[63270]_  = ~A302 & ~A301;
  assign \new_[63271]_  = \new_[63270]_  & \new_[63267]_ ;
  assign \new_[63272]_  = \new_[63271]_  & \new_[63264]_ ;
  assign \new_[63276]_  = A167 & ~A168;
  assign \new_[63277]_  = A169 & \new_[63276]_ ;
  assign \new_[63280]_  = A199 & ~A166;
  assign \new_[63283]_  = A201 & ~A200;
  assign \new_[63284]_  = \new_[63283]_  & \new_[63280]_ ;
  assign \new_[63285]_  = \new_[63284]_  & \new_[63277]_ ;
  assign \new_[63288]_  = ~A232 & A202;
  assign \new_[63291]_  = ~A266 & ~A233;
  assign \new_[63292]_  = \new_[63291]_  & \new_[63288]_ ;
  assign \new_[63295]_  = ~A269 & ~A268;
  assign \new_[63298]_  = A299 & ~A298;
  assign \new_[63299]_  = \new_[63298]_  & \new_[63295]_ ;
  assign \new_[63300]_  = \new_[63299]_  & \new_[63292]_ ;
  assign \new_[63304]_  = A167 & ~A168;
  assign \new_[63305]_  = A169 & \new_[63304]_ ;
  assign \new_[63308]_  = A199 & ~A166;
  assign \new_[63311]_  = A201 & ~A200;
  assign \new_[63312]_  = \new_[63311]_  & \new_[63308]_ ;
  assign \new_[63313]_  = \new_[63312]_  & \new_[63305]_ ;
  assign \new_[63316]_  = A232 & A203;
  assign \new_[63319]_  = A265 & A233;
  assign \new_[63320]_  = \new_[63319]_  & \new_[63316]_ ;
  assign \new_[63323]_  = ~A269 & ~A268;
  assign \new_[63326]_  = A299 & ~A298;
  assign \new_[63327]_  = \new_[63326]_  & \new_[63323]_ ;
  assign \new_[63328]_  = \new_[63327]_  & \new_[63320]_ ;
  assign \new_[63332]_  = A167 & ~A168;
  assign \new_[63333]_  = A169 & \new_[63332]_ ;
  assign \new_[63336]_  = A199 & ~A166;
  assign \new_[63339]_  = A201 & ~A200;
  assign \new_[63340]_  = \new_[63339]_  & \new_[63336]_ ;
  assign \new_[63341]_  = \new_[63340]_  & \new_[63333]_ ;
  assign \new_[63344]_  = ~A233 & A203;
  assign \new_[63347]_  = ~A236 & ~A235;
  assign \new_[63348]_  = \new_[63347]_  & \new_[63344]_ ;
  assign \new_[63351]_  = A266 & A265;
  assign \new_[63354]_  = A299 & ~A298;
  assign \new_[63355]_  = \new_[63354]_  & \new_[63351]_ ;
  assign \new_[63356]_  = \new_[63355]_  & \new_[63348]_ ;
  assign \new_[63360]_  = A167 & ~A168;
  assign \new_[63361]_  = A169 & \new_[63360]_ ;
  assign \new_[63364]_  = A199 & ~A166;
  assign \new_[63367]_  = A201 & ~A200;
  assign \new_[63368]_  = \new_[63367]_  & \new_[63364]_ ;
  assign \new_[63369]_  = \new_[63368]_  & \new_[63361]_ ;
  assign \new_[63372]_  = ~A233 & A203;
  assign \new_[63375]_  = ~A236 & ~A235;
  assign \new_[63376]_  = \new_[63375]_  & \new_[63372]_ ;
  assign \new_[63379]_  = ~A267 & ~A266;
  assign \new_[63382]_  = A299 & ~A298;
  assign \new_[63383]_  = \new_[63382]_  & \new_[63379]_ ;
  assign \new_[63384]_  = \new_[63383]_  & \new_[63376]_ ;
  assign \new_[63388]_  = A167 & ~A168;
  assign \new_[63389]_  = A169 & \new_[63388]_ ;
  assign \new_[63392]_  = A199 & ~A166;
  assign \new_[63395]_  = A201 & ~A200;
  assign \new_[63396]_  = \new_[63395]_  & \new_[63392]_ ;
  assign \new_[63397]_  = \new_[63396]_  & \new_[63389]_ ;
  assign \new_[63400]_  = ~A233 & A203;
  assign \new_[63403]_  = ~A236 & ~A235;
  assign \new_[63404]_  = \new_[63403]_  & \new_[63400]_ ;
  assign \new_[63407]_  = ~A266 & ~A265;
  assign \new_[63410]_  = A299 & ~A298;
  assign \new_[63411]_  = \new_[63410]_  & \new_[63407]_ ;
  assign \new_[63412]_  = \new_[63411]_  & \new_[63404]_ ;
  assign \new_[63416]_  = A167 & ~A168;
  assign \new_[63417]_  = A169 & \new_[63416]_ ;
  assign \new_[63420]_  = A199 & ~A166;
  assign \new_[63423]_  = A201 & ~A200;
  assign \new_[63424]_  = \new_[63423]_  & \new_[63420]_ ;
  assign \new_[63425]_  = \new_[63424]_  & \new_[63417]_ ;
  assign \new_[63428]_  = ~A233 & A203;
  assign \new_[63431]_  = ~A266 & ~A234;
  assign \new_[63432]_  = \new_[63431]_  & \new_[63428]_ ;
  assign \new_[63435]_  = ~A269 & ~A268;
  assign \new_[63438]_  = A299 & ~A298;
  assign \new_[63439]_  = \new_[63438]_  & \new_[63435]_ ;
  assign \new_[63440]_  = \new_[63439]_  & \new_[63432]_ ;
  assign \new_[63444]_  = A167 & ~A168;
  assign \new_[63445]_  = A169 & \new_[63444]_ ;
  assign \new_[63448]_  = A199 & ~A166;
  assign \new_[63451]_  = A201 & ~A200;
  assign \new_[63452]_  = \new_[63451]_  & \new_[63448]_ ;
  assign \new_[63453]_  = \new_[63452]_  & \new_[63445]_ ;
  assign \new_[63456]_  = A232 & A203;
  assign \new_[63459]_  = A234 & ~A233;
  assign \new_[63460]_  = \new_[63459]_  & \new_[63456]_ ;
  assign \new_[63463]_  = A298 & A235;
  assign \new_[63466]_  = ~A302 & ~A301;
  assign \new_[63467]_  = \new_[63466]_  & \new_[63463]_ ;
  assign \new_[63468]_  = \new_[63467]_  & \new_[63460]_ ;
  assign \new_[63472]_  = A167 & ~A168;
  assign \new_[63473]_  = A169 & \new_[63472]_ ;
  assign \new_[63476]_  = A199 & ~A166;
  assign \new_[63479]_  = A201 & ~A200;
  assign \new_[63480]_  = \new_[63479]_  & \new_[63476]_ ;
  assign \new_[63481]_  = \new_[63480]_  & \new_[63473]_ ;
  assign \new_[63484]_  = A232 & A203;
  assign \new_[63487]_  = A234 & ~A233;
  assign \new_[63488]_  = \new_[63487]_  & \new_[63484]_ ;
  assign \new_[63491]_  = A298 & A236;
  assign \new_[63494]_  = ~A302 & ~A301;
  assign \new_[63495]_  = \new_[63494]_  & \new_[63491]_ ;
  assign \new_[63496]_  = \new_[63495]_  & \new_[63488]_ ;
  assign \new_[63500]_  = A167 & ~A168;
  assign \new_[63501]_  = A169 & \new_[63500]_ ;
  assign \new_[63504]_  = A199 & ~A166;
  assign \new_[63507]_  = A201 & ~A200;
  assign \new_[63508]_  = \new_[63507]_  & \new_[63504]_ ;
  assign \new_[63509]_  = \new_[63508]_  & \new_[63501]_ ;
  assign \new_[63512]_  = ~A232 & A203;
  assign \new_[63515]_  = ~A266 & ~A233;
  assign \new_[63516]_  = \new_[63515]_  & \new_[63512]_ ;
  assign \new_[63519]_  = ~A269 & ~A268;
  assign \new_[63522]_  = A299 & ~A298;
  assign \new_[63523]_  = \new_[63522]_  & \new_[63519]_ ;
  assign \new_[63524]_  = \new_[63523]_  & \new_[63516]_ ;
  assign \new_[63528]_  = ~A167 & ~A168;
  assign \new_[63529]_  = A169 & \new_[63528]_ ;
  assign \new_[63532]_  = ~A199 & A166;
  assign \new_[63535]_  = A232 & A200;
  assign \new_[63536]_  = \new_[63535]_  & \new_[63532]_ ;
  assign \new_[63537]_  = \new_[63536]_  & \new_[63529]_ ;
  assign \new_[63540]_  = A265 & A233;
  assign \new_[63543]_  = ~A269 & ~A268;
  assign \new_[63544]_  = \new_[63543]_  & \new_[63540]_ ;
  assign \new_[63547]_  = ~A299 & A298;
  assign \new_[63550]_  = A301 & A300;
  assign \new_[63551]_  = \new_[63550]_  & \new_[63547]_ ;
  assign \new_[63552]_  = \new_[63551]_  & \new_[63544]_ ;
  assign \new_[63556]_  = ~A167 & ~A168;
  assign \new_[63557]_  = A169 & \new_[63556]_ ;
  assign \new_[63560]_  = ~A199 & A166;
  assign \new_[63563]_  = A232 & A200;
  assign \new_[63564]_  = \new_[63563]_  & \new_[63560]_ ;
  assign \new_[63565]_  = \new_[63564]_  & \new_[63557]_ ;
  assign \new_[63568]_  = A265 & A233;
  assign \new_[63571]_  = ~A269 & ~A268;
  assign \new_[63572]_  = \new_[63571]_  & \new_[63568]_ ;
  assign \new_[63575]_  = ~A299 & A298;
  assign \new_[63578]_  = A302 & A300;
  assign \new_[63579]_  = \new_[63578]_  & \new_[63575]_ ;
  assign \new_[63580]_  = \new_[63579]_  & \new_[63572]_ ;
  assign \new_[63584]_  = ~A167 & ~A168;
  assign \new_[63585]_  = A169 & \new_[63584]_ ;
  assign \new_[63588]_  = ~A199 & A166;
  assign \new_[63591]_  = ~A233 & A200;
  assign \new_[63592]_  = \new_[63591]_  & \new_[63588]_ ;
  assign \new_[63593]_  = \new_[63592]_  & \new_[63585]_ ;
  assign \new_[63596]_  = ~A236 & ~A235;
  assign \new_[63599]_  = A266 & A265;
  assign \new_[63600]_  = \new_[63599]_  & \new_[63596]_ ;
  assign \new_[63603]_  = ~A299 & A298;
  assign \new_[63606]_  = A301 & A300;
  assign \new_[63607]_  = \new_[63606]_  & \new_[63603]_ ;
  assign \new_[63608]_  = \new_[63607]_  & \new_[63600]_ ;
  assign \new_[63612]_  = ~A167 & ~A168;
  assign \new_[63613]_  = A169 & \new_[63612]_ ;
  assign \new_[63616]_  = ~A199 & A166;
  assign \new_[63619]_  = ~A233 & A200;
  assign \new_[63620]_  = \new_[63619]_  & \new_[63616]_ ;
  assign \new_[63621]_  = \new_[63620]_  & \new_[63613]_ ;
  assign \new_[63624]_  = ~A236 & ~A235;
  assign \new_[63627]_  = A266 & A265;
  assign \new_[63628]_  = \new_[63627]_  & \new_[63624]_ ;
  assign \new_[63631]_  = ~A299 & A298;
  assign \new_[63634]_  = A302 & A300;
  assign \new_[63635]_  = \new_[63634]_  & \new_[63631]_ ;
  assign \new_[63636]_  = \new_[63635]_  & \new_[63628]_ ;
  assign \new_[63640]_  = ~A167 & ~A168;
  assign \new_[63641]_  = A169 & \new_[63640]_ ;
  assign \new_[63644]_  = ~A199 & A166;
  assign \new_[63647]_  = ~A233 & A200;
  assign \new_[63648]_  = \new_[63647]_  & \new_[63644]_ ;
  assign \new_[63649]_  = \new_[63648]_  & \new_[63641]_ ;
  assign \new_[63652]_  = ~A236 & ~A235;
  assign \new_[63655]_  = ~A267 & ~A266;
  assign \new_[63656]_  = \new_[63655]_  & \new_[63652]_ ;
  assign \new_[63659]_  = ~A299 & A298;
  assign \new_[63662]_  = A301 & A300;
  assign \new_[63663]_  = \new_[63662]_  & \new_[63659]_ ;
  assign \new_[63664]_  = \new_[63663]_  & \new_[63656]_ ;
  assign \new_[63668]_  = ~A167 & ~A168;
  assign \new_[63669]_  = A169 & \new_[63668]_ ;
  assign \new_[63672]_  = ~A199 & A166;
  assign \new_[63675]_  = ~A233 & A200;
  assign \new_[63676]_  = \new_[63675]_  & \new_[63672]_ ;
  assign \new_[63677]_  = \new_[63676]_  & \new_[63669]_ ;
  assign \new_[63680]_  = ~A236 & ~A235;
  assign \new_[63683]_  = ~A267 & ~A266;
  assign \new_[63684]_  = \new_[63683]_  & \new_[63680]_ ;
  assign \new_[63687]_  = ~A299 & A298;
  assign \new_[63690]_  = A302 & A300;
  assign \new_[63691]_  = \new_[63690]_  & \new_[63687]_ ;
  assign \new_[63692]_  = \new_[63691]_  & \new_[63684]_ ;
  assign \new_[63696]_  = ~A167 & ~A168;
  assign \new_[63697]_  = A169 & \new_[63696]_ ;
  assign \new_[63700]_  = ~A199 & A166;
  assign \new_[63703]_  = ~A233 & A200;
  assign \new_[63704]_  = \new_[63703]_  & \new_[63700]_ ;
  assign \new_[63705]_  = \new_[63704]_  & \new_[63697]_ ;
  assign \new_[63708]_  = ~A236 & ~A235;
  assign \new_[63711]_  = ~A266 & ~A265;
  assign \new_[63712]_  = \new_[63711]_  & \new_[63708]_ ;
  assign \new_[63715]_  = ~A299 & A298;
  assign \new_[63718]_  = A301 & A300;
  assign \new_[63719]_  = \new_[63718]_  & \new_[63715]_ ;
  assign \new_[63720]_  = \new_[63719]_  & \new_[63712]_ ;
  assign \new_[63724]_  = ~A167 & ~A168;
  assign \new_[63725]_  = A169 & \new_[63724]_ ;
  assign \new_[63728]_  = ~A199 & A166;
  assign \new_[63731]_  = ~A233 & A200;
  assign \new_[63732]_  = \new_[63731]_  & \new_[63728]_ ;
  assign \new_[63733]_  = \new_[63732]_  & \new_[63725]_ ;
  assign \new_[63736]_  = ~A236 & ~A235;
  assign \new_[63739]_  = ~A266 & ~A265;
  assign \new_[63740]_  = \new_[63739]_  & \new_[63736]_ ;
  assign \new_[63743]_  = ~A299 & A298;
  assign \new_[63746]_  = A302 & A300;
  assign \new_[63747]_  = \new_[63746]_  & \new_[63743]_ ;
  assign \new_[63748]_  = \new_[63747]_  & \new_[63740]_ ;
  assign \new_[63752]_  = ~A167 & ~A168;
  assign \new_[63753]_  = A169 & \new_[63752]_ ;
  assign \new_[63756]_  = ~A199 & A166;
  assign \new_[63759]_  = ~A233 & A200;
  assign \new_[63760]_  = \new_[63759]_  & \new_[63756]_ ;
  assign \new_[63761]_  = \new_[63760]_  & \new_[63753]_ ;
  assign \new_[63764]_  = ~A266 & ~A234;
  assign \new_[63767]_  = ~A269 & ~A268;
  assign \new_[63768]_  = \new_[63767]_  & \new_[63764]_ ;
  assign \new_[63771]_  = ~A299 & A298;
  assign \new_[63774]_  = A301 & A300;
  assign \new_[63775]_  = \new_[63774]_  & \new_[63771]_ ;
  assign \new_[63776]_  = \new_[63775]_  & \new_[63768]_ ;
  assign \new_[63780]_  = ~A167 & ~A168;
  assign \new_[63781]_  = A169 & \new_[63780]_ ;
  assign \new_[63784]_  = ~A199 & A166;
  assign \new_[63787]_  = ~A233 & A200;
  assign \new_[63788]_  = \new_[63787]_  & \new_[63784]_ ;
  assign \new_[63789]_  = \new_[63788]_  & \new_[63781]_ ;
  assign \new_[63792]_  = ~A266 & ~A234;
  assign \new_[63795]_  = ~A269 & ~A268;
  assign \new_[63796]_  = \new_[63795]_  & \new_[63792]_ ;
  assign \new_[63799]_  = ~A299 & A298;
  assign \new_[63802]_  = A302 & A300;
  assign \new_[63803]_  = \new_[63802]_  & \new_[63799]_ ;
  assign \new_[63804]_  = \new_[63803]_  & \new_[63796]_ ;
  assign \new_[63808]_  = ~A167 & ~A168;
  assign \new_[63809]_  = A169 & \new_[63808]_ ;
  assign \new_[63812]_  = ~A199 & A166;
  assign \new_[63815]_  = ~A232 & A200;
  assign \new_[63816]_  = \new_[63815]_  & \new_[63812]_ ;
  assign \new_[63817]_  = \new_[63816]_  & \new_[63809]_ ;
  assign \new_[63820]_  = ~A266 & ~A233;
  assign \new_[63823]_  = ~A269 & ~A268;
  assign \new_[63824]_  = \new_[63823]_  & \new_[63820]_ ;
  assign \new_[63827]_  = ~A299 & A298;
  assign \new_[63830]_  = A301 & A300;
  assign \new_[63831]_  = \new_[63830]_  & \new_[63827]_ ;
  assign \new_[63832]_  = \new_[63831]_  & \new_[63824]_ ;
  assign \new_[63836]_  = ~A167 & ~A168;
  assign \new_[63837]_  = A169 & \new_[63836]_ ;
  assign \new_[63840]_  = ~A199 & A166;
  assign \new_[63843]_  = ~A232 & A200;
  assign \new_[63844]_  = \new_[63843]_  & \new_[63840]_ ;
  assign \new_[63845]_  = \new_[63844]_  & \new_[63837]_ ;
  assign \new_[63848]_  = ~A266 & ~A233;
  assign \new_[63851]_  = ~A269 & ~A268;
  assign \new_[63852]_  = \new_[63851]_  & \new_[63848]_ ;
  assign \new_[63855]_  = ~A299 & A298;
  assign \new_[63858]_  = A302 & A300;
  assign \new_[63859]_  = \new_[63858]_  & \new_[63855]_ ;
  assign \new_[63860]_  = \new_[63859]_  & \new_[63852]_ ;
  assign \new_[63864]_  = ~A167 & ~A168;
  assign \new_[63865]_  = A169 & \new_[63864]_ ;
  assign \new_[63868]_  = A199 & A166;
  assign \new_[63871]_  = A201 & ~A200;
  assign \new_[63872]_  = \new_[63871]_  & \new_[63868]_ ;
  assign \new_[63873]_  = \new_[63872]_  & \new_[63865]_ ;
  assign \new_[63876]_  = A232 & A202;
  assign \new_[63879]_  = A265 & A233;
  assign \new_[63880]_  = \new_[63879]_  & \new_[63876]_ ;
  assign \new_[63883]_  = ~A269 & ~A268;
  assign \new_[63886]_  = A299 & ~A298;
  assign \new_[63887]_  = \new_[63886]_  & \new_[63883]_ ;
  assign \new_[63888]_  = \new_[63887]_  & \new_[63880]_ ;
  assign \new_[63892]_  = ~A167 & ~A168;
  assign \new_[63893]_  = A169 & \new_[63892]_ ;
  assign \new_[63896]_  = A199 & A166;
  assign \new_[63899]_  = A201 & ~A200;
  assign \new_[63900]_  = \new_[63899]_  & \new_[63896]_ ;
  assign \new_[63901]_  = \new_[63900]_  & \new_[63893]_ ;
  assign \new_[63904]_  = ~A233 & A202;
  assign \new_[63907]_  = ~A236 & ~A235;
  assign \new_[63908]_  = \new_[63907]_  & \new_[63904]_ ;
  assign \new_[63911]_  = A266 & A265;
  assign \new_[63914]_  = A299 & ~A298;
  assign \new_[63915]_  = \new_[63914]_  & \new_[63911]_ ;
  assign \new_[63916]_  = \new_[63915]_  & \new_[63908]_ ;
  assign \new_[63920]_  = ~A167 & ~A168;
  assign \new_[63921]_  = A169 & \new_[63920]_ ;
  assign \new_[63924]_  = A199 & A166;
  assign \new_[63927]_  = A201 & ~A200;
  assign \new_[63928]_  = \new_[63927]_  & \new_[63924]_ ;
  assign \new_[63929]_  = \new_[63928]_  & \new_[63921]_ ;
  assign \new_[63932]_  = ~A233 & A202;
  assign \new_[63935]_  = ~A236 & ~A235;
  assign \new_[63936]_  = \new_[63935]_  & \new_[63932]_ ;
  assign \new_[63939]_  = ~A267 & ~A266;
  assign \new_[63942]_  = A299 & ~A298;
  assign \new_[63943]_  = \new_[63942]_  & \new_[63939]_ ;
  assign \new_[63944]_  = \new_[63943]_  & \new_[63936]_ ;
  assign \new_[63948]_  = ~A167 & ~A168;
  assign \new_[63949]_  = A169 & \new_[63948]_ ;
  assign \new_[63952]_  = A199 & A166;
  assign \new_[63955]_  = A201 & ~A200;
  assign \new_[63956]_  = \new_[63955]_  & \new_[63952]_ ;
  assign \new_[63957]_  = \new_[63956]_  & \new_[63949]_ ;
  assign \new_[63960]_  = ~A233 & A202;
  assign \new_[63963]_  = ~A236 & ~A235;
  assign \new_[63964]_  = \new_[63963]_  & \new_[63960]_ ;
  assign \new_[63967]_  = ~A266 & ~A265;
  assign \new_[63970]_  = A299 & ~A298;
  assign \new_[63971]_  = \new_[63970]_  & \new_[63967]_ ;
  assign \new_[63972]_  = \new_[63971]_  & \new_[63964]_ ;
  assign \new_[63976]_  = ~A167 & ~A168;
  assign \new_[63977]_  = A169 & \new_[63976]_ ;
  assign \new_[63980]_  = A199 & A166;
  assign \new_[63983]_  = A201 & ~A200;
  assign \new_[63984]_  = \new_[63983]_  & \new_[63980]_ ;
  assign \new_[63985]_  = \new_[63984]_  & \new_[63977]_ ;
  assign \new_[63988]_  = ~A233 & A202;
  assign \new_[63991]_  = ~A266 & ~A234;
  assign \new_[63992]_  = \new_[63991]_  & \new_[63988]_ ;
  assign \new_[63995]_  = ~A269 & ~A268;
  assign \new_[63998]_  = A299 & ~A298;
  assign \new_[63999]_  = \new_[63998]_  & \new_[63995]_ ;
  assign \new_[64000]_  = \new_[63999]_  & \new_[63992]_ ;
  assign \new_[64004]_  = ~A167 & ~A168;
  assign \new_[64005]_  = A169 & \new_[64004]_ ;
  assign \new_[64008]_  = A199 & A166;
  assign \new_[64011]_  = A201 & ~A200;
  assign \new_[64012]_  = \new_[64011]_  & \new_[64008]_ ;
  assign \new_[64013]_  = \new_[64012]_  & \new_[64005]_ ;
  assign \new_[64016]_  = A232 & A202;
  assign \new_[64019]_  = A234 & ~A233;
  assign \new_[64020]_  = \new_[64019]_  & \new_[64016]_ ;
  assign \new_[64023]_  = A298 & A235;
  assign \new_[64026]_  = ~A302 & ~A301;
  assign \new_[64027]_  = \new_[64026]_  & \new_[64023]_ ;
  assign \new_[64028]_  = \new_[64027]_  & \new_[64020]_ ;
  assign \new_[64032]_  = ~A167 & ~A168;
  assign \new_[64033]_  = A169 & \new_[64032]_ ;
  assign \new_[64036]_  = A199 & A166;
  assign \new_[64039]_  = A201 & ~A200;
  assign \new_[64040]_  = \new_[64039]_  & \new_[64036]_ ;
  assign \new_[64041]_  = \new_[64040]_  & \new_[64033]_ ;
  assign \new_[64044]_  = A232 & A202;
  assign \new_[64047]_  = A234 & ~A233;
  assign \new_[64048]_  = \new_[64047]_  & \new_[64044]_ ;
  assign \new_[64051]_  = A298 & A236;
  assign \new_[64054]_  = ~A302 & ~A301;
  assign \new_[64055]_  = \new_[64054]_  & \new_[64051]_ ;
  assign \new_[64056]_  = \new_[64055]_  & \new_[64048]_ ;
  assign \new_[64060]_  = ~A167 & ~A168;
  assign \new_[64061]_  = A169 & \new_[64060]_ ;
  assign \new_[64064]_  = A199 & A166;
  assign \new_[64067]_  = A201 & ~A200;
  assign \new_[64068]_  = \new_[64067]_  & \new_[64064]_ ;
  assign \new_[64069]_  = \new_[64068]_  & \new_[64061]_ ;
  assign \new_[64072]_  = ~A232 & A202;
  assign \new_[64075]_  = ~A266 & ~A233;
  assign \new_[64076]_  = \new_[64075]_  & \new_[64072]_ ;
  assign \new_[64079]_  = ~A269 & ~A268;
  assign \new_[64082]_  = A299 & ~A298;
  assign \new_[64083]_  = \new_[64082]_  & \new_[64079]_ ;
  assign \new_[64084]_  = \new_[64083]_  & \new_[64076]_ ;
  assign \new_[64088]_  = ~A167 & ~A168;
  assign \new_[64089]_  = A169 & \new_[64088]_ ;
  assign \new_[64092]_  = A199 & A166;
  assign \new_[64095]_  = A201 & ~A200;
  assign \new_[64096]_  = \new_[64095]_  & \new_[64092]_ ;
  assign \new_[64097]_  = \new_[64096]_  & \new_[64089]_ ;
  assign \new_[64100]_  = A232 & A203;
  assign \new_[64103]_  = A265 & A233;
  assign \new_[64104]_  = \new_[64103]_  & \new_[64100]_ ;
  assign \new_[64107]_  = ~A269 & ~A268;
  assign \new_[64110]_  = A299 & ~A298;
  assign \new_[64111]_  = \new_[64110]_  & \new_[64107]_ ;
  assign \new_[64112]_  = \new_[64111]_  & \new_[64104]_ ;
  assign \new_[64116]_  = ~A167 & ~A168;
  assign \new_[64117]_  = A169 & \new_[64116]_ ;
  assign \new_[64120]_  = A199 & A166;
  assign \new_[64123]_  = A201 & ~A200;
  assign \new_[64124]_  = \new_[64123]_  & \new_[64120]_ ;
  assign \new_[64125]_  = \new_[64124]_  & \new_[64117]_ ;
  assign \new_[64128]_  = ~A233 & A203;
  assign \new_[64131]_  = ~A236 & ~A235;
  assign \new_[64132]_  = \new_[64131]_  & \new_[64128]_ ;
  assign \new_[64135]_  = A266 & A265;
  assign \new_[64138]_  = A299 & ~A298;
  assign \new_[64139]_  = \new_[64138]_  & \new_[64135]_ ;
  assign \new_[64140]_  = \new_[64139]_  & \new_[64132]_ ;
  assign \new_[64144]_  = ~A167 & ~A168;
  assign \new_[64145]_  = A169 & \new_[64144]_ ;
  assign \new_[64148]_  = A199 & A166;
  assign \new_[64151]_  = A201 & ~A200;
  assign \new_[64152]_  = \new_[64151]_  & \new_[64148]_ ;
  assign \new_[64153]_  = \new_[64152]_  & \new_[64145]_ ;
  assign \new_[64156]_  = ~A233 & A203;
  assign \new_[64159]_  = ~A236 & ~A235;
  assign \new_[64160]_  = \new_[64159]_  & \new_[64156]_ ;
  assign \new_[64163]_  = ~A267 & ~A266;
  assign \new_[64166]_  = A299 & ~A298;
  assign \new_[64167]_  = \new_[64166]_  & \new_[64163]_ ;
  assign \new_[64168]_  = \new_[64167]_  & \new_[64160]_ ;
  assign \new_[64172]_  = ~A167 & ~A168;
  assign \new_[64173]_  = A169 & \new_[64172]_ ;
  assign \new_[64176]_  = A199 & A166;
  assign \new_[64179]_  = A201 & ~A200;
  assign \new_[64180]_  = \new_[64179]_  & \new_[64176]_ ;
  assign \new_[64181]_  = \new_[64180]_  & \new_[64173]_ ;
  assign \new_[64184]_  = ~A233 & A203;
  assign \new_[64187]_  = ~A236 & ~A235;
  assign \new_[64188]_  = \new_[64187]_  & \new_[64184]_ ;
  assign \new_[64191]_  = ~A266 & ~A265;
  assign \new_[64194]_  = A299 & ~A298;
  assign \new_[64195]_  = \new_[64194]_  & \new_[64191]_ ;
  assign \new_[64196]_  = \new_[64195]_  & \new_[64188]_ ;
  assign \new_[64200]_  = ~A167 & ~A168;
  assign \new_[64201]_  = A169 & \new_[64200]_ ;
  assign \new_[64204]_  = A199 & A166;
  assign \new_[64207]_  = A201 & ~A200;
  assign \new_[64208]_  = \new_[64207]_  & \new_[64204]_ ;
  assign \new_[64209]_  = \new_[64208]_  & \new_[64201]_ ;
  assign \new_[64212]_  = ~A233 & A203;
  assign \new_[64215]_  = ~A266 & ~A234;
  assign \new_[64216]_  = \new_[64215]_  & \new_[64212]_ ;
  assign \new_[64219]_  = ~A269 & ~A268;
  assign \new_[64222]_  = A299 & ~A298;
  assign \new_[64223]_  = \new_[64222]_  & \new_[64219]_ ;
  assign \new_[64224]_  = \new_[64223]_  & \new_[64216]_ ;
  assign \new_[64228]_  = ~A167 & ~A168;
  assign \new_[64229]_  = A169 & \new_[64228]_ ;
  assign \new_[64232]_  = A199 & A166;
  assign \new_[64235]_  = A201 & ~A200;
  assign \new_[64236]_  = \new_[64235]_  & \new_[64232]_ ;
  assign \new_[64237]_  = \new_[64236]_  & \new_[64229]_ ;
  assign \new_[64240]_  = A232 & A203;
  assign \new_[64243]_  = A234 & ~A233;
  assign \new_[64244]_  = \new_[64243]_  & \new_[64240]_ ;
  assign \new_[64247]_  = A298 & A235;
  assign \new_[64250]_  = ~A302 & ~A301;
  assign \new_[64251]_  = \new_[64250]_  & \new_[64247]_ ;
  assign \new_[64252]_  = \new_[64251]_  & \new_[64244]_ ;
  assign \new_[64256]_  = ~A167 & ~A168;
  assign \new_[64257]_  = A169 & \new_[64256]_ ;
  assign \new_[64260]_  = A199 & A166;
  assign \new_[64263]_  = A201 & ~A200;
  assign \new_[64264]_  = \new_[64263]_  & \new_[64260]_ ;
  assign \new_[64265]_  = \new_[64264]_  & \new_[64257]_ ;
  assign \new_[64268]_  = A232 & A203;
  assign \new_[64271]_  = A234 & ~A233;
  assign \new_[64272]_  = \new_[64271]_  & \new_[64268]_ ;
  assign \new_[64275]_  = A298 & A236;
  assign \new_[64278]_  = ~A302 & ~A301;
  assign \new_[64279]_  = \new_[64278]_  & \new_[64275]_ ;
  assign \new_[64280]_  = \new_[64279]_  & \new_[64272]_ ;
  assign \new_[64284]_  = ~A167 & ~A168;
  assign \new_[64285]_  = A169 & \new_[64284]_ ;
  assign \new_[64288]_  = A199 & A166;
  assign \new_[64291]_  = A201 & ~A200;
  assign \new_[64292]_  = \new_[64291]_  & \new_[64288]_ ;
  assign \new_[64293]_  = \new_[64292]_  & \new_[64285]_ ;
  assign \new_[64296]_  = ~A232 & A203;
  assign \new_[64299]_  = ~A266 & ~A233;
  assign \new_[64300]_  = \new_[64299]_  & \new_[64296]_ ;
  assign \new_[64303]_  = ~A269 & ~A268;
  assign \new_[64306]_  = A299 & ~A298;
  assign \new_[64307]_  = \new_[64306]_  & \new_[64303]_ ;
  assign \new_[64308]_  = \new_[64307]_  & \new_[64300]_ ;
  assign \new_[64312]_  = ~A168 & A169;
  assign \new_[64313]_  = A170 & \new_[64312]_ ;
  assign \new_[64316]_  = ~A200 & A199;
  assign \new_[64319]_  = A202 & A201;
  assign \new_[64320]_  = \new_[64319]_  & \new_[64316]_ ;
  assign \new_[64321]_  = \new_[64320]_  & \new_[64313]_ ;
  assign \new_[64324]_  = A233 & A232;
  assign \new_[64327]_  = ~A267 & A265;
  assign \new_[64328]_  = \new_[64327]_  & \new_[64324]_ ;
  assign \new_[64331]_  = ~A299 & A298;
  assign \new_[64334]_  = A301 & A300;
  assign \new_[64335]_  = \new_[64334]_  & \new_[64331]_ ;
  assign \new_[64336]_  = \new_[64335]_  & \new_[64328]_ ;
  assign \new_[64340]_  = ~A168 & A169;
  assign \new_[64341]_  = A170 & \new_[64340]_ ;
  assign \new_[64344]_  = ~A200 & A199;
  assign \new_[64347]_  = A202 & A201;
  assign \new_[64348]_  = \new_[64347]_  & \new_[64344]_ ;
  assign \new_[64349]_  = \new_[64348]_  & \new_[64341]_ ;
  assign \new_[64352]_  = A233 & A232;
  assign \new_[64355]_  = ~A267 & A265;
  assign \new_[64356]_  = \new_[64355]_  & \new_[64352]_ ;
  assign \new_[64359]_  = ~A299 & A298;
  assign \new_[64362]_  = A302 & A300;
  assign \new_[64363]_  = \new_[64362]_  & \new_[64359]_ ;
  assign \new_[64364]_  = \new_[64363]_  & \new_[64356]_ ;
  assign \new_[64368]_  = ~A168 & A169;
  assign \new_[64369]_  = A170 & \new_[64368]_ ;
  assign \new_[64372]_  = ~A200 & A199;
  assign \new_[64375]_  = A202 & A201;
  assign \new_[64376]_  = \new_[64375]_  & \new_[64372]_ ;
  assign \new_[64377]_  = \new_[64376]_  & \new_[64369]_ ;
  assign \new_[64380]_  = A233 & A232;
  assign \new_[64383]_  = A266 & A265;
  assign \new_[64384]_  = \new_[64383]_  & \new_[64380]_ ;
  assign \new_[64387]_  = ~A299 & A298;
  assign \new_[64390]_  = A301 & A300;
  assign \new_[64391]_  = \new_[64390]_  & \new_[64387]_ ;
  assign \new_[64392]_  = \new_[64391]_  & \new_[64384]_ ;
  assign \new_[64396]_  = ~A168 & A169;
  assign \new_[64397]_  = A170 & \new_[64396]_ ;
  assign \new_[64400]_  = ~A200 & A199;
  assign \new_[64403]_  = A202 & A201;
  assign \new_[64404]_  = \new_[64403]_  & \new_[64400]_ ;
  assign \new_[64405]_  = \new_[64404]_  & \new_[64397]_ ;
  assign \new_[64408]_  = A233 & A232;
  assign \new_[64411]_  = A266 & A265;
  assign \new_[64412]_  = \new_[64411]_  & \new_[64408]_ ;
  assign \new_[64415]_  = ~A299 & A298;
  assign \new_[64418]_  = A302 & A300;
  assign \new_[64419]_  = \new_[64418]_  & \new_[64415]_ ;
  assign \new_[64420]_  = \new_[64419]_  & \new_[64412]_ ;
  assign \new_[64424]_  = ~A168 & A169;
  assign \new_[64425]_  = A170 & \new_[64424]_ ;
  assign \new_[64428]_  = ~A200 & A199;
  assign \new_[64431]_  = A202 & A201;
  assign \new_[64432]_  = \new_[64431]_  & \new_[64428]_ ;
  assign \new_[64433]_  = \new_[64432]_  & \new_[64425]_ ;
  assign \new_[64436]_  = A233 & A232;
  assign \new_[64439]_  = ~A266 & ~A265;
  assign \new_[64440]_  = \new_[64439]_  & \new_[64436]_ ;
  assign \new_[64443]_  = ~A299 & A298;
  assign \new_[64446]_  = A301 & A300;
  assign \new_[64447]_  = \new_[64446]_  & \new_[64443]_ ;
  assign \new_[64448]_  = \new_[64447]_  & \new_[64440]_ ;
  assign \new_[64452]_  = ~A168 & A169;
  assign \new_[64453]_  = A170 & \new_[64452]_ ;
  assign \new_[64456]_  = ~A200 & A199;
  assign \new_[64459]_  = A202 & A201;
  assign \new_[64460]_  = \new_[64459]_  & \new_[64456]_ ;
  assign \new_[64461]_  = \new_[64460]_  & \new_[64453]_ ;
  assign \new_[64464]_  = A233 & A232;
  assign \new_[64467]_  = ~A266 & ~A265;
  assign \new_[64468]_  = \new_[64467]_  & \new_[64464]_ ;
  assign \new_[64471]_  = ~A299 & A298;
  assign \new_[64474]_  = A302 & A300;
  assign \new_[64475]_  = \new_[64474]_  & \new_[64471]_ ;
  assign \new_[64476]_  = \new_[64475]_  & \new_[64468]_ ;
  assign \new_[64480]_  = ~A168 & A169;
  assign \new_[64481]_  = A170 & \new_[64480]_ ;
  assign \new_[64484]_  = ~A200 & A199;
  assign \new_[64487]_  = A202 & A201;
  assign \new_[64488]_  = \new_[64487]_  & \new_[64484]_ ;
  assign \new_[64489]_  = \new_[64488]_  & \new_[64481]_ ;
  assign \new_[64492]_  = ~A235 & ~A233;
  assign \new_[64495]_  = ~A266 & ~A236;
  assign \new_[64496]_  = \new_[64495]_  & \new_[64492]_ ;
  assign \new_[64499]_  = ~A269 & ~A268;
  assign \new_[64502]_  = A299 & ~A298;
  assign \new_[64503]_  = \new_[64502]_  & \new_[64499]_ ;
  assign \new_[64504]_  = \new_[64503]_  & \new_[64496]_ ;
  assign \new_[64508]_  = ~A168 & A169;
  assign \new_[64509]_  = A170 & \new_[64508]_ ;
  assign \new_[64512]_  = ~A200 & A199;
  assign \new_[64515]_  = A202 & A201;
  assign \new_[64516]_  = \new_[64515]_  & \new_[64512]_ ;
  assign \new_[64517]_  = \new_[64516]_  & \new_[64509]_ ;
  assign \new_[64520]_  = ~A234 & ~A233;
  assign \new_[64523]_  = A266 & A265;
  assign \new_[64524]_  = \new_[64523]_  & \new_[64520]_ ;
  assign \new_[64527]_  = ~A299 & A298;
  assign \new_[64530]_  = A301 & A300;
  assign \new_[64531]_  = \new_[64530]_  & \new_[64527]_ ;
  assign \new_[64532]_  = \new_[64531]_  & \new_[64524]_ ;
  assign \new_[64536]_  = ~A168 & A169;
  assign \new_[64537]_  = A170 & \new_[64536]_ ;
  assign \new_[64540]_  = ~A200 & A199;
  assign \new_[64543]_  = A202 & A201;
  assign \new_[64544]_  = \new_[64543]_  & \new_[64540]_ ;
  assign \new_[64545]_  = \new_[64544]_  & \new_[64537]_ ;
  assign \new_[64548]_  = ~A234 & ~A233;
  assign \new_[64551]_  = A266 & A265;
  assign \new_[64552]_  = \new_[64551]_  & \new_[64548]_ ;
  assign \new_[64555]_  = ~A299 & A298;
  assign \new_[64558]_  = A302 & A300;
  assign \new_[64559]_  = \new_[64558]_  & \new_[64555]_ ;
  assign \new_[64560]_  = \new_[64559]_  & \new_[64552]_ ;
  assign \new_[64564]_  = ~A168 & A169;
  assign \new_[64565]_  = A170 & \new_[64564]_ ;
  assign \new_[64568]_  = ~A200 & A199;
  assign \new_[64571]_  = A202 & A201;
  assign \new_[64572]_  = \new_[64571]_  & \new_[64568]_ ;
  assign \new_[64573]_  = \new_[64572]_  & \new_[64565]_ ;
  assign \new_[64576]_  = ~A233 & A232;
  assign \new_[64579]_  = A235 & A234;
  assign \new_[64580]_  = \new_[64579]_  & \new_[64576]_ ;
  assign \new_[64583]_  = ~A266 & A265;
  assign \new_[64586]_  = A268 & A267;
  assign \new_[64587]_  = \new_[64586]_  & \new_[64583]_ ;
  assign \new_[64588]_  = \new_[64587]_  & \new_[64580]_ ;
  assign \new_[64592]_  = ~A168 & A169;
  assign \new_[64593]_  = A170 & \new_[64592]_ ;
  assign \new_[64596]_  = ~A200 & A199;
  assign \new_[64599]_  = A202 & A201;
  assign \new_[64600]_  = \new_[64599]_  & \new_[64596]_ ;
  assign \new_[64601]_  = \new_[64600]_  & \new_[64593]_ ;
  assign \new_[64604]_  = ~A233 & A232;
  assign \new_[64607]_  = A235 & A234;
  assign \new_[64608]_  = \new_[64607]_  & \new_[64604]_ ;
  assign \new_[64611]_  = ~A266 & A265;
  assign \new_[64614]_  = A269 & A267;
  assign \new_[64615]_  = \new_[64614]_  & \new_[64611]_ ;
  assign \new_[64616]_  = \new_[64615]_  & \new_[64608]_ ;
  assign \new_[64620]_  = ~A168 & A169;
  assign \new_[64621]_  = A170 & \new_[64620]_ ;
  assign \new_[64624]_  = ~A200 & A199;
  assign \new_[64627]_  = A202 & A201;
  assign \new_[64628]_  = \new_[64627]_  & \new_[64624]_ ;
  assign \new_[64629]_  = \new_[64628]_  & \new_[64621]_ ;
  assign \new_[64632]_  = ~A233 & A232;
  assign \new_[64635]_  = A236 & A234;
  assign \new_[64636]_  = \new_[64635]_  & \new_[64632]_ ;
  assign \new_[64639]_  = ~A266 & A265;
  assign \new_[64642]_  = A268 & A267;
  assign \new_[64643]_  = \new_[64642]_  & \new_[64639]_ ;
  assign \new_[64644]_  = \new_[64643]_  & \new_[64636]_ ;
  assign \new_[64648]_  = ~A168 & A169;
  assign \new_[64649]_  = A170 & \new_[64648]_ ;
  assign \new_[64652]_  = ~A200 & A199;
  assign \new_[64655]_  = A202 & A201;
  assign \new_[64656]_  = \new_[64655]_  & \new_[64652]_ ;
  assign \new_[64657]_  = \new_[64656]_  & \new_[64649]_ ;
  assign \new_[64660]_  = ~A233 & A232;
  assign \new_[64663]_  = A236 & A234;
  assign \new_[64664]_  = \new_[64663]_  & \new_[64660]_ ;
  assign \new_[64667]_  = ~A266 & A265;
  assign \new_[64670]_  = A269 & A267;
  assign \new_[64671]_  = \new_[64670]_  & \new_[64667]_ ;
  assign \new_[64672]_  = \new_[64671]_  & \new_[64664]_ ;
  assign \new_[64676]_  = ~A168 & A169;
  assign \new_[64677]_  = A170 & \new_[64676]_ ;
  assign \new_[64680]_  = ~A200 & A199;
  assign \new_[64683]_  = A202 & A201;
  assign \new_[64684]_  = \new_[64683]_  & \new_[64680]_ ;
  assign \new_[64685]_  = \new_[64684]_  & \new_[64677]_ ;
  assign \new_[64688]_  = ~A233 & ~A232;
  assign \new_[64691]_  = A266 & A265;
  assign \new_[64692]_  = \new_[64691]_  & \new_[64688]_ ;
  assign \new_[64695]_  = ~A299 & A298;
  assign \new_[64698]_  = A301 & A300;
  assign \new_[64699]_  = \new_[64698]_  & \new_[64695]_ ;
  assign \new_[64700]_  = \new_[64699]_  & \new_[64692]_ ;
  assign \new_[64704]_  = ~A168 & A169;
  assign \new_[64705]_  = A170 & \new_[64704]_ ;
  assign \new_[64708]_  = ~A200 & A199;
  assign \new_[64711]_  = A202 & A201;
  assign \new_[64712]_  = \new_[64711]_  & \new_[64708]_ ;
  assign \new_[64713]_  = \new_[64712]_  & \new_[64705]_ ;
  assign \new_[64716]_  = ~A233 & ~A232;
  assign \new_[64719]_  = A266 & A265;
  assign \new_[64720]_  = \new_[64719]_  & \new_[64716]_ ;
  assign \new_[64723]_  = ~A299 & A298;
  assign \new_[64726]_  = A302 & A300;
  assign \new_[64727]_  = \new_[64726]_  & \new_[64723]_ ;
  assign \new_[64728]_  = \new_[64727]_  & \new_[64720]_ ;
  assign \new_[64732]_  = ~A168 & A169;
  assign \new_[64733]_  = A170 & \new_[64732]_ ;
  assign \new_[64736]_  = ~A200 & A199;
  assign \new_[64739]_  = A203 & A201;
  assign \new_[64740]_  = \new_[64739]_  & \new_[64736]_ ;
  assign \new_[64741]_  = \new_[64740]_  & \new_[64733]_ ;
  assign \new_[64744]_  = A233 & A232;
  assign \new_[64747]_  = ~A267 & A265;
  assign \new_[64748]_  = \new_[64747]_  & \new_[64744]_ ;
  assign \new_[64751]_  = ~A299 & A298;
  assign \new_[64754]_  = A301 & A300;
  assign \new_[64755]_  = \new_[64754]_  & \new_[64751]_ ;
  assign \new_[64756]_  = \new_[64755]_  & \new_[64748]_ ;
  assign \new_[64760]_  = ~A168 & A169;
  assign \new_[64761]_  = A170 & \new_[64760]_ ;
  assign \new_[64764]_  = ~A200 & A199;
  assign \new_[64767]_  = A203 & A201;
  assign \new_[64768]_  = \new_[64767]_  & \new_[64764]_ ;
  assign \new_[64769]_  = \new_[64768]_  & \new_[64761]_ ;
  assign \new_[64772]_  = A233 & A232;
  assign \new_[64775]_  = ~A267 & A265;
  assign \new_[64776]_  = \new_[64775]_  & \new_[64772]_ ;
  assign \new_[64779]_  = ~A299 & A298;
  assign \new_[64782]_  = A302 & A300;
  assign \new_[64783]_  = \new_[64782]_  & \new_[64779]_ ;
  assign \new_[64784]_  = \new_[64783]_  & \new_[64776]_ ;
  assign \new_[64788]_  = ~A168 & A169;
  assign \new_[64789]_  = A170 & \new_[64788]_ ;
  assign \new_[64792]_  = ~A200 & A199;
  assign \new_[64795]_  = A203 & A201;
  assign \new_[64796]_  = \new_[64795]_  & \new_[64792]_ ;
  assign \new_[64797]_  = \new_[64796]_  & \new_[64789]_ ;
  assign \new_[64800]_  = A233 & A232;
  assign \new_[64803]_  = A266 & A265;
  assign \new_[64804]_  = \new_[64803]_  & \new_[64800]_ ;
  assign \new_[64807]_  = ~A299 & A298;
  assign \new_[64810]_  = A301 & A300;
  assign \new_[64811]_  = \new_[64810]_  & \new_[64807]_ ;
  assign \new_[64812]_  = \new_[64811]_  & \new_[64804]_ ;
  assign \new_[64816]_  = ~A168 & A169;
  assign \new_[64817]_  = A170 & \new_[64816]_ ;
  assign \new_[64820]_  = ~A200 & A199;
  assign \new_[64823]_  = A203 & A201;
  assign \new_[64824]_  = \new_[64823]_  & \new_[64820]_ ;
  assign \new_[64825]_  = \new_[64824]_  & \new_[64817]_ ;
  assign \new_[64828]_  = A233 & A232;
  assign \new_[64831]_  = A266 & A265;
  assign \new_[64832]_  = \new_[64831]_  & \new_[64828]_ ;
  assign \new_[64835]_  = ~A299 & A298;
  assign \new_[64838]_  = A302 & A300;
  assign \new_[64839]_  = \new_[64838]_  & \new_[64835]_ ;
  assign \new_[64840]_  = \new_[64839]_  & \new_[64832]_ ;
  assign \new_[64844]_  = ~A168 & A169;
  assign \new_[64845]_  = A170 & \new_[64844]_ ;
  assign \new_[64848]_  = ~A200 & A199;
  assign \new_[64851]_  = A203 & A201;
  assign \new_[64852]_  = \new_[64851]_  & \new_[64848]_ ;
  assign \new_[64853]_  = \new_[64852]_  & \new_[64845]_ ;
  assign \new_[64856]_  = A233 & A232;
  assign \new_[64859]_  = ~A266 & ~A265;
  assign \new_[64860]_  = \new_[64859]_  & \new_[64856]_ ;
  assign \new_[64863]_  = ~A299 & A298;
  assign \new_[64866]_  = A301 & A300;
  assign \new_[64867]_  = \new_[64866]_  & \new_[64863]_ ;
  assign \new_[64868]_  = \new_[64867]_  & \new_[64860]_ ;
  assign \new_[64872]_  = ~A168 & A169;
  assign \new_[64873]_  = A170 & \new_[64872]_ ;
  assign \new_[64876]_  = ~A200 & A199;
  assign \new_[64879]_  = A203 & A201;
  assign \new_[64880]_  = \new_[64879]_  & \new_[64876]_ ;
  assign \new_[64881]_  = \new_[64880]_  & \new_[64873]_ ;
  assign \new_[64884]_  = A233 & A232;
  assign \new_[64887]_  = ~A266 & ~A265;
  assign \new_[64888]_  = \new_[64887]_  & \new_[64884]_ ;
  assign \new_[64891]_  = ~A299 & A298;
  assign \new_[64894]_  = A302 & A300;
  assign \new_[64895]_  = \new_[64894]_  & \new_[64891]_ ;
  assign \new_[64896]_  = \new_[64895]_  & \new_[64888]_ ;
  assign \new_[64900]_  = ~A168 & A169;
  assign \new_[64901]_  = A170 & \new_[64900]_ ;
  assign \new_[64904]_  = ~A200 & A199;
  assign \new_[64907]_  = A203 & A201;
  assign \new_[64908]_  = \new_[64907]_  & \new_[64904]_ ;
  assign \new_[64909]_  = \new_[64908]_  & \new_[64901]_ ;
  assign \new_[64912]_  = ~A235 & ~A233;
  assign \new_[64915]_  = ~A266 & ~A236;
  assign \new_[64916]_  = \new_[64915]_  & \new_[64912]_ ;
  assign \new_[64919]_  = ~A269 & ~A268;
  assign \new_[64922]_  = A299 & ~A298;
  assign \new_[64923]_  = \new_[64922]_  & \new_[64919]_ ;
  assign \new_[64924]_  = \new_[64923]_  & \new_[64916]_ ;
  assign \new_[64928]_  = ~A168 & A169;
  assign \new_[64929]_  = A170 & \new_[64928]_ ;
  assign \new_[64932]_  = ~A200 & A199;
  assign \new_[64935]_  = A203 & A201;
  assign \new_[64936]_  = \new_[64935]_  & \new_[64932]_ ;
  assign \new_[64937]_  = \new_[64936]_  & \new_[64929]_ ;
  assign \new_[64940]_  = ~A234 & ~A233;
  assign \new_[64943]_  = A266 & A265;
  assign \new_[64944]_  = \new_[64943]_  & \new_[64940]_ ;
  assign \new_[64947]_  = ~A299 & A298;
  assign \new_[64950]_  = A301 & A300;
  assign \new_[64951]_  = \new_[64950]_  & \new_[64947]_ ;
  assign \new_[64952]_  = \new_[64951]_  & \new_[64944]_ ;
  assign \new_[64956]_  = ~A168 & A169;
  assign \new_[64957]_  = A170 & \new_[64956]_ ;
  assign \new_[64960]_  = ~A200 & A199;
  assign \new_[64963]_  = A203 & A201;
  assign \new_[64964]_  = \new_[64963]_  & \new_[64960]_ ;
  assign \new_[64965]_  = \new_[64964]_  & \new_[64957]_ ;
  assign \new_[64968]_  = ~A234 & ~A233;
  assign \new_[64971]_  = A266 & A265;
  assign \new_[64972]_  = \new_[64971]_  & \new_[64968]_ ;
  assign \new_[64975]_  = ~A299 & A298;
  assign \new_[64978]_  = A302 & A300;
  assign \new_[64979]_  = \new_[64978]_  & \new_[64975]_ ;
  assign \new_[64980]_  = \new_[64979]_  & \new_[64972]_ ;
  assign \new_[64984]_  = ~A168 & A169;
  assign \new_[64985]_  = A170 & \new_[64984]_ ;
  assign \new_[64988]_  = ~A200 & A199;
  assign \new_[64991]_  = A203 & A201;
  assign \new_[64992]_  = \new_[64991]_  & \new_[64988]_ ;
  assign \new_[64993]_  = \new_[64992]_  & \new_[64985]_ ;
  assign \new_[64996]_  = ~A233 & A232;
  assign \new_[64999]_  = A235 & A234;
  assign \new_[65000]_  = \new_[64999]_  & \new_[64996]_ ;
  assign \new_[65003]_  = ~A266 & A265;
  assign \new_[65006]_  = A268 & A267;
  assign \new_[65007]_  = \new_[65006]_  & \new_[65003]_ ;
  assign \new_[65008]_  = \new_[65007]_  & \new_[65000]_ ;
  assign \new_[65012]_  = ~A168 & A169;
  assign \new_[65013]_  = A170 & \new_[65012]_ ;
  assign \new_[65016]_  = ~A200 & A199;
  assign \new_[65019]_  = A203 & A201;
  assign \new_[65020]_  = \new_[65019]_  & \new_[65016]_ ;
  assign \new_[65021]_  = \new_[65020]_  & \new_[65013]_ ;
  assign \new_[65024]_  = ~A233 & A232;
  assign \new_[65027]_  = A235 & A234;
  assign \new_[65028]_  = \new_[65027]_  & \new_[65024]_ ;
  assign \new_[65031]_  = ~A266 & A265;
  assign \new_[65034]_  = A269 & A267;
  assign \new_[65035]_  = \new_[65034]_  & \new_[65031]_ ;
  assign \new_[65036]_  = \new_[65035]_  & \new_[65028]_ ;
  assign \new_[65040]_  = ~A168 & A169;
  assign \new_[65041]_  = A170 & \new_[65040]_ ;
  assign \new_[65044]_  = ~A200 & A199;
  assign \new_[65047]_  = A203 & A201;
  assign \new_[65048]_  = \new_[65047]_  & \new_[65044]_ ;
  assign \new_[65049]_  = \new_[65048]_  & \new_[65041]_ ;
  assign \new_[65052]_  = ~A233 & A232;
  assign \new_[65055]_  = A236 & A234;
  assign \new_[65056]_  = \new_[65055]_  & \new_[65052]_ ;
  assign \new_[65059]_  = ~A266 & A265;
  assign \new_[65062]_  = A268 & A267;
  assign \new_[65063]_  = \new_[65062]_  & \new_[65059]_ ;
  assign \new_[65064]_  = \new_[65063]_  & \new_[65056]_ ;
  assign \new_[65068]_  = ~A168 & A169;
  assign \new_[65069]_  = A170 & \new_[65068]_ ;
  assign \new_[65072]_  = ~A200 & A199;
  assign \new_[65075]_  = A203 & A201;
  assign \new_[65076]_  = \new_[65075]_  & \new_[65072]_ ;
  assign \new_[65077]_  = \new_[65076]_  & \new_[65069]_ ;
  assign \new_[65080]_  = ~A233 & A232;
  assign \new_[65083]_  = A236 & A234;
  assign \new_[65084]_  = \new_[65083]_  & \new_[65080]_ ;
  assign \new_[65087]_  = ~A266 & A265;
  assign \new_[65090]_  = A269 & A267;
  assign \new_[65091]_  = \new_[65090]_  & \new_[65087]_ ;
  assign \new_[65092]_  = \new_[65091]_  & \new_[65084]_ ;
  assign \new_[65096]_  = ~A168 & A169;
  assign \new_[65097]_  = A170 & \new_[65096]_ ;
  assign \new_[65100]_  = ~A200 & A199;
  assign \new_[65103]_  = A203 & A201;
  assign \new_[65104]_  = \new_[65103]_  & \new_[65100]_ ;
  assign \new_[65105]_  = \new_[65104]_  & \new_[65097]_ ;
  assign \new_[65108]_  = ~A233 & ~A232;
  assign \new_[65111]_  = A266 & A265;
  assign \new_[65112]_  = \new_[65111]_  & \new_[65108]_ ;
  assign \new_[65115]_  = ~A299 & A298;
  assign \new_[65118]_  = A301 & A300;
  assign \new_[65119]_  = \new_[65118]_  & \new_[65115]_ ;
  assign \new_[65120]_  = \new_[65119]_  & \new_[65112]_ ;
  assign \new_[65124]_  = ~A168 & A169;
  assign \new_[65125]_  = A170 & \new_[65124]_ ;
  assign \new_[65128]_  = ~A200 & A199;
  assign \new_[65131]_  = A203 & A201;
  assign \new_[65132]_  = \new_[65131]_  & \new_[65128]_ ;
  assign \new_[65133]_  = \new_[65132]_  & \new_[65125]_ ;
  assign \new_[65136]_  = ~A233 & ~A232;
  assign \new_[65139]_  = A266 & A265;
  assign \new_[65140]_  = \new_[65139]_  & \new_[65136]_ ;
  assign \new_[65143]_  = ~A299 & A298;
  assign \new_[65146]_  = A302 & A300;
  assign \new_[65147]_  = \new_[65146]_  & \new_[65143]_ ;
  assign \new_[65148]_  = \new_[65147]_  & \new_[65140]_ ;
  assign \new_[65152]_  = A167 & A169;
  assign \new_[65153]_  = ~A170 & \new_[65152]_ ;
  assign \new_[65156]_  = A199 & A166;
  assign \new_[65159]_  = A232 & A200;
  assign \new_[65160]_  = \new_[65159]_  & \new_[65156]_ ;
  assign \new_[65161]_  = \new_[65160]_  & \new_[65153]_ ;
  assign \new_[65164]_  = A265 & A233;
  assign \new_[65167]_  = ~A269 & ~A268;
  assign \new_[65168]_  = \new_[65167]_  & \new_[65164]_ ;
  assign \new_[65171]_  = ~A299 & A298;
  assign \new_[65174]_  = A301 & A300;
  assign \new_[65175]_  = \new_[65174]_  & \new_[65171]_ ;
  assign \new_[65176]_  = \new_[65175]_  & \new_[65168]_ ;
  assign \new_[65180]_  = A167 & A169;
  assign \new_[65181]_  = ~A170 & \new_[65180]_ ;
  assign \new_[65184]_  = A199 & A166;
  assign \new_[65187]_  = A232 & A200;
  assign \new_[65188]_  = \new_[65187]_  & \new_[65184]_ ;
  assign \new_[65189]_  = \new_[65188]_  & \new_[65181]_ ;
  assign \new_[65192]_  = A265 & A233;
  assign \new_[65195]_  = ~A269 & ~A268;
  assign \new_[65196]_  = \new_[65195]_  & \new_[65192]_ ;
  assign \new_[65199]_  = ~A299 & A298;
  assign \new_[65202]_  = A302 & A300;
  assign \new_[65203]_  = \new_[65202]_  & \new_[65199]_ ;
  assign \new_[65204]_  = \new_[65203]_  & \new_[65196]_ ;
  assign \new_[65208]_  = A167 & A169;
  assign \new_[65209]_  = ~A170 & \new_[65208]_ ;
  assign \new_[65212]_  = A199 & A166;
  assign \new_[65215]_  = ~A233 & A200;
  assign \new_[65216]_  = \new_[65215]_  & \new_[65212]_ ;
  assign \new_[65217]_  = \new_[65216]_  & \new_[65209]_ ;
  assign \new_[65220]_  = ~A236 & ~A235;
  assign \new_[65223]_  = A266 & A265;
  assign \new_[65224]_  = \new_[65223]_  & \new_[65220]_ ;
  assign \new_[65227]_  = ~A299 & A298;
  assign \new_[65230]_  = A301 & A300;
  assign \new_[65231]_  = \new_[65230]_  & \new_[65227]_ ;
  assign \new_[65232]_  = \new_[65231]_  & \new_[65224]_ ;
  assign \new_[65236]_  = A167 & A169;
  assign \new_[65237]_  = ~A170 & \new_[65236]_ ;
  assign \new_[65240]_  = A199 & A166;
  assign \new_[65243]_  = ~A233 & A200;
  assign \new_[65244]_  = \new_[65243]_  & \new_[65240]_ ;
  assign \new_[65245]_  = \new_[65244]_  & \new_[65237]_ ;
  assign \new_[65248]_  = ~A236 & ~A235;
  assign \new_[65251]_  = A266 & A265;
  assign \new_[65252]_  = \new_[65251]_  & \new_[65248]_ ;
  assign \new_[65255]_  = ~A299 & A298;
  assign \new_[65258]_  = A302 & A300;
  assign \new_[65259]_  = \new_[65258]_  & \new_[65255]_ ;
  assign \new_[65260]_  = \new_[65259]_  & \new_[65252]_ ;
  assign \new_[65264]_  = A167 & A169;
  assign \new_[65265]_  = ~A170 & \new_[65264]_ ;
  assign \new_[65268]_  = A199 & A166;
  assign \new_[65271]_  = ~A233 & A200;
  assign \new_[65272]_  = \new_[65271]_  & \new_[65268]_ ;
  assign \new_[65273]_  = \new_[65272]_  & \new_[65265]_ ;
  assign \new_[65276]_  = ~A236 & ~A235;
  assign \new_[65279]_  = ~A267 & ~A266;
  assign \new_[65280]_  = \new_[65279]_  & \new_[65276]_ ;
  assign \new_[65283]_  = ~A299 & A298;
  assign \new_[65286]_  = A301 & A300;
  assign \new_[65287]_  = \new_[65286]_  & \new_[65283]_ ;
  assign \new_[65288]_  = \new_[65287]_  & \new_[65280]_ ;
  assign \new_[65292]_  = A167 & A169;
  assign \new_[65293]_  = ~A170 & \new_[65292]_ ;
  assign \new_[65296]_  = A199 & A166;
  assign \new_[65299]_  = ~A233 & A200;
  assign \new_[65300]_  = \new_[65299]_  & \new_[65296]_ ;
  assign \new_[65301]_  = \new_[65300]_  & \new_[65293]_ ;
  assign \new_[65304]_  = ~A236 & ~A235;
  assign \new_[65307]_  = ~A267 & ~A266;
  assign \new_[65308]_  = \new_[65307]_  & \new_[65304]_ ;
  assign \new_[65311]_  = ~A299 & A298;
  assign \new_[65314]_  = A302 & A300;
  assign \new_[65315]_  = \new_[65314]_  & \new_[65311]_ ;
  assign \new_[65316]_  = \new_[65315]_  & \new_[65308]_ ;
  assign \new_[65320]_  = A167 & A169;
  assign \new_[65321]_  = ~A170 & \new_[65320]_ ;
  assign \new_[65324]_  = A199 & A166;
  assign \new_[65327]_  = ~A233 & A200;
  assign \new_[65328]_  = \new_[65327]_  & \new_[65324]_ ;
  assign \new_[65329]_  = \new_[65328]_  & \new_[65321]_ ;
  assign \new_[65332]_  = ~A236 & ~A235;
  assign \new_[65335]_  = ~A266 & ~A265;
  assign \new_[65336]_  = \new_[65335]_  & \new_[65332]_ ;
  assign \new_[65339]_  = ~A299 & A298;
  assign \new_[65342]_  = A301 & A300;
  assign \new_[65343]_  = \new_[65342]_  & \new_[65339]_ ;
  assign \new_[65344]_  = \new_[65343]_  & \new_[65336]_ ;
  assign \new_[65348]_  = A167 & A169;
  assign \new_[65349]_  = ~A170 & \new_[65348]_ ;
  assign \new_[65352]_  = A199 & A166;
  assign \new_[65355]_  = ~A233 & A200;
  assign \new_[65356]_  = \new_[65355]_  & \new_[65352]_ ;
  assign \new_[65357]_  = \new_[65356]_  & \new_[65349]_ ;
  assign \new_[65360]_  = ~A236 & ~A235;
  assign \new_[65363]_  = ~A266 & ~A265;
  assign \new_[65364]_  = \new_[65363]_  & \new_[65360]_ ;
  assign \new_[65367]_  = ~A299 & A298;
  assign \new_[65370]_  = A302 & A300;
  assign \new_[65371]_  = \new_[65370]_  & \new_[65367]_ ;
  assign \new_[65372]_  = \new_[65371]_  & \new_[65364]_ ;
  assign \new_[65376]_  = A167 & A169;
  assign \new_[65377]_  = ~A170 & \new_[65376]_ ;
  assign \new_[65380]_  = A199 & A166;
  assign \new_[65383]_  = ~A233 & A200;
  assign \new_[65384]_  = \new_[65383]_  & \new_[65380]_ ;
  assign \new_[65385]_  = \new_[65384]_  & \new_[65377]_ ;
  assign \new_[65388]_  = ~A266 & ~A234;
  assign \new_[65391]_  = ~A269 & ~A268;
  assign \new_[65392]_  = \new_[65391]_  & \new_[65388]_ ;
  assign \new_[65395]_  = ~A299 & A298;
  assign \new_[65398]_  = A301 & A300;
  assign \new_[65399]_  = \new_[65398]_  & \new_[65395]_ ;
  assign \new_[65400]_  = \new_[65399]_  & \new_[65392]_ ;
  assign \new_[65404]_  = A167 & A169;
  assign \new_[65405]_  = ~A170 & \new_[65404]_ ;
  assign \new_[65408]_  = A199 & A166;
  assign \new_[65411]_  = ~A233 & A200;
  assign \new_[65412]_  = \new_[65411]_  & \new_[65408]_ ;
  assign \new_[65413]_  = \new_[65412]_  & \new_[65405]_ ;
  assign \new_[65416]_  = ~A266 & ~A234;
  assign \new_[65419]_  = ~A269 & ~A268;
  assign \new_[65420]_  = \new_[65419]_  & \new_[65416]_ ;
  assign \new_[65423]_  = ~A299 & A298;
  assign \new_[65426]_  = A302 & A300;
  assign \new_[65427]_  = \new_[65426]_  & \new_[65423]_ ;
  assign \new_[65428]_  = \new_[65427]_  & \new_[65420]_ ;
  assign \new_[65432]_  = A167 & A169;
  assign \new_[65433]_  = ~A170 & \new_[65432]_ ;
  assign \new_[65436]_  = A199 & A166;
  assign \new_[65439]_  = ~A232 & A200;
  assign \new_[65440]_  = \new_[65439]_  & \new_[65436]_ ;
  assign \new_[65441]_  = \new_[65440]_  & \new_[65433]_ ;
  assign \new_[65444]_  = ~A266 & ~A233;
  assign \new_[65447]_  = ~A269 & ~A268;
  assign \new_[65448]_  = \new_[65447]_  & \new_[65444]_ ;
  assign \new_[65451]_  = ~A299 & A298;
  assign \new_[65454]_  = A301 & A300;
  assign \new_[65455]_  = \new_[65454]_  & \new_[65451]_ ;
  assign \new_[65456]_  = \new_[65455]_  & \new_[65448]_ ;
  assign \new_[65460]_  = A167 & A169;
  assign \new_[65461]_  = ~A170 & \new_[65460]_ ;
  assign \new_[65464]_  = A199 & A166;
  assign \new_[65467]_  = ~A232 & A200;
  assign \new_[65468]_  = \new_[65467]_  & \new_[65464]_ ;
  assign \new_[65469]_  = \new_[65468]_  & \new_[65461]_ ;
  assign \new_[65472]_  = ~A266 & ~A233;
  assign \new_[65475]_  = ~A269 & ~A268;
  assign \new_[65476]_  = \new_[65475]_  & \new_[65472]_ ;
  assign \new_[65479]_  = ~A299 & A298;
  assign \new_[65482]_  = A302 & A300;
  assign \new_[65483]_  = \new_[65482]_  & \new_[65479]_ ;
  assign \new_[65484]_  = \new_[65483]_  & \new_[65476]_ ;
  assign \new_[65488]_  = A167 & A169;
  assign \new_[65489]_  = ~A170 & \new_[65488]_ ;
  assign \new_[65492]_  = ~A200 & A166;
  assign \new_[65495]_  = ~A203 & ~A202;
  assign \new_[65496]_  = \new_[65495]_  & \new_[65492]_ ;
  assign \new_[65497]_  = \new_[65496]_  & \new_[65489]_ ;
  assign \new_[65500]_  = A233 & A232;
  assign \new_[65503]_  = ~A267 & A265;
  assign \new_[65504]_  = \new_[65503]_  & \new_[65500]_ ;
  assign \new_[65507]_  = ~A299 & A298;
  assign \new_[65510]_  = A301 & A300;
  assign \new_[65511]_  = \new_[65510]_  & \new_[65507]_ ;
  assign \new_[65512]_  = \new_[65511]_  & \new_[65504]_ ;
  assign \new_[65516]_  = A167 & A169;
  assign \new_[65517]_  = ~A170 & \new_[65516]_ ;
  assign \new_[65520]_  = ~A200 & A166;
  assign \new_[65523]_  = ~A203 & ~A202;
  assign \new_[65524]_  = \new_[65523]_  & \new_[65520]_ ;
  assign \new_[65525]_  = \new_[65524]_  & \new_[65517]_ ;
  assign \new_[65528]_  = A233 & A232;
  assign \new_[65531]_  = ~A267 & A265;
  assign \new_[65532]_  = \new_[65531]_  & \new_[65528]_ ;
  assign \new_[65535]_  = ~A299 & A298;
  assign \new_[65538]_  = A302 & A300;
  assign \new_[65539]_  = \new_[65538]_  & \new_[65535]_ ;
  assign \new_[65540]_  = \new_[65539]_  & \new_[65532]_ ;
  assign \new_[65544]_  = A167 & A169;
  assign \new_[65545]_  = ~A170 & \new_[65544]_ ;
  assign \new_[65548]_  = ~A200 & A166;
  assign \new_[65551]_  = ~A203 & ~A202;
  assign \new_[65552]_  = \new_[65551]_  & \new_[65548]_ ;
  assign \new_[65553]_  = \new_[65552]_  & \new_[65545]_ ;
  assign \new_[65556]_  = A233 & A232;
  assign \new_[65559]_  = A266 & A265;
  assign \new_[65560]_  = \new_[65559]_  & \new_[65556]_ ;
  assign \new_[65563]_  = ~A299 & A298;
  assign \new_[65566]_  = A301 & A300;
  assign \new_[65567]_  = \new_[65566]_  & \new_[65563]_ ;
  assign \new_[65568]_  = \new_[65567]_  & \new_[65560]_ ;
  assign \new_[65572]_  = A167 & A169;
  assign \new_[65573]_  = ~A170 & \new_[65572]_ ;
  assign \new_[65576]_  = ~A200 & A166;
  assign \new_[65579]_  = ~A203 & ~A202;
  assign \new_[65580]_  = \new_[65579]_  & \new_[65576]_ ;
  assign \new_[65581]_  = \new_[65580]_  & \new_[65573]_ ;
  assign \new_[65584]_  = A233 & A232;
  assign \new_[65587]_  = A266 & A265;
  assign \new_[65588]_  = \new_[65587]_  & \new_[65584]_ ;
  assign \new_[65591]_  = ~A299 & A298;
  assign \new_[65594]_  = A302 & A300;
  assign \new_[65595]_  = \new_[65594]_  & \new_[65591]_ ;
  assign \new_[65596]_  = \new_[65595]_  & \new_[65588]_ ;
  assign \new_[65600]_  = A167 & A169;
  assign \new_[65601]_  = ~A170 & \new_[65600]_ ;
  assign \new_[65604]_  = ~A200 & A166;
  assign \new_[65607]_  = ~A203 & ~A202;
  assign \new_[65608]_  = \new_[65607]_  & \new_[65604]_ ;
  assign \new_[65609]_  = \new_[65608]_  & \new_[65601]_ ;
  assign \new_[65612]_  = A233 & A232;
  assign \new_[65615]_  = ~A266 & ~A265;
  assign \new_[65616]_  = \new_[65615]_  & \new_[65612]_ ;
  assign \new_[65619]_  = ~A299 & A298;
  assign \new_[65622]_  = A301 & A300;
  assign \new_[65623]_  = \new_[65622]_  & \new_[65619]_ ;
  assign \new_[65624]_  = \new_[65623]_  & \new_[65616]_ ;
  assign \new_[65628]_  = A167 & A169;
  assign \new_[65629]_  = ~A170 & \new_[65628]_ ;
  assign \new_[65632]_  = ~A200 & A166;
  assign \new_[65635]_  = ~A203 & ~A202;
  assign \new_[65636]_  = \new_[65635]_  & \new_[65632]_ ;
  assign \new_[65637]_  = \new_[65636]_  & \new_[65629]_ ;
  assign \new_[65640]_  = A233 & A232;
  assign \new_[65643]_  = ~A266 & ~A265;
  assign \new_[65644]_  = \new_[65643]_  & \new_[65640]_ ;
  assign \new_[65647]_  = ~A299 & A298;
  assign \new_[65650]_  = A302 & A300;
  assign \new_[65651]_  = \new_[65650]_  & \new_[65647]_ ;
  assign \new_[65652]_  = \new_[65651]_  & \new_[65644]_ ;
  assign \new_[65656]_  = A167 & A169;
  assign \new_[65657]_  = ~A170 & \new_[65656]_ ;
  assign \new_[65660]_  = ~A200 & A166;
  assign \new_[65663]_  = ~A203 & ~A202;
  assign \new_[65664]_  = \new_[65663]_  & \new_[65660]_ ;
  assign \new_[65665]_  = \new_[65664]_  & \new_[65657]_ ;
  assign \new_[65668]_  = ~A235 & ~A233;
  assign \new_[65671]_  = ~A266 & ~A236;
  assign \new_[65672]_  = \new_[65671]_  & \new_[65668]_ ;
  assign \new_[65675]_  = ~A269 & ~A268;
  assign \new_[65678]_  = A299 & ~A298;
  assign \new_[65679]_  = \new_[65678]_  & \new_[65675]_ ;
  assign \new_[65680]_  = \new_[65679]_  & \new_[65672]_ ;
  assign \new_[65684]_  = A167 & A169;
  assign \new_[65685]_  = ~A170 & \new_[65684]_ ;
  assign \new_[65688]_  = ~A200 & A166;
  assign \new_[65691]_  = ~A203 & ~A202;
  assign \new_[65692]_  = \new_[65691]_  & \new_[65688]_ ;
  assign \new_[65693]_  = \new_[65692]_  & \new_[65685]_ ;
  assign \new_[65696]_  = ~A234 & ~A233;
  assign \new_[65699]_  = A266 & A265;
  assign \new_[65700]_  = \new_[65699]_  & \new_[65696]_ ;
  assign \new_[65703]_  = ~A299 & A298;
  assign \new_[65706]_  = A301 & A300;
  assign \new_[65707]_  = \new_[65706]_  & \new_[65703]_ ;
  assign \new_[65708]_  = \new_[65707]_  & \new_[65700]_ ;
  assign \new_[65712]_  = A167 & A169;
  assign \new_[65713]_  = ~A170 & \new_[65712]_ ;
  assign \new_[65716]_  = ~A200 & A166;
  assign \new_[65719]_  = ~A203 & ~A202;
  assign \new_[65720]_  = \new_[65719]_  & \new_[65716]_ ;
  assign \new_[65721]_  = \new_[65720]_  & \new_[65713]_ ;
  assign \new_[65724]_  = ~A234 & ~A233;
  assign \new_[65727]_  = A266 & A265;
  assign \new_[65728]_  = \new_[65727]_  & \new_[65724]_ ;
  assign \new_[65731]_  = ~A299 & A298;
  assign \new_[65734]_  = A302 & A300;
  assign \new_[65735]_  = \new_[65734]_  & \new_[65731]_ ;
  assign \new_[65736]_  = \new_[65735]_  & \new_[65728]_ ;
  assign \new_[65740]_  = A167 & A169;
  assign \new_[65741]_  = ~A170 & \new_[65740]_ ;
  assign \new_[65744]_  = ~A200 & A166;
  assign \new_[65747]_  = ~A203 & ~A202;
  assign \new_[65748]_  = \new_[65747]_  & \new_[65744]_ ;
  assign \new_[65749]_  = \new_[65748]_  & \new_[65741]_ ;
  assign \new_[65752]_  = ~A234 & ~A233;
  assign \new_[65755]_  = ~A267 & ~A266;
  assign \new_[65756]_  = \new_[65755]_  & \new_[65752]_ ;
  assign \new_[65759]_  = ~A299 & A298;
  assign \new_[65762]_  = A301 & A300;
  assign \new_[65763]_  = \new_[65762]_  & \new_[65759]_ ;
  assign \new_[65764]_  = \new_[65763]_  & \new_[65756]_ ;
  assign \new_[65768]_  = A167 & A169;
  assign \new_[65769]_  = ~A170 & \new_[65768]_ ;
  assign \new_[65772]_  = ~A200 & A166;
  assign \new_[65775]_  = ~A203 & ~A202;
  assign \new_[65776]_  = \new_[65775]_  & \new_[65772]_ ;
  assign \new_[65777]_  = \new_[65776]_  & \new_[65769]_ ;
  assign \new_[65780]_  = ~A234 & ~A233;
  assign \new_[65783]_  = ~A267 & ~A266;
  assign \new_[65784]_  = \new_[65783]_  & \new_[65780]_ ;
  assign \new_[65787]_  = ~A299 & A298;
  assign \new_[65790]_  = A302 & A300;
  assign \new_[65791]_  = \new_[65790]_  & \new_[65787]_ ;
  assign \new_[65792]_  = \new_[65791]_  & \new_[65784]_ ;
  assign \new_[65796]_  = A167 & A169;
  assign \new_[65797]_  = ~A170 & \new_[65796]_ ;
  assign \new_[65800]_  = ~A200 & A166;
  assign \new_[65803]_  = ~A203 & ~A202;
  assign \new_[65804]_  = \new_[65803]_  & \new_[65800]_ ;
  assign \new_[65805]_  = \new_[65804]_  & \new_[65797]_ ;
  assign \new_[65808]_  = ~A234 & ~A233;
  assign \new_[65811]_  = ~A266 & ~A265;
  assign \new_[65812]_  = \new_[65811]_  & \new_[65808]_ ;
  assign \new_[65815]_  = ~A299 & A298;
  assign \new_[65818]_  = A301 & A300;
  assign \new_[65819]_  = \new_[65818]_  & \new_[65815]_ ;
  assign \new_[65820]_  = \new_[65819]_  & \new_[65812]_ ;
  assign \new_[65824]_  = A167 & A169;
  assign \new_[65825]_  = ~A170 & \new_[65824]_ ;
  assign \new_[65828]_  = ~A200 & A166;
  assign \new_[65831]_  = ~A203 & ~A202;
  assign \new_[65832]_  = \new_[65831]_  & \new_[65828]_ ;
  assign \new_[65833]_  = \new_[65832]_  & \new_[65825]_ ;
  assign \new_[65836]_  = ~A234 & ~A233;
  assign \new_[65839]_  = ~A266 & ~A265;
  assign \new_[65840]_  = \new_[65839]_  & \new_[65836]_ ;
  assign \new_[65843]_  = ~A299 & A298;
  assign \new_[65846]_  = A302 & A300;
  assign \new_[65847]_  = \new_[65846]_  & \new_[65843]_ ;
  assign \new_[65848]_  = \new_[65847]_  & \new_[65840]_ ;
  assign \new_[65852]_  = A167 & A169;
  assign \new_[65853]_  = ~A170 & \new_[65852]_ ;
  assign \new_[65856]_  = ~A200 & A166;
  assign \new_[65859]_  = ~A203 & ~A202;
  assign \new_[65860]_  = \new_[65859]_  & \new_[65856]_ ;
  assign \new_[65861]_  = \new_[65860]_  & \new_[65853]_ ;
  assign \new_[65864]_  = ~A233 & A232;
  assign \new_[65867]_  = A235 & A234;
  assign \new_[65868]_  = \new_[65867]_  & \new_[65864]_ ;
  assign \new_[65871]_  = ~A266 & A265;
  assign \new_[65874]_  = A268 & A267;
  assign \new_[65875]_  = \new_[65874]_  & \new_[65871]_ ;
  assign \new_[65876]_  = \new_[65875]_  & \new_[65868]_ ;
  assign \new_[65880]_  = A167 & A169;
  assign \new_[65881]_  = ~A170 & \new_[65880]_ ;
  assign \new_[65884]_  = ~A200 & A166;
  assign \new_[65887]_  = ~A203 & ~A202;
  assign \new_[65888]_  = \new_[65887]_  & \new_[65884]_ ;
  assign \new_[65889]_  = \new_[65888]_  & \new_[65881]_ ;
  assign \new_[65892]_  = ~A233 & A232;
  assign \new_[65895]_  = A235 & A234;
  assign \new_[65896]_  = \new_[65895]_  & \new_[65892]_ ;
  assign \new_[65899]_  = ~A266 & A265;
  assign \new_[65902]_  = A269 & A267;
  assign \new_[65903]_  = \new_[65902]_  & \new_[65899]_ ;
  assign \new_[65904]_  = \new_[65903]_  & \new_[65896]_ ;
  assign \new_[65908]_  = A167 & A169;
  assign \new_[65909]_  = ~A170 & \new_[65908]_ ;
  assign \new_[65912]_  = ~A200 & A166;
  assign \new_[65915]_  = ~A203 & ~A202;
  assign \new_[65916]_  = \new_[65915]_  & \new_[65912]_ ;
  assign \new_[65917]_  = \new_[65916]_  & \new_[65909]_ ;
  assign \new_[65920]_  = ~A233 & A232;
  assign \new_[65923]_  = A236 & A234;
  assign \new_[65924]_  = \new_[65923]_  & \new_[65920]_ ;
  assign \new_[65927]_  = ~A266 & A265;
  assign \new_[65930]_  = A268 & A267;
  assign \new_[65931]_  = \new_[65930]_  & \new_[65927]_ ;
  assign \new_[65932]_  = \new_[65931]_  & \new_[65924]_ ;
  assign \new_[65936]_  = A167 & A169;
  assign \new_[65937]_  = ~A170 & \new_[65936]_ ;
  assign \new_[65940]_  = ~A200 & A166;
  assign \new_[65943]_  = ~A203 & ~A202;
  assign \new_[65944]_  = \new_[65943]_  & \new_[65940]_ ;
  assign \new_[65945]_  = \new_[65944]_  & \new_[65937]_ ;
  assign \new_[65948]_  = ~A233 & A232;
  assign \new_[65951]_  = A236 & A234;
  assign \new_[65952]_  = \new_[65951]_  & \new_[65948]_ ;
  assign \new_[65955]_  = ~A266 & A265;
  assign \new_[65958]_  = A269 & A267;
  assign \new_[65959]_  = \new_[65958]_  & \new_[65955]_ ;
  assign \new_[65960]_  = \new_[65959]_  & \new_[65952]_ ;
  assign \new_[65964]_  = A167 & A169;
  assign \new_[65965]_  = ~A170 & \new_[65964]_ ;
  assign \new_[65968]_  = ~A200 & A166;
  assign \new_[65971]_  = ~A203 & ~A202;
  assign \new_[65972]_  = \new_[65971]_  & \new_[65968]_ ;
  assign \new_[65973]_  = \new_[65972]_  & \new_[65965]_ ;
  assign \new_[65976]_  = ~A233 & ~A232;
  assign \new_[65979]_  = A266 & A265;
  assign \new_[65980]_  = \new_[65979]_  & \new_[65976]_ ;
  assign \new_[65983]_  = ~A299 & A298;
  assign \new_[65986]_  = A301 & A300;
  assign \new_[65987]_  = \new_[65986]_  & \new_[65983]_ ;
  assign \new_[65988]_  = \new_[65987]_  & \new_[65980]_ ;
  assign \new_[65992]_  = A167 & A169;
  assign \new_[65993]_  = ~A170 & \new_[65992]_ ;
  assign \new_[65996]_  = ~A200 & A166;
  assign \new_[65999]_  = ~A203 & ~A202;
  assign \new_[66000]_  = \new_[65999]_  & \new_[65996]_ ;
  assign \new_[66001]_  = \new_[66000]_  & \new_[65993]_ ;
  assign \new_[66004]_  = ~A233 & ~A232;
  assign \new_[66007]_  = A266 & A265;
  assign \new_[66008]_  = \new_[66007]_  & \new_[66004]_ ;
  assign \new_[66011]_  = ~A299 & A298;
  assign \new_[66014]_  = A302 & A300;
  assign \new_[66015]_  = \new_[66014]_  & \new_[66011]_ ;
  assign \new_[66016]_  = \new_[66015]_  & \new_[66008]_ ;
  assign \new_[66020]_  = A167 & A169;
  assign \new_[66021]_  = ~A170 & \new_[66020]_ ;
  assign \new_[66024]_  = ~A200 & A166;
  assign \new_[66027]_  = ~A203 & ~A202;
  assign \new_[66028]_  = \new_[66027]_  & \new_[66024]_ ;
  assign \new_[66029]_  = \new_[66028]_  & \new_[66021]_ ;
  assign \new_[66032]_  = ~A233 & ~A232;
  assign \new_[66035]_  = ~A267 & ~A266;
  assign \new_[66036]_  = \new_[66035]_  & \new_[66032]_ ;
  assign \new_[66039]_  = ~A299 & A298;
  assign \new_[66042]_  = A301 & A300;
  assign \new_[66043]_  = \new_[66042]_  & \new_[66039]_ ;
  assign \new_[66044]_  = \new_[66043]_  & \new_[66036]_ ;
  assign \new_[66048]_  = A167 & A169;
  assign \new_[66049]_  = ~A170 & \new_[66048]_ ;
  assign \new_[66052]_  = ~A200 & A166;
  assign \new_[66055]_  = ~A203 & ~A202;
  assign \new_[66056]_  = \new_[66055]_  & \new_[66052]_ ;
  assign \new_[66057]_  = \new_[66056]_  & \new_[66049]_ ;
  assign \new_[66060]_  = ~A233 & ~A232;
  assign \new_[66063]_  = ~A267 & ~A266;
  assign \new_[66064]_  = \new_[66063]_  & \new_[66060]_ ;
  assign \new_[66067]_  = ~A299 & A298;
  assign \new_[66070]_  = A302 & A300;
  assign \new_[66071]_  = \new_[66070]_  & \new_[66067]_ ;
  assign \new_[66072]_  = \new_[66071]_  & \new_[66064]_ ;
  assign \new_[66076]_  = A167 & A169;
  assign \new_[66077]_  = ~A170 & \new_[66076]_ ;
  assign \new_[66080]_  = ~A200 & A166;
  assign \new_[66083]_  = ~A203 & ~A202;
  assign \new_[66084]_  = \new_[66083]_  & \new_[66080]_ ;
  assign \new_[66085]_  = \new_[66084]_  & \new_[66077]_ ;
  assign \new_[66088]_  = ~A233 & ~A232;
  assign \new_[66091]_  = ~A266 & ~A265;
  assign \new_[66092]_  = \new_[66091]_  & \new_[66088]_ ;
  assign \new_[66095]_  = ~A299 & A298;
  assign \new_[66098]_  = A301 & A300;
  assign \new_[66099]_  = \new_[66098]_  & \new_[66095]_ ;
  assign \new_[66100]_  = \new_[66099]_  & \new_[66092]_ ;
  assign \new_[66104]_  = A167 & A169;
  assign \new_[66105]_  = ~A170 & \new_[66104]_ ;
  assign \new_[66108]_  = ~A200 & A166;
  assign \new_[66111]_  = ~A203 & ~A202;
  assign \new_[66112]_  = \new_[66111]_  & \new_[66108]_ ;
  assign \new_[66113]_  = \new_[66112]_  & \new_[66105]_ ;
  assign \new_[66116]_  = ~A233 & ~A232;
  assign \new_[66119]_  = ~A266 & ~A265;
  assign \new_[66120]_  = \new_[66119]_  & \new_[66116]_ ;
  assign \new_[66123]_  = ~A299 & A298;
  assign \new_[66126]_  = A302 & A300;
  assign \new_[66127]_  = \new_[66126]_  & \new_[66123]_ ;
  assign \new_[66128]_  = \new_[66127]_  & \new_[66120]_ ;
  assign \new_[66132]_  = A167 & A169;
  assign \new_[66133]_  = ~A170 & \new_[66132]_ ;
  assign \new_[66136]_  = ~A200 & A166;
  assign \new_[66139]_  = A232 & ~A201;
  assign \new_[66140]_  = \new_[66139]_  & \new_[66136]_ ;
  assign \new_[66141]_  = \new_[66140]_  & \new_[66133]_ ;
  assign \new_[66144]_  = A265 & A233;
  assign \new_[66147]_  = ~A269 & ~A268;
  assign \new_[66148]_  = \new_[66147]_  & \new_[66144]_ ;
  assign \new_[66151]_  = ~A299 & A298;
  assign \new_[66154]_  = A301 & A300;
  assign \new_[66155]_  = \new_[66154]_  & \new_[66151]_ ;
  assign \new_[66156]_  = \new_[66155]_  & \new_[66148]_ ;
  assign \new_[66160]_  = A167 & A169;
  assign \new_[66161]_  = ~A170 & \new_[66160]_ ;
  assign \new_[66164]_  = ~A200 & A166;
  assign \new_[66167]_  = A232 & ~A201;
  assign \new_[66168]_  = \new_[66167]_  & \new_[66164]_ ;
  assign \new_[66169]_  = \new_[66168]_  & \new_[66161]_ ;
  assign \new_[66172]_  = A265 & A233;
  assign \new_[66175]_  = ~A269 & ~A268;
  assign \new_[66176]_  = \new_[66175]_  & \new_[66172]_ ;
  assign \new_[66179]_  = ~A299 & A298;
  assign \new_[66182]_  = A302 & A300;
  assign \new_[66183]_  = \new_[66182]_  & \new_[66179]_ ;
  assign \new_[66184]_  = \new_[66183]_  & \new_[66176]_ ;
  assign \new_[66188]_  = A167 & A169;
  assign \new_[66189]_  = ~A170 & \new_[66188]_ ;
  assign \new_[66192]_  = ~A200 & A166;
  assign \new_[66195]_  = ~A233 & ~A201;
  assign \new_[66196]_  = \new_[66195]_  & \new_[66192]_ ;
  assign \new_[66197]_  = \new_[66196]_  & \new_[66189]_ ;
  assign \new_[66200]_  = ~A236 & ~A235;
  assign \new_[66203]_  = A266 & A265;
  assign \new_[66204]_  = \new_[66203]_  & \new_[66200]_ ;
  assign \new_[66207]_  = ~A299 & A298;
  assign \new_[66210]_  = A301 & A300;
  assign \new_[66211]_  = \new_[66210]_  & \new_[66207]_ ;
  assign \new_[66212]_  = \new_[66211]_  & \new_[66204]_ ;
  assign \new_[66216]_  = A167 & A169;
  assign \new_[66217]_  = ~A170 & \new_[66216]_ ;
  assign \new_[66220]_  = ~A200 & A166;
  assign \new_[66223]_  = ~A233 & ~A201;
  assign \new_[66224]_  = \new_[66223]_  & \new_[66220]_ ;
  assign \new_[66225]_  = \new_[66224]_  & \new_[66217]_ ;
  assign \new_[66228]_  = ~A236 & ~A235;
  assign \new_[66231]_  = A266 & A265;
  assign \new_[66232]_  = \new_[66231]_  & \new_[66228]_ ;
  assign \new_[66235]_  = ~A299 & A298;
  assign \new_[66238]_  = A302 & A300;
  assign \new_[66239]_  = \new_[66238]_  & \new_[66235]_ ;
  assign \new_[66240]_  = \new_[66239]_  & \new_[66232]_ ;
  assign \new_[66244]_  = A167 & A169;
  assign \new_[66245]_  = ~A170 & \new_[66244]_ ;
  assign \new_[66248]_  = ~A200 & A166;
  assign \new_[66251]_  = ~A233 & ~A201;
  assign \new_[66252]_  = \new_[66251]_  & \new_[66248]_ ;
  assign \new_[66253]_  = \new_[66252]_  & \new_[66245]_ ;
  assign \new_[66256]_  = ~A236 & ~A235;
  assign \new_[66259]_  = ~A267 & ~A266;
  assign \new_[66260]_  = \new_[66259]_  & \new_[66256]_ ;
  assign \new_[66263]_  = ~A299 & A298;
  assign \new_[66266]_  = A301 & A300;
  assign \new_[66267]_  = \new_[66266]_  & \new_[66263]_ ;
  assign \new_[66268]_  = \new_[66267]_  & \new_[66260]_ ;
  assign \new_[66272]_  = A167 & A169;
  assign \new_[66273]_  = ~A170 & \new_[66272]_ ;
  assign \new_[66276]_  = ~A200 & A166;
  assign \new_[66279]_  = ~A233 & ~A201;
  assign \new_[66280]_  = \new_[66279]_  & \new_[66276]_ ;
  assign \new_[66281]_  = \new_[66280]_  & \new_[66273]_ ;
  assign \new_[66284]_  = ~A236 & ~A235;
  assign \new_[66287]_  = ~A267 & ~A266;
  assign \new_[66288]_  = \new_[66287]_  & \new_[66284]_ ;
  assign \new_[66291]_  = ~A299 & A298;
  assign \new_[66294]_  = A302 & A300;
  assign \new_[66295]_  = \new_[66294]_  & \new_[66291]_ ;
  assign \new_[66296]_  = \new_[66295]_  & \new_[66288]_ ;
  assign \new_[66300]_  = A167 & A169;
  assign \new_[66301]_  = ~A170 & \new_[66300]_ ;
  assign \new_[66304]_  = ~A200 & A166;
  assign \new_[66307]_  = ~A233 & ~A201;
  assign \new_[66308]_  = \new_[66307]_  & \new_[66304]_ ;
  assign \new_[66309]_  = \new_[66308]_  & \new_[66301]_ ;
  assign \new_[66312]_  = ~A236 & ~A235;
  assign \new_[66315]_  = ~A266 & ~A265;
  assign \new_[66316]_  = \new_[66315]_  & \new_[66312]_ ;
  assign \new_[66319]_  = ~A299 & A298;
  assign \new_[66322]_  = A301 & A300;
  assign \new_[66323]_  = \new_[66322]_  & \new_[66319]_ ;
  assign \new_[66324]_  = \new_[66323]_  & \new_[66316]_ ;
  assign \new_[66328]_  = A167 & A169;
  assign \new_[66329]_  = ~A170 & \new_[66328]_ ;
  assign \new_[66332]_  = ~A200 & A166;
  assign \new_[66335]_  = ~A233 & ~A201;
  assign \new_[66336]_  = \new_[66335]_  & \new_[66332]_ ;
  assign \new_[66337]_  = \new_[66336]_  & \new_[66329]_ ;
  assign \new_[66340]_  = ~A236 & ~A235;
  assign \new_[66343]_  = ~A266 & ~A265;
  assign \new_[66344]_  = \new_[66343]_  & \new_[66340]_ ;
  assign \new_[66347]_  = ~A299 & A298;
  assign \new_[66350]_  = A302 & A300;
  assign \new_[66351]_  = \new_[66350]_  & \new_[66347]_ ;
  assign \new_[66352]_  = \new_[66351]_  & \new_[66344]_ ;
  assign \new_[66356]_  = A167 & A169;
  assign \new_[66357]_  = ~A170 & \new_[66356]_ ;
  assign \new_[66360]_  = ~A200 & A166;
  assign \new_[66363]_  = ~A233 & ~A201;
  assign \new_[66364]_  = \new_[66363]_  & \new_[66360]_ ;
  assign \new_[66365]_  = \new_[66364]_  & \new_[66357]_ ;
  assign \new_[66368]_  = ~A266 & ~A234;
  assign \new_[66371]_  = ~A269 & ~A268;
  assign \new_[66372]_  = \new_[66371]_  & \new_[66368]_ ;
  assign \new_[66375]_  = ~A299 & A298;
  assign \new_[66378]_  = A301 & A300;
  assign \new_[66379]_  = \new_[66378]_  & \new_[66375]_ ;
  assign \new_[66380]_  = \new_[66379]_  & \new_[66372]_ ;
  assign \new_[66384]_  = A167 & A169;
  assign \new_[66385]_  = ~A170 & \new_[66384]_ ;
  assign \new_[66388]_  = ~A200 & A166;
  assign \new_[66391]_  = ~A233 & ~A201;
  assign \new_[66392]_  = \new_[66391]_  & \new_[66388]_ ;
  assign \new_[66393]_  = \new_[66392]_  & \new_[66385]_ ;
  assign \new_[66396]_  = ~A266 & ~A234;
  assign \new_[66399]_  = ~A269 & ~A268;
  assign \new_[66400]_  = \new_[66399]_  & \new_[66396]_ ;
  assign \new_[66403]_  = ~A299 & A298;
  assign \new_[66406]_  = A302 & A300;
  assign \new_[66407]_  = \new_[66406]_  & \new_[66403]_ ;
  assign \new_[66408]_  = \new_[66407]_  & \new_[66400]_ ;
  assign \new_[66412]_  = A167 & A169;
  assign \new_[66413]_  = ~A170 & \new_[66412]_ ;
  assign \new_[66416]_  = ~A200 & A166;
  assign \new_[66419]_  = ~A232 & ~A201;
  assign \new_[66420]_  = \new_[66419]_  & \new_[66416]_ ;
  assign \new_[66421]_  = \new_[66420]_  & \new_[66413]_ ;
  assign \new_[66424]_  = ~A266 & ~A233;
  assign \new_[66427]_  = ~A269 & ~A268;
  assign \new_[66428]_  = \new_[66427]_  & \new_[66424]_ ;
  assign \new_[66431]_  = ~A299 & A298;
  assign \new_[66434]_  = A301 & A300;
  assign \new_[66435]_  = \new_[66434]_  & \new_[66431]_ ;
  assign \new_[66436]_  = \new_[66435]_  & \new_[66428]_ ;
  assign \new_[66440]_  = A167 & A169;
  assign \new_[66441]_  = ~A170 & \new_[66440]_ ;
  assign \new_[66444]_  = ~A200 & A166;
  assign \new_[66447]_  = ~A232 & ~A201;
  assign \new_[66448]_  = \new_[66447]_  & \new_[66444]_ ;
  assign \new_[66449]_  = \new_[66448]_  & \new_[66441]_ ;
  assign \new_[66452]_  = ~A266 & ~A233;
  assign \new_[66455]_  = ~A269 & ~A268;
  assign \new_[66456]_  = \new_[66455]_  & \new_[66452]_ ;
  assign \new_[66459]_  = ~A299 & A298;
  assign \new_[66462]_  = A302 & A300;
  assign \new_[66463]_  = \new_[66462]_  & \new_[66459]_ ;
  assign \new_[66464]_  = \new_[66463]_  & \new_[66456]_ ;
  assign \new_[66468]_  = A167 & A169;
  assign \new_[66469]_  = ~A170 & \new_[66468]_ ;
  assign \new_[66472]_  = ~A199 & A166;
  assign \new_[66475]_  = A232 & ~A200;
  assign \new_[66476]_  = \new_[66475]_  & \new_[66472]_ ;
  assign \new_[66477]_  = \new_[66476]_  & \new_[66469]_ ;
  assign \new_[66480]_  = A265 & A233;
  assign \new_[66483]_  = ~A269 & ~A268;
  assign \new_[66484]_  = \new_[66483]_  & \new_[66480]_ ;
  assign \new_[66487]_  = ~A299 & A298;
  assign \new_[66490]_  = A301 & A300;
  assign \new_[66491]_  = \new_[66490]_  & \new_[66487]_ ;
  assign \new_[66492]_  = \new_[66491]_  & \new_[66484]_ ;
  assign \new_[66496]_  = A167 & A169;
  assign \new_[66497]_  = ~A170 & \new_[66496]_ ;
  assign \new_[66500]_  = ~A199 & A166;
  assign \new_[66503]_  = A232 & ~A200;
  assign \new_[66504]_  = \new_[66503]_  & \new_[66500]_ ;
  assign \new_[66505]_  = \new_[66504]_  & \new_[66497]_ ;
  assign \new_[66508]_  = A265 & A233;
  assign \new_[66511]_  = ~A269 & ~A268;
  assign \new_[66512]_  = \new_[66511]_  & \new_[66508]_ ;
  assign \new_[66515]_  = ~A299 & A298;
  assign \new_[66518]_  = A302 & A300;
  assign \new_[66519]_  = \new_[66518]_  & \new_[66515]_ ;
  assign \new_[66520]_  = \new_[66519]_  & \new_[66512]_ ;
  assign \new_[66524]_  = A167 & A169;
  assign \new_[66525]_  = ~A170 & \new_[66524]_ ;
  assign \new_[66528]_  = ~A199 & A166;
  assign \new_[66531]_  = ~A233 & ~A200;
  assign \new_[66532]_  = \new_[66531]_  & \new_[66528]_ ;
  assign \new_[66533]_  = \new_[66532]_  & \new_[66525]_ ;
  assign \new_[66536]_  = ~A236 & ~A235;
  assign \new_[66539]_  = A266 & A265;
  assign \new_[66540]_  = \new_[66539]_  & \new_[66536]_ ;
  assign \new_[66543]_  = ~A299 & A298;
  assign \new_[66546]_  = A301 & A300;
  assign \new_[66547]_  = \new_[66546]_  & \new_[66543]_ ;
  assign \new_[66548]_  = \new_[66547]_  & \new_[66540]_ ;
  assign \new_[66552]_  = A167 & A169;
  assign \new_[66553]_  = ~A170 & \new_[66552]_ ;
  assign \new_[66556]_  = ~A199 & A166;
  assign \new_[66559]_  = ~A233 & ~A200;
  assign \new_[66560]_  = \new_[66559]_  & \new_[66556]_ ;
  assign \new_[66561]_  = \new_[66560]_  & \new_[66553]_ ;
  assign \new_[66564]_  = ~A236 & ~A235;
  assign \new_[66567]_  = A266 & A265;
  assign \new_[66568]_  = \new_[66567]_  & \new_[66564]_ ;
  assign \new_[66571]_  = ~A299 & A298;
  assign \new_[66574]_  = A302 & A300;
  assign \new_[66575]_  = \new_[66574]_  & \new_[66571]_ ;
  assign \new_[66576]_  = \new_[66575]_  & \new_[66568]_ ;
  assign \new_[66580]_  = A167 & A169;
  assign \new_[66581]_  = ~A170 & \new_[66580]_ ;
  assign \new_[66584]_  = ~A199 & A166;
  assign \new_[66587]_  = ~A233 & ~A200;
  assign \new_[66588]_  = \new_[66587]_  & \new_[66584]_ ;
  assign \new_[66589]_  = \new_[66588]_  & \new_[66581]_ ;
  assign \new_[66592]_  = ~A236 & ~A235;
  assign \new_[66595]_  = ~A267 & ~A266;
  assign \new_[66596]_  = \new_[66595]_  & \new_[66592]_ ;
  assign \new_[66599]_  = ~A299 & A298;
  assign \new_[66602]_  = A301 & A300;
  assign \new_[66603]_  = \new_[66602]_  & \new_[66599]_ ;
  assign \new_[66604]_  = \new_[66603]_  & \new_[66596]_ ;
  assign \new_[66608]_  = A167 & A169;
  assign \new_[66609]_  = ~A170 & \new_[66608]_ ;
  assign \new_[66612]_  = ~A199 & A166;
  assign \new_[66615]_  = ~A233 & ~A200;
  assign \new_[66616]_  = \new_[66615]_  & \new_[66612]_ ;
  assign \new_[66617]_  = \new_[66616]_  & \new_[66609]_ ;
  assign \new_[66620]_  = ~A236 & ~A235;
  assign \new_[66623]_  = ~A267 & ~A266;
  assign \new_[66624]_  = \new_[66623]_  & \new_[66620]_ ;
  assign \new_[66627]_  = ~A299 & A298;
  assign \new_[66630]_  = A302 & A300;
  assign \new_[66631]_  = \new_[66630]_  & \new_[66627]_ ;
  assign \new_[66632]_  = \new_[66631]_  & \new_[66624]_ ;
  assign \new_[66636]_  = A167 & A169;
  assign \new_[66637]_  = ~A170 & \new_[66636]_ ;
  assign \new_[66640]_  = ~A199 & A166;
  assign \new_[66643]_  = ~A233 & ~A200;
  assign \new_[66644]_  = \new_[66643]_  & \new_[66640]_ ;
  assign \new_[66645]_  = \new_[66644]_  & \new_[66637]_ ;
  assign \new_[66648]_  = ~A236 & ~A235;
  assign \new_[66651]_  = ~A266 & ~A265;
  assign \new_[66652]_  = \new_[66651]_  & \new_[66648]_ ;
  assign \new_[66655]_  = ~A299 & A298;
  assign \new_[66658]_  = A301 & A300;
  assign \new_[66659]_  = \new_[66658]_  & \new_[66655]_ ;
  assign \new_[66660]_  = \new_[66659]_  & \new_[66652]_ ;
  assign \new_[66664]_  = A167 & A169;
  assign \new_[66665]_  = ~A170 & \new_[66664]_ ;
  assign \new_[66668]_  = ~A199 & A166;
  assign \new_[66671]_  = ~A233 & ~A200;
  assign \new_[66672]_  = \new_[66671]_  & \new_[66668]_ ;
  assign \new_[66673]_  = \new_[66672]_  & \new_[66665]_ ;
  assign \new_[66676]_  = ~A236 & ~A235;
  assign \new_[66679]_  = ~A266 & ~A265;
  assign \new_[66680]_  = \new_[66679]_  & \new_[66676]_ ;
  assign \new_[66683]_  = ~A299 & A298;
  assign \new_[66686]_  = A302 & A300;
  assign \new_[66687]_  = \new_[66686]_  & \new_[66683]_ ;
  assign \new_[66688]_  = \new_[66687]_  & \new_[66680]_ ;
  assign \new_[66692]_  = A167 & A169;
  assign \new_[66693]_  = ~A170 & \new_[66692]_ ;
  assign \new_[66696]_  = ~A199 & A166;
  assign \new_[66699]_  = ~A233 & ~A200;
  assign \new_[66700]_  = \new_[66699]_  & \new_[66696]_ ;
  assign \new_[66701]_  = \new_[66700]_  & \new_[66693]_ ;
  assign \new_[66704]_  = ~A266 & ~A234;
  assign \new_[66707]_  = ~A269 & ~A268;
  assign \new_[66708]_  = \new_[66707]_  & \new_[66704]_ ;
  assign \new_[66711]_  = ~A299 & A298;
  assign \new_[66714]_  = A301 & A300;
  assign \new_[66715]_  = \new_[66714]_  & \new_[66711]_ ;
  assign \new_[66716]_  = \new_[66715]_  & \new_[66708]_ ;
  assign \new_[66720]_  = A167 & A169;
  assign \new_[66721]_  = ~A170 & \new_[66720]_ ;
  assign \new_[66724]_  = ~A199 & A166;
  assign \new_[66727]_  = ~A233 & ~A200;
  assign \new_[66728]_  = \new_[66727]_  & \new_[66724]_ ;
  assign \new_[66729]_  = \new_[66728]_  & \new_[66721]_ ;
  assign \new_[66732]_  = ~A266 & ~A234;
  assign \new_[66735]_  = ~A269 & ~A268;
  assign \new_[66736]_  = \new_[66735]_  & \new_[66732]_ ;
  assign \new_[66739]_  = ~A299 & A298;
  assign \new_[66742]_  = A302 & A300;
  assign \new_[66743]_  = \new_[66742]_  & \new_[66739]_ ;
  assign \new_[66744]_  = \new_[66743]_  & \new_[66736]_ ;
  assign \new_[66748]_  = A167 & A169;
  assign \new_[66749]_  = ~A170 & \new_[66748]_ ;
  assign \new_[66752]_  = ~A199 & A166;
  assign \new_[66755]_  = ~A232 & ~A200;
  assign \new_[66756]_  = \new_[66755]_  & \new_[66752]_ ;
  assign \new_[66757]_  = \new_[66756]_  & \new_[66749]_ ;
  assign \new_[66760]_  = ~A266 & ~A233;
  assign \new_[66763]_  = ~A269 & ~A268;
  assign \new_[66764]_  = \new_[66763]_  & \new_[66760]_ ;
  assign \new_[66767]_  = ~A299 & A298;
  assign \new_[66770]_  = A301 & A300;
  assign \new_[66771]_  = \new_[66770]_  & \new_[66767]_ ;
  assign \new_[66772]_  = \new_[66771]_  & \new_[66764]_ ;
  assign \new_[66776]_  = A167 & A169;
  assign \new_[66777]_  = ~A170 & \new_[66776]_ ;
  assign \new_[66780]_  = ~A199 & A166;
  assign \new_[66783]_  = ~A232 & ~A200;
  assign \new_[66784]_  = \new_[66783]_  & \new_[66780]_ ;
  assign \new_[66785]_  = \new_[66784]_  & \new_[66777]_ ;
  assign \new_[66788]_  = ~A266 & ~A233;
  assign \new_[66791]_  = ~A269 & ~A268;
  assign \new_[66792]_  = \new_[66791]_  & \new_[66788]_ ;
  assign \new_[66795]_  = ~A299 & A298;
  assign \new_[66798]_  = A302 & A300;
  assign \new_[66799]_  = \new_[66798]_  & \new_[66795]_ ;
  assign \new_[66800]_  = \new_[66799]_  & \new_[66792]_ ;
  assign \new_[66804]_  = ~A167 & A169;
  assign \new_[66805]_  = ~A170 & \new_[66804]_ ;
  assign \new_[66808]_  = A199 & ~A166;
  assign \new_[66811]_  = A232 & A200;
  assign \new_[66812]_  = \new_[66811]_  & \new_[66808]_ ;
  assign \new_[66813]_  = \new_[66812]_  & \new_[66805]_ ;
  assign \new_[66816]_  = A265 & A233;
  assign \new_[66819]_  = ~A269 & ~A268;
  assign \new_[66820]_  = \new_[66819]_  & \new_[66816]_ ;
  assign \new_[66823]_  = ~A299 & A298;
  assign \new_[66826]_  = A301 & A300;
  assign \new_[66827]_  = \new_[66826]_  & \new_[66823]_ ;
  assign \new_[66828]_  = \new_[66827]_  & \new_[66820]_ ;
  assign \new_[66832]_  = ~A167 & A169;
  assign \new_[66833]_  = ~A170 & \new_[66832]_ ;
  assign \new_[66836]_  = A199 & ~A166;
  assign \new_[66839]_  = A232 & A200;
  assign \new_[66840]_  = \new_[66839]_  & \new_[66836]_ ;
  assign \new_[66841]_  = \new_[66840]_  & \new_[66833]_ ;
  assign \new_[66844]_  = A265 & A233;
  assign \new_[66847]_  = ~A269 & ~A268;
  assign \new_[66848]_  = \new_[66847]_  & \new_[66844]_ ;
  assign \new_[66851]_  = ~A299 & A298;
  assign \new_[66854]_  = A302 & A300;
  assign \new_[66855]_  = \new_[66854]_  & \new_[66851]_ ;
  assign \new_[66856]_  = \new_[66855]_  & \new_[66848]_ ;
  assign \new_[66860]_  = ~A167 & A169;
  assign \new_[66861]_  = ~A170 & \new_[66860]_ ;
  assign \new_[66864]_  = A199 & ~A166;
  assign \new_[66867]_  = ~A233 & A200;
  assign \new_[66868]_  = \new_[66867]_  & \new_[66864]_ ;
  assign \new_[66869]_  = \new_[66868]_  & \new_[66861]_ ;
  assign \new_[66872]_  = ~A236 & ~A235;
  assign \new_[66875]_  = A266 & A265;
  assign \new_[66876]_  = \new_[66875]_  & \new_[66872]_ ;
  assign \new_[66879]_  = ~A299 & A298;
  assign \new_[66882]_  = A301 & A300;
  assign \new_[66883]_  = \new_[66882]_  & \new_[66879]_ ;
  assign \new_[66884]_  = \new_[66883]_  & \new_[66876]_ ;
  assign \new_[66888]_  = ~A167 & A169;
  assign \new_[66889]_  = ~A170 & \new_[66888]_ ;
  assign \new_[66892]_  = A199 & ~A166;
  assign \new_[66895]_  = ~A233 & A200;
  assign \new_[66896]_  = \new_[66895]_  & \new_[66892]_ ;
  assign \new_[66897]_  = \new_[66896]_  & \new_[66889]_ ;
  assign \new_[66900]_  = ~A236 & ~A235;
  assign \new_[66903]_  = A266 & A265;
  assign \new_[66904]_  = \new_[66903]_  & \new_[66900]_ ;
  assign \new_[66907]_  = ~A299 & A298;
  assign \new_[66910]_  = A302 & A300;
  assign \new_[66911]_  = \new_[66910]_  & \new_[66907]_ ;
  assign \new_[66912]_  = \new_[66911]_  & \new_[66904]_ ;
  assign \new_[66916]_  = ~A167 & A169;
  assign \new_[66917]_  = ~A170 & \new_[66916]_ ;
  assign \new_[66920]_  = A199 & ~A166;
  assign \new_[66923]_  = ~A233 & A200;
  assign \new_[66924]_  = \new_[66923]_  & \new_[66920]_ ;
  assign \new_[66925]_  = \new_[66924]_  & \new_[66917]_ ;
  assign \new_[66928]_  = ~A236 & ~A235;
  assign \new_[66931]_  = ~A267 & ~A266;
  assign \new_[66932]_  = \new_[66931]_  & \new_[66928]_ ;
  assign \new_[66935]_  = ~A299 & A298;
  assign \new_[66938]_  = A301 & A300;
  assign \new_[66939]_  = \new_[66938]_  & \new_[66935]_ ;
  assign \new_[66940]_  = \new_[66939]_  & \new_[66932]_ ;
  assign \new_[66944]_  = ~A167 & A169;
  assign \new_[66945]_  = ~A170 & \new_[66944]_ ;
  assign \new_[66948]_  = A199 & ~A166;
  assign \new_[66951]_  = ~A233 & A200;
  assign \new_[66952]_  = \new_[66951]_  & \new_[66948]_ ;
  assign \new_[66953]_  = \new_[66952]_  & \new_[66945]_ ;
  assign \new_[66956]_  = ~A236 & ~A235;
  assign \new_[66959]_  = ~A267 & ~A266;
  assign \new_[66960]_  = \new_[66959]_  & \new_[66956]_ ;
  assign \new_[66963]_  = ~A299 & A298;
  assign \new_[66966]_  = A302 & A300;
  assign \new_[66967]_  = \new_[66966]_  & \new_[66963]_ ;
  assign \new_[66968]_  = \new_[66967]_  & \new_[66960]_ ;
  assign \new_[66972]_  = ~A167 & A169;
  assign \new_[66973]_  = ~A170 & \new_[66972]_ ;
  assign \new_[66976]_  = A199 & ~A166;
  assign \new_[66979]_  = ~A233 & A200;
  assign \new_[66980]_  = \new_[66979]_  & \new_[66976]_ ;
  assign \new_[66981]_  = \new_[66980]_  & \new_[66973]_ ;
  assign \new_[66984]_  = ~A236 & ~A235;
  assign \new_[66987]_  = ~A266 & ~A265;
  assign \new_[66988]_  = \new_[66987]_  & \new_[66984]_ ;
  assign \new_[66991]_  = ~A299 & A298;
  assign \new_[66994]_  = A301 & A300;
  assign \new_[66995]_  = \new_[66994]_  & \new_[66991]_ ;
  assign \new_[66996]_  = \new_[66995]_  & \new_[66988]_ ;
  assign \new_[67000]_  = ~A167 & A169;
  assign \new_[67001]_  = ~A170 & \new_[67000]_ ;
  assign \new_[67004]_  = A199 & ~A166;
  assign \new_[67007]_  = ~A233 & A200;
  assign \new_[67008]_  = \new_[67007]_  & \new_[67004]_ ;
  assign \new_[67009]_  = \new_[67008]_  & \new_[67001]_ ;
  assign \new_[67012]_  = ~A236 & ~A235;
  assign \new_[67015]_  = ~A266 & ~A265;
  assign \new_[67016]_  = \new_[67015]_  & \new_[67012]_ ;
  assign \new_[67019]_  = ~A299 & A298;
  assign \new_[67022]_  = A302 & A300;
  assign \new_[67023]_  = \new_[67022]_  & \new_[67019]_ ;
  assign \new_[67024]_  = \new_[67023]_  & \new_[67016]_ ;
  assign \new_[67028]_  = ~A167 & A169;
  assign \new_[67029]_  = ~A170 & \new_[67028]_ ;
  assign \new_[67032]_  = A199 & ~A166;
  assign \new_[67035]_  = ~A233 & A200;
  assign \new_[67036]_  = \new_[67035]_  & \new_[67032]_ ;
  assign \new_[67037]_  = \new_[67036]_  & \new_[67029]_ ;
  assign \new_[67040]_  = ~A266 & ~A234;
  assign \new_[67043]_  = ~A269 & ~A268;
  assign \new_[67044]_  = \new_[67043]_  & \new_[67040]_ ;
  assign \new_[67047]_  = ~A299 & A298;
  assign \new_[67050]_  = A301 & A300;
  assign \new_[67051]_  = \new_[67050]_  & \new_[67047]_ ;
  assign \new_[67052]_  = \new_[67051]_  & \new_[67044]_ ;
  assign \new_[67056]_  = ~A167 & A169;
  assign \new_[67057]_  = ~A170 & \new_[67056]_ ;
  assign \new_[67060]_  = A199 & ~A166;
  assign \new_[67063]_  = ~A233 & A200;
  assign \new_[67064]_  = \new_[67063]_  & \new_[67060]_ ;
  assign \new_[67065]_  = \new_[67064]_  & \new_[67057]_ ;
  assign \new_[67068]_  = ~A266 & ~A234;
  assign \new_[67071]_  = ~A269 & ~A268;
  assign \new_[67072]_  = \new_[67071]_  & \new_[67068]_ ;
  assign \new_[67075]_  = ~A299 & A298;
  assign \new_[67078]_  = A302 & A300;
  assign \new_[67079]_  = \new_[67078]_  & \new_[67075]_ ;
  assign \new_[67080]_  = \new_[67079]_  & \new_[67072]_ ;
  assign \new_[67084]_  = ~A167 & A169;
  assign \new_[67085]_  = ~A170 & \new_[67084]_ ;
  assign \new_[67088]_  = A199 & ~A166;
  assign \new_[67091]_  = ~A232 & A200;
  assign \new_[67092]_  = \new_[67091]_  & \new_[67088]_ ;
  assign \new_[67093]_  = \new_[67092]_  & \new_[67085]_ ;
  assign \new_[67096]_  = ~A266 & ~A233;
  assign \new_[67099]_  = ~A269 & ~A268;
  assign \new_[67100]_  = \new_[67099]_  & \new_[67096]_ ;
  assign \new_[67103]_  = ~A299 & A298;
  assign \new_[67106]_  = A301 & A300;
  assign \new_[67107]_  = \new_[67106]_  & \new_[67103]_ ;
  assign \new_[67108]_  = \new_[67107]_  & \new_[67100]_ ;
  assign \new_[67112]_  = ~A167 & A169;
  assign \new_[67113]_  = ~A170 & \new_[67112]_ ;
  assign \new_[67116]_  = A199 & ~A166;
  assign \new_[67119]_  = ~A232 & A200;
  assign \new_[67120]_  = \new_[67119]_  & \new_[67116]_ ;
  assign \new_[67121]_  = \new_[67120]_  & \new_[67113]_ ;
  assign \new_[67124]_  = ~A266 & ~A233;
  assign \new_[67127]_  = ~A269 & ~A268;
  assign \new_[67128]_  = \new_[67127]_  & \new_[67124]_ ;
  assign \new_[67131]_  = ~A299 & A298;
  assign \new_[67134]_  = A302 & A300;
  assign \new_[67135]_  = \new_[67134]_  & \new_[67131]_ ;
  assign \new_[67136]_  = \new_[67135]_  & \new_[67128]_ ;
  assign \new_[67140]_  = ~A167 & A169;
  assign \new_[67141]_  = ~A170 & \new_[67140]_ ;
  assign \new_[67144]_  = ~A200 & ~A166;
  assign \new_[67147]_  = ~A203 & ~A202;
  assign \new_[67148]_  = \new_[67147]_  & \new_[67144]_ ;
  assign \new_[67149]_  = \new_[67148]_  & \new_[67141]_ ;
  assign \new_[67152]_  = A233 & A232;
  assign \new_[67155]_  = ~A267 & A265;
  assign \new_[67156]_  = \new_[67155]_  & \new_[67152]_ ;
  assign \new_[67159]_  = ~A299 & A298;
  assign \new_[67162]_  = A301 & A300;
  assign \new_[67163]_  = \new_[67162]_  & \new_[67159]_ ;
  assign \new_[67164]_  = \new_[67163]_  & \new_[67156]_ ;
  assign \new_[67168]_  = ~A167 & A169;
  assign \new_[67169]_  = ~A170 & \new_[67168]_ ;
  assign \new_[67172]_  = ~A200 & ~A166;
  assign \new_[67175]_  = ~A203 & ~A202;
  assign \new_[67176]_  = \new_[67175]_  & \new_[67172]_ ;
  assign \new_[67177]_  = \new_[67176]_  & \new_[67169]_ ;
  assign \new_[67180]_  = A233 & A232;
  assign \new_[67183]_  = ~A267 & A265;
  assign \new_[67184]_  = \new_[67183]_  & \new_[67180]_ ;
  assign \new_[67187]_  = ~A299 & A298;
  assign \new_[67190]_  = A302 & A300;
  assign \new_[67191]_  = \new_[67190]_  & \new_[67187]_ ;
  assign \new_[67192]_  = \new_[67191]_  & \new_[67184]_ ;
  assign \new_[67196]_  = ~A167 & A169;
  assign \new_[67197]_  = ~A170 & \new_[67196]_ ;
  assign \new_[67200]_  = ~A200 & ~A166;
  assign \new_[67203]_  = ~A203 & ~A202;
  assign \new_[67204]_  = \new_[67203]_  & \new_[67200]_ ;
  assign \new_[67205]_  = \new_[67204]_  & \new_[67197]_ ;
  assign \new_[67208]_  = A233 & A232;
  assign \new_[67211]_  = A266 & A265;
  assign \new_[67212]_  = \new_[67211]_  & \new_[67208]_ ;
  assign \new_[67215]_  = ~A299 & A298;
  assign \new_[67218]_  = A301 & A300;
  assign \new_[67219]_  = \new_[67218]_  & \new_[67215]_ ;
  assign \new_[67220]_  = \new_[67219]_  & \new_[67212]_ ;
  assign \new_[67224]_  = ~A167 & A169;
  assign \new_[67225]_  = ~A170 & \new_[67224]_ ;
  assign \new_[67228]_  = ~A200 & ~A166;
  assign \new_[67231]_  = ~A203 & ~A202;
  assign \new_[67232]_  = \new_[67231]_  & \new_[67228]_ ;
  assign \new_[67233]_  = \new_[67232]_  & \new_[67225]_ ;
  assign \new_[67236]_  = A233 & A232;
  assign \new_[67239]_  = A266 & A265;
  assign \new_[67240]_  = \new_[67239]_  & \new_[67236]_ ;
  assign \new_[67243]_  = ~A299 & A298;
  assign \new_[67246]_  = A302 & A300;
  assign \new_[67247]_  = \new_[67246]_  & \new_[67243]_ ;
  assign \new_[67248]_  = \new_[67247]_  & \new_[67240]_ ;
  assign \new_[67252]_  = ~A167 & A169;
  assign \new_[67253]_  = ~A170 & \new_[67252]_ ;
  assign \new_[67256]_  = ~A200 & ~A166;
  assign \new_[67259]_  = ~A203 & ~A202;
  assign \new_[67260]_  = \new_[67259]_  & \new_[67256]_ ;
  assign \new_[67261]_  = \new_[67260]_  & \new_[67253]_ ;
  assign \new_[67264]_  = A233 & A232;
  assign \new_[67267]_  = ~A266 & ~A265;
  assign \new_[67268]_  = \new_[67267]_  & \new_[67264]_ ;
  assign \new_[67271]_  = ~A299 & A298;
  assign \new_[67274]_  = A301 & A300;
  assign \new_[67275]_  = \new_[67274]_  & \new_[67271]_ ;
  assign \new_[67276]_  = \new_[67275]_  & \new_[67268]_ ;
  assign \new_[67280]_  = ~A167 & A169;
  assign \new_[67281]_  = ~A170 & \new_[67280]_ ;
  assign \new_[67284]_  = ~A200 & ~A166;
  assign \new_[67287]_  = ~A203 & ~A202;
  assign \new_[67288]_  = \new_[67287]_  & \new_[67284]_ ;
  assign \new_[67289]_  = \new_[67288]_  & \new_[67281]_ ;
  assign \new_[67292]_  = A233 & A232;
  assign \new_[67295]_  = ~A266 & ~A265;
  assign \new_[67296]_  = \new_[67295]_  & \new_[67292]_ ;
  assign \new_[67299]_  = ~A299 & A298;
  assign \new_[67302]_  = A302 & A300;
  assign \new_[67303]_  = \new_[67302]_  & \new_[67299]_ ;
  assign \new_[67304]_  = \new_[67303]_  & \new_[67296]_ ;
  assign \new_[67308]_  = ~A167 & A169;
  assign \new_[67309]_  = ~A170 & \new_[67308]_ ;
  assign \new_[67312]_  = ~A200 & ~A166;
  assign \new_[67315]_  = ~A203 & ~A202;
  assign \new_[67316]_  = \new_[67315]_  & \new_[67312]_ ;
  assign \new_[67317]_  = \new_[67316]_  & \new_[67309]_ ;
  assign \new_[67320]_  = ~A235 & ~A233;
  assign \new_[67323]_  = ~A266 & ~A236;
  assign \new_[67324]_  = \new_[67323]_  & \new_[67320]_ ;
  assign \new_[67327]_  = ~A269 & ~A268;
  assign \new_[67330]_  = A299 & ~A298;
  assign \new_[67331]_  = \new_[67330]_  & \new_[67327]_ ;
  assign \new_[67332]_  = \new_[67331]_  & \new_[67324]_ ;
  assign \new_[67336]_  = ~A167 & A169;
  assign \new_[67337]_  = ~A170 & \new_[67336]_ ;
  assign \new_[67340]_  = ~A200 & ~A166;
  assign \new_[67343]_  = ~A203 & ~A202;
  assign \new_[67344]_  = \new_[67343]_  & \new_[67340]_ ;
  assign \new_[67345]_  = \new_[67344]_  & \new_[67337]_ ;
  assign \new_[67348]_  = ~A234 & ~A233;
  assign \new_[67351]_  = A266 & A265;
  assign \new_[67352]_  = \new_[67351]_  & \new_[67348]_ ;
  assign \new_[67355]_  = ~A299 & A298;
  assign \new_[67358]_  = A301 & A300;
  assign \new_[67359]_  = \new_[67358]_  & \new_[67355]_ ;
  assign \new_[67360]_  = \new_[67359]_  & \new_[67352]_ ;
  assign \new_[67364]_  = ~A167 & A169;
  assign \new_[67365]_  = ~A170 & \new_[67364]_ ;
  assign \new_[67368]_  = ~A200 & ~A166;
  assign \new_[67371]_  = ~A203 & ~A202;
  assign \new_[67372]_  = \new_[67371]_  & \new_[67368]_ ;
  assign \new_[67373]_  = \new_[67372]_  & \new_[67365]_ ;
  assign \new_[67376]_  = ~A234 & ~A233;
  assign \new_[67379]_  = A266 & A265;
  assign \new_[67380]_  = \new_[67379]_  & \new_[67376]_ ;
  assign \new_[67383]_  = ~A299 & A298;
  assign \new_[67386]_  = A302 & A300;
  assign \new_[67387]_  = \new_[67386]_  & \new_[67383]_ ;
  assign \new_[67388]_  = \new_[67387]_  & \new_[67380]_ ;
  assign \new_[67392]_  = ~A167 & A169;
  assign \new_[67393]_  = ~A170 & \new_[67392]_ ;
  assign \new_[67396]_  = ~A200 & ~A166;
  assign \new_[67399]_  = ~A203 & ~A202;
  assign \new_[67400]_  = \new_[67399]_  & \new_[67396]_ ;
  assign \new_[67401]_  = \new_[67400]_  & \new_[67393]_ ;
  assign \new_[67404]_  = ~A234 & ~A233;
  assign \new_[67407]_  = ~A267 & ~A266;
  assign \new_[67408]_  = \new_[67407]_  & \new_[67404]_ ;
  assign \new_[67411]_  = ~A299 & A298;
  assign \new_[67414]_  = A301 & A300;
  assign \new_[67415]_  = \new_[67414]_  & \new_[67411]_ ;
  assign \new_[67416]_  = \new_[67415]_  & \new_[67408]_ ;
  assign \new_[67420]_  = ~A167 & A169;
  assign \new_[67421]_  = ~A170 & \new_[67420]_ ;
  assign \new_[67424]_  = ~A200 & ~A166;
  assign \new_[67427]_  = ~A203 & ~A202;
  assign \new_[67428]_  = \new_[67427]_  & \new_[67424]_ ;
  assign \new_[67429]_  = \new_[67428]_  & \new_[67421]_ ;
  assign \new_[67432]_  = ~A234 & ~A233;
  assign \new_[67435]_  = ~A267 & ~A266;
  assign \new_[67436]_  = \new_[67435]_  & \new_[67432]_ ;
  assign \new_[67439]_  = ~A299 & A298;
  assign \new_[67442]_  = A302 & A300;
  assign \new_[67443]_  = \new_[67442]_  & \new_[67439]_ ;
  assign \new_[67444]_  = \new_[67443]_  & \new_[67436]_ ;
  assign \new_[67448]_  = ~A167 & A169;
  assign \new_[67449]_  = ~A170 & \new_[67448]_ ;
  assign \new_[67452]_  = ~A200 & ~A166;
  assign \new_[67455]_  = ~A203 & ~A202;
  assign \new_[67456]_  = \new_[67455]_  & \new_[67452]_ ;
  assign \new_[67457]_  = \new_[67456]_  & \new_[67449]_ ;
  assign \new_[67460]_  = ~A234 & ~A233;
  assign \new_[67463]_  = ~A266 & ~A265;
  assign \new_[67464]_  = \new_[67463]_  & \new_[67460]_ ;
  assign \new_[67467]_  = ~A299 & A298;
  assign \new_[67470]_  = A301 & A300;
  assign \new_[67471]_  = \new_[67470]_  & \new_[67467]_ ;
  assign \new_[67472]_  = \new_[67471]_  & \new_[67464]_ ;
  assign \new_[67476]_  = ~A167 & A169;
  assign \new_[67477]_  = ~A170 & \new_[67476]_ ;
  assign \new_[67480]_  = ~A200 & ~A166;
  assign \new_[67483]_  = ~A203 & ~A202;
  assign \new_[67484]_  = \new_[67483]_  & \new_[67480]_ ;
  assign \new_[67485]_  = \new_[67484]_  & \new_[67477]_ ;
  assign \new_[67488]_  = ~A234 & ~A233;
  assign \new_[67491]_  = ~A266 & ~A265;
  assign \new_[67492]_  = \new_[67491]_  & \new_[67488]_ ;
  assign \new_[67495]_  = ~A299 & A298;
  assign \new_[67498]_  = A302 & A300;
  assign \new_[67499]_  = \new_[67498]_  & \new_[67495]_ ;
  assign \new_[67500]_  = \new_[67499]_  & \new_[67492]_ ;
  assign \new_[67504]_  = ~A167 & A169;
  assign \new_[67505]_  = ~A170 & \new_[67504]_ ;
  assign \new_[67508]_  = ~A200 & ~A166;
  assign \new_[67511]_  = ~A203 & ~A202;
  assign \new_[67512]_  = \new_[67511]_  & \new_[67508]_ ;
  assign \new_[67513]_  = \new_[67512]_  & \new_[67505]_ ;
  assign \new_[67516]_  = ~A233 & A232;
  assign \new_[67519]_  = A235 & A234;
  assign \new_[67520]_  = \new_[67519]_  & \new_[67516]_ ;
  assign \new_[67523]_  = ~A266 & A265;
  assign \new_[67526]_  = A268 & A267;
  assign \new_[67527]_  = \new_[67526]_  & \new_[67523]_ ;
  assign \new_[67528]_  = \new_[67527]_  & \new_[67520]_ ;
  assign \new_[67532]_  = ~A167 & A169;
  assign \new_[67533]_  = ~A170 & \new_[67532]_ ;
  assign \new_[67536]_  = ~A200 & ~A166;
  assign \new_[67539]_  = ~A203 & ~A202;
  assign \new_[67540]_  = \new_[67539]_  & \new_[67536]_ ;
  assign \new_[67541]_  = \new_[67540]_  & \new_[67533]_ ;
  assign \new_[67544]_  = ~A233 & A232;
  assign \new_[67547]_  = A235 & A234;
  assign \new_[67548]_  = \new_[67547]_  & \new_[67544]_ ;
  assign \new_[67551]_  = ~A266 & A265;
  assign \new_[67554]_  = A269 & A267;
  assign \new_[67555]_  = \new_[67554]_  & \new_[67551]_ ;
  assign \new_[67556]_  = \new_[67555]_  & \new_[67548]_ ;
  assign \new_[67560]_  = ~A167 & A169;
  assign \new_[67561]_  = ~A170 & \new_[67560]_ ;
  assign \new_[67564]_  = ~A200 & ~A166;
  assign \new_[67567]_  = ~A203 & ~A202;
  assign \new_[67568]_  = \new_[67567]_  & \new_[67564]_ ;
  assign \new_[67569]_  = \new_[67568]_  & \new_[67561]_ ;
  assign \new_[67572]_  = ~A233 & A232;
  assign \new_[67575]_  = A236 & A234;
  assign \new_[67576]_  = \new_[67575]_  & \new_[67572]_ ;
  assign \new_[67579]_  = ~A266 & A265;
  assign \new_[67582]_  = A268 & A267;
  assign \new_[67583]_  = \new_[67582]_  & \new_[67579]_ ;
  assign \new_[67584]_  = \new_[67583]_  & \new_[67576]_ ;
  assign \new_[67588]_  = ~A167 & A169;
  assign \new_[67589]_  = ~A170 & \new_[67588]_ ;
  assign \new_[67592]_  = ~A200 & ~A166;
  assign \new_[67595]_  = ~A203 & ~A202;
  assign \new_[67596]_  = \new_[67595]_  & \new_[67592]_ ;
  assign \new_[67597]_  = \new_[67596]_  & \new_[67589]_ ;
  assign \new_[67600]_  = ~A233 & A232;
  assign \new_[67603]_  = A236 & A234;
  assign \new_[67604]_  = \new_[67603]_  & \new_[67600]_ ;
  assign \new_[67607]_  = ~A266 & A265;
  assign \new_[67610]_  = A269 & A267;
  assign \new_[67611]_  = \new_[67610]_  & \new_[67607]_ ;
  assign \new_[67612]_  = \new_[67611]_  & \new_[67604]_ ;
  assign \new_[67616]_  = ~A167 & A169;
  assign \new_[67617]_  = ~A170 & \new_[67616]_ ;
  assign \new_[67620]_  = ~A200 & ~A166;
  assign \new_[67623]_  = ~A203 & ~A202;
  assign \new_[67624]_  = \new_[67623]_  & \new_[67620]_ ;
  assign \new_[67625]_  = \new_[67624]_  & \new_[67617]_ ;
  assign \new_[67628]_  = ~A233 & ~A232;
  assign \new_[67631]_  = A266 & A265;
  assign \new_[67632]_  = \new_[67631]_  & \new_[67628]_ ;
  assign \new_[67635]_  = ~A299 & A298;
  assign \new_[67638]_  = A301 & A300;
  assign \new_[67639]_  = \new_[67638]_  & \new_[67635]_ ;
  assign \new_[67640]_  = \new_[67639]_  & \new_[67632]_ ;
  assign \new_[67644]_  = ~A167 & A169;
  assign \new_[67645]_  = ~A170 & \new_[67644]_ ;
  assign \new_[67648]_  = ~A200 & ~A166;
  assign \new_[67651]_  = ~A203 & ~A202;
  assign \new_[67652]_  = \new_[67651]_  & \new_[67648]_ ;
  assign \new_[67653]_  = \new_[67652]_  & \new_[67645]_ ;
  assign \new_[67656]_  = ~A233 & ~A232;
  assign \new_[67659]_  = A266 & A265;
  assign \new_[67660]_  = \new_[67659]_  & \new_[67656]_ ;
  assign \new_[67663]_  = ~A299 & A298;
  assign \new_[67666]_  = A302 & A300;
  assign \new_[67667]_  = \new_[67666]_  & \new_[67663]_ ;
  assign \new_[67668]_  = \new_[67667]_  & \new_[67660]_ ;
  assign \new_[67672]_  = ~A167 & A169;
  assign \new_[67673]_  = ~A170 & \new_[67672]_ ;
  assign \new_[67676]_  = ~A200 & ~A166;
  assign \new_[67679]_  = ~A203 & ~A202;
  assign \new_[67680]_  = \new_[67679]_  & \new_[67676]_ ;
  assign \new_[67681]_  = \new_[67680]_  & \new_[67673]_ ;
  assign \new_[67684]_  = ~A233 & ~A232;
  assign \new_[67687]_  = ~A267 & ~A266;
  assign \new_[67688]_  = \new_[67687]_  & \new_[67684]_ ;
  assign \new_[67691]_  = ~A299 & A298;
  assign \new_[67694]_  = A301 & A300;
  assign \new_[67695]_  = \new_[67694]_  & \new_[67691]_ ;
  assign \new_[67696]_  = \new_[67695]_  & \new_[67688]_ ;
  assign \new_[67700]_  = ~A167 & A169;
  assign \new_[67701]_  = ~A170 & \new_[67700]_ ;
  assign \new_[67704]_  = ~A200 & ~A166;
  assign \new_[67707]_  = ~A203 & ~A202;
  assign \new_[67708]_  = \new_[67707]_  & \new_[67704]_ ;
  assign \new_[67709]_  = \new_[67708]_  & \new_[67701]_ ;
  assign \new_[67712]_  = ~A233 & ~A232;
  assign \new_[67715]_  = ~A267 & ~A266;
  assign \new_[67716]_  = \new_[67715]_  & \new_[67712]_ ;
  assign \new_[67719]_  = ~A299 & A298;
  assign \new_[67722]_  = A302 & A300;
  assign \new_[67723]_  = \new_[67722]_  & \new_[67719]_ ;
  assign \new_[67724]_  = \new_[67723]_  & \new_[67716]_ ;
  assign \new_[67728]_  = ~A167 & A169;
  assign \new_[67729]_  = ~A170 & \new_[67728]_ ;
  assign \new_[67732]_  = ~A200 & ~A166;
  assign \new_[67735]_  = ~A203 & ~A202;
  assign \new_[67736]_  = \new_[67735]_  & \new_[67732]_ ;
  assign \new_[67737]_  = \new_[67736]_  & \new_[67729]_ ;
  assign \new_[67740]_  = ~A233 & ~A232;
  assign \new_[67743]_  = ~A266 & ~A265;
  assign \new_[67744]_  = \new_[67743]_  & \new_[67740]_ ;
  assign \new_[67747]_  = ~A299 & A298;
  assign \new_[67750]_  = A301 & A300;
  assign \new_[67751]_  = \new_[67750]_  & \new_[67747]_ ;
  assign \new_[67752]_  = \new_[67751]_  & \new_[67744]_ ;
  assign \new_[67756]_  = ~A167 & A169;
  assign \new_[67757]_  = ~A170 & \new_[67756]_ ;
  assign \new_[67760]_  = ~A200 & ~A166;
  assign \new_[67763]_  = ~A203 & ~A202;
  assign \new_[67764]_  = \new_[67763]_  & \new_[67760]_ ;
  assign \new_[67765]_  = \new_[67764]_  & \new_[67757]_ ;
  assign \new_[67768]_  = ~A233 & ~A232;
  assign \new_[67771]_  = ~A266 & ~A265;
  assign \new_[67772]_  = \new_[67771]_  & \new_[67768]_ ;
  assign \new_[67775]_  = ~A299 & A298;
  assign \new_[67778]_  = A302 & A300;
  assign \new_[67779]_  = \new_[67778]_  & \new_[67775]_ ;
  assign \new_[67780]_  = \new_[67779]_  & \new_[67772]_ ;
  assign \new_[67784]_  = ~A167 & A169;
  assign \new_[67785]_  = ~A170 & \new_[67784]_ ;
  assign \new_[67788]_  = ~A200 & ~A166;
  assign \new_[67791]_  = A232 & ~A201;
  assign \new_[67792]_  = \new_[67791]_  & \new_[67788]_ ;
  assign \new_[67793]_  = \new_[67792]_  & \new_[67785]_ ;
  assign \new_[67796]_  = A265 & A233;
  assign \new_[67799]_  = ~A269 & ~A268;
  assign \new_[67800]_  = \new_[67799]_  & \new_[67796]_ ;
  assign \new_[67803]_  = ~A299 & A298;
  assign \new_[67806]_  = A301 & A300;
  assign \new_[67807]_  = \new_[67806]_  & \new_[67803]_ ;
  assign \new_[67808]_  = \new_[67807]_  & \new_[67800]_ ;
  assign \new_[67812]_  = ~A167 & A169;
  assign \new_[67813]_  = ~A170 & \new_[67812]_ ;
  assign \new_[67816]_  = ~A200 & ~A166;
  assign \new_[67819]_  = A232 & ~A201;
  assign \new_[67820]_  = \new_[67819]_  & \new_[67816]_ ;
  assign \new_[67821]_  = \new_[67820]_  & \new_[67813]_ ;
  assign \new_[67824]_  = A265 & A233;
  assign \new_[67827]_  = ~A269 & ~A268;
  assign \new_[67828]_  = \new_[67827]_  & \new_[67824]_ ;
  assign \new_[67831]_  = ~A299 & A298;
  assign \new_[67834]_  = A302 & A300;
  assign \new_[67835]_  = \new_[67834]_  & \new_[67831]_ ;
  assign \new_[67836]_  = \new_[67835]_  & \new_[67828]_ ;
  assign \new_[67840]_  = ~A167 & A169;
  assign \new_[67841]_  = ~A170 & \new_[67840]_ ;
  assign \new_[67844]_  = ~A200 & ~A166;
  assign \new_[67847]_  = ~A233 & ~A201;
  assign \new_[67848]_  = \new_[67847]_  & \new_[67844]_ ;
  assign \new_[67849]_  = \new_[67848]_  & \new_[67841]_ ;
  assign \new_[67852]_  = ~A236 & ~A235;
  assign \new_[67855]_  = A266 & A265;
  assign \new_[67856]_  = \new_[67855]_  & \new_[67852]_ ;
  assign \new_[67859]_  = ~A299 & A298;
  assign \new_[67862]_  = A301 & A300;
  assign \new_[67863]_  = \new_[67862]_  & \new_[67859]_ ;
  assign \new_[67864]_  = \new_[67863]_  & \new_[67856]_ ;
  assign \new_[67868]_  = ~A167 & A169;
  assign \new_[67869]_  = ~A170 & \new_[67868]_ ;
  assign \new_[67872]_  = ~A200 & ~A166;
  assign \new_[67875]_  = ~A233 & ~A201;
  assign \new_[67876]_  = \new_[67875]_  & \new_[67872]_ ;
  assign \new_[67877]_  = \new_[67876]_  & \new_[67869]_ ;
  assign \new_[67880]_  = ~A236 & ~A235;
  assign \new_[67883]_  = A266 & A265;
  assign \new_[67884]_  = \new_[67883]_  & \new_[67880]_ ;
  assign \new_[67887]_  = ~A299 & A298;
  assign \new_[67890]_  = A302 & A300;
  assign \new_[67891]_  = \new_[67890]_  & \new_[67887]_ ;
  assign \new_[67892]_  = \new_[67891]_  & \new_[67884]_ ;
  assign \new_[67896]_  = ~A167 & A169;
  assign \new_[67897]_  = ~A170 & \new_[67896]_ ;
  assign \new_[67900]_  = ~A200 & ~A166;
  assign \new_[67903]_  = ~A233 & ~A201;
  assign \new_[67904]_  = \new_[67903]_  & \new_[67900]_ ;
  assign \new_[67905]_  = \new_[67904]_  & \new_[67897]_ ;
  assign \new_[67908]_  = ~A236 & ~A235;
  assign \new_[67911]_  = ~A267 & ~A266;
  assign \new_[67912]_  = \new_[67911]_  & \new_[67908]_ ;
  assign \new_[67915]_  = ~A299 & A298;
  assign \new_[67918]_  = A301 & A300;
  assign \new_[67919]_  = \new_[67918]_  & \new_[67915]_ ;
  assign \new_[67920]_  = \new_[67919]_  & \new_[67912]_ ;
  assign \new_[67924]_  = ~A167 & A169;
  assign \new_[67925]_  = ~A170 & \new_[67924]_ ;
  assign \new_[67928]_  = ~A200 & ~A166;
  assign \new_[67931]_  = ~A233 & ~A201;
  assign \new_[67932]_  = \new_[67931]_  & \new_[67928]_ ;
  assign \new_[67933]_  = \new_[67932]_  & \new_[67925]_ ;
  assign \new_[67936]_  = ~A236 & ~A235;
  assign \new_[67939]_  = ~A267 & ~A266;
  assign \new_[67940]_  = \new_[67939]_  & \new_[67936]_ ;
  assign \new_[67943]_  = ~A299 & A298;
  assign \new_[67946]_  = A302 & A300;
  assign \new_[67947]_  = \new_[67946]_  & \new_[67943]_ ;
  assign \new_[67948]_  = \new_[67947]_  & \new_[67940]_ ;
  assign \new_[67952]_  = ~A167 & A169;
  assign \new_[67953]_  = ~A170 & \new_[67952]_ ;
  assign \new_[67956]_  = ~A200 & ~A166;
  assign \new_[67959]_  = ~A233 & ~A201;
  assign \new_[67960]_  = \new_[67959]_  & \new_[67956]_ ;
  assign \new_[67961]_  = \new_[67960]_  & \new_[67953]_ ;
  assign \new_[67964]_  = ~A236 & ~A235;
  assign \new_[67967]_  = ~A266 & ~A265;
  assign \new_[67968]_  = \new_[67967]_  & \new_[67964]_ ;
  assign \new_[67971]_  = ~A299 & A298;
  assign \new_[67974]_  = A301 & A300;
  assign \new_[67975]_  = \new_[67974]_  & \new_[67971]_ ;
  assign \new_[67976]_  = \new_[67975]_  & \new_[67968]_ ;
  assign \new_[67980]_  = ~A167 & A169;
  assign \new_[67981]_  = ~A170 & \new_[67980]_ ;
  assign \new_[67984]_  = ~A200 & ~A166;
  assign \new_[67987]_  = ~A233 & ~A201;
  assign \new_[67988]_  = \new_[67987]_  & \new_[67984]_ ;
  assign \new_[67989]_  = \new_[67988]_  & \new_[67981]_ ;
  assign \new_[67992]_  = ~A236 & ~A235;
  assign \new_[67995]_  = ~A266 & ~A265;
  assign \new_[67996]_  = \new_[67995]_  & \new_[67992]_ ;
  assign \new_[67999]_  = ~A299 & A298;
  assign \new_[68002]_  = A302 & A300;
  assign \new_[68003]_  = \new_[68002]_  & \new_[67999]_ ;
  assign \new_[68004]_  = \new_[68003]_  & \new_[67996]_ ;
  assign \new_[68008]_  = ~A167 & A169;
  assign \new_[68009]_  = ~A170 & \new_[68008]_ ;
  assign \new_[68012]_  = ~A200 & ~A166;
  assign \new_[68015]_  = ~A233 & ~A201;
  assign \new_[68016]_  = \new_[68015]_  & \new_[68012]_ ;
  assign \new_[68017]_  = \new_[68016]_  & \new_[68009]_ ;
  assign \new_[68020]_  = ~A266 & ~A234;
  assign \new_[68023]_  = ~A269 & ~A268;
  assign \new_[68024]_  = \new_[68023]_  & \new_[68020]_ ;
  assign \new_[68027]_  = ~A299 & A298;
  assign \new_[68030]_  = A301 & A300;
  assign \new_[68031]_  = \new_[68030]_  & \new_[68027]_ ;
  assign \new_[68032]_  = \new_[68031]_  & \new_[68024]_ ;
  assign \new_[68036]_  = ~A167 & A169;
  assign \new_[68037]_  = ~A170 & \new_[68036]_ ;
  assign \new_[68040]_  = ~A200 & ~A166;
  assign \new_[68043]_  = ~A233 & ~A201;
  assign \new_[68044]_  = \new_[68043]_  & \new_[68040]_ ;
  assign \new_[68045]_  = \new_[68044]_  & \new_[68037]_ ;
  assign \new_[68048]_  = ~A266 & ~A234;
  assign \new_[68051]_  = ~A269 & ~A268;
  assign \new_[68052]_  = \new_[68051]_  & \new_[68048]_ ;
  assign \new_[68055]_  = ~A299 & A298;
  assign \new_[68058]_  = A302 & A300;
  assign \new_[68059]_  = \new_[68058]_  & \new_[68055]_ ;
  assign \new_[68060]_  = \new_[68059]_  & \new_[68052]_ ;
  assign \new_[68064]_  = ~A167 & A169;
  assign \new_[68065]_  = ~A170 & \new_[68064]_ ;
  assign \new_[68068]_  = ~A200 & ~A166;
  assign \new_[68071]_  = ~A232 & ~A201;
  assign \new_[68072]_  = \new_[68071]_  & \new_[68068]_ ;
  assign \new_[68073]_  = \new_[68072]_  & \new_[68065]_ ;
  assign \new_[68076]_  = ~A266 & ~A233;
  assign \new_[68079]_  = ~A269 & ~A268;
  assign \new_[68080]_  = \new_[68079]_  & \new_[68076]_ ;
  assign \new_[68083]_  = ~A299 & A298;
  assign \new_[68086]_  = A301 & A300;
  assign \new_[68087]_  = \new_[68086]_  & \new_[68083]_ ;
  assign \new_[68088]_  = \new_[68087]_  & \new_[68080]_ ;
  assign \new_[68092]_  = ~A167 & A169;
  assign \new_[68093]_  = ~A170 & \new_[68092]_ ;
  assign \new_[68096]_  = ~A200 & ~A166;
  assign \new_[68099]_  = ~A232 & ~A201;
  assign \new_[68100]_  = \new_[68099]_  & \new_[68096]_ ;
  assign \new_[68101]_  = \new_[68100]_  & \new_[68093]_ ;
  assign \new_[68104]_  = ~A266 & ~A233;
  assign \new_[68107]_  = ~A269 & ~A268;
  assign \new_[68108]_  = \new_[68107]_  & \new_[68104]_ ;
  assign \new_[68111]_  = ~A299 & A298;
  assign \new_[68114]_  = A302 & A300;
  assign \new_[68115]_  = \new_[68114]_  & \new_[68111]_ ;
  assign \new_[68116]_  = \new_[68115]_  & \new_[68108]_ ;
  assign \new_[68120]_  = ~A167 & A169;
  assign \new_[68121]_  = ~A170 & \new_[68120]_ ;
  assign \new_[68124]_  = ~A199 & ~A166;
  assign \new_[68127]_  = A232 & ~A200;
  assign \new_[68128]_  = \new_[68127]_  & \new_[68124]_ ;
  assign \new_[68129]_  = \new_[68128]_  & \new_[68121]_ ;
  assign \new_[68132]_  = A265 & A233;
  assign \new_[68135]_  = ~A269 & ~A268;
  assign \new_[68136]_  = \new_[68135]_  & \new_[68132]_ ;
  assign \new_[68139]_  = ~A299 & A298;
  assign \new_[68142]_  = A301 & A300;
  assign \new_[68143]_  = \new_[68142]_  & \new_[68139]_ ;
  assign \new_[68144]_  = \new_[68143]_  & \new_[68136]_ ;
  assign \new_[68148]_  = ~A167 & A169;
  assign \new_[68149]_  = ~A170 & \new_[68148]_ ;
  assign \new_[68152]_  = ~A199 & ~A166;
  assign \new_[68155]_  = A232 & ~A200;
  assign \new_[68156]_  = \new_[68155]_  & \new_[68152]_ ;
  assign \new_[68157]_  = \new_[68156]_  & \new_[68149]_ ;
  assign \new_[68160]_  = A265 & A233;
  assign \new_[68163]_  = ~A269 & ~A268;
  assign \new_[68164]_  = \new_[68163]_  & \new_[68160]_ ;
  assign \new_[68167]_  = ~A299 & A298;
  assign \new_[68170]_  = A302 & A300;
  assign \new_[68171]_  = \new_[68170]_  & \new_[68167]_ ;
  assign \new_[68172]_  = \new_[68171]_  & \new_[68164]_ ;
  assign \new_[68176]_  = ~A167 & A169;
  assign \new_[68177]_  = ~A170 & \new_[68176]_ ;
  assign \new_[68180]_  = ~A199 & ~A166;
  assign \new_[68183]_  = ~A233 & ~A200;
  assign \new_[68184]_  = \new_[68183]_  & \new_[68180]_ ;
  assign \new_[68185]_  = \new_[68184]_  & \new_[68177]_ ;
  assign \new_[68188]_  = ~A236 & ~A235;
  assign \new_[68191]_  = A266 & A265;
  assign \new_[68192]_  = \new_[68191]_  & \new_[68188]_ ;
  assign \new_[68195]_  = ~A299 & A298;
  assign \new_[68198]_  = A301 & A300;
  assign \new_[68199]_  = \new_[68198]_  & \new_[68195]_ ;
  assign \new_[68200]_  = \new_[68199]_  & \new_[68192]_ ;
  assign \new_[68204]_  = ~A167 & A169;
  assign \new_[68205]_  = ~A170 & \new_[68204]_ ;
  assign \new_[68208]_  = ~A199 & ~A166;
  assign \new_[68211]_  = ~A233 & ~A200;
  assign \new_[68212]_  = \new_[68211]_  & \new_[68208]_ ;
  assign \new_[68213]_  = \new_[68212]_  & \new_[68205]_ ;
  assign \new_[68216]_  = ~A236 & ~A235;
  assign \new_[68219]_  = A266 & A265;
  assign \new_[68220]_  = \new_[68219]_  & \new_[68216]_ ;
  assign \new_[68223]_  = ~A299 & A298;
  assign \new_[68226]_  = A302 & A300;
  assign \new_[68227]_  = \new_[68226]_  & \new_[68223]_ ;
  assign \new_[68228]_  = \new_[68227]_  & \new_[68220]_ ;
  assign \new_[68232]_  = ~A167 & A169;
  assign \new_[68233]_  = ~A170 & \new_[68232]_ ;
  assign \new_[68236]_  = ~A199 & ~A166;
  assign \new_[68239]_  = ~A233 & ~A200;
  assign \new_[68240]_  = \new_[68239]_  & \new_[68236]_ ;
  assign \new_[68241]_  = \new_[68240]_  & \new_[68233]_ ;
  assign \new_[68244]_  = ~A236 & ~A235;
  assign \new_[68247]_  = ~A267 & ~A266;
  assign \new_[68248]_  = \new_[68247]_  & \new_[68244]_ ;
  assign \new_[68251]_  = ~A299 & A298;
  assign \new_[68254]_  = A301 & A300;
  assign \new_[68255]_  = \new_[68254]_  & \new_[68251]_ ;
  assign \new_[68256]_  = \new_[68255]_  & \new_[68248]_ ;
  assign \new_[68260]_  = ~A167 & A169;
  assign \new_[68261]_  = ~A170 & \new_[68260]_ ;
  assign \new_[68264]_  = ~A199 & ~A166;
  assign \new_[68267]_  = ~A233 & ~A200;
  assign \new_[68268]_  = \new_[68267]_  & \new_[68264]_ ;
  assign \new_[68269]_  = \new_[68268]_  & \new_[68261]_ ;
  assign \new_[68272]_  = ~A236 & ~A235;
  assign \new_[68275]_  = ~A267 & ~A266;
  assign \new_[68276]_  = \new_[68275]_  & \new_[68272]_ ;
  assign \new_[68279]_  = ~A299 & A298;
  assign \new_[68282]_  = A302 & A300;
  assign \new_[68283]_  = \new_[68282]_  & \new_[68279]_ ;
  assign \new_[68284]_  = \new_[68283]_  & \new_[68276]_ ;
  assign \new_[68288]_  = ~A167 & A169;
  assign \new_[68289]_  = ~A170 & \new_[68288]_ ;
  assign \new_[68292]_  = ~A199 & ~A166;
  assign \new_[68295]_  = ~A233 & ~A200;
  assign \new_[68296]_  = \new_[68295]_  & \new_[68292]_ ;
  assign \new_[68297]_  = \new_[68296]_  & \new_[68289]_ ;
  assign \new_[68300]_  = ~A236 & ~A235;
  assign \new_[68303]_  = ~A266 & ~A265;
  assign \new_[68304]_  = \new_[68303]_  & \new_[68300]_ ;
  assign \new_[68307]_  = ~A299 & A298;
  assign \new_[68310]_  = A301 & A300;
  assign \new_[68311]_  = \new_[68310]_  & \new_[68307]_ ;
  assign \new_[68312]_  = \new_[68311]_  & \new_[68304]_ ;
  assign \new_[68316]_  = ~A167 & A169;
  assign \new_[68317]_  = ~A170 & \new_[68316]_ ;
  assign \new_[68320]_  = ~A199 & ~A166;
  assign \new_[68323]_  = ~A233 & ~A200;
  assign \new_[68324]_  = \new_[68323]_  & \new_[68320]_ ;
  assign \new_[68325]_  = \new_[68324]_  & \new_[68317]_ ;
  assign \new_[68328]_  = ~A236 & ~A235;
  assign \new_[68331]_  = ~A266 & ~A265;
  assign \new_[68332]_  = \new_[68331]_  & \new_[68328]_ ;
  assign \new_[68335]_  = ~A299 & A298;
  assign \new_[68338]_  = A302 & A300;
  assign \new_[68339]_  = \new_[68338]_  & \new_[68335]_ ;
  assign \new_[68340]_  = \new_[68339]_  & \new_[68332]_ ;
  assign \new_[68344]_  = ~A167 & A169;
  assign \new_[68345]_  = ~A170 & \new_[68344]_ ;
  assign \new_[68348]_  = ~A199 & ~A166;
  assign \new_[68351]_  = ~A233 & ~A200;
  assign \new_[68352]_  = \new_[68351]_  & \new_[68348]_ ;
  assign \new_[68353]_  = \new_[68352]_  & \new_[68345]_ ;
  assign \new_[68356]_  = ~A266 & ~A234;
  assign \new_[68359]_  = ~A269 & ~A268;
  assign \new_[68360]_  = \new_[68359]_  & \new_[68356]_ ;
  assign \new_[68363]_  = ~A299 & A298;
  assign \new_[68366]_  = A301 & A300;
  assign \new_[68367]_  = \new_[68366]_  & \new_[68363]_ ;
  assign \new_[68368]_  = \new_[68367]_  & \new_[68360]_ ;
  assign \new_[68372]_  = ~A167 & A169;
  assign \new_[68373]_  = ~A170 & \new_[68372]_ ;
  assign \new_[68376]_  = ~A199 & ~A166;
  assign \new_[68379]_  = ~A233 & ~A200;
  assign \new_[68380]_  = \new_[68379]_  & \new_[68376]_ ;
  assign \new_[68381]_  = \new_[68380]_  & \new_[68373]_ ;
  assign \new_[68384]_  = ~A266 & ~A234;
  assign \new_[68387]_  = ~A269 & ~A268;
  assign \new_[68388]_  = \new_[68387]_  & \new_[68384]_ ;
  assign \new_[68391]_  = ~A299 & A298;
  assign \new_[68394]_  = A302 & A300;
  assign \new_[68395]_  = \new_[68394]_  & \new_[68391]_ ;
  assign \new_[68396]_  = \new_[68395]_  & \new_[68388]_ ;
  assign \new_[68400]_  = ~A167 & A169;
  assign \new_[68401]_  = ~A170 & \new_[68400]_ ;
  assign \new_[68404]_  = ~A199 & ~A166;
  assign \new_[68407]_  = ~A232 & ~A200;
  assign \new_[68408]_  = \new_[68407]_  & \new_[68404]_ ;
  assign \new_[68409]_  = \new_[68408]_  & \new_[68401]_ ;
  assign \new_[68412]_  = ~A266 & ~A233;
  assign \new_[68415]_  = ~A269 & ~A268;
  assign \new_[68416]_  = \new_[68415]_  & \new_[68412]_ ;
  assign \new_[68419]_  = ~A299 & A298;
  assign \new_[68422]_  = A301 & A300;
  assign \new_[68423]_  = \new_[68422]_  & \new_[68419]_ ;
  assign \new_[68424]_  = \new_[68423]_  & \new_[68416]_ ;
  assign \new_[68428]_  = ~A167 & A169;
  assign \new_[68429]_  = ~A170 & \new_[68428]_ ;
  assign \new_[68432]_  = ~A199 & ~A166;
  assign \new_[68435]_  = ~A232 & ~A200;
  assign \new_[68436]_  = \new_[68435]_  & \new_[68432]_ ;
  assign \new_[68437]_  = \new_[68436]_  & \new_[68429]_ ;
  assign \new_[68440]_  = ~A266 & ~A233;
  assign \new_[68443]_  = ~A269 & ~A268;
  assign \new_[68444]_  = \new_[68443]_  & \new_[68440]_ ;
  assign \new_[68447]_  = ~A299 & A298;
  assign \new_[68450]_  = A302 & A300;
  assign \new_[68451]_  = \new_[68450]_  & \new_[68447]_ ;
  assign \new_[68452]_  = \new_[68451]_  & \new_[68444]_ ;
  assign \new_[68456]_  = ~A166 & ~A167;
  assign \new_[68457]_  = ~A169 & \new_[68456]_ ;
  assign \new_[68460]_  = A200 & ~A199;
  assign \new_[68463]_  = ~A235 & ~A233;
  assign \new_[68464]_  = \new_[68463]_  & \new_[68460]_ ;
  assign \new_[68465]_  = \new_[68464]_  & \new_[68457]_ ;
  assign \new_[68468]_  = ~A266 & ~A236;
  assign \new_[68471]_  = ~A269 & ~A268;
  assign \new_[68472]_  = \new_[68471]_  & \new_[68468]_ ;
  assign \new_[68475]_  = ~A299 & A298;
  assign \new_[68478]_  = A301 & A300;
  assign \new_[68479]_  = \new_[68478]_  & \new_[68475]_ ;
  assign \new_[68480]_  = \new_[68479]_  & \new_[68472]_ ;
  assign \new_[68484]_  = ~A166 & ~A167;
  assign \new_[68485]_  = ~A169 & \new_[68484]_ ;
  assign \new_[68488]_  = A200 & ~A199;
  assign \new_[68491]_  = ~A235 & ~A233;
  assign \new_[68492]_  = \new_[68491]_  & \new_[68488]_ ;
  assign \new_[68493]_  = \new_[68492]_  & \new_[68485]_ ;
  assign \new_[68496]_  = ~A266 & ~A236;
  assign \new_[68499]_  = ~A269 & ~A268;
  assign \new_[68500]_  = \new_[68499]_  & \new_[68496]_ ;
  assign \new_[68503]_  = ~A299 & A298;
  assign \new_[68506]_  = A302 & A300;
  assign \new_[68507]_  = \new_[68506]_  & \new_[68503]_ ;
  assign \new_[68508]_  = \new_[68507]_  & \new_[68500]_ ;
  assign \new_[68512]_  = ~A166 & ~A167;
  assign \new_[68513]_  = ~A169 & \new_[68512]_ ;
  assign \new_[68516]_  = ~A200 & A199;
  assign \new_[68519]_  = A202 & A201;
  assign \new_[68520]_  = \new_[68519]_  & \new_[68516]_ ;
  assign \new_[68521]_  = \new_[68520]_  & \new_[68513]_ ;
  assign \new_[68524]_  = A233 & A232;
  assign \new_[68527]_  = ~A267 & A265;
  assign \new_[68528]_  = \new_[68527]_  & \new_[68524]_ ;
  assign \new_[68531]_  = ~A299 & A298;
  assign \new_[68534]_  = A301 & A300;
  assign \new_[68535]_  = \new_[68534]_  & \new_[68531]_ ;
  assign \new_[68536]_  = \new_[68535]_  & \new_[68528]_ ;
  assign \new_[68540]_  = ~A166 & ~A167;
  assign \new_[68541]_  = ~A169 & \new_[68540]_ ;
  assign \new_[68544]_  = ~A200 & A199;
  assign \new_[68547]_  = A202 & A201;
  assign \new_[68548]_  = \new_[68547]_  & \new_[68544]_ ;
  assign \new_[68549]_  = \new_[68548]_  & \new_[68541]_ ;
  assign \new_[68552]_  = A233 & A232;
  assign \new_[68555]_  = ~A267 & A265;
  assign \new_[68556]_  = \new_[68555]_  & \new_[68552]_ ;
  assign \new_[68559]_  = ~A299 & A298;
  assign \new_[68562]_  = A302 & A300;
  assign \new_[68563]_  = \new_[68562]_  & \new_[68559]_ ;
  assign \new_[68564]_  = \new_[68563]_  & \new_[68556]_ ;
  assign \new_[68568]_  = ~A166 & ~A167;
  assign \new_[68569]_  = ~A169 & \new_[68568]_ ;
  assign \new_[68572]_  = ~A200 & A199;
  assign \new_[68575]_  = A202 & A201;
  assign \new_[68576]_  = \new_[68575]_  & \new_[68572]_ ;
  assign \new_[68577]_  = \new_[68576]_  & \new_[68569]_ ;
  assign \new_[68580]_  = A233 & A232;
  assign \new_[68583]_  = A266 & A265;
  assign \new_[68584]_  = \new_[68583]_  & \new_[68580]_ ;
  assign \new_[68587]_  = ~A299 & A298;
  assign \new_[68590]_  = A301 & A300;
  assign \new_[68591]_  = \new_[68590]_  & \new_[68587]_ ;
  assign \new_[68592]_  = \new_[68591]_  & \new_[68584]_ ;
  assign \new_[68596]_  = ~A166 & ~A167;
  assign \new_[68597]_  = ~A169 & \new_[68596]_ ;
  assign \new_[68600]_  = ~A200 & A199;
  assign \new_[68603]_  = A202 & A201;
  assign \new_[68604]_  = \new_[68603]_  & \new_[68600]_ ;
  assign \new_[68605]_  = \new_[68604]_  & \new_[68597]_ ;
  assign \new_[68608]_  = A233 & A232;
  assign \new_[68611]_  = A266 & A265;
  assign \new_[68612]_  = \new_[68611]_  & \new_[68608]_ ;
  assign \new_[68615]_  = ~A299 & A298;
  assign \new_[68618]_  = A302 & A300;
  assign \new_[68619]_  = \new_[68618]_  & \new_[68615]_ ;
  assign \new_[68620]_  = \new_[68619]_  & \new_[68612]_ ;
  assign \new_[68624]_  = ~A166 & ~A167;
  assign \new_[68625]_  = ~A169 & \new_[68624]_ ;
  assign \new_[68628]_  = ~A200 & A199;
  assign \new_[68631]_  = A202 & A201;
  assign \new_[68632]_  = \new_[68631]_  & \new_[68628]_ ;
  assign \new_[68633]_  = \new_[68632]_  & \new_[68625]_ ;
  assign \new_[68636]_  = A233 & A232;
  assign \new_[68639]_  = ~A266 & ~A265;
  assign \new_[68640]_  = \new_[68639]_  & \new_[68636]_ ;
  assign \new_[68643]_  = ~A299 & A298;
  assign \new_[68646]_  = A301 & A300;
  assign \new_[68647]_  = \new_[68646]_  & \new_[68643]_ ;
  assign \new_[68648]_  = \new_[68647]_  & \new_[68640]_ ;
  assign \new_[68652]_  = ~A166 & ~A167;
  assign \new_[68653]_  = ~A169 & \new_[68652]_ ;
  assign \new_[68656]_  = ~A200 & A199;
  assign \new_[68659]_  = A202 & A201;
  assign \new_[68660]_  = \new_[68659]_  & \new_[68656]_ ;
  assign \new_[68661]_  = \new_[68660]_  & \new_[68653]_ ;
  assign \new_[68664]_  = A233 & A232;
  assign \new_[68667]_  = ~A266 & ~A265;
  assign \new_[68668]_  = \new_[68667]_  & \new_[68664]_ ;
  assign \new_[68671]_  = ~A299 & A298;
  assign \new_[68674]_  = A302 & A300;
  assign \new_[68675]_  = \new_[68674]_  & \new_[68671]_ ;
  assign \new_[68676]_  = \new_[68675]_  & \new_[68668]_ ;
  assign \new_[68680]_  = ~A166 & ~A167;
  assign \new_[68681]_  = ~A169 & \new_[68680]_ ;
  assign \new_[68684]_  = ~A200 & A199;
  assign \new_[68687]_  = A202 & A201;
  assign \new_[68688]_  = \new_[68687]_  & \new_[68684]_ ;
  assign \new_[68689]_  = \new_[68688]_  & \new_[68681]_ ;
  assign \new_[68692]_  = ~A235 & ~A233;
  assign \new_[68695]_  = ~A266 & ~A236;
  assign \new_[68696]_  = \new_[68695]_  & \new_[68692]_ ;
  assign \new_[68699]_  = ~A269 & ~A268;
  assign \new_[68702]_  = A299 & ~A298;
  assign \new_[68703]_  = \new_[68702]_  & \new_[68699]_ ;
  assign \new_[68704]_  = \new_[68703]_  & \new_[68696]_ ;
  assign \new_[68708]_  = ~A166 & ~A167;
  assign \new_[68709]_  = ~A169 & \new_[68708]_ ;
  assign \new_[68712]_  = ~A200 & A199;
  assign \new_[68715]_  = A202 & A201;
  assign \new_[68716]_  = \new_[68715]_  & \new_[68712]_ ;
  assign \new_[68717]_  = \new_[68716]_  & \new_[68709]_ ;
  assign \new_[68720]_  = ~A234 & ~A233;
  assign \new_[68723]_  = A266 & A265;
  assign \new_[68724]_  = \new_[68723]_  & \new_[68720]_ ;
  assign \new_[68727]_  = ~A299 & A298;
  assign \new_[68730]_  = A301 & A300;
  assign \new_[68731]_  = \new_[68730]_  & \new_[68727]_ ;
  assign \new_[68732]_  = \new_[68731]_  & \new_[68724]_ ;
  assign \new_[68736]_  = ~A166 & ~A167;
  assign \new_[68737]_  = ~A169 & \new_[68736]_ ;
  assign \new_[68740]_  = ~A200 & A199;
  assign \new_[68743]_  = A202 & A201;
  assign \new_[68744]_  = \new_[68743]_  & \new_[68740]_ ;
  assign \new_[68745]_  = \new_[68744]_  & \new_[68737]_ ;
  assign \new_[68748]_  = ~A234 & ~A233;
  assign \new_[68751]_  = A266 & A265;
  assign \new_[68752]_  = \new_[68751]_  & \new_[68748]_ ;
  assign \new_[68755]_  = ~A299 & A298;
  assign \new_[68758]_  = A302 & A300;
  assign \new_[68759]_  = \new_[68758]_  & \new_[68755]_ ;
  assign \new_[68760]_  = \new_[68759]_  & \new_[68752]_ ;
  assign \new_[68764]_  = ~A166 & ~A167;
  assign \new_[68765]_  = ~A169 & \new_[68764]_ ;
  assign \new_[68768]_  = ~A200 & A199;
  assign \new_[68771]_  = A202 & A201;
  assign \new_[68772]_  = \new_[68771]_  & \new_[68768]_ ;
  assign \new_[68773]_  = \new_[68772]_  & \new_[68765]_ ;
  assign \new_[68776]_  = ~A234 & ~A233;
  assign \new_[68779]_  = ~A267 & ~A266;
  assign \new_[68780]_  = \new_[68779]_  & \new_[68776]_ ;
  assign \new_[68783]_  = ~A299 & A298;
  assign \new_[68786]_  = A301 & A300;
  assign \new_[68787]_  = \new_[68786]_  & \new_[68783]_ ;
  assign \new_[68788]_  = \new_[68787]_  & \new_[68780]_ ;
  assign \new_[68792]_  = ~A166 & ~A167;
  assign \new_[68793]_  = ~A169 & \new_[68792]_ ;
  assign \new_[68796]_  = ~A200 & A199;
  assign \new_[68799]_  = A202 & A201;
  assign \new_[68800]_  = \new_[68799]_  & \new_[68796]_ ;
  assign \new_[68801]_  = \new_[68800]_  & \new_[68793]_ ;
  assign \new_[68804]_  = ~A234 & ~A233;
  assign \new_[68807]_  = ~A267 & ~A266;
  assign \new_[68808]_  = \new_[68807]_  & \new_[68804]_ ;
  assign \new_[68811]_  = ~A299 & A298;
  assign \new_[68814]_  = A302 & A300;
  assign \new_[68815]_  = \new_[68814]_  & \new_[68811]_ ;
  assign \new_[68816]_  = \new_[68815]_  & \new_[68808]_ ;
  assign \new_[68820]_  = ~A166 & ~A167;
  assign \new_[68821]_  = ~A169 & \new_[68820]_ ;
  assign \new_[68824]_  = ~A200 & A199;
  assign \new_[68827]_  = A202 & A201;
  assign \new_[68828]_  = \new_[68827]_  & \new_[68824]_ ;
  assign \new_[68829]_  = \new_[68828]_  & \new_[68821]_ ;
  assign \new_[68832]_  = ~A234 & ~A233;
  assign \new_[68835]_  = ~A266 & ~A265;
  assign \new_[68836]_  = \new_[68835]_  & \new_[68832]_ ;
  assign \new_[68839]_  = ~A299 & A298;
  assign \new_[68842]_  = A301 & A300;
  assign \new_[68843]_  = \new_[68842]_  & \new_[68839]_ ;
  assign \new_[68844]_  = \new_[68843]_  & \new_[68836]_ ;
  assign \new_[68848]_  = ~A166 & ~A167;
  assign \new_[68849]_  = ~A169 & \new_[68848]_ ;
  assign \new_[68852]_  = ~A200 & A199;
  assign \new_[68855]_  = A202 & A201;
  assign \new_[68856]_  = \new_[68855]_  & \new_[68852]_ ;
  assign \new_[68857]_  = \new_[68856]_  & \new_[68849]_ ;
  assign \new_[68860]_  = ~A234 & ~A233;
  assign \new_[68863]_  = ~A266 & ~A265;
  assign \new_[68864]_  = \new_[68863]_  & \new_[68860]_ ;
  assign \new_[68867]_  = ~A299 & A298;
  assign \new_[68870]_  = A302 & A300;
  assign \new_[68871]_  = \new_[68870]_  & \new_[68867]_ ;
  assign \new_[68872]_  = \new_[68871]_  & \new_[68864]_ ;
  assign \new_[68876]_  = ~A166 & ~A167;
  assign \new_[68877]_  = ~A169 & \new_[68876]_ ;
  assign \new_[68880]_  = ~A200 & A199;
  assign \new_[68883]_  = A202 & A201;
  assign \new_[68884]_  = \new_[68883]_  & \new_[68880]_ ;
  assign \new_[68885]_  = \new_[68884]_  & \new_[68877]_ ;
  assign \new_[68888]_  = ~A233 & A232;
  assign \new_[68891]_  = A235 & A234;
  assign \new_[68892]_  = \new_[68891]_  & \new_[68888]_ ;
  assign \new_[68895]_  = ~A266 & A265;
  assign \new_[68898]_  = A268 & A267;
  assign \new_[68899]_  = \new_[68898]_  & \new_[68895]_ ;
  assign \new_[68900]_  = \new_[68899]_  & \new_[68892]_ ;
  assign \new_[68904]_  = ~A166 & ~A167;
  assign \new_[68905]_  = ~A169 & \new_[68904]_ ;
  assign \new_[68908]_  = ~A200 & A199;
  assign \new_[68911]_  = A202 & A201;
  assign \new_[68912]_  = \new_[68911]_  & \new_[68908]_ ;
  assign \new_[68913]_  = \new_[68912]_  & \new_[68905]_ ;
  assign \new_[68916]_  = ~A233 & A232;
  assign \new_[68919]_  = A235 & A234;
  assign \new_[68920]_  = \new_[68919]_  & \new_[68916]_ ;
  assign \new_[68923]_  = ~A266 & A265;
  assign \new_[68926]_  = A269 & A267;
  assign \new_[68927]_  = \new_[68926]_  & \new_[68923]_ ;
  assign \new_[68928]_  = \new_[68927]_  & \new_[68920]_ ;
  assign \new_[68932]_  = ~A166 & ~A167;
  assign \new_[68933]_  = ~A169 & \new_[68932]_ ;
  assign \new_[68936]_  = ~A200 & A199;
  assign \new_[68939]_  = A202 & A201;
  assign \new_[68940]_  = \new_[68939]_  & \new_[68936]_ ;
  assign \new_[68941]_  = \new_[68940]_  & \new_[68933]_ ;
  assign \new_[68944]_  = ~A233 & A232;
  assign \new_[68947]_  = A236 & A234;
  assign \new_[68948]_  = \new_[68947]_  & \new_[68944]_ ;
  assign \new_[68951]_  = ~A266 & A265;
  assign \new_[68954]_  = A268 & A267;
  assign \new_[68955]_  = \new_[68954]_  & \new_[68951]_ ;
  assign \new_[68956]_  = \new_[68955]_  & \new_[68948]_ ;
  assign \new_[68960]_  = ~A166 & ~A167;
  assign \new_[68961]_  = ~A169 & \new_[68960]_ ;
  assign \new_[68964]_  = ~A200 & A199;
  assign \new_[68967]_  = A202 & A201;
  assign \new_[68968]_  = \new_[68967]_  & \new_[68964]_ ;
  assign \new_[68969]_  = \new_[68968]_  & \new_[68961]_ ;
  assign \new_[68972]_  = ~A233 & A232;
  assign \new_[68975]_  = A236 & A234;
  assign \new_[68976]_  = \new_[68975]_  & \new_[68972]_ ;
  assign \new_[68979]_  = ~A266 & A265;
  assign \new_[68982]_  = A269 & A267;
  assign \new_[68983]_  = \new_[68982]_  & \new_[68979]_ ;
  assign \new_[68984]_  = \new_[68983]_  & \new_[68976]_ ;
  assign \new_[68988]_  = ~A166 & ~A167;
  assign \new_[68989]_  = ~A169 & \new_[68988]_ ;
  assign \new_[68992]_  = ~A200 & A199;
  assign \new_[68995]_  = A202 & A201;
  assign \new_[68996]_  = \new_[68995]_  & \new_[68992]_ ;
  assign \new_[68997]_  = \new_[68996]_  & \new_[68989]_ ;
  assign \new_[69000]_  = ~A233 & ~A232;
  assign \new_[69003]_  = A266 & A265;
  assign \new_[69004]_  = \new_[69003]_  & \new_[69000]_ ;
  assign \new_[69007]_  = ~A299 & A298;
  assign \new_[69010]_  = A301 & A300;
  assign \new_[69011]_  = \new_[69010]_  & \new_[69007]_ ;
  assign \new_[69012]_  = \new_[69011]_  & \new_[69004]_ ;
  assign \new_[69016]_  = ~A166 & ~A167;
  assign \new_[69017]_  = ~A169 & \new_[69016]_ ;
  assign \new_[69020]_  = ~A200 & A199;
  assign \new_[69023]_  = A202 & A201;
  assign \new_[69024]_  = \new_[69023]_  & \new_[69020]_ ;
  assign \new_[69025]_  = \new_[69024]_  & \new_[69017]_ ;
  assign \new_[69028]_  = ~A233 & ~A232;
  assign \new_[69031]_  = A266 & A265;
  assign \new_[69032]_  = \new_[69031]_  & \new_[69028]_ ;
  assign \new_[69035]_  = ~A299 & A298;
  assign \new_[69038]_  = A302 & A300;
  assign \new_[69039]_  = \new_[69038]_  & \new_[69035]_ ;
  assign \new_[69040]_  = \new_[69039]_  & \new_[69032]_ ;
  assign \new_[69044]_  = ~A166 & ~A167;
  assign \new_[69045]_  = ~A169 & \new_[69044]_ ;
  assign \new_[69048]_  = ~A200 & A199;
  assign \new_[69051]_  = A202 & A201;
  assign \new_[69052]_  = \new_[69051]_  & \new_[69048]_ ;
  assign \new_[69053]_  = \new_[69052]_  & \new_[69045]_ ;
  assign \new_[69056]_  = ~A233 & ~A232;
  assign \new_[69059]_  = ~A267 & ~A266;
  assign \new_[69060]_  = \new_[69059]_  & \new_[69056]_ ;
  assign \new_[69063]_  = ~A299 & A298;
  assign \new_[69066]_  = A301 & A300;
  assign \new_[69067]_  = \new_[69066]_  & \new_[69063]_ ;
  assign \new_[69068]_  = \new_[69067]_  & \new_[69060]_ ;
  assign \new_[69072]_  = ~A166 & ~A167;
  assign \new_[69073]_  = ~A169 & \new_[69072]_ ;
  assign \new_[69076]_  = ~A200 & A199;
  assign \new_[69079]_  = A202 & A201;
  assign \new_[69080]_  = \new_[69079]_  & \new_[69076]_ ;
  assign \new_[69081]_  = \new_[69080]_  & \new_[69073]_ ;
  assign \new_[69084]_  = ~A233 & ~A232;
  assign \new_[69087]_  = ~A267 & ~A266;
  assign \new_[69088]_  = \new_[69087]_  & \new_[69084]_ ;
  assign \new_[69091]_  = ~A299 & A298;
  assign \new_[69094]_  = A302 & A300;
  assign \new_[69095]_  = \new_[69094]_  & \new_[69091]_ ;
  assign \new_[69096]_  = \new_[69095]_  & \new_[69088]_ ;
  assign \new_[69100]_  = ~A166 & ~A167;
  assign \new_[69101]_  = ~A169 & \new_[69100]_ ;
  assign \new_[69104]_  = ~A200 & A199;
  assign \new_[69107]_  = A202 & A201;
  assign \new_[69108]_  = \new_[69107]_  & \new_[69104]_ ;
  assign \new_[69109]_  = \new_[69108]_  & \new_[69101]_ ;
  assign \new_[69112]_  = ~A233 & ~A232;
  assign \new_[69115]_  = ~A266 & ~A265;
  assign \new_[69116]_  = \new_[69115]_  & \new_[69112]_ ;
  assign \new_[69119]_  = ~A299 & A298;
  assign \new_[69122]_  = A301 & A300;
  assign \new_[69123]_  = \new_[69122]_  & \new_[69119]_ ;
  assign \new_[69124]_  = \new_[69123]_  & \new_[69116]_ ;
  assign \new_[69128]_  = ~A166 & ~A167;
  assign \new_[69129]_  = ~A169 & \new_[69128]_ ;
  assign \new_[69132]_  = ~A200 & A199;
  assign \new_[69135]_  = A202 & A201;
  assign \new_[69136]_  = \new_[69135]_  & \new_[69132]_ ;
  assign \new_[69137]_  = \new_[69136]_  & \new_[69129]_ ;
  assign \new_[69140]_  = ~A233 & ~A232;
  assign \new_[69143]_  = ~A266 & ~A265;
  assign \new_[69144]_  = \new_[69143]_  & \new_[69140]_ ;
  assign \new_[69147]_  = ~A299 & A298;
  assign \new_[69150]_  = A302 & A300;
  assign \new_[69151]_  = \new_[69150]_  & \new_[69147]_ ;
  assign \new_[69152]_  = \new_[69151]_  & \new_[69144]_ ;
  assign \new_[69156]_  = ~A166 & ~A167;
  assign \new_[69157]_  = ~A169 & \new_[69156]_ ;
  assign \new_[69160]_  = ~A200 & A199;
  assign \new_[69163]_  = A203 & A201;
  assign \new_[69164]_  = \new_[69163]_  & \new_[69160]_ ;
  assign \new_[69165]_  = \new_[69164]_  & \new_[69157]_ ;
  assign \new_[69168]_  = A233 & A232;
  assign \new_[69171]_  = ~A267 & A265;
  assign \new_[69172]_  = \new_[69171]_  & \new_[69168]_ ;
  assign \new_[69175]_  = ~A299 & A298;
  assign \new_[69178]_  = A301 & A300;
  assign \new_[69179]_  = \new_[69178]_  & \new_[69175]_ ;
  assign \new_[69180]_  = \new_[69179]_  & \new_[69172]_ ;
  assign \new_[69184]_  = ~A166 & ~A167;
  assign \new_[69185]_  = ~A169 & \new_[69184]_ ;
  assign \new_[69188]_  = ~A200 & A199;
  assign \new_[69191]_  = A203 & A201;
  assign \new_[69192]_  = \new_[69191]_  & \new_[69188]_ ;
  assign \new_[69193]_  = \new_[69192]_  & \new_[69185]_ ;
  assign \new_[69196]_  = A233 & A232;
  assign \new_[69199]_  = ~A267 & A265;
  assign \new_[69200]_  = \new_[69199]_  & \new_[69196]_ ;
  assign \new_[69203]_  = ~A299 & A298;
  assign \new_[69206]_  = A302 & A300;
  assign \new_[69207]_  = \new_[69206]_  & \new_[69203]_ ;
  assign \new_[69208]_  = \new_[69207]_  & \new_[69200]_ ;
  assign \new_[69212]_  = ~A166 & ~A167;
  assign \new_[69213]_  = ~A169 & \new_[69212]_ ;
  assign \new_[69216]_  = ~A200 & A199;
  assign \new_[69219]_  = A203 & A201;
  assign \new_[69220]_  = \new_[69219]_  & \new_[69216]_ ;
  assign \new_[69221]_  = \new_[69220]_  & \new_[69213]_ ;
  assign \new_[69224]_  = A233 & A232;
  assign \new_[69227]_  = A266 & A265;
  assign \new_[69228]_  = \new_[69227]_  & \new_[69224]_ ;
  assign \new_[69231]_  = ~A299 & A298;
  assign \new_[69234]_  = A301 & A300;
  assign \new_[69235]_  = \new_[69234]_  & \new_[69231]_ ;
  assign \new_[69236]_  = \new_[69235]_  & \new_[69228]_ ;
  assign \new_[69240]_  = ~A166 & ~A167;
  assign \new_[69241]_  = ~A169 & \new_[69240]_ ;
  assign \new_[69244]_  = ~A200 & A199;
  assign \new_[69247]_  = A203 & A201;
  assign \new_[69248]_  = \new_[69247]_  & \new_[69244]_ ;
  assign \new_[69249]_  = \new_[69248]_  & \new_[69241]_ ;
  assign \new_[69252]_  = A233 & A232;
  assign \new_[69255]_  = A266 & A265;
  assign \new_[69256]_  = \new_[69255]_  & \new_[69252]_ ;
  assign \new_[69259]_  = ~A299 & A298;
  assign \new_[69262]_  = A302 & A300;
  assign \new_[69263]_  = \new_[69262]_  & \new_[69259]_ ;
  assign \new_[69264]_  = \new_[69263]_  & \new_[69256]_ ;
  assign \new_[69268]_  = ~A166 & ~A167;
  assign \new_[69269]_  = ~A169 & \new_[69268]_ ;
  assign \new_[69272]_  = ~A200 & A199;
  assign \new_[69275]_  = A203 & A201;
  assign \new_[69276]_  = \new_[69275]_  & \new_[69272]_ ;
  assign \new_[69277]_  = \new_[69276]_  & \new_[69269]_ ;
  assign \new_[69280]_  = A233 & A232;
  assign \new_[69283]_  = ~A266 & ~A265;
  assign \new_[69284]_  = \new_[69283]_  & \new_[69280]_ ;
  assign \new_[69287]_  = ~A299 & A298;
  assign \new_[69290]_  = A301 & A300;
  assign \new_[69291]_  = \new_[69290]_  & \new_[69287]_ ;
  assign \new_[69292]_  = \new_[69291]_  & \new_[69284]_ ;
  assign \new_[69296]_  = ~A166 & ~A167;
  assign \new_[69297]_  = ~A169 & \new_[69296]_ ;
  assign \new_[69300]_  = ~A200 & A199;
  assign \new_[69303]_  = A203 & A201;
  assign \new_[69304]_  = \new_[69303]_  & \new_[69300]_ ;
  assign \new_[69305]_  = \new_[69304]_  & \new_[69297]_ ;
  assign \new_[69308]_  = A233 & A232;
  assign \new_[69311]_  = ~A266 & ~A265;
  assign \new_[69312]_  = \new_[69311]_  & \new_[69308]_ ;
  assign \new_[69315]_  = ~A299 & A298;
  assign \new_[69318]_  = A302 & A300;
  assign \new_[69319]_  = \new_[69318]_  & \new_[69315]_ ;
  assign \new_[69320]_  = \new_[69319]_  & \new_[69312]_ ;
  assign \new_[69324]_  = ~A166 & ~A167;
  assign \new_[69325]_  = ~A169 & \new_[69324]_ ;
  assign \new_[69328]_  = ~A200 & A199;
  assign \new_[69331]_  = A203 & A201;
  assign \new_[69332]_  = \new_[69331]_  & \new_[69328]_ ;
  assign \new_[69333]_  = \new_[69332]_  & \new_[69325]_ ;
  assign \new_[69336]_  = ~A235 & ~A233;
  assign \new_[69339]_  = ~A266 & ~A236;
  assign \new_[69340]_  = \new_[69339]_  & \new_[69336]_ ;
  assign \new_[69343]_  = ~A269 & ~A268;
  assign \new_[69346]_  = A299 & ~A298;
  assign \new_[69347]_  = \new_[69346]_  & \new_[69343]_ ;
  assign \new_[69348]_  = \new_[69347]_  & \new_[69340]_ ;
  assign \new_[69352]_  = ~A166 & ~A167;
  assign \new_[69353]_  = ~A169 & \new_[69352]_ ;
  assign \new_[69356]_  = ~A200 & A199;
  assign \new_[69359]_  = A203 & A201;
  assign \new_[69360]_  = \new_[69359]_  & \new_[69356]_ ;
  assign \new_[69361]_  = \new_[69360]_  & \new_[69353]_ ;
  assign \new_[69364]_  = ~A234 & ~A233;
  assign \new_[69367]_  = A266 & A265;
  assign \new_[69368]_  = \new_[69367]_  & \new_[69364]_ ;
  assign \new_[69371]_  = ~A299 & A298;
  assign \new_[69374]_  = A301 & A300;
  assign \new_[69375]_  = \new_[69374]_  & \new_[69371]_ ;
  assign \new_[69376]_  = \new_[69375]_  & \new_[69368]_ ;
  assign \new_[69380]_  = ~A166 & ~A167;
  assign \new_[69381]_  = ~A169 & \new_[69380]_ ;
  assign \new_[69384]_  = ~A200 & A199;
  assign \new_[69387]_  = A203 & A201;
  assign \new_[69388]_  = \new_[69387]_  & \new_[69384]_ ;
  assign \new_[69389]_  = \new_[69388]_  & \new_[69381]_ ;
  assign \new_[69392]_  = ~A234 & ~A233;
  assign \new_[69395]_  = A266 & A265;
  assign \new_[69396]_  = \new_[69395]_  & \new_[69392]_ ;
  assign \new_[69399]_  = ~A299 & A298;
  assign \new_[69402]_  = A302 & A300;
  assign \new_[69403]_  = \new_[69402]_  & \new_[69399]_ ;
  assign \new_[69404]_  = \new_[69403]_  & \new_[69396]_ ;
  assign \new_[69408]_  = ~A166 & ~A167;
  assign \new_[69409]_  = ~A169 & \new_[69408]_ ;
  assign \new_[69412]_  = ~A200 & A199;
  assign \new_[69415]_  = A203 & A201;
  assign \new_[69416]_  = \new_[69415]_  & \new_[69412]_ ;
  assign \new_[69417]_  = \new_[69416]_  & \new_[69409]_ ;
  assign \new_[69420]_  = ~A234 & ~A233;
  assign \new_[69423]_  = ~A267 & ~A266;
  assign \new_[69424]_  = \new_[69423]_  & \new_[69420]_ ;
  assign \new_[69427]_  = ~A299 & A298;
  assign \new_[69430]_  = A301 & A300;
  assign \new_[69431]_  = \new_[69430]_  & \new_[69427]_ ;
  assign \new_[69432]_  = \new_[69431]_  & \new_[69424]_ ;
  assign \new_[69436]_  = ~A166 & ~A167;
  assign \new_[69437]_  = ~A169 & \new_[69436]_ ;
  assign \new_[69440]_  = ~A200 & A199;
  assign \new_[69443]_  = A203 & A201;
  assign \new_[69444]_  = \new_[69443]_  & \new_[69440]_ ;
  assign \new_[69445]_  = \new_[69444]_  & \new_[69437]_ ;
  assign \new_[69448]_  = ~A234 & ~A233;
  assign \new_[69451]_  = ~A267 & ~A266;
  assign \new_[69452]_  = \new_[69451]_  & \new_[69448]_ ;
  assign \new_[69455]_  = ~A299 & A298;
  assign \new_[69458]_  = A302 & A300;
  assign \new_[69459]_  = \new_[69458]_  & \new_[69455]_ ;
  assign \new_[69460]_  = \new_[69459]_  & \new_[69452]_ ;
  assign \new_[69464]_  = ~A166 & ~A167;
  assign \new_[69465]_  = ~A169 & \new_[69464]_ ;
  assign \new_[69468]_  = ~A200 & A199;
  assign \new_[69471]_  = A203 & A201;
  assign \new_[69472]_  = \new_[69471]_  & \new_[69468]_ ;
  assign \new_[69473]_  = \new_[69472]_  & \new_[69465]_ ;
  assign \new_[69476]_  = ~A234 & ~A233;
  assign \new_[69479]_  = ~A266 & ~A265;
  assign \new_[69480]_  = \new_[69479]_  & \new_[69476]_ ;
  assign \new_[69483]_  = ~A299 & A298;
  assign \new_[69486]_  = A301 & A300;
  assign \new_[69487]_  = \new_[69486]_  & \new_[69483]_ ;
  assign \new_[69488]_  = \new_[69487]_  & \new_[69480]_ ;
  assign \new_[69492]_  = ~A166 & ~A167;
  assign \new_[69493]_  = ~A169 & \new_[69492]_ ;
  assign \new_[69496]_  = ~A200 & A199;
  assign \new_[69499]_  = A203 & A201;
  assign \new_[69500]_  = \new_[69499]_  & \new_[69496]_ ;
  assign \new_[69501]_  = \new_[69500]_  & \new_[69493]_ ;
  assign \new_[69504]_  = ~A234 & ~A233;
  assign \new_[69507]_  = ~A266 & ~A265;
  assign \new_[69508]_  = \new_[69507]_  & \new_[69504]_ ;
  assign \new_[69511]_  = ~A299 & A298;
  assign \new_[69514]_  = A302 & A300;
  assign \new_[69515]_  = \new_[69514]_  & \new_[69511]_ ;
  assign \new_[69516]_  = \new_[69515]_  & \new_[69508]_ ;
  assign \new_[69520]_  = ~A166 & ~A167;
  assign \new_[69521]_  = ~A169 & \new_[69520]_ ;
  assign \new_[69524]_  = ~A200 & A199;
  assign \new_[69527]_  = A203 & A201;
  assign \new_[69528]_  = \new_[69527]_  & \new_[69524]_ ;
  assign \new_[69529]_  = \new_[69528]_  & \new_[69521]_ ;
  assign \new_[69532]_  = ~A233 & A232;
  assign \new_[69535]_  = A235 & A234;
  assign \new_[69536]_  = \new_[69535]_  & \new_[69532]_ ;
  assign \new_[69539]_  = ~A266 & A265;
  assign \new_[69542]_  = A268 & A267;
  assign \new_[69543]_  = \new_[69542]_  & \new_[69539]_ ;
  assign \new_[69544]_  = \new_[69543]_  & \new_[69536]_ ;
  assign \new_[69548]_  = ~A166 & ~A167;
  assign \new_[69549]_  = ~A169 & \new_[69548]_ ;
  assign \new_[69552]_  = ~A200 & A199;
  assign \new_[69555]_  = A203 & A201;
  assign \new_[69556]_  = \new_[69555]_  & \new_[69552]_ ;
  assign \new_[69557]_  = \new_[69556]_  & \new_[69549]_ ;
  assign \new_[69560]_  = ~A233 & A232;
  assign \new_[69563]_  = A235 & A234;
  assign \new_[69564]_  = \new_[69563]_  & \new_[69560]_ ;
  assign \new_[69567]_  = ~A266 & A265;
  assign \new_[69570]_  = A269 & A267;
  assign \new_[69571]_  = \new_[69570]_  & \new_[69567]_ ;
  assign \new_[69572]_  = \new_[69571]_  & \new_[69564]_ ;
  assign \new_[69576]_  = ~A166 & ~A167;
  assign \new_[69577]_  = ~A169 & \new_[69576]_ ;
  assign \new_[69580]_  = ~A200 & A199;
  assign \new_[69583]_  = A203 & A201;
  assign \new_[69584]_  = \new_[69583]_  & \new_[69580]_ ;
  assign \new_[69585]_  = \new_[69584]_  & \new_[69577]_ ;
  assign \new_[69588]_  = ~A233 & A232;
  assign \new_[69591]_  = A236 & A234;
  assign \new_[69592]_  = \new_[69591]_  & \new_[69588]_ ;
  assign \new_[69595]_  = ~A266 & A265;
  assign \new_[69598]_  = A268 & A267;
  assign \new_[69599]_  = \new_[69598]_  & \new_[69595]_ ;
  assign \new_[69600]_  = \new_[69599]_  & \new_[69592]_ ;
  assign \new_[69604]_  = ~A166 & ~A167;
  assign \new_[69605]_  = ~A169 & \new_[69604]_ ;
  assign \new_[69608]_  = ~A200 & A199;
  assign \new_[69611]_  = A203 & A201;
  assign \new_[69612]_  = \new_[69611]_  & \new_[69608]_ ;
  assign \new_[69613]_  = \new_[69612]_  & \new_[69605]_ ;
  assign \new_[69616]_  = ~A233 & A232;
  assign \new_[69619]_  = A236 & A234;
  assign \new_[69620]_  = \new_[69619]_  & \new_[69616]_ ;
  assign \new_[69623]_  = ~A266 & A265;
  assign \new_[69626]_  = A269 & A267;
  assign \new_[69627]_  = \new_[69626]_  & \new_[69623]_ ;
  assign \new_[69628]_  = \new_[69627]_  & \new_[69620]_ ;
  assign \new_[69632]_  = ~A166 & ~A167;
  assign \new_[69633]_  = ~A169 & \new_[69632]_ ;
  assign \new_[69636]_  = ~A200 & A199;
  assign \new_[69639]_  = A203 & A201;
  assign \new_[69640]_  = \new_[69639]_  & \new_[69636]_ ;
  assign \new_[69641]_  = \new_[69640]_  & \new_[69633]_ ;
  assign \new_[69644]_  = ~A233 & ~A232;
  assign \new_[69647]_  = A266 & A265;
  assign \new_[69648]_  = \new_[69647]_  & \new_[69644]_ ;
  assign \new_[69651]_  = ~A299 & A298;
  assign \new_[69654]_  = A301 & A300;
  assign \new_[69655]_  = \new_[69654]_  & \new_[69651]_ ;
  assign \new_[69656]_  = \new_[69655]_  & \new_[69648]_ ;
  assign \new_[69660]_  = ~A166 & ~A167;
  assign \new_[69661]_  = ~A169 & \new_[69660]_ ;
  assign \new_[69664]_  = ~A200 & A199;
  assign \new_[69667]_  = A203 & A201;
  assign \new_[69668]_  = \new_[69667]_  & \new_[69664]_ ;
  assign \new_[69669]_  = \new_[69668]_  & \new_[69661]_ ;
  assign \new_[69672]_  = ~A233 & ~A232;
  assign \new_[69675]_  = A266 & A265;
  assign \new_[69676]_  = \new_[69675]_  & \new_[69672]_ ;
  assign \new_[69679]_  = ~A299 & A298;
  assign \new_[69682]_  = A302 & A300;
  assign \new_[69683]_  = \new_[69682]_  & \new_[69679]_ ;
  assign \new_[69684]_  = \new_[69683]_  & \new_[69676]_ ;
  assign \new_[69688]_  = ~A166 & ~A167;
  assign \new_[69689]_  = ~A169 & \new_[69688]_ ;
  assign \new_[69692]_  = ~A200 & A199;
  assign \new_[69695]_  = A203 & A201;
  assign \new_[69696]_  = \new_[69695]_  & \new_[69692]_ ;
  assign \new_[69697]_  = \new_[69696]_  & \new_[69689]_ ;
  assign \new_[69700]_  = ~A233 & ~A232;
  assign \new_[69703]_  = ~A267 & ~A266;
  assign \new_[69704]_  = \new_[69703]_  & \new_[69700]_ ;
  assign \new_[69707]_  = ~A299 & A298;
  assign \new_[69710]_  = A301 & A300;
  assign \new_[69711]_  = \new_[69710]_  & \new_[69707]_ ;
  assign \new_[69712]_  = \new_[69711]_  & \new_[69704]_ ;
  assign \new_[69716]_  = ~A166 & ~A167;
  assign \new_[69717]_  = ~A169 & \new_[69716]_ ;
  assign \new_[69720]_  = ~A200 & A199;
  assign \new_[69723]_  = A203 & A201;
  assign \new_[69724]_  = \new_[69723]_  & \new_[69720]_ ;
  assign \new_[69725]_  = \new_[69724]_  & \new_[69717]_ ;
  assign \new_[69728]_  = ~A233 & ~A232;
  assign \new_[69731]_  = ~A267 & ~A266;
  assign \new_[69732]_  = \new_[69731]_  & \new_[69728]_ ;
  assign \new_[69735]_  = ~A299 & A298;
  assign \new_[69738]_  = A302 & A300;
  assign \new_[69739]_  = \new_[69738]_  & \new_[69735]_ ;
  assign \new_[69740]_  = \new_[69739]_  & \new_[69732]_ ;
  assign \new_[69744]_  = ~A166 & ~A167;
  assign \new_[69745]_  = ~A169 & \new_[69744]_ ;
  assign \new_[69748]_  = ~A200 & A199;
  assign \new_[69751]_  = A203 & A201;
  assign \new_[69752]_  = \new_[69751]_  & \new_[69748]_ ;
  assign \new_[69753]_  = \new_[69752]_  & \new_[69745]_ ;
  assign \new_[69756]_  = ~A233 & ~A232;
  assign \new_[69759]_  = ~A266 & ~A265;
  assign \new_[69760]_  = \new_[69759]_  & \new_[69756]_ ;
  assign \new_[69763]_  = ~A299 & A298;
  assign \new_[69766]_  = A301 & A300;
  assign \new_[69767]_  = \new_[69766]_  & \new_[69763]_ ;
  assign \new_[69768]_  = \new_[69767]_  & \new_[69760]_ ;
  assign \new_[69772]_  = ~A166 & ~A167;
  assign \new_[69773]_  = ~A169 & \new_[69772]_ ;
  assign \new_[69776]_  = ~A200 & A199;
  assign \new_[69779]_  = A203 & A201;
  assign \new_[69780]_  = \new_[69779]_  & \new_[69776]_ ;
  assign \new_[69781]_  = \new_[69780]_  & \new_[69773]_ ;
  assign \new_[69784]_  = ~A233 & ~A232;
  assign \new_[69787]_  = ~A266 & ~A265;
  assign \new_[69788]_  = \new_[69787]_  & \new_[69784]_ ;
  assign \new_[69791]_  = ~A299 & A298;
  assign \new_[69794]_  = A302 & A300;
  assign \new_[69795]_  = \new_[69794]_  & \new_[69791]_ ;
  assign \new_[69796]_  = \new_[69795]_  & \new_[69788]_ ;
  assign \new_[69800]_  = A167 & ~A168;
  assign \new_[69801]_  = ~A169 & \new_[69800]_ ;
  assign \new_[69804]_  = ~A199 & A166;
  assign \new_[69807]_  = A232 & A200;
  assign \new_[69808]_  = \new_[69807]_  & \new_[69804]_ ;
  assign \new_[69809]_  = \new_[69808]_  & \new_[69801]_ ;
  assign \new_[69812]_  = A265 & A233;
  assign \new_[69815]_  = ~A269 & ~A268;
  assign \new_[69816]_  = \new_[69815]_  & \new_[69812]_ ;
  assign \new_[69819]_  = ~A299 & A298;
  assign \new_[69822]_  = A301 & A300;
  assign \new_[69823]_  = \new_[69822]_  & \new_[69819]_ ;
  assign \new_[69824]_  = \new_[69823]_  & \new_[69816]_ ;
  assign \new_[69828]_  = A167 & ~A168;
  assign \new_[69829]_  = ~A169 & \new_[69828]_ ;
  assign \new_[69832]_  = ~A199 & A166;
  assign \new_[69835]_  = A232 & A200;
  assign \new_[69836]_  = \new_[69835]_  & \new_[69832]_ ;
  assign \new_[69837]_  = \new_[69836]_  & \new_[69829]_ ;
  assign \new_[69840]_  = A265 & A233;
  assign \new_[69843]_  = ~A269 & ~A268;
  assign \new_[69844]_  = \new_[69843]_  & \new_[69840]_ ;
  assign \new_[69847]_  = ~A299 & A298;
  assign \new_[69850]_  = A302 & A300;
  assign \new_[69851]_  = \new_[69850]_  & \new_[69847]_ ;
  assign \new_[69852]_  = \new_[69851]_  & \new_[69844]_ ;
  assign \new_[69856]_  = A167 & ~A168;
  assign \new_[69857]_  = ~A169 & \new_[69856]_ ;
  assign \new_[69860]_  = ~A199 & A166;
  assign \new_[69863]_  = ~A233 & A200;
  assign \new_[69864]_  = \new_[69863]_  & \new_[69860]_ ;
  assign \new_[69865]_  = \new_[69864]_  & \new_[69857]_ ;
  assign \new_[69868]_  = ~A236 & ~A235;
  assign \new_[69871]_  = A266 & A265;
  assign \new_[69872]_  = \new_[69871]_  & \new_[69868]_ ;
  assign \new_[69875]_  = ~A299 & A298;
  assign \new_[69878]_  = A301 & A300;
  assign \new_[69879]_  = \new_[69878]_  & \new_[69875]_ ;
  assign \new_[69880]_  = \new_[69879]_  & \new_[69872]_ ;
  assign \new_[69884]_  = A167 & ~A168;
  assign \new_[69885]_  = ~A169 & \new_[69884]_ ;
  assign \new_[69888]_  = ~A199 & A166;
  assign \new_[69891]_  = ~A233 & A200;
  assign \new_[69892]_  = \new_[69891]_  & \new_[69888]_ ;
  assign \new_[69893]_  = \new_[69892]_  & \new_[69885]_ ;
  assign \new_[69896]_  = ~A236 & ~A235;
  assign \new_[69899]_  = A266 & A265;
  assign \new_[69900]_  = \new_[69899]_  & \new_[69896]_ ;
  assign \new_[69903]_  = ~A299 & A298;
  assign \new_[69906]_  = A302 & A300;
  assign \new_[69907]_  = \new_[69906]_  & \new_[69903]_ ;
  assign \new_[69908]_  = \new_[69907]_  & \new_[69900]_ ;
  assign \new_[69912]_  = A167 & ~A168;
  assign \new_[69913]_  = ~A169 & \new_[69912]_ ;
  assign \new_[69916]_  = ~A199 & A166;
  assign \new_[69919]_  = ~A233 & A200;
  assign \new_[69920]_  = \new_[69919]_  & \new_[69916]_ ;
  assign \new_[69921]_  = \new_[69920]_  & \new_[69913]_ ;
  assign \new_[69924]_  = ~A236 & ~A235;
  assign \new_[69927]_  = ~A267 & ~A266;
  assign \new_[69928]_  = \new_[69927]_  & \new_[69924]_ ;
  assign \new_[69931]_  = ~A299 & A298;
  assign \new_[69934]_  = A301 & A300;
  assign \new_[69935]_  = \new_[69934]_  & \new_[69931]_ ;
  assign \new_[69936]_  = \new_[69935]_  & \new_[69928]_ ;
  assign \new_[69940]_  = A167 & ~A168;
  assign \new_[69941]_  = ~A169 & \new_[69940]_ ;
  assign \new_[69944]_  = ~A199 & A166;
  assign \new_[69947]_  = ~A233 & A200;
  assign \new_[69948]_  = \new_[69947]_  & \new_[69944]_ ;
  assign \new_[69949]_  = \new_[69948]_  & \new_[69941]_ ;
  assign \new_[69952]_  = ~A236 & ~A235;
  assign \new_[69955]_  = ~A267 & ~A266;
  assign \new_[69956]_  = \new_[69955]_  & \new_[69952]_ ;
  assign \new_[69959]_  = ~A299 & A298;
  assign \new_[69962]_  = A302 & A300;
  assign \new_[69963]_  = \new_[69962]_  & \new_[69959]_ ;
  assign \new_[69964]_  = \new_[69963]_  & \new_[69956]_ ;
  assign \new_[69968]_  = A167 & ~A168;
  assign \new_[69969]_  = ~A169 & \new_[69968]_ ;
  assign \new_[69972]_  = ~A199 & A166;
  assign \new_[69975]_  = ~A233 & A200;
  assign \new_[69976]_  = \new_[69975]_  & \new_[69972]_ ;
  assign \new_[69977]_  = \new_[69976]_  & \new_[69969]_ ;
  assign \new_[69980]_  = ~A236 & ~A235;
  assign \new_[69983]_  = ~A266 & ~A265;
  assign \new_[69984]_  = \new_[69983]_  & \new_[69980]_ ;
  assign \new_[69987]_  = ~A299 & A298;
  assign \new_[69990]_  = A301 & A300;
  assign \new_[69991]_  = \new_[69990]_  & \new_[69987]_ ;
  assign \new_[69992]_  = \new_[69991]_  & \new_[69984]_ ;
  assign \new_[69996]_  = A167 & ~A168;
  assign \new_[69997]_  = ~A169 & \new_[69996]_ ;
  assign \new_[70000]_  = ~A199 & A166;
  assign \new_[70003]_  = ~A233 & A200;
  assign \new_[70004]_  = \new_[70003]_  & \new_[70000]_ ;
  assign \new_[70005]_  = \new_[70004]_  & \new_[69997]_ ;
  assign \new_[70008]_  = ~A236 & ~A235;
  assign \new_[70011]_  = ~A266 & ~A265;
  assign \new_[70012]_  = \new_[70011]_  & \new_[70008]_ ;
  assign \new_[70015]_  = ~A299 & A298;
  assign \new_[70018]_  = A302 & A300;
  assign \new_[70019]_  = \new_[70018]_  & \new_[70015]_ ;
  assign \new_[70020]_  = \new_[70019]_  & \new_[70012]_ ;
  assign \new_[70024]_  = A167 & ~A168;
  assign \new_[70025]_  = ~A169 & \new_[70024]_ ;
  assign \new_[70028]_  = ~A199 & A166;
  assign \new_[70031]_  = ~A233 & A200;
  assign \new_[70032]_  = \new_[70031]_  & \new_[70028]_ ;
  assign \new_[70033]_  = \new_[70032]_  & \new_[70025]_ ;
  assign \new_[70036]_  = ~A266 & ~A234;
  assign \new_[70039]_  = ~A269 & ~A268;
  assign \new_[70040]_  = \new_[70039]_  & \new_[70036]_ ;
  assign \new_[70043]_  = ~A299 & A298;
  assign \new_[70046]_  = A301 & A300;
  assign \new_[70047]_  = \new_[70046]_  & \new_[70043]_ ;
  assign \new_[70048]_  = \new_[70047]_  & \new_[70040]_ ;
  assign \new_[70052]_  = A167 & ~A168;
  assign \new_[70053]_  = ~A169 & \new_[70052]_ ;
  assign \new_[70056]_  = ~A199 & A166;
  assign \new_[70059]_  = ~A233 & A200;
  assign \new_[70060]_  = \new_[70059]_  & \new_[70056]_ ;
  assign \new_[70061]_  = \new_[70060]_  & \new_[70053]_ ;
  assign \new_[70064]_  = ~A266 & ~A234;
  assign \new_[70067]_  = ~A269 & ~A268;
  assign \new_[70068]_  = \new_[70067]_  & \new_[70064]_ ;
  assign \new_[70071]_  = ~A299 & A298;
  assign \new_[70074]_  = A302 & A300;
  assign \new_[70075]_  = \new_[70074]_  & \new_[70071]_ ;
  assign \new_[70076]_  = \new_[70075]_  & \new_[70068]_ ;
  assign \new_[70080]_  = A167 & ~A168;
  assign \new_[70081]_  = ~A169 & \new_[70080]_ ;
  assign \new_[70084]_  = ~A199 & A166;
  assign \new_[70087]_  = ~A232 & A200;
  assign \new_[70088]_  = \new_[70087]_  & \new_[70084]_ ;
  assign \new_[70089]_  = \new_[70088]_  & \new_[70081]_ ;
  assign \new_[70092]_  = ~A266 & ~A233;
  assign \new_[70095]_  = ~A269 & ~A268;
  assign \new_[70096]_  = \new_[70095]_  & \new_[70092]_ ;
  assign \new_[70099]_  = ~A299 & A298;
  assign \new_[70102]_  = A301 & A300;
  assign \new_[70103]_  = \new_[70102]_  & \new_[70099]_ ;
  assign \new_[70104]_  = \new_[70103]_  & \new_[70096]_ ;
  assign \new_[70108]_  = A167 & ~A168;
  assign \new_[70109]_  = ~A169 & \new_[70108]_ ;
  assign \new_[70112]_  = ~A199 & A166;
  assign \new_[70115]_  = ~A232 & A200;
  assign \new_[70116]_  = \new_[70115]_  & \new_[70112]_ ;
  assign \new_[70117]_  = \new_[70116]_  & \new_[70109]_ ;
  assign \new_[70120]_  = ~A266 & ~A233;
  assign \new_[70123]_  = ~A269 & ~A268;
  assign \new_[70124]_  = \new_[70123]_  & \new_[70120]_ ;
  assign \new_[70127]_  = ~A299 & A298;
  assign \new_[70130]_  = A302 & A300;
  assign \new_[70131]_  = \new_[70130]_  & \new_[70127]_ ;
  assign \new_[70132]_  = \new_[70131]_  & \new_[70124]_ ;
  assign \new_[70136]_  = A167 & ~A168;
  assign \new_[70137]_  = ~A169 & \new_[70136]_ ;
  assign \new_[70140]_  = A199 & A166;
  assign \new_[70143]_  = A201 & ~A200;
  assign \new_[70144]_  = \new_[70143]_  & \new_[70140]_ ;
  assign \new_[70145]_  = \new_[70144]_  & \new_[70137]_ ;
  assign \new_[70148]_  = A232 & A202;
  assign \new_[70151]_  = A265 & A233;
  assign \new_[70152]_  = \new_[70151]_  & \new_[70148]_ ;
  assign \new_[70155]_  = ~A269 & ~A268;
  assign \new_[70158]_  = A299 & ~A298;
  assign \new_[70159]_  = \new_[70158]_  & \new_[70155]_ ;
  assign \new_[70160]_  = \new_[70159]_  & \new_[70152]_ ;
  assign \new_[70164]_  = A167 & ~A168;
  assign \new_[70165]_  = ~A169 & \new_[70164]_ ;
  assign \new_[70168]_  = A199 & A166;
  assign \new_[70171]_  = A201 & ~A200;
  assign \new_[70172]_  = \new_[70171]_  & \new_[70168]_ ;
  assign \new_[70173]_  = \new_[70172]_  & \new_[70165]_ ;
  assign \new_[70176]_  = ~A233 & A202;
  assign \new_[70179]_  = ~A236 & ~A235;
  assign \new_[70180]_  = \new_[70179]_  & \new_[70176]_ ;
  assign \new_[70183]_  = A266 & A265;
  assign \new_[70186]_  = A299 & ~A298;
  assign \new_[70187]_  = \new_[70186]_  & \new_[70183]_ ;
  assign \new_[70188]_  = \new_[70187]_  & \new_[70180]_ ;
  assign \new_[70192]_  = A167 & ~A168;
  assign \new_[70193]_  = ~A169 & \new_[70192]_ ;
  assign \new_[70196]_  = A199 & A166;
  assign \new_[70199]_  = A201 & ~A200;
  assign \new_[70200]_  = \new_[70199]_  & \new_[70196]_ ;
  assign \new_[70201]_  = \new_[70200]_  & \new_[70193]_ ;
  assign \new_[70204]_  = ~A233 & A202;
  assign \new_[70207]_  = ~A236 & ~A235;
  assign \new_[70208]_  = \new_[70207]_  & \new_[70204]_ ;
  assign \new_[70211]_  = ~A267 & ~A266;
  assign \new_[70214]_  = A299 & ~A298;
  assign \new_[70215]_  = \new_[70214]_  & \new_[70211]_ ;
  assign \new_[70216]_  = \new_[70215]_  & \new_[70208]_ ;
  assign \new_[70220]_  = A167 & ~A168;
  assign \new_[70221]_  = ~A169 & \new_[70220]_ ;
  assign \new_[70224]_  = A199 & A166;
  assign \new_[70227]_  = A201 & ~A200;
  assign \new_[70228]_  = \new_[70227]_  & \new_[70224]_ ;
  assign \new_[70229]_  = \new_[70228]_  & \new_[70221]_ ;
  assign \new_[70232]_  = ~A233 & A202;
  assign \new_[70235]_  = ~A236 & ~A235;
  assign \new_[70236]_  = \new_[70235]_  & \new_[70232]_ ;
  assign \new_[70239]_  = ~A266 & ~A265;
  assign \new_[70242]_  = A299 & ~A298;
  assign \new_[70243]_  = \new_[70242]_  & \new_[70239]_ ;
  assign \new_[70244]_  = \new_[70243]_  & \new_[70236]_ ;
  assign \new_[70248]_  = A167 & ~A168;
  assign \new_[70249]_  = ~A169 & \new_[70248]_ ;
  assign \new_[70252]_  = A199 & A166;
  assign \new_[70255]_  = A201 & ~A200;
  assign \new_[70256]_  = \new_[70255]_  & \new_[70252]_ ;
  assign \new_[70257]_  = \new_[70256]_  & \new_[70249]_ ;
  assign \new_[70260]_  = ~A233 & A202;
  assign \new_[70263]_  = ~A266 & ~A234;
  assign \new_[70264]_  = \new_[70263]_  & \new_[70260]_ ;
  assign \new_[70267]_  = ~A269 & ~A268;
  assign \new_[70270]_  = A299 & ~A298;
  assign \new_[70271]_  = \new_[70270]_  & \new_[70267]_ ;
  assign \new_[70272]_  = \new_[70271]_  & \new_[70264]_ ;
  assign \new_[70276]_  = A167 & ~A168;
  assign \new_[70277]_  = ~A169 & \new_[70276]_ ;
  assign \new_[70280]_  = A199 & A166;
  assign \new_[70283]_  = A201 & ~A200;
  assign \new_[70284]_  = \new_[70283]_  & \new_[70280]_ ;
  assign \new_[70285]_  = \new_[70284]_  & \new_[70277]_ ;
  assign \new_[70288]_  = A232 & A202;
  assign \new_[70291]_  = A234 & ~A233;
  assign \new_[70292]_  = \new_[70291]_  & \new_[70288]_ ;
  assign \new_[70295]_  = A298 & A235;
  assign \new_[70298]_  = ~A302 & ~A301;
  assign \new_[70299]_  = \new_[70298]_  & \new_[70295]_ ;
  assign \new_[70300]_  = \new_[70299]_  & \new_[70292]_ ;
  assign \new_[70304]_  = A167 & ~A168;
  assign \new_[70305]_  = ~A169 & \new_[70304]_ ;
  assign \new_[70308]_  = A199 & A166;
  assign \new_[70311]_  = A201 & ~A200;
  assign \new_[70312]_  = \new_[70311]_  & \new_[70308]_ ;
  assign \new_[70313]_  = \new_[70312]_  & \new_[70305]_ ;
  assign \new_[70316]_  = A232 & A202;
  assign \new_[70319]_  = A234 & ~A233;
  assign \new_[70320]_  = \new_[70319]_  & \new_[70316]_ ;
  assign \new_[70323]_  = A298 & A236;
  assign \new_[70326]_  = ~A302 & ~A301;
  assign \new_[70327]_  = \new_[70326]_  & \new_[70323]_ ;
  assign \new_[70328]_  = \new_[70327]_  & \new_[70320]_ ;
  assign \new_[70332]_  = A167 & ~A168;
  assign \new_[70333]_  = ~A169 & \new_[70332]_ ;
  assign \new_[70336]_  = A199 & A166;
  assign \new_[70339]_  = A201 & ~A200;
  assign \new_[70340]_  = \new_[70339]_  & \new_[70336]_ ;
  assign \new_[70341]_  = \new_[70340]_  & \new_[70333]_ ;
  assign \new_[70344]_  = ~A232 & A202;
  assign \new_[70347]_  = ~A266 & ~A233;
  assign \new_[70348]_  = \new_[70347]_  & \new_[70344]_ ;
  assign \new_[70351]_  = ~A269 & ~A268;
  assign \new_[70354]_  = A299 & ~A298;
  assign \new_[70355]_  = \new_[70354]_  & \new_[70351]_ ;
  assign \new_[70356]_  = \new_[70355]_  & \new_[70348]_ ;
  assign \new_[70360]_  = A167 & ~A168;
  assign \new_[70361]_  = ~A169 & \new_[70360]_ ;
  assign \new_[70364]_  = A199 & A166;
  assign \new_[70367]_  = A201 & ~A200;
  assign \new_[70368]_  = \new_[70367]_  & \new_[70364]_ ;
  assign \new_[70369]_  = \new_[70368]_  & \new_[70361]_ ;
  assign \new_[70372]_  = A232 & A203;
  assign \new_[70375]_  = A265 & A233;
  assign \new_[70376]_  = \new_[70375]_  & \new_[70372]_ ;
  assign \new_[70379]_  = ~A269 & ~A268;
  assign \new_[70382]_  = A299 & ~A298;
  assign \new_[70383]_  = \new_[70382]_  & \new_[70379]_ ;
  assign \new_[70384]_  = \new_[70383]_  & \new_[70376]_ ;
  assign \new_[70388]_  = A167 & ~A168;
  assign \new_[70389]_  = ~A169 & \new_[70388]_ ;
  assign \new_[70392]_  = A199 & A166;
  assign \new_[70395]_  = A201 & ~A200;
  assign \new_[70396]_  = \new_[70395]_  & \new_[70392]_ ;
  assign \new_[70397]_  = \new_[70396]_  & \new_[70389]_ ;
  assign \new_[70400]_  = ~A233 & A203;
  assign \new_[70403]_  = ~A236 & ~A235;
  assign \new_[70404]_  = \new_[70403]_  & \new_[70400]_ ;
  assign \new_[70407]_  = A266 & A265;
  assign \new_[70410]_  = A299 & ~A298;
  assign \new_[70411]_  = \new_[70410]_  & \new_[70407]_ ;
  assign \new_[70412]_  = \new_[70411]_  & \new_[70404]_ ;
  assign \new_[70416]_  = A167 & ~A168;
  assign \new_[70417]_  = ~A169 & \new_[70416]_ ;
  assign \new_[70420]_  = A199 & A166;
  assign \new_[70423]_  = A201 & ~A200;
  assign \new_[70424]_  = \new_[70423]_  & \new_[70420]_ ;
  assign \new_[70425]_  = \new_[70424]_  & \new_[70417]_ ;
  assign \new_[70428]_  = ~A233 & A203;
  assign \new_[70431]_  = ~A236 & ~A235;
  assign \new_[70432]_  = \new_[70431]_  & \new_[70428]_ ;
  assign \new_[70435]_  = ~A267 & ~A266;
  assign \new_[70438]_  = A299 & ~A298;
  assign \new_[70439]_  = \new_[70438]_  & \new_[70435]_ ;
  assign \new_[70440]_  = \new_[70439]_  & \new_[70432]_ ;
  assign \new_[70444]_  = A167 & ~A168;
  assign \new_[70445]_  = ~A169 & \new_[70444]_ ;
  assign \new_[70448]_  = A199 & A166;
  assign \new_[70451]_  = A201 & ~A200;
  assign \new_[70452]_  = \new_[70451]_  & \new_[70448]_ ;
  assign \new_[70453]_  = \new_[70452]_  & \new_[70445]_ ;
  assign \new_[70456]_  = ~A233 & A203;
  assign \new_[70459]_  = ~A236 & ~A235;
  assign \new_[70460]_  = \new_[70459]_  & \new_[70456]_ ;
  assign \new_[70463]_  = ~A266 & ~A265;
  assign \new_[70466]_  = A299 & ~A298;
  assign \new_[70467]_  = \new_[70466]_  & \new_[70463]_ ;
  assign \new_[70468]_  = \new_[70467]_  & \new_[70460]_ ;
  assign \new_[70472]_  = A167 & ~A168;
  assign \new_[70473]_  = ~A169 & \new_[70472]_ ;
  assign \new_[70476]_  = A199 & A166;
  assign \new_[70479]_  = A201 & ~A200;
  assign \new_[70480]_  = \new_[70479]_  & \new_[70476]_ ;
  assign \new_[70481]_  = \new_[70480]_  & \new_[70473]_ ;
  assign \new_[70484]_  = ~A233 & A203;
  assign \new_[70487]_  = ~A266 & ~A234;
  assign \new_[70488]_  = \new_[70487]_  & \new_[70484]_ ;
  assign \new_[70491]_  = ~A269 & ~A268;
  assign \new_[70494]_  = A299 & ~A298;
  assign \new_[70495]_  = \new_[70494]_  & \new_[70491]_ ;
  assign \new_[70496]_  = \new_[70495]_  & \new_[70488]_ ;
  assign \new_[70500]_  = A167 & ~A168;
  assign \new_[70501]_  = ~A169 & \new_[70500]_ ;
  assign \new_[70504]_  = A199 & A166;
  assign \new_[70507]_  = A201 & ~A200;
  assign \new_[70508]_  = \new_[70507]_  & \new_[70504]_ ;
  assign \new_[70509]_  = \new_[70508]_  & \new_[70501]_ ;
  assign \new_[70512]_  = A232 & A203;
  assign \new_[70515]_  = A234 & ~A233;
  assign \new_[70516]_  = \new_[70515]_  & \new_[70512]_ ;
  assign \new_[70519]_  = A298 & A235;
  assign \new_[70522]_  = ~A302 & ~A301;
  assign \new_[70523]_  = \new_[70522]_  & \new_[70519]_ ;
  assign \new_[70524]_  = \new_[70523]_  & \new_[70516]_ ;
  assign \new_[70528]_  = A167 & ~A168;
  assign \new_[70529]_  = ~A169 & \new_[70528]_ ;
  assign \new_[70532]_  = A199 & A166;
  assign \new_[70535]_  = A201 & ~A200;
  assign \new_[70536]_  = \new_[70535]_  & \new_[70532]_ ;
  assign \new_[70537]_  = \new_[70536]_  & \new_[70529]_ ;
  assign \new_[70540]_  = A232 & A203;
  assign \new_[70543]_  = A234 & ~A233;
  assign \new_[70544]_  = \new_[70543]_  & \new_[70540]_ ;
  assign \new_[70547]_  = A298 & A236;
  assign \new_[70550]_  = ~A302 & ~A301;
  assign \new_[70551]_  = \new_[70550]_  & \new_[70547]_ ;
  assign \new_[70552]_  = \new_[70551]_  & \new_[70544]_ ;
  assign \new_[70556]_  = A167 & ~A168;
  assign \new_[70557]_  = ~A169 & \new_[70556]_ ;
  assign \new_[70560]_  = A199 & A166;
  assign \new_[70563]_  = A201 & ~A200;
  assign \new_[70564]_  = \new_[70563]_  & \new_[70560]_ ;
  assign \new_[70565]_  = \new_[70564]_  & \new_[70557]_ ;
  assign \new_[70568]_  = ~A232 & A203;
  assign \new_[70571]_  = ~A266 & ~A233;
  assign \new_[70572]_  = \new_[70571]_  & \new_[70568]_ ;
  assign \new_[70575]_  = ~A269 & ~A268;
  assign \new_[70578]_  = A299 & ~A298;
  assign \new_[70579]_  = \new_[70578]_  & \new_[70575]_ ;
  assign \new_[70580]_  = \new_[70579]_  & \new_[70572]_ ;
  assign \new_[70584]_  = A167 & ~A169;
  assign \new_[70585]_  = A170 & \new_[70584]_ ;
  assign \new_[70588]_  = A199 & ~A166;
  assign \new_[70591]_  = A232 & A200;
  assign \new_[70592]_  = \new_[70591]_  & \new_[70588]_ ;
  assign \new_[70593]_  = \new_[70592]_  & \new_[70585]_ ;
  assign \new_[70596]_  = A265 & A233;
  assign \new_[70599]_  = ~A269 & ~A268;
  assign \new_[70600]_  = \new_[70599]_  & \new_[70596]_ ;
  assign \new_[70603]_  = ~A299 & A298;
  assign \new_[70606]_  = A301 & A300;
  assign \new_[70607]_  = \new_[70606]_  & \new_[70603]_ ;
  assign \new_[70608]_  = \new_[70607]_  & \new_[70600]_ ;
  assign \new_[70612]_  = A167 & ~A169;
  assign \new_[70613]_  = A170 & \new_[70612]_ ;
  assign \new_[70616]_  = A199 & ~A166;
  assign \new_[70619]_  = A232 & A200;
  assign \new_[70620]_  = \new_[70619]_  & \new_[70616]_ ;
  assign \new_[70621]_  = \new_[70620]_  & \new_[70613]_ ;
  assign \new_[70624]_  = A265 & A233;
  assign \new_[70627]_  = ~A269 & ~A268;
  assign \new_[70628]_  = \new_[70627]_  & \new_[70624]_ ;
  assign \new_[70631]_  = ~A299 & A298;
  assign \new_[70634]_  = A302 & A300;
  assign \new_[70635]_  = \new_[70634]_  & \new_[70631]_ ;
  assign \new_[70636]_  = \new_[70635]_  & \new_[70628]_ ;
  assign \new_[70640]_  = A167 & ~A169;
  assign \new_[70641]_  = A170 & \new_[70640]_ ;
  assign \new_[70644]_  = A199 & ~A166;
  assign \new_[70647]_  = ~A233 & A200;
  assign \new_[70648]_  = \new_[70647]_  & \new_[70644]_ ;
  assign \new_[70649]_  = \new_[70648]_  & \new_[70641]_ ;
  assign \new_[70652]_  = ~A236 & ~A235;
  assign \new_[70655]_  = A266 & A265;
  assign \new_[70656]_  = \new_[70655]_  & \new_[70652]_ ;
  assign \new_[70659]_  = ~A299 & A298;
  assign \new_[70662]_  = A301 & A300;
  assign \new_[70663]_  = \new_[70662]_  & \new_[70659]_ ;
  assign \new_[70664]_  = \new_[70663]_  & \new_[70656]_ ;
  assign \new_[70668]_  = A167 & ~A169;
  assign \new_[70669]_  = A170 & \new_[70668]_ ;
  assign \new_[70672]_  = A199 & ~A166;
  assign \new_[70675]_  = ~A233 & A200;
  assign \new_[70676]_  = \new_[70675]_  & \new_[70672]_ ;
  assign \new_[70677]_  = \new_[70676]_  & \new_[70669]_ ;
  assign \new_[70680]_  = ~A236 & ~A235;
  assign \new_[70683]_  = A266 & A265;
  assign \new_[70684]_  = \new_[70683]_  & \new_[70680]_ ;
  assign \new_[70687]_  = ~A299 & A298;
  assign \new_[70690]_  = A302 & A300;
  assign \new_[70691]_  = \new_[70690]_  & \new_[70687]_ ;
  assign \new_[70692]_  = \new_[70691]_  & \new_[70684]_ ;
  assign \new_[70696]_  = A167 & ~A169;
  assign \new_[70697]_  = A170 & \new_[70696]_ ;
  assign \new_[70700]_  = A199 & ~A166;
  assign \new_[70703]_  = ~A233 & A200;
  assign \new_[70704]_  = \new_[70703]_  & \new_[70700]_ ;
  assign \new_[70705]_  = \new_[70704]_  & \new_[70697]_ ;
  assign \new_[70708]_  = ~A236 & ~A235;
  assign \new_[70711]_  = ~A267 & ~A266;
  assign \new_[70712]_  = \new_[70711]_  & \new_[70708]_ ;
  assign \new_[70715]_  = ~A299 & A298;
  assign \new_[70718]_  = A301 & A300;
  assign \new_[70719]_  = \new_[70718]_  & \new_[70715]_ ;
  assign \new_[70720]_  = \new_[70719]_  & \new_[70712]_ ;
  assign \new_[70724]_  = A167 & ~A169;
  assign \new_[70725]_  = A170 & \new_[70724]_ ;
  assign \new_[70728]_  = A199 & ~A166;
  assign \new_[70731]_  = ~A233 & A200;
  assign \new_[70732]_  = \new_[70731]_  & \new_[70728]_ ;
  assign \new_[70733]_  = \new_[70732]_  & \new_[70725]_ ;
  assign \new_[70736]_  = ~A236 & ~A235;
  assign \new_[70739]_  = ~A267 & ~A266;
  assign \new_[70740]_  = \new_[70739]_  & \new_[70736]_ ;
  assign \new_[70743]_  = ~A299 & A298;
  assign \new_[70746]_  = A302 & A300;
  assign \new_[70747]_  = \new_[70746]_  & \new_[70743]_ ;
  assign \new_[70748]_  = \new_[70747]_  & \new_[70740]_ ;
  assign \new_[70752]_  = A167 & ~A169;
  assign \new_[70753]_  = A170 & \new_[70752]_ ;
  assign \new_[70756]_  = A199 & ~A166;
  assign \new_[70759]_  = ~A233 & A200;
  assign \new_[70760]_  = \new_[70759]_  & \new_[70756]_ ;
  assign \new_[70761]_  = \new_[70760]_  & \new_[70753]_ ;
  assign \new_[70764]_  = ~A236 & ~A235;
  assign \new_[70767]_  = ~A266 & ~A265;
  assign \new_[70768]_  = \new_[70767]_  & \new_[70764]_ ;
  assign \new_[70771]_  = ~A299 & A298;
  assign \new_[70774]_  = A301 & A300;
  assign \new_[70775]_  = \new_[70774]_  & \new_[70771]_ ;
  assign \new_[70776]_  = \new_[70775]_  & \new_[70768]_ ;
  assign \new_[70780]_  = A167 & ~A169;
  assign \new_[70781]_  = A170 & \new_[70780]_ ;
  assign \new_[70784]_  = A199 & ~A166;
  assign \new_[70787]_  = ~A233 & A200;
  assign \new_[70788]_  = \new_[70787]_  & \new_[70784]_ ;
  assign \new_[70789]_  = \new_[70788]_  & \new_[70781]_ ;
  assign \new_[70792]_  = ~A236 & ~A235;
  assign \new_[70795]_  = ~A266 & ~A265;
  assign \new_[70796]_  = \new_[70795]_  & \new_[70792]_ ;
  assign \new_[70799]_  = ~A299 & A298;
  assign \new_[70802]_  = A302 & A300;
  assign \new_[70803]_  = \new_[70802]_  & \new_[70799]_ ;
  assign \new_[70804]_  = \new_[70803]_  & \new_[70796]_ ;
  assign \new_[70808]_  = A167 & ~A169;
  assign \new_[70809]_  = A170 & \new_[70808]_ ;
  assign \new_[70812]_  = A199 & ~A166;
  assign \new_[70815]_  = ~A233 & A200;
  assign \new_[70816]_  = \new_[70815]_  & \new_[70812]_ ;
  assign \new_[70817]_  = \new_[70816]_  & \new_[70809]_ ;
  assign \new_[70820]_  = ~A266 & ~A234;
  assign \new_[70823]_  = ~A269 & ~A268;
  assign \new_[70824]_  = \new_[70823]_  & \new_[70820]_ ;
  assign \new_[70827]_  = ~A299 & A298;
  assign \new_[70830]_  = A301 & A300;
  assign \new_[70831]_  = \new_[70830]_  & \new_[70827]_ ;
  assign \new_[70832]_  = \new_[70831]_  & \new_[70824]_ ;
  assign \new_[70836]_  = A167 & ~A169;
  assign \new_[70837]_  = A170 & \new_[70836]_ ;
  assign \new_[70840]_  = A199 & ~A166;
  assign \new_[70843]_  = ~A233 & A200;
  assign \new_[70844]_  = \new_[70843]_  & \new_[70840]_ ;
  assign \new_[70845]_  = \new_[70844]_  & \new_[70837]_ ;
  assign \new_[70848]_  = ~A266 & ~A234;
  assign \new_[70851]_  = ~A269 & ~A268;
  assign \new_[70852]_  = \new_[70851]_  & \new_[70848]_ ;
  assign \new_[70855]_  = ~A299 & A298;
  assign \new_[70858]_  = A302 & A300;
  assign \new_[70859]_  = \new_[70858]_  & \new_[70855]_ ;
  assign \new_[70860]_  = \new_[70859]_  & \new_[70852]_ ;
  assign \new_[70864]_  = A167 & ~A169;
  assign \new_[70865]_  = A170 & \new_[70864]_ ;
  assign \new_[70868]_  = A199 & ~A166;
  assign \new_[70871]_  = ~A232 & A200;
  assign \new_[70872]_  = \new_[70871]_  & \new_[70868]_ ;
  assign \new_[70873]_  = \new_[70872]_  & \new_[70865]_ ;
  assign \new_[70876]_  = ~A266 & ~A233;
  assign \new_[70879]_  = ~A269 & ~A268;
  assign \new_[70880]_  = \new_[70879]_  & \new_[70876]_ ;
  assign \new_[70883]_  = ~A299 & A298;
  assign \new_[70886]_  = A301 & A300;
  assign \new_[70887]_  = \new_[70886]_  & \new_[70883]_ ;
  assign \new_[70888]_  = \new_[70887]_  & \new_[70880]_ ;
  assign \new_[70892]_  = A167 & ~A169;
  assign \new_[70893]_  = A170 & \new_[70892]_ ;
  assign \new_[70896]_  = A199 & ~A166;
  assign \new_[70899]_  = ~A232 & A200;
  assign \new_[70900]_  = \new_[70899]_  & \new_[70896]_ ;
  assign \new_[70901]_  = \new_[70900]_  & \new_[70893]_ ;
  assign \new_[70904]_  = ~A266 & ~A233;
  assign \new_[70907]_  = ~A269 & ~A268;
  assign \new_[70908]_  = \new_[70907]_  & \new_[70904]_ ;
  assign \new_[70911]_  = ~A299 & A298;
  assign \new_[70914]_  = A302 & A300;
  assign \new_[70915]_  = \new_[70914]_  & \new_[70911]_ ;
  assign \new_[70916]_  = \new_[70915]_  & \new_[70908]_ ;
  assign \new_[70920]_  = A167 & ~A169;
  assign \new_[70921]_  = A170 & \new_[70920]_ ;
  assign \new_[70924]_  = ~A200 & ~A166;
  assign \new_[70927]_  = ~A203 & ~A202;
  assign \new_[70928]_  = \new_[70927]_  & \new_[70924]_ ;
  assign \new_[70929]_  = \new_[70928]_  & \new_[70921]_ ;
  assign \new_[70932]_  = A233 & A232;
  assign \new_[70935]_  = ~A267 & A265;
  assign \new_[70936]_  = \new_[70935]_  & \new_[70932]_ ;
  assign \new_[70939]_  = ~A299 & A298;
  assign \new_[70942]_  = A301 & A300;
  assign \new_[70943]_  = \new_[70942]_  & \new_[70939]_ ;
  assign \new_[70944]_  = \new_[70943]_  & \new_[70936]_ ;
  assign \new_[70948]_  = A167 & ~A169;
  assign \new_[70949]_  = A170 & \new_[70948]_ ;
  assign \new_[70952]_  = ~A200 & ~A166;
  assign \new_[70955]_  = ~A203 & ~A202;
  assign \new_[70956]_  = \new_[70955]_  & \new_[70952]_ ;
  assign \new_[70957]_  = \new_[70956]_  & \new_[70949]_ ;
  assign \new_[70960]_  = A233 & A232;
  assign \new_[70963]_  = ~A267 & A265;
  assign \new_[70964]_  = \new_[70963]_  & \new_[70960]_ ;
  assign \new_[70967]_  = ~A299 & A298;
  assign \new_[70970]_  = A302 & A300;
  assign \new_[70971]_  = \new_[70970]_  & \new_[70967]_ ;
  assign \new_[70972]_  = \new_[70971]_  & \new_[70964]_ ;
  assign \new_[70976]_  = A167 & ~A169;
  assign \new_[70977]_  = A170 & \new_[70976]_ ;
  assign \new_[70980]_  = ~A200 & ~A166;
  assign \new_[70983]_  = ~A203 & ~A202;
  assign \new_[70984]_  = \new_[70983]_  & \new_[70980]_ ;
  assign \new_[70985]_  = \new_[70984]_  & \new_[70977]_ ;
  assign \new_[70988]_  = A233 & A232;
  assign \new_[70991]_  = A266 & A265;
  assign \new_[70992]_  = \new_[70991]_  & \new_[70988]_ ;
  assign \new_[70995]_  = ~A299 & A298;
  assign \new_[70998]_  = A301 & A300;
  assign \new_[70999]_  = \new_[70998]_  & \new_[70995]_ ;
  assign \new_[71000]_  = \new_[70999]_  & \new_[70992]_ ;
  assign \new_[71004]_  = A167 & ~A169;
  assign \new_[71005]_  = A170 & \new_[71004]_ ;
  assign \new_[71008]_  = ~A200 & ~A166;
  assign \new_[71011]_  = ~A203 & ~A202;
  assign \new_[71012]_  = \new_[71011]_  & \new_[71008]_ ;
  assign \new_[71013]_  = \new_[71012]_  & \new_[71005]_ ;
  assign \new_[71016]_  = A233 & A232;
  assign \new_[71019]_  = A266 & A265;
  assign \new_[71020]_  = \new_[71019]_  & \new_[71016]_ ;
  assign \new_[71023]_  = ~A299 & A298;
  assign \new_[71026]_  = A302 & A300;
  assign \new_[71027]_  = \new_[71026]_  & \new_[71023]_ ;
  assign \new_[71028]_  = \new_[71027]_  & \new_[71020]_ ;
  assign \new_[71032]_  = A167 & ~A169;
  assign \new_[71033]_  = A170 & \new_[71032]_ ;
  assign \new_[71036]_  = ~A200 & ~A166;
  assign \new_[71039]_  = ~A203 & ~A202;
  assign \new_[71040]_  = \new_[71039]_  & \new_[71036]_ ;
  assign \new_[71041]_  = \new_[71040]_  & \new_[71033]_ ;
  assign \new_[71044]_  = A233 & A232;
  assign \new_[71047]_  = ~A266 & ~A265;
  assign \new_[71048]_  = \new_[71047]_  & \new_[71044]_ ;
  assign \new_[71051]_  = ~A299 & A298;
  assign \new_[71054]_  = A301 & A300;
  assign \new_[71055]_  = \new_[71054]_  & \new_[71051]_ ;
  assign \new_[71056]_  = \new_[71055]_  & \new_[71048]_ ;
  assign \new_[71060]_  = A167 & ~A169;
  assign \new_[71061]_  = A170 & \new_[71060]_ ;
  assign \new_[71064]_  = ~A200 & ~A166;
  assign \new_[71067]_  = ~A203 & ~A202;
  assign \new_[71068]_  = \new_[71067]_  & \new_[71064]_ ;
  assign \new_[71069]_  = \new_[71068]_  & \new_[71061]_ ;
  assign \new_[71072]_  = A233 & A232;
  assign \new_[71075]_  = ~A266 & ~A265;
  assign \new_[71076]_  = \new_[71075]_  & \new_[71072]_ ;
  assign \new_[71079]_  = ~A299 & A298;
  assign \new_[71082]_  = A302 & A300;
  assign \new_[71083]_  = \new_[71082]_  & \new_[71079]_ ;
  assign \new_[71084]_  = \new_[71083]_  & \new_[71076]_ ;
  assign \new_[71088]_  = A167 & ~A169;
  assign \new_[71089]_  = A170 & \new_[71088]_ ;
  assign \new_[71092]_  = ~A200 & ~A166;
  assign \new_[71095]_  = ~A203 & ~A202;
  assign \new_[71096]_  = \new_[71095]_  & \new_[71092]_ ;
  assign \new_[71097]_  = \new_[71096]_  & \new_[71089]_ ;
  assign \new_[71100]_  = ~A235 & ~A233;
  assign \new_[71103]_  = ~A266 & ~A236;
  assign \new_[71104]_  = \new_[71103]_  & \new_[71100]_ ;
  assign \new_[71107]_  = ~A269 & ~A268;
  assign \new_[71110]_  = A299 & ~A298;
  assign \new_[71111]_  = \new_[71110]_  & \new_[71107]_ ;
  assign \new_[71112]_  = \new_[71111]_  & \new_[71104]_ ;
  assign \new_[71116]_  = A167 & ~A169;
  assign \new_[71117]_  = A170 & \new_[71116]_ ;
  assign \new_[71120]_  = ~A200 & ~A166;
  assign \new_[71123]_  = ~A203 & ~A202;
  assign \new_[71124]_  = \new_[71123]_  & \new_[71120]_ ;
  assign \new_[71125]_  = \new_[71124]_  & \new_[71117]_ ;
  assign \new_[71128]_  = ~A234 & ~A233;
  assign \new_[71131]_  = A266 & A265;
  assign \new_[71132]_  = \new_[71131]_  & \new_[71128]_ ;
  assign \new_[71135]_  = ~A299 & A298;
  assign \new_[71138]_  = A301 & A300;
  assign \new_[71139]_  = \new_[71138]_  & \new_[71135]_ ;
  assign \new_[71140]_  = \new_[71139]_  & \new_[71132]_ ;
  assign \new_[71144]_  = A167 & ~A169;
  assign \new_[71145]_  = A170 & \new_[71144]_ ;
  assign \new_[71148]_  = ~A200 & ~A166;
  assign \new_[71151]_  = ~A203 & ~A202;
  assign \new_[71152]_  = \new_[71151]_  & \new_[71148]_ ;
  assign \new_[71153]_  = \new_[71152]_  & \new_[71145]_ ;
  assign \new_[71156]_  = ~A234 & ~A233;
  assign \new_[71159]_  = A266 & A265;
  assign \new_[71160]_  = \new_[71159]_  & \new_[71156]_ ;
  assign \new_[71163]_  = ~A299 & A298;
  assign \new_[71166]_  = A302 & A300;
  assign \new_[71167]_  = \new_[71166]_  & \new_[71163]_ ;
  assign \new_[71168]_  = \new_[71167]_  & \new_[71160]_ ;
  assign \new_[71172]_  = A167 & ~A169;
  assign \new_[71173]_  = A170 & \new_[71172]_ ;
  assign \new_[71176]_  = ~A200 & ~A166;
  assign \new_[71179]_  = ~A203 & ~A202;
  assign \new_[71180]_  = \new_[71179]_  & \new_[71176]_ ;
  assign \new_[71181]_  = \new_[71180]_  & \new_[71173]_ ;
  assign \new_[71184]_  = ~A234 & ~A233;
  assign \new_[71187]_  = ~A267 & ~A266;
  assign \new_[71188]_  = \new_[71187]_  & \new_[71184]_ ;
  assign \new_[71191]_  = ~A299 & A298;
  assign \new_[71194]_  = A301 & A300;
  assign \new_[71195]_  = \new_[71194]_  & \new_[71191]_ ;
  assign \new_[71196]_  = \new_[71195]_  & \new_[71188]_ ;
  assign \new_[71200]_  = A167 & ~A169;
  assign \new_[71201]_  = A170 & \new_[71200]_ ;
  assign \new_[71204]_  = ~A200 & ~A166;
  assign \new_[71207]_  = ~A203 & ~A202;
  assign \new_[71208]_  = \new_[71207]_  & \new_[71204]_ ;
  assign \new_[71209]_  = \new_[71208]_  & \new_[71201]_ ;
  assign \new_[71212]_  = ~A234 & ~A233;
  assign \new_[71215]_  = ~A267 & ~A266;
  assign \new_[71216]_  = \new_[71215]_  & \new_[71212]_ ;
  assign \new_[71219]_  = ~A299 & A298;
  assign \new_[71222]_  = A302 & A300;
  assign \new_[71223]_  = \new_[71222]_  & \new_[71219]_ ;
  assign \new_[71224]_  = \new_[71223]_  & \new_[71216]_ ;
  assign \new_[71228]_  = A167 & ~A169;
  assign \new_[71229]_  = A170 & \new_[71228]_ ;
  assign \new_[71232]_  = ~A200 & ~A166;
  assign \new_[71235]_  = ~A203 & ~A202;
  assign \new_[71236]_  = \new_[71235]_  & \new_[71232]_ ;
  assign \new_[71237]_  = \new_[71236]_  & \new_[71229]_ ;
  assign \new_[71240]_  = ~A234 & ~A233;
  assign \new_[71243]_  = ~A266 & ~A265;
  assign \new_[71244]_  = \new_[71243]_  & \new_[71240]_ ;
  assign \new_[71247]_  = ~A299 & A298;
  assign \new_[71250]_  = A301 & A300;
  assign \new_[71251]_  = \new_[71250]_  & \new_[71247]_ ;
  assign \new_[71252]_  = \new_[71251]_  & \new_[71244]_ ;
  assign \new_[71256]_  = A167 & ~A169;
  assign \new_[71257]_  = A170 & \new_[71256]_ ;
  assign \new_[71260]_  = ~A200 & ~A166;
  assign \new_[71263]_  = ~A203 & ~A202;
  assign \new_[71264]_  = \new_[71263]_  & \new_[71260]_ ;
  assign \new_[71265]_  = \new_[71264]_  & \new_[71257]_ ;
  assign \new_[71268]_  = ~A234 & ~A233;
  assign \new_[71271]_  = ~A266 & ~A265;
  assign \new_[71272]_  = \new_[71271]_  & \new_[71268]_ ;
  assign \new_[71275]_  = ~A299 & A298;
  assign \new_[71278]_  = A302 & A300;
  assign \new_[71279]_  = \new_[71278]_  & \new_[71275]_ ;
  assign \new_[71280]_  = \new_[71279]_  & \new_[71272]_ ;
  assign \new_[71284]_  = A167 & ~A169;
  assign \new_[71285]_  = A170 & \new_[71284]_ ;
  assign \new_[71288]_  = ~A200 & ~A166;
  assign \new_[71291]_  = ~A203 & ~A202;
  assign \new_[71292]_  = \new_[71291]_  & \new_[71288]_ ;
  assign \new_[71293]_  = \new_[71292]_  & \new_[71285]_ ;
  assign \new_[71296]_  = ~A233 & A232;
  assign \new_[71299]_  = A235 & A234;
  assign \new_[71300]_  = \new_[71299]_  & \new_[71296]_ ;
  assign \new_[71303]_  = ~A266 & A265;
  assign \new_[71306]_  = A268 & A267;
  assign \new_[71307]_  = \new_[71306]_  & \new_[71303]_ ;
  assign \new_[71308]_  = \new_[71307]_  & \new_[71300]_ ;
  assign \new_[71312]_  = A167 & ~A169;
  assign \new_[71313]_  = A170 & \new_[71312]_ ;
  assign \new_[71316]_  = ~A200 & ~A166;
  assign \new_[71319]_  = ~A203 & ~A202;
  assign \new_[71320]_  = \new_[71319]_  & \new_[71316]_ ;
  assign \new_[71321]_  = \new_[71320]_  & \new_[71313]_ ;
  assign \new_[71324]_  = ~A233 & A232;
  assign \new_[71327]_  = A235 & A234;
  assign \new_[71328]_  = \new_[71327]_  & \new_[71324]_ ;
  assign \new_[71331]_  = ~A266 & A265;
  assign \new_[71334]_  = A269 & A267;
  assign \new_[71335]_  = \new_[71334]_  & \new_[71331]_ ;
  assign \new_[71336]_  = \new_[71335]_  & \new_[71328]_ ;
  assign \new_[71340]_  = A167 & ~A169;
  assign \new_[71341]_  = A170 & \new_[71340]_ ;
  assign \new_[71344]_  = ~A200 & ~A166;
  assign \new_[71347]_  = ~A203 & ~A202;
  assign \new_[71348]_  = \new_[71347]_  & \new_[71344]_ ;
  assign \new_[71349]_  = \new_[71348]_  & \new_[71341]_ ;
  assign \new_[71352]_  = ~A233 & A232;
  assign \new_[71355]_  = A236 & A234;
  assign \new_[71356]_  = \new_[71355]_  & \new_[71352]_ ;
  assign \new_[71359]_  = ~A266 & A265;
  assign \new_[71362]_  = A268 & A267;
  assign \new_[71363]_  = \new_[71362]_  & \new_[71359]_ ;
  assign \new_[71364]_  = \new_[71363]_  & \new_[71356]_ ;
  assign \new_[71368]_  = A167 & ~A169;
  assign \new_[71369]_  = A170 & \new_[71368]_ ;
  assign \new_[71372]_  = ~A200 & ~A166;
  assign \new_[71375]_  = ~A203 & ~A202;
  assign \new_[71376]_  = \new_[71375]_  & \new_[71372]_ ;
  assign \new_[71377]_  = \new_[71376]_  & \new_[71369]_ ;
  assign \new_[71380]_  = ~A233 & A232;
  assign \new_[71383]_  = A236 & A234;
  assign \new_[71384]_  = \new_[71383]_  & \new_[71380]_ ;
  assign \new_[71387]_  = ~A266 & A265;
  assign \new_[71390]_  = A269 & A267;
  assign \new_[71391]_  = \new_[71390]_  & \new_[71387]_ ;
  assign \new_[71392]_  = \new_[71391]_  & \new_[71384]_ ;
  assign \new_[71396]_  = A167 & ~A169;
  assign \new_[71397]_  = A170 & \new_[71396]_ ;
  assign \new_[71400]_  = ~A200 & ~A166;
  assign \new_[71403]_  = ~A203 & ~A202;
  assign \new_[71404]_  = \new_[71403]_  & \new_[71400]_ ;
  assign \new_[71405]_  = \new_[71404]_  & \new_[71397]_ ;
  assign \new_[71408]_  = ~A233 & ~A232;
  assign \new_[71411]_  = A266 & A265;
  assign \new_[71412]_  = \new_[71411]_  & \new_[71408]_ ;
  assign \new_[71415]_  = ~A299 & A298;
  assign \new_[71418]_  = A301 & A300;
  assign \new_[71419]_  = \new_[71418]_  & \new_[71415]_ ;
  assign \new_[71420]_  = \new_[71419]_  & \new_[71412]_ ;
  assign \new_[71424]_  = A167 & ~A169;
  assign \new_[71425]_  = A170 & \new_[71424]_ ;
  assign \new_[71428]_  = ~A200 & ~A166;
  assign \new_[71431]_  = ~A203 & ~A202;
  assign \new_[71432]_  = \new_[71431]_  & \new_[71428]_ ;
  assign \new_[71433]_  = \new_[71432]_  & \new_[71425]_ ;
  assign \new_[71436]_  = ~A233 & ~A232;
  assign \new_[71439]_  = A266 & A265;
  assign \new_[71440]_  = \new_[71439]_  & \new_[71436]_ ;
  assign \new_[71443]_  = ~A299 & A298;
  assign \new_[71446]_  = A302 & A300;
  assign \new_[71447]_  = \new_[71446]_  & \new_[71443]_ ;
  assign \new_[71448]_  = \new_[71447]_  & \new_[71440]_ ;
  assign \new_[71452]_  = A167 & ~A169;
  assign \new_[71453]_  = A170 & \new_[71452]_ ;
  assign \new_[71456]_  = ~A200 & ~A166;
  assign \new_[71459]_  = ~A203 & ~A202;
  assign \new_[71460]_  = \new_[71459]_  & \new_[71456]_ ;
  assign \new_[71461]_  = \new_[71460]_  & \new_[71453]_ ;
  assign \new_[71464]_  = ~A233 & ~A232;
  assign \new_[71467]_  = ~A267 & ~A266;
  assign \new_[71468]_  = \new_[71467]_  & \new_[71464]_ ;
  assign \new_[71471]_  = ~A299 & A298;
  assign \new_[71474]_  = A301 & A300;
  assign \new_[71475]_  = \new_[71474]_  & \new_[71471]_ ;
  assign \new_[71476]_  = \new_[71475]_  & \new_[71468]_ ;
  assign \new_[71480]_  = A167 & ~A169;
  assign \new_[71481]_  = A170 & \new_[71480]_ ;
  assign \new_[71484]_  = ~A200 & ~A166;
  assign \new_[71487]_  = ~A203 & ~A202;
  assign \new_[71488]_  = \new_[71487]_  & \new_[71484]_ ;
  assign \new_[71489]_  = \new_[71488]_  & \new_[71481]_ ;
  assign \new_[71492]_  = ~A233 & ~A232;
  assign \new_[71495]_  = ~A267 & ~A266;
  assign \new_[71496]_  = \new_[71495]_  & \new_[71492]_ ;
  assign \new_[71499]_  = ~A299 & A298;
  assign \new_[71502]_  = A302 & A300;
  assign \new_[71503]_  = \new_[71502]_  & \new_[71499]_ ;
  assign \new_[71504]_  = \new_[71503]_  & \new_[71496]_ ;
  assign \new_[71508]_  = A167 & ~A169;
  assign \new_[71509]_  = A170 & \new_[71508]_ ;
  assign \new_[71512]_  = ~A200 & ~A166;
  assign \new_[71515]_  = ~A203 & ~A202;
  assign \new_[71516]_  = \new_[71515]_  & \new_[71512]_ ;
  assign \new_[71517]_  = \new_[71516]_  & \new_[71509]_ ;
  assign \new_[71520]_  = ~A233 & ~A232;
  assign \new_[71523]_  = ~A266 & ~A265;
  assign \new_[71524]_  = \new_[71523]_  & \new_[71520]_ ;
  assign \new_[71527]_  = ~A299 & A298;
  assign \new_[71530]_  = A301 & A300;
  assign \new_[71531]_  = \new_[71530]_  & \new_[71527]_ ;
  assign \new_[71532]_  = \new_[71531]_  & \new_[71524]_ ;
  assign \new_[71536]_  = A167 & ~A169;
  assign \new_[71537]_  = A170 & \new_[71536]_ ;
  assign \new_[71540]_  = ~A200 & ~A166;
  assign \new_[71543]_  = ~A203 & ~A202;
  assign \new_[71544]_  = \new_[71543]_  & \new_[71540]_ ;
  assign \new_[71545]_  = \new_[71544]_  & \new_[71537]_ ;
  assign \new_[71548]_  = ~A233 & ~A232;
  assign \new_[71551]_  = ~A266 & ~A265;
  assign \new_[71552]_  = \new_[71551]_  & \new_[71548]_ ;
  assign \new_[71555]_  = ~A299 & A298;
  assign \new_[71558]_  = A302 & A300;
  assign \new_[71559]_  = \new_[71558]_  & \new_[71555]_ ;
  assign \new_[71560]_  = \new_[71559]_  & \new_[71552]_ ;
  assign \new_[71564]_  = A167 & ~A169;
  assign \new_[71565]_  = A170 & \new_[71564]_ ;
  assign \new_[71568]_  = ~A200 & ~A166;
  assign \new_[71571]_  = A232 & ~A201;
  assign \new_[71572]_  = \new_[71571]_  & \new_[71568]_ ;
  assign \new_[71573]_  = \new_[71572]_  & \new_[71565]_ ;
  assign \new_[71576]_  = A265 & A233;
  assign \new_[71579]_  = ~A269 & ~A268;
  assign \new_[71580]_  = \new_[71579]_  & \new_[71576]_ ;
  assign \new_[71583]_  = ~A299 & A298;
  assign \new_[71586]_  = A301 & A300;
  assign \new_[71587]_  = \new_[71586]_  & \new_[71583]_ ;
  assign \new_[71588]_  = \new_[71587]_  & \new_[71580]_ ;
  assign \new_[71592]_  = A167 & ~A169;
  assign \new_[71593]_  = A170 & \new_[71592]_ ;
  assign \new_[71596]_  = ~A200 & ~A166;
  assign \new_[71599]_  = A232 & ~A201;
  assign \new_[71600]_  = \new_[71599]_  & \new_[71596]_ ;
  assign \new_[71601]_  = \new_[71600]_  & \new_[71593]_ ;
  assign \new_[71604]_  = A265 & A233;
  assign \new_[71607]_  = ~A269 & ~A268;
  assign \new_[71608]_  = \new_[71607]_  & \new_[71604]_ ;
  assign \new_[71611]_  = ~A299 & A298;
  assign \new_[71614]_  = A302 & A300;
  assign \new_[71615]_  = \new_[71614]_  & \new_[71611]_ ;
  assign \new_[71616]_  = \new_[71615]_  & \new_[71608]_ ;
  assign \new_[71620]_  = A167 & ~A169;
  assign \new_[71621]_  = A170 & \new_[71620]_ ;
  assign \new_[71624]_  = ~A200 & ~A166;
  assign \new_[71627]_  = ~A233 & ~A201;
  assign \new_[71628]_  = \new_[71627]_  & \new_[71624]_ ;
  assign \new_[71629]_  = \new_[71628]_  & \new_[71621]_ ;
  assign \new_[71632]_  = ~A236 & ~A235;
  assign \new_[71635]_  = A266 & A265;
  assign \new_[71636]_  = \new_[71635]_  & \new_[71632]_ ;
  assign \new_[71639]_  = ~A299 & A298;
  assign \new_[71642]_  = A301 & A300;
  assign \new_[71643]_  = \new_[71642]_  & \new_[71639]_ ;
  assign \new_[71644]_  = \new_[71643]_  & \new_[71636]_ ;
  assign \new_[71648]_  = A167 & ~A169;
  assign \new_[71649]_  = A170 & \new_[71648]_ ;
  assign \new_[71652]_  = ~A200 & ~A166;
  assign \new_[71655]_  = ~A233 & ~A201;
  assign \new_[71656]_  = \new_[71655]_  & \new_[71652]_ ;
  assign \new_[71657]_  = \new_[71656]_  & \new_[71649]_ ;
  assign \new_[71660]_  = ~A236 & ~A235;
  assign \new_[71663]_  = A266 & A265;
  assign \new_[71664]_  = \new_[71663]_  & \new_[71660]_ ;
  assign \new_[71667]_  = ~A299 & A298;
  assign \new_[71670]_  = A302 & A300;
  assign \new_[71671]_  = \new_[71670]_  & \new_[71667]_ ;
  assign \new_[71672]_  = \new_[71671]_  & \new_[71664]_ ;
  assign \new_[71676]_  = A167 & ~A169;
  assign \new_[71677]_  = A170 & \new_[71676]_ ;
  assign \new_[71680]_  = ~A200 & ~A166;
  assign \new_[71683]_  = ~A233 & ~A201;
  assign \new_[71684]_  = \new_[71683]_  & \new_[71680]_ ;
  assign \new_[71685]_  = \new_[71684]_  & \new_[71677]_ ;
  assign \new_[71688]_  = ~A236 & ~A235;
  assign \new_[71691]_  = ~A267 & ~A266;
  assign \new_[71692]_  = \new_[71691]_  & \new_[71688]_ ;
  assign \new_[71695]_  = ~A299 & A298;
  assign \new_[71698]_  = A301 & A300;
  assign \new_[71699]_  = \new_[71698]_  & \new_[71695]_ ;
  assign \new_[71700]_  = \new_[71699]_  & \new_[71692]_ ;
  assign \new_[71704]_  = A167 & ~A169;
  assign \new_[71705]_  = A170 & \new_[71704]_ ;
  assign \new_[71708]_  = ~A200 & ~A166;
  assign \new_[71711]_  = ~A233 & ~A201;
  assign \new_[71712]_  = \new_[71711]_  & \new_[71708]_ ;
  assign \new_[71713]_  = \new_[71712]_  & \new_[71705]_ ;
  assign \new_[71716]_  = ~A236 & ~A235;
  assign \new_[71719]_  = ~A267 & ~A266;
  assign \new_[71720]_  = \new_[71719]_  & \new_[71716]_ ;
  assign \new_[71723]_  = ~A299 & A298;
  assign \new_[71726]_  = A302 & A300;
  assign \new_[71727]_  = \new_[71726]_  & \new_[71723]_ ;
  assign \new_[71728]_  = \new_[71727]_  & \new_[71720]_ ;
  assign \new_[71732]_  = A167 & ~A169;
  assign \new_[71733]_  = A170 & \new_[71732]_ ;
  assign \new_[71736]_  = ~A200 & ~A166;
  assign \new_[71739]_  = ~A233 & ~A201;
  assign \new_[71740]_  = \new_[71739]_  & \new_[71736]_ ;
  assign \new_[71741]_  = \new_[71740]_  & \new_[71733]_ ;
  assign \new_[71744]_  = ~A236 & ~A235;
  assign \new_[71747]_  = ~A266 & ~A265;
  assign \new_[71748]_  = \new_[71747]_  & \new_[71744]_ ;
  assign \new_[71751]_  = ~A299 & A298;
  assign \new_[71754]_  = A301 & A300;
  assign \new_[71755]_  = \new_[71754]_  & \new_[71751]_ ;
  assign \new_[71756]_  = \new_[71755]_  & \new_[71748]_ ;
  assign \new_[71760]_  = A167 & ~A169;
  assign \new_[71761]_  = A170 & \new_[71760]_ ;
  assign \new_[71764]_  = ~A200 & ~A166;
  assign \new_[71767]_  = ~A233 & ~A201;
  assign \new_[71768]_  = \new_[71767]_  & \new_[71764]_ ;
  assign \new_[71769]_  = \new_[71768]_  & \new_[71761]_ ;
  assign \new_[71772]_  = ~A236 & ~A235;
  assign \new_[71775]_  = ~A266 & ~A265;
  assign \new_[71776]_  = \new_[71775]_  & \new_[71772]_ ;
  assign \new_[71779]_  = ~A299 & A298;
  assign \new_[71782]_  = A302 & A300;
  assign \new_[71783]_  = \new_[71782]_  & \new_[71779]_ ;
  assign \new_[71784]_  = \new_[71783]_  & \new_[71776]_ ;
  assign \new_[71788]_  = A167 & ~A169;
  assign \new_[71789]_  = A170 & \new_[71788]_ ;
  assign \new_[71792]_  = ~A200 & ~A166;
  assign \new_[71795]_  = ~A233 & ~A201;
  assign \new_[71796]_  = \new_[71795]_  & \new_[71792]_ ;
  assign \new_[71797]_  = \new_[71796]_  & \new_[71789]_ ;
  assign \new_[71800]_  = ~A266 & ~A234;
  assign \new_[71803]_  = ~A269 & ~A268;
  assign \new_[71804]_  = \new_[71803]_  & \new_[71800]_ ;
  assign \new_[71807]_  = ~A299 & A298;
  assign \new_[71810]_  = A301 & A300;
  assign \new_[71811]_  = \new_[71810]_  & \new_[71807]_ ;
  assign \new_[71812]_  = \new_[71811]_  & \new_[71804]_ ;
  assign \new_[71816]_  = A167 & ~A169;
  assign \new_[71817]_  = A170 & \new_[71816]_ ;
  assign \new_[71820]_  = ~A200 & ~A166;
  assign \new_[71823]_  = ~A233 & ~A201;
  assign \new_[71824]_  = \new_[71823]_  & \new_[71820]_ ;
  assign \new_[71825]_  = \new_[71824]_  & \new_[71817]_ ;
  assign \new_[71828]_  = ~A266 & ~A234;
  assign \new_[71831]_  = ~A269 & ~A268;
  assign \new_[71832]_  = \new_[71831]_  & \new_[71828]_ ;
  assign \new_[71835]_  = ~A299 & A298;
  assign \new_[71838]_  = A302 & A300;
  assign \new_[71839]_  = \new_[71838]_  & \new_[71835]_ ;
  assign \new_[71840]_  = \new_[71839]_  & \new_[71832]_ ;
  assign \new_[71844]_  = A167 & ~A169;
  assign \new_[71845]_  = A170 & \new_[71844]_ ;
  assign \new_[71848]_  = ~A200 & ~A166;
  assign \new_[71851]_  = ~A232 & ~A201;
  assign \new_[71852]_  = \new_[71851]_  & \new_[71848]_ ;
  assign \new_[71853]_  = \new_[71852]_  & \new_[71845]_ ;
  assign \new_[71856]_  = ~A266 & ~A233;
  assign \new_[71859]_  = ~A269 & ~A268;
  assign \new_[71860]_  = \new_[71859]_  & \new_[71856]_ ;
  assign \new_[71863]_  = ~A299 & A298;
  assign \new_[71866]_  = A301 & A300;
  assign \new_[71867]_  = \new_[71866]_  & \new_[71863]_ ;
  assign \new_[71868]_  = \new_[71867]_  & \new_[71860]_ ;
  assign \new_[71872]_  = A167 & ~A169;
  assign \new_[71873]_  = A170 & \new_[71872]_ ;
  assign \new_[71876]_  = ~A200 & ~A166;
  assign \new_[71879]_  = ~A232 & ~A201;
  assign \new_[71880]_  = \new_[71879]_  & \new_[71876]_ ;
  assign \new_[71881]_  = \new_[71880]_  & \new_[71873]_ ;
  assign \new_[71884]_  = ~A266 & ~A233;
  assign \new_[71887]_  = ~A269 & ~A268;
  assign \new_[71888]_  = \new_[71887]_  & \new_[71884]_ ;
  assign \new_[71891]_  = ~A299 & A298;
  assign \new_[71894]_  = A302 & A300;
  assign \new_[71895]_  = \new_[71894]_  & \new_[71891]_ ;
  assign \new_[71896]_  = \new_[71895]_  & \new_[71888]_ ;
  assign \new_[71900]_  = A167 & ~A169;
  assign \new_[71901]_  = A170 & \new_[71900]_ ;
  assign \new_[71904]_  = ~A199 & ~A166;
  assign \new_[71907]_  = A232 & ~A200;
  assign \new_[71908]_  = \new_[71907]_  & \new_[71904]_ ;
  assign \new_[71909]_  = \new_[71908]_  & \new_[71901]_ ;
  assign \new_[71912]_  = A265 & A233;
  assign \new_[71915]_  = ~A269 & ~A268;
  assign \new_[71916]_  = \new_[71915]_  & \new_[71912]_ ;
  assign \new_[71919]_  = ~A299 & A298;
  assign \new_[71922]_  = A301 & A300;
  assign \new_[71923]_  = \new_[71922]_  & \new_[71919]_ ;
  assign \new_[71924]_  = \new_[71923]_  & \new_[71916]_ ;
  assign \new_[71928]_  = A167 & ~A169;
  assign \new_[71929]_  = A170 & \new_[71928]_ ;
  assign \new_[71932]_  = ~A199 & ~A166;
  assign \new_[71935]_  = A232 & ~A200;
  assign \new_[71936]_  = \new_[71935]_  & \new_[71932]_ ;
  assign \new_[71937]_  = \new_[71936]_  & \new_[71929]_ ;
  assign \new_[71940]_  = A265 & A233;
  assign \new_[71943]_  = ~A269 & ~A268;
  assign \new_[71944]_  = \new_[71943]_  & \new_[71940]_ ;
  assign \new_[71947]_  = ~A299 & A298;
  assign \new_[71950]_  = A302 & A300;
  assign \new_[71951]_  = \new_[71950]_  & \new_[71947]_ ;
  assign \new_[71952]_  = \new_[71951]_  & \new_[71944]_ ;
  assign \new_[71956]_  = A167 & ~A169;
  assign \new_[71957]_  = A170 & \new_[71956]_ ;
  assign \new_[71960]_  = ~A199 & ~A166;
  assign \new_[71963]_  = ~A233 & ~A200;
  assign \new_[71964]_  = \new_[71963]_  & \new_[71960]_ ;
  assign \new_[71965]_  = \new_[71964]_  & \new_[71957]_ ;
  assign \new_[71968]_  = ~A236 & ~A235;
  assign \new_[71971]_  = A266 & A265;
  assign \new_[71972]_  = \new_[71971]_  & \new_[71968]_ ;
  assign \new_[71975]_  = ~A299 & A298;
  assign \new_[71978]_  = A301 & A300;
  assign \new_[71979]_  = \new_[71978]_  & \new_[71975]_ ;
  assign \new_[71980]_  = \new_[71979]_  & \new_[71972]_ ;
  assign \new_[71984]_  = A167 & ~A169;
  assign \new_[71985]_  = A170 & \new_[71984]_ ;
  assign \new_[71988]_  = ~A199 & ~A166;
  assign \new_[71991]_  = ~A233 & ~A200;
  assign \new_[71992]_  = \new_[71991]_  & \new_[71988]_ ;
  assign \new_[71993]_  = \new_[71992]_  & \new_[71985]_ ;
  assign \new_[71996]_  = ~A236 & ~A235;
  assign \new_[71999]_  = A266 & A265;
  assign \new_[72000]_  = \new_[71999]_  & \new_[71996]_ ;
  assign \new_[72003]_  = ~A299 & A298;
  assign \new_[72006]_  = A302 & A300;
  assign \new_[72007]_  = \new_[72006]_  & \new_[72003]_ ;
  assign \new_[72008]_  = \new_[72007]_  & \new_[72000]_ ;
  assign \new_[72012]_  = A167 & ~A169;
  assign \new_[72013]_  = A170 & \new_[72012]_ ;
  assign \new_[72016]_  = ~A199 & ~A166;
  assign \new_[72019]_  = ~A233 & ~A200;
  assign \new_[72020]_  = \new_[72019]_  & \new_[72016]_ ;
  assign \new_[72021]_  = \new_[72020]_  & \new_[72013]_ ;
  assign \new_[72024]_  = ~A236 & ~A235;
  assign \new_[72027]_  = ~A267 & ~A266;
  assign \new_[72028]_  = \new_[72027]_  & \new_[72024]_ ;
  assign \new_[72031]_  = ~A299 & A298;
  assign \new_[72034]_  = A301 & A300;
  assign \new_[72035]_  = \new_[72034]_  & \new_[72031]_ ;
  assign \new_[72036]_  = \new_[72035]_  & \new_[72028]_ ;
  assign \new_[72040]_  = A167 & ~A169;
  assign \new_[72041]_  = A170 & \new_[72040]_ ;
  assign \new_[72044]_  = ~A199 & ~A166;
  assign \new_[72047]_  = ~A233 & ~A200;
  assign \new_[72048]_  = \new_[72047]_  & \new_[72044]_ ;
  assign \new_[72049]_  = \new_[72048]_  & \new_[72041]_ ;
  assign \new_[72052]_  = ~A236 & ~A235;
  assign \new_[72055]_  = ~A267 & ~A266;
  assign \new_[72056]_  = \new_[72055]_  & \new_[72052]_ ;
  assign \new_[72059]_  = ~A299 & A298;
  assign \new_[72062]_  = A302 & A300;
  assign \new_[72063]_  = \new_[72062]_  & \new_[72059]_ ;
  assign \new_[72064]_  = \new_[72063]_  & \new_[72056]_ ;
  assign \new_[72068]_  = A167 & ~A169;
  assign \new_[72069]_  = A170 & \new_[72068]_ ;
  assign \new_[72072]_  = ~A199 & ~A166;
  assign \new_[72075]_  = ~A233 & ~A200;
  assign \new_[72076]_  = \new_[72075]_  & \new_[72072]_ ;
  assign \new_[72077]_  = \new_[72076]_  & \new_[72069]_ ;
  assign \new_[72080]_  = ~A236 & ~A235;
  assign \new_[72083]_  = ~A266 & ~A265;
  assign \new_[72084]_  = \new_[72083]_  & \new_[72080]_ ;
  assign \new_[72087]_  = ~A299 & A298;
  assign \new_[72090]_  = A301 & A300;
  assign \new_[72091]_  = \new_[72090]_  & \new_[72087]_ ;
  assign \new_[72092]_  = \new_[72091]_  & \new_[72084]_ ;
  assign \new_[72096]_  = A167 & ~A169;
  assign \new_[72097]_  = A170 & \new_[72096]_ ;
  assign \new_[72100]_  = ~A199 & ~A166;
  assign \new_[72103]_  = ~A233 & ~A200;
  assign \new_[72104]_  = \new_[72103]_  & \new_[72100]_ ;
  assign \new_[72105]_  = \new_[72104]_  & \new_[72097]_ ;
  assign \new_[72108]_  = ~A236 & ~A235;
  assign \new_[72111]_  = ~A266 & ~A265;
  assign \new_[72112]_  = \new_[72111]_  & \new_[72108]_ ;
  assign \new_[72115]_  = ~A299 & A298;
  assign \new_[72118]_  = A302 & A300;
  assign \new_[72119]_  = \new_[72118]_  & \new_[72115]_ ;
  assign \new_[72120]_  = \new_[72119]_  & \new_[72112]_ ;
  assign \new_[72124]_  = A167 & ~A169;
  assign \new_[72125]_  = A170 & \new_[72124]_ ;
  assign \new_[72128]_  = ~A199 & ~A166;
  assign \new_[72131]_  = ~A233 & ~A200;
  assign \new_[72132]_  = \new_[72131]_  & \new_[72128]_ ;
  assign \new_[72133]_  = \new_[72132]_  & \new_[72125]_ ;
  assign \new_[72136]_  = ~A266 & ~A234;
  assign \new_[72139]_  = ~A269 & ~A268;
  assign \new_[72140]_  = \new_[72139]_  & \new_[72136]_ ;
  assign \new_[72143]_  = ~A299 & A298;
  assign \new_[72146]_  = A301 & A300;
  assign \new_[72147]_  = \new_[72146]_  & \new_[72143]_ ;
  assign \new_[72148]_  = \new_[72147]_  & \new_[72140]_ ;
  assign \new_[72152]_  = A167 & ~A169;
  assign \new_[72153]_  = A170 & \new_[72152]_ ;
  assign \new_[72156]_  = ~A199 & ~A166;
  assign \new_[72159]_  = ~A233 & ~A200;
  assign \new_[72160]_  = \new_[72159]_  & \new_[72156]_ ;
  assign \new_[72161]_  = \new_[72160]_  & \new_[72153]_ ;
  assign \new_[72164]_  = ~A266 & ~A234;
  assign \new_[72167]_  = ~A269 & ~A268;
  assign \new_[72168]_  = \new_[72167]_  & \new_[72164]_ ;
  assign \new_[72171]_  = ~A299 & A298;
  assign \new_[72174]_  = A302 & A300;
  assign \new_[72175]_  = \new_[72174]_  & \new_[72171]_ ;
  assign \new_[72176]_  = \new_[72175]_  & \new_[72168]_ ;
  assign \new_[72180]_  = A167 & ~A169;
  assign \new_[72181]_  = A170 & \new_[72180]_ ;
  assign \new_[72184]_  = ~A199 & ~A166;
  assign \new_[72187]_  = ~A232 & ~A200;
  assign \new_[72188]_  = \new_[72187]_  & \new_[72184]_ ;
  assign \new_[72189]_  = \new_[72188]_  & \new_[72181]_ ;
  assign \new_[72192]_  = ~A266 & ~A233;
  assign \new_[72195]_  = ~A269 & ~A268;
  assign \new_[72196]_  = \new_[72195]_  & \new_[72192]_ ;
  assign \new_[72199]_  = ~A299 & A298;
  assign \new_[72202]_  = A301 & A300;
  assign \new_[72203]_  = \new_[72202]_  & \new_[72199]_ ;
  assign \new_[72204]_  = \new_[72203]_  & \new_[72196]_ ;
  assign \new_[72208]_  = A167 & ~A169;
  assign \new_[72209]_  = A170 & \new_[72208]_ ;
  assign \new_[72212]_  = ~A199 & ~A166;
  assign \new_[72215]_  = ~A232 & ~A200;
  assign \new_[72216]_  = \new_[72215]_  & \new_[72212]_ ;
  assign \new_[72217]_  = \new_[72216]_  & \new_[72209]_ ;
  assign \new_[72220]_  = ~A266 & ~A233;
  assign \new_[72223]_  = ~A269 & ~A268;
  assign \new_[72224]_  = \new_[72223]_  & \new_[72220]_ ;
  assign \new_[72227]_  = ~A299 & A298;
  assign \new_[72230]_  = A302 & A300;
  assign \new_[72231]_  = \new_[72230]_  & \new_[72227]_ ;
  assign \new_[72232]_  = \new_[72231]_  & \new_[72224]_ ;
  assign \new_[72236]_  = ~A167 & ~A169;
  assign \new_[72237]_  = A170 & \new_[72236]_ ;
  assign \new_[72240]_  = A199 & A166;
  assign \new_[72243]_  = A232 & A200;
  assign \new_[72244]_  = \new_[72243]_  & \new_[72240]_ ;
  assign \new_[72245]_  = \new_[72244]_  & \new_[72237]_ ;
  assign \new_[72248]_  = A265 & A233;
  assign \new_[72251]_  = ~A269 & ~A268;
  assign \new_[72252]_  = \new_[72251]_  & \new_[72248]_ ;
  assign \new_[72255]_  = ~A299 & A298;
  assign \new_[72258]_  = A301 & A300;
  assign \new_[72259]_  = \new_[72258]_  & \new_[72255]_ ;
  assign \new_[72260]_  = \new_[72259]_  & \new_[72252]_ ;
  assign \new_[72264]_  = ~A167 & ~A169;
  assign \new_[72265]_  = A170 & \new_[72264]_ ;
  assign \new_[72268]_  = A199 & A166;
  assign \new_[72271]_  = A232 & A200;
  assign \new_[72272]_  = \new_[72271]_  & \new_[72268]_ ;
  assign \new_[72273]_  = \new_[72272]_  & \new_[72265]_ ;
  assign \new_[72276]_  = A265 & A233;
  assign \new_[72279]_  = ~A269 & ~A268;
  assign \new_[72280]_  = \new_[72279]_  & \new_[72276]_ ;
  assign \new_[72283]_  = ~A299 & A298;
  assign \new_[72286]_  = A302 & A300;
  assign \new_[72287]_  = \new_[72286]_  & \new_[72283]_ ;
  assign \new_[72288]_  = \new_[72287]_  & \new_[72280]_ ;
  assign \new_[72292]_  = ~A167 & ~A169;
  assign \new_[72293]_  = A170 & \new_[72292]_ ;
  assign \new_[72296]_  = A199 & A166;
  assign \new_[72299]_  = ~A233 & A200;
  assign \new_[72300]_  = \new_[72299]_  & \new_[72296]_ ;
  assign \new_[72301]_  = \new_[72300]_  & \new_[72293]_ ;
  assign \new_[72304]_  = ~A236 & ~A235;
  assign \new_[72307]_  = A266 & A265;
  assign \new_[72308]_  = \new_[72307]_  & \new_[72304]_ ;
  assign \new_[72311]_  = ~A299 & A298;
  assign \new_[72314]_  = A301 & A300;
  assign \new_[72315]_  = \new_[72314]_  & \new_[72311]_ ;
  assign \new_[72316]_  = \new_[72315]_  & \new_[72308]_ ;
  assign \new_[72320]_  = ~A167 & ~A169;
  assign \new_[72321]_  = A170 & \new_[72320]_ ;
  assign \new_[72324]_  = A199 & A166;
  assign \new_[72327]_  = ~A233 & A200;
  assign \new_[72328]_  = \new_[72327]_  & \new_[72324]_ ;
  assign \new_[72329]_  = \new_[72328]_  & \new_[72321]_ ;
  assign \new_[72332]_  = ~A236 & ~A235;
  assign \new_[72335]_  = A266 & A265;
  assign \new_[72336]_  = \new_[72335]_  & \new_[72332]_ ;
  assign \new_[72339]_  = ~A299 & A298;
  assign \new_[72342]_  = A302 & A300;
  assign \new_[72343]_  = \new_[72342]_  & \new_[72339]_ ;
  assign \new_[72344]_  = \new_[72343]_  & \new_[72336]_ ;
  assign \new_[72348]_  = ~A167 & ~A169;
  assign \new_[72349]_  = A170 & \new_[72348]_ ;
  assign \new_[72352]_  = A199 & A166;
  assign \new_[72355]_  = ~A233 & A200;
  assign \new_[72356]_  = \new_[72355]_  & \new_[72352]_ ;
  assign \new_[72357]_  = \new_[72356]_  & \new_[72349]_ ;
  assign \new_[72360]_  = ~A236 & ~A235;
  assign \new_[72363]_  = ~A267 & ~A266;
  assign \new_[72364]_  = \new_[72363]_  & \new_[72360]_ ;
  assign \new_[72367]_  = ~A299 & A298;
  assign \new_[72370]_  = A301 & A300;
  assign \new_[72371]_  = \new_[72370]_  & \new_[72367]_ ;
  assign \new_[72372]_  = \new_[72371]_  & \new_[72364]_ ;
  assign \new_[72376]_  = ~A167 & ~A169;
  assign \new_[72377]_  = A170 & \new_[72376]_ ;
  assign \new_[72380]_  = A199 & A166;
  assign \new_[72383]_  = ~A233 & A200;
  assign \new_[72384]_  = \new_[72383]_  & \new_[72380]_ ;
  assign \new_[72385]_  = \new_[72384]_  & \new_[72377]_ ;
  assign \new_[72388]_  = ~A236 & ~A235;
  assign \new_[72391]_  = ~A267 & ~A266;
  assign \new_[72392]_  = \new_[72391]_  & \new_[72388]_ ;
  assign \new_[72395]_  = ~A299 & A298;
  assign \new_[72398]_  = A302 & A300;
  assign \new_[72399]_  = \new_[72398]_  & \new_[72395]_ ;
  assign \new_[72400]_  = \new_[72399]_  & \new_[72392]_ ;
  assign \new_[72404]_  = ~A167 & ~A169;
  assign \new_[72405]_  = A170 & \new_[72404]_ ;
  assign \new_[72408]_  = A199 & A166;
  assign \new_[72411]_  = ~A233 & A200;
  assign \new_[72412]_  = \new_[72411]_  & \new_[72408]_ ;
  assign \new_[72413]_  = \new_[72412]_  & \new_[72405]_ ;
  assign \new_[72416]_  = ~A236 & ~A235;
  assign \new_[72419]_  = ~A266 & ~A265;
  assign \new_[72420]_  = \new_[72419]_  & \new_[72416]_ ;
  assign \new_[72423]_  = ~A299 & A298;
  assign \new_[72426]_  = A301 & A300;
  assign \new_[72427]_  = \new_[72426]_  & \new_[72423]_ ;
  assign \new_[72428]_  = \new_[72427]_  & \new_[72420]_ ;
  assign \new_[72432]_  = ~A167 & ~A169;
  assign \new_[72433]_  = A170 & \new_[72432]_ ;
  assign \new_[72436]_  = A199 & A166;
  assign \new_[72439]_  = ~A233 & A200;
  assign \new_[72440]_  = \new_[72439]_  & \new_[72436]_ ;
  assign \new_[72441]_  = \new_[72440]_  & \new_[72433]_ ;
  assign \new_[72444]_  = ~A236 & ~A235;
  assign \new_[72447]_  = ~A266 & ~A265;
  assign \new_[72448]_  = \new_[72447]_  & \new_[72444]_ ;
  assign \new_[72451]_  = ~A299 & A298;
  assign \new_[72454]_  = A302 & A300;
  assign \new_[72455]_  = \new_[72454]_  & \new_[72451]_ ;
  assign \new_[72456]_  = \new_[72455]_  & \new_[72448]_ ;
  assign \new_[72460]_  = ~A167 & ~A169;
  assign \new_[72461]_  = A170 & \new_[72460]_ ;
  assign \new_[72464]_  = A199 & A166;
  assign \new_[72467]_  = ~A233 & A200;
  assign \new_[72468]_  = \new_[72467]_  & \new_[72464]_ ;
  assign \new_[72469]_  = \new_[72468]_  & \new_[72461]_ ;
  assign \new_[72472]_  = ~A266 & ~A234;
  assign \new_[72475]_  = ~A269 & ~A268;
  assign \new_[72476]_  = \new_[72475]_  & \new_[72472]_ ;
  assign \new_[72479]_  = ~A299 & A298;
  assign \new_[72482]_  = A301 & A300;
  assign \new_[72483]_  = \new_[72482]_  & \new_[72479]_ ;
  assign \new_[72484]_  = \new_[72483]_  & \new_[72476]_ ;
  assign \new_[72488]_  = ~A167 & ~A169;
  assign \new_[72489]_  = A170 & \new_[72488]_ ;
  assign \new_[72492]_  = A199 & A166;
  assign \new_[72495]_  = ~A233 & A200;
  assign \new_[72496]_  = \new_[72495]_  & \new_[72492]_ ;
  assign \new_[72497]_  = \new_[72496]_  & \new_[72489]_ ;
  assign \new_[72500]_  = ~A266 & ~A234;
  assign \new_[72503]_  = ~A269 & ~A268;
  assign \new_[72504]_  = \new_[72503]_  & \new_[72500]_ ;
  assign \new_[72507]_  = ~A299 & A298;
  assign \new_[72510]_  = A302 & A300;
  assign \new_[72511]_  = \new_[72510]_  & \new_[72507]_ ;
  assign \new_[72512]_  = \new_[72511]_  & \new_[72504]_ ;
  assign \new_[72516]_  = ~A167 & ~A169;
  assign \new_[72517]_  = A170 & \new_[72516]_ ;
  assign \new_[72520]_  = A199 & A166;
  assign \new_[72523]_  = ~A232 & A200;
  assign \new_[72524]_  = \new_[72523]_  & \new_[72520]_ ;
  assign \new_[72525]_  = \new_[72524]_  & \new_[72517]_ ;
  assign \new_[72528]_  = ~A266 & ~A233;
  assign \new_[72531]_  = ~A269 & ~A268;
  assign \new_[72532]_  = \new_[72531]_  & \new_[72528]_ ;
  assign \new_[72535]_  = ~A299 & A298;
  assign \new_[72538]_  = A301 & A300;
  assign \new_[72539]_  = \new_[72538]_  & \new_[72535]_ ;
  assign \new_[72540]_  = \new_[72539]_  & \new_[72532]_ ;
  assign \new_[72544]_  = ~A167 & ~A169;
  assign \new_[72545]_  = A170 & \new_[72544]_ ;
  assign \new_[72548]_  = A199 & A166;
  assign \new_[72551]_  = ~A232 & A200;
  assign \new_[72552]_  = \new_[72551]_  & \new_[72548]_ ;
  assign \new_[72553]_  = \new_[72552]_  & \new_[72545]_ ;
  assign \new_[72556]_  = ~A266 & ~A233;
  assign \new_[72559]_  = ~A269 & ~A268;
  assign \new_[72560]_  = \new_[72559]_  & \new_[72556]_ ;
  assign \new_[72563]_  = ~A299 & A298;
  assign \new_[72566]_  = A302 & A300;
  assign \new_[72567]_  = \new_[72566]_  & \new_[72563]_ ;
  assign \new_[72568]_  = \new_[72567]_  & \new_[72560]_ ;
  assign \new_[72572]_  = ~A167 & ~A169;
  assign \new_[72573]_  = A170 & \new_[72572]_ ;
  assign \new_[72576]_  = ~A200 & A166;
  assign \new_[72579]_  = ~A203 & ~A202;
  assign \new_[72580]_  = \new_[72579]_  & \new_[72576]_ ;
  assign \new_[72581]_  = \new_[72580]_  & \new_[72573]_ ;
  assign \new_[72584]_  = A233 & A232;
  assign \new_[72587]_  = ~A267 & A265;
  assign \new_[72588]_  = \new_[72587]_  & \new_[72584]_ ;
  assign \new_[72591]_  = ~A299 & A298;
  assign \new_[72594]_  = A301 & A300;
  assign \new_[72595]_  = \new_[72594]_  & \new_[72591]_ ;
  assign \new_[72596]_  = \new_[72595]_  & \new_[72588]_ ;
  assign \new_[72600]_  = ~A167 & ~A169;
  assign \new_[72601]_  = A170 & \new_[72600]_ ;
  assign \new_[72604]_  = ~A200 & A166;
  assign \new_[72607]_  = ~A203 & ~A202;
  assign \new_[72608]_  = \new_[72607]_  & \new_[72604]_ ;
  assign \new_[72609]_  = \new_[72608]_  & \new_[72601]_ ;
  assign \new_[72612]_  = A233 & A232;
  assign \new_[72615]_  = ~A267 & A265;
  assign \new_[72616]_  = \new_[72615]_  & \new_[72612]_ ;
  assign \new_[72619]_  = ~A299 & A298;
  assign \new_[72622]_  = A302 & A300;
  assign \new_[72623]_  = \new_[72622]_  & \new_[72619]_ ;
  assign \new_[72624]_  = \new_[72623]_  & \new_[72616]_ ;
  assign \new_[72628]_  = ~A167 & ~A169;
  assign \new_[72629]_  = A170 & \new_[72628]_ ;
  assign \new_[72632]_  = ~A200 & A166;
  assign \new_[72635]_  = ~A203 & ~A202;
  assign \new_[72636]_  = \new_[72635]_  & \new_[72632]_ ;
  assign \new_[72637]_  = \new_[72636]_  & \new_[72629]_ ;
  assign \new_[72640]_  = A233 & A232;
  assign \new_[72643]_  = A266 & A265;
  assign \new_[72644]_  = \new_[72643]_  & \new_[72640]_ ;
  assign \new_[72647]_  = ~A299 & A298;
  assign \new_[72650]_  = A301 & A300;
  assign \new_[72651]_  = \new_[72650]_  & \new_[72647]_ ;
  assign \new_[72652]_  = \new_[72651]_  & \new_[72644]_ ;
  assign \new_[72656]_  = ~A167 & ~A169;
  assign \new_[72657]_  = A170 & \new_[72656]_ ;
  assign \new_[72660]_  = ~A200 & A166;
  assign \new_[72663]_  = ~A203 & ~A202;
  assign \new_[72664]_  = \new_[72663]_  & \new_[72660]_ ;
  assign \new_[72665]_  = \new_[72664]_  & \new_[72657]_ ;
  assign \new_[72668]_  = A233 & A232;
  assign \new_[72671]_  = A266 & A265;
  assign \new_[72672]_  = \new_[72671]_  & \new_[72668]_ ;
  assign \new_[72675]_  = ~A299 & A298;
  assign \new_[72678]_  = A302 & A300;
  assign \new_[72679]_  = \new_[72678]_  & \new_[72675]_ ;
  assign \new_[72680]_  = \new_[72679]_  & \new_[72672]_ ;
  assign \new_[72684]_  = ~A167 & ~A169;
  assign \new_[72685]_  = A170 & \new_[72684]_ ;
  assign \new_[72688]_  = ~A200 & A166;
  assign \new_[72691]_  = ~A203 & ~A202;
  assign \new_[72692]_  = \new_[72691]_  & \new_[72688]_ ;
  assign \new_[72693]_  = \new_[72692]_  & \new_[72685]_ ;
  assign \new_[72696]_  = A233 & A232;
  assign \new_[72699]_  = ~A266 & ~A265;
  assign \new_[72700]_  = \new_[72699]_  & \new_[72696]_ ;
  assign \new_[72703]_  = ~A299 & A298;
  assign \new_[72706]_  = A301 & A300;
  assign \new_[72707]_  = \new_[72706]_  & \new_[72703]_ ;
  assign \new_[72708]_  = \new_[72707]_  & \new_[72700]_ ;
  assign \new_[72712]_  = ~A167 & ~A169;
  assign \new_[72713]_  = A170 & \new_[72712]_ ;
  assign \new_[72716]_  = ~A200 & A166;
  assign \new_[72719]_  = ~A203 & ~A202;
  assign \new_[72720]_  = \new_[72719]_  & \new_[72716]_ ;
  assign \new_[72721]_  = \new_[72720]_  & \new_[72713]_ ;
  assign \new_[72724]_  = A233 & A232;
  assign \new_[72727]_  = ~A266 & ~A265;
  assign \new_[72728]_  = \new_[72727]_  & \new_[72724]_ ;
  assign \new_[72731]_  = ~A299 & A298;
  assign \new_[72734]_  = A302 & A300;
  assign \new_[72735]_  = \new_[72734]_  & \new_[72731]_ ;
  assign \new_[72736]_  = \new_[72735]_  & \new_[72728]_ ;
  assign \new_[72740]_  = ~A167 & ~A169;
  assign \new_[72741]_  = A170 & \new_[72740]_ ;
  assign \new_[72744]_  = ~A200 & A166;
  assign \new_[72747]_  = ~A203 & ~A202;
  assign \new_[72748]_  = \new_[72747]_  & \new_[72744]_ ;
  assign \new_[72749]_  = \new_[72748]_  & \new_[72741]_ ;
  assign \new_[72752]_  = ~A235 & ~A233;
  assign \new_[72755]_  = ~A266 & ~A236;
  assign \new_[72756]_  = \new_[72755]_  & \new_[72752]_ ;
  assign \new_[72759]_  = ~A269 & ~A268;
  assign \new_[72762]_  = A299 & ~A298;
  assign \new_[72763]_  = \new_[72762]_  & \new_[72759]_ ;
  assign \new_[72764]_  = \new_[72763]_  & \new_[72756]_ ;
  assign \new_[72768]_  = ~A167 & ~A169;
  assign \new_[72769]_  = A170 & \new_[72768]_ ;
  assign \new_[72772]_  = ~A200 & A166;
  assign \new_[72775]_  = ~A203 & ~A202;
  assign \new_[72776]_  = \new_[72775]_  & \new_[72772]_ ;
  assign \new_[72777]_  = \new_[72776]_  & \new_[72769]_ ;
  assign \new_[72780]_  = ~A234 & ~A233;
  assign \new_[72783]_  = A266 & A265;
  assign \new_[72784]_  = \new_[72783]_  & \new_[72780]_ ;
  assign \new_[72787]_  = ~A299 & A298;
  assign \new_[72790]_  = A301 & A300;
  assign \new_[72791]_  = \new_[72790]_  & \new_[72787]_ ;
  assign \new_[72792]_  = \new_[72791]_  & \new_[72784]_ ;
  assign \new_[72796]_  = ~A167 & ~A169;
  assign \new_[72797]_  = A170 & \new_[72796]_ ;
  assign \new_[72800]_  = ~A200 & A166;
  assign \new_[72803]_  = ~A203 & ~A202;
  assign \new_[72804]_  = \new_[72803]_  & \new_[72800]_ ;
  assign \new_[72805]_  = \new_[72804]_  & \new_[72797]_ ;
  assign \new_[72808]_  = ~A234 & ~A233;
  assign \new_[72811]_  = A266 & A265;
  assign \new_[72812]_  = \new_[72811]_  & \new_[72808]_ ;
  assign \new_[72815]_  = ~A299 & A298;
  assign \new_[72818]_  = A302 & A300;
  assign \new_[72819]_  = \new_[72818]_  & \new_[72815]_ ;
  assign \new_[72820]_  = \new_[72819]_  & \new_[72812]_ ;
  assign \new_[72824]_  = ~A167 & ~A169;
  assign \new_[72825]_  = A170 & \new_[72824]_ ;
  assign \new_[72828]_  = ~A200 & A166;
  assign \new_[72831]_  = ~A203 & ~A202;
  assign \new_[72832]_  = \new_[72831]_  & \new_[72828]_ ;
  assign \new_[72833]_  = \new_[72832]_  & \new_[72825]_ ;
  assign \new_[72836]_  = ~A234 & ~A233;
  assign \new_[72839]_  = ~A267 & ~A266;
  assign \new_[72840]_  = \new_[72839]_  & \new_[72836]_ ;
  assign \new_[72843]_  = ~A299 & A298;
  assign \new_[72846]_  = A301 & A300;
  assign \new_[72847]_  = \new_[72846]_  & \new_[72843]_ ;
  assign \new_[72848]_  = \new_[72847]_  & \new_[72840]_ ;
  assign \new_[72852]_  = ~A167 & ~A169;
  assign \new_[72853]_  = A170 & \new_[72852]_ ;
  assign \new_[72856]_  = ~A200 & A166;
  assign \new_[72859]_  = ~A203 & ~A202;
  assign \new_[72860]_  = \new_[72859]_  & \new_[72856]_ ;
  assign \new_[72861]_  = \new_[72860]_  & \new_[72853]_ ;
  assign \new_[72864]_  = ~A234 & ~A233;
  assign \new_[72867]_  = ~A267 & ~A266;
  assign \new_[72868]_  = \new_[72867]_  & \new_[72864]_ ;
  assign \new_[72871]_  = ~A299 & A298;
  assign \new_[72874]_  = A302 & A300;
  assign \new_[72875]_  = \new_[72874]_  & \new_[72871]_ ;
  assign \new_[72876]_  = \new_[72875]_  & \new_[72868]_ ;
  assign \new_[72880]_  = ~A167 & ~A169;
  assign \new_[72881]_  = A170 & \new_[72880]_ ;
  assign \new_[72884]_  = ~A200 & A166;
  assign \new_[72887]_  = ~A203 & ~A202;
  assign \new_[72888]_  = \new_[72887]_  & \new_[72884]_ ;
  assign \new_[72889]_  = \new_[72888]_  & \new_[72881]_ ;
  assign \new_[72892]_  = ~A234 & ~A233;
  assign \new_[72895]_  = ~A266 & ~A265;
  assign \new_[72896]_  = \new_[72895]_  & \new_[72892]_ ;
  assign \new_[72899]_  = ~A299 & A298;
  assign \new_[72902]_  = A301 & A300;
  assign \new_[72903]_  = \new_[72902]_  & \new_[72899]_ ;
  assign \new_[72904]_  = \new_[72903]_  & \new_[72896]_ ;
  assign \new_[72908]_  = ~A167 & ~A169;
  assign \new_[72909]_  = A170 & \new_[72908]_ ;
  assign \new_[72912]_  = ~A200 & A166;
  assign \new_[72915]_  = ~A203 & ~A202;
  assign \new_[72916]_  = \new_[72915]_  & \new_[72912]_ ;
  assign \new_[72917]_  = \new_[72916]_  & \new_[72909]_ ;
  assign \new_[72920]_  = ~A234 & ~A233;
  assign \new_[72923]_  = ~A266 & ~A265;
  assign \new_[72924]_  = \new_[72923]_  & \new_[72920]_ ;
  assign \new_[72927]_  = ~A299 & A298;
  assign \new_[72930]_  = A302 & A300;
  assign \new_[72931]_  = \new_[72930]_  & \new_[72927]_ ;
  assign \new_[72932]_  = \new_[72931]_  & \new_[72924]_ ;
  assign \new_[72936]_  = ~A167 & ~A169;
  assign \new_[72937]_  = A170 & \new_[72936]_ ;
  assign \new_[72940]_  = ~A200 & A166;
  assign \new_[72943]_  = ~A203 & ~A202;
  assign \new_[72944]_  = \new_[72943]_  & \new_[72940]_ ;
  assign \new_[72945]_  = \new_[72944]_  & \new_[72937]_ ;
  assign \new_[72948]_  = ~A233 & A232;
  assign \new_[72951]_  = A235 & A234;
  assign \new_[72952]_  = \new_[72951]_  & \new_[72948]_ ;
  assign \new_[72955]_  = ~A266 & A265;
  assign \new_[72958]_  = A268 & A267;
  assign \new_[72959]_  = \new_[72958]_  & \new_[72955]_ ;
  assign \new_[72960]_  = \new_[72959]_  & \new_[72952]_ ;
  assign \new_[72964]_  = ~A167 & ~A169;
  assign \new_[72965]_  = A170 & \new_[72964]_ ;
  assign \new_[72968]_  = ~A200 & A166;
  assign \new_[72971]_  = ~A203 & ~A202;
  assign \new_[72972]_  = \new_[72971]_  & \new_[72968]_ ;
  assign \new_[72973]_  = \new_[72972]_  & \new_[72965]_ ;
  assign \new_[72976]_  = ~A233 & A232;
  assign \new_[72979]_  = A235 & A234;
  assign \new_[72980]_  = \new_[72979]_  & \new_[72976]_ ;
  assign \new_[72983]_  = ~A266 & A265;
  assign \new_[72986]_  = A269 & A267;
  assign \new_[72987]_  = \new_[72986]_  & \new_[72983]_ ;
  assign \new_[72988]_  = \new_[72987]_  & \new_[72980]_ ;
  assign \new_[72992]_  = ~A167 & ~A169;
  assign \new_[72993]_  = A170 & \new_[72992]_ ;
  assign \new_[72996]_  = ~A200 & A166;
  assign \new_[72999]_  = ~A203 & ~A202;
  assign \new_[73000]_  = \new_[72999]_  & \new_[72996]_ ;
  assign \new_[73001]_  = \new_[73000]_  & \new_[72993]_ ;
  assign \new_[73004]_  = ~A233 & A232;
  assign \new_[73007]_  = A236 & A234;
  assign \new_[73008]_  = \new_[73007]_  & \new_[73004]_ ;
  assign \new_[73011]_  = ~A266 & A265;
  assign \new_[73014]_  = A268 & A267;
  assign \new_[73015]_  = \new_[73014]_  & \new_[73011]_ ;
  assign \new_[73016]_  = \new_[73015]_  & \new_[73008]_ ;
  assign \new_[73020]_  = ~A167 & ~A169;
  assign \new_[73021]_  = A170 & \new_[73020]_ ;
  assign \new_[73024]_  = ~A200 & A166;
  assign \new_[73027]_  = ~A203 & ~A202;
  assign \new_[73028]_  = \new_[73027]_  & \new_[73024]_ ;
  assign \new_[73029]_  = \new_[73028]_  & \new_[73021]_ ;
  assign \new_[73032]_  = ~A233 & A232;
  assign \new_[73035]_  = A236 & A234;
  assign \new_[73036]_  = \new_[73035]_  & \new_[73032]_ ;
  assign \new_[73039]_  = ~A266 & A265;
  assign \new_[73042]_  = A269 & A267;
  assign \new_[73043]_  = \new_[73042]_  & \new_[73039]_ ;
  assign \new_[73044]_  = \new_[73043]_  & \new_[73036]_ ;
  assign \new_[73048]_  = ~A167 & ~A169;
  assign \new_[73049]_  = A170 & \new_[73048]_ ;
  assign \new_[73052]_  = ~A200 & A166;
  assign \new_[73055]_  = ~A203 & ~A202;
  assign \new_[73056]_  = \new_[73055]_  & \new_[73052]_ ;
  assign \new_[73057]_  = \new_[73056]_  & \new_[73049]_ ;
  assign \new_[73060]_  = ~A233 & ~A232;
  assign \new_[73063]_  = A266 & A265;
  assign \new_[73064]_  = \new_[73063]_  & \new_[73060]_ ;
  assign \new_[73067]_  = ~A299 & A298;
  assign \new_[73070]_  = A301 & A300;
  assign \new_[73071]_  = \new_[73070]_  & \new_[73067]_ ;
  assign \new_[73072]_  = \new_[73071]_  & \new_[73064]_ ;
  assign \new_[73076]_  = ~A167 & ~A169;
  assign \new_[73077]_  = A170 & \new_[73076]_ ;
  assign \new_[73080]_  = ~A200 & A166;
  assign \new_[73083]_  = ~A203 & ~A202;
  assign \new_[73084]_  = \new_[73083]_  & \new_[73080]_ ;
  assign \new_[73085]_  = \new_[73084]_  & \new_[73077]_ ;
  assign \new_[73088]_  = ~A233 & ~A232;
  assign \new_[73091]_  = A266 & A265;
  assign \new_[73092]_  = \new_[73091]_  & \new_[73088]_ ;
  assign \new_[73095]_  = ~A299 & A298;
  assign \new_[73098]_  = A302 & A300;
  assign \new_[73099]_  = \new_[73098]_  & \new_[73095]_ ;
  assign \new_[73100]_  = \new_[73099]_  & \new_[73092]_ ;
  assign \new_[73104]_  = ~A167 & ~A169;
  assign \new_[73105]_  = A170 & \new_[73104]_ ;
  assign \new_[73108]_  = ~A200 & A166;
  assign \new_[73111]_  = ~A203 & ~A202;
  assign \new_[73112]_  = \new_[73111]_  & \new_[73108]_ ;
  assign \new_[73113]_  = \new_[73112]_  & \new_[73105]_ ;
  assign \new_[73116]_  = ~A233 & ~A232;
  assign \new_[73119]_  = ~A267 & ~A266;
  assign \new_[73120]_  = \new_[73119]_  & \new_[73116]_ ;
  assign \new_[73123]_  = ~A299 & A298;
  assign \new_[73126]_  = A301 & A300;
  assign \new_[73127]_  = \new_[73126]_  & \new_[73123]_ ;
  assign \new_[73128]_  = \new_[73127]_  & \new_[73120]_ ;
  assign \new_[73132]_  = ~A167 & ~A169;
  assign \new_[73133]_  = A170 & \new_[73132]_ ;
  assign \new_[73136]_  = ~A200 & A166;
  assign \new_[73139]_  = ~A203 & ~A202;
  assign \new_[73140]_  = \new_[73139]_  & \new_[73136]_ ;
  assign \new_[73141]_  = \new_[73140]_  & \new_[73133]_ ;
  assign \new_[73144]_  = ~A233 & ~A232;
  assign \new_[73147]_  = ~A267 & ~A266;
  assign \new_[73148]_  = \new_[73147]_  & \new_[73144]_ ;
  assign \new_[73151]_  = ~A299 & A298;
  assign \new_[73154]_  = A302 & A300;
  assign \new_[73155]_  = \new_[73154]_  & \new_[73151]_ ;
  assign \new_[73156]_  = \new_[73155]_  & \new_[73148]_ ;
  assign \new_[73160]_  = ~A167 & ~A169;
  assign \new_[73161]_  = A170 & \new_[73160]_ ;
  assign \new_[73164]_  = ~A200 & A166;
  assign \new_[73167]_  = ~A203 & ~A202;
  assign \new_[73168]_  = \new_[73167]_  & \new_[73164]_ ;
  assign \new_[73169]_  = \new_[73168]_  & \new_[73161]_ ;
  assign \new_[73172]_  = ~A233 & ~A232;
  assign \new_[73175]_  = ~A266 & ~A265;
  assign \new_[73176]_  = \new_[73175]_  & \new_[73172]_ ;
  assign \new_[73179]_  = ~A299 & A298;
  assign \new_[73182]_  = A301 & A300;
  assign \new_[73183]_  = \new_[73182]_  & \new_[73179]_ ;
  assign \new_[73184]_  = \new_[73183]_  & \new_[73176]_ ;
  assign \new_[73188]_  = ~A167 & ~A169;
  assign \new_[73189]_  = A170 & \new_[73188]_ ;
  assign \new_[73192]_  = ~A200 & A166;
  assign \new_[73195]_  = ~A203 & ~A202;
  assign \new_[73196]_  = \new_[73195]_  & \new_[73192]_ ;
  assign \new_[73197]_  = \new_[73196]_  & \new_[73189]_ ;
  assign \new_[73200]_  = ~A233 & ~A232;
  assign \new_[73203]_  = ~A266 & ~A265;
  assign \new_[73204]_  = \new_[73203]_  & \new_[73200]_ ;
  assign \new_[73207]_  = ~A299 & A298;
  assign \new_[73210]_  = A302 & A300;
  assign \new_[73211]_  = \new_[73210]_  & \new_[73207]_ ;
  assign \new_[73212]_  = \new_[73211]_  & \new_[73204]_ ;
  assign \new_[73216]_  = ~A167 & ~A169;
  assign \new_[73217]_  = A170 & \new_[73216]_ ;
  assign \new_[73220]_  = ~A200 & A166;
  assign \new_[73223]_  = A232 & ~A201;
  assign \new_[73224]_  = \new_[73223]_  & \new_[73220]_ ;
  assign \new_[73225]_  = \new_[73224]_  & \new_[73217]_ ;
  assign \new_[73228]_  = A265 & A233;
  assign \new_[73231]_  = ~A269 & ~A268;
  assign \new_[73232]_  = \new_[73231]_  & \new_[73228]_ ;
  assign \new_[73235]_  = ~A299 & A298;
  assign \new_[73238]_  = A301 & A300;
  assign \new_[73239]_  = \new_[73238]_  & \new_[73235]_ ;
  assign \new_[73240]_  = \new_[73239]_  & \new_[73232]_ ;
  assign \new_[73244]_  = ~A167 & ~A169;
  assign \new_[73245]_  = A170 & \new_[73244]_ ;
  assign \new_[73248]_  = ~A200 & A166;
  assign \new_[73251]_  = A232 & ~A201;
  assign \new_[73252]_  = \new_[73251]_  & \new_[73248]_ ;
  assign \new_[73253]_  = \new_[73252]_  & \new_[73245]_ ;
  assign \new_[73256]_  = A265 & A233;
  assign \new_[73259]_  = ~A269 & ~A268;
  assign \new_[73260]_  = \new_[73259]_  & \new_[73256]_ ;
  assign \new_[73263]_  = ~A299 & A298;
  assign \new_[73266]_  = A302 & A300;
  assign \new_[73267]_  = \new_[73266]_  & \new_[73263]_ ;
  assign \new_[73268]_  = \new_[73267]_  & \new_[73260]_ ;
  assign \new_[73272]_  = ~A167 & ~A169;
  assign \new_[73273]_  = A170 & \new_[73272]_ ;
  assign \new_[73276]_  = ~A200 & A166;
  assign \new_[73279]_  = ~A233 & ~A201;
  assign \new_[73280]_  = \new_[73279]_  & \new_[73276]_ ;
  assign \new_[73281]_  = \new_[73280]_  & \new_[73273]_ ;
  assign \new_[73284]_  = ~A236 & ~A235;
  assign \new_[73287]_  = A266 & A265;
  assign \new_[73288]_  = \new_[73287]_  & \new_[73284]_ ;
  assign \new_[73291]_  = ~A299 & A298;
  assign \new_[73294]_  = A301 & A300;
  assign \new_[73295]_  = \new_[73294]_  & \new_[73291]_ ;
  assign \new_[73296]_  = \new_[73295]_  & \new_[73288]_ ;
  assign \new_[73300]_  = ~A167 & ~A169;
  assign \new_[73301]_  = A170 & \new_[73300]_ ;
  assign \new_[73304]_  = ~A200 & A166;
  assign \new_[73307]_  = ~A233 & ~A201;
  assign \new_[73308]_  = \new_[73307]_  & \new_[73304]_ ;
  assign \new_[73309]_  = \new_[73308]_  & \new_[73301]_ ;
  assign \new_[73312]_  = ~A236 & ~A235;
  assign \new_[73315]_  = A266 & A265;
  assign \new_[73316]_  = \new_[73315]_  & \new_[73312]_ ;
  assign \new_[73319]_  = ~A299 & A298;
  assign \new_[73322]_  = A302 & A300;
  assign \new_[73323]_  = \new_[73322]_  & \new_[73319]_ ;
  assign \new_[73324]_  = \new_[73323]_  & \new_[73316]_ ;
  assign \new_[73328]_  = ~A167 & ~A169;
  assign \new_[73329]_  = A170 & \new_[73328]_ ;
  assign \new_[73332]_  = ~A200 & A166;
  assign \new_[73335]_  = ~A233 & ~A201;
  assign \new_[73336]_  = \new_[73335]_  & \new_[73332]_ ;
  assign \new_[73337]_  = \new_[73336]_  & \new_[73329]_ ;
  assign \new_[73340]_  = ~A236 & ~A235;
  assign \new_[73343]_  = ~A267 & ~A266;
  assign \new_[73344]_  = \new_[73343]_  & \new_[73340]_ ;
  assign \new_[73347]_  = ~A299 & A298;
  assign \new_[73350]_  = A301 & A300;
  assign \new_[73351]_  = \new_[73350]_  & \new_[73347]_ ;
  assign \new_[73352]_  = \new_[73351]_  & \new_[73344]_ ;
  assign \new_[73356]_  = ~A167 & ~A169;
  assign \new_[73357]_  = A170 & \new_[73356]_ ;
  assign \new_[73360]_  = ~A200 & A166;
  assign \new_[73363]_  = ~A233 & ~A201;
  assign \new_[73364]_  = \new_[73363]_  & \new_[73360]_ ;
  assign \new_[73365]_  = \new_[73364]_  & \new_[73357]_ ;
  assign \new_[73368]_  = ~A236 & ~A235;
  assign \new_[73371]_  = ~A267 & ~A266;
  assign \new_[73372]_  = \new_[73371]_  & \new_[73368]_ ;
  assign \new_[73375]_  = ~A299 & A298;
  assign \new_[73378]_  = A302 & A300;
  assign \new_[73379]_  = \new_[73378]_  & \new_[73375]_ ;
  assign \new_[73380]_  = \new_[73379]_  & \new_[73372]_ ;
  assign \new_[73384]_  = ~A167 & ~A169;
  assign \new_[73385]_  = A170 & \new_[73384]_ ;
  assign \new_[73388]_  = ~A200 & A166;
  assign \new_[73391]_  = ~A233 & ~A201;
  assign \new_[73392]_  = \new_[73391]_  & \new_[73388]_ ;
  assign \new_[73393]_  = \new_[73392]_  & \new_[73385]_ ;
  assign \new_[73396]_  = ~A236 & ~A235;
  assign \new_[73399]_  = ~A266 & ~A265;
  assign \new_[73400]_  = \new_[73399]_  & \new_[73396]_ ;
  assign \new_[73403]_  = ~A299 & A298;
  assign \new_[73406]_  = A301 & A300;
  assign \new_[73407]_  = \new_[73406]_  & \new_[73403]_ ;
  assign \new_[73408]_  = \new_[73407]_  & \new_[73400]_ ;
  assign \new_[73412]_  = ~A167 & ~A169;
  assign \new_[73413]_  = A170 & \new_[73412]_ ;
  assign \new_[73416]_  = ~A200 & A166;
  assign \new_[73419]_  = ~A233 & ~A201;
  assign \new_[73420]_  = \new_[73419]_  & \new_[73416]_ ;
  assign \new_[73421]_  = \new_[73420]_  & \new_[73413]_ ;
  assign \new_[73424]_  = ~A236 & ~A235;
  assign \new_[73427]_  = ~A266 & ~A265;
  assign \new_[73428]_  = \new_[73427]_  & \new_[73424]_ ;
  assign \new_[73431]_  = ~A299 & A298;
  assign \new_[73434]_  = A302 & A300;
  assign \new_[73435]_  = \new_[73434]_  & \new_[73431]_ ;
  assign \new_[73436]_  = \new_[73435]_  & \new_[73428]_ ;
  assign \new_[73440]_  = ~A167 & ~A169;
  assign \new_[73441]_  = A170 & \new_[73440]_ ;
  assign \new_[73444]_  = ~A200 & A166;
  assign \new_[73447]_  = ~A233 & ~A201;
  assign \new_[73448]_  = \new_[73447]_  & \new_[73444]_ ;
  assign \new_[73449]_  = \new_[73448]_  & \new_[73441]_ ;
  assign \new_[73452]_  = ~A266 & ~A234;
  assign \new_[73455]_  = ~A269 & ~A268;
  assign \new_[73456]_  = \new_[73455]_  & \new_[73452]_ ;
  assign \new_[73459]_  = ~A299 & A298;
  assign \new_[73462]_  = A301 & A300;
  assign \new_[73463]_  = \new_[73462]_  & \new_[73459]_ ;
  assign \new_[73464]_  = \new_[73463]_  & \new_[73456]_ ;
  assign \new_[73468]_  = ~A167 & ~A169;
  assign \new_[73469]_  = A170 & \new_[73468]_ ;
  assign \new_[73472]_  = ~A200 & A166;
  assign \new_[73475]_  = ~A233 & ~A201;
  assign \new_[73476]_  = \new_[73475]_  & \new_[73472]_ ;
  assign \new_[73477]_  = \new_[73476]_  & \new_[73469]_ ;
  assign \new_[73480]_  = ~A266 & ~A234;
  assign \new_[73483]_  = ~A269 & ~A268;
  assign \new_[73484]_  = \new_[73483]_  & \new_[73480]_ ;
  assign \new_[73487]_  = ~A299 & A298;
  assign \new_[73490]_  = A302 & A300;
  assign \new_[73491]_  = \new_[73490]_  & \new_[73487]_ ;
  assign \new_[73492]_  = \new_[73491]_  & \new_[73484]_ ;
  assign \new_[73496]_  = ~A167 & ~A169;
  assign \new_[73497]_  = A170 & \new_[73496]_ ;
  assign \new_[73500]_  = ~A200 & A166;
  assign \new_[73503]_  = ~A232 & ~A201;
  assign \new_[73504]_  = \new_[73503]_  & \new_[73500]_ ;
  assign \new_[73505]_  = \new_[73504]_  & \new_[73497]_ ;
  assign \new_[73508]_  = ~A266 & ~A233;
  assign \new_[73511]_  = ~A269 & ~A268;
  assign \new_[73512]_  = \new_[73511]_  & \new_[73508]_ ;
  assign \new_[73515]_  = ~A299 & A298;
  assign \new_[73518]_  = A301 & A300;
  assign \new_[73519]_  = \new_[73518]_  & \new_[73515]_ ;
  assign \new_[73520]_  = \new_[73519]_  & \new_[73512]_ ;
  assign \new_[73524]_  = ~A167 & ~A169;
  assign \new_[73525]_  = A170 & \new_[73524]_ ;
  assign \new_[73528]_  = ~A200 & A166;
  assign \new_[73531]_  = ~A232 & ~A201;
  assign \new_[73532]_  = \new_[73531]_  & \new_[73528]_ ;
  assign \new_[73533]_  = \new_[73532]_  & \new_[73525]_ ;
  assign \new_[73536]_  = ~A266 & ~A233;
  assign \new_[73539]_  = ~A269 & ~A268;
  assign \new_[73540]_  = \new_[73539]_  & \new_[73536]_ ;
  assign \new_[73543]_  = ~A299 & A298;
  assign \new_[73546]_  = A302 & A300;
  assign \new_[73547]_  = \new_[73546]_  & \new_[73543]_ ;
  assign \new_[73548]_  = \new_[73547]_  & \new_[73540]_ ;
  assign \new_[73552]_  = ~A167 & ~A169;
  assign \new_[73553]_  = A170 & \new_[73552]_ ;
  assign \new_[73556]_  = ~A199 & A166;
  assign \new_[73559]_  = A232 & ~A200;
  assign \new_[73560]_  = \new_[73559]_  & \new_[73556]_ ;
  assign \new_[73561]_  = \new_[73560]_  & \new_[73553]_ ;
  assign \new_[73564]_  = A265 & A233;
  assign \new_[73567]_  = ~A269 & ~A268;
  assign \new_[73568]_  = \new_[73567]_  & \new_[73564]_ ;
  assign \new_[73571]_  = ~A299 & A298;
  assign \new_[73574]_  = A301 & A300;
  assign \new_[73575]_  = \new_[73574]_  & \new_[73571]_ ;
  assign \new_[73576]_  = \new_[73575]_  & \new_[73568]_ ;
  assign \new_[73580]_  = ~A167 & ~A169;
  assign \new_[73581]_  = A170 & \new_[73580]_ ;
  assign \new_[73584]_  = ~A199 & A166;
  assign \new_[73587]_  = A232 & ~A200;
  assign \new_[73588]_  = \new_[73587]_  & \new_[73584]_ ;
  assign \new_[73589]_  = \new_[73588]_  & \new_[73581]_ ;
  assign \new_[73592]_  = A265 & A233;
  assign \new_[73595]_  = ~A269 & ~A268;
  assign \new_[73596]_  = \new_[73595]_  & \new_[73592]_ ;
  assign \new_[73599]_  = ~A299 & A298;
  assign \new_[73602]_  = A302 & A300;
  assign \new_[73603]_  = \new_[73602]_  & \new_[73599]_ ;
  assign \new_[73604]_  = \new_[73603]_  & \new_[73596]_ ;
  assign \new_[73608]_  = ~A167 & ~A169;
  assign \new_[73609]_  = A170 & \new_[73608]_ ;
  assign \new_[73612]_  = ~A199 & A166;
  assign \new_[73615]_  = ~A233 & ~A200;
  assign \new_[73616]_  = \new_[73615]_  & \new_[73612]_ ;
  assign \new_[73617]_  = \new_[73616]_  & \new_[73609]_ ;
  assign \new_[73620]_  = ~A236 & ~A235;
  assign \new_[73623]_  = A266 & A265;
  assign \new_[73624]_  = \new_[73623]_  & \new_[73620]_ ;
  assign \new_[73627]_  = ~A299 & A298;
  assign \new_[73630]_  = A301 & A300;
  assign \new_[73631]_  = \new_[73630]_  & \new_[73627]_ ;
  assign \new_[73632]_  = \new_[73631]_  & \new_[73624]_ ;
  assign \new_[73636]_  = ~A167 & ~A169;
  assign \new_[73637]_  = A170 & \new_[73636]_ ;
  assign \new_[73640]_  = ~A199 & A166;
  assign \new_[73643]_  = ~A233 & ~A200;
  assign \new_[73644]_  = \new_[73643]_  & \new_[73640]_ ;
  assign \new_[73645]_  = \new_[73644]_  & \new_[73637]_ ;
  assign \new_[73648]_  = ~A236 & ~A235;
  assign \new_[73651]_  = A266 & A265;
  assign \new_[73652]_  = \new_[73651]_  & \new_[73648]_ ;
  assign \new_[73655]_  = ~A299 & A298;
  assign \new_[73658]_  = A302 & A300;
  assign \new_[73659]_  = \new_[73658]_  & \new_[73655]_ ;
  assign \new_[73660]_  = \new_[73659]_  & \new_[73652]_ ;
  assign \new_[73664]_  = ~A167 & ~A169;
  assign \new_[73665]_  = A170 & \new_[73664]_ ;
  assign \new_[73668]_  = ~A199 & A166;
  assign \new_[73671]_  = ~A233 & ~A200;
  assign \new_[73672]_  = \new_[73671]_  & \new_[73668]_ ;
  assign \new_[73673]_  = \new_[73672]_  & \new_[73665]_ ;
  assign \new_[73676]_  = ~A236 & ~A235;
  assign \new_[73679]_  = ~A267 & ~A266;
  assign \new_[73680]_  = \new_[73679]_  & \new_[73676]_ ;
  assign \new_[73683]_  = ~A299 & A298;
  assign \new_[73686]_  = A301 & A300;
  assign \new_[73687]_  = \new_[73686]_  & \new_[73683]_ ;
  assign \new_[73688]_  = \new_[73687]_  & \new_[73680]_ ;
  assign \new_[73692]_  = ~A167 & ~A169;
  assign \new_[73693]_  = A170 & \new_[73692]_ ;
  assign \new_[73696]_  = ~A199 & A166;
  assign \new_[73699]_  = ~A233 & ~A200;
  assign \new_[73700]_  = \new_[73699]_  & \new_[73696]_ ;
  assign \new_[73701]_  = \new_[73700]_  & \new_[73693]_ ;
  assign \new_[73704]_  = ~A236 & ~A235;
  assign \new_[73707]_  = ~A267 & ~A266;
  assign \new_[73708]_  = \new_[73707]_  & \new_[73704]_ ;
  assign \new_[73711]_  = ~A299 & A298;
  assign \new_[73714]_  = A302 & A300;
  assign \new_[73715]_  = \new_[73714]_  & \new_[73711]_ ;
  assign \new_[73716]_  = \new_[73715]_  & \new_[73708]_ ;
  assign \new_[73720]_  = ~A167 & ~A169;
  assign \new_[73721]_  = A170 & \new_[73720]_ ;
  assign \new_[73724]_  = ~A199 & A166;
  assign \new_[73727]_  = ~A233 & ~A200;
  assign \new_[73728]_  = \new_[73727]_  & \new_[73724]_ ;
  assign \new_[73729]_  = \new_[73728]_  & \new_[73721]_ ;
  assign \new_[73732]_  = ~A236 & ~A235;
  assign \new_[73735]_  = ~A266 & ~A265;
  assign \new_[73736]_  = \new_[73735]_  & \new_[73732]_ ;
  assign \new_[73739]_  = ~A299 & A298;
  assign \new_[73742]_  = A301 & A300;
  assign \new_[73743]_  = \new_[73742]_  & \new_[73739]_ ;
  assign \new_[73744]_  = \new_[73743]_  & \new_[73736]_ ;
  assign \new_[73748]_  = ~A167 & ~A169;
  assign \new_[73749]_  = A170 & \new_[73748]_ ;
  assign \new_[73752]_  = ~A199 & A166;
  assign \new_[73755]_  = ~A233 & ~A200;
  assign \new_[73756]_  = \new_[73755]_  & \new_[73752]_ ;
  assign \new_[73757]_  = \new_[73756]_  & \new_[73749]_ ;
  assign \new_[73760]_  = ~A236 & ~A235;
  assign \new_[73763]_  = ~A266 & ~A265;
  assign \new_[73764]_  = \new_[73763]_  & \new_[73760]_ ;
  assign \new_[73767]_  = ~A299 & A298;
  assign \new_[73770]_  = A302 & A300;
  assign \new_[73771]_  = \new_[73770]_  & \new_[73767]_ ;
  assign \new_[73772]_  = \new_[73771]_  & \new_[73764]_ ;
  assign \new_[73776]_  = ~A167 & ~A169;
  assign \new_[73777]_  = A170 & \new_[73776]_ ;
  assign \new_[73780]_  = ~A199 & A166;
  assign \new_[73783]_  = ~A233 & ~A200;
  assign \new_[73784]_  = \new_[73783]_  & \new_[73780]_ ;
  assign \new_[73785]_  = \new_[73784]_  & \new_[73777]_ ;
  assign \new_[73788]_  = ~A266 & ~A234;
  assign \new_[73791]_  = ~A269 & ~A268;
  assign \new_[73792]_  = \new_[73791]_  & \new_[73788]_ ;
  assign \new_[73795]_  = ~A299 & A298;
  assign \new_[73798]_  = A301 & A300;
  assign \new_[73799]_  = \new_[73798]_  & \new_[73795]_ ;
  assign \new_[73800]_  = \new_[73799]_  & \new_[73792]_ ;
  assign \new_[73804]_  = ~A167 & ~A169;
  assign \new_[73805]_  = A170 & \new_[73804]_ ;
  assign \new_[73808]_  = ~A199 & A166;
  assign \new_[73811]_  = ~A233 & ~A200;
  assign \new_[73812]_  = \new_[73811]_  & \new_[73808]_ ;
  assign \new_[73813]_  = \new_[73812]_  & \new_[73805]_ ;
  assign \new_[73816]_  = ~A266 & ~A234;
  assign \new_[73819]_  = ~A269 & ~A268;
  assign \new_[73820]_  = \new_[73819]_  & \new_[73816]_ ;
  assign \new_[73823]_  = ~A299 & A298;
  assign \new_[73826]_  = A302 & A300;
  assign \new_[73827]_  = \new_[73826]_  & \new_[73823]_ ;
  assign \new_[73828]_  = \new_[73827]_  & \new_[73820]_ ;
  assign \new_[73832]_  = ~A167 & ~A169;
  assign \new_[73833]_  = A170 & \new_[73832]_ ;
  assign \new_[73836]_  = ~A199 & A166;
  assign \new_[73839]_  = ~A232 & ~A200;
  assign \new_[73840]_  = \new_[73839]_  & \new_[73836]_ ;
  assign \new_[73841]_  = \new_[73840]_  & \new_[73833]_ ;
  assign \new_[73844]_  = ~A266 & ~A233;
  assign \new_[73847]_  = ~A269 & ~A268;
  assign \new_[73848]_  = \new_[73847]_  & \new_[73844]_ ;
  assign \new_[73851]_  = ~A299 & A298;
  assign \new_[73854]_  = A301 & A300;
  assign \new_[73855]_  = \new_[73854]_  & \new_[73851]_ ;
  assign \new_[73856]_  = \new_[73855]_  & \new_[73848]_ ;
  assign \new_[73860]_  = ~A167 & ~A169;
  assign \new_[73861]_  = A170 & \new_[73860]_ ;
  assign \new_[73864]_  = ~A199 & A166;
  assign \new_[73867]_  = ~A232 & ~A200;
  assign \new_[73868]_  = \new_[73867]_  & \new_[73864]_ ;
  assign \new_[73869]_  = \new_[73868]_  & \new_[73861]_ ;
  assign \new_[73872]_  = ~A266 & ~A233;
  assign \new_[73875]_  = ~A269 & ~A268;
  assign \new_[73876]_  = \new_[73875]_  & \new_[73872]_ ;
  assign \new_[73879]_  = ~A299 & A298;
  assign \new_[73882]_  = A302 & A300;
  assign \new_[73883]_  = \new_[73882]_  & \new_[73879]_ ;
  assign \new_[73884]_  = \new_[73883]_  & \new_[73876]_ ;
  assign \new_[73888]_  = ~A168 & ~A169;
  assign \new_[73889]_  = ~A170 & \new_[73888]_ ;
  assign \new_[73892]_  = ~A200 & A199;
  assign \new_[73895]_  = A202 & A201;
  assign \new_[73896]_  = \new_[73895]_  & \new_[73892]_ ;
  assign \new_[73897]_  = \new_[73896]_  & \new_[73889]_ ;
  assign \new_[73900]_  = A233 & A232;
  assign \new_[73903]_  = ~A267 & A265;
  assign \new_[73904]_  = \new_[73903]_  & \new_[73900]_ ;
  assign \new_[73907]_  = ~A299 & A298;
  assign \new_[73910]_  = A301 & A300;
  assign \new_[73911]_  = \new_[73910]_  & \new_[73907]_ ;
  assign \new_[73912]_  = \new_[73911]_  & \new_[73904]_ ;
  assign \new_[73916]_  = ~A168 & ~A169;
  assign \new_[73917]_  = ~A170 & \new_[73916]_ ;
  assign \new_[73920]_  = ~A200 & A199;
  assign \new_[73923]_  = A202 & A201;
  assign \new_[73924]_  = \new_[73923]_  & \new_[73920]_ ;
  assign \new_[73925]_  = \new_[73924]_  & \new_[73917]_ ;
  assign \new_[73928]_  = A233 & A232;
  assign \new_[73931]_  = ~A267 & A265;
  assign \new_[73932]_  = \new_[73931]_  & \new_[73928]_ ;
  assign \new_[73935]_  = ~A299 & A298;
  assign \new_[73938]_  = A302 & A300;
  assign \new_[73939]_  = \new_[73938]_  & \new_[73935]_ ;
  assign \new_[73940]_  = \new_[73939]_  & \new_[73932]_ ;
  assign \new_[73944]_  = ~A168 & ~A169;
  assign \new_[73945]_  = ~A170 & \new_[73944]_ ;
  assign \new_[73948]_  = ~A200 & A199;
  assign \new_[73951]_  = A202 & A201;
  assign \new_[73952]_  = \new_[73951]_  & \new_[73948]_ ;
  assign \new_[73953]_  = \new_[73952]_  & \new_[73945]_ ;
  assign \new_[73956]_  = A233 & A232;
  assign \new_[73959]_  = A266 & A265;
  assign \new_[73960]_  = \new_[73959]_  & \new_[73956]_ ;
  assign \new_[73963]_  = ~A299 & A298;
  assign \new_[73966]_  = A301 & A300;
  assign \new_[73967]_  = \new_[73966]_  & \new_[73963]_ ;
  assign \new_[73968]_  = \new_[73967]_  & \new_[73960]_ ;
  assign \new_[73972]_  = ~A168 & ~A169;
  assign \new_[73973]_  = ~A170 & \new_[73972]_ ;
  assign \new_[73976]_  = ~A200 & A199;
  assign \new_[73979]_  = A202 & A201;
  assign \new_[73980]_  = \new_[73979]_  & \new_[73976]_ ;
  assign \new_[73981]_  = \new_[73980]_  & \new_[73973]_ ;
  assign \new_[73984]_  = A233 & A232;
  assign \new_[73987]_  = A266 & A265;
  assign \new_[73988]_  = \new_[73987]_  & \new_[73984]_ ;
  assign \new_[73991]_  = ~A299 & A298;
  assign \new_[73994]_  = A302 & A300;
  assign \new_[73995]_  = \new_[73994]_  & \new_[73991]_ ;
  assign \new_[73996]_  = \new_[73995]_  & \new_[73988]_ ;
  assign \new_[74000]_  = ~A168 & ~A169;
  assign \new_[74001]_  = ~A170 & \new_[74000]_ ;
  assign \new_[74004]_  = ~A200 & A199;
  assign \new_[74007]_  = A202 & A201;
  assign \new_[74008]_  = \new_[74007]_  & \new_[74004]_ ;
  assign \new_[74009]_  = \new_[74008]_  & \new_[74001]_ ;
  assign \new_[74012]_  = A233 & A232;
  assign \new_[74015]_  = ~A266 & ~A265;
  assign \new_[74016]_  = \new_[74015]_  & \new_[74012]_ ;
  assign \new_[74019]_  = ~A299 & A298;
  assign \new_[74022]_  = A301 & A300;
  assign \new_[74023]_  = \new_[74022]_  & \new_[74019]_ ;
  assign \new_[74024]_  = \new_[74023]_  & \new_[74016]_ ;
  assign \new_[74028]_  = ~A168 & ~A169;
  assign \new_[74029]_  = ~A170 & \new_[74028]_ ;
  assign \new_[74032]_  = ~A200 & A199;
  assign \new_[74035]_  = A202 & A201;
  assign \new_[74036]_  = \new_[74035]_  & \new_[74032]_ ;
  assign \new_[74037]_  = \new_[74036]_  & \new_[74029]_ ;
  assign \new_[74040]_  = A233 & A232;
  assign \new_[74043]_  = ~A266 & ~A265;
  assign \new_[74044]_  = \new_[74043]_  & \new_[74040]_ ;
  assign \new_[74047]_  = ~A299 & A298;
  assign \new_[74050]_  = A302 & A300;
  assign \new_[74051]_  = \new_[74050]_  & \new_[74047]_ ;
  assign \new_[74052]_  = \new_[74051]_  & \new_[74044]_ ;
  assign \new_[74056]_  = ~A168 & ~A169;
  assign \new_[74057]_  = ~A170 & \new_[74056]_ ;
  assign \new_[74060]_  = ~A200 & A199;
  assign \new_[74063]_  = A202 & A201;
  assign \new_[74064]_  = \new_[74063]_  & \new_[74060]_ ;
  assign \new_[74065]_  = \new_[74064]_  & \new_[74057]_ ;
  assign \new_[74068]_  = ~A235 & ~A233;
  assign \new_[74071]_  = ~A266 & ~A236;
  assign \new_[74072]_  = \new_[74071]_  & \new_[74068]_ ;
  assign \new_[74075]_  = ~A269 & ~A268;
  assign \new_[74078]_  = A299 & ~A298;
  assign \new_[74079]_  = \new_[74078]_  & \new_[74075]_ ;
  assign \new_[74080]_  = \new_[74079]_  & \new_[74072]_ ;
  assign \new_[74084]_  = ~A168 & ~A169;
  assign \new_[74085]_  = ~A170 & \new_[74084]_ ;
  assign \new_[74088]_  = ~A200 & A199;
  assign \new_[74091]_  = A202 & A201;
  assign \new_[74092]_  = \new_[74091]_  & \new_[74088]_ ;
  assign \new_[74093]_  = \new_[74092]_  & \new_[74085]_ ;
  assign \new_[74096]_  = ~A234 & ~A233;
  assign \new_[74099]_  = A266 & A265;
  assign \new_[74100]_  = \new_[74099]_  & \new_[74096]_ ;
  assign \new_[74103]_  = ~A299 & A298;
  assign \new_[74106]_  = A301 & A300;
  assign \new_[74107]_  = \new_[74106]_  & \new_[74103]_ ;
  assign \new_[74108]_  = \new_[74107]_  & \new_[74100]_ ;
  assign \new_[74112]_  = ~A168 & ~A169;
  assign \new_[74113]_  = ~A170 & \new_[74112]_ ;
  assign \new_[74116]_  = ~A200 & A199;
  assign \new_[74119]_  = A202 & A201;
  assign \new_[74120]_  = \new_[74119]_  & \new_[74116]_ ;
  assign \new_[74121]_  = \new_[74120]_  & \new_[74113]_ ;
  assign \new_[74124]_  = ~A234 & ~A233;
  assign \new_[74127]_  = A266 & A265;
  assign \new_[74128]_  = \new_[74127]_  & \new_[74124]_ ;
  assign \new_[74131]_  = ~A299 & A298;
  assign \new_[74134]_  = A302 & A300;
  assign \new_[74135]_  = \new_[74134]_  & \new_[74131]_ ;
  assign \new_[74136]_  = \new_[74135]_  & \new_[74128]_ ;
  assign \new_[74140]_  = ~A168 & ~A169;
  assign \new_[74141]_  = ~A170 & \new_[74140]_ ;
  assign \new_[74144]_  = ~A200 & A199;
  assign \new_[74147]_  = A202 & A201;
  assign \new_[74148]_  = \new_[74147]_  & \new_[74144]_ ;
  assign \new_[74149]_  = \new_[74148]_  & \new_[74141]_ ;
  assign \new_[74152]_  = ~A234 & ~A233;
  assign \new_[74155]_  = ~A267 & ~A266;
  assign \new_[74156]_  = \new_[74155]_  & \new_[74152]_ ;
  assign \new_[74159]_  = ~A299 & A298;
  assign \new_[74162]_  = A301 & A300;
  assign \new_[74163]_  = \new_[74162]_  & \new_[74159]_ ;
  assign \new_[74164]_  = \new_[74163]_  & \new_[74156]_ ;
  assign \new_[74168]_  = ~A168 & ~A169;
  assign \new_[74169]_  = ~A170 & \new_[74168]_ ;
  assign \new_[74172]_  = ~A200 & A199;
  assign \new_[74175]_  = A202 & A201;
  assign \new_[74176]_  = \new_[74175]_  & \new_[74172]_ ;
  assign \new_[74177]_  = \new_[74176]_  & \new_[74169]_ ;
  assign \new_[74180]_  = ~A234 & ~A233;
  assign \new_[74183]_  = ~A267 & ~A266;
  assign \new_[74184]_  = \new_[74183]_  & \new_[74180]_ ;
  assign \new_[74187]_  = ~A299 & A298;
  assign \new_[74190]_  = A302 & A300;
  assign \new_[74191]_  = \new_[74190]_  & \new_[74187]_ ;
  assign \new_[74192]_  = \new_[74191]_  & \new_[74184]_ ;
  assign \new_[74196]_  = ~A168 & ~A169;
  assign \new_[74197]_  = ~A170 & \new_[74196]_ ;
  assign \new_[74200]_  = ~A200 & A199;
  assign \new_[74203]_  = A202 & A201;
  assign \new_[74204]_  = \new_[74203]_  & \new_[74200]_ ;
  assign \new_[74205]_  = \new_[74204]_  & \new_[74197]_ ;
  assign \new_[74208]_  = ~A234 & ~A233;
  assign \new_[74211]_  = ~A266 & ~A265;
  assign \new_[74212]_  = \new_[74211]_  & \new_[74208]_ ;
  assign \new_[74215]_  = ~A299 & A298;
  assign \new_[74218]_  = A301 & A300;
  assign \new_[74219]_  = \new_[74218]_  & \new_[74215]_ ;
  assign \new_[74220]_  = \new_[74219]_  & \new_[74212]_ ;
  assign \new_[74224]_  = ~A168 & ~A169;
  assign \new_[74225]_  = ~A170 & \new_[74224]_ ;
  assign \new_[74228]_  = ~A200 & A199;
  assign \new_[74231]_  = A202 & A201;
  assign \new_[74232]_  = \new_[74231]_  & \new_[74228]_ ;
  assign \new_[74233]_  = \new_[74232]_  & \new_[74225]_ ;
  assign \new_[74236]_  = ~A234 & ~A233;
  assign \new_[74239]_  = ~A266 & ~A265;
  assign \new_[74240]_  = \new_[74239]_  & \new_[74236]_ ;
  assign \new_[74243]_  = ~A299 & A298;
  assign \new_[74246]_  = A302 & A300;
  assign \new_[74247]_  = \new_[74246]_  & \new_[74243]_ ;
  assign \new_[74248]_  = \new_[74247]_  & \new_[74240]_ ;
  assign \new_[74252]_  = ~A168 & ~A169;
  assign \new_[74253]_  = ~A170 & \new_[74252]_ ;
  assign \new_[74256]_  = ~A200 & A199;
  assign \new_[74259]_  = A202 & A201;
  assign \new_[74260]_  = \new_[74259]_  & \new_[74256]_ ;
  assign \new_[74261]_  = \new_[74260]_  & \new_[74253]_ ;
  assign \new_[74264]_  = ~A233 & A232;
  assign \new_[74267]_  = A235 & A234;
  assign \new_[74268]_  = \new_[74267]_  & \new_[74264]_ ;
  assign \new_[74271]_  = ~A266 & A265;
  assign \new_[74274]_  = A268 & A267;
  assign \new_[74275]_  = \new_[74274]_  & \new_[74271]_ ;
  assign \new_[74276]_  = \new_[74275]_  & \new_[74268]_ ;
  assign \new_[74280]_  = ~A168 & ~A169;
  assign \new_[74281]_  = ~A170 & \new_[74280]_ ;
  assign \new_[74284]_  = ~A200 & A199;
  assign \new_[74287]_  = A202 & A201;
  assign \new_[74288]_  = \new_[74287]_  & \new_[74284]_ ;
  assign \new_[74289]_  = \new_[74288]_  & \new_[74281]_ ;
  assign \new_[74292]_  = ~A233 & A232;
  assign \new_[74295]_  = A235 & A234;
  assign \new_[74296]_  = \new_[74295]_  & \new_[74292]_ ;
  assign \new_[74299]_  = ~A266 & A265;
  assign \new_[74302]_  = A269 & A267;
  assign \new_[74303]_  = \new_[74302]_  & \new_[74299]_ ;
  assign \new_[74304]_  = \new_[74303]_  & \new_[74296]_ ;
  assign \new_[74308]_  = ~A168 & ~A169;
  assign \new_[74309]_  = ~A170 & \new_[74308]_ ;
  assign \new_[74312]_  = ~A200 & A199;
  assign \new_[74315]_  = A202 & A201;
  assign \new_[74316]_  = \new_[74315]_  & \new_[74312]_ ;
  assign \new_[74317]_  = \new_[74316]_  & \new_[74309]_ ;
  assign \new_[74320]_  = ~A233 & A232;
  assign \new_[74323]_  = A236 & A234;
  assign \new_[74324]_  = \new_[74323]_  & \new_[74320]_ ;
  assign \new_[74327]_  = ~A266 & A265;
  assign \new_[74330]_  = A268 & A267;
  assign \new_[74331]_  = \new_[74330]_  & \new_[74327]_ ;
  assign \new_[74332]_  = \new_[74331]_  & \new_[74324]_ ;
  assign \new_[74336]_  = ~A168 & ~A169;
  assign \new_[74337]_  = ~A170 & \new_[74336]_ ;
  assign \new_[74340]_  = ~A200 & A199;
  assign \new_[74343]_  = A202 & A201;
  assign \new_[74344]_  = \new_[74343]_  & \new_[74340]_ ;
  assign \new_[74345]_  = \new_[74344]_  & \new_[74337]_ ;
  assign \new_[74348]_  = ~A233 & A232;
  assign \new_[74351]_  = A236 & A234;
  assign \new_[74352]_  = \new_[74351]_  & \new_[74348]_ ;
  assign \new_[74355]_  = ~A266 & A265;
  assign \new_[74358]_  = A269 & A267;
  assign \new_[74359]_  = \new_[74358]_  & \new_[74355]_ ;
  assign \new_[74360]_  = \new_[74359]_  & \new_[74352]_ ;
  assign \new_[74364]_  = ~A168 & ~A169;
  assign \new_[74365]_  = ~A170 & \new_[74364]_ ;
  assign \new_[74368]_  = ~A200 & A199;
  assign \new_[74371]_  = A202 & A201;
  assign \new_[74372]_  = \new_[74371]_  & \new_[74368]_ ;
  assign \new_[74373]_  = \new_[74372]_  & \new_[74365]_ ;
  assign \new_[74376]_  = ~A233 & ~A232;
  assign \new_[74379]_  = A266 & A265;
  assign \new_[74380]_  = \new_[74379]_  & \new_[74376]_ ;
  assign \new_[74383]_  = ~A299 & A298;
  assign \new_[74386]_  = A301 & A300;
  assign \new_[74387]_  = \new_[74386]_  & \new_[74383]_ ;
  assign \new_[74388]_  = \new_[74387]_  & \new_[74380]_ ;
  assign \new_[74392]_  = ~A168 & ~A169;
  assign \new_[74393]_  = ~A170 & \new_[74392]_ ;
  assign \new_[74396]_  = ~A200 & A199;
  assign \new_[74399]_  = A202 & A201;
  assign \new_[74400]_  = \new_[74399]_  & \new_[74396]_ ;
  assign \new_[74401]_  = \new_[74400]_  & \new_[74393]_ ;
  assign \new_[74404]_  = ~A233 & ~A232;
  assign \new_[74407]_  = A266 & A265;
  assign \new_[74408]_  = \new_[74407]_  & \new_[74404]_ ;
  assign \new_[74411]_  = ~A299 & A298;
  assign \new_[74414]_  = A302 & A300;
  assign \new_[74415]_  = \new_[74414]_  & \new_[74411]_ ;
  assign \new_[74416]_  = \new_[74415]_  & \new_[74408]_ ;
  assign \new_[74420]_  = ~A168 & ~A169;
  assign \new_[74421]_  = ~A170 & \new_[74420]_ ;
  assign \new_[74424]_  = ~A200 & A199;
  assign \new_[74427]_  = A202 & A201;
  assign \new_[74428]_  = \new_[74427]_  & \new_[74424]_ ;
  assign \new_[74429]_  = \new_[74428]_  & \new_[74421]_ ;
  assign \new_[74432]_  = ~A233 & ~A232;
  assign \new_[74435]_  = ~A267 & ~A266;
  assign \new_[74436]_  = \new_[74435]_  & \new_[74432]_ ;
  assign \new_[74439]_  = ~A299 & A298;
  assign \new_[74442]_  = A301 & A300;
  assign \new_[74443]_  = \new_[74442]_  & \new_[74439]_ ;
  assign \new_[74444]_  = \new_[74443]_  & \new_[74436]_ ;
  assign \new_[74448]_  = ~A168 & ~A169;
  assign \new_[74449]_  = ~A170 & \new_[74448]_ ;
  assign \new_[74452]_  = ~A200 & A199;
  assign \new_[74455]_  = A202 & A201;
  assign \new_[74456]_  = \new_[74455]_  & \new_[74452]_ ;
  assign \new_[74457]_  = \new_[74456]_  & \new_[74449]_ ;
  assign \new_[74460]_  = ~A233 & ~A232;
  assign \new_[74463]_  = ~A267 & ~A266;
  assign \new_[74464]_  = \new_[74463]_  & \new_[74460]_ ;
  assign \new_[74467]_  = ~A299 & A298;
  assign \new_[74470]_  = A302 & A300;
  assign \new_[74471]_  = \new_[74470]_  & \new_[74467]_ ;
  assign \new_[74472]_  = \new_[74471]_  & \new_[74464]_ ;
  assign \new_[74476]_  = ~A168 & ~A169;
  assign \new_[74477]_  = ~A170 & \new_[74476]_ ;
  assign \new_[74480]_  = ~A200 & A199;
  assign \new_[74483]_  = A202 & A201;
  assign \new_[74484]_  = \new_[74483]_  & \new_[74480]_ ;
  assign \new_[74485]_  = \new_[74484]_  & \new_[74477]_ ;
  assign \new_[74488]_  = ~A233 & ~A232;
  assign \new_[74491]_  = ~A266 & ~A265;
  assign \new_[74492]_  = \new_[74491]_  & \new_[74488]_ ;
  assign \new_[74495]_  = ~A299 & A298;
  assign \new_[74498]_  = A301 & A300;
  assign \new_[74499]_  = \new_[74498]_  & \new_[74495]_ ;
  assign \new_[74500]_  = \new_[74499]_  & \new_[74492]_ ;
  assign \new_[74504]_  = ~A168 & ~A169;
  assign \new_[74505]_  = ~A170 & \new_[74504]_ ;
  assign \new_[74508]_  = ~A200 & A199;
  assign \new_[74511]_  = A202 & A201;
  assign \new_[74512]_  = \new_[74511]_  & \new_[74508]_ ;
  assign \new_[74513]_  = \new_[74512]_  & \new_[74505]_ ;
  assign \new_[74516]_  = ~A233 & ~A232;
  assign \new_[74519]_  = ~A266 & ~A265;
  assign \new_[74520]_  = \new_[74519]_  & \new_[74516]_ ;
  assign \new_[74523]_  = ~A299 & A298;
  assign \new_[74526]_  = A302 & A300;
  assign \new_[74527]_  = \new_[74526]_  & \new_[74523]_ ;
  assign \new_[74528]_  = \new_[74527]_  & \new_[74520]_ ;
  assign \new_[74532]_  = ~A168 & ~A169;
  assign \new_[74533]_  = ~A170 & \new_[74532]_ ;
  assign \new_[74536]_  = ~A200 & A199;
  assign \new_[74539]_  = A203 & A201;
  assign \new_[74540]_  = \new_[74539]_  & \new_[74536]_ ;
  assign \new_[74541]_  = \new_[74540]_  & \new_[74533]_ ;
  assign \new_[74544]_  = A233 & A232;
  assign \new_[74547]_  = ~A267 & A265;
  assign \new_[74548]_  = \new_[74547]_  & \new_[74544]_ ;
  assign \new_[74551]_  = ~A299 & A298;
  assign \new_[74554]_  = A301 & A300;
  assign \new_[74555]_  = \new_[74554]_  & \new_[74551]_ ;
  assign \new_[74556]_  = \new_[74555]_  & \new_[74548]_ ;
  assign \new_[74560]_  = ~A168 & ~A169;
  assign \new_[74561]_  = ~A170 & \new_[74560]_ ;
  assign \new_[74564]_  = ~A200 & A199;
  assign \new_[74567]_  = A203 & A201;
  assign \new_[74568]_  = \new_[74567]_  & \new_[74564]_ ;
  assign \new_[74569]_  = \new_[74568]_  & \new_[74561]_ ;
  assign \new_[74572]_  = A233 & A232;
  assign \new_[74575]_  = ~A267 & A265;
  assign \new_[74576]_  = \new_[74575]_  & \new_[74572]_ ;
  assign \new_[74579]_  = ~A299 & A298;
  assign \new_[74582]_  = A302 & A300;
  assign \new_[74583]_  = \new_[74582]_  & \new_[74579]_ ;
  assign \new_[74584]_  = \new_[74583]_  & \new_[74576]_ ;
  assign \new_[74588]_  = ~A168 & ~A169;
  assign \new_[74589]_  = ~A170 & \new_[74588]_ ;
  assign \new_[74592]_  = ~A200 & A199;
  assign \new_[74595]_  = A203 & A201;
  assign \new_[74596]_  = \new_[74595]_  & \new_[74592]_ ;
  assign \new_[74597]_  = \new_[74596]_  & \new_[74589]_ ;
  assign \new_[74600]_  = A233 & A232;
  assign \new_[74603]_  = A266 & A265;
  assign \new_[74604]_  = \new_[74603]_  & \new_[74600]_ ;
  assign \new_[74607]_  = ~A299 & A298;
  assign \new_[74610]_  = A301 & A300;
  assign \new_[74611]_  = \new_[74610]_  & \new_[74607]_ ;
  assign \new_[74612]_  = \new_[74611]_  & \new_[74604]_ ;
  assign \new_[74616]_  = ~A168 & ~A169;
  assign \new_[74617]_  = ~A170 & \new_[74616]_ ;
  assign \new_[74620]_  = ~A200 & A199;
  assign \new_[74623]_  = A203 & A201;
  assign \new_[74624]_  = \new_[74623]_  & \new_[74620]_ ;
  assign \new_[74625]_  = \new_[74624]_  & \new_[74617]_ ;
  assign \new_[74628]_  = A233 & A232;
  assign \new_[74631]_  = A266 & A265;
  assign \new_[74632]_  = \new_[74631]_  & \new_[74628]_ ;
  assign \new_[74635]_  = ~A299 & A298;
  assign \new_[74638]_  = A302 & A300;
  assign \new_[74639]_  = \new_[74638]_  & \new_[74635]_ ;
  assign \new_[74640]_  = \new_[74639]_  & \new_[74632]_ ;
  assign \new_[74644]_  = ~A168 & ~A169;
  assign \new_[74645]_  = ~A170 & \new_[74644]_ ;
  assign \new_[74648]_  = ~A200 & A199;
  assign \new_[74651]_  = A203 & A201;
  assign \new_[74652]_  = \new_[74651]_  & \new_[74648]_ ;
  assign \new_[74653]_  = \new_[74652]_  & \new_[74645]_ ;
  assign \new_[74656]_  = A233 & A232;
  assign \new_[74659]_  = ~A266 & ~A265;
  assign \new_[74660]_  = \new_[74659]_  & \new_[74656]_ ;
  assign \new_[74663]_  = ~A299 & A298;
  assign \new_[74666]_  = A301 & A300;
  assign \new_[74667]_  = \new_[74666]_  & \new_[74663]_ ;
  assign \new_[74668]_  = \new_[74667]_  & \new_[74660]_ ;
  assign \new_[74672]_  = ~A168 & ~A169;
  assign \new_[74673]_  = ~A170 & \new_[74672]_ ;
  assign \new_[74676]_  = ~A200 & A199;
  assign \new_[74679]_  = A203 & A201;
  assign \new_[74680]_  = \new_[74679]_  & \new_[74676]_ ;
  assign \new_[74681]_  = \new_[74680]_  & \new_[74673]_ ;
  assign \new_[74684]_  = A233 & A232;
  assign \new_[74687]_  = ~A266 & ~A265;
  assign \new_[74688]_  = \new_[74687]_  & \new_[74684]_ ;
  assign \new_[74691]_  = ~A299 & A298;
  assign \new_[74694]_  = A302 & A300;
  assign \new_[74695]_  = \new_[74694]_  & \new_[74691]_ ;
  assign \new_[74696]_  = \new_[74695]_  & \new_[74688]_ ;
  assign \new_[74700]_  = ~A168 & ~A169;
  assign \new_[74701]_  = ~A170 & \new_[74700]_ ;
  assign \new_[74704]_  = ~A200 & A199;
  assign \new_[74707]_  = A203 & A201;
  assign \new_[74708]_  = \new_[74707]_  & \new_[74704]_ ;
  assign \new_[74709]_  = \new_[74708]_  & \new_[74701]_ ;
  assign \new_[74712]_  = ~A235 & ~A233;
  assign \new_[74715]_  = ~A266 & ~A236;
  assign \new_[74716]_  = \new_[74715]_  & \new_[74712]_ ;
  assign \new_[74719]_  = ~A269 & ~A268;
  assign \new_[74722]_  = A299 & ~A298;
  assign \new_[74723]_  = \new_[74722]_  & \new_[74719]_ ;
  assign \new_[74724]_  = \new_[74723]_  & \new_[74716]_ ;
  assign \new_[74728]_  = ~A168 & ~A169;
  assign \new_[74729]_  = ~A170 & \new_[74728]_ ;
  assign \new_[74732]_  = ~A200 & A199;
  assign \new_[74735]_  = A203 & A201;
  assign \new_[74736]_  = \new_[74735]_  & \new_[74732]_ ;
  assign \new_[74737]_  = \new_[74736]_  & \new_[74729]_ ;
  assign \new_[74740]_  = ~A234 & ~A233;
  assign \new_[74743]_  = A266 & A265;
  assign \new_[74744]_  = \new_[74743]_  & \new_[74740]_ ;
  assign \new_[74747]_  = ~A299 & A298;
  assign \new_[74750]_  = A301 & A300;
  assign \new_[74751]_  = \new_[74750]_  & \new_[74747]_ ;
  assign \new_[74752]_  = \new_[74751]_  & \new_[74744]_ ;
  assign \new_[74756]_  = ~A168 & ~A169;
  assign \new_[74757]_  = ~A170 & \new_[74756]_ ;
  assign \new_[74760]_  = ~A200 & A199;
  assign \new_[74763]_  = A203 & A201;
  assign \new_[74764]_  = \new_[74763]_  & \new_[74760]_ ;
  assign \new_[74765]_  = \new_[74764]_  & \new_[74757]_ ;
  assign \new_[74768]_  = ~A234 & ~A233;
  assign \new_[74771]_  = A266 & A265;
  assign \new_[74772]_  = \new_[74771]_  & \new_[74768]_ ;
  assign \new_[74775]_  = ~A299 & A298;
  assign \new_[74778]_  = A302 & A300;
  assign \new_[74779]_  = \new_[74778]_  & \new_[74775]_ ;
  assign \new_[74780]_  = \new_[74779]_  & \new_[74772]_ ;
  assign \new_[74784]_  = ~A168 & ~A169;
  assign \new_[74785]_  = ~A170 & \new_[74784]_ ;
  assign \new_[74788]_  = ~A200 & A199;
  assign \new_[74791]_  = A203 & A201;
  assign \new_[74792]_  = \new_[74791]_  & \new_[74788]_ ;
  assign \new_[74793]_  = \new_[74792]_  & \new_[74785]_ ;
  assign \new_[74796]_  = ~A234 & ~A233;
  assign \new_[74799]_  = ~A267 & ~A266;
  assign \new_[74800]_  = \new_[74799]_  & \new_[74796]_ ;
  assign \new_[74803]_  = ~A299 & A298;
  assign \new_[74806]_  = A301 & A300;
  assign \new_[74807]_  = \new_[74806]_  & \new_[74803]_ ;
  assign \new_[74808]_  = \new_[74807]_  & \new_[74800]_ ;
  assign \new_[74812]_  = ~A168 & ~A169;
  assign \new_[74813]_  = ~A170 & \new_[74812]_ ;
  assign \new_[74816]_  = ~A200 & A199;
  assign \new_[74819]_  = A203 & A201;
  assign \new_[74820]_  = \new_[74819]_  & \new_[74816]_ ;
  assign \new_[74821]_  = \new_[74820]_  & \new_[74813]_ ;
  assign \new_[74824]_  = ~A234 & ~A233;
  assign \new_[74827]_  = ~A267 & ~A266;
  assign \new_[74828]_  = \new_[74827]_  & \new_[74824]_ ;
  assign \new_[74831]_  = ~A299 & A298;
  assign \new_[74834]_  = A302 & A300;
  assign \new_[74835]_  = \new_[74834]_  & \new_[74831]_ ;
  assign \new_[74836]_  = \new_[74835]_  & \new_[74828]_ ;
  assign \new_[74840]_  = ~A168 & ~A169;
  assign \new_[74841]_  = ~A170 & \new_[74840]_ ;
  assign \new_[74844]_  = ~A200 & A199;
  assign \new_[74847]_  = A203 & A201;
  assign \new_[74848]_  = \new_[74847]_  & \new_[74844]_ ;
  assign \new_[74849]_  = \new_[74848]_  & \new_[74841]_ ;
  assign \new_[74852]_  = ~A234 & ~A233;
  assign \new_[74855]_  = ~A266 & ~A265;
  assign \new_[74856]_  = \new_[74855]_  & \new_[74852]_ ;
  assign \new_[74859]_  = ~A299 & A298;
  assign \new_[74862]_  = A301 & A300;
  assign \new_[74863]_  = \new_[74862]_  & \new_[74859]_ ;
  assign \new_[74864]_  = \new_[74863]_  & \new_[74856]_ ;
  assign \new_[74868]_  = ~A168 & ~A169;
  assign \new_[74869]_  = ~A170 & \new_[74868]_ ;
  assign \new_[74872]_  = ~A200 & A199;
  assign \new_[74875]_  = A203 & A201;
  assign \new_[74876]_  = \new_[74875]_  & \new_[74872]_ ;
  assign \new_[74877]_  = \new_[74876]_  & \new_[74869]_ ;
  assign \new_[74880]_  = ~A234 & ~A233;
  assign \new_[74883]_  = ~A266 & ~A265;
  assign \new_[74884]_  = \new_[74883]_  & \new_[74880]_ ;
  assign \new_[74887]_  = ~A299 & A298;
  assign \new_[74890]_  = A302 & A300;
  assign \new_[74891]_  = \new_[74890]_  & \new_[74887]_ ;
  assign \new_[74892]_  = \new_[74891]_  & \new_[74884]_ ;
  assign \new_[74896]_  = ~A168 & ~A169;
  assign \new_[74897]_  = ~A170 & \new_[74896]_ ;
  assign \new_[74900]_  = ~A200 & A199;
  assign \new_[74903]_  = A203 & A201;
  assign \new_[74904]_  = \new_[74903]_  & \new_[74900]_ ;
  assign \new_[74905]_  = \new_[74904]_  & \new_[74897]_ ;
  assign \new_[74908]_  = ~A233 & A232;
  assign \new_[74911]_  = A235 & A234;
  assign \new_[74912]_  = \new_[74911]_  & \new_[74908]_ ;
  assign \new_[74915]_  = ~A266 & A265;
  assign \new_[74918]_  = A268 & A267;
  assign \new_[74919]_  = \new_[74918]_  & \new_[74915]_ ;
  assign \new_[74920]_  = \new_[74919]_  & \new_[74912]_ ;
  assign \new_[74924]_  = ~A168 & ~A169;
  assign \new_[74925]_  = ~A170 & \new_[74924]_ ;
  assign \new_[74928]_  = ~A200 & A199;
  assign \new_[74931]_  = A203 & A201;
  assign \new_[74932]_  = \new_[74931]_  & \new_[74928]_ ;
  assign \new_[74933]_  = \new_[74932]_  & \new_[74925]_ ;
  assign \new_[74936]_  = ~A233 & A232;
  assign \new_[74939]_  = A235 & A234;
  assign \new_[74940]_  = \new_[74939]_  & \new_[74936]_ ;
  assign \new_[74943]_  = ~A266 & A265;
  assign \new_[74946]_  = A269 & A267;
  assign \new_[74947]_  = \new_[74946]_  & \new_[74943]_ ;
  assign \new_[74948]_  = \new_[74947]_  & \new_[74940]_ ;
  assign \new_[74952]_  = ~A168 & ~A169;
  assign \new_[74953]_  = ~A170 & \new_[74952]_ ;
  assign \new_[74956]_  = ~A200 & A199;
  assign \new_[74959]_  = A203 & A201;
  assign \new_[74960]_  = \new_[74959]_  & \new_[74956]_ ;
  assign \new_[74961]_  = \new_[74960]_  & \new_[74953]_ ;
  assign \new_[74964]_  = ~A233 & A232;
  assign \new_[74967]_  = A236 & A234;
  assign \new_[74968]_  = \new_[74967]_  & \new_[74964]_ ;
  assign \new_[74971]_  = ~A266 & A265;
  assign \new_[74974]_  = A268 & A267;
  assign \new_[74975]_  = \new_[74974]_  & \new_[74971]_ ;
  assign \new_[74976]_  = \new_[74975]_  & \new_[74968]_ ;
  assign \new_[74980]_  = ~A168 & ~A169;
  assign \new_[74981]_  = ~A170 & \new_[74980]_ ;
  assign \new_[74984]_  = ~A200 & A199;
  assign \new_[74987]_  = A203 & A201;
  assign \new_[74988]_  = \new_[74987]_  & \new_[74984]_ ;
  assign \new_[74989]_  = \new_[74988]_  & \new_[74981]_ ;
  assign \new_[74992]_  = ~A233 & A232;
  assign \new_[74995]_  = A236 & A234;
  assign \new_[74996]_  = \new_[74995]_  & \new_[74992]_ ;
  assign \new_[74999]_  = ~A266 & A265;
  assign \new_[75002]_  = A269 & A267;
  assign \new_[75003]_  = \new_[75002]_  & \new_[74999]_ ;
  assign \new_[75004]_  = \new_[75003]_  & \new_[74996]_ ;
  assign \new_[75008]_  = ~A168 & ~A169;
  assign \new_[75009]_  = ~A170 & \new_[75008]_ ;
  assign \new_[75012]_  = ~A200 & A199;
  assign \new_[75015]_  = A203 & A201;
  assign \new_[75016]_  = \new_[75015]_  & \new_[75012]_ ;
  assign \new_[75017]_  = \new_[75016]_  & \new_[75009]_ ;
  assign \new_[75020]_  = ~A233 & ~A232;
  assign \new_[75023]_  = A266 & A265;
  assign \new_[75024]_  = \new_[75023]_  & \new_[75020]_ ;
  assign \new_[75027]_  = ~A299 & A298;
  assign \new_[75030]_  = A301 & A300;
  assign \new_[75031]_  = \new_[75030]_  & \new_[75027]_ ;
  assign \new_[75032]_  = \new_[75031]_  & \new_[75024]_ ;
  assign \new_[75036]_  = ~A168 & ~A169;
  assign \new_[75037]_  = ~A170 & \new_[75036]_ ;
  assign \new_[75040]_  = ~A200 & A199;
  assign \new_[75043]_  = A203 & A201;
  assign \new_[75044]_  = \new_[75043]_  & \new_[75040]_ ;
  assign \new_[75045]_  = \new_[75044]_  & \new_[75037]_ ;
  assign \new_[75048]_  = ~A233 & ~A232;
  assign \new_[75051]_  = A266 & A265;
  assign \new_[75052]_  = \new_[75051]_  & \new_[75048]_ ;
  assign \new_[75055]_  = ~A299 & A298;
  assign \new_[75058]_  = A302 & A300;
  assign \new_[75059]_  = \new_[75058]_  & \new_[75055]_ ;
  assign \new_[75060]_  = \new_[75059]_  & \new_[75052]_ ;
  assign \new_[75064]_  = ~A168 & ~A169;
  assign \new_[75065]_  = ~A170 & \new_[75064]_ ;
  assign \new_[75068]_  = ~A200 & A199;
  assign \new_[75071]_  = A203 & A201;
  assign \new_[75072]_  = \new_[75071]_  & \new_[75068]_ ;
  assign \new_[75073]_  = \new_[75072]_  & \new_[75065]_ ;
  assign \new_[75076]_  = ~A233 & ~A232;
  assign \new_[75079]_  = ~A267 & ~A266;
  assign \new_[75080]_  = \new_[75079]_  & \new_[75076]_ ;
  assign \new_[75083]_  = ~A299 & A298;
  assign \new_[75086]_  = A301 & A300;
  assign \new_[75087]_  = \new_[75086]_  & \new_[75083]_ ;
  assign \new_[75088]_  = \new_[75087]_  & \new_[75080]_ ;
  assign \new_[75092]_  = ~A168 & ~A169;
  assign \new_[75093]_  = ~A170 & \new_[75092]_ ;
  assign \new_[75096]_  = ~A200 & A199;
  assign \new_[75099]_  = A203 & A201;
  assign \new_[75100]_  = \new_[75099]_  & \new_[75096]_ ;
  assign \new_[75101]_  = \new_[75100]_  & \new_[75093]_ ;
  assign \new_[75104]_  = ~A233 & ~A232;
  assign \new_[75107]_  = ~A267 & ~A266;
  assign \new_[75108]_  = \new_[75107]_  & \new_[75104]_ ;
  assign \new_[75111]_  = ~A299 & A298;
  assign \new_[75114]_  = A302 & A300;
  assign \new_[75115]_  = \new_[75114]_  & \new_[75111]_ ;
  assign \new_[75116]_  = \new_[75115]_  & \new_[75108]_ ;
  assign \new_[75120]_  = ~A168 & ~A169;
  assign \new_[75121]_  = ~A170 & \new_[75120]_ ;
  assign \new_[75124]_  = ~A200 & A199;
  assign \new_[75127]_  = A203 & A201;
  assign \new_[75128]_  = \new_[75127]_  & \new_[75124]_ ;
  assign \new_[75129]_  = \new_[75128]_  & \new_[75121]_ ;
  assign \new_[75132]_  = ~A233 & ~A232;
  assign \new_[75135]_  = ~A266 & ~A265;
  assign \new_[75136]_  = \new_[75135]_  & \new_[75132]_ ;
  assign \new_[75139]_  = ~A299 & A298;
  assign \new_[75142]_  = A301 & A300;
  assign \new_[75143]_  = \new_[75142]_  & \new_[75139]_ ;
  assign \new_[75144]_  = \new_[75143]_  & \new_[75136]_ ;
  assign \new_[75148]_  = ~A168 & ~A169;
  assign \new_[75149]_  = ~A170 & \new_[75148]_ ;
  assign \new_[75152]_  = ~A200 & A199;
  assign \new_[75155]_  = A203 & A201;
  assign \new_[75156]_  = \new_[75155]_  & \new_[75152]_ ;
  assign \new_[75157]_  = \new_[75156]_  & \new_[75149]_ ;
  assign \new_[75160]_  = ~A233 & ~A232;
  assign \new_[75163]_  = ~A266 & ~A265;
  assign \new_[75164]_  = \new_[75163]_  & \new_[75160]_ ;
  assign \new_[75167]_  = ~A299 & A298;
  assign \new_[75170]_  = A302 & A300;
  assign \new_[75171]_  = \new_[75170]_  & \new_[75167]_ ;
  assign \new_[75172]_  = \new_[75171]_  & \new_[75164]_ ;
  assign \new_[75175]_  = ~A167 & A170;
  assign \new_[75178]_  = A199 & ~A166;
  assign \new_[75179]_  = \new_[75178]_  & \new_[75175]_ ;
  assign \new_[75182]_  = A201 & ~A200;
  assign \new_[75185]_  = A232 & A202;
  assign \new_[75186]_  = \new_[75185]_  & \new_[75182]_ ;
  assign \new_[75187]_  = \new_[75186]_  & \new_[75179]_ ;
  assign \new_[75190]_  = A265 & A233;
  assign \new_[75193]_  = ~A269 & ~A268;
  assign \new_[75194]_  = \new_[75193]_  & \new_[75190]_ ;
  assign \new_[75197]_  = ~A299 & A298;
  assign \new_[75200]_  = A301 & A300;
  assign \new_[75201]_  = \new_[75200]_  & \new_[75197]_ ;
  assign \new_[75202]_  = \new_[75201]_  & \new_[75194]_ ;
  assign \new_[75205]_  = ~A167 & A170;
  assign \new_[75208]_  = A199 & ~A166;
  assign \new_[75209]_  = \new_[75208]_  & \new_[75205]_ ;
  assign \new_[75212]_  = A201 & ~A200;
  assign \new_[75215]_  = A232 & A202;
  assign \new_[75216]_  = \new_[75215]_  & \new_[75212]_ ;
  assign \new_[75217]_  = \new_[75216]_  & \new_[75209]_ ;
  assign \new_[75220]_  = A265 & A233;
  assign \new_[75223]_  = ~A269 & ~A268;
  assign \new_[75224]_  = \new_[75223]_  & \new_[75220]_ ;
  assign \new_[75227]_  = ~A299 & A298;
  assign \new_[75230]_  = A302 & A300;
  assign \new_[75231]_  = \new_[75230]_  & \new_[75227]_ ;
  assign \new_[75232]_  = \new_[75231]_  & \new_[75224]_ ;
  assign \new_[75235]_  = ~A167 & A170;
  assign \new_[75238]_  = A199 & ~A166;
  assign \new_[75239]_  = \new_[75238]_  & \new_[75235]_ ;
  assign \new_[75242]_  = A201 & ~A200;
  assign \new_[75245]_  = ~A233 & A202;
  assign \new_[75246]_  = \new_[75245]_  & \new_[75242]_ ;
  assign \new_[75247]_  = \new_[75246]_  & \new_[75239]_ ;
  assign \new_[75250]_  = ~A236 & ~A235;
  assign \new_[75253]_  = A266 & A265;
  assign \new_[75254]_  = \new_[75253]_  & \new_[75250]_ ;
  assign \new_[75257]_  = ~A299 & A298;
  assign \new_[75260]_  = A301 & A300;
  assign \new_[75261]_  = \new_[75260]_  & \new_[75257]_ ;
  assign \new_[75262]_  = \new_[75261]_  & \new_[75254]_ ;
  assign \new_[75265]_  = ~A167 & A170;
  assign \new_[75268]_  = A199 & ~A166;
  assign \new_[75269]_  = \new_[75268]_  & \new_[75265]_ ;
  assign \new_[75272]_  = A201 & ~A200;
  assign \new_[75275]_  = ~A233 & A202;
  assign \new_[75276]_  = \new_[75275]_  & \new_[75272]_ ;
  assign \new_[75277]_  = \new_[75276]_  & \new_[75269]_ ;
  assign \new_[75280]_  = ~A236 & ~A235;
  assign \new_[75283]_  = A266 & A265;
  assign \new_[75284]_  = \new_[75283]_  & \new_[75280]_ ;
  assign \new_[75287]_  = ~A299 & A298;
  assign \new_[75290]_  = A302 & A300;
  assign \new_[75291]_  = \new_[75290]_  & \new_[75287]_ ;
  assign \new_[75292]_  = \new_[75291]_  & \new_[75284]_ ;
  assign \new_[75295]_  = ~A167 & A170;
  assign \new_[75298]_  = A199 & ~A166;
  assign \new_[75299]_  = \new_[75298]_  & \new_[75295]_ ;
  assign \new_[75302]_  = A201 & ~A200;
  assign \new_[75305]_  = ~A233 & A202;
  assign \new_[75306]_  = \new_[75305]_  & \new_[75302]_ ;
  assign \new_[75307]_  = \new_[75306]_  & \new_[75299]_ ;
  assign \new_[75310]_  = ~A236 & ~A235;
  assign \new_[75313]_  = ~A267 & ~A266;
  assign \new_[75314]_  = \new_[75313]_  & \new_[75310]_ ;
  assign \new_[75317]_  = ~A299 & A298;
  assign \new_[75320]_  = A301 & A300;
  assign \new_[75321]_  = \new_[75320]_  & \new_[75317]_ ;
  assign \new_[75322]_  = \new_[75321]_  & \new_[75314]_ ;
  assign \new_[75325]_  = ~A167 & A170;
  assign \new_[75328]_  = A199 & ~A166;
  assign \new_[75329]_  = \new_[75328]_  & \new_[75325]_ ;
  assign \new_[75332]_  = A201 & ~A200;
  assign \new_[75335]_  = ~A233 & A202;
  assign \new_[75336]_  = \new_[75335]_  & \new_[75332]_ ;
  assign \new_[75337]_  = \new_[75336]_  & \new_[75329]_ ;
  assign \new_[75340]_  = ~A236 & ~A235;
  assign \new_[75343]_  = ~A267 & ~A266;
  assign \new_[75344]_  = \new_[75343]_  & \new_[75340]_ ;
  assign \new_[75347]_  = ~A299 & A298;
  assign \new_[75350]_  = A302 & A300;
  assign \new_[75351]_  = \new_[75350]_  & \new_[75347]_ ;
  assign \new_[75352]_  = \new_[75351]_  & \new_[75344]_ ;
  assign \new_[75355]_  = ~A167 & A170;
  assign \new_[75358]_  = A199 & ~A166;
  assign \new_[75359]_  = \new_[75358]_  & \new_[75355]_ ;
  assign \new_[75362]_  = A201 & ~A200;
  assign \new_[75365]_  = ~A233 & A202;
  assign \new_[75366]_  = \new_[75365]_  & \new_[75362]_ ;
  assign \new_[75367]_  = \new_[75366]_  & \new_[75359]_ ;
  assign \new_[75370]_  = ~A236 & ~A235;
  assign \new_[75373]_  = ~A266 & ~A265;
  assign \new_[75374]_  = \new_[75373]_  & \new_[75370]_ ;
  assign \new_[75377]_  = ~A299 & A298;
  assign \new_[75380]_  = A301 & A300;
  assign \new_[75381]_  = \new_[75380]_  & \new_[75377]_ ;
  assign \new_[75382]_  = \new_[75381]_  & \new_[75374]_ ;
  assign \new_[75385]_  = ~A167 & A170;
  assign \new_[75388]_  = A199 & ~A166;
  assign \new_[75389]_  = \new_[75388]_  & \new_[75385]_ ;
  assign \new_[75392]_  = A201 & ~A200;
  assign \new_[75395]_  = ~A233 & A202;
  assign \new_[75396]_  = \new_[75395]_  & \new_[75392]_ ;
  assign \new_[75397]_  = \new_[75396]_  & \new_[75389]_ ;
  assign \new_[75400]_  = ~A236 & ~A235;
  assign \new_[75403]_  = ~A266 & ~A265;
  assign \new_[75404]_  = \new_[75403]_  & \new_[75400]_ ;
  assign \new_[75407]_  = ~A299 & A298;
  assign \new_[75410]_  = A302 & A300;
  assign \new_[75411]_  = \new_[75410]_  & \new_[75407]_ ;
  assign \new_[75412]_  = \new_[75411]_  & \new_[75404]_ ;
  assign \new_[75415]_  = ~A167 & A170;
  assign \new_[75418]_  = A199 & ~A166;
  assign \new_[75419]_  = \new_[75418]_  & \new_[75415]_ ;
  assign \new_[75422]_  = A201 & ~A200;
  assign \new_[75425]_  = ~A233 & A202;
  assign \new_[75426]_  = \new_[75425]_  & \new_[75422]_ ;
  assign \new_[75427]_  = \new_[75426]_  & \new_[75419]_ ;
  assign \new_[75430]_  = ~A266 & ~A234;
  assign \new_[75433]_  = ~A269 & ~A268;
  assign \new_[75434]_  = \new_[75433]_  & \new_[75430]_ ;
  assign \new_[75437]_  = ~A299 & A298;
  assign \new_[75440]_  = A301 & A300;
  assign \new_[75441]_  = \new_[75440]_  & \new_[75437]_ ;
  assign \new_[75442]_  = \new_[75441]_  & \new_[75434]_ ;
  assign \new_[75445]_  = ~A167 & A170;
  assign \new_[75448]_  = A199 & ~A166;
  assign \new_[75449]_  = \new_[75448]_  & \new_[75445]_ ;
  assign \new_[75452]_  = A201 & ~A200;
  assign \new_[75455]_  = ~A233 & A202;
  assign \new_[75456]_  = \new_[75455]_  & \new_[75452]_ ;
  assign \new_[75457]_  = \new_[75456]_  & \new_[75449]_ ;
  assign \new_[75460]_  = ~A266 & ~A234;
  assign \new_[75463]_  = ~A269 & ~A268;
  assign \new_[75464]_  = \new_[75463]_  & \new_[75460]_ ;
  assign \new_[75467]_  = ~A299 & A298;
  assign \new_[75470]_  = A302 & A300;
  assign \new_[75471]_  = \new_[75470]_  & \new_[75467]_ ;
  assign \new_[75472]_  = \new_[75471]_  & \new_[75464]_ ;
  assign \new_[75475]_  = ~A167 & A170;
  assign \new_[75478]_  = A199 & ~A166;
  assign \new_[75479]_  = \new_[75478]_  & \new_[75475]_ ;
  assign \new_[75482]_  = A201 & ~A200;
  assign \new_[75485]_  = ~A232 & A202;
  assign \new_[75486]_  = \new_[75485]_  & \new_[75482]_ ;
  assign \new_[75487]_  = \new_[75486]_  & \new_[75479]_ ;
  assign \new_[75490]_  = ~A266 & ~A233;
  assign \new_[75493]_  = ~A269 & ~A268;
  assign \new_[75494]_  = \new_[75493]_  & \new_[75490]_ ;
  assign \new_[75497]_  = ~A299 & A298;
  assign \new_[75500]_  = A301 & A300;
  assign \new_[75501]_  = \new_[75500]_  & \new_[75497]_ ;
  assign \new_[75502]_  = \new_[75501]_  & \new_[75494]_ ;
  assign \new_[75505]_  = ~A167 & A170;
  assign \new_[75508]_  = A199 & ~A166;
  assign \new_[75509]_  = \new_[75508]_  & \new_[75505]_ ;
  assign \new_[75512]_  = A201 & ~A200;
  assign \new_[75515]_  = ~A232 & A202;
  assign \new_[75516]_  = \new_[75515]_  & \new_[75512]_ ;
  assign \new_[75517]_  = \new_[75516]_  & \new_[75509]_ ;
  assign \new_[75520]_  = ~A266 & ~A233;
  assign \new_[75523]_  = ~A269 & ~A268;
  assign \new_[75524]_  = \new_[75523]_  & \new_[75520]_ ;
  assign \new_[75527]_  = ~A299 & A298;
  assign \new_[75530]_  = A302 & A300;
  assign \new_[75531]_  = \new_[75530]_  & \new_[75527]_ ;
  assign \new_[75532]_  = \new_[75531]_  & \new_[75524]_ ;
  assign \new_[75535]_  = ~A167 & A170;
  assign \new_[75538]_  = A199 & ~A166;
  assign \new_[75539]_  = \new_[75538]_  & \new_[75535]_ ;
  assign \new_[75542]_  = A201 & ~A200;
  assign \new_[75545]_  = A232 & A203;
  assign \new_[75546]_  = \new_[75545]_  & \new_[75542]_ ;
  assign \new_[75547]_  = \new_[75546]_  & \new_[75539]_ ;
  assign \new_[75550]_  = A265 & A233;
  assign \new_[75553]_  = ~A269 & ~A268;
  assign \new_[75554]_  = \new_[75553]_  & \new_[75550]_ ;
  assign \new_[75557]_  = ~A299 & A298;
  assign \new_[75560]_  = A301 & A300;
  assign \new_[75561]_  = \new_[75560]_  & \new_[75557]_ ;
  assign \new_[75562]_  = \new_[75561]_  & \new_[75554]_ ;
  assign \new_[75565]_  = ~A167 & A170;
  assign \new_[75568]_  = A199 & ~A166;
  assign \new_[75569]_  = \new_[75568]_  & \new_[75565]_ ;
  assign \new_[75572]_  = A201 & ~A200;
  assign \new_[75575]_  = A232 & A203;
  assign \new_[75576]_  = \new_[75575]_  & \new_[75572]_ ;
  assign \new_[75577]_  = \new_[75576]_  & \new_[75569]_ ;
  assign \new_[75580]_  = A265 & A233;
  assign \new_[75583]_  = ~A269 & ~A268;
  assign \new_[75584]_  = \new_[75583]_  & \new_[75580]_ ;
  assign \new_[75587]_  = ~A299 & A298;
  assign \new_[75590]_  = A302 & A300;
  assign \new_[75591]_  = \new_[75590]_  & \new_[75587]_ ;
  assign \new_[75592]_  = \new_[75591]_  & \new_[75584]_ ;
  assign \new_[75595]_  = ~A167 & A170;
  assign \new_[75598]_  = A199 & ~A166;
  assign \new_[75599]_  = \new_[75598]_  & \new_[75595]_ ;
  assign \new_[75602]_  = A201 & ~A200;
  assign \new_[75605]_  = ~A233 & A203;
  assign \new_[75606]_  = \new_[75605]_  & \new_[75602]_ ;
  assign \new_[75607]_  = \new_[75606]_  & \new_[75599]_ ;
  assign \new_[75610]_  = ~A236 & ~A235;
  assign \new_[75613]_  = A266 & A265;
  assign \new_[75614]_  = \new_[75613]_  & \new_[75610]_ ;
  assign \new_[75617]_  = ~A299 & A298;
  assign \new_[75620]_  = A301 & A300;
  assign \new_[75621]_  = \new_[75620]_  & \new_[75617]_ ;
  assign \new_[75622]_  = \new_[75621]_  & \new_[75614]_ ;
  assign \new_[75625]_  = ~A167 & A170;
  assign \new_[75628]_  = A199 & ~A166;
  assign \new_[75629]_  = \new_[75628]_  & \new_[75625]_ ;
  assign \new_[75632]_  = A201 & ~A200;
  assign \new_[75635]_  = ~A233 & A203;
  assign \new_[75636]_  = \new_[75635]_  & \new_[75632]_ ;
  assign \new_[75637]_  = \new_[75636]_  & \new_[75629]_ ;
  assign \new_[75640]_  = ~A236 & ~A235;
  assign \new_[75643]_  = A266 & A265;
  assign \new_[75644]_  = \new_[75643]_  & \new_[75640]_ ;
  assign \new_[75647]_  = ~A299 & A298;
  assign \new_[75650]_  = A302 & A300;
  assign \new_[75651]_  = \new_[75650]_  & \new_[75647]_ ;
  assign \new_[75652]_  = \new_[75651]_  & \new_[75644]_ ;
  assign \new_[75655]_  = ~A167 & A170;
  assign \new_[75658]_  = A199 & ~A166;
  assign \new_[75659]_  = \new_[75658]_  & \new_[75655]_ ;
  assign \new_[75662]_  = A201 & ~A200;
  assign \new_[75665]_  = ~A233 & A203;
  assign \new_[75666]_  = \new_[75665]_  & \new_[75662]_ ;
  assign \new_[75667]_  = \new_[75666]_  & \new_[75659]_ ;
  assign \new_[75670]_  = ~A236 & ~A235;
  assign \new_[75673]_  = ~A267 & ~A266;
  assign \new_[75674]_  = \new_[75673]_  & \new_[75670]_ ;
  assign \new_[75677]_  = ~A299 & A298;
  assign \new_[75680]_  = A301 & A300;
  assign \new_[75681]_  = \new_[75680]_  & \new_[75677]_ ;
  assign \new_[75682]_  = \new_[75681]_  & \new_[75674]_ ;
  assign \new_[75685]_  = ~A167 & A170;
  assign \new_[75688]_  = A199 & ~A166;
  assign \new_[75689]_  = \new_[75688]_  & \new_[75685]_ ;
  assign \new_[75692]_  = A201 & ~A200;
  assign \new_[75695]_  = ~A233 & A203;
  assign \new_[75696]_  = \new_[75695]_  & \new_[75692]_ ;
  assign \new_[75697]_  = \new_[75696]_  & \new_[75689]_ ;
  assign \new_[75700]_  = ~A236 & ~A235;
  assign \new_[75703]_  = ~A267 & ~A266;
  assign \new_[75704]_  = \new_[75703]_  & \new_[75700]_ ;
  assign \new_[75707]_  = ~A299 & A298;
  assign \new_[75710]_  = A302 & A300;
  assign \new_[75711]_  = \new_[75710]_  & \new_[75707]_ ;
  assign \new_[75712]_  = \new_[75711]_  & \new_[75704]_ ;
  assign \new_[75715]_  = ~A167 & A170;
  assign \new_[75718]_  = A199 & ~A166;
  assign \new_[75719]_  = \new_[75718]_  & \new_[75715]_ ;
  assign \new_[75722]_  = A201 & ~A200;
  assign \new_[75725]_  = ~A233 & A203;
  assign \new_[75726]_  = \new_[75725]_  & \new_[75722]_ ;
  assign \new_[75727]_  = \new_[75726]_  & \new_[75719]_ ;
  assign \new_[75730]_  = ~A236 & ~A235;
  assign \new_[75733]_  = ~A266 & ~A265;
  assign \new_[75734]_  = \new_[75733]_  & \new_[75730]_ ;
  assign \new_[75737]_  = ~A299 & A298;
  assign \new_[75740]_  = A301 & A300;
  assign \new_[75741]_  = \new_[75740]_  & \new_[75737]_ ;
  assign \new_[75742]_  = \new_[75741]_  & \new_[75734]_ ;
  assign \new_[75745]_  = ~A167 & A170;
  assign \new_[75748]_  = A199 & ~A166;
  assign \new_[75749]_  = \new_[75748]_  & \new_[75745]_ ;
  assign \new_[75752]_  = A201 & ~A200;
  assign \new_[75755]_  = ~A233 & A203;
  assign \new_[75756]_  = \new_[75755]_  & \new_[75752]_ ;
  assign \new_[75757]_  = \new_[75756]_  & \new_[75749]_ ;
  assign \new_[75760]_  = ~A236 & ~A235;
  assign \new_[75763]_  = ~A266 & ~A265;
  assign \new_[75764]_  = \new_[75763]_  & \new_[75760]_ ;
  assign \new_[75767]_  = ~A299 & A298;
  assign \new_[75770]_  = A302 & A300;
  assign \new_[75771]_  = \new_[75770]_  & \new_[75767]_ ;
  assign \new_[75772]_  = \new_[75771]_  & \new_[75764]_ ;
  assign \new_[75775]_  = ~A167 & A170;
  assign \new_[75778]_  = A199 & ~A166;
  assign \new_[75779]_  = \new_[75778]_  & \new_[75775]_ ;
  assign \new_[75782]_  = A201 & ~A200;
  assign \new_[75785]_  = ~A233 & A203;
  assign \new_[75786]_  = \new_[75785]_  & \new_[75782]_ ;
  assign \new_[75787]_  = \new_[75786]_  & \new_[75779]_ ;
  assign \new_[75790]_  = ~A266 & ~A234;
  assign \new_[75793]_  = ~A269 & ~A268;
  assign \new_[75794]_  = \new_[75793]_  & \new_[75790]_ ;
  assign \new_[75797]_  = ~A299 & A298;
  assign \new_[75800]_  = A301 & A300;
  assign \new_[75801]_  = \new_[75800]_  & \new_[75797]_ ;
  assign \new_[75802]_  = \new_[75801]_  & \new_[75794]_ ;
  assign \new_[75805]_  = ~A167 & A170;
  assign \new_[75808]_  = A199 & ~A166;
  assign \new_[75809]_  = \new_[75808]_  & \new_[75805]_ ;
  assign \new_[75812]_  = A201 & ~A200;
  assign \new_[75815]_  = ~A233 & A203;
  assign \new_[75816]_  = \new_[75815]_  & \new_[75812]_ ;
  assign \new_[75817]_  = \new_[75816]_  & \new_[75809]_ ;
  assign \new_[75820]_  = ~A266 & ~A234;
  assign \new_[75823]_  = ~A269 & ~A268;
  assign \new_[75824]_  = \new_[75823]_  & \new_[75820]_ ;
  assign \new_[75827]_  = ~A299 & A298;
  assign \new_[75830]_  = A302 & A300;
  assign \new_[75831]_  = \new_[75830]_  & \new_[75827]_ ;
  assign \new_[75832]_  = \new_[75831]_  & \new_[75824]_ ;
  assign \new_[75835]_  = ~A167 & A170;
  assign \new_[75838]_  = A199 & ~A166;
  assign \new_[75839]_  = \new_[75838]_  & \new_[75835]_ ;
  assign \new_[75842]_  = A201 & ~A200;
  assign \new_[75845]_  = ~A232 & A203;
  assign \new_[75846]_  = \new_[75845]_  & \new_[75842]_ ;
  assign \new_[75847]_  = \new_[75846]_  & \new_[75839]_ ;
  assign \new_[75850]_  = ~A266 & ~A233;
  assign \new_[75853]_  = ~A269 & ~A268;
  assign \new_[75854]_  = \new_[75853]_  & \new_[75850]_ ;
  assign \new_[75857]_  = ~A299 & A298;
  assign \new_[75860]_  = A301 & A300;
  assign \new_[75861]_  = \new_[75860]_  & \new_[75857]_ ;
  assign \new_[75862]_  = \new_[75861]_  & \new_[75854]_ ;
  assign \new_[75865]_  = ~A167 & A170;
  assign \new_[75868]_  = A199 & ~A166;
  assign \new_[75869]_  = \new_[75868]_  & \new_[75865]_ ;
  assign \new_[75872]_  = A201 & ~A200;
  assign \new_[75875]_  = ~A232 & A203;
  assign \new_[75876]_  = \new_[75875]_  & \new_[75872]_ ;
  assign \new_[75877]_  = \new_[75876]_  & \new_[75869]_ ;
  assign \new_[75880]_  = ~A266 & ~A233;
  assign \new_[75883]_  = ~A269 & ~A268;
  assign \new_[75884]_  = \new_[75883]_  & \new_[75880]_ ;
  assign \new_[75887]_  = ~A299 & A298;
  assign \new_[75890]_  = A302 & A300;
  assign \new_[75891]_  = \new_[75890]_  & \new_[75887]_ ;
  assign \new_[75892]_  = \new_[75891]_  & \new_[75884]_ ;
  assign \new_[75895]_  = ~A168 & A170;
  assign \new_[75898]_  = A166 & A167;
  assign \new_[75899]_  = \new_[75898]_  & \new_[75895]_ ;
  assign \new_[75902]_  = A200 & ~A199;
  assign \new_[75905]_  = ~A235 & ~A233;
  assign \new_[75906]_  = \new_[75905]_  & \new_[75902]_ ;
  assign \new_[75907]_  = \new_[75906]_  & \new_[75899]_ ;
  assign \new_[75910]_  = ~A266 & ~A236;
  assign \new_[75913]_  = ~A269 & ~A268;
  assign \new_[75914]_  = \new_[75913]_  & \new_[75910]_ ;
  assign \new_[75917]_  = ~A299 & A298;
  assign \new_[75920]_  = A301 & A300;
  assign \new_[75921]_  = \new_[75920]_  & \new_[75917]_ ;
  assign \new_[75922]_  = \new_[75921]_  & \new_[75914]_ ;
  assign \new_[75925]_  = ~A168 & A170;
  assign \new_[75928]_  = A166 & A167;
  assign \new_[75929]_  = \new_[75928]_  & \new_[75925]_ ;
  assign \new_[75932]_  = A200 & ~A199;
  assign \new_[75935]_  = ~A235 & ~A233;
  assign \new_[75936]_  = \new_[75935]_  & \new_[75932]_ ;
  assign \new_[75937]_  = \new_[75936]_  & \new_[75929]_ ;
  assign \new_[75940]_  = ~A266 & ~A236;
  assign \new_[75943]_  = ~A269 & ~A268;
  assign \new_[75944]_  = \new_[75943]_  & \new_[75940]_ ;
  assign \new_[75947]_  = ~A299 & A298;
  assign \new_[75950]_  = A302 & A300;
  assign \new_[75951]_  = \new_[75950]_  & \new_[75947]_ ;
  assign \new_[75952]_  = \new_[75951]_  & \new_[75944]_ ;
  assign \new_[75955]_  = ~A168 & ~A170;
  assign \new_[75958]_  = ~A166 & A167;
  assign \new_[75959]_  = \new_[75958]_  & \new_[75955]_ ;
  assign \new_[75962]_  = A200 & ~A199;
  assign \new_[75965]_  = ~A235 & ~A233;
  assign \new_[75966]_  = \new_[75965]_  & \new_[75962]_ ;
  assign \new_[75967]_  = \new_[75966]_  & \new_[75959]_ ;
  assign \new_[75970]_  = ~A266 & ~A236;
  assign \new_[75973]_  = ~A269 & ~A268;
  assign \new_[75974]_  = \new_[75973]_  & \new_[75970]_ ;
  assign \new_[75977]_  = ~A299 & A298;
  assign \new_[75980]_  = A301 & A300;
  assign \new_[75981]_  = \new_[75980]_  & \new_[75977]_ ;
  assign \new_[75982]_  = \new_[75981]_  & \new_[75974]_ ;
  assign \new_[75985]_  = ~A168 & ~A170;
  assign \new_[75988]_  = ~A166 & A167;
  assign \new_[75989]_  = \new_[75988]_  & \new_[75985]_ ;
  assign \new_[75992]_  = A200 & ~A199;
  assign \new_[75995]_  = ~A235 & ~A233;
  assign \new_[75996]_  = \new_[75995]_  & \new_[75992]_ ;
  assign \new_[75997]_  = \new_[75996]_  & \new_[75989]_ ;
  assign \new_[76000]_  = ~A266 & ~A236;
  assign \new_[76003]_  = ~A269 & ~A268;
  assign \new_[76004]_  = \new_[76003]_  & \new_[76000]_ ;
  assign \new_[76007]_  = ~A299 & A298;
  assign \new_[76010]_  = A302 & A300;
  assign \new_[76011]_  = \new_[76010]_  & \new_[76007]_ ;
  assign \new_[76012]_  = \new_[76011]_  & \new_[76004]_ ;
  assign \new_[76015]_  = ~A168 & ~A170;
  assign \new_[76018]_  = A166 & ~A167;
  assign \new_[76019]_  = \new_[76018]_  & \new_[76015]_ ;
  assign \new_[76022]_  = A200 & ~A199;
  assign \new_[76025]_  = ~A235 & ~A233;
  assign \new_[76026]_  = \new_[76025]_  & \new_[76022]_ ;
  assign \new_[76027]_  = \new_[76026]_  & \new_[76019]_ ;
  assign \new_[76030]_  = ~A266 & ~A236;
  assign \new_[76033]_  = ~A269 & ~A268;
  assign \new_[76034]_  = \new_[76033]_  & \new_[76030]_ ;
  assign \new_[76037]_  = ~A299 & A298;
  assign \new_[76040]_  = A301 & A300;
  assign \new_[76041]_  = \new_[76040]_  & \new_[76037]_ ;
  assign \new_[76042]_  = \new_[76041]_  & \new_[76034]_ ;
  assign \new_[76045]_  = ~A168 & ~A170;
  assign \new_[76048]_  = A166 & ~A167;
  assign \new_[76049]_  = \new_[76048]_  & \new_[76045]_ ;
  assign \new_[76052]_  = A200 & ~A199;
  assign \new_[76055]_  = ~A235 & ~A233;
  assign \new_[76056]_  = \new_[76055]_  & \new_[76052]_ ;
  assign \new_[76057]_  = \new_[76056]_  & \new_[76049]_ ;
  assign \new_[76060]_  = ~A266 & ~A236;
  assign \new_[76063]_  = ~A269 & ~A268;
  assign \new_[76064]_  = \new_[76063]_  & \new_[76060]_ ;
  assign \new_[76067]_  = ~A299 & A298;
  assign \new_[76070]_  = A302 & A300;
  assign \new_[76071]_  = \new_[76070]_  & \new_[76067]_ ;
  assign \new_[76072]_  = \new_[76071]_  & \new_[76064]_ ;
  assign \new_[76075]_  = ~A168 & A169;
  assign \new_[76078]_  = ~A166 & A167;
  assign \new_[76079]_  = \new_[76078]_  & \new_[76075]_ ;
  assign \new_[76082]_  = A200 & ~A199;
  assign \new_[76085]_  = ~A235 & ~A233;
  assign \new_[76086]_  = \new_[76085]_  & \new_[76082]_ ;
  assign \new_[76087]_  = \new_[76086]_  & \new_[76079]_ ;
  assign \new_[76090]_  = ~A266 & ~A236;
  assign \new_[76093]_  = ~A269 & ~A268;
  assign \new_[76094]_  = \new_[76093]_  & \new_[76090]_ ;
  assign \new_[76097]_  = ~A299 & A298;
  assign \new_[76100]_  = A301 & A300;
  assign \new_[76101]_  = \new_[76100]_  & \new_[76097]_ ;
  assign \new_[76102]_  = \new_[76101]_  & \new_[76094]_ ;
  assign \new_[76105]_  = ~A168 & A169;
  assign \new_[76108]_  = ~A166 & A167;
  assign \new_[76109]_  = \new_[76108]_  & \new_[76105]_ ;
  assign \new_[76112]_  = A200 & ~A199;
  assign \new_[76115]_  = ~A235 & ~A233;
  assign \new_[76116]_  = \new_[76115]_  & \new_[76112]_ ;
  assign \new_[76117]_  = \new_[76116]_  & \new_[76109]_ ;
  assign \new_[76120]_  = ~A266 & ~A236;
  assign \new_[76123]_  = ~A269 & ~A268;
  assign \new_[76124]_  = \new_[76123]_  & \new_[76120]_ ;
  assign \new_[76127]_  = ~A299 & A298;
  assign \new_[76130]_  = A302 & A300;
  assign \new_[76131]_  = \new_[76130]_  & \new_[76127]_ ;
  assign \new_[76132]_  = \new_[76131]_  & \new_[76124]_ ;
  assign \new_[76135]_  = ~A168 & A169;
  assign \new_[76138]_  = ~A166 & A167;
  assign \new_[76139]_  = \new_[76138]_  & \new_[76135]_ ;
  assign \new_[76142]_  = ~A200 & A199;
  assign \new_[76145]_  = A202 & A201;
  assign \new_[76146]_  = \new_[76145]_  & \new_[76142]_ ;
  assign \new_[76147]_  = \new_[76146]_  & \new_[76139]_ ;
  assign \new_[76150]_  = A233 & A232;
  assign \new_[76153]_  = ~A267 & A265;
  assign \new_[76154]_  = \new_[76153]_  & \new_[76150]_ ;
  assign \new_[76157]_  = ~A299 & A298;
  assign \new_[76160]_  = A301 & A300;
  assign \new_[76161]_  = \new_[76160]_  & \new_[76157]_ ;
  assign \new_[76162]_  = \new_[76161]_  & \new_[76154]_ ;
  assign \new_[76165]_  = ~A168 & A169;
  assign \new_[76168]_  = ~A166 & A167;
  assign \new_[76169]_  = \new_[76168]_  & \new_[76165]_ ;
  assign \new_[76172]_  = ~A200 & A199;
  assign \new_[76175]_  = A202 & A201;
  assign \new_[76176]_  = \new_[76175]_  & \new_[76172]_ ;
  assign \new_[76177]_  = \new_[76176]_  & \new_[76169]_ ;
  assign \new_[76180]_  = A233 & A232;
  assign \new_[76183]_  = ~A267 & A265;
  assign \new_[76184]_  = \new_[76183]_  & \new_[76180]_ ;
  assign \new_[76187]_  = ~A299 & A298;
  assign \new_[76190]_  = A302 & A300;
  assign \new_[76191]_  = \new_[76190]_  & \new_[76187]_ ;
  assign \new_[76192]_  = \new_[76191]_  & \new_[76184]_ ;
  assign \new_[76195]_  = ~A168 & A169;
  assign \new_[76198]_  = ~A166 & A167;
  assign \new_[76199]_  = \new_[76198]_  & \new_[76195]_ ;
  assign \new_[76202]_  = ~A200 & A199;
  assign \new_[76205]_  = A202 & A201;
  assign \new_[76206]_  = \new_[76205]_  & \new_[76202]_ ;
  assign \new_[76207]_  = \new_[76206]_  & \new_[76199]_ ;
  assign \new_[76210]_  = A233 & A232;
  assign \new_[76213]_  = A266 & A265;
  assign \new_[76214]_  = \new_[76213]_  & \new_[76210]_ ;
  assign \new_[76217]_  = ~A299 & A298;
  assign \new_[76220]_  = A301 & A300;
  assign \new_[76221]_  = \new_[76220]_  & \new_[76217]_ ;
  assign \new_[76222]_  = \new_[76221]_  & \new_[76214]_ ;
  assign \new_[76225]_  = ~A168 & A169;
  assign \new_[76228]_  = ~A166 & A167;
  assign \new_[76229]_  = \new_[76228]_  & \new_[76225]_ ;
  assign \new_[76232]_  = ~A200 & A199;
  assign \new_[76235]_  = A202 & A201;
  assign \new_[76236]_  = \new_[76235]_  & \new_[76232]_ ;
  assign \new_[76237]_  = \new_[76236]_  & \new_[76229]_ ;
  assign \new_[76240]_  = A233 & A232;
  assign \new_[76243]_  = A266 & A265;
  assign \new_[76244]_  = \new_[76243]_  & \new_[76240]_ ;
  assign \new_[76247]_  = ~A299 & A298;
  assign \new_[76250]_  = A302 & A300;
  assign \new_[76251]_  = \new_[76250]_  & \new_[76247]_ ;
  assign \new_[76252]_  = \new_[76251]_  & \new_[76244]_ ;
  assign \new_[76255]_  = ~A168 & A169;
  assign \new_[76258]_  = ~A166 & A167;
  assign \new_[76259]_  = \new_[76258]_  & \new_[76255]_ ;
  assign \new_[76262]_  = ~A200 & A199;
  assign \new_[76265]_  = A202 & A201;
  assign \new_[76266]_  = \new_[76265]_  & \new_[76262]_ ;
  assign \new_[76267]_  = \new_[76266]_  & \new_[76259]_ ;
  assign \new_[76270]_  = A233 & A232;
  assign \new_[76273]_  = ~A266 & ~A265;
  assign \new_[76274]_  = \new_[76273]_  & \new_[76270]_ ;
  assign \new_[76277]_  = ~A299 & A298;
  assign \new_[76280]_  = A301 & A300;
  assign \new_[76281]_  = \new_[76280]_  & \new_[76277]_ ;
  assign \new_[76282]_  = \new_[76281]_  & \new_[76274]_ ;
  assign \new_[76285]_  = ~A168 & A169;
  assign \new_[76288]_  = ~A166 & A167;
  assign \new_[76289]_  = \new_[76288]_  & \new_[76285]_ ;
  assign \new_[76292]_  = ~A200 & A199;
  assign \new_[76295]_  = A202 & A201;
  assign \new_[76296]_  = \new_[76295]_  & \new_[76292]_ ;
  assign \new_[76297]_  = \new_[76296]_  & \new_[76289]_ ;
  assign \new_[76300]_  = A233 & A232;
  assign \new_[76303]_  = ~A266 & ~A265;
  assign \new_[76304]_  = \new_[76303]_  & \new_[76300]_ ;
  assign \new_[76307]_  = ~A299 & A298;
  assign \new_[76310]_  = A302 & A300;
  assign \new_[76311]_  = \new_[76310]_  & \new_[76307]_ ;
  assign \new_[76312]_  = \new_[76311]_  & \new_[76304]_ ;
  assign \new_[76315]_  = ~A168 & A169;
  assign \new_[76318]_  = ~A166 & A167;
  assign \new_[76319]_  = \new_[76318]_  & \new_[76315]_ ;
  assign \new_[76322]_  = ~A200 & A199;
  assign \new_[76325]_  = A202 & A201;
  assign \new_[76326]_  = \new_[76325]_  & \new_[76322]_ ;
  assign \new_[76327]_  = \new_[76326]_  & \new_[76319]_ ;
  assign \new_[76330]_  = ~A235 & ~A233;
  assign \new_[76333]_  = ~A266 & ~A236;
  assign \new_[76334]_  = \new_[76333]_  & \new_[76330]_ ;
  assign \new_[76337]_  = ~A269 & ~A268;
  assign \new_[76340]_  = A299 & ~A298;
  assign \new_[76341]_  = \new_[76340]_  & \new_[76337]_ ;
  assign \new_[76342]_  = \new_[76341]_  & \new_[76334]_ ;
  assign \new_[76345]_  = ~A168 & A169;
  assign \new_[76348]_  = ~A166 & A167;
  assign \new_[76349]_  = \new_[76348]_  & \new_[76345]_ ;
  assign \new_[76352]_  = ~A200 & A199;
  assign \new_[76355]_  = A202 & A201;
  assign \new_[76356]_  = \new_[76355]_  & \new_[76352]_ ;
  assign \new_[76357]_  = \new_[76356]_  & \new_[76349]_ ;
  assign \new_[76360]_  = ~A234 & ~A233;
  assign \new_[76363]_  = A266 & A265;
  assign \new_[76364]_  = \new_[76363]_  & \new_[76360]_ ;
  assign \new_[76367]_  = ~A299 & A298;
  assign \new_[76370]_  = A301 & A300;
  assign \new_[76371]_  = \new_[76370]_  & \new_[76367]_ ;
  assign \new_[76372]_  = \new_[76371]_  & \new_[76364]_ ;
  assign \new_[76375]_  = ~A168 & A169;
  assign \new_[76378]_  = ~A166 & A167;
  assign \new_[76379]_  = \new_[76378]_  & \new_[76375]_ ;
  assign \new_[76382]_  = ~A200 & A199;
  assign \new_[76385]_  = A202 & A201;
  assign \new_[76386]_  = \new_[76385]_  & \new_[76382]_ ;
  assign \new_[76387]_  = \new_[76386]_  & \new_[76379]_ ;
  assign \new_[76390]_  = ~A234 & ~A233;
  assign \new_[76393]_  = A266 & A265;
  assign \new_[76394]_  = \new_[76393]_  & \new_[76390]_ ;
  assign \new_[76397]_  = ~A299 & A298;
  assign \new_[76400]_  = A302 & A300;
  assign \new_[76401]_  = \new_[76400]_  & \new_[76397]_ ;
  assign \new_[76402]_  = \new_[76401]_  & \new_[76394]_ ;
  assign \new_[76405]_  = ~A168 & A169;
  assign \new_[76408]_  = ~A166 & A167;
  assign \new_[76409]_  = \new_[76408]_  & \new_[76405]_ ;
  assign \new_[76412]_  = ~A200 & A199;
  assign \new_[76415]_  = A202 & A201;
  assign \new_[76416]_  = \new_[76415]_  & \new_[76412]_ ;
  assign \new_[76417]_  = \new_[76416]_  & \new_[76409]_ ;
  assign \new_[76420]_  = ~A234 & ~A233;
  assign \new_[76423]_  = ~A267 & ~A266;
  assign \new_[76424]_  = \new_[76423]_  & \new_[76420]_ ;
  assign \new_[76427]_  = ~A299 & A298;
  assign \new_[76430]_  = A301 & A300;
  assign \new_[76431]_  = \new_[76430]_  & \new_[76427]_ ;
  assign \new_[76432]_  = \new_[76431]_  & \new_[76424]_ ;
  assign \new_[76435]_  = ~A168 & A169;
  assign \new_[76438]_  = ~A166 & A167;
  assign \new_[76439]_  = \new_[76438]_  & \new_[76435]_ ;
  assign \new_[76442]_  = ~A200 & A199;
  assign \new_[76445]_  = A202 & A201;
  assign \new_[76446]_  = \new_[76445]_  & \new_[76442]_ ;
  assign \new_[76447]_  = \new_[76446]_  & \new_[76439]_ ;
  assign \new_[76450]_  = ~A234 & ~A233;
  assign \new_[76453]_  = ~A267 & ~A266;
  assign \new_[76454]_  = \new_[76453]_  & \new_[76450]_ ;
  assign \new_[76457]_  = ~A299 & A298;
  assign \new_[76460]_  = A302 & A300;
  assign \new_[76461]_  = \new_[76460]_  & \new_[76457]_ ;
  assign \new_[76462]_  = \new_[76461]_  & \new_[76454]_ ;
  assign \new_[76465]_  = ~A168 & A169;
  assign \new_[76468]_  = ~A166 & A167;
  assign \new_[76469]_  = \new_[76468]_  & \new_[76465]_ ;
  assign \new_[76472]_  = ~A200 & A199;
  assign \new_[76475]_  = A202 & A201;
  assign \new_[76476]_  = \new_[76475]_  & \new_[76472]_ ;
  assign \new_[76477]_  = \new_[76476]_  & \new_[76469]_ ;
  assign \new_[76480]_  = ~A234 & ~A233;
  assign \new_[76483]_  = ~A266 & ~A265;
  assign \new_[76484]_  = \new_[76483]_  & \new_[76480]_ ;
  assign \new_[76487]_  = ~A299 & A298;
  assign \new_[76490]_  = A301 & A300;
  assign \new_[76491]_  = \new_[76490]_  & \new_[76487]_ ;
  assign \new_[76492]_  = \new_[76491]_  & \new_[76484]_ ;
  assign \new_[76495]_  = ~A168 & A169;
  assign \new_[76498]_  = ~A166 & A167;
  assign \new_[76499]_  = \new_[76498]_  & \new_[76495]_ ;
  assign \new_[76502]_  = ~A200 & A199;
  assign \new_[76505]_  = A202 & A201;
  assign \new_[76506]_  = \new_[76505]_  & \new_[76502]_ ;
  assign \new_[76507]_  = \new_[76506]_  & \new_[76499]_ ;
  assign \new_[76510]_  = ~A234 & ~A233;
  assign \new_[76513]_  = ~A266 & ~A265;
  assign \new_[76514]_  = \new_[76513]_  & \new_[76510]_ ;
  assign \new_[76517]_  = ~A299 & A298;
  assign \new_[76520]_  = A302 & A300;
  assign \new_[76521]_  = \new_[76520]_  & \new_[76517]_ ;
  assign \new_[76522]_  = \new_[76521]_  & \new_[76514]_ ;
  assign \new_[76525]_  = ~A168 & A169;
  assign \new_[76528]_  = ~A166 & A167;
  assign \new_[76529]_  = \new_[76528]_  & \new_[76525]_ ;
  assign \new_[76532]_  = ~A200 & A199;
  assign \new_[76535]_  = A202 & A201;
  assign \new_[76536]_  = \new_[76535]_  & \new_[76532]_ ;
  assign \new_[76537]_  = \new_[76536]_  & \new_[76529]_ ;
  assign \new_[76540]_  = ~A233 & A232;
  assign \new_[76543]_  = A235 & A234;
  assign \new_[76544]_  = \new_[76543]_  & \new_[76540]_ ;
  assign \new_[76547]_  = ~A266 & A265;
  assign \new_[76550]_  = A268 & A267;
  assign \new_[76551]_  = \new_[76550]_  & \new_[76547]_ ;
  assign \new_[76552]_  = \new_[76551]_  & \new_[76544]_ ;
  assign \new_[76555]_  = ~A168 & A169;
  assign \new_[76558]_  = ~A166 & A167;
  assign \new_[76559]_  = \new_[76558]_  & \new_[76555]_ ;
  assign \new_[76562]_  = ~A200 & A199;
  assign \new_[76565]_  = A202 & A201;
  assign \new_[76566]_  = \new_[76565]_  & \new_[76562]_ ;
  assign \new_[76567]_  = \new_[76566]_  & \new_[76559]_ ;
  assign \new_[76570]_  = ~A233 & A232;
  assign \new_[76573]_  = A235 & A234;
  assign \new_[76574]_  = \new_[76573]_  & \new_[76570]_ ;
  assign \new_[76577]_  = ~A266 & A265;
  assign \new_[76580]_  = A269 & A267;
  assign \new_[76581]_  = \new_[76580]_  & \new_[76577]_ ;
  assign \new_[76582]_  = \new_[76581]_  & \new_[76574]_ ;
  assign \new_[76585]_  = ~A168 & A169;
  assign \new_[76588]_  = ~A166 & A167;
  assign \new_[76589]_  = \new_[76588]_  & \new_[76585]_ ;
  assign \new_[76592]_  = ~A200 & A199;
  assign \new_[76595]_  = A202 & A201;
  assign \new_[76596]_  = \new_[76595]_  & \new_[76592]_ ;
  assign \new_[76597]_  = \new_[76596]_  & \new_[76589]_ ;
  assign \new_[76600]_  = ~A233 & A232;
  assign \new_[76603]_  = A236 & A234;
  assign \new_[76604]_  = \new_[76603]_  & \new_[76600]_ ;
  assign \new_[76607]_  = ~A266 & A265;
  assign \new_[76610]_  = A268 & A267;
  assign \new_[76611]_  = \new_[76610]_  & \new_[76607]_ ;
  assign \new_[76612]_  = \new_[76611]_  & \new_[76604]_ ;
  assign \new_[76615]_  = ~A168 & A169;
  assign \new_[76618]_  = ~A166 & A167;
  assign \new_[76619]_  = \new_[76618]_  & \new_[76615]_ ;
  assign \new_[76622]_  = ~A200 & A199;
  assign \new_[76625]_  = A202 & A201;
  assign \new_[76626]_  = \new_[76625]_  & \new_[76622]_ ;
  assign \new_[76627]_  = \new_[76626]_  & \new_[76619]_ ;
  assign \new_[76630]_  = ~A233 & A232;
  assign \new_[76633]_  = A236 & A234;
  assign \new_[76634]_  = \new_[76633]_  & \new_[76630]_ ;
  assign \new_[76637]_  = ~A266 & A265;
  assign \new_[76640]_  = A269 & A267;
  assign \new_[76641]_  = \new_[76640]_  & \new_[76637]_ ;
  assign \new_[76642]_  = \new_[76641]_  & \new_[76634]_ ;
  assign \new_[76645]_  = ~A168 & A169;
  assign \new_[76648]_  = ~A166 & A167;
  assign \new_[76649]_  = \new_[76648]_  & \new_[76645]_ ;
  assign \new_[76652]_  = ~A200 & A199;
  assign \new_[76655]_  = A202 & A201;
  assign \new_[76656]_  = \new_[76655]_  & \new_[76652]_ ;
  assign \new_[76657]_  = \new_[76656]_  & \new_[76649]_ ;
  assign \new_[76660]_  = ~A233 & ~A232;
  assign \new_[76663]_  = A266 & A265;
  assign \new_[76664]_  = \new_[76663]_  & \new_[76660]_ ;
  assign \new_[76667]_  = ~A299 & A298;
  assign \new_[76670]_  = A301 & A300;
  assign \new_[76671]_  = \new_[76670]_  & \new_[76667]_ ;
  assign \new_[76672]_  = \new_[76671]_  & \new_[76664]_ ;
  assign \new_[76675]_  = ~A168 & A169;
  assign \new_[76678]_  = ~A166 & A167;
  assign \new_[76679]_  = \new_[76678]_  & \new_[76675]_ ;
  assign \new_[76682]_  = ~A200 & A199;
  assign \new_[76685]_  = A202 & A201;
  assign \new_[76686]_  = \new_[76685]_  & \new_[76682]_ ;
  assign \new_[76687]_  = \new_[76686]_  & \new_[76679]_ ;
  assign \new_[76690]_  = ~A233 & ~A232;
  assign \new_[76693]_  = A266 & A265;
  assign \new_[76694]_  = \new_[76693]_  & \new_[76690]_ ;
  assign \new_[76697]_  = ~A299 & A298;
  assign \new_[76700]_  = A302 & A300;
  assign \new_[76701]_  = \new_[76700]_  & \new_[76697]_ ;
  assign \new_[76702]_  = \new_[76701]_  & \new_[76694]_ ;
  assign \new_[76705]_  = ~A168 & A169;
  assign \new_[76708]_  = ~A166 & A167;
  assign \new_[76709]_  = \new_[76708]_  & \new_[76705]_ ;
  assign \new_[76712]_  = ~A200 & A199;
  assign \new_[76715]_  = A202 & A201;
  assign \new_[76716]_  = \new_[76715]_  & \new_[76712]_ ;
  assign \new_[76717]_  = \new_[76716]_  & \new_[76709]_ ;
  assign \new_[76720]_  = ~A233 & ~A232;
  assign \new_[76723]_  = ~A267 & ~A266;
  assign \new_[76724]_  = \new_[76723]_  & \new_[76720]_ ;
  assign \new_[76727]_  = ~A299 & A298;
  assign \new_[76730]_  = A301 & A300;
  assign \new_[76731]_  = \new_[76730]_  & \new_[76727]_ ;
  assign \new_[76732]_  = \new_[76731]_  & \new_[76724]_ ;
  assign \new_[76735]_  = ~A168 & A169;
  assign \new_[76738]_  = ~A166 & A167;
  assign \new_[76739]_  = \new_[76738]_  & \new_[76735]_ ;
  assign \new_[76742]_  = ~A200 & A199;
  assign \new_[76745]_  = A202 & A201;
  assign \new_[76746]_  = \new_[76745]_  & \new_[76742]_ ;
  assign \new_[76747]_  = \new_[76746]_  & \new_[76739]_ ;
  assign \new_[76750]_  = ~A233 & ~A232;
  assign \new_[76753]_  = ~A267 & ~A266;
  assign \new_[76754]_  = \new_[76753]_  & \new_[76750]_ ;
  assign \new_[76757]_  = ~A299 & A298;
  assign \new_[76760]_  = A302 & A300;
  assign \new_[76761]_  = \new_[76760]_  & \new_[76757]_ ;
  assign \new_[76762]_  = \new_[76761]_  & \new_[76754]_ ;
  assign \new_[76765]_  = ~A168 & A169;
  assign \new_[76768]_  = ~A166 & A167;
  assign \new_[76769]_  = \new_[76768]_  & \new_[76765]_ ;
  assign \new_[76772]_  = ~A200 & A199;
  assign \new_[76775]_  = A202 & A201;
  assign \new_[76776]_  = \new_[76775]_  & \new_[76772]_ ;
  assign \new_[76777]_  = \new_[76776]_  & \new_[76769]_ ;
  assign \new_[76780]_  = ~A233 & ~A232;
  assign \new_[76783]_  = ~A266 & ~A265;
  assign \new_[76784]_  = \new_[76783]_  & \new_[76780]_ ;
  assign \new_[76787]_  = ~A299 & A298;
  assign \new_[76790]_  = A301 & A300;
  assign \new_[76791]_  = \new_[76790]_  & \new_[76787]_ ;
  assign \new_[76792]_  = \new_[76791]_  & \new_[76784]_ ;
  assign \new_[76795]_  = ~A168 & A169;
  assign \new_[76798]_  = ~A166 & A167;
  assign \new_[76799]_  = \new_[76798]_  & \new_[76795]_ ;
  assign \new_[76802]_  = ~A200 & A199;
  assign \new_[76805]_  = A202 & A201;
  assign \new_[76806]_  = \new_[76805]_  & \new_[76802]_ ;
  assign \new_[76807]_  = \new_[76806]_  & \new_[76799]_ ;
  assign \new_[76810]_  = ~A233 & ~A232;
  assign \new_[76813]_  = ~A266 & ~A265;
  assign \new_[76814]_  = \new_[76813]_  & \new_[76810]_ ;
  assign \new_[76817]_  = ~A299 & A298;
  assign \new_[76820]_  = A302 & A300;
  assign \new_[76821]_  = \new_[76820]_  & \new_[76817]_ ;
  assign \new_[76822]_  = \new_[76821]_  & \new_[76814]_ ;
  assign \new_[76825]_  = ~A168 & A169;
  assign \new_[76828]_  = ~A166 & A167;
  assign \new_[76829]_  = \new_[76828]_  & \new_[76825]_ ;
  assign \new_[76832]_  = ~A200 & A199;
  assign \new_[76835]_  = A203 & A201;
  assign \new_[76836]_  = \new_[76835]_  & \new_[76832]_ ;
  assign \new_[76837]_  = \new_[76836]_  & \new_[76829]_ ;
  assign \new_[76840]_  = A233 & A232;
  assign \new_[76843]_  = ~A267 & A265;
  assign \new_[76844]_  = \new_[76843]_  & \new_[76840]_ ;
  assign \new_[76847]_  = ~A299 & A298;
  assign \new_[76850]_  = A301 & A300;
  assign \new_[76851]_  = \new_[76850]_  & \new_[76847]_ ;
  assign \new_[76852]_  = \new_[76851]_  & \new_[76844]_ ;
  assign \new_[76855]_  = ~A168 & A169;
  assign \new_[76858]_  = ~A166 & A167;
  assign \new_[76859]_  = \new_[76858]_  & \new_[76855]_ ;
  assign \new_[76862]_  = ~A200 & A199;
  assign \new_[76865]_  = A203 & A201;
  assign \new_[76866]_  = \new_[76865]_  & \new_[76862]_ ;
  assign \new_[76867]_  = \new_[76866]_  & \new_[76859]_ ;
  assign \new_[76870]_  = A233 & A232;
  assign \new_[76873]_  = ~A267 & A265;
  assign \new_[76874]_  = \new_[76873]_  & \new_[76870]_ ;
  assign \new_[76877]_  = ~A299 & A298;
  assign \new_[76880]_  = A302 & A300;
  assign \new_[76881]_  = \new_[76880]_  & \new_[76877]_ ;
  assign \new_[76882]_  = \new_[76881]_  & \new_[76874]_ ;
  assign \new_[76885]_  = ~A168 & A169;
  assign \new_[76888]_  = ~A166 & A167;
  assign \new_[76889]_  = \new_[76888]_  & \new_[76885]_ ;
  assign \new_[76892]_  = ~A200 & A199;
  assign \new_[76895]_  = A203 & A201;
  assign \new_[76896]_  = \new_[76895]_  & \new_[76892]_ ;
  assign \new_[76897]_  = \new_[76896]_  & \new_[76889]_ ;
  assign \new_[76900]_  = A233 & A232;
  assign \new_[76903]_  = A266 & A265;
  assign \new_[76904]_  = \new_[76903]_  & \new_[76900]_ ;
  assign \new_[76907]_  = ~A299 & A298;
  assign \new_[76910]_  = A301 & A300;
  assign \new_[76911]_  = \new_[76910]_  & \new_[76907]_ ;
  assign \new_[76912]_  = \new_[76911]_  & \new_[76904]_ ;
  assign \new_[76915]_  = ~A168 & A169;
  assign \new_[76918]_  = ~A166 & A167;
  assign \new_[76919]_  = \new_[76918]_  & \new_[76915]_ ;
  assign \new_[76922]_  = ~A200 & A199;
  assign \new_[76925]_  = A203 & A201;
  assign \new_[76926]_  = \new_[76925]_  & \new_[76922]_ ;
  assign \new_[76927]_  = \new_[76926]_  & \new_[76919]_ ;
  assign \new_[76930]_  = A233 & A232;
  assign \new_[76933]_  = A266 & A265;
  assign \new_[76934]_  = \new_[76933]_  & \new_[76930]_ ;
  assign \new_[76937]_  = ~A299 & A298;
  assign \new_[76940]_  = A302 & A300;
  assign \new_[76941]_  = \new_[76940]_  & \new_[76937]_ ;
  assign \new_[76942]_  = \new_[76941]_  & \new_[76934]_ ;
  assign \new_[76945]_  = ~A168 & A169;
  assign \new_[76948]_  = ~A166 & A167;
  assign \new_[76949]_  = \new_[76948]_  & \new_[76945]_ ;
  assign \new_[76952]_  = ~A200 & A199;
  assign \new_[76955]_  = A203 & A201;
  assign \new_[76956]_  = \new_[76955]_  & \new_[76952]_ ;
  assign \new_[76957]_  = \new_[76956]_  & \new_[76949]_ ;
  assign \new_[76960]_  = A233 & A232;
  assign \new_[76963]_  = ~A266 & ~A265;
  assign \new_[76964]_  = \new_[76963]_  & \new_[76960]_ ;
  assign \new_[76967]_  = ~A299 & A298;
  assign \new_[76970]_  = A301 & A300;
  assign \new_[76971]_  = \new_[76970]_  & \new_[76967]_ ;
  assign \new_[76972]_  = \new_[76971]_  & \new_[76964]_ ;
  assign \new_[76975]_  = ~A168 & A169;
  assign \new_[76978]_  = ~A166 & A167;
  assign \new_[76979]_  = \new_[76978]_  & \new_[76975]_ ;
  assign \new_[76982]_  = ~A200 & A199;
  assign \new_[76985]_  = A203 & A201;
  assign \new_[76986]_  = \new_[76985]_  & \new_[76982]_ ;
  assign \new_[76987]_  = \new_[76986]_  & \new_[76979]_ ;
  assign \new_[76990]_  = A233 & A232;
  assign \new_[76993]_  = ~A266 & ~A265;
  assign \new_[76994]_  = \new_[76993]_  & \new_[76990]_ ;
  assign \new_[76997]_  = ~A299 & A298;
  assign \new_[77000]_  = A302 & A300;
  assign \new_[77001]_  = \new_[77000]_  & \new_[76997]_ ;
  assign \new_[77002]_  = \new_[77001]_  & \new_[76994]_ ;
  assign \new_[77005]_  = ~A168 & A169;
  assign \new_[77008]_  = ~A166 & A167;
  assign \new_[77009]_  = \new_[77008]_  & \new_[77005]_ ;
  assign \new_[77012]_  = ~A200 & A199;
  assign \new_[77015]_  = A203 & A201;
  assign \new_[77016]_  = \new_[77015]_  & \new_[77012]_ ;
  assign \new_[77017]_  = \new_[77016]_  & \new_[77009]_ ;
  assign \new_[77020]_  = ~A235 & ~A233;
  assign \new_[77023]_  = ~A266 & ~A236;
  assign \new_[77024]_  = \new_[77023]_  & \new_[77020]_ ;
  assign \new_[77027]_  = ~A269 & ~A268;
  assign \new_[77030]_  = A299 & ~A298;
  assign \new_[77031]_  = \new_[77030]_  & \new_[77027]_ ;
  assign \new_[77032]_  = \new_[77031]_  & \new_[77024]_ ;
  assign \new_[77035]_  = ~A168 & A169;
  assign \new_[77038]_  = ~A166 & A167;
  assign \new_[77039]_  = \new_[77038]_  & \new_[77035]_ ;
  assign \new_[77042]_  = ~A200 & A199;
  assign \new_[77045]_  = A203 & A201;
  assign \new_[77046]_  = \new_[77045]_  & \new_[77042]_ ;
  assign \new_[77047]_  = \new_[77046]_  & \new_[77039]_ ;
  assign \new_[77050]_  = ~A234 & ~A233;
  assign \new_[77053]_  = A266 & A265;
  assign \new_[77054]_  = \new_[77053]_  & \new_[77050]_ ;
  assign \new_[77057]_  = ~A299 & A298;
  assign \new_[77060]_  = A301 & A300;
  assign \new_[77061]_  = \new_[77060]_  & \new_[77057]_ ;
  assign \new_[77062]_  = \new_[77061]_  & \new_[77054]_ ;
  assign \new_[77065]_  = ~A168 & A169;
  assign \new_[77068]_  = ~A166 & A167;
  assign \new_[77069]_  = \new_[77068]_  & \new_[77065]_ ;
  assign \new_[77072]_  = ~A200 & A199;
  assign \new_[77075]_  = A203 & A201;
  assign \new_[77076]_  = \new_[77075]_  & \new_[77072]_ ;
  assign \new_[77077]_  = \new_[77076]_  & \new_[77069]_ ;
  assign \new_[77080]_  = ~A234 & ~A233;
  assign \new_[77083]_  = A266 & A265;
  assign \new_[77084]_  = \new_[77083]_  & \new_[77080]_ ;
  assign \new_[77087]_  = ~A299 & A298;
  assign \new_[77090]_  = A302 & A300;
  assign \new_[77091]_  = \new_[77090]_  & \new_[77087]_ ;
  assign \new_[77092]_  = \new_[77091]_  & \new_[77084]_ ;
  assign \new_[77095]_  = ~A168 & A169;
  assign \new_[77098]_  = ~A166 & A167;
  assign \new_[77099]_  = \new_[77098]_  & \new_[77095]_ ;
  assign \new_[77102]_  = ~A200 & A199;
  assign \new_[77105]_  = A203 & A201;
  assign \new_[77106]_  = \new_[77105]_  & \new_[77102]_ ;
  assign \new_[77107]_  = \new_[77106]_  & \new_[77099]_ ;
  assign \new_[77110]_  = ~A234 & ~A233;
  assign \new_[77113]_  = ~A267 & ~A266;
  assign \new_[77114]_  = \new_[77113]_  & \new_[77110]_ ;
  assign \new_[77117]_  = ~A299 & A298;
  assign \new_[77120]_  = A301 & A300;
  assign \new_[77121]_  = \new_[77120]_  & \new_[77117]_ ;
  assign \new_[77122]_  = \new_[77121]_  & \new_[77114]_ ;
  assign \new_[77125]_  = ~A168 & A169;
  assign \new_[77128]_  = ~A166 & A167;
  assign \new_[77129]_  = \new_[77128]_  & \new_[77125]_ ;
  assign \new_[77132]_  = ~A200 & A199;
  assign \new_[77135]_  = A203 & A201;
  assign \new_[77136]_  = \new_[77135]_  & \new_[77132]_ ;
  assign \new_[77137]_  = \new_[77136]_  & \new_[77129]_ ;
  assign \new_[77140]_  = ~A234 & ~A233;
  assign \new_[77143]_  = ~A267 & ~A266;
  assign \new_[77144]_  = \new_[77143]_  & \new_[77140]_ ;
  assign \new_[77147]_  = ~A299 & A298;
  assign \new_[77150]_  = A302 & A300;
  assign \new_[77151]_  = \new_[77150]_  & \new_[77147]_ ;
  assign \new_[77152]_  = \new_[77151]_  & \new_[77144]_ ;
  assign \new_[77155]_  = ~A168 & A169;
  assign \new_[77158]_  = ~A166 & A167;
  assign \new_[77159]_  = \new_[77158]_  & \new_[77155]_ ;
  assign \new_[77162]_  = ~A200 & A199;
  assign \new_[77165]_  = A203 & A201;
  assign \new_[77166]_  = \new_[77165]_  & \new_[77162]_ ;
  assign \new_[77167]_  = \new_[77166]_  & \new_[77159]_ ;
  assign \new_[77170]_  = ~A234 & ~A233;
  assign \new_[77173]_  = ~A266 & ~A265;
  assign \new_[77174]_  = \new_[77173]_  & \new_[77170]_ ;
  assign \new_[77177]_  = ~A299 & A298;
  assign \new_[77180]_  = A301 & A300;
  assign \new_[77181]_  = \new_[77180]_  & \new_[77177]_ ;
  assign \new_[77182]_  = \new_[77181]_  & \new_[77174]_ ;
  assign \new_[77185]_  = ~A168 & A169;
  assign \new_[77188]_  = ~A166 & A167;
  assign \new_[77189]_  = \new_[77188]_  & \new_[77185]_ ;
  assign \new_[77192]_  = ~A200 & A199;
  assign \new_[77195]_  = A203 & A201;
  assign \new_[77196]_  = \new_[77195]_  & \new_[77192]_ ;
  assign \new_[77197]_  = \new_[77196]_  & \new_[77189]_ ;
  assign \new_[77200]_  = ~A234 & ~A233;
  assign \new_[77203]_  = ~A266 & ~A265;
  assign \new_[77204]_  = \new_[77203]_  & \new_[77200]_ ;
  assign \new_[77207]_  = ~A299 & A298;
  assign \new_[77210]_  = A302 & A300;
  assign \new_[77211]_  = \new_[77210]_  & \new_[77207]_ ;
  assign \new_[77212]_  = \new_[77211]_  & \new_[77204]_ ;
  assign \new_[77215]_  = ~A168 & A169;
  assign \new_[77218]_  = ~A166 & A167;
  assign \new_[77219]_  = \new_[77218]_  & \new_[77215]_ ;
  assign \new_[77222]_  = ~A200 & A199;
  assign \new_[77225]_  = A203 & A201;
  assign \new_[77226]_  = \new_[77225]_  & \new_[77222]_ ;
  assign \new_[77227]_  = \new_[77226]_  & \new_[77219]_ ;
  assign \new_[77230]_  = ~A233 & A232;
  assign \new_[77233]_  = A235 & A234;
  assign \new_[77234]_  = \new_[77233]_  & \new_[77230]_ ;
  assign \new_[77237]_  = ~A266 & A265;
  assign \new_[77240]_  = A268 & A267;
  assign \new_[77241]_  = \new_[77240]_  & \new_[77237]_ ;
  assign \new_[77242]_  = \new_[77241]_  & \new_[77234]_ ;
  assign \new_[77245]_  = ~A168 & A169;
  assign \new_[77248]_  = ~A166 & A167;
  assign \new_[77249]_  = \new_[77248]_  & \new_[77245]_ ;
  assign \new_[77252]_  = ~A200 & A199;
  assign \new_[77255]_  = A203 & A201;
  assign \new_[77256]_  = \new_[77255]_  & \new_[77252]_ ;
  assign \new_[77257]_  = \new_[77256]_  & \new_[77249]_ ;
  assign \new_[77260]_  = ~A233 & A232;
  assign \new_[77263]_  = A235 & A234;
  assign \new_[77264]_  = \new_[77263]_  & \new_[77260]_ ;
  assign \new_[77267]_  = ~A266 & A265;
  assign \new_[77270]_  = A269 & A267;
  assign \new_[77271]_  = \new_[77270]_  & \new_[77267]_ ;
  assign \new_[77272]_  = \new_[77271]_  & \new_[77264]_ ;
  assign \new_[77275]_  = ~A168 & A169;
  assign \new_[77278]_  = ~A166 & A167;
  assign \new_[77279]_  = \new_[77278]_  & \new_[77275]_ ;
  assign \new_[77282]_  = ~A200 & A199;
  assign \new_[77285]_  = A203 & A201;
  assign \new_[77286]_  = \new_[77285]_  & \new_[77282]_ ;
  assign \new_[77287]_  = \new_[77286]_  & \new_[77279]_ ;
  assign \new_[77290]_  = ~A233 & A232;
  assign \new_[77293]_  = A236 & A234;
  assign \new_[77294]_  = \new_[77293]_  & \new_[77290]_ ;
  assign \new_[77297]_  = ~A266 & A265;
  assign \new_[77300]_  = A268 & A267;
  assign \new_[77301]_  = \new_[77300]_  & \new_[77297]_ ;
  assign \new_[77302]_  = \new_[77301]_  & \new_[77294]_ ;
  assign \new_[77305]_  = ~A168 & A169;
  assign \new_[77308]_  = ~A166 & A167;
  assign \new_[77309]_  = \new_[77308]_  & \new_[77305]_ ;
  assign \new_[77312]_  = ~A200 & A199;
  assign \new_[77315]_  = A203 & A201;
  assign \new_[77316]_  = \new_[77315]_  & \new_[77312]_ ;
  assign \new_[77317]_  = \new_[77316]_  & \new_[77309]_ ;
  assign \new_[77320]_  = ~A233 & A232;
  assign \new_[77323]_  = A236 & A234;
  assign \new_[77324]_  = \new_[77323]_  & \new_[77320]_ ;
  assign \new_[77327]_  = ~A266 & A265;
  assign \new_[77330]_  = A269 & A267;
  assign \new_[77331]_  = \new_[77330]_  & \new_[77327]_ ;
  assign \new_[77332]_  = \new_[77331]_  & \new_[77324]_ ;
  assign \new_[77335]_  = ~A168 & A169;
  assign \new_[77338]_  = ~A166 & A167;
  assign \new_[77339]_  = \new_[77338]_  & \new_[77335]_ ;
  assign \new_[77342]_  = ~A200 & A199;
  assign \new_[77345]_  = A203 & A201;
  assign \new_[77346]_  = \new_[77345]_  & \new_[77342]_ ;
  assign \new_[77347]_  = \new_[77346]_  & \new_[77339]_ ;
  assign \new_[77350]_  = ~A233 & ~A232;
  assign \new_[77353]_  = A266 & A265;
  assign \new_[77354]_  = \new_[77353]_  & \new_[77350]_ ;
  assign \new_[77357]_  = ~A299 & A298;
  assign \new_[77360]_  = A301 & A300;
  assign \new_[77361]_  = \new_[77360]_  & \new_[77357]_ ;
  assign \new_[77362]_  = \new_[77361]_  & \new_[77354]_ ;
  assign \new_[77365]_  = ~A168 & A169;
  assign \new_[77368]_  = ~A166 & A167;
  assign \new_[77369]_  = \new_[77368]_  & \new_[77365]_ ;
  assign \new_[77372]_  = ~A200 & A199;
  assign \new_[77375]_  = A203 & A201;
  assign \new_[77376]_  = \new_[77375]_  & \new_[77372]_ ;
  assign \new_[77377]_  = \new_[77376]_  & \new_[77369]_ ;
  assign \new_[77380]_  = ~A233 & ~A232;
  assign \new_[77383]_  = A266 & A265;
  assign \new_[77384]_  = \new_[77383]_  & \new_[77380]_ ;
  assign \new_[77387]_  = ~A299 & A298;
  assign \new_[77390]_  = A302 & A300;
  assign \new_[77391]_  = \new_[77390]_  & \new_[77387]_ ;
  assign \new_[77392]_  = \new_[77391]_  & \new_[77384]_ ;
  assign \new_[77395]_  = ~A168 & A169;
  assign \new_[77398]_  = ~A166 & A167;
  assign \new_[77399]_  = \new_[77398]_  & \new_[77395]_ ;
  assign \new_[77402]_  = ~A200 & A199;
  assign \new_[77405]_  = A203 & A201;
  assign \new_[77406]_  = \new_[77405]_  & \new_[77402]_ ;
  assign \new_[77407]_  = \new_[77406]_  & \new_[77399]_ ;
  assign \new_[77410]_  = ~A233 & ~A232;
  assign \new_[77413]_  = ~A267 & ~A266;
  assign \new_[77414]_  = \new_[77413]_  & \new_[77410]_ ;
  assign \new_[77417]_  = ~A299 & A298;
  assign \new_[77420]_  = A301 & A300;
  assign \new_[77421]_  = \new_[77420]_  & \new_[77417]_ ;
  assign \new_[77422]_  = \new_[77421]_  & \new_[77414]_ ;
  assign \new_[77425]_  = ~A168 & A169;
  assign \new_[77428]_  = ~A166 & A167;
  assign \new_[77429]_  = \new_[77428]_  & \new_[77425]_ ;
  assign \new_[77432]_  = ~A200 & A199;
  assign \new_[77435]_  = A203 & A201;
  assign \new_[77436]_  = \new_[77435]_  & \new_[77432]_ ;
  assign \new_[77437]_  = \new_[77436]_  & \new_[77429]_ ;
  assign \new_[77440]_  = ~A233 & ~A232;
  assign \new_[77443]_  = ~A267 & ~A266;
  assign \new_[77444]_  = \new_[77443]_  & \new_[77440]_ ;
  assign \new_[77447]_  = ~A299 & A298;
  assign \new_[77450]_  = A302 & A300;
  assign \new_[77451]_  = \new_[77450]_  & \new_[77447]_ ;
  assign \new_[77452]_  = \new_[77451]_  & \new_[77444]_ ;
  assign \new_[77455]_  = ~A168 & A169;
  assign \new_[77458]_  = ~A166 & A167;
  assign \new_[77459]_  = \new_[77458]_  & \new_[77455]_ ;
  assign \new_[77462]_  = ~A200 & A199;
  assign \new_[77465]_  = A203 & A201;
  assign \new_[77466]_  = \new_[77465]_  & \new_[77462]_ ;
  assign \new_[77467]_  = \new_[77466]_  & \new_[77459]_ ;
  assign \new_[77470]_  = ~A233 & ~A232;
  assign \new_[77473]_  = ~A266 & ~A265;
  assign \new_[77474]_  = \new_[77473]_  & \new_[77470]_ ;
  assign \new_[77477]_  = ~A299 & A298;
  assign \new_[77480]_  = A301 & A300;
  assign \new_[77481]_  = \new_[77480]_  & \new_[77477]_ ;
  assign \new_[77482]_  = \new_[77481]_  & \new_[77474]_ ;
  assign \new_[77485]_  = ~A168 & A169;
  assign \new_[77488]_  = ~A166 & A167;
  assign \new_[77489]_  = \new_[77488]_  & \new_[77485]_ ;
  assign \new_[77492]_  = ~A200 & A199;
  assign \new_[77495]_  = A203 & A201;
  assign \new_[77496]_  = \new_[77495]_  & \new_[77492]_ ;
  assign \new_[77497]_  = \new_[77496]_  & \new_[77489]_ ;
  assign \new_[77500]_  = ~A233 & ~A232;
  assign \new_[77503]_  = ~A266 & ~A265;
  assign \new_[77504]_  = \new_[77503]_  & \new_[77500]_ ;
  assign \new_[77507]_  = ~A299 & A298;
  assign \new_[77510]_  = A302 & A300;
  assign \new_[77511]_  = \new_[77510]_  & \new_[77507]_ ;
  assign \new_[77512]_  = \new_[77511]_  & \new_[77504]_ ;
  assign \new_[77515]_  = ~A168 & A169;
  assign \new_[77518]_  = A166 & ~A167;
  assign \new_[77519]_  = \new_[77518]_  & \new_[77515]_ ;
  assign \new_[77522]_  = A200 & ~A199;
  assign \new_[77525]_  = ~A235 & ~A233;
  assign \new_[77526]_  = \new_[77525]_  & \new_[77522]_ ;
  assign \new_[77527]_  = \new_[77526]_  & \new_[77519]_ ;
  assign \new_[77530]_  = ~A266 & ~A236;
  assign \new_[77533]_  = ~A269 & ~A268;
  assign \new_[77534]_  = \new_[77533]_  & \new_[77530]_ ;
  assign \new_[77537]_  = ~A299 & A298;
  assign \new_[77540]_  = A301 & A300;
  assign \new_[77541]_  = \new_[77540]_  & \new_[77537]_ ;
  assign \new_[77542]_  = \new_[77541]_  & \new_[77534]_ ;
  assign \new_[77545]_  = ~A168 & A169;
  assign \new_[77548]_  = A166 & ~A167;
  assign \new_[77549]_  = \new_[77548]_  & \new_[77545]_ ;
  assign \new_[77552]_  = A200 & ~A199;
  assign \new_[77555]_  = ~A235 & ~A233;
  assign \new_[77556]_  = \new_[77555]_  & \new_[77552]_ ;
  assign \new_[77557]_  = \new_[77556]_  & \new_[77549]_ ;
  assign \new_[77560]_  = ~A266 & ~A236;
  assign \new_[77563]_  = ~A269 & ~A268;
  assign \new_[77564]_  = \new_[77563]_  & \new_[77560]_ ;
  assign \new_[77567]_  = ~A299 & A298;
  assign \new_[77570]_  = A302 & A300;
  assign \new_[77571]_  = \new_[77570]_  & \new_[77567]_ ;
  assign \new_[77572]_  = \new_[77571]_  & \new_[77564]_ ;
  assign \new_[77575]_  = ~A168 & A169;
  assign \new_[77578]_  = A166 & ~A167;
  assign \new_[77579]_  = \new_[77578]_  & \new_[77575]_ ;
  assign \new_[77582]_  = ~A200 & A199;
  assign \new_[77585]_  = A202 & A201;
  assign \new_[77586]_  = \new_[77585]_  & \new_[77582]_ ;
  assign \new_[77587]_  = \new_[77586]_  & \new_[77579]_ ;
  assign \new_[77590]_  = A233 & A232;
  assign \new_[77593]_  = ~A267 & A265;
  assign \new_[77594]_  = \new_[77593]_  & \new_[77590]_ ;
  assign \new_[77597]_  = ~A299 & A298;
  assign \new_[77600]_  = A301 & A300;
  assign \new_[77601]_  = \new_[77600]_  & \new_[77597]_ ;
  assign \new_[77602]_  = \new_[77601]_  & \new_[77594]_ ;
  assign \new_[77605]_  = ~A168 & A169;
  assign \new_[77608]_  = A166 & ~A167;
  assign \new_[77609]_  = \new_[77608]_  & \new_[77605]_ ;
  assign \new_[77612]_  = ~A200 & A199;
  assign \new_[77615]_  = A202 & A201;
  assign \new_[77616]_  = \new_[77615]_  & \new_[77612]_ ;
  assign \new_[77617]_  = \new_[77616]_  & \new_[77609]_ ;
  assign \new_[77620]_  = A233 & A232;
  assign \new_[77623]_  = ~A267 & A265;
  assign \new_[77624]_  = \new_[77623]_  & \new_[77620]_ ;
  assign \new_[77627]_  = ~A299 & A298;
  assign \new_[77630]_  = A302 & A300;
  assign \new_[77631]_  = \new_[77630]_  & \new_[77627]_ ;
  assign \new_[77632]_  = \new_[77631]_  & \new_[77624]_ ;
  assign \new_[77635]_  = ~A168 & A169;
  assign \new_[77638]_  = A166 & ~A167;
  assign \new_[77639]_  = \new_[77638]_  & \new_[77635]_ ;
  assign \new_[77642]_  = ~A200 & A199;
  assign \new_[77645]_  = A202 & A201;
  assign \new_[77646]_  = \new_[77645]_  & \new_[77642]_ ;
  assign \new_[77647]_  = \new_[77646]_  & \new_[77639]_ ;
  assign \new_[77650]_  = A233 & A232;
  assign \new_[77653]_  = A266 & A265;
  assign \new_[77654]_  = \new_[77653]_  & \new_[77650]_ ;
  assign \new_[77657]_  = ~A299 & A298;
  assign \new_[77660]_  = A301 & A300;
  assign \new_[77661]_  = \new_[77660]_  & \new_[77657]_ ;
  assign \new_[77662]_  = \new_[77661]_  & \new_[77654]_ ;
  assign \new_[77665]_  = ~A168 & A169;
  assign \new_[77668]_  = A166 & ~A167;
  assign \new_[77669]_  = \new_[77668]_  & \new_[77665]_ ;
  assign \new_[77672]_  = ~A200 & A199;
  assign \new_[77675]_  = A202 & A201;
  assign \new_[77676]_  = \new_[77675]_  & \new_[77672]_ ;
  assign \new_[77677]_  = \new_[77676]_  & \new_[77669]_ ;
  assign \new_[77680]_  = A233 & A232;
  assign \new_[77683]_  = A266 & A265;
  assign \new_[77684]_  = \new_[77683]_  & \new_[77680]_ ;
  assign \new_[77687]_  = ~A299 & A298;
  assign \new_[77690]_  = A302 & A300;
  assign \new_[77691]_  = \new_[77690]_  & \new_[77687]_ ;
  assign \new_[77692]_  = \new_[77691]_  & \new_[77684]_ ;
  assign \new_[77695]_  = ~A168 & A169;
  assign \new_[77698]_  = A166 & ~A167;
  assign \new_[77699]_  = \new_[77698]_  & \new_[77695]_ ;
  assign \new_[77702]_  = ~A200 & A199;
  assign \new_[77705]_  = A202 & A201;
  assign \new_[77706]_  = \new_[77705]_  & \new_[77702]_ ;
  assign \new_[77707]_  = \new_[77706]_  & \new_[77699]_ ;
  assign \new_[77710]_  = A233 & A232;
  assign \new_[77713]_  = ~A266 & ~A265;
  assign \new_[77714]_  = \new_[77713]_  & \new_[77710]_ ;
  assign \new_[77717]_  = ~A299 & A298;
  assign \new_[77720]_  = A301 & A300;
  assign \new_[77721]_  = \new_[77720]_  & \new_[77717]_ ;
  assign \new_[77722]_  = \new_[77721]_  & \new_[77714]_ ;
  assign \new_[77725]_  = ~A168 & A169;
  assign \new_[77728]_  = A166 & ~A167;
  assign \new_[77729]_  = \new_[77728]_  & \new_[77725]_ ;
  assign \new_[77732]_  = ~A200 & A199;
  assign \new_[77735]_  = A202 & A201;
  assign \new_[77736]_  = \new_[77735]_  & \new_[77732]_ ;
  assign \new_[77737]_  = \new_[77736]_  & \new_[77729]_ ;
  assign \new_[77740]_  = A233 & A232;
  assign \new_[77743]_  = ~A266 & ~A265;
  assign \new_[77744]_  = \new_[77743]_  & \new_[77740]_ ;
  assign \new_[77747]_  = ~A299 & A298;
  assign \new_[77750]_  = A302 & A300;
  assign \new_[77751]_  = \new_[77750]_  & \new_[77747]_ ;
  assign \new_[77752]_  = \new_[77751]_  & \new_[77744]_ ;
  assign \new_[77755]_  = ~A168 & A169;
  assign \new_[77758]_  = A166 & ~A167;
  assign \new_[77759]_  = \new_[77758]_  & \new_[77755]_ ;
  assign \new_[77762]_  = ~A200 & A199;
  assign \new_[77765]_  = A202 & A201;
  assign \new_[77766]_  = \new_[77765]_  & \new_[77762]_ ;
  assign \new_[77767]_  = \new_[77766]_  & \new_[77759]_ ;
  assign \new_[77770]_  = ~A235 & ~A233;
  assign \new_[77773]_  = ~A266 & ~A236;
  assign \new_[77774]_  = \new_[77773]_  & \new_[77770]_ ;
  assign \new_[77777]_  = ~A269 & ~A268;
  assign \new_[77780]_  = A299 & ~A298;
  assign \new_[77781]_  = \new_[77780]_  & \new_[77777]_ ;
  assign \new_[77782]_  = \new_[77781]_  & \new_[77774]_ ;
  assign \new_[77785]_  = ~A168 & A169;
  assign \new_[77788]_  = A166 & ~A167;
  assign \new_[77789]_  = \new_[77788]_  & \new_[77785]_ ;
  assign \new_[77792]_  = ~A200 & A199;
  assign \new_[77795]_  = A202 & A201;
  assign \new_[77796]_  = \new_[77795]_  & \new_[77792]_ ;
  assign \new_[77797]_  = \new_[77796]_  & \new_[77789]_ ;
  assign \new_[77800]_  = ~A234 & ~A233;
  assign \new_[77803]_  = A266 & A265;
  assign \new_[77804]_  = \new_[77803]_  & \new_[77800]_ ;
  assign \new_[77807]_  = ~A299 & A298;
  assign \new_[77810]_  = A301 & A300;
  assign \new_[77811]_  = \new_[77810]_  & \new_[77807]_ ;
  assign \new_[77812]_  = \new_[77811]_  & \new_[77804]_ ;
  assign \new_[77815]_  = ~A168 & A169;
  assign \new_[77818]_  = A166 & ~A167;
  assign \new_[77819]_  = \new_[77818]_  & \new_[77815]_ ;
  assign \new_[77822]_  = ~A200 & A199;
  assign \new_[77825]_  = A202 & A201;
  assign \new_[77826]_  = \new_[77825]_  & \new_[77822]_ ;
  assign \new_[77827]_  = \new_[77826]_  & \new_[77819]_ ;
  assign \new_[77830]_  = ~A234 & ~A233;
  assign \new_[77833]_  = A266 & A265;
  assign \new_[77834]_  = \new_[77833]_  & \new_[77830]_ ;
  assign \new_[77837]_  = ~A299 & A298;
  assign \new_[77840]_  = A302 & A300;
  assign \new_[77841]_  = \new_[77840]_  & \new_[77837]_ ;
  assign \new_[77842]_  = \new_[77841]_  & \new_[77834]_ ;
  assign \new_[77845]_  = ~A168 & A169;
  assign \new_[77848]_  = A166 & ~A167;
  assign \new_[77849]_  = \new_[77848]_  & \new_[77845]_ ;
  assign \new_[77852]_  = ~A200 & A199;
  assign \new_[77855]_  = A202 & A201;
  assign \new_[77856]_  = \new_[77855]_  & \new_[77852]_ ;
  assign \new_[77857]_  = \new_[77856]_  & \new_[77849]_ ;
  assign \new_[77860]_  = ~A234 & ~A233;
  assign \new_[77863]_  = ~A267 & ~A266;
  assign \new_[77864]_  = \new_[77863]_  & \new_[77860]_ ;
  assign \new_[77867]_  = ~A299 & A298;
  assign \new_[77870]_  = A301 & A300;
  assign \new_[77871]_  = \new_[77870]_  & \new_[77867]_ ;
  assign \new_[77872]_  = \new_[77871]_  & \new_[77864]_ ;
  assign \new_[77875]_  = ~A168 & A169;
  assign \new_[77878]_  = A166 & ~A167;
  assign \new_[77879]_  = \new_[77878]_  & \new_[77875]_ ;
  assign \new_[77882]_  = ~A200 & A199;
  assign \new_[77885]_  = A202 & A201;
  assign \new_[77886]_  = \new_[77885]_  & \new_[77882]_ ;
  assign \new_[77887]_  = \new_[77886]_  & \new_[77879]_ ;
  assign \new_[77890]_  = ~A234 & ~A233;
  assign \new_[77893]_  = ~A267 & ~A266;
  assign \new_[77894]_  = \new_[77893]_  & \new_[77890]_ ;
  assign \new_[77897]_  = ~A299 & A298;
  assign \new_[77900]_  = A302 & A300;
  assign \new_[77901]_  = \new_[77900]_  & \new_[77897]_ ;
  assign \new_[77902]_  = \new_[77901]_  & \new_[77894]_ ;
  assign \new_[77905]_  = ~A168 & A169;
  assign \new_[77908]_  = A166 & ~A167;
  assign \new_[77909]_  = \new_[77908]_  & \new_[77905]_ ;
  assign \new_[77912]_  = ~A200 & A199;
  assign \new_[77915]_  = A202 & A201;
  assign \new_[77916]_  = \new_[77915]_  & \new_[77912]_ ;
  assign \new_[77917]_  = \new_[77916]_  & \new_[77909]_ ;
  assign \new_[77920]_  = ~A234 & ~A233;
  assign \new_[77923]_  = ~A266 & ~A265;
  assign \new_[77924]_  = \new_[77923]_  & \new_[77920]_ ;
  assign \new_[77927]_  = ~A299 & A298;
  assign \new_[77930]_  = A301 & A300;
  assign \new_[77931]_  = \new_[77930]_  & \new_[77927]_ ;
  assign \new_[77932]_  = \new_[77931]_  & \new_[77924]_ ;
  assign \new_[77935]_  = ~A168 & A169;
  assign \new_[77938]_  = A166 & ~A167;
  assign \new_[77939]_  = \new_[77938]_  & \new_[77935]_ ;
  assign \new_[77942]_  = ~A200 & A199;
  assign \new_[77945]_  = A202 & A201;
  assign \new_[77946]_  = \new_[77945]_  & \new_[77942]_ ;
  assign \new_[77947]_  = \new_[77946]_  & \new_[77939]_ ;
  assign \new_[77950]_  = ~A234 & ~A233;
  assign \new_[77953]_  = ~A266 & ~A265;
  assign \new_[77954]_  = \new_[77953]_  & \new_[77950]_ ;
  assign \new_[77957]_  = ~A299 & A298;
  assign \new_[77960]_  = A302 & A300;
  assign \new_[77961]_  = \new_[77960]_  & \new_[77957]_ ;
  assign \new_[77962]_  = \new_[77961]_  & \new_[77954]_ ;
  assign \new_[77965]_  = ~A168 & A169;
  assign \new_[77968]_  = A166 & ~A167;
  assign \new_[77969]_  = \new_[77968]_  & \new_[77965]_ ;
  assign \new_[77972]_  = ~A200 & A199;
  assign \new_[77975]_  = A202 & A201;
  assign \new_[77976]_  = \new_[77975]_  & \new_[77972]_ ;
  assign \new_[77977]_  = \new_[77976]_  & \new_[77969]_ ;
  assign \new_[77980]_  = ~A233 & A232;
  assign \new_[77983]_  = A235 & A234;
  assign \new_[77984]_  = \new_[77983]_  & \new_[77980]_ ;
  assign \new_[77987]_  = ~A266 & A265;
  assign \new_[77990]_  = A268 & A267;
  assign \new_[77991]_  = \new_[77990]_  & \new_[77987]_ ;
  assign \new_[77992]_  = \new_[77991]_  & \new_[77984]_ ;
  assign \new_[77995]_  = ~A168 & A169;
  assign \new_[77998]_  = A166 & ~A167;
  assign \new_[77999]_  = \new_[77998]_  & \new_[77995]_ ;
  assign \new_[78002]_  = ~A200 & A199;
  assign \new_[78005]_  = A202 & A201;
  assign \new_[78006]_  = \new_[78005]_  & \new_[78002]_ ;
  assign \new_[78007]_  = \new_[78006]_  & \new_[77999]_ ;
  assign \new_[78010]_  = ~A233 & A232;
  assign \new_[78013]_  = A235 & A234;
  assign \new_[78014]_  = \new_[78013]_  & \new_[78010]_ ;
  assign \new_[78017]_  = ~A266 & A265;
  assign \new_[78020]_  = A269 & A267;
  assign \new_[78021]_  = \new_[78020]_  & \new_[78017]_ ;
  assign \new_[78022]_  = \new_[78021]_  & \new_[78014]_ ;
  assign \new_[78025]_  = ~A168 & A169;
  assign \new_[78028]_  = A166 & ~A167;
  assign \new_[78029]_  = \new_[78028]_  & \new_[78025]_ ;
  assign \new_[78032]_  = ~A200 & A199;
  assign \new_[78035]_  = A202 & A201;
  assign \new_[78036]_  = \new_[78035]_  & \new_[78032]_ ;
  assign \new_[78037]_  = \new_[78036]_  & \new_[78029]_ ;
  assign \new_[78040]_  = ~A233 & A232;
  assign \new_[78043]_  = A236 & A234;
  assign \new_[78044]_  = \new_[78043]_  & \new_[78040]_ ;
  assign \new_[78047]_  = ~A266 & A265;
  assign \new_[78050]_  = A268 & A267;
  assign \new_[78051]_  = \new_[78050]_  & \new_[78047]_ ;
  assign \new_[78052]_  = \new_[78051]_  & \new_[78044]_ ;
  assign \new_[78055]_  = ~A168 & A169;
  assign \new_[78058]_  = A166 & ~A167;
  assign \new_[78059]_  = \new_[78058]_  & \new_[78055]_ ;
  assign \new_[78062]_  = ~A200 & A199;
  assign \new_[78065]_  = A202 & A201;
  assign \new_[78066]_  = \new_[78065]_  & \new_[78062]_ ;
  assign \new_[78067]_  = \new_[78066]_  & \new_[78059]_ ;
  assign \new_[78070]_  = ~A233 & A232;
  assign \new_[78073]_  = A236 & A234;
  assign \new_[78074]_  = \new_[78073]_  & \new_[78070]_ ;
  assign \new_[78077]_  = ~A266 & A265;
  assign \new_[78080]_  = A269 & A267;
  assign \new_[78081]_  = \new_[78080]_  & \new_[78077]_ ;
  assign \new_[78082]_  = \new_[78081]_  & \new_[78074]_ ;
  assign \new_[78085]_  = ~A168 & A169;
  assign \new_[78088]_  = A166 & ~A167;
  assign \new_[78089]_  = \new_[78088]_  & \new_[78085]_ ;
  assign \new_[78092]_  = ~A200 & A199;
  assign \new_[78095]_  = A202 & A201;
  assign \new_[78096]_  = \new_[78095]_  & \new_[78092]_ ;
  assign \new_[78097]_  = \new_[78096]_  & \new_[78089]_ ;
  assign \new_[78100]_  = ~A233 & ~A232;
  assign \new_[78103]_  = A266 & A265;
  assign \new_[78104]_  = \new_[78103]_  & \new_[78100]_ ;
  assign \new_[78107]_  = ~A299 & A298;
  assign \new_[78110]_  = A301 & A300;
  assign \new_[78111]_  = \new_[78110]_  & \new_[78107]_ ;
  assign \new_[78112]_  = \new_[78111]_  & \new_[78104]_ ;
  assign \new_[78115]_  = ~A168 & A169;
  assign \new_[78118]_  = A166 & ~A167;
  assign \new_[78119]_  = \new_[78118]_  & \new_[78115]_ ;
  assign \new_[78122]_  = ~A200 & A199;
  assign \new_[78125]_  = A202 & A201;
  assign \new_[78126]_  = \new_[78125]_  & \new_[78122]_ ;
  assign \new_[78127]_  = \new_[78126]_  & \new_[78119]_ ;
  assign \new_[78130]_  = ~A233 & ~A232;
  assign \new_[78133]_  = A266 & A265;
  assign \new_[78134]_  = \new_[78133]_  & \new_[78130]_ ;
  assign \new_[78137]_  = ~A299 & A298;
  assign \new_[78140]_  = A302 & A300;
  assign \new_[78141]_  = \new_[78140]_  & \new_[78137]_ ;
  assign \new_[78142]_  = \new_[78141]_  & \new_[78134]_ ;
  assign \new_[78145]_  = ~A168 & A169;
  assign \new_[78148]_  = A166 & ~A167;
  assign \new_[78149]_  = \new_[78148]_  & \new_[78145]_ ;
  assign \new_[78152]_  = ~A200 & A199;
  assign \new_[78155]_  = A202 & A201;
  assign \new_[78156]_  = \new_[78155]_  & \new_[78152]_ ;
  assign \new_[78157]_  = \new_[78156]_  & \new_[78149]_ ;
  assign \new_[78160]_  = ~A233 & ~A232;
  assign \new_[78163]_  = ~A267 & ~A266;
  assign \new_[78164]_  = \new_[78163]_  & \new_[78160]_ ;
  assign \new_[78167]_  = ~A299 & A298;
  assign \new_[78170]_  = A301 & A300;
  assign \new_[78171]_  = \new_[78170]_  & \new_[78167]_ ;
  assign \new_[78172]_  = \new_[78171]_  & \new_[78164]_ ;
  assign \new_[78175]_  = ~A168 & A169;
  assign \new_[78178]_  = A166 & ~A167;
  assign \new_[78179]_  = \new_[78178]_  & \new_[78175]_ ;
  assign \new_[78182]_  = ~A200 & A199;
  assign \new_[78185]_  = A202 & A201;
  assign \new_[78186]_  = \new_[78185]_  & \new_[78182]_ ;
  assign \new_[78187]_  = \new_[78186]_  & \new_[78179]_ ;
  assign \new_[78190]_  = ~A233 & ~A232;
  assign \new_[78193]_  = ~A267 & ~A266;
  assign \new_[78194]_  = \new_[78193]_  & \new_[78190]_ ;
  assign \new_[78197]_  = ~A299 & A298;
  assign \new_[78200]_  = A302 & A300;
  assign \new_[78201]_  = \new_[78200]_  & \new_[78197]_ ;
  assign \new_[78202]_  = \new_[78201]_  & \new_[78194]_ ;
  assign \new_[78205]_  = ~A168 & A169;
  assign \new_[78208]_  = A166 & ~A167;
  assign \new_[78209]_  = \new_[78208]_  & \new_[78205]_ ;
  assign \new_[78212]_  = ~A200 & A199;
  assign \new_[78215]_  = A202 & A201;
  assign \new_[78216]_  = \new_[78215]_  & \new_[78212]_ ;
  assign \new_[78217]_  = \new_[78216]_  & \new_[78209]_ ;
  assign \new_[78220]_  = ~A233 & ~A232;
  assign \new_[78223]_  = ~A266 & ~A265;
  assign \new_[78224]_  = \new_[78223]_  & \new_[78220]_ ;
  assign \new_[78227]_  = ~A299 & A298;
  assign \new_[78230]_  = A301 & A300;
  assign \new_[78231]_  = \new_[78230]_  & \new_[78227]_ ;
  assign \new_[78232]_  = \new_[78231]_  & \new_[78224]_ ;
  assign \new_[78235]_  = ~A168 & A169;
  assign \new_[78238]_  = A166 & ~A167;
  assign \new_[78239]_  = \new_[78238]_  & \new_[78235]_ ;
  assign \new_[78242]_  = ~A200 & A199;
  assign \new_[78245]_  = A202 & A201;
  assign \new_[78246]_  = \new_[78245]_  & \new_[78242]_ ;
  assign \new_[78247]_  = \new_[78246]_  & \new_[78239]_ ;
  assign \new_[78250]_  = ~A233 & ~A232;
  assign \new_[78253]_  = ~A266 & ~A265;
  assign \new_[78254]_  = \new_[78253]_  & \new_[78250]_ ;
  assign \new_[78257]_  = ~A299 & A298;
  assign \new_[78260]_  = A302 & A300;
  assign \new_[78261]_  = \new_[78260]_  & \new_[78257]_ ;
  assign \new_[78262]_  = \new_[78261]_  & \new_[78254]_ ;
  assign \new_[78265]_  = ~A168 & A169;
  assign \new_[78268]_  = A166 & ~A167;
  assign \new_[78269]_  = \new_[78268]_  & \new_[78265]_ ;
  assign \new_[78272]_  = ~A200 & A199;
  assign \new_[78275]_  = A203 & A201;
  assign \new_[78276]_  = \new_[78275]_  & \new_[78272]_ ;
  assign \new_[78277]_  = \new_[78276]_  & \new_[78269]_ ;
  assign \new_[78280]_  = A233 & A232;
  assign \new_[78283]_  = ~A267 & A265;
  assign \new_[78284]_  = \new_[78283]_  & \new_[78280]_ ;
  assign \new_[78287]_  = ~A299 & A298;
  assign \new_[78290]_  = A301 & A300;
  assign \new_[78291]_  = \new_[78290]_  & \new_[78287]_ ;
  assign \new_[78292]_  = \new_[78291]_  & \new_[78284]_ ;
  assign \new_[78295]_  = ~A168 & A169;
  assign \new_[78298]_  = A166 & ~A167;
  assign \new_[78299]_  = \new_[78298]_  & \new_[78295]_ ;
  assign \new_[78302]_  = ~A200 & A199;
  assign \new_[78305]_  = A203 & A201;
  assign \new_[78306]_  = \new_[78305]_  & \new_[78302]_ ;
  assign \new_[78307]_  = \new_[78306]_  & \new_[78299]_ ;
  assign \new_[78310]_  = A233 & A232;
  assign \new_[78313]_  = ~A267 & A265;
  assign \new_[78314]_  = \new_[78313]_  & \new_[78310]_ ;
  assign \new_[78317]_  = ~A299 & A298;
  assign \new_[78320]_  = A302 & A300;
  assign \new_[78321]_  = \new_[78320]_  & \new_[78317]_ ;
  assign \new_[78322]_  = \new_[78321]_  & \new_[78314]_ ;
  assign \new_[78325]_  = ~A168 & A169;
  assign \new_[78328]_  = A166 & ~A167;
  assign \new_[78329]_  = \new_[78328]_  & \new_[78325]_ ;
  assign \new_[78332]_  = ~A200 & A199;
  assign \new_[78335]_  = A203 & A201;
  assign \new_[78336]_  = \new_[78335]_  & \new_[78332]_ ;
  assign \new_[78337]_  = \new_[78336]_  & \new_[78329]_ ;
  assign \new_[78340]_  = A233 & A232;
  assign \new_[78343]_  = A266 & A265;
  assign \new_[78344]_  = \new_[78343]_  & \new_[78340]_ ;
  assign \new_[78347]_  = ~A299 & A298;
  assign \new_[78350]_  = A301 & A300;
  assign \new_[78351]_  = \new_[78350]_  & \new_[78347]_ ;
  assign \new_[78352]_  = \new_[78351]_  & \new_[78344]_ ;
  assign \new_[78355]_  = ~A168 & A169;
  assign \new_[78358]_  = A166 & ~A167;
  assign \new_[78359]_  = \new_[78358]_  & \new_[78355]_ ;
  assign \new_[78362]_  = ~A200 & A199;
  assign \new_[78365]_  = A203 & A201;
  assign \new_[78366]_  = \new_[78365]_  & \new_[78362]_ ;
  assign \new_[78367]_  = \new_[78366]_  & \new_[78359]_ ;
  assign \new_[78370]_  = A233 & A232;
  assign \new_[78373]_  = A266 & A265;
  assign \new_[78374]_  = \new_[78373]_  & \new_[78370]_ ;
  assign \new_[78377]_  = ~A299 & A298;
  assign \new_[78380]_  = A302 & A300;
  assign \new_[78381]_  = \new_[78380]_  & \new_[78377]_ ;
  assign \new_[78382]_  = \new_[78381]_  & \new_[78374]_ ;
  assign \new_[78385]_  = ~A168 & A169;
  assign \new_[78388]_  = A166 & ~A167;
  assign \new_[78389]_  = \new_[78388]_  & \new_[78385]_ ;
  assign \new_[78392]_  = ~A200 & A199;
  assign \new_[78395]_  = A203 & A201;
  assign \new_[78396]_  = \new_[78395]_  & \new_[78392]_ ;
  assign \new_[78397]_  = \new_[78396]_  & \new_[78389]_ ;
  assign \new_[78400]_  = A233 & A232;
  assign \new_[78403]_  = ~A266 & ~A265;
  assign \new_[78404]_  = \new_[78403]_  & \new_[78400]_ ;
  assign \new_[78407]_  = ~A299 & A298;
  assign \new_[78410]_  = A301 & A300;
  assign \new_[78411]_  = \new_[78410]_  & \new_[78407]_ ;
  assign \new_[78412]_  = \new_[78411]_  & \new_[78404]_ ;
  assign \new_[78415]_  = ~A168 & A169;
  assign \new_[78418]_  = A166 & ~A167;
  assign \new_[78419]_  = \new_[78418]_  & \new_[78415]_ ;
  assign \new_[78422]_  = ~A200 & A199;
  assign \new_[78425]_  = A203 & A201;
  assign \new_[78426]_  = \new_[78425]_  & \new_[78422]_ ;
  assign \new_[78427]_  = \new_[78426]_  & \new_[78419]_ ;
  assign \new_[78430]_  = A233 & A232;
  assign \new_[78433]_  = ~A266 & ~A265;
  assign \new_[78434]_  = \new_[78433]_  & \new_[78430]_ ;
  assign \new_[78437]_  = ~A299 & A298;
  assign \new_[78440]_  = A302 & A300;
  assign \new_[78441]_  = \new_[78440]_  & \new_[78437]_ ;
  assign \new_[78442]_  = \new_[78441]_  & \new_[78434]_ ;
  assign \new_[78445]_  = ~A168 & A169;
  assign \new_[78448]_  = A166 & ~A167;
  assign \new_[78449]_  = \new_[78448]_  & \new_[78445]_ ;
  assign \new_[78452]_  = ~A200 & A199;
  assign \new_[78455]_  = A203 & A201;
  assign \new_[78456]_  = \new_[78455]_  & \new_[78452]_ ;
  assign \new_[78457]_  = \new_[78456]_  & \new_[78449]_ ;
  assign \new_[78460]_  = ~A235 & ~A233;
  assign \new_[78463]_  = ~A266 & ~A236;
  assign \new_[78464]_  = \new_[78463]_  & \new_[78460]_ ;
  assign \new_[78467]_  = ~A269 & ~A268;
  assign \new_[78470]_  = A299 & ~A298;
  assign \new_[78471]_  = \new_[78470]_  & \new_[78467]_ ;
  assign \new_[78472]_  = \new_[78471]_  & \new_[78464]_ ;
  assign \new_[78475]_  = ~A168 & A169;
  assign \new_[78478]_  = A166 & ~A167;
  assign \new_[78479]_  = \new_[78478]_  & \new_[78475]_ ;
  assign \new_[78482]_  = ~A200 & A199;
  assign \new_[78485]_  = A203 & A201;
  assign \new_[78486]_  = \new_[78485]_  & \new_[78482]_ ;
  assign \new_[78487]_  = \new_[78486]_  & \new_[78479]_ ;
  assign \new_[78490]_  = ~A234 & ~A233;
  assign \new_[78493]_  = A266 & A265;
  assign \new_[78494]_  = \new_[78493]_  & \new_[78490]_ ;
  assign \new_[78497]_  = ~A299 & A298;
  assign \new_[78500]_  = A301 & A300;
  assign \new_[78501]_  = \new_[78500]_  & \new_[78497]_ ;
  assign \new_[78502]_  = \new_[78501]_  & \new_[78494]_ ;
  assign \new_[78505]_  = ~A168 & A169;
  assign \new_[78508]_  = A166 & ~A167;
  assign \new_[78509]_  = \new_[78508]_  & \new_[78505]_ ;
  assign \new_[78512]_  = ~A200 & A199;
  assign \new_[78515]_  = A203 & A201;
  assign \new_[78516]_  = \new_[78515]_  & \new_[78512]_ ;
  assign \new_[78517]_  = \new_[78516]_  & \new_[78509]_ ;
  assign \new_[78520]_  = ~A234 & ~A233;
  assign \new_[78523]_  = A266 & A265;
  assign \new_[78524]_  = \new_[78523]_  & \new_[78520]_ ;
  assign \new_[78527]_  = ~A299 & A298;
  assign \new_[78530]_  = A302 & A300;
  assign \new_[78531]_  = \new_[78530]_  & \new_[78527]_ ;
  assign \new_[78532]_  = \new_[78531]_  & \new_[78524]_ ;
  assign \new_[78535]_  = ~A168 & A169;
  assign \new_[78538]_  = A166 & ~A167;
  assign \new_[78539]_  = \new_[78538]_  & \new_[78535]_ ;
  assign \new_[78542]_  = ~A200 & A199;
  assign \new_[78545]_  = A203 & A201;
  assign \new_[78546]_  = \new_[78545]_  & \new_[78542]_ ;
  assign \new_[78547]_  = \new_[78546]_  & \new_[78539]_ ;
  assign \new_[78550]_  = ~A234 & ~A233;
  assign \new_[78553]_  = ~A267 & ~A266;
  assign \new_[78554]_  = \new_[78553]_  & \new_[78550]_ ;
  assign \new_[78557]_  = ~A299 & A298;
  assign \new_[78560]_  = A301 & A300;
  assign \new_[78561]_  = \new_[78560]_  & \new_[78557]_ ;
  assign \new_[78562]_  = \new_[78561]_  & \new_[78554]_ ;
  assign \new_[78565]_  = ~A168 & A169;
  assign \new_[78568]_  = A166 & ~A167;
  assign \new_[78569]_  = \new_[78568]_  & \new_[78565]_ ;
  assign \new_[78572]_  = ~A200 & A199;
  assign \new_[78575]_  = A203 & A201;
  assign \new_[78576]_  = \new_[78575]_  & \new_[78572]_ ;
  assign \new_[78577]_  = \new_[78576]_  & \new_[78569]_ ;
  assign \new_[78580]_  = ~A234 & ~A233;
  assign \new_[78583]_  = ~A267 & ~A266;
  assign \new_[78584]_  = \new_[78583]_  & \new_[78580]_ ;
  assign \new_[78587]_  = ~A299 & A298;
  assign \new_[78590]_  = A302 & A300;
  assign \new_[78591]_  = \new_[78590]_  & \new_[78587]_ ;
  assign \new_[78592]_  = \new_[78591]_  & \new_[78584]_ ;
  assign \new_[78595]_  = ~A168 & A169;
  assign \new_[78598]_  = A166 & ~A167;
  assign \new_[78599]_  = \new_[78598]_  & \new_[78595]_ ;
  assign \new_[78602]_  = ~A200 & A199;
  assign \new_[78605]_  = A203 & A201;
  assign \new_[78606]_  = \new_[78605]_  & \new_[78602]_ ;
  assign \new_[78607]_  = \new_[78606]_  & \new_[78599]_ ;
  assign \new_[78610]_  = ~A234 & ~A233;
  assign \new_[78613]_  = ~A266 & ~A265;
  assign \new_[78614]_  = \new_[78613]_  & \new_[78610]_ ;
  assign \new_[78617]_  = ~A299 & A298;
  assign \new_[78620]_  = A301 & A300;
  assign \new_[78621]_  = \new_[78620]_  & \new_[78617]_ ;
  assign \new_[78622]_  = \new_[78621]_  & \new_[78614]_ ;
  assign \new_[78625]_  = ~A168 & A169;
  assign \new_[78628]_  = A166 & ~A167;
  assign \new_[78629]_  = \new_[78628]_  & \new_[78625]_ ;
  assign \new_[78632]_  = ~A200 & A199;
  assign \new_[78635]_  = A203 & A201;
  assign \new_[78636]_  = \new_[78635]_  & \new_[78632]_ ;
  assign \new_[78637]_  = \new_[78636]_  & \new_[78629]_ ;
  assign \new_[78640]_  = ~A234 & ~A233;
  assign \new_[78643]_  = ~A266 & ~A265;
  assign \new_[78644]_  = \new_[78643]_  & \new_[78640]_ ;
  assign \new_[78647]_  = ~A299 & A298;
  assign \new_[78650]_  = A302 & A300;
  assign \new_[78651]_  = \new_[78650]_  & \new_[78647]_ ;
  assign \new_[78652]_  = \new_[78651]_  & \new_[78644]_ ;
  assign \new_[78655]_  = ~A168 & A169;
  assign \new_[78658]_  = A166 & ~A167;
  assign \new_[78659]_  = \new_[78658]_  & \new_[78655]_ ;
  assign \new_[78662]_  = ~A200 & A199;
  assign \new_[78665]_  = A203 & A201;
  assign \new_[78666]_  = \new_[78665]_  & \new_[78662]_ ;
  assign \new_[78667]_  = \new_[78666]_  & \new_[78659]_ ;
  assign \new_[78670]_  = ~A233 & A232;
  assign \new_[78673]_  = A235 & A234;
  assign \new_[78674]_  = \new_[78673]_  & \new_[78670]_ ;
  assign \new_[78677]_  = ~A266 & A265;
  assign \new_[78680]_  = A268 & A267;
  assign \new_[78681]_  = \new_[78680]_  & \new_[78677]_ ;
  assign \new_[78682]_  = \new_[78681]_  & \new_[78674]_ ;
  assign \new_[78685]_  = ~A168 & A169;
  assign \new_[78688]_  = A166 & ~A167;
  assign \new_[78689]_  = \new_[78688]_  & \new_[78685]_ ;
  assign \new_[78692]_  = ~A200 & A199;
  assign \new_[78695]_  = A203 & A201;
  assign \new_[78696]_  = \new_[78695]_  & \new_[78692]_ ;
  assign \new_[78697]_  = \new_[78696]_  & \new_[78689]_ ;
  assign \new_[78700]_  = ~A233 & A232;
  assign \new_[78703]_  = A235 & A234;
  assign \new_[78704]_  = \new_[78703]_  & \new_[78700]_ ;
  assign \new_[78707]_  = ~A266 & A265;
  assign \new_[78710]_  = A269 & A267;
  assign \new_[78711]_  = \new_[78710]_  & \new_[78707]_ ;
  assign \new_[78712]_  = \new_[78711]_  & \new_[78704]_ ;
  assign \new_[78715]_  = ~A168 & A169;
  assign \new_[78718]_  = A166 & ~A167;
  assign \new_[78719]_  = \new_[78718]_  & \new_[78715]_ ;
  assign \new_[78722]_  = ~A200 & A199;
  assign \new_[78725]_  = A203 & A201;
  assign \new_[78726]_  = \new_[78725]_  & \new_[78722]_ ;
  assign \new_[78727]_  = \new_[78726]_  & \new_[78719]_ ;
  assign \new_[78730]_  = ~A233 & A232;
  assign \new_[78733]_  = A236 & A234;
  assign \new_[78734]_  = \new_[78733]_  & \new_[78730]_ ;
  assign \new_[78737]_  = ~A266 & A265;
  assign \new_[78740]_  = A268 & A267;
  assign \new_[78741]_  = \new_[78740]_  & \new_[78737]_ ;
  assign \new_[78742]_  = \new_[78741]_  & \new_[78734]_ ;
  assign \new_[78745]_  = ~A168 & A169;
  assign \new_[78748]_  = A166 & ~A167;
  assign \new_[78749]_  = \new_[78748]_  & \new_[78745]_ ;
  assign \new_[78752]_  = ~A200 & A199;
  assign \new_[78755]_  = A203 & A201;
  assign \new_[78756]_  = \new_[78755]_  & \new_[78752]_ ;
  assign \new_[78757]_  = \new_[78756]_  & \new_[78749]_ ;
  assign \new_[78760]_  = ~A233 & A232;
  assign \new_[78763]_  = A236 & A234;
  assign \new_[78764]_  = \new_[78763]_  & \new_[78760]_ ;
  assign \new_[78767]_  = ~A266 & A265;
  assign \new_[78770]_  = A269 & A267;
  assign \new_[78771]_  = \new_[78770]_  & \new_[78767]_ ;
  assign \new_[78772]_  = \new_[78771]_  & \new_[78764]_ ;
  assign \new_[78775]_  = ~A168 & A169;
  assign \new_[78778]_  = A166 & ~A167;
  assign \new_[78779]_  = \new_[78778]_  & \new_[78775]_ ;
  assign \new_[78782]_  = ~A200 & A199;
  assign \new_[78785]_  = A203 & A201;
  assign \new_[78786]_  = \new_[78785]_  & \new_[78782]_ ;
  assign \new_[78787]_  = \new_[78786]_  & \new_[78779]_ ;
  assign \new_[78790]_  = ~A233 & ~A232;
  assign \new_[78793]_  = A266 & A265;
  assign \new_[78794]_  = \new_[78793]_  & \new_[78790]_ ;
  assign \new_[78797]_  = ~A299 & A298;
  assign \new_[78800]_  = A301 & A300;
  assign \new_[78801]_  = \new_[78800]_  & \new_[78797]_ ;
  assign \new_[78802]_  = \new_[78801]_  & \new_[78794]_ ;
  assign \new_[78805]_  = ~A168 & A169;
  assign \new_[78808]_  = A166 & ~A167;
  assign \new_[78809]_  = \new_[78808]_  & \new_[78805]_ ;
  assign \new_[78812]_  = ~A200 & A199;
  assign \new_[78815]_  = A203 & A201;
  assign \new_[78816]_  = \new_[78815]_  & \new_[78812]_ ;
  assign \new_[78817]_  = \new_[78816]_  & \new_[78809]_ ;
  assign \new_[78820]_  = ~A233 & ~A232;
  assign \new_[78823]_  = A266 & A265;
  assign \new_[78824]_  = \new_[78823]_  & \new_[78820]_ ;
  assign \new_[78827]_  = ~A299 & A298;
  assign \new_[78830]_  = A302 & A300;
  assign \new_[78831]_  = \new_[78830]_  & \new_[78827]_ ;
  assign \new_[78832]_  = \new_[78831]_  & \new_[78824]_ ;
  assign \new_[78835]_  = ~A168 & A169;
  assign \new_[78838]_  = A166 & ~A167;
  assign \new_[78839]_  = \new_[78838]_  & \new_[78835]_ ;
  assign \new_[78842]_  = ~A200 & A199;
  assign \new_[78845]_  = A203 & A201;
  assign \new_[78846]_  = \new_[78845]_  & \new_[78842]_ ;
  assign \new_[78847]_  = \new_[78846]_  & \new_[78839]_ ;
  assign \new_[78850]_  = ~A233 & ~A232;
  assign \new_[78853]_  = ~A267 & ~A266;
  assign \new_[78854]_  = \new_[78853]_  & \new_[78850]_ ;
  assign \new_[78857]_  = ~A299 & A298;
  assign \new_[78860]_  = A301 & A300;
  assign \new_[78861]_  = \new_[78860]_  & \new_[78857]_ ;
  assign \new_[78862]_  = \new_[78861]_  & \new_[78854]_ ;
  assign \new_[78865]_  = ~A168 & A169;
  assign \new_[78868]_  = A166 & ~A167;
  assign \new_[78869]_  = \new_[78868]_  & \new_[78865]_ ;
  assign \new_[78872]_  = ~A200 & A199;
  assign \new_[78875]_  = A203 & A201;
  assign \new_[78876]_  = \new_[78875]_  & \new_[78872]_ ;
  assign \new_[78877]_  = \new_[78876]_  & \new_[78869]_ ;
  assign \new_[78880]_  = ~A233 & ~A232;
  assign \new_[78883]_  = ~A267 & ~A266;
  assign \new_[78884]_  = \new_[78883]_  & \new_[78880]_ ;
  assign \new_[78887]_  = ~A299 & A298;
  assign \new_[78890]_  = A302 & A300;
  assign \new_[78891]_  = \new_[78890]_  & \new_[78887]_ ;
  assign \new_[78892]_  = \new_[78891]_  & \new_[78884]_ ;
  assign \new_[78895]_  = ~A168 & A169;
  assign \new_[78898]_  = A166 & ~A167;
  assign \new_[78899]_  = \new_[78898]_  & \new_[78895]_ ;
  assign \new_[78902]_  = ~A200 & A199;
  assign \new_[78905]_  = A203 & A201;
  assign \new_[78906]_  = \new_[78905]_  & \new_[78902]_ ;
  assign \new_[78907]_  = \new_[78906]_  & \new_[78899]_ ;
  assign \new_[78910]_  = ~A233 & ~A232;
  assign \new_[78913]_  = ~A266 & ~A265;
  assign \new_[78914]_  = \new_[78913]_  & \new_[78910]_ ;
  assign \new_[78917]_  = ~A299 & A298;
  assign \new_[78920]_  = A301 & A300;
  assign \new_[78921]_  = \new_[78920]_  & \new_[78917]_ ;
  assign \new_[78922]_  = \new_[78921]_  & \new_[78914]_ ;
  assign \new_[78925]_  = ~A168 & A169;
  assign \new_[78928]_  = A166 & ~A167;
  assign \new_[78929]_  = \new_[78928]_  & \new_[78925]_ ;
  assign \new_[78932]_  = ~A200 & A199;
  assign \new_[78935]_  = A203 & A201;
  assign \new_[78936]_  = \new_[78935]_  & \new_[78932]_ ;
  assign \new_[78937]_  = \new_[78936]_  & \new_[78929]_ ;
  assign \new_[78940]_  = ~A233 & ~A232;
  assign \new_[78943]_  = ~A266 & ~A265;
  assign \new_[78944]_  = \new_[78943]_  & \new_[78940]_ ;
  assign \new_[78947]_  = ~A299 & A298;
  assign \new_[78950]_  = A302 & A300;
  assign \new_[78951]_  = \new_[78950]_  & \new_[78947]_ ;
  assign \new_[78952]_  = \new_[78951]_  & \new_[78944]_ ;
  assign \new_[78955]_  = A169 & A170;
  assign \new_[78958]_  = A199 & ~A168;
  assign \new_[78959]_  = \new_[78958]_  & \new_[78955]_ ;
  assign \new_[78962]_  = A201 & ~A200;
  assign \new_[78965]_  = A232 & A202;
  assign \new_[78966]_  = \new_[78965]_  & \new_[78962]_ ;
  assign \new_[78967]_  = \new_[78966]_  & \new_[78959]_ ;
  assign \new_[78970]_  = A265 & A233;
  assign \new_[78973]_  = ~A269 & ~A268;
  assign \new_[78974]_  = \new_[78973]_  & \new_[78970]_ ;
  assign \new_[78977]_  = ~A299 & A298;
  assign \new_[78980]_  = A301 & A300;
  assign \new_[78981]_  = \new_[78980]_  & \new_[78977]_ ;
  assign \new_[78982]_  = \new_[78981]_  & \new_[78974]_ ;
  assign \new_[78985]_  = A169 & A170;
  assign \new_[78988]_  = A199 & ~A168;
  assign \new_[78989]_  = \new_[78988]_  & \new_[78985]_ ;
  assign \new_[78992]_  = A201 & ~A200;
  assign \new_[78995]_  = A232 & A202;
  assign \new_[78996]_  = \new_[78995]_  & \new_[78992]_ ;
  assign \new_[78997]_  = \new_[78996]_  & \new_[78989]_ ;
  assign \new_[79000]_  = A265 & A233;
  assign \new_[79003]_  = ~A269 & ~A268;
  assign \new_[79004]_  = \new_[79003]_  & \new_[79000]_ ;
  assign \new_[79007]_  = ~A299 & A298;
  assign \new_[79010]_  = A302 & A300;
  assign \new_[79011]_  = \new_[79010]_  & \new_[79007]_ ;
  assign \new_[79012]_  = \new_[79011]_  & \new_[79004]_ ;
  assign \new_[79015]_  = A169 & A170;
  assign \new_[79018]_  = A199 & ~A168;
  assign \new_[79019]_  = \new_[79018]_  & \new_[79015]_ ;
  assign \new_[79022]_  = A201 & ~A200;
  assign \new_[79025]_  = ~A233 & A202;
  assign \new_[79026]_  = \new_[79025]_  & \new_[79022]_ ;
  assign \new_[79027]_  = \new_[79026]_  & \new_[79019]_ ;
  assign \new_[79030]_  = ~A236 & ~A235;
  assign \new_[79033]_  = A266 & A265;
  assign \new_[79034]_  = \new_[79033]_  & \new_[79030]_ ;
  assign \new_[79037]_  = ~A299 & A298;
  assign \new_[79040]_  = A301 & A300;
  assign \new_[79041]_  = \new_[79040]_  & \new_[79037]_ ;
  assign \new_[79042]_  = \new_[79041]_  & \new_[79034]_ ;
  assign \new_[79045]_  = A169 & A170;
  assign \new_[79048]_  = A199 & ~A168;
  assign \new_[79049]_  = \new_[79048]_  & \new_[79045]_ ;
  assign \new_[79052]_  = A201 & ~A200;
  assign \new_[79055]_  = ~A233 & A202;
  assign \new_[79056]_  = \new_[79055]_  & \new_[79052]_ ;
  assign \new_[79057]_  = \new_[79056]_  & \new_[79049]_ ;
  assign \new_[79060]_  = ~A236 & ~A235;
  assign \new_[79063]_  = A266 & A265;
  assign \new_[79064]_  = \new_[79063]_  & \new_[79060]_ ;
  assign \new_[79067]_  = ~A299 & A298;
  assign \new_[79070]_  = A302 & A300;
  assign \new_[79071]_  = \new_[79070]_  & \new_[79067]_ ;
  assign \new_[79072]_  = \new_[79071]_  & \new_[79064]_ ;
  assign \new_[79075]_  = A169 & A170;
  assign \new_[79078]_  = A199 & ~A168;
  assign \new_[79079]_  = \new_[79078]_  & \new_[79075]_ ;
  assign \new_[79082]_  = A201 & ~A200;
  assign \new_[79085]_  = ~A233 & A202;
  assign \new_[79086]_  = \new_[79085]_  & \new_[79082]_ ;
  assign \new_[79087]_  = \new_[79086]_  & \new_[79079]_ ;
  assign \new_[79090]_  = ~A236 & ~A235;
  assign \new_[79093]_  = ~A267 & ~A266;
  assign \new_[79094]_  = \new_[79093]_  & \new_[79090]_ ;
  assign \new_[79097]_  = ~A299 & A298;
  assign \new_[79100]_  = A301 & A300;
  assign \new_[79101]_  = \new_[79100]_  & \new_[79097]_ ;
  assign \new_[79102]_  = \new_[79101]_  & \new_[79094]_ ;
  assign \new_[79105]_  = A169 & A170;
  assign \new_[79108]_  = A199 & ~A168;
  assign \new_[79109]_  = \new_[79108]_  & \new_[79105]_ ;
  assign \new_[79112]_  = A201 & ~A200;
  assign \new_[79115]_  = ~A233 & A202;
  assign \new_[79116]_  = \new_[79115]_  & \new_[79112]_ ;
  assign \new_[79117]_  = \new_[79116]_  & \new_[79109]_ ;
  assign \new_[79120]_  = ~A236 & ~A235;
  assign \new_[79123]_  = ~A267 & ~A266;
  assign \new_[79124]_  = \new_[79123]_  & \new_[79120]_ ;
  assign \new_[79127]_  = ~A299 & A298;
  assign \new_[79130]_  = A302 & A300;
  assign \new_[79131]_  = \new_[79130]_  & \new_[79127]_ ;
  assign \new_[79132]_  = \new_[79131]_  & \new_[79124]_ ;
  assign \new_[79135]_  = A169 & A170;
  assign \new_[79138]_  = A199 & ~A168;
  assign \new_[79139]_  = \new_[79138]_  & \new_[79135]_ ;
  assign \new_[79142]_  = A201 & ~A200;
  assign \new_[79145]_  = ~A233 & A202;
  assign \new_[79146]_  = \new_[79145]_  & \new_[79142]_ ;
  assign \new_[79147]_  = \new_[79146]_  & \new_[79139]_ ;
  assign \new_[79150]_  = ~A236 & ~A235;
  assign \new_[79153]_  = ~A266 & ~A265;
  assign \new_[79154]_  = \new_[79153]_  & \new_[79150]_ ;
  assign \new_[79157]_  = ~A299 & A298;
  assign \new_[79160]_  = A301 & A300;
  assign \new_[79161]_  = \new_[79160]_  & \new_[79157]_ ;
  assign \new_[79162]_  = \new_[79161]_  & \new_[79154]_ ;
  assign \new_[79165]_  = A169 & A170;
  assign \new_[79168]_  = A199 & ~A168;
  assign \new_[79169]_  = \new_[79168]_  & \new_[79165]_ ;
  assign \new_[79172]_  = A201 & ~A200;
  assign \new_[79175]_  = ~A233 & A202;
  assign \new_[79176]_  = \new_[79175]_  & \new_[79172]_ ;
  assign \new_[79177]_  = \new_[79176]_  & \new_[79169]_ ;
  assign \new_[79180]_  = ~A236 & ~A235;
  assign \new_[79183]_  = ~A266 & ~A265;
  assign \new_[79184]_  = \new_[79183]_  & \new_[79180]_ ;
  assign \new_[79187]_  = ~A299 & A298;
  assign \new_[79190]_  = A302 & A300;
  assign \new_[79191]_  = \new_[79190]_  & \new_[79187]_ ;
  assign \new_[79192]_  = \new_[79191]_  & \new_[79184]_ ;
  assign \new_[79195]_  = A169 & A170;
  assign \new_[79198]_  = A199 & ~A168;
  assign \new_[79199]_  = \new_[79198]_  & \new_[79195]_ ;
  assign \new_[79202]_  = A201 & ~A200;
  assign \new_[79205]_  = A232 & A203;
  assign \new_[79206]_  = \new_[79205]_  & \new_[79202]_ ;
  assign \new_[79207]_  = \new_[79206]_  & \new_[79199]_ ;
  assign \new_[79210]_  = A265 & A233;
  assign \new_[79213]_  = ~A269 & ~A268;
  assign \new_[79214]_  = \new_[79213]_  & \new_[79210]_ ;
  assign \new_[79217]_  = ~A299 & A298;
  assign \new_[79220]_  = A301 & A300;
  assign \new_[79221]_  = \new_[79220]_  & \new_[79217]_ ;
  assign \new_[79222]_  = \new_[79221]_  & \new_[79214]_ ;
  assign \new_[79225]_  = A169 & A170;
  assign \new_[79228]_  = A199 & ~A168;
  assign \new_[79229]_  = \new_[79228]_  & \new_[79225]_ ;
  assign \new_[79232]_  = A201 & ~A200;
  assign \new_[79235]_  = A232 & A203;
  assign \new_[79236]_  = \new_[79235]_  & \new_[79232]_ ;
  assign \new_[79237]_  = \new_[79236]_  & \new_[79229]_ ;
  assign \new_[79240]_  = A265 & A233;
  assign \new_[79243]_  = ~A269 & ~A268;
  assign \new_[79244]_  = \new_[79243]_  & \new_[79240]_ ;
  assign \new_[79247]_  = ~A299 & A298;
  assign \new_[79250]_  = A302 & A300;
  assign \new_[79251]_  = \new_[79250]_  & \new_[79247]_ ;
  assign \new_[79252]_  = \new_[79251]_  & \new_[79244]_ ;
  assign \new_[79255]_  = A169 & A170;
  assign \new_[79258]_  = A199 & ~A168;
  assign \new_[79259]_  = \new_[79258]_  & \new_[79255]_ ;
  assign \new_[79262]_  = A201 & ~A200;
  assign \new_[79265]_  = ~A233 & A203;
  assign \new_[79266]_  = \new_[79265]_  & \new_[79262]_ ;
  assign \new_[79267]_  = \new_[79266]_  & \new_[79259]_ ;
  assign \new_[79270]_  = ~A236 & ~A235;
  assign \new_[79273]_  = A266 & A265;
  assign \new_[79274]_  = \new_[79273]_  & \new_[79270]_ ;
  assign \new_[79277]_  = ~A299 & A298;
  assign \new_[79280]_  = A301 & A300;
  assign \new_[79281]_  = \new_[79280]_  & \new_[79277]_ ;
  assign \new_[79282]_  = \new_[79281]_  & \new_[79274]_ ;
  assign \new_[79285]_  = A169 & A170;
  assign \new_[79288]_  = A199 & ~A168;
  assign \new_[79289]_  = \new_[79288]_  & \new_[79285]_ ;
  assign \new_[79292]_  = A201 & ~A200;
  assign \new_[79295]_  = ~A233 & A203;
  assign \new_[79296]_  = \new_[79295]_  & \new_[79292]_ ;
  assign \new_[79297]_  = \new_[79296]_  & \new_[79289]_ ;
  assign \new_[79300]_  = ~A236 & ~A235;
  assign \new_[79303]_  = A266 & A265;
  assign \new_[79304]_  = \new_[79303]_  & \new_[79300]_ ;
  assign \new_[79307]_  = ~A299 & A298;
  assign \new_[79310]_  = A302 & A300;
  assign \new_[79311]_  = \new_[79310]_  & \new_[79307]_ ;
  assign \new_[79312]_  = \new_[79311]_  & \new_[79304]_ ;
  assign \new_[79315]_  = A169 & A170;
  assign \new_[79318]_  = A199 & ~A168;
  assign \new_[79319]_  = \new_[79318]_  & \new_[79315]_ ;
  assign \new_[79322]_  = A201 & ~A200;
  assign \new_[79325]_  = ~A233 & A203;
  assign \new_[79326]_  = \new_[79325]_  & \new_[79322]_ ;
  assign \new_[79327]_  = \new_[79326]_  & \new_[79319]_ ;
  assign \new_[79330]_  = ~A236 & ~A235;
  assign \new_[79333]_  = ~A267 & ~A266;
  assign \new_[79334]_  = \new_[79333]_  & \new_[79330]_ ;
  assign \new_[79337]_  = ~A299 & A298;
  assign \new_[79340]_  = A301 & A300;
  assign \new_[79341]_  = \new_[79340]_  & \new_[79337]_ ;
  assign \new_[79342]_  = \new_[79341]_  & \new_[79334]_ ;
  assign \new_[79345]_  = A169 & A170;
  assign \new_[79348]_  = A199 & ~A168;
  assign \new_[79349]_  = \new_[79348]_  & \new_[79345]_ ;
  assign \new_[79352]_  = A201 & ~A200;
  assign \new_[79355]_  = ~A233 & A203;
  assign \new_[79356]_  = \new_[79355]_  & \new_[79352]_ ;
  assign \new_[79357]_  = \new_[79356]_  & \new_[79349]_ ;
  assign \new_[79360]_  = ~A236 & ~A235;
  assign \new_[79363]_  = ~A267 & ~A266;
  assign \new_[79364]_  = \new_[79363]_  & \new_[79360]_ ;
  assign \new_[79367]_  = ~A299 & A298;
  assign \new_[79370]_  = A302 & A300;
  assign \new_[79371]_  = \new_[79370]_  & \new_[79367]_ ;
  assign \new_[79372]_  = \new_[79371]_  & \new_[79364]_ ;
  assign \new_[79375]_  = A169 & A170;
  assign \new_[79378]_  = A199 & ~A168;
  assign \new_[79379]_  = \new_[79378]_  & \new_[79375]_ ;
  assign \new_[79382]_  = A201 & ~A200;
  assign \new_[79385]_  = ~A233 & A203;
  assign \new_[79386]_  = \new_[79385]_  & \new_[79382]_ ;
  assign \new_[79387]_  = \new_[79386]_  & \new_[79379]_ ;
  assign \new_[79390]_  = ~A236 & ~A235;
  assign \new_[79393]_  = ~A266 & ~A265;
  assign \new_[79394]_  = \new_[79393]_  & \new_[79390]_ ;
  assign \new_[79397]_  = ~A299 & A298;
  assign \new_[79400]_  = A301 & A300;
  assign \new_[79401]_  = \new_[79400]_  & \new_[79397]_ ;
  assign \new_[79402]_  = \new_[79401]_  & \new_[79394]_ ;
  assign \new_[79405]_  = A169 & A170;
  assign \new_[79408]_  = A199 & ~A168;
  assign \new_[79409]_  = \new_[79408]_  & \new_[79405]_ ;
  assign \new_[79412]_  = A201 & ~A200;
  assign \new_[79415]_  = ~A233 & A203;
  assign \new_[79416]_  = \new_[79415]_  & \new_[79412]_ ;
  assign \new_[79417]_  = \new_[79416]_  & \new_[79409]_ ;
  assign \new_[79420]_  = ~A236 & ~A235;
  assign \new_[79423]_  = ~A266 & ~A265;
  assign \new_[79424]_  = \new_[79423]_  & \new_[79420]_ ;
  assign \new_[79427]_  = ~A299 & A298;
  assign \new_[79430]_  = A302 & A300;
  assign \new_[79431]_  = \new_[79430]_  & \new_[79427]_ ;
  assign \new_[79432]_  = \new_[79431]_  & \new_[79424]_ ;
  assign \new_[79435]_  = A169 & A170;
  assign \new_[79438]_  = A166 & ~A168;
  assign \new_[79439]_  = \new_[79438]_  & \new_[79435]_ ;
  assign \new_[79442]_  = ~A200 & A199;
  assign \new_[79445]_  = A202 & A201;
  assign \new_[79446]_  = \new_[79445]_  & \new_[79442]_ ;
  assign \new_[79447]_  = \new_[79446]_  & \new_[79439]_ ;
  assign \new_[79450]_  = ~A234 & ~A233;
  assign \new_[79453]_  = ~A267 & ~A266;
  assign \new_[79454]_  = \new_[79453]_  & \new_[79450]_ ;
  assign \new_[79457]_  = ~A299 & A298;
  assign \new_[79460]_  = A301 & A300;
  assign \new_[79461]_  = \new_[79460]_  & \new_[79457]_ ;
  assign \new_[79462]_  = \new_[79461]_  & \new_[79454]_ ;
  assign \new_[79465]_  = A169 & A170;
  assign \new_[79468]_  = A166 & ~A168;
  assign \new_[79469]_  = \new_[79468]_  & \new_[79465]_ ;
  assign \new_[79472]_  = ~A200 & A199;
  assign \new_[79475]_  = A202 & A201;
  assign \new_[79476]_  = \new_[79475]_  & \new_[79472]_ ;
  assign \new_[79477]_  = \new_[79476]_  & \new_[79469]_ ;
  assign \new_[79480]_  = ~A234 & ~A233;
  assign \new_[79483]_  = ~A267 & ~A266;
  assign \new_[79484]_  = \new_[79483]_  & \new_[79480]_ ;
  assign \new_[79487]_  = ~A299 & A298;
  assign \new_[79490]_  = A302 & A300;
  assign \new_[79491]_  = \new_[79490]_  & \new_[79487]_ ;
  assign \new_[79492]_  = \new_[79491]_  & \new_[79484]_ ;
  assign \new_[79495]_  = A169 & A170;
  assign \new_[79498]_  = A166 & ~A168;
  assign \new_[79499]_  = \new_[79498]_  & \new_[79495]_ ;
  assign \new_[79502]_  = ~A200 & A199;
  assign \new_[79505]_  = A202 & A201;
  assign \new_[79506]_  = \new_[79505]_  & \new_[79502]_ ;
  assign \new_[79507]_  = \new_[79506]_  & \new_[79499]_ ;
  assign \new_[79510]_  = ~A234 & ~A233;
  assign \new_[79513]_  = ~A266 & ~A265;
  assign \new_[79514]_  = \new_[79513]_  & \new_[79510]_ ;
  assign \new_[79517]_  = ~A299 & A298;
  assign \new_[79520]_  = A301 & A300;
  assign \new_[79521]_  = \new_[79520]_  & \new_[79517]_ ;
  assign \new_[79522]_  = \new_[79521]_  & \new_[79514]_ ;
  assign \new_[79525]_  = A169 & A170;
  assign \new_[79528]_  = A166 & ~A168;
  assign \new_[79529]_  = \new_[79528]_  & \new_[79525]_ ;
  assign \new_[79532]_  = ~A200 & A199;
  assign \new_[79535]_  = A202 & A201;
  assign \new_[79536]_  = \new_[79535]_  & \new_[79532]_ ;
  assign \new_[79537]_  = \new_[79536]_  & \new_[79529]_ ;
  assign \new_[79540]_  = ~A234 & ~A233;
  assign \new_[79543]_  = ~A266 & ~A265;
  assign \new_[79544]_  = \new_[79543]_  & \new_[79540]_ ;
  assign \new_[79547]_  = ~A299 & A298;
  assign \new_[79550]_  = A302 & A300;
  assign \new_[79551]_  = \new_[79550]_  & \new_[79547]_ ;
  assign \new_[79552]_  = \new_[79551]_  & \new_[79544]_ ;
  assign \new_[79555]_  = A169 & A170;
  assign \new_[79558]_  = A166 & ~A168;
  assign \new_[79559]_  = \new_[79558]_  & \new_[79555]_ ;
  assign \new_[79562]_  = ~A200 & A199;
  assign \new_[79565]_  = A202 & A201;
  assign \new_[79566]_  = \new_[79565]_  & \new_[79562]_ ;
  assign \new_[79567]_  = \new_[79566]_  & \new_[79559]_ ;
  assign \new_[79570]_  = ~A233 & ~A232;
  assign \new_[79573]_  = ~A267 & ~A266;
  assign \new_[79574]_  = \new_[79573]_  & \new_[79570]_ ;
  assign \new_[79577]_  = ~A299 & A298;
  assign \new_[79580]_  = A301 & A300;
  assign \new_[79581]_  = \new_[79580]_  & \new_[79577]_ ;
  assign \new_[79582]_  = \new_[79581]_  & \new_[79574]_ ;
  assign \new_[79585]_  = A169 & A170;
  assign \new_[79588]_  = A166 & ~A168;
  assign \new_[79589]_  = \new_[79588]_  & \new_[79585]_ ;
  assign \new_[79592]_  = ~A200 & A199;
  assign \new_[79595]_  = A202 & A201;
  assign \new_[79596]_  = \new_[79595]_  & \new_[79592]_ ;
  assign \new_[79597]_  = \new_[79596]_  & \new_[79589]_ ;
  assign \new_[79600]_  = ~A233 & ~A232;
  assign \new_[79603]_  = ~A267 & ~A266;
  assign \new_[79604]_  = \new_[79603]_  & \new_[79600]_ ;
  assign \new_[79607]_  = ~A299 & A298;
  assign \new_[79610]_  = A302 & A300;
  assign \new_[79611]_  = \new_[79610]_  & \new_[79607]_ ;
  assign \new_[79612]_  = \new_[79611]_  & \new_[79604]_ ;
  assign \new_[79615]_  = A169 & A170;
  assign \new_[79618]_  = A166 & ~A168;
  assign \new_[79619]_  = \new_[79618]_  & \new_[79615]_ ;
  assign \new_[79622]_  = ~A200 & A199;
  assign \new_[79625]_  = A202 & A201;
  assign \new_[79626]_  = \new_[79625]_  & \new_[79622]_ ;
  assign \new_[79627]_  = \new_[79626]_  & \new_[79619]_ ;
  assign \new_[79630]_  = ~A233 & ~A232;
  assign \new_[79633]_  = ~A266 & ~A265;
  assign \new_[79634]_  = \new_[79633]_  & \new_[79630]_ ;
  assign \new_[79637]_  = ~A299 & A298;
  assign \new_[79640]_  = A301 & A300;
  assign \new_[79641]_  = \new_[79640]_  & \new_[79637]_ ;
  assign \new_[79642]_  = \new_[79641]_  & \new_[79634]_ ;
  assign \new_[79645]_  = A169 & A170;
  assign \new_[79648]_  = A166 & ~A168;
  assign \new_[79649]_  = \new_[79648]_  & \new_[79645]_ ;
  assign \new_[79652]_  = ~A200 & A199;
  assign \new_[79655]_  = A202 & A201;
  assign \new_[79656]_  = \new_[79655]_  & \new_[79652]_ ;
  assign \new_[79657]_  = \new_[79656]_  & \new_[79649]_ ;
  assign \new_[79660]_  = ~A233 & ~A232;
  assign \new_[79663]_  = ~A266 & ~A265;
  assign \new_[79664]_  = \new_[79663]_  & \new_[79660]_ ;
  assign \new_[79667]_  = ~A299 & A298;
  assign \new_[79670]_  = A302 & A300;
  assign \new_[79671]_  = \new_[79670]_  & \new_[79667]_ ;
  assign \new_[79672]_  = \new_[79671]_  & \new_[79664]_ ;
  assign \new_[79675]_  = A169 & A170;
  assign \new_[79678]_  = A166 & ~A168;
  assign \new_[79679]_  = \new_[79678]_  & \new_[79675]_ ;
  assign \new_[79682]_  = ~A200 & A199;
  assign \new_[79685]_  = A203 & A201;
  assign \new_[79686]_  = \new_[79685]_  & \new_[79682]_ ;
  assign \new_[79687]_  = \new_[79686]_  & \new_[79679]_ ;
  assign \new_[79690]_  = ~A234 & ~A233;
  assign \new_[79693]_  = ~A267 & ~A266;
  assign \new_[79694]_  = \new_[79693]_  & \new_[79690]_ ;
  assign \new_[79697]_  = ~A299 & A298;
  assign \new_[79700]_  = A301 & A300;
  assign \new_[79701]_  = \new_[79700]_  & \new_[79697]_ ;
  assign \new_[79702]_  = \new_[79701]_  & \new_[79694]_ ;
  assign \new_[79705]_  = A169 & A170;
  assign \new_[79708]_  = A166 & ~A168;
  assign \new_[79709]_  = \new_[79708]_  & \new_[79705]_ ;
  assign \new_[79712]_  = ~A200 & A199;
  assign \new_[79715]_  = A203 & A201;
  assign \new_[79716]_  = \new_[79715]_  & \new_[79712]_ ;
  assign \new_[79717]_  = \new_[79716]_  & \new_[79709]_ ;
  assign \new_[79720]_  = ~A234 & ~A233;
  assign \new_[79723]_  = ~A267 & ~A266;
  assign \new_[79724]_  = \new_[79723]_  & \new_[79720]_ ;
  assign \new_[79727]_  = ~A299 & A298;
  assign \new_[79730]_  = A302 & A300;
  assign \new_[79731]_  = \new_[79730]_  & \new_[79727]_ ;
  assign \new_[79732]_  = \new_[79731]_  & \new_[79724]_ ;
  assign \new_[79735]_  = A169 & A170;
  assign \new_[79738]_  = A166 & ~A168;
  assign \new_[79739]_  = \new_[79738]_  & \new_[79735]_ ;
  assign \new_[79742]_  = ~A200 & A199;
  assign \new_[79745]_  = A203 & A201;
  assign \new_[79746]_  = \new_[79745]_  & \new_[79742]_ ;
  assign \new_[79747]_  = \new_[79746]_  & \new_[79739]_ ;
  assign \new_[79750]_  = ~A234 & ~A233;
  assign \new_[79753]_  = ~A266 & ~A265;
  assign \new_[79754]_  = \new_[79753]_  & \new_[79750]_ ;
  assign \new_[79757]_  = ~A299 & A298;
  assign \new_[79760]_  = A301 & A300;
  assign \new_[79761]_  = \new_[79760]_  & \new_[79757]_ ;
  assign \new_[79762]_  = \new_[79761]_  & \new_[79754]_ ;
  assign \new_[79765]_  = A169 & A170;
  assign \new_[79768]_  = A166 & ~A168;
  assign \new_[79769]_  = \new_[79768]_  & \new_[79765]_ ;
  assign \new_[79772]_  = ~A200 & A199;
  assign \new_[79775]_  = A203 & A201;
  assign \new_[79776]_  = \new_[79775]_  & \new_[79772]_ ;
  assign \new_[79777]_  = \new_[79776]_  & \new_[79769]_ ;
  assign \new_[79780]_  = ~A234 & ~A233;
  assign \new_[79783]_  = ~A266 & ~A265;
  assign \new_[79784]_  = \new_[79783]_  & \new_[79780]_ ;
  assign \new_[79787]_  = ~A299 & A298;
  assign \new_[79790]_  = A302 & A300;
  assign \new_[79791]_  = \new_[79790]_  & \new_[79787]_ ;
  assign \new_[79792]_  = \new_[79791]_  & \new_[79784]_ ;
  assign \new_[79795]_  = A169 & A170;
  assign \new_[79798]_  = A166 & ~A168;
  assign \new_[79799]_  = \new_[79798]_  & \new_[79795]_ ;
  assign \new_[79802]_  = ~A200 & A199;
  assign \new_[79805]_  = A203 & A201;
  assign \new_[79806]_  = \new_[79805]_  & \new_[79802]_ ;
  assign \new_[79807]_  = \new_[79806]_  & \new_[79799]_ ;
  assign \new_[79810]_  = ~A233 & ~A232;
  assign \new_[79813]_  = ~A267 & ~A266;
  assign \new_[79814]_  = \new_[79813]_  & \new_[79810]_ ;
  assign \new_[79817]_  = ~A299 & A298;
  assign \new_[79820]_  = A301 & A300;
  assign \new_[79821]_  = \new_[79820]_  & \new_[79817]_ ;
  assign \new_[79822]_  = \new_[79821]_  & \new_[79814]_ ;
  assign \new_[79825]_  = A169 & A170;
  assign \new_[79828]_  = A166 & ~A168;
  assign \new_[79829]_  = \new_[79828]_  & \new_[79825]_ ;
  assign \new_[79832]_  = ~A200 & A199;
  assign \new_[79835]_  = A203 & A201;
  assign \new_[79836]_  = \new_[79835]_  & \new_[79832]_ ;
  assign \new_[79837]_  = \new_[79836]_  & \new_[79829]_ ;
  assign \new_[79840]_  = ~A233 & ~A232;
  assign \new_[79843]_  = ~A267 & ~A266;
  assign \new_[79844]_  = \new_[79843]_  & \new_[79840]_ ;
  assign \new_[79847]_  = ~A299 & A298;
  assign \new_[79850]_  = A302 & A300;
  assign \new_[79851]_  = \new_[79850]_  & \new_[79847]_ ;
  assign \new_[79852]_  = \new_[79851]_  & \new_[79844]_ ;
  assign \new_[79855]_  = A169 & A170;
  assign \new_[79858]_  = A166 & ~A168;
  assign \new_[79859]_  = \new_[79858]_  & \new_[79855]_ ;
  assign \new_[79862]_  = ~A200 & A199;
  assign \new_[79865]_  = A203 & A201;
  assign \new_[79866]_  = \new_[79865]_  & \new_[79862]_ ;
  assign \new_[79867]_  = \new_[79866]_  & \new_[79859]_ ;
  assign \new_[79870]_  = ~A233 & ~A232;
  assign \new_[79873]_  = ~A266 & ~A265;
  assign \new_[79874]_  = \new_[79873]_  & \new_[79870]_ ;
  assign \new_[79877]_  = ~A299 & A298;
  assign \new_[79880]_  = A301 & A300;
  assign \new_[79881]_  = \new_[79880]_  & \new_[79877]_ ;
  assign \new_[79882]_  = \new_[79881]_  & \new_[79874]_ ;
  assign \new_[79885]_  = A169 & A170;
  assign \new_[79888]_  = A166 & ~A168;
  assign \new_[79889]_  = \new_[79888]_  & \new_[79885]_ ;
  assign \new_[79892]_  = ~A200 & A199;
  assign \new_[79895]_  = A203 & A201;
  assign \new_[79896]_  = \new_[79895]_  & \new_[79892]_ ;
  assign \new_[79897]_  = \new_[79896]_  & \new_[79889]_ ;
  assign \new_[79900]_  = ~A233 & ~A232;
  assign \new_[79903]_  = ~A266 & ~A265;
  assign \new_[79904]_  = \new_[79903]_  & \new_[79900]_ ;
  assign \new_[79907]_  = ~A299 & A298;
  assign \new_[79910]_  = A302 & A300;
  assign \new_[79911]_  = \new_[79910]_  & \new_[79907]_ ;
  assign \new_[79912]_  = \new_[79911]_  & \new_[79904]_ ;
  assign \new_[79915]_  = A169 & ~A170;
  assign \new_[79918]_  = A166 & A167;
  assign \new_[79919]_  = \new_[79918]_  & \new_[79915]_ ;
  assign \new_[79922]_  = A200 & A199;
  assign \new_[79925]_  = ~A235 & ~A233;
  assign \new_[79926]_  = \new_[79925]_  & \new_[79922]_ ;
  assign \new_[79927]_  = \new_[79926]_  & \new_[79919]_ ;
  assign \new_[79930]_  = ~A266 & ~A236;
  assign \new_[79933]_  = ~A269 & ~A268;
  assign \new_[79934]_  = \new_[79933]_  & \new_[79930]_ ;
  assign \new_[79937]_  = ~A299 & A298;
  assign \new_[79940]_  = A301 & A300;
  assign \new_[79941]_  = \new_[79940]_  & \new_[79937]_ ;
  assign \new_[79942]_  = \new_[79941]_  & \new_[79934]_ ;
  assign \new_[79945]_  = A169 & ~A170;
  assign \new_[79948]_  = A166 & A167;
  assign \new_[79949]_  = \new_[79948]_  & \new_[79945]_ ;
  assign \new_[79952]_  = A200 & A199;
  assign \new_[79955]_  = ~A235 & ~A233;
  assign \new_[79956]_  = \new_[79955]_  & \new_[79952]_ ;
  assign \new_[79957]_  = \new_[79956]_  & \new_[79949]_ ;
  assign \new_[79960]_  = ~A266 & ~A236;
  assign \new_[79963]_  = ~A269 & ~A268;
  assign \new_[79964]_  = \new_[79963]_  & \new_[79960]_ ;
  assign \new_[79967]_  = ~A299 & A298;
  assign \new_[79970]_  = A302 & A300;
  assign \new_[79971]_  = \new_[79970]_  & \new_[79967]_ ;
  assign \new_[79972]_  = \new_[79971]_  & \new_[79964]_ ;
  assign \new_[79975]_  = A169 & ~A170;
  assign \new_[79978]_  = A166 & A167;
  assign \new_[79979]_  = \new_[79978]_  & \new_[79975]_ ;
  assign \new_[79982]_  = ~A202 & ~A200;
  assign \new_[79985]_  = A232 & ~A203;
  assign \new_[79986]_  = \new_[79985]_  & \new_[79982]_ ;
  assign \new_[79987]_  = \new_[79986]_  & \new_[79979]_ ;
  assign \new_[79990]_  = A265 & A233;
  assign \new_[79993]_  = ~A269 & ~A268;
  assign \new_[79994]_  = \new_[79993]_  & \new_[79990]_ ;
  assign \new_[79997]_  = ~A299 & A298;
  assign \new_[80000]_  = A301 & A300;
  assign \new_[80001]_  = \new_[80000]_  & \new_[79997]_ ;
  assign \new_[80002]_  = \new_[80001]_  & \new_[79994]_ ;
  assign \new_[80005]_  = A169 & ~A170;
  assign \new_[80008]_  = A166 & A167;
  assign \new_[80009]_  = \new_[80008]_  & \new_[80005]_ ;
  assign \new_[80012]_  = ~A202 & ~A200;
  assign \new_[80015]_  = A232 & ~A203;
  assign \new_[80016]_  = \new_[80015]_  & \new_[80012]_ ;
  assign \new_[80017]_  = \new_[80016]_  & \new_[80009]_ ;
  assign \new_[80020]_  = A265 & A233;
  assign \new_[80023]_  = ~A269 & ~A268;
  assign \new_[80024]_  = \new_[80023]_  & \new_[80020]_ ;
  assign \new_[80027]_  = ~A299 & A298;
  assign \new_[80030]_  = A302 & A300;
  assign \new_[80031]_  = \new_[80030]_  & \new_[80027]_ ;
  assign \new_[80032]_  = \new_[80031]_  & \new_[80024]_ ;
  assign \new_[80035]_  = A169 & ~A170;
  assign \new_[80038]_  = A166 & A167;
  assign \new_[80039]_  = \new_[80038]_  & \new_[80035]_ ;
  assign \new_[80042]_  = ~A202 & ~A200;
  assign \new_[80045]_  = ~A233 & ~A203;
  assign \new_[80046]_  = \new_[80045]_  & \new_[80042]_ ;
  assign \new_[80047]_  = \new_[80046]_  & \new_[80039]_ ;
  assign \new_[80050]_  = ~A236 & ~A235;
  assign \new_[80053]_  = A266 & A265;
  assign \new_[80054]_  = \new_[80053]_  & \new_[80050]_ ;
  assign \new_[80057]_  = ~A299 & A298;
  assign \new_[80060]_  = A301 & A300;
  assign \new_[80061]_  = \new_[80060]_  & \new_[80057]_ ;
  assign \new_[80062]_  = \new_[80061]_  & \new_[80054]_ ;
  assign \new_[80065]_  = A169 & ~A170;
  assign \new_[80068]_  = A166 & A167;
  assign \new_[80069]_  = \new_[80068]_  & \new_[80065]_ ;
  assign \new_[80072]_  = ~A202 & ~A200;
  assign \new_[80075]_  = ~A233 & ~A203;
  assign \new_[80076]_  = \new_[80075]_  & \new_[80072]_ ;
  assign \new_[80077]_  = \new_[80076]_  & \new_[80069]_ ;
  assign \new_[80080]_  = ~A236 & ~A235;
  assign \new_[80083]_  = A266 & A265;
  assign \new_[80084]_  = \new_[80083]_  & \new_[80080]_ ;
  assign \new_[80087]_  = ~A299 & A298;
  assign \new_[80090]_  = A302 & A300;
  assign \new_[80091]_  = \new_[80090]_  & \new_[80087]_ ;
  assign \new_[80092]_  = \new_[80091]_  & \new_[80084]_ ;
  assign \new_[80095]_  = A169 & ~A170;
  assign \new_[80098]_  = A166 & A167;
  assign \new_[80099]_  = \new_[80098]_  & \new_[80095]_ ;
  assign \new_[80102]_  = ~A202 & ~A200;
  assign \new_[80105]_  = ~A233 & ~A203;
  assign \new_[80106]_  = \new_[80105]_  & \new_[80102]_ ;
  assign \new_[80107]_  = \new_[80106]_  & \new_[80099]_ ;
  assign \new_[80110]_  = ~A236 & ~A235;
  assign \new_[80113]_  = ~A267 & ~A266;
  assign \new_[80114]_  = \new_[80113]_  & \new_[80110]_ ;
  assign \new_[80117]_  = ~A299 & A298;
  assign \new_[80120]_  = A301 & A300;
  assign \new_[80121]_  = \new_[80120]_  & \new_[80117]_ ;
  assign \new_[80122]_  = \new_[80121]_  & \new_[80114]_ ;
  assign \new_[80125]_  = A169 & ~A170;
  assign \new_[80128]_  = A166 & A167;
  assign \new_[80129]_  = \new_[80128]_  & \new_[80125]_ ;
  assign \new_[80132]_  = ~A202 & ~A200;
  assign \new_[80135]_  = ~A233 & ~A203;
  assign \new_[80136]_  = \new_[80135]_  & \new_[80132]_ ;
  assign \new_[80137]_  = \new_[80136]_  & \new_[80129]_ ;
  assign \new_[80140]_  = ~A236 & ~A235;
  assign \new_[80143]_  = ~A267 & ~A266;
  assign \new_[80144]_  = \new_[80143]_  & \new_[80140]_ ;
  assign \new_[80147]_  = ~A299 & A298;
  assign \new_[80150]_  = A302 & A300;
  assign \new_[80151]_  = \new_[80150]_  & \new_[80147]_ ;
  assign \new_[80152]_  = \new_[80151]_  & \new_[80144]_ ;
  assign \new_[80155]_  = A169 & ~A170;
  assign \new_[80158]_  = A166 & A167;
  assign \new_[80159]_  = \new_[80158]_  & \new_[80155]_ ;
  assign \new_[80162]_  = ~A202 & ~A200;
  assign \new_[80165]_  = ~A233 & ~A203;
  assign \new_[80166]_  = \new_[80165]_  & \new_[80162]_ ;
  assign \new_[80167]_  = \new_[80166]_  & \new_[80159]_ ;
  assign \new_[80170]_  = ~A236 & ~A235;
  assign \new_[80173]_  = ~A266 & ~A265;
  assign \new_[80174]_  = \new_[80173]_  & \new_[80170]_ ;
  assign \new_[80177]_  = ~A299 & A298;
  assign \new_[80180]_  = A301 & A300;
  assign \new_[80181]_  = \new_[80180]_  & \new_[80177]_ ;
  assign \new_[80182]_  = \new_[80181]_  & \new_[80174]_ ;
  assign \new_[80185]_  = A169 & ~A170;
  assign \new_[80188]_  = A166 & A167;
  assign \new_[80189]_  = \new_[80188]_  & \new_[80185]_ ;
  assign \new_[80192]_  = ~A202 & ~A200;
  assign \new_[80195]_  = ~A233 & ~A203;
  assign \new_[80196]_  = \new_[80195]_  & \new_[80192]_ ;
  assign \new_[80197]_  = \new_[80196]_  & \new_[80189]_ ;
  assign \new_[80200]_  = ~A236 & ~A235;
  assign \new_[80203]_  = ~A266 & ~A265;
  assign \new_[80204]_  = \new_[80203]_  & \new_[80200]_ ;
  assign \new_[80207]_  = ~A299 & A298;
  assign \new_[80210]_  = A302 & A300;
  assign \new_[80211]_  = \new_[80210]_  & \new_[80207]_ ;
  assign \new_[80212]_  = \new_[80211]_  & \new_[80204]_ ;
  assign \new_[80215]_  = A169 & ~A170;
  assign \new_[80218]_  = A166 & A167;
  assign \new_[80219]_  = \new_[80218]_  & \new_[80215]_ ;
  assign \new_[80222]_  = ~A202 & ~A200;
  assign \new_[80225]_  = ~A233 & ~A203;
  assign \new_[80226]_  = \new_[80225]_  & \new_[80222]_ ;
  assign \new_[80227]_  = \new_[80226]_  & \new_[80219]_ ;
  assign \new_[80230]_  = ~A266 & ~A234;
  assign \new_[80233]_  = ~A269 & ~A268;
  assign \new_[80234]_  = \new_[80233]_  & \new_[80230]_ ;
  assign \new_[80237]_  = ~A299 & A298;
  assign \new_[80240]_  = A301 & A300;
  assign \new_[80241]_  = \new_[80240]_  & \new_[80237]_ ;
  assign \new_[80242]_  = \new_[80241]_  & \new_[80234]_ ;
  assign \new_[80245]_  = A169 & ~A170;
  assign \new_[80248]_  = A166 & A167;
  assign \new_[80249]_  = \new_[80248]_  & \new_[80245]_ ;
  assign \new_[80252]_  = ~A202 & ~A200;
  assign \new_[80255]_  = ~A233 & ~A203;
  assign \new_[80256]_  = \new_[80255]_  & \new_[80252]_ ;
  assign \new_[80257]_  = \new_[80256]_  & \new_[80249]_ ;
  assign \new_[80260]_  = ~A266 & ~A234;
  assign \new_[80263]_  = ~A269 & ~A268;
  assign \new_[80264]_  = \new_[80263]_  & \new_[80260]_ ;
  assign \new_[80267]_  = ~A299 & A298;
  assign \new_[80270]_  = A302 & A300;
  assign \new_[80271]_  = \new_[80270]_  & \new_[80267]_ ;
  assign \new_[80272]_  = \new_[80271]_  & \new_[80264]_ ;
  assign \new_[80275]_  = A169 & ~A170;
  assign \new_[80278]_  = A166 & A167;
  assign \new_[80279]_  = \new_[80278]_  & \new_[80275]_ ;
  assign \new_[80282]_  = ~A202 & ~A200;
  assign \new_[80285]_  = ~A232 & ~A203;
  assign \new_[80286]_  = \new_[80285]_  & \new_[80282]_ ;
  assign \new_[80287]_  = \new_[80286]_  & \new_[80279]_ ;
  assign \new_[80290]_  = ~A266 & ~A233;
  assign \new_[80293]_  = ~A269 & ~A268;
  assign \new_[80294]_  = \new_[80293]_  & \new_[80290]_ ;
  assign \new_[80297]_  = ~A299 & A298;
  assign \new_[80300]_  = A301 & A300;
  assign \new_[80301]_  = \new_[80300]_  & \new_[80297]_ ;
  assign \new_[80302]_  = \new_[80301]_  & \new_[80294]_ ;
  assign \new_[80305]_  = A169 & ~A170;
  assign \new_[80308]_  = A166 & A167;
  assign \new_[80309]_  = \new_[80308]_  & \new_[80305]_ ;
  assign \new_[80312]_  = ~A202 & ~A200;
  assign \new_[80315]_  = ~A232 & ~A203;
  assign \new_[80316]_  = \new_[80315]_  & \new_[80312]_ ;
  assign \new_[80317]_  = \new_[80316]_  & \new_[80309]_ ;
  assign \new_[80320]_  = ~A266 & ~A233;
  assign \new_[80323]_  = ~A269 & ~A268;
  assign \new_[80324]_  = \new_[80323]_  & \new_[80320]_ ;
  assign \new_[80327]_  = ~A299 & A298;
  assign \new_[80330]_  = A302 & A300;
  assign \new_[80331]_  = \new_[80330]_  & \new_[80327]_ ;
  assign \new_[80332]_  = \new_[80331]_  & \new_[80324]_ ;
  assign \new_[80335]_  = A169 & ~A170;
  assign \new_[80338]_  = A166 & A167;
  assign \new_[80339]_  = \new_[80338]_  & \new_[80335]_ ;
  assign \new_[80342]_  = ~A201 & ~A200;
  assign \new_[80345]_  = ~A235 & ~A233;
  assign \new_[80346]_  = \new_[80345]_  & \new_[80342]_ ;
  assign \new_[80347]_  = \new_[80346]_  & \new_[80339]_ ;
  assign \new_[80350]_  = ~A266 & ~A236;
  assign \new_[80353]_  = ~A269 & ~A268;
  assign \new_[80354]_  = \new_[80353]_  & \new_[80350]_ ;
  assign \new_[80357]_  = ~A299 & A298;
  assign \new_[80360]_  = A301 & A300;
  assign \new_[80361]_  = \new_[80360]_  & \new_[80357]_ ;
  assign \new_[80362]_  = \new_[80361]_  & \new_[80354]_ ;
  assign \new_[80365]_  = A169 & ~A170;
  assign \new_[80368]_  = A166 & A167;
  assign \new_[80369]_  = \new_[80368]_  & \new_[80365]_ ;
  assign \new_[80372]_  = ~A201 & ~A200;
  assign \new_[80375]_  = ~A235 & ~A233;
  assign \new_[80376]_  = \new_[80375]_  & \new_[80372]_ ;
  assign \new_[80377]_  = \new_[80376]_  & \new_[80369]_ ;
  assign \new_[80380]_  = ~A266 & ~A236;
  assign \new_[80383]_  = ~A269 & ~A268;
  assign \new_[80384]_  = \new_[80383]_  & \new_[80380]_ ;
  assign \new_[80387]_  = ~A299 & A298;
  assign \new_[80390]_  = A302 & A300;
  assign \new_[80391]_  = \new_[80390]_  & \new_[80387]_ ;
  assign \new_[80392]_  = \new_[80391]_  & \new_[80384]_ ;
  assign \new_[80395]_  = A169 & ~A170;
  assign \new_[80398]_  = A166 & A167;
  assign \new_[80399]_  = \new_[80398]_  & \new_[80395]_ ;
  assign \new_[80402]_  = ~A200 & ~A199;
  assign \new_[80405]_  = ~A235 & ~A233;
  assign \new_[80406]_  = \new_[80405]_  & \new_[80402]_ ;
  assign \new_[80407]_  = \new_[80406]_  & \new_[80399]_ ;
  assign \new_[80410]_  = ~A266 & ~A236;
  assign \new_[80413]_  = ~A269 & ~A268;
  assign \new_[80414]_  = \new_[80413]_  & \new_[80410]_ ;
  assign \new_[80417]_  = ~A299 & A298;
  assign \new_[80420]_  = A301 & A300;
  assign \new_[80421]_  = \new_[80420]_  & \new_[80417]_ ;
  assign \new_[80422]_  = \new_[80421]_  & \new_[80414]_ ;
  assign \new_[80425]_  = A169 & ~A170;
  assign \new_[80428]_  = A166 & A167;
  assign \new_[80429]_  = \new_[80428]_  & \new_[80425]_ ;
  assign \new_[80432]_  = ~A200 & ~A199;
  assign \new_[80435]_  = ~A235 & ~A233;
  assign \new_[80436]_  = \new_[80435]_  & \new_[80432]_ ;
  assign \new_[80437]_  = \new_[80436]_  & \new_[80429]_ ;
  assign \new_[80440]_  = ~A266 & ~A236;
  assign \new_[80443]_  = ~A269 & ~A268;
  assign \new_[80444]_  = \new_[80443]_  & \new_[80440]_ ;
  assign \new_[80447]_  = ~A299 & A298;
  assign \new_[80450]_  = A302 & A300;
  assign \new_[80451]_  = \new_[80450]_  & \new_[80447]_ ;
  assign \new_[80452]_  = \new_[80451]_  & \new_[80444]_ ;
  assign \new_[80455]_  = A169 & ~A170;
  assign \new_[80458]_  = ~A166 & ~A167;
  assign \new_[80459]_  = \new_[80458]_  & \new_[80455]_ ;
  assign \new_[80462]_  = A200 & A199;
  assign \new_[80465]_  = ~A235 & ~A233;
  assign \new_[80466]_  = \new_[80465]_  & \new_[80462]_ ;
  assign \new_[80467]_  = \new_[80466]_  & \new_[80459]_ ;
  assign \new_[80470]_  = ~A266 & ~A236;
  assign \new_[80473]_  = ~A269 & ~A268;
  assign \new_[80474]_  = \new_[80473]_  & \new_[80470]_ ;
  assign \new_[80477]_  = ~A299 & A298;
  assign \new_[80480]_  = A301 & A300;
  assign \new_[80481]_  = \new_[80480]_  & \new_[80477]_ ;
  assign \new_[80482]_  = \new_[80481]_  & \new_[80474]_ ;
  assign \new_[80485]_  = A169 & ~A170;
  assign \new_[80488]_  = ~A166 & ~A167;
  assign \new_[80489]_  = \new_[80488]_  & \new_[80485]_ ;
  assign \new_[80492]_  = A200 & A199;
  assign \new_[80495]_  = ~A235 & ~A233;
  assign \new_[80496]_  = \new_[80495]_  & \new_[80492]_ ;
  assign \new_[80497]_  = \new_[80496]_  & \new_[80489]_ ;
  assign \new_[80500]_  = ~A266 & ~A236;
  assign \new_[80503]_  = ~A269 & ~A268;
  assign \new_[80504]_  = \new_[80503]_  & \new_[80500]_ ;
  assign \new_[80507]_  = ~A299 & A298;
  assign \new_[80510]_  = A302 & A300;
  assign \new_[80511]_  = \new_[80510]_  & \new_[80507]_ ;
  assign \new_[80512]_  = \new_[80511]_  & \new_[80504]_ ;
  assign \new_[80515]_  = A169 & ~A170;
  assign \new_[80518]_  = ~A166 & ~A167;
  assign \new_[80519]_  = \new_[80518]_  & \new_[80515]_ ;
  assign \new_[80522]_  = ~A202 & ~A200;
  assign \new_[80525]_  = A232 & ~A203;
  assign \new_[80526]_  = \new_[80525]_  & \new_[80522]_ ;
  assign \new_[80527]_  = \new_[80526]_  & \new_[80519]_ ;
  assign \new_[80530]_  = A265 & A233;
  assign \new_[80533]_  = ~A269 & ~A268;
  assign \new_[80534]_  = \new_[80533]_  & \new_[80530]_ ;
  assign \new_[80537]_  = ~A299 & A298;
  assign \new_[80540]_  = A301 & A300;
  assign \new_[80541]_  = \new_[80540]_  & \new_[80537]_ ;
  assign \new_[80542]_  = \new_[80541]_  & \new_[80534]_ ;
  assign \new_[80545]_  = A169 & ~A170;
  assign \new_[80548]_  = ~A166 & ~A167;
  assign \new_[80549]_  = \new_[80548]_  & \new_[80545]_ ;
  assign \new_[80552]_  = ~A202 & ~A200;
  assign \new_[80555]_  = A232 & ~A203;
  assign \new_[80556]_  = \new_[80555]_  & \new_[80552]_ ;
  assign \new_[80557]_  = \new_[80556]_  & \new_[80549]_ ;
  assign \new_[80560]_  = A265 & A233;
  assign \new_[80563]_  = ~A269 & ~A268;
  assign \new_[80564]_  = \new_[80563]_  & \new_[80560]_ ;
  assign \new_[80567]_  = ~A299 & A298;
  assign \new_[80570]_  = A302 & A300;
  assign \new_[80571]_  = \new_[80570]_  & \new_[80567]_ ;
  assign \new_[80572]_  = \new_[80571]_  & \new_[80564]_ ;
  assign \new_[80575]_  = A169 & ~A170;
  assign \new_[80578]_  = ~A166 & ~A167;
  assign \new_[80579]_  = \new_[80578]_  & \new_[80575]_ ;
  assign \new_[80582]_  = ~A202 & ~A200;
  assign \new_[80585]_  = ~A233 & ~A203;
  assign \new_[80586]_  = \new_[80585]_  & \new_[80582]_ ;
  assign \new_[80587]_  = \new_[80586]_  & \new_[80579]_ ;
  assign \new_[80590]_  = ~A236 & ~A235;
  assign \new_[80593]_  = A266 & A265;
  assign \new_[80594]_  = \new_[80593]_  & \new_[80590]_ ;
  assign \new_[80597]_  = ~A299 & A298;
  assign \new_[80600]_  = A301 & A300;
  assign \new_[80601]_  = \new_[80600]_  & \new_[80597]_ ;
  assign \new_[80602]_  = \new_[80601]_  & \new_[80594]_ ;
  assign \new_[80605]_  = A169 & ~A170;
  assign \new_[80608]_  = ~A166 & ~A167;
  assign \new_[80609]_  = \new_[80608]_  & \new_[80605]_ ;
  assign \new_[80612]_  = ~A202 & ~A200;
  assign \new_[80615]_  = ~A233 & ~A203;
  assign \new_[80616]_  = \new_[80615]_  & \new_[80612]_ ;
  assign \new_[80617]_  = \new_[80616]_  & \new_[80609]_ ;
  assign \new_[80620]_  = ~A236 & ~A235;
  assign \new_[80623]_  = A266 & A265;
  assign \new_[80624]_  = \new_[80623]_  & \new_[80620]_ ;
  assign \new_[80627]_  = ~A299 & A298;
  assign \new_[80630]_  = A302 & A300;
  assign \new_[80631]_  = \new_[80630]_  & \new_[80627]_ ;
  assign \new_[80632]_  = \new_[80631]_  & \new_[80624]_ ;
  assign \new_[80635]_  = A169 & ~A170;
  assign \new_[80638]_  = ~A166 & ~A167;
  assign \new_[80639]_  = \new_[80638]_  & \new_[80635]_ ;
  assign \new_[80642]_  = ~A202 & ~A200;
  assign \new_[80645]_  = ~A233 & ~A203;
  assign \new_[80646]_  = \new_[80645]_  & \new_[80642]_ ;
  assign \new_[80647]_  = \new_[80646]_  & \new_[80639]_ ;
  assign \new_[80650]_  = ~A236 & ~A235;
  assign \new_[80653]_  = ~A267 & ~A266;
  assign \new_[80654]_  = \new_[80653]_  & \new_[80650]_ ;
  assign \new_[80657]_  = ~A299 & A298;
  assign \new_[80660]_  = A301 & A300;
  assign \new_[80661]_  = \new_[80660]_  & \new_[80657]_ ;
  assign \new_[80662]_  = \new_[80661]_  & \new_[80654]_ ;
  assign \new_[80665]_  = A169 & ~A170;
  assign \new_[80668]_  = ~A166 & ~A167;
  assign \new_[80669]_  = \new_[80668]_  & \new_[80665]_ ;
  assign \new_[80672]_  = ~A202 & ~A200;
  assign \new_[80675]_  = ~A233 & ~A203;
  assign \new_[80676]_  = \new_[80675]_  & \new_[80672]_ ;
  assign \new_[80677]_  = \new_[80676]_  & \new_[80669]_ ;
  assign \new_[80680]_  = ~A236 & ~A235;
  assign \new_[80683]_  = ~A267 & ~A266;
  assign \new_[80684]_  = \new_[80683]_  & \new_[80680]_ ;
  assign \new_[80687]_  = ~A299 & A298;
  assign \new_[80690]_  = A302 & A300;
  assign \new_[80691]_  = \new_[80690]_  & \new_[80687]_ ;
  assign \new_[80692]_  = \new_[80691]_  & \new_[80684]_ ;
  assign \new_[80695]_  = A169 & ~A170;
  assign \new_[80698]_  = ~A166 & ~A167;
  assign \new_[80699]_  = \new_[80698]_  & \new_[80695]_ ;
  assign \new_[80702]_  = ~A202 & ~A200;
  assign \new_[80705]_  = ~A233 & ~A203;
  assign \new_[80706]_  = \new_[80705]_  & \new_[80702]_ ;
  assign \new_[80707]_  = \new_[80706]_  & \new_[80699]_ ;
  assign \new_[80710]_  = ~A236 & ~A235;
  assign \new_[80713]_  = ~A266 & ~A265;
  assign \new_[80714]_  = \new_[80713]_  & \new_[80710]_ ;
  assign \new_[80717]_  = ~A299 & A298;
  assign \new_[80720]_  = A301 & A300;
  assign \new_[80721]_  = \new_[80720]_  & \new_[80717]_ ;
  assign \new_[80722]_  = \new_[80721]_  & \new_[80714]_ ;
  assign \new_[80725]_  = A169 & ~A170;
  assign \new_[80728]_  = ~A166 & ~A167;
  assign \new_[80729]_  = \new_[80728]_  & \new_[80725]_ ;
  assign \new_[80732]_  = ~A202 & ~A200;
  assign \new_[80735]_  = ~A233 & ~A203;
  assign \new_[80736]_  = \new_[80735]_  & \new_[80732]_ ;
  assign \new_[80737]_  = \new_[80736]_  & \new_[80729]_ ;
  assign \new_[80740]_  = ~A236 & ~A235;
  assign \new_[80743]_  = ~A266 & ~A265;
  assign \new_[80744]_  = \new_[80743]_  & \new_[80740]_ ;
  assign \new_[80747]_  = ~A299 & A298;
  assign \new_[80750]_  = A302 & A300;
  assign \new_[80751]_  = \new_[80750]_  & \new_[80747]_ ;
  assign \new_[80752]_  = \new_[80751]_  & \new_[80744]_ ;
  assign \new_[80755]_  = A169 & ~A170;
  assign \new_[80758]_  = ~A166 & ~A167;
  assign \new_[80759]_  = \new_[80758]_  & \new_[80755]_ ;
  assign \new_[80762]_  = ~A202 & ~A200;
  assign \new_[80765]_  = ~A233 & ~A203;
  assign \new_[80766]_  = \new_[80765]_  & \new_[80762]_ ;
  assign \new_[80767]_  = \new_[80766]_  & \new_[80759]_ ;
  assign \new_[80770]_  = ~A266 & ~A234;
  assign \new_[80773]_  = ~A269 & ~A268;
  assign \new_[80774]_  = \new_[80773]_  & \new_[80770]_ ;
  assign \new_[80777]_  = ~A299 & A298;
  assign \new_[80780]_  = A301 & A300;
  assign \new_[80781]_  = \new_[80780]_  & \new_[80777]_ ;
  assign \new_[80782]_  = \new_[80781]_  & \new_[80774]_ ;
  assign \new_[80785]_  = A169 & ~A170;
  assign \new_[80788]_  = ~A166 & ~A167;
  assign \new_[80789]_  = \new_[80788]_  & \new_[80785]_ ;
  assign \new_[80792]_  = ~A202 & ~A200;
  assign \new_[80795]_  = ~A233 & ~A203;
  assign \new_[80796]_  = \new_[80795]_  & \new_[80792]_ ;
  assign \new_[80797]_  = \new_[80796]_  & \new_[80789]_ ;
  assign \new_[80800]_  = ~A266 & ~A234;
  assign \new_[80803]_  = ~A269 & ~A268;
  assign \new_[80804]_  = \new_[80803]_  & \new_[80800]_ ;
  assign \new_[80807]_  = ~A299 & A298;
  assign \new_[80810]_  = A302 & A300;
  assign \new_[80811]_  = \new_[80810]_  & \new_[80807]_ ;
  assign \new_[80812]_  = \new_[80811]_  & \new_[80804]_ ;
  assign \new_[80815]_  = A169 & ~A170;
  assign \new_[80818]_  = ~A166 & ~A167;
  assign \new_[80819]_  = \new_[80818]_  & \new_[80815]_ ;
  assign \new_[80822]_  = ~A202 & ~A200;
  assign \new_[80825]_  = ~A232 & ~A203;
  assign \new_[80826]_  = \new_[80825]_  & \new_[80822]_ ;
  assign \new_[80827]_  = \new_[80826]_  & \new_[80819]_ ;
  assign \new_[80830]_  = ~A266 & ~A233;
  assign \new_[80833]_  = ~A269 & ~A268;
  assign \new_[80834]_  = \new_[80833]_  & \new_[80830]_ ;
  assign \new_[80837]_  = ~A299 & A298;
  assign \new_[80840]_  = A301 & A300;
  assign \new_[80841]_  = \new_[80840]_  & \new_[80837]_ ;
  assign \new_[80842]_  = \new_[80841]_  & \new_[80834]_ ;
  assign \new_[80845]_  = A169 & ~A170;
  assign \new_[80848]_  = ~A166 & ~A167;
  assign \new_[80849]_  = \new_[80848]_  & \new_[80845]_ ;
  assign \new_[80852]_  = ~A202 & ~A200;
  assign \new_[80855]_  = ~A232 & ~A203;
  assign \new_[80856]_  = \new_[80855]_  & \new_[80852]_ ;
  assign \new_[80857]_  = \new_[80856]_  & \new_[80849]_ ;
  assign \new_[80860]_  = ~A266 & ~A233;
  assign \new_[80863]_  = ~A269 & ~A268;
  assign \new_[80864]_  = \new_[80863]_  & \new_[80860]_ ;
  assign \new_[80867]_  = ~A299 & A298;
  assign \new_[80870]_  = A302 & A300;
  assign \new_[80871]_  = \new_[80870]_  & \new_[80867]_ ;
  assign \new_[80872]_  = \new_[80871]_  & \new_[80864]_ ;
  assign \new_[80875]_  = A169 & ~A170;
  assign \new_[80878]_  = ~A166 & ~A167;
  assign \new_[80879]_  = \new_[80878]_  & \new_[80875]_ ;
  assign \new_[80882]_  = ~A201 & ~A200;
  assign \new_[80885]_  = ~A235 & ~A233;
  assign \new_[80886]_  = \new_[80885]_  & \new_[80882]_ ;
  assign \new_[80887]_  = \new_[80886]_  & \new_[80879]_ ;
  assign \new_[80890]_  = ~A266 & ~A236;
  assign \new_[80893]_  = ~A269 & ~A268;
  assign \new_[80894]_  = \new_[80893]_  & \new_[80890]_ ;
  assign \new_[80897]_  = ~A299 & A298;
  assign \new_[80900]_  = A301 & A300;
  assign \new_[80901]_  = \new_[80900]_  & \new_[80897]_ ;
  assign \new_[80902]_  = \new_[80901]_  & \new_[80894]_ ;
  assign \new_[80905]_  = A169 & ~A170;
  assign \new_[80908]_  = ~A166 & ~A167;
  assign \new_[80909]_  = \new_[80908]_  & \new_[80905]_ ;
  assign \new_[80912]_  = ~A201 & ~A200;
  assign \new_[80915]_  = ~A235 & ~A233;
  assign \new_[80916]_  = \new_[80915]_  & \new_[80912]_ ;
  assign \new_[80917]_  = \new_[80916]_  & \new_[80909]_ ;
  assign \new_[80920]_  = ~A266 & ~A236;
  assign \new_[80923]_  = ~A269 & ~A268;
  assign \new_[80924]_  = \new_[80923]_  & \new_[80920]_ ;
  assign \new_[80927]_  = ~A299 & A298;
  assign \new_[80930]_  = A302 & A300;
  assign \new_[80931]_  = \new_[80930]_  & \new_[80927]_ ;
  assign \new_[80932]_  = \new_[80931]_  & \new_[80924]_ ;
  assign \new_[80935]_  = A169 & ~A170;
  assign \new_[80938]_  = ~A166 & ~A167;
  assign \new_[80939]_  = \new_[80938]_  & \new_[80935]_ ;
  assign \new_[80942]_  = ~A200 & ~A199;
  assign \new_[80945]_  = ~A235 & ~A233;
  assign \new_[80946]_  = \new_[80945]_  & \new_[80942]_ ;
  assign \new_[80947]_  = \new_[80946]_  & \new_[80939]_ ;
  assign \new_[80950]_  = ~A266 & ~A236;
  assign \new_[80953]_  = ~A269 & ~A268;
  assign \new_[80954]_  = \new_[80953]_  & \new_[80950]_ ;
  assign \new_[80957]_  = ~A299 & A298;
  assign \new_[80960]_  = A301 & A300;
  assign \new_[80961]_  = \new_[80960]_  & \new_[80957]_ ;
  assign \new_[80962]_  = \new_[80961]_  & \new_[80954]_ ;
  assign \new_[80965]_  = A169 & ~A170;
  assign \new_[80968]_  = ~A166 & ~A167;
  assign \new_[80969]_  = \new_[80968]_  & \new_[80965]_ ;
  assign \new_[80972]_  = ~A200 & ~A199;
  assign \new_[80975]_  = ~A235 & ~A233;
  assign \new_[80976]_  = \new_[80975]_  & \new_[80972]_ ;
  assign \new_[80977]_  = \new_[80976]_  & \new_[80969]_ ;
  assign \new_[80980]_  = ~A266 & ~A236;
  assign \new_[80983]_  = ~A269 & ~A268;
  assign \new_[80984]_  = \new_[80983]_  & \new_[80980]_ ;
  assign \new_[80987]_  = ~A299 & A298;
  assign \new_[80990]_  = A302 & A300;
  assign \new_[80991]_  = \new_[80990]_  & \new_[80987]_ ;
  assign \new_[80992]_  = \new_[80991]_  & \new_[80984]_ ;
  assign \new_[80995]_  = ~A167 & ~A169;
  assign \new_[80998]_  = A199 & ~A166;
  assign \new_[80999]_  = \new_[80998]_  & \new_[80995]_ ;
  assign \new_[81002]_  = A201 & ~A200;
  assign \new_[81005]_  = A232 & A202;
  assign \new_[81006]_  = \new_[81005]_  & \new_[81002]_ ;
  assign \new_[81007]_  = \new_[81006]_  & \new_[80999]_ ;
  assign \new_[81010]_  = A265 & A233;
  assign \new_[81013]_  = ~A269 & ~A268;
  assign \new_[81014]_  = \new_[81013]_  & \new_[81010]_ ;
  assign \new_[81017]_  = ~A299 & A298;
  assign \new_[81020]_  = A301 & A300;
  assign \new_[81021]_  = \new_[81020]_  & \new_[81017]_ ;
  assign \new_[81022]_  = \new_[81021]_  & \new_[81014]_ ;
  assign \new_[81025]_  = ~A167 & ~A169;
  assign \new_[81028]_  = A199 & ~A166;
  assign \new_[81029]_  = \new_[81028]_  & \new_[81025]_ ;
  assign \new_[81032]_  = A201 & ~A200;
  assign \new_[81035]_  = A232 & A202;
  assign \new_[81036]_  = \new_[81035]_  & \new_[81032]_ ;
  assign \new_[81037]_  = \new_[81036]_  & \new_[81029]_ ;
  assign \new_[81040]_  = A265 & A233;
  assign \new_[81043]_  = ~A269 & ~A268;
  assign \new_[81044]_  = \new_[81043]_  & \new_[81040]_ ;
  assign \new_[81047]_  = ~A299 & A298;
  assign \new_[81050]_  = A302 & A300;
  assign \new_[81051]_  = \new_[81050]_  & \new_[81047]_ ;
  assign \new_[81052]_  = \new_[81051]_  & \new_[81044]_ ;
  assign \new_[81055]_  = ~A167 & ~A169;
  assign \new_[81058]_  = A199 & ~A166;
  assign \new_[81059]_  = \new_[81058]_  & \new_[81055]_ ;
  assign \new_[81062]_  = A201 & ~A200;
  assign \new_[81065]_  = ~A233 & A202;
  assign \new_[81066]_  = \new_[81065]_  & \new_[81062]_ ;
  assign \new_[81067]_  = \new_[81066]_  & \new_[81059]_ ;
  assign \new_[81070]_  = ~A236 & ~A235;
  assign \new_[81073]_  = A266 & A265;
  assign \new_[81074]_  = \new_[81073]_  & \new_[81070]_ ;
  assign \new_[81077]_  = ~A299 & A298;
  assign \new_[81080]_  = A301 & A300;
  assign \new_[81081]_  = \new_[81080]_  & \new_[81077]_ ;
  assign \new_[81082]_  = \new_[81081]_  & \new_[81074]_ ;
  assign \new_[81085]_  = ~A167 & ~A169;
  assign \new_[81088]_  = A199 & ~A166;
  assign \new_[81089]_  = \new_[81088]_  & \new_[81085]_ ;
  assign \new_[81092]_  = A201 & ~A200;
  assign \new_[81095]_  = ~A233 & A202;
  assign \new_[81096]_  = \new_[81095]_  & \new_[81092]_ ;
  assign \new_[81097]_  = \new_[81096]_  & \new_[81089]_ ;
  assign \new_[81100]_  = ~A236 & ~A235;
  assign \new_[81103]_  = A266 & A265;
  assign \new_[81104]_  = \new_[81103]_  & \new_[81100]_ ;
  assign \new_[81107]_  = ~A299 & A298;
  assign \new_[81110]_  = A302 & A300;
  assign \new_[81111]_  = \new_[81110]_  & \new_[81107]_ ;
  assign \new_[81112]_  = \new_[81111]_  & \new_[81104]_ ;
  assign \new_[81115]_  = ~A167 & ~A169;
  assign \new_[81118]_  = A199 & ~A166;
  assign \new_[81119]_  = \new_[81118]_  & \new_[81115]_ ;
  assign \new_[81122]_  = A201 & ~A200;
  assign \new_[81125]_  = ~A233 & A202;
  assign \new_[81126]_  = \new_[81125]_  & \new_[81122]_ ;
  assign \new_[81127]_  = \new_[81126]_  & \new_[81119]_ ;
  assign \new_[81130]_  = ~A236 & ~A235;
  assign \new_[81133]_  = ~A267 & ~A266;
  assign \new_[81134]_  = \new_[81133]_  & \new_[81130]_ ;
  assign \new_[81137]_  = ~A299 & A298;
  assign \new_[81140]_  = A301 & A300;
  assign \new_[81141]_  = \new_[81140]_  & \new_[81137]_ ;
  assign \new_[81142]_  = \new_[81141]_  & \new_[81134]_ ;
  assign \new_[81145]_  = ~A167 & ~A169;
  assign \new_[81148]_  = A199 & ~A166;
  assign \new_[81149]_  = \new_[81148]_  & \new_[81145]_ ;
  assign \new_[81152]_  = A201 & ~A200;
  assign \new_[81155]_  = ~A233 & A202;
  assign \new_[81156]_  = \new_[81155]_  & \new_[81152]_ ;
  assign \new_[81157]_  = \new_[81156]_  & \new_[81149]_ ;
  assign \new_[81160]_  = ~A236 & ~A235;
  assign \new_[81163]_  = ~A267 & ~A266;
  assign \new_[81164]_  = \new_[81163]_  & \new_[81160]_ ;
  assign \new_[81167]_  = ~A299 & A298;
  assign \new_[81170]_  = A302 & A300;
  assign \new_[81171]_  = \new_[81170]_  & \new_[81167]_ ;
  assign \new_[81172]_  = \new_[81171]_  & \new_[81164]_ ;
  assign \new_[81175]_  = ~A167 & ~A169;
  assign \new_[81178]_  = A199 & ~A166;
  assign \new_[81179]_  = \new_[81178]_  & \new_[81175]_ ;
  assign \new_[81182]_  = A201 & ~A200;
  assign \new_[81185]_  = ~A233 & A202;
  assign \new_[81186]_  = \new_[81185]_  & \new_[81182]_ ;
  assign \new_[81187]_  = \new_[81186]_  & \new_[81179]_ ;
  assign \new_[81190]_  = ~A236 & ~A235;
  assign \new_[81193]_  = ~A266 & ~A265;
  assign \new_[81194]_  = \new_[81193]_  & \new_[81190]_ ;
  assign \new_[81197]_  = ~A299 & A298;
  assign \new_[81200]_  = A301 & A300;
  assign \new_[81201]_  = \new_[81200]_  & \new_[81197]_ ;
  assign \new_[81202]_  = \new_[81201]_  & \new_[81194]_ ;
  assign \new_[81205]_  = ~A167 & ~A169;
  assign \new_[81208]_  = A199 & ~A166;
  assign \new_[81209]_  = \new_[81208]_  & \new_[81205]_ ;
  assign \new_[81212]_  = A201 & ~A200;
  assign \new_[81215]_  = ~A233 & A202;
  assign \new_[81216]_  = \new_[81215]_  & \new_[81212]_ ;
  assign \new_[81217]_  = \new_[81216]_  & \new_[81209]_ ;
  assign \new_[81220]_  = ~A236 & ~A235;
  assign \new_[81223]_  = ~A266 & ~A265;
  assign \new_[81224]_  = \new_[81223]_  & \new_[81220]_ ;
  assign \new_[81227]_  = ~A299 & A298;
  assign \new_[81230]_  = A302 & A300;
  assign \new_[81231]_  = \new_[81230]_  & \new_[81227]_ ;
  assign \new_[81232]_  = \new_[81231]_  & \new_[81224]_ ;
  assign \new_[81235]_  = ~A167 & ~A169;
  assign \new_[81238]_  = A199 & ~A166;
  assign \new_[81239]_  = \new_[81238]_  & \new_[81235]_ ;
  assign \new_[81242]_  = A201 & ~A200;
  assign \new_[81245]_  = ~A233 & A202;
  assign \new_[81246]_  = \new_[81245]_  & \new_[81242]_ ;
  assign \new_[81247]_  = \new_[81246]_  & \new_[81239]_ ;
  assign \new_[81250]_  = ~A266 & ~A234;
  assign \new_[81253]_  = ~A269 & ~A268;
  assign \new_[81254]_  = \new_[81253]_  & \new_[81250]_ ;
  assign \new_[81257]_  = ~A299 & A298;
  assign \new_[81260]_  = A301 & A300;
  assign \new_[81261]_  = \new_[81260]_  & \new_[81257]_ ;
  assign \new_[81262]_  = \new_[81261]_  & \new_[81254]_ ;
  assign \new_[81265]_  = ~A167 & ~A169;
  assign \new_[81268]_  = A199 & ~A166;
  assign \new_[81269]_  = \new_[81268]_  & \new_[81265]_ ;
  assign \new_[81272]_  = A201 & ~A200;
  assign \new_[81275]_  = ~A233 & A202;
  assign \new_[81276]_  = \new_[81275]_  & \new_[81272]_ ;
  assign \new_[81277]_  = \new_[81276]_  & \new_[81269]_ ;
  assign \new_[81280]_  = ~A266 & ~A234;
  assign \new_[81283]_  = ~A269 & ~A268;
  assign \new_[81284]_  = \new_[81283]_  & \new_[81280]_ ;
  assign \new_[81287]_  = ~A299 & A298;
  assign \new_[81290]_  = A302 & A300;
  assign \new_[81291]_  = \new_[81290]_  & \new_[81287]_ ;
  assign \new_[81292]_  = \new_[81291]_  & \new_[81284]_ ;
  assign \new_[81295]_  = ~A167 & ~A169;
  assign \new_[81298]_  = A199 & ~A166;
  assign \new_[81299]_  = \new_[81298]_  & \new_[81295]_ ;
  assign \new_[81302]_  = A201 & ~A200;
  assign \new_[81305]_  = ~A232 & A202;
  assign \new_[81306]_  = \new_[81305]_  & \new_[81302]_ ;
  assign \new_[81307]_  = \new_[81306]_  & \new_[81299]_ ;
  assign \new_[81310]_  = ~A266 & ~A233;
  assign \new_[81313]_  = ~A269 & ~A268;
  assign \new_[81314]_  = \new_[81313]_  & \new_[81310]_ ;
  assign \new_[81317]_  = ~A299 & A298;
  assign \new_[81320]_  = A301 & A300;
  assign \new_[81321]_  = \new_[81320]_  & \new_[81317]_ ;
  assign \new_[81322]_  = \new_[81321]_  & \new_[81314]_ ;
  assign \new_[81325]_  = ~A167 & ~A169;
  assign \new_[81328]_  = A199 & ~A166;
  assign \new_[81329]_  = \new_[81328]_  & \new_[81325]_ ;
  assign \new_[81332]_  = A201 & ~A200;
  assign \new_[81335]_  = ~A232 & A202;
  assign \new_[81336]_  = \new_[81335]_  & \new_[81332]_ ;
  assign \new_[81337]_  = \new_[81336]_  & \new_[81329]_ ;
  assign \new_[81340]_  = ~A266 & ~A233;
  assign \new_[81343]_  = ~A269 & ~A268;
  assign \new_[81344]_  = \new_[81343]_  & \new_[81340]_ ;
  assign \new_[81347]_  = ~A299 & A298;
  assign \new_[81350]_  = A302 & A300;
  assign \new_[81351]_  = \new_[81350]_  & \new_[81347]_ ;
  assign \new_[81352]_  = \new_[81351]_  & \new_[81344]_ ;
  assign \new_[81355]_  = ~A167 & ~A169;
  assign \new_[81358]_  = A199 & ~A166;
  assign \new_[81359]_  = \new_[81358]_  & \new_[81355]_ ;
  assign \new_[81362]_  = A201 & ~A200;
  assign \new_[81365]_  = A232 & A203;
  assign \new_[81366]_  = \new_[81365]_  & \new_[81362]_ ;
  assign \new_[81367]_  = \new_[81366]_  & \new_[81359]_ ;
  assign \new_[81370]_  = A265 & A233;
  assign \new_[81373]_  = ~A269 & ~A268;
  assign \new_[81374]_  = \new_[81373]_  & \new_[81370]_ ;
  assign \new_[81377]_  = ~A299 & A298;
  assign \new_[81380]_  = A301 & A300;
  assign \new_[81381]_  = \new_[81380]_  & \new_[81377]_ ;
  assign \new_[81382]_  = \new_[81381]_  & \new_[81374]_ ;
  assign \new_[81385]_  = ~A167 & ~A169;
  assign \new_[81388]_  = A199 & ~A166;
  assign \new_[81389]_  = \new_[81388]_  & \new_[81385]_ ;
  assign \new_[81392]_  = A201 & ~A200;
  assign \new_[81395]_  = A232 & A203;
  assign \new_[81396]_  = \new_[81395]_  & \new_[81392]_ ;
  assign \new_[81397]_  = \new_[81396]_  & \new_[81389]_ ;
  assign \new_[81400]_  = A265 & A233;
  assign \new_[81403]_  = ~A269 & ~A268;
  assign \new_[81404]_  = \new_[81403]_  & \new_[81400]_ ;
  assign \new_[81407]_  = ~A299 & A298;
  assign \new_[81410]_  = A302 & A300;
  assign \new_[81411]_  = \new_[81410]_  & \new_[81407]_ ;
  assign \new_[81412]_  = \new_[81411]_  & \new_[81404]_ ;
  assign \new_[81415]_  = ~A167 & ~A169;
  assign \new_[81418]_  = A199 & ~A166;
  assign \new_[81419]_  = \new_[81418]_  & \new_[81415]_ ;
  assign \new_[81422]_  = A201 & ~A200;
  assign \new_[81425]_  = ~A233 & A203;
  assign \new_[81426]_  = \new_[81425]_  & \new_[81422]_ ;
  assign \new_[81427]_  = \new_[81426]_  & \new_[81419]_ ;
  assign \new_[81430]_  = ~A236 & ~A235;
  assign \new_[81433]_  = A266 & A265;
  assign \new_[81434]_  = \new_[81433]_  & \new_[81430]_ ;
  assign \new_[81437]_  = ~A299 & A298;
  assign \new_[81440]_  = A301 & A300;
  assign \new_[81441]_  = \new_[81440]_  & \new_[81437]_ ;
  assign \new_[81442]_  = \new_[81441]_  & \new_[81434]_ ;
  assign \new_[81445]_  = ~A167 & ~A169;
  assign \new_[81448]_  = A199 & ~A166;
  assign \new_[81449]_  = \new_[81448]_  & \new_[81445]_ ;
  assign \new_[81452]_  = A201 & ~A200;
  assign \new_[81455]_  = ~A233 & A203;
  assign \new_[81456]_  = \new_[81455]_  & \new_[81452]_ ;
  assign \new_[81457]_  = \new_[81456]_  & \new_[81449]_ ;
  assign \new_[81460]_  = ~A236 & ~A235;
  assign \new_[81463]_  = A266 & A265;
  assign \new_[81464]_  = \new_[81463]_  & \new_[81460]_ ;
  assign \new_[81467]_  = ~A299 & A298;
  assign \new_[81470]_  = A302 & A300;
  assign \new_[81471]_  = \new_[81470]_  & \new_[81467]_ ;
  assign \new_[81472]_  = \new_[81471]_  & \new_[81464]_ ;
  assign \new_[81475]_  = ~A167 & ~A169;
  assign \new_[81478]_  = A199 & ~A166;
  assign \new_[81479]_  = \new_[81478]_  & \new_[81475]_ ;
  assign \new_[81482]_  = A201 & ~A200;
  assign \new_[81485]_  = ~A233 & A203;
  assign \new_[81486]_  = \new_[81485]_  & \new_[81482]_ ;
  assign \new_[81487]_  = \new_[81486]_  & \new_[81479]_ ;
  assign \new_[81490]_  = ~A236 & ~A235;
  assign \new_[81493]_  = ~A267 & ~A266;
  assign \new_[81494]_  = \new_[81493]_  & \new_[81490]_ ;
  assign \new_[81497]_  = ~A299 & A298;
  assign \new_[81500]_  = A301 & A300;
  assign \new_[81501]_  = \new_[81500]_  & \new_[81497]_ ;
  assign \new_[81502]_  = \new_[81501]_  & \new_[81494]_ ;
  assign \new_[81505]_  = ~A167 & ~A169;
  assign \new_[81508]_  = A199 & ~A166;
  assign \new_[81509]_  = \new_[81508]_  & \new_[81505]_ ;
  assign \new_[81512]_  = A201 & ~A200;
  assign \new_[81515]_  = ~A233 & A203;
  assign \new_[81516]_  = \new_[81515]_  & \new_[81512]_ ;
  assign \new_[81517]_  = \new_[81516]_  & \new_[81509]_ ;
  assign \new_[81520]_  = ~A236 & ~A235;
  assign \new_[81523]_  = ~A267 & ~A266;
  assign \new_[81524]_  = \new_[81523]_  & \new_[81520]_ ;
  assign \new_[81527]_  = ~A299 & A298;
  assign \new_[81530]_  = A302 & A300;
  assign \new_[81531]_  = \new_[81530]_  & \new_[81527]_ ;
  assign \new_[81532]_  = \new_[81531]_  & \new_[81524]_ ;
  assign \new_[81535]_  = ~A167 & ~A169;
  assign \new_[81538]_  = A199 & ~A166;
  assign \new_[81539]_  = \new_[81538]_  & \new_[81535]_ ;
  assign \new_[81542]_  = A201 & ~A200;
  assign \new_[81545]_  = ~A233 & A203;
  assign \new_[81546]_  = \new_[81545]_  & \new_[81542]_ ;
  assign \new_[81547]_  = \new_[81546]_  & \new_[81539]_ ;
  assign \new_[81550]_  = ~A236 & ~A235;
  assign \new_[81553]_  = ~A266 & ~A265;
  assign \new_[81554]_  = \new_[81553]_  & \new_[81550]_ ;
  assign \new_[81557]_  = ~A299 & A298;
  assign \new_[81560]_  = A301 & A300;
  assign \new_[81561]_  = \new_[81560]_  & \new_[81557]_ ;
  assign \new_[81562]_  = \new_[81561]_  & \new_[81554]_ ;
  assign \new_[81565]_  = ~A167 & ~A169;
  assign \new_[81568]_  = A199 & ~A166;
  assign \new_[81569]_  = \new_[81568]_  & \new_[81565]_ ;
  assign \new_[81572]_  = A201 & ~A200;
  assign \new_[81575]_  = ~A233 & A203;
  assign \new_[81576]_  = \new_[81575]_  & \new_[81572]_ ;
  assign \new_[81577]_  = \new_[81576]_  & \new_[81569]_ ;
  assign \new_[81580]_  = ~A236 & ~A235;
  assign \new_[81583]_  = ~A266 & ~A265;
  assign \new_[81584]_  = \new_[81583]_  & \new_[81580]_ ;
  assign \new_[81587]_  = ~A299 & A298;
  assign \new_[81590]_  = A302 & A300;
  assign \new_[81591]_  = \new_[81590]_  & \new_[81587]_ ;
  assign \new_[81592]_  = \new_[81591]_  & \new_[81584]_ ;
  assign \new_[81595]_  = ~A167 & ~A169;
  assign \new_[81598]_  = A199 & ~A166;
  assign \new_[81599]_  = \new_[81598]_  & \new_[81595]_ ;
  assign \new_[81602]_  = A201 & ~A200;
  assign \new_[81605]_  = ~A233 & A203;
  assign \new_[81606]_  = \new_[81605]_  & \new_[81602]_ ;
  assign \new_[81607]_  = \new_[81606]_  & \new_[81599]_ ;
  assign \new_[81610]_  = ~A266 & ~A234;
  assign \new_[81613]_  = ~A269 & ~A268;
  assign \new_[81614]_  = \new_[81613]_  & \new_[81610]_ ;
  assign \new_[81617]_  = ~A299 & A298;
  assign \new_[81620]_  = A301 & A300;
  assign \new_[81621]_  = \new_[81620]_  & \new_[81617]_ ;
  assign \new_[81622]_  = \new_[81621]_  & \new_[81614]_ ;
  assign \new_[81625]_  = ~A167 & ~A169;
  assign \new_[81628]_  = A199 & ~A166;
  assign \new_[81629]_  = \new_[81628]_  & \new_[81625]_ ;
  assign \new_[81632]_  = A201 & ~A200;
  assign \new_[81635]_  = ~A233 & A203;
  assign \new_[81636]_  = \new_[81635]_  & \new_[81632]_ ;
  assign \new_[81637]_  = \new_[81636]_  & \new_[81629]_ ;
  assign \new_[81640]_  = ~A266 & ~A234;
  assign \new_[81643]_  = ~A269 & ~A268;
  assign \new_[81644]_  = \new_[81643]_  & \new_[81640]_ ;
  assign \new_[81647]_  = ~A299 & A298;
  assign \new_[81650]_  = A302 & A300;
  assign \new_[81651]_  = \new_[81650]_  & \new_[81647]_ ;
  assign \new_[81652]_  = \new_[81651]_  & \new_[81644]_ ;
  assign \new_[81655]_  = ~A167 & ~A169;
  assign \new_[81658]_  = A199 & ~A166;
  assign \new_[81659]_  = \new_[81658]_  & \new_[81655]_ ;
  assign \new_[81662]_  = A201 & ~A200;
  assign \new_[81665]_  = ~A232 & A203;
  assign \new_[81666]_  = \new_[81665]_  & \new_[81662]_ ;
  assign \new_[81667]_  = \new_[81666]_  & \new_[81659]_ ;
  assign \new_[81670]_  = ~A266 & ~A233;
  assign \new_[81673]_  = ~A269 & ~A268;
  assign \new_[81674]_  = \new_[81673]_  & \new_[81670]_ ;
  assign \new_[81677]_  = ~A299 & A298;
  assign \new_[81680]_  = A301 & A300;
  assign \new_[81681]_  = \new_[81680]_  & \new_[81677]_ ;
  assign \new_[81682]_  = \new_[81681]_  & \new_[81674]_ ;
  assign \new_[81685]_  = ~A167 & ~A169;
  assign \new_[81688]_  = A199 & ~A166;
  assign \new_[81689]_  = \new_[81688]_  & \new_[81685]_ ;
  assign \new_[81692]_  = A201 & ~A200;
  assign \new_[81695]_  = ~A232 & A203;
  assign \new_[81696]_  = \new_[81695]_  & \new_[81692]_ ;
  assign \new_[81697]_  = \new_[81696]_  & \new_[81689]_ ;
  assign \new_[81700]_  = ~A266 & ~A233;
  assign \new_[81703]_  = ~A269 & ~A268;
  assign \new_[81704]_  = \new_[81703]_  & \new_[81700]_ ;
  assign \new_[81707]_  = ~A299 & A298;
  assign \new_[81710]_  = A302 & A300;
  assign \new_[81711]_  = \new_[81710]_  & \new_[81707]_ ;
  assign \new_[81712]_  = \new_[81711]_  & \new_[81704]_ ;
  assign \new_[81715]_  = ~A168 & ~A169;
  assign \new_[81718]_  = A166 & A167;
  assign \new_[81719]_  = \new_[81718]_  & \new_[81715]_ ;
  assign \new_[81722]_  = A200 & ~A199;
  assign \new_[81725]_  = ~A235 & ~A233;
  assign \new_[81726]_  = \new_[81725]_  & \new_[81722]_ ;
  assign \new_[81727]_  = \new_[81726]_  & \new_[81719]_ ;
  assign \new_[81730]_  = ~A266 & ~A236;
  assign \new_[81733]_  = ~A269 & ~A268;
  assign \new_[81734]_  = \new_[81733]_  & \new_[81730]_ ;
  assign \new_[81737]_  = ~A299 & A298;
  assign \new_[81740]_  = A301 & A300;
  assign \new_[81741]_  = \new_[81740]_  & \new_[81737]_ ;
  assign \new_[81742]_  = \new_[81741]_  & \new_[81734]_ ;
  assign \new_[81745]_  = ~A168 & ~A169;
  assign \new_[81748]_  = A166 & A167;
  assign \new_[81749]_  = \new_[81748]_  & \new_[81745]_ ;
  assign \new_[81752]_  = A200 & ~A199;
  assign \new_[81755]_  = ~A235 & ~A233;
  assign \new_[81756]_  = \new_[81755]_  & \new_[81752]_ ;
  assign \new_[81757]_  = \new_[81756]_  & \new_[81749]_ ;
  assign \new_[81760]_  = ~A266 & ~A236;
  assign \new_[81763]_  = ~A269 & ~A268;
  assign \new_[81764]_  = \new_[81763]_  & \new_[81760]_ ;
  assign \new_[81767]_  = ~A299 & A298;
  assign \new_[81770]_  = A302 & A300;
  assign \new_[81771]_  = \new_[81770]_  & \new_[81767]_ ;
  assign \new_[81772]_  = \new_[81771]_  & \new_[81764]_ ;
  assign \new_[81775]_  = ~A168 & ~A169;
  assign \new_[81778]_  = A166 & A167;
  assign \new_[81779]_  = \new_[81778]_  & \new_[81775]_ ;
  assign \new_[81782]_  = ~A200 & A199;
  assign \new_[81785]_  = A202 & A201;
  assign \new_[81786]_  = \new_[81785]_  & \new_[81782]_ ;
  assign \new_[81787]_  = \new_[81786]_  & \new_[81779]_ ;
  assign \new_[81790]_  = A233 & A232;
  assign \new_[81793]_  = ~A267 & A265;
  assign \new_[81794]_  = \new_[81793]_  & \new_[81790]_ ;
  assign \new_[81797]_  = ~A299 & A298;
  assign \new_[81800]_  = A301 & A300;
  assign \new_[81801]_  = \new_[81800]_  & \new_[81797]_ ;
  assign \new_[81802]_  = \new_[81801]_  & \new_[81794]_ ;
  assign \new_[81805]_  = ~A168 & ~A169;
  assign \new_[81808]_  = A166 & A167;
  assign \new_[81809]_  = \new_[81808]_  & \new_[81805]_ ;
  assign \new_[81812]_  = ~A200 & A199;
  assign \new_[81815]_  = A202 & A201;
  assign \new_[81816]_  = \new_[81815]_  & \new_[81812]_ ;
  assign \new_[81817]_  = \new_[81816]_  & \new_[81809]_ ;
  assign \new_[81820]_  = A233 & A232;
  assign \new_[81823]_  = ~A267 & A265;
  assign \new_[81824]_  = \new_[81823]_  & \new_[81820]_ ;
  assign \new_[81827]_  = ~A299 & A298;
  assign \new_[81830]_  = A302 & A300;
  assign \new_[81831]_  = \new_[81830]_  & \new_[81827]_ ;
  assign \new_[81832]_  = \new_[81831]_  & \new_[81824]_ ;
  assign \new_[81835]_  = ~A168 & ~A169;
  assign \new_[81838]_  = A166 & A167;
  assign \new_[81839]_  = \new_[81838]_  & \new_[81835]_ ;
  assign \new_[81842]_  = ~A200 & A199;
  assign \new_[81845]_  = A202 & A201;
  assign \new_[81846]_  = \new_[81845]_  & \new_[81842]_ ;
  assign \new_[81847]_  = \new_[81846]_  & \new_[81839]_ ;
  assign \new_[81850]_  = A233 & A232;
  assign \new_[81853]_  = A266 & A265;
  assign \new_[81854]_  = \new_[81853]_  & \new_[81850]_ ;
  assign \new_[81857]_  = ~A299 & A298;
  assign \new_[81860]_  = A301 & A300;
  assign \new_[81861]_  = \new_[81860]_  & \new_[81857]_ ;
  assign \new_[81862]_  = \new_[81861]_  & \new_[81854]_ ;
  assign \new_[81865]_  = ~A168 & ~A169;
  assign \new_[81868]_  = A166 & A167;
  assign \new_[81869]_  = \new_[81868]_  & \new_[81865]_ ;
  assign \new_[81872]_  = ~A200 & A199;
  assign \new_[81875]_  = A202 & A201;
  assign \new_[81876]_  = \new_[81875]_  & \new_[81872]_ ;
  assign \new_[81877]_  = \new_[81876]_  & \new_[81869]_ ;
  assign \new_[81880]_  = A233 & A232;
  assign \new_[81883]_  = A266 & A265;
  assign \new_[81884]_  = \new_[81883]_  & \new_[81880]_ ;
  assign \new_[81887]_  = ~A299 & A298;
  assign \new_[81890]_  = A302 & A300;
  assign \new_[81891]_  = \new_[81890]_  & \new_[81887]_ ;
  assign \new_[81892]_  = \new_[81891]_  & \new_[81884]_ ;
  assign \new_[81895]_  = ~A168 & ~A169;
  assign \new_[81898]_  = A166 & A167;
  assign \new_[81899]_  = \new_[81898]_  & \new_[81895]_ ;
  assign \new_[81902]_  = ~A200 & A199;
  assign \new_[81905]_  = A202 & A201;
  assign \new_[81906]_  = \new_[81905]_  & \new_[81902]_ ;
  assign \new_[81907]_  = \new_[81906]_  & \new_[81899]_ ;
  assign \new_[81910]_  = A233 & A232;
  assign \new_[81913]_  = ~A266 & ~A265;
  assign \new_[81914]_  = \new_[81913]_  & \new_[81910]_ ;
  assign \new_[81917]_  = ~A299 & A298;
  assign \new_[81920]_  = A301 & A300;
  assign \new_[81921]_  = \new_[81920]_  & \new_[81917]_ ;
  assign \new_[81922]_  = \new_[81921]_  & \new_[81914]_ ;
  assign \new_[81925]_  = ~A168 & ~A169;
  assign \new_[81928]_  = A166 & A167;
  assign \new_[81929]_  = \new_[81928]_  & \new_[81925]_ ;
  assign \new_[81932]_  = ~A200 & A199;
  assign \new_[81935]_  = A202 & A201;
  assign \new_[81936]_  = \new_[81935]_  & \new_[81932]_ ;
  assign \new_[81937]_  = \new_[81936]_  & \new_[81929]_ ;
  assign \new_[81940]_  = A233 & A232;
  assign \new_[81943]_  = ~A266 & ~A265;
  assign \new_[81944]_  = \new_[81943]_  & \new_[81940]_ ;
  assign \new_[81947]_  = ~A299 & A298;
  assign \new_[81950]_  = A302 & A300;
  assign \new_[81951]_  = \new_[81950]_  & \new_[81947]_ ;
  assign \new_[81952]_  = \new_[81951]_  & \new_[81944]_ ;
  assign \new_[81955]_  = ~A168 & ~A169;
  assign \new_[81958]_  = A166 & A167;
  assign \new_[81959]_  = \new_[81958]_  & \new_[81955]_ ;
  assign \new_[81962]_  = ~A200 & A199;
  assign \new_[81965]_  = A202 & A201;
  assign \new_[81966]_  = \new_[81965]_  & \new_[81962]_ ;
  assign \new_[81967]_  = \new_[81966]_  & \new_[81959]_ ;
  assign \new_[81970]_  = ~A235 & ~A233;
  assign \new_[81973]_  = ~A266 & ~A236;
  assign \new_[81974]_  = \new_[81973]_  & \new_[81970]_ ;
  assign \new_[81977]_  = ~A269 & ~A268;
  assign \new_[81980]_  = A299 & ~A298;
  assign \new_[81981]_  = \new_[81980]_  & \new_[81977]_ ;
  assign \new_[81982]_  = \new_[81981]_  & \new_[81974]_ ;
  assign \new_[81985]_  = ~A168 & ~A169;
  assign \new_[81988]_  = A166 & A167;
  assign \new_[81989]_  = \new_[81988]_  & \new_[81985]_ ;
  assign \new_[81992]_  = ~A200 & A199;
  assign \new_[81995]_  = A202 & A201;
  assign \new_[81996]_  = \new_[81995]_  & \new_[81992]_ ;
  assign \new_[81997]_  = \new_[81996]_  & \new_[81989]_ ;
  assign \new_[82000]_  = ~A234 & ~A233;
  assign \new_[82003]_  = A266 & A265;
  assign \new_[82004]_  = \new_[82003]_  & \new_[82000]_ ;
  assign \new_[82007]_  = ~A299 & A298;
  assign \new_[82010]_  = A301 & A300;
  assign \new_[82011]_  = \new_[82010]_  & \new_[82007]_ ;
  assign \new_[82012]_  = \new_[82011]_  & \new_[82004]_ ;
  assign \new_[82015]_  = ~A168 & ~A169;
  assign \new_[82018]_  = A166 & A167;
  assign \new_[82019]_  = \new_[82018]_  & \new_[82015]_ ;
  assign \new_[82022]_  = ~A200 & A199;
  assign \new_[82025]_  = A202 & A201;
  assign \new_[82026]_  = \new_[82025]_  & \new_[82022]_ ;
  assign \new_[82027]_  = \new_[82026]_  & \new_[82019]_ ;
  assign \new_[82030]_  = ~A234 & ~A233;
  assign \new_[82033]_  = A266 & A265;
  assign \new_[82034]_  = \new_[82033]_  & \new_[82030]_ ;
  assign \new_[82037]_  = ~A299 & A298;
  assign \new_[82040]_  = A302 & A300;
  assign \new_[82041]_  = \new_[82040]_  & \new_[82037]_ ;
  assign \new_[82042]_  = \new_[82041]_  & \new_[82034]_ ;
  assign \new_[82045]_  = ~A168 & ~A169;
  assign \new_[82048]_  = A166 & A167;
  assign \new_[82049]_  = \new_[82048]_  & \new_[82045]_ ;
  assign \new_[82052]_  = ~A200 & A199;
  assign \new_[82055]_  = A202 & A201;
  assign \new_[82056]_  = \new_[82055]_  & \new_[82052]_ ;
  assign \new_[82057]_  = \new_[82056]_  & \new_[82049]_ ;
  assign \new_[82060]_  = ~A234 & ~A233;
  assign \new_[82063]_  = ~A267 & ~A266;
  assign \new_[82064]_  = \new_[82063]_  & \new_[82060]_ ;
  assign \new_[82067]_  = ~A299 & A298;
  assign \new_[82070]_  = A301 & A300;
  assign \new_[82071]_  = \new_[82070]_  & \new_[82067]_ ;
  assign \new_[82072]_  = \new_[82071]_  & \new_[82064]_ ;
  assign \new_[82075]_  = ~A168 & ~A169;
  assign \new_[82078]_  = A166 & A167;
  assign \new_[82079]_  = \new_[82078]_  & \new_[82075]_ ;
  assign \new_[82082]_  = ~A200 & A199;
  assign \new_[82085]_  = A202 & A201;
  assign \new_[82086]_  = \new_[82085]_  & \new_[82082]_ ;
  assign \new_[82087]_  = \new_[82086]_  & \new_[82079]_ ;
  assign \new_[82090]_  = ~A234 & ~A233;
  assign \new_[82093]_  = ~A267 & ~A266;
  assign \new_[82094]_  = \new_[82093]_  & \new_[82090]_ ;
  assign \new_[82097]_  = ~A299 & A298;
  assign \new_[82100]_  = A302 & A300;
  assign \new_[82101]_  = \new_[82100]_  & \new_[82097]_ ;
  assign \new_[82102]_  = \new_[82101]_  & \new_[82094]_ ;
  assign \new_[82105]_  = ~A168 & ~A169;
  assign \new_[82108]_  = A166 & A167;
  assign \new_[82109]_  = \new_[82108]_  & \new_[82105]_ ;
  assign \new_[82112]_  = ~A200 & A199;
  assign \new_[82115]_  = A202 & A201;
  assign \new_[82116]_  = \new_[82115]_  & \new_[82112]_ ;
  assign \new_[82117]_  = \new_[82116]_  & \new_[82109]_ ;
  assign \new_[82120]_  = ~A234 & ~A233;
  assign \new_[82123]_  = ~A266 & ~A265;
  assign \new_[82124]_  = \new_[82123]_  & \new_[82120]_ ;
  assign \new_[82127]_  = ~A299 & A298;
  assign \new_[82130]_  = A301 & A300;
  assign \new_[82131]_  = \new_[82130]_  & \new_[82127]_ ;
  assign \new_[82132]_  = \new_[82131]_  & \new_[82124]_ ;
  assign \new_[82135]_  = ~A168 & ~A169;
  assign \new_[82138]_  = A166 & A167;
  assign \new_[82139]_  = \new_[82138]_  & \new_[82135]_ ;
  assign \new_[82142]_  = ~A200 & A199;
  assign \new_[82145]_  = A202 & A201;
  assign \new_[82146]_  = \new_[82145]_  & \new_[82142]_ ;
  assign \new_[82147]_  = \new_[82146]_  & \new_[82139]_ ;
  assign \new_[82150]_  = ~A234 & ~A233;
  assign \new_[82153]_  = ~A266 & ~A265;
  assign \new_[82154]_  = \new_[82153]_  & \new_[82150]_ ;
  assign \new_[82157]_  = ~A299 & A298;
  assign \new_[82160]_  = A302 & A300;
  assign \new_[82161]_  = \new_[82160]_  & \new_[82157]_ ;
  assign \new_[82162]_  = \new_[82161]_  & \new_[82154]_ ;
  assign \new_[82165]_  = ~A168 & ~A169;
  assign \new_[82168]_  = A166 & A167;
  assign \new_[82169]_  = \new_[82168]_  & \new_[82165]_ ;
  assign \new_[82172]_  = ~A200 & A199;
  assign \new_[82175]_  = A202 & A201;
  assign \new_[82176]_  = \new_[82175]_  & \new_[82172]_ ;
  assign \new_[82177]_  = \new_[82176]_  & \new_[82169]_ ;
  assign \new_[82180]_  = ~A233 & A232;
  assign \new_[82183]_  = A235 & A234;
  assign \new_[82184]_  = \new_[82183]_  & \new_[82180]_ ;
  assign \new_[82187]_  = ~A266 & A265;
  assign \new_[82190]_  = A268 & A267;
  assign \new_[82191]_  = \new_[82190]_  & \new_[82187]_ ;
  assign \new_[82192]_  = \new_[82191]_  & \new_[82184]_ ;
  assign \new_[82195]_  = ~A168 & ~A169;
  assign \new_[82198]_  = A166 & A167;
  assign \new_[82199]_  = \new_[82198]_  & \new_[82195]_ ;
  assign \new_[82202]_  = ~A200 & A199;
  assign \new_[82205]_  = A202 & A201;
  assign \new_[82206]_  = \new_[82205]_  & \new_[82202]_ ;
  assign \new_[82207]_  = \new_[82206]_  & \new_[82199]_ ;
  assign \new_[82210]_  = ~A233 & A232;
  assign \new_[82213]_  = A235 & A234;
  assign \new_[82214]_  = \new_[82213]_  & \new_[82210]_ ;
  assign \new_[82217]_  = ~A266 & A265;
  assign \new_[82220]_  = A269 & A267;
  assign \new_[82221]_  = \new_[82220]_  & \new_[82217]_ ;
  assign \new_[82222]_  = \new_[82221]_  & \new_[82214]_ ;
  assign \new_[82225]_  = ~A168 & ~A169;
  assign \new_[82228]_  = A166 & A167;
  assign \new_[82229]_  = \new_[82228]_  & \new_[82225]_ ;
  assign \new_[82232]_  = ~A200 & A199;
  assign \new_[82235]_  = A202 & A201;
  assign \new_[82236]_  = \new_[82235]_  & \new_[82232]_ ;
  assign \new_[82237]_  = \new_[82236]_  & \new_[82229]_ ;
  assign \new_[82240]_  = ~A233 & A232;
  assign \new_[82243]_  = A236 & A234;
  assign \new_[82244]_  = \new_[82243]_  & \new_[82240]_ ;
  assign \new_[82247]_  = ~A266 & A265;
  assign \new_[82250]_  = A268 & A267;
  assign \new_[82251]_  = \new_[82250]_  & \new_[82247]_ ;
  assign \new_[82252]_  = \new_[82251]_  & \new_[82244]_ ;
  assign \new_[82255]_  = ~A168 & ~A169;
  assign \new_[82258]_  = A166 & A167;
  assign \new_[82259]_  = \new_[82258]_  & \new_[82255]_ ;
  assign \new_[82262]_  = ~A200 & A199;
  assign \new_[82265]_  = A202 & A201;
  assign \new_[82266]_  = \new_[82265]_  & \new_[82262]_ ;
  assign \new_[82267]_  = \new_[82266]_  & \new_[82259]_ ;
  assign \new_[82270]_  = ~A233 & A232;
  assign \new_[82273]_  = A236 & A234;
  assign \new_[82274]_  = \new_[82273]_  & \new_[82270]_ ;
  assign \new_[82277]_  = ~A266 & A265;
  assign \new_[82280]_  = A269 & A267;
  assign \new_[82281]_  = \new_[82280]_  & \new_[82277]_ ;
  assign \new_[82282]_  = \new_[82281]_  & \new_[82274]_ ;
  assign \new_[82285]_  = ~A168 & ~A169;
  assign \new_[82288]_  = A166 & A167;
  assign \new_[82289]_  = \new_[82288]_  & \new_[82285]_ ;
  assign \new_[82292]_  = ~A200 & A199;
  assign \new_[82295]_  = A202 & A201;
  assign \new_[82296]_  = \new_[82295]_  & \new_[82292]_ ;
  assign \new_[82297]_  = \new_[82296]_  & \new_[82289]_ ;
  assign \new_[82300]_  = ~A233 & ~A232;
  assign \new_[82303]_  = A266 & A265;
  assign \new_[82304]_  = \new_[82303]_  & \new_[82300]_ ;
  assign \new_[82307]_  = ~A299 & A298;
  assign \new_[82310]_  = A301 & A300;
  assign \new_[82311]_  = \new_[82310]_  & \new_[82307]_ ;
  assign \new_[82312]_  = \new_[82311]_  & \new_[82304]_ ;
  assign \new_[82315]_  = ~A168 & ~A169;
  assign \new_[82318]_  = A166 & A167;
  assign \new_[82319]_  = \new_[82318]_  & \new_[82315]_ ;
  assign \new_[82322]_  = ~A200 & A199;
  assign \new_[82325]_  = A202 & A201;
  assign \new_[82326]_  = \new_[82325]_  & \new_[82322]_ ;
  assign \new_[82327]_  = \new_[82326]_  & \new_[82319]_ ;
  assign \new_[82330]_  = ~A233 & ~A232;
  assign \new_[82333]_  = A266 & A265;
  assign \new_[82334]_  = \new_[82333]_  & \new_[82330]_ ;
  assign \new_[82337]_  = ~A299 & A298;
  assign \new_[82340]_  = A302 & A300;
  assign \new_[82341]_  = \new_[82340]_  & \new_[82337]_ ;
  assign \new_[82342]_  = \new_[82341]_  & \new_[82334]_ ;
  assign \new_[82345]_  = ~A168 & ~A169;
  assign \new_[82348]_  = A166 & A167;
  assign \new_[82349]_  = \new_[82348]_  & \new_[82345]_ ;
  assign \new_[82352]_  = ~A200 & A199;
  assign \new_[82355]_  = A202 & A201;
  assign \new_[82356]_  = \new_[82355]_  & \new_[82352]_ ;
  assign \new_[82357]_  = \new_[82356]_  & \new_[82349]_ ;
  assign \new_[82360]_  = ~A233 & ~A232;
  assign \new_[82363]_  = ~A267 & ~A266;
  assign \new_[82364]_  = \new_[82363]_  & \new_[82360]_ ;
  assign \new_[82367]_  = ~A299 & A298;
  assign \new_[82370]_  = A301 & A300;
  assign \new_[82371]_  = \new_[82370]_  & \new_[82367]_ ;
  assign \new_[82372]_  = \new_[82371]_  & \new_[82364]_ ;
  assign \new_[82375]_  = ~A168 & ~A169;
  assign \new_[82378]_  = A166 & A167;
  assign \new_[82379]_  = \new_[82378]_  & \new_[82375]_ ;
  assign \new_[82382]_  = ~A200 & A199;
  assign \new_[82385]_  = A202 & A201;
  assign \new_[82386]_  = \new_[82385]_  & \new_[82382]_ ;
  assign \new_[82387]_  = \new_[82386]_  & \new_[82379]_ ;
  assign \new_[82390]_  = ~A233 & ~A232;
  assign \new_[82393]_  = ~A267 & ~A266;
  assign \new_[82394]_  = \new_[82393]_  & \new_[82390]_ ;
  assign \new_[82397]_  = ~A299 & A298;
  assign \new_[82400]_  = A302 & A300;
  assign \new_[82401]_  = \new_[82400]_  & \new_[82397]_ ;
  assign \new_[82402]_  = \new_[82401]_  & \new_[82394]_ ;
  assign \new_[82405]_  = ~A168 & ~A169;
  assign \new_[82408]_  = A166 & A167;
  assign \new_[82409]_  = \new_[82408]_  & \new_[82405]_ ;
  assign \new_[82412]_  = ~A200 & A199;
  assign \new_[82415]_  = A202 & A201;
  assign \new_[82416]_  = \new_[82415]_  & \new_[82412]_ ;
  assign \new_[82417]_  = \new_[82416]_  & \new_[82409]_ ;
  assign \new_[82420]_  = ~A233 & ~A232;
  assign \new_[82423]_  = ~A266 & ~A265;
  assign \new_[82424]_  = \new_[82423]_  & \new_[82420]_ ;
  assign \new_[82427]_  = ~A299 & A298;
  assign \new_[82430]_  = A301 & A300;
  assign \new_[82431]_  = \new_[82430]_  & \new_[82427]_ ;
  assign \new_[82432]_  = \new_[82431]_  & \new_[82424]_ ;
  assign \new_[82435]_  = ~A168 & ~A169;
  assign \new_[82438]_  = A166 & A167;
  assign \new_[82439]_  = \new_[82438]_  & \new_[82435]_ ;
  assign \new_[82442]_  = ~A200 & A199;
  assign \new_[82445]_  = A202 & A201;
  assign \new_[82446]_  = \new_[82445]_  & \new_[82442]_ ;
  assign \new_[82447]_  = \new_[82446]_  & \new_[82439]_ ;
  assign \new_[82450]_  = ~A233 & ~A232;
  assign \new_[82453]_  = ~A266 & ~A265;
  assign \new_[82454]_  = \new_[82453]_  & \new_[82450]_ ;
  assign \new_[82457]_  = ~A299 & A298;
  assign \new_[82460]_  = A302 & A300;
  assign \new_[82461]_  = \new_[82460]_  & \new_[82457]_ ;
  assign \new_[82462]_  = \new_[82461]_  & \new_[82454]_ ;
  assign \new_[82465]_  = ~A168 & ~A169;
  assign \new_[82468]_  = A166 & A167;
  assign \new_[82469]_  = \new_[82468]_  & \new_[82465]_ ;
  assign \new_[82472]_  = ~A200 & A199;
  assign \new_[82475]_  = A203 & A201;
  assign \new_[82476]_  = \new_[82475]_  & \new_[82472]_ ;
  assign \new_[82477]_  = \new_[82476]_  & \new_[82469]_ ;
  assign \new_[82480]_  = A233 & A232;
  assign \new_[82483]_  = ~A267 & A265;
  assign \new_[82484]_  = \new_[82483]_  & \new_[82480]_ ;
  assign \new_[82487]_  = ~A299 & A298;
  assign \new_[82490]_  = A301 & A300;
  assign \new_[82491]_  = \new_[82490]_  & \new_[82487]_ ;
  assign \new_[82492]_  = \new_[82491]_  & \new_[82484]_ ;
  assign \new_[82495]_  = ~A168 & ~A169;
  assign \new_[82498]_  = A166 & A167;
  assign \new_[82499]_  = \new_[82498]_  & \new_[82495]_ ;
  assign \new_[82502]_  = ~A200 & A199;
  assign \new_[82505]_  = A203 & A201;
  assign \new_[82506]_  = \new_[82505]_  & \new_[82502]_ ;
  assign \new_[82507]_  = \new_[82506]_  & \new_[82499]_ ;
  assign \new_[82510]_  = A233 & A232;
  assign \new_[82513]_  = ~A267 & A265;
  assign \new_[82514]_  = \new_[82513]_  & \new_[82510]_ ;
  assign \new_[82517]_  = ~A299 & A298;
  assign \new_[82520]_  = A302 & A300;
  assign \new_[82521]_  = \new_[82520]_  & \new_[82517]_ ;
  assign \new_[82522]_  = \new_[82521]_  & \new_[82514]_ ;
  assign \new_[82525]_  = ~A168 & ~A169;
  assign \new_[82528]_  = A166 & A167;
  assign \new_[82529]_  = \new_[82528]_  & \new_[82525]_ ;
  assign \new_[82532]_  = ~A200 & A199;
  assign \new_[82535]_  = A203 & A201;
  assign \new_[82536]_  = \new_[82535]_  & \new_[82532]_ ;
  assign \new_[82537]_  = \new_[82536]_  & \new_[82529]_ ;
  assign \new_[82540]_  = A233 & A232;
  assign \new_[82543]_  = A266 & A265;
  assign \new_[82544]_  = \new_[82543]_  & \new_[82540]_ ;
  assign \new_[82547]_  = ~A299 & A298;
  assign \new_[82550]_  = A301 & A300;
  assign \new_[82551]_  = \new_[82550]_  & \new_[82547]_ ;
  assign \new_[82552]_  = \new_[82551]_  & \new_[82544]_ ;
  assign \new_[82555]_  = ~A168 & ~A169;
  assign \new_[82558]_  = A166 & A167;
  assign \new_[82559]_  = \new_[82558]_  & \new_[82555]_ ;
  assign \new_[82562]_  = ~A200 & A199;
  assign \new_[82565]_  = A203 & A201;
  assign \new_[82566]_  = \new_[82565]_  & \new_[82562]_ ;
  assign \new_[82567]_  = \new_[82566]_  & \new_[82559]_ ;
  assign \new_[82570]_  = A233 & A232;
  assign \new_[82573]_  = A266 & A265;
  assign \new_[82574]_  = \new_[82573]_  & \new_[82570]_ ;
  assign \new_[82577]_  = ~A299 & A298;
  assign \new_[82580]_  = A302 & A300;
  assign \new_[82581]_  = \new_[82580]_  & \new_[82577]_ ;
  assign \new_[82582]_  = \new_[82581]_  & \new_[82574]_ ;
  assign \new_[82585]_  = ~A168 & ~A169;
  assign \new_[82588]_  = A166 & A167;
  assign \new_[82589]_  = \new_[82588]_  & \new_[82585]_ ;
  assign \new_[82592]_  = ~A200 & A199;
  assign \new_[82595]_  = A203 & A201;
  assign \new_[82596]_  = \new_[82595]_  & \new_[82592]_ ;
  assign \new_[82597]_  = \new_[82596]_  & \new_[82589]_ ;
  assign \new_[82600]_  = A233 & A232;
  assign \new_[82603]_  = ~A266 & ~A265;
  assign \new_[82604]_  = \new_[82603]_  & \new_[82600]_ ;
  assign \new_[82607]_  = ~A299 & A298;
  assign \new_[82610]_  = A301 & A300;
  assign \new_[82611]_  = \new_[82610]_  & \new_[82607]_ ;
  assign \new_[82612]_  = \new_[82611]_  & \new_[82604]_ ;
  assign \new_[82615]_  = ~A168 & ~A169;
  assign \new_[82618]_  = A166 & A167;
  assign \new_[82619]_  = \new_[82618]_  & \new_[82615]_ ;
  assign \new_[82622]_  = ~A200 & A199;
  assign \new_[82625]_  = A203 & A201;
  assign \new_[82626]_  = \new_[82625]_  & \new_[82622]_ ;
  assign \new_[82627]_  = \new_[82626]_  & \new_[82619]_ ;
  assign \new_[82630]_  = A233 & A232;
  assign \new_[82633]_  = ~A266 & ~A265;
  assign \new_[82634]_  = \new_[82633]_  & \new_[82630]_ ;
  assign \new_[82637]_  = ~A299 & A298;
  assign \new_[82640]_  = A302 & A300;
  assign \new_[82641]_  = \new_[82640]_  & \new_[82637]_ ;
  assign \new_[82642]_  = \new_[82641]_  & \new_[82634]_ ;
  assign \new_[82645]_  = ~A168 & ~A169;
  assign \new_[82648]_  = A166 & A167;
  assign \new_[82649]_  = \new_[82648]_  & \new_[82645]_ ;
  assign \new_[82652]_  = ~A200 & A199;
  assign \new_[82655]_  = A203 & A201;
  assign \new_[82656]_  = \new_[82655]_  & \new_[82652]_ ;
  assign \new_[82657]_  = \new_[82656]_  & \new_[82649]_ ;
  assign \new_[82660]_  = ~A235 & ~A233;
  assign \new_[82663]_  = ~A266 & ~A236;
  assign \new_[82664]_  = \new_[82663]_  & \new_[82660]_ ;
  assign \new_[82667]_  = ~A269 & ~A268;
  assign \new_[82670]_  = A299 & ~A298;
  assign \new_[82671]_  = \new_[82670]_  & \new_[82667]_ ;
  assign \new_[82672]_  = \new_[82671]_  & \new_[82664]_ ;
  assign \new_[82675]_  = ~A168 & ~A169;
  assign \new_[82678]_  = A166 & A167;
  assign \new_[82679]_  = \new_[82678]_  & \new_[82675]_ ;
  assign \new_[82682]_  = ~A200 & A199;
  assign \new_[82685]_  = A203 & A201;
  assign \new_[82686]_  = \new_[82685]_  & \new_[82682]_ ;
  assign \new_[82687]_  = \new_[82686]_  & \new_[82679]_ ;
  assign \new_[82690]_  = ~A234 & ~A233;
  assign \new_[82693]_  = A266 & A265;
  assign \new_[82694]_  = \new_[82693]_  & \new_[82690]_ ;
  assign \new_[82697]_  = ~A299 & A298;
  assign \new_[82700]_  = A301 & A300;
  assign \new_[82701]_  = \new_[82700]_  & \new_[82697]_ ;
  assign \new_[82702]_  = \new_[82701]_  & \new_[82694]_ ;
  assign \new_[82705]_  = ~A168 & ~A169;
  assign \new_[82708]_  = A166 & A167;
  assign \new_[82709]_  = \new_[82708]_  & \new_[82705]_ ;
  assign \new_[82712]_  = ~A200 & A199;
  assign \new_[82715]_  = A203 & A201;
  assign \new_[82716]_  = \new_[82715]_  & \new_[82712]_ ;
  assign \new_[82717]_  = \new_[82716]_  & \new_[82709]_ ;
  assign \new_[82720]_  = ~A234 & ~A233;
  assign \new_[82723]_  = A266 & A265;
  assign \new_[82724]_  = \new_[82723]_  & \new_[82720]_ ;
  assign \new_[82727]_  = ~A299 & A298;
  assign \new_[82730]_  = A302 & A300;
  assign \new_[82731]_  = \new_[82730]_  & \new_[82727]_ ;
  assign \new_[82732]_  = \new_[82731]_  & \new_[82724]_ ;
  assign \new_[82735]_  = ~A168 & ~A169;
  assign \new_[82738]_  = A166 & A167;
  assign \new_[82739]_  = \new_[82738]_  & \new_[82735]_ ;
  assign \new_[82742]_  = ~A200 & A199;
  assign \new_[82745]_  = A203 & A201;
  assign \new_[82746]_  = \new_[82745]_  & \new_[82742]_ ;
  assign \new_[82747]_  = \new_[82746]_  & \new_[82739]_ ;
  assign \new_[82750]_  = ~A234 & ~A233;
  assign \new_[82753]_  = ~A267 & ~A266;
  assign \new_[82754]_  = \new_[82753]_  & \new_[82750]_ ;
  assign \new_[82757]_  = ~A299 & A298;
  assign \new_[82760]_  = A301 & A300;
  assign \new_[82761]_  = \new_[82760]_  & \new_[82757]_ ;
  assign \new_[82762]_  = \new_[82761]_  & \new_[82754]_ ;
  assign \new_[82765]_  = ~A168 & ~A169;
  assign \new_[82768]_  = A166 & A167;
  assign \new_[82769]_  = \new_[82768]_  & \new_[82765]_ ;
  assign \new_[82772]_  = ~A200 & A199;
  assign \new_[82775]_  = A203 & A201;
  assign \new_[82776]_  = \new_[82775]_  & \new_[82772]_ ;
  assign \new_[82777]_  = \new_[82776]_  & \new_[82769]_ ;
  assign \new_[82780]_  = ~A234 & ~A233;
  assign \new_[82783]_  = ~A267 & ~A266;
  assign \new_[82784]_  = \new_[82783]_  & \new_[82780]_ ;
  assign \new_[82787]_  = ~A299 & A298;
  assign \new_[82790]_  = A302 & A300;
  assign \new_[82791]_  = \new_[82790]_  & \new_[82787]_ ;
  assign \new_[82792]_  = \new_[82791]_  & \new_[82784]_ ;
  assign \new_[82795]_  = ~A168 & ~A169;
  assign \new_[82798]_  = A166 & A167;
  assign \new_[82799]_  = \new_[82798]_  & \new_[82795]_ ;
  assign \new_[82802]_  = ~A200 & A199;
  assign \new_[82805]_  = A203 & A201;
  assign \new_[82806]_  = \new_[82805]_  & \new_[82802]_ ;
  assign \new_[82807]_  = \new_[82806]_  & \new_[82799]_ ;
  assign \new_[82810]_  = ~A234 & ~A233;
  assign \new_[82813]_  = ~A266 & ~A265;
  assign \new_[82814]_  = \new_[82813]_  & \new_[82810]_ ;
  assign \new_[82817]_  = ~A299 & A298;
  assign \new_[82820]_  = A301 & A300;
  assign \new_[82821]_  = \new_[82820]_  & \new_[82817]_ ;
  assign \new_[82822]_  = \new_[82821]_  & \new_[82814]_ ;
  assign \new_[82825]_  = ~A168 & ~A169;
  assign \new_[82828]_  = A166 & A167;
  assign \new_[82829]_  = \new_[82828]_  & \new_[82825]_ ;
  assign \new_[82832]_  = ~A200 & A199;
  assign \new_[82835]_  = A203 & A201;
  assign \new_[82836]_  = \new_[82835]_  & \new_[82832]_ ;
  assign \new_[82837]_  = \new_[82836]_  & \new_[82829]_ ;
  assign \new_[82840]_  = ~A234 & ~A233;
  assign \new_[82843]_  = ~A266 & ~A265;
  assign \new_[82844]_  = \new_[82843]_  & \new_[82840]_ ;
  assign \new_[82847]_  = ~A299 & A298;
  assign \new_[82850]_  = A302 & A300;
  assign \new_[82851]_  = \new_[82850]_  & \new_[82847]_ ;
  assign \new_[82852]_  = \new_[82851]_  & \new_[82844]_ ;
  assign \new_[82855]_  = ~A168 & ~A169;
  assign \new_[82858]_  = A166 & A167;
  assign \new_[82859]_  = \new_[82858]_  & \new_[82855]_ ;
  assign \new_[82862]_  = ~A200 & A199;
  assign \new_[82865]_  = A203 & A201;
  assign \new_[82866]_  = \new_[82865]_  & \new_[82862]_ ;
  assign \new_[82867]_  = \new_[82866]_  & \new_[82859]_ ;
  assign \new_[82870]_  = ~A233 & A232;
  assign \new_[82873]_  = A235 & A234;
  assign \new_[82874]_  = \new_[82873]_  & \new_[82870]_ ;
  assign \new_[82877]_  = ~A266 & A265;
  assign \new_[82880]_  = A268 & A267;
  assign \new_[82881]_  = \new_[82880]_  & \new_[82877]_ ;
  assign \new_[82882]_  = \new_[82881]_  & \new_[82874]_ ;
  assign \new_[82885]_  = ~A168 & ~A169;
  assign \new_[82888]_  = A166 & A167;
  assign \new_[82889]_  = \new_[82888]_  & \new_[82885]_ ;
  assign \new_[82892]_  = ~A200 & A199;
  assign \new_[82895]_  = A203 & A201;
  assign \new_[82896]_  = \new_[82895]_  & \new_[82892]_ ;
  assign \new_[82897]_  = \new_[82896]_  & \new_[82889]_ ;
  assign \new_[82900]_  = ~A233 & A232;
  assign \new_[82903]_  = A235 & A234;
  assign \new_[82904]_  = \new_[82903]_  & \new_[82900]_ ;
  assign \new_[82907]_  = ~A266 & A265;
  assign \new_[82910]_  = A269 & A267;
  assign \new_[82911]_  = \new_[82910]_  & \new_[82907]_ ;
  assign \new_[82912]_  = \new_[82911]_  & \new_[82904]_ ;
  assign \new_[82915]_  = ~A168 & ~A169;
  assign \new_[82918]_  = A166 & A167;
  assign \new_[82919]_  = \new_[82918]_  & \new_[82915]_ ;
  assign \new_[82922]_  = ~A200 & A199;
  assign \new_[82925]_  = A203 & A201;
  assign \new_[82926]_  = \new_[82925]_  & \new_[82922]_ ;
  assign \new_[82927]_  = \new_[82926]_  & \new_[82919]_ ;
  assign \new_[82930]_  = ~A233 & A232;
  assign \new_[82933]_  = A236 & A234;
  assign \new_[82934]_  = \new_[82933]_  & \new_[82930]_ ;
  assign \new_[82937]_  = ~A266 & A265;
  assign \new_[82940]_  = A268 & A267;
  assign \new_[82941]_  = \new_[82940]_  & \new_[82937]_ ;
  assign \new_[82942]_  = \new_[82941]_  & \new_[82934]_ ;
  assign \new_[82945]_  = ~A168 & ~A169;
  assign \new_[82948]_  = A166 & A167;
  assign \new_[82949]_  = \new_[82948]_  & \new_[82945]_ ;
  assign \new_[82952]_  = ~A200 & A199;
  assign \new_[82955]_  = A203 & A201;
  assign \new_[82956]_  = \new_[82955]_  & \new_[82952]_ ;
  assign \new_[82957]_  = \new_[82956]_  & \new_[82949]_ ;
  assign \new_[82960]_  = ~A233 & A232;
  assign \new_[82963]_  = A236 & A234;
  assign \new_[82964]_  = \new_[82963]_  & \new_[82960]_ ;
  assign \new_[82967]_  = ~A266 & A265;
  assign \new_[82970]_  = A269 & A267;
  assign \new_[82971]_  = \new_[82970]_  & \new_[82967]_ ;
  assign \new_[82972]_  = \new_[82971]_  & \new_[82964]_ ;
  assign \new_[82975]_  = ~A168 & ~A169;
  assign \new_[82978]_  = A166 & A167;
  assign \new_[82979]_  = \new_[82978]_  & \new_[82975]_ ;
  assign \new_[82982]_  = ~A200 & A199;
  assign \new_[82985]_  = A203 & A201;
  assign \new_[82986]_  = \new_[82985]_  & \new_[82982]_ ;
  assign \new_[82987]_  = \new_[82986]_  & \new_[82979]_ ;
  assign \new_[82990]_  = ~A233 & ~A232;
  assign \new_[82993]_  = A266 & A265;
  assign \new_[82994]_  = \new_[82993]_  & \new_[82990]_ ;
  assign \new_[82997]_  = ~A299 & A298;
  assign \new_[83000]_  = A301 & A300;
  assign \new_[83001]_  = \new_[83000]_  & \new_[82997]_ ;
  assign \new_[83002]_  = \new_[83001]_  & \new_[82994]_ ;
  assign \new_[83005]_  = ~A168 & ~A169;
  assign \new_[83008]_  = A166 & A167;
  assign \new_[83009]_  = \new_[83008]_  & \new_[83005]_ ;
  assign \new_[83012]_  = ~A200 & A199;
  assign \new_[83015]_  = A203 & A201;
  assign \new_[83016]_  = \new_[83015]_  & \new_[83012]_ ;
  assign \new_[83017]_  = \new_[83016]_  & \new_[83009]_ ;
  assign \new_[83020]_  = ~A233 & ~A232;
  assign \new_[83023]_  = A266 & A265;
  assign \new_[83024]_  = \new_[83023]_  & \new_[83020]_ ;
  assign \new_[83027]_  = ~A299 & A298;
  assign \new_[83030]_  = A302 & A300;
  assign \new_[83031]_  = \new_[83030]_  & \new_[83027]_ ;
  assign \new_[83032]_  = \new_[83031]_  & \new_[83024]_ ;
  assign \new_[83035]_  = ~A168 & ~A169;
  assign \new_[83038]_  = A166 & A167;
  assign \new_[83039]_  = \new_[83038]_  & \new_[83035]_ ;
  assign \new_[83042]_  = ~A200 & A199;
  assign \new_[83045]_  = A203 & A201;
  assign \new_[83046]_  = \new_[83045]_  & \new_[83042]_ ;
  assign \new_[83047]_  = \new_[83046]_  & \new_[83039]_ ;
  assign \new_[83050]_  = ~A233 & ~A232;
  assign \new_[83053]_  = ~A267 & ~A266;
  assign \new_[83054]_  = \new_[83053]_  & \new_[83050]_ ;
  assign \new_[83057]_  = ~A299 & A298;
  assign \new_[83060]_  = A301 & A300;
  assign \new_[83061]_  = \new_[83060]_  & \new_[83057]_ ;
  assign \new_[83062]_  = \new_[83061]_  & \new_[83054]_ ;
  assign \new_[83065]_  = ~A168 & ~A169;
  assign \new_[83068]_  = A166 & A167;
  assign \new_[83069]_  = \new_[83068]_  & \new_[83065]_ ;
  assign \new_[83072]_  = ~A200 & A199;
  assign \new_[83075]_  = A203 & A201;
  assign \new_[83076]_  = \new_[83075]_  & \new_[83072]_ ;
  assign \new_[83077]_  = \new_[83076]_  & \new_[83069]_ ;
  assign \new_[83080]_  = ~A233 & ~A232;
  assign \new_[83083]_  = ~A267 & ~A266;
  assign \new_[83084]_  = \new_[83083]_  & \new_[83080]_ ;
  assign \new_[83087]_  = ~A299 & A298;
  assign \new_[83090]_  = A302 & A300;
  assign \new_[83091]_  = \new_[83090]_  & \new_[83087]_ ;
  assign \new_[83092]_  = \new_[83091]_  & \new_[83084]_ ;
  assign \new_[83095]_  = ~A168 & ~A169;
  assign \new_[83098]_  = A166 & A167;
  assign \new_[83099]_  = \new_[83098]_  & \new_[83095]_ ;
  assign \new_[83102]_  = ~A200 & A199;
  assign \new_[83105]_  = A203 & A201;
  assign \new_[83106]_  = \new_[83105]_  & \new_[83102]_ ;
  assign \new_[83107]_  = \new_[83106]_  & \new_[83099]_ ;
  assign \new_[83110]_  = ~A233 & ~A232;
  assign \new_[83113]_  = ~A266 & ~A265;
  assign \new_[83114]_  = \new_[83113]_  & \new_[83110]_ ;
  assign \new_[83117]_  = ~A299 & A298;
  assign \new_[83120]_  = A301 & A300;
  assign \new_[83121]_  = \new_[83120]_  & \new_[83117]_ ;
  assign \new_[83122]_  = \new_[83121]_  & \new_[83114]_ ;
  assign \new_[83125]_  = ~A168 & ~A169;
  assign \new_[83128]_  = A166 & A167;
  assign \new_[83129]_  = \new_[83128]_  & \new_[83125]_ ;
  assign \new_[83132]_  = ~A200 & A199;
  assign \new_[83135]_  = A203 & A201;
  assign \new_[83136]_  = \new_[83135]_  & \new_[83132]_ ;
  assign \new_[83137]_  = \new_[83136]_  & \new_[83129]_ ;
  assign \new_[83140]_  = ~A233 & ~A232;
  assign \new_[83143]_  = ~A266 & ~A265;
  assign \new_[83144]_  = \new_[83143]_  & \new_[83140]_ ;
  assign \new_[83147]_  = ~A299 & A298;
  assign \new_[83150]_  = A302 & A300;
  assign \new_[83151]_  = \new_[83150]_  & \new_[83147]_ ;
  assign \new_[83152]_  = \new_[83151]_  & \new_[83144]_ ;
  assign \new_[83155]_  = ~A169 & A170;
  assign \new_[83158]_  = ~A166 & A167;
  assign \new_[83159]_  = \new_[83158]_  & \new_[83155]_ ;
  assign \new_[83162]_  = A200 & A199;
  assign \new_[83165]_  = ~A235 & ~A233;
  assign \new_[83166]_  = \new_[83165]_  & \new_[83162]_ ;
  assign \new_[83167]_  = \new_[83166]_  & \new_[83159]_ ;
  assign \new_[83170]_  = ~A266 & ~A236;
  assign \new_[83173]_  = ~A269 & ~A268;
  assign \new_[83174]_  = \new_[83173]_  & \new_[83170]_ ;
  assign \new_[83177]_  = ~A299 & A298;
  assign \new_[83180]_  = A301 & A300;
  assign \new_[83181]_  = \new_[83180]_  & \new_[83177]_ ;
  assign \new_[83182]_  = \new_[83181]_  & \new_[83174]_ ;
  assign \new_[83185]_  = ~A169 & A170;
  assign \new_[83188]_  = ~A166 & A167;
  assign \new_[83189]_  = \new_[83188]_  & \new_[83185]_ ;
  assign \new_[83192]_  = A200 & A199;
  assign \new_[83195]_  = ~A235 & ~A233;
  assign \new_[83196]_  = \new_[83195]_  & \new_[83192]_ ;
  assign \new_[83197]_  = \new_[83196]_  & \new_[83189]_ ;
  assign \new_[83200]_  = ~A266 & ~A236;
  assign \new_[83203]_  = ~A269 & ~A268;
  assign \new_[83204]_  = \new_[83203]_  & \new_[83200]_ ;
  assign \new_[83207]_  = ~A299 & A298;
  assign \new_[83210]_  = A302 & A300;
  assign \new_[83211]_  = \new_[83210]_  & \new_[83207]_ ;
  assign \new_[83212]_  = \new_[83211]_  & \new_[83204]_ ;
  assign \new_[83215]_  = ~A169 & A170;
  assign \new_[83218]_  = ~A166 & A167;
  assign \new_[83219]_  = \new_[83218]_  & \new_[83215]_ ;
  assign \new_[83222]_  = ~A202 & ~A200;
  assign \new_[83225]_  = A232 & ~A203;
  assign \new_[83226]_  = \new_[83225]_  & \new_[83222]_ ;
  assign \new_[83227]_  = \new_[83226]_  & \new_[83219]_ ;
  assign \new_[83230]_  = A265 & A233;
  assign \new_[83233]_  = ~A269 & ~A268;
  assign \new_[83234]_  = \new_[83233]_  & \new_[83230]_ ;
  assign \new_[83237]_  = ~A299 & A298;
  assign \new_[83240]_  = A301 & A300;
  assign \new_[83241]_  = \new_[83240]_  & \new_[83237]_ ;
  assign \new_[83242]_  = \new_[83241]_  & \new_[83234]_ ;
  assign \new_[83245]_  = ~A169 & A170;
  assign \new_[83248]_  = ~A166 & A167;
  assign \new_[83249]_  = \new_[83248]_  & \new_[83245]_ ;
  assign \new_[83252]_  = ~A202 & ~A200;
  assign \new_[83255]_  = A232 & ~A203;
  assign \new_[83256]_  = \new_[83255]_  & \new_[83252]_ ;
  assign \new_[83257]_  = \new_[83256]_  & \new_[83249]_ ;
  assign \new_[83260]_  = A265 & A233;
  assign \new_[83263]_  = ~A269 & ~A268;
  assign \new_[83264]_  = \new_[83263]_  & \new_[83260]_ ;
  assign \new_[83267]_  = ~A299 & A298;
  assign \new_[83270]_  = A302 & A300;
  assign \new_[83271]_  = \new_[83270]_  & \new_[83267]_ ;
  assign \new_[83272]_  = \new_[83271]_  & \new_[83264]_ ;
  assign \new_[83275]_  = ~A169 & A170;
  assign \new_[83278]_  = ~A166 & A167;
  assign \new_[83279]_  = \new_[83278]_  & \new_[83275]_ ;
  assign \new_[83282]_  = ~A202 & ~A200;
  assign \new_[83285]_  = ~A233 & ~A203;
  assign \new_[83286]_  = \new_[83285]_  & \new_[83282]_ ;
  assign \new_[83287]_  = \new_[83286]_  & \new_[83279]_ ;
  assign \new_[83290]_  = ~A236 & ~A235;
  assign \new_[83293]_  = A266 & A265;
  assign \new_[83294]_  = \new_[83293]_  & \new_[83290]_ ;
  assign \new_[83297]_  = ~A299 & A298;
  assign \new_[83300]_  = A301 & A300;
  assign \new_[83301]_  = \new_[83300]_  & \new_[83297]_ ;
  assign \new_[83302]_  = \new_[83301]_  & \new_[83294]_ ;
  assign \new_[83305]_  = ~A169 & A170;
  assign \new_[83308]_  = ~A166 & A167;
  assign \new_[83309]_  = \new_[83308]_  & \new_[83305]_ ;
  assign \new_[83312]_  = ~A202 & ~A200;
  assign \new_[83315]_  = ~A233 & ~A203;
  assign \new_[83316]_  = \new_[83315]_  & \new_[83312]_ ;
  assign \new_[83317]_  = \new_[83316]_  & \new_[83309]_ ;
  assign \new_[83320]_  = ~A236 & ~A235;
  assign \new_[83323]_  = A266 & A265;
  assign \new_[83324]_  = \new_[83323]_  & \new_[83320]_ ;
  assign \new_[83327]_  = ~A299 & A298;
  assign \new_[83330]_  = A302 & A300;
  assign \new_[83331]_  = \new_[83330]_  & \new_[83327]_ ;
  assign \new_[83332]_  = \new_[83331]_  & \new_[83324]_ ;
  assign \new_[83335]_  = ~A169 & A170;
  assign \new_[83338]_  = ~A166 & A167;
  assign \new_[83339]_  = \new_[83338]_  & \new_[83335]_ ;
  assign \new_[83342]_  = ~A202 & ~A200;
  assign \new_[83345]_  = ~A233 & ~A203;
  assign \new_[83346]_  = \new_[83345]_  & \new_[83342]_ ;
  assign \new_[83347]_  = \new_[83346]_  & \new_[83339]_ ;
  assign \new_[83350]_  = ~A236 & ~A235;
  assign \new_[83353]_  = ~A267 & ~A266;
  assign \new_[83354]_  = \new_[83353]_  & \new_[83350]_ ;
  assign \new_[83357]_  = ~A299 & A298;
  assign \new_[83360]_  = A301 & A300;
  assign \new_[83361]_  = \new_[83360]_  & \new_[83357]_ ;
  assign \new_[83362]_  = \new_[83361]_  & \new_[83354]_ ;
  assign \new_[83365]_  = ~A169 & A170;
  assign \new_[83368]_  = ~A166 & A167;
  assign \new_[83369]_  = \new_[83368]_  & \new_[83365]_ ;
  assign \new_[83372]_  = ~A202 & ~A200;
  assign \new_[83375]_  = ~A233 & ~A203;
  assign \new_[83376]_  = \new_[83375]_  & \new_[83372]_ ;
  assign \new_[83377]_  = \new_[83376]_  & \new_[83369]_ ;
  assign \new_[83380]_  = ~A236 & ~A235;
  assign \new_[83383]_  = ~A267 & ~A266;
  assign \new_[83384]_  = \new_[83383]_  & \new_[83380]_ ;
  assign \new_[83387]_  = ~A299 & A298;
  assign \new_[83390]_  = A302 & A300;
  assign \new_[83391]_  = \new_[83390]_  & \new_[83387]_ ;
  assign \new_[83392]_  = \new_[83391]_  & \new_[83384]_ ;
  assign \new_[83395]_  = ~A169 & A170;
  assign \new_[83398]_  = ~A166 & A167;
  assign \new_[83399]_  = \new_[83398]_  & \new_[83395]_ ;
  assign \new_[83402]_  = ~A202 & ~A200;
  assign \new_[83405]_  = ~A233 & ~A203;
  assign \new_[83406]_  = \new_[83405]_  & \new_[83402]_ ;
  assign \new_[83407]_  = \new_[83406]_  & \new_[83399]_ ;
  assign \new_[83410]_  = ~A236 & ~A235;
  assign \new_[83413]_  = ~A266 & ~A265;
  assign \new_[83414]_  = \new_[83413]_  & \new_[83410]_ ;
  assign \new_[83417]_  = ~A299 & A298;
  assign \new_[83420]_  = A301 & A300;
  assign \new_[83421]_  = \new_[83420]_  & \new_[83417]_ ;
  assign \new_[83422]_  = \new_[83421]_  & \new_[83414]_ ;
  assign \new_[83425]_  = ~A169 & A170;
  assign \new_[83428]_  = ~A166 & A167;
  assign \new_[83429]_  = \new_[83428]_  & \new_[83425]_ ;
  assign \new_[83432]_  = ~A202 & ~A200;
  assign \new_[83435]_  = ~A233 & ~A203;
  assign \new_[83436]_  = \new_[83435]_  & \new_[83432]_ ;
  assign \new_[83437]_  = \new_[83436]_  & \new_[83429]_ ;
  assign \new_[83440]_  = ~A236 & ~A235;
  assign \new_[83443]_  = ~A266 & ~A265;
  assign \new_[83444]_  = \new_[83443]_  & \new_[83440]_ ;
  assign \new_[83447]_  = ~A299 & A298;
  assign \new_[83450]_  = A302 & A300;
  assign \new_[83451]_  = \new_[83450]_  & \new_[83447]_ ;
  assign \new_[83452]_  = \new_[83451]_  & \new_[83444]_ ;
  assign \new_[83455]_  = ~A169 & A170;
  assign \new_[83458]_  = ~A166 & A167;
  assign \new_[83459]_  = \new_[83458]_  & \new_[83455]_ ;
  assign \new_[83462]_  = ~A202 & ~A200;
  assign \new_[83465]_  = ~A233 & ~A203;
  assign \new_[83466]_  = \new_[83465]_  & \new_[83462]_ ;
  assign \new_[83467]_  = \new_[83466]_  & \new_[83459]_ ;
  assign \new_[83470]_  = ~A266 & ~A234;
  assign \new_[83473]_  = ~A269 & ~A268;
  assign \new_[83474]_  = \new_[83473]_  & \new_[83470]_ ;
  assign \new_[83477]_  = ~A299 & A298;
  assign \new_[83480]_  = A301 & A300;
  assign \new_[83481]_  = \new_[83480]_  & \new_[83477]_ ;
  assign \new_[83482]_  = \new_[83481]_  & \new_[83474]_ ;
  assign \new_[83485]_  = ~A169 & A170;
  assign \new_[83488]_  = ~A166 & A167;
  assign \new_[83489]_  = \new_[83488]_  & \new_[83485]_ ;
  assign \new_[83492]_  = ~A202 & ~A200;
  assign \new_[83495]_  = ~A233 & ~A203;
  assign \new_[83496]_  = \new_[83495]_  & \new_[83492]_ ;
  assign \new_[83497]_  = \new_[83496]_  & \new_[83489]_ ;
  assign \new_[83500]_  = ~A266 & ~A234;
  assign \new_[83503]_  = ~A269 & ~A268;
  assign \new_[83504]_  = \new_[83503]_  & \new_[83500]_ ;
  assign \new_[83507]_  = ~A299 & A298;
  assign \new_[83510]_  = A302 & A300;
  assign \new_[83511]_  = \new_[83510]_  & \new_[83507]_ ;
  assign \new_[83512]_  = \new_[83511]_  & \new_[83504]_ ;
  assign \new_[83515]_  = ~A169 & A170;
  assign \new_[83518]_  = ~A166 & A167;
  assign \new_[83519]_  = \new_[83518]_  & \new_[83515]_ ;
  assign \new_[83522]_  = ~A202 & ~A200;
  assign \new_[83525]_  = ~A232 & ~A203;
  assign \new_[83526]_  = \new_[83525]_  & \new_[83522]_ ;
  assign \new_[83527]_  = \new_[83526]_  & \new_[83519]_ ;
  assign \new_[83530]_  = ~A266 & ~A233;
  assign \new_[83533]_  = ~A269 & ~A268;
  assign \new_[83534]_  = \new_[83533]_  & \new_[83530]_ ;
  assign \new_[83537]_  = ~A299 & A298;
  assign \new_[83540]_  = A301 & A300;
  assign \new_[83541]_  = \new_[83540]_  & \new_[83537]_ ;
  assign \new_[83542]_  = \new_[83541]_  & \new_[83534]_ ;
  assign \new_[83545]_  = ~A169 & A170;
  assign \new_[83548]_  = ~A166 & A167;
  assign \new_[83549]_  = \new_[83548]_  & \new_[83545]_ ;
  assign \new_[83552]_  = ~A202 & ~A200;
  assign \new_[83555]_  = ~A232 & ~A203;
  assign \new_[83556]_  = \new_[83555]_  & \new_[83552]_ ;
  assign \new_[83557]_  = \new_[83556]_  & \new_[83549]_ ;
  assign \new_[83560]_  = ~A266 & ~A233;
  assign \new_[83563]_  = ~A269 & ~A268;
  assign \new_[83564]_  = \new_[83563]_  & \new_[83560]_ ;
  assign \new_[83567]_  = ~A299 & A298;
  assign \new_[83570]_  = A302 & A300;
  assign \new_[83571]_  = \new_[83570]_  & \new_[83567]_ ;
  assign \new_[83572]_  = \new_[83571]_  & \new_[83564]_ ;
  assign \new_[83575]_  = ~A169 & A170;
  assign \new_[83578]_  = ~A166 & A167;
  assign \new_[83579]_  = \new_[83578]_  & \new_[83575]_ ;
  assign \new_[83582]_  = ~A201 & ~A200;
  assign \new_[83585]_  = ~A235 & ~A233;
  assign \new_[83586]_  = \new_[83585]_  & \new_[83582]_ ;
  assign \new_[83587]_  = \new_[83586]_  & \new_[83579]_ ;
  assign \new_[83590]_  = ~A266 & ~A236;
  assign \new_[83593]_  = ~A269 & ~A268;
  assign \new_[83594]_  = \new_[83593]_  & \new_[83590]_ ;
  assign \new_[83597]_  = ~A299 & A298;
  assign \new_[83600]_  = A301 & A300;
  assign \new_[83601]_  = \new_[83600]_  & \new_[83597]_ ;
  assign \new_[83602]_  = \new_[83601]_  & \new_[83594]_ ;
  assign \new_[83605]_  = ~A169 & A170;
  assign \new_[83608]_  = ~A166 & A167;
  assign \new_[83609]_  = \new_[83608]_  & \new_[83605]_ ;
  assign \new_[83612]_  = ~A201 & ~A200;
  assign \new_[83615]_  = ~A235 & ~A233;
  assign \new_[83616]_  = \new_[83615]_  & \new_[83612]_ ;
  assign \new_[83617]_  = \new_[83616]_  & \new_[83609]_ ;
  assign \new_[83620]_  = ~A266 & ~A236;
  assign \new_[83623]_  = ~A269 & ~A268;
  assign \new_[83624]_  = \new_[83623]_  & \new_[83620]_ ;
  assign \new_[83627]_  = ~A299 & A298;
  assign \new_[83630]_  = A302 & A300;
  assign \new_[83631]_  = \new_[83630]_  & \new_[83627]_ ;
  assign \new_[83632]_  = \new_[83631]_  & \new_[83624]_ ;
  assign \new_[83635]_  = ~A169 & A170;
  assign \new_[83638]_  = ~A166 & A167;
  assign \new_[83639]_  = \new_[83638]_  & \new_[83635]_ ;
  assign \new_[83642]_  = ~A200 & ~A199;
  assign \new_[83645]_  = ~A235 & ~A233;
  assign \new_[83646]_  = \new_[83645]_  & \new_[83642]_ ;
  assign \new_[83647]_  = \new_[83646]_  & \new_[83639]_ ;
  assign \new_[83650]_  = ~A266 & ~A236;
  assign \new_[83653]_  = ~A269 & ~A268;
  assign \new_[83654]_  = \new_[83653]_  & \new_[83650]_ ;
  assign \new_[83657]_  = ~A299 & A298;
  assign \new_[83660]_  = A301 & A300;
  assign \new_[83661]_  = \new_[83660]_  & \new_[83657]_ ;
  assign \new_[83662]_  = \new_[83661]_  & \new_[83654]_ ;
  assign \new_[83665]_  = ~A169 & A170;
  assign \new_[83668]_  = ~A166 & A167;
  assign \new_[83669]_  = \new_[83668]_  & \new_[83665]_ ;
  assign \new_[83672]_  = ~A200 & ~A199;
  assign \new_[83675]_  = ~A235 & ~A233;
  assign \new_[83676]_  = \new_[83675]_  & \new_[83672]_ ;
  assign \new_[83677]_  = \new_[83676]_  & \new_[83669]_ ;
  assign \new_[83680]_  = ~A266 & ~A236;
  assign \new_[83683]_  = ~A269 & ~A268;
  assign \new_[83684]_  = \new_[83683]_  & \new_[83680]_ ;
  assign \new_[83687]_  = ~A299 & A298;
  assign \new_[83690]_  = A302 & A300;
  assign \new_[83691]_  = \new_[83690]_  & \new_[83687]_ ;
  assign \new_[83692]_  = \new_[83691]_  & \new_[83684]_ ;
  assign \new_[83695]_  = ~A169 & A170;
  assign \new_[83698]_  = A166 & ~A167;
  assign \new_[83699]_  = \new_[83698]_  & \new_[83695]_ ;
  assign \new_[83702]_  = A200 & A199;
  assign \new_[83705]_  = ~A235 & ~A233;
  assign \new_[83706]_  = \new_[83705]_  & \new_[83702]_ ;
  assign \new_[83707]_  = \new_[83706]_  & \new_[83699]_ ;
  assign \new_[83710]_  = ~A266 & ~A236;
  assign \new_[83713]_  = ~A269 & ~A268;
  assign \new_[83714]_  = \new_[83713]_  & \new_[83710]_ ;
  assign \new_[83717]_  = ~A299 & A298;
  assign \new_[83720]_  = A301 & A300;
  assign \new_[83721]_  = \new_[83720]_  & \new_[83717]_ ;
  assign \new_[83722]_  = \new_[83721]_  & \new_[83714]_ ;
  assign \new_[83725]_  = ~A169 & A170;
  assign \new_[83728]_  = A166 & ~A167;
  assign \new_[83729]_  = \new_[83728]_  & \new_[83725]_ ;
  assign \new_[83732]_  = A200 & A199;
  assign \new_[83735]_  = ~A235 & ~A233;
  assign \new_[83736]_  = \new_[83735]_  & \new_[83732]_ ;
  assign \new_[83737]_  = \new_[83736]_  & \new_[83729]_ ;
  assign \new_[83740]_  = ~A266 & ~A236;
  assign \new_[83743]_  = ~A269 & ~A268;
  assign \new_[83744]_  = \new_[83743]_  & \new_[83740]_ ;
  assign \new_[83747]_  = ~A299 & A298;
  assign \new_[83750]_  = A302 & A300;
  assign \new_[83751]_  = \new_[83750]_  & \new_[83747]_ ;
  assign \new_[83752]_  = \new_[83751]_  & \new_[83744]_ ;
  assign \new_[83755]_  = ~A169 & A170;
  assign \new_[83758]_  = A166 & ~A167;
  assign \new_[83759]_  = \new_[83758]_  & \new_[83755]_ ;
  assign \new_[83762]_  = ~A202 & ~A200;
  assign \new_[83765]_  = A232 & ~A203;
  assign \new_[83766]_  = \new_[83765]_  & \new_[83762]_ ;
  assign \new_[83767]_  = \new_[83766]_  & \new_[83759]_ ;
  assign \new_[83770]_  = A265 & A233;
  assign \new_[83773]_  = ~A269 & ~A268;
  assign \new_[83774]_  = \new_[83773]_  & \new_[83770]_ ;
  assign \new_[83777]_  = ~A299 & A298;
  assign \new_[83780]_  = A301 & A300;
  assign \new_[83781]_  = \new_[83780]_  & \new_[83777]_ ;
  assign \new_[83782]_  = \new_[83781]_  & \new_[83774]_ ;
  assign \new_[83785]_  = ~A169 & A170;
  assign \new_[83788]_  = A166 & ~A167;
  assign \new_[83789]_  = \new_[83788]_  & \new_[83785]_ ;
  assign \new_[83792]_  = ~A202 & ~A200;
  assign \new_[83795]_  = A232 & ~A203;
  assign \new_[83796]_  = \new_[83795]_  & \new_[83792]_ ;
  assign \new_[83797]_  = \new_[83796]_  & \new_[83789]_ ;
  assign \new_[83800]_  = A265 & A233;
  assign \new_[83803]_  = ~A269 & ~A268;
  assign \new_[83804]_  = \new_[83803]_  & \new_[83800]_ ;
  assign \new_[83807]_  = ~A299 & A298;
  assign \new_[83810]_  = A302 & A300;
  assign \new_[83811]_  = \new_[83810]_  & \new_[83807]_ ;
  assign \new_[83812]_  = \new_[83811]_  & \new_[83804]_ ;
  assign \new_[83815]_  = ~A169 & A170;
  assign \new_[83818]_  = A166 & ~A167;
  assign \new_[83819]_  = \new_[83818]_  & \new_[83815]_ ;
  assign \new_[83822]_  = ~A202 & ~A200;
  assign \new_[83825]_  = ~A233 & ~A203;
  assign \new_[83826]_  = \new_[83825]_  & \new_[83822]_ ;
  assign \new_[83827]_  = \new_[83826]_  & \new_[83819]_ ;
  assign \new_[83830]_  = ~A236 & ~A235;
  assign \new_[83833]_  = A266 & A265;
  assign \new_[83834]_  = \new_[83833]_  & \new_[83830]_ ;
  assign \new_[83837]_  = ~A299 & A298;
  assign \new_[83840]_  = A301 & A300;
  assign \new_[83841]_  = \new_[83840]_  & \new_[83837]_ ;
  assign \new_[83842]_  = \new_[83841]_  & \new_[83834]_ ;
  assign \new_[83845]_  = ~A169 & A170;
  assign \new_[83848]_  = A166 & ~A167;
  assign \new_[83849]_  = \new_[83848]_  & \new_[83845]_ ;
  assign \new_[83852]_  = ~A202 & ~A200;
  assign \new_[83855]_  = ~A233 & ~A203;
  assign \new_[83856]_  = \new_[83855]_  & \new_[83852]_ ;
  assign \new_[83857]_  = \new_[83856]_  & \new_[83849]_ ;
  assign \new_[83860]_  = ~A236 & ~A235;
  assign \new_[83863]_  = A266 & A265;
  assign \new_[83864]_  = \new_[83863]_  & \new_[83860]_ ;
  assign \new_[83867]_  = ~A299 & A298;
  assign \new_[83870]_  = A302 & A300;
  assign \new_[83871]_  = \new_[83870]_  & \new_[83867]_ ;
  assign \new_[83872]_  = \new_[83871]_  & \new_[83864]_ ;
  assign \new_[83875]_  = ~A169 & A170;
  assign \new_[83878]_  = A166 & ~A167;
  assign \new_[83879]_  = \new_[83878]_  & \new_[83875]_ ;
  assign \new_[83882]_  = ~A202 & ~A200;
  assign \new_[83885]_  = ~A233 & ~A203;
  assign \new_[83886]_  = \new_[83885]_  & \new_[83882]_ ;
  assign \new_[83887]_  = \new_[83886]_  & \new_[83879]_ ;
  assign \new_[83890]_  = ~A236 & ~A235;
  assign \new_[83893]_  = ~A267 & ~A266;
  assign \new_[83894]_  = \new_[83893]_  & \new_[83890]_ ;
  assign \new_[83897]_  = ~A299 & A298;
  assign \new_[83900]_  = A301 & A300;
  assign \new_[83901]_  = \new_[83900]_  & \new_[83897]_ ;
  assign \new_[83902]_  = \new_[83901]_  & \new_[83894]_ ;
  assign \new_[83905]_  = ~A169 & A170;
  assign \new_[83908]_  = A166 & ~A167;
  assign \new_[83909]_  = \new_[83908]_  & \new_[83905]_ ;
  assign \new_[83912]_  = ~A202 & ~A200;
  assign \new_[83915]_  = ~A233 & ~A203;
  assign \new_[83916]_  = \new_[83915]_  & \new_[83912]_ ;
  assign \new_[83917]_  = \new_[83916]_  & \new_[83909]_ ;
  assign \new_[83920]_  = ~A236 & ~A235;
  assign \new_[83923]_  = ~A267 & ~A266;
  assign \new_[83924]_  = \new_[83923]_  & \new_[83920]_ ;
  assign \new_[83927]_  = ~A299 & A298;
  assign \new_[83930]_  = A302 & A300;
  assign \new_[83931]_  = \new_[83930]_  & \new_[83927]_ ;
  assign \new_[83932]_  = \new_[83931]_  & \new_[83924]_ ;
  assign \new_[83935]_  = ~A169 & A170;
  assign \new_[83938]_  = A166 & ~A167;
  assign \new_[83939]_  = \new_[83938]_  & \new_[83935]_ ;
  assign \new_[83942]_  = ~A202 & ~A200;
  assign \new_[83945]_  = ~A233 & ~A203;
  assign \new_[83946]_  = \new_[83945]_  & \new_[83942]_ ;
  assign \new_[83947]_  = \new_[83946]_  & \new_[83939]_ ;
  assign \new_[83950]_  = ~A236 & ~A235;
  assign \new_[83953]_  = ~A266 & ~A265;
  assign \new_[83954]_  = \new_[83953]_  & \new_[83950]_ ;
  assign \new_[83957]_  = ~A299 & A298;
  assign \new_[83960]_  = A301 & A300;
  assign \new_[83961]_  = \new_[83960]_  & \new_[83957]_ ;
  assign \new_[83962]_  = \new_[83961]_  & \new_[83954]_ ;
  assign \new_[83965]_  = ~A169 & A170;
  assign \new_[83968]_  = A166 & ~A167;
  assign \new_[83969]_  = \new_[83968]_  & \new_[83965]_ ;
  assign \new_[83972]_  = ~A202 & ~A200;
  assign \new_[83975]_  = ~A233 & ~A203;
  assign \new_[83976]_  = \new_[83975]_  & \new_[83972]_ ;
  assign \new_[83977]_  = \new_[83976]_  & \new_[83969]_ ;
  assign \new_[83980]_  = ~A236 & ~A235;
  assign \new_[83983]_  = ~A266 & ~A265;
  assign \new_[83984]_  = \new_[83983]_  & \new_[83980]_ ;
  assign \new_[83987]_  = ~A299 & A298;
  assign \new_[83990]_  = A302 & A300;
  assign \new_[83991]_  = \new_[83990]_  & \new_[83987]_ ;
  assign \new_[83992]_  = \new_[83991]_  & \new_[83984]_ ;
  assign \new_[83995]_  = ~A169 & A170;
  assign \new_[83998]_  = A166 & ~A167;
  assign \new_[83999]_  = \new_[83998]_  & \new_[83995]_ ;
  assign \new_[84002]_  = ~A202 & ~A200;
  assign \new_[84005]_  = ~A233 & ~A203;
  assign \new_[84006]_  = \new_[84005]_  & \new_[84002]_ ;
  assign \new_[84007]_  = \new_[84006]_  & \new_[83999]_ ;
  assign \new_[84010]_  = ~A266 & ~A234;
  assign \new_[84013]_  = ~A269 & ~A268;
  assign \new_[84014]_  = \new_[84013]_  & \new_[84010]_ ;
  assign \new_[84017]_  = ~A299 & A298;
  assign \new_[84020]_  = A301 & A300;
  assign \new_[84021]_  = \new_[84020]_  & \new_[84017]_ ;
  assign \new_[84022]_  = \new_[84021]_  & \new_[84014]_ ;
  assign \new_[84025]_  = ~A169 & A170;
  assign \new_[84028]_  = A166 & ~A167;
  assign \new_[84029]_  = \new_[84028]_  & \new_[84025]_ ;
  assign \new_[84032]_  = ~A202 & ~A200;
  assign \new_[84035]_  = ~A233 & ~A203;
  assign \new_[84036]_  = \new_[84035]_  & \new_[84032]_ ;
  assign \new_[84037]_  = \new_[84036]_  & \new_[84029]_ ;
  assign \new_[84040]_  = ~A266 & ~A234;
  assign \new_[84043]_  = ~A269 & ~A268;
  assign \new_[84044]_  = \new_[84043]_  & \new_[84040]_ ;
  assign \new_[84047]_  = ~A299 & A298;
  assign \new_[84050]_  = A302 & A300;
  assign \new_[84051]_  = \new_[84050]_  & \new_[84047]_ ;
  assign \new_[84052]_  = \new_[84051]_  & \new_[84044]_ ;
  assign \new_[84055]_  = ~A169 & A170;
  assign \new_[84058]_  = A166 & ~A167;
  assign \new_[84059]_  = \new_[84058]_  & \new_[84055]_ ;
  assign \new_[84062]_  = ~A202 & ~A200;
  assign \new_[84065]_  = ~A232 & ~A203;
  assign \new_[84066]_  = \new_[84065]_  & \new_[84062]_ ;
  assign \new_[84067]_  = \new_[84066]_  & \new_[84059]_ ;
  assign \new_[84070]_  = ~A266 & ~A233;
  assign \new_[84073]_  = ~A269 & ~A268;
  assign \new_[84074]_  = \new_[84073]_  & \new_[84070]_ ;
  assign \new_[84077]_  = ~A299 & A298;
  assign \new_[84080]_  = A301 & A300;
  assign \new_[84081]_  = \new_[84080]_  & \new_[84077]_ ;
  assign \new_[84082]_  = \new_[84081]_  & \new_[84074]_ ;
  assign \new_[84085]_  = ~A169 & A170;
  assign \new_[84088]_  = A166 & ~A167;
  assign \new_[84089]_  = \new_[84088]_  & \new_[84085]_ ;
  assign \new_[84092]_  = ~A202 & ~A200;
  assign \new_[84095]_  = ~A232 & ~A203;
  assign \new_[84096]_  = \new_[84095]_  & \new_[84092]_ ;
  assign \new_[84097]_  = \new_[84096]_  & \new_[84089]_ ;
  assign \new_[84100]_  = ~A266 & ~A233;
  assign \new_[84103]_  = ~A269 & ~A268;
  assign \new_[84104]_  = \new_[84103]_  & \new_[84100]_ ;
  assign \new_[84107]_  = ~A299 & A298;
  assign \new_[84110]_  = A302 & A300;
  assign \new_[84111]_  = \new_[84110]_  & \new_[84107]_ ;
  assign \new_[84112]_  = \new_[84111]_  & \new_[84104]_ ;
  assign \new_[84115]_  = ~A169 & A170;
  assign \new_[84118]_  = A166 & ~A167;
  assign \new_[84119]_  = \new_[84118]_  & \new_[84115]_ ;
  assign \new_[84122]_  = ~A201 & ~A200;
  assign \new_[84125]_  = ~A235 & ~A233;
  assign \new_[84126]_  = \new_[84125]_  & \new_[84122]_ ;
  assign \new_[84127]_  = \new_[84126]_  & \new_[84119]_ ;
  assign \new_[84130]_  = ~A266 & ~A236;
  assign \new_[84133]_  = ~A269 & ~A268;
  assign \new_[84134]_  = \new_[84133]_  & \new_[84130]_ ;
  assign \new_[84137]_  = ~A299 & A298;
  assign \new_[84140]_  = A301 & A300;
  assign \new_[84141]_  = \new_[84140]_  & \new_[84137]_ ;
  assign \new_[84142]_  = \new_[84141]_  & \new_[84134]_ ;
  assign \new_[84145]_  = ~A169 & A170;
  assign \new_[84148]_  = A166 & ~A167;
  assign \new_[84149]_  = \new_[84148]_  & \new_[84145]_ ;
  assign \new_[84152]_  = ~A201 & ~A200;
  assign \new_[84155]_  = ~A235 & ~A233;
  assign \new_[84156]_  = \new_[84155]_  & \new_[84152]_ ;
  assign \new_[84157]_  = \new_[84156]_  & \new_[84149]_ ;
  assign \new_[84160]_  = ~A266 & ~A236;
  assign \new_[84163]_  = ~A269 & ~A268;
  assign \new_[84164]_  = \new_[84163]_  & \new_[84160]_ ;
  assign \new_[84167]_  = ~A299 & A298;
  assign \new_[84170]_  = A302 & A300;
  assign \new_[84171]_  = \new_[84170]_  & \new_[84167]_ ;
  assign \new_[84172]_  = \new_[84171]_  & \new_[84164]_ ;
  assign \new_[84175]_  = ~A169 & A170;
  assign \new_[84178]_  = A166 & ~A167;
  assign \new_[84179]_  = \new_[84178]_  & \new_[84175]_ ;
  assign \new_[84182]_  = ~A200 & ~A199;
  assign \new_[84185]_  = ~A235 & ~A233;
  assign \new_[84186]_  = \new_[84185]_  & \new_[84182]_ ;
  assign \new_[84187]_  = \new_[84186]_  & \new_[84179]_ ;
  assign \new_[84190]_  = ~A266 & ~A236;
  assign \new_[84193]_  = ~A269 & ~A268;
  assign \new_[84194]_  = \new_[84193]_  & \new_[84190]_ ;
  assign \new_[84197]_  = ~A299 & A298;
  assign \new_[84200]_  = A301 & A300;
  assign \new_[84201]_  = \new_[84200]_  & \new_[84197]_ ;
  assign \new_[84202]_  = \new_[84201]_  & \new_[84194]_ ;
  assign \new_[84205]_  = ~A169 & A170;
  assign \new_[84208]_  = A166 & ~A167;
  assign \new_[84209]_  = \new_[84208]_  & \new_[84205]_ ;
  assign \new_[84212]_  = ~A200 & ~A199;
  assign \new_[84215]_  = ~A235 & ~A233;
  assign \new_[84216]_  = \new_[84215]_  & \new_[84212]_ ;
  assign \new_[84217]_  = \new_[84216]_  & \new_[84209]_ ;
  assign \new_[84220]_  = ~A266 & ~A236;
  assign \new_[84223]_  = ~A269 & ~A268;
  assign \new_[84224]_  = \new_[84223]_  & \new_[84220]_ ;
  assign \new_[84227]_  = ~A299 & A298;
  assign \new_[84230]_  = A302 & A300;
  assign \new_[84231]_  = \new_[84230]_  & \new_[84227]_ ;
  assign \new_[84232]_  = \new_[84231]_  & \new_[84224]_ ;
  assign \new_[84235]_  = ~A169 & ~A170;
  assign \new_[84238]_  = A199 & ~A168;
  assign \new_[84239]_  = \new_[84238]_  & \new_[84235]_ ;
  assign \new_[84242]_  = A201 & ~A200;
  assign \new_[84245]_  = A232 & A202;
  assign \new_[84246]_  = \new_[84245]_  & \new_[84242]_ ;
  assign \new_[84247]_  = \new_[84246]_  & \new_[84239]_ ;
  assign \new_[84250]_  = A265 & A233;
  assign \new_[84253]_  = ~A269 & ~A268;
  assign \new_[84254]_  = \new_[84253]_  & \new_[84250]_ ;
  assign \new_[84257]_  = ~A299 & A298;
  assign \new_[84260]_  = A301 & A300;
  assign \new_[84261]_  = \new_[84260]_  & \new_[84257]_ ;
  assign \new_[84262]_  = \new_[84261]_  & \new_[84254]_ ;
  assign \new_[84265]_  = ~A169 & ~A170;
  assign \new_[84268]_  = A199 & ~A168;
  assign \new_[84269]_  = \new_[84268]_  & \new_[84265]_ ;
  assign \new_[84272]_  = A201 & ~A200;
  assign \new_[84275]_  = A232 & A202;
  assign \new_[84276]_  = \new_[84275]_  & \new_[84272]_ ;
  assign \new_[84277]_  = \new_[84276]_  & \new_[84269]_ ;
  assign \new_[84280]_  = A265 & A233;
  assign \new_[84283]_  = ~A269 & ~A268;
  assign \new_[84284]_  = \new_[84283]_  & \new_[84280]_ ;
  assign \new_[84287]_  = ~A299 & A298;
  assign \new_[84290]_  = A302 & A300;
  assign \new_[84291]_  = \new_[84290]_  & \new_[84287]_ ;
  assign \new_[84292]_  = \new_[84291]_  & \new_[84284]_ ;
  assign \new_[84295]_  = ~A169 & ~A170;
  assign \new_[84298]_  = A199 & ~A168;
  assign \new_[84299]_  = \new_[84298]_  & \new_[84295]_ ;
  assign \new_[84302]_  = A201 & ~A200;
  assign \new_[84305]_  = ~A233 & A202;
  assign \new_[84306]_  = \new_[84305]_  & \new_[84302]_ ;
  assign \new_[84307]_  = \new_[84306]_  & \new_[84299]_ ;
  assign \new_[84310]_  = ~A236 & ~A235;
  assign \new_[84313]_  = A266 & A265;
  assign \new_[84314]_  = \new_[84313]_  & \new_[84310]_ ;
  assign \new_[84317]_  = ~A299 & A298;
  assign \new_[84320]_  = A301 & A300;
  assign \new_[84321]_  = \new_[84320]_  & \new_[84317]_ ;
  assign \new_[84322]_  = \new_[84321]_  & \new_[84314]_ ;
  assign \new_[84325]_  = ~A169 & ~A170;
  assign \new_[84328]_  = A199 & ~A168;
  assign \new_[84329]_  = \new_[84328]_  & \new_[84325]_ ;
  assign \new_[84332]_  = A201 & ~A200;
  assign \new_[84335]_  = ~A233 & A202;
  assign \new_[84336]_  = \new_[84335]_  & \new_[84332]_ ;
  assign \new_[84337]_  = \new_[84336]_  & \new_[84329]_ ;
  assign \new_[84340]_  = ~A236 & ~A235;
  assign \new_[84343]_  = A266 & A265;
  assign \new_[84344]_  = \new_[84343]_  & \new_[84340]_ ;
  assign \new_[84347]_  = ~A299 & A298;
  assign \new_[84350]_  = A302 & A300;
  assign \new_[84351]_  = \new_[84350]_  & \new_[84347]_ ;
  assign \new_[84352]_  = \new_[84351]_  & \new_[84344]_ ;
  assign \new_[84355]_  = ~A169 & ~A170;
  assign \new_[84358]_  = A199 & ~A168;
  assign \new_[84359]_  = \new_[84358]_  & \new_[84355]_ ;
  assign \new_[84362]_  = A201 & ~A200;
  assign \new_[84365]_  = ~A233 & A202;
  assign \new_[84366]_  = \new_[84365]_  & \new_[84362]_ ;
  assign \new_[84367]_  = \new_[84366]_  & \new_[84359]_ ;
  assign \new_[84370]_  = ~A236 & ~A235;
  assign \new_[84373]_  = ~A267 & ~A266;
  assign \new_[84374]_  = \new_[84373]_  & \new_[84370]_ ;
  assign \new_[84377]_  = ~A299 & A298;
  assign \new_[84380]_  = A301 & A300;
  assign \new_[84381]_  = \new_[84380]_  & \new_[84377]_ ;
  assign \new_[84382]_  = \new_[84381]_  & \new_[84374]_ ;
  assign \new_[84385]_  = ~A169 & ~A170;
  assign \new_[84388]_  = A199 & ~A168;
  assign \new_[84389]_  = \new_[84388]_  & \new_[84385]_ ;
  assign \new_[84392]_  = A201 & ~A200;
  assign \new_[84395]_  = ~A233 & A202;
  assign \new_[84396]_  = \new_[84395]_  & \new_[84392]_ ;
  assign \new_[84397]_  = \new_[84396]_  & \new_[84389]_ ;
  assign \new_[84400]_  = ~A236 & ~A235;
  assign \new_[84403]_  = ~A267 & ~A266;
  assign \new_[84404]_  = \new_[84403]_  & \new_[84400]_ ;
  assign \new_[84407]_  = ~A299 & A298;
  assign \new_[84410]_  = A302 & A300;
  assign \new_[84411]_  = \new_[84410]_  & \new_[84407]_ ;
  assign \new_[84412]_  = \new_[84411]_  & \new_[84404]_ ;
  assign \new_[84415]_  = ~A169 & ~A170;
  assign \new_[84418]_  = A199 & ~A168;
  assign \new_[84419]_  = \new_[84418]_  & \new_[84415]_ ;
  assign \new_[84422]_  = A201 & ~A200;
  assign \new_[84425]_  = ~A233 & A202;
  assign \new_[84426]_  = \new_[84425]_  & \new_[84422]_ ;
  assign \new_[84427]_  = \new_[84426]_  & \new_[84419]_ ;
  assign \new_[84430]_  = ~A236 & ~A235;
  assign \new_[84433]_  = ~A266 & ~A265;
  assign \new_[84434]_  = \new_[84433]_  & \new_[84430]_ ;
  assign \new_[84437]_  = ~A299 & A298;
  assign \new_[84440]_  = A301 & A300;
  assign \new_[84441]_  = \new_[84440]_  & \new_[84437]_ ;
  assign \new_[84442]_  = \new_[84441]_  & \new_[84434]_ ;
  assign \new_[84445]_  = ~A169 & ~A170;
  assign \new_[84448]_  = A199 & ~A168;
  assign \new_[84449]_  = \new_[84448]_  & \new_[84445]_ ;
  assign \new_[84452]_  = A201 & ~A200;
  assign \new_[84455]_  = ~A233 & A202;
  assign \new_[84456]_  = \new_[84455]_  & \new_[84452]_ ;
  assign \new_[84457]_  = \new_[84456]_  & \new_[84449]_ ;
  assign \new_[84460]_  = ~A236 & ~A235;
  assign \new_[84463]_  = ~A266 & ~A265;
  assign \new_[84464]_  = \new_[84463]_  & \new_[84460]_ ;
  assign \new_[84467]_  = ~A299 & A298;
  assign \new_[84470]_  = A302 & A300;
  assign \new_[84471]_  = \new_[84470]_  & \new_[84467]_ ;
  assign \new_[84472]_  = \new_[84471]_  & \new_[84464]_ ;
  assign \new_[84475]_  = ~A169 & ~A170;
  assign \new_[84478]_  = A199 & ~A168;
  assign \new_[84479]_  = \new_[84478]_  & \new_[84475]_ ;
  assign \new_[84482]_  = A201 & ~A200;
  assign \new_[84485]_  = ~A233 & A202;
  assign \new_[84486]_  = \new_[84485]_  & \new_[84482]_ ;
  assign \new_[84487]_  = \new_[84486]_  & \new_[84479]_ ;
  assign \new_[84490]_  = ~A266 & ~A234;
  assign \new_[84493]_  = ~A269 & ~A268;
  assign \new_[84494]_  = \new_[84493]_  & \new_[84490]_ ;
  assign \new_[84497]_  = ~A299 & A298;
  assign \new_[84500]_  = A301 & A300;
  assign \new_[84501]_  = \new_[84500]_  & \new_[84497]_ ;
  assign \new_[84502]_  = \new_[84501]_  & \new_[84494]_ ;
  assign \new_[84505]_  = ~A169 & ~A170;
  assign \new_[84508]_  = A199 & ~A168;
  assign \new_[84509]_  = \new_[84508]_  & \new_[84505]_ ;
  assign \new_[84512]_  = A201 & ~A200;
  assign \new_[84515]_  = ~A233 & A202;
  assign \new_[84516]_  = \new_[84515]_  & \new_[84512]_ ;
  assign \new_[84517]_  = \new_[84516]_  & \new_[84509]_ ;
  assign \new_[84520]_  = ~A266 & ~A234;
  assign \new_[84523]_  = ~A269 & ~A268;
  assign \new_[84524]_  = \new_[84523]_  & \new_[84520]_ ;
  assign \new_[84527]_  = ~A299 & A298;
  assign \new_[84530]_  = A302 & A300;
  assign \new_[84531]_  = \new_[84530]_  & \new_[84527]_ ;
  assign \new_[84532]_  = \new_[84531]_  & \new_[84524]_ ;
  assign \new_[84535]_  = ~A169 & ~A170;
  assign \new_[84538]_  = A199 & ~A168;
  assign \new_[84539]_  = \new_[84538]_  & \new_[84535]_ ;
  assign \new_[84542]_  = A201 & ~A200;
  assign \new_[84545]_  = ~A232 & A202;
  assign \new_[84546]_  = \new_[84545]_  & \new_[84542]_ ;
  assign \new_[84547]_  = \new_[84546]_  & \new_[84539]_ ;
  assign \new_[84550]_  = ~A266 & ~A233;
  assign \new_[84553]_  = ~A269 & ~A268;
  assign \new_[84554]_  = \new_[84553]_  & \new_[84550]_ ;
  assign \new_[84557]_  = ~A299 & A298;
  assign \new_[84560]_  = A301 & A300;
  assign \new_[84561]_  = \new_[84560]_  & \new_[84557]_ ;
  assign \new_[84562]_  = \new_[84561]_  & \new_[84554]_ ;
  assign \new_[84565]_  = ~A169 & ~A170;
  assign \new_[84568]_  = A199 & ~A168;
  assign \new_[84569]_  = \new_[84568]_  & \new_[84565]_ ;
  assign \new_[84572]_  = A201 & ~A200;
  assign \new_[84575]_  = ~A232 & A202;
  assign \new_[84576]_  = \new_[84575]_  & \new_[84572]_ ;
  assign \new_[84577]_  = \new_[84576]_  & \new_[84569]_ ;
  assign \new_[84580]_  = ~A266 & ~A233;
  assign \new_[84583]_  = ~A269 & ~A268;
  assign \new_[84584]_  = \new_[84583]_  & \new_[84580]_ ;
  assign \new_[84587]_  = ~A299 & A298;
  assign \new_[84590]_  = A302 & A300;
  assign \new_[84591]_  = \new_[84590]_  & \new_[84587]_ ;
  assign \new_[84592]_  = \new_[84591]_  & \new_[84584]_ ;
  assign \new_[84595]_  = ~A169 & ~A170;
  assign \new_[84598]_  = A199 & ~A168;
  assign \new_[84599]_  = \new_[84598]_  & \new_[84595]_ ;
  assign \new_[84602]_  = A201 & ~A200;
  assign \new_[84605]_  = A232 & A203;
  assign \new_[84606]_  = \new_[84605]_  & \new_[84602]_ ;
  assign \new_[84607]_  = \new_[84606]_  & \new_[84599]_ ;
  assign \new_[84610]_  = A265 & A233;
  assign \new_[84613]_  = ~A269 & ~A268;
  assign \new_[84614]_  = \new_[84613]_  & \new_[84610]_ ;
  assign \new_[84617]_  = ~A299 & A298;
  assign \new_[84620]_  = A301 & A300;
  assign \new_[84621]_  = \new_[84620]_  & \new_[84617]_ ;
  assign \new_[84622]_  = \new_[84621]_  & \new_[84614]_ ;
  assign \new_[84625]_  = ~A169 & ~A170;
  assign \new_[84628]_  = A199 & ~A168;
  assign \new_[84629]_  = \new_[84628]_  & \new_[84625]_ ;
  assign \new_[84632]_  = A201 & ~A200;
  assign \new_[84635]_  = A232 & A203;
  assign \new_[84636]_  = \new_[84635]_  & \new_[84632]_ ;
  assign \new_[84637]_  = \new_[84636]_  & \new_[84629]_ ;
  assign \new_[84640]_  = A265 & A233;
  assign \new_[84643]_  = ~A269 & ~A268;
  assign \new_[84644]_  = \new_[84643]_  & \new_[84640]_ ;
  assign \new_[84647]_  = ~A299 & A298;
  assign \new_[84650]_  = A302 & A300;
  assign \new_[84651]_  = \new_[84650]_  & \new_[84647]_ ;
  assign \new_[84652]_  = \new_[84651]_  & \new_[84644]_ ;
  assign \new_[84655]_  = ~A169 & ~A170;
  assign \new_[84658]_  = A199 & ~A168;
  assign \new_[84659]_  = \new_[84658]_  & \new_[84655]_ ;
  assign \new_[84662]_  = A201 & ~A200;
  assign \new_[84665]_  = ~A233 & A203;
  assign \new_[84666]_  = \new_[84665]_  & \new_[84662]_ ;
  assign \new_[84667]_  = \new_[84666]_  & \new_[84659]_ ;
  assign \new_[84670]_  = ~A236 & ~A235;
  assign \new_[84673]_  = A266 & A265;
  assign \new_[84674]_  = \new_[84673]_  & \new_[84670]_ ;
  assign \new_[84677]_  = ~A299 & A298;
  assign \new_[84680]_  = A301 & A300;
  assign \new_[84681]_  = \new_[84680]_  & \new_[84677]_ ;
  assign \new_[84682]_  = \new_[84681]_  & \new_[84674]_ ;
  assign \new_[84685]_  = ~A169 & ~A170;
  assign \new_[84688]_  = A199 & ~A168;
  assign \new_[84689]_  = \new_[84688]_  & \new_[84685]_ ;
  assign \new_[84692]_  = A201 & ~A200;
  assign \new_[84695]_  = ~A233 & A203;
  assign \new_[84696]_  = \new_[84695]_  & \new_[84692]_ ;
  assign \new_[84697]_  = \new_[84696]_  & \new_[84689]_ ;
  assign \new_[84700]_  = ~A236 & ~A235;
  assign \new_[84703]_  = A266 & A265;
  assign \new_[84704]_  = \new_[84703]_  & \new_[84700]_ ;
  assign \new_[84707]_  = ~A299 & A298;
  assign \new_[84710]_  = A302 & A300;
  assign \new_[84711]_  = \new_[84710]_  & \new_[84707]_ ;
  assign \new_[84712]_  = \new_[84711]_  & \new_[84704]_ ;
  assign \new_[84715]_  = ~A169 & ~A170;
  assign \new_[84718]_  = A199 & ~A168;
  assign \new_[84719]_  = \new_[84718]_  & \new_[84715]_ ;
  assign \new_[84722]_  = A201 & ~A200;
  assign \new_[84725]_  = ~A233 & A203;
  assign \new_[84726]_  = \new_[84725]_  & \new_[84722]_ ;
  assign \new_[84727]_  = \new_[84726]_  & \new_[84719]_ ;
  assign \new_[84730]_  = ~A236 & ~A235;
  assign \new_[84733]_  = ~A267 & ~A266;
  assign \new_[84734]_  = \new_[84733]_  & \new_[84730]_ ;
  assign \new_[84737]_  = ~A299 & A298;
  assign \new_[84740]_  = A301 & A300;
  assign \new_[84741]_  = \new_[84740]_  & \new_[84737]_ ;
  assign \new_[84742]_  = \new_[84741]_  & \new_[84734]_ ;
  assign \new_[84745]_  = ~A169 & ~A170;
  assign \new_[84748]_  = A199 & ~A168;
  assign \new_[84749]_  = \new_[84748]_  & \new_[84745]_ ;
  assign \new_[84752]_  = A201 & ~A200;
  assign \new_[84755]_  = ~A233 & A203;
  assign \new_[84756]_  = \new_[84755]_  & \new_[84752]_ ;
  assign \new_[84757]_  = \new_[84756]_  & \new_[84749]_ ;
  assign \new_[84760]_  = ~A236 & ~A235;
  assign \new_[84763]_  = ~A267 & ~A266;
  assign \new_[84764]_  = \new_[84763]_  & \new_[84760]_ ;
  assign \new_[84767]_  = ~A299 & A298;
  assign \new_[84770]_  = A302 & A300;
  assign \new_[84771]_  = \new_[84770]_  & \new_[84767]_ ;
  assign \new_[84772]_  = \new_[84771]_  & \new_[84764]_ ;
  assign \new_[84775]_  = ~A169 & ~A170;
  assign \new_[84778]_  = A199 & ~A168;
  assign \new_[84779]_  = \new_[84778]_  & \new_[84775]_ ;
  assign \new_[84782]_  = A201 & ~A200;
  assign \new_[84785]_  = ~A233 & A203;
  assign \new_[84786]_  = \new_[84785]_  & \new_[84782]_ ;
  assign \new_[84787]_  = \new_[84786]_  & \new_[84779]_ ;
  assign \new_[84790]_  = ~A236 & ~A235;
  assign \new_[84793]_  = ~A266 & ~A265;
  assign \new_[84794]_  = \new_[84793]_  & \new_[84790]_ ;
  assign \new_[84797]_  = ~A299 & A298;
  assign \new_[84800]_  = A301 & A300;
  assign \new_[84801]_  = \new_[84800]_  & \new_[84797]_ ;
  assign \new_[84802]_  = \new_[84801]_  & \new_[84794]_ ;
  assign \new_[84805]_  = ~A169 & ~A170;
  assign \new_[84808]_  = A199 & ~A168;
  assign \new_[84809]_  = \new_[84808]_  & \new_[84805]_ ;
  assign \new_[84812]_  = A201 & ~A200;
  assign \new_[84815]_  = ~A233 & A203;
  assign \new_[84816]_  = \new_[84815]_  & \new_[84812]_ ;
  assign \new_[84817]_  = \new_[84816]_  & \new_[84809]_ ;
  assign \new_[84820]_  = ~A236 & ~A235;
  assign \new_[84823]_  = ~A266 & ~A265;
  assign \new_[84824]_  = \new_[84823]_  & \new_[84820]_ ;
  assign \new_[84827]_  = ~A299 & A298;
  assign \new_[84830]_  = A302 & A300;
  assign \new_[84831]_  = \new_[84830]_  & \new_[84827]_ ;
  assign \new_[84832]_  = \new_[84831]_  & \new_[84824]_ ;
  assign \new_[84835]_  = ~A169 & ~A170;
  assign \new_[84838]_  = A199 & ~A168;
  assign \new_[84839]_  = \new_[84838]_  & \new_[84835]_ ;
  assign \new_[84842]_  = A201 & ~A200;
  assign \new_[84845]_  = ~A233 & A203;
  assign \new_[84846]_  = \new_[84845]_  & \new_[84842]_ ;
  assign \new_[84847]_  = \new_[84846]_  & \new_[84839]_ ;
  assign \new_[84850]_  = ~A266 & ~A234;
  assign \new_[84853]_  = ~A269 & ~A268;
  assign \new_[84854]_  = \new_[84853]_  & \new_[84850]_ ;
  assign \new_[84857]_  = ~A299 & A298;
  assign \new_[84860]_  = A301 & A300;
  assign \new_[84861]_  = \new_[84860]_  & \new_[84857]_ ;
  assign \new_[84862]_  = \new_[84861]_  & \new_[84854]_ ;
  assign \new_[84865]_  = ~A169 & ~A170;
  assign \new_[84868]_  = A199 & ~A168;
  assign \new_[84869]_  = \new_[84868]_  & \new_[84865]_ ;
  assign \new_[84872]_  = A201 & ~A200;
  assign \new_[84875]_  = ~A233 & A203;
  assign \new_[84876]_  = \new_[84875]_  & \new_[84872]_ ;
  assign \new_[84877]_  = \new_[84876]_  & \new_[84869]_ ;
  assign \new_[84880]_  = ~A266 & ~A234;
  assign \new_[84883]_  = ~A269 & ~A268;
  assign \new_[84884]_  = \new_[84883]_  & \new_[84880]_ ;
  assign \new_[84887]_  = ~A299 & A298;
  assign \new_[84890]_  = A302 & A300;
  assign \new_[84891]_  = \new_[84890]_  & \new_[84887]_ ;
  assign \new_[84892]_  = \new_[84891]_  & \new_[84884]_ ;
  assign \new_[84895]_  = ~A169 & ~A170;
  assign \new_[84898]_  = A199 & ~A168;
  assign \new_[84899]_  = \new_[84898]_  & \new_[84895]_ ;
  assign \new_[84902]_  = A201 & ~A200;
  assign \new_[84905]_  = ~A232 & A203;
  assign \new_[84906]_  = \new_[84905]_  & \new_[84902]_ ;
  assign \new_[84907]_  = \new_[84906]_  & \new_[84899]_ ;
  assign \new_[84910]_  = ~A266 & ~A233;
  assign \new_[84913]_  = ~A269 & ~A268;
  assign \new_[84914]_  = \new_[84913]_  & \new_[84910]_ ;
  assign \new_[84917]_  = ~A299 & A298;
  assign \new_[84920]_  = A301 & A300;
  assign \new_[84921]_  = \new_[84920]_  & \new_[84917]_ ;
  assign \new_[84922]_  = \new_[84921]_  & \new_[84914]_ ;
  assign \new_[84925]_  = ~A169 & ~A170;
  assign \new_[84928]_  = A199 & ~A168;
  assign \new_[84929]_  = \new_[84928]_  & \new_[84925]_ ;
  assign \new_[84932]_  = A201 & ~A200;
  assign \new_[84935]_  = ~A232 & A203;
  assign \new_[84936]_  = \new_[84935]_  & \new_[84932]_ ;
  assign \new_[84937]_  = \new_[84936]_  & \new_[84929]_ ;
  assign \new_[84940]_  = ~A266 & ~A233;
  assign \new_[84943]_  = ~A269 & ~A268;
  assign \new_[84944]_  = \new_[84943]_  & \new_[84940]_ ;
  assign \new_[84947]_  = ~A299 & A298;
  assign \new_[84950]_  = A302 & A300;
  assign \new_[84951]_  = \new_[84950]_  & \new_[84947]_ ;
  assign \new_[84952]_  = \new_[84951]_  & \new_[84944]_ ;
  assign \new_[84955]_  = ~A167 & A170;
  assign \new_[84958]_  = A199 & ~A166;
  assign \new_[84959]_  = \new_[84958]_  & \new_[84955]_ ;
  assign \new_[84962]_  = A201 & ~A200;
  assign \new_[84965]_  = ~A233 & A202;
  assign \new_[84966]_  = \new_[84965]_  & \new_[84962]_ ;
  assign \new_[84967]_  = \new_[84966]_  & \new_[84959]_ ;
  assign \new_[84970]_  = ~A236 & ~A235;
  assign \new_[84973]_  = ~A268 & ~A266;
  assign \new_[84974]_  = \new_[84973]_  & \new_[84970]_ ;
  assign \new_[84977]_  = A298 & ~A269;
  assign \new_[84981]_  = A301 & A300;
  assign \new_[84982]_  = ~A299 & \new_[84981]_ ;
  assign \new_[84983]_  = \new_[84982]_  & \new_[84977]_ ;
  assign \new_[84984]_  = \new_[84983]_  & \new_[84974]_ ;
  assign \new_[84987]_  = ~A167 & A170;
  assign \new_[84990]_  = A199 & ~A166;
  assign \new_[84991]_  = \new_[84990]_  & \new_[84987]_ ;
  assign \new_[84994]_  = A201 & ~A200;
  assign \new_[84997]_  = ~A233 & A202;
  assign \new_[84998]_  = \new_[84997]_  & \new_[84994]_ ;
  assign \new_[84999]_  = \new_[84998]_  & \new_[84991]_ ;
  assign \new_[85002]_  = ~A236 & ~A235;
  assign \new_[85005]_  = ~A268 & ~A266;
  assign \new_[85006]_  = \new_[85005]_  & \new_[85002]_ ;
  assign \new_[85009]_  = A298 & ~A269;
  assign \new_[85013]_  = A302 & A300;
  assign \new_[85014]_  = ~A299 & \new_[85013]_ ;
  assign \new_[85015]_  = \new_[85014]_  & \new_[85009]_ ;
  assign \new_[85016]_  = \new_[85015]_  & \new_[85006]_ ;
  assign \new_[85019]_  = ~A167 & A170;
  assign \new_[85022]_  = A199 & ~A166;
  assign \new_[85023]_  = \new_[85022]_  & \new_[85019]_ ;
  assign \new_[85026]_  = A201 & ~A200;
  assign \new_[85029]_  = ~A233 & A203;
  assign \new_[85030]_  = \new_[85029]_  & \new_[85026]_ ;
  assign \new_[85031]_  = \new_[85030]_  & \new_[85023]_ ;
  assign \new_[85034]_  = ~A236 & ~A235;
  assign \new_[85037]_  = ~A268 & ~A266;
  assign \new_[85038]_  = \new_[85037]_  & \new_[85034]_ ;
  assign \new_[85041]_  = A298 & ~A269;
  assign \new_[85045]_  = A301 & A300;
  assign \new_[85046]_  = ~A299 & \new_[85045]_ ;
  assign \new_[85047]_  = \new_[85046]_  & \new_[85041]_ ;
  assign \new_[85048]_  = \new_[85047]_  & \new_[85038]_ ;
  assign \new_[85051]_  = ~A167 & A170;
  assign \new_[85054]_  = A199 & ~A166;
  assign \new_[85055]_  = \new_[85054]_  & \new_[85051]_ ;
  assign \new_[85058]_  = A201 & ~A200;
  assign \new_[85061]_  = ~A233 & A203;
  assign \new_[85062]_  = \new_[85061]_  & \new_[85058]_ ;
  assign \new_[85063]_  = \new_[85062]_  & \new_[85055]_ ;
  assign \new_[85066]_  = ~A236 & ~A235;
  assign \new_[85069]_  = ~A268 & ~A266;
  assign \new_[85070]_  = \new_[85069]_  & \new_[85066]_ ;
  assign \new_[85073]_  = A298 & ~A269;
  assign \new_[85077]_  = A302 & A300;
  assign \new_[85078]_  = ~A299 & \new_[85077]_ ;
  assign \new_[85079]_  = \new_[85078]_  & \new_[85073]_ ;
  assign \new_[85080]_  = \new_[85079]_  & \new_[85070]_ ;
  assign \new_[85083]_  = ~A168 & A169;
  assign \new_[85086]_  = ~A166 & A167;
  assign \new_[85087]_  = \new_[85086]_  & \new_[85083]_ ;
  assign \new_[85090]_  = ~A200 & A199;
  assign \new_[85093]_  = A202 & A201;
  assign \new_[85094]_  = \new_[85093]_  & \new_[85090]_ ;
  assign \new_[85095]_  = \new_[85094]_  & \new_[85087]_ ;
  assign \new_[85098]_  = A233 & A232;
  assign \new_[85101]_  = ~A268 & A265;
  assign \new_[85102]_  = \new_[85101]_  & \new_[85098]_ ;
  assign \new_[85105]_  = A298 & ~A269;
  assign \new_[85109]_  = A301 & A300;
  assign \new_[85110]_  = ~A299 & \new_[85109]_ ;
  assign \new_[85111]_  = \new_[85110]_  & \new_[85105]_ ;
  assign \new_[85112]_  = \new_[85111]_  & \new_[85102]_ ;
  assign \new_[85115]_  = ~A168 & A169;
  assign \new_[85118]_  = ~A166 & A167;
  assign \new_[85119]_  = \new_[85118]_  & \new_[85115]_ ;
  assign \new_[85122]_  = ~A200 & A199;
  assign \new_[85125]_  = A202 & A201;
  assign \new_[85126]_  = \new_[85125]_  & \new_[85122]_ ;
  assign \new_[85127]_  = \new_[85126]_  & \new_[85119]_ ;
  assign \new_[85130]_  = A233 & A232;
  assign \new_[85133]_  = ~A268 & A265;
  assign \new_[85134]_  = \new_[85133]_  & \new_[85130]_ ;
  assign \new_[85137]_  = A298 & ~A269;
  assign \new_[85141]_  = A302 & A300;
  assign \new_[85142]_  = ~A299 & \new_[85141]_ ;
  assign \new_[85143]_  = \new_[85142]_  & \new_[85137]_ ;
  assign \new_[85144]_  = \new_[85143]_  & \new_[85134]_ ;
  assign \new_[85147]_  = ~A168 & A169;
  assign \new_[85150]_  = ~A166 & A167;
  assign \new_[85151]_  = \new_[85150]_  & \new_[85147]_ ;
  assign \new_[85154]_  = ~A200 & A199;
  assign \new_[85157]_  = A202 & A201;
  assign \new_[85158]_  = \new_[85157]_  & \new_[85154]_ ;
  assign \new_[85159]_  = \new_[85158]_  & \new_[85151]_ ;
  assign \new_[85162]_  = ~A235 & ~A233;
  assign \new_[85165]_  = A265 & ~A236;
  assign \new_[85166]_  = \new_[85165]_  & \new_[85162]_ ;
  assign \new_[85169]_  = A298 & A266;
  assign \new_[85173]_  = A301 & A300;
  assign \new_[85174]_  = ~A299 & \new_[85173]_ ;
  assign \new_[85175]_  = \new_[85174]_  & \new_[85169]_ ;
  assign \new_[85176]_  = \new_[85175]_  & \new_[85166]_ ;
  assign \new_[85179]_  = ~A168 & A169;
  assign \new_[85182]_  = ~A166 & A167;
  assign \new_[85183]_  = \new_[85182]_  & \new_[85179]_ ;
  assign \new_[85186]_  = ~A200 & A199;
  assign \new_[85189]_  = A202 & A201;
  assign \new_[85190]_  = \new_[85189]_  & \new_[85186]_ ;
  assign \new_[85191]_  = \new_[85190]_  & \new_[85183]_ ;
  assign \new_[85194]_  = ~A235 & ~A233;
  assign \new_[85197]_  = A265 & ~A236;
  assign \new_[85198]_  = \new_[85197]_  & \new_[85194]_ ;
  assign \new_[85201]_  = A298 & A266;
  assign \new_[85205]_  = A302 & A300;
  assign \new_[85206]_  = ~A299 & \new_[85205]_ ;
  assign \new_[85207]_  = \new_[85206]_  & \new_[85201]_ ;
  assign \new_[85208]_  = \new_[85207]_  & \new_[85198]_ ;
  assign \new_[85211]_  = ~A168 & A169;
  assign \new_[85214]_  = ~A166 & A167;
  assign \new_[85215]_  = \new_[85214]_  & \new_[85211]_ ;
  assign \new_[85218]_  = ~A200 & A199;
  assign \new_[85221]_  = A202 & A201;
  assign \new_[85222]_  = \new_[85221]_  & \new_[85218]_ ;
  assign \new_[85223]_  = \new_[85222]_  & \new_[85215]_ ;
  assign \new_[85226]_  = ~A235 & ~A233;
  assign \new_[85229]_  = ~A266 & ~A236;
  assign \new_[85230]_  = \new_[85229]_  & \new_[85226]_ ;
  assign \new_[85233]_  = A298 & ~A267;
  assign \new_[85237]_  = A301 & A300;
  assign \new_[85238]_  = ~A299 & \new_[85237]_ ;
  assign \new_[85239]_  = \new_[85238]_  & \new_[85233]_ ;
  assign \new_[85240]_  = \new_[85239]_  & \new_[85230]_ ;
  assign \new_[85243]_  = ~A168 & A169;
  assign \new_[85246]_  = ~A166 & A167;
  assign \new_[85247]_  = \new_[85246]_  & \new_[85243]_ ;
  assign \new_[85250]_  = ~A200 & A199;
  assign \new_[85253]_  = A202 & A201;
  assign \new_[85254]_  = \new_[85253]_  & \new_[85250]_ ;
  assign \new_[85255]_  = \new_[85254]_  & \new_[85247]_ ;
  assign \new_[85258]_  = ~A235 & ~A233;
  assign \new_[85261]_  = ~A266 & ~A236;
  assign \new_[85262]_  = \new_[85261]_  & \new_[85258]_ ;
  assign \new_[85265]_  = A298 & ~A267;
  assign \new_[85269]_  = A302 & A300;
  assign \new_[85270]_  = ~A299 & \new_[85269]_ ;
  assign \new_[85271]_  = \new_[85270]_  & \new_[85265]_ ;
  assign \new_[85272]_  = \new_[85271]_  & \new_[85262]_ ;
  assign \new_[85275]_  = ~A168 & A169;
  assign \new_[85278]_  = ~A166 & A167;
  assign \new_[85279]_  = \new_[85278]_  & \new_[85275]_ ;
  assign \new_[85282]_  = ~A200 & A199;
  assign \new_[85285]_  = A202 & A201;
  assign \new_[85286]_  = \new_[85285]_  & \new_[85282]_ ;
  assign \new_[85287]_  = \new_[85286]_  & \new_[85279]_ ;
  assign \new_[85290]_  = ~A235 & ~A233;
  assign \new_[85293]_  = ~A265 & ~A236;
  assign \new_[85294]_  = \new_[85293]_  & \new_[85290]_ ;
  assign \new_[85297]_  = A298 & ~A266;
  assign \new_[85301]_  = A301 & A300;
  assign \new_[85302]_  = ~A299 & \new_[85301]_ ;
  assign \new_[85303]_  = \new_[85302]_  & \new_[85297]_ ;
  assign \new_[85304]_  = \new_[85303]_  & \new_[85294]_ ;
  assign \new_[85307]_  = ~A168 & A169;
  assign \new_[85310]_  = ~A166 & A167;
  assign \new_[85311]_  = \new_[85310]_  & \new_[85307]_ ;
  assign \new_[85314]_  = ~A200 & A199;
  assign \new_[85317]_  = A202 & A201;
  assign \new_[85318]_  = \new_[85317]_  & \new_[85314]_ ;
  assign \new_[85319]_  = \new_[85318]_  & \new_[85311]_ ;
  assign \new_[85322]_  = ~A235 & ~A233;
  assign \new_[85325]_  = ~A265 & ~A236;
  assign \new_[85326]_  = \new_[85325]_  & \new_[85322]_ ;
  assign \new_[85329]_  = A298 & ~A266;
  assign \new_[85333]_  = A302 & A300;
  assign \new_[85334]_  = ~A299 & \new_[85333]_ ;
  assign \new_[85335]_  = \new_[85334]_  & \new_[85329]_ ;
  assign \new_[85336]_  = \new_[85335]_  & \new_[85326]_ ;
  assign \new_[85339]_  = ~A168 & A169;
  assign \new_[85342]_  = ~A166 & A167;
  assign \new_[85343]_  = \new_[85342]_  & \new_[85339]_ ;
  assign \new_[85346]_  = ~A200 & A199;
  assign \new_[85349]_  = A202 & A201;
  assign \new_[85350]_  = \new_[85349]_  & \new_[85346]_ ;
  assign \new_[85351]_  = \new_[85350]_  & \new_[85343]_ ;
  assign \new_[85354]_  = ~A234 & ~A233;
  assign \new_[85357]_  = ~A268 & ~A266;
  assign \new_[85358]_  = \new_[85357]_  & \new_[85354]_ ;
  assign \new_[85361]_  = A298 & ~A269;
  assign \new_[85365]_  = A301 & A300;
  assign \new_[85366]_  = ~A299 & \new_[85365]_ ;
  assign \new_[85367]_  = \new_[85366]_  & \new_[85361]_ ;
  assign \new_[85368]_  = \new_[85367]_  & \new_[85358]_ ;
  assign \new_[85371]_  = ~A168 & A169;
  assign \new_[85374]_  = ~A166 & A167;
  assign \new_[85375]_  = \new_[85374]_  & \new_[85371]_ ;
  assign \new_[85378]_  = ~A200 & A199;
  assign \new_[85381]_  = A202 & A201;
  assign \new_[85382]_  = \new_[85381]_  & \new_[85378]_ ;
  assign \new_[85383]_  = \new_[85382]_  & \new_[85375]_ ;
  assign \new_[85386]_  = ~A234 & ~A233;
  assign \new_[85389]_  = ~A268 & ~A266;
  assign \new_[85390]_  = \new_[85389]_  & \new_[85386]_ ;
  assign \new_[85393]_  = A298 & ~A269;
  assign \new_[85397]_  = A302 & A300;
  assign \new_[85398]_  = ~A299 & \new_[85397]_ ;
  assign \new_[85399]_  = \new_[85398]_  & \new_[85393]_ ;
  assign \new_[85400]_  = \new_[85399]_  & \new_[85390]_ ;
  assign \new_[85403]_  = ~A168 & A169;
  assign \new_[85406]_  = ~A166 & A167;
  assign \new_[85407]_  = \new_[85406]_  & \new_[85403]_ ;
  assign \new_[85410]_  = ~A200 & A199;
  assign \new_[85413]_  = A202 & A201;
  assign \new_[85414]_  = \new_[85413]_  & \new_[85410]_ ;
  assign \new_[85415]_  = \new_[85414]_  & \new_[85407]_ ;
  assign \new_[85418]_  = ~A233 & ~A232;
  assign \new_[85421]_  = ~A268 & ~A266;
  assign \new_[85422]_  = \new_[85421]_  & \new_[85418]_ ;
  assign \new_[85425]_  = A298 & ~A269;
  assign \new_[85429]_  = A301 & A300;
  assign \new_[85430]_  = ~A299 & \new_[85429]_ ;
  assign \new_[85431]_  = \new_[85430]_  & \new_[85425]_ ;
  assign \new_[85432]_  = \new_[85431]_  & \new_[85422]_ ;
  assign \new_[85435]_  = ~A168 & A169;
  assign \new_[85438]_  = ~A166 & A167;
  assign \new_[85439]_  = \new_[85438]_  & \new_[85435]_ ;
  assign \new_[85442]_  = ~A200 & A199;
  assign \new_[85445]_  = A202 & A201;
  assign \new_[85446]_  = \new_[85445]_  & \new_[85442]_ ;
  assign \new_[85447]_  = \new_[85446]_  & \new_[85439]_ ;
  assign \new_[85450]_  = ~A233 & ~A232;
  assign \new_[85453]_  = ~A268 & ~A266;
  assign \new_[85454]_  = \new_[85453]_  & \new_[85450]_ ;
  assign \new_[85457]_  = A298 & ~A269;
  assign \new_[85461]_  = A302 & A300;
  assign \new_[85462]_  = ~A299 & \new_[85461]_ ;
  assign \new_[85463]_  = \new_[85462]_  & \new_[85457]_ ;
  assign \new_[85464]_  = \new_[85463]_  & \new_[85454]_ ;
  assign \new_[85467]_  = ~A168 & A169;
  assign \new_[85470]_  = ~A166 & A167;
  assign \new_[85471]_  = \new_[85470]_  & \new_[85467]_ ;
  assign \new_[85474]_  = ~A200 & A199;
  assign \new_[85477]_  = A203 & A201;
  assign \new_[85478]_  = \new_[85477]_  & \new_[85474]_ ;
  assign \new_[85479]_  = \new_[85478]_  & \new_[85471]_ ;
  assign \new_[85482]_  = A233 & A232;
  assign \new_[85485]_  = ~A268 & A265;
  assign \new_[85486]_  = \new_[85485]_  & \new_[85482]_ ;
  assign \new_[85489]_  = A298 & ~A269;
  assign \new_[85493]_  = A301 & A300;
  assign \new_[85494]_  = ~A299 & \new_[85493]_ ;
  assign \new_[85495]_  = \new_[85494]_  & \new_[85489]_ ;
  assign \new_[85496]_  = \new_[85495]_  & \new_[85486]_ ;
  assign \new_[85499]_  = ~A168 & A169;
  assign \new_[85502]_  = ~A166 & A167;
  assign \new_[85503]_  = \new_[85502]_  & \new_[85499]_ ;
  assign \new_[85506]_  = ~A200 & A199;
  assign \new_[85509]_  = A203 & A201;
  assign \new_[85510]_  = \new_[85509]_  & \new_[85506]_ ;
  assign \new_[85511]_  = \new_[85510]_  & \new_[85503]_ ;
  assign \new_[85514]_  = A233 & A232;
  assign \new_[85517]_  = ~A268 & A265;
  assign \new_[85518]_  = \new_[85517]_  & \new_[85514]_ ;
  assign \new_[85521]_  = A298 & ~A269;
  assign \new_[85525]_  = A302 & A300;
  assign \new_[85526]_  = ~A299 & \new_[85525]_ ;
  assign \new_[85527]_  = \new_[85526]_  & \new_[85521]_ ;
  assign \new_[85528]_  = \new_[85527]_  & \new_[85518]_ ;
  assign \new_[85531]_  = ~A168 & A169;
  assign \new_[85534]_  = ~A166 & A167;
  assign \new_[85535]_  = \new_[85534]_  & \new_[85531]_ ;
  assign \new_[85538]_  = ~A200 & A199;
  assign \new_[85541]_  = A203 & A201;
  assign \new_[85542]_  = \new_[85541]_  & \new_[85538]_ ;
  assign \new_[85543]_  = \new_[85542]_  & \new_[85535]_ ;
  assign \new_[85546]_  = ~A235 & ~A233;
  assign \new_[85549]_  = A265 & ~A236;
  assign \new_[85550]_  = \new_[85549]_  & \new_[85546]_ ;
  assign \new_[85553]_  = A298 & A266;
  assign \new_[85557]_  = A301 & A300;
  assign \new_[85558]_  = ~A299 & \new_[85557]_ ;
  assign \new_[85559]_  = \new_[85558]_  & \new_[85553]_ ;
  assign \new_[85560]_  = \new_[85559]_  & \new_[85550]_ ;
  assign \new_[85563]_  = ~A168 & A169;
  assign \new_[85566]_  = ~A166 & A167;
  assign \new_[85567]_  = \new_[85566]_  & \new_[85563]_ ;
  assign \new_[85570]_  = ~A200 & A199;
  assign \new_[85573]_  = A203 & A201;
  assign \new_[85574]_  = \new_[85573]_  & \new_[85570]_ ;
  assign \new_[85575]_  = \new_[85574]_  & \new_[85567]_ ;
  assign \new_[85578]_  = ~A235 & ~A233;
  assign \new_[85581]_  = A265 & ~A236;
  assign \new_[85582]_  = \new_[85581]_  & \new_[85578]_ ;
  assign \new_[85585]_  = A298 & A266;
  assign \new_[85589]_  = A302 & A300;
  assign \new_[85590]_  = ~A299 & \new_[85589]_ ;
  assign \new_[85591]_  = \new_[85590]_  & \new_[85585]_ ;
  assign \new_[85592]_  = \new_[85591]_  & \new_[85582]_ ;
  assign \new_[85595]_  = ~A168 & A169;
  assign \new_[85598]_  = ~A166 & A167;
  assign \new_[85599]_  = \new_[85598]_  & \new_[85595]_ ;
  assign \new_[85602]_  = ~A200 & A199;
  assign \new_[85605]_  = A203 & A201;
  assign \new_[85606]_  = \new_[85605]_  & \new_[85602]_ ;
  assign \new_[85607]_  = \new_[85606]_  & \new_[85599]_ ;
  assign \new_[85610]_  = ~A235 & ~A233;
  assign \new_[85613]_  = ~A266 & ~A236;
  assign \new_[85614]_  = \new_[85613]_  & \new_[85610]_ ;
  assign \new_[85617]_  = A298 & ~A267;
  assign \new_[85621]_  = A301 & A300;
  assign \new_[85622]_  = ~A299 & \new_[85621]_ ;
  assign \new_[85623]_  = \new_[85622]_  & \new_[85617]_ ;
  assign \new_[85624]_  = \new_[85623]_  & \new_[85614]_ ;
  assign \new_[85627]_  = ~A168 & A169;
  assign \new_[85630]_  = ~A166 & A167;
  assign \new_[85631]_  = \new_[85630]_  & \new_[85627]_ ;
  assign \new_[85634]_  = ~A200 & A199;
  assign \new_[85637]_  = A203 & A201;
  assign \new_[85638]_  = \new_[85637]_  & \new_[85634]_ ;
  assign \new_[85639]_  = \new_[85638]_  & \new_[85631]_ ;
  assign \new_[85642]_  = ~A235 & ~A233;
  assign \new_[85645]_  = ~A266 & ~A236;
  assign \new_[85646]_  = \new_[85645]_  & \new_[85642]_ ;
  assign \new_[85649]_  = A298 & ~A267;
  assign \new_[85653]_  = A302 & A300;
  assign \new_[85654]_  = ~A299 & \new_[85653]_ ;
  assign \new_[85655]_  = \new_[85654]_  & \new_[85649]_ ;
  assign \new_[85656]_  = \new_[85655]_  & \new_[85646]_ ;
  assign \new_[85659]_  = ~A168 & A169;
  assign \new_[85662]_  = ~A166 & A167;
  assign \new_[85663]_  = \new_[85662]_  & \new_[85659]_ ;
  assign \new_[85666]_  = ~A200 & A199;
  assign \new_[85669]_  = A203 & A201;
  assign \new_[85670]_  = \new_[85669]_  & \new_[85666]_ ;
  assign \new_[85671]_  = \new_[85670]_  & \new_[85663]_ ;
  assign \new_[85674]_  = ~A235 & ~A233;
  assign \new_[85677]_  = ~A265 & ~A236;
  assign \new_[85678]_  = \new_[85677]_  & \new_[85674]_ ;
  assign \new_[85681]_  = A298 & ~A266;
  assign \new_[85685]_  = A301 & A300;
  assign \new_[85686]_  = ~A299 & \new_[85685]_ ;
  assign \new_[85687]_  = \new_[85686]_  & \new_[85681]_ ;
  assign \new_[85688]_  = \new_[85687]_  & \new_[85678]_ ;
  assign \new_[85691]_  = ~A168 & A169;
  assign \new_[85694]_  = ~A166 & A167;
  assign \new_[85695]_  = \new_[85694]_  & \new_[85691]_ ;
  assign \new_[85698]_  = ~A200 & A199;
  assign \new_[85701]_  = A203 & A201;
  assign \new_[85702]_  = \new_[85701]_  & \new_[85698]_ ;
  assign \new_[85703]_  = \new_[85702]_  & \new_[85695]_ ;
  assign \new_[85706]_  = ~A235 & ~A233;
  assign \new_[85709]_  = ~A265 & ~A236;
  assign \new_[85710]_  = \new_[85709]_  & \new_[85706]_ ;
  assign \new_[85713]_  = A298 & ~A266;
  assign \new_[85717]_  = A302 & A300;
  assign \new_[85718]_  = ~A299 & \new_[85717]_ ;
  assign \new_[85719]_  = \new_[85718]_  & \new_[85713]_ ;
  assign \new_[85720]_  = \new_[85719]_  & \new_[85710]_ ;
  assign \new_[85723]_  = ~A168 & A169;
  assign \new_[85726]_  = ~A166 & A167;
  assign \new_[85727]_  = \new_[85726]_  & \new_[85723]_ ;
  assign \new_[85730]_  = ~A200 & A199;
  assign \new_[85733]_  = A203 & A201;
  assign \new_[85734]_  = \new_[85733]_  & \new_[85730]_ ;
  assign \new_[85735]_  = \new_[85734]_  & \new_[85727]_ ;
  assign \new_[85738]_  = ~A234 & ~A233;
  assign \new_[85741]_  = ~A268 & ~A266;
  assign \new_[85742]_  = \new_[85741]_  & \new_[85738]_ ;
  assign \new_[85745]_  = A298 & ~A269;
  assign \new_[85749]_  = A301 & A300;
  assign \new_[85750]_  = ~A299 & \new_[85749]_ ;
  assign \new_[85751]_  = \new_[85750]_  & \new_[85745]_ ;
  assign \new_[85752]_  = \new_[85751]_  & \new_[85742]_ ;
  assign \new_[85755]_  = ~A168 & A169;
  assign \new_[85758]_  = ~A166 & A167;
  assign \new_[85759]_  = \new_[85758]_  & \new_[85755]_ ;
  assign \new_[85762]_  = ~A200 & A199;
  assign \new_[85765]_  = A203 & A201;
  assign \new_[85766]_  = \new_[85765]_  & \new_[85762]_ ;
  assign \new_[85767]_  = \new_[85766]_  & \new_[85759]_ ;
  assign \new_[85770]_  = ~A234 & ~A233;
  assign \new_[85773]_  = ~A268 & ~A266;
  assign \new_[85774]_  = \new_[85773]_  & \new_[85770]_ ;
  assign \new_[85777]_  = A298 & ~A269;
  assign \new_[85781]_  = A302 & A300;
  assign \new_[85782]_  = ~A299 & \new_[85781]_ ;
  assign \new_[85783]_  = \new_[85782]_  & \new_[85777]_ ;
  assign \new_[85784]_  = \new_[85783]_  & \new_[85774]_ ;
  assign \new_[85787]_  = ~A168 & A169;
  assign \new_[85790]_  = ~A166 & A167;
  assign \new_[85791]_  = \new_[85790]_  & \new_[85787]_ ;
  assign \new_[85794]_  = ~A200 & A199;
  assign \new_[85797]_  = A203 & A201;
  assign \new_[85798]_  = \new_[85797]_  & \new_[85794]_ ;
  assign \new_[85799]_  = \new_[85798]_  & \new_[85791]_ ;
  assign \new_[85802]_  = ~A233 & ~A232;
  assign \new_[85805]_  = ~A268 & ~A266;
  assign \new_[85806]_  = \new_[85805]_  & \new_[85802]_ ;
  assign \new_[85809]_  = A298 & ~A269;
  assign \new_[85813]_  = A301 & A300;
  assign \new_[85814]_  = ~A299 & \new_[85813]_ ;
  assign \new_[85815]_  = \new_[85814]_  & \new_[85809]_ ;
  assign \new_[85816]_  = \new_[85815]_  & \new_[85806]_ ;
  assign \new_[85819]_  = ~A168 & A169;
  assign \new_[85822]_  = ~A166 & A167;
  assign \new_[85823]_  = \new_[85822]_  & \new_[85819]_ ;
  assign \new_[85826]_  = ~A200 & A199;
  assign \new_[85829]_  = A203 & A201;
  assign \new_[85830]_  = \new_[85829]_  & \new_[85826]_ ;
  assign \new_[85831]_  = \new_[85830]_  & \new_[85823]_ ;
  assign \new_[85834]_  = ~A233 & ~A232;
  assign \new_[85837]_  = ~A268 & ~A266;
  assign \new_[85838]_  = \new_[85837]_  & \new_[85834]_ ;
  assign \new_[85841]_  = A298 & ~A269;
  assign \new_[85845]_  = A302 & A300;
  assign \new_[85846]_  = ~A299 & \new_[85845]_ ;
  assign \new_[85847]_  = \new_[85846]_  & \new_[85841]_ ;
  assign \new_[85848]_  = \new_[85847]_  & \new_[85838]_ ;
  assign \new_[85851]_  = ~A168 & A169;
  assign \new_[85854]_  = A166 & ~A167;
  assign \new_[85855]_  = \new_[85854]_  & \new_[85851]_ ;
  assign \new_[85858]_  = ~A200 & A199;
  assign \new_[85861]_  = A202 & A201;
  assign \new_[85862]_  = \new_[85861]_  & \new_[85858]_ ;
  assign \new_[85863]_  = \new_[85862]_  & \new_[85855]_ ;
  assign \new_[85866]_  = A233 & A232;
  assign \new_[85869]_  = ~A268 & A265;
  assign \new_[85870]_  = \new_[85869]_  & \new_[85866]_ ;
  assign \new_[85873]_  = A298 & ~A269;
  assign \new_[85877]_  = A301 & A300;
  assign \new_[85878]_  = ~A299 & \new_[85877]_ ;
  assign \new_[85879]_  = \new_[85878]_  & \new_[85873]_ ;
  assign \new_[85880]_  = \new_[85879]_  & \new_[85870]_ ;
  assign \new_[85883]_  = ~A168 & A169;
  assign \new_[85886]_  = A166 & ~A167;
  assign \new_[85887]_  = \new_[85886]_  & \new_[85883]_ ;
  assign \new_[85890]_  = ~A200 & A199;
  assign \new_[85893]_  = A202 & A201;
  assign \new_[85894]_  = \new_[85893]_  & \new_[85890]_ ;
  assign \new_[85895]_  = \new_[85894]_  & \new_[85887]_ ;
  assign \new_[85898]_  = A233 & A232;
  assign \new_[85901]_  = ~A268 & A265;
  assign \new_[85902]_  = \new_[85901]_  & \new_[85898]_ ;
  assign \new_[85905]_  = A298 & ~A269;
  assign \new_[85909]_  = A302 & A300;
  assign \new_[85910]_  = ~A299 & \new_[85909]_ ;
  assign \new_[85911]_  = \new_[85910]_  & \new_[85905]_ ;
  assign \new_[85912]_  = \new_[85911]_  & \new_[85902]_ ;
  assign \new_[85915]_  = ~A168 & A169;
  assign \new_[85918]_  = A166 & ~A167;
  assign \new_[85919]_  = \new_[85918]_  & \new_[85915]_ ;
  assign \new_[85922]_  = ~A200 & A199;
  assign \new_[85925]_  = A202 & A201;
  assign \new_[85926]_  = \new_[85925]_  & \new_[85922]_ ;
  assign \new_[85927]_  = \new_[85926]_  & \new_[85919]_ ;
  assign \new_[85930]_  = ~A235 & ~A233;
  assign \new_[85933]_  = A265 & ~A236;
  assign \new_[85934]_  = \new_[85933]_  & \new_[85930]_ ;
  assign \new_[85937]_  = A298 & A266;
  assign \new_[85941]_  = A301 & A300;
  assign \new_[85942]_  = ~A299 & \new_[85941]_ ;
  assign \new_[85943]_  = \new_[85942]_  & \new_[85937]_ ;
  assign \new_[85944]_  = \new_[85943]_  & \new_[85934]_ ;
  assign \new_[85947]_  = ~A168 & A169;
  assign \new_[85950]_  = A166 & ~A167;
  assign \new_[85951]_  = \new_[85950]_  & \new_[85947]_ ;
  assign \new_[85954]_  = ~A200 & A199;
  assign \new_[85957]_  = A202 & A201;
  assign \new_[85958]_  = \new_[85957]_  & \new_[85954]_ ;
  assign \new_[85959]_  = \new_[85958]_  & \new_[85951]_ ;
  assign \new_[85962]_  = ~A235 & ~A233;
  assign \new_[85965]_  = A265 & ~A236;
  assign \new_[85966]_  = \new_[85965]_  & \new_[85962]_ ;
  assign \new_[85969]_  = A298 & A266;
  assign \new_[85973]_  = A302 & A300;
  assign \new_[85974]_  = ~A299 & \new_[85973]_ ;
  assign \new_[85975]_  = \new_[85974]_  & \new_[85969]_ ;
  assign \new_[85976]_  = \new_[85975]_  & \new_[85966]_ ;
  assign \new_[85979]_  = ~A168 & A169;
  assign \new_[85982]_  = A166 & ~A167;
  assign \new_[85983]_  = \new_[85982]_  & \new_[85979]_ ;
  assign \new_[85986]_  = ~A200 & A199;
  assign \new_[85989]_  = A202 & A201;
  assign \new_[85990]_  = \new_[85989]_  & \new_[85986]_ ;
  assign \new_[85991]_  = \new_[85990]_  & \new_[85983]_ ;
  assign \new_[85994]_  = ~A235 & ~A233;
  assign \new_[85997]_  = ~A266 & ~A236;
  assign \new_[85998]_  = \new_[85997]_  & \new_[85994]_ ;
  assign \new_[86001]_  = A298 & ~A267;
  assign \new_[86005]_  = A301 & A300;
  assign \new_[86006]_  = ~A299 & \new_[86005]_ ;
  assign \new_[86007]_  = \new_[86006]_  & \new_[86001]_ ;
  assign \new_[86008]_  = \new_[86007]_  & \new_[85998]_ ;
  assign \new_[86011]_  = ~A168 & A169;
  assign \new_[86014]_  = A166 & ~A167;
  assign \new_[86015]_  = \new_[86014]_  & \new_[86011]_ ;
  assign \new_[86018]_  = ~A200 & A199;
  assign \new_[86021]_  = A202 & A201;
  assign \new_[86022]_  = \new_[86021]_  & \new_[86018]_ ;
  assign \new_[86023]_  = \new_[86022]_  & \new_[86015]_ ;
  assign \new_[86026]_  = ~A235 & ~A233;
  assign \new_[86029]_  = ~A266 & ~A236;
  assign \new_[86030]_  = \new_[86029]_  & \new_[86026]_ ;
  assign \new_[86033]_  = A298 & ~A267;
  assign \new_[86037]_  = A302 & A300;
  assign \new_[86038]_  = ~A299 & \new_[86037]_ ;
  assign \new_[86039]_  = \new_[86038]_  & \new_[86033]_ ;
  assign \new_[86040]_  = \new_[86039]_  & \new_[86030]_ ;
  assign \new_[86043]_  = ~A168 & A169;
  assign \new_[86046]_  = A166 & ~A167;
  assign \new_[86047]_  = \new_[86046]_  & \new_[86043]_ ;
  assign \new_[86050]_  = ~A200 & A199;
  assign \new_[86053]_  = A202 & A201;
  assign \new_[86054]_  = \new_[86053]_  & \new_[86050]_ ;
  assign \new_[86055]_  = \new_[86054]_  & \new_[86047]_ ;
  assign \new_[86058]_  = ~A235 & ~A233;
  assign \new_[86061]_  = ~A265 & ~A236;
  assign \new_[86062]_  = \new_[86061]_  & \new_[86058]_ ;
  assign \new_[86065]_  = A298 & ~A266;
  assign \new_[86069]_  = A301 & A300;
  assign \new_[86070]_  = ~A299 & \new_[86069]_ ;
  assign \new_[86071]_  = \new_[86070]_  & \new_[86065]_ ;
  assign \new_[86072]_  = \new_[86071]_  & \new_[86062]_ ;
  assign \new_[86075]_  = ~A168 & A169;
  assign \new_[86078]_  = A166 & ~A167;
  assign \new_[86079]_  = \new_[86078]_  & \new_[86075]_ ;
  assign \new_[86082]_  = ~A200 & A199;
  assign \new_[86085]_  = A202 & A201;
  assign \new_[86086]_  = \new_[86085]_  & \new_[86082]_ ;
  assign \new_[86087]_  = \new_[86086]_  & \new_[86079]_ ;
  assign \new_[86090]_  = ~A235 & ~A233;
  assign \new_[86093]_  = ~A265 & ~A236;
  assign \new_[86094]_  = \new_[86093]_  & \new_[86090]_ ;
  assign \new_[86097]_  = A298 & ~A266;
  assign \new_[86101]_  = A302 & A300;
  assign \new_[86102]_  = ~A299 & \new_[86101]_ ;
  assign \new_[86103]_  = \new_[86102]_  & \new_[86097]_ ;
  assign \new_[86104]_  = \new_[86103]_  & \new_[86094]_ ;
  assign \new_[86107]_  = ~A168 & A169;
  assign \new_[86110]_  = A166 & ~A167;
  assign \new_[86111]_  = \new_[86110]_  & \new_[86107]_ ;
  assign \new_[86114]_  = ~A200 & A199;
  assign \new_[86117]_  = A202 & A201;
  assign \new_[86118]_  = \new_[86117]_  & \new_[86114]_ ;
  assign \new_[86119]_  = \new_[86118]_  & \new_[86111]_ ;
  assign \new_[86122]_  = ~A234 & ~A233;
  assign \new_[86125]_  = ~A268 & ~A266;
  assign \new_[86126]_  = \new_[86125]_  & \new_[86122]_ ;
  assign \new_[86129]_  = A298 & ~A269;
  assign \new_[86133]_  = A301 & A300;
  assign \new_[86134]_  = ~A299 & \new_[86133]_ ;
  assign \new_[86135]_  = \new_[86134]_  & \new_[86129]_ ;
  assign \new_[86136]_  = \new_[86135]_  & \new_[86126]_ ;
  assign \new_[86139]_  = ~A168 & A169;
  assign \new_[86142]_  = A166 & ~A167;
  assign \new_[86143]_  = \new_[86142]_  & \new_[86139]_ ;
  assign \new_[86146]_  = ~A200 & A199;
  assign \new_[86149]_  = A202 & A201;
  assign \new_[86150]_  = \new_[86149]_  & \new_[86146]_ ;
  assign \new_[86151]_  = \new_[86150]_  & \new_[86143]_ ;
  assign \new_[86154]_  = ~A234 & ~A233;
  assign \new_[86157]_  = ~A268 & ~A266;
  assign \new_[86158]_  = \new_[86157]_  & \new_[86154]_ ;
  assign \new_[86161]_  = A298 & ~A269;
  assign \new_[86165]_  = A302 & A300;
  assign \new_[86166]_  = ~A299 & \new_[86165]_ ;
  assign \new_[86167]_  = \new_[86166]_  & \new_[86161]_ ;
  assign \new_[86168]_  = \new_[86167]_  & \new_[86158]_ ;
  assign \new_[86171]_  = ~A168 & A169;
  assign \new_[86174]_  = A166 & ~A167;
  assign \new_[86175]_  = \new_[86174]_  & \new_[86171]_ ;
  assign \new_[86178]_  = ~A200 & A199;
  assign \new_[86181]_  = A202 & A201;
  assign \new_[86182]_  = \new_[86181]_  & \new_[86178]_ ;
  assign \new_[86183]_  = \new_[86182]_  & \new_[86175]_ ;
  assign \new_[86186]_  = ~A233 & ~A232;
  assign \new_[86189]_  = ~A268 & ~A266;
  assign \new_[86190]_  = \new_[86189]_  & \new_[86186]_ ;
  assign \new_[86193]_  = A298 & ~A269;
  assign \new_[86197]_  = A301 & A300;
  assign \new_[86198]_  = ~A299 & \new_[86197]_ ;
  assign \new_[86199]_  = \new_[86198]_  & \new_[86193]_ ;
  assign \new_[86200]_  = \new_[86199]_  & \new_[86190]_ ;
  assign \new_[86203]_  = ~A168 & A169;
  assign \new_[86206]_  = A166 & ~A167;
  assign \new_[86207]_  = \new_[86206]_  & \new_[86203]_ ;
  assign \new_[86210]_  = ~A200 & A199;
  assign \new_[86213]_  = A202 & A201;
  assign \new_[86214]_  = \new_[86213]_  & \new_[86210]_ ;
  assign \new_[86215]_  = \new_[86214]_  & \new_[86207]_ ;
  assign \new_[86218]_  = ~A233 & ~A232;
  assign \new_[86221]_  = ~A268 & ~A266;
  assign \new_[86222]_  = \new_[86221]_  & \new_[86218]_ ;
  assign \new_[86225]_  = A298 & ~A269;
  assign \new_[86229]_  = A302 & A300;
  assign \new_[86230]_  = ~A299 & \new_[86229]_ ;
  assign \new_[86231]_  = \new_[86230]_  & \new_[86225]_ ;
  assign \new_[86232]_  = \new_[86231]_  & \new_[86222]_ ;
  assign \new_[86235]_  = ~A168 & A169;
  assign \new_[86238]_  = A166 & ~A167;
  assign \new_[86239]_  = \new_[86238]_  & \new_[86235]_ ;
  assign \new_[86242]_  = ~A200 & A199;
  assign \new_[86245]_  = A203 & A201;
  assign \new_[86246]_  = \new_[86245]_  & \new_[86242]_ ;
  assign \new_[86247]_  = \new_[86246]_  & \new_[86239]_ ;
  assign \new_[86250]_  = A233 & A232;
  assign \new_[86253]_  = ~A268 & A265;
  assign \new_[86254]_  = \new_[86253]_  & \new_[86250]_ ;
  assign \new_[86257]_  = A298 & ~A269;
  assign \new_[86261]_  = A301 & A300;
  assign \new_[86262]_  = ~A299 & \new_[86261]_ ;
  assign \new_[86263]_  = \new_[86262]_  & \new_[86257]_ ;
  assign \new_[86264]_  = \new_[86263]_  & \new_[86254]_ ;
  assign \new_[86267]_  = ~A168 & A169;
  assign \new_[86270]_  = A166 & ~A167;
  assign \new_[86271]_  = \new_[86270]_  & \new_[86267]_ ;
  assign \new_[86274]_  = ~A200 & A199;
  assign \new_[86277]_  = A203 & A201;
  assign \new_[86278]_  = \new_[86277]_  & \new_[86274]_ ;
  assign \new_[86279]_  = \new_[86278]_  & \new_[86271]_ ;
  assign \new_[86282]_  = A233 & A232;
  assign \new_[86285]_  = ~A268 & A265;
  assign \new_[86286]_  = \new_[86285]_  & \new_[86282]_ ;
  assign \new_[86289]_  = A298 & ~A269;
  assign \new_[86293]_  = A302 & A300;
  assign \new_[86294]_  = ~A299 & \new_[86293]_ ;
  assign \new_[86295]_  = \new_[86294]_  & \new_[86289]_ ;
  assign \new_[86296]_  = \new_[86295]_  & \new_[86286]_ ;
  assign \new_[86299]_  = ~A168 & A169;
  assign \new_[86302]_  = A166 & ~A167;
  assign \new_[86303]_  = \new_[86302]_  & \new_[86299]_ ;
  assign \new_[86306]_  = ~A200 & A199;
  assign \new_[86309]_  = A203 & A201;
  assign \new_[86310]_  = \new_[86309]_  & \new_[86306]_ ;
  assign \new_[86311]_  = \new_[86310]_  & \new_[86303]_ ;
  assign \new_[86314]_  = ~A235 & ~A233;
  assign \new_[86317]_  = A265 & ~A236;
  assign \new_[86318]_  = \new_[86317]_  & \new_[86314]_ ;
  assign \new_[86321]_  = A298 & A266;
  assign \new_[86325]_  = A301 & A300;
  assign \new_[86326]_  = ~A299 & \new_[86325]_ ;
  assign \new_[86327]_  = \new_[86326]_  & \new_[86321]_ ;
  assign \new_[86328]_  = \new_[86327]_  & \new_[86318]_ ;
  assign \new_[86331]_  = ~A168 & A169;
  assign \new_[86334]_  = A166 & ~A167;
  assign \new_[86335]_  = \new_[86334]_  & \new_[86331]_ ;
  assign \new_[86338]_  = ~A200 & A199;
  assign \new_[86341]_  = A203 & A201;
  assign \new_[86342]_  = \new_[86341]_  & \new_[86338]_ ;
  assign \new_[86343]_  = \new_[86342]_  & \new_[86335]_ ;
  assign \new_[86346]_  = ~A235 & ~A233;
  assign \new_[86349]_  = A265 & ~A236;
  assign \new_[86350]_  = \new_[86349]_  & \new_[86346]_ ;
  assign \new_[86353]_  = A298 & A266;
  assign \new_[86357]_  = A302 & A300;
  assign \new_[86358]_  = ~A299 & \new_[86357]_ ;
  assign \new_[86359]_  = \new_[86358]_  & \new_[86353]_ ;
  assign \new_[86360]_  = \new_[86359]_  & \new_[86350]_ ;
  assign \new_[86363]_  = ~A168 & A169;
  assign \new_[86366]_  = A166 & ~A167;
  assign \new_[86367]_  = \new_[86366]_  & \new_[86363]_ ;
  assign \new_[86370]_  = ~A200 & A199;
  assign \new_[86373]_  = A203 & A201;
  assign \new_[86374]_  = \new_[86373]_  & \new_[86370]_ ;
  assign \new_[86375]_  = \new_[86374]_  & \new_[86367]_ ;
  assign \new_[86378]_  = ~A235 & ~A233;
  assign \new_[86381]_  = ~A266 & ~A236;
  assign \new_[86382]_  = \new_[86381]_  & \new_[86378]_ ;
  assign \new_[86385]_  = A298 & ~A267;
  assign \new_[86389]_  = A301 & A300;
  assign \new_[86390]_  = ~A299 & \new_[86389]_ ;
  assign \new_[86391]_  = \new_[86390]_  & \new_[86385]_ ;
  assign \new_[86392]_  = \new_[86391]_  & \new_[86382]_ ;
  assign \new_[86395]_  = ~A168 & A169;
  assign \new_[86398]_  = A166 & ~A167;
  assign \new_[86399]_  = \new_[86398]_  & \new_[86395]_ ;
  assign \new_[86402]_  = ~A200 & A199;
  assign \new_[86405]_  = A203 & A201;
  assign \new_[86406]_  = \new_[86405]_  & \new_[86402]_ ;
  assign \new_[86407]_  = \new_[86406]_  & \new_[86399]_ ;
  assign \new_[86410]_  = ~A235 & ~A233;
  assign \new_[86413]_  = ~A266 & ~A236;
  assign \new_[86414]_  = \new_[86413]_  & \new_[86410]_ ;
  assign \new_[86417]_  = A298 & ~A267;
  assign \new_[86421]_  = A302 & A300;
  assign \new_[86422]_  = ~A299 & \new_[86421]_ ;
  assign \new_[86423]_  = \new_[86422]_  & \new_[86417]_ ;
  assign \new_[86424]_  = \new_[86423]_  & \new_[86414]_ ;
  assign \new_[86427]_  = ~A168 & A169;
  assign \new_[86430]_  = A166 & ~A167;
  assign \new_[86431]_  = \new_[86430]_  & \new_[86427]_ ;
  assign \new_[86434]_  = ~A200 & A199;
  assign \new_[86437]_  = A203 & A201;
  assign \new_[86438]_  = \new_[86437]_  & \new_[86434]_ ;
  assign \new_[86439]_  = \new_[86438]_  & \new_[86431]_ ;
  assign \new_[86442]_  = ~A235 & ~A233;
  assign \new_[86445]_  = ~A265 & ~A236;
  assign \new_[86446]_  = \new_[86445]_  & \new_[86442]_ ;
  assign \new_[86449]_  = A298 & ~A266;
  assign \new_[86453]_  = A301 & A300;
  assign \new_[86454]_  = ~A299 & \new_[86453]_ ;
  assign \new_[86455]_  = \new_[86454]_  & \new_[86449]_ ;
  assign \new_[86456]_  = \new_[86455]_  & \new_[86446]_ ;
  assign \new_[86459]_  = ~A168 & A169;
  assign \new_[86462]_  = A166 & ~A167;
  assign \new_[86463]_  = \new_[86462]_  & \new_[86459]_ ;
  assign \new_[86466]_  = ~A200 & A199;
  assign \new_[86469]_  = A203 & A201;
  assign \new_[86470]_  = \new_[86469]_  & \new_[86466]_ ;
  assign \new_[86471]_  = \new_[86470]_  & \new_[86463]_ ;
  assign \new_[86474]_  = ~A235 & ~A233;
  assign \new_[86477]_  = ~A265 & ~A236;
  assign \new_[86478]_  = \new_[86477]_  & \new_[86474]_ ;
  assign \new_[86481]_  = A298 & ~A266;
  assign \new_[86485]_  = A302 & A300;
  assign \new_[86486]_  = ~A299 & \new_[86485]_ ;
  assign \new_[86487]_  = \new_[86486]_  & \new_[86481]_ ;
  assign \new_[86488]_  = \new_[86487]_  & \new_[86478]_ ;
  assign \new_[86491]_  = ~A168 & A169;
  assign \new_[86494]_  = A166 & ~A167;
  assign \new_[86495]_  = \new_[86494]_  & \new_[86491]_ ;
  assign \new_[86498]_  = ~A200 & A199;
  assign \new_[86501]_  = A203 & A201;
  assign \new_[86502]_  = \new_[86501]_  & \new_[86498]_ ;
  assign \new_[86503]_  = \new_[86502]_  & \new_[86495]_ ;
  assign \new_[86506]_  = ~A234 & ~A233;
  assign \new_[86509]_  = ~A268 & ~A266;
  assign \new_[86510]_  = \new_[86509]_  & \new_[86506]_ ;
  assign \new_[86513]_  = A298 & ~A269;
  assign \new_[86517]_  = A301 & A300;
  assign \new_[86518]_  = ~A299 & \new_[86517]_ ;
  assign \new_[86519]_  = \new_[86518]_  & \new_[86513]_ ;
  assign \new_[86520]_  = \new_[86519]_  & \new_[86510]_ ;
  assign \new_[86523]_  = ~A168 & A169;
  assign \new_[86526]_  = A166 & ~A167;
  assign \new_[86527]_  = \new_[86526]_  & \new_[86523]_ ;
  assign \new_[86530]_  = ~A200 & A199;
  assign \new_[86533]_  = A203 & A201;
  assign \new_[86534]_  = \new_[86533]_  & \new_[86530]_ ;
  assign \new_[86535]_  = \new_[86534]_  & \new_[86527]_ ;
  assign \new_[86538]_  = ~A234 & ~A233;
  assign \new_[86541]_  = ~A268 & ~A266;
  assign \new_[86542]_  = \new_[86541]_  & \new_[86538]_ ;
  assign \new_[86545]_  = A298 & ~A269;
  assign \new_[86549]_  = A302 & A300;
  assign \new_[86550]_  = ~A299 & \new_[86549]_ ;
  assign \new_[86551]_  = \new_[86550]_  & \new_[86545]_ ;
  assign \new_[86552]_  = \new_[86551]_  & \new_[86542]_ ;
  assign \new_[86555]_  = ~A168 & A169;
  assign \new_[86558]_  = A166 & ~A167;
  assign \new_[86559]_  = \new_[86558]_  & \new_[86555]_ ;
  assign \new_[86562]_  = ~A200 & A199;
  assign \new_[86565]_  = A203 & A201;
  assign \new_[86566]_  = \new_[86565]_  & \new_[86562]_ ;
  assign \new_[86567]_  = \new_[86566]_  & \new_[86559]_ ;
  assign \new_[86570]_  = ~A233 & ~A232;
  assign \new_[86573]_  = ~A268 & ~A266;
  assign \new_[86574]_  = \new_[86573]_  & \new_[86570]_ ;
  assign \new_[86577]_  = A298 & ~A269;
  assign \new_[86581]_  = A301 & A300;
  assign \new_[86582]_  = ~A299 & \new_[86581]_ ;
  assign \new_[86583]_  = \new_[86582]_  & \new_[86577]_ ;
  assign \new_[86584]_  = \new_[86583]_  & \new_[86574]_ ;
  assign \new_[86587]_  = ~A168 & A169;
  assign \new_[86590]_  = A166 & ~A167;
  assign \new_[86591]_  = \new_[86590]_  & \new_[86587]_ ;
  assign \new_[86594]_  = ~A200 & A199;
  assign \new_[86597]_  = A203 & A201;
  assign \new_[86598]_  = \new_[86597]_  & \new_[86594]_ ;
  assign \new_[86599]_  = \new_[86598]_  & \new_[86591]_ ;
  assign \new_[86602]_  = ~A233 & ~A232;
  assign \new_[86605]_  = ~A268 & ~A266;
  assign \new_[86606]_  = \new_[86605]_  & \new_[86602]_ ;
  assign \new_[86609]_  = A298 & ~A269;
  assign \new_[86613]_  = A302 & A300;
  assign \new_[86614]_  = ~A299 & \new_[86613]_ ;
  assign \new_[86615]_  = \new_[86614]_  & \new_[86609]_ ;
  assign \new_[86616]_  = \new_[86615]_  & \new_[86606]_ ;
  assign \new_[86619]_  = A169 & A170;
  assign \new_[86622]_  = A199 & ~A168;
  assign \new_[86623]_  = \new_[86622]_  & \new_[86619]_ ;
  assign \new_[86626]_  = A201 & ~A200;
  assign \new_[86629]_  = ~A233 & A202;
  assign \new_[86630]_  = \new_[86629]_  & \new_[86626]_ ;
  assign \new_[86631]_  = \new_[86630]_  & \new_[86623]_ ;
  assign \new_[86634]_  = ~A236 & ~A235;
  assign \new_[86637]_  = ~A268 & ~A266;
  assign \new_[86638]_  = \new_[86637]_  & \new_[86634]_ ;
  assign \new_[86641]_  = A298 & ~A269;
  assign \new_[86645]_  = A301 & A300;
  assign \new_[86646]_  = ~A299 & \new_[86645]_ ;
  assign \new_[86647]_  = \new_[86646]_  & \new_[86641]_ ;
  assign \new_[86648]_  = \new_[86647]_  & \new_[86638]_ ;
  assign \new_[86651]_  = A169 & A170;
  assign \new_[86654]_  = A199 & ~A168;
  assign \new_[86655]_  = \new_[86654]_  & \new_[86651]_ ;
  assign \new_[86658]_  = A201 & ~A200;
  assign \new_[86661]_  = ~A233 & A202;
  assign \new_[86662]_  = \new_[86661]_  & \new_[86658]_ ;
  assign \new_[86663]_  = \new_[86662]_  & \new_[86655]_ ;
  assign \new_[86666]_  = ~A236 & ~A235;
  assign \new_[86669]_  = ~A268 & ~A266;
  assign \new_[86670]_  = \new_[86669]_  & \new_[86666]_ ;
  assign \new_[86673]_  = A298 & ~A269;
  assign \new_[86677]_  = A302 & A300;
  assign \new_[86678]_  = ~A299 & \new_[86677]_ ;
  assign \new_[86679]_  = \new_[86678]_  & \new_[86673]_ ;
  assign \new_[86680]_  = \new_[86679]_  & \new_[86670]_ ;
  assign \new_[86683]_  = A169 & A170;
  assign \new_[86686]_  = A199 & ~A168;
  assign \new_[86687]_  = \new_[86686]_  & \new_[86683]_ ;
  assign \new_[86690]_  = A201 & ~A200;
  assign \new_[86693]_  = ~A233 & A203;
  assign \new_[86694]_  = \new_[86693]_  & \new_[86690]_ ;
  assign \new_[86695]_  = \new_[86694]_  & \new_[86687]_ ;
  assign \new_[86698]_  = ~A236 & ~A235;
  assign \new_[86701]_  = ~A268 & ~A266;
  assign \new_[86702]_  = \new_[86701]_  & \new_[86698]_ ;
  assign \new_[86705]_  = A298 & ~A269;
  assign \new_[86709]_  = A301 & A300;
  assign \new_[86710]_  = ~A299 & \new_[86709]_ ;
  assign \new_[86711]_  = \new_[86710]_  & \new_[86705]_ ;
  assign \new_[86712]_  = \new_[86711]_  & \new_[86702]_ ;
  assign \new_[86715]_  = A169 & A170;
  assign \new_[86718]_  = A199 & ~A168;
  assign \new_[86719]_  = \new_[86718]_  & \new_[86715]_ ;
  assign \new_[86722]_  = A201 & ~A200;
  assign \new_[86725]_  = ~A233 & A203;
  assign \new_[86726]_  = \new_[86725]_  & \new_[86722]_ ;
  assign \new_[86727]_  = \new_[86726]_  & \new_[86719]_ ;
  assign \new_[86730]_  = ~A236 & ~A235;
  assign \new_[86733]_  = ~A268 & ~A266;
  assign \new_[86734]_  = \new_[86733]_  & \new_[86730]_ ;
  assign \new_[86737]_  = A298 & ~A269;
  assign \new_[86741]_  = A302 & A300;
  assign \new_[86742]_  = ~A299 & \new_[86741]_ ;
  assign \new_[86743]_  = \new_[86742]_  & \new_[86737]_ ;
  assign \new_[86744]_  = \new_[86743]_  & \new_[86734]_ ;
  assign \new_[86747]_  = A169 & A170;
  assign \new_[86750]_  = A166 & ~A168;
  assign \new_[86751]_  = \new_[86750]_  & \new_[86747]_ ;
  assign \new_[86754]_  = ~A200 & A199;
  assign \new_[86757]_  = A202 & A201;
  assign \new_[86758]_  = \new_[86757]_  & \new_[86754]_ ;
  assign \new_[86759]_  = \new_[86758]_  & \new_[86751]_ ;
  assign \new_[86762]_  = ~A234 & ~A233;
  assign \new_[86765]_  = ~A268 & ~A266;
  assign \new_[86766]_  = \new_[86765]_  & \new_[86762]_ ;
  assign \new_[86769]_  = A298 & ~A269;
  assign \new_[86773]_  = A301 & A300;
  assign \new_[86774]_  = ~A299 & \new_[86773]_ ;
  assign \new_[86775]_  = \new_[86774]_  & \new_[86769]_ ;
  assign \new_[86776]_  = \new_[86775]_  & \new_[86766]_ ;
  assign \new_[86779]_  = A169 & A170;
  assign \new_[86782]_  = A166 & ~A168;
  assign \new_[86783]_  = \new_[86782]_  & \new_[86779]_ ;
  assign \new_[86786]_  = ~A200 & A199;
  assign \new_[86789]_  = A202 & A201;
  assign \new_[86790]_  = \new_[86789]_  & \new_[86786]_ ;
  assign \new_[86791]_  = \new_[86790]_  & \new_[86783]_ ;
  assign \new_[86794]_  = ~A234 & ~A233;
  assign \new_[86797]_  = ~A268 & ~A266;
  assign \new_[86798]_  = \new_[86797]_  & \new_[86794]_ ;
  assign \new_[86801]_  = A298 & ~A269;
  assign \new_[86805]_  = A302 & A300;
  assign \new_[86806]_  = ~A299 & \new_[86805]_ ;
  assign \new_[86807]_  = \new_[86806]_  & \new_[86801]_ ;
  assign \new_[86808]_  = \new_[86807]_  & \new_[86798]_ ;
  assign \new_[86811]_  = A169 & A170;
  assign \new_[86814]_  = A166 & ~A168;
  assign \new_[86815]_  = \new_[86814]_  & \new_[86811]_ ;
  assign \new_[86818]_  = ~A200 & A199;
  assign \new_[86821]_  = A202 & A201;
  assign \new_[86822]_  = \new_[86821]_  & \new_[86818]_ ;
  assign \new_[86823]_  = \new_[86822]_  & \new_[86815]_ ;
  assign \new_[86826]_  = ~A233 & ~A232;
  assign \new_[86829]_  = ~A268 & ~A266;
  assign \new_[86830]_  = \new_[86829]_  & \new_[86826]_ ;
  assign \new_[86833]_  = A298 & ~A269;
  assign \new_[86837]_  = A301 & A300;
  assign \new_[86838]_  = ~A299 & \new_[86837]_ ;
  assign \new_[86839]_  = \new_[86838]_  & \new_[86833]_ ;
  assign \new_[86840]_  = \new_[86839]_  & \new_[86830]_ ;
  assign \new_[86843]_  = A169 & A170;
  assign \new_[86846]_  = A166 & ~A168;
  assign \new_[86847]_  = \new_[86846]_  & \new_[86843]_ ;
  assign \new_[86850]_  = ~A200 & A199;
  assign \new_[86853]_  = A202 & A201;
  assign \new_[86854]_  = \new_[86853]_  & \new_[86850]_ ;
  assign \new_[86855]_  = \new_[86854]_  & \new_[86847]_ ;
  assign \new_[86858]_  = ~A233 & ~A232;
  assign \new_[86861]_  = ~A268 & ~A266;
  assign \new_[86862]_  = \new_[86861]_  & \new_[86858]_ ;
  assign \new_[86865]_  = A298 & ~A269;
  assign \new_[86869]_  = A302 & A300;
  assign \new_[86870]_  = ~A299 & \new_[86869]_ ;
  assign \new_[86871]_  = \new_[86870]_  & \new_[86865]_ ;
  assign \new_[86872]_  = \new_[86871]_  & \new_[86862]_ ;
  assign \new_[86875]_  = A169 & A170;
  assign \new_[86878]_  = A166 & ~A168;
  assign \new_[86879]_  = \new_[86878]_  & \new_[86875]_ ;
  assign \new_[86882]_  = ~A200 & A199;
  assign \new_[86885]_  = A203 & A201;
  assign \new_[86886]_  = \new_[86885]_  & \new_[86882]_ ;
  assign \new_[86887]_  = \new_[86886]_  & \new_[86879]_ ;
  assign \new_[86890]_  = ~A234 & ~A233;
  assign \new_[86893]_  = ~A268 & ~A266;
  assign \new_[86894]_  = \new_[86893]_  & \new_[86890]_ ;
  assign \new_[86897]_  = A298 & ~A269;
  assign \new_[86901]_  = A301 & A300;
  assign \new_[86902]_  = ~A299 & \new_[86901]_ ;
  assign \new_[86903]_  = \new_[86902]_  & \new_[86897]_ ;
  assign \new_[86904]_  = \new_[86903]_  & \new_[86894]_ ;
  assign \new_[86907]_  = A169 & A170;
  assign \new_[86910]_  = A166 & ~A168;
  assign \new_[86911]_  = \new_[86910]_  & \new_[86907]_ ;
  assign \new_[86914]_  = ~A200 & A199;
  assign \new_[86917]_  = A203 & A201;
  assign \new_[86918]_  = \new_[86917]_  & \new_[86914]_ ;
  assign \new_[86919]_  = \new_[86918]_  & \new_[86911]_ ;
  assign \new_[86922]_  = ~A234 & ~A233;
  assign \new_[86925]_  = ~A268 & ~A266;
  assign \new_[86926]_  = \new_[86925]_  & \new_[86922]_ ;
  assign \new_[86929]_  = A298 & ~A269;
  assign \new_[86933]_  = A302 & A300;
  assign \new_[86934]_  = ~A299 & \new_[86933]_ ;
  assign \new_[86935]_  = \new_[86934]_  & \new_[86929]_ ;
  assign \new_[86936]_  = \new_[86935]_  & \new_[86926]_ ;
  assign \new_[86939]_  = A169 & A170;
  assign \new_[86942]_  = A166 & ~A168;
  assign \new_[86943]_  = \new_[86942]_  & \new_[86939]_ ;
  assign \new_[86946]_  = ~A200 & A199;
  assign \new_[86949]_  = A203 & A201;
  assign \new_[86950]_  = \new_[86949]_  & \new_[86946]_ ;
  assign \new_[86951]_  = \new_[86950]_  & \new_[86943]_ ;
  assign \new_[86954]_  = ~A233 & ~A232;
  assign \new_[86957]_  = ~A268 & ~A266;
  assign \new_[86958]_  = \new_[86957]_  & \new_[86954]_ ;
  assign \new_[86961]_  = A298 & ~A269;
  assign \new_[86965]_  = A301 & A300;
  assign \new_[86966]_  = ~A299 & \new_[86965]_ ;
  assign \new_[86967]_  = \new_[86966]_  & \new_[86961]_ ;
  assign \new_[86968]_  = \new_[86967]_  & \new_[86958]_ ;
  assign \new_[86971]_  = A169 & A170;
  assign \new_[86974]_  = A166 & ~A168;
  assign \new_[86975]_  = \new_[86974]_  & \new_[86971]_ ;
  assign \new_[86978]_  = ~A200 & A199;
  assign \new_[86981]_  = A203 & A201;
  assign \new_[86982]_  = \new_[86981]_  & \new_[86978]_ ;
  assign \new_[86983]_  = \new_[86982]_  & \new_[86975]_ ;
  assign \new_[86986]_  = ~A233 & ~A232;
  assign \new_[86989]_  = ~A268 & ~A266;
  assign \new_[86990]_  = \new_[86989]_  & \new_[86986]_ ;
  assign \new_[86993]_  = A298 & ~A269;
  assign \new_[86997]_  = A302 & A300;
  assign \new_[86998]_  = ~A299 & \new_[86997]_ ;
  assign \new_[86999]_  = \new_[86998]_  & \new_[86993]_ ;
  assign \new_[87000]_  = \new_[86999]_  & \new_[86990]_ ;
  assign \new_[87003]_  = A169 & ~A170;
  assign \new_[87006]_  = A166 & A167;
  assign \new_[87007]_  = \new_[87006]_  & \new_[87003]_ ;
  assign \new_[87010]_  = ~A202 & ~A200;
  assign \new_[87013]_  = ~A233 & ~A203;
  assign \new_[87014]_  = \new_[87013]_  & \new_[87010]_ ;
  assign \new_[87015]_  = \new_[87014]_  & \new_[87007]_ ;
  assign \new_[87018]_  = ~A236 & ~A235;
  assign \new_[87021]_  = ~A268 & ~A266;
  assign \new_[87022]_  = \new_[87021]_  & \new_[87018]_ ;
  assign \new_[87025]_  = A298 & ~A269;
  assign \new_[87029]_  = A301 & A300;
  assign \new_[87030]_  = ~A299 & \new_[87029]_ ;
  assign \new_[87031]_  = \new_[87030]_  & \new_[87025]_ ;
  assign \new_[87032]_  = \new_[87031]_  & \new_[87022]_ ;
  assign \new_[87035]_  = A169 & ~A170;
  assign \new_[87038]_  = A166 & A167;
  assign \new_[87039]_  = \new_[87038]_  & \new_[87035]_ ;
  assign \new_[87042]_  = ~A202 & ~A200;
  assign \new_[87045]_  = ~A233 & ~A203;
  assign \new_[87046]_  = \new_[87045]_  & \new_[87042]_ ;
  assign \new_[87047]_  = \new_[87046]_  & \new_[87039]_ ;
  assign \new_[87050]_  = ~A236 & ~A235;
  assign \new_[87053]_  = ~A268 & ~A266;
  assign \new_[87054]_  = \new_[87053]_  & \new_[87050]_ ;
  assign \new_[87057]_  = A298 & ~A269;
  assign \new_[87061]_  = A302 & A300;
  assign \new_[87062]_  = ~A299 & \new_[87061]_ ;
  assign \new_[87063]_  = \new_[87062]_  & \new_[87057]_ ;
  assign \new_[87064]_  = \new_[87063]_  & \new_[87054]_ ;
  assign \new_[87067]_  = A169 & ~A170;
  assign \new_[87070]_  = ~A166 & ~A167;
  assign \new_[87071]_  = \new_[87070]_  & \new_[87067]_ ;
  assign \new_[87074]_  = ~A202 & ~A200;
  assign \new_[87077]_  = ~A233 & ~A203;
  assign \new_[87078]_  = \new_[87077]_  & \new_[87074]_ ;
  assign \new_[87079]_  = \new_[87078]_  & \new_[87071]_ ;
  assign \new_[87082]_  = ~A236 & ~A235;
  assign \new_[87085]_  = ~A268 & ~A266;
  assign \new_[87086]_  = \new_[87085]_  & \new_[87082]_ ;
  assign \new_[87089]_  = A298 & ~A269;
  assign \new_[87093]_  = A301 & A300;
  assign \new_[87094]_  = ~A299 & \new_[87093]_ ;
  assign \new_[87095]_  = \new_[87094]_  & \new_[87089]_ ;
  assign \new_[87096]_  = \new_[87095]_  & \new_[87086]_ ;
  assign \new_[87099]_  = A169 & ~A170;
  assign \new_[87102]_  = ~A166 & ~A167;
  assign \new_[87103]_  = \new_[87102]_  & \new_[87099]_ ;
  assign \new_[87106]_  = ~A202 & ~A200;
  assign \new_[87109]_  = ~A233 & ~A203;
  assign \new_[87110]_  = \new_[87109]_  & \new_[87106]_ ;
  assign \new_[87111]_  = \new_[87110]_  & \new_[87103]_ ;
  assign \new_[87114]_  = ~A236 & ~A235;
  assign \new_[87117]_  = ~A268 & ~A266;
  assign \new_[87118]_  = \new_[87117]_  & \new_[87114]_ ;
  assign \new_[87121]_  = A298 & ~A269;
  assign \new_[87125]_  = A302 & A300;
  assign \new_[87126]_  = ~A299 & \new_[87125]_ ;
  assign \new_[87127]_  = \new_[87126]_  & \new_[87121]_ ;
  assign \new_[87128]_  = \new_[87127]_  & \new_[87118]_ ;
  assign \new_[87131]_  = ~A167 & ~A169;
  assign \new_[87134]_  = A199 & ~A166;
  assign \new_[87135]_  = \new_[87134]_  & \new_[87131]_ ;
  assign \new_[87138]_  = A201 & ~A200;
  assign \new_[87141]_  = ~A233 & A202;
  assign \new_[87142]_  = \new_[87141]_  & \new_[87138]_ ;
  assign \new_[87143]_  = \new_[87142]_  & \new_[87135]_ ;
  assign \new_[87146]_  = ~A236 & ~A235;
  assign \new_[87149]_  = ~A268 & ~A266;
  assign \new_[87150]_  = \new_[87149]_  & \new_[87146]_ ;
  assign \new_[87153]_  = A298 & ~A269;
  assign \new_[87157]_  = A301 & A300;
  assign \new_[87158]_  = ~A299 & \new_[87157]_ ;
  assign \new_[87159]_  = \new_[87158]_  & \new_[87153]_ ;
  assign \new_[87160]_  = \new_[87159]_  & \new_[87150]_ ;
  assign \new_[87163]_  = ~A167 & ~A169;
  assign \new_[87166]_  = A199 & ~A166;
  assign \new_[87167]_  = \new_[87166]_  & \new_[87163]_ ;
  assign \new_[87170]_  = A201 & ~A200;
  assign \new_[87173]_  = ~A233 & A202;
  assign \new_[87174]_  = \new_[87173]_  & \new_[87170]_ ;
  assign \new_[87175]_  = \new_[87174]_  & \new_[87167]_ ;
  assign \new_[87178]_  = ~A236 & ~A235;
  assign \new_[87181]_  = ~A268 & ~A266;
  assign \new_[87182]_  = \new_[87181]_  & \new_[87178]_ ;
  assign \new_[87185]_  = A298 & ~A269;
  assign \new_[87189]_  = A302 & A300;
  assign \new_[87190]_  = ~A299 & \new_[87189]_ ;
  assign \new_[87191]_  = \new_[87190]_  & \new_[87185]_ ;
  assign \new_[87192]_  = \new_[87191]_  & \new_[87182]_ ;
  assign \new_[87195]_  = ~A167 & ~A169;
  assign \new_[87198]_  = A199 & ~A166;
  assign \new_[87199]_  = \new_[87198]_  & \new_[87195]_ ;
  assign \new_[87202]_  = A201 & ~A200;
  assign \new_[87205]_  = ~A233 & A203;
  assign \new_[87206]_  = \new_[87205]_  & \new_[87202]_ ;
  assign \new_[87207]_  = \new_[87206]_  & \new_[87199]_ ;
  assign \new_[87210]_  = ~A236 & ~A235;
  assign \new_[87213]_  = ~A268 & ~A266;
  assign \new_[87214]_  = \new_[87213]_  & \new_[87210]_ ;
  assign \new_[87217]_  = A298 & ~A269;
  assign \new_[87221]_  = A301 & A300;
  assign \new_[87222]_  = ~A299 & \new_[87221]_ ;
  assign \new_[87223]_  = \new_[87222]_  & \new_[87217]_ ;
  assign \new_[87224]_  = \new_[87223]_  & \new_[87214]_ ;
  assign \new_[87227]_  = ~A167 & ~A169;
  assign \new_[87230]_  = A199 & ~A166;
  assign \new_[87231]_  = \new_[87230]_  & \new_[87227]_ ;
  assign \new_[87234]_  = A201 & ~A200;
  assign \new_[87237]_  = ~A233 & A203;
  assign \new_[87238]_  = \new_[87237]_  & \new_[87234]_ ;
  assign \new_[87239]_  = \new_[87238]_  & \new_[87231]_ ;
  assign \new_[87242]_  = ~A236 & ~A235;
  assign \new_[87245]_  = ~A268 & ~A266;
  assign \new_[87246]_  = \new_[87245]_  & \new_[87242]_ ;
  assign \new_[87249]_  = A298 & ~A269;
  assign \new_[87253]_  = A302 & A300;
  assign \new_[87254]_  = ~A299 & \new_[87253]_ ;
  assign \new_[87255]_  = \new_[87254]_  & \new_[87249]_ ;
  assign \new_[87256]_  = \new_[87255]_  & \new_[87246]_ ;
  assign \new_[87259]_  = ~A168 & ~A169;
  assign \new_[87262]_  = A166 & A167;
  assign \new_[87263]_  = \new_[87262]_  & \new_[87259]_ ;
  assign \new_[87266]_  = ~A200 & A199;
  assign \new_[87269]_  = A202 & A201;
  assign \new_[87270]_  = \new_[87269]_  & \new_[87266]_ ;
  assign \new_[87271]_  = \new_[87270]_  & \new_[87263]_ ;
  assign \new_[87274]_  = A233 & A232;
  assign \new_[87277]_  = ~A268 & A265;
  assign \new_[87278]_  = \new_[87277]_  & \new_[87274]_ ;
  assign \new_[87281]_  = A298 & ~A269;
  assign \new_[87285]_  = A301 & A300;
  assign \new_[87286]_  = ~A299 & \new_[87285]_ ;
  assign \new_[87287]_  = \new_[87286]_  & \new_[87281]_ ;
  assign \new_[87288]_  = \new_[87287]_  & \new_[87278]_ ;
  assign \new_[87291]_  = ~A168 & ~A169;
  assign \new_[87294]_  = A166 & A167;
  assign \new_[87295]_  = \new_[87294]_  & \new_[87291]_ ;
  assign \new_[87298]_  = ~A200 & A199;
  assign \new_[87301]_  = A202 & A201;
  assign \new_[87302]_  = \new_[87301]_  & \new_[87298]_ ;
  assign \new_[87303]_  = \new_[87302]_  & \new_[87295]_ ;
  assign \new_[87306]_  = A233 & A232;
  assign \new_[87309]_  = ~A268 & A265;
  assign \new_[87310]_  = \new_[87309]_  & \new_[87306]_ ;
  assign \new_[87313]_  = A298 & ~A269;
  assign \new_[87317]_  = A302 & A300;
  assign \new_[87318]_  = ~A299 & \new_[87317]_ ;
  assign \new_[87319]_  = \new_[87318]_  & \new_[87313]_ ;
  assign \new_[87320]_  = \new_[87319]_  & \new_[87310]_ ;
  assign \new_[87323]_  = ~A168 & ~A169;
  assign \new_[87326]_  = A166 & A167;
  assign \new_[87327]_  = \new_[87326]_  & \new_[87323]_ ;
  assign \new_[87330]_  = ~A200 & A199;
  assign \new_[87333]_  = A202 & A201;
  assign \new_[87334]_  = \new_[87333]_  & \new_[87330]_ ;
  assign \new_[87335]_  = \new_[87334]_  & \new_[87327]_ ;
  assign \new_[87338]_  = ~A235 & ~A233;
  assign \new_[87341]_  = A265 & ~A236;
  assign \new_[87342]_  = \new_[87341]_  & \new_[87338]_ ;
  assign \new_[87345]_  = A298 & A266;
  assign \new_[87349]_  = A301 & A300;
  assign \new_[87350]_  = ~A299 & \new_[87349]_ ;
  assign \new_[87351]_  = \new_[87350]_  & \new_[87345]_ ;
  assign \new_[87352]_  = \new_[87351]_  & \new_[87342]_ ;
  assign \new_[87355]_  = ~A168 & ~A169;
  assign \new_[87358]_  = A166 & A167;
  assign \new_[87359]_  = \new_[87358]_  & \new_[87355]_ ;
  assign \new_[87362]_  = ~A200 & A199;
  assign \new_[87365]_  = A202 & A201;
  assign \new_[87366]_  = \new_[87365]_  & \new_[87362]_ ;
  assign \new_[87367]_  = \new_[87366]_  & \new_[87359]_ ;
  assign \new_[87370]_  = ~A235 & ~A233;
  assign \new_[87373]_  = A265 & ~A236;
  assign \new_[87374]_  = \new_[87373]_  & \new_[87370]_ ;
  assign \new_[87377]_  = A298 & A266;
  assign \new_[87381]_  = A302 & A300;
  assign \new_[87382]_  = ~A299 & \new_[87381]_ ;
  assign \new_[87383]_  = \new_[87382]_  & \new_[87377]_ ;
  assign \new_[87384]_  = \new_[87383]_  & \new_[87374]_ ;
  assign \new_[87387]_  = ~A168 & ~A169;
  assign \new_[87390]_  = A166 & A167;
  assign \new_[87391]_  = \new_[87390]_  & \new_[87387]_ ;
  assign \new_[87394]_  = ~A200 & A199;
  assign \new_[87397]_  = A202 & A201;
  assign \new_[87398]_  = \new_[87397]_  & \new_[87394]_ ;
  assign \new_[87399]_  = \new_[87398]_  & \new_[87391]_ ;
  assign \new_[87402]_  = ~A235 & ~A233;
  assign \new_[87405]_  = ~A266 & ~A236;
  assign \new_[87406]_  = \new_[87405]_  & \new_[87402]_ ;
  assign \new_[87409]_  = A298 & ~A267;
  assign \new_[87413]_  = A301 & A300;
  assign \new_[87414]_  = ~A299 & \new_[87413]_ ;
  assign \new_[87415]_  = \new_[87414]_  & \new_[87409]_ ;
  assign \new_[87416]_  = \new_[87415]_  & \new_[87406]_ ;
  assign \new_[87419]_  = ~A168 & ~A169;
  assign \new_[87422]_  = A166 & A167;
  assign \new_[87423]_  = \new_[87422]_  & \new_[87419]_ ;
  assign \new_[87426]_  = ~A200 & A199;
  assign \new_[87429]_  = A202 & A201;
  assign \new_[87430]_  = \new_[87429]_  & \new_[87426]_ ;
  assign \new_[87431]_  = \new_[87430]_  & \new_[87423]_ ;
  assign \new_[87434]_  = ~A235 & ~A233;
  assign \new_[87437]_  = ~A266 & ~A236;
  assign \new_[87438]_  = \new_[87437]_  & \new_[87434]_ ;
  assign \new_[87441]_  = A298 & ~A267;
  assign \new_[87445]_  = A302 & A300;
  assign \new_[87446]_  = ~A299 & \new_[87445]_ ;
  assign \new_[87447]_  = \new_[87446]_  & \new_[87441]_ ;
  assign \new_[87448]_  = \new_[87447]_  & \new_[87438]_ ;
  assign \new_[87451]_  = ~A168 & ~A169;
  assign \new_[87454]_  = A166 & A167;
  assign \new_[87455]_  = \new_[87454]_  & \new_[87451]_ ;
  assign \new_[87458]_  = ~A200 & A199;
  assign \new_[87461]_  = A202 & A201;
  assign \new_[87462]_  = \new_[87461]_  & \new_[87458]_ ;
  assign \new_[87463]_  = \new_[87462]_  & \new_[87455]_ ;
  assign \new_[87466]_  = ~A235 & ~A233;
  assign \new_[87469]_  = ~A265 & ~A236;
  assign \new_[87470]_  = \new_[87469]_  & \new_[87466]_ ;
  assign \new_[87473]_  = A298 & ~A266;
  assign \new_[87477]_  = A301 & A300;
  assign \new_[87478]_  = ~A299 & \new_[87477]_ ;
  assign \new_[87479]_  = \new_[87478]_  & \new_[87473]_ ;
  assign \new_[87480]_  = \new_[87479]_  & \new_[87470]_ ;
  assign \new_[87483]_  = ~A168 & ~A169;
  assign \new_[87486]_  = A166 & A167;
  assign \new_[87487]_  = \new_[87486]_  & \new_[87483]_ ;
  assign \new_[87490]_  = ~A200 & A199;
  assign \new_[87493]_  = A202 & A201;
  assign \new_[87494]_  = \new_[87493]_  & \new_[87490]_ ;
  assign \new_[87495]_  = \new_[87494]_  & \new_[87487]_ ;
  assign \new_[87498]_  = ~A235 & ~A233;
  assign \new_[87501]_  = ~A265 & ~A236;
  assign \new_[87502]_  = \new_[87501]_  & \new_[87498]_ ;
  assign \new_[87505]_  = A298 & ~A266;
  assign \new_[87509]_  = A302 & A300;
  assign \new_[87510]_  = ~A299 & \new_[87509]_ ;
  assign \new_[87511]_  = \new_[87510]_  & \new_[87505]_ ;
  assign \new_[87512]_  = \new_[87511]_  & \new_[87502]_ ;
  assign \new_[87515]_  = ~A168 & ~A169;
  assign \new_[87518]_  = A166 & A167;
  assign \new_[87519]_  = \new_[87518]_  & \new_[87515]_ ;
  assign \new_[87522]_  = ~A200 & A199;
  assign \new_[87525]_  = A202 & A201;
  assign \new_[87526]_  = \new_[87525]_  & \new_[87522]_ ;
  assign \new_[87527]_  = \new_[87526]_  & \new_[87519]_ ;
  assign \new_[87530]_  = ~A234 & ~A233;
  assign \new_[87533]_  = ~A268 & ~A266;
  assign \new_[87534]_  = \new_[87533]_  & \new_[87530]_ ;
  assign \new_[87537]_  = A298 & ~A269;
  assign \new_[87541]_  = A301 & A300;
  assign \new_[87542]_  = ~A299 & \new_[87541]_ ;
  assign \new_[87543]_  = \new_[87542]_  & \new_[87537]_ ;
  assign \new_[87544]_  = \new_[87543]_  & \new_[87534]_ ;
  assign \new_[87547]_  = ~A168 & ~A169;
  assign \new_[87550]_  = A166 & A167;
  assign \new_[87551]_  = \new_[87550]_  & \new_[87547]_ ;
  assign \new_[87554]_  = ~A200 & A199;
  assign \new_[87557]_  = A202 & A201;
  assign \new_[87558]_  = \new_[87557]_  & \new_[87554]_ ;
  assign \new_[87559]_  = \new_[87558]_  & \new_[87551]_ ;
  assign \new_[87562]_  = ~A234 & ~A233;
  assign \new_[87565]_  = ~A268 & ~A266;
  assign \new_[87566]_  = \new_[87565]_  & \new_[87562]_ ;
  assign \new_[87569]_  = A298 & ~A269;
  assign \new_[87573]_  = A302 & A300;
  assign \new_[87574]_  = ~A299 & \new_[87573]_ ;
  assign \new_[87575]_  = \new_[87574]_  & \new_[87569]_ ;
  assign \new_[87576]_  = \new_[87575]_  & \new_[87566]_ ;
  assign \new_[87579]_  = ~A168 & ~A169;
  assign \new_[87582]_  = A166 & A167;
  assign \new_[87583]_  = \new_[87582]_  & \new_[87579]_ ;
  assign \new_[87586]_  = ~A200 & A199;
  assign \new_[87589]_  = A202 & A201;
  assign \new_[87590]_  = \new_[87589]_  & \new_[87586]_ ;
  assign \new_[87591]_  = \new_[87590]_  & \new_[87583]_ ;
  assign \new_[87594]_  = ~A233 & ~A232;
  assign \new_[87597]_  = ~A268 & ~A266;
  assign \new_[87598]_  = \new_[87597]_  & \new_[87594]_ ;
  assign \new_[87601]_  = A298 & ~A269;
  assign \new_[87605]_  = A301 & A300;
  assign \new_[87606]_  = ~A299 & \new_[87605]_ ;
  assign \new_[87607]_  = \new_[87606]_  & \new_[87601]_ ;
  assign \new_[87608]_  = \new_[87607]_  & \new_[87598]_ ;
  assign \new_[87611]_  = ~A168 & ~A169;
  assign \new_[87614]_  = A166 & A167;
  assign \new_[87615]_  = \new_[87614]_  & \new_[87611]_ ;
  assign \new_[87618]_  = ~A200 & A199;
  assign \new_[87621]_  = A202 & A201;
  assign \new_[87622]_  = \new_[87621]_  & \new_[87618]_ ;
  assign \new_[87623]_  = \new_[87622]_  & \new_[87615]_ ;
  assign \new_[87626]_  = ~A233 & ~A232;
  assign \new_[87629]_  = ~A268 & ~A266;
  assign \new_[87630]_  = \new_[87629]_  & \new_[87626]_ ;
  assign \new_[87633]_  = A298 & ~A269;
  assign \new_[87637]_  = A302 & A300;
  assign \new_[87638]_  = ~A299 & \new_[87637]_ ;
  assign \new_[87639]_  = \new_[87638]_  & \new_[87633]_ ;
  assign \new_[87640]_  = \new_[87639]_  & \new_[87630]_ ;
  assign \new_[87643]_  = ~A168 & ~A169;
  assign \new_[87646]_  = A166 & A167;
  assign \new_[87647]_  = \new_[87646]_  & \new_[87643]_ ;
  assign \new_[87650]_  = ~A200 & A199;
  assign \new_[87653]_  = A203 & A201;
  assign \new_[87654]_  = \new_[87653]_  & \new_[87650]_ ;
  assign \new_[87655]_  = \new_[87654]_  & \new_[87647]_ ;
  assign \new_[87658]_  = A233 & A232;
  assign \new_[87661]_  = ~A268 & A265;
  assign \new_[87662]_  = \new_[87661]_  & \new_[87658]_ ;
  assign \new_[87665]_  = A298 & ~A269;
  assign \new_[87669]_  = A301 & A300;
  assign \new_[87670]_  = ~A299 & \new_[87669]_ ;
  assign \new_[87671]_  = \new_[87670]_  & \new_[87665]_ ;
  assign \new_[87672]_  = \new_[87671]_  & \new_[87662]_ ;
  assign \new_[87675]_  = ~A168 & ~A169;
  assign \new_[87678]_  = A166 & A167;
  assign \new_[87679]_  = \new_[87678]_  & \new_[87675]_ ;
  assign \new_[87682]_  = ~A200 & A199;
  assign \new_[87685]_  = A203 & A201;
  assign \new_[87686]_  = \new_[87685]_  & \new_[87682]_ ;
  assign \new_[87687]_  = \new_[87686]_  & \new_[87679]_ ;
  assign \new_[87690]_  = A233 & A232;
  assign \new_[87693]_  = ~A268 & A265;
  assign \new_[87694]_  = \new_[87693]_  & \new_[87690]_ ;
  assign \new_[87697]_  = A298 & ~A269;
  assign \new_[87701]_  = A302 & A300;
  assign \new_[87702]_  = ~A299 & \new_[87701]_ ;
  assign \new_[87703]_  = \new_[87702]_  & \new_[87697]_ ;
  assign \new_[87704]_  = \new_[87703]_  & \new_[87694]_ ;
  assign \new_[87707]_  = ~A168 & ~A169;
  assign \new_[87710]_  = A166 & A167;
  assign \new_[87711]_  = \new_[87710]_  & \new_[87707]_ ;
  assign \new_[87714]_  = ~A200 & A199;
  assign \new_[87717]_  = A203 & A201;
  assign \new_[87718]_  = \new_[87717]_  & \new_[87714]_ ;
  assign \new_[87719]_  = \new_[87718]_  & \new_[87711]_ ;
  assign \new_[87722]_  = ~A235 & ~A233;
  assign \new_[87725]_  = A265 & ~A236;
  assign \new_[87726]_  = \new_[87725]_  & \new_[87722]_ ;
  assign \new_[87729]_  = A298 & A266;
  assign \new_[87733]_  = A301 & A300;
  assign \new_[87734]_  = ~A299 & \new_[87733]_ ;
  assign \new_[87735]_  = \new_[87734]_  & \new_[87729]_ ;
  assign \new_[87736]_  = \new_[87735]_  & \new_[87726]_ ;
  assign \new_[87739]_  = ~A168 & ~A169;
  assign \new_[87742]_  = A166 & A167;
  assign \new_[87743]_  = \new_[87742]_  & \new_[87739]_ ;
  assign \new_[87746]_  = ~A200 & A199;
  assign \new_[87749]_  = A203 & A201;
  assign \new_[87750]_  = \new_[87749]_  & \new_[87746]_ ;
  assign \new_[87751]_  = \new_[87750]_  & \new_[87743]_ ;
  assign \new_[87754]_  = ~A235 & ~A233;
  assign \new_[87757]_  = A265 & ~A236;
  assign \new_[87758]_  = \new_[87757]_  & \new_[87754]_ ;
  assign \new_[87761]_  = A298 & A266;
  assign \new_[87765]_  = A302 & A300;
  assign \new_[87766]_  = ~A299 & \new_[87765]_ ;
  assign \new_[87767]_  = \new_[87766]_  & \new_[87761]_ ;
  assign \new_[87768]_  = \new_[87767]_  & \new_[87758]_ ;
  assign \new_[87771]_  = ~A168 & ~A169;
  assign \new_[87774]_  = A166 & A167;
  assign \new_[87775]_  = \new_[87774]_  & \new_[87771]_ ;
  assign \new_[87778]_  = ~A200 & A199;
  assign \new_[87781]_  = A203 & A201;
  assign \new_[87782]_  = \new_[87781]_  & \new_[87778]_ ;
  assign \new_[87783]_  = \new_[87782]_  & \new_[87775]_ ;
  assign \new_[87786]_  = ~A235 & ~A233;
  assign \new_[87789]_  = ~A266 & ~A236;
  assign \new_[87790]_  = \new_[87789]_  & \new_[87786]_ ;
  assign \new_[87793]_  = A298 & ~A267;
  assign \new_[87797]_  = A301 & A300;
  assign \new_[87798]_  = ~A299 & \new_[87797]_ ;
  assign \new_[87799]_  = \new_[87798]_  & \new_[87793]_ ;
  assign \new_[87800]_  = \new_[87799]_  & \new_[87790]_ ;
  assign \new_[87803]_  = ~A168 & ~A169;
  assign \new_[87806]_  = A166 & A167;
  assign \new_[87807]_  = \new_[87806]_  & \new_[87803]_ ;
  assign \new_[87810]_  = ~A200 & A199;
  assign \new_[87813]_  = A203 & A201;
  assign \new_[87814]_  = \new_[87813]_  & \new_[87810]_ ;
  assign \new_[87815]_  = \new_[87814]_  & \new_[87807]_ ;
  assign \new_[87818]_  = ~A235 & ~A233;
  assign \new_[87821]_  = ~A266 & ~A236;
  assign \new_[87822]_  = \new_[87821]_  & \new_[87818]_ ;
  assign \new_[87825]_  = A298 & ~A267;
  assign \new_[87829]_  = A302 & A300;
  assign \new_[87830]_  = ~A299 & \new_[87829]_ ;
  assign \new_[87831]_  = \new_[87830]_  & \new_[87825]_ ;
  assign \new_[87832]_  = \new_[87831]_  & \new_[87822]_ ;
  assign \new_[87835]_  = ~A168 & ~A169;
  assign \new_[87838]_  = A166 & A167;
  assign \new_[87839]_  = \new_[87838]_  & \new_[87835]_ ;
  assign \new_[87842]_  = ~A200 & A199;
  assign \new_[87845]_  = A203 & A201;
  assign \new_[87846]_  = \new_[87845]_  & \new_[87842]_ ;
  assign \new_[87847]_  = \new_[87846]_  & \new_[87839]_ ;
  assign \new_[87850]_  = ~A235 & ~A233;
  assign \new_[87853]_  = ~A265 & ~A236;
  assign \new_[87854]_  = \new_[87853]_  & \new_[87850]_ ;
  assign \new_[87857]_  = A298 & ~A266;
  assign \new_[87861]_  = A301 & A300;
  assign \new_[87862]_  = ~A299 & \new_[87861]_ ;
  assign \new_[87863]_  = \new_[87862]_  & \new_[87857]_ ;
  assign \new_[87864]_  = \new_[87863]_  & \new_[87854]_ ;
  assign \new_[87867]_  = ~A168 & ~A169;
  assign \new_[87870]_  = A166 & A167;
  assign \new_[87871]_  = \new_[87870]_  & \new_[87867]_ ;
  assign \new_[87874]_  = ~A200 & A199;
  assign \new_[87877]_  = A203 & A201;
  assign \new_[87878]_  = \new_[87877]_  & \new_[87874]_ ;
  assign \new_[87879]_  = \new_[87878]_  & \new_[87871]_ ;
  assign \new_[87882]_  = ~A235 & ~A233;
  assign \new_[87885]_  = ~A265 & ~A236;
  assign \new_[87886]_  = \new_[87885]_  & \new_[87882]_ ;
  assign \new_[87889]_  = A298 & ~A266;
  assign \new_[87893]_  = A302 & A300;
  assign \new_[87894]_  = ~A299 & \new_[87893]_ ;
  assign \new_[87895]_  = \new_[87894]_  & \new_[87889]_ ;
  assign \new_[87896]_  = \new_[87895]_  & \new_[87886]_ ;
  assign \new_[87899]_  = ~A168 & ~A169;
  assign \new_[87902]_  = A166 & A167;
  assign \new_[87903]_  = \new_[87902]_  & \new_[87899]_ ;
  assign \new_[87906]_  = ~A200 & A199;
  assign \new_[87909]_  = A203 & A201;
  assign \new_[87910]_  = \new_[87909]_  & \new_[87906]_ ;
  assign \new_[87911]_  = \new_[87910]_  & \new_[87903]_ ;
  assign \new_[87914]_  = ~A234 & ~A233;
  assign \new_[87917]_  = ~A268 & ~A266;
  assign \new_[87918]_  = \new_[87917]_  & \new_[87914]_ ;
  assign \new_[87921]_  = A298 & ~A269;
  assign \new_[87925]_  = A301 & A300;
  assign \new_[87926]_  = ~A299 & \new_[87925]_ ;
  assign \new_[87927]_  = \new_[87926]_  & \new_[87921]_ ;
  assign \new_[87928]_  = \new_[87927]_  & \new_[87918]_ ;
  assign \new_[87931]_  = ~A168 & ~A169;
  assign \new_[87934]_  = A166 & A167;
  assign \new_[87935]_  = \new_[87934]_  & \new_[87931]_ ;
  assign \new_[87938]_  = ~A200 & A199;
  assign \new_[87941]_  = A203 & A201;
  assign \new_[87942]_  = \new_[87941]_  & \new_[87938]_ ;
  assign \new_[87943]_  = \new_[87942]_  & \new_[87935]_ ;
  assign \new_[87946]_  = ~A234 & ~A233;
  assign \new_[87949]_  = ~A268 & ~A266;
  assign \new_[87950]_  = \new_[87949]_  & \new_[87946]_ ;
  assign \new_[87953]_  = A298 & ~A269;
  assign \new_[87957]_  = A302 & A300;
  assign \new_[87958]_  = ~A299 & \new_[87957]_ ;
  assign \new_[87959]_  = \new_[87958]_  & \new_[87953]_ ;
  assign \new_[87960]_  = \new_[87959]_  & \new_[87950]_ ;
  assign \new_[87963]_  = ~A168 & ~A169;
  assign \new_[87966]_  = A166 & A167;
  assign \new_[87967]_  = \new_[87966]_  & \new_[87963]_ ;
  assign \new_[87970]_  = ~A200 & A199;
  assign \new_[87973]_  = A203 & A201;
  assign \new_[87974]_  = \new_[87973]_  & \new_[87970]_ ;
  assign \new_[87975]_  = \new_[87974]_  & \new_[87967]_ ;
  assign \new_[87978]_  = ~A233 & ~A232;
  assign \new_[87981]_  = ~A268 & ~A266;
  assign \new_[87982]_  = \new_[87981]_  & \new_[87978]_ ;
  assign \new_[87985]_  = A298 & ~A269;
  assign \new_[87989]_  = A301 & A300;
  assign \new_[87990]_  = ~A299 & \new_[87989]_ ;
  assign \new_[87991]_  = \new_[87990]_  & \new_[87985]_ ;
  assign \new_[87992]_  = \new_[87991]_  & \new_[87982]_ ;
  assign \new_[87995]_  = ~A168 & ~A169;
  assign \new_[87998]_  = A166 & A167;
  assign \new_[87999]_  = \new_[87998]_  & \new_[87995]_ ;
  assign \new_[88002]_  = ~A200 & A199;
  assign \new_[88005]_  = A203 & A201;
  assign \new_[88006]_  = \new_[88005]_  & \new_[88002]_ ;
  assign \new_[88007]_  = \new_[88006]_  & \new_[87999]_ ;
  assign \new_[88010]_  = ~A233 & ~A232;
  assign \new_[88013]_  = ~A268 & ~A266;
  assign \new_[88014]_  = \new_[88013]_  & \new_[88010]_ ;
  assign \new_[88017]_  = A298 & ~A269;
  assign \new_[88021]_  = A302 & A300;
  assign \new_[88022]_  = ~A299 & \new_[88021]_ ;
  assign \new_[88023]_  = \new_[88022]_  & \new_[88017]_ ;
  assign \new_[88024]_  = \new_[88023]_  & \new_[88014]_ ;
  assign \new_[88027]_  = ~A169 & A170;
  assign \new_[88030]_  = ~A166 & A167;
  assign \new_[88031]_  = \new_[88030]_  & \new_[88027]_ ;
  assign \new_[88034]_  = ~A202 & ~A200;
  assign \new_[88037]_  = ~A233 & ~A203;
  assign \new_[88038]_  = \new_[88037]_  & \new_[88034]_ ;
  assign \new_[88039]_  = \new_[88038]_  & \new_[88031]_ ;
  assign \new_[88042]_  = ~A236 & ~A235;
  assign \new_[88045]_  = ~A268 & ~A266;
  assign \new_[88046]_  = \new_[88045]_  & \new_[88042]_ ;
  assign \new_[88049]_  = A298 & ~A269;
  assign \new_[88053]_  = A301 & A300;
  assign \new_[88054]_  = ~A299 & \new_[88053]_ ;
  assign \new_[88055]_  = \new_[88054]_  & \new_[88049]_ ;
  assign \new_[88056]_  = \new_[88055]_  & \new_[88046]_ ;
  assign \new_[88059]_  = ~A169 & A170;
  assign \new_[88062]_  = ~A166 & A167;
  assign \new_[88063]_  = \new_[88062]_  & \new_[88059]_ ;
  assign \new_[88066]_  = ~A202 & ~A200;
  assign \new_[88069]_  = ~A233 & ~A203;
  assign \new_[88070]_  = \new_[88069]_  & \new_[88066]_ ;
  assign \new_[88071]_  = \new_[88070]_  & \new_[88063]_ ;
  assign \new_[88074]_  = ~A236 & ~A235;
  assign \new_[88077]_  = ~A268 & ~A266;
  assign \new_[88078]_  = \new_[88077]_  & \new_[88074]_ ;
  assign \new_[88081]_  = A298 & ~A269;
  assign \new_[88085]_  = A302 & A300;
  assign \new_[88086]_  = ~A299 & \new_[88085]_ ;
  assign \new_[88087]_  = \new_[88086]_  & \new_[88081]_ ;
  assign \new_[88088]_  = \new_[88087]_  & \new_[88078]_ ;
  assign \new_[88091]_  = ~A169 & A170;
  assign \new_[88094]_  = A166 & ~A167;
  assign \new_[88095]_  = \new_[88094]_  & \new_[88091]_ ;
  assign \new_[88098]_  = ~A202 & ~A200;
  assign \new_[88101]_  = ~A233 & ~A203;
  assign \new_[88102]_  = \new_[88101]_  & \new_[88098]_ ;
  assign \new_[88103]_  = \new_[88102]_  & \new_[88095]_ ;
  assign \new_[88106]_  = ~A236 & ~A235;
  assign \new_[88109]_  = ~A268 & ~A266;
  assign \new_[88110]_  = \new_[88109]_  & \new_[88106]_ ;
  assign \new_[88113]_  = A298 & ~A269;
  assign \new_[88117]_  = A301 & A300;
  assign \new_[88118]_  = ~A299 & \new_[88117]_ ;
  assign \new_[88119]_  = \new_[88118]_  & \new_[88113]_ ;
  assign \new_[88120]_  = \new_[88119]_  & \new_[88110]_ ;
  assign \new_[88123]_  = ~A169 & A170;
  assign \new_[88126]_  = A166 & ~A167;
  assign \new_[88127]_  = \new_[88126]_  & \new_[88123]_ ;
  assign \new_[88130]_  = ~A202 & ~A200;
  assign \new_[88133]_  = ~A233 & ~A203;
  assign \new_[88134]_  = \new_[88133]_  & \new_[88130]_ ;
  assign \new_[88135]_  = \new_[88134]_  & \new_[88127]_ ;
  assign \new_[88138]_  = ~A236 & ~A235;
  assign \new_[88141]_  = ~A268 & ~A266;
  assign \new_[88142]_  = \new_[88141]_  & \new_[88138]_ ;
  assign \new_[88145]_  = A298 & ~A269;
  assign \new_[88149]_  = A302 & A300;
  assign \new_[88150]_  = ~A299 & \new_[88149]_ ;
  assign \new_[88151]_  = \new_[88150]_  & \new_[88145]_ ;
  assign \new_[88152]_  = \new_[88151]_  & \new_[88142]_ ;
  assign \new_[88155]_  = ~A169 & ~A170;
  assign \new_[88158]_  = A199 & ~A168;
  assign \new_[88159]_  = \new_[88158]_  & \new_[88155]_ ;
  assign \new_[88162]_  = A201 & ~A200;
  assign \new_[88165]_  = ~A233 & A202;
  assign \new_[88166]_  = \new_[88165]_  & \new_[88162]_ ;
  assign \new_[88167]_  = \new_[88166]_  & \new_[88159]_ ;
  assign \new_[88170]_  = ~A236 & ~A235;
  assign \new_[88173]_  = ~A268 & ~A266;
  assign \new_[88174]_  = \new_[88173]_  & \new_[88170]_ ;
  assign \new_[88177]_  = A298 & ~A269;
  assign \new_[88181]_  = A301 & A300;
  assign \new_[88182]_  = ~A299 & \new_[88181]_ ;
  assign \new_[88183]_  = \new_[88182]_  & \new_[88177]_ ;
  assign \new_[88184]_  = \new_[88183]_  & \new_[88174]_ ;
  assign \new_[88187]_  = ~A169 & ~A170;
  assign \new_[88190]_  = A199 & ~A168;
  assign \new_[88191]_  = \new_[88190]_  & \new_[88187]_ ;
  assign \new_[88194]_  = A201 & ~A200;
  assign \new_[88197]_  = ~A233 & A202;
  assign \new_[88198]_  = \new_[88197]_  & \new_[88194]_ ;
  assign \new_[88199]_  = \new_[88198]_  & \new_[88191]_ ;
  assign \new_[88202]_  = ~A236 & ~A235;
  assign \new_[88205]_  = ~A268 & ~A266;
  assign \new_[88206]_  = \new_[88205]_  & \new_[88202]_ ;
  assign \new_[88209]_  = A298 & ~A269;
  assign \new_[88213]_  = A302 & A300;
  assign \new_[88214]_  = ~A299 & \new_[88213]_ ;
  assign \new_[88215]_  = \new_[88214]_  & \new_[88209]_ ;
  assign \new_[88216]_  = \new_[88215]_  & \new_[88206]_ ;
  assign \new_[88219]_  = ~A169 & ~A170;
  assign \new_[88222]_  = A199 & ~A168;
  assign \new_[88223]_  = \new_[88222]_  & \new_[88219]_ ;
  assign \new_[88226]_  = A201 & ~A200;
  assign \new_[88229]_  = ~A233 & A203;
  assign \new_[88230]_  = \new_[88229]_  & \new_[88226]_ ;
  assign \new_[88231]_  = \new_[88230]_  & \new_[88223]_ ;
  assign \new_[88234]_  = ~A236 & ~A235;
  assign \new_[88237]_  = ~A268 & ~A266;
  assign \new_[88238]_  = \new_[88237]_  & \new_[88234]_ ;
  assign \new_[88241]_  = A298 & ~A269;
  assign \new_[88245]_  = A301 & A300;
  assign \new_[88246]_  = ~A299 & \new_[88245]_ ;
  assign \new_[88247]_  = \new_[88246]_  & \new_[88241]_ ;
  assign \new_[88248]_  = \new_[88247]_  & \new_[88238]_ ;
  assign \new_[88251]_  = ~A169 & ~A170;
  assign \new_[88254]_  = A199 & ~A168;
  assign \new_[88255]_  = \new_[88254]_  & \new_[88251]_ ;
  assign \new_[88258]_  = A201 & ~A200;
  assign \new_[88261]_  = ~A233 & A203;
  assign \new_[88262]_  = \new_[88261]_  & \new_[88258]_ ;
  assign \new_[88263]_  = \new_[88262]_  & \new_[88255]_ ;
  assign \new_[88266]_  = ~A236 & ~A235;
  assign \new_[88269]_  = ~A268 & ~A266;
  assign \new_[88270]_  = \new_[88269]_  & \new_[88266]_ ;
  assign \new_[88273]_  = A298 & ~A269;
  assign \new_[88277]_  = A302 & A300;
  assign \new_[88278]_  = ~A299 & \new_[88277]_ ;
  assign \new_[88279]_  = \new_[88278]_  & \new_[88273]_ ;
  assign \new_[88280]_  = \new_[88279]_  & \new_[88270]_ ;
  assign \new_[88283]_  = ~A168 & A169;
  assign \new_[88286]_  = ~A166 & A167;
  assign \new_[88287]_  = \new_[88286]_  & \new_[88283]_ ;
  assign \new_[88290]_  = ~A200 & A199;
  assign \new_[88294]_  = ~A233 & A202;
  assign \new_[88295]_  = A201 & \new_[88294]_ ;
  assign \new_[88296]_  = \new_[88295]_  & \new_[88290]_ ;
  assign \new_[88297]_  = \new_[88296]_  & \new_[88287]_ ;
  assign \new_[88300]_  = ~A236 & ~A235;
  assign \new_[88303]_  = ~A268 & ~A266;
  assign \new_[88304]_  = \new_[88303]_  & \new_[88300]_ ;
  assign \new_[88307]_  = A298 & ~A269;
  assign \new_[88311]_  = A301 & A300;
  assign \new_[88312]_  = ~A299 & \new_[88311]_ ;
  assign \new_[88313]_  = \new_[88312]_  & \new_[88307]_ ;
  assign \new_[88314]_  = \new_[88313]_  & \new_[88304]_ ;
  assign \new_[88317]_  = ~A168 & A169;
  assign \new_[88320]_  = ~A166 & A167;
  assign \new_[88321]_  = \new_[88320]_  & \new_[88317]_ ;
  assign \new_[88324]_  = ~A200 & A199;
  assign \new_[88328]_  = ~A233 & A202;
  assign \new_[88329]_  = A201 & \new_[88328]_ ;
  assign \new_[88330]_  = \new_[88329]_  & \new_[88324]_ ;
  assign \new_[88331]_  = \new_[88330]_  & \new_[88321]_ ;
  assign \new_[88334]_  = ~A236 & ~A235;
  assign \new_[88337]_  = ~A268 & ~A266;
  assign \new_[88338]_  = \new_[88337]_  & \new_[88334]_ ;
  assign \new_[88341]_  = A298 & ~A269;
  assign \new_[88345]_  = A302 & A300;
  assign \new_[88346]_  = ~A299 & \new_[88345]_ ;
  assign \new_[88347]_  = \new_[88346]_  & \new_[88341]_ ;
  assign \new_[88348]_  = \new_[88347]_  & \new_[88338]_ ;
  assign \new_[88351]_  = ~A168 & A169;
  assign \new_[88354]_  = ~A166 & A167;
  assign \new_[88355]_  = \new_[88354]_  & \new_[88351]_ ;
  assign \new_[88358]_  = ~A200 & A199;
  assign \new_[88362]_  = ~A233 & A203;
  assign \new_[88363]_  = A201 & \new_[88362]_ ;
  assign \new_[88364]_  = \new_[88363]_  & \new_[88358]_ ;
  assign \new_[88365]_  = \new_[88364]_  & \new_[88355]_ ;
  assign \new_[88368]_  = ~A236 & ~A235;
  assign \new_[88371]_  = ~A268 & ~A266;
  assign \new_[88372]_  = \new_[88371]_  & \new_[88368]_ ;
  assign \new_[88375]_  = A298 & ~A269;
  assign \new_[88379]_  = A301 & A300;
  assign \new_[88380]_  = ~A299 & \new_[88379]_ ;
  assign \new_[88381]_  = \new_[88380]_  & \new_[88375]_ ;
  assign \new_[88382]_  = \new_[88381]_  & \new_[88372]_ ;
  assign \new_[88385]_  = ~A168 & A169;
  assign \new_[88388]_  = ~A166 & A167;
  assign \new_[88389]_  = \new_[88388]_  & \new_[88385]_ ;
  assign \new_[88392]_  = ~A200 & A199;
  assign \new_[88396]_  = ~A233 & A203;
  assign \new_[88397]_  = A201 & \new_[88396]_ ;
  assign \new_[88398]_  = \new_[88397]_  & \new_[88392]_ ;
  assign \new_[88399]_  = \new_[88398]_  & \new_[88389]_ ;
  assign \new_[88402]_  = ~A236 & ~A235;
  assign \new_[88405]_  = ~A268 & ~A266;
  assign \new_[88406]_  = \new_[88405]_  & \new_[88402]_ ;
  assign \new_[88409]_  = A298 & ~A269;
  assign \new_[88413]_  = A302 & A300;
  assign \new_[88414]_  = ~A299 & \new_[88413]_ ;
  assign \new_[88415]_  = \new_[88414]_  & \new_[88409]_ ;
  assign \new_[88416]_  = \new_[88415]_  & \new_[88406]_ ;
  assign \new_[88419]_  = ~A168 & A169;
  assign \new_[88422]_  = A166 & ~A167;
  assign \new_[88423]_  = \new_[88422]_  & \new_[88419]_ ;
  assign \new_[88426]_  = ~A200 & A199;
  assign \new_[88430]_  = ~A233 & A202;
  assign \new_[88431]_  = A201 & \new_[88430]_ ;
  assign \new_[88432]_  = \new_[88431]_  & \new_[88426]_ ;
  assign \new_[88433]_  = \new_[88432]_  & \new_[88423]_ ;
  assign \new_[88436]_  = ~A236 & ~A235;
  assign \new_[88439]_  = ~A268 & ~A266;
  assign \new_[88440]_  = \new_[88439]_  & \new_[88436]_ ;
  assign \new_[88443]_  = A298 & ~A269;
  assign \new_[88447]_  = A301 & A300;
  assign \new_[88448]_  = ~A299 & \new_[88447]_ ;
  assign \new_[88449]_  = \new_[88448]_  & \new_[88443]_ ;
  assign \new_[88450]_  = \new_[88449]_  & \new_[88440]_ ;
  assign \new_[88453]_  = ~A168 & A169;
  assign \new_[88456]_  = A166 & ~A167;
  assign \new_[88457]_  = \new_[88456]_  & \new_[88453]_ ;
  assign \new_[88460]_  = ~A200 & A199;
  assign \new_[88464]_  = ~A233 & A202;
  assign \new_[88465]_  = A201 & \new_[88464]_ ;
  assign \new_[88466]_  = \new_[88465]_  & \new_[88460]_ ;
  assign \new_[88467]_  = \new_[88466]_  & \new_[88457]_ ;
  assign \new_[88470]_  = ~A236 & ~A235;
  assign \new_[88473]_  = ~A268 & ~A266;
  assign \new_[88474]_  = \new_[88473]_  & \new_[88470]_ ;
  assign \new_[88477]_  = A298 & ~A269;
  assign \new_[88481]_  = A302 & A300;
  assign \new_[88482]_  = ~A299 & \new_[88481]_ ;
  assign \new_[88483]_  = \new_[88482]_  & \new_[88477]_ ;
  assign \new_[88484]_  = \new_[88483]_  & \new_[88474]_ ;
  assign \new_[88487]_  = ~A168 & A169;
  assign \new_[88490]_  = A166 & ~A167;
  assign \new_[88491]_  = \new_[88490]_  & \new_[88487]_ ;
  assign \new_[88494]_  = ~A200 & A199;
  assign \new_[88498]_  = ~A233 & A203;
  assign \new_[88499]_  = A201 & \new_[88498]_ ;
  assign \new_[88500]_  = \new_[88499]_  & \new_[88494]_ ;
  assign \new_[88501]_  = \new_[88500]_  & \new_[88491]_ ;
  assign \new_[88504]_  = ~A236 & ~A235;
  assign \new_[88507]_  = ~A268 & ~A266;
  assign \new_[88508]_  = \new_[88507]_  & \new_[88504]_ ;
  assign \new_[88511]_  = A298 & ~A269;
  assign \new_[88515]_  = A301 & A300;
  assign \new_[88516]_  = ~A299 & \new_[88515]_ ;
  assign \new_[88517]_  = \new_[88516]_  & \new_[88511]_ ;
  assign \new_[88518]_  = \new_[88517]_  & \new_[88508]_ ;
  assign \new_[88521]_  = ~A168 & A169;
  assign \new_[88524]_  = A166 & ~A167;
  assign \new_[88525]_  = \new_[88524]_  & \new_[88521]_ ;
  assign \new_[88528]_  = ~A200 & A199;
  assign \new_[88532]_  = ~A233 & A203;
  assign \new_[88533]_  = A201 & \new_[88532]_ ;
  assign \new_[88534]_  = \new_[88533]_  & \new_[88528]_ ;
  assign \new_[88535]_  = \new_[88534]_  & \new_[88525]_ ;
  assign \new_[88538]_  = ~A236 & ~A235;
  assign \new_[88541]_  = ~A268 & ~A266;
  assign \new_[88542]_  = \new_[88541]_  & \new_[88538]_ ;
  assign \new_[88545]_  = A298 & ~A269;
  assign \new_[88549]_  = A302 & A300;
  assign \new_[88550]_  = ~A299 & \new_[88549]_ ;
  assign \new_[88551]_  = \new_[88550]_  & \new_[88545]_ ;
  assign \new_[88552]_  = \new_[88551]_  & \new_[88542]_ ;
  assign \new_[88555]_  = ~A168 & ~A169;
  assign \new_[88558]_  = A166 & A167;
  assign \new_[88559]_  = \new_[88558]_  & \new_[88555]_ ;
  assign \new_[88562]_  = ~A200 & A199;
  assign \new_[88566]_  = ~A233 & A202;
  assign \new_[88567]_  = A201 & \new_[88566]_ ;
  assign \new_[88568]_  = \new_[88567]_  & \new_[88562]_ ;
  assign \new_[88569]_  = \new_[88568]_  & \new_[88559]_ ;
  assign \new_[88572]_  = ~A236 & ~A235;
  assign \new_[88575]_  = ~A268 & ~A266;
  assign \new_[88576]_  = \new_[88575]_  & \new_[88572]_ ;
  assign \new_[88579]_  = A298 & ~A269;
  assign \new_[88583]_  = A301 & A300;
  assign \new_[88584]_  = ~A299 & \new_[88583]_ ;
  assign \new_[88585]_  = \new_[88584]_  & \new_[88579]_ ;
  assign \new_[88586]_  = \new_[88585]_  & \new_[88576]_ ;
  assign \new_[88589]_  = ~A168 & ~A169;
  assign \new_[88592]_  = A166 & A167;
  assign \new_[88593]_  = \new_[88592]_  & \new_[88589]_ ;
  assign \new_[88596]_  = ~A200 & A199;
  assign \new_[88600]_  = ~A233 & A202;
  assign \new_[88601]_  = A201 & \new_[88600]_ ;
  assign \new_[88602]_  = \new_[88601]_  & \new_[88596]_ ;
  assign \new_[88603]_  = \new_[88602]_  & \new_[88593]_ ;
  assign \new_[88606]_  = ~A236 & ~A235;
  assign \new_[88609]_  = ~A268 & ~A266;
  assign \new_[88610]_  = \new_[88609]_  & \new_[88606]_ ;
  assign \new_[88613]_  = A298 & ~A269;
  assign \new_[88617]_  = A302 & A300;
  assign \new_[88618]_  = ~A299 & \new_[88617]_ ;
  assign \new_[88619]_  = \new_[88618]_  & \new_[88613]_ ;
  assign \new_[88620]_  = \new_[88619]_  & \new_[88610]_ ;
  assign \new_[88623]_  = ~A168 & ~A169;
  assign \new_[88626]_  = A166 & A167;
  assign \new_[88627]_  = \new_[88626]_  & \new_[88623]_ ;
  assign \new_[88630]_  = ~A200 & A199;
  assign \new_[88634]_  = ~A233 & A203;
  assign \new_[88635]_  = A201 & \new_[88634]_ ;
  assign \new_[88636]_  = \new_[88635]_  & \new_[88630]_ ;
  assign \new_[88637]_  = \new_[88636]_  & \new_[88627]_ ;
  assign \new_[88640]_  = ~A236 & ~A235;
  assign \new_[88643]_  = ~A268 & ~A266;
  assign \new_[88644]_  = \new_[88643]_  & \new_[88640]_ ;
  assign \new_[88647]_  = A298 & ~A269;
  assign \new_[88651]_  = A301 & A300;
  assign \new_[88652]_  = ~A299 & \new_[88651]_ ;
  assign \new_[88653]_  = \new_[88652]_  & \new_[88647]_ ;
  assign \new_[88654]_  = \new_[88653]_  & \new_[88644]_ ;
  assign \new_[88657]_  = ~A168 & ~A169;
  assign \new_[88660]_  = A166 & A167;
  assign \new_[88661]_  = \new_[88660]_  & \new_[88657]_ ;
  assign \new_[88664]_  = ~A200 & A199;
  assign \new_[88668]_  = ~A233 & A203;
  assign \new_[88669]_  = A201 & \new_[88668]_ ;
  assign \new_[88670]_  = \new_[88669]_  & \new_[88664]_ ;
  assign \new_[88671]_  = \new_[88670]_  & \new_[88661]_ ;
  assign \new_[88674]_  = ~A236 & ~A235;
  assign \new_[88677]_  = ~A268 & ~A266;
  assign \new_[88678]_  = \new_[88677]_  & \new_[88674]_ ;
  assign \new_[88681]_  = A298 & ~A269;
  assign \new_[88685]_  = A302 & A300;
  assign \new_[88686]_  = ~A299 & \new_[88685]_ ;
  assign \new_[88687]_  = \new_[88686]_  & \new_[88681]_ ;
  assign \new_[88688]_  = \new_[88687]_  & \new_[88678]_ ;
endmodule


