module top ( 
    _128_9_, _113_4_, _469_24_, _101_0_, _210_16_, _224_20_, _214_17_,
    _116_5_, _104_1_, _137_12_, _234_22_, _217_18_, _107_2_, _134_11_,
    _952_31_, _110_3_, _221_19_, _131_10_, _227_21_, _953_32_, _472_25_,
    _900_29_, _478_27_, _140_13_, _122_7_, _119_6_, _237_23_, _898_28_,
    _146_15_, _125_8_, _475_26_, _143_14_, _902_30_,
    _36_854_, _12_862_, _42_852_, _39_853_, _63_902_, _33_855_, _75_866_,
    _66_903_, _69_908_, _72_909_, _18_860_, _48_850_, _51_899_, _30_856_,
    _57_912_, _60_901_, _27_857_, _54_900_, _9_863_, _21_859_, _24_858_,
    _45_851_, _3_865_, _15_861_, _6_864_  );
  input  _128_9_, _113_4_, _469_24_, _101_0_, _210_16_, _224_20_,
    _214_17_, _116_5_, _104_1_, _137_12_, _234_22_, _217_18_, _107_2_,
    _134_11_, _952_31_, _110_3_, _221_19_, _131_10_, _227_21_, _953_32_,
    _472_25_, _900_29_, _478_27_, _140_13_, _122_7_, _119_6_, _237_23_,
    _898_28_, _146_15_, _125_8_, _475_26_, _143_14_, _902_30_;
  output _36_854_, _12_862_, _42_852_, _39_853_, _63_902_, _33_855_, _75_866_,
    _66_903_, _69_908_, _72_909_, _18_860_, _48_850_, _51_899_, _30_856_,
    _57_912_, _60_901_, _27_857_, _54_900_, _9_863_, _21_859_, _24_858_,
    _45_851_, _3_865_, _15_861_, _6_864_;
  wire new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n330_, new_n331_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n411_, new_n412_, new_n414_, new_n415_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n425_,
    new_n426_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n441_, new_n442_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n449_, new_n450_, new_n452_, new_n453_, new_n455_, new_n456_,
    new_n458_, new_n459_, new_n461_, new_n462_, new_n464_, new_n465_,
    new_n467_, new_n468_;
  assign new_n59_ = ~_140_13_ & _125_8_;
  assign new_n60_ = _140_13_ & ~_125_8_;
  assign new_n61_ = ~new_n59_ & ~new_n60_;
  assign new_n62_ = ~_146_15_ & new_n61_;
  assign new_n63_ = _146_15_ & ~new_n61_;
  assign new_n64_ = ~new_n62_ & ~new_n63_;
  assign new_n65_ = ~_953_32_ & ~_237_23_;
  assign new_n66_ = _214_17_ & new_n65_;
  assign new_n67_ = _143_14_ & new_n66_;
  assign new_n68_ = ~_143_14_ & ~new_n66_;
  assign new_n69_ = ~new_n67_ & ~new_n68_;
  assign new_n70_ = ~_131_10_ & new_n69_;
  assign new_n71_ = _131_10_ & ~new_n69_;
  assign new_n72_ = ~new_n70_ & ~new_n71_;
  assign new_n73_ = new_n64_ & ~new_n72_;
  assign new_n74_ = ~new_n64_ & new_n72_;
  assign new_n75_ = ~new_n73_ & ~new_n74_;
  assign new_n76_ = ~_113_4_ & _122_7_;
  assign new_n77_ = _113_4_ & ~_122_7_;
  assign new_n78_ = ~new_n76_ & ~new_n77_;
  assign new_n79_ = ~_104_1_ & new_n78_;
  assign new_n80_ = _104_1_ & ~new_n78_;
  assign new_n81_ = ~new_n79_ & ~new_n80_;
  assign new_n82_ = new_n75_ & ~new_n81_;
  assign new_n83_ = ~new_n75_ & new_n81_;
  assign new_n84_ = ~new_n82_ & ~new_n83_;
  assign new_n85_ = ~_902_30_ & ~new_n84_;
  assign new_n86_ = ~_475_26_ & new_n85_;
  assign new_n87_ = _475_26_ & ~new_n85_;
  assign new_n88_ = ~new_n86_ & ~new_n87_;
  assign new_n89_ = ~_116_5_ & _122_7_;
  assign new_n90_ = _116_5_ & ~_122_7_;
  assign new_n91_ = ~new_n89_ & ~new_n90_;
  assign new_n92_ = ~_107_2_ & new_n91_;
  assign new_n93_ = _107_2_ & ~new_n91_;
  assign new_n94_ = ~new_n92_ & ~new_n93_;
  assign new_n95_ = ~_128_9_ & _143_14_;
  assign new_n96_ = _128_9_ & ~_143_14_;
  assign new_n97_ = ~new_n95_ & ~new_n96_;
  assign new_n98_ = ~_134_11_ & new_n97_;
  assign new_n99_ = _134_11_ & ~new_n97_;
  assign new_n100_ = ~new_n98_ & ~new_n99_;
  assign new_n101_ = new_n94_ & ~new_n100_;
  assign new_n102_ = ~new_n94_ & new_n100_;
  assign new_n103_ = ~new_n101_ & ~new_n102_;
  assign new_n104_ = _234_22_ & ~_953_32_;
  assign new_n105_ = _217_18_ & new_n104_;
  assign new_n106_ = new_n103_ & new_n105_;
  assign new_n107_ = ~new_n103_ & ~new_n105_;
  assign new_n108_ = ~new_n106_ & ~new_n107_;
  assign new_n109_ = ~_902_30_ & ~new_n108_;
  assign new_n110_ = ~_478_27_ & new_n109_;
  assign new_n111_ = _478_27_ & ~new_n109_;
  assign new_n112_ = ~new_n110_ & ~new_n111_;
  assign new_n113_ = new_n88_ & ~new_n112_;
  assign new_n114_ = _234_22_ & _237_23_;
  assign new_n115_ = ~_953_32_ & ~new_n114_;
  assign new_n116_ = _952_31_ & new_n115_;
  assign new_n117_ = _902_30_ & ~new_n114_;
  assign new_n118_ = _953_32_ & new_n117_;
  assign new_n119_ = ~_900_29_ & new_n118_;
  assign new_n120_ = ~new_n116_ & ~new_n119_;
  assign new_n121_ = _110_3_ & ~_140_13_;
  assign new_n122_ = ~_110_3_ & _140_13_;
  assign new_n123_ = ~new_n121_ & ~new_n122_;
  assign new_n124_ = _227_21_ & ~_953_32_;
  assign new_n125_ = new_n123_ & new_n124_;
  assign new_n126_ = ~new_n123_ & ~new_n124_;
  assign new_n127_ = ~new_n125_ & ~new_n126_;
  assign new_n128_ = ~_104_1_ & _107_2_;
  assign new_n129_ = _104_1_ & ~_107_2_;
  assign new_n130_ = ~new_n128_ & ~new_n129_;
  assign new_n131_ = ~_101_0_ & new_n130_;
  assign new_n132_ = _101_0_ & ~new_n130_;
  assign new_n133_ = ~new_n131_ & ~new_n132_;
  assign new_n134_ = _146_15_ & ~_143_14_;
  assign new_n135_ = ~_146_15_ & _143_14_;
  assign new_n136_ = ~new_n134_ & ~new_n135_;
  assign new_n137_ = ~_128_9_ & new_n136_;
  assign new_n138_ = _128_9_ & ~new_n136_;
  assign new_n139_ = ~new_n137_ & ~new_n138_;
  assign new_n140_ = new_n133_ & new_n139_;
  assign new_n141_ = ~new_n133_ & ~new_n139_;
  assign new_n142_ = ~new_n140_ & ~new_n141_;
  assign new_n143_ = _137_12_ & ~_134_11_;
  assign new_n144_ = ~_137_12_ & _134_11_;
  assign new_n145_ = ~new_n143_ & ~new_n144_;
  assign new_n146_ = ~_131_10_ & new_n145_;
  assign new_n147_ = _131_10_ & ~new_n145_;
  assign new_n148_ = ~new_n146_ & ~new_n147_;
  assign new_n149_ = new_n142_ & new_n148_;
  assign new_n150_ = ~new_n142_ & ~new_n148_;
  assign new_n151_ = ~new_n149_ & ~new_n150_;
  assign new_n152_ = new_n127_ & new_n151_;
  assign new_n153_ = ~new_n127_ & ~new_n151_;
  assign new_n154_ = ~new_n152_ & ~new_n153_;
  assign new_n155_ = ~_902_30_ & ~new_n154_;
  assign new_n156_ = ~_469_24_ & new_n155_;
  assign new_n157_ = _469_24_ & ~new_n155_;
  assign new_n158_ = ~new_n156_ & ~new_n157_;
  assign new_n159_ = _234_22_ & ~_902_30_;
  assign new_n160_ = _221_19_ & ~new_n159_;
  assign new_n161_ = ~new_n158_ & ~new_n160_;
  assign new_n162_ = _210_16_ & new_n65_;
  assign new_n163_ = _101_0_ & new_n162_;
  assign new_n164_ = ~_101_0_ & ~new_n162_;
  assign new_n165_ = ~new_n163_ & ~new_n164_;
  assign new_n166_ = ~new_n139_ & ~new_n148_;
  assign new_n167_ = new_n139_ & new_n148_;
  assign new_n168_ = ~new_n166_ & ~new_n167_;
  assign new_n169_ = ~_116_5_ & _119_6_;
  assign new_n170_ = _116_5_ & ~_119_6_;
  assign new_n171_ = ~new_n169_ & ~new_n170_;
  assign new_n172_ = ~_113_4_ & new_n171_;
  assign new_n173_ = _113_4_ & ~new_n171_;
  assign new_n174_ = ~new_n172_ & ~new_n173_;
  assign new_n175_ = new_n168_ & new_n174_;
  assign new_n176_ = ~new_n168_ & ~new_n174_;
  assign new_n177_ = ~new_n175_ & ~new_n176_;
  assign new_n178_ = ~new_n165_ & new_n177_;
  assign new_n179_ = new_n165_ & ~new_n177_;
  assign new_n180_ = ~new_n178_ & ~new_n179_;
  assign new_n181_ = ~_902_30_ & ~new_n180_;
  assign new_n182_ = ~_472_25_ & new_n181_;
  assign new_n183_ = _472_25_ & ~new_n181_;
  assign new_n184_ = ~new_n182_ & ~new_n183_;
  assign new_n185_ = _128_9_ & ~_119_6_;
  assign new_n186_ = ~_128_9_ & _119_6_;
  assign new_n187_ = ~new_n185_ & ~new_n186_;
  assign new_n188_ = ~_110_3_ & new_n187_;
  assign new_n189_ = _110_3_ & ~new_n187_;
  assign new_n190_ = ~new_n188_ & ~new_n189_;
  assign new_n191_ = ~new_n64_ & new_n190_;
  assign new_n192_ = new_n64_ & ~new_n190_;
  assign new_n193_ = ~new_n191_ & ~new_n192_;
  assign new_n194_ = _221_19_ & new_n104_;
  assign new_n195_ = ~_137_12_ & ~new_n194_;
  assign new_n196_ = _137_12_ & new_n194_;
  assign new_n197_ = ~new_n195_ & ~new_n196_;
  assign new_n198_ = new_n193_ & new_n197_;
  assign new_n199_ = ~new_n193_ & ~new_n197_;
  assign new_n200_ = ~new_n198_ & ~new_n199_;
  assign new_n201_ = ~_902_30_ & ~new_n200_;
  assign new_n202_ = _217_18_ & ~new_n159_;
  assign new_n203_ = new_n201_ & ~new_n202_;
  assign new_n204_ = ~new_n201_ & new_n202_;
  assign new_n205_ = ~new_n203_ & ~new_n204_;
  assign new_n206_ = ~new_n184_ & new_n205_;
  assign new_n207_ = ~_125_8_ & new_n139_;
  assign new_n208_ = _125_8_ & ~new_n139_;
  assign new_n209_ = ~new_n207_ & ~new_n208_;
  assign new_n210_ = _224_20_ & ~_953_32_;
  assign new_n211_ = new_n209_ & new_n210_;
  assign new_n212_ = ~new_n209_ & ~new_n210_;
  assign new_n213_ = ~new_n211_ & ~new_n212_;
  assign new_n214_ = ~new_n133_ & ~new_n174_;
  assign new_n215_ = new_n133_ & new_n174_;
  assign new_n216_ = ~new_n214_ & ~new_n215_;
  assign new_n217_ = ~_110_3_ & _122_7_;
  assign new_n218_ = _110_3_ & ~_122_7_;
  assign new_n219_ = ~new_n217_ & ~new_n218_;
  assign new_n220_ = new_n216_ & new_n219_;
  assign new_n221_ = ~new_n216_ & ~new_n219_;
  assign new_n222_ = ~new_n220_ & ~new_n221_;
  assign new_n223_ = ~new_n213_ & ~new_n222_;
  assign new_n224_ = new_n213_ & new_n222_;
  assign new_n225_ = ~new_n223_ & ~new_n224_;
  assign new_n226_ = ~_902_30_ & new_n225_;
  assign new_n227_ = ~_237_23_ & ~_902_30_;
  assign new_n228_ = _210_16_ & ~new_n227_;
  assign new_n229_ = new_n226_ & ~new_n228_;
  assign new_n230_ = ~new_n226_ & new_n228_;
  assign new_n231_ = ~new_n229_ & ~new_n230_;
  assign new_n232_ = _214_17_ & ~new_n227_;
  assign new_n233_ = new_n231_ & ~new_n232_;
  assign new_n234_ = new_n113_ & ~new_n120_;
  assign new_n235_ = new_n161_ & new_n234_;
  assign new_n236_ = new_n206_ & new_n235_;
  assign new_n237_ = new_n233_ & new_n236_;
  assign new_n238_ = _134_11_ & ~new_n237_;
  assign new_n239_ = ~_134_11_ & new_n237_;
  assign _36_854_ = new_n238_ | new_n239_;
  assign new_n241_ = new_n88_ & new_n112_;
  assign new_n242_ = ~_898_28_ & new_n118_;
  assign new_n243_ = ~new_n116_ & ~new_n242_;
  assign new_n244_ = new_n184_ & ~new_n205_;
  assign new_n245_ = ~new_n231_ & ~new_n232_;
  assign new_n246_ = new_n241_ & ~new_n243_;
  assign new_n247_ = new_n161_ & new_n246_;
  assign new_n248_ = new_n244_ & new_n247_;
  assign new_n249_ = new_n245_ & new_n248_;
  assign new_n250_ = _110_3_ & ~new_n249_;
  assign new_n251_ = ~_110_3_ & new_n249_;
  assign _12_862_ = new_n250_ | new_n251_;
  assign new_n253_ = ~new_n88_ & new_n112_;
  assign new_n254_ = ~new_n120_ & new_n253_;
  assign new_n255_ = new_n161_ & new_n254_;
  assign new_n256_ = new_n244_ & new_n255_;
  assign new_n257_ = new_n233_ & new_n256_;
  assign new_n258_ = _140_13_ & ~new_n257_;
  assign new_n259_ = ~_140_13_ & new_n257_;
  assign _42_852_ = new_n258_ | new_n259_;
  assign new_n261_ = ~new_n184_ & ~new_n205_;
  assign new_n262_ = ~new_n120_ & new_n241_;
  assign new_n263_ = new_n161_ & new_n262_;
  assign new_n264_ = new_n261_ & new_n263_;
  assign new_n265_ = new_n233_ & new_n264_;
  assign new_n266_ = _137_12_ & ~new_n265_;
  assign new_n267_ = ~_137_12_ & new_n265_;
  assign _39_853_ = new_n266_ | new_n267_;
  assign new_n269_ = ~_952_31_ & _953_32_;
  assign new_n270_ = new_n235_ & new_n261_;
  assign new_n271_ = new_n245_ & new_n270_;
  assign new_n272_ = new_n206_ & new_n255_;
  assign new_n273_ = new_n233_ & new_n272_;
  assign new_n274_ = new_n158_ & ~new_n160_;
  assign new_n275_ = new_n254_ & new_n274_;
  assign new_n276_ = new_n244_ & new_n275_;
  assign new_n277_ = new_n245_ & new_n276_;
  assign new_n278_ = new_n255_ & new_n261_;
  assign new_n279_ = new_n245_ & new_n278_;
  assign new_n280_ = ~new_n88_ & ~new_n112_;
  assign new_n281_ = ~new_n120_ & new_n280_;
  assign new_n282_ = new_n161_ & new_n281_;
  assign new_n283_ = new_n206_ & new_n282_;
  assign new_n284_ = new_n245_ & new_n283_;
  assign new_n285_ = ~new_n237_ & ~new_n265_;
  assign new_n286_ = ~new_n271_ & new_n285_;
  assign new_n287_ = ~new_n273_ & new_n286_;
  assign new_n288_ = ~new_n277_ & new_n287_;
  assign new_n289_ = ~new_n279_ & new_n288_;
  assign new_n290_ = ~new_n257_ & new_n289_;
  assign new_n291_ = ~new_n284_ & new_n290_;
  assign new_n292_ = ~new_n243_ & new_n253_;
  assign new_n293_ = new_n274_ & new_n292_;
  assign new_n294_ = new_n206_ & new_n293_;
  assign new_n295_ = new_n245_ & new_n294_;
  assign new_n296_ = new_n184_ & new_n205_;
  assign new_n297_ = new_n161_ & new_n292_;
  assign new_n298_ = new_n296_ & new_n297_;
  assign new_n299_ = new_n245_ & new_n298_;
  assign new_n300_ = new_n113_ & ~new_n243_;
  assign new_n301_ = new_n161_ & new_n300_;
  assign new_n302_ = new_n296_ & new_n301_;
  assign new_n303_ = new_n245_ & new_n302_;
  assign new_n304_ = new_n206_ & new_n247_;
  assign new_n305_ = new_n245_ & new_n304_;
  assign new_n306_ = ~new_n243_ & new_n280_;
  assign new_n307_ = new_n274_ & new_n306_;
  assign new_n308_ = new_n296_ & new_n307_;
  assign new_n309_ = new_n245_ & new_n308_;
  assign new_n310_ = new_n274_ & new_n300_;
  assign new_n311_ = new_n206_ & new_n310_;
  assign new_n312_ = new_n245_ & new_n311_;
  assign new_n313_ = new_n246_ & new_n274_;
  assign new_n314_ = new_n261_ & new_n313_;
  assign new_n315_ = new_n245_ & new_n314_;
  assign new_n316_ = ~new_n249_ & ~new_n295_;
  assign new_n317_ = ~new_n299_ & new_n316_;
  assign new_n318_ = ~new_n303_ & new_n317_;
  assign new_n319_ = ~new_n305_ & new_n318_;
  assign new_n320_ = ~new_n309_ & new_n319_;
  assign new_n321_ = ~new_n312_ & new_n320_;
  assign new_n322_ = ~new_n315_ & new_n321_;
  assign new_n323_ = new_n291_ & new_n322_;
  assign new_n324_ = _902_30_ & ~new_n323_;
  assign new_n325_ = _478_27_ & new_n324_;
  assign new_n326_ = new_n108_ & new_n325_;
  assign new_n327_ = ~new_n108_ & ~new_n325_;
  assign new_n328_ = ~new_n326_ & ~new_n327_;
  assign _63_902_ = ~new_n269_ & ~new_n328_;
  assign new_n330_ = _131_10_ & ~new_n273_;
  assign new_n331_ = ~_131_10_ & new_n273_;
  assign _33_855_ = new_n330_ | new_n331_;
  assign new_n333_ = new_n116_ & new_n253_;
  assign new_n334_ = new_n274_ & new_n333_;
  assign new_n335_ = new_n296_ & new_n334_;
  assign new_n336_ = new_n233_ & new_n335_;
  assign new_n337_ = new_n113_ & new_n116_;
  assign new_n338_ = new_n274_ & new_n337_;
  assign new_n339_ = new_n296_ & new_n338_;
  assign new_n340_ = new_n233_ & new_n339_;
  assign new_n341_ = new_n116_ & new_n241_;
  assign new_n342_ = new_n161_ & new_n341_;
  assign new_n343_ = new_n296_ & new_n342_;
  assign new_n344_ = new_n233_ & new_n343_;
  assign new_n345_ = new_n274_ & new_n341_;
  assign new_n346_ = new_n206_ & new_n345_;
  assign new_n347_ = new_n233_ & new_n346_;
  assign new_n348_ = new_n296_ & new_n345_;
  assign new_n349_ = new_n245_ & new_n348_;
  assign new_n350_ = new_n231_ & new_n232_;
  assign new_n351_ = new_n348_ & new_n350_;
  assign new_n352_ = new_n244_ & new_n345_;
  assign new_n353_ = new_n233_ & new_n352_;
  assign new_n354_ = new_n158_ & new_n160_;
  assign new_n355_ = new_n341_ & new_n354_;
  assign new_n356_ = new_n296_ & new_n355_;
  assign new_n357_ = new_n233_ & new_n356_;
  assign new_n358_ = ~new_n336_ & ~new_n340_;
  assign new_n359_ = ~new_n344_ & new_n358_;
  assign new_n360_ = ~new_n347_ & new_n359_;
  assign new_n361_ = ~new_n349_ & new_n360_;
  assign new_n362_ = ~new_n351_ & new_n361_;
  assign new_n363_ = ~new_n353_ & new_n362_;
  assign new_n364_ = ~new_n357_ & new_n363_;
  assign new_n365_ = new_n291_ & new_n364_;
  assign new_n366_ = new_n322_ & new_n365_;
  assign new_n367_ = new_n184_ & ~new_n232_;
  assign new_n368_ = new_n112_ & new_n367_;
  assign new_n369_ = new_n88_ & new_n368_;
  assign new_n370_ = new_n205_ & new_n369_;
  assign new_n371_ = ~new_n160_ & new_n370_;
  assign new_n372_ = new_n158_ & new_n371_;
  assign new_n373_ = new_n231_ & new_n372_;
  assign new_n374_ = new_n366_ & ~new_n373_;
  assign new_n375_ = _952_31_ & new_n374_;
  assign new_n376_ = ~_953_32_ & new_n375_;
  assign new_n377_ = ~_952_31_ & ~new_n373_;
  assign new_n378_ = ~_952_31_ & new_n377_;
  assign new_n379_ = ~_953_32_ & new_n378_;
  assign _75_866_ = ~new_n376_ & ~new_n379_;
  assign new_n381_ = new_n202_ & new_n324_;
  assign new_n382_ = new_n200_ & new_n381_;
  assign new_n383_ = ~new_n200_ & ~new_n381_;
  assign new_n384_ = ~new_n382_ & ~new_n383_;
  assign _66_903_ = ~new_n269_ & ~new_n384_;
  assign new_n386_ = ~_953_32_ & ~new_n322_;
  assign new_n387_ = _953_32_ & ~_898_28_;
  assign new_n388_ = new_n222_ & ~new_n387_;
  assign new_n389_ = ~new_n386_ & new_n388_;
  assign new_n390_ = new_n386_ & ~new_n388_;
  assign new_n391_ = ~new_n389_ & ~new_n390_;
  assign new_n392_ = _224_20_ & _898_28_;
  assign new_n393_ = _953_32_ & ~new_n392_;
  assign new_n394_ = new_n391_ & new_n393_;
  assign new_n395_ = ~new_n391_ & ~new_n393_;
  assign _69_908_ = new_n394_ | new_n395_;
  assign new_n397_ = ~_953_32_ & ~new_n291_;
  assign new_n398_ = new_n61_ & new_n168_;
  assign new_n399_ = ~new_n61_ & ~new_n168_;
  assign new_n400_ = ~new_n398_ & ~new_n399_;
  assign new_n401_ = _953_32_ & ~_900_29_;
  assign new_n402_ = new_n400_ & ~new_n401_;
  assign new_n403_ = ~new_n397_ & new_n402_;
  assign new_n404_ = new_n397_ & ~new_n402_;
  assign new_n405_ = ~new_n403_ & ~new_n404_;
  assign new_n406_ = _227_21_ & _900_29_;
  assign new_n407_ = _953_32_ & ~new_n406_;
  assign new_n408_ = new_n405_ & new_n407_;
  assign new_n409_ = ~new_n405_ & ~new_n407_;
  assign _72_909_ = new_n408_ | new_n409_;
  assign new_n411_ = _116_5_ & ~new_n312_;
  assign new_n412_ = ~_116_5_ & new_n312_;
  assign _18_860_ = new_n411_ | new_n412_;
  assign new_n414_ = _146_15_ & ~new_n279_;
  assign new_n415_ = ~_146_15_ & new_n279_;
  assign _48_850_ = new_n414_ | new_n415_;
  assign new_n417_ = new_n213_ & ~new_n222_;
  assign new_n418_ = ~new_n213_ & new_n222_;
  assign new_n419_ = ~new_n417_ & ~new_n418_;
  assign new_n420_ = new_n228_ & new_n324_;
  assign new_n421_ = new_n419_ & new_n420_;
  assign new_n422_ = ~new_n419_ & ~new_n420_;
  assign new_n423_ = ~new_n421_ & ~new_n422_;
  assign _51_899_ = ~new_n269_ & ~new_n423_;
  assign new_n425_ = _128_9_ & ~new_n271_;
  assign new_n426_ = ~_128_9_ & new_n271_;
  assign _30_856_ = new_n425_ | new_n426_;
  assign new_n428_ = _472_25_ & new_n324_;
  assign new_n429_ = new_n177_ & new_n428_;
  assign new_n430_ = ~new_n177_ & ~new_n428_;
  assign new_n431_ = ~new_n429_ & ~new_n430_;
  assign new_n432_ = ~new_n165_ & new_n431_;
  assign new_n433_ = new_n165_ & ~new_n431_;
  assign new_n434_ = ~new_n432_ & ~new_n433_;
  assign _57_912_ = ~new_n269_ & ~new_n434_;
  assign new_n436_ = _475_26_ & new_n324_;
  assign new_n437_ = new_n84_ & new_n436_;
  assign new_n438_ = ~new_n84_ & ~new_n436_;
  assign new_n439_ = ~new_n437_ & ~new_n438_;
  assign _60_901_ = ~new_n269_ & ~new_n439_;
  assign new_n441_ = _125_8_ & ~new_n277_;
  assign new_n442_ = ~_125_8_ & new_n277_;
  assign _27_857_ = new_n441_ | new_n442_;
  assign new_n444_ = _469_24_ & new_n324_;
  assign new_n445_ = new_n154_ & new_n444_;
  assign new_n446_ = ~new_n154_ & ~new_n444_;
  assign new_n447_ = ~new_n445_ & ~new_n446_;
  assign _54_900_ = ~new_n269_ & ~new_n447_;
  assign new_n449_ = _107_2_ & ~new_n303_;
  assign new_n450_ = ~_107_2_ & new_n303_;
  assign _9_863_ = new_n449_ | new_n450_;
  assign new_n452_ = _119_6_ & ~new_n315_;
  assign new_n453_ = ~_119_6_ & new_n315_;
  assign _21_859_ = new_n452_ | new_n453_;
  assign new_n455_ = _122_7_ & ~new_n309_;
  assign new_n456_ = ~_122_7_ & new_n309_;
  assign _24_858_ = new_n455_ | new_n456_;
  assign new_n458_ = _143_14_ & ~new_n284_;
  assign new_n459_ = ~_143_14_ & new_n284_;
  assign _45_851_ = new_n458_ | new_n459_;
  assign new_n461_ = _101_0_ & ~new_n305_;
  assign new_n462_ = ~_101_0_ & new_n305_;
  assign _3_865_ = new_n461_ | new_n462_;
  assign new_n464_ = _113_4_ & ~new_n295_;
  assign new_n465_ = ~_113_4_ & new_n295_;
  assign _15_861_ = new_n464_ | new_n465_;
  assign new_n467_ = _104_1_ & ~new_n299_;
  assign new_n468_ = ~_104_1_ & new_n299_;
  assign _6_864_ = new_n467_ | new_n468_;
endmodule

