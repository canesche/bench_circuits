module top ( 
    pp, pq, pr, ps, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn,
    po,
    pa0, pb0, pt, pu, pv, pw, px, py, pz  );
  input  pp, pq, pr, ps, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk, pl,
    pm, pn, po;
  output pa0, pb0, pt, pu, pv, pw, px, py, pz;
  wire new_n29_, new_n30_, new_n31_, new_n32_, new_n33_, new_n34_, new_n35_,
    new_n36_, new_n37_, new_n38_, new_n39_, new_n40_, new_n41_, new_n43_,
    new_n44_, new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n51_,
    new_n53_, new_n54_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_,
    new_n61_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_,
    new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n77_,
    new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n89_;
  assign new_n29_ = pl & pm;
  assign new_n30_ = pn & new_n29_;
  assign new_n31_ = po & new_n30_;
  assign new_n32_ = pp & new_n31_;
  assign new_n33_ = pq & new_n32_;
  assign new_n34_ = pj & ~pk;
  assign new_n35_ = ~pi & new_n34_;
  assign new_n36_ = ~pr & new_n33_;
  assign new_n37_ = new_n35_ & new_n36_;
  assign new_n38_ = pr & ~new_n33_;
  assign new_n39_ = new_n35_ & new_n38_;
  assign new_n40_ = pg & pi;
  assign new_n41_ = ~new_n37_ & ~new_n39_;
  assign pa0 = new_n40_ | ~new_n41_;
  assign new_n43_ = pr & new_n33_;
  assign new_n44_ = ~ps & new_n43_;
  assign new_n45_ = new_n35_ & new_n44_;
  assign new_n46_ = ps & ~new_n43_;
  assign new_n47_ = new_n35_ & new_n46_;
  assign new_n48_ = ph & pi;
  assign new_n49_ = ~new_n45_ & ~new_n47_;
  assign pb0 = new_n48_ | ~new_n49_;
  assign new_n51_ = new_n35_ & new_n43_;
  assign pt = ps & new_n51_;
  assign new_n53_ = ~pl & new_n35_;
  assign new_n54_ = pa & pi;
  assign pu = new_n53_ | new_n54_;
  assign new_n56_ = ~pl & pm;
  assign new_n57_ = new_n35_ & new_n56_;
  assign new_n58_ = pl & ~pm;
  assign new_n59_ = new_n35_ & new_n58_;
  assign new_n60_ = pb & pi;
  assign new_n61_ = ~new_n57_ & ~new_n59_;
  assign pv = new_n60_ | ~new_n61_;
  assign new_n63_ = ~pn & new_n29_;
  assign new_n64_ = new_n35_ & new_n63_;
  assign new_n65_ = pn & ~new_n29_;
  assign new_n66_ = new_n35_ & new_n65_;
  assign new_n67_ = pc & pi;
  assign new_n68_ = ~new_n64_ & ~new_n66_;
  assign pw = new_n67_ | ~new_n68_;
  assign new_n70_ = ~po & new_n30_;
  assign new_n71_ = new_n35_ & new_n70_;
  assign new_n72_ = po & ~new_n30_;
  assign new_n73_ = new_n35_ & new_n72_;
  assign new_n74_ = pd & pi;
  assign new_n75_ = ~new_n71_ & ~new_n73_;
  assign px = new_n74_ | ~new_n75_;
  assign new_n77_ = ~pp & new_n31_;
  assign new_n78_ = new_n35_ & new_n77_;
  assign new_n79_ = pp & ~new_n31_;
  assign new_n80_ = new_n35_ & new_n79_;
  assign new_n81_ = pe & pi;
  assign new_n82_ = ~new_n78_ & ~new_n80_;
  assign py = new_n81_ | ~new_n82_;
  assign new_n84_ = ~pq & new_n32_;
  assign new_n85_ = new_n35_ & new_n84_;
  assign new_n86_ = pq & ~new_n32_;
  assign new_n87_ = new_n35_ & new_n86_;
  assign new_n88_ = pf & pi;
  assign new_n89_ = ~new_n85_ & ~new_n87_;
  assign pz = new_n88_ | ~new_n89_;
endmodule

