module MultiplierB_32 ( clock, 
    \1 , 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20,
    21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33,
    98  );
  input  clock;
  input  \1 , 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18,
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33;
  output 98;
  reg 34, 2, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51,
    52, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69,
    70, 71, 72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87,
    88, 89, 90, 91, 92, 93, 94, 95;
  wire new_n220_, new_n221_, new_n222_, new_n223_1_, new_n224_, new_n225_,
    new_n228_1_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_1_,
    new_n235_, new_n236_, new_n237_, new_n238_1_, new_n239_, new_n240_,
    new_n242_, new_n243_1_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_1_, new_n254_,
    new_n256_, new_n257_, new_n258_1_, new_n259_, new_n260_, new_n261_,
    new_n263_1_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_1_,
    new_n270_, new_n271_, new_n272_, new_n273_1_, new_n274_, new_n275_,
    new_n277_, new_n278_1_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_1_, new_n289_,
    new_n291_, new_n292_, new_n293_1_, new_n294_, new_n295_, new_n296_,
    new_n298_1_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_1_,
    new_n305_, new_n306_, new_n307_, new_n308_1_, new_n309_, new_n310_,
    new_n312_, new_n313_1_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_1_, new_n324_,
    new_n326_, new_n327_, new_n328_1_, new_n329_, new_n330_, new_n331_,
    new_n333_1_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_1_,
    new_n340_, new_n341_, new_n342_, new_n343_1_, new_n344_, new_n345_,
    new_n347_, new_n348_1_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_1_, new_n359_,
    new_n361_, new_n362_, new_n363_1_, new_n364_, new_n365_, new_n366_,
    new_n368_1_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_1_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n431_, new_n432_, new_n433_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n440_, new_n441_, new_n442_, new_n443_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n455_, new_n456_, new_n457_, new_n458_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n470_, new_n471_, new_n472_, new_n473_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n485_, new_n486_, new_n487_, new_n488_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n500_, new_n501_, new_n502_, new_n503_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n515_, new_n516_, new_n517_, new_n518_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n530_, new_n531_, new_n532_, new_n533_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n545_, new_n546_, new_n547_, new_n548_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n560_, new_n561_, new_n562_, new_n563_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n575_, new_n576_, new_n577_, new_n578_, new_n580_,
    new_n581_, new_n582_, new_n583_, n68, n73, n78, n83, n88, n93, n98,
    n103, n108, n113, n118, n123, n128, n133, n138, n143, n148, n153, n158,
    n163, n168, n173, n178, n183, n188, n193, n198, n203, n208, n213, n218,
    n223, n228, n233, n238, n243, n248, n253, n258, n263, n268, n273, n278,
    n283, n288, n293, n298, n303, n308, n313, n318, n323, n328, n333, n338,
    n343, n348, n353, n358, n363, n368, n373;
  assign new_n220_ = \1  & 3;
  assign new_n221_ = ~36 & 66;
  assign new_n222_ = 36 & ~66;
  assign new_n223_1_ = ~new_n221_ & ~new_n222_;
  assign new_n224_ = new_n220_ & new_n223_1_;
  assign new_n225_ = ~new_n220_ & ~new_n223_1_;
  assign 98 = new_n224_ | new_n225_;
  assign n68 = \1  & 34;
  assign new_n228_1_ = \1  & 4;
  assign new_n229_ = ~37 & 67;
  assign new_n230_ = 37 & ~67;
  assign new_n231_ = ~new_n229_ & ~new_n230_;
  assign new_n232_ = new_n228_1_ & new_n231_;
  assign new_n233_1_ = ~new_n228_1_ & ~new_n231_;
  assign n73 = new_n232_ | new_n233_1_;
  assign new_n235_ = \1  & 5;
  assign new_n236_ = ~38 & 68;
  assign new_n237_ = 38 & ~68;
  assign new_n238_1_ = ~new_n236_ & ~new_n237_;
  assign new_n239_ = new_n235_ & new_n238_1_;
  assign new_n240_ = ~new_n235_ & ~new_n238_1_;
  assign n78 = new_n239_ | new_n240_;
  assign new_n242_ = \1  & 6;
  assign new_n243_1_ = ~39 & 69;
  assign new_n244_ = 39 & ~69;
  assign new_n245_ = ~new_n243_1_ & ~new_n244_;
  assign new_n246_ = new_n242_ & new_n245_;
  assign new_n247_ = ~new_n242_ & ~new_n245_;
  assign n83 = new_n246_ | new_n247_;
  assign new_n249_ = \1  & 7;
  assign new_n250_ = ~40 & 70;
  assign new_n251_ = 40 & ~70;
  assign new_n252_ = ~new_n250_ & ~new_n251_;
  assign new_n253_1_ = new_n249_ & new_n252_;
  assign new_n254_ = ~new_n249_ & ~new_n252_;
  assign n88 = new_n253_1_ | new_n254_;
  assign new_n256_ = \1  & 8;
  assign new_n257_ = ~41 & 71;
  assign new_n258_1_ = 41 & ~71;
  assign new_n259_ = ~new_n257_ & ~new_n258_1_;
  assign new_n260_ = new_n256_ & new_n259_;
  assign new_n261_ = ~new_n256_ & ~new_n259_;
  assign n93 = new_n260_ | new_n261_;
  assign new_n263_1_ = \1  & 9;
  assign new_n264_ = ~42 & 72;
  assign new_n265_ = 42 & ~72;
  assign new_n266_ = ~new_n264_ & ~new_n265_;
  assign new_n267_ = new_n263_1_ & new_n266_;
  assign new_n268_1_ = ~new_n263_1_ & ~new_n266_;
  assign n98 = new_n267_ | new_n268_1_;
  assign new_n270_ = \1  & 10;
  assign new_n271_ = ~43 & 73;
  assign new_n272_ = 43 & ~73;
  assign new_n273_1_ = ~new_n271_ & ~new_n272_;
  assign new_n274_ = new_n270_ & new_n273_1_;
  assign new_n275_ = ~new_n270_ & ~new_n273_1_;
  assign n103 = new_n274_ | new_n275_;
  assign new_n277_ = \1  & 11;
  assign new_n278_1_ = ~44 & 74;
  assign new_n279_ = 44 & ~74;
  assign new_n280_ = ~new_n278_1_ & ~new_n279_;
  assign new_n281_ = new_n277_ & new_n280_;
  assign new_n282_ = ~new_n277_ & ~new_n280_;
  assign n108 = new_n281_ | new_n282_;
  assign new_n284_ = \1  & 12;
  assign new_n285_ = ~45 & 75;
  assign new_n286_ = 45 & ~75;
  assign new_n287_ = ~new_n285_ & ~new_n286_;
  assign new_n288_1_ = new_n284_ & new_n287_;
  assign new_n289_ = ~new_n284_ & ~new_n287_;
  assign n113 = new_n288_1_ | new_n289_;
  assign new_n291_ = \1  & 13;
  assign new_n292_ = ~46 & 76;
  assign new_n293_1_ = 46 & ~76;
  assign new_n294_ = ~new_n292_ & ~new_n293_1_;
  assign new_n295_ = new_n291_ & new_n294_;
  assign new_n296_ = ~new_n291_ & ~new_n294_;
  assign n118 = new_n295_ | new_n296_;
  assign new_n298_1_ = \1  & 14;
  assign new_n299_ = ~47 & 77;
  assign new_n300_ = 47 & ~77;
  assign new_n301_ = ~new_n299_ & ~new_n300_;
  assign new_n302_ = new_n298_1_ & new_n301_;
  assign new_n303_1_ = ~new_n298_1_ & ~new_n301_;
  assign n123 = new_n302_ | new_n303_1_;
  assign new_n305_ = \1  & 15;
  assign new_n306_ = ~48 & 78;
  assign new_n307_ = 48 & ~78;
  assign new_n308_1_ = ~new_n306_ & ~new_n307_;
  assign new_n309_ = new_n305_ & new_n308_1_;
  assign new_n310_ = ~new_n305_ & ~new_n308_1_;
  assign n128 = new_n309_ | new_n310_;
  assign new_n312_ = \1  & 16;
  assign new_n313_1_ = ~49 & 79;
  assign new_n314_ = 49 & ~79;
  assign new_n315_ = ~new_n313_1_ & ~new_n314_;
  assign new_n316_ = new_n312_ & new_n315_;
  assign new_n317_ = ~new_n312_ & ~new_n315_;
  assign n133 = new_n316_ | new_n317_;
  assign new_n319_ = \1  & 17;
  assign new_n320_ = ~50 & 80;
  assign new_n321_ = 50 & ~80;
  assign new_n322_ = ~new_n320_ & ~new_n321_;
  assign new_n323_1_ = new_n319_ & new_n322_;
  assign new_n324_ = ~new_n319_ & ~new_n322_;
  assign n138 = new_n323_1_ | new_n324_;
  assign new_n326_ = \1  & 18;
  assign new_n327_ = ~51 & 81;
  assign new_n328_1_ = 51 & ~81;
  assign new_n329_ = ~new_n327_ & ~new_n328_1_;
  assign new_n330_ = new_n326_ & new_n329_;
  assign new_n331_ = ~new_n326_ & ~new_n329_;
  assign n143 = new_n330_ | new_n331_;
  assign new_n333_1_ = \1  & 19;
  assign new_n334_ = ~52 & 82;
  assign new_n335_ = 52 & ~82;
  assign new_n336_ = ~new_n334_ & ~new_n335_;
  assign new_n337_ = new_n333_1_ & new_n336_;
  assign new_n338_1_ = ~new_n333_1_ & ~new_n336_;
  assign n148 = new_n337_ | new_n338_1_;
  assign new_n340_ = \1  & 20;
  assign new_n341_ = ~53 & 83;
  assign new_n342_ = 53 & ~83;
  assign new_n343_1_ = ~new_n341_ & ~new_n342_;
  assign new_n344_ = new_n340_ & new_n343_1_;
  assign new_n345_ = ~new_n340_ & ~new_n343_1_;
  assign n153 = new_n344_ | new_n345_;
  assign new_n347_ = \1  & 21;
  assign new_n348_1_ = ~54 & 84;
  assign new_n349_ = 54 & ~84;
  assign new_n350_ = ~new_n348_1_ & ~new_n349_;
  assign new_n351_ = new_n347_ & new_n350_;
  assign new_n352_ = ~new_n347_ & ~new_n350_;
  assign n158 = new_n351_ | new_n352_;
  assign new_n354_ = \1  & 22;
  assign new_n355_ = ~55 & 85;
  assign new_n356_ = 55 & ~85;
  assign new_n357_ = ~new_n355_ & ~new_n356_;
  assign new_n358_1_ = new_n354_ & new_n357_;
  assign new_n359_ = ~new_n354_ & ~new_n357_;
  assign n163 = new_n358_1_ | new_n359_;
  assign new_n361_ = \1  & 23;
  assign new_n362_ = ~56 & 86;
  assign new_n363_1_ = 56 & ~86;
  assign new_n364_ = ~new_n362_ & ~new_n363_1_;
  assign new_n365_ = new_n361_ & new_n364_;
  assign new_n366_ = ~new_n361_ & ~new_n364_;
  assign n168 = new_n365_ | new_n366_;
  assign new_n368_1_ = \1  & 24;
  assign new_n369_ = ~57 & 87;
  assign new_n370_ = 57 & ~87;
  assign new_n371_ = ~new_n369_ & ~new_n370_;
  assign new_n372_ = new_n368_1_ & new_n371_;
  assign new_n373_1_ = ~new_n368_1_ & ~new_n371_;
  assign n173 = new_n372_ | new_n373_1_;
  assign new_n375_ = \1  & 25;
  assign new_n376_ = ~58 & 88;
  assign new_n377_ = 58 & ~88;
  assign new_n378_ = ~new_n376_ & ~new_n377_;
  assign new_n379_ = new_n375_ & new_n378_;
  assign new_n380_ = ~new_n375_ & ~new_n378_;
  assign n178 = new_n379_ | new_n380_;
  assign new_n382_ = \1  & 26;
  assign new_n383_ = ~59 & 89;
  assign new_n384_ = 59 & ~89;
  assign new_n385_ = ~new_n383_ & ~new_n384_;
  assign new_n386_ = new_n382_ & new_n385_;
  assign new_n387_ = ~new_n382_ & ~new_n385_;
  assign n183 = new_n386_ | new_n387_;
  assign new_n389_ = \1  & 27;
  assign new_n390_ = ~60 & 90;
  assign new_n391_ = 60 & ~90;
  assign new_n392_ = ~new_n390_ & ~new_n391_;
  assign new_n393_ = new_n389_ & new_n392_;
  assign new_n394_ = ~new_n389_ & ~new_n392_;
  assign n188 = new_n393_ | new_n394_;
  assign new_n396_ = \1  & 28;
  assign new_n397_ = ~61 & 91;
  assign new_n398_ = 61 & ~91;
  assign new_n399_ = ~new_n397_ & ~new_n398_;
  assign new_n400_ = new_n396_ & new_n399_;
  assign new_n401_ = ~new_n396_ & ~new_n399_;
  assign n193 = new_n400_ | new_n401_;
  assign new_n403_ = \1  & 29;
  assign new_n404_ = ~62 & 92;
  assign new_n405_ = 62 & ~92;
  assign new_n406_ = ~new_n404_ & ~new_n405_;
  assign new_n407_ = new_n403_ & new_n406_;
  assign new_n408_ = ~new_n403_ & ~new_n406_;
  assign n198 = new_n407_ | new_n408_;
  assign new_n410_ = \1  & 30;
  assign new_n411_ = ~63 & 93;
  assign new_n412_ = 63 & ~93;
  assign new_n413_ = ~new_n411_ & ~new_n412_;
  assign new_n414_ = new_n410_ & new_n413_;
  assign new_n415_ = ~new_n410_ & ~new_n413_;
  assign n203 = new_n414_ | new_n415_;
  assign new_n417_ = \1  & 31;
  assign new_n418_ = ~64 & 94;
  assign new_n419_ = 64 & ~94;
  assign new_n420_ = ~new_n418_ & ~new_n419_;
  assign new_n421_ = new_n417_ & new_n420_;
  assign new_n422_ = ~new_n417_ & ~new_n420_;
  assign n208 = new_n421_ | new_n422_;
  assign new_n424_ = \1  & 32;
  assign new_n425_ = ~65 & 95;
  assign new_n426_ = 65 & ~95;
  assign new_n427_ = ~new_n425_ & ~new_n426_;
  assign new_n428_ = new_n424_ & new_n427_;
  assign new_n429_ = ~new_n424_ & ~new_n427_;
  assign n213 = new_n428_ | new_n429_;
  assign new_n431_ = \1  & 33;
  assign new_n432_ = ~2 & new_n431_;
  assign new_n433_ = 2 & ~new_n431_;
  assign n218 = new_n432_ | new_n433_;
  assign new_n435_ = 36 & 66;
  assign new_n436_ = 36 & new_n220_;
  assign new_n437_ = 66 & new_n220_;
  assign new_n438_ = ~new_n436_ & ~new_n437_;
  assign n223 = new_n435_ | ~new_n438_;
  assign new_n440_ = 37 & 67;
  assign new_n441_ = 37 & new_n228_1_;
  assign new_n442_ = 67 & new_n228_1_;
  assign new_n443_ = ~new_n441_ & ~new_n442_;
  assign n228 = new_n440_ | ~new_n443_;
  assign new_n445_ = 38 & 68;
  assign new_n446_ = 38 & new_n235_;
  assign new_n447_ = 68 & new_n235_;
  assign new_n448_ = ~new_n446_ & ~new_n447_;
  assign n233 = new_n445_ | ~new_n448_;
  assign new_n450_ = 39 & 69;
  assign new_n451_ = 39 & new_n242_;
  assign new_n452_ = 69 & new_n242_;
  assign new_n453_ = ~new_n451_ & ~new_n452_;
  assign n238 = new_n450_ | ~new_n453_;
  assign new_n455_ = 40 & 70;
  assign new_n456_ = 40 & new_n249_;
  assign new_n457_ = 70 & new_n249_;
  assign new_n458_ = ~new_n456_ & ~new_n457_;
  assign n243 = new_n455_ | ~new_n458_;
  assign new_n460_ = 41 & 71;
  assign new_n461_ = 41 & new_n256_;
  assign new_n462_ = 71 & new_n256_;
  assign new_n463_ = ~new_n461_ & ~new_n462_;
  assign n248 = new_n460_ | ~new_n463_;
  assign new_n465_ = 42 & 72;
  assign new_n466_ = 42 & new_n263_1_;
  assign new_n467_ = 72 & new_n263_1_;
  assign new_n468_ = ~new_n466_ & ~new_n467_;
  assign n253 = new_n465_ | ~new_n468_;
  assign new_n470_ = 43 & 73;
  assign new_n471_ = 43 & new_n270_;
  assign new_n472_ = 73 & new_n270_;
  assign new_n473_ = ~new_n471_ & ~new_n472_;
  assign n258 = new_n470_ | ~new_n473_;
  assign new_n475_ = 44 & 74;
  assign new_n476_ = 44 & new_n277_;
  assign new_n477_ = 74 & new_n277_;
  assign new_n478_ = ~new_n476_ & ~new_n477_;
  assign n263 = new_n475_ | ~new_n478_;
  assign new_n480_ = 45 & 75;
  assign new_n481_ = 45 & new_n284_;
  assign new_n482_ = 75 & new_n284_;
  assign new_n483_ = ~new_n481_ & ~new_n482_;
  assign n268 = new_n480_ | ~new_n483_;
  assign new_n485_ = 46 & 76;
  assign new_n486_ = 46 & new_n291_;
  assign new_n487_ = 76 & new_n291_;
  assign new_n488_ = ~new_n486_ & ~new_n487_;
  assign n273 = new_n485_ | ~new_n488_;
  assign new_n490_ = 47 & 77;
  assign new_n491_ = 47 & new_n298_1_;
  assign new_n492_ = 77 & new_n298_1_;
  assign new_n493_ = ~new_n491_ & ~new_n492_;
  assign n278 = new_n490_ | ~new_n493_;
  assign new_n495_ = 48 & 78;
  assign new_n496_ = 48 & new_n305_;
  assign new_n497_ = 78 & new_n305_;
  assign new_n498_ = ~new_n496_ & ~new_n497_;
  assign n283 = new_n495_ | ~new_n498_;
  assign new_n500_ = 49 & 79;
  assign new_n501_ = 49 & new_n312_;
  assign new_n502_ = 79 & new_n312_;
  assign new_n503_ = ~new_n501_ & ~new_n502_;
  assign n288 = new_n500_ | ~new_n503_;
  assign new_n505_ = 50 & 80;
  assign new_n506_ = 50 & new_n319_;
  assign new_n507_ = 80 & new_n319_;
  assign new_n508_ = ~new_n506_ & ~new_n507_;
  assign n293 = new_n505_ | ~new_n508_;
  assign new_n510_ = 51 & 81;
  assign new_n511_ = 51 & new_n326_;
  assign new_n512_ = 81 & new_n326_;
  assign new_n513_ = ~new_n511_ & ~new_n512_;
  assign n298 = new_n510_ | ~new_n513_;
  assign new_n515_ = 52 & 82;
  assign new_n516_ = 52 & new_n333_1_;
  assign new_n517_ = 82 & new_n333_1_;
  assign new_n518_ = ~new_n516_ & ~new_n517_;
  assign n303 = new_n515_ | ~new_n518_;
  assign new_n520_ = 53 & 83;
  assign new_n521_ = 53 & new_n340_;
  assign new_n522_ = 83 & new_n340_;
  assign new_n523_ = ~new_n521_ & ~new_n522_;
  assign n308 = new_n520_ | ~new_n523_;
  assign new_n525_ = 54 & 84;
  assign new_n526_ = 54 & new_n347_;
  assign new_n527_ = 84 & new_n347_;
  assign new_n528_ = ~new_n526_ & ~new_n527_;
  assign n313 = new_n525_ | ~new_n528_;
  assign new_n530_ = 55 & 85;
  assign new_n531_ = 55 & new_n354_;
  assign new_n532_ = 85 & new_n354_;
  assign new_n533_ = ~new_n531_ & ~new_n532_;
  assign n318 = new_n530_ | ~new_n533_;
  assign new_n535_ = 56 & 86;
  assign new_n536_ = 56 & new_n361_;
  assign new_n537_ = 86 & new_n361_;
  assign new_n538_ = ~new_n536_ & ~new_n537_;
  assign n323 = new_n535_ | ~new_n538_;
  assign new_n540_ = 57 & 87;
  assign new_n541_ = 57 & new_n368_1_;
  assign new_n542_ = 87 & new_n368_1_;
  assign new_n543_ = ~new_n541_ & ~new_n542_;
  assign n328 = new_n540_ | ~new_n543_;
  assign new_n545_ = 58 & 88;
  assign new_n546_ = 58 & new_n375_;
  assign new_n547_ = 88 & new_n375_;
  assign new_n548_ = ~new_n546_ & ~new_n547_;
  assign n333 = new_n545_ | ~new_n548_;
  assign new_n550_ = 59 & 89;
  assign new_n551_ = 59 & new_n382_;
  assign new_n552_ = 89 & new_n382_;
  assign new_n553_ = ~new_n551_ & ~new_n552_;
  assign n338 = new_n550_ | ~new_n553_;
  assign new_n555_ = 60 & 90;
  assign new_n556_ = 60 & new_n389_;
  assign new_n557_ = 90 & new_n389_;
  assign new_n558_ = ~new_n556_ & ~new_n557_;
  assign n343 = new_n555_ | ~new_n558_;
  assign new_n560_ = 61 & 91;
  assign new_n561_ = 61 & new_n396_;
  assign new_n562_ = 91 & new_n396_;
  assign new_n563_ = ~new_n561_ & ~new_n562_;
  assign n348 = new_n560_ | ~new_n563_;
  assign new_n565_ = 62 & 92;
  assign new_n566_ = 62 & new_n403_;
  assign new_n567_ = 92 & new_n403_;
  assign new_n568_ = ~new_n566_ & ~new_n567_;
  assign n353 = new_n565_ | ~new_n568_;
  assign new_n570_ = 63 & 93;
  assign new_n571_ = 63 & new_n410_;
  assign new_n572_ = 93 & new_n410_;
  assign new_n573_ = ~new_n571_ & ~new_n572_;
  assign n358 = new_n570_ | ~new_n573_;
  assign new_n575_ = 64 & 94;
  assign new_n576_ = 64 & new_n417_;
  assign new_n577_ = 94 & new_n417_;
  assign new_n578_ = ~new_n576_ & ~new_n577_;
  assign n363 = new_n575_ | ~new_n578_;
  assign new_n580_ = 65 & 95;
  assign new_n581_ = 65 & new_n424_;
  assign new_n582_ = 95 & new_n424_;
  assign new_n583_ = ~new_n581_ & ~new_n582_;
  assign n368 = new_n580_ | ~new_n583_;
  assign n373 = 2 & new_n431_;
  always @ (posedge clock) begin
    34 <= n68;
    2 <= n73;
    36 <= n78;
    37 <= n83;
    38 <= n88;
    39 <= n93;
    40 <= n98;
    41 <= n103;
    42 <= n108;
    43 <= n113;
    44 <= n118;
    45 <= n123;
    46 <= n128;
    47 <= n133;
    48 <= n138;
    49 <= n143;
    50 <= n148;
    51 <= n153;
    52 <= n158;
    53 <= n163;
    54 <= n168;
    55 <= n173;
    56 <= n178;
    57 <= n183;
    58 <= n188;
    59 <= n193;
    60 <= n198;
    61 <= n203;
    62 <= n208;
    63 <= n213;
    64 <= n218;
    65 <= n223;
    66 <= n228;
    67 <= n233;
    68 <= n238;
    69 <= n243;
    70 <= n248;
    71 <= n253;
    72 <= n258;
    73 <= n263;
    74 <= n268;
    75 <= n273;
    76 <= n278;
    77 <= n283;
    78 <= n288;
    79 <= n293;
    80 <= n298;
    81 <= n303;
    82 <= n308;
    83 <= n313;
    84 <= n318;
    85 <= n323;
    86 <= n328;
    87 <= n333;
    88 <= n338;
    89 <= n343;
    90 <= n348;
    91 <= n353;
    92 <= n358;
    93 <= n363;
    94 <= n368;
    95 <= n373;
  end
  initial begin
    34 <= 1'b0;
    2 <= 1'b0;
    36 <= 1'b0;
    37 <= 1'b0;
    38 <= 1'b0;
    39 <= 1'b0;
    40 <= 1'b0;
    41 <= 1'b0;
    42 <= 1'b0;
    43 <= 1'b0;
    44 <= 1'b0;
    45 <= 1'b0;
    46 <= 1'b0;
    47 <= 1'b0;
    48 <= 1'b0;
    49 <= 1'b0;
    50 <= 1'b0;
    51 <= 1'b0;
    52 <= 1'b0;
    53 <= 1'b0;
    54 <= 1'b0;
    55 <= 1'b0;
    56 <= 1'b0;
    57 <= 1'b0;
    58 <= 1'b0;
    59 <= 1'b0;
    60 <= 1'b0;
    61 <= 1'b0;
    62 <= 1'b0;
    63 <= 1'b0;
    64 <= 1'b0;
    65 <= 1'b0;
    66 <= 1'b0;
    67 <= 1'b0;
    68 <= 1'b0;
    69 <= 1'b0;
    70 <= 1'b0;
    71 <= 1'b0;
    72 <= 1'b0;
    73 <= 1'b0;
    74 <= 1'b0;
    75 <= 1'b0;
    76 <= 1'b0;
    77 <= 1'b0;
    78 <= 1'b0;
    79 <= 1'b0;
    80 <= 1'b0;
    81 <= 1'b0;
    82 <= 1'b0;
    83 <= 1'b0;
    84 <= 1'b0;
    85 <= 1'b0;
    86 <= 1'b0;
    87 <= 1'b0;
    88 <= 1'b0;
    89 <= 1'b0;
    90 <= 1'b0;
    91 <= 1'b0;
    92 <= 1'b0;
    93 <= 1'b0;
    94 <= 1'b0;
    95 <= 1'b0;
  end
endmodule

