module MultiplierA_32 ( clock, 
    \1 , 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20,
    21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34,
    68  );
  input  clock;
  input  \1 , 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18,
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34;
  output 68;
  reg 2, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52,
    53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66;
  wire new_n131_, new_n132_, new_n133_, new_n135_1_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_1_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_1_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_1_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_1_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_1_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_1_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_1_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_1_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_1_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_1_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_1_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_1_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_1_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_1_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_1_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_1_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_1_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_1_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, n70, n75, n80, n85, n90, n95, n100, n105, n110, n115, n120,
    n125, n130, n135, n140, n145, n150, n155, n160, n165, n170, n175, n180,
    n185, n190, n195, n200, n205, n210, n215, n220, n225;
  assign new_n131_ = \1  & 3;
  assign new_n132_ = 36 & ~new_n131_;
  assign new_n133_ = ~36 & new_n131_;
  assign 68 = new_n132_ | new_n133_;
  assign new_n135_1_ = \1  & 34;
  assign new_n136_ = 2 & new_n135_1_;
  assign new_n137_ = 36 & new_n131_;
  assign new_n138_ = \1  & 4;
  assign new_n139_ = ~new_n137_ & ~new_n138_;
  assign new_n140_1_ = 37 & ~new_n139_;
  assign new_n141_ = new_n137_ & new_n138_;
  assign new_n142_ = ~new_n140_1_ & ~new_n141_;
  assign new_n143_ = \1  & 5;
  assign new_n144_ = new_n142_ & ~new_n143_;
  assign new_n145_1_ = 38 & ~new_n144_;
  assign new_n146_ = ~new_n142_ & new_n143_;
  assign new_n147_ = ~new_n145_1_ & ~new_n146_;
  assign new_n148_ = \1  & 6;
  assign new_n149_ = new_n147_ & ~new_n148_;
  assign new_n150_1_ = 39 & ~new_n149_;
  assign new_n151_ = ~new_n147_ & new_n148_;
  assign new_n152_ = ~new_n150_1_ & ~new_n151_;
  assign new_n153_ = \1  & 7;
  assign new_n154_ = new_n152_ & ~new_n153_;
  assign new_n155_1_ = 40 & ~new_n154_;
  assign new_n156_ = ~new_n152_ & new_n153_;
  assign new_n157_ = ~new_n155_1_ & ~new_n156_;
  assign new_n158_ = \1  & 8;
  assign new_n159_ = new_n157_ & ~new_n158_;
  assign new_n160_1_ = 41 & ~new_n159_;
  assign new_n161_ = ~new_n157_ & new_n158_;
  assign new_n162_ = ~new_n160_1_ & ~new_n161_;
  assign new_n163_ = \1  & 9;
  assign new_n164_ = new_n162_ & ~new_n163_;
  assign new_n165_1_ = 42 & ~new_n164_;
  assign new_n166_ = ~new_n162_ & new_n163_;
  assign new_n167_ = ~new_n165_1_ & ~new_n166_;
  assign new_n168_ = \1  & 10;
  assign new_n169_ = new_n167_ & ~new_n168_;
  assign new_n170_1_ = 43 & ~new_n169_;
  assign new_n171_ = ~new_n167_ & new_n168_;
  assign new_n172_ = ~new_n170_1_ & ~new_n171_;
  assign new_n173_ = \1  & 11;
  assign new_n174_ = new_n172_ & ~new_n173_;
  assign new_n175_1_ = 44 & ~new_n174_;
  assign new_n176_ = ~new_n172_ & new_n173_;
  assign new_n177_ = ~new_n175_1_ & ~new_n176_;
  assign new_n178_ = \1  & 12;
  assign new_n179_ = new_n177_ & ~new_n178_;
  assign new_n180_1_ = 45 & ~new_n179_;
  assign new_n181_ = ~new_n177_ & new_n178_;
  assign new_n182_ = ~new_n180_1_ & ~new_n181_;
  assign new_n183_ = \1  & 13;
  assign new_n184_ = new_n182_ & ~new_n183_;
  assign new_n185_1_ = 46 & ~new_n184_;
  assign new_n186_ = ~new_n182_ & new_n183_;
  assign new_n187_ = ~new_n185_1_ & ~new_n186_;
  assign new_n188_ = \1  & 14;
  assign new_n189_ = new_n187_ & ~new_n188_;
  assign new_n190_1_ = 47 & ~new_n189_;
  assign new_n191_ = ~new_n187_ & new_n188_;
  assign new_n192_ = ~new_n190_1_ & ~new_n191_;
  assign new_n193_ = \1  & 15;
  assign new_n194_ = new_n192_ & ~new_n193_;
  assign new_n195_1_ = 48 & ~new_n194_;
  assign new_n196_ = ~new_n192_ & new_n193_;
  assign new_n197_ = ~new_n195_1_ & ~new_n196_;
  assign new_n198_ = \1  & 16;
  assign new_n199_ = new_n197_ & ~new_n198_;
  assign new_n200_1_ = 49 & ~new_n199_;
  assign new_n201_ = ~new_n197_ & new_n198_;
  assign new_n202_ = ~new_n200_1_ & ~new_n201_;
  assign new_n203_ = \1  & 17;
  assign new_n204_ = new_n202_ & ~new_n203_;
  assign new_n205_1_ = 50 & ~new_n204_;
  assign new_n206_ = ~new_n202_ & new_n203_;
  assign new_n207_ = ~new_n205_1_ & ~new_n206_;
  assign new_n208_ = \1  & 18;
  assign new_n209_ = new_n207_ & ~new_n208_;
  assign new_n210_1_ = 51 & ~new_n209_;
  assign new_n211_ = ~new_n207_ & new_n208_;
  assign new_n212_ = ~new_n210_1_ & ~new_n211_;
  assign new_n213_ = \1  & 19;
  assign new_n214_ = new_n212_ & ~new_n213_;
  assign new_n215_1_ = 52 & ~new_n214_;
  assign new_n216_ = ~new_n212_ & new_n213_;
  assign new_n217_ = ~new_n215_1_ & ~new_n216_;
  assign new_n218_ = \1  & 20;
  assign new_n219_ = new_n217_ & ~new_n218_;
  assign new_n220_1_ = 53 & ~new_n219_;
  assign new_n221_ = ~new_n217_ & new_n218_;
  assign new_n222_ = ~new_n220_1_ & ~new_n221_;
  assign new_n223_ = \1  & 21;
  assign new_n224_ = new_n222_ & ~new_n223_;
  assign new_n225_1_ = 54 & ~new_n224_;
  assign new_n226_ = ~new_n222_ & new_n223_;
  assign new_n227_ = ~new_n225_1_ & ~new_n226_;
  assign new_n228_ = \1  & 22;
  assign new_n229_ = new_n227_ & ~new_n228_;
  assign new_n230_ = 55 & ~new_n229_;
  assign new_n231_ = ~new_n227_ & new_n228_;
  assign new_n232_ = ~new_n230_ & ~new_n231_;
  assign new_n233_ = \1  & 23;
  assign new_n234_ = new_n232_ & ~new_n233_;
  assign new_n235_ = 56 & ~new_n234_;
  assign new_n236_ = ~new_n232_ & new_n233_;
  assign new_n237_ = ~new_n235_ & ~new_n236_;
  assign new_n238_ = \1  & 24;
  assign new_n239_ = new_n237_ & ~new_n238_;
  assign new_n240_ = 57 & ~new_n239_;
  assign new_n241_ = ~new_n237_ & new_n238_;
  assign new_n242_ = ~new_n240_ & ~new_n241_;
  assign new_n243_ = \1  & 25;
  assign new_n244_ = new_n242_ & ~new_n243_;
  assign new_n245_ = 58 & ~new_n244_;
  assign new_n246_ = ~new_n242_ & new_n243_;
  assign new_n247_ = ~new_n245_ & ~new_n246_;
  assign new_n248_ = \1  & 26;
  assign new_n249_ = new_n247_ & ~new_n248_;
  assign new_n250_ = 59 & ~new_n249_;
  assign new_n251_ = ~new_n247_ & new_n248_;
  assign new_n252_ = ~new_n250_ & ~new_n251_;
  assign new_n253_ = \1  & 27;
  assign new_n254_ = new_n252_ & ~new_n253_;
  assign new_n255_ = 60 & ~new_n254_;
  assign new_n256_ = ~new_n252_ & new_n253_;
  assign new_n257_ = ~new_n255_ & ~new_n256_;
  assign new_n258_ = \1  & 28;
  assign new_n259_ = new_n257_ & ~new_n258_;
  assign new_n260_ = 61 & ~new_n259_;
  assign new_n261_ = ~new_n257_ & new_n258_;
  assign new_n262_ = ~new_n260_ & ~new_n261_;
  assign new_n263_ = \1  & 29;
  assign new_n264_ = new_n262_ & ~new_n263_;
  assign new_n265_ = 62 & ~new_n264_;
  assign new_n266_ = ~new_n262_ & new_n263_;
  assign new_n267_ = ~new_n265_ & ~new_n266_;
  assign new_n268_ = \1  & 30;
  assign new_n269_ = new_n267_ & ~new_n268_;
  assign new_n270_ = 63 & ~new_n269_;
  assign new_n271_ = ~new_n267_ & new_n268_;
  assign new_n272_ = ~new_n270_ & ~new_n271_;
  assign new_n273_ = \1  & 31;
  assign new_n274_ = new_n272_ & ~new_n273_;
  assign new_n275_ = 64 & ~new_n274_;
  assign new_n276_ = ~new_n272_ & new_n273_;
  assign new_n277_ = ~new_n275_ & ~new_n276_;
  assign new_n278_ = \1  & 32;
  assign new_n279_ = new_n277_ & ~new_n278_;
  assign new_n280_ = 65 & ~new_n279_;
  assign new_n281_ = ~new_n277_ & new_n278_;
  assign new_n282_ = ~new_n280_ & ~new_n281_;
  assign new_n283_ = \1  & 33;
  assign new_n284_ = new_n282_ & ~new_n283_;
  assign new_n285_ = 66 & ~new_n284_;
  assign new_n286_ = ~new_n282_ & new_n283_;
  assign new_n287_ = ~new_n285_ & ~new_n286_;
  assign new_n288_ = new_n136_ & new_n287_;
  assign new_n289_ = 2 & ~new_n135_1_;
  assign new_n290_ = ~new_n287_ & new_n289_;
  assign new_n291_ = ~new_n288_ & ~new_n290_;
  assign new_n292_ = ~2 & new_n135_1_;
  assign new_n293_ = ~new_n287_ & new_n292_;
  assign new_n294_ = new_n136_ & ~new_n287_;
  assign new_n295_ = ~new_n293_ & ~new_n294_;
  assign n70 = ~new_n291_ | ~new_n295_;
  assign new_n297_ = ~new_n139_ & ~new_n141_;
  assign new_n298_ = 37 & ~new_n297_;
  assign new_n299_ = ~new_n137_ & new_n138_;
  assign new_n300_ = new_n137_ & ~new_n138_;
  assign new_n301_ = ~new_n299_ & ~new_n300_;
  assign new_n302_ = ~37 & ~new_n301_;
  assign n75 = new_n298_ | new_n302_;
  assign new_n304_ = ~new_n144_ & ~new_n146_;
  assign new_n305_ = 38 & ~new_n304_;
  assign new_n306_ = new_n142_ & new_n143_;
  assign new_n307_ = ~new_n142_ & ~new_n143_;
  assign new_n308_ = ~new_n306_ & ~new_n307_;
  assign new_n309_ = ~38 & ~new_n308_;
  assign n80 = new_n305_ | new_n309_;
  assign new_n311_ = ~new_n149_ & ~new_n151_;
  assign new_n312_ = 39 & ~new_n311_;
  assign new_n313_ = new_n147_ & new_n148_;
  assign new_n314_ = ~new_n147_ & ~new_n148_;
  assign new_n315_ = ~new_n313_ & ~new_n314_;
  assign new_n316_ = ~39 & ~new_n315_;
  assign n85 = new_n312_ | new_n316_;
  assign new_n318_ = ~new_n154_ & ~new_n156_;
  assign new_n319_ = 40 & ~new_n318_;
  assign new_n320_ = new_n152_ & new_n153_;
  assign new_n321_ = ~new_n152_ & ~new_n153_;
  assign new_n322_ = ~new_n320_ & ~new_n321_;
  assign new_n323_ = ~40 & ~new_n322_;
  assign n90 = new_n319_ | new_n323_;
  assign new_n325_ = ~new_n159_ & ~new_n161_;
  assign new_n326_ = 41 & ~new_n325_;
  assign new_n327_ = new_n157_ & new_n158_;
  assign new_n328_ = ~new_n157_ & ~new_n158_;
  assign new_n329_ = ~new_n327_ & ~new_n328_;
  assign new_n330_ = ~41 & ~new_n329_;
  assign n95 = new_n326_ | new_n330_;
  assign new_n332_ = ~new_n164_ & ~new_n166_;
  assign new_n333_ = 42 & ~new_n332_;
  assign new_n334_ = new_n162_ & new_n163_;
  assign new_n335_ = ~new_n162_ & ~new_n163_;
  assign new_n336_ = ~new_n334_ & ~new_n335_;
  assign new_n337_ = ~42 & ~new_n336_;
  assign n100 = new_n333_ | new_n337_;
  assign new_n339_ = ~new_n169_ & ~new_n171_;
  assign new_n340_ = 43 & ~new_n339_;
  assign new_n341_ = new_n167_ & new_n168_;
  assign new_n342_ = ~new_n167_ & ~new_n168_;
  assign new_n343_ = ~new_n341_ & ~new_n342_;
  assign new_n344_ = ~43 & ~new_n343_;
  assign n105 = new_n340_ | new_n344_;
  assign new_n346_ = ~new_n174_ & ~new_n176_;
  assign new_n347_ = 44 & ~new_n346_;
  assign new_n348_ = new_n172_ & new_n173_;
  assign new_n349_ = ~new_n172_ & ~new_n173_;
  assign new_n350_ = ~new_n348_ & ~new_n349_;
  assign new_n351_ = ~44 & ~new_n350_;
  assign n110 = new_n347_ | new_n351_;
  assign new_n353_ = ~new_n179_ & ~new_n181_;
  assign new_n354_ = 45 & ~new_n353_;
  assign new_n355_ = new_n177_ & new_n178_;
  assign new_n356_ = ~new_n177_ & ~new_n178_;
  assign new_n357_ = ~new_n355_ & ~new_n356_;
  assign new_n358_ = ~45 & ~new_n357_;
  assign n115 = new_n354_ | new_n358_;
  assign new_n360_ = ~new_n184_ & ~new_n186_;
  assign new_n361_ = 46 & ~new_n360_;
  assign new_n362_ = new_n182_ & new_n183_;
  assign new_n363_ = ~new_n182_ & ~new_n183_;
  assign new_n364_ = ~new_n362_ & ~new_n363_;
  assign new_n365_ = ~46 & ~new_n364_;
  assign n120 = new_n361_ | new_n365_;
  assign new_n367_ = ~new_n189_ & ~new_n191_;
  assign new_n368_ = 47 & ~new_n367_;
  assign new_n369_ = new_n187_ & new_n188_;
  assign new_n370_ = ~new_n187_ & ~new_n188_;
  assign new_n371_ = ~new_n369_ & ~new_n370_;
  assign new_n372_ = ~47 & ~new_n371_;
  assign n125 = new_n368_ | new_n372_;
  assign new_n374_ = ~new_n194_ & ~new_n196_;
  assign new_n375_ = 48 & ~new_n374_;
  assign new_n376_ = new_n192_ & new_n193_;
  assign new_n377_ = ~new_n192_ & ~new_n193_;
  assign new_n378_ = ~new_n376_ & ~new_n377_;
  assign new_n379_ = ~48 & ~new_n378_;
  assign n130 = new_n375_ | new_n379_;
  assign new_n381_ = ~new_n199_ & ~new_n201_;
  assign new_n382_ = 49 & ~new_n381_;
  assign new_n383_ = new_n197_ & new_n198_;
  assign new_n384_ = ~new_n197_ & ~new_n198_;
  assign new_n385_ = ~new_n383_ & ~new_n384_;
  assign new_n386_ = ~49 & ~new_n385_;
  assign n135 = new_n382_ | new_n386_;
  assign new_n388_ = ~new_n204_ & ~new_n206_;
  assign new_n389_ = 50 & ~new_n388_;
  assign new_n390_ = new_n202_ & new_n203_;
  assign new_n391_ = ~new_n202_ & ~new_n203_;
  assign new_n392_ = ~new_n390_ & ~new_n391_;
  assign new_n393_ = ~50 & ~new_n392_;
  assign n140 = new_n389_ | new_n393_;
  assign new_n395_ = ~new_n209_ & ~new_n211_;
  assign new_n396_ = 51 & ~new_n395_;
  assign new_n397_ = new_n207_ & new_n208_;
  assign new_n398_ = ~new_n207_ & ~new_n208_;
  assign new_n399_ = ~new_n397_ & ~new_n398_;
  assign new_n400_ = ~51 & ~new_n399_;
  assign n145 = new_n396_ | new_n400_;
  assign new_n402_ = ~new_n214_ & ~new_n216_;
  assign new_n403_ = 52 & ~new_n402_;
  assign new_n404_ = new_n212_ & new_n213_;
  assign new_n405_ = ~new_n212_ & ~new_n213_;
  assign new_n406_ = ~new_n404_ & ~new_n405_;
  assign new_n407_ = ~52 & ~new_n406_;
  assign n150 = new_n403_ | new_n407_;
  assign new_n409_ = ~new_n219_ & ~new_n221_;
  assign new_n410_ = 53 & ~new_n409_;
  assign new_n411_ = new_n217_ & new_n218_;
  assign new_n412_ = ~new_n217_ & ~new_n218_;
  assign new_n413_ = ~new_n411_ & ~new_n412_;
  assign new_n414_ = ~53 & ~new_n413_;
  assign n155 = new_n410_ | new_n414_;
  assign new_n416_ = ~new_n224_ & ~new_n226_;
  assign new_n417_ = 54 & ~new_n416_;
  assign new_n418_ = new_n222_ & new_n223_;
  assign new_n419_ = ~new_n222_ & ~new_n223_;
  assign new_n420_ = ~new_n418_ & ~new_n419_;
  assign new_n421_ = ~54 & ~new_n420_;
  assign n160 = new_n417_ | new_n421_;
  assign new_n423_ = ~new_n229_ & ~new_n231_;
  assign new_n424_ = 55 & ~new_n423_;
  assign new_n425_ = new_n227_ & new_n228_;
  assign new_n426_ = ~new_n227_ & ~new_n228_;
  assign new_n427_ = ~new_n425_ & ~new_n426_;
  assign new_n428_ = ~55 & ~new_n427_;
  assign n165 = new_n424_ | new_n428_;
  assign new_n430_ = ~new_n234_ & ~new_n236_;
  assign new_n431_ = 56 & ~new_n430_;
  assign new_n432_ = new_n232_ & new_n233_;
  assign new_n433_ = ~new_n232_ & ~new_n233_;
  assign new_n434_ = ~new_n432_ & ~new_n433_;
  assign new_n435_ = ~56 & ~new_n434_;
  assign n170 = new_n431_ | new_n435_;
  assign new_n437_ = ~new_n239_ & ~new_n241_;
  assign new_n438_ = 57 & ~new_n437_;
  assign new_n439_ = new_n237_ & new_n238_;
  assign new_n440_ = ~new_n237_ & ~new_n238_;
  assign new_n441_ = ~new_n439_ & ~new_n440_;
  assign new_n442_ = ~57 & ~new_n441_;
  assign n175 = new_n438_ | new_n442_;
  assign new_n444_ = ~new_n244_ & ~new_n246_;
  assign new_n445_ = 58 & ~new_n444_;
  assign new_n446_ = new_n242_ & new_n243_;
  assign new_n447_ = ~new_n242_ & ~new_n243_;
  assign new_n448_ = ~new_n446_ & ~new_n447_;
  assign new_n449_ = ~58 & ~new_n448_;
  assign n180 = new_n445_ | new_n449_;
  assign new_n451_ = ~new_n249_ & ~new_n251_;
  assign new_n452_ = 59 & ~new_n451_;
  assign new_n453_ = new_n247_ & new_n248_;
  assign new_n454_ = ~new_n247_ & ~new_n248_;
  assign new_n455_ = ~new_n453_ & ~new_n454_;
  assign new_n456_ = ~59 & ~new_n455_;
  assign n185 = new_n452_ | new_n456_;
  assign new_n458_ = ~new_n254_ & ~new_n256_;
  assign new_n459_ = 60 & ~new_n458_;
  assign new_n460_ = new_n252_ & new_n253_;
  assign new_n461_ = ~new_n252_ & ~new_n253_;
  assign new_n462_ = ~new_n460_ & ~new_n461_;
  assign new_n463_ = ~60 & ~new_n462_;
  assign n190 = new_n459_ | new_n463_;
  assign new_n465_ = ~new_n259_ & ~new_n261_;
  assign new_n466_ = 61 & ~new_n465_;
  assign new_n467_ = new_n257_ & new_n258_;
  assign new_n468_ = ~new_n257_ & ~new_n258_;
  assign new_n469_ = ~new_n467_ & ~new_n468_;
  assign new_n470_ = ~61 & ~new_n469_;
  assign n195 = new_n466_ | new_n470_;
  assign new_n472_ = ~new_n264_ & ~new_n266_;
  assign new_n473_ = 62 & ~new_n472_;
  assign new_n474_ = new_n262_ & new_n263_;
  assign new_n475_ = ~new_n262_ & ~new_n263_;
  assign new_n476_ = ~new_n474_ & ~new_n475_;
  assign new_n477_ = ~62 & ~new_n476_;
  assign n200 = new_n473_ | new_n477_;
  assign new_n479_ = ~new_n269_ & ~new_n271_;
  assign new_n480_ = 63 & ~new_n479_;
  assign new_n481_ = new_n267_ & new_n268_;
  assign new_n482_ = ~new_n267_ & ~new_n268_;
  assign new_n483_ = ~new_n481_ & ~new_n482_;
  assign new_n484_ = ~63 & ~new_n483_;
  assign n205 = new_n480_ | new_n484_;
  assign new_n486_ = ~new_n274_ & ~new_n276_;
  assign new_n487_ = 64 & ~new_n486_;
  assign new_n488_ = new_n272_ & new_n273_;
  assign new_n489_ = ~new_n272_ & ~new_n273_;
  assign new_n490_ = ~new_n488_ & ~new_n489_;
  assign new_n491_ = ~64 & ~new_n490_;
  assign n210 = new_n487_ | new_n491_;
  assign new_n493_ = ~new_n279_ & ~new_n281_;
  assign new_n494_ = 65 & ~new_n493_;
  assign new_n495_ = new_n277_ & new_n278_;
  assign new_n496_ = ~new_n277_ & ~new_n278_;
  assign new_n497_ = ~new_n495_ & ~new_n496_;
  assign new_n498_ = ~65 & ~new_n497_;
  assign n215 = new_n494_ | new_n498_;
  assign new_n500_ = ~new_n284_ & ~new_n286_;
  assign new_n501_ = 66 & ~new_n500_;
  assign new_n502_ = new_n282_ & new_n283_;
  assign new_n503_ = ~new_n282_ & ~new_n283_;
  assign new_n504_ = ~new_n502_ & ~new_n503_;
  assign new_n505_ = ~66 & ~new_n504_;
  assign n220 = new_n501_ | new_n505_;
  assign new_n507_ = ~new_n135_1_ & ~new_n287_;
  assign new_n508_ = new_n135_1_ & new_n287_;
  assign new_n509_ = ~new_n507_ & ~new_n508_;
  assign new_n510_ = 2 & new_n509_;
  assign new_n511_ = ~2 & ~new_n509_;
  assign n225 = new_n510_ | new_n511_;
  always @ (posedge clock) begin
    2 <= n70;
    36 <= n75;
    37 <= n80;
    38 <= n85;
    39 <= n90;
    40 <= n95;
    41 <= n100;
    42 <= n105;
    43 <= n110;
    44 <= n115;
    45 <= n120;
    46 <= n125;
    47 <= n130;
    48 <= n135;
    49 <= n140;
    50 <= n145;
    51 <= n150;
    52 <= n155;
    53 <= n160;
    54 <= n165;
    55 <= n170;
    56 <= n175;
    57 <= n180;
    58 <= n185;
    59 <= n190;
    60 <= n195;
    61 <= n200;
    62 <= n205;
    63 <= n210;
    64 <= n215;
    65 <= n220;
    66 <= n225;
  end
  initial begin
    2 <= 1'b0;
    36 <= 1'b0;
    37 <= 1'b0;
    38 <= 1'b0;
    39 <= 1'b0;
    40 <= 1'b0;
    41 <= 1'b0;
    42 <= 1'b0;
    43 <= 1'b0;
    44 <= 1'b0;
    45 <= 1'b0;
    46 <= 1'b0;
    47 <= 1'b0;
    48 <= 1'b0;
    49 <= 1'b0;
    50 <= 1'b0;
    51 <= 1'b0;
    52 <= 1'b0;
    53 <= 1'b0;
    54 <= 1'b0;
    55 <= 1'b0;
    56 <= 1'b0;
    57 <= 1'b0;
    58 <= 1'b0;
    59 <= 1'b0;
    60 <= 1'b0;
    61 <= 1'b0;
    62 <= 1'b0;
    63 <= 1'b0;
    64 <= 1'b0;
    65 <= 1'b0;
    66 <= 1'b0;
  end
endmodule

