// Benchmark "testing" written by ABC on Thu Oct  8 22:16:58 2020

module testing ( 
    A2777, A2776, A2775, A2774, A2773, A2744, A2743, A2742, A2741, A2740,
    A2711, A2710, A2709, A2708, A2707, A2678, A2677, A2676, A2675, A2674,
    A2645, A2644, A2643, A2642, A2641, A2612, A2611, A2610, A2609, A2608,
    A2579, A2578, A2577, A2576, A2575, A2546, A2545, A2544, A2543, A2542,
    A2513, A2512, A2511, A2510, A2509, A2480, A2479, A2478, A2477, A2476,
    A2447, A2446, A2445, A2444, A2443, A2414, A2413, A2412, A2411, A2410,
    A2381, A2380, A2379, A2378, A2377, A2348, A2347, A2346, A2345, A2344,
    A2315, A2314, A2313, A2312, A2311, A2282, A2281, A2280, A2279, A2278,
    A2249, A2248, A2247, A2246, A2245, A2216, A2215, A2214, A2213, A2212,
    A2183, A2182, A2181, A2180, A2179, A2150, A2149, A2148, A2147, A2146,
    A2117, A2116, A2115, A2114, A2113, A2084, A2083, A2082, A2081, A2080,
    A2051, A2050, A2049, A2048, A2047, A2018, A2017, A2016, A2015, A2014,
    A1981, A1982, A1983, A1984, A1985,
    A1132, A1131, A1130, A1129, A1128, A1099, A1098, A1097, A1096, A1095,
    A1066, A1065, A1064, A1063, A1062, A1033, A1032, A1031, A1030, A1029,
    A1000, A999, A998, A997, A996, A967, A966, A965, A964, A963, A934,
    A933, A932, A931, A930, A901, A900, A899, A898, A897, A868, A867, A866,
    A865, A864, A835, A834, A833, A832, A831, A802, A801, A800, A799, A798,
    A769, A768, A767, A766, A765, A736, A735, A734, A733, A732, A703, A702,
    A701, A700, A699, A670, A669, A668, A667, A666, A637, A636, A635, A634,
    A633, A604, A603, A602, A601, A600, A571, A570, A569, A568, A567, A538,
    A537, A536, A535, A534, A505, A504, A503, A502, A501, A472, A471, A470,
    A469, A468, A439, A438, A437, A436, A435, A406, A405, A404, A403, A402,
    A373, A372, A371, A370, A369, A336, A337, A338, A339, A340  );
  input  A2777, A2776, A2775, A2774, A2773, A2744, A2743, A2742, A2741,
    A2740, A2711, A2710, A2709, A2708, A2707, A2678, A2677, A2676, A2675,
    A2674, A2645, A2644, A2643, A2642, A2641, A2612, A2611, A2610, A2609,
    A2608, A2579, A2578, A2577, A2576, A2575, A2546, A2545, A2544, A2543,
    A2542, A2513, A2512, A2511, A2510, A2509, A2480, A2479, A2478, A2477,
    A2476, A2447, A2446, A2445, A2444, A2443, A2414, A2413, A2412, A2411,
    A2410, A2381, A2380, A2379, A2378, A2377, A2348, A2347, A2346, A2345,
    A2344, A2315, A2314, A2313, A2312, A2311, A2282, A2281, A2280, A2279,
    A2278, A2249, A2248, A2247, A2246, A2245, A2216, A2215, A2214, A2213,
    A2212, A2183, A2182, A2181, A2180, A2179, A2150, A2149, A2148, A2147,
    A2146, A2117, A2116, A2115, A2114, A2113, A2084, A2083, A2082, A2081,
    A2080, A2051, A2050, A2049, A2048, A2047, A2018, A2017, A2016, A2015,
    A2014, A1981, A1982, A1983, A1984, A1985;
  output A1132, A1131, A1130, A1129, A1128, A1099, A1098, A1097, A1096, A1095,
    A1066, A1065, A1064, A1063, A1062, A1033, A1032, A1031, A1030, A1029,
    A1000, A999, A998, A997, A996, A967, A966, A965, A964, A963, A934,
    A933, A932, A931, A930, A901, A900, A899, A898, A897, A868, A867, A866,
    A865, A864, A835, A834, A833, A832, A831, A802, A801, A800, A799, A798,
    A769, A768, A767, A766, A765, A736, A735, A734, A733, A732, A703, A702,
    A701, A700, A699, A670, A669, A668, A667, A666, A637, A636, A635, A634,
    A633, A604, A603, A602, A601, A600, A571, A570, A569, A568, A567, A538,
    A537, A536, A535, A534, A505, A504, A503, A502, A501, A472, A471, A470,
    A469, A468, A439, A438, A437, A436, A435, A406, A405, A404, A403, A402,
    A373, A372, A371, A370, A369, A336, A337, A338, A339, A340;
  wire new_A2013_, new_A2012_, new_A2011_, new_A2010_, new_A2009_,
    new_A2008_, new_A2007_, new_A2006_, new_A2005_, new_A2004_, new_A2003_,
    new_A2002_, new_A2001_, new_A2000_, new_A1999_, new_A1998_, new_A1997_,
    new_A1996_, new_A1995_, new_A1994_, new_A1993_, new_A1992_, new_A1991_,
    new_A1990_, new_A1989_, new_A1988_, new_A1987_, new_A1986_, new_A2019_,
    new_A2020_, new_A2021_, new_A2022_, new_A2023_, new_A2024_, new_A2025_,
    new_A2026_, new_A2027_, new_A2028_, new_A2029_, new_A2030_, new_A2031_,
    new_A2032_, new_A2033_, new_A2034_, new_A2035_, new_A2036_, new_A2037_,
    new_A2038_, new_A2039_, new_A2040_, new_A2041_, new_A2042_, new_A2043_,
    new_A2044_, new_A2045_, new_A2046_, new_A2052_, new_A2053_, new_A2054_,
    new_A2055_, new_A2056_, new_A2057_, new_A2058_, new_A2059_, new_A2060_,
    new_A2061_, new_A2062_, new_A2063_, new_A2064_, new_A2065_, new_A2066_,
    new_A2067_, new_A2068_, new_A2069_, new_A2070_, new_A2071_, new_A2072_,
    new_A2073_, new_A2074_, new_A2075_, new_A2076_, new_A2077_, new_A2078_,
    new_A2079_, new_A2085_, new_A2086_, new_A2087_, new_A2088_, new_A2089_,
    new_A2090_, new_A2091_, new_A2092_, new_A2093_, new_A2094_, new_A2095_,
    new_A2096_, new_A2097_, new_A2098_, new_A2099_, new_A2100_, new_A2101_,
    new_A2102_, new_A2103_, new_A2104_, new_A2105_, new_A2106_, new_A2107_,
    new_A2108_, new_A2109_, new_A2110_, new_A2111_, new_A2112_, new_A2118_,
    new_A2119_, new_A2120_, new_A2121_, new_A2122_, new_A2123_, new_A2124_,
    new_A2125_, new_A2126_, new_A2127_, new_A2128_, new_A2129_, new_A2130_,
    new_A2131_, new_A2132_, new_A2133_, new_A2134_, new_A2135_, new_A2136_,
    new_A2137_, new_A2138_, new_A2139_, new_A2140_, new_A2141_, new_A2142_,
    new_A2143_, new_A2144_, new_A2145_, new_A2151_, new_A2152_, new_A2153_,
    new_A2154_, new_A2155_, new_A2156_, new_A2157_, new_A2158_, new_A2159_,
    new_A2160_, new_A2161_, new_A2162_, new_A2163_, new_A2164_, new_A2165_,
    new_A2166_, new_A2167_, new_A2168_, new_A2169_, new_A2170_, new_A2171_,
    new_A2172_, new_A2173_, new_A2174_, new_A2175_, new_A2176_, new_A2177_,
    new_A2178_, new_A2184_, new_A2185_, new_A2186_, new_A2187_, new_A2188_,
    new_A2189_, new_A2190_, new_A2191_, new_A2192_, new_A2193_, new_A2194_,
    new_A2195_, new_A2196_, new_A2197_, new_A2198_, new_A2199_, new_A2200_,
    new_A2201_, new_A2202_, new_A2203_, new_A2204_, new_A2205_, new_A2206_,
    new_A2207_, new_A2208_, new_A2209_, new_A2210_, new_A2211_, new_A2217_,
    new_A2218_, new_A2219_, new_A2220_, new_A2221_, new_A2222_, new_A2223_,
    new_A2224_, new_A2225_, new_A2226_, new_A2227_, new_A2228_, new_A2229_,
    new_A2230_, new_A2231_, new_A2232_, new_A2233_, new_A2234_, new_A2235_,
    new_A2236_, new_A2237_, new_A2238_, new_A2239_, new_A2240_, new_A2241_,
    new_A2242_, new_A2243_, new_A2244_, new_A2250_, new_A2251_, new_A2252_,
    new_A2253_, new_A2254_, new_A2255_, new_A2256_, new_A2257_, new_A2258_,
    new_A2259_, new_A2260_, new_A2261_, new_A2262_, new_A2263_, new_A2264_,
    new_A2265_, new_A2266_, new_A2267_, new_A2268_, new_A2269_, new_A2270_,
    new_A2271_, new_A2272_, new_A2273_, new_A2274_, new_A2275_, new_A2276_,
    new_A2277_, new_A2283_, new_A2284_, new_A2285_, new_A2286_, new_A2287_,
    new_A2288_, new_A2289_, new_A2290_, new_A2291_, new_A2292_, new_A2293_,
    new_A2294_, new_A2295_, new_A2296_, new_A2297_, new_A2298_, new_A2299_,
    new_A2300_, new_A2301_, new_A2302_, new_A2303_, new_A2304_, new_A2305_,
    new_A2306_, new_A2307_, new_A2308_, new_A2309_, new_A2310_, new_A2316_,
    new_A2317_, new_A2318_, new_A2319_, new_A2320_, new_A2321_, new_A2322_,
    new_A2323_, new_A2324_, new_A2325_, new_A2326_, new_A2327_, new_A2328_,
    new_A2329_, new_A2330_, new_A2331_, new_A2332_, new_A2333_, new_A2334_,
    new_A2335_, new_A2336_, new_A2337_, new_A2338_, new_A2339_, new_A2340_,
    new_A2341_, new_A2342_, new_A2343_, new_A2349_, new_A2350_, new_A2351_,
    new_A2352_, new_A2353_, new_A2354_, new_A2355_, new_A2356_, new_A2357_,
    new_A2358_, new_A2359_, new_A2360_, new_A2361_, new_A2362_, new_A2363_,
    new_A2364_, new_A2365_, new_A2366_, new_A2367_, new_A2368_, new_A2369_,
    new_A2370_, new_A2371_, new_A2372_, new_A2373_, new_A2374_, new_A2375_,
    new_A2376_, new_A2382_, new_A2383_, new_A2384_, new_A2385_, new_A2386_,
    new_A2387_, new_A2388_, new_A2389_, new_A2390_, new_A2391_, new_A2392_,
    new_A2393_, new_A2394_, new_A2395_, new_A2396_, new_A2397_, new_A2398_,
    new_A2399_, new_A2400_, new_A2401_, new_A2402_, new_A2403_, new_A2404_,
    new_A2405_, new_A2406_, new_A2407_, new_A2408_, new_A2409_, new_A2415_,
    new_A2416_, new_A2417_, new_A2418_, new_A2419_, new_A2420_, new_A2421_,
    new_A2422_, new_A2423_, new_A2424_, new_A2425_, new_A2426_, new_A2427_,
    new_A2428_, new_A2429_, new_A2430_, new_A2431_, new_A2432_, new_A2433_,
    new_A2434_, new_A2435_, new_A2436_, new_A2437_, new_A2438_, new_A2439_,
    new_A2440_, new_A2441_, new_A2442_, new_A2448_, new_A2449_, new_A2450_,
    new_A2451_, new_A2452_, new_A2453_, new_A2454_, new_A2455_, new_A2456_,
    new_A2457_, new_A2458_, new_A2459_, new_A2460_, new_A2461_, new_A2462_,
    new_A2463_, new_A2464_, new_A2465_, new_A2466_, new_A2467_, new_A2468_,
    new_A2469_, new_A2470_, new_A2471_, new_A2472_, new_A2473_, new_A2474_,
    new_A2475_, new_A2481_, new_A2482_, new_A2483_, new_A2484_, new_A2485_,
    new_A2486_, new_A2487_, new_A2488_, new_A2489_, new_A2490_, new_A2491_,
    new_A2492_, new_A2493_, new_A2494_, new_A2495_, new_A2496_, new_A2497_,
    new_A2498_, new_A2499_, new_A2500_, new_A2501_, new_A2502_, new_A2503_,
    new_A2504_, new_A2505_, new_A2506_, new_A2507_, new_A2508_, new_A2514_,
    new_A2515_, new_A2516_, new_A2517_, new_A2518_, new_A2519_, new_A2520_,
    new_A2521_, new_A2522_, new_A2523_, new_A2524_, new_A2525_, new_A2526_,
    new_A2527_, new_A2528_, new_A2529_, new_A2530_, new_A2531_, new_A2532_,
    new_A2533_, new_A2534_, new_A2535_, new_A2536_, new_A2537_, new_A2538_,
    new_A2539_, new_A2540_, new_A2541_, new_A2547_, new_A2548_, new_A2549_,
    new_A2550_, new_A2551_, new_A2552_, new_A2553_, new_A2554_, new_A2555_,
    new_A2556_, new_A2557_, new_A2558_, new_A2559_, new_A2560_, new_A2561_,
    new_A2562_, new_A2563_, new_A2564_, new_A2565_, new_A2566_, new_A2567_,
    new_A2568_, new_A2569_, new_A2570_, new_A2571_, new_A2572_, new_A2573_,
    new_A2574_, new_A2580_, new_A2581_, new_A2582_, new_A2583_, new_A2584_,
    new_A2585_, new_A2586_, new_A2587_, new_A2588_, new_A2589_, new_A2590_,
    new_A2591_, new_A2592_, new_A2593_, new_A2594_, new_A2595_, new_A2596_,
    new_A2597_, new_A2598_, new_A2599_, new_A2600_, new_A2601_, new_A2602_,
    new_A2603_, new_A2604_, new_A2605_, new_A2606_, new_A2607_, new_A2613_,
    new_A2614_, new_A2615_, new_A2616_, new_A2617_, new_A2618_, new_A2619_,
    new_A2620_, new_A2621_, new_A2622_, new_A2623_, new_A2624_, new_A2625_,
    new_A2626_, new_A2627_, new_A2628_, new_A2629_, new_A2630_, new_A2631_,
    new_A2632_, new_A2633_, new_A2634_, new_A2635_, new_A2636_, new_A2637_,
    new_A2638_, new_A2639_, new_A2640_, new_A2646_, new_A2647_, new_A2648_,
    new_A2649_, new_A2650_, new_A2651_, new_A2652_, new_A2653_, new_A2654_,
    new_A2655_, new_A2656_, new_A2657_, new_A2658_, new_A2659_, new_A2660_,
    new_A2661_, new_A2662_, new_A2663_, new_A2664_, new_A2665_, new_A2666_,
    new_A2667_, new_A2668_, new_A2669_, new_A2670_, new_A2671_, new_A2672_,
    new_A2673_, new_A2679_, new_A2680_, new_A2681_, new_A2682_, new_A2683_,
    new_A2684_, new_A2685_, new_A2686_, new_A2687_, new_A2688_, new_A2689_,
    new_A2690_, new_A2691_, new_A2692_, new_A2693_, new_A2694_, new_A2695_,
    new_A2696_, new_A2697_, new_A2698_, new_A2699_, new_A2700_, new_A2701_,
    new_A2702_, new_A2703_, new_A2704_, new_A2705_, new_A2706_, new_A2712_,
    new_A2713_, new_A2714_, new_A2715_, new_A2716_, new_A2717_, new_A2718_,
    new_A2719_, new_A2720_, new_A2721_, new_A2722_, new_A2723_, new_A2724_,
    new_A2725_, new_A2726_, new_A2727_, new_A2728_, new_A2729_, new_A2730_,
    new_A2731_, new_A2732_, new_A2733_, new_A2734_, new_A2735_, new_A2736_,
    new_A2737_, new_A2738_, new_A2739_, new_A2745_, new_A2746_, new_A2747_,
    new_A2748_, new_A2749_, new_A2750_, new_A2751_, new_A2752_, new_A2753_,
    new_A2754_, new_A2755_, new_A2756_, new_A2757_, new_A2758_, new_A2759_,
    new_A2760_, new_A2761_, new_A2762_, new_A2763_, new_A2764_, new_A2765_,
    new_A2766_, new_A2767_, new_A2768_, new_A2769_, new_A2770_, new_A2771_,
    new_A2772_, new_A2778_, new_A2779_, new_A2780_, new_A2781_, new_A2782_,
    new_A2783_, new_A2784_, new_A2785_, new_A2786_, new_A2787_, new_A2788_,
    new_A2789_, new_A2790_, new_A2791_, new_A2792_, new_A2793_, new_A2794_,
    new_A2795_, new_A2796_, new_A2797_, new_A2798_, new_A2799_, new_A2800_,
    new_A2801_, new_A2802_, new_A2803_, new_A2804_, new_A2805_, new_A1188_,
    new_A1187_, new_A1186_, new_A1185_, new_A1184_, new_A1183_, new_A1182_,
    new_A1181_, new_A1180_, new_A1179_, new_A1178_, new_A1177_, new_A1176_,
    new_A1175_, new_A1174_, new_A1173_, new_A1172_, new_A1171_, new_A1170_,
    new_A1169_, new_A1168_, new_A1167_, new_A1166_, new_A1165_, new_A1164_,
    new_A1163_, new_A1162_, new_A1161_, new_A1160_, new_A1159_, new_A1158_,
    new_A1157_, new_A1156_, new_A1189_, new_A1190_, new_A1191_, new_A1192_,
    new_A1193_, new_A1194_, new_A1195_, new_A1196_, new_A1197_, new_A1198_,
    new_A1199_, new_A1200_, new_A1201_, new_A1202_, new_A1203_, new_A1204_,
    new_A1205_, new_A1206_, new_A1207_, new_A1208_, new_A1209_, new_A1210_,
    new_A1211_, new_A1212_, new_A1213_, new_A1214_, new_A1215_, new_A1216_,
    new_A1217_, new_A1218_, new_A1219_, new_A1220_, new_A1221_, new_A1222_,
    new_A1223_, new_A1224_, new_A1225_, new_A1226_, new_A1227_, new_A1228_,
    new_A1229_, new_A1230_, new_A1231_, new_A1232_, new_A1233_, new_A1234_,
    new_A1235_, new_A1236_, new_A1237_, new_A1238_, new_A1239_, new_A1240_,
    new_A1241_, new_A1242_, new_A1243_, new_A1244_, new_A1245_, new_A1246_,
    new_A1247_, new_A1248_, new_A1249_, new_A1250_, new_A1251_, new_A1252_,
    new_A1253_, new_A1254_, new_A1255_, new_A1256_, new_A1257_, new_A1258_,
    new_A1259_, new_A1260_, new_A1261_, new_A1262_, new_A1263_, new_A1264_,
    new_A1265_, new_A1266_, new_A1267_, new_A1268_, new_A1269_, new_A1270_,
    new_A1271_, new_A1272_, new_A1273_, new_A1274_, new_A1275_, new_A1276_,
    new_A1277_, new_A1278_, new_A1279_, new_A1280_, new_A1281_, new_A1282_,
    new_A1283_, new_A1284_, new_A1285_, new_A1286_, new_A1287_, new_A1288_,
    new_A1289_, new_A1290_, new_A1291_, new_A1292_, new_A1293_, new_A1294_,
    new_A1295_, new_A1296_, new_A1297_, new_A1298_, new_A1299_, new_A1300_,
    new_A1301_, new_A1302_, new_A1303_, new_A1304_, new_A1305_, new_A1306_,
    new_A1307_, new_A1308_, new_A1309_, new_A1310_, new_A1311_, new_A1312_,
    new_A1313_, new_A1314_, new_A1315_, new_A1316_, new_A1317_, new_A1318_,
    new_A1319_, new_A1320_, new_A1321_, new_A1322_, new_A1323_, new_A1324_,
    new_A1325_, new_A1326_, new_A1327_, new_A1328_, new_A1329_, new_A1330_,
    new_A1331_, new_A1332_, new_A1333_, new_A1334_, new_A1335_, new_A1336_,
    new_A1337_, new_A1338_, new_A1339_, new_A1340_, new_A1341_, new_A1342_,
    new_A1343_, new_A1344_, new_A1345_, new_A1346_, new_A1347_, new_A1348_,
    new_A1349_, new_A1350_, new_A1351_, new_A1352_, new_A1353_, new_A1354_,
    new_A1355_, new_A1356_, new_A1357_, new_A1358_, new_A1359_, new_A1360_,
    new_A1361_, new_A1362_, new_A1363_, new_A1364_, new_A1365_, new_A1366_,
    new_A1367_, new_A1368_, new_A1369_, new_A1370_, new_A1371_, new_A1372_,
    new_A1373_, new_A1374_, new_A1375_, new_A1376_, new_A1377_, new_A1378_,
    new_A1379_, new_A1380_, new_A1381_, new_A1382_, new_A1383_, new_A1384_,
    new_A1385_, new_A1386_, new_A1387_, new_A1388_, new_A1389_, new_A1390_,
    new_A1391_, new_A1392_, new_A1393_, new_A1394_, new_A1395_, new_A1396_,
    new_A1397_, new_A1398_, new_A1399_, new_A1400_, new_A1401_, new_A1402_,
    new_A1403_, new_A1404_, new_A1405_, new_A1406_, new_A1407_, new_A1408_,
    new_A1409_, new_A1410_, new_A1411_, new_A1412_, new_A1413_, new_A1414_,
    new_A1415_, new_A1416_, new_A1417_, new_A1418_, new_A1419_, new_A1420_,
    new_A1421_, new_A1422_, new_A1423_, new_A1424_, new_A1425_, new_A1426_,
    new_A1427_, new_A1428_, new_A1429_, new_A1430_, new_A1431_, new_A1432_,
    new_A1433_, new_A1434_, new_A1435_, new_A1436_, new_A1437_, new_A1438_,
    new_A1439_, new_A1440_, new_A1441_, new_A1442_, new_A1443_, new_A1444_,
    new_A1445_, new_A1446_, new_A1447_, new_A1448_, new_A1449_, new_A1450_,
    new_A1451_, new_A1452_, new_A1453_, new_A1454_, new_A1455_, new_A1456_,
    new_A1457_, new_A1458_, new_A1459_, new_A1460_, new_A1461_, new_A1462_,
    new_A1463_, new_A1464_, new_A1465_, new_A1466_, new_A1467_, new_A1468_,
    new_A1469_, new_A1470_, new_A1471_, new_A1472_, new_A1473_, new_A1474_,
    new_A1475_, new_A1476_, new_A1477_, new_A1478_, new_A1479_, new_A1480_,
    new_A1481_, new_A1482_, new_A1483_, new_A1484_, new_A1485_, new_A1486_,
    new_A1487_, new_A1488_, new_A1489_, new_A1490_, new_A1491_, new_A1492_,
    new_A1493_, new_A1494_, new_A1495_, new_A1496_, new_A1497_, new_A1498_,
    new_A1499_, new_A1500_, new_A1501_, new_A1502_, new_A1503_, new_A1504_,
    new_A1505_, new_A1506_, new_A1507_, new_A1508_, new_A1509_, new_A1510_,
    new_A1511_, new_A1512_, new_A1513_, new_A1514_, new_A1515_, new_A1516_,
    new_A1517_, new_A1518_, new_A1519_, new_A1520_, new_A1521_, new_A1522_,
    new_A1523_, new_A1524_, new_A1525_, new_A1526_, new_A1527_, new_A1528_,
    new_A1529_, new_A1530_, new_A1531_, new_A1532_, new_A1533_, new_A1534_,
    new_A1535_, new_A1536_, new_A1537_, new_A1538_, new_A1539_, new_A1540_,
    new_A1541_, new_A1542_, new_A1543_, new_A1544_, new_A1545_, new_A1546_,
    new_A1547_, new_A1548_, new_A1549_, new_A1550_, new_A1551_, new_A1552_,
    new_A1553_, new_A1554_, new_A1555_, new_A1556_, new_A1557_, new_A1558_,
    new_A1559_, new_A1560_, new_A1561_, new_A1562_, new_A1563_, new_A1564_,
    new_A1565_, new_A1566_, new_A1567_, new_A1568_, new_A1569_, new_A1570_,
    new_A1571_, new_A1572_, new_A1573_, new_A1574_, new_A1575_, new_A1576_,
    new_A1577_, new_A1578_, new_A1579_, new_A1580_, new_A1581_, new_A1582_,
    new_A1583_, new_A1584_, new_A1585_, new_A1586_, new_A1587_, new_A1588_,
    new_A1589_, new_A1590_, new_A1591_, new_A1592_, new_A1593_, new_A1594_,
    new_A1595_, new_A1596_, new_A1597_, new_A1598_, new_A1599_, new_A1600_,
    new_A1601_, new_A1602_, new_A1603_, new_A1604_, new_A1605_, new_A1606_,
    new_A1607_, new_A1608_, new_A1609_, new_A1610_, new_A1611_, new_A1612_,
    new_A1613_, new_A1614_, new_A1615_, new_A1616_, new_A1617_, new_A1618_,
    new_A1619_, new_A1620_, new_A1621_, new_A1622_, new_A1623_, new_A1624_,
    new_A1625_, new_A1626_, new_A1627_, new_A1628_, new_A1629_, new_A1630_,
    new_A1631_, new_A1632_, new_A1633_, new_A1634_, new_A1635_, new_A1636_,
    new_A1637_, new_A1638_, new_A1639_, new_A1640_, new_A1641_, new_A1642_,
    new_A1643_, new_A1644_, new_A1645_, new_A1646_, new_A1647_, new_A1648_,
    new_A1649_, new_A1650_, new_A1651_, new_A1652_, new_A1653_, new_A1654_,
    new_A1655_, new_A1656_, new_A1657_, new_A1658_, new_A1659_, new_A1660_,
    new_A1661_, new_A1662_, new_A1663_, new_A1664_, new_A1665_, new_A1666_,
    new_A1667_, new_A1668_, new_A1669_, new_A1670_, new_A1671_, new_A1672_,
    new_A1673_, new_A1674_, new_A1675_, new_A1676_, new_A1677_, new_A1678_,
    new_A1679_, new_A1680_, new_A1681_, new_A1682_, new_A1683_, new_A1684_,
    new_A1685_, new_A1686_, new_A1687_, new_A1688_, new_A1689_, new_A1690_,
    new_A1691_, new_A1692_, new_A1693_, new_A1694_, new_A1695_, new_A1696_,
    new_A1697_, new_A1698_, new_A1699_, new_A1700_, new_A1701_, new_A1702_,
    new_A1703_, new_A1704_, new_A1705_, new_A1706_, new_A1707_, new_A1708_,
    new_A1709_, new_A1710_, new_A1711_, new_A1712_, new_A1713_, new_A1714_,
    new_A1715_, new_A1716_, new_A1717_, new_A1718_, new_A1719_, new_A1720_,
    new_A1721_, new_A1722_, new_A1723_, new_A1724_, new_A1725_, new_A1726_,
    new_A1727_, new_A1728_, new_A1729_, new_A1730_, new_A1731_, new_A1732_,
    new_A1733_, new_A1734_, new_A1735_, new_A1736_, new_A1737_, new_A1738_,
    new_A1739_, new_A1740_, new_A1741_, new_A1742_, new_A1743_, new_A1744_,
    new_A1745_, new_A1746_, new_A1747_, new_A1748_, new_A1749_, new_A1750_,
    new_A1751_, new_A1752_, new_A1753_, new_A1754_, new_A1755_, new_A1756_,
    new_A1757_, new_A1758_, new_A1759_, new_A1760_, new_A1761_, new_A1762_,
    new_A1763_, new_A1764_, new_A1765_, new_A1766_, new_A1767_, new_A1768_,
    new_A1769_, new_A1770_, new_A1771_, new_A1772_, new_A1773_, new_A1774_,
    new_A1775_, new_A1776_, new_A1777_, new_A1778_, new_A1779_, new_A1780_,
    new_A1781_, new_A1782_, new_A1783_, new_A1784_, new_A1785_, new_A1786_,
    new_A1787_, new_A1788_, new_A1789_, new_A1790_, new_A1791_, new_A1792_,
    new_A1793_, new_A1794_, new_A1795_, new_A1796_, new_A1797_, new_A1798_,
    new_A1799_, new_A1800_, new_A1801_, new_A1802_, new_A1803_, new_A1804_,
    new_A1805_, new_A1806_, new_A1807_, new_A1808_, new_A1809_, new_A1810_,
    new_A1811_, new_A1812_, new_A1813_, new_A1814_, new_A1815_, new_A1816_,
    new_A1817_, new_A1818_, new_A1819_, new_A1820_, new_A1821_, new_A1822_,
    new_A1823_, new_A1824_, new_A1825_, new_A1826_, new_A1827_, new_A1828_,
    new_A1829_, new_A1830_, new_A1831_, new_A1832_, new_A1833_, new_A1834_,
    new_A1835_, new_A1836_, new_A1837_, new_A1838_, new_A1839_, new_A1840_,
    new_A1841_, new_A1842_, new_A1843_, new_A1844_, new_A1845_, new_A1846_,
    new_A1847_, new_A1848_, new_A1849_, new_A1850_, new_A1851_, new_A1852_,
    new_A1853_, new_A1854_, new_A1855_, new_A1856_, new_A1857_, new_A1858_,
    new_A1859_, new_A1860_, new_A1861_, new_A1862_, new_A1863_, new_A1864_,
    new_A1865_, new_A1866_, new_A1867_, new_A1868_, new_A1869_, new_A1870_,
    new_A1871_, new_A1872_, new_A1873_, new_A1874_, new_A1875_, new_A1876_,
    new_A1877_, new_A1878_, new_A1879_, new_A1880_, new_A1881_, new_A1882_,
    new_A1883_, new_A1884_, new_A1885_, new_A1886_, new_A1887_, new_A1888_,
    new_A1889_, new_A1890_, new_A1891_, new_A1892_, new_A1893_, new_A1894_,
    new_A1895_, new_A1896_, new_A1897_, new_A1898_, new_A1899_, new_A1900_,
    new_A1901_, new_A1902_, new_A1903_, new_A1904_, new_A1905_, new_A1906_,
    new_A1907_, new_A1908_, new_A1909_, new_A1910_, new_A1911_, new_A1912_,
    new_A1913_, new_A1914_, new_A1915_, new_A1916_, new_A1917_, new_A1918_,
    new_A1919_, new_A1920_, new_A1921_, new_A1922_, new_A1923_, new_A1924_,
    new_A1925_, new_A1926_, new_A1927_, new_A1928_, new_A1929_, new_A1930_,
    new_A1931_, new_A1932_, new_A1933_, new_A1934_, new_A1935_, new_A1936_,
    new_A1937_, new_A1938_, new_A1939_, new_A1940_, new_A1941_, new_A1942_,
    new_A1943_, new_A1944_, new_A1945_, new_A1946_, new_A1947_, new_A1948_,
    new_A1949_, new_A1950_, new_A1951_, new_A1952_, new_A1953_, new_A1954_,
    new_A1955_, new_A1956_, new_A1957_, new_A1958_, new_A1959_, new_A1960_,
    new_A1961_, new_A1962_, new_A1963_, new_A1964_, new_A1965_, new_A1966_,
    new_A1967_, new_A1968_, new_A1969_, new_A1970_, new_A1971_, new_A1972_,
    new_A1973_, new_A1974_, new_A1975_, new_A1976_, new_A1977_, new_A1978_,
    new_A1979_, new_A1980_, new_A1155_, new_A1154_, new_A1153_, new_A1152_,
    new_A1151_, new_A1150_, new_A1149_, new_A1148_, new_A1147_, new_A1146_,
    new_A1145_, new_A1144_, new_A1143_, new_A1142_, new_A1141_, new_A1140_,
    new_A1139_, new_A1138_, new_A1137_, new_A1136_, new_A1135_, new_A1134_,
    new_A1133_, new_A1127_, new_A1126_, new_A1125_, new_A1124_, new_A1123_,
    new_A1122_, new_A1121_, new_A1120_, new_A1119_, new_A1118_, new_A1117_,
    new_A1116_, new_A1115_, new_A1114_, new_A1113_, new_A1112_, new_A1111_,
    new_A1110_, new_A1109_, new_A1108_, new_A1107_, new_A1106_, new_A1105_,
    new_A1104_, new_A1103_, new_A1102_, new_A1101_, new_A1100_, new_A1094_,
    new_A1093_, new_A1092_, new_A1091_, new_A1090_, new_A1089_, new_A1088_,
    new_A1087_, new_A1086_, new_A1085_, new_A1084_, new_A1083_, new_A1082_,
    new_A1081_, new_A1080_, new_A1079_, new_A1078_, new_A1077_, new_A1076_,
    new_A1075_, new_A1074_, new_A1073_, new_A1072_, new_A1071_, new_A1070_,
    new_A1069_, new_A1068_, new_A1067_, new_A1061_, new_A1060_, new_A1059_,
    new_A1058_, new_A1057_, new_A1056_, new_A1055_, new_A1054_, new_A1053_,
    new_A1052_, new_A1051_, new_A1050_, new_A1049_, new_A1048_, new_A1047_,
    new_A1046_, new_A1045_, new_A1044_, new_A1043_, new_A1042_, new_A1041_,
    new_A1040_, new_A1039_, new_A1038_, new_A1037_, new_A1036_, new_A1035_,
    new_A1034_, new_A1028_, new_A1027_, new_A1026_, new_A1025_, new_A1024_,
    new_A1023_, new_A1022_, new_A1021_, new_A1020_, new_A1019_, new_A1018_,
    new_A1017_, new_A1016_, new_A1015_, new_A1014_, new_A1013_, new_A1012_,
    new_A1011_, new_A1010_, new_A1009_, new_A1008_, new_A1007_, new_A1006_,
    new_A1005_, new_A1004_, new_A1003_, new_A1002_, new_A1001_, new_A995_,
    new_A994_, new_A993_, new_A992_, new_A991_, new_A990_, new_A989_,
    new_A988_, new_A987_, new_A986_, new_A985_, new_A984_, new_A983_,
    new_A982_, new_A981_, new_A980_, new_A979_, new_A978_, new_A977_,
    new_A976_, new_A975_, new_A974_, new_A973_, new_A972_, new_A971_,
    new_A970_, new_A969_, new_A968_, new_A962_, new_A961_, new_A960_,
    new_A959_, new_A958_, new_A957_, new_A956_, new_A955_, new_A954_,
    new_A953_, new_A952_, new_A951_, new_A950_, new_A949_, new_A948_,
    new_A947_, new_A946_, new_A945_, new_A944_, new_A943_, new_A942_,
    new_A941_, new_A940_, new_A939_, new_A938_, new_A937_, new_A936_,
    new_A935_, new_A929_, new_A928_, new_A927_, new_A926_, new_A925_,
    new_A924_, new_A923_, new_A922_, new_A921_, new_A920_, new_A919_,
    new_A918_, new_A917_, new_A916_, new_A915_, new_A914_, new_A913_,
    new_A912_, new_A911_, new_A910_, new_A909_, new_A908_, new_A907_,
    new_A906_, new_A905_, new_A904_, new_A903_, new_A902_, new_A896_,
    new_A895_, new_A894_, new_A893_, new_A892_, new_A891_, new_A890_,
    new_A889_, new_A888_, new_A887_, new_A886_, new_A885_, new_A884_,
    new_A883_, new_A882_, new_A881_, new_A880_, new_A879_, new_A878_,
    new_A877_, new_A876_, new_A875_, new_A874_, new_A873_, new_A872_,
    new_A871_, new_A870_, new_A869_, new_A863_, new_A862_, new_A861_,
    new_A860_, new_A859_, new_A858_, new_A857_, new_A856_, new_A855_,
    new_A854_, new_A853_, new_A852_, new_A851_, new_A850_, new_A849_,
    new_A848_, new_A847_, new_A846_, new_A845_, new_A844_, new_A843_,
    new_A842_, new_A841_, new_A840_, new_A839_, new_A838_, new_A837_,
    new_A836_, new_A830_, new_A829_, new_A828_, new_A827_, new_A826_,
    new_A825_, new_A824_, new_A823_, new_A822_, new_A821_, new_A820_,
    new_A819_, new_A818_, new_A817_, new_A816_, new_A815_, new_A814_,
    new_A813_, new_A812_, new_A811_, new_A810_, new_A809_, new_A808_,
    new_A807_, new_A806_, new_A805_, new_A804_, new_A803_, new_A797_,
    new_A796_, new_A795_, new_A794_, new_A793_, new_A792_, new_A791_,
    new_A790_, new_A789_, new_A788_, new_A787_, new_A786_, new_A785_,
    new_A784_, new_A783_, new_A782_, new_A781_, new_A780_, new_A779_,
    new_A778_, new_A777_, new_A776_, new_A775_, new_A774_, new_A773_,
    new_A772_, new_A771_, new_A770_, new_A764_, new_A763_, new_A762_,
    new_A761_, new_A760_, new_A759_, new_A758_, new_A757_, new_A756_,
    new_A755_, new_A754_, new_A753_, new_A752_, new_A751_, new_A750_,
    new_A749_, new_A748_, new_A747_, new_A746_, new_A745_, new_A744_,
    new_A743_, new_A742_, new_A741_, new_A740_, new_A739_, new_A738_,
    new_A737_, new_A731_, new_A730_, new_A729_, new_A728_, new_A727_,
    new_A726_, new_A725_, new_A724_, new_A723_, new_A722_, new_A721_,
    new_A720_, new_A719_, new_A718_, new_A717_, new_A716_, new_A715_,
    new_A714_, new_A713_, new_A712_, new_A711_, new_A710_, new_A709_,
    new_A708_, new_A707_, new_A706_, new_A705_, new_A704_, new_A698_,
    new_A697_, new_A696_, new_A695_, new_A694_, new_A693_, new_A692_,
    new_A691_, new_A690_, new_A689_, new_A688_, new_A687_, new_A686_,
    new_A685_, new_A684_, new_A683_, new_A682_, new_A681_, new_A680_,
    new_A679_, new_A678_, new_A677_, new_A676_, new_A675_, new_A674_,
    new_A673_, new_A672_, new_A671_, new_A665_, new_A664_, new_A663_,
    new_A662_, new_A661_, new_A660_, new_A659_, new_A658_, new_A657_,
    new_A656_, new_A655_, new_A654_, new_A653_, new_A652_, new_A651_,
    new_A650_, new_A649_, new_A648_, new_A647_, new_A646_, new_A645_,
    new_A644_, new_A643_, new_A642_, new_A641_, new_A640_, new_A639_,
    new_A638_, new_A632_, new_A631_, new_A630_, new_A629_, new_A628_,
    new_A627_, new_A626_, new_A625_, new_A624_, new_A623_, new_A622_,
    new_A621_, new_A620_, new_A619_, new_A618_, new_A617_, new_A616_,
    new_A615_, new_A614_, new_A613_, new_A612_, new_A611_, new_A610_,
    new_A609_, new_A608_, new_A607_, new_A606_, new_A605_, new_A599_,
    new_A598_, new_A597_, new_A596_, new_A595_, new_A594_, new_A593_,
    new_A592_, new_A591_, new_A590_, new_A589_, new_A588_, new_A587_,
    new_A586_, new_A585_, new_A584_, new_A583_, new_A582_, new_A581_,
    new_A580_, new_A579_, new_A578_, new_A577_, new_A576_, new_A575_,
    new_A574_, new_A573_, new_A572_, new_A566_, new_A565_, new_A564_,
    new_A563_, new_A562_, new_A561_, new_A560_, new_A559_, new_A558_,
    new_A557_, new_A556_, new_A555_, new_A554_, new_A553_, new_A552_,
    new_A551_, new_A550_, new_A549_, new_A548_, new_A547_, new_A546_,
    new_A545_, new_A544_, new_A543_, new_A542_, new_A541_, new_A540_,
    new_A539_, new_A533_, new_A532_, new_A531_, new_A530_, new_A529_,
    new_A528_, new_A527_, new_A526_, new_A525_, new_A524_, new_A523_,
    new_A522_, new_A521_, new_A520_, new_A519_, new_A518_, new_A517_,
    new_A516_, new_A515_, new_A514_, new_A513_, new_A512_, new_A511_,
    new_A510_, new_A509_, new_A508_, new_A507_, new_A506_, new_A500_,
    new_A499_, new_A498_, new_A497_, new_A496_, new_A495_, new_A494_,
    new_A493_, new_A492_, new_A491_, new_A490_, new_A489_, new_A488_,
    new_A487_, new_A486_, new_A485_, new_A484_, new_A483_, new_A482_,
    new_A481_, new_A480_, new_A479_, new_A478_, new_A477_, new_A476_,
    new_A475_, new_A474_, new_A473_, new_A467_, new_A466_, new_A465_,
    new_A464_, new_A463_, new_A462_, new_A461_, new_A460_, new_A459_,
    new_A458_, new_A457_, new_A456_, new_A455_, new_A454_, new_A453_,
    new_A452_, new_A451_, new_A450_, new_A449_, new_A448_, new_A447_,
    new_A446_, new_A445_, new_A444_, new_A443_, new_A442_, new_A441_,
    new_A440_, new_A434_, new_A433_, new_A432_, new_A431_, new_A430_,
    new_A429_, new_A428_, new_A427_, new_A426_, new_A425_, new_A424_,
    new_A423_, new_A422_, new_A421_, new_A420_, new_A419_, new_A418_,
    new_A417_, new_A416_, new_A415_, new_A414_, new_A413_, new_A412_,
    new_A411_, new_A410_, new_A409_, new_A408_, new_A407_, new_A401_,
    new_A400_, new_A399_, new_A398_, new_A397_, new_A396_, new_A395_,
    new_A394_, new_A393_, new_A392_, new_A391_, new_A390_, new_A389_,
    new_A388_, new_A387_, new_A386_, new_A385_, new_A384_, new_A383_,
    new_A382_, new_A381_, new_A380_, new_A379_, new_A378_, new_A377_,
    new_A376_, new_A375_, new_A374_, new_A368_, new_A367_, new_A366_,
    new_A365_, new_A364_, new_A331_, new_A332_, new_A333_, new_A334_,
    new_A335_, new_A341_, new_A342_, new_A343_, new_A344_, new_A345_,
    new_A346_, new_A347_, new_A348_, new_A349_, new_A350_, new_A351_,
    new_A352_, new_A353_, new_A354_, new_A355_, new_A356_, new_A357_,
    new_A358_, new_A359_, new_A360_, new_A361_, new_A362_, new_A363_;
  assign new_A2013_ = new_A1991_ & new_A2006_;
  assign new_A2012_ = ~new_A1991_ & ~new_A2013_;
  assign new_A2011_ = new_A1991_ | new_A2006_;
  assign new_A2010_ = ~A1984 | ~A1985;
  assign new_A2009_ = new_A1991_ | new_A2006_;
  assign new_A2008_ = ~new_A2007_ & ~new_A1991_;
  assign new_A2007_ = new_A1991_ & new_A2006_;
  assign new_A2006_ = ~A1982 | ~A1983;
  assign new_A2005_ = A1983 & new_A1995_;
  assign new_A2004_ = A1984 | new_A1991_;
  assign new_A2003_ = A1984 | A1985;
  assign new_A2002_ = ~new_A2012_ | ~new_A2011_;
  assign new_A2001_ = new_A2010_ & new_A2003_;
  assign new_A2000_ = A1984 ^ new_A1991_;
  assign new_A1999_ = ~new_A2008_ | ~new_A2009_;
  assign new_A1998_ = ~A1983 ^ new_A1995_;
  assign new_A1997_ = new_A2005_ | A1982;
  assign new_A1996_ = new_A2002_ & A1983;
  assign new_A1995_ = new_A2004_ & new_A2003_;
  assign new_A1994_ = new_A1999_ & A1983;
  assign new_A1993_ = new_A2001_ & new_A2000_;
  assign new_A1992_ = new_A1993_ ^ A1983;
  assign new_A1991_ = A1981 ^ A1982;
  assign new_A1990_ = new_A1991_ & new_A1998_;
  assign new_A1989_ = new_A1991_ & new_A1997_;
  assign new_A1988_ = new_A1996_ | new_A1995_;
  assign new_A1987_ = new_A1994_ | new_A1993_;
  assign new_A1986_ = new_A1992_ & new_A1991_;
  assign new_A2019_ = new_A2025_ & new_A2024_;
  assign new_A2020_ = new_A2027_ | new_A2026_;
  assign new_A2021_ = new_A2029_ | new_A2028_;
  assign new_A2022_ = new_A2024_ & new_A2030_;
  assign new_A2023_ = new_A2024_ & new_A2031_;
  assign new_A2024_ = A2014 ^ A2015;
  assign new_A2025_ = new_A2026_ ^ A2016;
  assign new_A2026_ = new_A2034_ & new_A2033_;
  assign new_A2027_ = new_A2032_ & A2016;
  assign new_A2028_ = new_A2037_ & new_A2036_;
  assign new_A2029_ = new_A2035_ & A2016;
  assign new_A2030_ = new_A2038_ | A2015;
  assign new_A2031_ = ~A2016 ^ new_A2028_;
  assign new_A2032_ = ~new_A2041_ | ~new_A2042_;
  assign new_A2033_ = A2017 ^ new_A2024_;
  assign new_A2034_ = new_A2043_ & new_A2036_;
  assign new_A2035_ = ~new_A2045_ | ~new_A2044_;
  assign new_A2036_ = A2017 | A2018;
  assign new_A2037_ = A2017 | new_A2024_;
  assign new_A2038_ = A2016 & new_A2028_;
  assign new_A2039_ = ~A2015 | ~A2016;
  assign new_A2040_ = new_A2024_ & new_A2039_;
  assign new_A2041_ = ~new_A2040_ & ~new_A2024_;
  assign new_A2042_ = new_A2024_ | new_A2039_;
  assign new_A2043_ = ~A2017 | ~A2018;
  assign new_A2044_ = new_A2024_ | new_A2039_;
  assign new_A2045_ = ~new_A2024_ & ~new_A2046_;
  assign new_A2046_ = new_A2024_ & new_A2039_;
  assign new_A2052_ = new_A2058_ & new_A2057_;
  assign new_A2053_ = new_A2060_ | new_A2059_;
  assign new_A2054_ = new_A2062_ | new_A2061_;
  assign new_A2055_ = new_A2057_ & new_A2063_;
  assign new_A2056_ = new_A2057_ & new_A2064_;
  assign new_A2057_ = A2047 ^ A2048;
  assign new_A2058_ = new_A2059_ ^ A2049;
  assign new_A2059_ = new_A2067_ & new_A2066_;
  assign new_A2060_ = new_A2065_ & A2049;
  assign new_A2061_ = new_A2070_ & new_A2069_;
  assign new_A2062_ = new_A2068_ & A2049;
  assign new_A2063_ = new_A2071_ | A2048;
  assign new_A2064_ = ~A2049 ^ new_A2061_;
  assign new_A2065_ = ~new_A2074_ | ~new_A2075_;
  assign new_A2066_ = A2050 ^ new_A2057_;
  assign new_A2067_ = new_A2076_ & new_A2069_;
  assign new_A2068_ = ~new_A2078_ | ~new_A2077_;
  assign new_A2069_ = A2050 | A2051;
  assign new_A2070_ = A2050 | new_A2057_;
  assign new_A2071_ = A2049 & new_A2061_;
  assign new_A2072_ = ~A2048 | ~A2049;
  assign new_A2073_ = new_A2057_ & new_A2072_;
  assign new_A2074_ = ~new_A2073_ & ~new_A2057_;
  assign new_A2075_ = new_A2057_ | new_A2072_;
  assign new_A2076_ = ~A2050 | ~A2051;
  assign new_A2077_ = new_A2057_ | new_A2072_;
  assign new_A2078_ = ~new_A2057_ & ~new_A2079_;
  assign new_A2079_ = new_A2057_ & new_A2072_;
  assign new_A2085_ = new_A2091_ & new_A2090_;
  assign new_A2086_ = new_A2093_ | new_A2092_;
  assign new_A2087_ = new_A2095_ | new_A2094_;
  assign new_A2088_ = new_A2090_ & new_A2096_;
  assign new_A2089_ = new_A2090_ & new_A2097_;
  assign new_A2090_ = A2080 ^ A2081;
  assign new_A2091_ = new_A2092_ ^ A2082;
  assign new_A2092_ = new_A2100_ & new_A2099_;
  assign new_A2093_ = new_A2098_ & A2082;
  assign new_A2094_ = new_A2103_ & new_A2102_;
  assign new_A2095_ = new_A2101_ & A2082;
  assign new_A2096_ = new_A2104_ | A2081;
  assign new_A2097_ = ~A2082 ^ new_A2094_;
  assign new_A2098_ = ~new_A2107_ | ~new_A2108_;
  assign new_A2099_ = A2083 ^ new_A2090_;
  assign new_A2100_ = new_A2109_ & new_A2102_;
  assign new_A2101_ = ~new_A2111_ | ~new_A2110_;
  assign new_A2102_ = A2083 | A2084;
  assign new_A2103_ = A2083 | new_A2090_;
  assign new_A2104_ = A2082 & new_A2094_;
  assign new_A2105_ = ~A2081 | ~A2082;
  assign new_A2106_ = new_A2090_ & new_A2105_;
  assign new_A2107_ = ~new_A2106_ & ~new_A2090_;
  assign new_A2108_ = new_A2090_ | new_A2105_;
  assign new_A2109_ = ~A2083 | ~A2084;
  assign new_A2110_ = new_A2090_ | new_A2105_;
  assign new_A2111_ = ~new_A2090_ & ~new_A2112_;
  assign new_A2112_ = new_A2090_ & new_A2105_;
  assign new_A2118_ = new_A2124_ & new_A2123_;
  assign new_A2119_ = new_A2126_ | new_A2125_;
  assign new_A2120_ = new_A2128_ | new_A2127_;
  assign new_A2121_ = new_A2123_ & new_A2129_;
  assign new_A2122_ = new_A2123_ & new_A2130_;
  assign new_A2123_ = A2113 ^ A2114;
  assign new_A2124_ = new_A2125_ ^ A2115;
  assign new_A2125_ = new_A2133_ & new_A2132_;
  assign new_A2126_ = new_A2131_ & A2115;
  assign new_A2127_ = new_A2136_ & new_A2135_;
  assign new_A2128_ = new_A2134_ & A2115;
  assign new_A2129_ = new_A2137_ | A2114;
  assign new_A2130_ = ~A2115 ^ new_A2127_;
  assign new_A2131_ = ~new_A2140_ | ~new_A2141_;
  assign new_A2132_ = A2116 ^ new_A2123_;
  assign new_A2133_ = new_A2142_ & new_A2135_;
  assign new_A2134_ = ~new_A2144_ | ~new_A2143_;
  assign new_A2135_ = A2116 | A2117;
  assign new_A2136_ = A2116 | new_A2123_;
  assign new_A2137_ = A2115 & new_A2127_;
  assign new_A2138_ = ~A2114 | ~A2115;
  assign new_A2139_ = new_A2123_ & new_A2138_;
  assign new_A2140_ = ~new_A2139_ & ~new_A2123_;
  assign new_A2141_ = new_A2123_ | new_A2138_;
  assign new_A2142_ = ~A2116 | ~A2117;
  assign new_A2143_ = new_A2123_ | new_A2138_;
  assign new_A2144_ = ~new_A2123_ & ~new_A2145_;
  assign new_A2145_ = new_A2123_ & new_A2138_;
  assign new_A2151_ = new_A2157_ & new_A2156_;
  assign new_A2152_ = new_A2159_ | new_A2158_;
  assign new_A2153_ = new_A2161_ | new_A2160_;
  assign new_A2154_ = new_A2156_ & new_A2162_;
  assign new_A2155_ = new_A2156_ & new_A2163_;
  assign new_A2156_ = A2146 ^ A2147;
  assign new_A2157_ = new_A2158_ ^ A2148;
  assign new_A2158_ = new_A2166_ & new_A2165_;
  assign new_A2159_ = new_A2164_ & A2148;
  assign new_A2160_ = new_A2169_ & new_A2168_;
  assign new_A2161_ = new_A2167_ & A2148;
  assign new_A2162_ = new_A2170_ | A2147;
  assign new_A2163_ = ~A2148 ^ new_A2160_;
  assign new_A2164_ = ~new_A2173_ | ~new_A2174_;
  assign new_A2165_ = A2149 ^ new_A2156_;
  assign new_A2166_ = new_A2175_ & new_A2168_;
  assign new_A2167_ = ~new_A2177_ | ~new_A2176_;
  assign new_A2168_ = A2149 | A2150;
  assign new_A2169_ = A2149 | new_A2156_;
  assign new_A2170_ = A2148 & new_A2160_;
  assign new_A2171_ = ~A2147 | ~A2148;
  assign new_A2172_ = new_A2156_ & new_A2171_;
  assign new_A2173_ = ~new_A2172_ & ~new_A2156_;
  assign new_A2174_ = new_A2156_ | new_A2171_;
  assign new_A2175_ = ~A2149 | ~A2150;
  assign new_A2176_ = new_A2156_ | new_A2171_;
  assign new_A2177_ = ~new_A2156_ & ~new_A2178_;
  assign new_A2178_ = new_A2156_ & new_A2171_;
  assign new_A2184_ = new_A2190_ & new_A2189_;
  assign new_A2185_ = new_A2192_ | new_A2191_;
  assign new_A2186_ = new_A2194_ | new_A2193_;
  assign new_A2187_ = new_A2189_ & new_A2195_;
  assign new_A2188_ = new_A2189_ & new_A2196_;
  assign new_A2189_ = A2179 ^ A2180;
  assign new_A2190_ = new_A2191_ ^ A2181;
  assign new_A2191_ = new_A2199_ & new_A2198_;
  assign new_A2192_ = new_A2197_ & A2181;
  assign new_A2193_ = new_A2202_ & new_A2201_;
  assign new_A2194_ = new_A2200_ & A2181;
  assign new_A2195_ = new_A2203_ | A2180;
  assign new_A2196_ = ~A2181 ^ new_A2193_;
  assign new_A2197_ = ~new_A2206_ | ~new_A2207_;
  assign new_A2198_ = A2182 ^ new_A2189_;
  assign new_A2199_ = new_A2208_ & new_A2201_;
  assign new_A2200_ = ~new_A2210_ | ~new_A2209_;
  assign new_A2201_ = A2182 | A2183;
  assign new_A2202_ = A2182 | new_A2189_;
  assign new_A2203_ = A2181 & new_A2193_;
  assign new_A2204_ = ~A2180 | ~A2181;
  assign new_A2205_ = new_A2189_ & new_A2204_;
  assign new_A2206_ = ~new_A2205_ & ~new_A2189_;
  assign new_A2207_ = new_A2189_ | new_A2204_;
  assign new_A2208_ = ~A2182 | ~A2183;
  assign new_A2209_ = new_A2189_ | new_A2204_;
  assign new_A2210_ = ~new_A2189_ & ~new_A2211_;
  assign new_A2211_ = new_A2189_ & new_A2204_;
  assign new_A2217_ = new_A2223_ & new_A2222_;
  assign new_A2218_ = new_A2225_ | new_A2224_;
  assign new_A2219_ = new_A2227_ | new_A2226_;
  assign new_A2220_ = new_A2222_ & new_A2228_;
  assign new_A2221_ = new_A2222_ & new_A2229_;
  assign new_A2222_ = A2212 ^ A2213;
  assign new_A2223_ = new_A2224_ ^ A2214;
  assign new_A2224_ = new_A2232_ & new_A2231_;
  assign new_A2225_ = new_A2230_ & A2214;
  assign new_A2226_ = new_A2235_ & new_A2234_;
  assign new_A2227_ = new_A2233_ & A2214;
  assign new_A2228_ = new_A2236_ | A2213;
  assign new_A2229_ = ~A2214 ^ new_A2226_;
  assign new_A2230_ = ~new_A2239_ | ~new_A2240_;
  assign new_A2231_ = A2215 ^ new_A2222_;
  assign new_A2232_ = new_A2241_ & new_A2234_;
  assign new_A2233_ = ~new_A2243_ | ~new_A2242_;
  assign new_A2234_ = A2215 | A2216;
  assign new_A2235_ = A2215 | new_A2222_;
  assign new_A2236_ = A2214 & new_A2226_;
  assign new_A2237_ = ~A2213 | ~A2214;
  assign new_A2238_ = new_A2222_ & new_A2237_;
  assign new_A2239_ = ~new_A2238_ & ~new_A2222_;
  assign new_A2240_ = new_A2222_ | new_A2237_;
  assign new_A2241_ = ~A2215 | ~A2216;
  assign new_A2242_ = new_A2222_ | new_A2237_;
  assign new_A2243_ = ~new_A2222_ & ~new_A2244_;
  assign new_A2244_ = new_A2222_ & new_A2237_;
  assign new_A2250_ = new_A2256_ & new_A2255_;
  assign new_A2251_ = new_A2258_ | new_A2257_;
  assign new_A2252_ = new_A2260_ | new_A2259_;
  assign new_A2253_ = new_A2255_ & new_A2261_;
  assign new_A2254_ = new_A2255_ & new_A2262_;
  assign new_A2255_ = A2245 ^ A2246;
  assign new_A2256_ = new_A2257_ ^ A2247;
  assign new_A2257_ = new_A2265_ & new_A2264_;
  assign new_A2258_ = new_A2263_ & A2247;
  assign new_A2259_ = new_A2268_ & new_A2267_;
  assign new_A2260_ = new_A2266_ & A2247;
  assign new_A2261_ = new_A2269_ | A2246;
  assign new_A2262_ = ~A2247 ^ new_A2259_;
  assign new_A2263_ = ~new_A2272_ | ~new_A2273_;
  assign new_A2264_ = A2248 ^ new_A2255_;
  assign new_A2265_ = new_A2274_ & new_A2267_;
  assign new_A2266_ = ~new_A2276_ | ~new_A2275_;
  assign new_A2267_ = A2248 | A2249;
  assign new_A2268_ = A2248 | new_A2255_;
  assign new_A2269_ = A2247 & new_A2259_;
  assign new_A2270_ = ~A2246 | ~A2247;
  assign new_A2271_ = new_A2255_ & new_A2270_;
  assign new_A2272_ = ~new_A2271_ & ~new_A2255_;
  assign new_A2273_ = new_A2255_ | new_A2270_;
  assign new_A2274_ = ~A2248 | ~A2249;
  assign new_A2275_ = new_A2255_ | new_A2270_;
  assign new_A2276_ = ~new_A2255_ & ~new_A2277_;
  assign new_A2277_ = new_A2255_ & new_A2270_;
  assign new_A2283_ = new_A2289_ & new_A2288_;
  assign new_A2284_ = new_A2291_ | new_A2290_;
  assign new_A2285_ = new_A2293_ | new_A2292_;
  assign new_A2286_ = new_A2288_ & new_A2294_;
  assign new_A2287_ = new_A2288_ & new_A2295_;
  assign new_A2288_ = A2278 ^ A2279;
  assign new_A2289_ = new_A2290_ ^ A2280;
  assign new_A2290_ = new_A2298_ & new_A2297_;
  assign new_A2291_ = new_A2296_ & A2280;
  assign new_A2292_ = new_A2301_ & new_A2300_;
  assign new_A2293_ = new_A2299_ & A2280;
  assign new_A2294_ = new_A2302_ | A2279;
  assign new_A2295_ = ~A2280 ^ new_A2292_;
  assign new_A2296_ = ~new_A2305_ | ~new_A2306_;
  assign new_A2297_ = A2281 ^ new_A2288_;
  assign new_A2298_ = new_A2307_ & new_A2300_;
  assign new_A2299_ = ~new_A2309_ | ~new_A2308_;
  assign new_A2300_ = A2281 | A2282;
  assign new_A2301_ = A2281 | new_A2288_;
  assign new_A2302_ = A2280 & new_A2292_;
  assign new_A2303_ = ~A2279 | ~A2280;
  assign new_A2304_ = new_A2288_ & new_A2303_;
  assign new_A2305_ = ~new_A2304_ & ~new_A2288_;
  assign new_A2306_ = new_A2288_ | new_A2303_;
  assign new_A2307_ = ~A2281 | ~A2282;
  assign new_A2308_ = new_A2288_ | new_A2303_;
  assign new_A2309_ = ~new_A2288_ & ~new_A2310_;
  assign new_A2310_ = new_A2288_ & new_A2303_;
  assign new_A2316_ = new_A2322_ & new_A2321_;
  assign new_A2317_ = new_A2324_ | new_A2323_;
  assign new_A2318_ = new_A2326_ | new_A2325_;
  assign new_A2319_ = new_A2321_ & new_A2327_;
  assign new_A2320_ = new_A2321_ & new_A2328_;
  assign new_A2321_ = A2311 ^ A2312;
  assign new_A2322_ = new_A2323_ ^ A2313;
  assign new_A2323_ = new_A2331_ & new_A2330_;
  assign new_A2324_ = new_A2329_ & A2313;
  assign new_A2325_ = new_A2334_ & new_A2333_;
  assign new_A2326_ = new_A2332_ & A2313;
  assign new_A2327_ = new_A2335_ | A2312;
  assign new_A2328_ = ~A2313 ^ new_A2325_;
  assign new_A2329_ = ~new_A2338_ | ~new_A2339_;
  assign new_A2330_ = A2314 ^ new_A2321_;
  assign new_A2331_ = new_A2340_ & new_A2333_;
  assign new_A2332_ = ~new_A2342_ | ~new_A2341_;
  assign new_A2333_ = A2314 | A2315;
  assign new_A2334_ = A2314 | new_A2321_;
  assign new_A2335_ = A2313 & new_A2325_;
  assign new_A2336_ = ~A2312 | ~A2313;
  assign new_A2337_ = new_A2321_ & new_A2336_;
  assign new_A2338_ = ~new_A2337_ & ~new_A2321_;
  assign new_A2339_ = new_A2321_ | new_A2336_;
  assign new_A2340_ = ~A2314 | ~A2315;
  assign new_A2341_ = new_A2321_ | new_A2336_;
  assign new_A2342_ = ~new_A2321_ & ~new_A2343_;
  assign new_A2343_ = new_A2321_ & new_A2336_;
  assign new_A2349_ = new_A2355_ & new_A2354_;
  assign new_A2350_ = new_A2357_ | new_A2356_;
  assign new_A2351_ = new_A2359_ | new_A2358_;
  assign new_A2352_ = new_A2354_ & new_A2360_;
  assign new_A2353_ = new_A2354_ & new_A2361_;
  assign new_A2354_ = A2344 ^ A2345;
  assign new_A2355_ = new_A2356_ ^ A2346;
  assign new_A2356_ = new_A2364_ & new_A2363_;
  assign new_A2357_ = new_A2362_ & A2346;
  assign new_A2358_ = new_A2367_ & new_A2366_;
  assign new_A2359_ = new_A2365_ & A2346;
  assign new_A2360_ = new_A2368_ | A2345;
  assign new_A2361_ = ~A2346 ^ new_A2358_;
  assign new_A2362_ = ~new_A2371_ | ~new_A2372_;
  assign new_A2363_ = A2347 ^ new_A2354_;
  assign new_A2364_ = new_A2373_ & new_A2366_;
  assign new_A2365_ = ~new_A2375_ | ~new_A2374_;
  assign new_A2366_ = A2347 | A2348;
  assign new_A2367_ = A2347 | new_A2354_;
  assign new_A2368_ = A2346 & new_A2358_;
  assign new_A2369_ = ~A2345 | ~A2346;
  assign new_A2370_ = new_A2354_ & new_A2369_;
  assign new_A2371_ = ~new_A2370_ & ~new_A2354_;
  assign new_A2372_ = new_A2354_ | new_A2369_;
  assign new_A2373_ = ~A2347 | ~A2348;
  assign new_A2374_ = new_A2354_ | new_A2369_;
  assign new_A2375_ = ~new_A2354_ & ~new_A2376_;
  assign new_A2376_ = new_A2354_ & new_A2369_;
  assign new_A2382_ = new_A2388_ & new_A2387_;
  assign new_A2383_ = new_A2390_ | new_A2389_;
  assign new_A2384_ = new_A2392_ | new_A2391_;
  assign new_A2385_ = new_A2387_ & new_A2393_;
  assign new_A2386_ = new_A2387_ & new_A2394_;
  assign new_A2387_ = A2377 ^ A2378;
  assign new_A2388_ = new_A2389_ ^ A2379;
  assign new_A2389_ = new_A2397_ & new_A2396_;
  assign new_A2390_ = new_A2395_ & A2379;
  assign new_A2391_ = new_A2400_ & new_A2399_;
  assign new_A2392_ = new_A2398_ & A2379;
  assign new_A2393_ = new_A2401_ | A2378;
  assign new_A2394_ = ~A2379 ^ new_A2391_;
  assign new_A2395_ = ~new_A2404_ | ~new_A2405_;
  assign new_A2396_ = A2380 ^ new_A2387_;
  assign new_A2397_ = new_A2406_ & new_A2399_;
  assign new_A2398_ = ~new_A2408_ | ~new_A2407_;
  assign new_A2399_ = A2380 | A2381;
  assign new_A2400_ = A2380 | new_A2387_;
  assign new_A2401_ = A2379 & new_A2391_;
  assign new_A2402_ = ~A2378 | ~A2379;
  assign new_A2403_ = new_A2387_ & new_A2402_;
  assign new_A2404_ = ~new_A2403_ & ~new_A2387_;
  assign new_A2405_ = new_A2387_ | new_A2402_;
  assign new_A2406_ = ~A2380 | ~A2381;
  assign new_A2407_ = new_A2387_ | new_A2402_;
  assign new_A2408_ = ~new_A2387_ & ~new_A2409_;
  assign new_A2409_ = new_A2387_ & new_A2402_;
  assign new_A2415_ = new_A2421_ & new_A2420_;
  assign new_A2416_ = new_A2423_ | new_A2422_;
  assign new_A2417_ = new_A2425_ | new_A2424_;
  assign new_A2418_ = new_A2420_ & new_A2426_;
  assign new_A2419_ = new_A2420_ & new_A2427_;
  assign new_A2420_ = A2410 ^ A2411;
  assign new_A2421_ = new_A2422_ ^ A2412;
  assign new_A2422_ = new_A2430_ & new_A2429_;
  assign new_A2423_ = new_A2428_ & A2412;
  assign new_A2424_ = new_A2433_ & new_A2432_;
  assign new_A2425_ = new_A2431_ & A2412;
  assign new_A2426_ = new_A2434_ | A2411;
  assign new_A2427_ = ~A2412 ^ new_A2424_;
  assign new_A2428_ = ~new_A2437_ | ~new_A2438_;
  assign new_A2429_ = A2413 ^ new_A2420_;
  assign new_A2430_ = new_A2439_ & new_A2432_;
  assign new_A2431_ = ~new_A2441_ | ~new_A2440_;
  assign new_A2432_ = A2413 | A2414;
  assign new_A2433_ = A2413 | new_A2420_;
  assign new_A2434_ = A2412 & new_A2424_;
  assign new_A2435_ = ~A2411 | ~A2412;
  assign new_A2436_ = new_A2420_ & new_A2435_;
  assign new_A2437_ = ~new_A2436_ & ~new_A2420_;
  assign new_A2438_ = new_A2420_ | new_A2435_;
  assign new_A2439_ = ~A2413 | ~A2414;
  assign new_A2440_ = new_A2420_ | new_A2435_;
  assign new_A2441_ = ~new_A2420_ & ~new_A2442_;
  assign new_A2442_ = new_A2420_ & new_A2435_;
  assign new_A2448_ = new_A2454_ & new_A2453_;
  assign new_A2449_ = new_A2456_ | new_A2455_;
  assign new_A2450_ = new_A2458_ | new_A2457_;
  assign new_A2451_ = new_A2453_ & new_A2459_;
  assign new_A2452_ = new_A2453_ & new_A2460_;
  assign new_A2453_ = A2443 ^ A2444;
  assign new_A2454_ = new_A2455_ ^ A2445;
  assign new_A2455_ = new_A2463_ & new_A2462_;
  assign new_A2456_ = new_A2461_ & A2445;
  assign new_A2457_ = new_A2466_ & new_A2465_;
  assign new_A2458_ = new_A2464_ & A2445;
  assign new_A2459_ = new_A2467_ | A2444;
  assign new_A2460_ = ~A2445 ^ new_A2457_;
  assign new_A2461_ = ~new_A2470_ | ~new_A2471_;
  assign new_A2462_ = A2446 ^ new_A2453_;
  assign new_A2463_ = new_A2472_ & new_A2465_;
  assign new_A2464_ = ~new_A2474_ | ~new_A2473_;
  assign new_A2465_ = A2446 | A2447;
  assign new_A2466_ = A2446 | new_A2453_;
  assign new_A2467_ = A2445 & new_A2457_;
  assign new_A2468_ = ~A2444 | ~A2445;
  assign new_A2469_ = new_A2453_ & new_A2468_;
  assign new_A2470_ = ~new_A2469_ & ~new_A2453_;
  assign new_A2471_ = new_A2453_ | new_A2468_;
  assign new_A2472_ = ~A2446 | ~A2447;
  assign new_A2473_ = new_A2453_ | new_A2468_;
  assign new_A2474_ = ~new_A2453_ & ~new_A2475_;
  assign new_A2475_ = new_A2453_ & new_A2468_;
  assign new_A2481_ = new_A2487_ & new_A2486_;
  assign new_A2482_ = new_A2489_ | new_A2488_;
  assign new_A2483_ = new_A2491_ | new_A2490_;
  assign new_A2484_ = new_A2486_ & new_A2492_;
  assign new_A2485_ = new_A2486_ & new_A2493_;
  assign new_A2486_ = A2476 ^ A2477;
  assign new_A2487_ = new_A2488_ ^ A2478;
  assign new_A2488_ = new_A2496_ & new_A2495_;
  assign new_A2489_ = new_A2494_ & A2478;
  assign new_A2490_ = new_A2499_ & new_A2498_;
  assign new_A2491_ = new_A2497_ & A2478;
  assign new_A2492_ = new_A2500_ | A2477;
  assign new_A2493_ = ~A2478 ^ new_A2490_;
  assign new_A2494_ = ~new_A2503_ | ~new_A2504_;
  assign new_A2495_ = A2479 ^ new_A2486_;
  assign new_A2496_ = new_A2505_ & new_A2498_;
  assign new_A2497_ = ~new_A2507_ | ~new_A2506_;
  assign new_A2498_ = A2479 | A2480;
  assign new_A2499_ = A2479 | new_A2486_;
  assign new_A2500_ = A2478 & new_A2490_;
  assign new_A2501_ = ~A2477 | ~A2478;
  assign new_A2502_ = new_A2486_ & new_A2501_;
  assign new_A2503_ = ~new_A2502_ & ~new_A2486_;
  assign new_A2504_ = new_A2486_ | new_A2501_;
  assign new_A2505_ = ~A2479 | ~A2480;
  assign new_A2506_ = new_A2486_ | new_A2501_;
  assign new_A2507_ = ~new_A2486_ & ~new_A2508_;
  assign new_A2508_ = new_A2486_ & new_A2501_;
  assign new_A2514_ = new_A2520_ & new_A2519_;
  assign new_A2515_ = new_A2522_ | new_A2521_;
  assign new_A2516_ = new_A2524_ | new_A2523_;
  assign new_A2517_ = new_A2519_ & new_A2525_;
  assign new_A2518_ = new_A2519_ & new_A2526_;
  assign new_A2519_ = A2509 ^ A2510;
  assign new_A2520_ = new_A2521_ ^ A2511;
  assign new_A2521_ = new_A2529_ & new_A2528_;
  assign new_A2522_ = new_A2527_ & A2511;
  assign new_A2523_ = new_A2532_ & new_A2531_;
  assign new_A2524_ = new_A2530_ & A2511;
  assign new_A2525_ = new_A2533_ | A2510;
  assign new_A2526_ = ~A2511 ^ new_A2523_;
  assign new_A2527_ = ~new_A2536_ | ~new_A2537_;
  assign new_A2528_ = A2512 ^ new_A2519_;
  assign new_A2529_ = new_A2538_ & new_A2531_;
  assign new_A2530_ = ~new_A2540_ | ~new_A2539_;
  assign new_A2531_ = A2512 | A2513;
  assign new_A2532_ = A2512 | new_A2519_;
  assign new_A2533_ = A2511 & new_A2523_;
  assign new_A2534_ = ~A2510 | ~A2511;
  assign new_A2535_ = new_A2519_ & new_A2534_;
  assign new_A2536_ = ~new_A2535_ & ~new_A2519_;
  assign new_A2537_ = new_A2519_ | new_A2534_;
  assign new_A2538_ = ~A2512 | ~A2513;
  assign new_A2539_ = new_A2519_ | new_A2534_;
  assign new_A2540_ = ~new_A2519_ & ~new_A2541_;
  assign new_A2541_ = new_A2519_ & new_A2534_;
  assign new_A2547_ = new_A2553_ & new_A2552_;
  assign new_A2548_ = new_A2555_ | new_A2554_;
  assign new_A2549_ = new_A2557_ | new_A2556_;
  assign new_A2550_ = new_A2552_ & new_A2558_;
  assign new_A2551_ = new_A2552_ & new_A2559_;
  assign new_A2552_ = A2542 ^ A2543;
  assign new_A2553_ = new_A2554_ ^ A2544;
  assign new_A2554_ = new_A2562_ & new_A2561_;
  assign new_A2555_ = new_A2560_ & A2544;
  assign new_A2556_ = new_A2565_ & new_A2564_;
  assign new_A2557_ = new_A2563_ & A2544;
  assign new_A2558_ = new_A2566_ | A2543;
  assign new_A2559_ = ~A2544 ^ new_A2556_;
  assign new_A2560_ = ~new_A2569_ | ~new_A2570_;
  assign new_A2561_ = A2545 ^ new_A2552_;
  assign new_A2562_ = new_A2571_ & new_A2564_;
  assign new_A2563_ = ~new_A2573_ | ~new_A2572_;
  assign new_A2564_ = A2545 | A2546;
  assign new_A2565_ = A2545 | new_A2552_;
  assign new_A2566_ = A2544 & new_A2556_;
  assign new_A2567_ = ~A2543 | ~A2544;
  assign new_A2568_ = new_A2552_ & new_A2567_;
  assign new_A2569_ = ~new_A2568_ & ~new_A2552_;
  assign new_A2570_ = new_A2552_ | new_A2567_;
  assign new_A2571_ = ~A2545 | ~A2546;
  assign new_A2572_ = new_A2552_ | new_A2567_;
  assign new_A2573_ = ~new_A2552_ & ~new_A2574_;
  assign new_A2574_ = new_A2552_ & new_A2567_;
  assign new_A2580_ = new_A2586_ & new_A2585_;
  assign new_A2581_ = new_A2588_ | new_A2587_;
  assign new_A2582_ = new_A2590_ | new_A2589_;
  assign new_A2583_ = new_A2585_ & new_A2591_;
  assign new_A2584_ = new_A2585_ & new_A2592_;
  assign new_A2585_ = A2575 ^ A2576;
  assign new_A2586_ = new_A2587_ ^ A2577;
  assign new_A2587_ = new_A2595_ & new_A2594_;
  assign new_A2588_ = new_A2593_ & A2577;
  assign new_A2589_ = new_A2598_ & new_A2597_;
  assign new_A2590_ = new_A2596_ & A2577;
  assign new_A2591_ = new_A2599_ | A2576;
  assign new_A2592_ = ~A2577 ^ new_A2589_;
  assign new_A2593_ = ~new_A2602_ | ~new_A2603_;
  assign new_A2594_ = A2578 ^ new_A2585_;
  assign new_A2595_ = new_A2604_ & new_A2597_;
  assign new_A2596_ = ~new_A2606_ | ~new_A2605_;
  assign new_A2597_ = A2578 | A2579;
  assign new_A2598_ = A2578 | new_A2585_;
  assign new_A2599_ = A2577 & new_A2589_;
  assign new_A2600_ = ~A2576 | ~A2577;
  assign new_A2601_ = new_A2585_ & new_A2600_;
  assign new_A2602_ = ~new_A2601_ & ~new_A2585_;
  assign new_A2603_ = new_A2585_ | new_A2600_;
  assign new_A2604_ = ~A2578 | ~A2579;
  assign new_A2605_ = new_A2585_ | new_A2600_;
  assign new_A2606_ = ~new_A2585_ & ~new_A2607_;
  assign new_A2607_ = new_A2585_ & new_A2600_;
  assign new_A2613_ = new_A2619_ & new_A2618_;
  assign new_A2614_ = new_A2621_ | new_A2620_;
  assign new_A2615_ = new_A2623_ | new_A2622_;
  assign new_A2616_ = new_A2618_ & new_A2624_;
  assign new_A2617_ = new_A2618_ & new_A2625_;
  assign new_A2618_ = A2608 ^ A2609;
  assign new_A2619_ = new_A2620_ ^ A2610;
  assign new_A2620_ = new_A2628_ & new_A2627_;
  assign new_A2621_ = new_A2626_ & A2610;
  assign new_A2622_ = new_A2631_ & new_A2630_;
  assign new_A2623_ = new_A2629_ & A2610;
  assign new_A2624_ = new_A2632_ | A2609;
  assign new_A2625_ = ~A2610 ^ new_A2622_;
  assign new_A2626_ = ~new_A2635_ | ~new_A2636_;
  assign new_A2627_ = A2611 ^ new_A2618_;
  assign new_A2628_ = new_A2637_ & new_A2630_;
  assign new_A2629_ = ~new_A2639_ | ~new_A2638_;
  assign new_A2630_ = A2611 | A2612;
  assign new_A2631_ = A2611 | new_A2618_;
  assign new_A2632_ = A2610 & new_A2622_;
  assign new_A2633_ = ~A2609 | ~A2610;
  assign new_A2634_ = new_A2618_ & new_A2633_;
  assign new_A2635_ = ~new_A2634_ & ~new_A2618_;
  assign new_A2636_ = new_A2618_ | new_A2633_;
  assign new_A2637_ = ~A2611 | ~A2612;
  assign new_A2638_ = new_A2618_ | new_A2633_;
  assign new_A2639_ = ~new_A2618_ & ~new_A2640_;
  assign new_A2640_ = new_A2618_ & new_A2633_;
  assign new_A2646_ = new_A2652_ & new_A2651_;
  assign new_A2647_ = new_A2654_ | new_A2653_;
  assign new_A2648_ = new_A2656_ | new_A2655_;
  assign new_A2649_ = new_A2651_ & new_A2657_;
  assign new_A2650_ = new_A2651_ & new_A2658_;
  assign new_A2651_ = A2641 ^ A2642;
  assign new_A2652_ = new_A2653_ ^ A2643;
  assign new_A2653_ = new_A2661_ & new_A2660_;
  assign new_A2654_ = new_A2659_ & A2643;
  assign new_A2655_ = new_A2664_ & new_A2663_;
  assign new_A2656_ = new_A2662_ & A2643;
  assign new_A2657_ = new_A2665_ | A2642;
  assign new_A2658_ = ~A2643 ^ new_A2655_;
  assign new_A2659_ = ~new_A2668_ | ~new_A2669_;
  assign new_A2660_ = A2644 ^ new_A2651_;
  assign new_A2661_ = new_A2670_ & new_A2663_;
  assign new_A2662_ = ~new_A2672_ | ~new_A2671_;
  assign new_A2663_ = A2644 | A2645;
  assign new_A2664_ = A2644 | new_A2651_;
  assign new_A2665_ = A2643 & new_A2655_;
  assign new_A2666_ = ~A2642 | ~A2643;
  assign new_A2667_ = new_A2651_ & new_A2666_;
  assign new_A2668_ = ~new_A2667_ & ~new_A2651_;
  assign new_A2669_ = new_A2651_ | new_A2666_;
  assign new_A2670_ = ~A2644 | ~A2645;
  assign new_A2671_ = new_A2651_ | new_A2666_;
  assign new_A2672_ = ~new_A2651_ & ~new_A2673_;
  assign new_A2673_ = new_A2651_ & new_A2666_;
  assign new_A2679_ = new_A2685_ & new_A2684_;
  assign new_A2680_ = new_A2687_ | new_A2686_;
  assign new_A2681_ = new_A2689_ | new_A2688_;
  assign new_A2682_ = new_A2684_ & new_A2690_;
  assign new_A2683_ = new_A2684_ & new_A2691_;
  assign new_A2684_ = A2674 ^ A2675;
  assign new_A2685_ = new_A2686_ ^ A2676;
  assign new_A2686_ = new_A2694_ & new_A2693_;
  assign new_A2687_ = new_A2692_ & A2676;
  assign new_A2688_ = new_A2697_ & new_A2696_;
  assign new_A2689_ = new_A2695_ & A2676;
  assign new_A2690_ = new_A2698_ | A2675;
  assign new_A2691_ = ~A2676 ^ new_A2688_;
  assign new_A2692_ = ~new_A2701_ | ~new_A2702_;
  assign new_A2693_ = A2677 ^ new_A2684_;
  assign new_A2694_ = new_A2703_ & new_A2696_;
  assign new_A2695_ = ~new_A2705_ | ~new_A2704_;
  assign new_A2696_ = A2677 | A2678;
  assign new_A2697_ = A2677 | new_A2684_;
  assign new_A2698_ = A2676 & new_A2688_;
  assign new_A2699_ = ~A2675 | ~A2676;
  assign new_A2700_ = new_A2684_ & new_A2699_;
  assign new_A2701_ = ~new_A2700_ & ~new_A2684_;
  assign new_A2702_ = new_A2684_ | new_A2699_;
  assign new_A2703_ = ~A2677 | ~A2678;
  assign new_A2704_ = new_A2684_ | new_A2699_;
  assign new_A2705_ = ~new_A2684_ & ~new_A2706_;
  assign new_A2706_ = new_A2684_ & new_A2699_;
  assign new_A2712_ = new_A2718_ & new_A2717_;
  assign new_A2713_ = new_A2720_ | new_A2719_;
  assign new_A2714_ = new_A2722_ | new_A2721_;
  assign new_A2715_ = new_A2717_ & new_A2723_;
  assign new_A2716_ = new_A2717_ & new_A2724_;
  assign new_A2717_ = A2707 ^ A2708;
  assign new_A2718_ = new_A2719_ ^ A2709;
  assign new_A2719_ = new_A2727_ & new_A2726_;
  assign new_A2720_ = new_A2725_ & A2709;
  assign new_A2721_ = new_A2730_ & new_A2729_;
  assign new_A2722_ = new_A2728_ & A2709;
  assign new_A2723_ = new_A2731_ | A2708;
  assign new_A2724_ = ~A2709 ^ new_A2721_;
  assign new_A2725_ = ~new_A2734_ | ~new_A2735_;
  assign new_A2726_ = A2710 ^ new_A2717_;
  assign new_A2727_ = new_A2736_ & new_A2729_;
  assign new_A2728_ = ~new_A2738_ | ~new_A2737_;
  assign new_A2729_ = A2710 | A2711;
  assign new_A2730_ = A2710 | new_A2717_;
  assign new_A2731_ = A2709 & new_A2721_;
  assign new_A2732_ = ~A2708 | ~A2709;
  assign new_A2733_ = new_A2717_ & new_A2732_;
  assign new_A2734_ = ~new_A2733_ & ~new_A2717_;
  assign new_A2735_ = new_A2717_ | new_A2732_;
  assign new_A2736_ = ~A2710 | ~A2711;
  assign new_A2737_ = new_A2717_ | new_A2732_;
  assign new_A2738_ = ~new_A2717_ & ~new_A2739_;
  assign new_A2739_ = new_A2717_ & new_A2732_;
  assign new_A2745_ = new_A2751_ & new_A2750_;
  assign new_A2746_ = new_A2753_ | new_A2752_;
  assign new_A2747_ = new_A2755_ | new_A2754_;
  assign new_A2748_ = new_A2750_ & new_A2756_;
  assign new_A2749_ = new_A2750_ & new_A2757_;
  assign new_A2750_ = A2740 ^ A2741;
  assign new_A2751_ = new_A2752_ ^ A2742;
  assign new_A2752_ = new_A2760_ & new_A2759_;
  assign new_A2753_ = new_A2758_ & A2742;
  assign new_A2754_ = new_A2763_ & new_A2762_;
  assign new_A2755_ = new_A2761_ & A2742;
  assign new_A2756_ = new_A2764_ | A2741;
  assign new_A2757_ = ~A2742 ^ new_A2754_;
  assign new_A2758_ = ~new_A2767_ | ~new_A2768_;
  assign new_A2759_ = A2743 ^ new_A2750_;
  assign new_A2760_ = new_A2769_ & new_A2762_;
  assign new_A2761_ = ~new_A2771_ | ~new_A2770_;
  assign new_A2762_ = A2743 | A2744;
  assign new_A2763_ = A2743 | new_A2750_;
  assign new_A2764_ = A2742 & new_A2754_;
  assign new_A2765_ = ~A2741 | ~A2742;
  assign new_A2766_ = new_A2750_ & new_A2765_;
  assign new_A2767_ = ~new_A2766_ & ~new_A2750_;
  assign new_A2768_ = new_A2750_ | new_A2765_;
  assign new_A2769_ = ~A2743 | ~A2744;
  assign new_A2770_ = new_A2750_ | new_A2765_;
  assign new_A2771_ = ~new_A2750_ & ~new_A2772_;
  assign new_A2772_ = new_A2750_ & new_A2765_;
  assign new_A2778_ = new_A2784_ & new_A2783_;
  assign new_A2779_ = new_A2786_ | new_A2785_;
  assign new_A2780_ = new_A2788_ | new_A2787_;
  assign new_A2781_ = new_A2783_ & new_A2789_;
  assign new_A2782_ = new_A2783_ & new_A2790_;
  assign new_A2783_ = A2773 ^ A2774;
  assign new_A2784_ = new_A2785_ ^ A2775;
  assign new_A2785_ = new_A2793_ & new_A2792_;
  assign new_A2786_ = new_A2791_ & A2775;
  assign new_A2787_ = new_A2796_ & new_A2795_;
  assign new_A2788_ = new_A2794_ & A2775;
  assign new_A2789_ = new_A2797_ | A2774;
  assign new_A2790_ = ~A2775 ^ new_A2787_;
  assign new_A2791_ = ~new_A2800_ | ~new_A2801_;
  assign new_A2792_ = A2776 ^ new_A2783_;
  assign new_A2793_ = new_A2802_ & new_A2795_;
  assign new_A2794_ = ~new_A2804_ | ~new_A2803_;
  assign new_A2795_ = A2776 | A2777;
  assign new_A2796_ = A2776 | new_A2783_;
  assign new_A2797_ = A2775 & new_A2787_;
  assign new_A2798_ = ~A2774 | ~A2775;
  assign new_A2799_ = new_A2783_ & new_A2798_;
  assign new_A2800_ = ~new_A2799_ & ~new_A2783_;
  assign new_A2801_ = new_A2783_ | new_A2798_;
  assign new_A2802_ = ~A2776 | ~A2777;
  assign new_A2803_ = new_A2783_ | new_A2798_;
  assign new_A2804_ = ~new_A2783_ & ~new_A2805_;
  assign new_A2805_ = new_A2783_ & new_A2798_;
  assign new_A1188_ = new_A1166_ & new_A1181_;
  assign new_A1187_ = ~new_A1166_ & ~new_A1188_;
  assign new_A1186_ = new_A1166_ | new_A1181_;
  assign new_A1185_ = ~new_A1159_ | ~new_A1160_;
  assign new_A1184_ = new_A1166_ | new_A1181_;
  assign new_A1183_ = ~new_A1182_ & ~new_A1166_;
  assign new_A1182_ = new_A1166_ & new_A1181_;
  assign new_A1181_ = ~new_A1157_ | ~new_A1158_;
  assign new_A1180_ = new_A1158_ & new_A1170_;
  assign new_A1179_ = new_A1159_ | new_A1166_;
  assign new_A1178_ = new_A1159_ | new_A1160_;
  assign new_A1177_ = ~new_A1187_ | ~new_A1186_;
  assign new_A1176_ = new_A1185_ & new_A1178_;
  assign new_A1175_ = new_A1159_ ^ new_A1166_;
  assign new_A1174_ = ~new_A1183_ | ~new_A1184_;
  assign new_A1173_ = ~new_A1158_ ^ new_A1170_;
  assign new_A1172_ = new_A1180_ | new_A1157_;
  assign new_A1171_ = new_A1177_ & new_A1158_;
  assign new_A1170_ = new_A1179_ & new_A1178_;
  assign new_A1169_ = new_A1174_ & new_A1158_;
  assign new_A1168_ = new_A1176_ & new_A1175_;
  assign new_A1167_ = new_A1168_ ^ new_A1158_;
  assign new_A1166_ = new_A1156_ ^ new_A1157_;
  assign new_A1165_ = new_A1166_ & new_A1173_;
  assign new_A1164_ = new_A1166_ & new_A1172_;
  assign new_A1163_ = new_A1171_ | new_A1170_;
  assign new_A1162_ = new_A1169_ | new_A1168_;
  assign new_A1161_ = new_A1167_ & new_A1166_;
  assign new_A1160_ = new_A1990_;
  assign new_A1159_ = new_A2019_;
  assign new_A1158_ = new_A2052_;
  assign new_A1157_ = new_A2085_;
  assign new_A1156_ = new_A2118_;
  assign new_A1189_ = new_A2151_;
  assign new_A1190_ = new_A2184_;
  assign new_A1191_ = new_A2217_;
  assign new_A1192_ = new_A2250_;
  assign new_A1193_ = new_A2283_;
  assign new_A1194_ = new_A1200_ & new_A1199_;
  assign new_A1195_ = new_A1202_ | new_A1201_;
  assign new_A1196_ = new_A1204_ | new_A1203_;
  assign new_A1197_ = new_A1199_ & new_A1205_;
  assign new_A1198_ = new_A1199_ & new_A1206_;
  assign new_A1199_ = new_A1189_ ^ new_A1190_;
  assign new_A1200_ = new_A1201_ ^ new_A1191_;
  assign new_A1201_ = new_A1209_ & new_A1208_;
  assign new_A1202_ = new_A1207_ & new_A1191_;
  assign new_A1203_ = new_A1212_ & new_A1211_;
  assign new_A1204_ = new_A1210_ & new_A1191_;
  assign new_A1205_ = new_A1213_ | new_A1190_;
  assign new_A1206_ = ~new_A1191_ ^ new_A1203_;
  assign new_A1207_ = ~new_A1216_ | ~new_A1217_;
  assign new_A1208_ = new_A1192_ ^ new_A1199_;
  assign new_A1209_ = new_A1218_ & new_A1211_;
  assign new_A1210_ = ~new_A1220_ | ~new_A1219_;
  assign new_A1211_ = new_A1192_ | new_A1193_;
  assign new_A1212_ = new_A1192_ | new_A1199_;
  assign new_A1213_ = new_A1191_ & new_A1203_;
  assign new_A1214_ = ~new_A1190_ | ~new_A1191_;
  assign new_A1215_ = new_A1199_ & new_A1214_;
  assign new_A1216_ = ~new_A1215_ & ~new_A1199_;
  assign new_A1217_ = new_A1199_ | new_A1214_;
  assign new_A1218_ = ~new_A1192_ | ~new_A1193_;
  assign new_A1219_ = new_A1199_ | new_A1214_;
  assign new_A1220_ = ~new_A1199_ & ~new_A1221_;
  assign new_A1221_ = new_A1199_ & new_A1214_;
  assign new_A1222_ = new_A2316_;
  assign new_A1223_ = new_A2349_;
  assign new_A1224_ = new_A2382_;
  assign new_A1225_ = new_A2415_;
  assign new_A1226_ = new_A2448_;
  assign new_A1227_ = new_A1233_ & new_A1232_;
  assign new_A1228_ = new_A1235_ | new_A1234_;
  assign new_A1229_ = new_A1237_ | new_A1236_;
  assign new_A1230_ = new_A1232_ & new_A1238_;
  assign new_A1231_ = new_A1232_ & new_A1239_;
  assign new_A1232_ = new_A1222_ ^ new_A1223_;
  assign new_A1233_ = new_A1234_ ^ new_A1224_;
  assign new_A1234_ = new_A1242_ & new_A1241_;
  assign new_A1235_ = new_A1240_ & new_A1224_;
  assign new_A1236_ = new_A1245_ & new_A1244_;
  assign new_A1237_ = new_A1243_ & new_A1224_;
  assign new_A1238_ = new_A1246_ | new_A1223_;
  assign new_A1239_ = ~new_A1224_ ^ new_A1236_;
  assign new_A1240_ = ~new_A1249_ | ~new_A1250_;
  assign new_A1241_ = new_A1225_ ^ new_A1232_;
  assign new_A1242_ = new_A1251_ & new_A1244_;
  assign new_A1243_ = ~new_A1253_ | ~new_A1252_;
  assign new_A1244_ = new_A1225_ | new_A1226_;
  assign new_A1245_ = new_A1225_ | new_A1232_;
  assign new_A1246_ = new_A1224_ & new_A1236_;
  assign new_A1247_ = ~new_A1223_ | ~new_A1224_;
  assign new_A1248_ = new_A1232_ & new_A1247_;
  assign new_A1249_ = ~new_A1248_ & ~new_A1232_;
  assign new_A1250_ = new_A1232_ | new_A1247_;
  assign new_A1251_ = ~new_A1225_ | ~new_A1226_;
  assign new_A1252_ = new_A1232_ | new_A1247_;
  assign new_A1253_ = ~new_A1232_ & ~new_A1254_;
  assign new_A1254_ = new_A1232_ & new_A1247_;
  assign new_A1255_ = new_A2481_;
  assign new_A1256_ = new_A2514_;
  assign new_A1257_ = new_A2547_;
  assign new_A1258_ = new_A2580_;
  assign new_A1259_ = new_A2613_;
  assign new_A1260_ = new_A1266_ & new_A1265_;
  assign new_A1261_ = new_A1268_ | new_A1267_;
  assign new_A1262_ = new_A1270_ | new_A1269_;
  assign new_A1263_ = new_A1265_ & new_A1271_;
  assign new_A1264_ = new_A1265_ & new_A1272_;
  assign new_A1265_ = new_A1255_ ^ new_A1256_;
  assign new_A1266_ = new_A1267_ ^ new_A1257_;
  assign new_A1267_ = new_A1275_ & new_A1274_;
  assign new_A1268_ = new_A1273_ & new_A1257_;
  assign new_A1269_ = new_A1278_ & new_A1277_;
  assign new_A1270_ = new_A1276_ & new_A1257_;
  assign new_A1271_ = new_A1279_ | new_A1256_;
  assign new_A1272_ = ~new_A1257_ ^ new_A1269_;
  assign new_A1273_ = ~new_A1282_ | ~new_A1283_;
  assign new_A1274_ = new_A1258_ ^ new_A1265_;
  assign new_A1275_ = new_A1284_ & new_A1277_;
  assign new_A1276_ = ~new_A1286_ | ~new_A1285_;
  assign new_A1277_ = new_A1258_ | new_A1259_;
  assign new_A1278_ = new_A1258_ | new_A1265_;
  assign new_A1279_ = new_A1257_ & new_A1269_;
  assign new_A1280_ = ~new_A1256_ | ~new_A1257_;
  assign new_A1281_ = new_A1265_ & new_A1280_;
  assign new_A1282_ = ~new_A1281_ & ~new_A1265_;
  assign new_A1283_ = new_A1265_ | new_A1280_;
  assign new_A1284_ = ~new_A1258_ | ~new_A1259_;
  assign new_A1285_ = new_A1265_ | new_A1280_;
  assign new_A1286_ = ~new_A1265_ & ~new_A1287_;
  assign new_A1287_ = new_A1265_ & new_A1280_;
  assign new_A1288_ = new_A2646_;
  assign new_A1289_ = new_A2679_;
  assign new_A1290_ = new_A2712_;
  assign new_A1291_ = new_A2745_;
  assign new_A1292_ = new_A2778_;
  assign new_A1293_ = new_A1299_ & new_A1298_;
  assign new_A1294_ = new_A1301_ | new_A1300_;
  assign new_A1295_ = new_A1303_ | new_A1302_;
  assign new_A1296_ = new_A1298_ & new_A1304_;
  assign new_A1297_ = new_A1298_ & new_A1305_;
  assign new_A1298_ = new_A1288_ ^ new_A1289_;
  assign new_A1299_ = new_A1300_ ^ new_A1290_;
  assign new_A1300_ = new_A1308_ & new_A1307_;
  assign new_A1301_ = new_A1306_ & new_A1290_;
  assign new_A1302_ = new_A1311_ & new_A1310_;
  assign new_A1303_ = new_A1309_ & new_A1290_;
  assign new_A1304_ = new_A1312_ | new_A1289_;
  assign new_A1305_ = ~new_A1290_ ^ new_A1302_;
  assign new_A1306_ = ~new_A1315_ | ~new_A1316_;
  assign new_A1307_ = new_A1291_ ^ new_A1298_;
  assign new_A1308_ = new_A1317_ & new_A1310_;
  assign new_A1309_ = ~new_A1319_ | ~new_A1318_;
  assign new_A1310_ = new_A1291_ | new_A1292_;
  assign new_A1311_ = new_A1291_ | new_A1298_;
  assign new_A1312_ = new_A1290_ & new_A1302_;
  assign new_A1313_ = ~new_A1289_ | ~new_A1290_;
  assign new_A1314_ = new_A1298_ & new_A1313_;
  assign new_A1315_ = ~new_A1314_ & ~new_A1298_;
  assign new_A1316_ = new_A1298_ | new_A1313_;
  assign new_A1317_ = ~new_A1291_ | ~new_A1292_;
  assign new_A1318_ = new_A1298_ | new_A1313_;
  assign new_A1319_ = ~new_A1298_ & ~new_A1320_;
  assign new_A1320_ = new_A1298_ & new_A1313_;
  assign new_A1321_ = new_A1989_;
  assign new_A1322_ = new_A2020_;
  assign new_A1323_ = new_A2053_;
  assign new_A1324_ = new_A2086_;
  assign new_A1325_ = new_A2119_;
  assign new_A1326_ = new_A1332_ & new_A1331_;
  assign new_A1327_ = new_A1334_ | new_A1333_;
  assign new_A1328_ = new_A1336_ | new_A1335_;
  assign new_A1329_ = new_A1331_ & new_A1337_;
  assign new_A1330_ = new_A1331_ & new_A1338_;
  assign new_A1331_ = new_A1321_ ^ new_A1322_;
  assign new_A1332_ = new_A1333_ ^ new_A1323_;
  assign new_A1333_ = new_A1341_ & new_A1340_;
  assign new_A1334_ = new_A1339_ & new_A1323_;
  assign new_A1335_ = new_A1344_ & new_A1343_;
  assign new_A1336_ = new_A1342_ & new_A1323_;
  assign new_A1337_ = new_A1345_ | new_A1322_;
  assign new_A1338_ = ~new_A1323_ ^ new_A1335_;
  assign new_A1339_ = ~new_A1348_ | ~new_A1349_;
  assign new_A1340_ = new_A1324_ ^ new_A1331_;
  assign new_A1341_ = new_A1350_ & new_A1343_;
  assign new_A1342_ = ~new_A1352_ | ~new_A1351_;
  assign new_A1343_ = new_A1324_ | new_A1325_;
  assign new_A1344_ = new_A1324_ | new_A1331_;
  assign new_A1345_ = new_A1323_ & new_A1335_;
  assign new_A1346_ = ~new_A1322_ | ~new_A1323_;
  assign new_A1347_ = new_A1331_ & new_A1346_;
  assign new_A1348_ = ~new_A1347_ & ~new_A1331_;
  assign new_A1349_ = new_A1331_ | new_A1346_;
  assign new_A1350_ = ~new_A1324_ | ~new_A1325_;
  assign new_A1351_ = new_A1331_ | new_A1346_;
  assign new_A1352_ = ~new_A1331_ & ~new_A1353_;
  assign new_A1353_ = new_A1331_ & new_A1346_;
  assign new_A1354_ = new_A2152_;
  assign new_A1355_ = new_A2185_;
  assign new_A1356_ = new_A2218_;
  assign new_A1357_ = new_A2251_;
  assign new_A1358_ = new_A2284_;
  assign new_A1359_ = new_A1365_ & new_A1364_;
  assign new_A1360_ = new_A1367_ | new_A1366_;
  assign new_A1361_ = new_A1369_ | new_A1368_;
  assign new_A1362_ = new_A1364_ & new_A1370_;
  assign new_A1363_ = new_A1364_ & new_A1371_;
  assign new_A1364_ = new_A1354_ ^ new_A1355_;
  assign new_A1365_ = new_A1366_ ^ new_A1356_;
  assign new_A1366_ = new_A1374_ & new_A1373_;
  assign new_A1367_ = new_A1372_ & new_A1356_;
  assign new_A1368_ = new_A1377_ & new_A1376_;
  assign new_A1369_ = new_A1375_ & new_A1356_;
  assign new_A1370_ = new_A1378_ | new_A1355_;
  assign new_A1371_ = ~new_A1356_ ^ new_A1368_;
  assign new_A1372_ = ~new_A1381_ | ~new_A1382_;
  assign new_A1373_ = new_A1357_ ^ new_A1364_;
  assign new_A1374_ = new_A1383_ & new_A1376_;
  assign new_A1375_ = ~new_A1385_ | ~new_A1384_;
  assign new_A1376_ = new_A1357_ | new_A1358_;
  assign new_A1377_ = new_A1357_ | new_A1364_;
  assign new_A1378_ = new_A1356_ & new_A1368_;
  assign new_A1379_ = ~new_A1355_ | ~new_A1356_;
  assign new_A1380_ = new_A1364_ & new_A1379_;
  assign new_A1381_ = ~new_A1380_ & ~new_A1364_;
  assign new_A1382_ = new_A1364_ | new_A1379_;
  assign new_A1383_ = ~new_A1357_ | ~new_A1358_;
  assign new_A1384_ = new_A1364_ | new_A1379_;
  assign new_A1385_ = ~new_A1364_ & ~new_A1386_;
  assign new_A1386_ = new_A1364_ & new_A1379_;
  assign new_A1387_ = new_A2317_;
  assign new_A1388_ = new_A2350_;
  assign new_A1389_ = new_A2383_;
  assign new_A1390_ = new_A2416_;
  assign new_A1391_ = new_A2449_;
  assign new_A1392_ = new_A1398_ & new_A1397_;
  assign new_A1393_ = new_A1400_ | new_A1399_;
  assign new_A1394_ = new_A1402_ | new_A1401_;
  assign new_A1395_ = new_A1397_ & new_A1403_;
  assign new_A1396_ = new_A1397_ & new_A1404_;
  assign new_A1397_ = new_A1387_ ^ new_A1388_;
  assign new_A1398_ = new_A1399_ ^ new_A1389_;
  assign new_A1399_ = new_A1407_ & new_A1406_;
  assign new_A1400_ = new_A1405_ & new_A1389_;
  assign new_A1401_ = new_A1410_ & new_A1409_;
  assign new_A1402_ = new_A1408_ & new_A1389_;
  assign new_A1403_ = new_A1411_ | new_A1388_;
  assign new_A1404_ = ~new_A1389_ ^ new_A1401_;
  assign new_A1405_ = ~new_A1414_ | ~new_A1415_;
  assign new_A1406_ = new_A1390_ ^ new_A1397_;
  assign new_A1407_ = new_A1416_ & new_A1409_;
  assign new_A1408_ = ~new_A1418_ | ~new_A1417_;
  assign new_A1409_ = new_A1390_ | new_A1391_;
  assign new_A1410_ = new_A1390_ | new_A1397_;
  assign new_A1411_ = new_A1389_ & new_A1401_;
  assign new_A1412_ = ~new_A1388_ | ~new_A1389_;
  assign new_A1413_ = new_A1397_ & new_A1412_;
  assign new_A1414_ = ~new_A1413_ & ~new_A1397_;
  assign new_A1415_ = new_A1397_ | new_A1412_;
  assign new_A1416_ = ~new_A1390_ | ~new_A1391_;
  assign new_A1417_ = new_A1397_ | new_A1412_;
  assign new_A1418_ = ~new_A1397_ & ~new_A1419_;
  assign new_A1419_ = new_A1397_ & new_A1412_;
  assign new_A1420_ = new_A2482_;
  assign new_A1421_ = new_A2515_;
  assign new_A1422_ = new_A2548_;
  assign new_A1423_ = new_A2581_;
  assign new_A1424_ = new_A2614_;
  assign new_A1425_ = new_A1431_ & new_A1430_;
  assign new_A1426_ = new_A1433_ | new_A1432_;
  assign new_A1427_ = new_A1435_ | new_A1434_;
  assign new_A1428_ = new_A1430_ & new_A1436_;
  assign new_A1429_ = new_A1430_ & new_A1437_;
  assign new_A1430_ = new_A1420_ ^ new_A1421_;
  assign new_A1431_ = new_A1432_ ^ new_A1422_;
  assign new_A1432_ = new_A1440_ & new_A1439_;
  assign new_A1433_ = new_A1438_ & new_A1422_;
  assign new_A1434_ = new_A1443_ & new_A1442_;
  assign new_A1435_ = new_A1441_ & new_A1422_;
  assign new_A1436_ = new_A1444_ | new_A1421_;
  assign new_A1437_ = ~new_A1422_ ^ new_A1434_;
  assign new_A1438_ = ~new_A1447_ | ~new_A1448_;
  assign new_A1439_ = new_A1423_ ^ new_A1430_;
  assign new_A1440_ = new_A1449_ & new_A1442_;
  assign new_A1441_ = ~new_A1451_ | ~new_A1450_;
  assign new_A1442_ = new_A1423_ | new_A1424_;
  assign new_A1443_ = new_A1423_ | new_A1430_;
  assign new_A1444_ = new_A1422_ & new_A1434_;
  assign new_A1445_ = ~new_A1421_ | ~new_A1422_;
  assign new_A1446_ = new_A1430_ & new_A1445_;
  assign new_A1447_ = ~new_A1446_ & ~new_A1430_;
  assign new_A1448_ = new_A1430_ | new_A1445_;
  assign new_A1449_ = ~new_A1423_ | ~new_A1424_;
  assign new_A1450_ = new_A1430_ | new_A1445_;
  assign new_A1451_ = ~new_A1430_ & ~new_A1452_;
  assign new_A1452_ = new_A1430_ & new_A1445_;
  assign new_A1453_ = new_A2647_;
  assign new_A1454_ = new_A2680_;
  assign new_A1455_ = new_A2713_;
  assign new_A1456_ = new_A2746_;
  assign new_A1457_ = new_A2779_;
  assign new_A1458_ = new_A1464_ & new_A1463_;
  assign new_A1459_ = new_A1466_ | new_A1465_;
  assign new_A1460_ = new_A1468_ | new_A1467_;
  assign new_A1461_ = new_A1463_ & new_A1469_;
  assign new_A1462_ = new_A1463_ & new_A1470_;
  assign new_A1463_ = new_A1453_ ^ new_A1454_;
  assign new_A1464_ = new_A1465_ ^ new_A1455_;
  assign new_A1465_ = new_A1473_ & new_A1472_;
  assign new_A1466_ = new_A1471_ & new_A1455_;
  assign new_A1467_ = new_A1476_ & new_A1475_;
  assign new_A1468_ = new_A1474_ & new_A1455_;
  assign new_A1469_ = new_A1477_ | new_A1454_;
  assign new_A1470_ = ~new_A1455_ ^ new_A1467_;
  assign new_A1471_ = ~new_A1480_ | ~new_A1481_;
  assign new_A1472_ = new_A1456_ ^ new_A1463_;
  assign new_A1473_ = new_A1482_ & new_A1475_;
  assign new_A1474_ = ~new_A1484_ | ~new_A1483_;
  assign new_A1475_ = new_A1456_ | new_A1457_;
  assign new_A1476_ = new_A1456_ | new_A1463_;
  assign new_A1477_ = new_A1455_ & new_A1467_;
  assign new_A1478_ = ~new_A1454_ | ~new_A1455_;
  assign new_A1479_ = new_A1463_ & new_A1478_;
  assign new_A1480_ = ~new_A1479_ & ~new_A1463_;
  assign new_A1481_ = new_A1463_ | new_A1478_;
  assign new_A1482_ = ~new_A1456_ | ~new_A1457_;
  assign new_A1483_ = new_A1463_ | new_A1478_;
  assign new_A1484_ = ~new_A1463_ & ~new_A1485_;
  assign new_A1485_ = new_A1463_ & new_A1478_;
  assign new_A1486_ = new_A1988_;
  assign new_A1487_ = new_A2021_;
  assign new_A1488_ = new_A2054_;
  assign new_A1489_ = new_A2087_;
  assign new_A1490_ = new_A2120_;
  assign new_A1491_ = new_A1497_ & new_A1496_;
  assign new_A1492_ = new_A1499_ | new_A1498_;
  assign new_A1493_ = new_A1501_ | new_A1500_;
  assign new_A1494_ = new_A1496_ & new_A1502_;
  assign new_A1495_ = new_A1496_ & new_A1503_;
  assign new_A1496_ = new_A1486_ ^ new_A1487_;
  assign new_A1497_ = new_A1498_ ^ new_A1488_;
  assign new_A1498_ = new_A1506_ & new_A1505_;
  assign new_A1499_ = new_A1504_ & new_A1488_;
  assign new_A1500_ = new_A1509_ & new_A1508_;
  assign new_A1501_ = new_A1507_ & new_A1488_;
  assign new_A1502_ = new_A1510_ | new_A1487_;
  assign new_A1503_ = ~new_A1488_ ^ new_A1500_;
  assign new_A1504_ = ~new_A1513_ | ~new_A1514_;
  assign new_A1505_ = new_A1489_ ^ new_A1496_;
  assign new_A1506_ = new_A1515_ & new_A1508_;
  assign new_A1507_ = ~new_A1517_ | ~new_A1516_;
  assign new_A1508_ = new_A1489_ | new_A1490_;
  assign new_A1509_ = new_A1489_ | new_A1496_;
  assign new_A1510_ = new_A1488_ & new_A1500_;
  assign new_A1511_ = ~new_A1487_ | ~new_A1488_;
  assign new_A1512_ = new_A1496_ & new_A1511_;
  assign new_A1513_ = ~new_A1512_ & ~new_A1496_;
  assign new_A1514_ = new_A1496_ | new_A1511_;
  assign new_A1515_ = ~new_A1489_ | ~new_A1490_;
  assign new_A1516_ = new_A1496_ | new_A1511_;
  assign new_A1517_ = ~new_A1496_ & ~new_A1518_;
  assign new_A1518_ = new_A1496_ & new_A1511_;
  assign new_A1519_ = new_A2153_;
  assign new_A1520_ = new_A2186_;
  assign new_A1521_ = new_A2219_;
  assign new_A1522_ = new_A2252_;
  assign new_A1523_ = new_A2285_;
  assign new_A1524_ = new_A1530_ & new_A1529_;
  assign new_A1525_ = new_A1532_ | new_A1531_;
  assign new_A1526_ = new_A1534_ | new_A1533_;
  assign new_A1527_ = new_A1529_ & new_A1535_;
  assign new_A1528_ = new_A1529_ & new_A1536_;
  assign new_A1529_ = new_A1519_ ^ new_A1520_;
  assign new_A1530_ = new_A1531_ ^ new_A1521_;
  assign new_A1531_ = new_A1539_ & new_A1538_;
  assign new_A1532_ = new_A1537_ & new_A1521_;
  assign new_A1533_ = new_A1542_ & new_A1541_;
  assign new_A1534_ = new_A1540_ & new_A1521_;
  assign new_A1535_ = new_A1543_ | new_A1520_;
  assign new_A1536_ = ~new_A1521_ ^ new_A1533_;
  assign new_A1537_ = ~new_A1546_ | ~new_A1547_;
  assign new_A1538_ = new_A1522_ ^ new_A1529_;
  assign new_A1539_ = new_A1548_ & new_A1541_;
  assign new_A1540_ = ~new_A1550_ | ~new_A1549_;
  assign new_A1541_ = new_A1522_ | new_A1523_;
  assign new_A1542_ = new_A1522_ | new_A1529_;
  assign new_A1543_ = new_A1521_ & new_A1533_;
  assign new_A1544_ = ~new_A1520_ | ~new_A1521_;
  assign new_A1545_ = new_A1529_ & new_A1544_;
  assign new_A1546_ = ~new_A1545_ & ~new_A1529_;
  assign new_A1547_ = new_A1529_ | new_A1544_;
  assign new_A1548_ = ~new_A1522_ | ~new_A1523_;
  assign new_A1549_ = new_A1529_ | new_A1544_;
  assign new_A1550_ = ~new_A1529_ & ~new_A1551_;
  assign new_A1551_ = new_A1529_ & new_A1544_;
  assign new_A1552_ = new_A2318_;
  assign new_A1553_ = new_A2351_;
  assign new_A1554_ = new_A2384_;
  assign new_A1555_ = new_A2417_;
  assign new_A1556_ = new_A2450_;
  assign new_A1557_ = new_A1563_ & new_A1562_;
  assign new_A1558_ = new_A1565_ | new_A1564_;
  assign new_A1559_ = new_A1567_ | new_A1566_;
  assign new_A1560_ = new_A1562_ & new_A1568_;
  assign new_A1561_ = new_A1562_ & new_A1569_;
  assign new_A1562_ = new_A1552_ ^ new_A1553_;
  assign new_A1563_ = new_A1564_ ^ new_A1554_;
  assign new_A1564_ = new_A1572_ & new_A1571_;
  assign new_A1565_ = new_A1570_ & new_A1554_;
  assign new_A1566_ = new_A1575_ & new_A1574_;
  assign new_A1567_ = new_A1573_ & new_A1554_;
  assign new_A1568_ = new_A1576_ | new_A1553_;
  assign new_A1569_ = ~new_A1554_ ^ new_A1566_;
  assign new_A1570_ = ~new_A1579_ | ~new_A1580_;
  assign new_A1571_ = new_A1555_ ^ new_A1562_;
  assign new_A1572_ = new_A1581_ & new_A1574_;
  assign new_A1573_ = ~new_A1583_ | ~new_A1582_;
  assign new_A1574_ = new_A1555_ | new_A1556_;
  assign new_A1575_ = new_A1555_ | new_A1562_;
  assign new_A1576_ = new_A1554_ & new_A1566_;
  assign new_A1577_ = ~new_A1553_ | ~new_A1554_;
  assign new_A1578_ = new_A1562_ & new_A1577_;
  assign new_A1579_ = ~new_A1578_ & ~new_A1562_;
  assign new_A1580_ = new_A1562_ | new_A1577_;
  assign new_A1581_ = ~new_A1555_ | ~new_A1556_;
  assign new_A1582_ = new_A1562_ | new_A1577_;
  assign new_A1583_ = ~new_A1562_ & ~new_A1584_;
  assign new_A1584_ = new_A1562_ & new_A1577_;
  assign new_A1585_ = new_A2483_;
  assign new_A1586_ = new_A2516_;
  assign new_A1587_ = new_A2549_;
  assign new_A1588_ = new_A2582_;
  assign new_A1589_ = new_A2615_;
  assign new_A1590_ = new_A1596_ & new_A1595_;
  assign new_A1591_ = new_A1598_ | new_A1597_;
  assign new_A1592_ = new_A1600_ | new_A1599_;
  assign new_A1593_ = new_A1595_ & new_A1601_;
  assign new_A1594_ = new_A1595_ & new_A1602_;
  assign new_A1595_ = new_A1585_ ^ new_A1586_;
  assign new_A1596_ = new_A1597_ ^ new_A1587_;
  assign new_A1597_ = new_A1605_ & new_A1604_;
  assign new_A1598_ = new_A1603_ & new_A1587_;
  assign new_A1599_ = new_A1608_ & new_A1607_;
  assign new_A1600_ = new_A1606_ & new_A1587_;
  assign new_A1601_ = new_A1609_ | new_A1586_;
  assign new_A1602_ = ~new_A1587_ ^ new_A1599_;
  assign new_A1603_ = ~new_A1612_ | ~new_A1613_;
  assign new_A1604_ = new_A1588_ ^ new_A1595_;
  assign new_A1605_ = new_A1614_ & new_A1607_;
  assign new_A1606_ = ~new_A1616_ | ~new_A1615_;
  assign new_A1607_ = new_A1588_ | new_A1589_;
  assign new_A1608_ = new_A1588_ | new_A1595_;
  assign new_A1609_ = new_A1587_ & new_A1599_;
  assign new_A1610_ = ~new_A1586_ | ~new_A1587_;
  assign new_A1611_ = new_A1595_ & new_A1610_;
  assign new_A1612_ = ~new_A1611_ & ~new_A1595_;
  assign new_A1613_ = new_A1595_ | new_A1610_;
  assign new_A1614_ = ~new_A1588_ | ~new_A1589_;
  assign new_A1615_ = new_A1595_ | new_A1610_;
  assign new_A1616_ = ~new_A1595_ & ~new_A1617_;
  assign new_A1617_ = new_A1595_ & new_A1610_;
  assign new_A1618_ = new_A2648_;
  assign new_A1619_ = new_A2681_;
  assign new_A1620_ = new_A2714_;
  assign new_A1621_ = new_A2747_;
  assign new_A1622_ = new_A2780_;
  assign new_A1623_ = new_A1629_ & new_A1628_;
  assign new_A1624_ = new_A1631_ | new_A1630_;
  assign new_A1625_ = new_A1633_ | new_A1632_;
  assign new_A1626_ = new_A1628_ & new_A1634_;
  assign new_A1627_ = new_A1628_ & new_A1635_;
  assign new_A1628_ = new_A1618_ ^ new_A1619_;
  assign new_A1629_ = new_A1630_ ^ new_A1620_;
  assign new_A1630_ = new_A1638_ & new_A1637_;
  assign new_A1631_ = new_A1636_ & new_A1620_;
  assign new_A1632_ = new_A1641_ & new_A1640_;
  assign new_A1633_ = new_A1639_ & new_A1620_;
  assign new_A1634_ = new_A1642_ | new_A1619_;
  assign new_A1635_ = ~new_A1620_ ^ new_A1632_;
  assign new_A1636_ = ~new_A1645_ | ~new_A1646_;
  assign new_A1637_ = new_A1621_ ^ new_A1628_;
  assign new_A1638_ = new_A1647_ & new_A1640_;
  assign new_A1639_ = ~new_A1649_ | ~new_A1648_;
  assign new_A1640_ = new_A1621_ | new_A1622_;
  assign new_A1641_ = new_A1621_ | new_A1628_;
  assign new_A1642_ = new_A1620_ & new_A1632_;
  assign new_A1643_ = ~new_A1619_ | ~new_A1620_;
  assign new_A1644_ = new_A1628_ & new_A1643_;
  assign new_A1645_ = ~new_A1644_ & ~new_A1628_;
  assign new_A1646_ = new_A1628_ | new_A1643_;
  assign new_A1647_ = ~new_A1621_ | ~new_A1622_;
  assign new_A1648_ = new_A1628_ | new_A1643_;
  assign new_A1649_ = ~new_A1628_ & ~new_A1650_;
  assign new_A1650_ = new_A1628_ & new_A1643_;
  assign new_A1651_ = new_A1987_;
  assign new_A1652_ = new_A2022_;
  assign new_A1653_ = new_A2055_;
  assign new_A1654_ = new_A2088_;
  assign new_A1655_ = new_A2121_;
  assign new_A1656_ = new_A1662_ & new_A1661_;
  assign new_A1657_ = new_A1664_ | new_A1663_;
  assign new_A1658_ = new_A1666_ | new_A1665_;
  assign new_A1659_ = new_A1661_ & new_A1667_;
  assign new_A1660_ = new_A1661_ & new_A1668_;
  assign new_A1661_ = new_A1651_ ^ new_A1652_;
  assign new_A1662_ = new_A1663_ ^ new_A1653_;
  assign new_A1663_ = new_A1671_ & new_A1670_;
  assign new_A1664_ = new_A1669_ & new_A1653_;
  assign new_A1665_ = new_A1674_ & new_A1673_;
  assign new_A1666_ = new_A1672_ & new_A1653_;
  assign new_A1667_ = new_A1675_ | new_A1652_;
  assign new_A1668_ = ~new_A1653_ ^ new_A1665_;
  assign new_A1669_ = ~new_A1678_ | ~new_A1679_;
  assign new_A1670_ = new_A1654_ ^ new_A1661_;
  assign new_A1671_ = new_A1680_ & new_A1673_;
  assign new_A1672_ = ~new_A1682_ | ~new_A1681_;
  assign new_A1673_ = new_A1654_ | new_A1655_;
  assign new_A1674_ = new_A1654_ | new_A1661_;
  assign new_A1675_ = new_A1653_ & new_A1665_;
  assign new_A1676_ = ~new_A1652_ | ~new_A1653_;
  assign new_A1677_ = new_A1661_ & new_A1676_;
  assign new_A1678_ = ~new_A1677_ & ~new_A1661_;
  assign new_A1679_ = new_A1661_ | new_A1676_;
  assign new_A1680_ = ~new_A1654_ | ~new_A1655_;
  assign new_A1681_ = new_A1661_ | new_A1676_;
  assign new_A1682_ = ~new_A1661_ & ~new_A1683_;
  assign new_A1683_ = new_A1661_ & new_A1676_;
  assign new_A1684_ = new_A2154_;
  assign new_A1685_ = new_A2187_;
  assign new_A1686_ = new_A2220_;
  assign new_A1687_ = new_A2253_;
  assign new_A1688_ = new_A2286_;
  assign new_A1689_ = new_A1695_ & new_A1694_;
  assign new_A1690_ = new_A1697_ | new_A1696_;
  assign new_A1691_ = new_A1699_ | new_A1698_;
  assign new_A1692_ = new_A1694_ & new_A1700_;
  assign new_A1693_ = new_A1694_ & new_A1701_;
  assign new_A1694_ = new_A1684_ ^ new_A1685_;
  assign new_A1695_ = new_A1696_ ^ new_A1686_;
  assign new_A1696_ = new_A1704_ & new_A1703_;
  assign new_A1697_ = new_A1702_ & new_A1686_;
  assign new_A1698_ = new_A1707_ & new_A1706_;
  assign new_A1699_ = new_A1705_ & new_A1686_;
  assign new_A1700_ = new_A1708_ | new_A1685_;
  assign new_A1701_ = ~new_A1686_ ^ new_A1698_;
  assign new_A1702_ = ~new_A1711_ | ~new_A1712_;
  assign new_A1703_ = new_A1687_ ^ new_A1694_;
  assign new_A1704_ = new_A1713_ & new_A1706_;
  assign new_A1705_ = ~new_A1715_ | ~new_A1714_;
  assign new_A1706_ = new_A1687_ | new_A1688_;
  assign new_A1707_ = new_A1687_ | new_A1694_;
  assign new_A1708_ = new_A1686_ & new_A1698_;
  assign new_A1709_ = ~new_A1685_ | ~new_A1686_;
  assign new_A1710_ = new_A1694_ & new_A1709_;
  assign new_A1711_ = ~new_A1710_ & ~new_A1694_;
  assign new_A1712_ = new_A1694_ | new_A1709_;
  assign new_A1713_ = ~new_A1687_ | ~new_A1688_;
  assign new_A1714_ = new_A1694_ | new_A1709_;
  assign new_A1715_ = ~new_A1694_ & ~new_A1716_;
  assign new_A1716_ = new_A1694_ & new_A1709_;
  assign new_A1717_ = new_A2319_;
  assign new_A1718_ = new_A2352_;
  assign new_A1719_ = new_A2385_;
  assign new_A1720_ = new_A2418_;
  assign new_A1721_ = new_A2451_;
  assign new_A1722_ = new_A1728_ & new_A1727_;
  assign new_A1723_ = new_A1730_ | new_A1729_;
  assign new_A1724_ = new_A1732_ | new_A1731_;
  assign new_A1725_ = new_A1727_ & new_A1733_;
  assign new_A1726_ = new_A1727_ & new_A1734_;
  assign new_A1727_ = new_A1717_ ^ new_A1718_;
  assign new_A1728_ = new_A1729_ ^ new_A1719_;
  assign new_A1729_ = new_A1737_ & new_A1736_;
  assign new_A1730_ = new_A1735_ & new_A1719_;
  assign new_A1731_ = new_A1740_ & new_A1739_;
  assign new_A1732_ = new_A1738_ & new_A1719_;
  assign new_A1733_ = new_A1741_ | new_A1718_;
  assign new_A1734_ = ~new_A1719_ ^ new_A1731_;
  assign new_A1735_ = ~new_A1744_ | ~new_A1745_;
  assign new_A1736_ = new_A1720_ ^ new_A1727_;
  assign new_A1737_ = new_A1746_ & new_A1739_;
  assign new_A1738_ = ~new_A1748_ | ~new_A1747_;
  assign new_A1739_ = new_A1720_ | new_A1721_;
  assign new_A1740_ = new_A1720_ | new_A1727_;
  assign new_A1741_ = new_A1719_ & new_A1731_;
  assign new_A1742_ = ~new_A1718_ | ~new_A1719_;
  assign new_A1743_ = new_A1727_ & new_A1742_;
  assign new_A1744_ = ~new_A1743_ & ~new_A1727_;
  assign new_A1745_ = new_A1727_ | new_A1742_;
  assign new_A1746_ = ~new_A1720_ | ~new_A1721_;
  assign new_A1747_ = new_A1727_ | new_A1742_;
  assign new_A1748_ = ~new_A1727_ & ~new_A1749_;
  assign new_A1749_ = new_A1727_ & new_A1742_;
  assign new_A1750_ = new_A2484_;
  assign new_A1751_ = new_A2517_;
  assign new_A1752_ = new_A2550_;
  assign new_A1753_ = new_A2583_;
  assign new_A1754_ = new_A2616_;
  assign new_A1755_ = new_A1761_ & new_A1760_;
  assign new_A1756_ = new_A1763_ | new_A1762_;
  assign new_A1757_ = new_A1765_ | new_A1764_;
  assign new_A1758_ = new_A1760_ & new_A1766_;
  assign new_A1759_ = new_A1760_ & new_A1767_;
  assign new_A1760_ = new_A1750_ ^ new_A1751_;
  assign new_A1761_ = new_A1762_ ^ new_A1752_;
  assign new_A1762_ = new_A1770_ & new_A1769_;
  assign new_A1763_ = new_A1768_ & new_A1752_;
  assign new_A1764_ = new_A1773_ & new_A1772_;
  assign new_A1765_ = new_A1771_ & new_A1752_;
  assign new_A1766_ = new_A1774_ | new_A1751_;
  assign new_A1767_ = ~new_A1752_ ^ new_A1764_;
  assign new_A1768_ = ~new_A1777_ | ~new_A1778_;
  assign new_A1769_ = new_A1753_ ^ new_A1760_;
  assign new_A1770_ = new_A1779_ & new_A1772_;
  assign new_A1771_ = ~new_A1781_ | ~new_A1780_;
  assign new_A1772_ = new_A1753_ | new_A1754_;
  assign new_A1773_ = new_A1753_ | new_A1760_;
  assign new_A1774_ = new_A1752_ & new_A1764_;
  assign new_A1775_ = ~new_A1751_ | ~new_A1752_;
  assign new_A1776_ = new_A1760_ & new_A1775_;
  assign new_A1777_ = ~new_A1776_ & ~new_A1760_;
  assign new_A1778_ = new_A1760_ | new_A1775_;
  assign new_A1779_ = ~new_A1753_ | ~new_A1754_;
  assign new_A1780_ = new_A1760_ | new_A1775_;
  assign new_A1781_ = ~new_A1760_ & ~new_A1782_;
  assign new_A1782_ = new_A1760_ & new_A1775_;
  assign new_A1783_ = new_A2649_;
  assign new_A1784_ = new_A2682_;
  assign new_A1785_ = new_A2715_;
  assign new_A1786_ = new_A2748_;
  assign new_A1787_ = new_A2781_;
  assign new_A1788_ = new_A1794_ & new_A1793_;
  assign new_A1789_ = new_A1796_ | new_A1795_;
  assign new_A1790_ = new_A1798_ | new_A1797_;
  assign new_A1791_ = new_A1793_ & new_A1799_;
  assign new_A1792_ = new_A1793_ & new_A1800_;
  assign new_A1793_ = new_A1783_ ^ new_A1784_;
  assign new_A1794_ = new_A1795_ ^ new_A1785_;
  assign new_A1795_ = new_A1803_ & new_A1802_;
  assign new_A1796_ = new_A1801_ & new_A1785_;
  assign new_A1797_ = new_A1806_ & new_A1805_;
  assign new_A1798_ = new_A1804_ & new_A1785_;
  assign new_A1799_ = new_A1807_ | new_A1784_;
  assign new_A1800_ = ~new_A1785_ ^ new_A1797_;
  assign new_A1801_ = ~new_A1810_ | ~new_A1811_;
  assign new_A1802_ = new_A1786_ ^ new_A1793_;
  assign new_A1803_ = new_A1812_ & new_A1805_;
  assign new_A1804_ = ~new_A1814_ | ~new_A1813_;
  assign new_A1805_ = new_A1786_ | new_A1787_;
  assign new_A1806_ = new_A1786_ | new_A1793_;
  assign new_A1807_ = new_A1785_ & new_A1797_;
  assign new_A1808_ = ~new_A1784_ | ~new_A1785_;
  assign new_A1809_ = new_A1793_ & new_A1808_;
  assign new_A1810_ = ~new_A1809_ & ~new_A1793_;
  assign new_A1811_ = new_A1793_ | new_A1808_;
  assign new_A1812_ = ~new_A1786_ | ~new_A1787_;
  assign new_A1813_ = new_A1793_ | new_A1808_;
  assign new_A1814_ = ~new_A1793_ & ~new_A1815_;
  assign new_A1815_ = new_A1793_ & new_A1808_;
  assign new_A1816_ = new_A1986_;
  assign new_A1817_ = new_A2023_;
  assign new_A1818_ = new_A2056_;
  assign new_A1819_ = new_A2089_;
  assign new_A1820_ = new_A2122_;
  assign new_A1821_ = new_A1827_ & new_A1826_;
  assign new_A1822_ = new_A1829_ | new_A1828_;
  assign new_A1823_ = new_A1831_ | new_A1830_;
  assign new_A1824_ = new_A1826_ & new_A1832_;
  assign new_A1825_ = new_A1826_ & new_A1833_;
  assign new_A1826_ = new_A1816_ ^ new_A1817_;
  assign new_A1827_ = new_A1828_ ^ new_A1818_;
  assign new_A1828_ = new_A1836_ & new_A1835_;
  assign new_A1829_ = new_A1834_ & new_A1818_;
  assign new_A1830_ = new_A1839_ & new_A1838_;
  assign new_A1831_ = new_A1837_ & new_A1818_;
  assign new_A1832_ = new_A1840_ | new_A1817_;
  assign new_A1833_ = ~new_A1818_ ^ new_A1830_;
  assign new_A1834_ = ~new_A1843_ | ~new_A1844_;
  assign new_A1835_ = new_A1819_ ^ new_A1826_;
  assign new_A1836_ = new_A1845_ & new_A1838_;
  assign new_A1837_ = ~new_A1847_ | ~new_A1846_;
  assign new_A1838_ = new_A1819_ | new_A1820_;
  assign new_A1839_ = new_A1819_ | new_A1826_;
  assign new_A1840_ = new_A1818_ & new_A1830_;
  assign new_A1841_ = ~new_A1817_ | ~new_A1818_;
  assign new_A1842_ = new_A1826_ & new_A1841_;
  assign new_A1843_ = ~new_A1842_ & ~new_A1826_;
  assign new_A1844_ = new_A1826_ | new_A1841_;
  assign new_A1845_ = ~new_A1819_ | ~new_A1820_;
  assign new_A1846_ = new_A1826_ | new_A1841_;
  assign new_A1847_ = ~new_A1826_ & ~new_A1848_;
  assign new_A1848_ = new_A1826_ & new_A1841_;
  assign new_A1849_ = new_A2155_;
  assign new_A1850_ = new_A2188_;
  assign new_A1851_ = new_A2221_;
  assign new_A1852_ = new_A2254_;
  assign new_A1853_ = new_A2287_;
  assign new_A1854_ = new_A1860_ & new_A1859_;
  assign new_A1855_ = new_A1862_ | new_A1861_;
  assign new_A1856_ = new_A1864_ | new_A1863_;
  assign new_A1857_ = new_A1859_ & new_A1865_;
  assign new_A1858_ = new_A1859_ & new_A1866_;
  assign new_A1859_ = new_A1849_ ^ new_A1850_;
  assign new_A1860_ = new_A1861_ ^ new_A1851_;
  assign new_A1861_ = new_A1869_ & new_A1868_;
  assign new_A1862_ = new_A1867_ & new_A1851_;
  assign new_A1863_ = new_A1872_ & new_A1871_;
  assign new_A1864_ = new_A1870_ & new_A1851_;
  assign new_A1865_ = new_A1873_ | new_A1850_;
  assign new_A1866_ = ~new_A1851_ ^ new_A1863_;
  assign new_A1867_ = ~new_A1876_ | ~new_A1877_;
  assign new_A1868_ = new_A1852_ ^ new_A1859_;
  assign new_A1869_ = new_A1878_ & new_A1871_;
  assign new_A1870_ = ~new_A1880_ | ~new_A1879_;
  assign new_A1871_ = new_A1852_ | new_A1853_;
  assign new_A1872_ = new_A1852_ | new_A1859_;
  assign new_A1873_ = new_A1851_ & new_A1863_;
  assign new_A1874_ = ~new_A1850_ | ~new_A1851_;
  assign new_A1875_ = new_A1859_ & new_A1874_;
  assign new_A1876_ = ~new_A1875_ & ~new_A1859_;
  assign new_A1877_ = new_A1859_ | new_A1874_;
  assign new_A1878_ = ~new_A1852_ | ~new_A1853_;
  assign new_A1879_ = new_A1859_ | new_A1874_;
  assign new_A1880_ = ~new_A1859_ & ~new_A1881_;
  assign new_A1881_ = new_A1859_ & new_A1874_;
  assign new_A1882_ = new_A2320_;
  assign new_A1883_ = new_A2353_;
  assign new_A1884_ = new_A2386_;
  assign new_A1885_ = new_A2419_;
  assign new_A1886_ = new_A2452_;
  assign new_A1887_ = new_A1893_ & new_A1892_;
  assign new_A1888_ = new_A1895_ | new_A1894_;
  assign new_A1889_ = new_A1897_ | new_A1896_;
  assign new_A1890_ = new_A1892_ & new_A1898_;
  assign new_A1891_ = new_A1892_ & new_A1899_;
  assign new_A1892_ = new_A1882_ ^ new_A1883_;
  assign new_A1893_ = new_A1894_ ^ new_A1884_;
  assign new_A1894_ = new_A1902_ & new_A1901_;
  assign new_A1895_ = new_A1900_ & new_A1884_;
  assign new_A1896_ = new_A1905_ & new_A1904_;
  assign new_A1897_ = new_A1903_ & new_A1884_;
  assign new_A1898_ = new_A1906_ | new_A1883_;
  assign new_A1899_ = ~new_A1884_ ^ new_A1896_;
  assign new_A1900_ = ~new_A1909_ | ~new_A1910_;
  assign new_A1901_ = new_A1885_ ^ new_A1892_;
  assign new_A1902_ = new_A1911_ & new_A1904_;
  assign new_A1903_ = ~new_A1913_ | ~new_A1912_;
  assign new_A1904_ = new_A1885_ | new_A1886_;
  assign new_A1905_ = new_A1885_ | new_A1892_;
  assign new_A1906_ = new_A1884_ & new_A1896_;
  assign new_A1907_ = ~new_A1883_ | ~new_A1884_;
  assign new_A1908_ = new_A1892_ & new_A1907_;
  assign new_A1909_ = ~new_A1908_ & ~new_A1892_;
  assign new_A1910_ = new_A1892_ | new_A1907_;
  assign new_A1911_ = ~new_A1885_ | ~new_A1886_;
  assign new_A1912_ = new_A1892_ | new_A1907_;
  assign new_A1913_ = ~new_A1892_ & ~new_A1914_;
  assign new_A1914_ = new_A1892_ & new_A1907_;
  assign new_A1915_ = new_A2485_;
  assign new_A1916_ = new_A2518_;
  assign new_A1917_ = new_A2551_;
  assign new_A1918_ = new_A2584_;
  assign new_A1919_ = new_A2617_;
  assign new_A1920_ = new_A1926_ & new_A1925_;
  assign new_A1921_ = new_A1928_ | new_A1927_;
  assign new_A1922_ = new_A1930_ | new_A1929_;
  assign new_A1923_ = new_A1925_ & new_A1931_;
  assign new_A1924_ = new_A1925_ & new_A1932_;
  assign new_A1925_ = new_A1915_ ^ new_A1916_;
  assign new_A1926_ = new_A1927_ ^ new_A1917_;
  assign new_A1927_ = new_A1935_ & new_A1934_;
  assign new_A1928_ = new_A1933_ & new_A1917_;
  assign new_A1929_ = new_A1938_ & new_A1937_;
  assign new_A1930_ = new_A1936_ & new_A1917_;
  assign new_A1931_ = new_A1939_ | new_A1916_;
  assign new_A1932_ = ~new_A1917_ ^ new_A1929_;
  assign new_A1933_ = ~new_A1942_ | ~new_A1943_;
  assign new_A1934_ = new_A1918_ ^ new_A1925_;
  assign new_A1935_ = new_A1944_ & new_A1937_;
  assign new_A1936_ = ~new_A1946_ | ~new_A1945_;
  assign new_A1937_ = new_A1918_ | new_A1919_;
  assign new_A1938_ = new_A1918_ | new_A1925_;
  assign new_A1939_ = new_A1917_ & new_A1929_;
  assign new_A1940_ = ~new_A1916_ | ~new_A1917_;
  assign new_A1941_ = new_A1925_ & new_A1940_;
  assign new_A1942_ = ~new_A1941_ & ~new_A1925_;
  assign new_A1943_ = new_A1925_ | new_A1940_;
  assign new_A1944_ = ~new_A1918_ | ~new_A1919_;
  assign new_A1945_ = new_A1925_ | new_A1940_;
  assign new_A1946_ = ~new_A1925_ & ~new_A1947_;
  assign new_A1947_ = new_A1925_ & new_A1940_;
  assign new_A1948_ = new_A2650_;
  assign new_A1949_ = new_A2683_;
  assign new_A1950_ = new_A2716_;
  assign new_A1951_ = new_A2749_;
  assign new_A1952_ = new_A2782_;
  assign new_A1953_ = new_A1959_ & new_A1958_;
  assign new_A1954_ = new_A1961_ | new_A1960_;
  assign new_A1955_ = new_A1963_ | new_A1962_;
  assign new_A1956_ = new_A1958_ & new_A1964_;
  assign new_A1957_ = new_A1958_ & new_A1965_;
  assign new_A1958_ = new_A1948_ ^ new_A1949_;
  assign new_A1959_ = new_A1960_ ^ new_A1950_;
  assign new_A1960_ = new_A1968_ & new_A1967_;
  assign new_A1961_ = new_A1966_ & new_A1950_;
  assign new_A1962_ = new_A1971_ & new_A1970_;
  assign new_A1963_ = new_A1969_ & new_A1950_;
  assign new_A1964_ = new_A1972_ | new_A1949_;
  assign new_A1965_ = ~new_A1950_ ^ new_A1962_;
  assign new_A1966_ = ~new_A1975_ | ~new_A1976_;
  assign new_A1967_ = new_A1951_ ^ new_A1958_;
  assign new_A1968_ = new_A1977_ & new_A1970_;
  assign new_A1969_ = ~new_A1979_ | ~new_A1978_;
  assign new_A1970_ = new_A1951_ | new_A1952_;
  assign new_A1971_ = new_A1951_ | new_A1958_;
  assign new_A1972_ = new_A1950_ & new_A1962_;
  assign new_A1973_ = ~new_A1949_ | ~new_A1950_;
  assign new_A1974_ = new_A1958_ & new_A1973_;
  assign new_A1975_ = ~new_A1974_ & ~new_A1958_;
  assign new_A1976_ = new_A1958_ | new_A1973_;
  assign new_A1977_ = ~new_A1951_ | ~new_A1952_;
  assign new_A1978_ = new_A1958_ | new_A1973_;
  assign new_A1979_ = ~new_A1958_ & ~new_A1980_;
  assign new_A1980_ = new_A1958_ & new_A1973_;
  assign new_A1155_ = new_A1133_ & new_A1148_;
  assign new_A1154_ = ~new_A1133_ & ~new_A1155_;
  assign new_A1153_ = new_A1133_ | new_A1148_;
  assign new_A1152_ = ~new_A1126_ | ~new_A1127_;
  assign new_A1151_ = new_A1133_ | new_A1148_;
  assign new_A1150_ = ~new_A1149_ & ~new_A1133_;
  assign new_A1149_ = new_A1133_ & new_A1148_;
  assign new_A1148_ = ~new_A1124_ | ~new_A1125_;
  assign new_A1147_ = new_A1125_ & new_A1137_;
  assign new_A1146_ = new_A1126_ | new_A1133_;
  assign new_A1145_ = new_A1126_ | new_A1127_;
  assign new_A1144_ = ~new_A1154_ | ~new_A1153_;
  assign new_A1143_ = new_A1152_ & new_A1145_;
  assign new_A1142_ = new_A1126_ ^ new_A1133_;
  assign new_A1141_ = ~new_A1150_ | ~new_A1151_;
  assign new_A1140_ = ~new_A1125_ ^ new_A1137_;
  assign new_A1139_ = new_A1147_ | new_A1124_;
  assign new_A1138_ = new_A1144_ & new_A1125_;
  assign new_A1137_ = new_A1146_ & new_A1145_;
  assign new_A1136_ = new_A1141_ & new_A1125_;
  assign new_A1135_ = new_A1143_ & new_A1142_;
  assign new_A1134_ = new_A1135_ ^ new_A1125_;
  assign new_A1133_ = new_A1123_ ^ new_A1124_;
  assign A1132 = new_A1133_ & new_A1140_;
  assign A1131 = new_A1133_ & new_A1139_;
  assign A1130 = new_A1138_ | new_A1137_;
  assign A1129 = new_A1136_ | new_A1135_;
  assign A1128 = new_A1134_ & new_A1133_;
  assign new_A1127_ = new_A1957_;
  assign new_A1126_ = new_A1924_;
  assign new_A1125_ = new_A1891_;
  assign new_A1124_ = new_A1858_;
  assign new_A1123_ = new_A1825_;
  assign new_A1122_ = new_A1100_ & new_A1115_;
  assign new_A1121_ = ~new_A1100_ & ~new_A1122_;
  assign new_A1120_ = new_A1100_ | new_A1115_;
  assign new_A1119_ = ~new_A1093_ | ~new_A1094_;
  assign new_A1118_ = new_A1100_ | new_A1115_;
  assign new_A1117_ = ~new_A1116_ & ~new_A1100_;
  assign new_A1116_ = new_A1100_ & new_A1115_;
  assign new_A1115_ = ~new_A1091_ | ~new_A1092_;
  assign new_A1114_ = new_A1092_ & new_A1104_;
  assign new_A1113_ = new_A1093_ | new_A1100_;
  assign new_A1112_ = new_A1093_ | new_A1094_;
  assign new_A1111_ = ~new_A1121_ | ~new_A1120_;
  assign new_A1110_ = new_A1119_ & new_A1112_;
  assign new_A1109_ = new_A1093_ ^ new_A1100_;
  assign new_A1108_ = ~new_A1117_ | ~new_A1118_;
  assign new_A1107_ = ~new_A1092_ ^ new_A1104_;
  assign new_A1106_ = new_A1114_ | new_A1091_;
  assign new_A1105_ = new_A1111_ & new_A1092_;
  assign new_A1104_ = new_A1113_ & new_A1112_;
  assign new_A1103_ = new_A1108_ & new_A1092_;
  assign new_A1102_ = new_A1110_ & new_A1109_;
  assign new_A1101_ = new_A1102_ ^ new_A1092_;
  assign new_A1100_ = new_A1090_ ^ new_A1091_;
  assign A1099 = new_A1100_ & new_A1107_;
  assign A1098 = new_A1100_ & new_A1106_;
  assign A1097 = new_A1105_ | new_A1104_;
  assign A1096 = new_A1103_ | new_A1102_;
  assign A1095 = new_A1101_ & new_A1100_;
  assign new_A1094_ = new_A1792_;
  assign new_A1093_ = new_A1759_;
  assign new_A1092_ = new_A1726_;
  assign new_A1091_ = new_A1693_;
  assign new_A1090_ = new_A1660_;
  assign new_A1089_ = new_A1067_ & new_A1082_;
  assign new_A1088_ = ~new_A1067_ & ~new_A1089_;
  assign new_A1087_ = new_A1067_ | new_A1082_;
  assign new_A1086_ = ~new_A1060_ | ~new_A1061_;
  assign new_A1085_ = new_A1067_ | new_A1082_;
  assign new_A1084_ = ~new_A1083_ & ~new_A1067_;
  assign new_A1083_ = new_A1067_ & new_A1082_;
  assign new_A1082_ = ~new_A1058_ | ~new_A1059_;
  assign new_A1081_ = new_A1059_ & new_A1071_;
  assign new_A1080_ = new_A1060_ | new_A1067_;
  assign new_A1079_ = new_A1060_ | new_A1061_;
  assign new_A1078_ = ~new_A1088_ | ~new_A1087_;
  assign new_A1077_ = new_A1086_ & new_A1079_;
  assign new_A1076_ = new_A1060_ ^ new_A1067_;
  assign new_A1075_ = ~new_A1084_ | ~new_A1085_;
  assign new_A1074_ = ~new_A1059_ ^ new_A1071_;
  assign new_A1073_ = new_A1081_ | new_A1058_;
  assign new_A1072_ = new_A1078_ & new_A1059_;
  assign new_A1071_ = new_A1080_ & new_A1079_;
  assign new_A1070_ = new_A1075_ & new_A1059_;
  assign new_A1069_ = new_A1077_ & new_A1076_;
  assign new_A1068_ = new_A1069_ ^ new_A1059_;
  assign new_A1067_ = new_A1057_ ^ new_A1058_;
  assign A1066 = new_A1067_ & new_A1074_;
  assign A1065 = new_A1067_ & new_A1073_;
  assign A1064 = new_A1072_ | new_A1071_;
  assign A1063 = new_A1070_ | new_A1069_;
  assign A1062 = new_A1068_ & new_A1067_;
  assign new_A1061_ = new_A1627_;
  assign new_A1060_ = new_A1594_;
  assign new_A1059_ = new_A1561_;
  assign new_A1058_ = new_A1528_;
  assign new_A1057_ = new_A1495_;
  assign new_A1056_ = new_A1034_ & new_A1049_;
  assign new_A1055_ = ~new_A1034_ & ~new_A1056_;
  assign new_A1054_ = new_A1034_ | new_A1049_;
  assign new_A1053_ = ~new_A1027_ | ~new_A1028_;
  assign new_A1052_ = new_A1034_ | new_A1049_;
  assign new_A1051_ = ~new_A1050_ & ~new_A1034_;
  assign new_A1050_ = new_A1034_ & new_A1049_;
  assign new_A1049_ = ~new_A1025_ | ~new_A1026_;
  assign new_A1048_ = new_A1026_ & new_A1038_;
  assign new_A1047_ = new_A1027_ | new_A1034_;
  assign new_A1046_ = new_A1027_ | new_A1028_;
  assign new_A1045_ = ~new_A1055_ | ~new_A1054_;
  assign new_A1044_ = new_A1053_ & new_A1046_;
  assign new_A1043_ = new_A1027_ ^ new_A1034_;
  assign new_A1042_ = ~new_A1051_ | ~new_A1052_;
  assign new_A1041_ = ~new_A1026_ ^ new_A1038_;
  assign new_A1040_ = new_A1048_ | new_A1025_;
  assign new_A1039_ = new_A1045_ & new_A1026_;
  assign new_A1038_ = new_A1047_ & new_A1046_;
  assign new_A1037_ = new_A1042_ & new_A1026_;
  assign new_A1036_ = new_A1044_ & new_A1043_;
  assign new_A1035_ = new_A1036_ ^ new_A1026_;
  assign new_A1034_ = new_A1024_ ^ new_A1025_;
  assign A1033 = new_A1034_ & new_A1041_;
  assign A1032 = new_A1034_ & new_A1040_;
  assign A1031 = new_A1039_ | new_A1038_;
  assign A1030 = new_A1037_ | new_A1036_;
  assign A1029 = new_A1035_ & new_A1034_;
  assign new_A1028_ = new_A1462_;
  assign new_A1027_ = new_A1429_;
  assign new_A1026_ = new_A1396_;
  assign new_A1025_ = new_A1363_;
  assign new_A1024_ = new_A1330_;
  assign new_A1023_ = new_A1001_ & new_A1016_;
  assign new_A1022_ = ~new_A1001_ & ~new_A1023_;
  assign new_A1021_ = new_A1001_ | new_A1016_;
  assign new_A1020_ = ~new_A994_ | ~new_A995_;
  assign new_A1019_ = new_A1001_ | new_A1016_;
  assign new_A1018_ = ~new_A1017_ & ~new_A1001_;
  assign new_A1017_ = new_A1001_ & new_A1016_;
  assign new_A1016_ = ~new_A992_ | ~new_A993_;
  assign new_A1015_ = new_A993_ & new_A1005_;
  assign new_A1014_ = new_A994_ | new_A1001_;
  assign new_A1013_ = new_A994_ | new_A995_;
  assign new_A1012_ = ~new_A1022_ | ~new_A1021_;
  assign new_A1011_ = new_A1020_ & new_A1013_;
  assign new_A1010_ = new_A994_ ^ new_A1001_;
  assign new_A1009_ = ~new_A1018_ | ~new_A1019_;
  assign new_A1008_ = ~new_A993_ ^ new_A1005_;
  assign new_A1007_ = new_A1015_ | new_A992_;
  assign new_A1006_ = new_A1012_ & new_A993_;
  assign new_A1005_ = new_A1014_ & new_A1013_;
  assign new_A1004_ = new_A1009_ & new_A993_;
  assign new_A1003_ = new_A1011_ & new_A1010_;
  assign new_A1002_ = new_A1003_ ^ new_A993_;
  assign new_A1001_ = new_A991_ ^ new_A992_;
  assign A1000 = new_A1001_ & new_A1008_;
  assign A999 = new_A1001_ & new_A1007_;
  assign A998 = new_A1006_ | new_A1005_;
  assign A997 = new_A1004_ | new_A1003_;
  assign A996 = new_A1002_ & new_A1001_;
  assign new_A995_ = new_A1297_;
  assign new_A994_ = new_A1264_;
  assign new_A993_ = new_A1231_;
  assign new_A992_ = new_A1198_;
  assign new_A991_ = new_A1161_;
  assign new_A990_ = new_A968_ & new_A983_;
  assign new_A989_ = ~new_A968_ & ~new_A990_;
  assign new_A988_ = new_A968_ | new_A983_;
  assign new_A987_ = ~new_A961_ | ~new_A962_;
  assign new_A986_ = new_A968_ | new_A983_;
  assign new_A985_ = ~new_A984_ & ~new_A968_;
  assign new_A984_ = new_A968_ & new_A983_;
  assign new_A983_ = ~new_A959_ | ~new_A960_;
  assign new_A982_ = new_A960_ & new_A972_;
  assign new_A981_ = new_A961_ | new_A968_;
  assign new_A980_ = new_A961_ | new_A962_;
  assign new_A979_ = ~new_A989_ | ~new_A988_;
  assign new_A978_ = new_A987_ & new_A980_;
  assign new_A977_ = new_A961_ ^ new_A968_;
  assign new_A976_ = ~new_A985_ | ~new_A986_;
  assign new_A975_ = ~new_A960_ ^ new_A972_;
  assign new_A974_ = new_A982_ | new_A959_;
  assign new_A973_ = new_A979_ & new_A960_;
  assign new_A972_ = new_A981_ & new_A980_;
  assign new_A971_ = new_A976_ & new_A960_;
  assign new_A970_ = new_A978_ & new_A977_;
  assign new_A969_ = new_A970_ ^ new_A960_;
  assign new_A968_ = new_A958_ ^ new_A959_;
  assign A967 = new_A968_ & new_A975_;
  assign A966 = new_A968_ & new_A974_;
  assign A965 = new_A973_ | new_A972_;
  assign A964 = new_A971_ | new_A970_;
  assign A963 = new_A969_ & new_A968_;
  assign new_A962_ = new_A1956_;
  assign new_A961_ = new_A1923_;
  assign new_A960_ = new_A1890_;
  assign new_A959_ = new_A1857_;
  assign new_A958_ = new_A1824_;
  assign new_A957_ = new_A935_ & new_A950_;
  assign new_A956_ = ~new_A935_ & ~new_A957_;
  assign new_A955_ = new_A935_ | new_A950_;
  assign new_A954_ = ~new_A928_ | ~new_A929_;
  assign new_A953_ = new_A935_ | new_A950_;
  assign new_A952_ = ~new_A951_ & ~new_A935_;
  assign new_A951_ = new_A935_ & new_A950_;
  assign new_A950_ = ~new_A926_ | ~new_A927_;
  assign new_A949_ = new_A927_ & new_A939_;
  assign new_A948_ = new_A928_ | new_A935_;
  assign new_A947_ = new_A928_ | new_A929_;
  assign new_A946_ = ~new_A956_ | ~new_A955_;
  assign new_A945_ = new_A954_ & new_A947_;
  assign new_A944_ = new_A928_ ^ new_A935_;
  assign new_A943_ = ~new_A952_ | ~new_A953_;
  assign new_A942_ = ~new_A927_ ^ new_A939_;
  assign new_A941_ = new_A949_ | new_A926_;
  assign new_A940_ = new_A946_ & new_A927_;
  assign new_A939_ = new_A948_ & new_A947_;
  assign new_A938_ = new_A943_ & new_A927_;
  assign new_A937_ = new_A945_ & new_A944_;
  assign new_A936_ = new_A937_ ^ new_A927_;
  assign new_A935_ = new_A925_ ^ new_A926_;
  assign A934 = new_A935_ & new_A942_;
  assign A933 = new_A935_ & new_A941_;
  assign A932 = new_A940_ | new_A939_;
  assign A931 = new_A938_ | new_A937_;
  assign A930 = new_A936_ & new_A935_;
  assign new_A929_ = new_A1791_;
  assign new_A928_ = new_A1758_;
  assign new_A927_ = new_A1725_;
  assign new_A926_ = new_A1692_;
  assign new_A925_ = new_A1659_;
  assign new_A924_ = new_A902_ & new_A917_;
  assign new_A923_ = ~new_A902_ & ~new_A924_;
  assign new_A922_ = new_A902_ | new_A917_;
  assign new_A921_ = ~new_A895_ | ~new_A896_;
  assign new_A920_ = new_A902_ | new_A917_;
  assign new_A919_ = ~new_A918_ & ~new_A902_;
  assign new_A918_ = new_A902_ & new_A917_;
  assign new_A917_ = ~new_A893_ | ~new_A894_;
  assign new_A916_ = new_A894_ & new_A906_;
  assign new_A915_ = new_A895_ | new_A902_;
  assign new_A914_ = new_A895_ | new_A896_;
  assign new_A913_ = ~new_A923_ | ~new_A922_;
  assign new_A912_ = new_A921_ & new_A914_;
  assign new_A911_ = new_A895_ ^ new_A902_;
  assign new_A910_ = ~new_A919_ | ~new_A920_;
  assign new_A909_ = ~new_A894_ ^ new_A906_;
  assign new_A908_ = new_A916_ | new_A893_;
  assign new_A907_ = new_A913_ & new_A894_;
  assign new_A906_ = new_A915_ & new_A914_;
  assign new_A905_ = new_A910_ & new_A894_;
  assign new_A904_ = new_A912_ & new_A911_;
  assign new_A903_ = new_A904_ ^ new_A894_;
  assign new_A902_ = new_A892_ ^ new_A893_;
  assign A901 = new_A902_ & new_A909_;
  assign A900 = new_A902_ & new_A908_;
  assign A899 = new_A907_ | new_A906_;
  assign A898 = new_A905_ | new_A904_;
  assign A897 = new_A903_ & new_A902_;
  assign new_A896_ = new_A1626_;
  assign new_A895_ = new_A1593_;
  assign new_A894_ = new_A1560_;
  assign new_A893_ = new_A1527_;
  assign new_A892_ = new_A1494_;
  assign new_A891_ = new_A869_ & new_A884_;
  assign new_A890_ = ~new_A869_ & ~new_A891_;
  assign new_A889_ = new_A869_ | new_A884_;
  assign new_A888_ = ~new_A862_ | ~new_A863_;
  assign new_A887_ = new_A869_ | new_A884_;
  assign new_A886_ = ~new_A885_ & ~new_A869_;
  assign new_A885_ = new_A869_ & new_A884_;
  assign new_A884_ = ~new_A860_ | ~new_A861_;
  assign new_A883_ = new_A861_ & new_A873_;
  assign new_A882_ = new_A862_ | new_A869_;
  assign new_A881_ = new_A862_ | new_A863_;
  assign new_A880_ = ~new_A890_ | ~new_A889_;
  assign new_A879_ = new_A888_ & new_A881_;
  assign new_A878_ = new_A862_ ^ new_A869_;
  assign new_A877_ = ~new_A886_ | ~new_A887_;
  assign new_A876_ = ~new_A861_ ^ new_A873_;
  assign new_A875_ = new_A883_ | new_A860_;
  assign new_A874_ = new_A880_ & new_A861_;
  assign new_A873_ = new_A882_ & new_A881_;
  assign new_A872_ = new_A877_ & new_A861_;
  assign new_A871_ = new_A879_ & new_A878_;
  assign new_A870_ = new_A871_ ^ new_A861_;
  assign new_A869_ = new_A859_ ^ new_A860_;
  assign A868 = new_A869_ & new_A876_;
  assign A867 = new_A869_ & new_A875_;
  assign A866 = new_A874_ | new_A873_;
  assign A865 = new_A872_ | new_A871_;
  assign A864 = new_A870_ & new_A869_;
  assign new_A863_ = new_A1461_;
  assign new_A862_ = new_A1428_;
  assign new_A861_ = new_A1395_;
  assign new_A860_ = new_A1362_;
  assign new_A859_ = new_A1329_;
  assign new_A858_ = new_A836_ & new_A851_;
  assign new_A857_ = ~new_A836_ & ~new_A858_;
  assign new_A856_ = new_A836_ | new_A851_;
  assign new_A855_ = ~new_A829_ | ~new_A830_;
  assign new_A854_ = new_A836_ | new_A851_;
  assign new_A853_ = ~new_A852_ & ~new_A836_;
  assign new_A852_ = new_A836_ & new_A851_;
  assign new_A851_ = ~new_A827_ | ~new_A828_;
  assign new_A850_ = new_A828_ & new_A840_;
  assign new_A849_ = new_A829_ | new_A836_;
  assign new_A848_ = new_A829_ | new_A830_;
  assign new_A847_ = ~new_A857_ | ~new_A856_;
  assign new_A846_ = new_A855_ & new_A848_;
  assign new_A845_ = new_A829_ ^ new_A836_;
  assign new_A844_ = ~new_A853_ | ~new_A854_;
  assign new_A843_ = ~new_A828_ ^ new_A840_;
  assign new_A842_ = new_A850_ | new_A827_;
  assign new_A841_ = new_A847_ & new_A828_;
  assign new_A840_ = new_A849_ & new_A848_;
  assign new_A839_ = new_A844_ & new_A828_;
  assign new_A838_ = new_A846_ & new_A845_;
  assign new_A837_ = new_A838_ ^ new_A828_;
  assign new_A836_ = new_A826_ ^ new_A827_;
  assign A835 = new_A836_ & new_A843_;
  assign A834 = new_A836_ & new_A842_;
  assign A833 = new_A841_ | new_A840_;
  assign A832 = new_A839_ | new_A838_;
  assign A831 = new_A837_ & new_A836_;
  assign new_A830_ = new_A1296_;
  assign new_A829_ = new_A1263_;
  assign new_A828_ = new_A1230_;
  assign new_A827_ = new_A1197_;
  assign new_A826_ = new_A1162_;
  assign new_A825_ = new_A803_ & new_A818_;
  assign new_A824_ = ~new_A803_ & ~new_A825_;
  assign new_A823_ = new_A803_ | new_A818_;
  assign new_A822_ = ~new_A796_ | ~new_A797_;
  assign new_A821_ = new_A803_ | new_A818_;
  assign new_A820_ = ~new_A819_ & ~new_A803_;
  assign new_A819_ = new_A803_ & new_A818_;
  assign new_A818_ = ~new_A794_ | ~new_A795_;
  assign new_A817_ = new_A795_ & new_A807_;
  assign new_A816_ = new_A796_ | new_A803_;
  assign new_A815_ = new_A796_ | new_A797_;
  assign new_A814_ = ~new_A824_ | ~new_A823_;
  assign new_A813_ = new_A822_ & new_A815_;
  assign new_A812_ = new_A796_ ^ new_A803_;
  assign new_A811_ = ~new_A820_ | ~new_A821_;
  assign new_A810_ = ~new_A795_ ^ new_A807_;
  assign new_A809_ = new_A817_ | new_A794_;
  assign new_A808_ = new_A814_ & new_A795_;
  assign new_A807_ = new_A816_ & new_A815_;
  assign new_A806_ = new_A811_ & new_A795_;
  assign new_A805_ = new_A813_ & new_A812_;
  assign new_A804_ = new_A805_ ^ new_A795_;
  assign new_A803_ = new_A793_ ^ new_A794_;
  assign A802 = new_A803_ & new_A810_;
  assign A801 = new_A803_ & new_A809_;
  assign A800 = new_A808_ | new_A807_;
  assign A799 = new_A806_ | new_A805_;
  assign A798 = new_A804_ & new_A803_;
  assign new_A797_ = new_A1955_;
  assign new_A796_ = new_A1922_;
  assign new_A795_ = new_A1889_;
  assign new_A794_ = new_A1856_;
  assign new_A793_ = new_A1823_;
  assign new_A792_ = new_A770_ & new_A785_;
  assign new_A791_ = ~new_A770_ & ~new_A792_;
  assign new_A790_ = new_A770_ | new_A785_;
  assign new_A789_ = ~new_A763_ | ~new_A764_;
  assign new_A788_ = new_A770_ | new_A785_;
  assign new_A787_ = ~new_A786_ & ~new_A770_;
  assign new_A786_ = new_A770_ & new_A785_;
  assign new_A785_ = ~new_A761_ | ~new_A762_;
  assign new_A784_ = new_A762_ & new_A774_;
  assign new_A783_ = new_A763_ | new_A770_;
  assign new_A782_ = new_A763_ | new_A764_;
  assign new_A781_ = ~new_A791_ | ~new_A790_;
  assign new_A780_ = new_A789_ & new_A782_;
  assign new_A779_ = new_A763_ ^ new_A770_;
  assign new_A778_ = ~new_A787_ | ~new_A788_;
  assign new_A777_ = ~new_A762_ ^ new_A774_;
  assign new_A776_ = new_A784_ | new_A761_;
  assign new_A775_ = new_A781_ & new_A762_;
  assign new_A774_ = new_A783_ & new_A782_;
  assign new_A773_ = new_A778_ & new_A762_;
  assign new_A772_ = new_A780_ & new_A779_;
  assign new_A771_ = new_A772_ ^ new_A762_;
  assign new_A770_ = new_A760_ ^ new_A761_;
  assign A769 = new_A770_ & new_A777_;
  assign A768 = new_A770_ & new_A776_;
  assign A767 = new_A775_ | new_A774_;
  assign A766 = new_A773_ | new_A772_;
  assign A765 = new_A771_ & new_A770_;
  assign new_A764_ = new_A1790_;
  assign new_A763_ = new_A1757_;
  assign new_A762_ = new_A1724_;
  assign new_A761_ = new_A1691_;
  assign new_A760_ = new_A1658_;
  assign new_A759_ = new_A737_ & new_A752_;
  assign new_A758_ = ~new_A737_ & ~new_A759_;
  assign new_A757_ = new_A737_ | new_A752_;
  assign new_A756_ = ~new_A730_ | ~new_A731_;
  assign new_A755_ = new_A737_ | new_A752_;
  assign new_A754_ = ~new_A753_ & ~new_A737_;
  assign new_A753_ = new_A737_ & new_A752_;
  assign new_A752_ = ~new_A728_ | ~new_A729_;
  assign new_A751_ = new_A729_ & new_A741_;
  assign new_A750_ = new_A730_ | new_A737_;
  assign new_A749_ = new_A730_ | new_A731_;
  assign new_A748_ = ~new_A758_ | ~new_A757_;
  assign new_A747_ = new_A756_ & new_A749_;
  assign new_A746_ = new_A730_ ^ new_A737_;
  assign new_A745_ = ~new_A754_ | ~new_A755_;
  assign new_A744_ = ~new_A729_ ^ new_A741_;
  assign new_A743_ = new_A751_ | new_A728_;
  assign new_A742_ = new_A748_ & new_A729_;
  assign new_A741_ = new_A750_ & new_A749_;
  assign new_A740_ = new_A745_ & new_A729_;
  assign new_A739_ = new_A747_ & new_A746_;
  assign new_A738_ = new_A739_ ^ new_A729_;
  assign new_A737_ = new_A727_ ^ new_A728_;
  assign A736 = new_A737_ & new_A744_;
  assign A735 = new_A737_ & new_A743_;
  assign A734 = new_A742_ | new_A741_;
  assign A733 = new_A740_ | new_A739_;
  assign A732 = new_A738_ & new_A737_;
  assign new_A731_ = new_A1625_;
  assign new_A730_ = new_A1592_;
  assign new_A729_ = new_A1559_;
  assign new_A728_ = new_A1526_;
  assign new_A727_ = new_A1493_;
  assign new_A726_ = new_A704_ & new_A719_;
  assign new_A725_ = ~new_A704_ & ~new_A726_;
  assign new_A724_ = new_A704_ | new_A719_;
  assign new_A723_ = ~new_A697_ | ~new_A698_;
  assign new_A722_ = new_A704_ | new_A719_;
  assign new_A721_ = ~new_A720_ & ~new_A704_;
  assign new_A720_ = new_A704_ & new_A719_;
  assign new_A719_ = ~new_A695_ | ~new_A696_;
  assign new_A718_ = new_A696_ & new_A708_;
  assign new_A717_ = new_A697_ | new_A704_;
  assign new_A716_ = new_A697_ | new_A698_;
  assign new_A715_ = ~new_A725_ | ~new_A724_;
  assign new_A714_ = new_A723_ & new_A716_;
  assign new_A713_ = new_A697_ ^ new_A704_;
  assign new_A712_ = ~new_A721_ | ~new_A722_;
  assign new_A711_ = ~new_A696_ ^ new_A708_;
  assign new_A710_ = new_A718_ | new_A695_;
  assign new_A709_ = new_A715_ & new_A696_;
  assign new_A708_ = new_A717_ & new_A716_;
  assign new_A707_ = new_A712_ & new_A696_;
  assign new_A706_ = new_A714_ & new_A713_;
  assign new_A705_ = new_A706_ ^ new_A696_;
  assign new_A704_ = new_A694_ ^ new_A695_;
  assign A703 = new_A704_ & new_A711_;
  assign A702 = new_A704_ & new_A710_;
  assign A701 = new_A709_ | new_A708_;
  assign A700 = new_A707_ | new_A706_;
  assign A699 = new_A705_ & new_A704_;
  assign new_A698_ = new_A1460_;
  assign new_A697_ = new_A1427_;
  assign new_A696_ = new_A1394_;
  assign new_A695_ = new_A1361_;
  assign new_A694_ = new_A1328_;
  assign new_A693_ = new_A671_ & new_A686_;
  assign new_A692_ = ~new_A671_ & ~new_A693_;
  assign new_A691_ = new_A671_ | new_A686_;
  assign new_A690_ = ~new_A664_ | ~new_A665_;
  assign new_A689_ = new_A671_ | new_A686_;
  assign new_A688_ = ~new_A687_ & ~new_A671_;
  assign new_A687_ = new_A671_ & new_A686_;
  assign new_A686_ = ~new_A662_ | ~new_A663_;
  assign new_A685_ = new_A663_ & new_A675_;
  assign new_A684_ = new_A664_ | new_A671_;
  assign new_A683_ = new_A664_ | new_A665_;
  assign new_A682_ = ~new_A692_ | ~new_A691_;
  assign new_A681_ = new_A690_ & new_A683_;
  assign new_A680_ = new_A664_ ^ new_A671_;
  assign new_A679_ = ~new_A688_ | ~new_A689_;
  assign new_A678_ = ~new_A663_ ^ new_A675_;
  assign new_A677_ = new_A685_ | new_A662_;
  assign new_A676_ = new_A682_ & new_A663_;
  assign new_A675_ = new_A684_ & new_A683_;
  assign new_A674_ = new_A679_ & new_A663_;
  assign new_A673_ = new_A681_ & new_A680_;
  assign new_A672_ = new_A673_ ^ new_A663_;
  assign new_A671_ = new_A661_ ^ new_A662_;
  assign A670 = new_A671_ & new_A678_;
  assign A669 = new_A671_ & new_A677_;
  assign A668 = new_A676_ | new_A675_;
  assign A667 = new_A674_ | new_A673_;
  assign A666 = new_A672_ & new_A671_;
  assign new_A665_ = new_A1295_;
  assign new_A664_ = new_A1262_;
  assign new_A663_ = new_A1229_;
  assign new_A662_ = new_A1196_;
  assign new_A661_ = new_A1163_;
  assign new_A660_ = new_A638_ & new_A653_;
  assign new_A659_ = ~new_A638_ & ~new_A660_;
  assign new_A658_ = new_A638_ | new_A653_;
  assign new_A657_ = ~new_A631_ | ~new_A632_;
  assign new_A656_ = new_A638_ | new_A653_;
  assign new_A655_ = ~new_A654_ & ~new_A638_;
  assign new_A654_ = new_A638_ & new_A653_;
  assign new_A653_ = ~new_A629_ | ~new_A630_;
  assign new_A652_ = new_A630_ & new_A642_;
  assign new_A651_ = new_A631_ | new_A638_;
  assign new_A650_ = new_A631_ | new_A632_;
  assign new_A649_ = ~new_A659_ | ~new_A658_;
  assign new_A648_ = new_A657_ & new_A650_;
  assign new_A647_ = new_A631_ ^ new_A638_;
  assign new_A646_ = ~new_A655_ | ~new_A656_;
  assign new_A645_ = ~new_A630_ ^ new_A642_;
  assign new_A644_ = new_A652_ | new_A629_;
  assign new_A643_ = new_A649_ & new_A630_;
  assign new_A642_ = new_A651_ & new_A650_;
  assign new_A641_ = new_A646_ & new_A630_;
  assign new_A640_ = new_A648_ & new_A647_;
  assign new_A639_ = new_A640_ ^ new_A630_;
  assign new_A638_ = new_A628_ ^ new_A629_;
  assign A637 = new_A638_ & new_A645_;
  assign A636 = new_A638_ & new_A644_;
  assign A635 = new_A643_ | new_A642_;
  assign A634 = new_A641_ | new_A640_;
  assign A633 = new_A639_ & new_A638_;
  assign new_A632_ = new_A1954_;
  assign new_A631_ = new_A1921_;
  assign new_A630_ = new_A1888_;
  assign new_A629_ = new_A1855_;
  assign new_A628_ = new_A1822_;
  assign new_A627_ = new_A605_ & new_A620_;
  assign new_A626_ = ~new_A605_ & ~new_A627_;
  assign new_A625_ = new_A605_ | new_A620_;
  assign new_A624_ = ~new_A598_ | ~new_A599_;
  assign new_A623_ = new_A605_ | new_A620_;
  assign new_A622_ = ~new_A621_ & ~new_A605_;
  assign new_A621_ = new_A605_ & new_A620_;
  assign new_A620_ = ~new_A596_ | ~new_A597_;
  assign new_A619_ = new_A597_ & new_A609_;
  assign new_A618_ = new_A598_ | new_A605_;
  assign new_A617_ = new_A598_ | new_A599_;
  assign new_A616_ = ~new_A626_ | ~new_A625_;
  assign new_A615_ = new_A624_ & new_A617_;
  assign new_A614_ = new_A598_ ^ new_A605_;
  assign new_A613_ = ~new_A622_ | ~new_A623_;
  assign new_A612_ = ~new_A597_ ^ new_A609_;
  assign new_A611_ = new_A619_ | new_A596_;
  assign new_A610_ = new_A616_ & new_A597_;
  assign new_A609_ = new_A618_ & new_A617_;
  assign new_A608_ = new_A613_ & new_A597_;
  assign new_A607_ = new_A615_ & new_A614_;
  assign new_A606_ = new_A607_ ^ new_A597_;
  assign new_A605_ = new_A595_ ^ new_A596_;
  assign A604 = new_A605_ & new_A612_;
  assign A603 = new_A605_ & new_A611_;
  assign A602 = new_A610_ | new_A609_;
  assign A601 = new_A608_ | new_A607_;
  assign A600 = new_A606_ & new_A605_;
  assign new_A599_ = new_A1789_;
  assign new_A598_ = new_A1756_;
  assign new_A597_ = new_A1723_;
  assign new_A596_ = new_A1690_;
  assign new_A595_ = new_A1657_;
  assign new_A594_ = new_A572_ & new_A587_;
  assign new_A593_ = ~new_A572_ & ~new_A594_;
  assign new_A592_ = new_A572_ | new_A587_;
  assign new_A591_ = ~new_A565_ | ~new_A566_;
  assign new_A590_ = new_A572_ | new_A587_;
  assign new_A589_ = ~new_A588_ & ~new_A572_;
  assign new_A588_ = new_A572_ & new_A587_;
  assign new_A587_ = ~new_A563_ | ~new_A564_;
  assign new_A586_ = new_A564_ & new_A576_;
  assign new_A585_ = new_A565_ | new_A572_;
  assign new_A584_ = new_A565_ | new_A566_;
  assign new_A583_ = ~new_A593_ | ~new_A592_;
  assign new_A582_ = new_A591_ & new_A584_;
  assign new_A581_ = new_A565_ ^ new_A572_;
  assign new_A580_ = ~new_A589_ | ~new_A590_;
  assign new_A579_ = ~new_A564_ ^ new_A576_;
  assign new_A578_ = new_A586_ | new_A563_;
  assign new_A577_ = new_A583_ & new_A564_;
  assign new_A576_ = new_A585_ & new_A584_;
  assign new_A575_ = new_A580_ & new_A564_;
  assign new_A574_ = new_A582_ & new_A581_;
  assign new_A573_ = new_A574_ ^ new_A564_;
  assign new_A572_ = new_A562_ ^ new_A563_;
  assign A571 = new_A572_ & new_A579_;
  assign A570 = new_A572_ & new_A578_;
  assign A569 = new_A577_ | new_A576_;
  assign A568 = new_A575_ | new_A574_;
  assign A567 = new_A573_ & new_A572_;
  assign new_A566_ = new_A1624_;
  assign new_A565_ = new_A1591_;
  assign new_A564_ = new_A1558_;
  assign new_A563_ = new_A1525_;
  assign new_A562_ = new_A1492_;
  assign new_A561_ = new_A539_ & new_A554_;
  assign new_A560_ = ~new_A539_ & ~new_A561_;
  assign new_A559_ = new_A539_ | new_A554_;
  assign new_A558_ = ~new_A532_ | ~new_A533_;
  assign new_A557_ = new_A539_ | new_A554_;
  assign new_A556_ = ~new_A555_ & ~new_A539_;
  assign new_A555_ = new_A539_ & new_A554_;
  assign new_A554_ = ~new_A530_ | ~new_A531_;
  assign new_A553_ = new_A531_ & new_A543_;
  assign new_A552_ = new_A532_ | new_A539_;
  assign new_A551_ = new_A532_ | new_A533_;
  assign new_A550_ = ~new_A560_ | ~new_A559_;
  assign new_A549_ = new_A558_ & new_A551_;
  assign new_A548_ = new_A532_ ^ new_A539_;
  assign new_A547_ = ~new_A556_ | ~new_A557_;
  assign new_A546_ = ~new_A531_ ^ new_A543_;
  assign new_A545_ = new_A553_ | new_A530_;
  assign new_A544_ = new_A550_ & new_A531_;
  assign new_A543_ = new_A552_ & new_A551_;
  assign new_A542_ = new_A547_ & new_A531_;
  assign new_A541_ = new_A549_ & new_A548_;
  assign new_A540_ = new_A541_ ^ new_A531_;
  assign new_A539_ = new_A529_ ^ new_A530_;
  assign A538 = new_A539_ & new_A546_;
  assign A537 = new_A539_ & new_A545_;
  assign A536 = new_A544_ | new_A543_;
  assign A535 = new_A542_ | new_A541_;
  assign A534 = new_A540_ & new_A539_;
  assign new_A533_ = new_A1459_;
  assign new_A532_ = new_A1426_;
  assign new_A531_ = new_A1393_;
  assign new_A530_ = new_A1360_;
  assign new_A529_ = new_A1327_;
  assign new_A528_ = new_A506_ & new_A521_;
  assign new_A527_ = ~new_A506_ & ~new_A528_;
  assign new_A526_ = new_A506_ | new_A521_;
  assign new_A525_ = ~new_A499_ | ~new_A500_;
  assign new_A524_ = new_A506_ | new_A521_;
  assign new_A523_ = ~new_A522_ & ~new_A506_;
  assign new_A522_ = new_A506_ & new_A521_;
  assign new_A521_ = ~new_A497_ | ~new_A498_;
  assign new_A520_ = new_A498_ & new_A510_;
  assign new_A519_ = new_A499_ | new_A506_;
  assign new_A518_ = new_A499_ | new_A500_;
  assign new_A517_ = ~new_A527_ | ~new_A526_;
  assign new_A516_ = new_A525_ & new_A518_;
  assign new_A515_ = new_A499_ ^ new_A506_;
  assign new_A514_ = ~new_A523_ | ~new_A524_;
  assign new_A513_ = ~new_A498_ ^ new_A510_;
  assign new_A512_ = new_A520_ | new_A497_;
  assign new_A511_ = new_A517_ & new_A498_;
  assign new_A510_ = new_A519_ & new_A518_;
  assign new_A509_ = new_A514_ & new_A498_;
  assign new_A508_ = new_A516_ & new_A515_;
  assign new_A507_ = new_A508_ ^ new_A498_;
  assign new_A506_ = new_A496_ ^ new_A497_;
  assign A505 = new_A506_ & new_A513_;
  assign A504 = new_A506_ & new_A512_;
  assign A503 = new_A511_ | new_A510_;
  assign A502 = new_A509_ | new_A508_;
  assign A501 = new_A507_ & new_A506_;
  assign new_A500_ = new_A1294_;
  assign new_A499_ = new_A1261_;
  assign new_A498_ = new_A1228_;
  assign new_A497_ = new_A1195_;
  assign new_A496_ = new_A1164_;
  assign new_A495_ = new_A473_ & new_A488_;
  assign new_A494_ = ~new_A473_ & ~new_A495_;
  assign new_A493_ = new_A473_ | new_A488_;
  assign new_A492_ = ~new_A466_ | ~new_A467_;
  assign new_A491_ = new_A473_ | new_A488_;
  assign new_A490_ = ~new_A489_ & ~new_A473_;
  assign new_A489_ = new_A473_ & new_A488_;
  assign new_A488_ = ~new_A464_ | ~new_A465_;
  assign new_A487_ = new_A465_ & new_A477_;
  assign new_A486_ = new_A466_ | new_A473_;
  assign new_A485_ = new_A466_ | new_A467_;
  assign new_A484_ = ~new_A494_ | ~new_A493_;
  assign new_A483_ = new_A492_ & new_A485_;
  assign new_A482_ = new_A466_ ^ new_A473_;
  assign new_A481_ = ~new_A490_ | ~new_A491_;
  assign new_A480_ = ~new_A465_ ^ new_A477_;
  assign new_A479_ = new_A487_ | new_A464_;
  assign new_A478_ = new_A484_ & new_A465_;
  assign new_A477_ = new_A486_ & new_A485_;
  assign new_A476_ = new_A481_ & new_A465_;
  assign new_A475_ = new_A483_ & new_A482_;
  assign new_A474_ = new_A475_ ^ new_A465_;
  assign new_A473_ = new_A463_ ^ new_A464_;
  assign A472 = new_A473_ & new_A480_;
  assign A471 = new_A473_ & new_A479_;
  assign A470 = new_A478_ | new_A477_;
  assign A469 = new_A476_ | new_A475_;
  assign A468 = new_A474_ & new_A473_;
  assign new_A467_ = new_A1953_;
  assign new_A466_ = new_A1920_;
  assign new_A465_ = new_A1887_;
  assign new_A464_ = new_A1854_;
  assign new_A463_ = new_A1821_;
  assign new_A462_ = new_A440_ & new_A455_;
  assign new_A461_ = ~new_A440_ & ~new_A462_;
  assign new_A460_ = new_A440_ | new_A455_;
  assign new_A459_ = ~new_A433_ | ~new_A434_;
  assign new_A458_ = new_A440_ | new_A455_;
  assign new_A457_ = ~new_A456_ & ~new_A440_;
  assign new_A456_ = new_A440_ & new_A455_;
  assign new_A455_ = ~new_A431_ | ~new_A432_;
  assign new_A454_ = new_A432_ & new_A444_;
  assign new_A453_ = new_A433_ | new_A440_;
  assign new_A452_ = new_A433_ | new_A434_;
  assign new_A451_ = ~new_A461_ | ~new_A460_;
  assign new_A450_ = new_A459_ & new_A452_;
  assign new_A449_ = new_A433_ ^ new_A440_;
  assign new_A448_ = ~new_A457_ | ~new_A458_;
  assign new_A447_ = ~new_A432_ ^ new_A444_;
  assign new_A446_ = new_A454_ | new_A431_;
  assign new_A445_ = new_A451_ & new_A432_;
  assign new_A444_ = new_A453_ & new_A452_;
  assign new_A443_ = new_A448_ & new_A432_;
  assign new_A442_ = new_A450_ & new_A449_;
  assign new_A441_ = new_A442_ ^ new_A432_;
  assign new_A440_ = new_A430_ ^ new_A431_;
  assign A439 = new_A440_ & new_A447_;
  assign A438 = new_A440_ & new_A446_;
  assign A437 = new_A445_ | new_A444_;
  assign A436 = new_A443_ | new_A442_;
  assign A435 = new_A441_ & new_A440_;
  assign new_A434_ = new_A1788_;
  assign new_A433_ = new_A1755_;
  assign new_A432_ = new_A1722_;
  assign new_A431_ = new_A1689_;
  assign new_A430_ = new_A1656_;
  assign new_A429_ = new_A407_ & new_A422_;
  assign new_A428_ = ~new_A407_ & ~new_A429_;
  assign new_A427_ = new_A407_ | new_A422_;
  assign new_A426_ = ~new_A400_ | ~new_A401_;
  assign new_A425_ = new_A407_ | new_A422_;
  assign new_A424_ = ~new_A423_ & ~new_A407_;
  assign new_A423_ = new_A407_ & new_A422_;
  assign new_A422_ = ~new_A398_ | ~new_A399_;
  assign new_A421_ = new_A399_ & new_A411_;
  assign new_A420_ = new_A400_ | new_A407_;
  assign new_A419_ = new_A400_ | new_A401_;
  assign new_A418_ = ~new_A428_ | ~new_A427_;
  assign new_A417_ = new_A426_ & new_A419_;
  assign new_A416_ = new_A400_ ^ new_A407_;
  assign new_A415_ = ~new_A424_ | ~new_A425_;
  assign new_A414_ = ~new_A399_ ^ new_A411_;
  assign new_A413_ = new_A421_ | new_A398_;
  assign new_A412_ = new_A418_ & new_A399_;
  assign new_A411_ = new_A420_ & new_A419_;
  assign new_A410_ = new_A415_ & new_A399_;
  assign new_A409_ = new_A417_ & new_A416_;
  assign new_A408_ = new_A409_ ^ new_A399_;
  assign new_A407_ = new_A397_ ^ new_A398_;
  assign A406 = new_A407_ & new_A414_;
  assign A405 = new_A407_ & new_A413_;
  assign A404 = new_A412_ | new_A411_;
  assign A403 = new_A410_ | new_A409_;
  assign A402 = new_A408_ & new_A407_;
  assign new_A401_ = new_A1623_;
  assign new_A400_ = new_A1590_;
  assign new_A399_ = new_A1557_;
  assign new_A398_ = new_A1524_;
  assign new_A397_ = new_A1491_;
  assign new_A396_ = new_A374_ & new_A389_;
  assign new_A395_ = ~new_A374_ & ~new_A396_;
  assign new_A394_ = new_A374_ | new_A389_;
  assign new_A393_ = ~new_A367_ | ~new_A368_;
  assign new_A392_ = new_A374_ | new_A389_;
  assign new_A391_ = ~new_A390_ & ~new_A374_;
  assign new_A390_ = new_A374_ & new_A389_;
  assign new_A389_ = ~new_A365_ | ~new_A366_;
  assign new_A388_ = new_A366_ & new_A378_;
  assign new_A387_ = new_A367_ | new_A374_;
  assign new_A386_ = new_A367_ | new_A368_;
  assign new_A385_ = ~new_A395_ | ~new_A394_;
  assign new_A384_ = new_A393_ & new_A386_;
  assign new_A383_ = new_A367_ ^ new_A374_;
  assign new_A382_ = ~new_A391_ | ~new_A392_;
  assign new_A381_ = ~new_A366_ ^ new_A378_;
  assign new_A380_ = new_A388_ | new_A365_;
  assign new_A379_ = new_A385_ & new_A366_;
  assign new_A378_ = new_A387_ & new_A386_;
  assign new_A377_ = new_A382_ & new_A366_;
  assign new_A376_ = new_A384_ & new_A383_;
  assign new_A375_ = new_A376_ ^ new_A366_;
  assign new_A374_ = new_A364_ ^ new_A365_;
  assign A373 = new_A374_ & new_A381_;
  assign A372 = new_A374_ & new_A380_;
  assign A371 = new_A379_ | new_A378_;
  assign A370 = new_A377_ | new_A376_;
  assign A369 = new_A375_ & new_A374_;
  assign new_A368_ = new_A1458_;
  assign new_A367_ = new_A1425_;
  assign new_A366_ = new_A1392_;
  assign new_A365_ = new_A1359_;
  assign new_A364_ = new_A1326_;
  assign new_A331_ = new_A1293_;
  assign new_A332_ = new_A1260_;
  assign new_A333_ = new_A1227_;
  assign new_A334_ = new_A1194_;
  assign new_A335_ = new_A1165_;
  assign A336 = new_A342_ & new_A341_;
  assign A337 = new_A344_ | new_A343_;
  assign A338 = new_A346_ | new_A345_;
  assign A339 = new_A341_ & new_A347_;
  assign A340 = new_A341_ & new_A348_;
  assign new_A341_ = new_A331_ ^ new_A332_;
  assign new_A342_ = new_A343_ ^ new_A333_;
  assign new_A343_ = new_A351_ & new_A350_;
  assign new_A344_ = new_A349_ & new_A333_;
  assign new_A345_ = new_A354_ & new_A353_;
  assign new_A346_ = new_A352_ & new_A333_;
  assign new_A347_ = new_A355_ | new_A332_;
  assign new_A348_ = ~new_A333_ ^ new_A345_;
  assign new_A349_ = ~new_A358_ | ~new_A359_;
  assign new_A350_ = new_A334_ ^ new_A341_;
  assign new_A351_ = new_A360_ & new_A353_;
  assign new_A352_ = ~new_A362_ | ~new_A361_;
  assign new_A353_ = new_A334_ | new_A335_;
  assign new_A354_ = new_A334_ | new_A341_;
  assign new_A355_ = new_A333_ & new_A345_;
  assign new_A356_ = ~new_A332_ | ~new_A333_;
  assign new_A357_ = new_A341_ & new_A356_;
  assign new_A358_ = ~new_A357_ & ~new_A341_;
  assign new_A359_ = new_A341_ | new_A356_;
  assign new_A360_ = ~new_A334_ | ~new_A335_;
  assign new_A361_ = new_A341_ | new_A356_;
  assign new_A362_ = ~new_A341_ & ~new_A363_;
  assign new_A363_ = new_A341_ & new_A356_;
endmodule


