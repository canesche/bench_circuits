module DES ( 
    \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
    \data_in<2> , \data_in<1> , \data_in<0> , \reset<0> , \encrypt<0> ,
    \load_key<0> , \inreg<55> , \inreg<54> , \inreg<53> , \inreg<52> ,
    \inreg<51> , \inreg<50> , \inreg<49> , \inreg<48> , \inreg<47> ,
    \inreg<46> , \inreg<45> , \inreg<44> , \inreg<43> , \inreg<42> ,
    \inreg<41> , \inreg<40> , \inreg<39> , \inreg<38> , \inreg<37> ,
    \inreg<36> , \inreg<35> , \inreg<34> , \inreg<33> , \inreg<32> ,
    \inreg<31> , \inreg<30> , \inreg<29> , \inreg<28> , \inreg<27> ,
    \inreg<26> , \inreg<25> , \inreg<24> , \inreg<23> , \inreg<22> ,
    \inreg<21> , \inreg<20> , \inreg<19> , \inreg<18> , \inreg<17> ,
    \inreg<16> , \inreg<15> , \inreg<14> , \inreg<13> , \inreg<12> ,
    \inreg<11> , \inreg<10> , \inreg<9> , \inreg<8> , \inreg<7> ,
    \inreg<6> , \inreg<5> , \inreg<4> , \inreg<3> , \inreg<2> , \inreg<1> ,
    \inreg<0> , \outreg<63> , \outreg<62> , \outreg<61> , \outreg<60> ,
    \outreg<59> , \outreg<58> , \outreg<57> , \outreg<56> , \outreg<55> ,
    \outreg<54> , \outreg<53> , \outreg<52> , \outreg<51> , \outreg<50> ,
    \outreg<49> , \outreg<48> , \outreg<47> , \outreg<46> , \outreg<45> ,
    \outreg<44> , \outreg<43> , \outreg<42> , \outreg<41> , \outreg<40> ,
    \outreg<39> , \outreg<38> , \outreg<37> , \outreg<36> , \outreg<35> ,
    \outreg<34> , \outreg<33> , \outreg<32> , \outreg<31> , \outreg<30> ,
    \outreg<29> , \outreg<28> , \outreg<27> , \outreg<26> , \outreg<25> ,
    \outreg<24> , \outreg<23> , \outreg<22> , \outreg<21> , \outreg<20> ,
    \outreg<19> , \outreg<18> , \outreg<17> , \outreg<16> , \outreg<15> ,
    \outreg<14> , \outreg<13> , \outreg<12> , \outreg<11> , \outreg<10> ,
    \outreg<9> , \outreg<8> , \outreg<7> , \outreg<6> , \outreg<5> ,
    \outreg<4> , \outreg<3> , \outreg<2> , \outreg<1> , \outreg<0> ,
    \data<63> , \data<62> , \data<61> , \data<60> , \data<59> , \data<58> ,
    \data<57> , \data<56> , \data<55> , \data<54> , \data<53> , \data<52> ,
    \data<51> , \data<50> , \data<49> , \data<48> , \data<47> , \data<46> ,
    \data<45> , \data<44> , \data<43> , \data<42> , \data<41> , \data<40> ,
    \data<39> , \data<38> , \data<37> , \data<36> , \data<35> , \data<34> ,
    \data<33> , \data<32> , \data<31> , \data<30> , \data<29> , \data<28> ,
    \data<27> , \data<26> , \data<25> , \data<24> , \data<23> , \data<22> ,
    \data<21> , \data<20> , \data<19> , \data<18> , \data<17> , \data<16> ,
    \data<15> , \data<14> , \data<13> , \data<12> , \data<11> , \data<10> ,
    \data<9> , \data<8> , \data<7> , \data<6> , \data<5> , \data<4> ,
    \data<3> , \data<2> , \data<1> , \data<0> , \count<3> , \count<2> ,
    \count<1> , \count<0> , \C<27> , \C<26> , \C<25> , \C<24> , \C<23> ,
    \C<22> , \C<21> , \C<20> , \C<19> , \C<18> , \C<17> , \C<16> , \C<15> ,
    \C<14> , \C<13> , \C<12> , \C<11> , \C<10> , \C<9> , \C<8> , \C<7> ,
    \C<6> , \C<5> , \C<4> , \C<3> , \C<2> , \C<1> , \C<0> , \D<27> ,
    \D<26> , \D<25> , \D<24> , \D<23> , \D<22> , \D<21> , \D<20> , \D<19> ,
    \D<18> , \D<17> , \D<16> , \D<15> , \D<14> , \D<13> , \D<12> , \D<11> ,
    \D<10> , \D<9> , \D<8> , \D<7> , \D<6> , \D<5> , \D<4> , \D<3> ,
    \D<2> , \D<1> , \D<0> , \encrypt_mode<0> ,
    \inreg_new<55> , \inreg_new<54> , \inreg_new<53> , \inreg_new<52> ,
    \inreg_new<51> , \inreg_new<50> , \inreg_new<49> , \inreg_new<48> ,
    \inreg_new<47> , \inreg_new<46> , \inreg_new<45> , \inreg_new<44> ,
    \inreg_new<43> , \inreg_new<42> , \inreg_new<41> , \inreg_new<40> ,
    \inreg_new<39> , \inreg_new<38> , \inreg_new<37> , \inreg_new<36> ,
    \inreg_new<35> , \inreg_new<34> , \inreg_new<33> , \inreg_new<32> ,
    \inreg_new<31> , \inreg_new<30> , \inreg_new<29> , \inreg_new<28> ,
    \inreg_new<27> , \inreg_new<26> , \inreg_new<25> , \inreg_new<24> ,
    \inreg_new<23> , \inreg_new<22> , \inreg_new<21> , \inreg_new<20> ,
    \inreg_new<19> , \inreg_new<18> , \inreg_new<17> , \inreg_new<16> ,
    \inreg_new<15> , \inreg_new<14> , \inreg_new<13> , \inreg_new<12> ,
    \inreg_new<11> , \inreg_new<10> , \inreg_new<9> , \inreg_new<8> ,
    \inreg_new<7> , \inreg_new<6> , \inreg_new<5> , \inreg_new<4> ,
    \inreg_new<3> , \inreg_new<2> , \inreg_new<1> , \inreg_new<0> ,
    \outreg_new<63> , \outreg_new<62> , \outreg_new<61> , \outreg_new<60> ,
    \outreg_new<59> , \outreg_new<58> , \outreg_new<57> , \outreg_new<56> ,
    \outreg_new<55> , \outreg_new<54> , \outreg_new<53> , \outreg_new<52> ,
    \outreg_new<51> , \outreg_new<50> , \outreg_new<49> , \outreg_new<48> ,
    \outreg_new<47> , \outreg_new<46> , \outreg_new<45> , \outreg_new<44> ,
    \outreg_new<43> , \outreg_new<42> , \outreg_new<41> , \outreg_new<40> ,
    \outreg_new<39> , \outreg_new<38> , \outreg_new<37> , \outreg_new<36> ,
    \outreg_new<35> , \outreg_new<34> , \outreg_new<33> , \outreg_new<32> ,
    \outreg_new<31> , \outreg_new<30> , \outreg_new<29> , \outreg_new<28> ,
    \outreg_new<27> , \outreg_new<26> , \outreg_new<25> , \outreg_new<24> ,
    \outreg_new<23> , \outreg_new<22> , \outreg_new<21> , \outreg_new<20> ,
    \outreg_new<19> , \outreg_new<18> , \outreg_new<17> , \outreg_new<16> ,
    \outreg_new<15> , \outreg_new<14> , \outreg_new<13> , \outreg_new<12> ,
    \outreg_new<11> , \outreg_new<10> , \outreg_new<9> , \outreg_new<8> ,
    \outreg_new<7> , \outreg_new<6> , \outreg_new<5> , \outreg_new<4> ,
    \outreg_new<3> , \outreg_new<2> , \outreg_new<1> , \outreg_new<0> ,
    \data_new<63> , \data_new<62> , \data_new<61> , \data_new<60> ,
    \data_new<59> , \data_new<58> , \data_new<57> , \data_new<56> ,
    \data_new<55> , \data_new<54> , \data_new<53> , \data_new<52> ,
    \data_new<51> , \data_new<50> , \data_new<49> , \data_new<48> ,
    \data_new<47> , \data_new<46> , \data_new<45> , \data_new<44> ,
    \data_new<43> , \data_new<42> , \data_new<41> , \data_new<40> ,
    \data_new<39> , \data_new<38> , \data_new<37> , \data_new<36> ,
    \data_new<35> , \data_new<34> , \data_new<33> , \data_new<32> ,
    \data_new<31> , \data_new<30> , \data_new<29> , \data_new<28> ,
    \data_new<27> , \data_new<26> , \data_new<25> , \data_new<24> ,
    \data_new<23> , \data_new<22> , \data_new<21> , \data_new<20> ,
    \data_new<19> , \data_new<18> , \data_new<17> , \data_new<16> ,
    \data_new<15> , \data_new<14> , \data_new<13> , \data_new<12> ,
    \data_new<11> , \data_new<10> , \data_new<9> , \data_new<8> ,
    \data_new<7> , \data_new<6> , \data_new<5> , \data_new<4> ,
    \data_new<3> , \data_new<2> , \data_new<1> , \data_new<0> ,
    \count_new<3> , \count_new<2> , \count_new<1> , \count_new<0> ,
    \C_new<27> , \C_new<26> , \C_new<25> , \C_new<24> , \C_new<23> ,
    \C_new<22> , \C_new<21> , \C_new<20> , \C_new<19> , \C_new<18> ,
    \C_new<17> , \C_new<16> , \C_new<15> , \C_new<14> , \C_new<13> ,
    \C_new<12> , \C_new<11> , \C_new<10> , \C_new<9> , \C_new<8> ,
    \C_new<7> , \C_new<6> , \C_new<5> , \C_new<4> , \C_new<3> , \C_new<2> ,
    \C_new<1> , \C_new<0> , \D_new<27> , \D_new<26> , \D_new<25> ,
    \D_new<24> , \D_new<23> , \D_new<22> , \D_new<21> , \D_new<20> ,
    \D_new<19> , \D_new<18> , \D_new<17> , \D_new<16> , \D_new<15> ,
    \D_new<14> , \D_new<13> , \D_new<12> , \D_new<11> , \D_new<10> ,
    \D_new<9> , \D_new<8> , \D_new<7> , \D_new<6> , \D_new<5> , \D_new<4> ,
    \D_new<3> , \D_new<2> , \D_new<1> , \D_new<0> , \encrypt_mode_new<0>   );
  input  \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
    \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , \reset<0> ,
    \encrypt<0> , \load_key<0> , \inreg<55> , \inreg<54> , \inreg<53> ,
    \inreg<52> , \inreg<51> , \inreg<50> , \inreg<49> , \inreg<48> ,
    \inreg<47> , \inreg<46> , \inreg<45> , \inreg<44> , \inreg<43> ,
    \inreg<42> , \inreg<41> , \inreg<40> , \inreg<39> , \inreg<38> ,
    \inreg<37> , \inreg<36> , \inreg<35> , \inreg<34> , \inreg<33> ,
    \inreg<32> , \inreg<31> , \inreg<30> , \inreg<29> , \inreg<28> ,
    \inreg<27> , \inreg<26> , \inreg<25> , \inreg<24> , \inreg<23> ,
    \inreg<22> , \inreg<21> , \inreg<20> , \inreg<19> , \inreg<18> ,
    \inreg<17> , \inreg<16> , \inreg<15> , \inreg<14> , \inreg<13> ,
    \inreg<12> , \inreg<11> , \inreg<10> , \inreg<9> , \inreg<8> ,
    \inreg<7> , \inreg<6> , \inreg<5> , \inreg<4> , \inreg<3> , \inreg<2> ,
    \inreg<1> , \inreg<0> , \outreg<63> , \outreg<62> , \outreg<61> ,
    \outreg<60> , \outreg<59> , \outreg<58> , \outreg<57> , \outreg<56> ,
    \outreg<55> , \outreg<54> , \outreg<53> , \outreg<52> , \outreg<51> ,
    \outreg<50> , \outreg<49> , \outreg<48> , \outreg<47> , \outreg<46> ,
    \outreg<45> , \outreg<44> , \outreg<43> , \outreg<42> , \outreg<41> ,
    \outreg<40> , \outreg<39> , \outreg<38> , \outreg<37> , \outreg<36> ,
    \outreg<35> , \outreg<34> , \outreg<33> , \outreg<32> , \outreg<31> ,
    \outreg<30> , \outreg<29> , \outreg<28> , \outreg<27> , \outreg<26> ,
    \outreg<25> , \outreg<24> , \outreg<23> , \outreg<22> , \outreg<21> ,
    \outreg<20> , \outreg<19> , \outreg<18> , \outreg<17> , \outreg<16> ,
    \outreg<15> , \outreg<14> , \outreg<13> , \outreg<12> , \outreg<11> ,
    \outreg<10> , \outreg<9> , \outreg<8> , \outreg<7> , \outreg<6> ,
    \outreg<5> , \outreg<4> , \outreg<3> , \outreg<2> , \outreg<1> ,
    \outreg<0> , \data<63> , \data<62> , \data<61> , \data<60> ,
    \data<59> , \data<58> , \data<57> , \data<56> , \data<55> , \data<54> ,
    \data<53> , \data<52> , \data<51> , \data<50> , \data<49> , \data<48> ,
    \data<47> , \data<46> , \data<45> , \data<44> , \data<43> , \data<42> ,
    \data<41> , \data<40> , \data<39> , \data<38> , \data<37> , \data<36> ,
    \data<35> , \data<34> , \data<33> , \data<32> , \data<31> , \data<30> ,
    \data<29> , \data<28> , \data<27> , \data<26> , \data<25> , \data<24> ,
    \data<23> , \data<22> , \data<21> , \data<20> , \data<19> , \data<18> ,
    \data<17> , \data<16> , \data<15> , \data<14> , \data<13> , \data<12> ,
    \data<11> , \data<10> , \data<9> , \data<8> , \data<7> , \data<6> ,
    \data<5> , \data<4> , \data<3> , \data<2> , \data<1> , \data<0> ,
    \count<3> , \count<2> , \count<1> , \count<0> , \C<27> , \C<26> ,
    \C<25> , \C<24> , \C<23> , \C<22> , \C<21> , \C<20> , \C<19> , \C<18> ,
    \C<17> , \C<16> , \C<15> , \C<14> , \C<13> , \C<12> , \C<11> , \C<10> ,
    \C<9> , \C<8> , \C<7> , \C<6> , \C<5> , \C<4> , \C<3> , \C<2> , \C<1> ,
    \C<0> , \D<27> , \D<26> , \D<25> , \D<24> , \D<23> , \D<22> , \D<21> ,
    \D<20> , \D<19> , \D<18> , \D<17> , \D<16> , \D<15> , \D<14> , \D<13> ,
    \D<12> , \D<11> , \D<10> , \D<9> , \D<8> , \D<7> , \D<6> , \D<5> ,
    \D<4> , \D<3> , \D<2> , \D<1> , \D<0> , \encrypt_mode<0> ;
  output \inreg_new<55> , \inreg_new<54> , \inreg_new<53> , \inreg_new<52> ,
    \inreg_new<51> , \inreg_new<50> , \inreg_new<49> , \inreg_new<48> ,
    \inreg_new<47> , \inreg_new<46> , \inreg_new<45> , \inreg_new<44> ,
    \inreg_new<43> , \inreg_new<42> , \inreg_new<41> , \inreg_new<40> ,
    \inreg_new<39> , \inreg_new<38> , \inreg_new<37> , \inreg_new<36> ,
    \inreg_new<35> , \inreg_new<34> , \inreg_new<33> , \inreg_new<32> ,
    \inreg_new<31> , \inreg_new<30> , \inreg_new<29> , \inreg_new<28> ,
    \inreg_new<27> , \inreg_new<26> , \inreg_new<25> , \inreg_new<24> ,
    \inreg_new<23> , \inreg_new<22> , \inreg_new<21> , \inreg_new<20> ,
    \inreg_new<19> , \inreg_new<18> , \inreg_new<17> , \inreg_new<16> ,
    \inreg_new<15> , \inreg_new<14> , \inreg_new<13> , \inreg_new<12> ,
    \inreg_new<11> , \inreg_new<10> , \inreg_new<9> , \inreg_new<8> ,
    \inreg_new<7> , \inreg_new<6> , \inreg_new<5> , \inreg_new<4> ,
    \inreg_new<3> , \inreg_new<2> , \inreg_new<1> , \inreg_new<0> ,
    \outreg_new<63> , \outreg_new<62> , \outreg_new<61> , \outreg_new<60> ,
    \outreg_new<59> , \outreg_new<58> , \outreg_new<57> , \outreg_new<56> ,
    \outreg_new<55> , \outreg_new<54> , \outreg_new<53> , \outreg_new<52> ,
    \outreg_new<51> , \outreg_new<50> , \outreg_new<49> , \outreg_new<48> ,
    \outreg_new<47> , \outreg_new<46> , \outreg_new<45> , \outreg_new<44> ,
    \outreg_new<43> , \outreg_new<42> , \outreg_new<41> , \outreg_new<40> ,
    \outreg_new<39> , \outreg_new<38> , \outreg_new<37> , \outreg_new<36> ,
    \outreg_new<35> , \outreg_new<34> , \outreg_new<33> , \outreg_new<32> ,
    \outreg_new<31> , \outreg_new<30> , \outreg_new<29> , \outreg_new<28> ,
    \outreg_new<27> , \outreg_new<26> , \outreg_new<25> , \outreg_new<24> ,
    \outreg_new<23> , \outreg_new<22> , \outreg_new<21> , \outreg_new<20> ,
    \outreg_new<19> , \outreg_new<18> , \outreg_new<17> , \outreg_new<16> ,
    \outreg_new<15> , \outreg_new<14> , \outreg_new<13> , \outreg_new<12> ,
    \outreg_new<11> , \outreg_new<10> , \outreg_new<9> , \outreg_new<8> ,
    \outreg_new<7> , \outreg_new<6> , \outreg_new<5> , \outreg_new<4> ,
    \outreg_new<3> , \outreg_new<2> , \outreg_new<1> , \outreg_new<0> ,
    \data_new<63> , \data_new<62> , \data_new<61> , \data_new<60> ,
    \data_new<59> , \data_new<58> , \data_new<57> , \data_new<56> ,
    \data_new<55> , \data_new<54> , \data_new<53> , \data_new<52> ,
    \data_new<51> , \data_new<50> , \data_new<49> , \data_new<48> ,
    \data_new<47> , \data_new<46> , \data_new<45> , \data_new<44> ,
    \data_new<43> , \data_new<42> , \data_new<41> , \data_new<40> ,
    \data_new<39> , \data_new<38> , \data_new<37> , \data_new<36> ,
    \data_new<35> , \data_new<34> , \data_new<33> , \data_new<32> ,
    \data_new<31> , \data_new<30> , \data_new<29> , \data_new<28> ,
    \data_new<27> , \data_new<26> , \data_new<25> , \data_new<24> ,
    \data_new<23> , \data_new<22> , \data_new<21> , \data_new<20> ,
    \data_new<19> , \data_new<18> , \data_new<17> , \data_new<16> ,
    \data_new<15> , \data_new<14> , \data_new<13> , \data_new<12> ,
    \data_new<11> , \data_new<10> , \data_new<9> , \data_new<8> ,
    \data_new<7> , \data_new<6> , \data_new<5> , \data_new<4> ,
    \data_new<3> , \data_new<2> , \data_new<1> , \data_new<0> ,
    \count_new<3> , \count_new<2> , \count_new<1> , \count_new<0> ,
    \C_new<27> , \C_new<26> , \C_new<25> , \C_new<24> , \C_new<23> ,
    \C_new<22> , \C_new<21> , \C_new<20> , \C_new<19> , \C_new<18> ,
    \C_new<17> , \C_new<16> , \C_new<15> , \C_new<14> , \C_new<13> ,
    \C_new<12> , \C_new<11> , \C_new<10> , \C_new<9> , \C_new<8> ,
    \C_new<7> , \C_new<6> , \C_new<5> , \C_new<4> , \C_new<3> , \C_new<2> ,
    \C_new<1> , \C_new<0> , \D_new<27> , \D_new<26> , \D_new<25> ,
    \D_new<24> , \D_new<23> , \D_new<22> , \D_new<21> , \D_new<20> ,
    \D_new<19> , \D_new<18> , \D_new<17> , \D_new<16> , \D_new<15> ,
    \D_new<14> , \D_new<13> , \D_new<12> , \D_new<11> , \D_new<10> ,
    \D_new<9> , \D_new<8> , \D_new<7> , \D_new<6> , \D_new<5> , \D_new<4> ,
    \D_new<3> , \D_new<2> , \D_new<1> , \D_new<0> , \encrypt_mode_new<0> ;
  wire new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n509_, new_n510_, new_n511_, new_n513_, new_n514_, new_n515_,
    new_n517_, new_n518_, new_n519_, new_n521_, new_n522_, new_n523_,
    new_n525_, new_n526_, new_n527_, new_n529_, new_n530_, new_n531_,
    new_n533_, new_n534_, new_n535_, new_n537_, new_n538_, new_n539_,
    new_n541_, new_n542_, new_n543_, new_n545_, new_n546_, new_n547_,
    new_n549_, new_n550_, new_n551_, new_n553_, new_n554_, new_n555_,
    new_n557_, new_n558_, new_n559_, new_n561_, new_n562_, new_n563_,
    new_n565_, new_n566_, new_n567_, new_n569_, new_n570_, new_n571_,
    new_n573_, new_n574_, new_n575_, new_n577_, new_n578_, new_n579_,
    new_n581_, new_n582_, new_n583_, new_n585_, new_n586_, new_n587_,
    new_n589_, new_n590_, new_n591_, new_n593_, new_n594_, new_n595_,
    new_n597_, new_n598_, new_n599_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n613_, new_n614_, new_n615_, new_n617_, new_n618_, new_n619_,
    new_n621_, new_n622_, new_n623_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n645_, new_n646_, new_n647_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1022_,
    new_n1023_, new_n1024_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1088_, new_n1089_, new_n1090_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1235_, new_n1236_,
    new_n1237_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_,
    new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_,
    new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_,
    new_n1598_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_,
    new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_,
    new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_,
    new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_,
    new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_,
    new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_,
    new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_,
    new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_,
    new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_,
    new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_,
    new_n1756_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_,
    new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_,
    new_n1914_, new_n1915_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_,
    new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_,
    new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_,
    new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_,
    new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1989_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_,
    new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_,
    new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_,
    new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_,
    new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_,
    new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_,
    new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_,
    new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_,
    new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2124_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2168_,
    new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2174_, new_n2175_,
    new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_,
    new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_,
    new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_,
    new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_,
    new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_,
    new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_,
    new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_,
    new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_,
    new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_,
    new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_,
    new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_,
    new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_,
    new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_,
    new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_,
    new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_,
    new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_,
    new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_,
    new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_,
    new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_,
    new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_,
    new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_,
    new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_,
    new_n2314_, new_n2315_, new_n2316_, new_n2318_, new_n2319_, new_n2320_,
    new_n2321_, new_n2322_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_,
    new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_,
    new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_,
    new_n2376_, new_n2377_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_,
    new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_,
    new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_,
    new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_,
    new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_,
    new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_,
    new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_,
    new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2432_,
    new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2438_, new_n2439_,
    new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_,
    new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_,
    new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_,
    new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_,
    new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_,
    new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_,
    new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_,
    new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_,
    new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_,
    new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_,
    new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_,
    new_n2556_, new_n2557_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_,
    new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_,
    new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_,
    new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_,
    new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_,
    new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_,
    new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_,
    new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_,
    new_n2612_, new_n2613_, new_n2615_, new_n2616_, new_n2617_, new_n2618_,
    new_n2619_, new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_,
    new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_,
    new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_,
    new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_,
    new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_,
    new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_,
    new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_,
    new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_,
    new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_,
    new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_,
    new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_,
    new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_,
    new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_,
    new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_,
    new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_,
    new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_,
    new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_,
    new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_,
    new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_,
    new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_,
    new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_,
    new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_,
    new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_,
    new_n2764_, new_n2765_, new_n2766_, new_n2768_, new_n2769_, new_n2770_,
    new_n2771_, new_n2772_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2851_,
    new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_,
    new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_,
    new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_,
    new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_,
    new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_,
    new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_,
    new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_,
    new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_,
    new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_,
    new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2911_, new_n2912_,
    new_n2913_, new_n2914_, new_n2915_, new_n2917_, new_n2918_, new_n2919_,
    new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_,
    new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_,
    new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_,
    new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_,
    new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_,
    new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_,
    new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_,
    new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_,
    new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_,
    new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_,
    new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_,
    new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_,
    new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_,
    new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_,
    new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_,
    new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_,
    new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_,
    new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_,
    new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_,
    new_n3092_, new_n3093_, new_n3094_, new_n3096_, new_n3097_, new_n3098_,
    new_n3099_, new_n3100_, new_n3102_, new_n3103_, new_n3104_, new_n3105_,
    new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_,
    new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_,
    new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_,
    new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_,
    new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_,
    new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_,
    new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_,
    new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3154_,
    new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3214_, new_n3215_, new_n3216_,
    new_n3217_, new_n3218_, new_n3220_, new_n3221_, new_n3222_, new_n3223_,
    new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_,
    new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_,
    new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_,
    new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_,
    new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_,
    new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_,
    new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_,
    new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_,
    new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3326_, new_n3327_, new_n3328_,
    new_n3329_, new_n3330_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_,
    new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_,
    new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_,
    new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_,
    new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_,
    new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_,
    new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_,
    new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_,
    new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3434_,
    new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3440_, new_n3441_,
    new_n3443_, new_n3444_, new_n3446_, new_n3447_, new_n3449_, new_n3450_,
    new_n3452_, new_n3453_, new_n3455_, new_n3456_, new_n3458_, new_n3459_,
    new_n3461_, new_n3462_, new_n3464_, new_n3465_, new_n3467_, new_n3468_,
    new_n3470_, new_n3471_, new_n3473_, new_n3474_, new_n3476_, new_n3477_,
    new_n3479_, new_n3480_, new_n3482_, new_n3483_, new_n3485_, new_n3486_,
    new_n3488_, new_n3489_, new_n3491_, new_n3492_, new_n3494_, new_n3495_,
    new_n3497_, new_n3498_, new_n3500_, new_n3501_, new_n3503_, new_n3504_,
    new_n3506_, new_n3507_, new_n3509_, new_n3510_, new_n3512_, new_n3513_,
    new_n3515_, new_n3516_, new_n3518_, new_n3519_, new_n3521_, new_n3522_,
    new_n3524_, new_n3525_, new_n3527_, new_n3528_, new_n3530_, new_n3531_,
    new_n3533_, new_n3534_, new_n3536_, new_n3537_, new_n3539_, new_n3540_,
    new_n3542_, new_n3543_, new_n3545_, new_n3546_, new_n3548_, new_n3549_,
    new_n3551_, new_n3552_, new_n3554_, new_n3555_, new_n3557_, new_n3558_,
    new_n3560_, new_n3561_, new_n3563_, new_n3564_, new_n3566_, new_n3567_,
    new_n3569_, new_n3570_, new_n3572_, new_n3573_, new_n3575_, new_n3576_,
    new_n3578_, new_n3579_, new_n3581_, new_n3582_, new_n3584_, new_n3585_,
    new_n3587_, new_n3588_, new_n3590_, new_n3591_, new_n3593_, new_n3594_,
    new_n3596_, new_n3597_, new_n3599_, new_n3600_, new_n3602_, new_n3603_,
    new_n3605_, new_n3606_, new_n3608_, new_n3609_, new_n3611_, new_n3612_,
    new_n3614_, new_n3615_, new_n3617_, new_n3618_, new_n3620_, new_n3621_,
    new_n3623_, new_n3624_, new_n3626_, new_n3627_, new_n3629_, new_n3630_,
    new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_,
    new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3644_, new_n3645_,
    new_n3646_, new_n3647_, new_n3649_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_,
    new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_,
    new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_,
    new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_,
    new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_,
    new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3722_,
    new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_,
    new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_,
    new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3740_, new_n3741_,
    new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_,
    new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_,
    new_n3754_, new_n3755_, new_n3757_, new_n3758_, new_n3759_, new_n3760_,
    new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_,
    new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3791_, new_n3792_,
    new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_,
    new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_,
    new_n3805_, new_n3806_, new_n3808_, new_n3809_, new_n3810_, new_n3811_,
    new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_,
    new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_,
    new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_,
    new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_,
    new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3842_, new_n3843_,
    new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_,
    new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_,
    new_n3856_, new_n3857_, new_n3859_, new_n3860_, new_n3861_, new_n3862_,
    new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_,
    new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3893_, new_n3894_,
    new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_,
    new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_,
    new_n3907_, new_n3908_, new_n3910_, new_n3911_, new_n3912_, new_n3913_,
    new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_,
    new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_,
    new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_,
    new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_,
    new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3944_, new_n3945_,
    new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_,
    new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_,
    new_n3958_, new_n3959_, new_n3961_, new_n3962_, new_n3963_, new_n3964_,
    new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_,
    new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3995_, new_n3996_,
    new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_,
    new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_,
    new_n4009_, new_n4010_, new_n4012_, new_n4013_, new_n4014_, new_n4015_,
    new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_,
    new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_,
    new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_,
    new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_,
    new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4046_, new_n4047_,
    new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_,
    new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_,
    new_n4060_, new_n4061_, new_n4063_, new_n4064_, new_n4065_, new_n4066_,
    new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_,
    new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4096_, new_n4097_, new_n4098_,
    new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_,
    new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_,
    new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_, new_n4117_,
    new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_, new_n4123_,
    new_n4124_, new_n4125_, new_n4127_, new_n4128_, new_n4129_, new_n4130_,
    new_n4131_, new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_,
    new_n4137_, new_n4138_, new_n4139_, new_n4140_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_,
    new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_,
    new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4161_, new_n4162_,
    new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_,
    new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_,
    new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4180_, new_n4181_,
    new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_,
    new_n4213_, new_n4214_, new_n4216_, new_n4217_, new_n4218_, new_n4219_,
    new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_, new_n4225_,
    new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_,
    new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_,
    new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_,
    new_n4245_, new_n4246_, new_n4247_, new_n4248_, new_n4250_, new_n4251_,
    new_n4252_, new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_,
    new_n4258_, new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_,
    new_n4264_, new_n4265_, new_n4267_, new_n4268_, new_n4269_, new_n4270_,
    new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_,
    new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4301_, new_n4302_,
    new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_,
    new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_,
    new_n4315_, new_n4316_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_, new_n4340_,
    new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_,
    new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4352_, new_n4353_,
    new_n4354_, new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_,
    new_n4360_, new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_,
    new_n4366_, new_n4367_, new_n4369_, new_n4370_, new_n4371_, new_n4372_,
    new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_,
    new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4403_, new_n4404_,
    new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_,
    new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_,
    new_n4417_, new_n4418_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_, new_n4442_,
    new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_, new_n4448_,
    new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4454_, new_n4455_,
    new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_,
    new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_,
    new_n4468_, new_n4469_, new_n4471_, new_n4472_, new_n4473_, new_n4474_,
    new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_,
    new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4505_, new_n4506_,
    new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_,
    new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_,
    new_n4519_, new_n4520_, new_n4522_, new_n4523_, new_n4524_, new_n4525_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_,
    new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_,
    new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_,
    new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4556_, new_n4557_,
    new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_,
    new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_,
    new_n4570_, new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_,
    new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_,
    new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_,
    new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_,
    new_n4615_, new_n4616_, new_n4618_, new_n4619_, new_n4620_, new_n4621_,
    new_n4622_, new_n4623_;
  assign new_n502_ = \count<1>  & \count<0> ;
  assign new_n503_ = \count<2>  & new_n502_;
  assign new_n504_ = \count<3>  & new_n503_;
  assign new_n505_ = \inreg<47>  & \count<0> ;
  assign new_n506_ = \inreg<55>  & ~\count<0> ;
  assign new_n507_ = ~new_n505_ & ~new_n506_;
  assign \inreg_new<55>  = ~new_n504_ & ~new_n507_;
  assign new_n509_ = \inreg<46>  & \count<0> ;
  assign new_n510_ = \inreg<54>  & ~\count<0> ;
  assign new_n511_ = ~new_n509_ & ~new_n510_;
  assign \inreg_new<54>  = ~new_n504_ & ~new_n511_;
  assign new_n513_ = \inreg<45>  & \count<0> ;
  assign new_n514_ = \inreg<53>  & ~\count<0> ;
  assign new_n515_ = ~new_n513_ & ~new_n514_;
  assign \inreg_new<53>  = ~new_n504_ & ~new_n515_;
  assign new_n517_ = \inreg<44>  & \count<0> ;
  assign new_n518_ = \inreg<52>  & ~\count<0> ;
  assign new_n519_ = ~new_n517_ & ~new_n518_;
  assign \inreg_new<52>  = ~new_n504_ & ~new_n519_;
  assign new_n521_ = \inreg<43>  & \count<0> ;
  assign new_n522_ = \inreg<51>  & ~\count<0> ;
  assign new_n523_ = ~new_n521_ & ~new_n522_;
  assign \inreg_new<51>  = ~new_n504_ & ~new_n523_;
  assign new_n525_ = \inreg<42>  & \count<0> ;
  assign new_n526_ = \inreg<50>  & ~\count<0> ;
  assign new_n527_ = ~new_n525_ & ~new_n526_;
  assign \inreg_new<50>  = ~new_n504_ & ~new_n527_;
  assign new_n529_ = \inreg<41>  & \count<0> ;
  assign new_n530_ = \inreg<49>  & ~\count<0> ;
  assign new_n531_ = ~new_n529_ & ~new_n530_;
  assign \inreg_new<49>  = ~new_n504_ & ~new_n531_;
  assign new_n533_ = \inreg<40>  & \count<0> ;
  assign new_n534_ = \inreg<48>  & ~\count<0> ;
  assign new_n535_ = ~new_n533_ & ~new_n534_;
  assign \inreg_new<48>  = ~new_n504_ & ~new_n535_;
  assign new_n537_ = \inreg<39>  & \count<0> ;
  assign new_n538_ = \inreg<47>  & ~\count<0> ;
  assign new_n539_ = ~new_n537_ & ~new_n538_;
  assign \inreg_new<47>  = ~new_n504_ & ~new_n539_;
  assign new_n541_ = \inreg<38>  & \count<0> ;
  assign new_n542_ = \inreg<46>  & ~\count<0> ;
  assign new_n543_ = ~new_n541_ & ~new_n542_;
  assign \inreg_new<46>  = ~new_n504_ & ~new_n543_;
  assign new_n545_ = \inreg<37>  & \count<0> ;
  assign new_n546_ = \inreg<45>  & ~\count<0> ;
  assign new_n547_ = ~new_n545_ & ~new_n546_;
  assign \inreg_new<45>  = ~new_n504_ & ~new_n547_;
  assign new_n549_ = \inreg<36>  & \count<0> ;
  assign new_n550_ = \inreg<44>  & ~\count<0> ;
  assign new_n551_ = ~new_n549_ & ~new_n550_;
  assign \inreg_new<44>  = ~new_n504_ & ~new_n551_;
  assign new_n553_ = \inreg<35>  & \count<0> ;
  assign new_n554_ = \inreg<43>  & ~\count<0> ;
  assign new_n555_ = ~new_n553_ & ~new_n554_;
  assign \inreg_new<43>  = ~new_n504_ & ~new_n555_;
  assign new_n557_ = \inreg<34>  & \count<0> ;
  assign new_n558_ = \inreg<42>  & ~\count<0> ;
  assign new_n559_ = ~new_n557_ & ~new_n558_;
  assign \inreg_new<42>  = ~new_n504_ & ~new_n559_;
  assign new_n561_ = \inreg<33>  & \count<0> ;
  assign new_n562_ = \inreg<41>  & ~\count<0> ;
  assign new_n563_ = ~new_n561_ & ~new_n562_;
  assign \inreg_new<41>  = ~new_n504_ & ~new_n563_;
  assign new_n565_ = \inreg<32>  & \count<0> ;
  assign new_n566_ = \inreg<40>  & ~\count<0> ;
  assign new_n567_ = ~new_n565_ & ~new_n566_;
  assign \inreg_new<40>  = ~new_n504_ & ~new_n567_;
  assign new_n569_ = \inreg<31>  & \count<0> ;
  assign new_n570_ = \inreg<39>  & ~\count<0> ;
  assign new_n571_ = ~new_n569_ & ~new_n570_;
  assign \inreg_new<39>  = ~new_n504_ & ~new_n571_;
  assign new_n573_ = \inreg<30>  & \count<0> ;
  assign new_n574_ = \inreg<38>  & ~\count<0> ;
  assign new_n575_ = ~new_n573_ & ~new_n574_;
  assign \inreg_new<38>  = ~new_n504_ & ~new_n575_;
  assign new_n577_ = \inreg<29>  & \count<0> ;
  assign new_n578_ = \inreg<37>  & ~\count<0> ;
  assign new_n579_ = ~new_n577_ & ~new_n578_;
  assign \inreg_new<37>  = ~new_n504_ & ~new_n579_;
  assign new_n581_ = \inreg<28>  & \count<0> ;
  assign new_n582_ = \inreg<36>  & ~\count<0> ;
  assign new_n583_ = ~new_n581_ & ~new_n582_;
  assign \inreg_new<36>  = ~new_n504_ & ~new_n583_;
  assign new_n585_ = \inreg<27>  & \count<0> ;
  assign new_n586_ = \inreg<35>  & ~\count<0> ;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign \inreg_new<35>  = ~new_n504_ & ~new_n587_;
  assign new_n589_ = \inreg<26>  & \count<0> ;
  assign new_n590_ = \inreg<34>  & ~\count<0> ;
  assign new_n591_ = ~new_n589_ & ~new_n590_;
  assign \inreg_new<34>  = ~new_n504_ & ~new_n591_;
  assign new_n593_ = \inreg<25>  & \count<0> ;
  assign new_n594_ = \inreg<33>  & ~\count<0> ;
  assign new_n595_ = ~new_n593_ & ~new_n594_;
  assign \inreg_new<33>  = ~new_n504_ & ~new_n595_;
  assign new_n597_ = \inreg<24>  & \count<0> ;
  assign new_n598_ = \inreg<32>  & ~\count<0> ;
  assign new_n599_ = ~new_n597_ & ~new_n598_;
  assign \inreg_new<32>  = ~new_n504_ & ~new_n599_;
  assign new_n601_ = \inreg<23>  & \count<0> ;
  assign new_n602_ = \inreg<31>  & ~\count<0> ;
  assign new_n603_ = ~new_n601_ & ~new_n602_;
  assign \inreg_new<31>  = ~new_n504_ & ~new_n603_;
  assign new_n605_ = \inreg<22>  & \count<0> ;
  assign new_n606_ = \inreg<30>  & ~\count<0> ;
  assign new_n607_ = ~new_n605_ & ~new_n606_;
  assign \inreg_new<30>  = ~new_n504_ & ~new_n607_;
  assign new_n609_ = \inreg<21>  & \count<0> ;
  assign new_n610_ = \inreg<29>  & ~\count<0> ;
  assign new_n611_ = ~new_n609_ & ~new_n610_;
  assign \inreg_new<29>  = ~new_n504_ & ~new_n611_;
  assign new_n613_ = \inreg<20>  & \count<0> ;
  assign new_n614_ = \inreg<28>  & ~\count<0> ;
  assign new_n615_ = ~new_n613_ & ~new_n614_;
  assign \inreg_new<28>  = ~new_n504_ & ~new_n615_;
  assign new_n617_ = \inreg<19>  & \count<0> ;
  assign new_n618_ = \inreg<27>  & ~\count<0> ;
  assign new_n619_ = ~new_n617_ & ~new_n618_;
  assign \inreg_new<27>  = ~new_n504_ & ~new_n619_;
  assign new_n621_ = \inreg<18>  & \count<0> ;
  assign new_n622_ = \inreg<26>  & ~\count<0> ;
  assign new_n623_ = ~new_n621_ & ~new_n622_;
  assign \inreg_new<26>  = ~new_n504_ & ~new_n623_;
  assign new_n625_ = \inreg<17>  & \count<0> ;
  assign new_n626_ = \inreg<25>  & ~\count<0> ;
  assign new_n627_ = ~new_n625_ & ~new_n626_;
  assign \inreg_new<25>  = ~new_n504_ & ~new_n627_;
  assign new_n629_ = \inreg<16>  & \count<0> ;
  assign new_n630_ = \inreg<24>  & ~\count<0> ;
  assign new_n631_ = ~new_n629_ & ~new_n630_;
  assign \inreg_new<24>  = ~new_n504_ & ~new_n631_;
  assign new_n633_ = \inreg<15>  & \count<0> ;
  assign new_n634_ = \inreg<23>  & ~\count<0> ;
  assign new_n635_ = ~new_n633_ & ~new_n634_;
  assign \inreg_new<23>  = ~new_n504_ & ~new_n635_;
  assign new_n637_ = \inreg<14>  & \count<0> ;
  assign new_n638_ = \inreg<22>  & ~\count<0> ;
  assign new_n639_ = ~new_n637_ & ~new_n638_;
  assign \inreg_new<22>  = ~new_n504_ & ~new_n639_;
  assign new_n641_ = \inreg<13>  & \count<0> ;
  assign new_n642_ = \inreg<21>  & ~\count<0> ;
  assign new_n643_ = ~new_n641_ & ~new_n642_;
  assign \inreg_new<21>  = ~new_n504_ & ~new_n643_;
  assign new_n645_ = \inreg<12>  & \count<0> ;
  assign new_n646_ = \inreg<20>  & ~\count<0> ;
  assign new_n647_ = ~new_n645_ & ~new_n646_;
  assign \inreg_new<20>  = ~new_n504_ & ~new_n647_;
  assign new_n649_ = \inreg<11>  & \count<0> ;
  assign new_n650_ = \inreg<19>  & ~\count<0> ;
  assign new_n651_ = ~new_n649_ & ~new_n650_;
  assign \inreg_new<19>  = ~new_n504_ & ~new_n651_;
  assign new_n653_ = \inreg<10>  & \count<0> ;
  assign new_n654_ = \inreg<18>  & ~\count<0> ;
  assign new_n655_ = ~new_n653_ & ~new_n654_;
  assign \inreg_new<18>  = ~new_n504_ & ~new_n655_;
  assign new_n657_ = \inreg<17>  & ~\count<0> ;
  assign new_n658_ = \inreg<9>  & \count<0> ;
  assign new_n659_ = ~new_n657_ & ~new_n658_;
  assign \inreg_new<17>  = ~new_n504_ & ~new_n659_;
  assign new_n661_ = \inreg<16>  & ~\count<0> ;
  assign new_n662_ = \inreg<8>  & \count<0> ;
  assign new_n663_ = ~new_n661_ & ~new_n662_;
  assign \inreg_new<16>  = ~new_n504_ & ~new_n663_;
  assign new_n665_ = \inreg<15>  & ~\count<0> ;
  assign new_n666_ = \inreg<7>  & \count<0> ;
  assign new_n667_ = ~new_n665_ & ~new_n666_;
  assign \inreg_new<15>  = ~new_n504_ & ~new_n667_;
  assign new_n669_ = \inreg<14>  & ~\count<0> ;
  assign new_n670_ = \inreg<6>  & \count<0> ;
  assign new_n671_ = ~new_n669_ & ~new_n670_;
  assign \inreg_new<14>  = ~new_n504_ & ~new_n671_;
  assign new_n673_ = \inreg<13>  & ~\count<0> ;
  assign new_n674_ = \inreg<5>  & \count<0> ;
  assign new_n675_ = ~new_n673_ & ~new_n674_;
  assign \inreg_new<13>  = ~new_n504_ & ~new_n675_;
  assign new_n677_ = \inreg<12>  & ~\count<0> ;
  assign new_n678_ = \inreg<4>  & \count<0> ;
  assign new_n679_ = ~new_n677_ & ~new_n678_;
  assign \inreg_new<12>  = ~new_n504_ & ~new_n679_;
  assign new_n681_ = \inreg<11>  & ~\count<0> ;
  assign new_n682_ = \inreg<3>  & \count<0> ;
  assign new_n683_ = ~new_n681_ & ~new_n682_;
  assign \inreg_new<11>  = ~new_n504_ & ~new_n683_;
  assign new_n685_ = \inreg<10>  & ~\count<0> ;
  assign new_n686_ = \inreg<2>  & \count<0> ;
  assign new_n687_ = ~new_n685_ & ~new_n686_;
  assign \inreg_new<10>  = ~new_n504_ & ~new_n687_;
  assign new_n689_ = \inreg<1>  & \count<0> ;
  assign new_n690_ = \inreg<9>  & ~\count<0> ;
  assign new_n691_ = ~new_n689_ & ~new_n690_;
  assign \inreg_new<9>  = ~new_n504_ & ~new_n691_;
  assign new_n693_ = \inreg<0>  & \count<0> ;
  assign new_n694_ = \inreg<8>  & ~\count<0> ;
  assign new_n695_ = ~new_n693_ & ~new_n694_;
  assign \inreg_new<8>  = ~new_n504_ & ~new_n695_;
  assign new_n697_ = \data_in<7>  & \count<0> ;
  assign new_n698_ = \inreg<7>  & ~\count<0> ;
  assign new_n699_ = ~new_n697_ & ~new_n698_;
  assign \inreg_new<7>  = ~new_n504_ & ~new_n699_;
  assign new_n701_ = \data_in<6>  & \count<0> ;
  assign new_n702_ = \inreg<6>  & ~\count<0> ;
  assign new_n703_ = ~new_n701_ & ~new_n702_;
  assign \inreg_new<6>  = ~new_n504_ & ~new_n703_;
  assign new_n705_ = \data_in<5>  & \count<0> ;
  assign new_n706_ = \inreg<5>  & ~\count<0> ;
  assign new_n707_ = ~new_n705_ & ~new_n706_;
  assign \inreg_new<5>  = ~new_n504_ & ~new_n707_;
  assign new_n709_ = \data_in<4>  & \count<0> ;
  assign new_n710_ = \inreg<4>  & ~\count<0> ;
  assign new_n711_ = ~new_n709_ & ~new_n710_;
  assign \inreg_new<4>  = ~new_n504_ & ~new_n711_;
  assign new_n713_ = \data_in<3>  & \count<0> ;
  assign new_n714_ = \inreg<3>  & ~\count<0> ;
  assign new_n715_ = ~new_n713_ & ~new_n714_;
  assign \inreg_new<3>  = ~new_n504_ & ~new_n715_;
  assign new_n717_ = \data_in<2>  & \count<0> ;
  assign new_n718_ = \inreg<2>  & ~\count<0> ;
  assign new_n719_ = ~new_n717_ & ~new_n718_;
  assign \inreg_new<2>  = ~new_n504_ & ~new_n719_;
  assign new_n721_ = \data_in<1>  & \count<0> ;
  assign new_n722_ = \inreg<1>  & ~\count<0> ;
  assign new_n723_ = ~new_n721_ & ~new_n722_;
  assign \inreg_new<1>  = ~new_n504_ & ~new_n723_;
  assign new_n725_ = \data_in<0>  & \count<0> ;
  assign new_n726_ = \inreg<0>  & ~\count<0> ;
  assign new_n727_ = ~new_n725_ & ~new_n726_;
  assign \inreg_new<0>  = ~new_n504_ & ~new_n727_;
  assign new_n729_ = \data<47>  & ~\D<12> ;
  assign new_n730_ = ~\data<47>  & \D<12> ;
  assign new_n731_ = ~new_n729_ & ~new_n730_;
  assign new_n732_ = \data<48>  & ~\D<23> ;
  assign new_n733_ = ~\data<48>  & \D<23> ;
  assign new_n734_ = ~new_n732_ & ~new_n733_;
  assign new_n735_ = \data<49>  & ~\D<2> ;
  assign new_n736_ = ~\data<49>  & \D<2> ;
  assign new_n737_ = ~new_n735_ & ~new_n736_;
  assign new_n738_ = \data<50>  & ~\D<8> ;
  assign new_n739_ = ~\data<50>  & \D<8> ;
  assign new_n740_ = ~new_n738_ & ~new_n739_;
  assign new_n741_ = \data<51>  & ~\D<18> ;
  assign new_n742_ = ~\data<51>  & \D<18> ;
  assign new_n743_ = ~new_n741_ & ~new_n742_;
  assign new_n744_ = \data<52>  & ~\D<26> ;
  assign new_n745_ = ~\data<52>  & \D<26> ;
  assign new_n746_ = ~new_n744_ & ~new_n745_;
  assign new_n747_ = new_n731_ & new_n734_;
  assign new_n748_ = ~new_n737_ & new_n747_;
  assign new_n749_ = new_n740_ & new_n748_;
  assign new_n750_ = new_n743_ & new_n749_;
  assign new_n751_ = new_n746_ & new_n750_;
  assign new_n752_ = ~new_n743_ & new_n749_;
  assign new_n753_ = new_n746_ & new_n752_;
  assign new_n754_ = ~new_n740_ & new_n748_;
  assign new_n755_ = new_n743_ & new_n754_;
  assign new_n756_ = new_n746_ & new_n755_;
  assign new_n757_ = ~new_n743_ & new_n754_;
  assign new_n758_ = new_n746_ & new_n757_;
  assign new_n759_ = new_n731_ & ~new_n734_;
  assign new_n760_ = new_n737_ & new_n759_;
  assign new_n761_ = ~new_n740_ & new_n760_;
  assign new_n762_ = new_n743_ & new_n761_;
  assign new_n763_ = new_n746_ & new_n762_;
  assign new_n764_ = ~new_n743_ & new_n761_;
  assign new_n765_ = new_n746_ & new_n764_;
  assign new_n766_ = ~new_n737_ & new_n759_;
  assign new_n767_ = ~new_n740_ & new_n766_;
  assign new_n768_ = new_n743_ & new_n767_;
  assign new_n769_ = new_n746_ & new_n768_;
  assign new_n770_ = new_n737_ & new_n747_;
  assign new_n771_ = new_n740_ & new_n770_;
  assign new_n772_ = new_n743_ & new_n771_;
  assign new_n773_ = ~new_n746_ & new_n772_;
  assign new_n774_ = ~new_n743_ & new_n771_;
  assign new_n775_ = ~new_n746_ & new_n774_;
  assign new_n776_ = ~new_n746_ & new_n752_;
  assign new_n777_ = ~new_n746_ & new_n762_;
  assign new_n778_ = ~new_n746_ & new_n764_;
  assign new_n779_ = new_n740_ & new_n766_;
  assign new_n780_ = new_n743_ & new_n779_;
  assign new_n781_ = ~new_n746_ & new_n780_;
  assign new_n782_ = ~new_n743_ & new_n767_;
  assign new_n783_ = ~new_n746_ & new_n782_;
  assign new_n784_ = ~new_n731_ & new_n734_;
  assign new_n785_ = new_n737_ & new_n784_;
  assign new_n786_ = ~new_n740_ & new_n785_;
  assign new_n787_ = ~new_n743_ & new_n786_;
  assign new_n788_ = new_n746_ & new_n787_;
  assign new_n789_ = ~new_n737_ & new_n784_;
  assign new_n790_ = new_n740_ & new_n789_;
  assign new_n791_ = new_n743_ & new_n790_;
  assign new_n792_ = new_n746_ & new_n791_;
  assign new_n793_ = ~new_n740_ & new_n789_;
  assign new_n794_ = new_n743_ & new_n793_;
  assign new_n795_ = new_n746_ & new_n794_;
  assign new_n796_ = ~new_n731_ & ~new_n734_;
  assign new_n797_ = new_n737_ & new_n796_;
  assign new_n798_ = new_n740_ & new_n797_;
  assign new_n799_ = new_n743_ & new_n798_;
  assign new_n800_ = new_n746_ & new_n799_;
  assign new_n801_ = ~new_n737_ & new_n796_;
  assign new_n802_ = new_n740_ & new_n801_;
  assign new_n803_ = new_n743_ & new_n802_;
  assign new_n804_ = new_n746_ & new_n803_;
  assign new_n805_ = ~new_n743_ & new_n802_;
  assign new_n806_ = new_n746_ & new_n805_;
  assign new_n807_ = ~new_n740_ & new_n801_;
  assign new_n808_ = ~new_n743_ & new_n807_;
  assign new_n809_ = new_n746_ & new_n808_;
  assign new_n810_ = new_n740_ & new_n785_;
  assign new_n811_ = new_n743_ & new_n810_;
  assign new_n812_ = ~new_n746_ & new_n811_;
  assign new_n813_ = ~new_n746_ & new_n787_;
  assign new_n814_ = ~new_n743_ & new_n790_;
  assign new_n815_ = ~new_n746_ & new_n814_;
  assign new_n816_ = ~new_n746_ & new_n799_;
  assign new_n817_ = ~new_n743_ & new_n798_;
  assign new_n818_ = ~new_n746_ & new_n817_;
  assign new_n819_ = ~new_n746_ & new_n803_;
  assign new_n820_ = ~new_n746_ & new_n808_;
  assign new_n821_ = ~new_n753_ & ~new_n756_;
  assign new_n822_ = ~new_n751_ & new_n821_;
  assign new_n823_ = ~new_n758_ & ~new_n763_;
  assign new_n824_ = ~new_n765_ & ~new_n769_;
  assign new_n825_ = new_n823_ & new_n824_;
  assign new_n826_ = new_n822_ & new_n825_;
  assign new_n827_ = ~new_n775_ & ~new_n776_;
  assign new_n828_ = ~new_n773_ & new_n827_;
  assign new_n829_ = ~new_n777_ & ~new_n778_;
  assign new_n830_ = ~new_n781_ & ~new_n783_;
  assign new_n831_ = new_n829_ & new_n830_;
  assign new_n832_ = new_n828_ & new_n831_;
  assign new_n833_ = new_n826_ & new_n832_;
  assign new_n834_ = ~new_n792_ & ~new_n795_;
  assign new_n835_ = ~new_n788_ & new_n834_;
  assign new_n836_ = ~new_n800_ & ~new_n804_;
  assign new_n837_ = ~new_n806_ & ~new_n809_;
  assign new_n838_ = new_n836_ & new_n837_;
  assign new_n839_ = new_n835_ & new_n838_;
  assign new_n840_ = ~new_n813_ & ~new_n815_;
  assign new_n841_ = ~new_n812_ & new_n840_;
  assign new_n842_ = ~new_n816_ & ~new_n818_;
  assign new_n843_ = ~new_n819_ & ~new_n820_;
  assign new_n844_ = new_n842_ & new_n843_;
  assign new_n845_ = new_n841_ & new_n844_;
  assign new_n846_ = new_n839_ & new_n845_;
  assign new_n847_ = new_n833_ & new_n846_;
  assign new_n848_ = new_n743_ & ~new_n746_;
  assign new_n849_ = ~new_n737_ & ~new_n740_;
  assign new_n850_ = new_n848_ & new_n849_;
  assign new_n851_ = new_n737_ & new_n740_;
  assign new_n852_ = ~new_n743_ & new_n746_;
  assign new_n853_ = new_n851_ & new_n852_;
  assign new_n854_ = ~new_n850_ & ~new_n853_;
  assign new_n855_ = ~new_n731_ & ~new_n854_;
  assign new_n856_ = ~new_n740_ & ~new_n746_;
  assign new_n857_ = new_n740_ & new_n746_;
  assign new_n858_ = ~new_n856_ & ~new_n857_;
  assign new_n859_ = new_n743_ & ~new_n858_;
  assign new_n860_ = new_n737_ & new_n859_;
  assign new_n861_ = new_n731_ & new_n860_;
  assign new_n862_ = ~new_n855_ & ~new_n861_;
  assign new_n863_ = new_n734_ & ~new_n862_;
  assign new_n864_ = new_n847_ & ~new_n863_;
  assign new_n865_ = ~\data<24>  & ~new_n864_;
  assign new_n866_ = \data<24>  & new_n864_;
  assign new_n867_ = ~new_n865_ & ~new_n866_;
  assign new_n868_ = new_n504_ & ~new_n867_;
  assign new_n869_ = \outreg<63>  & ~\count<0> ;
  assign new_n870_ = ~new_n504_ & new_n869_;
  assign \outreg_new<63>  = new_n868_ | new_n870_;
  assign new_n872_ = \data<56>  & new_n504_;
  assign new_n873_ = \outreg<62>  & ~\count<0> ;
  assign new_n874_ = ~new_n504_ & new_n873_;
  assign \outreg_new<62>  = new_n872_ | new_n874_;
  assign new_n876_ = \data<63>  & ~\C<13> ;
  assign new_n877_ = ~\data<63>  & \C<13> ;
  assign new_n878_ = ~new_n876_ & ~new_n877_;
  assign new_n879_ = \data<32>  & ~\C<16> ;
  assign new_n880_ = ~\data<32>  & \C<16> ;
  assign new_n881_ = ~new_n879_ & ~new_n880_;
  assign new_n882_ = \data<33>  & ~\C<10> ;
  assign new_n883_ = ~\data<33>  & \C<10> ;
  assign new_n884_ = ~new_n882_ & ~new_n883_;
  assign new_n885_ = \data<34>  & ~\C<23> ;
  assign new_n886_ = ~\data<34>  & \C<23> ;
  assign new_n887_ = ~new_n885_ & ~new_n886_;
  assign new_n888_ = \data<35>  & ~\C<0> ;
  assign new_n889_ = ~\data<35>  & \C<0> ;
  assign new_n890_ = ~new_n888_ & ~new_n889_;
  assign new_n891_ = \data<36>  & ~\C<4> ;
  assign new_n892_ = ~\data<36>  & \C<4> ;
  assign new_n893_ = ~new_n891_ & ~new_n892_;
  assign new_n894_ = new_n878_ & new_n881_;
  assign new_n895_ = new_n884_ & new_n894_;
  assign new_n896_ = new_n887_ & new_n895_;
  assign new_n897_ = new_n890_ & new_n896_;
  assign new_n898_ = new_n893_ & new_n897_;
  assign new_n899_ = new_n878_ & ~new_n881_;
  assign new_n900_ = new_n884_ & new_n899_;
  assign new_n901_ = ~new_n887_ & new_n900_;
  assign new_n902_ = new_n890_ & new_n901_;
  assign new_n903_ = new_n893_ & new_n902_;
  assign new_n904_ = ~new_n890_ & new_n901_;
  assign new_n905_ = new_n893_ & new_n904_;
  assign new_n906_ = ~new_n884_ & new_n899_;
  assign new_n907_ = new_n887_ & new_n906_;
  assign new_n908_ = new_n890_ & new_n907_;
  assign new_n909_ = new_n893_ & new_n908_;
  assign new_n910_ = ~new_n887_ & new_n906_;
  assign new_n911_ = ~new_n890_ & new_n910_;
  assign new_n912_ = new_n893_ & new_n911_;
  assign new_n913_ = ~new_n890_ & new_n896_;
  assign new_n914_ = ~new_n893_ & new_n913_;
  assign new_n915_ = ~new_n887_ & new_n895_;
  assign new_n916_ = new_n890_ & new_n915_;
  assign new_n917_ = ~new_n893_ & new_n916_;
  assign new_n918_ = ~new_n884_ & new_n894_;
  assign new_n919_ = new_n887_ & new_n918_;
  assign new_n920_ = new_n890_ & new_n919_;
  assign new_n921_ = ~new_n893_ & new_n920_;
  assign new_n922_ = ~new_n887_ & new_n918_;
  assign new_n923_ = new_n890_ & new_n922_;
  assign new_n924_ = ~new_n893_ & new_n923_;
  assign new_n925_ = new_n887_ & new_n900_;
  assign new_n926_ = ~new_n890_ & new_n925_;
  assign new_n927_ = ~new_n893_ & new_n926_;
  assign new_n928_ = ~new_n893_ & new_n902_;
  assign new_n929_ = ~new_n890_ & new_n907_;
  assign new_n930_ = ~new_n893_ & new_n929_;
  assign new_n931_ = new_n893_ & new_n916_;
  assign new_n932_ = ~new_n878_ & new_n881_;
  assign new_n933_ = new_n884_ & new_n932_;
  assign new_n934_ = ~new_n887_ & new_n933_;
  assign new_n935_ = new_n890_ & new_n934_;
  assign new_n936_ = new_n893_ & new_n935_;
  assign new_n937_ = ~new_n884_ & new_n932_;
  assign new_n938_ = new_n887_ & new_n937_;
  assign new_n939_ = new_n890_ & new_n938_;
  assign new_n940_ = new_n893_ & new_n939_;
  assign new_n941_ = ~new_n890_ & new_n938_;
  assign new_n942_ = new_n893_ & new_n941_;
  assign new_n943_ = ~new_n878_ & ~new_n881_;
  assign new_n944_ = new_n884_ & new_n943_;
  assign new_n945_ = new_n887_ & new_n944_;
  assign new_n946_ = new_n890_ & new_n945_;
  assign new_n947_ = new_n893_ & new_n946_;
  assign new_n948_ = ~new_n890_ & new_n945_;
  assign new_n949_ = new_n893_ & new_n948_;
  assign new_n950_ = ~new_n887_ & new_n944_;
  assign new_n951_ = ~new_n890_ & new_n950_;
  assign new_n952_ = new_n893_ & new_n951_;
  assign new_n953_ = ~new_n884_ & new_n943_;
  assign new_n954_ = ~new_n887_ & new_n953_;
  assign new_n955_ = new_n890_ & new_n954_;
  assign new_n956_ = new_n893_ & new_n955_;
  assign new_n957_ = new_n887_ & new_n933_;
  assign new_n958_ = new_n890_ & new_n957_;
  assign new_n959_ = ~new_n893_ & new_n958_;
  assign new_n960_ = ~new_n890_ & new_n957_;
  assign new_n961_ = ~new_n893_ & new_n960_;
  assign new_n962_ = ~new_n887_ & new_n937_;
  assign new_n963_ = ~new_n890_ & new_n962_;
  assign new_n964_ = ~new_n893_ & new_n963_;
  assign new_n965_ = ~new_n893_ & new_n946_;
  assign new_n966_ = ~new_n893_ & new_n951_;
  assign new_n967_ = ~new_n890_ & new_n919_;
  assign new_n968_ = new_n893_ & new_n967_;
  assign new_n969_ = ~new_n893_ & new_n955_;
  assign new_n970_ = ~new_n890_ & new_n954_;
  assign new_n971_ = ~new_n893_ & new_n970_;
  assign new_n972_ = ~new_n903_ & ~new_n905_;
  assign new_n973_ = ~new_n898_ & new_n972_;
  assign new_n974_ = ~new_n909_ & ~new_n912_;
  assign new_n975_ = ~new_n914_ & ~new_n917_;
  assign new_n976_ = new_n974_ & new_n975_;
  assign new_n977_ = new_n973_ & new_n976_;
  assign new_n978_ = ~new_n924_ & ~new_n927_;
  assign new_n979_ = ~new_n921_ & new_n978_;
  assign new_n980_ = ~new_n928_ & ~new_n930_;
  assign new_n981_ = ~new_n931_ & ~new_n936_;
  assign new_n982_ = new_n980_ & new_n981_;
  assign new_n983_ = new_n979_ & new_n982_;
  assign new_n984_ = new_n977_ & new_n983_;
  assign new_n985_ = ~new_n942_ & ~new_n947_;
  assign new_n986_ = ~new_n940_ & new_n985_;
  assign new_n987_ = ~new_n949_ & ~new_n952_;
  assign new_n988_ = ~new_n956_ & ~new_n959_;
  assign new_n989_ = new_n987_ & new_n988_;
  assign new_n990_ = new_n986_ & new_n989_;
  assign new_n991_ = ~new_n964_ & ~new_n965_;
  assign new_n992_ = ~new_n961_ & new_n991_;
  assign new_n993_ = ~new_n966_ & ~new_n968_;
  assign new_n994_ = ~new_n969_ & ~new_n971_;
  assign new_n995_ = new_n993_ & new_n994_;
  assign new_n996_ = new_n992_ & new_n995_;
  assign new_n997_ = new_n990_ & new_n996_;
  assign new_n998_ = new_n984_ & new_n997_;
  assign new_n999_ = ~new_n884_ & ~new_n893_;
  assign new_n1000_ = new_n884_ & new_n893_;
  assign new_n1001_ = ~new_n999_ & ~new_n1000_;
  assign new_n1002_ = new_n890_ & ~new_n1001_;
  assign new_n1003_ = ~new_n878_ & new_n1002_;
  assign new_n1004_ = ~new_n890_ & new_n893_;
  assign new_n1005_ = new_n878_ & new_n884_;
  assign new_n1006_ = new_n1004_ & new_n1005_;
  assign new_n1007_ = ~new_n1003_ & ~new_n1006_;
  assign new_n1008_ = new_n887_ & ~new_n1007_;
  assign new_n1009_ = ~new_n890_ & ~new_n893_;
  assign new_n1010_ = ~new_n887_ & new_n1009_;
  assign new_n1011_ = new_n1005_ & new_n1010_;
  assign new_n1012_ = ~new_n1008_ & ~new_n1011_;
  assign new_n1013_ = new_n881_ & ~new_n1012_;
  assign new_n1014_ = new_n998_ & ~new_n1013_;
  assign new_n1015_ = ~\data<16>  & ~new_n1014_;
  assign new_n1016_ = \data<16>  & new_n1014_;
  assign new_n1017_ = ~new_n1015_ & ~new_n1016_;
  assign new_n1018_ = new_n504_ & ~new_n1017_;
  assign new_n1019_ = \outreg<61>  & ~\count<0> ;
  assign new_n1020_ = ~new_n504_ & new_n1019_;
  assign \outreg_new<61>  = new_n1018_ | new_n1020_;
  assign new_n1022_ = \data<48>  & new_n504_;
  assign new_n1023_ = \outreg<60>  & ~\count<0> ;
  assign new_n1024_ = ~new_n504_ & new_n1023_;
  assign \outreg_new<60>  = new_n1022_ | new_n1024_;
  assign new_n1026_ = new_n893_ & new_n929_;
  assign new_n1027_ = new_n890_ & new_n925_;
  assign new_n1028_ = ~new_n893_ & new_n1027_;
  assign new_n1029_ = ~new_n893_ & new_n904_;
  assign new_n1030_ = ~new_n893_ & new_n908_;
  assign new_n1031_ = new_n893_ & new_n963_;
  assign new_n1032_ = new_n890_ & new_n950_;
  assign new_n1033_ = new_n893_ & new_n1032_;
  assign new_n1034_ = new_n887_ & new_n953_;
  assign new_n1035_ = ~new_n890_ & new_n1034_;
  assign new_n1036_ = new_n893_ & new_n1035_;
  assign new_n1037_ = ~new_n893_ & new_n941_;
  assign new_n1038_ = ~new_n893_ & new_n948_;
  assign new_n1039_ = new_n890_ & new_n1034_;
  assign new_n1040_ = ~new_n893_ & new_n1039_;
  assign new_n1041_ = new_n893_ & new_n923_;
  assign new_n1042_ = new_n893_ & new_n926_;
  assign new_n1043_ = ~new_n905_ & ~new_n1026_;
  assign new_n1044_ = ~new_n898_ & new_n1043_;
  assign new_n1045_ = ~new_n914_ & ~new_n921_;
  assign new_n1046_ = ~new_n924_ & ~new_n1028_;
  assign new_n1047_ = new_n1045_ & new_n1046_;
  assign new_n1048_ = new_n1044_ & new_n1047_;
  assign new_n1049_ = ~new_n1029_ & ~new_n1030_;
  assign new_n1050_ = ~new_n928_ & new_n1049_;
  assign new_n1051_ = ~new_n940_ & ~new_n1031_;
  assign new_n1052_ = new_n981_ & new_n1051_;
  assign new_n1053_ = new_n1050_ & new_n1052_;
  assign new_n1054_ = new_n1048_ & new_n1053_;
  assign new_n1055_ = ~new_n949_ & ~new_n1033_;
  assign new_n1056_ = ~new_n947_ & new_n1055_;
  assign new_n1057_ = ~new_n959_ & ~new_n1036_;
  assign new_n1058_ = ~new_n961_ & ~new_n1037_;
  assign new_n1059_ = new_n1057_ & new_n1058_;
  assign new_n1060_ = new_n1056_ & new_n1059_;
  assign new_n1061_ = new_n993_ & ~new_n1038_;
  assign new_n1062_ = ~new_n971_ & ~new_n1040_;
  assign new_n1063_ = ~new_n1041_ & ~new_n1042_;
  assign new_n1064_ = new_n1062_ & new_n1063_;
  assign new_n1065_ = new_n1061_ & new_n1064_;
  assign new_n1066_ = new_n1060_ & new_n1065_;
  assign new_n1067_ = new_n1054_ & new_n1066_;
  assign new_n1068_ = new_n890_ & ~new_n893_;
  assign new_n1069_ = ~new_n1004_ & ~new_n1068_;
  assign new_n1070_ = new_n884_ & ~new_n1069_;
  assign new_n1071_ = ~new_n878_ & new_n1070_;
  assign new_n1072_ = new_n878_ & ~new_n884_;
  assign new_n1073_ = new_n1004_ & new_n1072_;
  assign new_n1074_ = ~new_n1071_ & ~new_n1073_;
  assign new_n1075_ = new_n881_ & ~new_n1074_;
  assign new_n1076_ = ~new_n884_ & new_n1009_;
  assign new_n1077_ = new_n899_ & new_n1076_;
  assign new_n1078_ = ~new_n1075_ & ~new_n1077_;
  assign new_n1079_ = ~new_n887_ & ~new_n1078_;
  assign new_n1080_ = new_n1067_ & ~new_n1079_;
  assign new_n1081_ = ~\data<8>  & ~new_n1080_;
  assign new_n1082_ = \data<8>  & new_n1080_;
  assign new_n1083_ = ~new_n1081_ & ~new_n1082_;
  assign new_n1084_ = new_n504_ & ~new_n1083_;
  assign new_n1085_ = \outreg<59>  & ~\count<0> ;
  assign new_n1086_ = ~new_n504_ & new_n1085_;
  assign \outreg_new<59>  = new_n1084_ | new_n1086_;
  assign new_n1088_ = \data<40>  & new_n504_;
  assign new_n1089_ = \outreg<58>  & ~\count<0> ;
  assign new_n1090_ = ~new_n504_ & new_n1089_;
  assign \outreg_new<58>  = new_n1088_ | new_n1090_;
  assign new_n1092_ = \data<43>  & ~\C<15> ;
  assign new_n1093_ = ~\data<43>  & \C<15> ;
  assign new_n1094_ = ~new_n1092_ & ~new_n1093_;
  assign new_n1095_ = \data<44>  & ~\C<6> ;
  assign new_n1096_ = ~\data<44>  & \C<6> ;
  assign new_n1097_ = ~new_n1095_ & ~new_n1096_;
  assign new_n1098_ = \data<45>  & ~\C<26> ;
  assign new_n1099_ = ~\data<45>  & \C<26> ;
  assign new_n1100_ = ~new_n1098_ & ~new_n1099_;
  assign new_n1101_ = \data<46>  & ~\C<19> ;
  assign new_n1102_ = ~\data<46>  & \C<19> ;
  assign new_n1103_ = ~new_n1101_ & ~new_n1102_;
  assign new_n1104_ = \data<47>  & ~\C<12> ;
  assign new_n1105_ = ~\data<47>  & \C<12> ;
  assign new_n1106_ = ~new_n1104_ & ~new_n1105_;
  assign new_n1107_ = \data<48>  & ~\C<1> ;
  assign new_n1108_ = ~\data<48>  & \C<1> ;
  assign new_n1109_ = ~new_n1107_ & ~new_n1108_;
  assign new_n1110_ = new_n1094_ & new_n1097_;
  assign new_n1111_ = new_n1100_ & new_n1110_;
  assign new_n1112_ = new_n1103_ & new_n1111_;
  assign new_n1113_ = new_n1106_ & new_n1112_;
  assign new_n1114_ = new_n1109_ & new_n1113_;
  assign new_n1115_ = ~new_n1106_ & new_n1112_;
  assign new_n1116_ = new_n1109_ & new_n1115_;
  assign new_n1117_ = ~new_n1103_ & new_n1111_;
  assign new_n1118_ = ~new_n1106_ & new_n1117_;
  assign new_n1119_ = new_n1109_ & new_n1118_;
  assign new_n1120_ = ~new_n1100_ & new_n1110_;
  assign new_n1121_ = ~new_n1103_ & new_n1120_;
  assign new_n1122_ = new_n1106_ & new_n1121_;
  assign new_n1123_ = new_n1109_ & new_n1122_;
  assign new_n1124_ = new_n1094_ & ~new_n1097_;
  assign new_n1125_ = new_n1100_ & new_n1124_;
  assign new_n1126_ = ~new_n1103_ & new_n1125_;
  assign new_n1127_ = ~new_n1106_ & new_n1126_;
  assign new_n1128_ = new_n1109_ & new_n1127_;
  assign new_n1129_ = ~new_n1100_ & new_n1124_;
  assign new_n1130_ = new_n1103_ & new_n1129_;
  assign new_n1131_ = new_n1106_ & new_n1130_;
  assign new_n1132_ = new_n1109_ & new_n1131_;
  assign new_n1133_ = ~new_n1103_ & new_n1129_;
  assign new_n1134_ = ~new_n1106_ & new_n1133_;
  assign new_n1135_ = new_n1109_ & new_n1134_;
  assign new_n1136_ = ~new_n1109_ & new_n1113_;
  assign new_n1137_ = new_n1106_ & new_n1117_;
  assign new_n1138_ = ~new_n1109_ & new_n1137_;
  assign new_n1139_ = ~new_n1109_ & new_n1118_;
  assign new_n1140_ = new_n1103_ & new_n1120_;
  assign new_n1141_ = ~new_n1106_ & new_n1140_;
  assign new_n1142_ = ~new_n1109_ & new_n1141_;
  assign new_n1143_ = ~new_n1106_ & new_n1121_;
  assign new_n1144_ = ~new_n1109_ & new_n1143_;
  assign new_n1145_ = new_n1103_ & new_n1125_;
  assign new_n1146_ = ~new_n1106_ & new_n1145_;
  assign new_n1147_ = ~new_n1109_ & new_n1146_;
  assign new_n1148_ = ~new_n1109_ & new_n1134_;
  assign new_n1149_ = ~new_n1094_ & new_n1097_;
  assign new_n1150_ = new_n1100_ & new_n1149_;
  assign new_n1151_ = ~new_n1103_ & new_n1150_;
  assign new_n1152_ = new_n1106_ & new_n1151_;
  assign new_n1153_ = new_n1109_ & new_n1152_;
  assign new_n1154_ = ~new_n1100_ & new_n1149_;
  assign new_n1155_ = new_n1103_ & new_n1154_;
  assign new_n1156_ = ~new_n1106_ & new_n1155_;
  assign new_n1157_ = new_n1109_ & new_n1156_;
  assign new_n1158_ = ~new_n1103_ & new_n1154_;
  assign new_n1159_ = new_n1106_ & new_n1158_;
  assign new_n1160_ = new_n1109_ & new_n1159_;
  assign new_n1161_ = ~new_n1106_ & new_n1158_;
  assign new_n1162_ = new_n1109_ & new_n1161_;
  assign new_n1163_ = ~new_n1094_ & ~new_n1097_;
  assign new_n1164_ = new_n1100_ & new_n1163_;
  assign new_n1165_ = new_n1103_ & new_n1164_;
  assign new_n1166_ = new_n1106_ & new_n1165_;
  assign new_n1167_ = new_n1109_ & new_n1166_;
  assign new_n1168_ = ~new_n1103_ & new_n1164_;
  assign new_n1169_ = new_n1106_ & new_n1168_;
  assign new_n1170_ = new_n1109_ & new_n1169_;
  assign new_n1171_ = ~new_n1100_ & new_n1163_;
  assign new_n1172_ = new_n1103_ & new_n1171_;
  assign new_n1173_ = new_n1106_ & new_n1172_;
  assign new_n1174_ = new_n1109_ & new_n1173_;
  assign new_n1175_ = new_n1103_ & new_n1150_;
  assign new_n1176_ = new_n1106_ & new_n1175_;
  assign new_n1177_ = ~new_n1109_ & new_n1176_;
  assign new_n1178_ = ~new_n1106_ & new_n1175_;
  assign new_n1179_ = ~new_n1109_ & new_n1178_;
  assign new_n1180_ = ~new_n1109_ & new_n1159_;
  assign new_n1181_ = ~new_n1109_ & new_n1166_;
  assign new_n1182_ = ~new_n1109_ & new_n1169_;
  assign new_n1183_ = ~new_n1106_ & new_n1168_;
  assign new_n1184_ = ~new_n1109_ & new_n1183_;
  assign new_n1185_ = ~new_n1106_ & new_n1172_;
  assign new_n1186_ = ~new_n1109_ & new_n1185_;
  assign new_n1187_ = ~new_n1116_ & ~new_n1119_;
  assign new_n1188_ = ~new_n1114_ & new_n1187_;
  assign new_n1189_ = ~new_n1123_ & ~new_n1128_;
  assign new_n1190_ = ~new_n1132_ & ~new_n1135_;
  assign new_n1191_ = new_n1189_ & new_n1190_;
  assign new_n1192_ = new_n1188_ & new_n1191_;
  assign new_n1193_ = ~new_n1138_ & ~new_n1139_;
  assign new_n1194_ = ~new_n1136_ & new_n1193_;
  assign new_n1195_ = ~new_n1142_ & ~new_n1144_;
  assign new_n1196_ = ~new_n1147_ & ~new_n1148_;
  assign new_n1197_ = new_n1195_ & new_n1196_;
  assign new_n1198_ = new_n1194_ & new_n1197_;
  assign new_n1199_ = new_n1192_ & new_n1198_;
  assign new_n1200_ = ~new_n1157_ & ~new_n1160_;
  assign new_n1201_ = ~new_n1153_ & new_n1200_;
  assign new_n1202_ = ~new_n1162_ & ~new_n1167_;
  assign new_n1203_ = ~new_n1170_ & ~new_n1174_;
  assign new_n1204_ = new_n1202_ & new_n1203_;
  assign new_n1205_ = new_n1201_ & new_n1204_;
  assign new_n1206_ = ~new_n1179_ & ~new_n1180_;
  assign new_n1207_ = ~new_n1177_ & new_n1206_;
  assign new_n1208_ = ~new_n1181_ & ~new_n1182_;
  assign new_n1209_ = ~new_n1184_ & ~new_n1186_;
  assign new_n1210_ = new_n1208_ & new_n1209_;
  assign new_n1211_ = new_n1207_ & new_n1210_;
  assign new_n1212_ = new_n1205_ & new_n1211_;
  assign new_n1213_ = new_n1199_ & new_n1212_;
  assign new_n1214_ = ~new_n1100_ & ~new_n1109_;
  assign new_n1215_ = new_n1097_ & new_n1214_;
  assign new_n1216_ = new_n1100_ & new_n1109_;
  assign new_n1217_ = ~new_n1097_ & new_n1216_;
  assign new_n1218_ = ~new_n1215_ & ~new_n1217_;
  assign new_n1219_ = ~new_n1106_ & ~new_n1218_;
  assign new_n1220_ = ~new_n1094_ & new_n1219_;
  assign new_n1221_ = ~new_n1214_ & ~new_n1216_;
  assign new_n1222_ = new_n1106_ & ~new_n1221_;
  assign new_n1223_ = ~new_n1097_ & new_n1222_;
  assign new_n1224_ = new_n1094_ & new_n1223_;
  assign new_n1225_ = ~new_n1220_ & ~new_n1224_;
  assign new_n1226_ = new_n1103_ & ~new_n1225_;
  assign new_n1227_ = new_n1213_ & ~new_n1226_;
  assign new_n1228_ = ~\data<0>  & ~new_n1227_;
  assign new_n1229_ = \data<0>  & new_n1227_;
  assign new_n1230_ = ~new_n1228_ & ~new_n1229_;
  assign new_n1231_ = new_n504_ & ~new_n1230_;
  assign new_n1232_ = \outreg<57>  & ~\count<0> ;
  assign new_n1233_ = ~new_n504_ & new_n1232_;
  assign \outreg_new<57>  = new_n1231_ | new_n1233_;
  assign new_n1235_ = \data<32>  & new_n504_;
  assign new_n1236_ = \outreg<56>  & ~\count<0> ;
  assign new_n1237_ = ~new_n504_ & new_n1236_;
  assign \outreg_new<56>  = new_n1235_ | new_n1237_;
  assign new_n1239_ = new_n1109_ & new_n1137_;
  assign new_n1240_ = new_n1109_ & new_n1143_;
  assign new_n1241_ = ~new_n1106_ & new_n1130_;
  assign new_n1242_ = new_n1109_ & new_n1241_;
  assign new_n1243_ = ~new_n1109_ & new_n1127_;
  assign new_n1244_ = ~new_n1109_ & new_n1241_;
  assign new_n1245_ = new_n1106_ & new_n1133_;
  assign new_n1246_ = ~new_n1109_ & new_n1245_;
  assign new_n1247_ = new_n1109_ & new_n1176_;
  assign new_n1248_ = new_n1106_ & new_n1155_;
  assign new_n1249_ = new_n1109_ & new_n1248_;
  assign new_n1250_ = new_n1109_ & new_n1183_;
  assign new_n1251_ = ~new_n1109_ & new_n1248_;
  assign new_n1252_ = ~new_n1109_ & new_n1173_;
  assign new_n1253_ = ~new_n1103_ & new_n1171_;
  assign new_n1254_ = ~new_n1106_ & new_n1253_;
  assign new_n1255_ = ~new_n1109_ & new_n1254_;
  assign new_n1256_ = ~new_n1106_ & ~new_n1109_;
  assign new_n1257_ = new_n1097_ & new_n1256_;
  assign new_n1258_ = new_n1106_ & new_n1109_;
  assign new_n1259_ = ~new_n1097_ & new_n1258_;
  assign new_n1260_ = ~new_n1257_ & ~new_n1259_;
  assign new_n1261_ = ~new_n1100_ & ~new_n1260_;
  assign new_n1262_ = ~new_n1094_ & new_n1261_;
  assign new_n1263_ = new_n1100_ & new_n1258_;
  assign new_n1264_ = new_n1124_ & new_n1263_;
  assign new_n1265_ = ~new_n1262_ & ~new_n1264_;
  assign new_n1266_ = ~new_n1103_ & ~new_n1265_;
  assign new_n1267_ = ~new_n1123_ & ~new_n1239_;
  assign new_n1268_ = ~new_n1116_ & new_n1267_;
  assign new_n1269_ = ~new_n1132_ & ~new_n1240_;
  assign new_n1270_ = ~new_n1135_ & ~new_n1242_;
  assign new_n1271_ = new_n1269_ & new_n1270_;
  assign new_n1272_ = new_n1268_ & new_n1271_;
  assign new_n1273_ = ~new_n1138_ & ~new_n1142_;
  assign new_n1274_ = ~new_n1136_ & new_n1273_;
  assign new_n1275_ = ~new_n1243_ & ~new_n1244_;
  assign new_n1276_ = ~new_n1148_ & ~new_n1246_;
  assign new_n1277_ = new_n1275_ & new_n1276_;
  assign new_n1278_ = new_n1274_ & new_n1277_;
  assign new_n1279_ = new_n1272_ & new_n1278_;
  assign new_n1280_ = ~new_n1153_ & ~new_n1249_;
  assign new_n1281_ = ~new_n1247_ & new_n1280_;
  assign new_n1282_ = ~new_n1157_ & ~new_n1162_;
  assign new_n1283_ = ~new_n1167_ & ~new_n1250_;
  assign new_n1284_ = new_n1282_ & new_n1283_;
  assign new_n1285_ = new_n1281_ & new_n1284_;
  assign new_n1286_ = ~new_n1179_ & ~new_n1251_;
  assign new_n1287_ = ~new_n1180_ & ~new_n1181_;
  assign new_n1288_ = new_n1286_ & new_n1287_;
  assign new_n1289_ = ~new_n1184_ & ~new_n1252_;
  assign new_n1290_ = new_n1097_ & new_n1100_;
  assign new_n1291_ = new_n1094_ & new_n1290_;
  assign new_n1292_ = new_n1103_ & new_n1256_;
  assign new_n1293_ = new_n1291_ & new_n1292_;
  assign new_n1294_ = ~new_n1255_ & ~new_n1293_;
  assign new_n1295_ = new_n1289_ & new_n1294_;
  assign new_n1296_ = new_n1288_ & new_n1295_;
  assign new_n1297_ = new_n1285_ & new_n1296_;
  assign new_n1298_ = new_n1279_ & new_n1297_;
  assign new_n1299_ = ~new_n1266_ & new_n1298_;
  assign new_n1300_ = ~\data<25>  & ~new_n1299_;
  assign new_n1301_ = \data<25>  & new_n1299_;
  assign new_n1302_ = ~new_n1300_ & ~new_n1301_;
  assign new_n1303_ = new_n504_ & ~new_n1302_;
  assign new_n1304_ = \outreg<55>  & ~\count<0> ;
  assign new_n1305_ = \outreg<63>  & \count<0> ;
  assign new_n1306_ = ~new_n1304_ & ~new_n1305_;
  assign new_n1307_ = ~new_n504_ & ~new_n1306_;
  assign \outreg_new<55>  = new_n1303_ | new_n1307_;
  assign new_n1309_ = \data<57>  & new_n504_;
  assign new_n1310_ = \outreg<54>  & ~\count<0> ;
  assign new_n1311_ = \outreg<62>  & \count<0> ;
  assign new_n1312_ = ~new_n1310_ & ~new_n1311_;
  assign new_n1313_ = ~new_n504_ & ~new_n1312_;
  assign \outreg_new<54>  = new_n1309_ | new_n1313_;
  assign new_n1315_ = \data<39>  & ~\C<20> ;
  assign new_n1316_ = ~\data<39>  & \C<20> ;
  assign new_n1317_ = ~new_n1315_ & ~new_n1316_;
  assign new_n1318_ = \data<40>  & ~\C<9> ;
  assign new_n1319_ = ~\data<40>  & \C<9> ;
  assign new_n1320_ = ~new_n1318_ & ~new_n1319_;
  assign new_n1321_ = \data<35>  & ~\C<2> ;
  assign new_n1322_ = ~\data<35>  & \C<2> ;
  assign new_n1323_ = ~new_n1321_ & ~new_n1322_;
  assign new_n1324_ = \data<36>  & ~\C<27> ;
  assign new_n1325_ = ~\data<36>  & \C<27> ;
  assign new_n1326_ = ~new_n1324_ & ~new_n1325_;
  assign new_n1327_ = \data<37>  & ~\C<14> ;
  assign new_n1328_ = ~\data<37>  & \C<14> ;
  assign new_n1329_ = ~new_n1327_ & ~new_n1328_;
  assign new_n1330_ = \data<38>  & ~\C<5> ;
  assign new_n1331_ = ~\data<38>  & \C<5> ;
  assign new_n1332_ = ~new_n1330_ & ~new_n1331_;
  assign new_n1333_ = ~new_n1317_ & new_n1320_;
  assign new_n1334_ = ~new_n1323_ & new_n1333_;
  assign new_n1335_ = new_n1326_ & new_n1334_;
  assign new_n1336_ = new_n1329_ & new_n1335_;
  assign new_n1337_ = ~new_n1332_ & new_n1336_;
  assign new_n1338_ = new_n1317_ & new_n1320_;
  assign new_n1339_ = ~new_n1323_ & new_n1338_;
  assign new_n1340_ = new_n1326_ & new_n1339_;
  assign new_n1341_ = ~new_n1329_ & new_n1340_;
  assign new_n1342_ = ~new_n1332_ & new_n1341_;
  assign new_n1343_ = ~new_n1326_ & new_n1339_;
  assign new_n1344_ = new_n1329_ & new_n1343_;
  assign new_n1345_ = new_n1332_ & new_n1344_;
  assign new_n1346_ = ~new_n1329_ & new_n1343_;
  assign new_n1347_ = new_n1332_ & new_n1346_;
  assign new_n1348_ = ~new_n1326_ & new_n1334_;
  assign new_n1349_ = ~new_n1329_ & new_n1348_;
  assign new_n1350_ = new_n1332_ & new_n1349_;
  assign new_n1351_ = ~new_n1332_ & new_n1349_;
  assign new_n1352_ = new_n1317_ & ~new_n1320_;
  assign new_n1353_ = ~new_n1323_ & new_n1352_;
  assign new_n1354_ = new_n1326_ & new_n1353_;
  assign new_n1355_ = new_n1329_ & new_n1354_;
  assign new_n1356_ = new_n1332_ & new_n1355_;
  assign new_n1357_ = ~new_n1329_ & new_n1354_;
  assign new_n1358_ = new_n1332_ & new_n1357_;
  assign new_n1359_ = ~new_n1317_ & ~new_n1320_;
  assign new_n1360_ = ~new_n1323_ & new_n1359_;
  assign new_n1361_ = new_n1326_ & new_n1360_;
  assign new_n1362_ = ~new_n1329_ & new_n1361_;
  assign new_n1363_ = new_n1332_ & new_n1362_;
  assign new_n1364_ = ~new_n1326_ & new_n1353_;
  assign new_n1365_ = new_n1329_ & new_n1364_;
  assign new_n1366_ = new_n1332_ & new_n1365_;
  assign new_n1367_ = ~new_n1332_ & new_n1365_;
  assign new_n1368_ = ~new_n1326_ & new_n1360_;
  assign new_n1369_ = ~new_n1329_ & new_n1368_;
  assign new_n1370_ = new_n1332_ & new_n1369_;
  assign new_n1371_ = ~new_n1332_ & new_n1369_;
  assign new_n1372_ = new_n1323_ & new_n1338_;
  assign new_n1373_ = new_n1326_ & new_n1372_;
  assign new_n1374_ = new_n1329_ & new_n1373_;
  assign new_n1375_ = new_n1332_ & new_n1374_;
  assign new_n1376_ = new_n1323_ & new_n1333_;
  assign new_n1377_ = new_n1326_ & new_n1376_;
  assign new_n1378_ = ~new_n1329_ & new_n1377_;
  assign new_n1379_ = new_n1332_ & new_n1378_;
  assign new_n1380_ = ~new_n1329_ & new_n1373_;
  assign new_n1381_ = ~new_n1332_ & new_n1380_;
  assign new_n1382_ = ~new_n1326_ & new_n1372_;
  assign new_n1383_ = new_n1329_ & new_n1382_;
  assign new_n1384_ = new_n1332_ & new_n1383_;
  assign new_n1385_ = ~new_n1326_ & new_n1376_;
  assign new_n1386_ = new_n1329_ & new_n1385_;
  assign new_n1387_ = new_n1332_ & new_n1386_;
  assign new_n1388_ = ~new_n1332_ & new_n1386_;
  assign new_n1389_ = ~new_n1329_ & new_n1382_;
  assign new_n1390_ = ~new_n1332_ & new_n1389_;
  assign new_n1391_ = new_n1323_ & new_n1352_;
  assign new_n1392_ = new_n1326_ & new_n1391_;
  assign new_n1393_ = new_n1329_ & new_n1392_;
  assign new_n1394_ = new_n1332_ & new_n1393_;
  assign new_n1395_ = new_n1323_ & new_n1359_;
  assign new_n1396_ = new_n1326_ & new_n1395_;
  assign new_n1397_ = new_n1329_ & new_n1396_;
  assign new_n1398_ = new_n1332_ & new_n1397_;
  assign new_n1399_ = ~new_n1332_ & new_n1397_;
  assign new_n1400_ = ~new_n1329_ & new_n1392_;
  assign new_n1401_ = new_n1332_ & new_n1400_;
  assign new_n1402_ = ~new_n1326_ & new_n1395_;
  assign new_n1403_ = ~new_n1329_ & new_n1402_;
  assign new_n1404_ = new_n1332_ & new_n1403_;
  assign new_n1405_ = ~new_n1326_ & new_n1391_;
  assign new_n1406_ = ~new_n1329_ & new_n1405_;
  assign new_n1407_ = ~new_n1332_ & new_n1406_;
  assign new_n1408_ = ~new_n1332_ & new_n1403_;
  assign new_n1409_ = new_n1329_ & new_n1340_;
  assign new_n1410_ = ~new_n1332_ & new_n1409_;
  assign new_n1411_ = ~new_n1323_ & ~new_n1332_;
  assign new_n1412_ = ~new_n1320_ & new_n1411_;
  assign new_n1413_ = new_n1323_ & new_n1332_;
  assign new_n1414_ = new_n1320_ & new_n1413_;
  assign new_n1415_ = ~new_n1412_ & ~new_n1414_;
  assign new_n1416_ = new_n1326_ & ~new_n1415_;
  assign new_n1417_ = ~new_n1317_ & new_n1416_;
  assign new_n1418_ = ~new_n1326_ & ~new_n1332_;
  assign new_n1419_ = new_n1323_ & new_n1418_;
  assign new_n1420_ = new_n1352_ & new_n1419_;
  assign new_n1421_ = ~new_n1417_ & ~new_n1420_;
  assign new_n1422_ = new_n1329_ & ~new_n1421_;
  assign new_n1423_ = ~new_n1342_ & ~new_n1345_;
  assign new_n1424_ = ~new_n1337_ & new_n1423_;
  assign new_n1425_ = ~new_n1347_ & ~new_n1350_;
  assign new_n1426_ = ~new_n1351_ & ~new_n1356_;
  assign new_n1427_ = new_n1425_ & new_n1426_;
  assign new_n1428_ = new_n1424_ & new_n1427_;
  assign new_n1429_ = ~new_n1363_ & ~new_n1366_;
  assign new_n1430_ = ~new_n1358_ & new_n1429_;
  assign new_n1431_ = ~new_n1367_ & ~new_n1370_;
  assign new_n1432_ = ~new_n1371_ & ~new_n1375_;
  assign new_n1433_ = new_n1431_ & new_n1432_;
  assign new_n1434_ = new_n1430_ & new_n1433_;
  assign new_n1435_ = new_n1428_ & new_n1434_;
  assign new_n1436_ = ~new_n1381_ & ~new_n1384_;
  assign new_n1437_ = ~new_n1379_ & new_n1436_;
  assign new_n1438_ = ~new_n1387_ & ~new_n1388_;
  assign new_n1439_ = ~new_n1390_ & ~new_n1394_;
  assign new_n1440_ = new_n1438_ & new_n1439_;
  assign new_n1441_ = new_n1437_ & new_n1440_;
  assign new_n1442_ = ~new_n1398_ & ~new_n1399_;
  assign new_n1443_ = ~new_n1401_ & ~new_n1404_;
  assign new_n1444_ = new_n1442_ & new_n1443_;
  assign new_n1445_ = ~new_n1407_ & ~new_n1408_;
  assign new_n1446_ = ~new_n1329_ & ~new_n1332_;
  assign new_n1447_ = new_n1326_ & new_n1446_;
  assign new_n1448_ = new_n1320_ & ~new_n1323_;
  assign new_n1449_ = ~new_n1317_ & new_n1448_;
  assign new_n1450_ = new_n1447_ & new_n1449_;
  assign new_n1451_ = ~new_n1410_ & ~new_n1450_;
  assign new_n1452_ = new_n1445_ & new_n1451_;
  assign new_n1453_ = new_n1444_ & new_n1452_;
  assign new_n1454_ = new_n1441_ & new_n1453_;
  assign new_n1455_ = new_n1435_ & new_n1454_;
  assign new_n1456_ = ~new_n1422_ & new_n1455_;
  assign new_n1457_ = ~\data<17>  & ~new_n1456_;
  assign new_n1458_ = \data<17>  & new_n1456_;
  assign new_n1459_ = ~new_n1457_ & ~new_n1458_;
  assign new_n1460_ = new_n504_ & ~new_n1459_;
  assign new_n1461_ = \outreg<53>  & ~\count<0> ;
  assign new_n1462_ = \outreg<61>  & \count<0> ;
  assign new_n1463_ = ~new_n1461_ & ~new_n1462_;
  assign new_n1464_ = ~new_n504_ & ~new_n1463_;
  assign \outreg_new<53>  = new_n1460_ | new_n1464_;
  assign new_n1466_ = \data<49>  & new_n504_;
  assign new_n1467_ = \outreg<52>  & ~\count<0> ;
  assign new_n1468_ = \outreg<60>  & \count<0> ;
  assign new_n1469_ = ~new_n1467_ & ~new_n1468_;
  assign new_n1470_ = ~new_n504_ & ~new_n1469_;
  assign \outreg_new<52>  = new_n1466_ | new_n1470_;
  assign new_n1472_ = new_n1109_ & new_n1141_;
  assign new_n1473_ = new_n1106_ & new_n1140_;
  assign new_n1474_ = ~new_n1109_ & new_n1473_;
  assign new_n1475_ = new_n1109_ & new_n1178_;
  assign new_n1476_ = ~new_n1106_ & new_n1151_;
  assign new_n1477_ = ~new_n1109_ & new_n1476_;
  assign new_n1478_ = ~new_n1119_ & ~new_n1239_;
  assign new_n1479_ = ~new_n1114_ & new_n1478_;
  assign new_n1480_ = ~new_n1240_ & ~new_n1472_;
  assign new_n1481_ = new_n1190_ & new_n1480_;
  assign new_n1482_ = new_n1479_ & new_n1481_;
  assign new_n1483_ = ~new_n1142_ & ~new_n1474_;
  assign new_n1484_ = ~new_n1138_ & new_n1483_;
  assign new_n1485_ = ~new_n1144_ & ~new_n1147_;
  assign new_n1486_ = ~new_n1244_ & ~new_n1246_;
  assign new_n1487_ = new_n1485_ & new_n1486_;
  assign new_n1488_ = new_n1484_ & new_n1487_;
  assign new_n1489_ = new_n1482_ & new_n1488_;
  assign new_n1490_ = ~new_n1157_ & ~new_n1475_;
  assign new_n1491_ = ~new_n1247_ & new_n1490_;
  assign new_n1492_ = ~new_n1160_ & ~new_n1167_;
  assign new_n1493_ = ~new_n1170_ & ~new_n1250_;
  assign new_n1494_ = new_n1492_ & new_n1493_;
  assign new_n1495_ = new_n1491_ & new_n1494_;
  assign new_n1496_ = ~new_n1179_ & ~new_n1477_;
  assign new_n1497_ = ~new_n1177_ & new_n1496_;
  assign new_n1498_ = ~new_n1184_ & ~new_n1251_;
  assign new_n1499_ = ~new_n1186_ & ~new_n1255_;
  assign new_n1500_ = new_n1498_ & new_n1499_;
  assign new_n1501_ = new_n1497_ & new_n1500_;
  assign new_n1502_ = new_n1495_ & new_n1501_;
  assign new_n1503_ = new_n1489_ & new_n1502_;
  assign new_n1504_ = ~new_n1106_ & new_n1109_;
  assign new_n1505_ = new_n1103_ & new_n1504_;
  assign new_n1506_ = new_n1106_ & ~new_n1109_;
  assign new_n1507_ = ~new_n1103_ & new_n1506_;
  assign new_n1508_ = ~new_n1505_ & ~new_n1507_;
  assign new_n1509_ = new_n1094_ & new_n1100_;
  assign new_n1510_ = ~new_n1094_ & ~new_n1100_;
  assign new_n1511_ = ~new_n1509_ & ~new_n1510_;
  assign new_n1512_ = ~new_n1508_ & ~new_n1511_;
  assign new_n1513_ = ~new_n1097_ & new_n1512_;
  assign new_n1514_ = new_n1503_ & ~new_n1513_;
  assign new_n1515_ = ~\data<9>  & ~new_n1514_;
  assign new_n1516_ = \data<9>  & new_n1514_;
  assign new_n1517_ = ~new_n1515_ & ~new_n1516_;
  assign new_n1518_ = new_n504_ & ~new_n1517_;
  assign new_n1519_ = \outreg<51>  & ~\count<0> ;
  assign new_n1520_ = \outreg<59>  & \count<0> ;
  assign new_n1521_ = ~new_n1519_ & ~new_n1520_;
  assign new_n1522_ = ~new_n504_ & ~new_n1521_;
  assign \outreg_new<51>  = new_n1518_ | new_n1522_;
  assign new_n1524_ = \data<41>  & new_n504_;
  assign new_n1525_ = \outreg<50>  & ~\count<0> ;
  assign new_n1526_ = \outreg<58>  & \count<0> ;
  assign new_n1527_ = ~new_n1525_ & ~new_n1526_;
  assign new_n1528_ = ~new_n504_ & ~new_n1527_;
  assign \outreg_new<50>  = new_n1524_ | new_n1528_;
  assign new_n1530_ = new_n1332_ & new_n1341_;
  assign new_n1531_ = new_n1329_ & new_n1348_;
  assign new_n1532_ = ~new_n1332_ & new_n1531_;
  assign new_n1533_ = ~new_n1332_ & new_n1355_;
  assign new_n1534_ = new_n1329_ & new_n1368_;
  assign new_n1535_ = new_n1332_ & new_n1534_;
  assign new_n1536_ = ~new_n1329_ & new_n1364_;
  assign new_n1537_ = ~new_n1332_ & new_n1536_;
  assign new_n1538_ = new_n1329_ & new_n1377_;
  assign new_n1539_ = ~new_n1332_ & new_n1538_;
  assign new_n1540_ = new_n1332_ & new_n1380_;
  assign new_n1541_ = ~new_n1329_ & new_n1385_;
  assign new_n1542_ = ~new_n1332_ & new_n1541_;
  assign new_n1543_ = ~new_n1329_ & new_n1396_;
  assign new_n1544_ = ~new_n1332_ & new_n1543_;
  assign new_n1545_ = new_n1329_ & new_n1402_;
  assign new_n1546_ = ~new_n1332_ & new_n1545_;
  assign new_n1547_ = new_n1332_ & new_n1406_;
  assign new_n1548_ = new_n1332_ & new_n1336_;
  assign new_n1549_ = ~new_n1411_ & ~new_n1413_;
  assign new_n1550_ = new_n1326_ & ~new_n1549_;
  assign new_n1551_ = ~new_n1320_ & new_n1550_;
  assign new_n1552_ = ~new_n1317_ & new_n1551_;
  assign new_n1553_ = ~new_n1323_ & new_n1418_;
  assign new_n1554_ = new_n1338_ & new_n1553_;
  assign new_n1555_ = ~new_n1552_ & ~new_n1554_;
  assign new_n1556_ = ~new_n1329_ & ~new_n1555_;
  assign new_n1557_ = ~new_n1530_ & ~new_n1532_;
  assign new_n1558_ = ~new_n1337_ & new_n1557_;
  assign new_n1559_ = ~new_n1350_ & ~new_n1351_;
  assign new_n1560_ = ~new_n1358_ & ~new_n1533_;
  assign new_n1561_ = new_n1559_ & new_n1560_;
  assign new_n1562_ = new_n1558_ & new_n1561_;
  assign new_n1563_ = ~new_n1366_ & ~new_n1535_;
  assign new_n1564_ = ~new_n1363_ & new_n1563_;
  assign new_n1565_ = ~new_n1367_ & ~new_n1537_;
  assign new_n1566_ = ~new_n1375_ & ~new_n1539_;
  assign new_n1567_ = new_n1565_ & new_n1566_;
  assign new_n1568_ = new_n1564_ & new_n1567_;
  assign new_n1569_ = new_n1562_ & new_n1568_;
  assign new_n1570_ = ~new_n1379_ & ~new_n1381_;
  assign new_n1571_ = ~new_n1540_ & new_n1570_;
  assign new_n1572_ = ~new_n1387_ & ~new_n1542_;
  assign new_n1573_ = ~new_n1394_ & ~new_n1399_;
  assign new_n1574_ = new_n1572_ & new_n1573_;
  assign new_n1575_ = new_n1571_ & new_n1574_;
  assign new_n1576_ = ~new_n1401_ & ~new_n1544_;
  assign new_n1577_ = ~new_n1546_ & ~new_n1547_;
  assign new_n1578_ = new_n1576_ & new_n1577_;
  assign new_n1579_ = ~new_n1407_ & ~new_n1548_;
  assign new_n1580_ = new_n1320_ & new_n1323_;
  assign new_n1581_ = new_n1317_ & new_n1580_;
  assign new_n1582_ = new_n1329_ & ~new_n1332_;
  assign new_n1583_ = ~new_n1326_ & new_n1582_;
  assign new_n1584_ = new_n1581_ & new_n1583_;
  assign new_n1585_ = ~new_n1410_ & ~new_n1584_;
  assign new_n1586_ = new_n1579_ & new_n1585_;
  assign new_n1587_ = new_n1578_ & new_n1586_;
  assign new_n1588_ = new_n1575_ & new_n1587_;
  assign new_n1589_ = new_n1569_ & new_n1588_;
  assign new_n1590_ = ~new_n1556_ & new_n1589_;
  assign new_n1591_ = ~\data<1>  & ~new_n1590_;
  assign new_n1592_ = \data<1>  & new_n1590_;
  assign new_n1593_ = ~new_n1591_ & ~new_n1592_;
  assign new_n1594_ = new_n504_ & ~new_n1593_;
  assign new_n1595_ = \outreg<49>  & ~\count<0> ;
  assign new_n1596_ = \outreg<57>  & \count<0> ;
  assign new_n1597_ = ~new_n1595_ & ~new_n1596_;
  assign new_n1598_ = ~new_n504_ & ~new_n1597_;
  assign \outreg_new<49>  = new_n1594_ | new_n1598_;
  assign new_n1600_ = \data<33>  & new_n504_;
  assign new_n1601_ = \outreg<48>  & ~\count<0> ;
  assign new_n1602_ = \outreg<56>  & \count<0> ;
  assign new_n1603_ = ~new_n1601_ & ~new_n1602_;
  assign new_n1604_ = ~new_n504_ & ~new_n1603_;
  assign \outreg_new<48>  = new_n1600_ | new_n1604_;
  assign new_n1606_ = \data<59>  & ~\D<17> ;
  assign new_n1607_ = ~\data<59>  & \D<17> ;
  assign new_n1608_ = ~new_n1606_ & ~new_n1607_;
  assign new_n1609_ = \data<60>  & ~\D<13> ;
  assign new_n1610_ = ~\data<60>  & \D<13> ;
  assign new_n1611_ = ~new_n1609_ & ~new_n1610_;
  assign new_n1612_ = \data<61>  & ~\D<21> ;
  assign new_n1613_ = ~\data<61>  & \D<21> ;
  assign new_n1614_ = ~new_n1612_ & ~new_n1613_;
  assign new_n1615_ = \data<62>  & ~\D<7> ;
  assign new_n1616_ = ~\data<62>  & \D<7> ;
  assign new_n1617_ = ~new_n1615_ & ~new_n1616_;
  assign new_n1618_ = \data<63>  & ~\D<0> ;
  assign new_n1619_ = ~\data<63>  & \D<0> ;
  assign new_n1620_ = ~new_n1618_ & ~new_n1619_;
  assign new_n1621_ = \data<32>  & ~\D<3> ;
  assign new_n1622_ = ~\data<32>  & \D<3> ;
  assign new_n1623_ = ~new_n1621_ & ~new_n1622_;
  assign new_n1624_ = new_n1608_ & new_n1611_;
  assign new_n1625_ = new_n1614_ & new_n1624_;
  assign new_n1626_ = new_n1617_ & new_n1625_;
  assign new_n1627_ = new_n1620_ & new_n1626_;
  assign new_n1628_ = new_n1623_ & new_n1627_;
  assign new_n1629_ = ~new_n1614_ & new_n1624_;
  assign new_n1630_ = new_n1617_ & new_n1629_;
  assign new_n1631_ = new_n1620_ & new_n1630_;
  assign new_n1632_ = new_n1623_ & new_n1631_;
  assign new_n1633_ = ~new_n1620_ & new_n1630_;
  assign new_n1634_ = new_n1623_ & new_n1633_;
  assign new_n1635_ = new_n1608_ & ~new_n1611_;
  assign new_n1636_ = new_n1614_ & new_n1635_;
  assign new_n1637_ = ~new_n1617_ & new_n1636_;
  assign new_n1638_ = ~new_n1620_ & new_n1637_;
  assign new_n1639_ = new_n1623_ & new_n1638_;
  assign new_n1640_ = ~new_n1614_ & new_n1635_;
  assign new_n1641_ = new_n1617_ & new_n1640_;
  assign new_n1642_ = new_n1620_ & new_n1641_;
  assign new_n1643_ = new_n1623_ & new_n1642_;
  assign new_n1644_ = ~new_n1617_ & new_n1640_;
  assign new_n1645_ = new_n1620_ & new_n1644_;
  assign new_n1646_ = new_n1623_ & new_n1645_;
  assign new_n1647_ = ~new_n1620_ & new_n1644_;
  assign new_n1648_ = new_n1623_ & new_n1647_;
  assign new_n1649_ = ~new_n1620_ & new_n1626_;
  assign new_n1650_ = ~new_n1623_ & new_n1649_;
  assign new_n1651_ = ~new_n1617_ & new_n1625_;
  assign new_n1652_ = new_n1620_ & new_n1651_;
  assign new_n1653_ = ~new_n1623_ & new_n1652_;
  assign new_n1654_ = ~new_n1617_ & new_n1629_;
  assign new_n1655_ = new_n1620_ & new_n1654_;
  assign new_n1656_ = ~new_n1623_ & new_n1655_;
  assign new_n1657_ = new_n1617_ & new_n1636_;
  assign new_n1658_ = new_n1620_ & new_n1657_;
  assign new_n1659_ = ~new_n1623_ & new_n1658_;
  assign new_n1660_ = ~new_n1620_ & new_n1657_;
  assign new_n1661_ = ~new_n1623_ & new_n1660_;
  assign new_n1662_ = new_n1620_ & new_n1637_;
  assign new_n1663_ = ~new_n1623_ & new_n1662_;
  assign new_n1664_ = ~new_n1620_ & new_n1641_;
  assign new_n1665_ = ~new_n1623_ & new_n1664_;
  assign new_n1666_ = ~new_n1608_ & new_n1611_;
  assign new_n1667_ = new_n1614_ & new_n1666_;
  assign new_n1668_ = new_n1617_ & new_n1667_;
  assign new_n1669_ = new_n1620_ & new_n1668_;
  assign new_n1670_ = new_n1623_ & new_n1669_;
  assign new_n1671_ = ~new_n1614_ & new_n1666_;
  assign new_n1672_ = new_n1617_ & new_n1671_;
  assign new_n1673_ = ~new_n1620_ & new_n1672_;
  assign new_n1674_ = new_n1623_ & new_n1673_;
  assign new_n1675_ = ~new_n1617_ & new_n1671_;
  assign new_n1676_ = new_n1620_ & new_n1675_;
  assign new_n1677_ = new_n1623_ & new_n1676_;
  assign new_n1678_ = ~new_n1608_ & ~new_n1611_;
  assign new_n1679_ = new_n1614_ & new_n1678_;
  assign new_n1680_ = new_n1617_ & new_n1679_;
  assign new_n1681_ = ~new_n1620_ & new_n1680_;
  assign new_n1682_ = new_n1623_ & new_n1681_;
  assign new_n1683_ = ~new_n1617_ & new_n1679_;
  assign new_n1684_ = ~new_n1620_ & new_n1683_;
  assign new_n1685_ = new_n1623_ & new_n1684_;
  assign new_n1686_ = ~new_n1614_ & new_n1678_;
  assign new_n1687_ = new_n1617_ & new_n1686_;
  assign new_n1688_ = new_n1620_ & new_n1687_;
  assign new_n1689_ = new_n1623_ & new_n1688_;
  assign new_n1690_ = ~new_n1617_ & new_n1686_;
  assign new_n1691_ = new_n1620_ & new_n1690_;
  assign new_n1692_ = new_n1623_ & new_n1691_;
  assign new_n1693_ = ~new_n1617_ & new_n1667_;
  assign new_n1694_ = new_n1620_ & new_n1693_;
  assign new_n1695_ = ~new_n1623_ & new_n1694_;
  assign new_n1696_ = ~new_n1620_ & new_n1693_;
  assign new_n1697_ = ~new_n1623_ & new_n1696_;
  assign new_n1698_ = ~new_n1620_ & new_n1675_;
  assign new_n1699_ = ~new_n1623_ & new_n1698_;
  assign new_n1700_ = new_n1620_ & new_n1680_;
  assign new_n1701_ = ~new_n1623_ & new_n1700_;
  assign new_n1702_ = ~new_n1623_ & new_n1681_;
  assign new_n1703_ = ~new_n1620_ & new_n1687_;
  assign new_n1704_ = ~new_n1623_ & new_n1703_;
  assign new_n1705_ = ~new_n1623_ & new_n1691_;
  assign new_n1706_ = new_n1617_ & ~new_n1623_;
  assign new_n1707_ = ~new_n1614_ & new_n1706_;
  assign new_n1708_ = ~new_n1617_ & new_n1623_;
  assign new_n1709_ = new_n1614_ & new_n1708_;
  assign new_n1710_ = ~new_n1707_ & ~new_n1709_;
  assign new_n1711_ = new_n1620_ & ~new_n1710_;
  assign new_n1712_ = ~new_n1608_ & new_n1711_;
  assign new_n1713_ = ~new_n1614_ & ~new_n1623_;
  assign new_n1714_ = new_n1614_ & new_n1623_;
  assign new_n1715_ = ~new_n1713_ & ~new_n1714_;
  assign new_n1716_ = ~new_n1620_ & ~new_n1715_;
  assign new_n1717_ = ~new_n1617_ & new_n1716_;
  assign new_n1718_ = new_n1608_ & new_n1717_;
  assign new_n1719_ = ~new_n1712_ & ~new_n1718_;
  assign new_n1720_ = new_n1611_ & ~new_n1719_;
  assign new_n1721_ = ~new_n1632_ & ~new_n1634_;
  assign new_n1722_ = ~new_n1628_ & new_n1721_;
  assign new_n1723_ = ~new_n1639_ & ~new_n1643_;
  assign new_n1724_ = ~new_n1646_ & ~new_n1648_;
  assign new_n1725_ = new_n1723_ & new_n1724_;
  assign new_n1726_ = new_n1722_ & new_n1725_;
  assign new_n1727_ = ~new_n1653_ & ~new_n1656_;
  assign new_n1728_ = ~new_n1650_ & new_n1727_;
  assign new_n1729_ = ~new_n1659_ & ~new_n1661_;
  assign new_n1730_ = ~new_n1663_ & ~new_n1665_;
  assign new_n1731_ = new_n1729_ & new_n1730_;
  assign new_n1732_ = new_n1728_ & new_n1731_;
  assign new_n1733_ = new_n1726_ & new_n1732_;
  assign new_n1734_ = ~new_n1674_ & ~new_n1677_;
  assign new_n1735_ = ~new_n1670_ & new_n1734_;
  assign new_n1736_ = ~new_n1682_ & ~new_n1685_;
  assign new_n1737_ = ~new_n1689_ & ~new_n1692_;
  assign new_n1738_ = new_n1736_ & new_n1737_;
  assign new_n1739_ = new_n1735_ & new_n1738_;
  assign new_n1740_ = ~new_n1697_ & ~new_n1699_;
  assign new_n1741_ = ~new_n1695_ & new_n1740_;
  assign new_n1742_ = ~new_n1701_ & ~new_n1702_;
  assign new_n1743_ = ~new_n1704_ & ~new_n1705_;
  assign new_n1744_ = new_n1742_ & new_n1743_;
  assign new_n1745_ = new_n1741_ & new_n1744_;
  assign new_n1746_ = new_n1739_ & new_n1745_;
  assign new_n1747_ = new_n1733_ & new_n1746_;
  assign new_n1748_ = ~new_n1720_ & new_n1747_;
  assign new_n1749_ = ~\data<26>  & ~new_n1748_;
  assign new_n1750_ = \data<26>  & new_n1748_;
  assign new_n1751_ = ~new_n1749_ & ~new_n1750_;
  assign new_n1752_ = new_n504_ & ~new_n1751_;
  assign new_n1753_ = \outreg<47>  & ~\count<0> ;
  assign new_n1754_ = \outreg<55>  & \count<0> ;
  assign new_n1755_ = ~new_n1753_ & ~new_n1754_;
  assign new_n1756_ = ~new_n504_ & ~new_n1755_;
  assign \outreg_new<47>  = new_n1752_ | new_n1756_;
  assign new_n1758_ = \data<58>  & new_n504_;
  assign new_n1759_ = \outreg<46>  & ~\count<0> ;
  assign new_n1760_ = \outreg<54>  & \count<0> ;
  assign new_n1761_ = ~new_n1759_ & ~new_n1760_;
  assign new_n1762_ = ~new_n504_ & ~new_n1761_;
  assign \outreg_new<46>  = new_n1758_ | new_n1762_;
  assign new_n1764_ = \data<51>  & ~\D<1> ;
  assign new_n1765_ = ~\data<51>  & \D<1> ;
  assign new_n1766_ = ~new_n1764_ & ~new_n1765_;
  assign new_n1767_ = \data<52>  & ~\D<11> ;
  assign new_n1768_ = ~\data<52>  & \D<11> ;
  assign new_n1769_ = ~new_n1767_ & ~new_n1768_;
  assign new_n1770_ = \data<53>  & ~\D<22> ;
  assign new_n1771_ = ~\data<53>  & \D<22> ;
  assign new_n1772_ = ~new_n1770_ & ~new_n1771_;
  assign new_n1773_ = \data<54>  & ~\D<16> ;
  assign new_n1774_ = ~\data<54>  & \D<16> ;
  assign new_n1775_ = ~new_n1773_ & ~new_n1774_;
  assign new_n1776_ = \data<55>  & ~\D<4> ;
  assign new_n1777_ = ~\data<55>  & \D<4> ;
  assign new_n1778_ = ~new_n1776_ & ~new_n1777_;
  assign new_n1779_ = \data<56>  & ~\D<19> ;
  assign new_n1780_ = ~\data<56>  & \D<19> ;
  assign new_n1781_ = ~new_n1779_ & ~new_n1780_;
  assign new_n1782_ = new_n1766_ & new_n1769_;
  assign new_n1783_ = new_n1772_ & new_n1782_;
  assign new_n1784_ = ~new_n1775_ & new_n1783_;
  assign new_n1785_ = ~new_n1778_ & new_n1784_;
  assign new_n1786_ = new_n1781_ & new_n1785_;
  assign new_n1787_ = ~new_n1772_ & new_n1782_;
  assign new_n1788_ = new_n1775_ & new_n1787_;
  assign new_n1789_ = new_n1778_ & new_n1788_;
  assign new_n1790_ = new_n1781_ & new_n1789_;
  assign new_n1791_ = new_n1766_ & ~new_n1769_;
  assign new_n1792_ = new_n1772_ & new_n1791_;
  assign new_n1793_ = new_n1775_ & new_n1792_;
  assign new_n1794_ = ~new_n1778_ & new_n1793_;
  assign new_n1795_ = new_n1781_ & new_n1794_;
  assign new_n1796_ = ~new_n1775_ & new_n1792_;
  assign new_n1797_ = new_n1778_ & new_n1796_;
  assign new_n1798_ = new_n1781_ & new_n1797_;
  assign new_n1799_ = ~new_n1772_ & new_n1791_;
  assign new_n1800_ = new_n1775_ & new_n1799_;
  assign new_n1801_ = ~new_n1778_ & new_n1800_;
  assign new_n1802_ = new_n1781_ & new_n1801_;
  assign new_n1803_ = ~new_n1775_ & new_n1799_;
  assign new_n1804_ = new_n1778_ & new_n1803_;
  assign new_n1805_ = new_n1781_ & new_n1804_;
  assign new_n1806_ = ~new_n1778_ & new_n1803_;
  assign new_n1807_ = new_n1781_ & new_n1806_;
  assign new_n1808_ = new_n1775_ & new_n1783_;
  assign new_n1809_ = ~new_n1778_ & new_n1808_;
  assign new_n1810_ = ~new_n1781_ & new_n1809_;
  assign new_n1811_ = ~new_n1781_ & new_n1789_;
  assign new_n1812_ = ~new_n1775_ & new_n1787_;
  assign new_n1813_ = new_n1778_ & new_n1812_;
  assign new_n1814_ = ~new_n1781_ & new_n1813_;
  assign new_n1815_ = ~new_n1778_ & new_n1812_;
  assign new_n1816_ = ~new_n1781_ & new_n1815_;
  assign new_n1817_ = ~new_n1781_ & new_n1797_;
  assign new_n1818_ = ~new_n1781_ & new_n1801_;
  assign new_n1819_ = ~new_n1781_ & new_n1804_;
  assign new_n1820_ = ~new_n1766_ & new_n1769_;
  assign new_n1821_ = new_n1772_ & new_n1820_;
  assign new_n1822_ = new_n1775_ & new_n1821_;
  assign new_n1823_ = new_n1778_ & new_n1822_;
  assign new_n1824_ = new_n1781_ & new_n1823_;
  assign new_n1825_ = ~new_n1775_ & new_n1821_;
  assign new_n1826_ = new_n1778_ & new_n1825_;
  assign new_n1827_ = new_n1781_ & new_n1826_;
  assign new_n1828_ = ~new_n1778_ & new_n1825_;
  assign new_n1829_ = new_n1781_ & new_n1828_;
  assign new_n1830_ = ~new_n1772_ & new_n1820_;
  assign new_n1831_ = ~new_n1775_ & new_n1830_;
  assign new_n1832_ = ~new_n1778_ & new_n1831_;
  assign new_n1833_ = new_n1781_ & new_n1832_;
  assign new_n1834_ = ~new_n1766_ & ~new_n1769_;
  assign new_n1835_ = new_n1772_ & new_n1834_;
  assign new_n1836_ = new_n1775_ & new_n1835_;
  assign new_n1837_ = new_n1778_ & new_n1836_;
  assign new_n1838_ = new_n1781_ & new_n1837_;
  assign new_n1839_ = ~new_n1772_ & new_n1834_;
  assign new_n1840_ = new_n1775_ & new_n1839_;
  assign new_n1841_ = ~new_n1778_ & new_n1840_;
  assign new_n1842_ = new_n1781_ & new_n1841_;
  assign new_n1843_ = ~new_n1775_ & new_n1839_;
  assign new_n1844_ = new_n1778_ & new_n1843_;
  assign new_n1845_ = new_n1781_ & new_n1844_;
  assign new_n1846_ = ~new_n1778_ & new_n1822_;
  assign new_n1847_ = ~new_n1781_ & new_n1846_;
  assign new_n1848_ = new_n1775_ & new_n1830_;
  assign new_n1849_ = new_n1778_ & new_n1848_;
  assign new_n1850_ = ~new_n1781_ & new_n1849_;
  assign new_n1851_ = ~new_n1778_ & new_n1848_;
  assign new_n1852_ = ~new_n1781_ & new_n1851_;
  assign new_n1853_ = new_n1778_ & new_n1831_;
  assign new_n1854_ = ~new_n1781_ & new_n1853_;
  assign new_n1855_ = ~new_n1781_ & new_n1837_;
  assign new_n1856_ = ~new_n1775_ & new_n1835_;
  assign new_n1857_ = ~new_n1778_ & new_n1856_;
  assign new_n1858_ = ~new_n1781_ & new_n1857_;
  assign new_n1859_ = ~new_n1778_ & new_n1843_;
  assign new_n1860_ = ~new_n1781_ & new_n1859_;
  assign new_n1861_ = ~new_n1775_ & ~new_n1781_;
  assign new_n1862_ = new_n1772_ & new_n1861_;
  assign new_n1863_ = new_n1775_ & new_n1781_;
  assign new_n1864_ = ~new_n1772_ & new_n1863_;
  assign new_n1865_ = ~new_n1862_ & ~new_n1864_;
  assign new_n1866_ = new_n1778_ & ~new_n1865_;
  assign new_n1867_ = ~new_n1766_ & new_n1866_;
  assign new_n1868_ = new_n1766_ & new_n1772_;
  assign new_n1869_ = ~new_n1778_ & ~new_n1781_;
  assign new_n1870_ = new_n1775_ & new_n1869_;
  assign new_n1871_ = new_n1868_ & new_n1870_;
  assign new_n1872_ = ~new_n1867_ & ~new_n1871_;
  assign new_n1873_ = ~new_n1769_ & ~new_n1872_;
  assign new_n1874_ = ~new_n1790_ & ~new_n1795_;
  assign new_n1875_ = ~new_n1786_ & new_n1874_;
  assign new_n1876_ = ~new_n1798_ & ~new_n1802_;
  assign new_n1877_ = ~new_n1805_ & ~new_n1807_;
  assign new_n1878_ = new_n1876_ & new_n1877_;
  assign new_n1879_ = new_n1875_ & new_n1878_;
  assign new_n1880_ = ~new_n1811_ & ~new_n1814_;
  assign new_n1881_ = ~new_n1810_ & new_n1880_;
  assign new_n1882_ = ~new_n1816_ & ~new_n1817_;
  assign new_n1883_ = ~new_n1818_ & ~new_n1819_;
  assign new_n1884_ = new_n1882_ & new_n1883_;
  assign new_n1885_ = new_n1881_ & new_n1884_;
  assign new_n1886_ = new_n1879_ & new_n1885_;
  assign new_n1887_ = ~new_n1827_ & ~new_n1829_;
  assign new_n1888_ = ~new_n1824_ & new_n1887_;
  assign new_n1889_ = ~new_n1833_ & ~new_n1838_;
  assign new_n1890_ = ~new_n1842_ & ~new_n1845_;
  assign new_n1891_ = new_n1889_ & new_n1890_;
  assign new_n1892_ = new_n1888_ & new_n1891_;
  assign new_n1893_ = ~new_n1847_ & ~new_n1850_;
  assign new_n1894_ = ~new_n1852_ & ~new_n1854_;
  assign new_n1895_ = new_n1893_ & new_n1894_;
  assign new_n1896_ = ~new_n1855_ & ~new_n1858_;
  assign new_n1897_ = ~new_n1778_ & new_n1781_;
  assign new_n1898_ = new_n1775_ & new_n1897_;
  assign new_n1899_ = new_n1769_ & new_n1772_;
  assign new_n1900_ = new_n1766_ & new_n1899_;
  assign new_n1901_ = new_n1898_ & new_n1900_;
  assign new_n1902_ = ~new_n1860_ & ~new_n1901_;
  assign new_n1903_ = new_n1896_ & new_n1902_;
  assign new_n1904_ = new_n1895_ & new_n1903_;
  assign new_n1905_ = new_n1892_ & new_n1904_;
  assign new_n1906_ = new_n1886_ & new_n1905_;
  assign new_n1907_ = ~new_n1873_ & new_n1906_;
  assign new_n1908_ = ~\data<18>  & ~new_n1907_;
  assign new_n1909_ = \data<18>  & new_n1907_;
  assign new_n1910_ = ~new_n1908_ & ~new_n1909_;
  assign new_n1911_ = new_n504_ & ~new_n1910_;
  assign new_n1912_ = \outreg<45>  & ~\count<0> ;
  assign new_n1913_ = \outreg<53>  & \count<0> ;
  assign new_n1914_ = ~new_n1912_ & ~new_n1913_;
  assign new_n1915_ = ~new_n504_ & ~new_n1914_;
  assign \outreg_new<45>  = new_n1911_ | new_n1915_;
  assign new_n1917_ = \data<50>  & new_n504_;
  assign new_n1918_ = \outreg<44>  & ~\count<0> ;
  assign new_n1919_ = \outreg<52>  & \count<0> ;
  assign new_n1920_ = ~new_n1918_ & ~new_n1919_;
  assign new_n1921_ = ~new_n504_ & ~new_n1920_;
  assign \outreg_new<44>  = new_n1917_ | new_n1921_;
  assign new_n1923_ = new_n1778_ & new_n1784_;
  assign new_n1924_ = new_n1781_ & new_n1923_;
  assign new_n1925_ = new_n1781_ & new_n1813_;
  assign new_n1926_ = new_n1778_ & new_n1800_;
  assign new_n1927_ = new_n1781_ & new_n1926_;
  assign new_n1928_ = new_n1778_ & new_n1808_;
  assign new_n1929_ = ~new_n1781_ & new_n1928_;
  assign new_n1930_ = new_n1778_ & new_n1793_;
  assign new_n1931_ = ~new_n1781_ & new_n1930_;
  assign new_n1932_ = ~new_n1778_ & new_n1796_;
  assign new_n1933_ = ~new_n1781_ & new_n1932_;
  assign new_n1934_ = new_n1781_ & new_n1846_;
  assign new_n1935_ = new_n1781_ & new_n1857_;
  assign new_n1936_ = new_n1781_ & new_n1859_;
  assign new_n1937_ = ~new_n1781_ & new_n1832_;
  assign new_n1938_ = ~new_n1778_ & new_n1836_;
  assign new_n1939_ = ~new_n1781_ & new_n1938_;
  assign new_n1940_ = new_n1778_ & new_n1840_;
  assign new_n1941_ = ~new_n1781_ & new_n1940_;
  assign new_n1942_ = ~new_n1786_ & ~new_n1925_;
  assign new_n1943_ = ~new_n1924_ & new_n1942_;
  assign new_n1944_ = ~new_n1798_ & ~new_n1927_;
  assign new_n1945_ = ~new_n1802_ & ~new_n1807_;
  assign new_n1946_ = new_n1944_ & new_n1945_;
  assign new_n1947_ = new_n1943_ & new_n1946_;
  assign new_n1948_ = ~new_n1810_ & ~new_n1811_;
  assign new_n1949_ = ~new_n1929_ & new_n1948_;
  assign new_n1950_ = ~new_n1931_ & ~new_n1933_;
  assign new_n1951_ = new_n1883_ & new_n1950_;
  assign new_n1952_ = new_n1949_ & new_n1951_;
  assign new_n1953_ = new_n1947_ & new_n1952_;
  assign new_n1954_ = ~new_n1827_ & ~new_n1833_;
  assign new_n1955_ = ~new_n1934_ & new_n1954_;
  assign new_n1956_ = ~new_n1838_ & ~new_n1935_;
  assign new_n1957_ = ~new_n1845_ & ~new_n1936_;
  assign new_n1958_ = new_n1956_ & new_n1957_;
  assign new_n1959_ = new_n1955_ & new_n1958_;
  assign new_n1960_ = ~new_n1854_ & ~new_n1937_;
  assign new_n1961_ = ~new_n1847_ & new_n1960_;
  assign new_n1962_ = ~new_n1855_ & ~new_n1939_;
  assign new_n1963_ = ~new_n1858_ & ~new_n1941_;
  assign new_n1964_ = new_n1962_ & new_n1963_;
  assign new_n1965_ = new_n1961_ & new_n1964_;
  assign new_n1966_ = new_n1959_ & new_n1965_;
  assign new_n1967_ = new_n1953_ & new_n1966_;
  assign new_n1968_ = new_n1766_ & ~new_n1778_;
  assign new_n1969_ = ~new_n1766_ & new_n1778_;
  assign new_n1970_ = ~new_n1968_ & ~new_n1969_;
  assign new_n1971_ = ~new_n1865_ & ~new_n1970_;
  assign new_n1972_ = new_n1769_ & new_n1971_;
  assign new_n1973_ = new_n1967_ & ~new_n1972_;
  assign new_n1974_ = ~\data<10>  & ~new_n1973_;
  assign new_n1975_ = \data<10>  & new_n1973_;
  assign new_n1976_ = ~new_n1974_ & ~new_n1975_;
  assign new_n1977_ = new_n504_ & ~new_n1976_;
  assign new_n1978_ = \outreg<43>  & ~\count<0> ;
  assign new_n1979_ = \outreg<51>  & \count<0> ;
  assign new_n1980_ = ~new_n1978_ & ~new_n1979_;
  assign new_n1981_ = ~new_n504_ & ~new_n1980_;
  assign \outreg_new<43>  = new_n1977_ | new_n1981_;
  assign new_n1983_ = \data<42>  & new_n504_;
  assign new_n1984_ = \outreg<42>  & ~\count<0> ;
  assign new_n1985_ = \outreg<50>  & \count<0> ;
  assign new_n1986_ = ~new_n1984_ & ~new_n1985_;
  assign new_n1987_ = ~new_n504_ & ~new_n1986_;
  assign \outreg_new<42>  = new_n1983_ | new_n1987_;
  assign new_n1989_ = new_n740_ & new_n760_;
  assign new_n1990_ = ~new_n743_ & new_n1989_;
  assign new_n1991_ = new_n746_ & new_n1990_;
  assign new_n1992_ = new_n746_ & new_n780_;
  assign new_n1993_ = new_n746_ & new_n782_;
  assign new_n1994_ = ~new_n746_ & new_n755_;
  assign new_n1995_ = new_n743_ & new_n1989_;
  assign new_n1996_ = ~new_n746_ & new_n1995_;
  assign new_n1997_ = ~new_n743_ & new_n779_;
  assign new_n1998_ = ~new_n746_ & new_n1997_;
  assign new_n1999_ = new_n746_ & new_n814_;
  assign new_n2000_ = new_n746_ & new_n817_;
  assign new_n2001_ = ~new_n740_ & new_n797_;
  assign new_n2002_ = ~new_n743_ & new_n2001_;
  assign new_n2003_ = new_n746_ & new_n2002_;
  assign new_n2004_ = ~new_n743_ & new_n793_;
  assign new_n2005_ = ~new_n746_ & new_n2004_;
  assign new_n2006_ = ~new_n746_ & new_n2002_;
  assign new_n2007_ = new_n743_ & new_n807_;
  assign new_n2008_ = ~new_n746_ & new_n2007_;
  assign new_n2009_ = new_n740_ & ~new_n746_;
  assign new_n2010_ = ~new_n737_ & new_n2009_;
  assign new_n2011_ = ~new_n740_ & new_n746_;
  assign new_n2012_ = new_n737_ & new_n2011_;
  assign new_n2013_ = ~new_n2010_ & ~new_n2012_;
  assign new_n2014_ = new_n743_ & ~new_n2013_;
  assign new_n2015_ = ~new_n731_ & new_n2014_;
  assign new_n2016_ = ~new_n737_ & ~new_n746_;
  assign new_n2017_ = new_n737_ & new_n746_;
  assign new_n2018_ = ~new_n2016_ & ~new_n2017_;
  assign new_n2019_ = ~new_n743_ & ~new_n2018_;
  assign new_n2020_ = ~new_n740_ & new_n2019_;
  assign new_n2021_ = new_n731_ & new_n2020_;
  assign new_n2022_ = ~new_n2015_ & ~new_n2021_;
  assign new_n2023_ = new_n734_ & ~new_n2022_;
  assign new_n2024_ = ~new_n756_ & ~new_n1991_;
  assign new_n2025_ = ~new_n751_ & new_n2024_;
  assign new_n2026_ = ~new_n763_ & ~new_n765_;
  assign new_n2027_ = ~new_n1992_ & ~new_n1993_;
  assign new_n2028_ = new_n2026_ & new_n2027_;
  assign new_n2029_ = new_n2025_ & new_n2028_;
  assign new_n2030_ = ~new_n776_ & ~new_n1994_;
  assign new_n2031_ = ~new_n775_ & new_n2030_;
  assign new_n2032_ = ~new_n777_ & ~new_n1996_;
  assign new_n2033_ = ~new_n781_ & ~new_n1998_;
  assign new_n2034_ = new_n2032_ & new_n2033_;
  assign new_n2035_ = new_n2031_ & new_n2034_;
  assign new_n2036_ = new_n2029_ & new_n2035_;
  assign new_n2037_ = ~new_n795_ & ~new_n1999_;
  assign new_n2038_ = ~new_n788_ & new_n2037_;
  assign new_n2039_ = ~new_n800_ & ~new_n2000_;
  assign new_n2040_ = ~new_n806_ & ~new_n2003_;
  assign new_n2041_ = new_n2039_ & new_n2040_;
  assign new_n2042_ = new_n2038_ & new_n2041_;
  assign new_n2043_ = ~new_n813_ & ~new_n2005_;
  assign new_n2044_ = ~new_n812_ & new_n2043_;
  assign new_n2045_ = ~new_n818_ & ~new_n2006_;
  assign new_n2046_ = ~new_n820_ & ~new_n2008_;
  assign new_n2047_ = new_n2045_ & new_n2046_;
  assign new_n2048_ = new_n2044_ & new_n2047_;
  assign new_n2049_ = new_n2042_ & new_n2048_;
  assign new_n2050_ = new_n2036_ & new_n2049_;
  assign new_n2051_ = ~new_n2023_ & new_n2050_;
  assign new_n2052_ = ~\data<2>  & ~new_n2051_;
  assign new_n2053_ = \data<2>  & new_n2051_;
  assign new_n2054_ = ~new_n2052_ & ~new_n2053_;
  assign new_n2055_ = new_n504_ & ~new_n2054_;
  assign new_n2056_ = \outreg<41>  & ~\count<0> ;
  assign new_n2057_ = \outreg<49>  & \count<0> ;
  assign new_n2058_ = ~new_n2056_ & ~new_n2057_;
  assign new_n2059_ = ~new_n504_ & ~new_n2058_;
  assign \outreg_new<41>  = new_n2055_ | new_n2059_;
  assign new_n2061_ = \data<34>  & new_n504_;
  assign new_n2062_ = \outreg<40>  & ~\count<0> ;
  assign new_n2063_ = \outreg<48>  & \count<0> ;
  assign new_n2064_ = ~new_n2062_ & ~new_n2063_;
  assign new_n2065_ = ~new_n504_ & ~new_n2064_;
  assign \outreg_new<40>  = new_n2061_ | new_n2065_;
  assign new_n2067_ = ~new_n1332_ & new_n1344_;
  assign new_n2068_ = ~new_n1332_ & new_n1534_;
  assign new_n2069_ = new_n1332_ & new_n1389_;
  assign new_n2070_ = new_n1329_ & new_n1405_;
  assign new_n2071_ = new_n1332_ & new_n2070_;
  assign new_n2072_ = ~new_n1345_ & ~new_n2067_;
  assign new_n2073_ = ~new_n1342_ & new_n2072_;
  assign new_n2074_ = ~new_n1351_ & ~new_n1532_;
  assign new_n2075_ = ~new_n1356_ & ~new_n1363_;
  assign new_n2076_ = new_n2074_ & new_n2075_;
  assign new_n2077_ = new_n2073_ & new_n2076_;
  assign new_n2078_ = ~new_n1367_ & ~new_n2068_;
  assign new_n2079_ = ~new_n1535_ & new_n2078_;
  assign new_n2080_ = ~new_n1370_ & ~new_n1537_;
  assign new_n2081_ = new_n1566_ & new_n2080_;
  assign new_n2082_ = new_n2079_ & new_n2081_;
  assign new_n2083_ = new_n2077_ & new_n2082_;
  assign new_n2084_ = new_n1438_ & ~new_n1540_;
  assign new_n2085_ = ~new_n1390_ & ~new_n2069_;
  assign new_n2086_ = new_n1442_ & new_n2085_;
  assign new_n2087_ = new_n2084_ & new_n2086_;
  assign new_n2088_ = ~new_n1544_ & ~new_n2071_;
  assign new_n2089_ = ~new_n1401_ & new_n2088_;
  assign new_n2090_ = ~new_n1408_ & ~new_n1547_;
  assign new_n2091_ = ~new_n1410_ & ~new_n1548_;
  assign new_n2092_ = new_n2090_ & new_n2091_;
  assign new_n2093_ = new_n2089_ & new_n2092_;
  assign new_n2094_ = new_n2087_ & new_n2093_;
  assign new_n2095_ = new_n2083_ & new_n2094_;
  assign new_n2096_ = ~new_n1323_ & new_n1332_;
  assign new_n2097_ = new_n1323_ & ~new_n1332_;
  assign new_n2098_ = ~new_n2096_ & ~new_n2097_;
  assign new_n2099_ = new_n1320_ & ~new_n2098_;
  assign new_n2100_ = ~new_n1317_ & new_n2099_;
  assign new_n2101_ = new_n1352_ & new_n1411_;
  assign new_n2102_ = ~new_n2100_ & ~new_n2101_;
  assign new_n2103_ = ~new_n1329_ & ~new_n2102_;
  assign new_n2104_ = new_n1323_ & new_n1582_;
  assign new_n2105_ = new_n1352_ & new_n2104_;
  assign new_n2106_ = ~new_n2103_ & ~new_n2105_;
  assign new_n2107_ = new_n1326_ & ~new_n2106_;
  assign new_n2108_ = new_n2095_ & ~new_n2107_;
  assign new_n2109_ = ~\data<27>  & ~new_n2108_;
  assign new_n2110_ = \data<27>  & new_n2108_;
  assign new_n2111_ = ~new_n2109_ & ~new_n2110_;
  assign new_n2112_ = new_n504_ & ~new_n2111_;
  assign new_n2113_ = \outreg<39>  & ~\count<0> ;
  assign new_n2114_ = \outreg<47>  & \count<0> ;
  assign new_n2115_ = ~new_n2113_ & ~new_n2114_;
  assign new_n2116_ = ~new_n504_ & ~new_n2115_;
  assign \outreg_new<39>  = new_n2112_ | new_n2116_;
  assign new_n2118_ = \data<59>  & new_n504_;
  assign new_n2119_ = \outreg<38>  & ~\count<0> ;
  assign new_n2120_ = \outreg<46>  & \count<0> ;
  assign new_n2121_ = ~new_n2119_ & ~new_n2120_;
  assign new_n2122_ = ~new_n504_ & ~new_n2121_;
  assign \outreg_new<38>  = new_n2118_ | new_n2122_;
  assign new_n2124_ = ~new_n1116_ & ~new_n1239_;
  assign new_n2125_ = ~new_n1114_ & new_n2124_;
  assign new_n2126_ = ~new_n1128_ & ~new_n1472_;
  assign new_n2127_ = new_n1270_ & new_n2126_;
  assign new_n2128_ = new_n2125_ & new_n2127_;
  assign new_n2129_ = ~new_n1139_ & ~new_n1474_;
  assign new_n2130_ = ~new_n1136_ & new_n2129_;
  assign new_n2131_ = ~new_n1142_ & ~new_n1147_;
  assign new_n2132_ = ~new_n1243_ & ~new_n1246_;
  assign new_n2133_ = new_n2131_ & new_n2132_;
  assign new_n2134_ = new_n2130_ & new_n2133_;
  assign new_n2135_ = new_n2128_ & new_n2134_;
  assign new_n2136_ = ~new_n1160_ & ~new_n1249_;
  assign new_n2137_ = ~new_n1475_ & new_n2136_;
  assign new_n2138_ = ~new_n1174_ & ~new_n1250_;
  assign new_n2139_ = new_n1202_ & new_n2138_;
  assign new_n2140_ = new_n2137_ & new_n2139_;
  assign new_n2141_ = ~new_n1180_ & ~new_n1477_;
  assign new_n2142_ = ~new_n1179_ & new_n2141_;
  assign new_n2143_ = ~new_n1182_ & ~new_n1252_;
  assign new_n2144_ = new_n1499_ & new_n2143_;
  assign new_n2145_ = new_n2142_ & new_n2144_;
  assign new_n2146_ = new_n2140_ & new_n2145_;
  assign new_n2147_ = new_n2135_ & new_n2146_;
  assign new_n2148_ = ~new_n1094_ & ~new_n1106_;
  assign new_n2149_ = new_n1094_ & new_n1106_;
  assign new_n2150_ = ~new_n2148_ & ~new_n2149_;
  assign new_n2151_ = new_n1103_ & ~new_n1109_;
  assign new_n2152_ = new_n1100_ & new_n2151_;
  assign new_n2153_ = ~new_n1103_ & new_n1109_;
  assign new_n2154_ = ~new_n1100_ & new_n2153_;
  assign new_n2155_ = ~new_n2152_ & ~new_n2154_;
  assign new_n2156_ = ~new_n2150_ & ~new_n2155_;
  assign new_n2157_ = ~new_n1097_ & new_n2156_;
  assign new_n2158_ = new_n2147_ & ~new_n2157_;
  assign new_n2159_ = ~\data<19>  & ~new_n2158_;
  assign new_n2160_ = \data<19>  & new_n2158_;
  assign new_n2161_ = ~new_n2159_ & ~new_n2160_;
  assign new_n2162_ = new_n504_ & ~new_n2161_;
  assign new_n2163_ = \outreg<37>  & ~\count<0> ;
  assign new_n2164_ = \outreg<45>  & \count<0> ;
  assign new_n2165_ = ~new_n2163_ & ~new_n2164_;
  assign new_n2166_ = ~new_n504_ & ~new_n2165_;
  assign \outreg_new<37>  = new_n2162_ | new_n2166_;
  assign new_n2168_ = \data<51>  & new_n504_;
  assign new_n2169_ = \outreg<36>  & ~\count<0> ;
  assign new_n2170_ = \outreg<44>  & \count<0> ;
  assign new_n2171_ = ~new_n2169_ & ~new_n2170_;
  assign new_n2172_ = ~new_n504_ & ~new_n2171_;
  assign \outreg_new<36>  = new_n2168_ | new_n2172_;
  assign new_n2174_ = \data<55>  & ~\D<15> ;
  assign new_n2175_ = ~\data<55>  & \D<15> ;
  assign new_n2176_ = ~new_n2174_ & ~new_n2175_;
  assign new_n2177_ = \data<56>  & ~\D<20> ;
  assign new_n2178_ = ~\data<56>  & \D<20> ;
  assign new_n2179_ = ~new_n2177_ & ~new_n2178_;
  assign new_n2180_ = \data<57>  & ~\D<10> ;
  assign new_n2181_ = ~\data<57>  & \D<10> ;
  assign new_n2182_ = ~new_n2180_ & ~new_n2181_;
  assign new_n2183_ = \data<58>  & ~\D<27> ;
  assign new_n2184_ = ~\data<58>  & \D<27> ;
  assign new_n2185_ = ~new_n2183_ & ~new_n2184_;
  assign new_n2186_ = \data<59>  & ~\D<5> ;
  assign new_n2187_ = ~\data<59>  & \D<5> ;
  assign new_n2188_ = ~new_n2186_ & ~new_n2187_;
  assign new_n2189_ = \data<60>  & ~\D<24> ;
  assign new_n2190_ = ~\data<60>  & \D<24> ;
  assign new_n2191_ = ~new_n2189_ & ~new_n2190_;
  assign new_n2192_ = new_n2176_ & new_n2179_;
  assign new_n2193_ = new_n2182_ & new_n2192_;
  assign new_n2194_ = ~new_n2185_ & new_n2193_;
  assign new_n2195_ = ~new_n2188_ & new_n2194_;
  assign new_n2196_ = new_n2191_ & new_n2195_;
  assign new_n2197_ = ~new_n2182_ & new_n2192_;
  assign new_n2198_ = new_n2185_ & new_n2197_;
  assign new_n2199_ = new_n2188_ & new_n2198_;
  assign new_n2200_ = new_n2191_ & new_n2199_;
  assign new_n2201_ = ~new_n2185_ & new_n2197_;
  assign new_n2202_ = ~new_n2188_ & new_n2201_;
  assign new_n2203_ = new_n2191_ & new_n2202_;
  assign new_n2204_ = new_n2176_ & ~new_n2179_;
  assign new_n2205_ = new_n2182_ & new_n2204_;
  assign new_n2206_ = new_n2185_ & new_n2205_;
  assign new_n2207_ = ~new_n2188_ & new_n2206_;
  assign new_n2208_ = new_n2191_ & new_n2207_;
  assign new_n2209_ = ~new_n2185_ & new_n2205_;
  assign new_n2210_ = ~new_n2188_ & new_n2209_;
  assign new_n2211_ = new_n2191_ & new_n2210_;
  assign new_n2212_ = ~new_n2182_ & new_n2204_;
  assign new_n2213_ = new_n2185_ & new_n2212_;
  assign new_n2214_ = new_n2188_ & new_n2213_;
  assign new_n2215_ = new_n2191_ & new_n2214_;
  assign new_n2216_ = ~new_n2185_ & new_n2212_;
  assign new_n2217_ = new_n2188_ & new_n2216_;
  assign new_n2218_ = new_n2191_ & new_n2217_;
  assign new_n2219_ = new_n2185_ & new_n2193_;
  assign new_n2220_ = new_n2188_ & new_n2219_;
  assign new_n2221_ = ~new_n2191_ & new_n2220_;
  assign new_n2222_ = ~new_n2191_ & new_n2195_;
  assign new_n2223_ = new_n2188_ & new_n2206_;
  assign new_n2224_ = ~new_n2191_ & new_n2223_;
  assign new_n2225_ = new_n2188_ & new_n2209_;
  assign new_n2226_ = ~new_n2191_ & new_n2225_;
  assign new_n2227_ = ~new_n2191_ & new_n2210_;
  assign new_n2228_ = ~new_n2188_ & new_n2213_;
  assign new_n2229_ = ~new_n2191_ & new_n2228_;
  assign new_n2230_ = ~new_n2188_ & new_n2216_;
  assign new_n2231_ = ~new_n2191_ & new_n2230_;
  assign new_n2232_ = ~new_n2176_ & new_n2179_;
  assign new_n2233_ = new_n2182_ & new_n2232_;
  assign new_n2234_ = ~new_n2185_ & new_n2233_;
  assign new_n2235_ = ~new_n2188_ & new_n2234_;
  assign new_n2236_ = new_n2191_ & new_n2235_;
  assign new_n2237_ = ~new_n2182_ & new_n2232_;
  assign new_n2238_ = new_n2185_ & new_n2237_;
  assign new_n2239_ = new_n2188_ & new_n2238_;
  assign new_n2240_ = new_n2191_ & new_n2239_;
  assign new_n2241_ = ~new_n2185_ & new_n2237_;
  assign new_n2242_ = new_n2188_ & new_n2241_;
  assign new_n2243_ = new_n2191_ & new_n2242_;
  assign new_n2244_ = ~new_n2188_ & new_n2241_;
  assign new_n2245_ = new_n2191_ & new_n2244_;
  assign new_n2246_ = ~new_n2176_ & ~new_n2179_;
  assign new_n2247_ = new_n2182_ & new_n2246_;
  assign new_n2248_ = new_n2185_ & new_n2247_;
  assign new_n2249_ = ~new_n2188_ & new_n2248_;
  assign new_n2250_ = new_n2191_ & new_n2249_;
  assign new_n2251_ = ~new_n2185_ & new_n2247_;
  assign new_n2252_ = new_n2188_ & new_n2251_;
  assign new_n2253_ = new_n2191_ & new_n2252_;
  assign new_n2254_ = ~new_n2182_ & new_n2246_;
  assign new_n2255_ = new_n2185_ & new_n2254_;
  assign new_n2256_ = ~new_n2188_ & new_n2255_;
  assign new_n2257_ = new_n2191_ & new_n2256_;
  assign new_n2258_ = new_n2185_ & new_n2233_;
  assign new_n2259_ = new_n2188_ & new_n2258_;
  assign new_n2260_ = ~new_n2191_ & new_n2259_;
  assign new_n2261_ = new_n2188_ & new_n2234_;
  assign new_n2262_ = ~new_n2191_ & new_n2261_;
  assign new_n2263_ = ~new_n2191_ & new_n2244_;
  assign new_n2264_ = ~new_n2191_ & new_n2249_;
  assign new_n2265_ = ~new_n2188_ & new_n2251_;
  assign new_n2266_ = ~new_n2191_ & new_n2265_;
  assign new_n2267_ = new_n2188_ & new_n2255_;
  assign new_n2268_ = ~new_n2191_ & new_n2267_;
  assign new_n2269_ = ~new_n2185_ & new_n2254_;
  assign new_n2270_ = ~new_n2188_ & new_n2269_;
  assign new_n2271_ = ~new_n2191_ & new_n2270_;
  assign new_n2272_ = ~new_n2200_ & ~new_n2203_;
  assign new_n2273_ = ~new_n2196_ & new_n2272_;
  assign new_n2274_ = ~new_n2208_ & ~new_n2211_;
  assign new_n2275_ = ~new_n2215_ & ~new_n2218_;
  assign new_n2276_ = new_n2274_ & new_n2275_;
  assign new_n2277_ = new_n2273_ & new_n2276_;
  assign new_n2278_ = ~new_n2222_ & ~new_n2224_;
  assign new_n2279_ = ~new_n2221_ & new_n2278_;
  assign new_n2280_ = ~new_n2226_ & ~new_n2227_;
  assign new_n2281_ = ~new_n2229_ & ~new_n2231_;
  assign new_n2282_ = new_n2280_ & new_n2281_;
  assign new_n2283_ = new_n2279_ & new_n2282_;
  assign new_n2284_ = new_n2277_ & new_n2283_;
  assign new_n2285_ = ~new_n2240_ & ~new_n2243_;
  assign new_n2286_ = ~new_n2236_ & new_n2285_;
  assign new_n2287_ = ~new_n2245_ & ~new_n2250_;
  assign new_n2288_ = ~new_n2253_ & ~new_n2257_;
  assign new_n2289_ = new_n2287_ & new_n2288_;
  assign new_n2290_ = new_n2286_ & new_n2289_;
  assign new_n2291_ = ~new_n2262_ & ~new_n2263_;
  assign new_n2292_ = ~new_n2260_ & new_n2291_;
  assign new_n2293_ = ~new_n2264_ & ~new_n2266_;
  assign new_n2294_ = ~new_n2268_ & ~new_n2271_;
  assign new_n2295_ = new_n2293_ & new_n2294_;
  assign new_n2296_ = new_n2292_ & new_n2295_;
  assign new_n2297_ = new_n2290_ & new_n2296_;
  assign new_n2298_ = new_n2284_ & new_n2297_;
  assign new_n2299_ = ~new_n2182_ & ~new_n2191_;
  assign new_n2300_ = new_n2182_ & new_n2191_;
  assign new_n2301_ = ~new_n2299_ & ~new_n2300_;
  assign new_n2302_ = ~new_n2176_ & ~new_n2188_;
  assign new_n2303_ = new_n2176_ & new_n2188_;
  assign new_n2304_ = ~new_n2302_ & ~new_n2303_;
  assign new_n2305_ = ~new_n2301_ & ~new_n2304_;
  assign new_n2306_ = new_n2185_ & new_n2305_;
  assign new_n2307_ = new_n2179_ & new_n2306_;
  assign new_n2308_ = new_n2298_ & ~new_n2307_;
  assign new_n2309_ = ~\data<11>  & ~new_n2308_;
  assign new_n2310_ = \data<11>  & new_n2308_;
  assign new_n2311_ = ~new_n2309_ & ~new_n2310_;
  assign new_n2312_ = new_n504_ & ~new_n2311_;
  assign new_n2313_ = \outreg<35>  & ~\count<0> ;
  assign new_n2314_ = \outreg<43>  & \count<0> ;
  assign new_n2315_ = ~new_n2313_ & ~new_n2314_;
  assign new_n2316_ = ~new_n504_ & ~new_n2315_;
  assign \outreg_new<35>  = new_n2312_ | new_n2316_;
  assign new_n2318_ = \data<43>  & new_n504_;
  assign new_n2319_ = \outreg<34>  & ~\count<0> ;
  assign new_n2320_ = \outreg<42>  & \count<0> ;
  assign new_n2321_ = ~new_n2319_ & ~new_n2320_;
  assign new_n2322_ = ~new_n504_ & ~new_n2321_;
  assign \outreg_new<34>  = new_n2318_ | new_n2322_;
  assign new_n2324_ = new_n1781_ & new_n1928_;
  assign new_n2325_ = ~new_n1778_ & new_n1788_;
  assign new_n2326_ = ~new_n1781_ & new_n2325_;
  assign new_n2327_ = new_n1781_ & new_n1853_;
  assign new_n2328_ = ~new_n1781_ & new_n1828_;
  assign new_n2329_ = ~new_n1786_ & ~new_n1924_;
  assign new_n2330_ = ~new_n2324_ & new_n2329_;
  assign new_n2331_ = ~new_n1807_ & ~new_n1927_;
  assign new_n2332_ = new_n1874_ & new_n2331_;
  assign new_n2333_ = new_n2330_ & new_n2332_;
  assign new_n2334_ = ~new_n1810_ & ~new_n2326_;
  assign new_n2335_ = ~new_n1929_ & new_n2334_;
  assign new_n2336_ = ~new_n1814_ & ~new_n1817_;
  assign new_n2337_ = ~new_n1818_ & ~new_n1933_;
  assign new_n2338_ = new_n2336_ & new_n2337_;
  assign new_n2339_ = new_n2335_ & new_n2338_;
  assign new_n2340_ = new_n2333_ & new_n2339_;
  assign new_n2341_ = ~new_n1827_ & ~new_n1934_;
  assign new_n2342_ = ~new_n1824_ & new_n2341_;
  assign new_n2343_ = ~new_n1935_ & ~new_n2327_;
  assign new_n2344_ = new_n1890_ & new_n2343_;
  assign new_n2345_ = new_n2342_ & new_n2344_;
  assign new_n2346_ = ~new_n1850_ & ~new_n1854_;
  assign new_n2347_ = ~new_n2328_ & new_n2346_;
  assign new_n2348_ = ~new_n1855_ & ~new_n1937_;
  assign new_n2349_ = ~new_n1860_ & ~new_n1939_;
  assign new_n2350_ = new_n2348_ & new_n2349_;
  assign new_n2351_ = new_n2347_ & new_n2350_;
  assign new_n2352_ = new_n2345_ & new_n2351_;
  assign new_n2353_ = new_n2340_ & new_n2352_;
  assign new_n2354_ = new_n1778_ & ~new_n1781_;
  assign new_n2355_ = ~new_n1769_ & ~new_n1775_;
  assign new_n2356_ = new_n2354_ & new_n2355_;
  assign new_n2357_ = new_n1769_ & new_n1775_;
  assign new_n2358_ = new_n1897_ & new_n2357_;
  assign new_n2359_ = ~new_n2356_ & ~new_n2358_;
  assign new_n2360_ = ~new_n1766_ & ~new_n2359_;
  assign new_n2361_ = ~new_n1769_ & ~new_n1781_;
  assign new_n2362_ = new_n1769_ & new_n1781_;
  assign new_n2363_ = ~new_n2361_ & ~new_n2362_;
  assign new_n2364_ = ~new_n1778_ & ~new_n2363_;
  assign new_n2365_ = ~new_n1775_ & new_n2364_;
  assign new_n2366_ = new_n1766_ & new_n2365_;
  assign new_n2367_ = ~new_n2360_ & ~new_n2366_;
  assign new_n2368_ = ~new_n1772_ & ~new_n2367_;
  assign new_n2369_ = new_n2353_ & ~new_n2368_;
  assign new_n2370_ = ~\data<3>  & ~new_n2369_;
  assign new_n2371_ = \data<3>  & new_n2369_;
  assign new_n2372_ = ~new_n2370_ & ~new_n2371_;
  assign new_n2373_ = new_n504_ & ~new_n2372_;
  assign new_n2374_ = \outreg<33>  & ~\count<0> ;
  assign new_n2375_ = \outreg<41>  & \count<0> ;
  assign new_n2376_ = ~new_n2374_ & ~new_n2375_;
  assign new_n2377_ = ~new_n504_ & ~new_n2376_;
  assign \outreg_new<33>  = new_n2373_ | new_n2377_;
  assign new_n2379_ = \data<35>  & new_n504_;
  assign new_n2380_ = \outreg<32>  & ~\count<0> ;
  assign new_n2381_ = \outreg<40>  & \count<0> ;
  assign new_n2382_ = ~new_n2380_ & ~new_n2381_;
  assign new_n2383_ = ~new_n504_ & ~new_n2382_;
  assign \outreg_new<32>  = new_n2379_ | new_n2383_;
  assign new_n2385_ = new_n1942_ & ~new_n2324_;
  assign new_n2386_ = ~new_n1795_ & ~new_n1927_;
  assign new_n2387_ = ~new_n1802_ & ~new_n1805_;
  assign new_n2388_ = new_n2386_ & new_n2387_;
  assign new_n2389_ = new_n2385_ & new_n2388_;
  assign new_n2390_ = ~new_n1811_ & ~new_n2326_;
  assign new_n2391_ = ~new_n1810_ & new_n2390_;
  assign new_n2392_ = ~new_n1816_ & ~new_n1931_;
  assign new_n2393_ = ~new_n1817_ & ~new_n1933_;
  assign new_n2394_ = new_n2392_ & new_n2393_;
  assign new_n2395_ = new_n2391_ & new_n2394_;
  assign new_n2396_ = new_n2389_ & new_n2395_;
  assign new_n2397_ = new_n1887_ & ~new_n1934_;
  assign new_n2398_ = ~new_n1838_ & ~new_n2327_;
  assign new_n2399_ = ~new_n1842_ & ~new_n1936_;
  assign new_n2400_ = new_n2398_ & new_n2399_;
  assign new_n2401_ = new_n2397_ & new_n2400_;
  assign new_n2402_ = new_n1894_ & ~new_n2328_;
  assign new_n2403_ = ~new_n1858_ & ~new_n1939_;
  assign new_n2404_ = ~new_n1860_ & ~new_n1941_;
  assign new_n2405_ = new_n2403_ & new_n2404_;
  assign new_n2406_ = new_n2402_ & new_n2405_;
  assign new_n2407_ = new_n2401_ & new_n2406_;
  assign new_n2408_ = new_n2396_ & new_n2407_;
  assign new_n2409_ = new_n1775_ & ~new_n1781_;
  assign new_n2410_ = new_n1769_ & new_n2409_;
  assign new_n2411_ = ~new_n1775_ & new_n1781_;
  assign new_n2412_ = ~new_n1769_ & new_n2411_;
  assign new_n2413_ = ~new_n2410_ & ~new_n2412_;
  assign new_n2414_ = ~new_n1766_ & ~new_n2413_;
  assign new_n2415_ = new_n1782_ & new_n1861_;
  assign new_n2416_ = ~new_n2414_ & ~new_n2415_;
  assign new_n2417_ = new_n1778_ & ~new_n2416_;
  assign new_n2418_ = ~new_n1775_ & new_n1897_;
  assign new_n2419_ = new_n1791_ & new_n2418_;
  assign new_n2420_ = ~new_n2417_ & ~new_n2419_;
  assign new_n2421_ = new_n1772_ & ~new_n2420_;
  assign new_n2422_ = new_n2408_ & ~new_n2421_;
  assign new_n2423_ = ~\data<28>  & ~new_n2422_;
  assign new_n2424_ = \data<28>  & new_n2422_;
  assign new_n2425_ = ~new_n2423_ & ~new_n2424_;
  assign new_n2426_ = new_n504_ & ~new_n2425_;
  assign new_n2427_ = \outreg<31>  & ~\count<0> ;
  assign new_n2428_ = \outreg<39>  & \count<0> ;
  assign new_n2429_ = ~new_n2427_ & ~new_n2428_;
  assign new_n2430_ = ~new_n504_ & ~new_n2429_;
  assign \outreg_new<31>  = new_n2426_ | new_n2430_;
  assign new_n2432_ = \data<60>  & new_n504_;
  assign new_n2433_ = \outreg<30>  & ~\count<0> ;
  assign new_n2434_ = \outreg<38>  & \count<0> ;
  assign new_n2435_ = ~new_n2433_ & ~new_n2434_;
  assign new_n2436_ = ~new_n504_ & ~new_n2435_;
  assign \outreg_new<30>  = new_n2432_ | new_n2436_;
  assign new_n2438_ = new_n1623_ & new_n1655_;
  assign new_n2439_ = new_n1623_ & new_n1660_;
  assign new_n2440_ = new_n1623_ & new_n1662_;
  assign new_n2441_ = ~new_n1623_ & new_n1633_;
  assign new_n2442_ = ~new_n1623_ & new_n1638_;
  assign new_n2443_ = ~new_n1623_ & new_n1645_;
  assign new_n2444_ = ~new_n1620_ & new_n1668_;
  assign new_n2445_ = new_n1623_ & new_n2444_;
  assign new_n2446_ = new_n1620_ & new_n1672_;
  assign new_n2447_ = new_n1623_ & new_n2446_;
  assign new_n2448_ = new_n1623_ & new_n1703_;
  assign new_n2449_ = new_n1620_ & new_n1683_;
  assign new_n2450_ = ~new_n1623_ & new_n2449_;
  assign new_n2451_ = ~new_n1623_ & new_n1688_;
  assign new_n2452_ = ~new_n1620_ & new_n1690_;
  assign new_n2453_ = ~new_n1623_ & new_n2452_;
  assign new_n2454_ = ~new_n1634_ & ~new_n2438_;
  assign new_n2455_ = ~new_n1628_ & new_n2454_;
  assign new_n2456_ = ~new_n2439_ & ~new_n2440_;
  assign new_n2457_ = ~new_n1643_ & ~new_n1648_;
  assign new_n2458_ = new_n2456_ & new_n2457_;
  assign new_n2459_ = new_n2455_ & new_n2458_;
  assign new_n2460_ = ~new_n1653_ & ~new_n2441_;
  assign new_n2461_ = ~new_n1650_ & new_n2460_;
  assign new_n2462_ = ~new_n1656_ & ~new_n1661_;
  assign new_n2463_ = ~new_n2442_ & ~new_n2443_;
  assign new_n2464_ = new_n2462_ & new_n2463_;
  assign new_n2465_ = new_n2461_ & new_n2464_;
  assign new_n2466_ = new_n2459_ & new_n2465_;
  assign new_n2467_ = ~new_n2445_ & ~new_n2447_;
  assign new_n2468_ = ~new_n1670_ & new_n2467_;
  assign new_n2469_ = ~new_n1685_ & ~new_n1689_;
  assign new_n2470_ = ~new_n1692_ & ~new_n2448_;
  assign new_n2471_ = new_n2469_ & new_n2470_;
  assign new_n2472_ = new_n2468_ & new_n2471_;
  assign new_n2473_ = ~new_n1699_ & ~new_n1701_;
  assign new_n2474_ = ~new_n1697_ & new_n2473_;
  assign new_n2475_ = ~new_n2450_ & ~new_n2451_;
  assign new_n2476_ = ~new_n1704_ & ~new_n2453_;
  assign new_n2477_ = new_n2475_ & new_n2476_;
  assign new_n2478_ = new_n2474_ & new_n2477_;
  assign new_n2479_ = new_n2472_ & new_n2478_;
  assign new_n2480_ = new_n2466_ & new_n2479_;
  assign new_n2481_ = ~new_n1706_ & ~new_n1708_;
  assign new_n2482_ = ~new_n1620_ & ~new_n2481_;
  assign new_n2483_ = ~new_n1608_ & new_n2482_;
  assign new_n2484_ = new_n1620_ & ~new_n1623_;
  assign new_n2485_ = new_n1608_ & new_n1617_;
  assign new_n2486_ = new_n2484_ & new_n2485_;
  assign new_n2487_ = ~new_n2483_ & ~new_n2486_;
  assign new_n2488_ = new_n1614_ & ~new_n2487_;
  assign new_n2489_ = new_n1608_ & ~new_n1614_;
  assign new_n2490_ = ~new_n1620_ & new_n1623_;
  assign new_n2491_ = ~new_n1617_ & new_n2490_;
  assign new_n2492_ = new_n2489_ & new_n2491_;
  assign new_n2493_ = ~new_n2488_ & ~new_n2492_;
  assign new_n2494_ = new_n1611_ & ~new_n2493_;
  assign new_n2495_ = new_n2480_ & ~new_n2494_;
  assign new_n2496_ = ~\data<20>  & ~new_n2495_;
  assign new_n2497_ = \data<20>  & new_n2495_;
  assign new_n2498_ = ~new_n2496_ & ~new_n2497_;
  assign new_n2499_ = new_n504_ & ~new_n2498_;
  assign new_n2500_ = \outreg<29>  & ~\count<0> ;
  assign new_n2501_ = \outreg<37>  & \count<0> ;
  assign new_n2502_ = ~new_n2500_ & ~new_n2501_;
  assign new_n2503_ = ~new_n504_ & ~new_n2502_;
  assign \outreg_new<29>  = new_n2499_ | new_n2503_;
  assign new_n2505_ = \data<52>  & new_n504_;
  assign new_n2506_ = \outreg<28>  & ~\count<0> ;
  assign new_n2507_ = \outreg<36>  & \count<0> ;
  assign new_n2508_ = ~new_n2506_ & ~new_n2507_;
  assign new_n2509_ = ~new_n504_ & ~new_n2508_;
  assign \outreg_new<28>  = new_n2505_ | new_n2509_;
  assign new_n2511_ = new_n1320_ & ~new_n1326_;
  assign new_n2512_ = ~new_n1320_ & new_n1326_;
  assign new_n2513_ = ~new_n2511_ & ~new_n2512_;
  assign new_n2514_ = new_n1332_ & ~new_n2513_;
  assign new_n2515_ = ~new_n1323_ & new_n2514_;
  assign new_n2516_ = ~new_n1317_ & new_n2515_;
  assign new_n2517_ = new_n1326_ & ~new_n1332_;
  assign new_n2518_ = new_n1323_ & new_n2517_;
  assign new_n2519_ = new_n1338_ & new_n2518_;
  assign new_n2520_ = ~new_n2516_ & ~new_n2519_;
  assign new_n2521_ = new_n1329_ & ~new_n2520_;
  assign new_n2522_ = ~new_n1342_ & ~new_n1530_;
  assign new_n2523_ = ~new_n1337_ & new_n2522_;
  assign new_n2524_ = ~new_n1347_ & ~new_n2067_;
  assign new_n2525_ = new_n1426_ & new_n2524_;
  assign new_n2526_ = new_n2523_ & new_n2525_;
  assign new_n2527_ = new_n1429_ & ~new_n1533_;
  assign new_n2528_ = ~new_n1537_ & ~new_n2068_;
  assign new_n2529_ = new_n1432_ & new_n2528_;
  assign new_n2530_ = new_n2527_ & new_n2529_;
  assign new_n2531_ = new_n2526_ & new_n2530_;
  assign new_n2532_ = ~new_n1379_ & ~new_n1384_;
  assign new_n2533_ = ~new_n1539_ & new_n2532_;
  assign new_n2534_ = ~new_n1388_ & ~new_n2069_;
  assign new_n2535_ = ~new_n1398_ & ~new_n1542_;
  assign new_n2536_ = new_n2534_ & new_n2535_;
  assign new_n2537_ = new_n2533_ & new_n2536_;
  assign new_n2538_ = ~new_n1546_ & ~new_n2071_;
  assign new_n2539_ = new_n1576_ & new_n2538_;
  assign new_n2540_ = ~new_n1404_ & ~new_n1407_;
  assign new_n2541_ = ~new_n1320_ & new_n1323_;
  assign new_n2542_ = new_n1317_ & new_n2541_;
  assign new_n2543_ = new_n1447_ & new_n2542_;
  assign new_n2544_ = ~new_n1548_ & ~new_n2543_;
  assign new_n2545_ = new_n2540_ & new_n2544_;
  assign new_n2546_ = new_n2539_ & new_n2545_;
  assign new_n2547_ = new_n2537_ & new_n2546_;
  assign new_n2548_ = new_n2531_ & new_n2547_;
  assign new_n2549_ = ~new_n2521_ & new_n2548_;
  assign new_n2550_ = ~\data<12>  & ~new_n2549_;
  assign new_n2551_ = \data<12>  & new_n2549_;
  assign new_n2552_ = ~new_n2550_ & ~new_n2551_;
  assign new_n2553_ = new_n504_ & ~new_n2552_;
  assign new_n2554_ = \outreg<27>  & ~\count<0> ;
  assign new_n2555_ = \outreg<35>  & \count<0> ;
  assign new_n2556_ = ~new_n2554_ & ~new_n2555_;
  assign new_n2557_ = ~new_n504_ & ~new_n2556_;
  assign \outreg_new<27>  = new_n2553_ | new_n2557_;
  assign new_n2559_ = \data<44>  & new_n504_;
  assign new_n2560_ = \outreg<26>  & ~\count<0> ;
  assign new_n2561_ = \outreg<34>  & \count<0> ;
  assign new_n2562_ = ~new_n2560_ & ~new_n2561_;
  assign new_n2563_ = ~new_n504_ & ~new_n2562_;
  assign \outreg_new<26>  = new_n2559_ | new_n2563_;
  assign new_n2565_ = new_n1623_ & new_n1658_;
  assign new_n2566_ = ~new_n1623_ & new_n1631_;
  assign new_n2567_ = new_n1623_ & new_n2449_;
  assign new_n2568_ = ~new_n1623_ & new_n1673_;
  assign new_n2569_ = ~new_n2439_ & ~new_n2565_;
  assign new_n2570_ = ~new_n1639_ & ~new_n1646_;
  assign new_n2571_ = new_n2569_ & new_n2570_;
  assign new_n2572_ = new_n2455_ & new_n2571_;
  assign new_n2573_ = ~new_n1653_ & ~new_n2566_;
  assign new_n2574_ = ~new_n1650_ & new_n2573_;
  assign new_n2575_ = ~new_n1659_ & ~new_n2442_;
  assign new_n2576_ = ~new_n1665_ & ~new_n2443_;
  assign new_n2577_ = new_n2575_ & new_n2576_;
  assign new_n2578_ = new_n2574_ & new_n2577_;
  assign new_n2579_ = new_n2572_ & new_n2578_;
  assign new_n2580_ = ~new_n1674_ & ~new_n2447_;
  assign new_n2581_ = ~new_n2445_ & new_n2580_;
  assign new_n2582_ = ~new_n1677_ & ~new_n2567_;
  assign new_n2583_ = new_n2469_ & new_n2582_;
  assign new_n2584_ = new_n2581_ & new_n2583_;
  assign new_n2585_ = ~new_n1699_ & ~new_n2568_;
  assign new_n2586_ = ~new_n1695_ & new_n2585_;
  assign new_n2587_ = ~new_n2450_ & ~new_n2453_;
  assign new_n2588_ = new_n1742_ & new_n2587_;
  assign new_n2589_ = new_n2586_ & new_n2588_;
  assign new_n2590_ = new_n2584_ & new_n2589_;
  assign new_n2591_ = new_n2579_ & new_n2590_;
  assign new_n2592_ = new_n1611_ & new_n2484_;
  assign new_n2593_ = ~new_n1611_ & new_n2490_;
  assign new_n2594_ = ~new_n2592_ & ~new_n2593_;
  assign new_n2595_ = ~new_n1614_ & ~new_n2594_;
  assign new_n2596_ = ~new_n1608_ & new_n2595_;
  assign new_n2597_ = ~new_n1620_ & ~new_n1623_;
  assign new_n2598_ = new_n1620_ & new_n1623_;
  assign new_n2599_ = ~new_n2597_ & ~new_n2598_;
  assign new_n2600_ = new_n1614_ & ~new_n2599_;
  assign new_n2601_ = new_n1611_ & new_n2600_;
  assign new_n2602_ = new_n1608_ & new_n2601_;
  assign new_n2603_ = ~new_n2596_ & ~new_n2602_;
  assign new_n2604_ = ~new_n1617_ & ~new_n2603_;
  assign new_n2605_ = new_n2591_ & ~new_n2604_;
  assign new_n2606_ = ~\data<4>  & ~new_n2605_;
  assign new_n2607_ = \data<4>  & new_n2605_;
  assign new_n2608_ = ~new_n2606_ & ~new_n2607_;
  assign new_n2609_ = new_n504_ & ~new_n2608_;
  assign new_n2610_ = \outreg<25>  & ~\count<0> ;
  assign new_n2611_ = \outreg<33>  & \count<0> ;
  assign new_n2612_ = ~new_n2610_ & ~new_n2611_;
  assign new_n2613_ = ~new_n504_ & ~new_n2612_;
  assign \outreg_new<25>  = new_n2609_ | new_n2613_;
  assign new_n2615_ = \data<36>  & new_n504_;
  assign new_n2616_ = \outreg<24>  & ~\count<0> ;
  assign new_n2617_ = \outreg<32>  & \count<0> ;
  assign new_n2618_ = ~new_n2616_ & ~new_n2617_;
  assign new_n2619_ = ~new_n504_ & ~new_n2618_;
  assign \outreg_new<24>  = new_n2615_ | new_n2619_;
  assign new_n2621_ = \data<39>  & ~\C<22> ;
  assign new_n2622_ = ~\data<39>  & \C<22> ;
  assign new_n2623_ = ~new_n2621_ & ~new_n2622_;
  assign new_n2624_ = \data<40>  & ~\C<18> ;
  assign new_n2625_ = ~\data<40>  & \C<18> ;
  assign new_n2626_ = ~new_n2624_ & ~new_n2625_;
  assign new_n2627_ = \data<41>  & ~\C<11> ;
  assign new_n2628_ = ~\data<41>  & \C<11> ;
  assign new_n2629_ = ~new_n2627_ & ~new_n2628_;
  assign new_n2630_ = \data<42>  & ~\C<3> ;
  assign new_n2631_ = ~\data<42>  & \C<3> ;
  assign new_n2632_ = ~new_n2630_ & ~new_n2631_;
  assign new_n2633_ = \data<43>  & ~\C<25> ;
  assign new_n2634_ = ~\data<43>  & \C<25> ;
  assign new_n2635_ = ~new_n2633_ & ~new_n2634_;
  assign new_n2636_ = \data<44>  & ~\C<7> ;
  assign new_n2637_ = ~\data<44>  & \C<7> ;
  assign new_n2638_ = ~new_n2636_ & ~new_n2637_;
  assign new_n2639_ = new_n2623_ & new_n2626_;
  assign new_n2640_ = new_n2629_ & new_n2639_;
  assign new_n2641_ = new_n2632_ & new_n2640_;
  assign new_n2642_ = new_n2635_ & new_n2641_;
  assign new_n2643_ = new_n2638_ & new_n2642_;
  assign new_n2644_ = ~new_n2632_ & new_n2640_;
  assign new_n2645_ = ~new_n2635_ & new_n2644_;
  assign new_n2646_ = new_n2638_ & new_n2645_;
  assign new_n2647_ = ~new_n2629_ & new_n2639_;
  assign new_n2648_ = new_n2632_ & new_n2647_;
  assign new_n2649_ = new_n2635_ & new_n2648_;
  assign new_n2650_ = new_n2638_ & new_n2649_;
  assign new_n2651_ = ~new_n2635_ & new_n2648_;
  assign new_n2652_ = new_n2638_ & new_n2651_;
  assign new_n2653_ = ~new_n2632_ & new_n2647_;
  assign new_n2654_ = new_n2635_ & new_n2653_;
  assign new_n2655_ = new_n2638_ & new_n2654_;
  assign new_n2656_ = new_n2623_ & ~new_n2626_;
  assign new_n2657_ = new_n2629_ & new_n2656_;
  assign new_n2658_ = ~new_n2632_ & new_n2657_;
  assign new_n2659_ = ~new_n2635_ & new_n2658_;
  assign new_n2660_ = new_n2638_ & new_n2659_;
  assign new_n2661_ = ~new_n2629_ & new_n2656_;
  assign new_n2662_ = new_n2632_ & new_n2661_;
  assign new_n2663_ = new_n2635_ & new_n2662_;
  assign new_n2664_ = new_n2638_ & new_n2663_;
  assign new_n2665_ = ~new_n2635_ & new_n2641_;
  assign new_n2666_ = ~new_n2638_ & new_n2665_;
  assign new_n2667_ = ~new_n2638_ & new_n2649_;
  assign new_n2668_ = ~new_n2638_ & new_n2654_;
  assign new_n2669_ = ~new_n2635_ & new_n2653_;
  assign new_n2670_ = ~new_n2638_ & new_n2669_;
  assign new_n2671_ = ~new_n2638_ & new_n2659_;
  assign new_n2672_ = ~new_n2635_ & new_n2662_;
  assign new_n2673_ = ~new_n2638_ & new_n2672_;
  assign new_n2674_ = ~new_n2632_ & new_n2661_;
  assign new_n2675_ = new_n2635_ & new_n2674_;
  assign new_n2676_ = ~new_n2638_ & new_n2675_;
  assign new_n2677_ = ~new_n2623_ & new_n2626_;
  assign new_n2678_ = new_n2629_ & new_n2677_;
  assign new_n2679_ = new_n2632_ & new_n2678_;
  assign new_n2680_ = ~new_n2635_ & new_n2679_;
  assign new_n2681_ = new_n2638_ & new_n2680_;
  assign new_n2682_ = ~new_n2629_ & new_n2677_;
  assign new_n2683_ = new_n2632_ & new_n2682_;
  assign new_n2684_ = ~new_n2635_ & new_n2683_;
  assign new_n2685_ = new_n2638_ & new_n2684_;
  assign new_n2686_ = ~new_n2632_ & new_n2682_;
  assign new_n2687_ = new_n2635_ & new_n2686_;
  assign new_n2688_ = new_n2638_ & new_n2687_;
  assign new_n2689_ = ~new_n2623_ & ~new_n2626_;
  assign new_n2690_ = new_n2629_ & new_n2689_;
  assign new_n2691_ = new_n2632_ & new_n2690_;
  assign new_n2692_ = new_n2635_ & new_n2691_;
  assign new_n2693_ = new_n2638_ & new_n2692_;
  assign new_n2694_ = ~new_n2629_ & new_n2689_;
  assign new_n2695_ = new_n2632_ & new_n2694_;
  assign new_n2696_ = ~new_n2635_ & new_n2695_;
  assign new_n2697_ = new_n2638_ & new_n2696_;
  assign new_n2698_ = ~new_n2632_ & new_n2694_;
  assign new_n2699_ = new_n2635_ & new_n2698_;
  assign new_n2700_ = new_n2638_ & new_n2699_;
  assign new_n2701_ = ~new_n2635_ & new_n2698_;
  assign new_n2702_ = new_n2638_ & new_n2701_;
  assign new_n2703_ = ~new_n2638_ & new_n2680_;
  assign new_n2704_ = new_n2635_ & new_n2683_;
  assign new_n2705_ = ~new_n2638_ & new_n2704_;
  assign new_n2706_ = ~new_n2635_ & new_n2686_;
  assign new_n2707_ = ~new_n2638_ & new_n2706_;
  assign new_n2708_ = ~new_n2635_ & new_n2691_;
  assign new_n2709_ = ~new_n2638_ & new_n2708_;
  assign new_n2710_ = ~new_n2632_ & new_n2690_;
  assign new_n2711_ = new_n2635_ & new_n2710_;
  assign new_n2712_ = ~new_n2638_ & new_n2711_;
  assign new_n2713_ = ~new_n2635_ & new_n2710_;
  assign new_n2714_ = ~new_n2638_ & new_n2713_;
  assign new_n2715_ = new_n2635_ & new_n2695_;
  assign new_n2716_ = ~new_n2638_ & new_n2715_;
  assign new_n2717_ = ~new_n2646_ & ~new_n2650_;
  assign new_n2718_ = ~new_n2643_ & new_n2717_;
  assign new_n2719_ = ~new_n2652_ & ~new_n2655_;
  assign new_n2720_ = ~new_n2660_ & ~new_n2664_;
  assign new_n2721_ = new_n2719_ & new_n2720_;
  assign new_n2722_ = new_n2718_ & new_n2721_;
  assign new_n2723_ = ~new_n2667_ & ~new_n2668_;
  assign new_n2724_ = ~new_n2666_ & new_n2723_;
  assign new_n2725_ = ~new_n2670_ & ~new_n2671_;
  assign new_n2726_ = ~new_n2673_ & ~new_n2676_;
  assign new_n2727_ = new_n2725_ & new_n2726_;
  assign new_n2728_ = new_n2724_ & new_n2727_;
  assign new_n2729_ = new_n2722_ & new_n2728_;
  assign new_n2730_ = ~new_n2685_ & ~new_n2688_;
  assign new_n2731_ = ~new_n2681_ & new_n2730_;
  assign new_n2732_ = ~new_n2693_ & ~new_n2697_;
  assign new_n2733_ = ~new_n2700_ & ~new_n2702_;
  assign new_n2734_ = new_n2732_ & new_n2733_;
  assign new_n2735_ = new_n2731_ & new_n2734_;
  assign new_n2736_ = ~new_n2705_ & ~new_n2707_;
  assign new_n2737_ = ~new_n2703_ & new_n2736_;
  assign new_n2738_ = ~new_n2709_ & ~new_n2712_;
  assign new_n2739_ = ~new_n2714_ & ~new_n2716_;
  assign new_n2740_ = new_n2738_ & new_n2739_;
  assign new_n2741_ = new_n2737_ & new_n2740_;
  assign new_n2742_ = new_n2735_ & new_n2741_;
  assign new_n2743_ = new_n2729_ & new_n2742_;
  assign new_n2744_ = ~new_n2629_ & ~new_n2638_;
  assign new_n2745_ = new_n2629_ & new_n2638_;
  assign new_n2746_ = ~new_n2744_ & ~new_n2745_;
  assign new_n2747_ = ~new_n2623_ & ~new_n2746_;
  assign new_n2748_ = ~new_n2629_ & new_n2638_;
  assign new_n2749_ = new_n2623_ & new_n2748_;
  assign new_n2750_ = ~new_n2747_ & ~new_n2749_;
  assign new_n2751_ = ~new_n2632_ & ~new_n2750_;
  assign new_n2752_ = new_n2632_ & ~new_n2638_;
  assign new_n2753_ = new_n2623_ & new_n2629_;
  assign new_n2754_ = new_n2752_ & new_n2753_;
  assign new_n2755_ = ~new_n2751_ & ~new_n2754_;
  assign new_n2756_ = new_n2635_ & ~new_n2755_;
  assign new_n2757_ = ~new_n2626_ & new_n2756_;
  assign new_n2758_ = new_n2743_ & ~new_n2757_;
  assign new_n2759_ = ~\data<29>  & ~new_n2758_;
  assign new_n2760_ = \data<29>  & new_n2758_;
  assign new_n2761_ = ~new_n2759_ & ~new_n2760_;
  assign new_n2762_ = new_n504_ & ~new_n2761_;
  assign new_n2763_ = \outreg<23>  & ~\count<0> ;
  assign new_n2764_ = \outreg<31>  & \count<0> ;
  assign new_n2765_ = ~new_n2763_ & ~new_n2764_;
  assign new_n2766_ = ~new_n504_ & ~new_n2765_;
  assign \outreg_new<23>  = new_n2762_ | new_n2766_;
  assign new_n2768_ = \data<61>  & new_n504_;
  assign new_n2769_ = \outreg<22>  & ~\count<0> ;
  assign new_n2770_ = \outreg<30>  & \count<0> ;
  assign new_n2771_ = ~new_n2769_ & ~new_n2770_;
  assign new_n2772_ = ~new_n504_ & ~new_n2771_;
  assign \outreg_new<22>  = new_n2768_ | new_n2772_;
  assign new_n2774_ = ~new_n2188_ & new_n2219_;
  assign new_n2775_ = new_n2191_ & new_n2774_;
  assign new_n2776_ = new_n2191_ & new_n2223_;
  assign new_n2777_ = new_n2191_ & new_n2228_;
  assign new_n2778_ = new_n2188_ & new_n2194_;
  assign new_n2779_ = ~new_n2191_ & new_n2778_;
  assign new_n2780_ = ~new_n2191_ & new_n2202_;
  assign new_n2781_ = ~new_n2191_ & new_n2207_;
  assign new_n2782_ = new_n2191_ & new_n2261_;
  assign new_n2783_ = ~new_n2188_ & new_n2238_;
  assign new_n2784_ = new_n2191_ & new_n2783_;
  assign new_n2785_ = new_n2188_ & new_n2248_;
  assign new_n2786_ = new_n2191_ & new_n2785_;
  assign new_n2787_ = ~new_n2188_ & new_n2258_;
  assign new_n2788_ = ~new_n2191_ & new_n2787_;
  assign new_n2789_ = ~new_n2191_ & new_n2242_;
  assign new_n2790_ = new_n2188_ & new_n2269_;
  assign new_n2791_ = ~new_n2191_ & new_n2790_;
  assign new_n2792_ = new_n2185_ & ~new_n2191_;
  assign new_n2793_ = ~new_n2185_ & new_n2191_;
  assign new_n2794_ = ~new_n2792_ & ~new_n2793_;
  assign new_n2795_ = ~new_n2188_ & ~new_n2794_;
  assign new_n2796_ = ~new_n2176_ & new_n2795_;
  assign new_n2797_ = new_n2188_ & ~new_n2191_;
  assign new_n2798_ = new_n2176_ & new_n2185_;
  assign new_n2799_ = new_n2797_ & new_n2798_;
  assign new_n2800_ = ~new_n2796_ & ~new_n2799_;
  assign new_n2801_ = ~new_n2182_ & ~new_n2800_;
  assign new_n2802_ = ~new_n2179_ & new_n2801_;
  assign new_n2803_ = ~new_n2196_ & ~new_n2200_;
  assign new_n2804_ = ~new_n2775_ & new_n2803_;
  assign new_n2805_ = ~new_n2211_ & ~new_n2776_;
  assign new_n2806_ = ~new_n2218_ & ~new_n2777_;
  assign new_n2807_ = new_n2805_ & new_n2806_;
  assign new_n2808_ = new_n2804_ & new_n2807_;
  assign new_n2809_ = ~new_n2222_ & ~new_n2780_;
  assign new_n2810_ = ~new_n2779_ & new_n2809_;
  assign new_n2811_ = ~new_n2224_ & ~new_n2781_;
  assign new_n2812_ = new_n2281_ & new_n2811_;
  assign new_n2813_ = new_n2810_ & new_n2812_;
  assign new_n2814_ = new_n2808_ & new_n2813_;
  assign new_n2815_ = ~new_n2243_ & ~new_n2784_;
  assign new_n2816_ = ~new_n2782_ & new_n2815_;
  assign new_n2817_ = ~new_n2245_ & ~new_n2786_;
  assign new_n2818_ = ~new_n2250_ & ~new_n2253_;
  assign new_n2819_ = new_n2817_ & new_n2818_;
  assign new_n2820_ = new_n2816_ & new_n2819_;
  assign new_n2821_ = ~new_n2260_ & ~new_n2788_;
  assign new_n2822_ = ~new_n2263_ & ~new_n2789_;
  assign new_n2823_ = new_n2821_ & new_n2822_;
  assign new_n2824_ = ~new_n2266_ & ~new_n2268_;
  assign new_n2825_ = new_n2179_ & new_n2182_;
  assign new_n2826_ = new_n2176_ & new_n2825_;
  assign new_n2827_ = new_n2188_ & new_n2191_;
  assign new_n2828_ = ~new_n2185_ & new_n2827_;
  assign new_n2829_ = new_n2826_ & new_n2828_;
  assign new_n2830_ = ~new_n2791_ & ~new_n2829_;
  assign new_n2831_ = new_n2824_ & new_n2830_;
  assign new_n2832_ = new_n2823_ & new_n2831_;
  assign new_n2833_ = new_n2820_ & new_n2832_;
  assign new_n2834_ = new_n2814_ & new_n2833_;
  assign new_n2835_ = ~new_n2802_ & new_n2834_;
  assign new_n2836_ = ~\data<21>  & ~new_n2835_;
  assign new_n2837_ = \data<21>  & new_n2835_;
  assign new_n2838_ = ~new_n2836_ & ~new_n2837_;
  assign new_n2839_ = new_n504_ & ~new_n2838_;
  assign new_n2840_ = \outreg<21>  & ~\count<0> ;
  assign new_n2841_ = \outreg<29>  & \count<0> ;
  assign new_n2842_ = ~new_n2840_ & ~new_n2841_;
  assign new_n2843_ = ~new_n504_ & ~new_n2842_;
  assign \outreg_new<21>  = new_n2839_ | new_n2843_;
  assign new_n2845_ = \data<53>  & new_n504_;
  assign new_n2846_ = \outreg<20>  & ~\count<0> ;
  assign new_n2847_ = \outreg<28>  & \count<0> ;
  assign new_n2848_ = ~new_n2846_ & ~new_n2847_;
  assign new_n2849_ = ~new_n504_ & ~new_n2848_;
  assign \outreg_new<20>  = new_n2845_ | new_n2849_;
  assign new_n2851_ = new_n746_ & new_n774_;
  assign new_n2852_ = ~new_n740_ & new_n770_;
  assign new_n2853_ = ~new_n743_ & new_n2852_;
  assign new_n2854_ = ~new_n746_ & new_n2853_;
  assign new_n2855_ = new_n743_ & new_n2001_;
  assign new_n2856_ = new_n746_ & new_n2855_;
  assign new_n2857_ = new_n743_ & new_n786_;
  assign new_n2858_ = ~new_n746_ & new_n2857_;
  assign new_n2859_ = ~new_n751_ & ~new_n758_;
  assign new_n2860_ = ~new_n2851_ & new_n2859_;
  assign new_n2861_ = ~new_n765_ & ~new_n1991_;
  assign new_n2862_ = ~new_n769_ & ~new_n1992_;
  assign new_n2863_ = new_n2861_ & new_n2862_;
  assign new_n2864_ = new_n2860_ & new_n2863_;
  assign new_n2865_ = ~new_n776_ & ~new_n2854_;
  assign new_n2866_ = ~new_n773_ & new_n2865_;
  assign new_n2867_ = ~new_n1994_ & ~new_n1996_;
  assign new_n2868_ = ~new_n777_ & ~new_n783_;
  assign new_n2869_ = new_n2867_ & new_n2868_;
  assign new_n2870_ = new_n2866_ & new_n2869_;
  assign new_n2871_ = new_n2864_ & new_n2870_;
  assign new_n2872_ = ~new_n795_ & ~new_n800_;
  assign new_n2873_ = ~new_n1999_ & new_n2872_;
  assign new_n2874_ = ~new_n2003_ & ~new_n2856_;
  assign new_n2875_ = ~new_n804_ & ~new_n809_;
  assign new_n2876_ = new_n2874_ & new_n2875_;
  assign new_n2877_ = new_n2873_ & new_n2876_;
  assign new_n2878_ = ~new_n813_ & ~new_n2858_;
  assign new_n2879_ = ~new_n815_ & ~new_n2005_;
  assign new_n2880_ = new_n2878_ & new_n2879_;
  assign new_n2881_ = new_n734_ & new_n737_;
  assign new_n2882_ = new_n731_ & new_n2881_;
  assign new_n2883_ = new_n743_ & new_n746_;
  assign new_n2884_ = ~new_n740_ & new_n2883_;
  assign new_n2885_ = new_n2882_ & new_n2884_;
  assign new_n2886_ = ~new_n2008_ & ~new_n2885_;
  assign new_n2887_ = new_n842_ & new_n2886_;
  assign new_n2888_ = new_n2880_ & new_n2887_;
  assign new_n2889_ = new_n2877_ & new_n2888_;
  assign new_n2890_ = new_n2871_ & new_n2889_;
  assign new_n2891_ = ~new_n734_ & ~new_n737_;
  assign new_n2892_ = ~new_n743_ & ~new_n746_;
  assign new_n2893_ = new_n2891_ & new_n2892_;
  assign new_n2894_ = new_n2881_ & new_n2883_;
  assign new_n2895_ = ~new_n2893_ & ~new_n2894_;
  assign new_n2896_ = ~new_n731_ & ~new_n2895_;
  assign new_n2897_ = ~new_n737_ & new_n848_;
  assign new_n2898_ = new_n747_ & new_n2897_;
  assign new_n2899_ = ~new_n2896_ & ~new_n2898_;
  assign new_n2900_ = new_n740_ & ~new_n2899_;
  assign new_n2901_ = new_n2890_ & ~new_n2900_;
  assign new_n2902_ = ~\data<13>  & ~new_n2901_;
  assign new_n2903_ = \data<13>  & new_n2901_;
  assign new_n2904_ = ~new_n2902_ & ~new_n2903_;
  assign new_n2905_ = new_n504_ & ~new_n2904_;
  assign new_n2906_ = \outreg<19>  & ~\count<0> ;
  assign new_n2907_ = \outreg<27>  & \count<0> ;
  assign new_n2908_ = ~new_n2906_ & ~new_n2907_;
  assign new_n2909_ = ~new_n504_ & ~new_n2908_;
  assign \outreg_new<19>  = new_n2905_ | new_n2909_;
  assign new_n2911_ = \data<45>  & new_n504_;
  assign new_n2912_ = \outreg<18>  & ~\count<0> ;
  assign new_n2913_ = \outreg<26>  & \count<0> ;
  assign new_n2914_ = ~new_n2912_ & ~new_n2913_;
  assign new_n2915_ = ~new_n504_ & ~new_n2914_;
  assign \outreg_new<18>  = new_n2911_ | new_n2915_;
  assign new_n2917_ = new_n2635_ & new_n2644_;
  assign new_n2918_ = new_n2638_ & new_n2917_;
  assign new_n2919_ = new_n2638_ & new_n2669_;
  assign new_n2920_ = new_n2632_ & new_n2657_;
  assign new_n2921_ = ~new_n2635_ & new_n2920_;
  assign new_n2922_ = new_n2638_ & new_n2921_;
  assign new_n2923_ = ~new_n2638_ & new_n2642_;
  assign new_n2924_ = ~new_n2638_ & new_n2645_;
  assign new_n2925_ = new_n2635_ & new_n2658_;
  assign new_n2926_ = ~new_n2638_ & new_n2925_;
  assign new_n2927_ = new_n2635_ & new_n2679_;
  assign new_n2928_ = new_n2638_ & new_n2927_;
  assign new_n2929_ = ~new_n2632_ & new_n2678_;
  assign new_n2930_ = ~new_n2635_ & new_n2929_;
  assign new_n2931_ = new_n2638_ & new_n2930_;
  assign new_n2932_ = new_n2638_ & new_n2715_;
  assign new_n2933_ = new_n2635_ & new_n2929_;
  assign new_n2934_ = ~new_n2638_ & new_n2933_;
  assign new_n2935_ = ~new_n2638_ & new_n2684_;
  assign new_n2936_ = ~new_n2638_ & new_n2696_;
  assign new_n2937_ = new_n2719_ & ~new_n2918_;
  assign new_n2938_ = ~new_n2919_ & ~new_n2922_;
  assign new_n2939_ = new_n2720_ & new_n2938_;
  assign new_n2940_ = new_n2937_ & new_n2939_;
  assign new_n2941_ = ~new_n2666_ & ~new_n2924_;
  assign new_n2942_ = ~new_n2923_ & new_n2941_;
  assign new_n2943_ = ~new_n2667_ & ~new_n2926_;
  assign new_n2944_ = new_n2726_ & new_n2943_;
  assign new_n2945_ = new_n2942_ & new_n2944_;
  assign new_n2946_ = new_n2940_ & new_n2945_;
  assign new_n2947_ = ~new_n2685_ & ~new_n2931_;
  assign new_n2948_ = ~new_n2928_ & new_n2947_;
  assign new_n2949_ = ~new_n2688_ & ~new_n2693_;
  assign new_n2950_ = ~new_n2702_ & ~new_n2932_;
  assign new_n2951_ = new_n2949_ & new_n2950_;
  assign new_n2952_ = new_n2948_ & new_n2951_;
  assign new_n2953_ = ~new_n2934_ & ~new_n2935_;
  assign new_n2954_ = ~new_n2707_ & ~new_n2709_;
  assign new_n2955_ = new_n2953_ & new_n2954_;
  assign new_n2956_ = ~new_n2626_ & ~new_n2629_;
  assign new_n2957_ = new_n2623_ & new_n2956_;
  assign new_n2958_ = ~new_n2635_ & ~new_n2638_;
  assign new_n2959_ = ~new_n2632_ & new_n2958_;
  assign new_n2960_ = new_n2957_ & new_n2959_;
  assign new_n2961_ = ~new_n2936_ & ~new_n2960_;
  assign new_n2962_ = new_n2739_ & new_n2961_;
  assign new_n2963_ = new_n2955_ & new_n2962_;
  assign new_n2964_ = new_n2952_ & new_n2963_;
  assign new_n2965_ = new_n2946_ & new_n2964_;
  assign new_n2966_ = new_n2635_ & ~new_n2638_;
  assign new_n2967_ = new_n2626_ & new_n2966_;
  assign new_n2968_ = ~new_n2635_ & new_n2638_;
  assign new_n2969_ = ~new_n2626_ & new_n2968_;
  assign new_n2970_ = ~new_n2967_ & ~new_n2969_;
  assign new_n2971_ = ~new_n2623_ & ~new_n2970_;
  assign new_n2972_ = new_n2635_ & new_n2638_;
  assign new_n2973_ = new_n2656_ & new_n2972_;
  assign new_n2974_ = ~new_n2971_ & ~new_n2973_;
  assign new_n2975_ = new_n2632_ & ~new_n2974_;
  assign new_n2976_ = new_n2629_ & new_n2975_;
  assign new_n2977_ = new_n2965_ & ~new_n2976_;
  assign new_n2978_ = ~\data<5>  & ~new_n2977_;
  assign new_n2979_ = \data<5>  & new_n2977_;
  assign new_n2980_ = ~new_n2978_ & ~new_n2979_;
  assign new_n2981_ = new_n504_ & ~new_n2980_;
  assign new_n2982_ = \outreg<17>  & ~\count<0> ;
  assign new_n2983_ = \outreg<25>  & \count<0> ;
  assign new_n2984_ = ~new_n2982_ & ~new_n2983_;
  assign new_n2985_ = ~new_n504_ & ~new_n2984_;
  assign \outreg_new<17>  = new_n2981_ | new_n2985_;
  assign new_n2987_ = \data<37>  & new_n504_;
  assign new_n2988_ = \outreg<16>  & ~\count<0> ;
  assign new_n2989_ = \outreg<24>  & \count<0> ;
  assign new_n2990_ = ~new_n2988_ & ~new_n2989_;
  assign new_n2991_ = ~new_n504_ & ~new_n2990_;
  assign \outreg_new<16>  = new_n2987_ | new_n2991_;
  assign new_n2993_ = new_n890_ & new_n910_;
  assign new_n2994_ = ~new_n893_ & new_n2993_;
  assign new_n2995_ = new_n893_ & new_n1039_;
  assign new_n2996_ = ~new_n893_ & new_n1032_;
  assign new_n2997_ = new_n893_ & new_n1027_;
  assign new_n2998_ = ~new_n912_ & ~new_n1026_;
  assign new_n2999_ = ~new_n909_ & new_n2998_;
  assign new_n3000_ = ~new_n924_ & ~new_n1029_;
  assign new_n3001_ = new_n975_ & new_n3000_;
  assign new_n3002_ = new_n2999_ & new_n3001_;
  assign new_n3003_ = ~new_n930_ & ~new_n931_;
  assign new_n3004_ = ~new_n1030_ & new_n3003_;
  assign new_n3005_ = ~new_n940_ & ~new_n2994_;
  assign new_n3006_ = ~new_n947_ & ~new_n1031_;
  assign new_n3007_ = new_n3005_ & new_n3006_;
  assign new_n3008_ = new_n3004_ & new_n3007_;
  assign new_n3009_ = new_n3002_ & new_n3008_;
  assign new_n3010_ = ~new_n952_ & ~new_n2995_;
  assign new_n3011_ = ~new_n1033_ & new_n3010_;
  assign new_n3012_ = ~new_n964_ & ~new_n1037_;
  assign new_n3013_ = new_n988_ & new_n3012_;
  assign new_n3014_ = new_n3011_ & new_n3013_;
  assign new_n3015_ = ~new_n1038_ & ~new_n2996_;
  assign new_n3016_ = ~new_n965_ & new_n3015_;
  assign new_n3017_ = ~new_n968_ & ~new_n971_;
  assign new_n3018_ = ~new_n1041_ & ~new_n2997_;
  assign new_n3019_ = new_n3017_ & new_n3018_;
  assign new_n3020_ = new_n3016_ & new_n3019_;
  assign new_n3021_ = new_n3014_ & new_n3020_;
  assign new_n3022_ = new_n3009_ & new_n3021_;
  assign new_n3023_ = ~new_n890_ & ~new_n1001_;
  assign new_n3024_ = ~new_n887_ & new_n3023_;
  assign new_n3025_ = new_n878_ & new_n3024_;
  assign new_n3026_ = ~new_n884_ & ~new_n887_;
  assign new_n3027_ = new_n1068_ & new_n3026_;
  assign new_n3028_ = new_n884_ & new_n887_;
  assign new_n3029_ = new_n1004_ & new_n3028_;
  assign new_n3030_ = ~new_n3027_ & ~new_n3029_;
  assign new_n3031_ = ~new_n878_ & ~new_n3030_;
  assign new_n3032_ = ~new_n3025_ & ~new_n3031_;
  assign new_n3033_ = new_n881_ & ~new_n3032_;
  assign new_n3034_ = new_n3022_ & ~new_n3033_;
  assign new_n3035_ = ~\data<30>  & ~new_n3034_;
  assign new_n3036_ = \data<30>  & new_n3034_;
  assign new_n3037_ = ~new_n3035_ & ~new_n3036_;
  assign new_n3038_ = new_n504_ & ~new_n3037_;
  assign new_n3039_ = \outreg<15>  & ~\count<0> ;
  assign new_n3040_ = \outreg<23>  & \count<0> ;
  assign new_n3041_ = ~new_n3039_ & ~new_n3040_;
  assign new_n3042_ = ~new_n504_ & ~new_n3041_;
  assign \outreg_new<15>  = new_n3038_ | new_n3042_;
  assign new_n3044_ = \data<62>  & new_n504_;
  assign new_n3045_ = \outreg<14>  & ~\count<0> ;
  assign new_n3046_ = \outreg<22>  & \count<0> ;
  assign new_n3047_ = ~new_n3045_ & ~new_n3046_;
  assign new_n3048_ = ~new_n504_ & ~new_n3047_;
  assign \outreg_new<14>  = new_n3044_ | new_n3048_;
  assign new_n3050_ = ~new_n903_ & ~new_n912_;
  assign new_n3051_ = ~new_n898_ & new_n3050_;
  assign new_n3052_ = ~new_n921_ & ~new_n1028_;
  assign new_n3053_ = new_n975_ & new_n3052_;
  assign new_n3054_ = new_n3051_ & new_n3053_;
  assign new_n3055_ = ~new_n1029_ & ~new_n2994_;
  assign new_n3056_ = ~new_n927_ & new_n3055_;
  assign new_n3057_ = ~new_n936_ & ~new_n942_;
  assign new_n3058_ = new_n3006_ & new_n3057_;
  assign new_n3059_ = new_n3056_ & new_n3058_;
  assign new_n3060_ = new_n3054_ & new_n3059_;
  assign new_n3061_ = ~new_n1036_ & ~new_n2995_;
  assign new_n3062_ = ~new_n952_ & new_n3061_;
  assign new_n3063_ = ~new_n959_ & ~new_n964_;
  assign new_n3064_ = new_n3015_ & new_n3063_;
  assign new_n3065_ = new_n3062_ & new_n3064_;
  assign new_n3066_ = ~new_n968_ & ~new_n1040_;
  assign new_n3067_ = ~new_n966_ & new_n3066_;
  assign new_n3068_ = ~new_n969_ & ~new_n1041_;
  assign new_n3069_ = ~new_n1042_ & ~new_n2997_;
  assign new_n3070_ = new_n3068_ & new_n3069_;
  assign new_n3071_ = new_n3067_ & new_n3070_;
  assign new_n3072_ = new_n3065_ & new_n3071_;
  assign new_n3073_ = new_n3060_ & new_n3072_;
  assign new_n3074_ = new_n884_ & new_n1009_;
  assign new_n3075_ = new_n890_ & new_n893_;
  assign new_n3076_ = ~new_n884_ & new_n3075_;
  assign new_n3077_ = ~new_n3074_ & ~new_n3076_;
  assign new_n3078_ = ~new_n887_ & ~new_n3077_;
  assign new_n3079_ = ~new_n878_ & new_n3078_;
  assign new_n3080_ = ~new_n1009_ & ~new_n3075_;
  assign new_n3081_ = new_n887_ & ~new_n3080_;
  assign new_n3082_ = ~new_n884_ & new_n3081_;
  assign new_n3083_ = new_n878_ & new_n3082_;
  assign new_n3084_ = ~new_n3079_ & ~new_n3083_;
  assign new_n3085_ = new_n881_ & ~new_n3084_;
  assign new_n3086_ = new_n3073_ & ~new_n3085_;
  assign new_n3087_ = ~\data<22>  & ~new_n3086_;
  assign new_n3088_ = \data<22>  & new_n3086_;
  assign new_n3089_ = ~new_n3087_ & ~new_n3088_;
  assign new_n3090_ = new_n504_ & ~new_n3089_;
  assign new_n3091_ = \outreg<13>  & ~\count<0> ;
  assign new_n3092_ = \outreg<21>  & \count<0> ;
  assign new_n3093_ = ~new_n3091_ & ~new_n3092_;
  assign new_n3094_ = ~new_n504_ & ~new_n3093_;
  assign \outreg_new<13>  = new_n3090_ | new_n3094_;
  assign new_n3096_ = \data<54>  & new_n504_;
  assign new_n3097_ = \outreg<12>  & ~\count<0> ;
  assign new_n3098_ = \outreg<20>  & \count<0> ;
  assign new_n3099_ = ~new_n3097_ & ~new_n3098_;
  assign new_n3100_ = ~new_n504_ & ~new_n3099_;
  assign \outreg_new<12>  = new_n3096_ | new_n3100_;
  assign new_n3102_ = new_n1614_ & new_n1617_;
  assign new_n3103_ = new_n2484_ & new_n3102_;
  assign new_n3104_ = ~new_n1614_ & ~new_n1617_;
  assign new_n3105_ = new_n2490_ & new_n3104_;
  assign new_n3106_ = ~new_n3103_ & ~new_n3105_;
  assign new_n3107_ = ~new_n1608_ & ~new_n3106_;
  assign new_n3108_ = new_n1608_ & new_n1614_;
  assign new_n3109_ = new_n1617_ & new_n2490_;
  assign new_n3110_ = new_n3108_ & new_n3109_;
  assign new_n3111_ = ~new_n3107_ & ~new_n3110_;
  assign new_n3112_ = new_n1611_ & ~new_n3111_;
  assign new_n3113_ = ~new_n1632_ & new_n2454_;
  assign new_n3114_ = ~new_n2440_ & ~new_n2565_;
  assign new_n3115_ = ~new_n1639_ & ~new_n1648_;
  assign new_n3116_ = new_n3114_ & new_n3115_;
  assign new_n3117_ = new_n3113_ & new_n3116_;
  assign new_n3118_ = ~new_n2441_ & ~new_n2566_;
  assign new_n3119_ = ~new_n1650_ & new_n3118_;
  assign new_n3120_ = ~new_n1656_ & ~new_n1663_;
  assign new_n3121_ = ~new_n1665_ & ~new_n2442_;
  assign new_n3122_ = new_n3120_ & new_n3121_;
  assign new_n3123_ = new_n3119_ & new_n3122_;
  assign new_n3124_ = new_n3117_ & new_n3123_;
  assign new_n3125_ = ~new_n1677_ & ~new_n2445_;
  assign new_n3126_ = ~new_n1670_ & new_n3125_;
  assign new_n3127_ = ~new_n1682_ & ~new_n2567_;
  assign new_n3128_ = ~new_n1689_ & ~new_n2448_;
  assign new_n3129_ = new_n3127_ & new_n3128_;
  assign new_n3130_ = new_n3126_ & new_n3129_;
  assign new_n3131_ = ~new_n1695_ & ~new_n1697_;
  assign new_n3132_ = ~new_n1701_ & ~new_n2568_;
  assign new_n3133_ = new_n3131_ & new_n3132_;
  assign new_n3134_ = ~new_n1705_ & ~new_n2451_;
  assign new_n3135_ = ~new_n1611_ & ~new_n1614_;
  assign new_n3136_ = new_n1608_ & new_n3135_;
  assign new_n3137_ = ~new_n1617_ & new_n2597_;
  assign new_n3138_ = new_n3136_ & new_n3137_;
  assign new_n3139_ = ~new_n2453_ & ~new_n3138_;
  assign new_n3140_ = new_n3134_ & new_n3139_;
  assign new_n3141_ = new_n3133_ & new_n3140_;
  assign new_n3142_ = new_n3130_ & new_n3141_;
  assign new_n3143_ = new_n3124_ & new_n3142_;
  assign new_n3144_ = ~new_n3112_ & new_n3143_;
  assign new_n3145_ = ~\data<14>  & ~new_n3144_;
  assign new_n3146_ = \data<14>  & new_n3144_;
  assign new_n3147_ = ~new_n3145_ & ~new_n3146_;
  assign new_n3148_ = new_n504_ & ~new_n3147_;
  assign new_n3149_ = \outreg<11>  & ~\count<0> ;
  assign new_n3150_ = \outreg<19>  & \count<0> ;
  assign new_n3151_ = ~new_n3149_ & ~new_n3150_;
  assign new_n3152_ = ~new_n504_ & ~new_n3151_;
  assign \outreg_new<11>  = new_n3148_ | new_n3152_;
  assign new_n3154_ = \data<46>  & new_n504_;
  assign new_n3155_ = \outreg<10>  & ~\count<0> ;
  assign new_n3156_ = \outreg<18>  & \count<0> ;
  assign new_n3157_ = ~new_n3155_ & ~new_n3156_;
  assign new_n3158_ = ~new_n504_ & ~new_n3157_;
  assign \outreg_new<10>  = new_n3154_ | new_n3158_;
  assign new_n3160_ = new_n2191_ & new_n2225_;
  assign new_n3161_ = ~new_n2188_ & new_n2198_;
  assign new_n3162_ = ~new_n2191_ & new_n3161_;
  assign new_n3163_ = new_n2191_ & new_n2790_;
  assign new_n3164_ = ~new_n2191_ & new_n2785_;
  assign new_n3165_ = new_n2185_ & ~new_n2301_;
  assign new_n3166_ = ~new_n2176_ & new_n3165_;
  assign new_n3167_ = new_n2176_ & ~new_n2182_;
  assign new_n3168_ = ~new_n2185_ & ~new_n2191_;
  assign new_n3169_ = new_n3167_ & new_n3168_;
  assign new_n3170_ = ~new_n3166_ & ~new_n3169_;
  assign new_n3171_ = new_n2188_ & ~new_n3170_;
  assign new_n3172_ = new_n2179_ & new_n3171_;
  assign new_n3173_ = new_n2272_ & ~new_n2775_;
  assign new_n3174_ = ~new_n2776_ & ~new_n3160_;
  assign new_n3175_ = ~new_n2211_ & ~new_n2215_;
  assign new_n3176_ = new_n3174_ & new_n3175_;
  assign new_n3177_ = new_n3173_ & new_n3176_;
  assign new_n3178_ = ~new_n2222_ & ~new_n2779_;
  assign new_n3179_ = ~new_n2221_ & new_n3178_;
  assign new_n3180_ = ~new_n2781_ & ~new_n3162_;
  assign new_n3181_ = ~new_n2226_ & ~new_n2229_;
  assign new_n3182_ = new_n3180_ & new_n3181_;
  assign new_n3183_ = new_n3179_ & new_n3182_;
  assign new_n3184_ = new_n3177_ & new_n3183_;
  assign new_n3185_ = ~new_n2236_ & ~new_n2784_;
  assign new_n3186_ = ~new_n2782_ & new_n3185_;
  assign new_n3187_ = ~new_n2243_ & ~new_n2250_;
  assign new_n3188_ = ~new_n2257_ & ~new_n3163_;
  assign new_n3189_ = new_n3187_ & new_n3188_;
  assign new_n3190_ = new_n3186_ & new_n3189_;
  assign new_n3191_ = ~new_n2262_ & ~new_n2788_;
  assign new_n3192_ = ~new_n2263_ & ~new_n3164_;
  assign new_n3193_ = new_n3191_ & new_n3192_;
  assign new_n3194_ = ~new_n2179_ & ~new_n2182_;
  assign new_n3195_ = new_n2176_ & new_n3194_;
  assign new_n3196_ = ~new_n2188_ & new_n2191_;
  assign new_n3197_ = ~new_n2185_ & new_n3196_;
  assign new_n3198_ = new_n3195_ & new_n3197_;
  assign new_n3199_ = ~new_n2791_ & ~new_n3198_;
  assign new_n3200_ = new_n2293_ & new_n3199_;
  assign new_n3201_ = new_n3193_ & new_n3200_;
  assign new_n3202_ = new_n3190_ & new_n3201_;
  assign new_n3203_ = new_n3184_ & new_n3202_;
  assign new_n3204_ = ~new_n3172_ & new_n3203_;
  assign new_n3205_ = ~\data<6>  & ~new_n3204_;
  assign new_n3206_ = \data<6>  & new_n3204_;
  assign new_n3207_ = ~new_n3205_ & ~new_n3206_;
  assign new_n3208_ = new_n504_ & ~new_n3207_;
  assign new_n3209_ = \outreg<17>  & \count<0> ;
  assign new_n3210_ = \outreg<9>  & ~\count<0> ;
  assign new_n3211_ = ~new_n3209_ & ~new_n3210_;
  assign new_n3212_ = ~new_n504_ & ~new_n3211_;
  assign \outreg_new<9>  = new_n3208_ | new_n3212_;
  assign new_n3214_ = \data<38>  & new_n504_;
  assign new_n3215_ = \outreg<16>  & \count<0> ;
  assign new_n3216_ = \outreg<8>  & ~\count<0> ;
  assign new_n3217_ = ~new_n3215_ & ~new_n3216_;
  assign new_n3218_ = ~new_n504_ & ~new_n3217_;
  assign \outreg_new<8>  = new_n3214_ | new_n3218_;
  assign new_n3220_ = ~new_n2203_ & ~new_n2208_;
  assign new_n3221_ = ~new_n2777_ & ~new_n3160_;
  assign new_n3222_ = new_n3220_ & new_n3221_;
  assign new_n3223_ = new_n2804_ & new_n3222_;
  assign new_n3224_ = ~new_n2779_ & ~new_n3162_;
  assign new_n3225_ = ~new_n2221_ & new_n3224_;
  assign new_n3226_ = ~new_n2224_ & ~new_n2780_;
  assign new_n3227_ = ~new_n2227_ & ~new_n2229_;
  assign new_n3228_ = new_n3226_ & new_n3227_;
  assign new_n3229_ = new_n3225_ & new_n3228_;
  assign new_n3230_ = new_n3223_ & new_n3229_;
  assign new_n3231_ = ~new_n2236_ & ~new_n2240_;
  assign new_n3232_ = ~new_n2782_ & new_n3231_;
  assign new_n3233_ = ~new_n2250_ & ~new_n3163_;
  assign new_n3234_ = new_n2817_ & new_n3233_;
  assign new_n3235_ = new_n3232_ & new_n3234_;
  assign new_n3236_ = ~new_n2262_ & ~new_n2789_;
  assign new_n3237_ = ~new_n2788_ & new_n3236_;
  assign new_n3238_ = ~new_n2266_ & ~new_n3164_;
  assign new_n3239_ = new_n2294_ & new_n3238_;
  assign new_n3240_ = new_n3237_ & new_n3239_;
  assign new_n3241_ = new_n3235_ & new_n3240_;
  assign new_n3242_ = new_n3230_ & new_n3241_;
  assign new_n3243_ = new_n2179_ & ~new_n2191_;
  assign new_n3244_ = ~new_n2179_ & new_n2191_;
  assign new_n3245_ = ~new_n3243_ & ~new_n3244_;
  assign new_n3246_ = ~new_n2188_ & ~new_n3245_;
  assign new_n3247_ = new_n2182_ & new_n3246_;
  assign new_n3248_ = ~new_n2176_ & new_n3247_;
  assign new_n3249_ = ~new_n2179_ & ~new_n2191_;
  assign new_n3250_ = new_n2179_ & new_n2191_;
  assign new_n3251_ = ~new_n3249_ & ~new_n3250_;
  assign new_n3252_ = new_n2188_ & ~new_n3251_;
  assign new_n3253_ = ~new_n2182_ & new_n3252_;
  assign new_n3254_ = new_n2176_ & new_n3253_;
  assign new_n3255_ = ~new_n3248_ & ~new_n3254_;
  assign new_n3256_ = ~new_n2185_ & ~new_n3255_;
  assign new_n3257_ = new_n3242_ & ~new_n3256_;
  assign new_n3258_ = ~\data<31>  & ~new_n3257_;
  assign new_n3259_ = \data<31>  & new_n3257_;
  assign new_n3260_ = ~new_n3258_ & ~new_n3259_;
  assign new_n3261_ = new_n504_ & ~new_n3260_;
  assign new_n3262_ = \outreg<15>  & \count<0> ;
  assign new_n3263_ = \outreg<7>  & ~\count<0> ;
  assign new_n3264_ = ~new_n3262_ & ~new_n3263_;
  assign new_n3265_ = ~new_n504_ & ~new_n3264_;
  assign \outreg_new<7>  = new_n3261_ | new_n3265_;
  assign new_n3267_ = \data<63>  & new_n504_;
  assign new_n3268_ = \outreg<14>  & \count<0> ;
  assign new_n3269_ = \outreg<6>  & ~\count<0> ;
  assign new_n3270_ = ~new_n3268_ & ~new_n3269_;
  assign new_n3271_ = ~new_n504_ & ~new_n3270_;
  assign \outreg_new<6>  = new_n3267_ | new_n3271_;
  assign new_n3273_ = new_n2638_ & new_n2925_;
  assign new_n3274_ = ~new_n2638_ & new_n2663_;
  assign new_n3275_ = new_n2638_ & new_n2713_;
  assign new_n3276_ = ~new_n2638_ & new_n2701_;
  assign new_n3277_ = ~new_n2646_ & ~new_n2918_;
  assign new_n3278_ = ~new_n2643_ & new_n3277_;
  assign new_n3279_ = ~new_n2655_ & ~new_n2922_;
  assign new_n3280_ = ~new_n2664_ & ~new_n3273_;
  assign new_n3281_ = new_n3279_ & new_n3280_;
  assign new_n3282_ = new_n3278_ & new_n3281_;
  assign new_n3283_ = ~new_n2670_ & ~new_n2924_;
  assign new_n3284_ = ~new_n2923_ & new_n3283_;
  assign new_n3285_ = ~new_n2671_ & ~new_n3274_;
  assign new_n3286_ = new_n2726_ & new_n3285_;
  assign new_n3287_ = new_n3284_ & new_n3286_;
  assign new_n3288_ = new_n3282_ & new_n3287_;
  assign new_n3289_ = ~new_n2693_ & ~new_n3275_;
  assign new_n3290_ = ~new_n2697_ & ~new_n2700_;
  assign new_n3291_ = new_n3289_ & new_n3290_;
  assign new_n3292_ = new_n2948_ & new_n3291_;
  assign new_n3293_ = ~new_n2703_ & ~new_n2934_;
  assign new_n3294_ = ~new_n2709_ & ~new_n2935_;
  assign new_n3295_ = new_n3293_ & new_n3294_;
  assign new_n3296_ = ~new_n2712_ & ~new_n2716_;
  assign new_n3297_ = new_n2632_ & new_n2958_;
  assign new_n3298_ = ~new_n2626_ & new_n2629_;
  assign new_n3299_ = new_n2623_ & new_n3298_;
  assign new_n3300_ = new_n3297_ & new_n3299_;
  assign new_n3301_ = ~new_n3276_ & ~new_n3300_;
  assign new_n3302_ = new_n3296_ & new_n3301_;
  assign new_n3303_ = new_n3295_ & new_n3302_;
  assign new_n3304_ = new_n3292_ & new_n3303_;
  assign new_n3305_ = new_n3288_ & new_n3304_;
  assign new_n3306_ = ~new_n2632_ & new_n2968_;
  assign new_n3307_ = new_n2656_ & new_n3306_;
  assign new_n3308_ = ~new_n2632_ & ~new_n2638_;
  assign new_n3309_ = new_n2632_ & new_n2638_;
  assign new_n3310_ = ~new_n3308_ & ~new_n3309_;
  assign new_n3311_ = new_n2635_ & ~new_n3310_;
  assign new_n3312_ = new_n2626_ & new_n3311_;
  assign new_n3313_ = ~new_n2623_ & new_n3312_;
  assign new_n3314_ = ~new_n3307_ & ~new_n3313_;
  assign new_n3315_ = ~new_n2629_ & ~new_n3314_;
  assign new_n3316_ = new_n3305_ & ~new_n3315_;
  assign new_n3317_ = ~\data<23>  & ~new_n3316_;
  assign new_n3318_ = \data<23>  & new_n3316_;
  assign new_n3319_ = ~new_n3317_ & ~new_n3318_;
  assign new_n3320_ = new_n504_ & ~new_n3319_;
  assign new_n3321_ = \outreg<13>  & \count<0> ;
  assign new_n3322_ = \outreg<5>  & ~\count<0> ;
  assign new_n3323_ = ~new_n3321_ & ~new_n3322_;
  assign new_n3324_ = ~new_n504_ & ~new_n3323_;
  assign \outreg_new<5>  = new_n3320_ | new_n3324_;
  assign new_n3326_ = \data<55>  & new_n504_;
  assign new_n3327_ = \outreg<12>  & \count<0> ;
  assign new_n3328_ = \outreg<4>  & ~\count<0> ;
  assign new_n3329_ = ~new_n3327_ & ~new_n3328_;
  assign new_n3330_ = ~new_n504_ & ~new_n3329_;
  assign \outreg_new<4>  = new_n3326_ | new_n3330_;
  assign new_n3332_ = ~new_n2626_ & new_n2752_;
  assign new_n3333_ = ~new_n2632_ & new_n2638_;
  assign new_n3334_ = new_n2626_ & new_n3333_;
  assign new_n3335_ = ~new_n3332_ & ~new_n3334_;
  assign new_n3336_ = new_n2635_ & ~new_n3335_;
  assign new_n3337_ = new_n2629_ & new_n3336_;
  assign new_n3338_ = ~new_n2623_ & new_n3337_;
  assign new_n3339_ = ~new_n2650_ & ~new_n2655_;
  assign new_n3340_ = ~new_n2646_ & new_n3339_;
  assign new_n3341_ = ~new_n2660_ & ~new_n3273_;
  assign new_n3342_ = new_n2938_ & new_n3341_;
  assign new_n3343_ = new_n3340_ & new_n3342_;
  assign new_n3344_ = ~new_n2666_ & ~new_n2668_;
  assign new_n3345_ = ~new_n2923_ & new_n3344_;
  assign new_n3346_ = ~new_n2671_ & ~new_n2926_;
  assign new_n3347_ = ~new_n2676_ & ~new_n3274_;
  assign new_n3348_ = new_n3346_ & new_n3347_;
  assign new_n3349_ = new_n3345_ & new_n3348_;
  assign new_n3350_ = new_n3343_ & new_n3349_;
  assign new_n3351_ = ~new_n2681_ & ~new_n2685_;
  assign new_n3352_ = ~new_n2928_ & new_n3351_;
  assign new_n3353_ = ~new_n2932_ & ~new_n3275_;
  assign new_n3354_ = new_n2733_ & new_n3353_;
  assign new_n3355_ = new_n3352_ & new_n3354_;
  assign new_n3356_ = new_n2736_ & ~new_n2934_;
  assign new_n3357_ = ~new_n2936_ & ~new_n3276_;
  assign new_n3358_ = new_n2738_ & new_n3357_;
  assign new_n3359_ = new_n3356_ & new_n3358_;
  assign new_n3360_ = new_n3355_ & new_n3359_;
  assign new_n3361_ = new_n3350_ & new_n3360_;
  assign new_n3362_ = new_n2626_ & ~new_n2638_;
  assign new_n3363_ = ~new_n2626_ & new_n2638_;
  assign new_n3364_ = ~new_n3362_ & ~new_n3363_;
  assign new_n3365_ = ~new_n2635_ & ~new_n3364_;
  assign new_n3366_ = new_n2632_ & new_n3365_;
  assign new_n3367_ = ~new_n2629_ & new_n3366_;
  assign new_n3368_ = new_n2623_ & new_n3367_;
  assign new_n3369_ = new_n3361_ & ~new_n3368_;
  assign new_n3370_ = ~new_n3338_ & new_n3369_;
  assign new_n3371_ = ~\data<15>  & ~new_n3370_;
  assign new_n3372_ = \data<15>  & new_n3370_;
  assign new_n3373_ = ~new_n3371_ & ~new_n3372_;
  assign new_n3374_ = new_n504_ & ~new_n3373_;
  assign new_n3375_ = \outreg<11>  & \count<0> ;
  assign new_n3376_ = \outreg<3>  & ~\count<0> ;
  assign new_n3377_ = ~new_n3375_ & ~new_n3376_;
  assign new_n3378_ = ~new_n504_ & ~new_n3377_;
  assign \outreg_new<3>  = new_n3374_ | new_n3378_;
  assign new_n3380_ = \data<47>  & new_n504_;
  assign new_n3381_ = \outreg<10>  & \count<0> ;
  assign new_n3382_ = \outreg<2>  & ~\count<0> ;
  assign new_n3383_ = ~new_n3381_ & ~new_n3382_;
  assign new_n3384_ = ~new_n504_ & ~new_n3383_;
  assign \outreg_new<2>  = new_n3380_ | new_n3384_;
  assign new_n3386_ = new_n737_ & new_n2009_;
  assign new_n3387_ = ~new_n737_ & new_n2011_;
  assign new_n3388_ = ~new_n3386_ & ~new_n3387_;
  assign new_n3389_ = ~new_n743_ & ~new_n3388_;
  assign new_n3390_ = new_n734_ & new_n3389_;
  assign new_n3391_ = ~new_n731_ & new_n3390_;
  assign new_n3392_ = new_n821_ & ~new_n2851_;
  assign new_n3393_ = ~new_n765_ & ~new_n1992_;
  assign new_n3394_ = ~new_n769_ & ~new_n1993_;
  assign new_n3395_ = new_n3393_ & new_n3394_;
  assign new_n3396_ = new_n3392_ & new_n3395_;
  assign new_n3397_ = ~new_n775_ & ~new_n2854_;
  assign new_n3398_ = ~new_n773_ & new_n3397_;
  assign new_n3399_ = ~new_n777_ & ~new_n1994_;
  assign new_n3400_ = ~new_n778_ & ~new_n1998_;
  assign new_n3401_ = new_n3399_ & new_n3400_;
  assign new_n3402_ = new_n3398_ & new_n3401_;
  assign new_n3403_ = new_n3396_ & new_n3402_;
  assign new_n3404_ = ~new_n792_ & ~new_n1999_;
  assign new_n3405_ = ~new_n788_ & new_n3404_;
  assign new_n3406_ = ~new_n809_ & ~new_n2856_;
  assign new_n3407_ = new_n2039_ & new_n3406_;
  assign new_n3408_ = new_n3405_ & new_n3407_;
  assign new_n3409_ = ~new_n815_ & ~new_n2858_;
  assign new_n3410_ = ~new_n812_ & new_n3409_;
  assign new_n3411_ = ~new_n818_ & ~new_n2005_;
  assign new_n3412_ = ~new_n819_ & ~new_n2006_;
  assign new_n3413_ = new_n3411_ & new_n3412_;
  assign new_n3414_ = new_n3410_ & new_n3413_;
  assign new_n3415_ = new_n3408_ & new_n3414_;
  assign new_n3416_ = new_n3403_ & new_n3415_;
  assign new_n3417_ = ~new_n737_ & new_n856_;
  assign new_n3418_ = new_n737_ & new_n857_;
  assign new_n3419_ = ~new_n3417_ & ~new_n3418_;
  assign new_n3420_ = new_n743_ & ~new_n3419_;
  assign new_n3421_ = ~new_n734_ & new_n3420_;
  assign new_n3422_ = new_n731_ & new_n3421_;
  assign new_n3423_ = new_n3416_ & ~new_n3422_;
  assign new_n3424_ = ~new_n3391_ & new_n3423_;
  assign new_n3425_ = ~\data<7>  & ~new_n3424_;
  assign new_n3426_ = \data<7>  & new_n3424_;
  assign new_n3427_ = ~new_n3425_ & ~new_n3426_;
  assign new_n3428_ = new_n504_ & ~new_n3427_;
  assign new_n3429_ = \outreg<1>  & ~\count<0> ;
  assign new_n3430_ = \outreg<9>  & \count<0> ;
  assign new_n3431_ = ~new_n3429_ & ~new_n3430_;
  assign new_n3432_ = ~new_n504_ & ~new_n3431_;
  assign \outreg_new<1>  = new_n3428_ | new_n3432_;
  assign new_n3434_ = \data<39>  & new_n504_;
  assign new_n3435_ = \outreg<0>  & ~\count<0> ;
  assign new_n3436_ = \outreg<8>  & \count<0> ;
  assign new_n3437_ = ~new_n3435_ & ~new_n3436_;
  assign new_n3438_ = ~new_n504_ & ~new_n3437_;
  assign \outreg_new<0>  = new_n3434_ | new_n3438_;
  assign new_n3440_ = ~new_n504_ & ~new_n3260_;
  assign new_n3441_ = \data_in<6>  & new_n504_;
  assign \data_new<63>  = new_n3440_ | new_n3441_;
  assign new_n3443_ = ~new_n504_ & ~new_n3037_;
  assign new_n3444_ = \inreg<6>  & new_n504_;
  assign \data_new<62>  = new_n3443_ | new_n3444_;
  assign new_n3446_ = ~new_n504_ & ~new_n2761_;
  assign new_n3447_ = \inreg<14>  & new_n504_;
  assign \data_new<61>  = new_n3446_ | new_n3447_;
  assign new_n3449_ = ~new_n504_ & ~new_n2425_;
  assign new_n3450_ = \inreg<22>  & new_n504_;
  assign \data_new<60>  = new_n3449_ | new_n3450_;
  assign new_n3452_ = ~new_n504_ & ~new_n2111_;
  assign new_n3453_ = \inreg<30>  & new_n504_;
  assign \data_new<59>  = new_n3452_ | new_n3453_;
  assign new_n3455_ = ~new_n504_ & ~new_n1751_;
  assign new_n3456_ = \inreg<38>  & new_n504_;
  assign \data_new<58>  = new_n3455_ | new_n3456_;
  assign new_n3458_ = ~new_n504_ & ~new_n1302_;
  assign new_n3459_ = \inreg<46>  & new_n504_;
  assign \data_new<57>  = new_n3458_ | new_n3459_;
  assign new_n3461_ = ~new_n504_ & ~new_n867_;
  assign new_n3462_ = \inreg<54>  & new_n504_;
  assign \data_new<56>  = new_n3461_ | new_n3462_;
  assign new_n3464_ = ~new_n504_ & ~new_n3319_;
  assign new_n3465_ = \data_in<4>  & new_n504_;
  assign \data_new<55>  = new_n3464_ | new_n3465_;
  assign new_n3467_ = ~new_n504_ & ~new_n3089_;
  assign new_n3468_ = \inreg<4>  & new_n504_;
  assign \data_new<54>  = new_n3467_ | new_n3468_;
  assign new_n3470_ = ~new_n504_ & ~new_n2838_;
  assign new_n3471_ = \inreg<12>  & new_n504_;
  assign \data_new<53>  = new_n3470_ | new_n3471_;
  assign new_n3473_ = ~new_n504_ & ~new_n2498_;
  assign new_n3474_ = \inreg<20>  & new_n504_;
  assign \data_new<52>  = new_n3473_ | new_n3474_;
  assign new_n3476_ = ~new_n504_ & ~new_n2161_;
  assign new_n3477_ = \inreg<28>  & new_n504_;
  assign \data_new<51>  = new_n3476_ | new_n3477_;
  assign new_n3479_ = ~new_n504_ & ~new_n1910_;
  assign new_n3480_ = \inreg<36>  & new_n504_;
  assign \data_new<50>  = new_n3479_ | new_n3480_;
  assign new_n3482_ = ~new_n504_ & ~new_n1459_;
  assign new_n3483_ = \inreg<44>  & new_n504_;
  assign \data_new<49>  = new_n3482_ | new_n3483_;
  assign new_n3485_ = ~new_n504_ & ~new_n1017_;
  assign new_n3486_ = \inreg<52>  & new_n504_;
  assign \data_new<48>  = new_n3485_ | new_n3486_;
  assign new_n3488_ = ~new_n504_ & ~new_n3373_;
  assign new_n3489_ = \data_in<2>  & new_n504_;
  assign \data_new<47>  = new_n3488_ | new_n3489_;
  assign new_n3491_ = ~new_n504_ & ~new_n3147_;
  assign new_n3492_ = \inreg<2>  & new_n504_;
  assign \data_new<46>  = new_n3491_ | new_n3492_;
  assign new_n3494_ = ~new_n504_ & ~new_n2904_;
  assign new_n3495_ = \inreg<10>  & new_n504_;
  assign \data_new<45>  = new_n3494_ | new_n3495_;
  assign new_n3497_ = ~new_n504_ & ~new_n2552_;
  assign new_n3498_ = \inreg<18>  & new_n504_;
  assign \data_new<44>  = new_n3497_ | new_n3498_;
  assign new_n3500_ = ~new_n504_ & ~new_n2311_;
  assign new_n3501_ = \inreg<26>  & new_n504_;
  assign \data_new<43>  = new_n3500_ | new_n3501_;
  assign new_n3503_ = ~new_n504_ & ~new_n1976_;
  assign new_n3504_ = \inreg<34>  & new_n504_;
  assign \data_new<42>  = new_n3503_ | new_n3504_;
  assign new_n3506_ = ~new_n504_ & ~new_n1517_;
  assign new_n3507_ = \inreg<42>  & new_n504_;
  assign \data_new<41>  = new_n3506_ | new_n3507_;
  assign new_n3509_ = ~new_n504_ & ~new_n1083_;
  assign new_n3510_ = \inreg<50>  & new_n504_;
  assign \data_new<40>  = new_n3509_ | new_n3510_;
  assign new_n3512_ = ~new_n504_ & ~new_n3427_;
  assign new_n3513_ = \data_in<0>  & new_n504_;
  assign \data_new<39>  = new_n3512_ | new_n3513_;
  assign new_n3515_ = ~new_n504_ & ~new_n3207_;
  assign new_n3516_ = \inreg<0>  & new_n504_;
  assign \data_new<38>  = new_n3515_ | new_n3516_;
  assign new_n3518_ = ~new_n504_ & ~new_n2980_;
  assign new_n3519_ = \inreg<8>  & new_n504_;
  assign \data_new<37>  = new_n3518_ | new_n3519_;
  assign new_n3521_ = ~new_n504_ & ~new_n2608_;
  assign new_n3522_ = \inreg<16>  & new_n504_;
  assign \data_new<36>  = new_n3521_ | new_n3522_;
  assign new_n3524_ = ~new_n504_ & ~new_n2372_;
  assign new_n3525_ = \inreg<24>  & new_n504_;
  assign \data_new<35>  = new_n3524_ | new_n3525_;
  assign new_n3527_ = ~new_n504_ & ~new_n2054_;
  assign new_n3528_ = \inreg<32>  & new_n504_;
  assign \data_new<34>  = new_n3527_ | new_n3528_;
  assign new_n3530_ = ~new_n504_ & ~new_n1593_;
  assign new_n3531_ = \inreg<40>  & new_n504_;
  assign \data_new<33>  = new_n3530_ | new_n3531_;
  assign new_n3533_ = ~new_n504_ & ~new_n1230_;
  assign new_n3534_ = \inreg<48>  & new_n504_;
  assign \data_new<32>  = new_n3533_ | new_n3534_;
  assign new_n3536_ = \data<63>  & ~new_n504_;
  assign new_n3537_ = \data_in<7>  & new_n504_;
  assign \data_new<31>  = new_n3536_ | new_n3537_;
  assign new_n3539_ = \data<62>  & ~new_n504_;
  assign new_n3540_ = \inreg<7>  & new_n504_;
  assign \data_new<30>  = new_n3539_ | new_n3540_;
  assign new_n3542_ = \data<61>  & ~new_n504_;
  assign new_n3543_ = \inreg<15>  & new_n504_;
  assign \data_new<29>  = new_n3542_ | new_n3543_;
  assign new_n3545_ = \data<60>  & ~new_n504_;
  assign new_n3546_ = \inreg<23>  & new_n504_;
  assign \data_new<28>  = new_n3545_ | new_n3546_;
  assign new_n3548_ = \data<59>  & ~new_n504_;
  assign new_n3549_ = \inreg<31>  & new_n504_;
  assign \data_new<27>  = new_n3548_ | new_n3549_;
  assign new_n3551_ = \data<58>  & ~new_n504_;
  assign new_n3552_ = \inreg<39>  & new_n504_;
  assign \data_new<26>  = new_n3551_ | new_n3552_;
  assign new_n3554_ = \data<57>  & ~new_n504_;
  assign new_n3555_ = \inreg<47>  & new_n504_;
  assign \data_new<25>  = new_n3554_ | new_n3555_;
  assign new_n3557_ = \data<56>  & ~new_n504_;
  assign new_n3558_ = \inreg<55>  & new_n504_;
  assign \data_new<24>  = new_n3557_ | new_n3558_;
  assign new_n3560_ = \data<55>  & ~new_n504_;
  assign new_n3561_ = \data_in<5>  & new_n504_;
  assign \data_new<23>  = new_n3560_ | new_n3561_;
  assign new_n3563_ = \data<54>  & ~new_n504_;
  assign new_n3564_ = \inreg<5>  & new_n504_;
  assign \data_new<22>  = new_n3563_ | new_n3564_;
  assign new_n3566_ = \data<53>  & ~new_n504_;
  assign new_n3567_ = \inreg<13>  & new_n504_;
  assign \data_new<21>  = new_n3566_ | new_n3567_;
  assign new_n3569_ = \data<52>  & ~new_n504_;
  assign new_n3570_ = \inreg<21>  & new_n504_;
  assign \data_new<20>  = new_n3569_ | new_n3570_;
  assign new_n3572_ = \data<51>  & ~new_n504_;
  assign new_n3573_ = \inreg<29>  & new_n504_;
  assign \data_new<19>  = new_n3572_ | new_n3573_;
  assign new_n3575_ = \data<50>  & ~new_n504_;
  assign new_n3576_ = \inreg<37>  & new_n504_;
  assign \data_new<18>  = new_n3575_ | new_n3576_;
  assign new_n3578_ = \data<49>  & ~new_n504_;
  assign new_n3579_ = \inreg<45>  & new_n504_;
  assign \data_new<17>  = new_n3578_ | new_n3579_;
  assign new_n3581_ = \data<48>  & ~new_n504_;
  assign new_n3582_ = \inreg<53>  & new_n504_;
  assign \data_new<16>  = new_n3581_ | new_n3582_;
  assign new_n3584_ = \data<47>  & ~new_n504_;
  assign new_n3585_ = \data_in<3>  & new_n504_;
  assign \data_new<15>  = new_n3584_ | new_n3585_;
  assign new_n3587_ = \data<46>  & ~new_n504_;
  assign new_n3588_ = \inreg<3>  & new_n504_;
  assign \data_new<14>  = new_n3587_ | new_n3588_;
  assign new_n3590_ = \data<45>  & ~new_n504_;
  assign new_n3591_ = \inreg<11>  & new_n504_;
  assign \data_new<13>  = new_n3590_ | new_n3591_;
  assign new_n3593_ = \data<44>  & ~new_n504_;
  assign new_n3594_ = \inreg<19>  & new_n504_;
  assign \data_new<12>  = new_n3593_ | new_n3594_;
  assign new_n3596_ = \data<43>  & ~new_n504_;
  assign new_n3597_ = \inreg<27>  & new_n504_;
  assign \data_new<11>  = new_n3596_ | new_n3597_;
  assign new_n3599_ = \data<42>  & ~new_n504_;
  assign new_n3600_ = \inreg<35>  & new_n504_;
  assign \data_new<10>  = new_n3599_ | new_n3600_;
  assign new_n3602_ = \data<41>  & ~new_n504_;
  assign new_n3603_ = \inreg<43>  & new_n504_;
  assign \data_new<9>  = new_n3602_ | new_n3603_;
  assign new_n3605_ = \data<40>  & ~new_n504_;
  assign new_n3606_ = \inreg<51>  & new_n504_;
  assign \data_new<8>  = new_n3605_ | new_n3606_;
  assign new_n3608_ = \data<39>  & ~new_n504_;
  assign new_n3609_ = \data_in<1>  & new_n504_;
  assign \data_new<7>  = new_n3608_ | new_n3609_;
  assign new_n3611_ = \data<38>  & ~new_n504_;
  assign new_n3612_ = \inreg<1>  & new_n504_;
  assign \data_new<6>  = new_n3611_ | new_n3612_;
  assign new_n3614_ = \data<37>  & ~new_n504_;
  assign new_n3615_ = \inreg<9>  & new_n504_;
  assign \data_new<5>  = new_n3614_ | new_n3615_;
  assign new_n3617_ = \data<36>  & ~new_n504_;
  assign new_n3618_ = \inreg<17>  & new_n504_;
  assign \data_new<4>  = new_n3617_ | new_n3618_;
  assign new_n3620_ = \data<35>  & ~new_n504_;
  assign new_n3621_ = \inreg<25>  & new_n504_;
  assign \data_new<3>  = new_n3620_ | new_n3621_;
  assign new_n3623_ = \data<34>  & ~new_n504_;
  assign new_n3624_ = \inreg<33>  & new_n504_;
  assign \data_new<2>  = new_n3623_ | new_n3624_;
  assign new_n3626_ = \data<33>  & ~new_n504_;
  assign new_n3627_ = \inreg<41>  & new_n504_;
  assign \data_new<1>  = new_n3626_ | new_n3627_;
  assign new_n3629_ = \data<32>  & ~new_n504_;
  assign new_n3630_ = \inreg<49>  & new_n504_;
  assign \data_new<0>  = new_n3629_ | new_n3630_;
  assign new_n3632_ = \load_key<0>  & new_n504_;
  assign new_n3633_ = \count<3>  & ~new_n503_;
  assign new_n3634_ = ~\count<3>  & \count<2> ;
  assign new_n3635_ = new_n502_ & new_n3634_;
  assign new_n3636_ = ~new_n3633_ & ~new_n3635_;
  assign new_n3637_ = ~\reset<0>  & ~new_n3636_;
  assign \count_new<3>  = ~new_n3632_ & new_n3637_;
  assign new_n3639_ = \count<2>  & ~new_n502_;
  assign new_n3640_ = ~\count<2>  & new_n502_;
  assign new_n3641_ = ~new_n3639_ & ~new_n3640_;
  assign new_n3642_ = ~\reset<0>  & ~new_n3641_;
  assign \count_new<2>  = ~new_n3632_ & new_n3642_;
  assign new_n3644_ = \count<1>  & ~\count<0> ;
  assign new_n3645_ = ~\count<1>  & \count<0> ;
  assign new_n3646_ = ~new_n3644_ & ~new_n3645_;
  assign new_n3647_ = ~\reset<0>  & ~new_n3646_;
  assign \count_new<1>  = ~new_n3632_ & new_n3647_;
  assign new_n3649_ = ~\reset<0>  & ~new_n3632_;
  assign \count_new<0>  = ~\count<0>  & new_n3649_;
  assign new_n3651_ = ~\encrypt<0>  & \encrypt_mode<0> ;
  assign new_n3652_ = \encrypt<0>  & ~\encrypt_mode<0> ;
  assign new_n3653_ = ~new_n3651_ & ~new_n3652_;
  assign new_n3654_ = \count<3>  & ~new_n3653_;
  assign new_n3655_ = \count<2>  & new_n3654_;
  assign new_n3656_ = \count<1>  & new_n3655_;
  assign new_n3657_ = \count<0>  & new_n3656_;
  assign new_n3658_ = \count<3>  & ~\count<0> ;
  assign new_n3659_ = ~\count<0>  & ~new_n3658_;
  assign new_n3660_ = \count<2>  & ~new_n3659_;
  assign new_n3661_ = \count<1>  & new_n3660_;
  assign new_n3662_ = ~\count<1>  & ~\count<0> ;
  assign new_n3663_ = ~\count<3>  & ~\count<2> ;
  assign new_n3664_ = new_n3662_ & new_n3663_;
  assign new_n3665_ = ~new_n3661_ & ~new_n3664_;
  assign new_n3666_ = ~\encrypt<0>  & \inreg<27> ;
  assign new_n3667_ = \encrypt<0>  & \inreg<48> ;
  assign new_n3668_ = ~new_n3666_ & ~new_n3667_;
  assign new_n3669_ = new_n3632_ & ~new_n3668_;
  assign new_n3670_ = \C<0>  & ~new_n3665_;
  assign new_n3671_ = \C<1>  & new_n3665_;
  assign new_n3672_ = ~new_n3670_ & ~new_n3671_;
  assign new_n3673_ = \encrypt_mode<0>  & ~new_n3672_;
  assign new_n3674_ = \C<26>  & ~new_n3665_;
  assign new_n3675_ = \C<25>  & new_n3665_;
  assign new_n3676_ = ~new_n3674_ & ~new_n3675_;
  assign new_n3677_ = ~\encrypt_mode<0>  & ~new_n3676_;
  assign new_n3678_ = ~new_n3673_ & ~new_n3677_;
  assign new_n3679_ = ~new_n3657_ & ~new_n3678_;
  assign new_n3680_ = \C<27>  & new_n3657_;
  assign new_n3681_ = ~new_n3679_ & ~new_n3680_;
  assign new_n3682_ = ~new_n3632_ & ~new_n3681_;
  assign new_n3683_ = ~new_n3669_ & ~new_n3682_;
  assign \C_new<27>  = ~\reset<0>  & ~new_n3683_;
  assign new_n3685_ = \encrypt<0>  & \inreg<27> ;
  assign new_n3686_ = ~\encrypt<0>  & \inreg<35> ;
  assign new_n3687_ = ~new_n3685_ & ~new_n3686_;
  assign new_n3688_ = new_n3632_ & ~new_n3687_;
  assign new_n3689_ = \C<27>  & ~new_n3665_;
  assign new_n3690_ = \C<0>  & new_n3665_;
  assign new_n3691_ = ~new_n3689_ & ~new_n3690_;
  assign new_n3692_ = \encrypt_mode<0>  & ~new_n3691_;
  assign new_n3693_ = \C<25>  & ~new_n3665_;
  assign new_n3694_ = \C<24>  & new_n3665_;
  assign new_n3695_ = ~new_n3693_ & ~new_n3694_;
  assign new_n3696_ = ~\encrypt_mode<0>  & ~new_n3695_;
  assign new_n3697_ = ~new_n3692_ & ~new_n3696_;
  assign new_n3698_ = ~new_n3657_ & ~new_n3697_;
  assign new_n3699_ = \C<26>  & new_n3657_;
  assign new_n3700_ = ~new_n3698_ & ~new_n3699_;
  assign new_n3701_ = ~new_n3632_ & ~new_n3700_;
  assign new_n3702_ = ~new_n3688_ & ~new_n3701_;
  assign \C_new<26>  = ~\reset<0>  & ~new_n3702_;
  assign new_n3704_ = \C<27>  & new_n3665_;
  assign new_n3705_ = ~new_n3674_ & ~new_n3704_;
  assign new_n3706_ = \encrypt_mode<0>  & ~new_n3705_;
  assign new_n3707_ = \C<24>  & ~new_n3665_;
  assign new_n3708_ = \C<23>  & new_n3665_;
  assign new_n3709_ = ~new_n3707_ & ~new_n3708_;
  assign new_n3710_ = ~\encrypt_mode<0>  & ~new_n3709_;
  assign new_n3711_ = ~new_n3706_ & ~new_n3710_;
  assign new_n3712_ = ~new_n3657_ & ~new_n3711_;
  assign new_n3713_ = \C<25>  & new_n3657_;
  assign new_n3714_ = ~new_n3712_ & ~new_n3713_;
  assign new_n3715_ = ~new_n3632_ & ~new_n3714_;
  assign new_n3716_ = \encrypt<0>  & \inreg<35> ;
  assign new_n3717_ = ~\encrypt<0>  & \inreg<43> ;
  assign new_n3718_ = ~new_n3716_ & ~new_n3717_;
  assign new_n3719_ = new_n3632_ & ~new_n3718_;
  assign new_n3720_ = ~new_n3715_ & ~new_n3719_;
  assign \C_new<25>  = ~\reset<0>  & ~new_n3720_;
  assign new_n3722_ = \C<26>  & new_n3665_;
  assign new_n3723_ = ~new_n3693_ & ~new_n3722_;
  assign new_n3724_ = \encrypt_mode<0>  & ~new_n3723_;
  assign new_n3725_ = \C<23>  & ~new_n3665_;
  assign new_n3726_ = \C<22>  & new_n3665_;
  assign new_n3727_ = ~new_n3725_ & ~new_n3726_;
  assign new_n3728_ = ~\encrypt_mode<0>  & ~new_n3727_;
  assign new_n3729_ = ~new_n3724_ & ~new_n3728_;
  assign new_n3730_ = ~new_n3657_ & ~new_n3729_;
  assign new_n3731_ = \C<24>  & new_n3657_;
  assign new_n3732_ = ~new_n3730_ & ~new_n3731_;
  assign new_n3733_ = ~new_n3632_ & ~new_n3732_;
  assign new_n3734_ = \encrypt<0>  & \inreg<43> ;
  assign new_n3735_ = ~\encrypt<0>  & \inreg<51> ;
  assign new_n3736_ = ~new_n3734_ & ~new_n3735_;
  assign new_n3737_ = new_n3632_ & ~new_n3736_;
  assign new_n3738_ = ~new_n3733_ & ~new_n3737_;
  assign \C_new<24>  = ~\reset<0>  & ~new_n3738_;
  assign new_n3740_ = \data_in<2>  & ~\encrypt<0> ;
  assign new_n3741_ = \encrypt<0>  & \inreg<51> ;
  assign new_n3742_ = ~new_n3740_ & ~new_n3741_;
  assign new_n3743_ = new_n3632_ & ~new_n3742_;
  assign new_n3744_ = ~new_n3675_ & ~new_n3707_;
  assign new_n3745_ = \encrypt_mode<0>  & ~new_n3744_;
  assign new_n3746_ = \C<21>  & new_n3665_;
  assign new_n3747_ = \C<22>  & ~new_n3665_;
  assign new_n3748_ = ~new_n3746_ & ~new_n3747_;
  assign new_n3749_ = ~\encrypt_mode<0>  & ~new_n3748_;
  assign new_n3750_ = ~new_n3745_ & ~new_n3749_;
  assign new_n3751_ = ~new_n3657_ & ~new_n3750_;
  assign new_n3752_ = \C<23>  & new_n3657_;
  assign new_n3753_ = ~new_n3751_ & ~new_n3752_;
  assign new_n3754_ = ~new_n3632_ & ~new_n3753_;
  assign new_n3755_ = ~new_n3743_ & ~new_n3754_;
  assign \C_new<23>  = ~\reset<0>  & ~new_n3755_;
  assign new_n3757_ = \data_in<2>  & \encrypt<0> ;
  assign new_n3758_ = ~\encrypt<0>  & \inreg<2> ;
  assign new_n3759_ = ~new_n3757_ & ~new_n3758_;
  assign new_n3760_ = new_n3632_ & ~new_n3759_;
  assign new_n3761_ = ~new_n3694_ & ~new_n3725_;
  assign new_n3762_ = \encrypt_mode<0>  & ~new_n3761_;
  assign new_n3763_ = \C<20>  & new_n3665_;
  assign new_n3764_ = \C<21>  & ~new_n3665_;
  assign new_n3765_ = ~new_n3763_ & ~new_n3764_;
  assign new_n3766_ = ~\encrypt_mode<0>  & ~new_n3765_;
  assign new_n3767_ = ~new_n3762_ & ~new_n3766_;
  assign new_n3768_ = ~new_n3657_ & ~new_n3767_;
  assign new_n3769_ = \C<22>  & new_n3657_;
  assign new_n3770_ = ~new_n3768_ & ~new_n3769_;
  assign new_n3771_ = ~new_n3632_ & ~new_n3770_;
  assign new_n3772_ = ~new_n3760_ & ~new_n3771_;
  assign \C_new<22>  = ~\reset<0>  & ~new_n3772_;
  assign new_n3774_ = ~\encrypt<0>  & \inreg<10> ;
  assign new_n3775_ = \encrypt<0>  & \inreg<2> ;
  assign new_n3776_ = ~new_n3774_ & ~new_n3775_;
  assign new_n3777_ = new_n3632_ & ~new_n3776_;
  assign new_n3778_ = ~new_n3708_ & ~new_n3747_;
  assign new_n3779_ = \encrypt_mode<0>  & ~new_n3778_;
  assign new_n3780_ = \C<20>  & ~new_n3665_;
  assign new_n3781_ = \C<19>  & new_n3665_;
  assign new_n3782_ = ~new_n3780_ & ~new_n3781_;
  assign new_n3783_ = ~\encrypt_mode<0>  & ~new_n3782_;
  assign new_n3784_ = ~new_n3779_ & ~new_n3783_;
  assign new_n3785_ = ~new_n3657_ & ~new_n3784_;
  assign new_n3786_ = \C<21>  & new_n3657_;
  assign new_n3787_ = ~new_n3785_ & ~new_n3786_;
  assign new_n3788_ = ~new_n3632_ & ~new_n3787_;
  assign new_n3789_ = ~new_n3777_ & ~new_n3788_;
  assign \C_new<21>  = ~\reset<0>  & ~new_n3789_;
  assign new_n3791_ = ~new_n3726_ & ~new_n3764_;
  assign new_n3792_ = \encrypt_mode<0>  & ~new_n3791_;
  assign new_n3793_ = \C<19>  & ~new_n3665_;
  assign new_n3794_ = \C<18>  & new_n3665_;
  assign new_n3795_ = ~new_n3793_ & ~new_n3794_;
  assign new_n3796_ = ~\encrypt_mode<0>  & ~new_n3795_;
  assign new_n3797_ = ~new_n3792_ & ~new_n3796_;
  assign new_n3798_ = ~new_n3657_ & ~new_n3797_;
  assign new_n3799_ = \C<20>  & new_n3657_;
  assign new_n3800_ = ~new_n3798_ & ~new_n3799_;
  assign new_n3801_ = ~new_n3632_ & ~new_n3800_;
  assign new_n3802_ = \encrypt<0>  & \inreg<10> ;
  assign new_n3803_ = ~\encrypt<0>  & \inreg<18> ;
  assign new_n3804_ = ~new_n3802_ & ~new_n3803_;
  assign new_n3805_ = new_n3632_ & ~new_n3804_;
  assign new_n3806_ = ~new_n3801_ & ~new_n3805_;
  assign \C_new<20>  = ~\reset<0>  & ~new_n3806_;
  assign new_n3808_ = ~new_n3746_ & ~new_n3780_;
  assign new_n3809_ = \encrypt_mode<0>  & ~new_n3808_;
  assign new_n3810_ = \C<18>  & ~new_n3665_;
  assign new_n3811_ = \C<17>  & new_n3665_;
  assign new_n3812_ = ~new_n3810_ & ~new_n3811_;
  assign new_n3813_ = ~\encrypt_mode<0>  & ~new_n3812_;
  assign new_n3814_ = ~new_n3809_ & ~new_n3813_;
  assign new_n3815_ = ~new_n3657_ & ~new_n3814_;
  assign new_n3816_ = \C<19>  & new_n3657_;
  assign new_n3817_ = ~new_n3815_ & ~new_n3816_;
  assign new_n3818_ = ~new_n3632_ & ~new_n3817_;
  assign new_n3819_ = \encrypt<0>  & \inreg<18> ;
  assign new_n3820_ = ~\encrypt<0>  & \inreg<26> ;
  assign new_n3821_ = ~new_n3819_ & ~new_n3820_;
  assign new_n3822_ = new_n3632_ & ~new_n3821_;
  assign new_n3823_ = ~new_n3818_ & ~new_n3822_;
  assign \C_new<19>  = ~\reset<0>  & ~new_n3823_;
  assign new_n3825_ = ~new_n3763_ & ~new_n3793_;
  assign new_n3826_ = \encrypt_mode<0>  & ~new_n3825_;
  assign new_n3827_ = \C<17>  & ~new_n3665_;
  assign new_n3828_ = \C<16>  & new_n3665_;
  assign new_n3829_ = ~new_n3827_ & ~new_n3828_;
  assign new_n3830_ = ~\encrypt_mode<0>  & ~new_n3829_;
  assign new_n3831_ = ~new_n3826_ & ~new_n3830_;
  assign new_n3832_ = ~new_n3657_ & ~new_n3831_;
  assign new_n3833_ = \C<18>  & new_n3657_;
  assign new_n3834_ = ~new_n3832_ & ~new_n3833_;
  assign new_n3835_ = ~new_n3632_ & ~new_n3834_;
  assign new_n3836_ = \encrypt<0>  & \inreg<26> ;
  assign new_n3837_ = ~\encrypt<0>  & \inreg<34> ;
  assign new_n3838_ = ~new_n3836_ & ~new_n3837_;
  assign new_n3839_ = new_n3632_ & ~new_n3838_;
  assign new_n3840_ = ~new_n3835_ & ~new_n3839_;
  assign \C_new<18>  = ~\reset<0>  & ~new_n3840_;
  assign new_n3842_ = ~new_n3781_ & ~new_n3810_;
  assign new_n3843_ = \encrypt_mode<0>  & ~new_n3842_;
  assign new_n3844_ = \C<16>  & ~new_n3665_;
  assign new_n3845_ = \C<15>  & new_n3665_;
  assign new_n3846_ = ~new_n3844_ & ~new_n3845_;
  assign new_n3847_ = ~\encrypt_mode<0>  & ~new_n3846_;
  assign new_n3848_ = ~new_n3843_ & ~new_n3847_;
  assign new_n3849_ = ~new_n3657_ & ~new_n3848_;
  assign new_n3850_ = \C<17>  & new_n3657_;
  assign new_n3851_ = ~new_n3849_ & ~new_n3850_;
  assign new_n3852_ = ~new_n3632_ & ~new_n3851_;
  assign new_n3853_ = \encrypt<0>  & \inreg<34> ;
  assign new_n3854_ = ~\encrypt<0>  & \inreg<42> ;
  assign new_n3855_ = ~new_n3853_ & ~new_n3854_;
  assign new_n3856_ = new_n3632_ & ~new_n3855_;
  assign new_n3857_ = ~new_n3852_ & ~new_n3856_;
  assign \C_new<17>  = ~\reset<0>  & ~new_n3857_;
  assign new_n3859_ = ~new_n3794_ & ~new_n3827_;
  assign new_n3860_ = \encrypt_mode<0>  & ~new_n3859_;
  assign new_n3861_ = \C<15>  & ~new_n3665_;
  assign new_n3862_ = \C<14>  & new_n3665_;
  assign new_n3863_ = ~new_n3861_ & ~new_n3862_;
  assign new_n3864_ = ~\encrypt_mode<0>  & ~new_n3863_;
  assign new_n3865_ = ~new_n3860_ & ~new_n3864_;
  assign new_n3866_ = ~new_n3657_ & ~new_n3865_;
  assign new_n3867_ = \C<16>  & new_n3657_;
  assign new_n3868_ = ~new_n3866_ & ~new_n3867_;
  assign new_n3869_ = ~new_n3632_ & ~new_n3868_;
  assign new_n3870_ = \encrypt<0>  & \inreg<42> ;
  assign new_n3871_ = ~\encrypt<0>  & \inreg<50> ;
  assign new_n3872_ = ~new_n3870_ & ~new_n3871_;
  assign new_n3873_ = new_n3632_ & ~new_n3872_;
  assign new_n3874_ = ~new_n3869_ & ~new_n3873_;
  assign \C_new<16>  = ~\reset<0>  & ~new_n3874_;
  assign new_n3876_ = \data_in<1>  & ~\encrypt<0> ;
  assign new_n3877_ = \encrypt<0>  & \inreg<50> ;
  assign new_n3878_ = ~new_n3876_ & ~new_n3877_;
  assign new_n3879_ = new_n3632_ & ~new_n3878_;
  assign new_n3880_ = ~new_n3811_ & ~new_n3844_;
  assign new_n3881_ = \encrypt_mode<0>  & ~new_n3880_;
  assign new_n3882_ = \C<13>  & new_n3665_;
  assign new_n3883_ = \C<14>  & ~new_n3665_;
  assign new_n3884_ = ~new_n3882_ & ~new_n3883_;
  assign new_n3885_ = ~\encrypt_mode<0>  & ~new_n3884_;
  assign new_n3886_ = ~new_n3881_ & ~new_n3885_;
  assign new_n3887_ = ~new_n3657_ & ~new_n3886_;
  assign new_n3888_ = \C<15>  & new_n3657_;
  assign new_n3889_ = ~new_n3887_ & ~new_n3888_;
  assign new_n3890_ = ~new_n3632_ & ~new_n3889_;
  assign new_n3891_ = ~new_n3879_ & ~new_n3890_;
  assign \C_new<15>  = ~\reset<0>  & ~new_n3891_;
  assign new_n3893_ = \data_in<1>  & \encrypt<0> ;
  assign new_n3894_ = ~\encrypt<0>  & \inreg<1> ;
  assign new_n3895_ = ~new_n3893_ & ~new_n3894_;
  assign new_n3896_ = new_n3632_ & ~new_n3895_;
  assign new_n3897_ = ~new_n3828_ & ~new_n3861_;
  assign new_n3898_ = \encrypt_mode<0>  & ~new_n3897_;
  assign new_n3899_ = \C<12>  & new_n3665_;
  assign new_n3900_ = \C<13>  & ~new_n3665_;
  assign new_n3901_ = ~new_n3899_ & ~new_n3900_;
  assign new_n3902_ = ~\encrypt_mode<0>  & ~new_n3901_;
  assign new_n3903_ = ~new_n3898_ & ~new_n3902_;
  assign new_n3904_ = ~new_n3657_ & ~new_n3903_;
  assign new_n3905_ = \C<14>  & new_n3657_;
  assign new_n3906_ = ~new_n3904_ & ~new_n3905_;
  assign new_n3907_ = ~new_n3632_ & ~new_n3906_;
  assign new_n3908_ = ~new_n3896_ & ~new_n3907_;
  assign \C_new<14>  = ~\reset<0>  & ~new_n3908_;
  assign new_n3910_ = ~new_n3845_ & ~new_n3883_;
  assign new_n3911_ = \encrypt_mode<0>  & ~new_n3910_;
  assign new_n3912_ = \C<12>  & ~new_n3665_;
  assign new_n3913_ = \C<11>  & new_n3665_;
  assign new_n3914_ = ~new_n3912_ & ~new_n3913_;
  assign new_n3915_ = ~\encrypt_mode<0>  & ~new_n3914_;
  assign new_n3916_ = ~new_n3911_ & ~new_n3915_;
  assign new_n3917_ = ~new_n3657_ & ~new_n3916_;
  assign new_n3918_ = \C<13>  & new_n3657_;
  assign new_n3919_ = ~new_n3917_ & ~new_n3918_;
  assign new_n3920_ = ~new_n3632_ & ~new_n3919_;
  assign new_n3921_ = \encrypt<0>  & \inreg<1> ;
  assign new_n3922_ = ~\encrypt<0>  & \inreg<9> ;
  assign new_n3923_ = ~new_n3921_ & ~new_n3922_;
  assign new_n3924_ = new_n3632_ & ~new_n3923_;
  assign new_n3925_ = ~new_n3920_ & ~new_n3924_;
  assign \C_new<13>  = ~\reset<0>  & ~new_n3925_;
  assign new_n3927_ = ~\encrypt<0>  & \inreg<17> ;
  assign new_n3928_ = \encrypt<0>  & \inreg<9> ;
  assign new_n3929_ = ~new_n3927_ & ~new_n3928_;
  assign new_n3930_ = new_n3632_ & ~new_n3929_;
  assign new_n3931_ = ~new_n3862_ & ~new_n3900_;
  assign new_n3932_ = \encrypt_mode<0>  & ~new_n3931_;
  assign new_n3933_ = \C<11>  & ~new_n3665_;
  assign new_n3934_ = \C<10>  & new_n3665_;
  assign new_n3935_ = ~new_n3933_ & ~new_n3934_;
  assign new_n3936_ = ~\encrypt_mode<0>  & ~new_n3935_;
  assign new_n3937_ = ~new_n3932_ & ~new_n3936_;
  assign new_n3938_ = ~new_n3657_ & ~new_n3937_;
  assign new_n3939_ = \C<12>  & new_n3657_;
  assign new_n3940_ = ~new_n3938_ & ~new_n3939_;
  assign new_n3941_ = ~new_n3632_ & ~new_n3940_;
  assign new_n3942_ = ~new_n3930_ & ~new_n3941_;
  assign \C_new<12>  = ~\reset<0>  & ~new_n3942_;
  assign new_n3944_ = \encrypt<0>  & \inreg<17> ;
  assign new_n3945_ = ~\encrypt<0>  & \inreg<25> ;
  assign new_n3946_ = ~new_n3944_ & ~new_n3945_;
  assign new_n3947_ = new_n3632_ & ~new_n3946_;
  assign new_n3948_ = ~new_n3882_ & ~new_n3912_;
  assign new_n3949_ = \encrypt_mode<0>  & ~new_n3948_;
  assign new_n3950_ = \C<9>  & new_n3665_;
  assign new_n3951_ = \C<10>  & ~new_n3665_;
  assign new_n3952_ = ~new_n3950_ & ~new_n3951_;
  assign new_n3953_ = ~\encrypt_mode<0>  & ~new_n3952_;
  assign new_n3954_ = ~new_n3949_ & ~new_n3953_;
  assign new_n3955_ = ~new_n3657_ & ~new_n3954_;
  assign new_n3956_ = \C<11>  & new_n3657_;
  assign new_n3957_ = ~new_n3955_ & ~new_n3956_;
  assign new_n3958_ = ~new_n3632_ & ~new_n3957_;
  assign new_n3959_ = ~new_n3947_ & ~new_n3958_;
  assign \C_new<11>  = ~\reset<0>  & ~new_n3959_;
  assign new_n3961_ = \encrypt<0>  & \inreg<25> ;
  assign new_n3962_ = ~\encrypt<0>  & \inreg<33> ;
  assign new_n3963_ = ~new_n3961_ & ~new_n3962_;
  assign new_n3964_ = new_n3632_ & ~new_n3963_;
  assign new_n3965_ = ~new_n3899_ & ~new_n3933_;
  assign new_n3966_ = \encrypt_mode<0>  & ~new_n3965_;
  assign new_n3967_ = \C<9>  & ~new_n3665_;
  assign new_n3968_ = \C<8>  & new_n3665_;
  assign new_n3969_ = ~new_n3967_ & ~new_n3968_;
  assign new_n3970_ = ~\encrypt_mode<0>  & ~new_n3969_;
  assign new_n3971_ = ~new_n3966_ & ~new_n3970_;
  assign new_n3972_ = ~new_n3657_ & ~new_n3971_;
  assign new_n3973_ = \C<10>  & new_n3657_;
  assign new_n3974_ = ~new_n3972_ & ~new_n3973_;
  assign new_n3975_ = ~new_n3632_ & ~new_n3974_;
  assign new_n3976_ = ~new_n3964_ & ~new_n3975_;
  assign \C_new<10>  = ~\reset<0>  & ~new_n3976_;
  assign new_n3978_ = \encrypt<0>  & \inreg<33> ;
  assign new_n3979_ = ~\encrypt<0>  & \inreg<41> ;
  assign new_n3980_ = ~new_n3978_ & ~new_n3979_;
  assign new_n3981_ = new_n3632_ & ~new_n3980_;
  assign new_n3982_ = ~new_n3913_ & ~new_n3951_;
  assign new_n3983_ = \encrypt_mode<0>  & ~new_n3982_;
  assign new_n3984_ = \C<8>  & ~new_n3665_;
  assign new_n3985_ = \C<7>  & new_n3665_;
  assign new_n3986_ = ~new_n3984_ & ~new_n3985_;
  assign new_n3987_ = ~\encrypt_mode<0>  & ~new_n3986_;
  assign new_n3988_ = ~new_n3983_ & ~new_n3987_;
  assign new_n3989_ = ~new_n3657_ & ~new_n3988_;
  assign new_n3990_ = \C<9>  & new_n3657_;
  assign new_n3991_ = ~new_n3989_ & ~new_n3990_;
  assign new_n3992_ = ~new_n3632_ & ~new_n3991_;
  assign new_n3993_ = ~new_n3981_ & ~new_n3992_;
  assign \C_new<9>  = ~\reset<0>  & ~new_n3993_;
  assign new_n3995_ = \encrypt<0>  & \inreg<41> ;
  assign new_n3996_ = ~\encrypt<0>  & \inreg<49> ;
  assign new_n3997_ = ~new_n3995_ & ~new_n3996_;
  assign new_n3998_ = new_n3632_ & ~new_n3997_;
  assign new_n3999_ = ~new_n3934_ & ~new_n3967_;
  assign new_n4000_ = \encrypt_mode<0>  & ~new_n3999_;
  assign new_n4001_ = \C<7>  & ~new_n3665_;
  assign new_n4002_ = \C<6>  & new_n3665_;
  assign new_n4003_ = ~new_n4001_ & ~new_n4002_;
  assign new_n4004_ = ~\encrypt_mode<0>  & ~new_n4003_;
  assign new_n4005_ = ~new_n4000_ & ~new_n4004_;
  assign new_n4006_ = ~new_n3657_ & ~new_n4005_;
  assign new_n4007_ = \C<8>  & new_n3657_;
  assign new_n4008_ = ~new_n4006_ & ~new_n4007_;
  assign new_n4009_ = ~new_n3632_ & ~new_n4008_;
  assign new_n4010_ = ~new_n3998_ & ~new_n4009_;
  assign \C_new<8>  = ~\reset<0>  & ~new_n4010_;
  assign new_n4012_ = \data_in<0>  & ~\encrypt<0> ;
  assign new_n4013_ = \encrypt<0>  & \inreg<49> ;
  assign new_n4014_ = ~new_n4012_ & ~new_n4013_;
  assign new_n4015_ = new_n3632_ & ~new_n4014_;
  assign new_n4016_ = ~new_n3950_ & ~new_n3984_;
  assign new_n4017_ = \encrypt_mode<0>  & ~new_n4016_;
  assign new_n4018_ = \C<5>  & new_n3665_;
  assign new_n4019_ = \C<6>  & ~new_n3665_;
  assign new_n4020_ = ~new_n4018_ & ~new_n4019_;
  assign new_n4021_ = ~\encrypt_mode<0>  & ~new_n4020_;
  assign new_n4022_ = ~new_n4017_ & ~new_n4021_;
  assign new_n4023_ = ~new_n3657_ & ~new_n4022_;
  assign new_n4024_ = \C<7>  & new_n3657_;
  assign new_n4025_ = ~new_n4023_ & ~new_n4024_;
  assign new_n4026_ = ~new_n3632_ & ~new_n4025_;
  assign new_n4027_ = ~new_n4015_ & ~new_n4026_;
  assign \C_new<7>  = ~\reset<0>  & ~new_n4027_;
  assign new_n4029_ = \data_in<0>  & \encrypt<0> ;
  assign new_n4030_ = ~\encrypt<0>  & \inreg<0> ;
  assign new_n4031_ = ~new_n4029_ & ~new_n4030_;
  assign new_n4032_ = new_n3632_ & ~new_n4031_;
  assign new_n4033_ = ~new_n3968_ & ~new_n4001_;
  assign new_n4034_ = \encrypt_mode<0>  & ~new_n4033_;
  assign new_n4035_ = \C<4>  & new_n3665_;
  assign new_n4036_ = \C<5>  & ~new_n3665_;
  assign new_n4037_ = ~new_n4035_ & ~new_n4036_;
  assign new_n4038_ = ~\encrypt_mode<0>  & ~new_n4037_;
  assign new_n4039_ = ~new_n4034_ & ~new_n4038_;
  assign new_n4040_ = ~new_n3657_ & ~new_n4039_;
  assign new_n4041_ = \C<6>  & new_n3657_;
  assign new_n4042_ = ~new_n4040_ & ~new_n4041_;
  assign new_n4043_ = ~new_n3632_ & ~new_n4042_;
  assign new_n4044_ = ~new_n4032_ & ~new_n4043_;
  assign \C_new<6>  = ~\reset<0>  & ~new_n4044_;
  assign new_n4046_ = ~new_n3985_ & ~new_n4019_;
  assign new_n4047_ = \encrypt_mode<0>  & ~new_n4046_;
  assign new_n4048_ = \C<4>  & ~new_n3665_;
  assign new_n4049_ = \C<3>  & new_n3665_;
  assign new_n4050_ = ~new_n4048_ & ~new_n4049_;
  assign new_n4051_ = ~\encrypt_mode<0>  & ~new_n4050_;
  assign new_n4052_ = ~new_n4047_ & ~new_n4051_;
  assign new_n4053_ = ~new_n3657_ & ~new_n4052_;
  assign new_n4054_ = \C<5>  & new_n3657_;
  assign new_n4055_ = ~new_n4053_ & ~new_n4054_;
  assign new_n4056_ = ~new_n3632_ & ~new_n4055_;
  assign new_n4057_ = \encrypt<0>  & \inreg<0> ;
  assign new_n4058_ = ~\encrypt<0>  & \inreg<8> ;
  assign new_n4059_ = ~new_n4057_ & ~new_n4058_;
  assign new_n4060_ = new_n3632_ & ~new_n4059_;
  assign new_n4061_ = ~new_n4056_ & ~new_n4060_;
  assign \C_new<5>  = ~\reset<0>  & ~new_n4061_;
  assign new_n4063_ = ~\encrypt<0>  & \inreg<16> ;
  assign new_n4064_ = \encrypt<0>  & \inreg<8> ;
  assign new_n4065_ = ~new_n4063_ & ~new_n4064_;
  assign new_n4066_ = new_n3632_ & ~new_n4065_;
  assign new_n4067_ = ~new_n4002_ & ~new_n4036_;
  assign new_n4068_ = \encrypt_mode<0>  & ~new_n4067_;
  assign new_n4069_ = \C<3>  & ~new_n3665_;
  assign new_n4070_ = \C<2>  & new_n3665_;
  assign new_n4071_ = ~new_n4069_ & ~new_n4070_;
  assign new_n4072_ = ~\encrypt_mode<0>  & ~new_n4071_;
  assign new_n4073_ = ~new_n4068_ & ~new_n4072_;
  assign new_n4074_ = ~new_n3657_ & ~new_n4073_;
  assign new_n4075_ = \C<4>  & new_n3657_;
  assign new_n4076_ = ~new_n4074_ & ~new_n4075_;
  assign new_n4077_ = ~new_n3632_ & ~new_n4076_;
  assign new_n4078_ = ~new_n4066_ & ~new_n4077_;
  assign \C_new<4>  = ~\reset<0>  & ~new_n4078_;
  assign new_n4080_ = ~new_n4018_ & ~new_n4048_;
  assign new_n4081_ = \encrypt_mode<0>  & ~new_n4080_;
  assign new_n4082_ = \C<2>  & ~new_n3665_;
  assign new_n4083_ = ~new_n3671_ & ~new_n4082_;
  assign new_n4084_ = ~\encrypt_mode<0>  & ~new_n4083_;
  assign new_n4085_ = ~new_n4081_ & ~new_n4084_;
  assign new_n4086_ = ~new_n3657_ & ~new_n4085_;
  assign new_n4087_ = \C<3>  & new_n3657_;
  assign new_n4088_ = ~new_n4086_ & ~new_n4087_;
  assign new_n4089_ = ~new_n3632_ & ~new_n4088_;
  assign new_n4090_ = \encrypt<0>  & \inreg<16> ;
  assign new_n4091_ = ~\encrypt<0>  & \inreg<24> ;
  assign new_n4092_ = ~new_n4090_ & ~new_n4091_;
  assign new_n4093_ = new_n3632_ & ~new_n4092_;
  assign new_n4094_ = ~new_n4089_ & ~new_n4093_;
  assign \C_new<3>  = ~\reset<0>  & ~new_n4094_;
  assign new_n4096_ = ~new_n4035_ & ~new_n4069_;
  assign new_n4097_ = \encrypt_mode<0>  & ~new_n4096_;
  assign new_n4098_ = \C<1>  & ~new_n3665_;
  assign new_n4099_ = ~new_n3690_ & ~new_n4098_;
  assign new_n4100_ = ~\encrypt_mode<0>  & ~new_n4099_;
  assign new_n4101_ = ~new_n4097_ & ~new_n4100_;
  assign new_n4102_ = ~new_n3657_ & ~new_n4101_;
  assign new_n4103_ = \C<2>  & new_n3657_;
  assign new_n4104_ = ~new_n4102_ & ~new_n4103_;
  assign new_n4105_ = ~new_n3632_ & ~new_n4104_;
  assign new_n4106_ = \encrypt<0>  & \inreg<24> ;
  assign new_n4107_ = ~\encrypt<0>  & \inreg<32> ;
  assign new_n4108_ = ~new_n4106_ & ~new_n4107_;
  assign new_n4109_ = new_n3632_ & ~new_n4108_;
  assign new_n4110_ = ~new_n4105_ & ~new_n4109_;
  assign \C_new<2>  = ~\reset<0>  & ~new_n4110_;
  assign new_n4112_ = \encrypt<0>  & \inreg<32> ;
  assign new_n4113_ = ~\encrypt<0>  & \inreg<40> ;
  assign new_n4114_ = ~new_n4112_ & ~new_n4113_;
  assign new_n4115_ = new_n3632_ & ~new_n4114_;
  assign new_n4116_ = \C<1>  & new_n3657_;
  assign new_n4117_ = ~new_n4049_ & ~new_n4082_;
  assign new_n4118_ = \encrypt_mode<0>  & ~new_n4117_;
  assign new_n4119_ = ~new_n3670_ & ~new_n3704_;
  assign new_n4120_ = ~\encrypt_mode<0>  & ~new_n4119_;
  assign new_n4121_ = ~new_n4118_ & ~new_n4120_;
  assign new_n4122_ = ~new_n3657_ & ~new_n4121_;
  assign new_n4123_ = ~new_n4116_ & ~new_n4122_;
  assign new_n4124_ = ~new_n3632_ & ~new_n4123_;
  assign new_n4125_ = ~new_n4115_ & ~new_n4124_;
  assign \C_new<1>  = ~\reset<0>  & ~new_n4125_;
  assign new_n4127_ = \encrypt<0>  & \inreg<40> ;
  assign new_n4128_ = ~\encrypt<0>  & \inreg<48> ;
  assign new_n4129_ = ~new_n4127_ & ~new_n4128_;
  assign new_n4130_ = new_n3632_ & ~new_n4129_;
  assign new_n4131_ = \C<0>  & new_n3657_;
  assign new_n4132_ = ~new_n3689_ & ~new_n3722_;
  assign new_n4133_ = ~\encrypt_mode<0>  & ~new_n4132_;
  assign new_n4134_ = ~new_n4070_ & ~new_n4098_;
  assign new_n4135_ = \encrypt_mode<0>  & ~new_n4134_;
  assign new_n4136_ = ~new_n4133_ & ~new_n4135_;
  assign new_n4137_ = ~new_n3657_ & ~new_n4136_;
  assign new_n4138_ = ~new_n4131_ & ~new_n4137_;
  assign new_n4139_ = ~new_n3632_ & ~new_n4138_;
  assign new_n4140_ = ~new_n4130_ & ~new_n4139_;
  assign \C_new<0>  = ~\reset<0>  & ~new_n4140_;
  assign new_n4142_ = \data_in<3>  & ~\encrypt<0> ;
  assign new_n4143_ = \encrypt<0>  & \inreg<54> ;
  assign new_n4144_ = ~new_n4142_ & ~new_n4143_;
  assign new_n4145_ = new_n3632_ & ~new_n4144_;
  assign new_n4146_ = \D<0>  & ~new_n3665_;
  assign new_n4147_ = \D<1>  & new_n3665_;
  assign new_n4148_ = ~new_n4146_ & ~new_n4147_;
  assign new_n4149_ = \encrypt_mode<0>  & ~new_n4148_;
  assign new_n4150_ = \D<26>  & ~new_n3665_;
  assign new_n4151_ = \D<25>  & new_n3665_;
  assign new_n4152_ = ~new_n4150_ & ~new_n4151_;
  assign new_n4153_ = ~\encrypt_mode<0>  & ~new_n4152_;
  assign new_n4154_ = ~new_n4149_ & ~new_n4153_;
  assign new_n4155_ = ~new_n3657_ & ~new_n4154_;
  assign new_n4156_ = \D<27>  & new_n3657_;
  assign new_n4157_ = ~new_n4155_ & ~new_n4156_;
  assign new_n4158_ = ~new_n3632_ & ~new_n4157_;
  assign new_n4159_ = ~new_n4145_ & ~new_n4158_;
  assign \D_new<27>  = ~\reset<0>  & ~new_n4159_;
  assign new_n4161_ = \data_in<3>  & \encrypt<0> ;
  assign new_n4162_ = ~\encrypt<0>  & \inreg<3> ;
  assign new_n4163_ = ~new_n4161_ & ~new_n4162_;
  assign new_n4164_ = new_n3632_ & ~new_n4163_;
  assign new_n4165_ = \D<27>  & ~new_n3665_;
  assign new_n4166_ = \D<0>  & new_n3665_;
  assign new_n4167_ = ~new_n4165_ & ~new_n4166_;
  assign new_n4168_ = \encrypt_mode<0>  & ~new_n4167_;
  assign new_n4169_ = \D<24>  & new_n3665_;
  assign new_n4170_ = \D<25>  & ~new_n3665_;
  assign new_n4171_ = ~new_n4169_ & ~new_n4170_;
  assign new_n4172_ = ~\encrypt_mode<0>  & ~new_n4171_;
  assign new_n4173_ = ~new_n4168_ & ~new_n4172_;
  assign new_n4174_ = ~new_n3657_ & ~new_n4173_;
  assign new_n4175_ = \D<26>  & new_n3657_;
  assign new_n4176_ = ~new_n4174_ & ~new_n4175_;
  assign new_n4177_ = ~new_n3632_ & ~new_n4176_;
  assign new_n4178_ = ~new_n4164_ & ~new_n4177_;
  assign \D_new<26>  = ~\reset<0>  & ~new_n4178_;
  assign new_n4180_ = ~\encrypt<0>  & \inreg<11> ;
  assign new_n4181_ = \encrypt<0>  & \inreg<3> ;
  assign new_n4182_ = ~new_n4180_ & ~new_n4181_;
  assign new_n4183_ = new_n3632_ & ~new_n4182_;
  assign new_n4184_ = \D<27>  & new_n3665_;
  assign new_n4185_ = ~new_n4150_ & ~new_n4184_;
  assign new_n4186_ = \encrypt_mode<0>  & ~new_n4185_;
  assign new_n4187_ = \D<24>  & ~new_n3665_;
  assign new_n4188_ = \D<23>  & new_n3665_;
  assign new_n4189_ = ~new_n4187_ & ~new_n4188_;
  assign new_n4190_ = ~\encrypt_mode<0>  & ~new_n4189_;
  assign new_n4191_ = ~new_n4186_ & ~new_n4190_;
  assign new_n4192_ = ~new_n3657_ & ~new_n4191_;
  assign new_n4193_ = \D<25>  & new_n3657_;
  assign new_n4194_ = ~new_n4192_ & ~new_n4193_;
  assign new_n4195_ = ~new_n3632_ & ~new_n4194_;
  assign new_n4196_ = ~new_n4183_ & ~new_n4195_;
  assign \D_new<25>  = ~\reset<0>  & ~new_n4196_;
  assign new_n4198_ = \D<26>  & new_n3665_;
  assign new_n4199_ = ~new_n4170_ & ~new_n4198_;
  assign new_n4200_ = \encrypt_mode<0>  & ~new_n4199_;
  assign new_n4201_ = \D<23>  & ~new_n3665_;
  assign new_n4202_ = \D<22>  & new_n3665_;
  assign new_n4203_ = ~new_n4201_ & ~new_n4202_;
  assign new_n4204_ = ~\encrypt_mode<0>  & ~new_n4203_;
  assign new_n4205_ = ~new_n4200_ & ~new_n4204_;
  assign new_n4206_ = ~new_n3657_ & ~new_n4205_;
  assign new_n4207_ = \D<24>  & new_n3657_;
  assign new_n4208_ = ~new_n4206_ & ~new_n4207_;
  assign new_n4209_ = ~new_n3632_ & ~new_n4208_;
  assign new_n4210_ = \encrypt<0>  & \inreg<11> ;
  assign new_n4211_ = ~\encrypt<0>  & \inreg<19> ;
  assign new_n4212_ = ~new_n4210_ & ~new_n4211_;
  assign new_n4213_ = new_n3632_ & ~new_n4212_;
  assign new_n4214_ = ~new_n4209_ & ~new_n4213_;
  assign \D_new<24>  = ~\reset<0>  & ~new_n4214_;
  assign new_n4216_ = \data_in<4>  & ~\encrypt<0> ;
  assign new_n4217_ = \encrypt<0>  & \inreg<19> ;
  assign new_n4218_ = ~new_n4216_ & ~new_n4217_;
  assign new_n4219_ = new_n3632_ & ~new_n4218_;
  assign new_n4220_ = ~new_n4151_ & ~new_n4187_;
  assign new_n4221_ = \encrypt_mode<0>  & ~new_n4220_;
  assign new_n4222_ = \D<21>  & new_n3665_;
  assign new_n4223_ = \D<22>  & ~new_n3665_;
  assign new_n4224_ = ~new_n4222_ & ~new_n4223_;
  assign new_n4225_ = ~\encrypt_mode<0>  & ~new_n4224_;
  assign new_n4226_ = ~new_n4221_ & ~new_n4225_;
  assign new_n4227_ = ~new_n3657_ & ~new_n4226_;
  assign new_n4228_ = \D<23>  & new_n3657_;
  assign new_n4229_ = ~new_n4227_ & ~new_n4228_;
  assign new_n4230_ = ~new_n3632_ & ~new_n4229_;
  assign new_n4231_ = ~new_n4219_ & ~new_n4230_;
  assign \D_new<23>  = ~\reset<0>  & ~new_n4231_;
  assign new_n4233_ = \data_in<4>  & \encrypt<0> ;
  assign new_n4234_ = ~\encrypt<0>  & \inreg<4> ;
  assign new_n4235_ = ~new_n4233_ & ~new_n4234_;
  assign new_n4236_ = new_n3632_ & ~new_n4235_;
  assign new_n4237_ = ~new_n4169_ & ~new_n4201_;
  assign new_n4238_ = \encrypt_mode<0>  & ~new_n4237_;
  assign new_n4239_ = \D<20>  & new_n3665_;
  assign new_n4240_ = \D<21>  & ~new_n3665_;
  assign new_n4241_ = ~new_n4239_ & ~new_n4240_;
  assign new_n4242_ = ~\encrypt_mode<0>  & ~new_n4241_;
  assign new_n4243_ = ~new_n4238_ & ~new_n4242_;
  assign new_n4244_ = ~new_n3657_ & ~new_n4243_;
  assign new_n4245_ = \D<22>  & new_n3657_;
  assign new_n4246_ = ~new_n4244_ & ~new_n4245_;
  assign new_n4247_ = ~new_n3632_ & ~new_n4246_;
  assign new_n4248_ = ~new_n4236_ & ~new_n4247_;
  assign \D_new<22>  = ~\reset<0>  & ~new_n4248_;
  assign new_n4250_ = ~\encrypt<0>  & \inreg<12> ;
  assign new_n4251_ = \encrypt<0>  & \inreg<4> ;
  assign new_n4252_ = ~new_n4250_ & ~new_n4251_;
  assign new_n4253_ = new_n3632_ & ~new_n4252_;
  assign new_n4254_ = ~new_n4188_ & ~new_n4223_;
  assign new_n4255_ = \encrypt_mode<0>  & ~new_n4254_;
  assign new_n4256_ = \D<20>  & ~new_n3665_;
  assign new_n4257_ = \D<19>  & new_n3665_;
  assign new_n4258_ = ~new_n4256_ & ~new_n4257_;
  assign new_n4259_ = ~\encrypt_mode<0>  & ~new_n4258_;
  assign new_n4260_ = ~new_n4255_ & ~new_n4259_;
  assign new_n4261_ = ~new_n3657_ & ~new_n4260_;
  assign new_n4262_ = \D<21>  & new_n3657_;
  assign new_n4263_ = ~new_n4261_ & ~new_n4262_;
  assign new_n4264_ = ~new_n3632_ & ~new_n4263_;
  assign new_n4265_ = ~new_n4253_ & ~new_n4264_;
  assign \D_new<21>  = ~\reset<0>  & ~new_n4265_;
  assign new_n4267_ = ~new_n4202_ & ~new_n4240_;
  assign new_n4268_ = \encrypt_mode<0>  & ~new_n4267_;
  assign new_n4269_ = \D<19>  & ~new_n3665_;
  assign new_n4270_ = \D<18>  & new_n3665_;
  assign new_n4271_ = ~new_n4269_ & ~new_n4270_;
  assign new_n4272_ = ~\encrypt_mode<0>  & ~new_n4271_;
  assign new_n4273_ = ~new_n4268_ & ~new_n4272_;
  assign new_n4274_ = ~new_n3657_ & ~new_n4273_;
  assign new_n4275_ = \D<20>  & new_n3657_;
  assign new_n4276_ = ~new_n4274_ & ~new_n4275_;
  assign new_n4277_ = ~new_n3632_ & ~new_n4276_;
  assign new_n4278_ = \encrypt<0>  & \inreg<12> ;
  assign new_n4279_ = ~\encrypt<0>  & \inreg<20> ;
  assign new_n4280_ = ~new_n4278_ & ~new_n4279_;
  assign new_n4281_ = new_n3632_ & ~new_n4280_;
  assign new_n4282_ = ~new_n4277_ & ~new_n4281_;
  assign \D_new<20>  = ~\reset<0>  & ~new_n4282_;
  assign new_n4284_ = ~new_n4222_ & ~new_n4256_;
  assign new_n4285_ = \encrypt_mode<0>  & ~new_n4284_;
  assign new_n4286_ = \D<18>  & ~new_n3665_;
  assign new_n4287_ = \D<17>  & new_n3665_;
  assign new_n4288_ = ~new_n4286_ & ~new_n4287_;
  assign new_n4289_ = ~\encrypt_mode<0>  & ~new_n4288_;
  assign new_n4290_ = ~new_n4285_ & ~new_n4289_;
  assign new_n4291_ = ~new_n3657_ & ~new_n4290_;
  assign new_n4292_ = \D<19>  & new_n3657_;
  assign new_n4293_ = ~new_n4291_ & ~new_n4292_;
  assign new_n4294_ = ~new_n3632_ & ~new_n4293_;
  assign new_n4295_ = \encrypt<0>  & \inreg<20> ;
  assign new_n4296_ = ~\encrypt<0>  & \inreg<28> ;
  assign new_n4297_ = ~new_n4295_ & ~new_n4296_;
  assign new_n4298_ = new_n3632_ & ~new_n4297_;
  assign new_n4299_ = ~new_n4294_ & ~new_n4298_;
  assign \D_new<19>  = ~\reset<0>  & ~new_n4299_;
  assign new_n4301_ = ~new_n4239_ & ~new_n4269_;
  assign new_n4302_ = \encrypt_mode<0>  & ~new_n4301_;
  assign new_n4303_ = \D<17>  & ~new_n3665_;
  assign new_n4304_ = \D<16>  & new_n3665_;
  assign new_n4305_ = ~new_n4303_ & ~new_n4304_;
  assign new_n4306_ = ~\encrypt_mode<0>  & ~new_n4305_;
  assign new_n4307_ = ~new_n4302_ & ~new_n4306_;
  assign new_n4308_ = ~new_n3657_ & ~new_n4307_;
  assign new_n4309_ = \D<18>  & new_n3657_;
  assign new_n4310_ = ~new_n4308_ & ~new_n4309_;
  assign new_n4311_ = ~new_n3632_ & ~new_n4310_;
  assign new_n4312_ = \encrypt<0>  & \inreg<28> ;
  assign new_n4313_ = ~\encrypt<0>  & \inreg<36> ;
  assign new_n4314_ = ~new_n4312_ & ~new_n4313_;
  assign new_n4315_ = new_n3632_ & ~new_n4314_;
  assign new_n4316_ = ~new_n4311_ & ~new_n4315_;
  assign \D_new<18>  = ~\reset<0>  & ~new_n4316_;
  assign new_n4318_ = ~new_n4257_ & ~new_n4286_;
  assign new_n4319_ = \encrypt_mode<0>  & ~new_n4318_;
  assign new_n4320_ = \D<16>  & ~new_n3665_;
  assign new_n4321_ = \D<15>  & new_n3665_;
  assign new_n4322_ = ~new_n4320_ & ~new_n4321_;
  assign new_n4323_ = ~\encrypt_mode<0>  & ~new_n4322_;
  assign new_n4324_ = ~new_n4319_ & ~new_n4323_;
  assign new_n4325_ = ~new_n3657_ & ~new_n4324_;
  assign new_n4326_ = \D<17>  & new_n3657_;
  assign new_n4327_ = ~new_n4325_ & ~new_n4326_;
  assign new_n4328_ = ~new_n3632_ & ~new_n4327_;
  assign new_n4329_ = \encrypt<0>  & \inreg<36> ;
  assign new_n4330_ = ~\encrypt<0>  & \inreg<44> ;
  assign new_n4331_ = ~new_n4329_ & ~new_n4330_;
  assign new_n4332_ = new_n3632_ & ~new_n4331_;
  assign new_n4333_ = ~new_n4328_ & ~new_n4332_;
  assign \D_new<17>  = ~\reset<0>  & ~new_n4333_;
  assign new_n4335_ = ~new_n4270_ & ~new_n4303_;
  assign new_n4336_ = \encrypt_mode<0>  & ~new_n4335_;
  assign new_n4337_ = \D<15>  & ~new_n3665_;
  assign new_n4338_ = \D<14>  & new_n3665_;
  assign new_n4339_ = ~new_n4337_ & ~new_n4338_;
  assign new_n4340_ = ~\encrypt_mode<0>  & ~new_n4339_;
  assign new_n4341_ = ~new_n4336_ & ~new_n4340_;
  assign new_n4342_ = ~new_n3657_ & ~new_n4341_;
  assign new_n4343_ = \D<16>  & new_n3657_;
  assign new_n4344_ = ~new_n4342_ & ~new_n4343_;
  assign new_n4345_ = ~new_n3632_ & ~new_n4344_;
  assign new_n4346_ = \encrypt<0>  & \inreg<44> ;
  assign new_n4347_ = ~\encrypt<0>  & \inreg<52> ;
  assign new_n4348_ = ~new_n4346_ & ~new_n4347_;
  assign new_n4349_ = new_n3632_ & ~new_n4348_;
  assign new_n4350_ = ~new_n4345_ & ~new_n4349_;
  assign \D_new<16>  = ~\reset<0>  & ~new_n4350_;
  assign new_n4352_ = \data_in<5>  & ~\encrypt<0> ;
  assign new_n4353_ = \encrypt<0>  & \inreg<52> ;
  assign new_n4354_ = ~new_n4352_ & ~new_n4353_;
  assign new_n4355_ = new_n3632_ & ~new_n4354_;
  assign new_n4356_ = ~new_n4287_ & ~new_n4320_;
  assign new_n4357_ = \encrypt_mode<0>  & ~new_n4356_;
  assign new_n4358_ = \D<13>  & new_n3665_;
  assign new_n4359_ = \D<14>  & ~new_n3665_;
  assign new_n4360_ = ~new_n4358_ & ~new_n4359_;
  assign new_n4361_ = ~\encrypt_mode<0>  & ~new_n4360_;
  assign new_n4362_ = ~new_n4357_ & ~new_n4361_;
  assign new_n4363_ = ~new_n3657_ & ~new_n4362_;
  assign new_n4364_ = \D<15>  & new_n3657_;
  assign new_n4365_ = ~new_n4363_ & ~new_n4364_;
  assign new_n4366_ = ~new_n3632_ & ~new_n4365_;
  assign new_n4367_ = ~new_n4355_ & ~new_n4366_;
  assign \D_new<15>  = ~\reset<0>  & ~new_n4367_;
  assign new_n4369_ = \data_in<5>  & \encrypt<0> ;
  assign new_n4370_ = ~\encrypt<0>  & \inreg<5> ;
  assign new_n4371_ = ~new_n4369_ & ~new_n4370_;
  assign new_n4372_ = new_n3632_ & ~new_n4371_;
  assign new_n4373_ = ~new_n4304_ & ~new_n4337_;
  assign new_n4374_ = \encrypt_mode<0>  & ~new_n4373_;
  assign new_n4375_ = \D<12>  & new_n3665_;
  assign new_n4376_ = \D<13>  & ~new_n3665_;
  assign new_n4377_ = ~new_n4375_ & ~new_n4376_;
  assign new_n4378_ = ~\encrypt_mode<0>  & ~new_n4377_;
  assign new_n4379_ = ~new_n4374_ & ~new_n4378_;
  assign new_n4380_ = ~new_n3657_ & ~new_n4379_;
  assign new_n4381_ = \D<14>  & new_n3657_;
  assign new_n4382_ = ~new_n4380_ & ~new_n4381_;
  assign new_n4383_ = ~new_n3632_ & ~new_n4382_;
  assign new_n4384_ = ~new_n4372_ & ~new_n4383_;
  assign \D_new<14>  = ~\reset<0>  & ~new_n4384_;
  assign new_n4386_ = ~\encrypt<0>  & \inreg<13> ;
  assign new_n4387_ = \encrypt<0>  & \inreg<5> ;
  assign new_n4388_ = ~new_n4386_ & ~new_n4387_;
  assign new_n4389_ = new_n3632_ & ~new_n4388_;
  assign new_n4390_ = ~new_n4321_ & ~new_n4359_;
  assign new_n4391_ = \encrypt_mode<0>  & ~new_n4390_;
  assign new_n4392_ = \D<12>  & ~new_n3665_;
  assign new_n4393_ = \D<11>  & new_n3665_;
  assign new_n4394_ = ~new_n4392_ & ~new_n4393_;
  assign new_n4395_ = ~\encrypt_mode<0>  & ~new_n4394_;
  assign new_n4396_ = ~new_n4391_ & ~new_n4395_;
  assign new_n4397_ = ~new_n3657_ & ~new_n4396_;
  assign new_n4398_ = \D<13>  & new_n3657_;
  assign new_n4399_ = ~new_n4397_ & ~new_n4398_;
  assign new_n4400_ = ~new_n3632_ & ~new_n4399_;
  assign new_n4401_ = ~new_n4389_ & ~new_n4400_;
  assign \D_new<13>  = ~\reset<0>  & ~new_n4401_;
  assign new_n4403_ = ~new_n4338_ & ~new_n4376_;
  assign new_n4404_ = \encrypt_mode<0>  & ~new_n4403_;
  assign new_n4405_ = \D<11>  & ~new_n3665_;
  assign new_n4406_ = \D<10>  & new_n3665_;
  assign new_n4407_ = ~new_n4405_ & ~new_n4406_;
  assign new_n4408_ = ~\encrypt_mode<0>  & ~new_n4407_;
  assign new_n4409_ = ~new_n4404_ & ~new_n4408_;
  assign new_n4410_ = ~new_n3657_ & ~new_n4409_;
  assign new_n4411_ = \D<12>  & new_n3657_;
  assign new_n4412_ = ~new_n4410_ & ~new_n4411_;
  assign new_n4413_ = ~new_n3632_ & ~new_n4412_;
  assign new_n4414_ = \encrypt<0>  & \inreg<13> ;
  assign new_n4415_ = ~\encrypt<0>  & \inreg<21> ;
  assign new_n4416_ = ~new_n4414_ & ~new_n4415_;
  assign new_n4417_ = new_n3632_ & ~new_n4416_;
  assign new_n4418_ = ~new_n4413_ & ~new_n4417_;
  assign \D_new<12>  = ~\reset<0>  & ~new_n4418_;
  assign new_n4420_ = \encrypt<0>  & \inreg<21> ;
  assign new_n4421_ = ~\encrypt<0>  & \inreg<29> ;
  assign new_n4422_ = ~new_n4420_ & ~new_n4421_;
  assign new_n4423_ = new_n3632_ & ~new_n4422_;
  assign new_n4424_ = ~new_n4358_ & ~new_n4392_;
  assign new_n4425_ = \encrypt_mode<0>  & ~new_n4424_;
  assign new_n4426_ = \D<9>  & new_n3665_;
  assign new_n4427_ = \D<10>  & ~new_n3665_;
  assign new_n4428_ = ~new_n4426_ & ~new_n4427_;
  assign new_n4429_ = ~\encrypt_mode<0>  & ~new_n4428_;
  assign new_n4430_ = ~new_n4425_ & ~new_n4429_;
  assign new_n4431_ = ~new_n3657_ & ~new_n4430_;
  assign new_n4432_ = \D<11>  & new_n3657_;
  assign new_n4433_ = ~new_n4431_ & ~new_n4432_;
  assign new_n4434_ = ~new_n3632_ & ~new_n4433_;
  assign new_n4435_ = ~new_n4423_ & ~new_n4434_;
  assign \D_new<11>  = ~\reset<0>  & ~new_n4435_;
  assign new_n4437_ = \encrypt<0>  & \inreg<29> ;
  assign new_n4438_ = ~\encrypt<0>  & \inreg<37> ;
  assign new_n4439_ = ~new_n4437_ & ~new_n4438_;
  assign new_n4440_ = new_n3632_ & ~new_n4439_;
  assign new_n4441_ = ~new_n4375_ & ~new_n4405_;
  assign new_n4442_ = \encrypt_mode<0>  & ~new_n4441_;
  assign new_n4443_ = \D<9>  & ~new_n3665_;
  assign new_n4444_ = \D<8>  & new_n3665_;
  assign new_n4445_ = ~new_n4443_ & ~new_n4444_;
  assign new_n4446_ = ~\encrypt_mode<0>  & ~new_n4445_;
  assign new_n4447_ = ~new_n4442_ & ~new_n4446_;
  assign new_n4448_ = ~new_n3657_ & ~new_n4447_;
  assign new_n4449_ = \D<10>  & new_n3657_;
  assign new_n4450_ = ~new_n4448_ & ~new_n4449_;
  assign new_n4451_ = ~new_n3632_ & ~new_n4450_;
  assign new_n4452_ = ~new_n4440_ & ~new_n4451_;
  assign \D_new<10>  = ~\reset<0>  & ~new_n4452_;
  assign new_n4454_ = \encrypt<0>  & \inreg<37> ;
  assign new_n4455_ = ~\encrypt<0>  & \inreg<45> ;
  assign new_n4456_ = ~new_n4454_ & ~new_n4455_;
  assign new_n4457_ = new_n3632_ & ~new_n4456_;
  assign new_n4458_ = ~new_n4393_ & ~new_n4427_;
  assign new_n4459_ = \encrypt_mode<0>  & ~new_n4458_;
  assign new_n4460_ = \D<8>  & ~new_n3665_;
  assign new_n4461_ = \D<7>  & new_n3665_;
  assign new_n4462_ = ~new_n4460_ & ~new_n4461_;
  assign new_n4463_ = ~\encrypt_mode<0>  & ~new_n4462_;
  assign new_n4464_ = ~new_n4459_ & ~new_n4463_;
  assign new_n4465_ = ~new_n3657_ & ~new_n4464_;
  assign new_n4466_ = \D<9>  & new_n3657_;
  assign new_n4467_ = ~new_n4465_ & ~new_n4466_;
  assign new_n4468_ = ~new_n3632_ & ~new_n4467_;
  assign new_n4469_ = ~new_n4457_ & ~new_n4468_;
  assign \D_new<9>  = ~\reset<0>  & ~new_n4469_;
  assign new_n4471_ = \encrypt<0>  & \inreg<45> ;
  assign new_n4472_ = ~\encrypt<0>  & \inreg<53> ;
  assign new_n4473_ = ~new_n4471_ & ~new_n4472_;
  assign new_n4474_ = new_n3632_ & ~new_n4473_;
  assign new_n4475_ = ~new_n4406_ & ~new_n4443_;
  assign new_n4476_ = \encrypt_mode<0>  & ~new_n4475_;
  assign new_n4477_ = \D<7>  & ~new_n3665_;
  assign new_n4478_ = \D<6>  & new_n3665_;
  assign new_n4479_ = ~new_n4477_ & ~new_n4478_;
  assign new_n4480_ = ~\encrypt_mode<0>  & ~new_n4479_;
  assign new_n4481_ = ~new_n4476_ & ~new_n4480_;
  assign new_n4482_ = ~new_n3657_ & ~new_n4481_;
  assign new_n4483_ = \D<8>  & new_n3657_;
  assign new_n4484_ = ~new_n4482_ & ~new_n4483_;
  assign new_n4485_ = ~new_n3632_ & ~new_n4484_;
  assign new_n4486_ = ~new_n4474_ & ~new_n4485_;
  assign \D_new<8>  = ~\reset<0>  & ~new_n4486_;
  assign new_n4488_ = \data_in<6>  & ~\encrypt<0> ;
  assign new_n4489_ = \encrypt<0>  & \inreg<53> ;
  assign new_n4490_ = ~new_n4488_ & ~new_n4489_;
  assign new_n4491_ = new_n3632_ & ~new_n4490_;
  assign new_n4492_ = ~new_n4426_ & ~new_n4460_;
  assign new_n4493_ = \encrypt_mode<0>  & ~new_n4492_;
  assign new_n4494_ = \D<5>  & new_n3665_;
  assign new_n4495_ = \D<6>  & ~new_n3665_;
  assign new_n4496_ = ~new_n4494_ & ~new_n4495_;
  assign new_n4497_ = ~\encrypt_mode<0>  & ~new_n4496_;
  assign new_n4498_ = ~new_n4493_ & ~new_n4497_;
  assign new_n4499_ = ~new_n3657_ & ~new_n4498_;
  assign new_n4500_ = \D<7>  & new_n3657_;
  assign new_n4501_ = ~new_n4499_ & ~new_n4500_;
  assign new_n4502_ = ~new_n3632_ & ~new_n4501_;
  assign new_n4503_ = ~new_n4491_ & ~new_n4502_;
  assign \D_new<7>  = ~\reset<0>  & ~new_n4503_;
  assign new_n4505_ = \data_in<6>  & \encrypt<0> ;
  assign new_n4506_ = ~\encrypt<0>  & \inreg<6> ;
  assign new_n4507_ = ~new_n4505_ & ~new_n4506_;
  assign new_n4508_ = new_n3632_ & ~new_n4507_;
  assign new_n4509_ = ~new_n4444_ & ~new_n4477_;
  assign new_n4510_ = \encrypt_mode<0>  & ~new_n4509_;
  assign new_n4511_ = \D<4>  & new_n3665_;
  assign new_n4512_ = \D<5>  & ~new_n3665_;
  assign new_n4513_ = ~new_n4511_ & ~new_n4512_;
  assign new_n4514_ = ~\encrypt_mode<0>  & ~new_n4513_;
  assign new_n4515_ = ~new_n4510_ & ~new_n4514_;
  assign new_n4516_ = ~new_n3657_ & ~new_n4515_;
  assign new_n4517_ = \D<6>  & new_n3657_;
  assign new_n4518_ = ~new_n4516_ & ~new_n4517_;
  assign new_n4519_ = ~new_n3632_ & ~new_n4518_;
  assign new_n4520_ = ~new_n4508_ & ~new_n4519_;
  assign \D_new<6>  = ~\reset<0>  & ~new_n4520_;
  assign new_n4522_ = ~\encrypt<0>  & \inreg<14> ;
  assign new_n4523_ = \encrypt<0>  & \inreg<6> ;
  assign new_n4524_ = ~new_n4522_ & ~new_n4523_;
  assign new_n4525_ = new_n3632_ & ~new_n4524_;
  assign new_n4526_ = ~new_n4461_ & ~new_n4495_;
  assign new_n4527_ = \encrypt_mode<0>  & ~new_n4526_;
  assign new_n4528_ = \D<4>  & ~new_n3665_;
  assign new_n4529_ = \D<3>  & new_n3665_;
  assign new_n4530_ = ~new_n4528_ & ~new_n4529_;
  assign new_n4531_ = ~\encrypt_mode<0>  & ~new_n4530_;
  assign new_n4532_ = ~new_n4527_ & ~new_n4531_;
  assign new_n4533_ = ~new_n3657_ & ~new_n4532_;
  assign new_n4534_ = \D<5>  & new_n3657_;
  assign new_n4535_ = ~new_n4533_ & ~new_n4534_;
  assign new_n4536_ = ~new_n3632_ & ~new_n4535_;
  assign new_n4537_ = ~new_n4525_ & ~new_n4536_;
  assign \D_new<5>  = ~\reset<0>  & ~new_n4537_;
  assign new_n4539_ = ~new_n4478_ & ~new_n4512_;
  assign new_n4540_ = \encrypt_mode<0>  & ~new_n4539_;
  assign new_n4541_ = \D<3>  & ~new_n3665_;
  assign new_n4542_ = \D<2>  & new_n3665_;
  assign new_n4543_ = ~new_n4541_ & ~new_n4542_;
  assign new_n4544_ = ~\encrypt_mode<0>  & ~new_n4543_;
  assign new_n4545_ = ~new_n4540_ & ~new_n4544_;
  assign new_n4546_ = ~new_n3657_ & ~new_n4545_;
  assign new_n4547_ = \D<4>  & new_n3657_;
  assign new_n4548_ = ~new_n4546_ & ~new_n4547_;
  assign new_n4549_ = ~new_n3632_ & ~new_n4548_;
  assign new_n4550_ = \encrypt<0>  & \inreg<14> ;
  assign new_n4551_ = ~\encrypt<0>  & \inreg<22> ;
  assign new_n4552_ = ~new_n4550_ & ~new_n4551_;
  assign new_n4553_ = new_n3632_ & ~new_n4552_;
  assign new_n4554_ = ~new_n4549_ & ~new_n4553_;
  assign \D_new<4>  = ~\reset<0>  & ~new_n4554_;
  assign new_n4556_ = ~new_n4494_ & ~new_n4528_;
  assign new_n4557_ = \encrypt_mode<0>  & ~new_n4556_;
  assign new_n4558_ = \D<2>  & ~new_n3665_;
  assign new_n4559_ = ~new_n4147_ & ~new_n4558_;
  assign new_n4560_ = ~\encrypt_mode<0>  & ~new_n4559_;
  assign new_n4561_ = ~new_n4557_ & ~new_n4560_;
  assign new_n4562_ = ~new_n3657_ & ~new_n4561_;
  assign new_n4563_ = \D<3>  & new_n3657_;
  assign new_n4564_ = ~new_n4562_ & ~new_n4563_;
  assign new_n4565_ = ~new_n3632_ & ~new_n4564_;
  assign new_n4566_ = \encrypt<0>  & \inreg<22> ;
  assign new_n4567_ = ~\encrypt<0>  & \inreg<30> ;
  assign new_n4568_ = ~new_n4566_ & ~new_n4567_;
  assign new_n4569_ = new_n3632_ & ~new_n4568_;
  assign new_n4570_ = ~new_n4565_ & ~new_n4569_;
  assign \D_new<3>  = ~\reset<0>  & ~new_n4570_;
  assign new_n4572_ = ~new_n4511_ & ~new_n4541_;
  assign new_n4573_ = \encrypt_mode<0>  & ~new_n4572_;
  assign new_n4574_ = \D<1>  & ~new_n3665_;
  assign new_n4575_ = ~new_n4166_ & ~new_n4574_;
  assign new_n4576_ = ~\encrypt_mode<0>  & ~new_n4575_;
  assign new_n4577_ = ~new_n4573_ & ~new_n4576_;
  assign new_n4578_ = ~new_n3657_ & ~new_n4577_;
  assign new_n4579_ = \D<2>  & new_n3657_;
  assign new_n4580_ = ~new_n4578_ & ~new_n4579_;
  assign new_n4581_ = ~new_n3632_ & ~new_n4580_;
  assign new_n4582_ = \encrypt<0>  & \inreg<30> ;
  assign new_n4583_ = ~\encrypt<0>  & \inreg<38> ;
  assign new_n4584_ = ~new_n4582_ & ~new_n4583_;
  assign new_n4585_ = new_n3632_ & ~new_n4584_;
  assign new_n4586_ = ~new_n4581_ & ~new_n4585_;
  assign \D_new<2>  = ~\reset<0>  & ~new_n4586_;
  assign new_n4588_ = \encrypt<0>  & \inreg<38> ;
  assign new_n4589_ = ~\encrypt<0>  & \inreg<46> ;
  assign new_n4590_ = ~new_n4588_ & ~new_n4589_;
  assign new_n4591_ = new_n3632_ & ~new_n4590_;
  assign new_n4592_ = \D<1>  & new_n3657_;
  assign new_n4593_ = ~new_n4529_ & ~new_n4558_;
  assign new_n4594_ = \encrypt_mode<0>  & ~new_n4593_;
  assign new_n4595_ = ~new_n4146_ & ~new_n4184_;
  assign new_n4596_ = ~\encrypt_mode<0>  & ~new_n4595_;
  assign new_n4597_ = ~new_n4594_ & ~new_n4596_;
  assign new_n4598_ = ~new_n3657_ & ~new_n4597_;
  assign new_n4599_ = ~new_n4592_ & ~new_n4598_;
  assign new_n4600_ = ~new_n3632_ & ~new_n4599_;
  assign new_n4601_ = ~new_n4591_ & ~new_n4600_;
  assign \D_new<1>  = ~\reset<0>  & ~new_n4601_;
  assign new_n4603_ = \encrypt<0>  & \inreg<46> ;
  assign new_n4604_ = ~\encrypt<0>  & \inreg<54> ;
  assign new_n4605_ = ~new_n4603_ & ~new_n4604_;
  assign new_n4606_ = new_n3632_ & ~new_n4605_;
  assign new_n4607_ = \D<0>  & new_n3657_;
  assign new_n4608_ = ~new_n4165_ & ~new_n4198_;
  assign new_n4609_ = ~\encrypt_mode<0>  & ~new_n4608_;
  assign new_n4610_ = ~new_n4542_ & ~new_n4574_;
  assign new_n4611_ = \encrypt_mode<0>  & ~new_n4610_;
  assign new_n4612_ = ~new_n4609_ & ~new_n4611_;
  assign new_n4613_ = ~new_n3657_ & ~new_n4612_;
  assign new_n4614_ = ~new_n4607_ & ~new_n4613_;
  assign new_n4615_ = ~new_n3632_ & ~new_n4614_;
  assign new_n4616_ = ~new_n4606_ & ~new_n4615_;
  assign \D_new<0>  = ~\reset<0>  & ~new_n4616_;
  assign new_n4618_ = \count<3>  & \count<2> ;
  assign new_n4619_ = new_n502_ & new_n4618_;
  assign new_n4620_ = \encrypt_mode<0>  & ~new_n4619_;
  assign new_n4621_ = \count<1>  & new_n4618_;
  assign new_n4622_ = \encrypt<0>  & \count<0> ;
  assign new_n4623_ = new_n4621_ & new_n4622_;
  assign \encrypt_mode_new<0>  = new_n4620_ | new_n4623_;
endmodule

