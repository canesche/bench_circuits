module top ( 
    pp, pa0, pq, pb0, pr, pc0, ps, pt, pu, pv, pw, px, py, pz, pa, pb, pc,
    pe, pf, pg, ph, pi, pj, pk, pl, pm, pn, po,
    pd0, pe0, pf0  );
  input  pp, pa0, pq, pb0, pr, pc0, ps, pt, pu, pv, pw, px, py, pz, pa,
    pb, pc, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn, po;
  output pd0, pe0, pf0;
  wire new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_, new_n38_,
    new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_, new_n45_,
    new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_,
    new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_,
    new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_,
    new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_,
    new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_;
  assign new_n32_ = pe & ~pi;
  assign new_n33_ = ~pj & new_n32_;
  assign new_n34_ = ~pc & new_n33_;
  assign new_n35_ = ~pi & ~pj;
  assign new_n36_ = pa & new_n35_;
  assign new_n37_ = ~pc & new_n36_;
  assign new_n38_ = ~pq & ~pv;
  assign new_n39_ = pe & new_n38_;
  assign new_n40_ = ~pr & new_n39_;
  assign new_n41_ = ~pc & new_n40_;
  assign new_n42_ = ~pm & new_n41_;
  assign new_n43_ = ~pu & new_n42_;
  assign new_n44_ = ~ps & new_n43_;
  assign new_n45_ = ~pt & new_n44_;
  assign new_n46_ = ~po & new_n45_;
  assign new_n47_ = ~pp & new_n46_;
  assign new_n48_ = pe & ~pg;
  assign new_n49_ = ~ph & new_n48_;
  assign new_n50_ = ~pc & new_n49_;
  assign new_n51_ = ~pq & pa;
  assign new_n52_ = ~pr & new_n51_;
  assign new_n53_ = ~pv & new_n52_;
  assign new_n54_ = ~pc & new_n53_;
  assign new_n55_ = ~pm & new_n54_;
  assign new_n56_ = ~pu & new_n55_;
  assign new_n57_ = ~ps & new_n56_;
  assign new_n58_ = ~pt & new_n57_;
  assign new_n59_ = ~po & new_n58_;
  assign new_n60_ = ~pp & new_n59_;
  assign new_n61_ = pa & ~ph;
  assign new_n62_ = ~pg & new_n61_;
  assign new_n63_ = ~pc & new_n62_;
  assign new_n64_ = ~pz & ~pk;
  assign new_n65_ = pe & new_n64_;
  assign new_n66_ = ~pr & new_n65_;
  assign new_n67_ = ~pc & new_n66_;
  assign new_n68_ = ~px & new_n67_;
  assign new_n69_ = ~pw & new_n68_;
  assign new_n70_ = ~po & new_n69_;
  assign new_n71_ = ~pp & new_n70_;
  assign new_n72_ = ~pq & new_n71_;
  assign new_n73_ = ~py & new_n72_;
  assign new_n74_ = ~pq & ~pk;
  assign new_n75_ = ~pr & new_n74_;
  assign new_n76_ = ~pz & new_n75_;
  assign new_n77_ = ~pc & new_n76_;
  assign new_n78_ = ~px & new_n77_;
  assign new_n79_ = ~pw & new_n78_;
  assign new_n80_ = ~po & new_n79_;
  assign new_n81_ = ~pp & new_n80_;
  assign new_n82_ = ~py & new_n81_;
  assign new_n83_ = pa & new_n82_;
  assign new_n84_ = ~pb & pc;
  assign new_n85_ = ~pr & ~pv;
  assign new_n86_ = pe & new_n85_;
  assign new_n87_ = ~ph & new_n86_;
  assign new_n88_ = ~pc & new_n87_;
  assign new_n89_ = ~px & new_n88_;
  assign new_n90_ = ~ps & new_n89_;
  assign new_n91_ = ~pt & new_n90_;
  assign new_n92_ = ~pz & new_n91_;
  assign new_n93_ = ~pp & new_n92_;
  assign new_n94_ = ~pv & ~pz;
  assign new_n95_ = ~ph & new_n94_;
  assign new_n96_ = ~pr & new_n95_;
  assign new_n97_ = ~pc & new_n96_;
  assign new_n98_ = ~px & new_n97_;
  assign new_n99_ = ~ps & new_n98_;
  assign new_n100_ = ~pt & new_n99_;
  assign new_n101_ = pa & new_n100_;
  assign new_n102_ = ~pp & new_n101_;
  assign new_n103_ = ~pp & ~ps;
  assign new_n104_ = pe & new_n103_;
  assign new_n105_ = ~po & new_n104_;
  assign new_n106_ = ~pc & new_n105_;
  assign new_n107_ = ~px & new_n106_;
  assign new_n108_ = ~pi & new_n107_;
  assign new_n109_ = ~pt & new_n108_;
  assign new_n110_ = ~pw & new_n109_;
  assign new_n111_ = ~pq & ~py;
  assign new_n112_ = ~pj & new_n111_;
  assign new_n113_ = ~pg & new_n112_;
  assign new_n114_ = ~pc & new_n113_;
  assign new_n115_ = pa & new_n114_;
  assign new_n116_ = ~pu & new_n115_;
  assign new_n117_ = ~px & ~pi;
  assign new_n118_ = pe & new_n117_;
  assign new_n119_ = ~ph & new_n118_;
  assign new_n120_ = ~pc & new_n119_;
  assign new_n121_ = ~pn & new_n120_;
  assign new_n122_ = ~py & ~pz;
  assign new_n123_ = pe & new_n122_;
  assign new_n124_ = ~pj & new_n123_;
  assign new_n125_ = ~pc & new_n124_;
  assign new_n126_ = ~pn & new_n125_;
  assign new_n127_ = ~pw & ~po;
  assign new_n128_ = pe & new_n127_;
  assign new_n129_ = ~pg & new_n128_;
  assign new_n130_ = ~pc & new_n129_;
  assign new_n131_ = ~pi & new_n130_;
  assign new_n132_ = pa & new_n103_;
  assign new_n133_ = ~po & new_n132_;
  assign new_n134_ = ~pc & new_n133_;
  assign new_n135_ = ~px & new_n134_;
  assign new_n136_ = ~pi & new_n135_;
  assign new_n137_ = ~pt & new_n136_;
  assign new_n138_ = ~pw & new_n137_;
  assign new_n139_ = ~pq & ~pg;
  assign new_n140_ = pe & new_n139_;
  assign new_n141_ = ~pj & new_n140_;
  assign new_n142_ = ~pc & new_n141_;
  assign new_n143_ = ~py & new_n142_;
  assign new_n144_ = ~pu & new_n143_;
  assign new_n145_ = ~ph & new_n117_;
  assign new_n146_ = pa & new_n145_;
  assign new_n147_ = ~pc & new_n146_;
  assign new_n148_ = ~pn & new_n147_;
  assign new_n149_ = ~pz & ~pj;
  assign new_n150_ = pe & new_n149_;
  assign new_n151_ = ~ph & new_n150_;
  assign new_n152_ = ~pc & new_n151_;
  assign new_n153_ = ~pn & new_n152_;
  assign new_n154_ = ~pg & new_n127_;
  assign new_n155_ = pa & new_n154_;
  assign new_n156_ = ~pc & new_n155_;
  assign new_n157_ = ~pi & new_n156_;
  assign new_n158_ = ~pq & ~pz;
  assign new_n159_ = ~pr & new_n158_;
  assign new_n160_ = ~pv & new_n159_;
  assign new_n161_ = ~pc & new_n160_;
  assign new_n162_ = ~pw & new_n161_;
  assign new_n163_ = ~px & new_n162_;
  assign new_n164_ = ~pt & new_n163_;
  assign new_n165_ = ~pu & new_n164_;
  assign new_n166_ = ~ps & new_n165_;
  assign new_n167_ = ~po & new_n166_;
  assign new_n168_ = ~pp & new_n167_;
  assign new_n169_ = ~py & new_n168_;
  assign new_n170_ = pa & new_n169_;
  assign new_n171_ = ~pt & new_n88_;
  assign new_n172_ = ~pm & new_n171_;
  assign new_n173_ = ~pp & new_n172_;
  assign new_n174_ = ~ps & new_n173_;
  assign new_n175_ = ~ph & new_n104_;
  assign new_n176_ = ~pc & new_n175_;
  assign new_n177_ = ~pi & new_n176_;
  assign new_n178_ = ~pt & new_n177_;
  assign new_n179_ = ~px & new_n178_;
  assign new_n180_ = ~pj & new_n74_;
  assign new_n181_ = ~pg & new_n180_;
  assign new_n182_ = ~pc & new_n181_;
  assign new_n183_ = ~py & new_n182_;
  assign new_n184_ = pa & new_n183_;
  assign new_n185_ = ~pw & ~pi;
  assign new_n186_ = pe & new_n185_;
  assign new_n187_ = ~pg & new_n186_;
  assign new_n188_ = ~pc & new_n187_;
  assign new_n189_ = ~pn & new_n188_;
  assign new_n190_ = ~pz & pa;
  assign new_n191_ = ~ph & new_n190_;
  assign new_n192_ = ~pj & new_n191_;
  assign new_n193_ = ~pc & new_n192_;
  assign new_n194_ = ~pn & new_n193_;
  assign new_n195_ = ~pm & ~po;
  assign new_n196_ = pe & new_n195_;
  assign new_n197_ = ~pg & new_n196_;
  assign new_n198_ = ~pc & new_n197_;
  assign new_n199_ = ~pi & new_n198_;
  assign new_n200_ = pe & new_n94_;
  assign new_n201_ = ~pr & new_n200_;
  assign new_n202_ = ~pc & new_n201_;
  assign new_n203_ = ~pw & new_n202_;
  assign new_n204_ = ~px & new_n203_;
  assign new_n205_ = ~pt & new_n204_;
  assign new_n206_ = ~pu & new_n205_;
  assign new_n207_ = ~ps & new_n206_;
  assign new_n208_ = ~po & new_n207_;
  assign new_n209_ = ~pp & new_n208_;
  assign new_n210_ = ~pq & new_n209_;
  assign new_n211_ = ~py & new_n210_;
  assign new_n212_ = ~pv & pa;
  assign new_n213_ = ~ph & new_n212_;
  assign new_n214_ = ~pr & new_n213_;
  assign new_n215_ = ~pc & new_n214_;
  assign new_n216_ = ~pt & new_n215_;
  assign new_n217_ = ~pm & new_n216_;
  assign new_n218_ = ~pp & new_n217_;
  assign new_n219_ = ~ps & new_n218_;
  assign new_n220_ = ~ph & new_n103_;
  assign new_n221_ = pa & new_n220_;
  assign new_n222_ = ~pc & new_n221_;
  assign new_n223_ = ~pi & new_n222_;
  assign new_n224_ = ~pt & new_n223_;
  assign new_n225_ = ~px & new_n224_;
  assign new_n226_ = ~pr & ~pz;
  assign new_n227_ = ~ph & new_n226_;
  assign new_n228_ = ~pj & new_n227_;
  assign new_n229_ = ~pc & new_n228_;
  assign new_n230_ = ~pk & new_n229_;
  assign new_n231_ = pa & new_n230_;
  assign new_n232_ = ~pg & new_n185_;
  assign new_n233_ = pa & new_n232_;
  assign new_n234_ = ~pc & new_n233_;
  assign new_n235_ = ~pn & new_n234_;
  assign new_n236_ = ~py & ~pg;
  assign new_n237_ = pe & new_n236_;
  assign new_n238_ = ~pj & new_n237_;
  assign new_n239_ = ~pc & new_n238_;
  assign new_n240_ = ~pn & new_n239_;
  assign new_n241_ = ~pg & new_n195_;
  assign new_n242_ = pa & new_n241_;
  assign new_n243_ = ~pc & new_n242_;
  assign new_n244_ = ~pi & new_n243_;
  assign new_n245_ = ~pg & new_n111_;
  assign new_n246_ = ~pk & new_n245_;
  assign new_n247_ = ~pc & new_n246_;
  assign new_n248_ = ~pw & new_n247_;
  assign new_n249_ = pa & new_n248_;
  assign new_n250_ = ~po & new_n249_;
  assign new_n251_ = ~pp & ~po;
  assign new_n252_ = pe & new_n251_;
  assign new_n253_ = ~pk & new_n252_;
  assign new_n254_ = ~pc & new_n253_;
  assign new_n255_ = ~pm & new_n254_;
  assign new_n256_ = ~pi & new_n255_;
  assign new_n257_ = ~ph & new_n85_;
  assign new_n258_ = ~pj & new_n257_;
  assign new_n259_ = ~pc & new_n258_;
  assign new_n260_ = ~pz & new_n259_;
  assign new_n261_ = pa & new_n260_;
  assign new_n262_ = ~px & ~pz;
  assign new_n263_ = pe & new_n262_;
  assign new_n264_ = ~ph & new_n263_;
  assign new_n265_ = ~pc & new_n264_;
  assign new_n266_ = ~pn & new_n265_;
  assign new_n267_ = ~pu & pa;
  assign new_n268_ = ~pj & new_n267_;
  assign new_n269_ = ~pv & new_n268_;
  assign new_n270_ = ~pc & new_n269_;
  assign new_n271_ = ~pl & new_n270_;
  assign new_n272_ = ~pu & ~pl;
  assign new_n273_ = pe & new_n272_;
  assign new_n274_ = ~pg & new_n273_;
  assign new_n275_ = ~pc & new_n274_;
  assign new_n276_ = pe & new_n74_;
  assign new_n277_ = ~pg & new_n276_;
  assign new_n278_ = ~pc & new_n277_;
  assign new_n279_ = ~pw & new_n278_;
  assign new_n280_ = ~py & new_n279_;
  assign new_n281_ = ~po & new_n280_;
  assign new_n282_ = ~pk & new_n251_;
  assign new_n283_ = pa & new_n282_;
  assign new_n284_ = ~pc & new_n283_;
  assign new_n285_ = ~pm & new_n284_;
  assign new_n286_ = ~pi & new_n285_;
  assign new_n287_ = ~pg & ~pk;
  assign new_n288_ = pe & new_n287_;
  assign new_n289_ = ~pj & new_n288_;
  assign new_n290_ = ~pc & new_n289_;
  assign new_n291_ = ~pq & new_n290_;
  assign new_n292_ = ~py & new_n291_;
  assign new_n293_ = ~px & pa;
  assign new_n294_ = ~ph & new_n293_;
  assign new_n295_ = ~pz & new_n294_;
  assign new_n296_ = ~pc & new_n295_;
  assign new_n297_ = ~pn & new_n296_;
  assign new_n298_ = ~pu & ~pv;
  assign new_n299_ = pe & new_n298_;
  assign new_n300_ = ~pj & new_n299_;
  assign new_n301_ = ~pc & new_n300_;
  assign new_n302_ = ~pl & new_n301_;
  assign new_n303_ = ~pg & new_n272_;
  assign new_n304_ = pa & new_n303_;
  assign new_n305_ = ~pc & new_n304_;
  assign new_n306_ = pa & ~pk;
  assign new_n307_ = ~ph & new_n306_;
  assign new_n308_ = ~pr & new_n307_;
  assign new_n309_ = ~pc & new_n308_;
  assign new_n310_ = ~pp & new_n309_;
  assign new_n311_ = ~pm & new_n310_;
  assign new_n312_ = ~pr & ~pj;
  assign new_n313_ = pe & new_n312_;
  assign new_n314_ = ~ph & new_n313_;
  assign new_n315_ = ~pc & new_n314_;
  assign new_n316_ = ~pv & new_n315_;
  assign new_n317_ = ~pm & new_n316_;
  assign new_n318_ = ~pz & new_n315_;
  assign new_n319_ = ~pk & new_n318_;
  assign new_n320_ = ~pw & ~py;
  assign new_n321_ = pe & new_n320_;
  assign new_n322_ = ~pg & new_n321_;
  assign new_n323_ = ~pc & new_n322_;
  assign new_n324_ = ~pn & new_n323_;
  assign new_n325_ = ~pt & ~pi;
  assign new_n326_ = pa & new_n325_;
  assign new_n327_ = ~ps & new_n326_;
  assign new_n328_ = ~pc & new_n327_;
  assign new_n329_ = ~pl & new_n328_;
  assign new_n330_ = ~pi & ~pl;
  assign new_n331_ = pe & new_n330_;
  assign new_n332_ = ~pg & new_n331_;
  assign new_n333_ = ~pc & new_n332_;
  assign new_n334_ = ~pr & ~pk;
  assign new_n335_ = pe & new_n334_;
  assign new_n336_ = ~ph & new_n335_;
  assign new_n337_ = ~pc & new_n336_;
  assign new_n338_ = ~pp & new_n337_;
  assign new_n339_ = ~pm & new_n338_;
  assign new_n340_ = ~pk & new_n315_;
  assign new_n341_ = ~pm & new_n340_;
  assign new_n342_ = ~pz & new_n316_;
  assign new_n343_ = ~pw & pa;
  assign new_n344_ = ~pg & new_n343_;
  assign new_n345_ = ~py & new_n344_;
  assign new_n346_ = ~pc & new_n345_;
  assign new_n347_ = ~pn & new_n346_;
  assign new_n348_ = pe & new_n325_;
  assign new_n349_ = ~ps & new_n348_;
  assign new_n350_ = ~pc & new_n349_;
  assign new_n351_ = ~pl & new_n350_;
  assign new_n352_ = ~pg & new_n330_;
  assign new_n353_ = pa & new_n352_;
  assign new_n354_ = ~pc & new_n353_;
  assign new_n355_ = ~pi & new_n106_;
  assign new_n356_ = ~pt & new_n355_;
  assign new_n357_ = ~pm & new_n356_;
  assign new_n358_ = ~ph & new_n64_;
  assign new_n359_ = ~pr & new_n358_;
  assign new_n360_ = ~pc & new_n359_;
  assign new_n361_ = ~px & new_n360_;
  assign new_n362_ = pa & new_n361_;
  assign new_n363_ = ~pp & new_n362_;
  assign new_n364_ = ~ps & ~pt;
  assign new_n365_ = pe & new_n364_;
  assign new_n366_ = ~pv & new_n365_;
  assign new_n367_ = ~pc & new_n366_;
  assign new_n368_ = ~pu & new_n367_;
  assign new_n369_ = ~pl & new_n368_;
  assign new_n370_ = ~pj & new_n51_;
  assign new_n371_ = ~pg & new_n370_;
  assign new_n372_ = ~pc & new_n371_;
  assign new_n373_ = ~pu & new_n372_;
  assign new_n374_ = ~pm & new_n373_;
  assign new_n375_ = ~pj & new_n335_;
  assign new_n376_ = ~pc & new_n375_;
  assign new_n377_ = ~pq & new_n376_;
  assign new_n378_ = ~pm & new_n377_;
  assign new_n379_ = pa & new_n117_;
  assign new_n380_ = ~pw & new_n379_;
  assign new_n381_ = ~pc & new_n380_;
  assign new_n382_ = ~pn & new_n381_;
  assign new_n383_ = ~py & pa;
  assign new_n384_ = ~pj & new_n383_;
  assign new_n385_ = ~pz & new_n384_;
  assign new_n386_ = ~pc & new_n385_;
  assign new_n387_ = ~pn & new_n386_;
  assign new_n388_ = ~pi & new_n134_;
  assign new_n389_ = ~pt & new_n388_;
  assign new_n390_ = ~pm & new_n389_;
  assign new_n391_ = pe & new_n226_;
  assign new_n392_ = ~ph & new_n391_;
  assign new_n393_ = ~pc & new_n392_;
  assign new_n394_ = ~px & new_n393_;
  assign new_n395_ = ~pk & new_n394_;
  assign new_n396_ = ~pp & new_n395_;
  assign new_n397_ = ~pv & new_n364_;
  assign new_n398_ = pa & new_n397_;
  assign new_n399_ = ~pc & new_n398_;
  assign new_n400_ = ~pu & new_n399_;
  assign new_n401_ = ~pl & new_n400_;
  assign new_n402_ = ~pu & new_n142_;
  assign new_n403_ = ~pm & new_n402_;
  assign new_n404_ = ~pm & new_n291_;
  assign new_n405_ = ~pw & new_n118_;
  assign new_n406_ = ~pc & new_n405_;
  assign new_n407_ = ~pn & new_n406_;
  assign new_n408_ = ~pg & new_n384_;
  assign new_n409_ = ~pc & new_n408_;
  assign new_n410_ = ~pn & new_n409_;
  assign new_n411_ = ~pj & new_n86_;
  assign new_n412_ = ~pc & new_n411_;
  assign new_n413_ = ~py & new_n412_;
  assign new_n414_ = ~pu & new_n413_;
  assign new_n415_ = ~pz & new_n414_;
  assign new_n416_ = ~pq & new_n415_;
  assign new_n417_ = ~pg & new_n383_;
  assign new_n418_ = ~pq & new_n417_;
  assign new_n419_ = ~pc & new_n418_;
  assign new_n420_ = ~pw & new_n419_;
  assign new_n421_ = ~po & new_n420_;
  assign new_n422_ = ~pu & new_n421_;
  assign new_n423_ = ~ps & ~pv;
  assign new_n424_ = pe & new_n423_;
  assign new_n425_ = ~ph & new_n424_;
  assign new_n426_ = ~pc & new_n425_;
  assign new_n427_ = ~pt & new_n426_;
  assign new_n428_ = ~pl & new_n427_;
  assign new_n429_ = pa & ~po;
  assign new_n430_ = ~pg & new_n429_;
  assign new_n431_ = ~pq & new_n430_;
  assign new_n432_ = ~pc & new_n431_;
  assign new_n433_ = ~pu & new_n432_;
  assign new_n434_ = ~pm & new_n433_;
  assign new_n435_ = pa & new_n259_;
  assign new_n436_ = ~pm & new_n435_;
  assign new_n437_ = ~pj & new_n213_;
  assign new_n438_ = ~pc & new_n437_;
  assign new_n439_ = ~pl & new_n438_;
  assign new_n440_ = pa & ~pn;
  assign new_n441_ = ~pl & new_n440_;
  assign new_n442_ = ~pc & new_n441_;
  assign new_n443_ = ~pj & new_n94_;
  assign new_n444_ = ~pr & new_n443_;
  assign new_n445_ = ~pc & new_n444_;
  assign new_n446_ = pa & new_n445_;
  assign new_n447_ = ~pu & new_n446_;
  assign new_n448_ = ~pq & new_n447_;
  assign new_n449_ = ~py & new_n448_;
  assign new_n450_ = pe & new_n111_;
  assign new_n451_ = ~pg & new_n450_;
  assign new_n452_ = ~pc & new_n451_;
  assign new_n453_ = ~pw & new_n452_;
  assign new_n454_ = ~po & new_n453_;
  assign new_n455_ = ~pu & new_n454_;
  assign new_n456_ = ~ps & pa;
  assign new_n457_ = ~ph & new_n456_;
  assign new_n458_ = ~pv & new_n457_;
  assign new_n459_ = ~pc & new_n458_;
  assign new_n460_ = ~pt & new_n459_;
  assign new_n461_ = ~pl & new_n460_;
  assign new_n462_ = ~pq & ~po;
  assign new_n463_ = pe & new_n462_;
  assign new_n464_ = ~pg & new_n463_;
  assign new_n465_ = ~pc & new_n464_;
  assign new_n466_ = ~pu & new_n465_;
  assign new_n467_ = ~pm & new_n466_;
  assign new_n468_ = ~ph & new_n334_;
  assign new_n469_ = ~pj & new_n468_;
  assign new_n470_ = ~pc & new_n469_;
  assign new_n471_ = pa & new_n470_;
  assign new_n472_ = ~pm & new_n471_;
  assign new_n473_ = ~pv & ~pj;
  assign new_n474_ = pe & new_n473_;
  assign new_n475_ = ~ph & new_n474_;
  assign new_n476_ = ~pc & new_n475_;
  assign new_n477_ = ~pl & new_n476_;
  assign new_n478_ = ~pc0 & ~pe;
  assign new_n479_ = ~pa & new_n478_;
  assign new_n480_ = ~pc & new_n479_;
  assign new_n481_ = ~pi & new_n254_;
  assign new_n482_ = ~pw & new_n481_;
  assign new_n483_ = ~px & new_n482_;
  assign new_n484_ = ~pj & new_n38_;
  assign new_n485_ = ~pr & new_n484_;
  assign new_n486_ = ~pc & new_n485_;
  assign new_n487_ = ~pm & new_n486_;
  assign new_n488_ = pa & new_n487_;
  assign new_n489_ = ~pu & new_n488_;
  assign new_n490_ = ~pj & new_n391_;
  assign new_n491_ = ~pc & new_n490_;
  assign new_n492_ = ~py & new_n491_;
  assign new_n493_ = ~pk & new_n492_;
  assign new_n494_ = ~pq & new_n493_;
  assign new_n495_ = ~pp & pa;
  assign new_n496_ = ~ph & new_n495_;
  assign new_n497_ = ~pk & new_n496_;
  assign new_n498_ = ~pc & new_n497_;
  assign new_n499_ = ~px & new_n498_;
  assign new_n500_ = ~pi & new_n499_;
  assign new_n501_ = ~pr & new_n180_;
  assign new_n502_ = ~pc & new_n501_;
  assign new_n503_ = pa & new_n502_;
  assign new_n504_ = ~pm & new_n503_;
  assign new_n505_ = ~pi & new_n284_;
  assign new_n506_ = ~pw & new_n505_;
  assign new_n507_ = ~px & new_n506_;
  assign new_n508_ = ~pm & new_n412_;
  assign new_n509_ = ~pq & new_n508_;
  assign new_n510_ = ~pu & new_n509_;
  assign new_n511_ = ~pj & new_n64_;
  assign new_n512_ = ~pr & new_n511_;
  assign new_n513_ = ~pc & new_n512_;
  assign new_n514_ = pa & new_n513_;
  assign new_n515_ = ~pq & new_n514_;
  assign new_n516_ = ~py & new_n515_;
  assign new_n517_ = ~pp & ~pk;
  assign new_n518_ = pe & new_n517_;
  assign new_n519_ = ~ph & new_n518_;
  assign new_n520_ = ~pc & new_n519_;
  assign new_n521_ = ~px & new_n520_;
  assign new_n522_ = ~pi & new_n521_;
  assign new_n523_ = pa & new_n182_;
  assign new_n524_ = ~pm & new_n523_;
  assign new_n525_ = ~pm & new_n178_;
  assign new_n526_ = ~pk & new_n52_;
  assign new_n527_ = ~pc & new_n526_;
  assign new_n528_ = ~pm & new_n527_;
  assign new_n529_ = ~po & new_n528_;
  assign new_n530_ = ~pp & new_n529_;
  assign new_n531_ = ~pz & new_n321_;
  assign new_n532_ = ~pc & new_n531_;
  assign new_n533_ = ~px & new_n532_;
  assign new_n534_ = ~pn & new_n533_;
  assign new_n535_ = ~pm & new_n498_;
  assign new_n536_ = ~pi & new_n535_;
  assign new_n537_ = ~po & new_n278_;
  assign new_n538_ = ~pm & new_n537_;
  assign new_n539_ = ~pm & new_n224_;
  assign new_n540_ = ~pr & new_n276_;
  assign new_n541_ = ~pc & new_n540_;
  assign new_n542_ = ~pm & new_n541_;
  assign new_n543_ = ~po & new_n542_;
  assign new_n544_ = ~pp & new_n543_;
  assign new_n545_ = ~pz & new_n343_;
  assign new_n546_ = ~py & new_n545_;
  assign new_n547_ = ~pc & new_n546_;
  assign new_n548_ = ~px & new_n547_;
  assign new_n549_ = ~pn & new_n548_;
  assign new_n550_ = ~pm & new_n520_;
  assign new_n551_ = ~pi & new_n550_;
  assign new_n552_ = ~pg & new_n51_;
  assign new_n553_ = ~pk & new_n552_;
  assign new_n554_ = ~pc & new_n553_;
  assign new_n555_ = ~po & new_n554_;
  assign new_n556_ = ~pm & new_n555_;
  assign new_n557_ = pe & ~pn;
  assign new_n558_ = ~pl & new_n557_;
  assign new_n559_ = ~pc & new_n558_;
  assign new_n560_ = ~pm & new_n557_;
  assign new_n561_ = ~pc & new_n560_;
  assign new_n562_ = ~pm & new_n440_;
  assign new_n563_ = ~pc & new_n562_;
  assign new_n564_ = pe & ~pl;
  assign new_n565_ = ~pk & new_n564_;
  assign new_n566_ = ~pc & new_n565_;
  assign new_n567_ = ~pk & ~pl;
  assign new_n568_ = pa & new_n567_;
  assign new_n569_ = ~pc & new_n568_;
  assign new_n570_ = ~new_n563_ & ~new_n566_;
  assign new_n571_ = ~new_n569_ & new_n570_;
  assign new_n572_ = ~new_n559_ & ~new_n561_;
  assign new_n573_ = ~new_n551_ & ~new_n556_;
  assign new_n574_ = new_n572_ & new_n573_;
  assign new_n575_ = new_n571_ & new_n574_;
  assign new_n576_ = ~new_n539_ & ~new_n544_;
  assign new_n577_ = ~new_n549_ & new_n576_;
  assign new_n578_ = ~new_n536_ & ~new_n538_;
  assign new_n579_ = ~new_n530_ & ~new_n534_;
  assign new_n580_ = new_n578_ & new_n579_;
  assign new_n581_ = new_n577_ & new_n580_;
  assign new_n582_ = new_n575_ & new_n581_;
  assign new_n583_ = ~new_n522_ & ~new_n524_;
  assign new_n584_ = ~new_n525_ & new_n583_;
  assign new_n585_ = ~new_n510_ & ~new_n516_;
  assign new_n586_ = ~new_n504_ & ~new_n507_;
  assign new_n587_ = new_n585_ & new_n586_;
  assign new_n588_ = new_n584_ & new_n587_;
  assign new_n589_ = ~new_n489_ & ~new_n494_;
  assign new_n590_ = ~new_n500_ & new_n589_;
  assign new_n591_ = ~new_n480_ & ~new_n483_;
  assign new_n592_ = ~new_n472_ & ~new_n477_;
  assign new_n593_ = new_n591_ & new_n592_;
  assign new_n594_ = new_n590_ & new_n593_;
  assign new_n595_ = new_n588_ & new_n594_;
  assign new_n596_ = new_n582_ & new_n595_;
  assign new_n597_ = ~new_n455_ & ~new_n461_;
  assign new_n598_ = ~new_n467_ & new_n597_;
  assign new_n599_ = ~new_n442_ & ~new_n449_;
  assign new_n600_ = ~new_n436_ & ~new_n439_;
  assign new_n601_ = new_n599_ & new_n600_;
  assign new_n602_ = new_n598_ & new_n601_;
  assign new_n603_ = ~new_n422_ & ~new_n428_;
  assign new_n604_ = ~new_n434_ & new_n603_;
  assign new_n605_ = ~new_n410_ & ~new_n416_;
  assign new_n606_ = ~new_n404_ & ~new_n407_;
  assign new_n607_ = new_n605_ & new_n606_;
  assign new_n608_ = new_n604_ & new_n607_;
  assign new_n609_ = new_n602_ & new_n608_;
  assign new_n610_ = ~new_n396_ & ~new_n401_;
  assign new_n611_ = ~new_n403_ & new_n610_;
  assign new_n612_ = ~new_n387_ & ~new_n390_;
  assign new_n613_ = ~new_n378_ & ~new_n382_;
  assign new_n614_ = new_n612_ & new_n613_;
  assign new_n615_ = new_n611_ & new_n614_;
  assign new_n616_ = ~new_n363_ & ~new_n369_;
  assign new_n617_ = ~new_n374_ & new_n616_;
  assign new_n618_ = ~new_n354_ & ~new_n357_;
  assign new_n619_ = ~new_n347_ & ~new_n351_;
  assign new_n620_ = new_n618_ & new_n619_;
  assign new_n621_ = new_n617_ & new_n620_;
  assign new_n622_ = new_n615_ & new_n621_;
  assign new_n623_ = new_n609_ & new_n622_;
  assign new_n624_ = new_n596_ & new_n623_;
  assign new_n625_ = ~new_n339_ & ~new_n341_;
  assign new_n626_ = ~new_n342_ & new_n625_;
  assign new_n627_ = ~new_n329_ & ~new_n333_;
  assign new_n628_ = ~new_n319_ & ~new_n324_;
  assign new_n629_ = new_n627_ & new_n628_;
  assign new_n630_ = new_n626_ & new_n629_;
  assign new_n631_ = ~new_n305_ & ~new_n311_;
  assign new_n632_ = ~new_n317_ & new_n631_;
  assign new_n633_ = ~new_n297_ & ~new_n302_;
  assign new_n634_ = ~new_n286_ & ~new_n292_;
  assign new_n635_ = new_n633_ & new_n634_;
  assign new_n636_ = new_n632_ & new_n635_;
  assign new_n637_ = new_n630_ & new_n636_;
  assign new_n638_ = ~new_n271_ & ~new_n275_;
  assign new_n639_ = ~new_n281_ & new_n638_;
  assign new_n640_ = ~new_n261_ & ~new_n266_;
  assign new_n641_ = ~new_n250_ & ~new_n256_;
  assign new_n642_ = new_n640_ & new_n641_;
  assign new_n643_ = new_n639_ & new_n642_;
  assign new_n644_ = ~new_n235_ & ~new_n240_;
  assign new_n645_ = ~new_n244_ & new_n644_;
  assign new_n646_ = ~new_n225_ & ~new_n231_;
  assign new_n647_ = ~new_n211_ & ~new_n219_;
  assign new_n648_ = new_n646_ & new_n647_;
  assign new_n649_ = new_n645_ & new_n648_;
  assign new_n650_ = new_n643_ & new_n649_;
  assign new_n651_ = new_n637_ & new_n650_;
  assign new_n652_ = ~new_n189_ & ~new_n194_;
  assign new_n653_ = ~new_n199_ & new_n652_;
  assign new_n654_ = ~new_n179_ & ~new_n184_;
  assign new_n655_ = ~new_n170_ & ~new_n174_;
  assign new_n656_ = new_n654_ & new_n655_;
  assign new_n657_ = new_n653_ & new_n656_;
  assign new_n658_ = ~new_n148_ & ~new_n153_;
  assign new_n659_ = ~new_n157_ & new_n658_;
  assign new_n660_ = ~new_n138_ & ~new_n144_;
  assign new_n661_ = ~new_n126_ & ~new_n131_;
  assign new_n662_ = new_n660_ & new_n661_;
  assign new_n663_ = new_n659_ & new_n662_;
  assign new_n664_ = new_n657_ & new_n663_;
  assign new_n665_ = ~new_n110_ & ~new_n116_;
  assign new_n666_ = ~new_n121_ & new_n665_;
  assign new_n667_ = ~new_n93_ & ~new_n102_;
  assign new_n668_ = ~new_n83_ & ~new_n84_;
  assign new_n669_ = new_n667_ & new_n668_;
  assign new_n670_ = new_n666_ & new_n669_;
  assign new_n671_ = ~new_n60_ & ~new_n63_;
  assign new_n672_ = ~new_n73_ & new_n671_;
  assign new_n673_ = ~new_n47_ & ~new_n50_;
  assign new_n674_ = ~new_n34_ & ~new_n37_;
  assign new_n675_ = new_n673_ & new_n674_;
  assign new_n676_ = new_n672_ & new_n675_;
  assign new_n677_ = new_n670_ & new_n676_;
  assign new_n678_ = new_n664_ & new_n677_;
  assign new_n679_ = new_n651_ & new_n678_;
  assign pd0 = ~new_n624_ | ~new_n679_;
  assign new_n681_ = pe & pf;
  assign new_n682_ = ~pa0 & pf;
  assign new_n683_ = ~pa & ~new_n682_;
  assign new_n684_ = ~pc & ~new_n681_;
  assign pe0 = ~new_n683_ | ~new_n684_;
  assign new_n686_ = ~pb0 & ~pe;
  assign new_n687_ = pc & ~pe;
  assign new_n688_ = pa & ~pe;
  assign new_n689_ = ~new_n686_ & ~new_n687_;
  assign pf0 = new_n688_ | ~new_n689_;
endmodule

