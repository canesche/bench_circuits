module term1 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x,
    y, z, a0, c0, d0, e0, f0, g0, h0, i0,
    j0, k0, l0, m0, n0, o0, p0, q0, r0, s0  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, x, y, z, a0, c0, d0, e0, f0, g0, h0, i0;
  output j0, k0, l0, m0, n0, o0, p0, q0, r0, s0;
  wire new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_,
    new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_,
    new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_,
    new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n118_, new_n119_, new_n120_, new_n121_,
    new_n122_, new_n123_, new_n124_, new_n125_, new_n126_, new_n127_,
    new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_,
    new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_,
    new_n140_, new_n141_, new_n142_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n165_,
    new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_;
  assign new_n45_ = c & ~i0;
  assign new_n46_ = ~c & i0;
  assign new_n47_ = ~d & ~new_n46_;
  assign new_n48_ = ~new_n45_ & ~new_n47_;
  assign new_n49_ = ~c & d;
  assign new_n50_ = ~h0 & new_n49_;
  assign new_n51_ = new_n48_ & ~new_n50_;
  assign new_n52_ = c & ~d;
  assign new_n53_ = h0 & new_n52_;
  assign k0 = ~new_n51_ & ~new_n53_;
  assign new_n55_ = i & ~j;
  assign new_n56_ = ~e & ~h;
  assign new_n57_ = e & h;
  assign new_n58_ = ~new_n56_ & ~new_n57_;
  assign new_n59_ = ~d & f;
  assign new_n60_ = e & ~new_n59_;
  assign new_n61_ = ~h & new_n60_;
  assign new_n62_ = ~d & ~new_n58_;
  assign new_n63_ = f & new_n62_;
  assign new_n64_ = ~e & ~new_n59_;
  assign new_n65_ = h & new_n64_;
  assign new_n66_ = ~new_n63_ & ~new_n65_;
  assign new_n67_ = ~new_n61_ & new_n66_;
  assign new_n68_ = ~c & g;
  assign new_n69_ = ~new_n58_ & ~new_n68_;
  assign new_n70_ = ~new_n56_ & ~new_n59_;
  assign new_n71_ = ~new_n68_ & new_n70_;
  assign new_n72_ = ~new_n57_ & new_n71_;
  assign new_n73_ = ~c & new_n67_;
  assign new_n74_ = g & new_n73_;
  assign new_n75_ = ~d & new_n69_;
  assign new_n76_ = f & new_n75_;
  assign new_n77_ = ~new_n74_ & ~new_n76_;
  assign new_n78_ = ~new_n72_ & new_n77_;
  assign new_n79_ = ~d & ~new_n56_;
  assign new_n80_ = ~new_n57_ & ~new_n79_;
  assign new_n81_ = d & ~e;
  assign new_n82_ = ~h & new_n81_;
  assign new_n83_ = new_n80_ & ~new_n82_;
  assign new_n84_ = ~d & e;
  assign new_n85_ = h & new_n84_;
  assign new_n86_ = ~new_n83_ & ~new_n85_;
  assign new_n87_ = d & ~new_n56_;
  assign new_n88_ = ~new_n57_ & ~new_n87_;
  assign new_n89_ = ~d & ~e;
  assign new_n90_ = ~h & new_n89_;
  assign new_n91_ = new_n88_ & ~new_n90_;
  assign new_n92_ = d & e;
  assign new_n93_ = h & new_n92_;
  assign new_n94_ = ~new_n91_ & ~new_n93_;
  assign new_n95_ = c & new_n94_;
  assign new_n96_ = ~new_n86_ & ~new_n95_;
  assign new_n97_ = c & ~new_n94_;
  assign new_n98_ = ~new_n96_ & ~new_n97_;
  assign new_n99_ = ~b & ~new_n78_;
  assign new_n100_ = b & ~new_n98_;
  assign new_n101_ = ~new_n99_ & ~new_n100_;
  assign l0 = new_n55_ & ~new_n101_;
  assign new_n103_ = ~a0 & ~c0;
  assign new_n104_ = z & new_n103_;
  assign new_n105_ = ~p & ~u;
  assign new_n106_ = ~q & ~v;
  assign new_n107_ = ~new_n105_ & ~new_n106_;
  assign new_n108_ = ~r & ~w;
  assign new_n109_ = new_n107_ & ~new_n108_;
  assign new_n110_ = ~s & ~x;
  assign new_n111_ = ~t & ~y;
  assign new_n112_ = ~new_n110_ & ~new_n111_;
  assign new_n113_ = new_n109_ & new_n112_;
  assign new_n114_ = c & d;
  assign new_n115_ = ~new_n113_ & ~new_n114_;
  assign new_n116_ = b & new_n104_;
  assign m0 = new_n115_ & new_n116_;
  assign new_n118_ = z & ~a0;
  assign new_n119_ = ~new_n105_ & ~new_n110_;
  assign new_n120_ = ~new_n108_ & new_n119_;
  assign new_n121_ = ~new_n106_ & ~new_n111_;
  assign new_n122_ = new_n120_ & new_n121_;
  assign new_n123_ = ~new_n106_ & ~new_n110_;
  assign new_n124_ = ~new_n108_ & new_n123_;
  assign new_n125_ = ~new_n105_ & ~new_n111_;
  assign new_n126_ = new_n124_ & new_n125_;
  assign new_n127_ = ~c & ~new_n122_;
  assign new_n128_ = ~d & ~new_n126_;
  assign new_n129_ = ~new_n127_ & ~new_n128_;
  assign new_n130_ = ~new_n110_ & new_n125_;
  assign new_n131_ = ~new_n106_ & ~new_n108_;
  assign new_n132_ = new_n130_ & new_n131_;
  assign new_n133_ = ~new_n114_ & ~new_n132_;
  assign new_n134_ = ~d0 & new_n133_;
  assign new_n135_ = ~c0 & ~new_n129_;
  assign new_n136_ = ~new_n134_ & ~new_n135_;
  assign new_n137_ = d0 & ~new_n129_;
  assign new_n138_ = ~c0 & ~new_n137_;
  assign new_n139_ = ~d0 & ~new_n133_;
  assign new_n140_ = ~new_n138_ & ~new_n139_;
  assign new_n141_ = ~new_n136_ & new_n140_;
  assign new_n142_ = b & new_n118_;
  assign n0 = new_n141_ & new_n142_;
  assign new_n144_ = d0 & ~e0;
  assign new_n145_ = new_n107_ & ~new_n110_;
  assign new_n146_ = ~new_n108_ & ~new_n111_;
  assign new_n147_ = new_n145_ & new_n146_;
  assign new_n148_ = ~c0 & ~new_n147_;
  assign new_n149_ = ~d0 & ~new_n122_;
  assign new_n150_ = ~new_n148_ & ~new_n149_;
  assign new_n151_ = ~new_n108_ & ~new_n110_;
  assign new_n152_ = ~new_n106_ & new_n151_;
  assign new_n153_ = new_n125_ & new_n152_;
  assign new_n154_ = ~d0 & ~new_n153_;
  assign new_n155_ = ~new_n148_ & ~new_n154_;
  assign new_n156_ = ~d & e0;
  assign new_n157_ = ~new_n155_ & new_n156_;
  assign new_n158_ = ~c & ~new_n150_;
  assign new_n159_ = e0 & new_n158_;
  assign new_n160_ = new_n133_ & new_n144_;
  assign new_n161_ = c0 & new_n160_;
  assign new_n162_ = ~new_n159_ & ~new_n161_;
  assign new_n163_ = ~new_n157_ & new_n162_;
  assign o0 = new_n142_ & ~new_n163_;
  assign new_n165_ = e0 & ~f0;
  assign new_n166_ = d0 & new_n165_;
  assign new_n167_ = d0 & e0;
  assign new_n168_ = c0 & new_n167_;
  assign new_n169_ = x & ~new_n111_;
  assign new_n170_ = w & new_n169_;
  assign new_n171_ = ~new_n168_ & ~new_n170_;
  assign new_n172_ = r & new_n112_;
  assign new_n173_ = s & ~new_n111_;
  assign new_n174_ = w & new_n173_;
  assign new_n175_ = ~new_n172_ & ~new_n174_;
  assign new_n176_ = new_n171_ & new_n175_;
  assign new_n177_ = ~new_n107_ & ~new_n168_;
  assign new_n178_ = ~new_n176_ & ~new_n177_;
  assign new_n179_ = ~d & f0;
  assign new_n180_ = ~new_n178_ & new_n179_;
  assign new_n181_ = ~c & ~new_n178_;
  assign new_n182_ = f0 & new_n181_;
  assign new_n183_ = new_n133_ & new_n166_;
  assign new_n184_ = c0 & new_n183_;
  assign new_n185_ = ~new_n182_ & ~new_n184_;
  assign new_n186_ = ~new_n180_ & new_n185_;
  assign p0 = new_n142_ & ~new_n186_;
  assign new_n188_ = ~new_n108_ & new_n112_;
  assign new_n189_ = w & ~new_n110_;
  assign new_n190_ = v & new_n189_;
  assign new_n191_ = ~new_n111_ & new_n190_;
  assign new_n192_ = v & new_n172_;
  assign new_n193_ = q & new_n188_;
  assign new_n194_ = ~new_n192_ & ~new_n193_;
  assign new_n195_ = ~new_n191_ & new_n194_;
  assign new_n196_ = e0 & f0;
  assign new_n197_ = c0 & d0;
  assign new_n198_ = new_n196_ & new_n197_;
  assign new_n199_ = f0 & ~g0;
  assign new_n200_ = new_n168_ & new_n199_;
  assign new_n201_ = ~new_n114_ & ~new_n200_;
  assign new_n202_ = ~a0 & new_n201_;
  assign new_n203_ = b & z;
  assign new_n204_ = new_n202_ & new_n203_;
  assign new_n205_ = u & new_n188_;
  assign new_n206_ = v & new_n205_;
  assign new_n207_ = g0 & ~new_n198_;
  assign new_n208_ = ~new_n206_ & ~new_n207_;
  assign new_n209_ = new_n204_ & new_n208_;
  assign new_n210_ = p & ~new_n195_;
  assign new_n211_ = u & new_n193_;
  assign new_n212_ = ~new_n210_ & ~new_n211_;
  assign q0 = ~new_n209_ | ~new_n212_;
  assign new_n214_ = s & t;
  assign new_n215_ = r & new_n214_;
  assign new_n216_ = ~p & q;
  assign new_n217_ = k & new_n216_;
  assign new_n218_ = ~c0 & ~d0;
  assign new_n219_ = e0 & ~new_n218_;
  assign new_n220_ = ~f0 & ~new_n219_;
  assign new_n221_ = f0 & new_n219_;
  assign new_n222_ = ~new_n220_ & ~new_n221_;
  assign new_n223_ = p & ~q;
  assign new_n224_ = l & new_n223_;
  assign new_n225_ = p & q;
  assign new_n226_ = m & new_n225_;
  assign new_n227_ = ~r & new_n214_;
  assign new_n228_ = n & new_n225_;
  assign new_n229_ = ~s & t;
  assign new_n230_ = r & new_n229_;
  assign new_n231_ = r & s;
  assign new_n232_ = q & new_n231_;
  assign new_n233_ = o & p;
  assign new_n234_ = new_n232_ & new_n233_;
  assign new_n235_ = ~f0 & new_n218_;
  assign new_n236_ = ~t & ~new_n235_;
  assign new_n237_ = new_n234_ & new_n236_;
  assign new_n238_ = f0 & ~new_n219_;
  assign new_n239_ = f0 & ~new_n218_;
  assign new_n240_ = e0 & ~new_n239_;
  assign new_n241_ = ~new_n238_ & ~new_n240_;
  assign new_n242_ = new_n237_ & ~new_n241_;
  assign new_n243_ = new_n226_ & new_n227_;
  assign new_n244_ = new_n228_ & new_n230_;
  assign new_n245_ = ~new_n243_ & ~new_n244_;
  assign new_n246_ = new_n222_ & ~new_n245_;
  assign new_n247_ = ~new_n242_ & ~new_n246_;
  assign new_n248_ = ~new_n217_ & ~new_n224_;
  assign new_n249_ = new_n222_ & ~new_n248_;
  assign new_n250_ = new_n215_ & new_n249_;
  assign new_n251_ = new_n247_ & ~new_n250_;
  assign new_n252_ = ~l & r;
  assign new_n253_ = new_n214_ & new_n252_;
  assign new_n254_ = ~m & new_n214_;
  assign new_n255_ = ~o & s;
  assign new_n256_ = n & ~s;
  assign new_n257_ = t & ~new_n256_;
  assign new_n258_ = ~new_n255_ & ~new_n257_;
  assign new_n259_ = ~q & ~new_n253_;
  assign new_n260_ = ~r & ~new_n254_;
  assign new_n261_ = ~new_n259_ & ~new_n260_;
  assign new_n262_ = ~new_n258_ & new_n261_;
  assign new_n263_ = q & r;
  assign new_n264_ = new_n214_ & new_n263_;
  assign new_n265_ = ~k & new_n263_;
  assign new_n266_ = new_n214_ & new_n265_;
  assign new_n267_ = ~r & ~t;
  assign new_n268_ = g0 & ~new_n267_;
  assign new_n269_ = ~new_n266_ & new_n268_;
  assign new_n270_ = r & t;
  assign new_n271_ = ~s & ~new_n270_;
  assign new_n272_ = new_n269_ & ~new_n271_;
  assign new_n273_ = ~new_n220_ & new_n272_;
  assign new_n274_ = ~q & ~new_n215_;
  assign new_n275_ = ~new_n221_ & ~new_n274_;
  assign new_n276_ = new_n273_ & new_n275_;
  assign new_n277_ = ~p & ~new_n264_;
  assign new_n278_ = p & new_n262_;
  assign new_n279_ = ~new_n277_ & ~new_n278_;
  assign new_n280_ = new_n276_ & new_n279_;
  assign new_n281_ = g0 & ~new_n251_;
  assign new_n282_ = h0 & ~new_n280_;
  assign new_n283_ = ~new_n281_ & ~new_n282_;
  assign new_n284_ = h0 & new_n280_;
  assign new_n285_ = ~new_n283_ & ~new_n284_;
  assign new_n286_ = a & ~a0;
  assign r0 = new_n285_ & new_n286_;
  assign new_n288_ = t & ~i0;
  assign new_n289_ = k & ~p;
  assign new_n290_ = new_n288_ & new_n289_;
  assign new_n291_ = f0 & g0;
  assign new_n292_ = ~g0 & new_n220_;
  assign new_n293_ = ~new_n218_ & new_n291_;
  assign new_n294_ = e0 & new_n293_;
  assign new_n295_ = ~new_n292_ & ~new_n294_;
  assign new_n296_ = ~new_n258_ & ~new_n260_;
  assign new_n297_ = ~l & new_n231_;
  assign new_n298_ = t & new_n297_;
  assign new_n299_ = ~r & ~new_n214_;
  assign new_n300_ = ~new_n298_ & ~new_n299_;
  assign new_n301_ = ~s & ~t;
  assign new_n302_ = ~new_n218_ & ~new_n301_;
  assign new_n303_ = new_n300_ & new_n302_;
  assign new_n304_ = q & new_n296_;
  assign new_n305_ = ~new_n274_ & ~new_n304_;
  assign new_n306_ = new_n303_ & new_n305_;
  assign new_n307_ = ~f0 & ~g0;
  assign new_n308_ = o & ~t;
  assign new_n309_ = ~n & t;
  assign new_n310_ = ~s & ~new_n309_;
  assign new_n311_ = ~new_n308_ & ~new_n310_;
  assign new_n312_ = r & ~new_n214_;
  assign new_n313_ = ~m & ~new_n312_;
  assign new_n314_ = ~new_n299_ & ~new_n313_;
  assign new_n315_ = c0 & e0;
  assign new_n316_ = ~new_n301_ & ~new_n315_;
  assign new_n317_ = new_n314_ & new_n316_;
  assign new_n318_ = r & new_n311_;
  assign new_n319_ = ~new_n167_ & ~new_n318_;
  assign new_n320_ = new_n317_ & new_n319_;
  assign new_n321_ = l & ~q;
  assign new_n322_ = new_n215_ & new_n321_;
  assign new_n323_ = ~new_n219_ & new_n322_;
  assign new_n324_ = new_n307_ & new_n323_;
  assign new_n325_ = new_n291_ & new_n306_;
  assign new_n326_ = e0 & new_n325_;
  assign new_n327_ = new_n307_ & new_n320_;
  assign new_n328_ = q & new_n327_;
  assign new_n329_ = ~new_n326_ & ~new_n328_;
  assign new_n330_ = ~new_n324_ & new_n329_;
  assign new_n331_ = new_n261_ & new_n311_;
  assign new_n332_ = e0 & new_n239_;
  assign new_n333_ = ~new_n307_ & ~new_n332_;
  assign new_n334_ = ~r & ~s;
  assign new_n335_ = ~k & new_n215_;
  assign new_n336_ = q & new_n335_;
  assign new_n337_ = ~new_n334_ & ~new_n336_;
  assign new_n338_ = ~new_n333_ & new_n337_;
  assign new_n339_ = ~t & ~new_n231_;
  assign new_n340_ = new_n338_ & ~new_n339_;
  assign new_n341_ = ~g0 & new_n219_;
  assign new_n342_ = ~new_n274_ & ~new_n341_;
  assign new_n343_ = new_n340_ & new_n342_;
  assign new_n344_ = ~p & new_n264_;
  assign new_n345_ = ~new_n277_ & ~new_n331_;
  assign new_n346_ = ~new_n344_ & ~new_n345_;
  assign new_n347_ = new_n343_ & ~new_n346_;
  assign new_n348_ = i0 & ~new_n347_;
  assign new_n349_ = new_n232_ & ~new_n295_;
  assign new_n350_ = new_n290_ & new_n349_;
  assign new_n351_ = p & ~new_n330_;
  assign new_n352_ = ~i0 & new_n351_;
  assign new_n353_ = ~new_n350_ & ~new_n352_;
  assign new_n354_ = ~new_n348_ & new_n353_;
  assign s0 = new_n286_ & ~new_n354_;
  assign j0 = ~h0;
endmodule

