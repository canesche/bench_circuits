module top ( 
    pv28_20_, pv56_12_, pv56_23_, pv88_6_, pv88_19_, pv120_16_, pv120_29_,
    pv28_10_, pv56_13_, pv56_22_, pv88_7_, pv88_29_, pv120_15_, pv56_14_,
    pv56_25_, pv88_8_, pv88_17_, pv88_28_, pv120_18_, pv56_15_, pv56_24_,
    pv88_9_, pv88_18_, pv88_27_, pv120_17_, pv88_2_, pv88_15_, pv88_26_,
    pv120_12_, pv88_3_, pv88_16_, pv88_25_, pv120_11_, pv56_10_, pv56_21_,
    pv88_4_, pv88_13_, pv88_24_, pv120_14_, pv126_5_, pv56_11_, pv56_20_,
    pv88_5_, pv88_14_, pv88_23_, pv120_13_, pv28_8_, pv56_5_, pv88_11_,
    pv88_22_, pv120_5_, pv132_0_, pv28_9_, pv56_4_, pv88_12_, pv88_21_,
    pv120_6_, pv28_6_, pv56_7_, pv88_20_, pv120_3_, pv120_10_, pv28_7_,
    pv56_6_, pv88_10_, pv120_4_, pv28_4_, pv56_9_, pv120_1_, pv28_5_,
    pv56_8_, pv120_2_, pv28_2_, pv28_3_, pv120_0_, pv28_0_, pv28_1_,
    pv132_5_, pv56_1_, pv120_9_, pv120_30_, pv132_4_, pv56_0_, pv88_30_,
    pv132_3_, pv28_19_, pv56_3_, pv88_31_, pv120_7_, pv132_2_, pv56_2_,
    pv120_8_, pv120_20_, pv132_1_, pv28_17_, pv120_21_, pv126_3_, pv28_18_,
    pv28_27_, pv120_22_, pv126_4_, pv28_15_, pv28_26_, pv88_0_, pv120_23_,
    pv126_1_, pv28_16_, pv28_25_, pv88_1_, pv120_24_, pv120_31_, pv126_2_,
    pv28_13_, pv28_24_, pv56_16_, pv56_27_, pv120_25_, pv28_14_, pv28_23_,
    pv56_17_, pv56_26_, pv120_19_, pv120_26_, pv126_0_, pv28_11_, pv28_22_,
    pv56_18_, pv120_27_, pv28_12_, pv28_21_, pv56_19_, pv120_28_,
    pv138_3_, pv138_2_, pv138_1_, pv138_0_, pv134_1_, pv134_0_  );
  input  pv28_20_, pv56_12_, pv56_23_, pv88_6_, pv88_19_, pv120_16_,
    pv120_29_, pv28_10_, pv56_13_, pv56_22_, pv88_7_, pv88_29_, pv120_15_,
    pv56_14_, pv56_25_, pv88_8_, pv88_17_, pv88_28_, pv120_18_, pv56_15_,
    pv56_24_, pv88_9_, pv88_18_, pv88_27_, pv120_17_, pv88_2_, pv88_15_,
    pv88_26_, pv120_12_, pv88_3_, pv88_16_, pv88_25_, pv120_11_, pv56_10_,
    pv56_21_, pv88_4_, pv88_13_, pv88_24_, pv120_14_, pv126_5_, pv56_11_,
    pv56_20_, pv88_5_, pv88_14_, pv88_23_, pv120_13_, pv28_8_, pv56_5_,
    pv88_11_, pv88_22_, pv120_5_, pv132_0_, pv28_9_, pv56_4_, pv88_12_,
    pv88_21_, pv120_6_, pv28_6_, pv56_7_, pv88_20_, pv120_3_, pv120_10_,
    pv28_7_, pv56_6_, pv88_10_, pv120_4_, pv28_4_, pv56_9_, pv120_1_,
    pv28_5_, pv56_8_, pv120_2_, pv28_2_, pv28_3_, pv120_0_, pv28_0_,
    pv28_1_, pv132_5_, pv56_1_, pv120_9_, pv120_30_, pv132_4_, pv56_0_,
    pv88_30_, pv132_3_, pv28_19_, pv56_3_, pv88_31_, pv120_7_, pv132_2_,
    pv56_2_, pv120_8_, pv120_20_, pv132_1_, pv28_17_, pv120_21_, pv126_3_,
    pv28_18_, pv28_27_, pv120_22_, pv126_4_, pv28_15_, pv28_26_, pv88_0_,
    pv120_23_, pv126_1_, pv28_16_, pv28_25_, pv88_1_, pv120_24_, pv120_31_,
    pv126_2_, pv28_13_, pv28_24_, pv56_16_, pv56_27_, pv120_25_, pv28_14_,
    pv28_23_, pv56_17_, pv56_26_, pv120_19_, pv120_26_, pv126_0_, pv28_11_,
    pv28_22_, pv56_18_, pv120_27_, pv28_12_, pv28_21_, pv56_19_, pv120_28_;
  output pv138_3_, pv138_2_, pv138_1_, pv138_0_, pv134_1_, pv134_0_;
  wire new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_;
  assign new_n139_ = ~pv132_3_ & ~pv126_3_;
  assign new_n140_ = ~pv88_25_ & ~pv120_25_;
  assign new_n141_ = ~pv132_4_ & ~pv126_4_;
  assign new_n142_ = ~pv132_2_ & ~pv126_2_;
  assign new_n143_ = ~pv126_5_ & ~pv132_5_;
  assign new_n144_ = ~pv88_31_ & ~pv120_31_;
  assign new_n145_ = ~pv120_30_ & ~pv88_30_;
  assign new_n146_ = ~pv132_0_ & ~pv126_0_;
  assign new_n147_ = ~pv132_1_ & ~pv126_1_;
  assign new_n148_ = ~pv88_27_ & ~pv120_27_;
  assign new_n149_ = ~pv120_29_ & ~pv88_29_;
  assign new_n150_ = ~pv88_26_ & ~pv120_26_;
  assign new_n151_ = ~pv88_23_ & ~pv120_23_;
  assign new_n152_ = ~pv88_28_ & ~pv120_28_;
  assign new_n153_ = ~pv88_24_ & ~pv120_24_;
  assign new_n154_ = ~pv88_22_ & ~pv120_22_;
  assign new_n155_ = ~new_n139_ & ~new_n140_;
  assign new_n156_ = ~new_n141_ & new_n155_;
  assign new_n157_ = ~new_n142_ & new_n156_;
  assign new_n158_ = ~new_n143_ & new_n157_;
  assign new_n159_ = ~new_n144_ & new_n158_;
  assign new_n160_ = ~new_n145_ & new_n159_;
  assign new_n161_ = ~new_n146_ & new_n160_;
  assign new_n162_ = ~new_n147_ & new_n161_;
  assign new_n163_ = ~new_n148_ & new_n162_;
  assign new_n164_ = ~new_n149_ & new_n163_;
  assign new_n165_ = ~new_n150_ & new_n164_;
  assign new_n166_ = ~new_n151_ & new_n165_;
  assign new_n167_ = ~new_n152_ & new_n166_;
  assign new_n168_ = ~new_n153_ & new_n167_;
  assign pv138_3_ = ~new_n154_ & new_n168_;
  assign new_n170_ = ~pv88_19_ & ~pv120_19_;
  assign new_n171_ = ~pv88_9_ & ~pv120_9_;
  assign new_n172_ = ~pv88_20_ & ~pv120_20_;
  assign new_n173_ = ~pv120_18_ & ~pv88_18_;
  assign new_n174_ = ~pv88_21_ & ~pv120_21_;
  assign new_n175_ = ~pv120_15_ & ~pv88_15_;
  assign new_n176_ = ~pv120_14_ & ~pv88_14_;
  assign new_n177_ = ~pv120_16_ & ~pv88_16_;
  assign new_n178_ = ~pv88_17_ & ~pv120_17_;
  assign new_n179_ = ~pv120_11_ & ~pv88_11_;
  assign new_n180_ = ~pv88_13_ & ~pv120_13_;
  assign new_n181_ = ~pv120_10_ & ~pv88_10_;
  assign new_n182_ = ~pv88_7_ & ~pv120_7_;
  assign new_n183_ = ~pv120_12_ & ~pv88_12_;
  assign new_n184_ = ~pv88_8_ & ~pv120_8_;
  assign new_n185_ = ~pv88_6_ & ~pv120_6_;
  assign new_n186_ = ~new_n170_ & ~new_n171_;
  assign new_n187_ = ~new_n172_ & new_n186_;
  assign new_n188_ = ~new_n173_ & new_n187_;
  assign new_n189_ = ~new_n174_ & new_n188_;
  assign new_n190_ = ~new_n175_ & new_n189_;
  assign new_n191_ = ~new_n176_ & new_n190_;
  assign new_n192_ = ~new_n177_ & new_n191_;
  assign new_n193_ = ~new_n178_ & new_n192_;
  assign new_n194_ = ~new_n179_ & new_n193_;
  assign new_n195_ = ~new_n180_ & new_n194_;
  assign new_n196_ = ~new_n181_ & new_n195_;
  assign new_n197_ = ~new_n182_ & new_n196_;
  assign new_n198_ = ~new_n183_ & new_n197_;
  assign new_n199_ = ~new_n184_ & new_n198_;
  assign pv138_2_ = ~new_n185_ & new_n199_;
  assign new_n201_ = ~pv88_3_ & ~pv120_3_;
  assign new_n202_ = ~pv56_21_ & ~pv28_21_;
  assign new_n203_ = ~pv88_4_ & ~pv120_4_;
  assign new_n204_ = ~pv88_2_ & ~pv120_2_;
  assign new_n205_ = ~pv88_5_ & ~pv120_5_;
  assign new_n206_ = ~pv28_27_ & ~pv56_27_;
  assign new_n207_ = ~pv28_26_ & ~pv56_26_;
  assign new_n208_ = ~pv120_0_ & ~pv88_0_;
  assign new_n209_ = ~pv120_1_ & ~pv88_1_;
  assign new_n210_ = ~pv56_23_ & ~pv28_23_;
  assign new_n211_ = ~pv56_25_ & ~pv28_25_;
  assign new_n212_ = ~pv56_22_ & ~pv28_22_;
  assign new_n213_ = ~pv28_19_ & ~pv56_19_;
  assign new_n214_ = ~pv56_24_ & ~pv28_24_;
  assign new_n215_ = ~pv28_20_ & ~pv56_20_;
  assign new_n216_ = ~pv28_18_ & ~pv56_18_;
  assign new_n217_ = ~new_n201_ & ~new_n202_;
  assign new_n218_ = ~new_n203_ & new_n217_;
  assign new_n219_ = ~new_n204_ & new_n218_;
  assign new_n220_ = ~new_n205_ & new_n219_;
  assign new_n221_ = ~new_n206_ & new_n220_;
  assign new_n222_ = ~new_n207_ & new_n221_;
  assign new_n223_ = ~new_n208_ & new_n222_;
  assign new_n224_ = ~new_n209_ & new_n223_;
  assign new_n225_ = ~new_n210_ & new_n224_;
  assign new_n226_ = ~new_n211_ & new_n225_;
  assign new_n227_ = ~new_n212_ & new_n226_;
  assign new_n228_ = ~new_n213_ & new_n227_;
  assign new_n229_ = ~new_n214_ & new_n228_;
  assign new_n230_ = ~new_n215_ & new_n229_;
  assign pv138_1_ = ~new_n216_ & new_n230_;
  assign new_n232_ = ~pv56_15_ & ~pv28_15_;
  assign new_n233_ = ~pv56_5_ & ~pv28_5_;
  assign new_n234_ = ~pv28_16_ & ~pv56_16_;
  assign new_n235_ = ~pv56_14_ & ~pv28_14_;
  assign new_n236_ = ~pv28_17_ & ~pv56_17_;
  assign new_n237_ = ~pv56_11_ & ~pv28_11_;
  assign new_n238_ = ~pv28_10_ & ~pv56_10_;
  assign new_n239_ = ~pv56_12_ & ~pv28_12_;
  assign new_n240_ = ~pv56_13_ & ~pv28_13_;
  assign new_n241_ = ~pv56_7_ & ~pv28_7_;
  assign new_n242_ = ~pv28_9_ & ~pv56_9_;
  assign new_n243_ = ~pv28_6_ & ~pv56_6_;
  assign new_n244_ = ~pv28_3_ & ~pv56_3_;
  assign new_n245_ = ~pv28_8_ & ~pv56_8_;
  assign new_n246_ = ~pv56_4_ & ~pv28_4_;
  assign new_n247_ = ~pv28_2_ & ~pv56_2_;
  assign new_n248_ = ~new_n232_ & ~new_n233_;
  assign new_n249_ = ~new_n234_ & new_n248_;
  assign new_n250_ = ~new_n235_ & new_n249_;
  assign new_n251_ = ~new_n236_ & new_n250_;
  assign new_n252_ = ~new_n237_ & new_n251_;
  assign new_n253_ = ~new_n238_ & new_n252_;
  assign new_n254_ = ~new_n239_ & new_n253_;
  assign new_n255_ = ~new_n240_ & new_n254_;
  assign new_n256_ = ~new_n241_ & new_n255_;
  assign new_n257_ = ~new_n242_ & new_n256_;
  assign new_n258_ = ~new_n243_ & new_n257_;
  assign new_n259_ = ~new_n244_ & new_n258_;
  assign new_n260_ = ~new_n245_ & new_n259_;
  assign new_n261_ = ~new_n246_ & new_n260_;
  assign pv138_0_ = ~new_n247_ & new_n261_;
  assign pv134_1_ = pv28_1_ | pv56_1_;
  assign pv134_0_ = pv28_0_ | pv56_0_;
endmodule

