module top ( 
    pp, pq, pr, ps, pt, pu, pv, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk,
    pl, pm, po,
    pa0, pb0, pc0, pd0, pe0, pf0, pg0, pw, ph0, px, pi0, py, pj0, pz, pk0,
    pl0, pm0, pn0, po0, pp0  );
  input  pp, pq, pr, ps, pt, pu, pv, pa, pb, pc, pd, pe, pf, pg, ph, pi,
    pj, pk, pl, pm, po;
  output pa0, pb0, pc0, pd0, pe0, pf0, pg0, pw, ph0, px, pi0, py, pj0, pz,
    pk0, pl0, pm0, pn0, po0, pp0;
  wire new_n44_, new_n45_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n56_, new_n57_, new_n58_, new_n60_,
    new_n61_, new_n62_, new_n63_, new_n64_, new_n66_, new_n67_, new_n68_,
    new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_,
    new_n77_, new_n78_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_,
    new_n86_, new_n87_, new_n88_, new_n89_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n96_, new_n97_, new_n98_, new_n99_, new_n101_, new_n102_,
    new_n103_, new_n104_;
  assign pf0 = pi & pj;
  assign pw = pv & pl;
  assign new_n44_ = ~pp & pi;
  assign new_n45_ = pk & new_n44_;
  assign px = pq & new_n45_;
  assign new_n47_ = ~pq & pi;
  assign new_n48_ = pk & new_n47_;
  assign new_n49_ = ~pa & new_n48_;
  assign new_n50_ = pm & ~new_n49_;
  assign new_n51_ = pi & pk;
  assign new_n52_ = ~pq & new_n51_;
  assign new_n53_ = new_n50_ & new_n52_;
  assign new_n54_ = po & new_n50_;
  assign pi0 = new_n53_ | new_n54_;
  assign new_n56_ = ~pl & pm;
  assign new_n57_ = new_n52_ & new_n56_;
  assign new_n58_ = pp & new_n56_;
  assign py = new_n57_ | new_n58_;
  assign new_n60_ = pb & new_n48_;
  assign new_n61_ = pm & ~new_n60_;
  assign new_n62_ = pq & new_n51_;
  assign new_n63_ = new_n61_ & new_n62_;
  assign new_n64_ = pp & new_n61_;
  assign pj0 = new_n63_ | new_n64_;
  assign new_n66_ = pi & pm;
  assign new_n67_ = ~pp & pk;
  assign new_n68_ = new_n66_ & new_n67_;
  assign pz = pq & new_n68_;
  assign new_n70_ = ~pq & ~pi;
  assign new_n71_ = ~pq & ~pk;
  assign new_n72_ = ~new_n70_ & ~new_n71_;
  assign new_n73_ = pm & new_n72_;
  assign new_n74_ = ~pi & new_n73_;
  assign new_n75_ = ~pq & pc;
  assign new_n76_ = new_n73_ & new_n75_;
  assign new_n77_ = ~pk & new_n73_;
  assign new_n78_ = ~new_n74_ & ~new_n76_;
  assign pk0 = new_n77_ | ~new_n78_;
  assign new_n80_ = ~pd & new_n48_;
  assign new_n81_ = pm & ~new_n80_;
  assign new_n82_ = pr & new_n81_;
  assign new_n83_ = ~pp & new_n82_;
  assign new_n84_ = new_n52_ & new_n81_;
  assign pl0 = new_n83_ | new_n84_;
  assign new_n86_ = ~pe & new_n48_;
  assign new_n87_ = pm & ~new_n86_;
  assign new_n88_ = new_n52_ & new_n87_;
  assign new_n89_ = ps & new_n87_;
  assign pm0 = new_n88_ | new_n89_;
  assign new_n91_ = ~pf & new_n48_;
  assign new_n92_ = pm & ~new_n91_;
  assign new_n93_ = new_n52_ & new_n92_;
  assign new_n94_ = pt & new_n92_;
  assign pn0 = new_n93_ | new_n94_;
  assign new_n96_ = ~pg & new_n48_;
  assign new_n97_ = pm & ~new_n96_;
  assign new_n98_ = new_n52_ & new_n97_;
  assign new_n99_ = pu & new_n97_;
  assign po0 = new_n98_ | new_n99_;
  assign new_n101_ = ~ph & new_n48_;
  assign new_n102_ = pm & ~new_n101_;
  assign new_n103_ = new_n52_ & new_n102_;
  assign new_n104_ = pv & new_n102_;
  assign pp0 = new_n103_ | new_n104_;
  assign pa0 = ~pt;
  assign pg0 = ~pf0;
  assign pb0 = pu;
  assign pc0 = pq;
  assign pd0 = ps;
  assign pe0 = pr;
  assign ph0 = pp;
endmodule

