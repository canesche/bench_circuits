module MultiplierA_16 ( clock, 
    \1 , 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18,
    36  );
  input  clock;
  input  \1 , 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18;
  output 36;
  reg 2, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34;
  wire new_n67_, new_n68_1_, new_n69_, new_n71_, new_n72_, new_n73_1_,
    new_n74_, new_n75_, new_n76_, new_n77_, new_n78_1_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_1_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_1_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_1_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_1_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_1_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_1_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_1_, new_n114_, new_n115_, new_n116_, new_n117_,
    new_n118_, new_n119_, new_n120_, new_n121_, new_n122_, new_n123_,
    new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_,
    new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_,
    new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_,
    new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_,
    new_n148_, new_n149_, new_n150_, new_n151_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, n38, n43, n48, n53, n58, n63, n68,
    n73, n78, n83, n88, n93, n98, n103, n108, n113;
  assign new_n67_ = \1  & 3;
  assign new_n68_1_ = 20 & ~new_n67_;
  assign new_n69_ = ~20 & new_n67_;
  assign 36 = new_n68_1_ | new_n69_;
  assign new_n71_ = \1  & 18;
  assign new_n72_ = 2 & new_n71_;
  assign new_n73_1_ = 20 & new_n67_;
  assign new_n74_ = \1  & 4;
  assign new_n75_ = ~new_n73_1_ & ~new_n74_;
  assign new_n76_ = 21 & ~new_n75_;
  assign new_n77_ = new_n73_1_ & new_n74_;
  assign new_n78_1_ = ~new_n76_ & ~new_n77_;
  assign new_n79_ = \1  & 5;
  assign new_n80_ = new_n78_1_ & ~new_n79_;
  assign new_n81_ = 22 & ~new_n80_;
  assign new_n82_ = ~new_n78_1_ & new_n79_;
  assign new_n83_1_ = ~new_n81_ & ~new_n82_;
  assign new_n84_ = \1  & 6;
  assign new_n85_ = new_n83_1_ & ~new_n84_;
  assign new_n86_ = 23 & ~new_n85_;
  assign new_n87_ = ~new_n83_1_ & new_n84_;
  assign new_n88_1_ = ~new_n86_ & ~new_n87_;
  assign new_n89_ = \1  & 7;
  assign new_n90_ = new_n88_1_ & ~new_n89_;
  assign new_n91_ = 24 & ~new_n90_;
  assign new_n92_ = ~new_n88_1_ & new_n89_;
  assign new_n93_1_ = ~new_n91_ & ~new_n92_;
  assign new_n94_ = \1  & 8;
  assign new_n95_ = new_n93_1_ & ~new_n94_;
  assign new_n96_ = 25 & ~new_n95_;
  assign new_n97_ = ~new_n93_1_ & new_n94_;
  assign new_n98_1_ = ~new_n96_ & ~new_n97_;
  assign new_n99_ = \1  & 9;
  assign new_n100_ = new_n98_1_ & ~new_n99_;
  assign new_n101_ = 26 & ~new_n100_;
  assign new_n102_ = ~new_n98_1_ & new_n99_;
  assign new_n103_1_ = ~new_n101_ & ~new_n102_;
  assign new_n104_ = \1  & 10;
  assign new_n105_ = new_n103_1_ & ~new_n104_;
  assign new_n106_ = 27 & ~new_n105_;
  assign new_n107_ = ~new_n103_1_ & new_n104_;
  assign new_n108_1_ = ~new_n106_ & ~new_n107_;
  assign new_n109_ = \1  & 11;
  assign new_n110_ = new_n108_1_ & ~new_n109_;
  assign new_n111_ = 28 & ~new_n110_;
  assign new_n112_ = ~new_n108_1_ & new_n109_;
  assign new_n113_1_ = ~new_n111_ & ~new_n112_;
  assign new_n114_ = \1  & 12;
  assign new_n115_ = new_n113_1_ & ~new_n114_;
  assign new_n116_ = 29 & ~new_n115_;
  assign new_n117_ = ~new_n113_1_ & new_n114_;
  assign new_n118_ = ~new_n116_ & ~new_n117_;
  assign new_n119_ = \1  & 13;
  assign new_n120_ = new_n118_ & ~new_n119_;
  assign new_n121_ = 30 & ~new_n120_;
  assign new_n122_ = ~new_n118_ & new_n119_;
  assign new_n123_ = ~new_n121_ & ~new_n122_;
  assign new_n124_ = \1  & 14;
  assign new_n125_ = new_n123_ & ~new_n124_;
  assign new_n126_ = 31 & ~new_n125_;
  assign new_n127_ = ~new_n123_ & new_n124_;
  assign new_n128_ = ~new_n126_ & ~new_n127_;
  assign new_n129_ = \1  & 15;
  assign new_n130_ = new_n128_ & ~new_n129_;
  assign new_n131_ = 32 & ~new_n130_;
  assign new_n132_ = ~new_n128_ & new_n129_;
  assign new_n133_ = ~new_n131_ & ~new_n132_;
  assign new_n134_ = \1  & 16;
  assign new_n135_ = new_n133_ & ~new_n134_;
  assign new_n136_ = 33 & ~new_n135_;
  assign new_n137_ = ~new_n133_ & new_n134_;
  assign new_n138_ = ~new_n136_ & ~new_n137_;
  assign new_n139_ = \1  & 17;
  assign new_n140_ = new_n138_ & ~new_n139_;
  assign new_n141_ = 34 & ~new_n140_;
  assign new_n142_ = ~new_n138_ & new_n139_;
  assign new_n143_ = ~new_n141_ & ~new_n142_;
  assign new_n144_ = new_n72_ & new_n143_;
  assign new_n145_ = 2 & ~new_n71_;
  assign new_n146_ = ~new_n143_ & new_n145_;
  assign new_n147_ = ~new_n144_ & ~new_n146_;
  assign new_n148_ = ~2 & new_n71_;
  assign new_n149_ = ~new_n143_ & new_n148_;
  assign new_n150_ = new_n72_ & ~new_n143_;
  assign new_n151_ = ~new_n149_ & ~new_n150_;
  assign n38 = ~new_n147_ | ~new_n151_;
  assign new_n153_ = ~new_n75_ & ~new_n77_;
  assign new_n154_ = 21 & ~new_n153_;
  assign new_n155_ = ~new_n73_1_ & new_n74_;
  assign new_n156_ = new_n73_1_ & ~new_n74_;
  assign new_n157_ = ~new_n155_ & ~new_n156_;
  assign new_n158_ = ~21 & ~new_n157_;
  assign n43 = new_n154_ | new_n158_;
  assign new_n160_ = ~new_n80_ & ~new_n82_;
  assign new_n161_ = 22 & ~new_n160_;
  assign new_n162_ = new_n78_1_ & new_n79_;
  assign new_n163_ = ~new_n78_1_ & ~new_n79_;
  assign new_n164_ = ~new_n162_ & ~new_n163_;
  assign new_n165_ = ~22 & ~new_n164_;
  assign n48 = new_n161_ | new_n165_;
  assign new_n167_ = ~new_n85_ & ~new_n87_;
  assign new_n168_ = 23 & ~new_n167_;
  assign new_n169_ = new_n83_1_ & new_n84_;
  assign new_n170_ = ~new_n83_1_ & ~new_n84_;
  assign new_n171_ = ~new_n169_ & ~new_n170_;
  assign new_n172_ = ~23 & ~new_n171_;
  assign n53 = new_n168_ | new_n172_;
  assign new_n174_ = ~new_n90_ & ~new_n92_;
  assign new_n175_ = 24 & ~new_n174_;
  assign new_n176_ = new_n88_1_ & new_n89_;
  assign new_n177_ = ~new_n88_1_ & ~new_n89_;
  assign new_n178_ = ~new_n176_ & ~new_n177_;
  assign new_n179_ = ~24 & ~new_n178_;
  assign n58 = new_n175_ | new_n179_;
  assign new_n181_ = ~new_n95_ & ~new_n97_;
  assign new_n182_ = 25 & ~new_n181_;
  assign new_n183_ = new_n93_1_ & new_n94_;
  assign new_n184_ = ~new_n93_1_ & ~new_n94_;
  assign new_n185_ = ~new_n183_ & ~new_n184_;
  assign new_n186_ = ~25 & ~new_n185_;
  assign n63 = new_n182_ | new_n186_;
  assign new_n188_ = ~new_n100_ & ~new_n102_;
  assign new_n189_ = 26 & ~new_n188_;
  assign new_n190_ = new_n98_1_ & new_n99_;
  assign new_n191_ = ~new_n98_1_ & ~new_n99_;
  assign new_n192_ = ~new_n190_ & ~new_n191_;
  assign new_n193_ = ~26 & ~new_n192_;
  assign n68 = new_n189_ | new_n193_;
  assign new_n195_ = ~new_n105_ & ~new_n107_;
  assign new_n196_ = 27 & ~new_n195_;
  assign new_n197_ = new_n103_1_ & new_n104_;
  assign new_n198_ = ~new_n103_1_ & ~new_n104_;
  assign new_n199_ = ~new_n197_ & ~new_n198_;
  assign new_n200_ = ~27 & ~new_n199_;
  assign n73 = new_n196_ | new_n200_;
  assign new_n202_ = ~new_n110_ & ~new_n112_;
  assign new_n203_ = 28 & ~new_n202_;
  assign new_n204_ = new_n108_1_ & new_n109_;
  assign new_n205_ = ~new_n108_1_ & ~new_n109_;
  assign new_n206_ = ~new_n204_ & ~new_n205_;
  assign new_n207_ = ~28 & ~new_n206_;
  assign n78 = new_n203_ | new_n207_;
  assign new_n209_ = ~new_n115_ & ~new_n117_;
  assign new_n210_ = 29 & ~new_n209_;
  assign new_n211_ = new_n113_1_ & new_n114_;
  assign new_n212_ = ~new_n113_1_ & ~new_n114_;
  assign new_n213_ = ~new_n211_ & ~new_n212_;
  assign new_n214_ = ~29 & ~new_n213_;
  assign n83 = new_n210_ | new_n214_;
  assign new_n216_ = ~new_n120_ & ~new_n122_;
  assign new_n217_ = 30 & ~new_n216_;
  assign new_n218_ = new_n118_ & new_n119_;
  assign new_n219_ = ~new_n118_ & ~new_n119_;
  assign new_n220_ = ~new_n218_ & ~new_n219_;
  assign new_n221_ = ~30 & ~new_n220_;
  assign n88 = new_n217_ | new_n221_;
  assign new_n223_ = ~new_n125_ & ~new_n127_;
  assign new_n224_ = 31 & ~new_n223_;
  assign new_n225_ = new_n123_ & new_n124_;
  assign new_n226_ = ~new_n123_ & ~new_n124_;
  assign new_n227_ = ~new_n225_ & ~new_n226_;
  assign new_n228_ = ~31 & ~new_n227_;
  assign n93 = new_n224_ | new_n228_;
  assign new_n230_ = ~new_n130_ & ~new_n132_;
  assign new_n231_ = 32 & ~new_n230_;
  assign new_n232_ = new_n128_ & new_n129_;
  assign new_n233_ = ~new_n128_ & ~new_n129_;
  assign new_n234_ = ~new_n232_ & ~new_n233_;
  assign new_n235_ = ~32 & ~new_n234_;
  assign n98 = new_n231_ | new_n235_;
  assign new_n237_ = ~new_n135_ & ~new_n137_;
  assign new_n238_ = 33 & ~new_n237_;
  assign new_n239_ = new_n133_ & new_n134_;
  assign new_n240_ = ~new_n133_ & ~new_n134_;
  assign new_n241_ = ~new_n239_ & ~new_n240_;
  assign new_n242_ = ~33 & ~new_n241_;
  assign n103 = new_n238_ | new_n242_;
  assign new_n244_ = ~new_n140_ & ~new_n142_;
  assign new_n245_ = 34 & ~new_n244_;
  assign new_n246_ = new_n138_ & new_n139_;
  assign new_n247_ = ~new_n138_ & ~new_n139_;
  assign new_n248_ = ~new_n246_ & ~new_n247_;
  assign new_n249_ = ~34 & ~new_n248_;
  assign n108 = new_n245_ | new_n249_;
  assign new_n251_ = ~new_n71_ & ~new_n143_;
  assign new_n252_ = new_n71_ & new_n143_;
  assign new_n253_ = ~new_n251_ & ~new_n252_;
  assign new_n254_ = 2 & new_n253_;
  assign new_n255_ = ~2 & ~new_n253_;
  assign n113 = new_n254_ | new_n255_;
  always @ (posedge clock) begin
    2 <= n38;
    20 <= n43;
    21 <= n48;
    22 <= n53;
    23 <= n58;
    24 <= n63;
    25 <= n68;
    26 <= n73;
    27 <= n78;
    28 <= n83;
    29 <= n88;
    30 <= n93;
    31 <= n98;
    32 <= n103;
    33 <= n108;
    34 <= n113;
  end
  initial begin
    2 <= 1'b0;
    20 <= 1'b0;
    21 <= 1'b0;
    22 <= 1'b0;
    23 <= 1'b0;
    24 <= 1'b0;
    25 <= 1'b0;
    26 <= 1'b0;
    27 <= 1'b0;
    28 <= 1'b0;
    29 <= 1'b0;
    30 <= 1'b0;
    31 <= 1'b0;
    32 <= 1'b0;
    33 <= 1'b0;
    34 <= 1'b0;
  end
endmodule

