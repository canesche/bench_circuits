module top ( clock, 
    pg7, pg6, pg5, pg4, pg3, pg2, pg1, pg0, pg9, pg8, pclk, pg10, pg12,
    pg11, pg14, pg13, pg16, pg15,
    pg701bf, pg702, pg726, pg727, pg729  );
  input  clock;
  input  pg7, pg6, pg5, pg4, pg3, pg2, pg1, pg0, pg9, pg8, pclk, pg10,
    pg12, pg11, pg14, pg13, pg16, pg15;
  output pg701bf, pg702, pg726, pg727, pg729;
  reg ng31, ng27, ng28, ng29, ng30, ng23, ng24, ng25, ng26, ng72, ng83,
    ng94, ng73, ng82, ng95, ng74, ng85, ng92, ng22, ng75, ng84, ng93, ng32,
    ng43, ng54, ng65, ng33, ng42, ng55, ng64, ng34, ng45, ng52, ng63, ng35,
    ng44, ng53, ng62, ng36, ng47, ng58, ng69, ng80, ng91, ng37, ng46, ng59,
    ng68, ng81, ng90, ng38, ng49, ng56, ng67, ng39, ng48, ng57, ng66, ng40,
    ng51, ng76, ng87, ng41, ng50, ng77, ng86, ng60, ng71, ng78, ng89, ng61,
    ng70, ng79, ng88;
  wire new_n246_, new_n247_, new_n248_1_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_1_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_1_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_1_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_1_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_1_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_1_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_1_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_1_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_1_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_1_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_1_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_1_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_1_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_1_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_1_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_1_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_1_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_1_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_1_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_1_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_1_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_1_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_1_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_1_, new_n374_, new_n375_, new_n376_, new_n378_1_, new_n379_,
    new_n381_, new_n382_, new_n384_, new_n385_, new_n387_, new_n388_1_,
    new_n390_, new_n391_, new_n393_1_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_1_, new_n399_, new_n400_, new_n401_, new_n403_1_,
    new_n404_, new_n405_, new_n407_, new_n408_1_, new_n410_, new_n411_,
    new_n413_1_, new_n414_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n445_,
    new_n446_, new_n447_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n455_, new_n456_, new_n457_, new_n458_, new_n460_,
    new_n461_, new_n463_, new_n464_, new_n465_, new_n467_, new_n468_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n477_,
    new_n478_, new_n479_, new_n481_, new_n482_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n509_, new_n510_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n527_, new_n529_, new_n530_, new_n532_, new_n533_,
    new_n535_, new_n536_, new_n537_, new_n539_, new_n540_, new_n541_,
    new_n543_, new_n544_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n557_,
    new_n560_, new_n561_, new_n563_, new_n564_, new_n565_, new_n567_,
    new_n568_, new_n570_, new_n571_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n594_, new_n595_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n605_,
    new_n606_, new_n607_, new_n609_, new_n610_, new_n612_, new_n613_,
    new_n615_, new_n616_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n636_, new_n637_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, n48, n53, n58, n63, n68, n73, n78,
    n83, n88, n93, n98, n103, n108, n113, n118, n123, n128, n133, n138,
    n143, n148, n153, n158, n163, n168, n173, n178, n183, n188, n193, n198,
    n203, n208, n213, n218, n223, n228, n233, n238, n243, n248, n253, n258,
    n263, n268, n273, n278, n283, n288, n293, n298, n303, n308, n313, n318,
    n323, n328, n333, n338, n343, n348, n353, n358, n363, n368, n373, n378,
    n383, n388, n393, n398, n403, n408, n413;
  assign new_n246_ = ~ng82 & ~ng80;
  assign new_n247_ = ~ng81 & new_n246_;
  assign new_n248_1_ = ~ng79 & new_n247_;
  assign new_n249_ = ~ng78 & ~new_n248_1_;
  assign new_n250_ = ng78 & new_n248_1_;
  assign new_n251_ = ~new_n249_ & ~new_n250_;
  assign new_n252_ = ~ng82 & ~ng77;
  assign new_n253_1_ = ng82 & ng77;
  assign new_n254_ = ~new_n252_ & ~new_n253_1_;
  assign new_n255_ = ~new_n251_ & ~new_n254_;
  assign new_n256_ = ~ng75 & ~ng80;
  assign new_n257_ = ng75 & ng80;
  assign new_n258_1_ = ~new_n256_ & ~new_n257_;
  assign new_n259_ = ~ng81 & ~ng76;
  assign new_n260_ = ng81 & ng76;
  assign new_n261_ = ~new_n259_ & ~new_n260_;
  assign new_n262_ = ~ng74 & ~ng79;
  assign new_n263_1_ = ng74 & ng79;
  assign new_n264_ = ~new_n262_ & ~new_n263_1_;
  assign new_n265_ = ~new_n258_1_ & ~new_n261_;
  assign new_n266_ = ~new_n264_ & new_n265_;
  assign new_n267_ = new_n255_ & new_n266_;
  assign new_n268_1_ = ~ng83 & new_n267_;
  assign new_n269_ = pg16 & ~ng66;
  assign new_n270_ = new_n268_1_ & new_n269_;
  assign new_n271_ = ng90 & ~new_n270_;
  assign new_n272_ = ~pg0 & ~ng90;
  assign new_n273_1_ = ~pg8 & ~ng90;
  assign new_n274_ = ng64 & ng90;
  assign new_n275_ = ~new_n273_1_ & ~new_n274_;
  assign new_n276_ = ~ng84 & new_n275_;
  assign new_n277_ = ~ng85 & ~new_n275_;
  assign new_n278_1_ = ~new_n276_ & ~new_n277_;
  assign new_n279_ = ng74 & new_n278_1_;
  assign new_n280_ = ng90 & new_n279_;
  assign new_n281_ = ~new_n272_ & ~new_n280_;
  assign new_n282_ = ~ng42 & ~new_n281_;
  assign new_n283_1_ = ng42 & new_n281_;
  assign new_n284_ = ~new_n282_ & ~new_n283_1_;
  assign new_n285_ = ~new_n282_ & ~new_n284_;
  assign new_n286_ = ~pg1 & ~ng90;
  assign new_n287_ = ng75 & new_n278_1_;
  assign new_n288_1_ = ng90 & new_n287_;
  assign new_n289_ = ~new_n286_ & ~new_n288_1_;
  assign new_n290_ = ~ng43 & ~new_n289_;
  assign new_n291_ = ng43 & new_n289_;
  assign new_n292_ = ~new_n290_ & ~new_n291_;
  assign new_n293_1_ = ~new_n285_ & new_n292_;
  assign new_n294_ = ~new_n290_ & ~new_n293_1_;
  assign new_n295_ = ~pg2 & ~ng90;
  assign new_n296_ = ng76 & new_n278_1_;
  assign new_n297_ = ng90 & new_n296_;
  assign new_n298_1_ = ~new_n295_ & ~new_n297_;
  assign new_n299_ = ~ng44 & ~new_n298_1_;
  assign new_n300_ = ng44 & new_n298_1_;
  assign new_n301_ = ~new_n299_ & ~new_n300_;
  assign new_n302_ = ~new_n294_ & new_n301_;
  assign new_n303_1_ = ~new_n299_ & ~new_n302_;
  assign new_n304_ = ~pg3 & ~ng90;
  assign new_n305_ = ng77 & new_n278_1_;
  assign new_n306_ = ng90 & new_n305_;
  assign new_n307_ = ~new_n304_ & ~new_n306_;
  assign new_n308_1_ = ~ng45 & ~new_n307_;
  assign new_n309_ = ng45 & new_n307_;
  assign new_n310_ = ~new_n308_1_ & ~new_n309_;
  assign new_n311_ = ~new_n303_1_ & new_n310_;
  assign new_n312_ = ~new_n308_1_ & ~new_n311_;
  assign new_n313_1_ = ~pg4 & ~ng90;
  assign new_n314_ = ng78 & new_n278_1_;
  assign new_n315_ = ng90 & new_n314_;
  assign new_n316_ = ~new_n313_1_ & ~new_n315_;
  assign new_n317_ = ~ng46 & ~new_n316_;
  assign new_n318_1_ = ng46 & new_n316_;
  assign new_n319_ = ~new_n317_ & ~new_n318_1_;
  assign new_n320_ = ~new_n312_ & new_n319_;
  assign new_n321_ = ~new_n317_ & ~new_n320_;
  assign new_n322_ = ~ng24 & ~new_n321_;
  assign new_n323_1_ = ng25 & new_n322_;
  assign new_n324_ = ng26 & new_n323_1_;
  assign new_n325_ = ~ng27 & new_n324_;
  assign new_n326_ = ng28 & new_n325_;
  assign new_n327_ = ng92 & ~new_n326_;
  assign new_n328_1_ = ~ng29 & ~new_n327_;
  assign new_n329_ = ng30 & new_n328_1_;
  assign new_n330_ = ng31 & new_n329_;
  assign new_n331_ = ng32 & new_n330_;
  assign new_n332_ = ng33 & new_n331_;
  assign new_n333_1_ = ~ng34 & new_n332_;
  assign new_n334_ = ng92 & ~new_n333_1_;
  assign new_n335_ = ~new_n271_ & new_n334_;
  assign new_n336_ = ~ng39 & ~new_n334_;
  assign new_n337_ = ~ng40 & new_n336_;
  assign new_n338_1_ = ng41 & new_n337_;
  assign new_n339_ = ng91 & ~new_n338_1_;
  assign new_n340_ = ~ng36 & ~new_n339_;
  assign new_n341_ = ng37 & new_n340_;
  assign new_n342_ = ng38 & new_n341_;
  assign new_n343_1_ = new_n271_ & ~new_n342_;
  assign new_n344_ = ~new_n335_ & ~new_n343_1_;
  assign new_n345_ = ng58 & new_n344_;
  assign new_n346_ = ng59 & new_n345_;
  assign new_n347_ = ng91 & ~new_n346_;
  assign new_n348_1_ = ng53 & ~new_n347_;
  assign new_n349_ = ng61 & new_n348_1_;
  assign new_n350_ = ng62 & new_n349_;
  assign new_n351_ = ng89 & new_n350_;
  assign new_n352_ = ng87 & new_n333_1_;
  assign new_n353_1_ = ng88 & new_n338_1_;
  assign new_n354_ = ~ng94 & new_n326_;
  assign new_n355_ = ~new_n351_ & ~new_n352_;
  assign new_n356_ = ~new_n353_1_ & new_n355_;
  assign new_n357_ = ~new_n354_ & new_n356_;
  assign pg702 = ~ng90 & new_n357_;
  assign new_n359_ = ~ng72 & ~ng73;
  assign new_n360_ = ~ng71 & new_n359_;
  assign new_n361_ = ~ng70 & ~new_n360_;
  assign new_n362_ = ng70 & new_n360_;
  assign new_n363_1_ = ~new_n361_ & ~new_n362_;
  assign new_n364_ = ~ng72 & ~ng68;
  assign new_n365_ = ng72 & ng68;
  assign new_n366_ = ~new_n364_ & ~new_n365_;
  assign new_n367_ = ~ng73 & ~ng69;
  assign new_n368_1_ = ng73 & ng69;
  assign new_n369_ = ~new_n367_ & ~new_n368_1_;
  assign new_n370_ = ~ng67 & ~ng71;
  assign new_n371_ = ng67 & ng71;
  assign new_n372_ = ~new_n370_ & ~new_n371_;
  assign new_n373_1_ = ~new_n363_1_ & ~new_n366_;
  assign new_n374_ = ~new_n369_ & ~new_n372_;
  assign new_n375_ = new_n373_1_ & new_n374_;
  assign new_n376_ = pg14 & ~new_n375_;
  assign pg727 = ~ng90 & ~new_n376_;
  assign new_n378_1_ = ~ng31 & ~new_n329_;
  assign new_n379_ = ~new_n330_ & ~new_n378_1_;
  assign n48 = pg14 & new_n379_;
  assign new_n381_ = ng27 & ~new_n324_;
  assign new_n382_ = ~new_n325_ & ~new_n381_;
  assign n53 = pg14 & ~new_n382_;
  assign new_n384_ = ~ng28 & ~new_n325_;
  assign new_n385_ = ~new_n326_ & ~new_n384_;
  assign n58 = pg14 & new_n385_;
  assign new_n387_ = ng29 & new_n327_;
  assign new_n388_1_ = ~new_n328_1_ & ~new_n387_;
  assign n63 = pg14 & ~new_n388_1_;
  assign new_n390_ = ~ng30 & ~new_n328_1_;
  assign new_n391_ = ~new_n329_ & ~new_n390_;
  assign n68 = pg14 & new_n391_;
  assign new_n393_1_ = ~ng47 & ~ng49;
  assign new_n394_ = ~ng48 & ~ng50;
  assign new_n395_ = new_n393_1_ & new_n394_;
  assign new_n396_ = ~pg15 & new_n395_;
  assign new_n397_ = ng22 & ~new_n396_;
  assign new_n398_1_ = ng47 & ng49;
  assign new_n399_ = ng48 & ng50;
  assign new_n400_ = new_n398_1_ & new_n399_;
  assign new_n401_ = ~pg15 & new_n400_;
  assign n138 = new_n397_ | new_n401_;
  assign new_n403_1_ = pg15 & n138;
  assign new_n404_ = ~ng23 & ~new_n403_1_;
  assign new_n405_ = pg15 & ~new_n397_;
  assign n73 = ~new_n404_ & ~new_n405_;
  assign new_n407_ = ng24 & new_n321_;
  assign new_n408_1_ = ~new_n322_ & ~new_n407_;
  assign n78 = pg14 & ~new_n408_1_;
  assign new_n410_ = ~ng25 & ~new_n322_;
  assign new_n411_ = ~new_n323_1_ & ~new_n410_;
  assign n83 = pg14 & new_n411_;
  assign new_n413_1_ = ~ng26 & ~new_n323_1_;
  assign new_n414_ = ~new_n324_ & ~new_n413_1_;
  assign n88 = pg14 & new_n414_;
  assign new_n416_ = ng90 & ~new_n376_;
  assign new_n417_ = pg14 & ~new_n416_;
  assign new_n418_ = ~pg1 & ~ng63;
  assign new_n419_ = ~pg4 & ng63;
  assign new_n420_ = ~new_n418_ & ~new_n419_;
  assign new_n421_ = ~new_n417_ & ~new_n420_;
  assign new_n422_ = ~ng72 & new_n417_;
  assign n93 = ~new_n421_ & ~new_n422_;
  assign new_n424_ = ~pg9 & ~ng90;
  assign new_n425_ = ng90 & new_n376_;
  assign new_n426_ = ~new_n424_ & ~new_n425_;
  assign new_n427_ = ng34 & new_n332_;
  assign new_n428_ = ng92 & ~new_n427_;
  assign new_n429_ = ~new_n271_ & new_n428_;
  assign new_n430_ = ~ng38 & new_n341_;
  assign new_n431_ = new_n271_ & ~new_n430_;
  assign new_n432_ = ~new_n429_ & ~new_n431_;
  assign new_n433_ = ~new_n267_ & new_n432_;
  assign new_n434_ = ~ng92 & ~ng35;
  assign new_n435_ = ng92 & ng34;
  assign new_n436_ = ~new_n434_ & ~new_n435_;
  assign new_n437_ = ~new_n271_ & ~new_n436_;
  assign new_n438_ = ~ng38 & new_n271_;
  assign new_n439_ = ~new_n437_ & ~new_n438_;
  assign new_n440_ = new_n267_ & ~new_n439_;
  assign new_n441_ = ~ng83 & ~new_n440_;
  assign new_n442_ = ~new_n440_ & ~new_n441_;
  assign new_n443_ = ~new_n433_ & ~new_n442_;
  assign n98 = ~new_n426_ & ~new_n443_;
  assign new_n445_ = ~pg11 & ~ng94;
  assign new_n446_ = pg11 & ng89;
  assign new_n447_ = ~new_n445_ & ~new_n446_;
  assign n103 = pg14 & new_n447_;
  assign new_n449_ = ~pg2 & ~ng63;
  assign new_n450_ = ~pg5 & ng63;
  assign new_n451_ = ~new_n449_ & ~new_n450_;
  assign new_n452_ = ~new_n417_ & ~new_n451_;
  assign new_n453_ = ~ng73 & new_n417_;
  assign n108 = ~new_n452_ & ~new_n453_;
  assign new_n455_ = ng91 & ~new_n376_;
  assign new_n456_ = pg14 & ~new_n455_;
  assign new_n457_ = ~pg9 & ~new_n456_;
  assign new_n458_ = ~ng82 & new_n456_;
  assign n113 = ~new_n457_ & ~new_n458_;
  assign new_n460_ = ng83 & new_n439_;
  assign new_n461_ = new_n278_1_ & new_n460_;
  assign n118 = pg14 & new_n461_;
  assign new_n463_ = ng74 & new_n433_;
  assign new_n464_ = ~ng74 & ~new_n433_;
  assign new_n465_ = ~new_n463_ & ~new_n464_;
  assign n123 = ~new_n426_ & new_n465_;
  assign new_n467_ = ~pg11 & ~new_n456_;
  assign new_n468_ = ~ng85 & new_n456_;
  assign n128 = ~new_n467_ & ~new_n468_;
  assign n373 = pg14 & pg13;
  assign new_n471_ = pg13 & ~ng86;
  assign new_n472_ = pg10 & ng91;
  assign new_n473_ = ~pg10 & ng92;
  assign new_n474_ = ~new_n472_ & ~new_n473_;
  assign new_n475_ = ~new_n471_ & ~new_n474_;
  assign n133 = ~n373 | new_n475_;
  assign new_n477_ = ng75 & new_n463_;
  assign new_n478_ = ~ng75 & ~new_n463_;
  assign new_n479_ = ~new_n477_ & ~new_n478_;
  assign n143 = ~new_n426_ & new_n479_;
  assign new_n481_ = ~pg10 & ~new_n456_;
  assign new_n482_ = ~ng84 & new_n456_;
  assign n148 = ~new_n481_ & ~new_n482_;
  assign new_n484_ = new_n284_ & new_n292_;
  assign new_n485_ = new_n301_ & new_n310_;
  assign new_n486_ = new_n319_ & new_n485_;
  assign new_n487_ = new_n484_ & new_n486_;
  assign new_n488_ = ~new_n321_ & ~new_n487_;
  assign new_n489_ = new_n439_ & ~new_n488_;
  assign new_n490_ = new_n487_ & new_n489_;
  assign new_n491_ = ~pg5 & ~ng90;
  assign new_n492_ = ng90 & new_n268_1_;
  assign new_n493_ = ~new_n491_ & ~new_n492_;
  assign new_n494_ = new_n439_ & new_n493_;
  assign new_n495_ = ~new_n490_ & ~new_n494_;
  assign new_n496_ = ~new_n321_ & new_n495_;
  assign new_n497_ = ~pg6 & ~ng90;
  assign new_n498_ = ~new_n271_ & ~new_n497_;
  assign new_n499_ = new_n496_ & ~new_n498_;
  assign new_n500_ = ~ng35 & ~ng90;
  assign new_n501_ = ~ng91 & ~ng59;
  assign new_n502_ = ~ng62 & ng91;
  assign new_n503_ = ~new_n501_ & ~new_n502_;
  assign new_n504_ = ng90 & ~new_n503_;
  assign new_n505_ = ~new_n500_ & ~new_n504_;
  assign new_n506_ = new_n498_ & new_n505_;
  assign new_n507_ = ~new_n499_ & ~new_n506_;
  assign n153 = pg14 & ~new_n507_;
  assign new_n509_ = ~ng32 & ~new_n330_;
  assign new_n510_ = ~new_n331_ & ~new_n509_;
  assign n158 = pg14 & new_n510_;
  assign new_n512_ = ~pg7 & ~ng90;
  assign new_n513_ = ~new_n425_ & ~new_n512_;
  assign new_n514_ = new_n400_ & ~n73;
  assign new_n515_ = ng42 & new_n514_;
  assign new_n516_ = ng43 & new_n515_;
  assign new_n517_ = ~ng43 & ~new_n515_;
  assign new_n518_ = ~new_n516_ & ~new_n517_;
  assign n163 = ~new_n513_ & new_n518_;
  assign new_n520_ = ng54 & ng56;
  assign new_n521_ = ~new_n334_ & new_n520_;
  assign new_n522_ = pg14 & ~new_n521_;
  assign new_n523_ = ng54 & ~new_n334_;
  assign new_n524_ = ~ng54 & new_n334_;
  assign new_n525_ = ~new_n523_ & ~new_n524_;
  assign n168 = new_n522_ & new_n525_;
  assign new_n527_ = ~ng65 & ~new_n375_;
  assign n173 = pg14 & ~new_n527_;
  assign new_n529_ = ~ng33 & ~new_n331_;
  assign new_n530_ = ~new_n332_ & ~new_n529_;
  assign n178 = pg14 & new_n530_;
  assign new_n532_ = ~ng42 & ~new_n514_;
  assign new_n533_ = ~new_n515_ & ~new_n532_;
  assign n183 = ~new_n513_ & new_n533_;
  assign new_n535_ = ng55 & new_n523_;
  assign new_n536_ = ~ng55 & ~new_n523_;
  assign new_n537_ = ~new_n535_ & ~new_n536_;
  assign n188 = new_n522_ & new_n537_;
  assign new_n539_ = ~ng64 & ~new_n375_;
  assign new_n540_ = ~ng63 & new_n375_;
  assign new_n541_ = ~new_n539_ & ~new_n540_;
  assign n193 = pg14 & new_n541_;
  assign new_n543_ = ng34 & ~new_n332_;
  assign new_n544_ = ~new_n333_1_ & ~new_n543_;
  assign n198 = pg14 & ~new_n544_;
  assign new_n546_ = ng44 & new_n516_;
  assign new_n547_ = ng45 & new_n546_;
  assign new_n548_ = ~ng45 & ~new_n546_;
  assign new_n549_ = ~new_n547_ & ~new_n548_;
  assign n203 = ~new_n513_ & new_n549_;
  assign new_n551_ = pg14 & ~new_n348_1_;
  assign new_n552_ = ng51 & ~new_n347_;
  assign new_n553_ = ng52 & new_n552_;
  assign new_n554_ = ~ng52 & ~new_n552_;
  assign new_n555_ = ~new_n553_ & ~new_n554_;
  assign n208 = new_n551_ & new_n555_;
  assign new_n557_ = ~ng63 & ~new_n439_;
  assign n213 = pg14 & ~new_n557_;
  assign n218 = pg14 & ~ng35;
  assign new_n560_ = ~ng44 & ~new_n516_;
  assign new_n561_ = ~new_n546_ & ~new_n560_;
  assign n223 = ~new_n513_ & new_n561_;
  assign new_n563_ = ng53 & new_n553_;
  assign new_n564_ = ~ng53 & ~new_n553_;
  assign new_n565_ = ~new_n563_ & ~new_n564_;
  assign n228 = new_n551_ & new_n565_;
  assign new_n567_ = ~ng62 & ~new_n349_;
  assign new_n568_ = ~new_n350_ & ~new_n567_;
  assign n233 = pg14 & new_n568_;
  assign new_n570_ = ng36 & new_n339_;
  assign new_n571_ = ~new_n340_ & ~new_n570_;
  assign n238 = pg14 & ~new_n571_;
  assign new_n573_ = ng91 & ~new_n521_;
  assign new_n574_ = ~pg12 & ~new_n573_;
  assign new_n575_ = ~ng47 & new_n573_;
  assign new_n576_ = ~new_n574_ & ~new_n575_;
  assign n243 = pg14 & new_n576_;
  assign new_n578_ = pg14 & ~new_n345_;
  assign new_n579_ = ng57 & new_n344_;
  assign new_n580_ = ng58 & new_n579_;
  assign new_n581_ = ~ng58 & ~new_n579_;
  assign new_n582_ = ~new_n580_ & ~new_n581_;
  assign n248 = new_n578_ & new_n582_;
  assign new_n584_ = ~ng91 & ~new_n346_;
  assign new_n585_ = ng91 & ~new_n350_;
  assign new_n586_ = ~new_n584_ & ~new_n585_;
  assign new_n587_ = ng90 & ~new_n586_;
  assign new_n588_ = ng67 & ~new_n587_;
  assign new_n589_ = ng68 & new_n588_;
  assign new_n590_ = ng69 & new_n589_;
  assign new_n591_ = ~ng69 & ~new_n589_;
  assign new_n592_ = ~new_n590_ & ~new_n591_;
  assign n253 = new_n376_ & new_n592_;
  assign new_n594_ = ~pg7 & ~new_n456_;
  assign new_n595_ = ~ng80 & new_n456_;
  assign n258 = ~new_n594_ & ~new_n595_;
  assign new_n597_ = pg10 & ng90;
  assign new_n598_ = ~pg10 & ng91;
  assign new_n599_ = ~new_n597_ & ~new_n598_;
  assign new_n600_ = ~new_n471_ & ~new_n599_;
  assign n263 = ~n373 | new_n600_;
  assign new_n602_ = ~ng37 & ~new_n340_;
  assign new_n603_ = ~new_n341_ & ~new_n602_;
  assign n268 = pg14 & new_n603_;
  assign new_n605_ = ng46 & new_n547_;
  assign new_n606_ = ~ng46 & ~new_n547_;
  assign new_n607_ = ~new_n605_ & ~new_n606_;
  assign n273 = ~new_n513_ & new_n607_;
  assign new_n609_ = ~ng59 & ~new_n345_;
  assign new_n610_ = ~new_n346_ & ~new_n609_;
  assign n278 = pg14 & new_n610_;
  assign new_n612_ = ~ng68 & ~new_n588_;
  assign new_n613_ = ~new_n589_ & ~new_n612_;
  assign n283 = new_n376_ & new_n613_;
  assign new_n615_ = ~pg8 & ~new_n456_;
  assign new_n616_ = ~ng81 & new_n456_;
  assign n288 = ~new_n615_ & ~new_n616_;
  assign new_n618_ = ~pg10 & ng90;
  assign new_n619_ = ~pg10 & ~new_n618_;
  assign new_n620_ = ~new_n471_ & ~new_n619_;
  assign n293 = ~n373 | new_n620_;
  assign new_n622_ = ~ng38 & ~new_n341_;
  assign new_n623_ = ~new_n342_ & ~new_n622_;
  assign n298 = pg14 & new_n623_;
  assign new_n625_ = ~ng48 & ~new_n573_;
  assign new_n626_ = ~ng49 & new_n573_;
  assign new_n627_ = ~new_n625_ & ~new_n626_;
  assign n303 = pg14 & new_n627_;
  assign new_n629_ = ng56 & new_n535_;
  assign new_n630_ = ~ng56 & ~new_n535_;
  assign new_n631_ = ~new_n629_ & ~new_n630_;
  assign n308 = new_n522_ & new_n631_;
  assign new_n633_ = ~ng67 & new_n587_;
  assign new_n634_ = ~new_n588_ & ~new_n633_;
  assign n313 = new_n376_ & new_n634_;
  assign new_n636_ = ng39 & new_n334_;
  assign new_n637_ = ~new_n336_ & ~new_n636_;
  assign n318 = pg14 & ~new_n637_;
  assign new_n639_ = ~ng47 & ~new_n573_;
  assign new_n640_ = ~ng48 & new_n573_;
  assign new_n641_ = ~new_n639_ & ~new_n640_;
  assign n323 = pg14 & new_n641_;
  assign new_n643_ = ~ng57 & ~new_n344_;
  assign new_n644_ = ~new_n579_ & ~new_n643_;
  assign n328 = new_n578_ & new_n644_;
  assign new_n646_ = ~ng66 & ~new_n375_;
  assign new_n647_ = ~ng65 & new_n375_;
  assign new_n648_ = ~new_n646_ & ~new_n647_;
  assign n333 = pg14 & new_n648_;
  assign new_n650_ = ng40 & ~new_n336_;
  assign new_n651_ = ~new_n337_ & ~new_n650_;
  assign n338 = pg14 & ~new_n651_;
  assign new_n653_ = ~ng51 & new_n347_;
  assign new_n654_ = ~new_n552_ & ~new_n653_;
  assign n343 = new_n551_ & new_n654_;
  assign new_n656_ = ng76 & new_n477_;
  assign new_n657_ = ~ng76 & ~new_n477_;
  assign new_n658_ = ~new_n656_ & ~new_n657_;
  assign n348 = ~new_n426_ & new_n658_;
  assign new_n660_ = pg11 & ng94;
  assign new_n661_ = ~pg11 & ~ng87;
  assign new_n662_ = ~new_n660_ & ~new_n661_;
  assign n353 = pg14 & new_n662_;
  assign new_n664_ = ~ng41 & ~new_n337_;
  assign new_n665_ = ~new_n338_1_ & ~new_n664_;
  assign n358 = pg14 & new_n665_;
  assign new_n667_ = ~ng49 & ~new_n573_;
  assign new_n668_ = ~ng50 & new_n573_;
  assign new_n669_ = ~new_n667_ & ~new_n668_;
  assign n363 = pg14 & new_n669_;
  assign new_n671_ = ng77 & new_n656_;
  assign new_n672_ = ~ng77 & ~new_n656_;
  assign new_n673_ = ~new_n671_ & ~new_n672_;
  assign n368 = ~new_n426_ & new_n673_;
  assign new_n675_ = pg14 & ~new_n349_;
  assign new_n676_ = ng60 & new_n348_1_;
  assign new_n677_ = ~ng60 & ~new_n348_1_;
  assign new_n678_ = ~new_n676_ & ~new_n677_;
  assign n378 = new_n675_ & new_n678_;
  assign new_n680_ = ~pg0 & ~ng63;
  assign new_n681_ = ~pg3 & ng63;
  assign new_n682_ = ~new_n680_ & ~new_n681_;
  assign new_n683_ = ~new_n417_ & ~new_n682_;
  assign new_n684_ = ~ng71 & new_n417_;
  assign n383 = ~new_n683_ & ~new_n684_;
  assign new_n686_ = ng78 & new_n671_;
  assign new_n687_ = ~ng78 & ~new_n671_;
  assign new_n688_ = ~new_n686_ & ~new_n687_;
  assign n388 = ~new_n426_ & new_n688_;
  assign new_n690_ = pg11 & ~ng88;
  assign new_n691_ = ~pg11 & ~ng89;
  assign new_n692_ = ~new_n690_ & ~new_n691_;
  assign n393 = pg14 & new_n692_;
  assign new_n694_ = ng61 & new_n676_;
  assign new_n695_ = ~ng61 & ~new_n676_;
  assign new_n696_ = ~new_n694_ & ~new_n695_;
  assign n398 = new_n675_ & new_n696_;
  assign new_n698_ = ng70 & new_n590_;
  assign new_n699_ = ~ng70 & ~new_n590_;
  assign new_n700_ = ~new_n698_ & ~new_n699_;
  assign n403 = new_n376_ & new_n700_;
  assign new_n702_ = ~pg6 & ~new_n456_;
  assign new_n703_ = ~ng79 & new_n456_;
  assign n408 = ~new_n702_ & ~new_n703_;
  assign new_n705_ = pg11 & ~ng87;
  assign new_n706_ = ~pg11 & ~ng88;
  assign new_n707_ = ~new_n705_ & ~new_n706_;
  assign n413 = pg14 & new_n707_;
  assign pg701bf = ~pg15;
  assign pg726 = ng93;
  assign pg729 = ng95;
  always @ (posedge clock) begin
    ng31 <= n48;
    ng27 <= n53;
    ng28 <= n58;
    ng29 <= n63;
    ng30 <= n68;
    ng23 <= n73;
    ng24 <= n78;
    ng25 <= n83;
    ng26 <= n88;
    ng72 <= n93;
    ng83 <= n98;
    ng94 <= n103;
    ng73 <= n108;
    ng82 <= n113;
    ng95 <= n118;
    ng74 <= n123;
    ng85 <= n128;
    ng92 <= n133;
    ng22 <= n138;
    ng75 <= n143;
    ng84 <= n148;
    ng93 <= n153;
    ng32 <= n158;
    ng43 <= n163;
    ng54 <= n168;
    ng65 <= n173;
    ng33 <= n178;
    ng42 <= n183;
    ng55 <= n188;
    ng64 <= n193;
    ng34 <= n198;
    ng45 <= n203;
    ng52 <= n208;
    ng63 <= n213;
    ng35 <= n218;
    ng44 <= n223;
    ng53 <= n228;
    ng62 <= n233;
    ng36 <= n238;
    ng47 <= n243;
    ng58 <= n248;
    ng69 <= n253;
    ng80 <= n258;
    ng91 <= n263;
    ng37 <= n268;
    ng46 <= n273;
    ng59 <= n278;
    ng68 <= n283;
    ng81 <= n288;
    ng90 <= n293;
    ng38 <= n298;
    ng49 <= n303;
    ng56 <= n308;
    ng67 <= n313;
    ng39 <= n318;
    ng48 <= n323;
    ng57 <= n328;
    ng66 <= n333;
    ng40 <= n338;
    ng51 <= n343;
    ng76 <= n348;
    ng87 <= n353;
    ng41 <= n358;
    ng50 <= n363;
    ng77 <= n368;
    ng86 <= n373;
    ng60 <= n378;
    ng71 <= n383;
    ng78 <= n388;
    ng89 <= n393;
    ng61 <= n398;
    ng70 <= n403;
    ng79 <= n408;
    ng88 <= n413;
  end
endmodule

