// Benchmark "wb_dma" written by ABC on Thu Oct  8 22:04:31 2020

module wb_dma ( clock, 
    clk_i, rst_i, wb0_we_i, wb0_cyc_i, wb0_stb_i, wb0_ack_i, wb0_err_i,
    wb0_rty_i, wb1_we_i, wb1_cyc_i, wb1_stb_i, wb1_ack_i, wb1_err_i,
    wb1_rty_i, \wb0s_data_i[0] , \wb0s_data_i[1] , \wb0s_data_i[2] ,
    \wb0s_data_i[3] , \wb0s_data_i[4] , \wb0s_data_i[5] , \wb0s_data_i[6] ,
    \wb0s_data_i[7] , \wb0s_data_i[8] , \wb0s_data_i[9] ,
    \wb0s_data_i[10] , \wb0s_data_i[11] , \wb0s_data_i[12] ,
    \wb0s_data_i[13] , \wb0s_data_i[14] , \wb0s_data_i[15] ,
    \wb0s_data_i[16] , \wb0s_data_i[17] , \wb0s_data_i[18] ,
    \wb0s_data_i[19] , \wb0s_data_i[20] , \wb0s_data_i[21] ,
    \wb0s_data_i[22] , \wb0s_data_i[23] , \wb0s_data_i[24] ,
    \wb0s_data_i[25] , \wb0s_data_i[26] , \wb0s_data_i[27] ,
    \wb0s_data_i[28] , \wb0s_data_i[29] , \wb0s_data_i[30] ,
    \wb0s_data_i[31] , \wb0_addr_i[0] , \wb0_addr_i[1] , \wb0_addr_i[2] ,
    \wb0_addr_i[3] , \wb0_addr_i[4] , \wb0_addr_i[5] , \wb0_addr_i[6] ,
    \wb0_addr_i[7] , \wb0_addr_i[8] , \wb0_addr_i[9] , \wb0_addr_i[10] ,
    \wb0_addr_i[11] , \wb0_addr_i[12] , \wb0_addr_i[13] , \wb0_addr_i[14] ,
    \wb0_addr_i[15] , \wb0_addr_i[16] , \wb0_addr_i[17] , \wb0_addr_i[18] ,
    \wb0_addr_i[19] , \wb0_addr_i[20] , \wb0_addr_i[21] , \wb0_addr_i[22] ,
    \wb0_addr_i[23] , \wb0_addr_i[24] , \wb0_addr_i[25] , \wb0_addr_i[26] ,
    \wb0_addr_i[27] , \wb0_addr_i[28] , \wb0_addr_i[29] , \wb0_addr_i[30] ,
    \wb0_addr_i[31] , \wb0m_data_i[0] , \wb0m_data_i[1] , \wb0m_data_i[2] ,
    \wb0m_data_i[3] , \wb0m_data_i[4] , \wb0m_data_i[5] , \wb0m_data_i[6] ,
    \wb0m_data_i[7] , \wb0m_data_i[8] , \wb0m_data_i[9] ,
    \wb0m_data_i[10] , \wb0m_data_i[11] , \wb0m_data_i[12] ,
    \wb0m_data_i[13] , \wb0m_data_i[14] , \wb0m_data_i[15] ,
    \wb0m_data_i[16] , \wb0m_data_i[17] , \wb0m_data_i[18] ,
    \wb0m_data_i[19] , \wb0m_data_i[20] , \wb0m_data_i[21] ,
    \wb0m_data_i[22] , \wb0m_data_i[23] , \wb0m_data_i[24] ,
    \wb0m_data_i[25] , \wb0m_data_i[26] , \wb0m_data_i[27] ,
    \wb0m_data_i[28] , \wb0m_data_i[29] , \wb0m_data_i[30] ,
    \wb0m_data_i[31] , \wb1s_data_i[0] , \wb1s_data_i[1] ,
    \wb1s_data_i[2] , \wb1s_data_i[3] , \wb1s_data_i[4] , \wb1s_data_i[5] ,
    \wb1s_data_i[6] , \wb1s_data_i[7] , \wb1s_data_i[8] , \wb1s_data_i[9] ,
    \wb1s_data_i[10] , \wb1s_data_i[11] , \wb1s_data_i[12] ,
    \wb1s_data_i[13] , \wb1s_data_i[14] , \wb1s_data_i[15] ,
    \wb1s_data_i[16] , \wb1s_data_i[17] , \wb1s_data_i[18] ,
    \wb1s_data_i[19] , \wb1s_data_i[20] , \wb1s_data_i[21] ,
    \wb1s_data_i[22] , \wb1s_data_i[23] , \wb1s_data_i[24] ,
    \wb1s_data_i[25] , \wb1s_data_i[26] , \wb1s_data_i[27] ,
    \wb1s_data_i[28] , \wb1s_data_i[29] , \wb1s_data_i[30] ,
    \wb1s_data_i[31] , \wb1_addr_i[0] , \wb1_addr_i[1] , \wb1_addr_i[2] ,
    \wb1_addr_i[3] , \wb1_addr_i[4] , \wb1_addr_i[5] , \wb1_addr_i[6] ,
    \wb1_addr_i[7] , \wb1_addr_i[8] , \wb1_addr_i[9] , \wb1_addr_i[10] ,
    \wb1_addr_i[11] , \wb1_addr_i[12] , \wb1_addr_i[13] , \wb1_addr_i[14] ,
    \wb1_addr_i[15] , \wb1_addr_i[16] , \wb1_addr_i[17] , \wb1_addr_i[18] ,
    \wb1_addr_i[19] , \wb1_addr_i[20] , \wb1_addr_i[21] , \wb1_addr_i[22] ,
    \wb1_addr_i[23] , \wb1_addr_i[24] , \wb1_addr_i[25] , \wb1_addr_i[26] ,
    \wb1_addr_i[27] , \wb1_addr_i[28] , \wb1_addr_i[29] , \wb1_addr_i[30] ,
    \wb1_addr_i[31] , \wb1m_data_i[0] , \wb1m_data_i[1] , \wb1m_data_i[2] ,
    \wb1m_data_i[3] , \wb1m_data_i[4] , \wb1m_data_i[5] , \wb1m_data_i[6] ,
    \wb1m_data_i[7] , \wb1m_data_i[8] , \wb1m_data_i[9] ,
    \wb1m_data_i[10] , \wb1m_data_i[11] , \wb1m_data_i[12] ,
    \wb1m_data_i[13] , \wb1m_data_i[14] , \wb1m_data_i[15] ,
    \wb1m_data_i[16] , \wb1m_data_i[17] , \wb1m_data_i[18] ,
    \wb1m_data_i[19] , \wb1m_data_i[20] , \wb1m_data_i[21] ,
    \wb1m_data_i[22] , \wb1m_data_i[23] , \wb1m_data_i[24] ,
    \wb1m_data_i[25] , \wb1m_data_i[26] , \wb1m_data_i[27] ,
    \wb1m_data_i[28] , \wb1m_data_i[29] , \wb1m_data_i[30] ,
    \wb1m_data_i[31] , \wb0_sel_i[0] , \wb0_sel_i[1] , \wb0_sel_i[2] ,
    \wb0_sel_i[3] , \wb1_sel_i[0] , \wb1_sel_i[1] , \wb1_sel_i[2] ,
    \wb1_sel_i[3] , dma_req_i, dma_nd_i, dma_rest_i,
    \wb0s_data_o[0] , \wb0s_data_o[1] , \wb0s_data_o[2] , \wb0s_data_o[3] ,
    \wb0s_data_o[4] , \wb0s_data_o[5] , \wb0s_data_o[6] , \wb0s_data_o[7] ,
    \wb0s_data_o[8] , \wb0s_data_o[9] , \wb0s_data_o[10] ,
    \wb0s_data_o[11] , \wb0s_data_o[12] , \wb0s_data_o[13] ,
    \wb0s_data_o[14] , \wb0s_data_o[15] , \wb0s_data_o[16] ,
    \wb0s_data_o[17] , \wb0s_data_o[18] , \wb0s_data_o[19] ,
    \wb0s_data_o[20] , \wb0s_data_o[21] , \wb0s_data_o[22] ,
    \wb0s_data_o[23] , \wb0s_data_o[24] , \wb0s_data_o[25] ,
    \wb0s_data_o[26] , \wb0s_data_o[27] , \wb0s_data_o[28] ,
    \wb0s_data_o[29] , \wb0s_data_o[30] , \wb0s_data_o[31] ,
    \wb0m_data_o[0] , \wb0m_data_o[1] , \wb0m_data_o[2] , \wb0m_data_o[3] ,
    \wb0m_data_o[4] , \wb0m_data_o[5] , \wb0m_data_o[6] , \wb0m_data_o[7] ,
    \wb0m_data_o[8] , \wb0m_data_o[9] , \wb0m_data_o[10] ,
    \wb0m_data_o[11] , \wb0m_data_o[12] , \wb0m_data_o[13] ,
    \wb0m_data_o[14] , \wb0m_data_o[15] , \wb0m_data_o[16] ,
    \wb0m_data_o[17] , \wb0m_data_o[18] , \wb0m_data_o[19] ,
    \wb0m_data_o[20] , \wb0m_data_o[21] , \wb0m_data_o[22] ,
    \wb0m_data_o[23] , \wb0m_data_o[24] , \wb0m_data_o[25] ,
    \wb0m_data_o[26] , \wb0m_data_o[27] , \wb0m_data_o[28] ,
    \wb0m_data_o[29] , \wb0m_data_o[30] , \wb0m_data_o[31] ,
    \wb0_addr_o[0] , \wb0_addr_o[1] , \wb0_addr_o[2] , \wb0_addr_o[3] ,
    \wb0_addr_o[4] , \wb0_addr_o[5] , \wb0_addr_o[6] , \wb0_addr_o[7] ,
    \wb0_addr_o[8] , \wb0_addr_o[9] , \wb0_addr_o[10] , \wb0_addr_o[11] ,
    \wb0_addr_o[12] , \wb0_addr_o[13] , \wb0_addr_o[14] , \wb0_addr_o[15] ,
    \wb0_addr_o[16] , \wb0_addr_o[17] , \wb0_addr_o[18] , \wb0_addr_o[19] ,
    \wb0_addr_o[20] , \wb0_addr_o[21] , \wb0_addr_o[22] , \wb0_addr_o[23] ,
    \wb0_addr_o[24] , \wb0_addr_o[25] , \wb0_addr_o[26] , \wb0_addr_o[27] ,
    \wb0_addr_o[28] , \wb0_addr_o[29] , \wb0_addr_o[30] , \wb0_addr_o[31] ,
    \wb1s_data_o[0] , \wb1s_data_o[1] , \wb1s_data_o[2] , \wb1s_data_o[3] ,
    \wb1s_data_o[4] , \wb1s_data_o[5] , \wb1s_data_o[6] , \wb1s_data_o[7] ,
    \wb1s_data_o[8] , \wb1s_data_o[9] , \wb1s_data_o[10] ,
    \wb1s_data_o[11] , \wb1s_data_o[12] , \wb1s_data_o[13] ,
    \wb1s_data_o[14] , \wb1s_data_o[15] , \wb1s_data_o[16] ,
    \wb1s_data_o[17] , \wb1s_data_o[18] , \wb1s_data_o[19] ,
    \wb1s_data_o[20] , \wb1s_data_o[21] , \wb1s_data_o[22] ,
    \wb1s_data_o[23] , \wb1s_data_o[24] , \wb1s_data_o[25] ,
    \wb1s_data_o[26] , \wb1s_data_o[27] , \wb1s_data_o[28] ,
    \wb1s_data_o[29] , \wb1s_data_o[30] , \wb1s_data_o[31] ,
    \wb1m_data_o[0] , \wb1m_data_o[1] , \wb1m_data_o[2] , \wb1m_data_o[3] ,
    \wb1m_data_o[4] , \wb1m_data_o[5] , \wb1m_data_o[6] , \wb1m_data_o[7] ,
    \wb1m_data_o[8] , \wb1m_data_o[9] , \wb1m_data_o[10] ,
    \wb1m_data_o[11] , \wb1m_data_o[12] , \wb1m_data_o[13] ,
    \wb1m_data_o[14] , \wb1m_data_o[15] , \wb1m_data_o[16] ,
    \wb1m_data_o[17] , \wb1m_data_o[18] , \wb1m_data_o[19] ,
    \wb1m_data_o[20] , \wb1m_data_o[21] , \wb1m_data_o[22] ,
    \wb1m_data_o[23] , \wb1m_data_o[24] , \wb1m_data_o[25] ,
    \wb1m_data_o[26] , \wb1m_data_o[27] , \wb1m_data_o[28] ,
    \wb1m_data_o[29] , \wb1m_data_o[30] , \wb1m_data_o[31] ,
    \wb1_addr_o[0] , \wb1_addr_o[1] , \wb1_addr_o[2] , \wb1_addr_o[3] ,
    \wb1_addr_o[4] , \wb1_addr_o[5] , \wb1_addr_o[6] , \wb1_addr_o[7] ,
    \wb1_addr_o[8] , \wb1_addr_o[9] , \wb1_addr_o[10] , \wb1_addr_o[11] ,
    \wb1_addr_o[12] , \wb1_addr_o[13] , \wb1_addr_o[14] , \wb1_addr_o[15] ,
    \wb1_addr_o[16] , \wb1_addr_o[17] , \wb1_addr_o[18] , \wb1_addr_o[19] ,
    \wb1_addr_o[20] , \wb1_addr_o[21] , \wb1_addr_o[22] , \wb1_addr_o[23] ,
    \wb1_addr_o[24] , \wb1_addr_o[25] , \wb1_addr_o[26] , \wb1_addr_o[27] ,
    \wb1_addr_o[28] , \wb1_addr_o[29] , \wb1_addr_o[30] , \wb1_addr_o[31] ,
    wb0_ack_o, wb0_err_o, wb0_rty_o, wb0_we_o, wb0_cyc_o, wb0_stb_o,
    wb1_ack_o, wb1_err_o, wb1_rty_o, wb1_we_o, wb1_cyc_o, wb1_stb_o,
    inta_o, intb_o, \wb0_sel_o[0] , \wb0_sel_o[1] , \wb0_sel_o[2] ,
    \wb0_sel_o[3] , \wb1_sel_o[0] , \wb1_sel_o[1] , \wb1_sel_o[2] ,
    \wb1_sel_o[3] , dma_ack_o  );
  input  clock;
  input  clk_i, rst_i, wb0_we_i, wb0_cyc_i, wb0_stb_i, wb0_ack_i,
    wb0_err_i, wb0_rty_i, wb1_we_i, wb1_cyc_i, wb1_stb_i, wb1_ack_i,
    wb1_err_i, wb1_rty_i, \wb0s_data_i[0] , \wb0s_data_i[1] ,
    \wb0s_data_i[2] , \wb0s_data_i[3] , \wb0s_data_i[4] , \wb0s_data_i[5] ,
    \wb0s_data_i[6] , \wb0s_data_i[7] , \wb0s_data_i[8] , \wb0s_data_i[9] ,
    \wb0s_data_i[10] , \wb0s_data_i[11] , \wb0s_data_i[12] ,
    \wb0s_data_i[13] , \wb0s_data_i[14] , \wb0s_data_i[15] ,
    \wb0s_data_i[16] , \wb0s_data_i[17] , \wb0s_data_i[18] ,
    \wb0s_data_i[19] , \wb0s_data_i[20] , \wb0s_data_i[21] ,
    \wb0s_data_i[22] , \wb0s_data_i[23] , \wb0s_data_i[24] ,
    \wb0s_data_i[25] , \wb0s_data_i[26] , \wb0s_data_i[27] ,
    \wb0s_data_i[28] , \wb0s_data_i[29] , \wb0s_data_i[30] ,
    \wb0s_data_i[31] , \wb0_addr_i[0] , \wb0_addr_i[1] , \wb0_addr_i[2] ,
    \wb0_addr_i[3] , \wb0_addr_i[4] , \wb0_addr_i[5] , \wb0_addr_i[6] ,
    \wb0_addr_i[7] , \wb0_addr_i[8] , \wb0_addr_i[9] , \wb0_addr_i[10] ,
    \wb0_addr_i[11] , \wb0_addr_i[12] , \wb0_addr_i[13] , \wb0_addr_i[14] ,
    \wb0_addr_i[15] , \wb0_addr_i[16] , \wb0_addr_i[17] , \wb0_addr_i[18] ,
    \wb0_addr_i[19] , \wb0_addr_i[20] , \wb0_addr_i[21] , \wb0_addr_i[22] ,
    \wb0_addr_i[23] , \wb0_addr_i[24] , \wb0_addr_i[25] , \wb0_addr_i[26] ,
    \wb0_addr_i[27] , \wb0_addr_i[28] , \wb0_addr_i[29] , \wb0_addr_i[30] ,
    \wb0_addr_i[31] , \wb0m_data_i[0] , \wb0m_data_i[1] , \wb0m_data_i[2] ,
    \wb0m_data_i[3] , \wb0m_data_i[4] , \wb0m_data_i[5] , \wb0m_data_i[6] ,
    \wb0m_data_i[7] , \wb0m_data_i[8] , \wb0m_data_i[9] ,
    \wb0m_data_i[10] , \wb0m_data_i[11] , \wb0m_data_i[12] ,
    \wb0m_data_i[13] , \wb0m_data_i[14] , \wb0m_data_i[15] ,
    \wb0m_data_i[16] , \wb0m_data_i[17] , \wb0m_data_i[18] ,
    \wb0m_data_i[19] , \wb0m_data_i[20] , \wb0m_data_i[21] ,
    \wb0m_data_i[22] , \wb0m_data_i[23] , \wb0m_data_i[24] ,
    \wb0m_data_i[25] , \wb0m_data_i[26] , \wb0m_data_i[27] ,
    \wb0m_data_i[28] , \wb0m_data_i[29] , \wb0m_data_i[30] ,
    \wb0m_data_i[31] , \wb1s_data_i[0] , \wb1s_data_i[1] ,
    \wb1s_data_i[2] , \wb1s_data_i[3] , \wb1s_data_i[4] , \wb1s_data_i[5] ,
    \wb1s_data_i[6] , \wb1s_data_i[7] , \wb1s_data_i[8] , \wb1s_data_i[9] ,
    \wb1s_data_i[10] , \wb1s_data_i[11] , \wb1s_data_i[12] ,
    \wb1s_data_i[13] , \wb1s_data_i[14] , \wb1s_data_i[15] ,
    \wb1s_data_i[16] , \wb1s_data_i[17] , \wb1s_data_i[18] ,
    \wb1s_data_i[19] , \wb1s_data_i[20] , \wb1s_data_i[21] ,
    \wb1s_data_i[22] , \wb1s_data_i[23] , \wb1s_data_i[24] ,
    \wb1s_data_i[25] , \wb1s_data_i[26] , \wb1s_data_i[27] ,
    \wb1s_data_i[28] , \wb1s_data_i[29] , \wb1s_data_i[30] ,
    \wb1s_data_i[31] , \wb1_addr_i[0] , \wb1_addr_i[1] , \wb1_addr_i[2] ,
    \wb1_addr_i[3] , \wb1_addr_i[4] , \wb1_addr_i[5] , \wb1_addr_i[6] ,
    \wb1_addr_i[7] , \wb1_addr_i[8] , \wb1_addr_i[9] , \wb1_addr_i[10] ,
    \wb1_addr_i[11] , \wb1_addr_i[12] , \wb1_addr_i[13] , \wb1_addr_i[14] ,
    \wb1_addr_i[15] , \wb1_addr_i[16] , \wb1_addr_i[17] , \wb1_addr_i[18] ,
    \wb1_addr_i[19] , \wb1_addr_i[20] , \wb1_addr_i[21] , \wb1_addr_i[22] ,
    \wb1_addr_i[23] , \wb1_addr_i[24] , \wb1_addr_i[25] , \wb1_addr_i[26] ,
    \wb1_addr_i[27] , \wb1_addr_i[28] , \wb1_addr_i[29] , \wb1_addr_i[30] ,
    \wb1_addr_i[31] , \wb1m_data_i[0] , \wb1m_data_i[1] , \wb1m_data_i[2] ,
    \wb1m_data_i[3] , \wb1m_data_i[4] , \wb1m_data_i[5] , \wb1m_data_i[6] ,
    \wb1m_data_i[7] , \wb1m_data_i[8] , \wb1m_data_i[9] ,
    \wb1m_data_i[10] , \wb1m_data_i[11] , \wb1m_data_i[12] ,
    \wb1m_data_i[13] , \wb1m_data_i[14] , \wb1m_data_i[15] ,
    \wb1m_data_i[16] , \wb1m_data_i[17] , \wb1m_data_i[18] ,
    \wb1m_data_i[19] , \wb1m_data_i[20] , \wb1m_data_i[21] ,
    \wb1m_data_i[22] , \wb1m_data_i[23] , \wb1m_data_i[24] ,
    \wb1m_data_i[25] , \wb1m_data_i[26] , \wb1m_data_i[27] ,
    \wb1m_data_i[28] , \wb1m_data_i[29] , \wb1m_data_i[30] ,
    \wb1m_data_i[31] , \wb0_sel_i[0] , \wb0_sel_i[1] , \wb0_sel_i[2] ,
    \wb0_sel_i[3] , \wb1_sel_i[0] , \wb1_sel_i[1] , \wb1_sel_i[2] ,
    \wb1_sel_i[3] , dma_req_i, dma_nd_i, dma_rest_i;
  output \wb0s_data_o[0] , \wb0s_data_o[1] , \wb0s_data_o[2] ,
    \wb0s_data_o[3] , \wb0s_data_o[4] , \wb0s_data_o[5] , \wb0s_data_o[6] ,
    \wb0s_data_o[7] , \wb0s_data_o[8] , \wb0s_data_o[9] ,
    \wb0s_data_o[10] , \wb0s_data_o[11] , \wb0s_data_o[12] ,
    \wb0s_data_o[13] , \wb0s_data_o[14] , \wb0s_data_o[15] ,
    \wb0s_data_o[16] , \wb0s_data_o[17] , \wb0s_data_o[18] ,
    \wb0s_data_o[19] , \wb0s_data_o[20] , \wb0s_data_o[21] ,
    \wb0s_data_o[22] , \wb0s_data_o[23] , \wb0s_data_o[24] ,
    \wb0s_data_o[25] , \wb0s_data_o[26] , \wb0s_data_o[27] ,
    \wb0s_data_o[28] , \wb0s_data_o[29] , \wb0s_data_o[30] ,
    \wb0s_data_o[31] , \wb0m_data_o[0] , \wb0m_data_o[1] ,
    \wb0m_data_o[2] , \wb0m_data_o[3] , \wb0m_data_o[4] , \wb0m_data_o[5] ,
    \wb0m_data_o[6] , \wb0m_data_o[7] , \wb0m_data_o[8] , \wb0m_data_o[9] ,
    \wb0m_data_o[10] , \wb0m_data_o[11] , \wb0m_data_o[12] ,
    \wb0m_data_o[13] , \wb0m_data_o[14] , \wb0m_data_o[15] ,
    \wb0m_data_o[16] , \wb0m_data_o[17] , \wb0m_data_o[18] ,
    \wb0m_data_o[19] , \wb0m_data_o[20] , \wb0m_data_o[21] ,
    \wb0m_data_o[22] , \wb0m_data_o[23] , \wb0m_data_o[24] ,
    \wb0m_data_o[25] , \wb0m_data_o[26] , \wb0m_data_o[27] ,
    \wb0m_data_o[28] , \wb0m_data_o[29] , \wb0m_data_o[30] ,
    \wb0m_data_o[31] , \wb0_addr_o[0] , \wb0_addr_o[1] , \wb0_addr_o[2] ,
    \wb0_addr_o[3] , \wb0_addr_o[4] , \wb0_addr_o[5] , \wb0_addr_o[6] ,
    \wb0_addr_o[7] , \wb0_addr_o[8] , \wb0_addr_o[9] , \wb0_addr_o[10] ,
    \wb0_addr_o[11] , \wb0_addr_o[12] , \wb0_addr_o[13] , \wb0_addr_o[14] ,
    \wb0_addr_o[15] , \wb0_addr_o[16] , \wb0_addr_o[17] , \wb0_addr_o[18] ,
    \wb0_addr_o[19] , \wb0_addr_o[20] , \wb0_addr_o[21] , \wb0_addr_o[22] ,
    \wb0_addr_o[23] , \wb0_addr_o[24] , \wb0_addr_o[25] , \wb0_addr_o[26] ,
    \wb0_addr_o[27] , \wb0_addr_o[28] , \wb0_addr_o[29] , \wb0_addr_o[30] ,
    \wb0_addr_o[31] , \wb1s_data_o[0] , \wb1s_data_o[1] , \wb1s_data_o[2] ,
    \wb1s_data_o[3] , \wb1s_data_o[4] , \wb1s_data_o[5] , \wb1s_data_o[6] ,
    \wb1s_data_o[7] , \wb1s_data_o[8] , \wb1s_data_o[9] ,
    \wb1s_data_o[10] , \wb1s_data_o[11] , \wb1s_data_o[12] ,
    \wb1s_data_o[13] , \wb1s_data_o[14] , \wb1s_data_o[15] ,
    \wb1s_data_o[16] , \wb1s_data_o[17] , \wb1s_data_o[18] ,
    \wb1s_data_o[19] , \wb1s_data_o[20] , \wb1s_data_o[21] ,
    \wb1s_data_o[22] , \wb1s_data_o[23] , \wb1s_data_o[24] ,
    \wb1s_data_o[25] , \wb1s_data_o[26] , \wb1s_data_o[27] ,
    \wb1s_data_o[28] , \wb1s_data_o[29] , \wb1s_data_o[30] ,
    \wb1s_data_o[31] , \wb1m_data_o[0] , \wb1m_data_o[1] ,
    \wb1m_data_o[2] , \wb1m_data_o[3] , \wb1m_data_o[4] , \wb1m_data_o[5] ,
    \wb1m_data_o[6] , \wb1m_data_o[7] , \wb1m_data_o[8] , \wb1m_data_o[9] ,
    \wb1m_data_o[10] , \wb1m_data_o[11] , \wb1m_data_o[12] ,
    \wb1m_data_o[13] , \wb1m_data_o[14] , \wb1m_data_o[15] ,
    \wb1m_data_o[16] , \wb1m_data_o[17] , \wb1m_data_o[18] ,
    \wb1m_data_o[19] , \wb1m_data_o[20] , \wb1m_data_o[21] ,
    \wb1m_data_o[22] , \wb1m_data_o[23] , \wb1m_data_o[24] ,
    \wb1m_data_o[25] , \wb1m_data_o[26] , \wb1m_data_o[27] ,
    \wb1m_data_o[28] , \wb1m_data_o[29] , \wb1m_data_o[30] ,
    \wb1m_data_o[31] , \wb1_addr_o[0] , \wb1_addr_o[1] , \wb1_addr_o[2] ,
    \wb1_addr_o[3] , \wb1_addr_o[4] , \wb1_addr_o[5] , \wb1_addr_o[6] ,
    \wb1_addr_o[7] , \wb1_addr_o[8] , \wb1_addr_o[9] , \wb1_addr_o[10] ,
    \wb1_addr_o[11] , \wb1_addr_o[12] , \wb1_addr_o[13] , \wb1_addr_o[14] ,
    \wb1_addr_o[15] , \wb1_addr_o[16] , \wb1_addr_o[17] , \wb1_addr_o[18] ,
    \wb1_addr_o[19] , \wb1_addr_o[20] , \wb1_addr_o[21] , \wb1_addr_o[22] ,
    \wb1_addr_o[23] , \wb1_addr_o[24] , \wb1_addr_o[25] , \wb1_addr_o[26] ,
    \wb1_addr_o[27] , \wb1_addr_o[28] , \wb1_addr_o[29] , \wb1_addr_o[30] ,
    \wb1_addr_o[31] , wb0_ack_o, wb0_err_o, wb0_rty_o, wb0_we_o, wb0_cyc_o,
    wb0_stb_o, wb1_ack_o, wb1_err_o, wb1_rty_o, wb1_we_o, wb1_cyc_o,
    wb1_stb_o, inta_o, intb_o, \wb0_sel_o[0] , \wb0_sel_o[1] ,
    \wb0_sel_o[2] , \wb0_sel_o[3] , \wb1_sel_o[0] , \wb1_sel_o[1] ,
    \wb1_sel_o[2] , \wb1_sel_o[3] , dma_ack_o;
  reg u3_u0_mast_stb_reg, u4_u0_mast_stb_reg, u3_u0_mast_cyc_reg,
    u4_u0_mast_cyc_reg, \\u2_mast0_adr_reg[3] , \\u2_mast0_adr_reg[2] ,
    \\u2_mast0_adr_reg[23] , \\u2_mast0_adr_reg[22] ,
    \\u2_mast0_adr_reg[21] , \\u2_mast0_adr_reg[25] ,
    \\u2_mast0_adr_reg[20] , \\u2_mast0_adr_reg[19] ,
    \\u2_mast0_adr_reg[18] , \\u2_mast0_adr_reg[16] ,
    \\u2_mast0_adr_reg[15] , \\u2_mast0_adr_reg[14] ,
    \\u2_mast0_adr_reg[13] , \\u2_mast0_adr_reg[12] ,
    \\u2_mast0_adr_reg[11] , \\u2_mast0_adr_reg[10] ,
    \\u2_mast0_adr_reg[9] , \\u2_mast0_adr_reg[6] , \\u2_mast0_adr_reg[5] ,
    \\u2_mast0_adr_reg[4] , \\u2_mast0_adr_reg[29] ,
    \\u2_mast0_adr_reg[28] , \\u2_mast0_adr_reg[27] ,
    \\u2_mast0_adr_reg[26] , \\u2_mast0_adr_reg[24] ,
    \\u2_mast0_adr_reg[17] , \\u2_mast0_adr_reg[7] ,
    \\u2_mast0_adr_reg[8] , \\u2_mast1_adr_reg[29] ,
    \\u2_mast1_adr_reg[28] , \\u2_mast1_adr_reg[27] ,
    \\u2_mast1_adr_reg[26] , \\u2_mast1_adr_reg[25] ,
    \\u2_mast1_adr_reg[24] , \\u2_mast1_adr_reg[22] ,
    \\u2_mast1_adr_reg[23] , \\u2_mast1_adr_reg[21] ,
    \\u2_mast1_adr_reg[20] , \\u2_mast1_adr_reg[19] ,
    \\u2_mast1_adr_reg[18] , \\u2_mast1_adr_reg[16] ,
    \\u2_mast1_adr_reg[15] , \\u2_mast1_adr_reg[13] ,
    \\u2_mast1_adr_reg[12] , \\u2_mast1_adr_reg[14] ,
    \\u2_mast1_adr_reg[11] , \\u2_mast1_adr_reg[10] ,
    \\u2_mast1_adr_reg[9] , \\u2_mast1_adr_reg[6] , \\u2_mast1_adr_reg[5] ,
    \\u2_mast1_adr_reg[4] , \\u2_mast0_adr_reg[31] ,
    \\u2_mast0_adr_reg[30] , \\u2_mast1_adr_reg[31] ,
    \\u2_mast1_adr_reg[30] , \\u2_mast1_adr_reg[17] ,
    \\u2_mast1_adr_reg[8] , \\u2_mast1_adr_reg[7] , \\u2_mast1_adr_reg[3] ,
    \\u2_mast1_adr_reg[2] , \\u2_state_reg[1] , \\u2_state_reg[3] ,
    u2_chunk_dec_reg, u2_tsz_dec_reg, \\u2_adr1_cnt_reg[28] ,
    \\u2_adr1_cnt_reg[27] , \\u2_adr1_cnt_reg[23] , \\u2_adr1_cnt_reg[24] ,
    \\u2_adr1_cnt_reg[20] , \\u2_adr1_cnt_reg[19] , \\u2_adr1_cnt_reg[18] ,
    \\u2_adr1_cnt_reg[25] , \\u2_adr1_cnt_reg[29] , \\u2_adr1_cnt_reg[17] ,
    \\u2_adr1_cnt_reg[21] , \\u2_adr1_cnt_reg[16] , \\u2_adr1_cnt_reg[2] ,
    \\u2_adr1_cnt_reg[3] , \\u2_adr1_cnt_reg[4] , \\u2_adr1_cnt_reg[5] ,
    \\u2_adr1_cnt_reg[6] , \\u2_adr1_cnt_reg[7] , \\u2_adr1_cnt_reg[8] ,
    \\u2_adr1_cnt_reg[9] , \\u2_adr1_cnt_reg[10] , \\u2_adr1_cnt_reg[11] ,
    \\u2_adr1_cnt_reg[13] , \\u2_adr1_cnt_reg[14] , \\u2_adr1_cnt_reg[15] ,
    u2_read_r_reg, \\u2_adr1_cnt_reg[26] , \\u2_adr1_cnt_reg[22] ,
    \\u2_adr1_cnt_reg[0] , \\u2_adr1_cnt_reg[12] , \\u2_adr1_cnt_reg[1] ,
    u2_write_hold_r_reg, u3_u0_mast_we_r_reg, \\u2_adr0_cnt_reg[16] ,
    \\u0_u0_int_src_r_reg[2] , \\u1_ack_o_reg[0] , u1_next_start_reg,
    \\u2_adr0_cnt_reg[9] , \\u2_adr0_cnt_reg[28] , \\u2_adr0_cnt_reg[27] ,
    \\u2_adr0_cnt_reg[24] , \\u2_adr0_cnt_reg[23] , \\u2_adr0_cnt_reg[26] ,
    \\u2_adr0_cnt_reg[20] , \\u2_adr0_cnt_reg[18] , \\u2_adr0_cnt_reg[10] ,
    \\u2_adr0_cnt_reg[11] , \\u2_adr0_cnt_reg[12] , \\u2_adr0_cnt_reg[13] ,
    \\u2_adr0_cnt_reg[17] , \\u2_adr0_cnt_reg[21] , \\u2_adr0_cnt_reg[25] ,
    \\u2_adr0_cnt_reg[2] , \\u2_adr0_cnt_reg[3] , \\u2_adr0_cnt_reg[5] ,
    \\u2_adr0_cnt_reg[6] , \\u2_adr0_cnt_reg[8] , \\u2_adr0_cnt_reg[7] ,
    \\u2_adr0_cnt_reg[4] , \\u0_u0_ch_csr_r_reg[0] ,
    \\u2_adr0_cnt_reg[14] , \\u2_adr0_cnt_reg[22] , \\u2_adr0_cnt_reg[19] ,
    \\u2_adr0_cnt_reg[29] , \\u2_adr0_cnt_reg[15] , u0_u0_ch_done_reg,
    u2_next_ch_reg, \\u0_u0_int_src_r_reg[1] , \\u2_state_reg[0] ,
    \\u2_state_reg[9] , \\u2_adr0_cnt_reg[0] , \\u2_adr0_cnt_reg[1] ,
    \\u2_tsz_cnt_reg[8] , \\u2_tsz_cnt_reg[2] , u4_u0_mast_we_r_reg,
    \\u0_wb_rf_dout_reg[10] , \\u2_state_reg[10] , \\u2_state_reg[4] ,
    \\u2_tsz_cnt_reg[0] , \\u2_tsz_cnt_reg[4] , \\u2_tsz_cnt_reg[5] ,
    \\u2_tsz_cnt_reg[6] , \\u2_tsz_cnt_reg[7] , \\u2_tsz_cnt_reg[10] ,
    \\u2_tsz_cnt_reg[11] , \\u2_tsz_cnt_reg[1] , \\u2_tsz_cnt_reg[3] ,
    \\u2_tsz_cnt_reg[9] , u2_chunk_0_reg, u2_write_r_reg,
    \\u2_state_reg[2] , \\u0_u0_ch_tot_sz_r_reg[0] ,
    \\u0_u0_ch_adr1_r_reg[25] , \\u0_u0_ch_adr0_r_reg[17] ,
    \\u0_u0_ch_adr0_r_reg[13] , \\u0_u0_ch_adr1_r_reg[29] ,
    \\u0_u0_ch_adr1_r_reg[21] , \\u0_u0_ch_adr1_r_reg[13] ,
    \\u0_u0_ch_adr1_r_reg[17] , \\u0_u0_ch_tot_sz_r_reg[1] ,
    \\u0_u0_ch_adr1_r_reg[10] , \\u0_u0_ch_adr1_r_reg[11] ,
    \\u0_u0_ch_adr1_r_reg[12] , \\u0_u0_ch_adr1_r_reg[14] ,
    \\u0_u0_ch_adr1_r_reg[15] , \\u0_u0_ch_adr1_r_reg[16] ,
    \\u0_u0_ch_adr1_r_reg[18] , \\u0_u0_ch_adr1_r_reg[19] ,
    \\u0_u0_ch_adr1_r_reg[20] , \\u0_u0_ch_adr1_r_reg[22] ,
    \\u0_u0_ch_adr1_r_reg[23] , \\u0_u0_ch_adr1_r_reg[24] ,
    \\u0_u0_ch_adr1_r_reg[26] , \\u0_u0_ch_adr1_r_reg[27] ,
    \\u0_u0_ch_adr1_r_reg[28] , \\u0_u0_ch_adr0_r_reg[10] ,
    \\u0_u0_ch_adr0_r_reg[11] , \\u0_u0_ch_adr0_r_reg[12] ,
    \\u0_u0_ch_adr0_r_reg[14] , \\u0_u0_ch_adr0_r_reg[15] ,
    \\u0_u0_ch_adr0_r_reg[16] , \\u0_u0_ch_adr0_r_reg[18] ,
    \\u0_u0_ch_adr0_r_reg[19] , \\u0_u0_ch_adr0_r_reg[20] ,
    \\u0_u0_ch_adr0_r_reg[22] , \\u0_u0_ch_adr0_r_reg[23] ,
    \\u0_u0_ch_adr0_r_reg[24] , \\u0_u0_ch_adr0_r_reg[26] ,
    \\u0_u0_ch_adr0_r_reg[27] , \\u0_u0_ch_adr0_r_reg[28] ,
    \\u0_u0_ch_adr0_r_reg[21] , \\u0_u0_ch_adr0_r_reg[29] ,
    \\u0_u0_ch_adr0_r_reg[25] , \\u0_u0_ch_tot_sz_r_reg[9] ,
    \\u0_u0_ch_tot_sz_r_reg[5] , \\u0_u0_ch_tot_sz_r_reg[10] ,
    \\u0_u0_ch_tot_sz_r_reg[11] , \\u0_u0_ch_tot_sz_r_reg[2] ,
    \\u0_u0_ch_tot_sz_r_reg[3] , \\u0_u0_ch_tot_sz_r_reg[4] ,
    \\u0_u0_ch_tot_sz_r_reg[6] , \\u0_u0_ch_tot_sz_r_reg[7] ,
    \\u0_u0_ch_tot_sz_r_reg[8] , \\u0_u0_ch_csr_r_reg[4] ,
    u0_u0_ch_err_reg, \\u0_u0_ch_csr_r_reg[1] , \\u0_u0_ch_csr_r_reg[2] ,
    \\u0_u0_ch_csr_r_reg[3] , \\u0_u0_ch_adr1_r_reg[0] ,
    \\u0_u0_ch_adr1_r_reg[1] , \\u0_u0_ch_adr1_r_reg[3] ,
    \\u0_u0_ch_adr1_r_reg[4] , \\u0_u0_ch_adr1_r_reg[5] ,
    \\u0_u0_ch_adr1_r_reg[7] , \\u0_u0_ch_adr1_r_reg[8] ,
    \\u0_u0_ch_adr1_r_reg[9] , \\u0_u0_ch_adr0_r_reg[9] ,
    \\u0_u0_ch_adr0_r_reg[0] , \\u0_u0_ch_adr0_r_reg[1] ,
    \\u0_u0_ch_adr0_r_reg[3] , \\u0_u0_ch_adr0_r_reg[4] ,
    \\u0_u0_ch_adr0_r_reg[5] , \\u0_u0_ch_adr0_r_reg[7] ,
    \\u0_u0_int_src_r_reg[0] , \\u0_u0_ch_adr0_r_reg[6] ,
    \\u0_u0_ch_adr0_r_reg[2] , \\u0_u0_ch_adr0_r_reg[8] ,
    \\u0_u0_ch_adr1_r_reg[6] , \\u0_u0_ch_adr1_r_reg[2] ,
    \\u2_chunk_cnt_reg[8] , \\u2_chunk_cnt_reg[7] , \\u2_chunk_cnt_reg[6] ,
    \\u1_ch_sel_r_reg[2] , \\u1_ch_sel_r_reg[1] , \\u1_ch_sel_r_reg[3] ,
    \\u1_ch_sel_r_reg[4] , \\u2_chunk_cnt_reg[1] , \\u2_chunk_cnt_reg[3] ,
    \\u2_chunk_cnt_reg[4] , \\u2_chunk_cnt_reg[0] , \\u2_chunk_cnt_reg[5] ,
    \\u2_chunk_cnt_reg[2] , \\u1_ch_sel_r_reg[0] ,
    \\u0_wb_rf_dout_reg[26] , \\u0_wb_rf_dout_reg[25] ,
    \\u0_wb_rf_dout_reg[24] , \\u0_wb_rf_dout_reg[23] ,
    \\u0_wb_rf_dout_reg[14] , \\u0_wb_rf_dout_reg[13] ,
    \\u0_wb_rf_dout_reg[12] , \\u0_wb_rf_dout_reg[3] ,
    \\u0_wb_rf_dout_reg[2] , \\u0_wb_rf_dout_reg[0] ,
    \\u0_wb_rf_dout_reg[22] , \\u0_wb_rf_dout_reg[21] ,
    \\u0_wb_rf_dout_reg[20] , \\u0_wb_rf_dout_reg[19] ,
    \\u0_wb_rf_dout_reg[18] , \\u0_wb_rf_dout_reg[17] ,
    \\u0_wb_rf_dout_reg[16] , \\u0_wb_rf_dout_reg[15] ,
    \\u0_wb_rf_dout_reg[11] , \\u0_wb_rf_dout_reg[8] ,
    \\u0_wb_rf_dout_reg[7] , \\u0_wb_rf_dout_reg[6] ,
    \\u0_wb_rf_dout_reg[5] , \\u0_wb_rf_dout_reg[4] , u0_u0_ch_busy_reg,
    \\u0_wb_rf_dout_reg[9] , \\u0_wb_rf_dout_reg[30] ,
    \\u0_wb_rf_dout_reg[29] , \\u0_wb_rf_dout_reg[28] ,
    \\u0_wb_rf_dout_reg[27] , \\u0_wb_rf_dout_reg[1] ,
    \\u0_wb_rf_dout_reg[31] , u2_tsz_cnt_is_0_r_reg, u2_dma_abort_r_reg,
    u1_de_start_r_reg, \\u2_state_reg[5] , \\u0_u0_ch_csr_r3_reg[2] ,
    \\u0_u0_ch_csr_r3_reg[0] , u0_u0_rest_en_reg, \\u0_u0_ch_csr_r_reg[7] ,
    \\u0_u0_ch_csr_r_reg[5] , \\u0_u0_ch_csr_r2_reg[2] ,
    \\u0_u0_ch_csr_r2_reg[1] , \\u0_u0_ch_csr_r2_reg[0] ,
    \\u0_u0_ch_csr_r3_reg[1] , \\u0_u0_ch_csr_r_reg[6] ,
    \\u0_u0_ch_csr_r_reg[8] , u0_u0_ch_stop_reg, u0_u0_ch_sz_inf_reg,
    \\u1_u1_state_reg[2] , \\u1_u1_state_reg[3] ,
    \\u0_u0_ch_chk_sz_r_reg[5] , \\u0_u0_ch_chk_sz_r_reg[3] ,
    \\u0_u0_ch_chk_sz_r_reg[7] , \\u0_u0_ch_chk_sz_r_reg[1] ,
    \\u0_u0_ch_chk_sz_r_reg[2] , \\u1_u1_state_reg[4] ,
    \\u0_u0_ch_chk_sz_r_reg[4] , \\u0_u0_ch_chk_sz_r_reg[6] ,
    \\u0_u0_ch_chk_sz_r_reg[0] , \\u1_u1_state_reg[0] ,
    \\u1_u1_state_reg[1] , u4_u1_rf_ack_reg, \\u0_u0_ch_chk_sz_r_reg[10] ,
    \\u0_u0_ch_chk_sz_r_reg[8] , \\u0_u0_ch_chk_sz_r_reg[9] ,
    \\u2_u0_out_r_reg[15] , \\u2_u1_out_r_reg[15] , \\u2_state_reg[8] ,
    \\u2_state_reg[7] , \\u2_state_reg[6] , \\u2_u0_out_r_reg[11] ,
    \\u2_u1_out_r_reg[11] , \\u2_u0_out_r_reg[12] , \\u2_u1_out_r_reg[12] ,
    \\u2_u0_out_r_reg[16] , \\u2_u1_out_r_reg[16] ,
    \\u0_int_maska_r_reg[11] , \\u0_csr_r_reg[0] ,
    \\u0_int_maska_r_reg[0] , \\u2_u0_out_r_reg[14] ,
    \\u2_u1_out_r_reg[14] , \\u0_int_maska_r_reg[10] ,
    \\u0_int_maska_r_reg[5] , \\u2_u1_out_r_reg[8] , \\u2_u0_out_r_reg[8] ,
    \\u0_int_maska_r_reg[6] , \\u0_int_maska_r_reg[7] ,
    \\u0_int_maska_r_reg[8] , \\u0_int_maska_r_reg[9] ,
    \\u0_int_maska_r_reg[2] , \\u0_int_maska_r_reg[4] ,
    \\u0_int_maska_r_reg[3] , \\u0_int_maska_r_reg[29] ,
    \\u0_int_maska_r_reg[26] , \\u0_int_maska_r_reg[27] ,
    \\u0_int_maska_r_reg[28] , \\u0_int_maska_r_reg[19] ,
    \\u0_int_maska_r_reg[22] , \\u0_int_maska_r_reg[24] ,
    \\u0_int_maska_r_reg[23] , \\u0_int_maska_r_reg[1] ,
    \\u0_int_maska_r_reg[20] , \\u0_int_maska_r_reg[16] ,
    \\u0_int_maska_r_reg[17] , \\u0_int_maska_r_reg[15] ,
    \\u0_int_maska_r_reg[12] , \\u0_int_maska_r_reg[13] ,
    \\u0_int_maska_r_reg[14] , \\u0_int_maskb_r_reg[6] ,
    \\u0_int_maskb_r_reg[9] , \\u2_u1_out_r_reg[7] , \\u2_u0_out_r_reg[7] ,
    \\u0_int_maska_r_reg[18] , \\u0_int_maska_r_reg[21] ,
    \\u0_int_maska_r_reg[25] , \\u0_int_maska_r_reg[30] ,
    \\u0_int_maskb_r_reg[0] , \\u0_int_maskb_r_reg[7] ,
    \\u0_int_maskb_r_reg[8] , \\u0_int_maskb_r_reg[5] ,
    \\u0_int_maskb_r_reg[11] , \\u0_int_maskb_r_reg[10] ,
    \\u0_int_maskb_r_reg[14] , \\u0_int_maskb_r_reg[17] ,
    \\u0_int_maskb_r_reg[20] , \\u0_int_maskb_r_reg[22] ,
    \\u0_int_maskb_r_reg[2] , \\u0_int_maskb_r_reg[12] ,
    \\u0_int_maskb_r_reg[18] , \\u0_int_maskb_r_reg[19] ,
    \\u0_int_maskb_r_reg[15] , \\u2_u0_out_r_reg[13] ,
    \\u2_u1_out_r_reg[13] , \\u0_int_maskb_r_reg[24] ,
    \\u0_int_maskb_r_reg[30] , \\u0_int_maskb_r_reg[3] ,
    \\u0_int_maskb_r_reg[4] , \\u0_int_maskb_r_reg[25] ,
    \\u0_int_maskb_r_reg[28] , \\u0_int_maskb_r_reg[29] ,
    \\u0_int_maskb_r_reg[26] , \\u0_int_maskb_r_reg[27] ,
    \\u0_int_maskb_r_reg[23] , \\u0_int_maskb_r_reg[1] ,
    \\u0_int_maskb_r_reg[21] , \\u0_int_maskb_r_reg[16] ,
    \\u0_int_maskb_r_reg[13] , u2_chunk_cnt_is_0_r_reg,
    \\u2_u1_out_r_reg[4] , \\u2_u0_out_r_reg[4] , \\u2_u1_out_r_reg[10] ,
    \\u2_u0_out_r_reg[10] , u4_u1_slv_we_reg, u3_u1_slv_re_reg,
    u4_u1_slv_re_reg, u3_u1_slv_we_reg, \\u3_u0_mast_dout_reg[4] ,
    \\u3_u0_mast_dout_reg[28] , \\u3_u0_mast_dout_reg[19] ,
    \\u3_u0_mast_dout_reg[29] , u0_inta_o_reg, \\u3_u0_mast_dout_reg[1] ,
    \\u3_u0_mast_dout_reg[8] , \\u3_u0_mast_dout_reg[30] ,
    \\u3_u0_mast_dout_reg[3] , \\u3_u0_mast_dout_reg[22] ,
    \\u3_u0_mast_dout_reg[18] , \\u3_u0_mast_dout_reg[10] ,
    \\u3_u0_mast_dout_reg[12] , \\u3_u0_mast_dout_reg[0] ,
    \\u3_u0_mast_dout_reg[15] , \\u3_u0_mast_dout_reg[20] ,
    \\u3_u0_mast_dout_reg[25] , \\u3_u0_mast_dout_reg[14] ,
    \\u3_u0_mast_dout_reg[9] , \\u3_u0_mast_dout_reg[13] ,
    \\u3_u0_mast_dout_reg[11] , \\u3_u0_mast_dout_reg[17] ,
    \\u3_u0_mast_dout_reg[2] , \\u2_u1_out_r_reg[3] ,
    \\u3_u0_mast_dout_reg[31] , \\u3_u0_mast_dout_reg[6] ,
    \\u3_u0_mast_dout_reg[27] , \\u3_u0_mast_dout_reg[23] ,
    \\u3_u0_mast_dout_reg[24] , u0_intb_o_reg, \\u2_u0_out_r_reg[3] ,
    \\u3_u0_mast_dout_reg[21] , \\u3_u0_mast_dout_reg[7] ,
    \\u2_u1_out_r_reg[6] , \\u2_u0_out_r_reg[6] ,
    \\u3_u0_mast_dout_reg[5] , \\u2_u1_out_r_reg[9] ,
    \\u2_u0_out_r_reg[9] , \\u3_u0_mast_dout_reg[26] ,
    \\u3_u0_mast_dout_reg[16] , \\u2_u0_out_r_reg[5] ,
    \\u2_u1_out_r_reg[5] , \\u2_u1_out_r_reg[2] , \\u2_u0_out_r_reg[2] ,
    u2_mast0_drdy_r_reg, u3_u1_rf_ack_reg, \\u4_u0_mast_dout_reg[23] ,
    \\u4_u0_mast_dout_reg[20] , \\u4_u0_mast_dout_reg[16] ,
    \\u4_u0_mast_dout_reg[22] , \\u4_u0_mast_dout_reg[5] ,
    \\u4_u0_mast_dout_reg[11] , \\u4_u0_mast_dout_reg[12] ,
    \\u4_u0_mast_dout_reg[7] , \\u4_u0_mast_dout_reg[3] ,
    \\u4_u0_mast_dout_reg[13] , \\u4_u0_mast_dout_reg[4] ,
    \\u4_u0_mast_dout_reg[27] , \\u4_u0_mast_dout_reg[1] ,
    \\u4_u0_mast_dout_reg[26] , \\u4_u0_mast_dout_reg[25] ,
    \\u4_u0_mast_dout_reg[21] , \\u4_u0_mast_dout_reg[2] ,
    \\u4_u0_mast_dout_reg[24] , \\u4_u0_mast_dout_reg[0] ,
    \\u4_u0_mast_dout_reg[17] , \\u4_u0_mast_dout_reg[31] ,
    \\u4_u0_mast_dout_reg[14] , \\u4_u0_mast_dout_reg[8] ,
    \\u4_u0_mast_dout_reg[28] , \\u4_u0_mast_dout_reg[10] ,
    \\u4_u0_mast_dout_reg[18] , \\u4_u0_mast_dout_reg[29] ,
    \\u4_u0_mast_dout_reg[6] , \\u4_u0_mast_dout_reg[9] ,
    \\u4_u0_mast_dout_reg[19] , \\u4_u0_mast_dout_reg[15] ,
    \\u4_u0_mast_dout_reg[30] , \\u2_u0_out_r_reg[1] ,
    \\u2_u1_out_r_reg[1] , \\u1_ndr_r_reg[2] , \\u1_ndr_r_reg[1] ,
    \\u1_ndr_r_reg[24] , \\u1_ndr_r_reg[10] , \\u1_ndr_r_reg[11] ,
    \\u1_ndr_r_reg[12] , \\u1_ndr_r_reg[29] , \\u1_ndr_r_reg[17] ,
    \\u1_ndr_r_reg[9] , \\u1_ndr_r_reg[22] , \\u1_ndr_r_reg[7] ,
    \\u1_ndr_r_reg[30] , \\u1_ndr_r_reg[23] , \\u1_ndr_r_reg[15] ,
    \\u1_ndr_r_reg[14] , \\u1_ndr_r_reg[28] , \\u1_ndr_r_reg[18] ,
    \\u1_ndr_r_reg[16] , \\u1_ndr_r_reg[8] , \\u1_ndr_r_reg[4] ,
    \\u1_ndr_r_reg[27] , \\u1_ndr_r_reg[20] , \\u1_ndr_r_reg[5] ,
    \\u1_ndr_r_reg[6] , \\u1_ndr_r_reg[19] , \\u1_ndr_r_reg[21] ,
    \\u1_ndr_r_reg[25] , \\u1_ndr_r_reg[13] , \\u1_ndr_r_reg[3] ,
    \\u1_ndr_r_reg[26] , \\u1_ndr_r_reg[0] , \\u1_ndnr_reg[0] ,
    \\u2_u0_out_r_reg[0] , \\u2_u1_out_r_reg[0] , \\u1_req_r_reg[0] ,
    \\u3_u1_slv_adr_reg[3] , \\u3_u1_slv_dout_reg[4] ,
    \\u3_u1_slv_dout_reg[0] , \\u3_u1_slv_dout_reg[18] ,
    \\u3_u1_slv_dout_reg[7] , \\u3_u1_slv_adr_reg[6] ,
    \\u3_u1_slv_dout_reg[5] , \\u3_u1_slv_dout_reg[24] ,
    \\u3_u1_slv_dout_reg[1] , \\u3_u1_slv_adr_reg[8] ,
    \\u3_u1_slv_dout_reg[19] , \\u3_u1_slv_dout_reg[31] ,
    \\u3_u1_slv_dout_reg[6] , \\u3_u1_slv_adr_reg[9] ,
    \\u3_u1_slv_dout_reg[20] , \\u3_u1_slv_adr_reg[4] ,
    \\u3_u1_slv_dout_reg[30] , \\u3_u1_slv_dout_reg[26] ,
    \\u3_u1_slv_dout_reg[29] , \\u3_u1_slv_dout_reg[28] ,
    \\u3_u1_slv_dout_reg[2] , \\u3_u1_slv_dout_reg[8] ,
    \\u3_u1_slv_adr_reg[7] , \\u3_u1_slv_adr_reg[2] ,
    \\u3_u1_slv_dout_reg[14] , \\u3_u1_slv_dout_reg[23] ,
    \\u3_u1_slv_dout_reg[9] , \\u3_u1_slv_dout_reg[21] ,
    \\u3_u1_slv_dout_reg[25] , \\u3_u1_slv_dout_reg[27] ,
    \\u3_u1_slv_dout_reg[3] , \\u3_u1_slv_dout_reg[12] ,
    \\u3_u1_slv_dout_reg[17] , \\u3_u1_slv_adr_reg[5] ,
    \\u3_u1_slv_dout_reg[11] , \\u3_u1_slv_dout_reg[15] ,
    \\u3_u1_slv_dout_reg[13] , \\u3_u1_slv_dout_reg[10] ,
    \\u3_u1_slv_dout_reg[16] , \\u3_u1_slv_dout_reg[22] ;
  wire \new_[1001]_ , \new_[1025]_ , \new_[1030]_ , \new_[1058]_ ,
    \new_[1060]_ , \new_[1061]_ , \new_[1067]_ , \new_[1068]_ ,
    \new_[1069]_ , \new_[1070]_ , \new_[1071]_ , \new_[1072]_ ,
    \new_[1073]_ , \new_[1074]_ , \new_[1075]_ , \new_[1076]_ ,
    \new_[1077]_ , \new_[1078]_ , \new_[1079]_ , \new_[1080]_ ,
    \new_[1081]_ , \new_[1082]_ , \new_[1083]_ , \new_[1084]_ ,
    \new_[1089]_ , \new_[1090]_ , \new_[1091]_ , \new_[1092]_ ,
    \new_[1093]_ , \new_[1094]_ , \new_[1095]_ , \new_[1096]_ ,
    \new_[1097]_ , \new_[1098]_ , \new_[1099]_ , \new_[1100]_ ,
    \new_[1101]_ , \new_[1102]_ , \new_[1103]_ , \new_[1104]_ ,
    \new_[1105]_ , \new_[1106]_ , \new_[1107]_ , \new_[1108]_ ,
    \new_[1109]_ , \new_[1110]_ , \new_[1111]_ , \new_[1112]_ ,
    \new_[1113]_ , \new_[1114]_ , \new_[1115]_ , \new_[1116]_ ,
    \new_[1117]_ , \new_[1118]_ , \new_[1119]_ , \new_[1120]_ ,
    \new_[1123]_ , \new_[1124]_ , \new_[1148]_ , \new_[1149]_ ,
    \new_[1150]_ , \new_[1151]_ , \new_[1152]_ , \new_[1157]_ ,
    \new_[1159]_ , \new_[1162]_ , \new_[1165]_ , \new_[1166]_ ,
    \new_[1167]_ , \new_[1168]_ , \new_[1189]_ , \new_[1190]_ ,
    \new_[1191]_ , \new_[1194]_ , \new_[1195]_ , \new_[1196]_ ,
    \new_[1197]_ , \new_[1198]_ , \new_[1199]_ , \new_[1200]_ ,
    \new_[1201]_ , \new_[1202]_ , \new_[1203]_ , \new_[1204]_ ,
    \new_[1205]_ , \new_[1206]_ , \new_[1207]_ , \new_[1209]_ ,
    \new_[1210]_ , \new_[1211]_ , \new_[1212]_ , \new_[1213]_ ,
    \new_[1214]_ , \new_[1215]_ , \new_[1216]_ , \new_[1217]_ ,
    \new_[1218]_ , \new_[1219]_ , \new_[1220]_ , \new_[1222]_ ,
    \new_[1224]_ , \new_[1225]_ , \new_[1226]_ , \new_[1227]_ ,
    \new_[1228]_ , \new_[1229]_ , \new_[1230]_ , \new_[1231]_ ,
    \new_[1232]_ , \new_[1233]_ , \new_[1234]_ , \new_[1235]_ ,
    \new_[1236]_ , \new_[1237]_ , \new_[1238]_ , \new_[1239]_ ,
    \new_[1240]_ , \new_[1241]_ , \new_[1242]_ , \new_[1243]_ ,
    \new_[1244]_ , \new_[1245]_ , \new_[1246]_ , \new_[1247]_ ,
    \new_[1248]_ , \new_[1249]_ , \new_[1250]_ , \new_[1251]_ ,
    \new_[1252]_ , \new_[1253]_ , \new_[1255]_ , \new_[1256]_ ,
    \new_[1258]_ , \new_[1259]_ , \new_[1260]_ , \new_[1261]_ ,
    \new_[1262]_ , \new_[1263]_ , \new_[1264]_ , \new_[1265]_ ,
    \new_[1266]_ , \new_[1267]_ , \new_[1268]_ , \new_[1269]_ ,
    \new_[1270]_ , \new_[1271]_ , \new_[1272]_ , \new_[1273]_ ,
    \new_[1274]_ , \new_[1275]_ , \new_[1276]_ , \new_[1277]_ ,
    \new_[1278]_ , \new_[1279]_ , \new_[1280]_ , \new_[1281]_ ,
    \new_[1282]_ , \new_[1284]_ , \new_[1285]_ , \new_[1287]_ ,
    \new_[1288]_ , \new_[1291]_ , \new_[1292]_ , \new_[1317]_ ,
    \new_[1318]_ , \new_[1319]_ , \new_[1320]_ , \new_[1324]_ ,
    \new_[1325]_ , \new_[1326]_ , \new_[1327]_ , \new_[1329]_ ,
    \new_[1331]_ , \new_[1332]_ , \new_[1333]_ , \new_[1334]_ ,
    \new_[1335]_ , \new_[1337]_ , \new_[1338]_ , \new_[1339]_ ,
    \new_[1340]_ , \new_[1342]_ , \new_[1343]_ , \new_[1344]_ ,
    \new_[1345]_ , \new_[1346]_ , \new_[1347]_ , \new_[1348]_ ,
    \new_[1349]_ , \new_[1350]_ , \new_[1351]_ , \new_[1352]_ ,
    \new_[1353]_ , \new_[1354]_ , \new_[1355]_ , \new_[1356]_ ,
    \new_[1357]_ , \new_[1358]_ , \new_[1359]_ , \new_[1360]_ ,
    \new_[1361]_ , \new_[1362]_ , \new_[1363]_ , \new_[1364]_ ,
    \new_[1365]_ , \new_[1366]_ , \new_[1367]_ , \new_[1368]_ ,
    \new_[1369]_ , \new_[1370]_ , \new_[1371]_ , \new_[1372]_ ,
    \new_[1373]_ , \new_[1374]_ , \new_[1375]_ , \new_[1376]_ ,
    \new_[1377]_ , \new_[1378]_ , \new_[1379]_ , \new_[1380]_ ,
    \new_[1381]_ , \new_[1382]_ , \new_[1383]_ , \new_[1384]_ ,
    \new_[1385]_ , \new_[1386]_ , \new_[1387]_ , \new_[1388]_ ,
    \new_[1389]_ , \new_[1390]_ , \new_[1403]_ , \new_[1404]_ ,
    \new_[1405]_ , \new_[1406]_ , \new_[1407]_ , \new_[1411]_ ,
    \new_[1412]_ , \new_[1413]_ , \new_[1414]_ , \new_[1415]_ ,
    \new_[1416]_ , \new_[1417]_ , \new_[1434]_ , \new_[1436]_ ,
    \new_[1437]_ , \new_[1439]_ , \new_[1440]_ , \new_[1443]_ ,
    \new_[1444]_ , \new_[1445]_ , \new_[1447]_ , \new_[1448]_ ,
    \new_[1449]_ , \new_[1450]_ , \new_[1451]_ , \new_[1452]_ ,
    \new_[1453]_ , \new_[1454]_ , \new_[1455]_ , \new_[1456]_ ,
    \new_[1458]_ , \new_[1459]_ , \new_[1460]_ , \new_[1461]_ ,
    \new_[1462]_ , \new_[1464]_ , \new_[1465]_ , \new_[1470]_ ,
    \new_[1471]_ , \new_[1488]_ , \new_[1490]_ , \new_[1491]_ ,
    \new_[1492]_ , \new_[1493]_ , \new_[1494]_ , \new_[1495]_ ,
    \new_[1496]_ , \new_[1498]_ , \new_[1499]_ , \new_[1500]_ ,
    \new_[1501]_ , \new_[1502]_ , \new_[1503]_ , \new_[1504]_ ,
    \new_[1505]_ , \new_[1506]_ , \new_[1507]_ , \new_[1508]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1512]_ ,
    \new_[1516]_ , \new_[1517]_ , \new_[1518]_ , \new_[1519]_ ,
    \new_[1520]_ , \new_[1521]_ , \new_[1522]_ , \new_[1523]_ ,
    \new_[1524]_ , \new_[1525]_ , \new_[1526]_ , \new_[1527]_ ,
    \new_[1528]_ , \new_[1529]_ , \new_[1530]_ , \new_[1531]_ ,
    \new_[1532]_ , \new_[1533]_ , \new_[1535]_ , \new_[1536]_ ,
    \new_[1537]_ , \new_[1538]_ , \new_[1539]_ , \new_[1540]_ ,
    \new_[1541]_ , \new_[1542]_ , \new_[1543]_ , \new_[1547]_ ,
    \new_[1548]_ , \new_[1549]_ , \new_[1550]_ , \new_[1551]_ ,
    \new_[1552]_ , \new_[1553]_ , \new_[1554]_ , \new_[1555]_ ,
    \new_[1556]_ , \new_[1557]_ , \new_[1558]_ , \new_[1559]_ ,
    \new_[1560]_ , \new_[1561]_ , \new_[1562]_ , \new_[1563]_ ,
    \new_[1564]_ , \new_[1565]_ , \new_[1566]_ , \new_[1567]_ ,
    \new_[1568]_ , \new_[1569]_ , \new_[1570]_ , \new_[1571]_ ,
    \new_[1572]_ , \new_[1573]_ , \new_[1574]_ , \new_[1575]_ ,
    \new_[1576]_ , \new_[1577]_ , \new_[1578]_ , \new_[1579]_ ,
    \new_[1580]_ , \new_[1581]_ , \new_[1583]_ , \new_[1584]_ ,
    \new_[1585]_ , \new_[1586]_ , \new_[1587]_ , \new_[1588]_ ,
    \new_[1589]_ , \new_[1590]_ , \new_[1592]_ , \new_[1593]_ ,
    \new_[1596]_ , \new_[1597]_ , \new_[1598]_ , \new_[1599]_ ,
    \new_[1600]_ , \new_[1601]_ , \new_[1602]_ , \new_[1603]_ ,
    \new_[1604]_ , \new_[1605]_ , \new_[1606]_ , \new_[1607]_ ,
    \new_[1608]_ , \new_[1609]_ , \new_[1610]_ , \new_[1611]_ ,
    \new_[1612]_ , \new_[1613]_ , \new_[1614]_ , \new_[1615]_ ,
    \new_[1616]_ , \new_[1617]_ , \new_[1618]_ , \new_[1619]_ ,
    \new_[1620]_ , \new_[1621]_ , \new_[1622]_ , \new_[1623]_ ,
    \new_[1624]_ , \new_[1625]_ , \new_[1626]_ , \new_[1627]_ ,
    \new_[1628]_ , \new_[1629]_ , \new_[1630]_ , \new_[1631]_ ,
    \new_[1632]_ , \new_[1633]_ , \new_[1634]_ , \new_[1635]_ ,
    \new_[1636]_ , \new_[1637]_ , \new_[1638]_ , \new_[1639]_ ,
    \new_[1640]_ , \new_[1641]_ , \new_[1642]_ , \new_[1643]_ ,
    \new_[1644]_ , \new_[1645]_ , \new_[1647]_ , \new_[1649]_ ,
    \new_[1650]_ , \new_[1651]_ , \new_[1652]_ , \new_[1653]_ ,
    \new_[1654]_ , \new_[1655]_ , \new_[1656]_ , \new_[1657]_ ,
    \new_[1658]_ , \new_[1659]_ , \new_[1660]_ , \new_[1661]_ ,
    \new_[1662]_ , \new_[1663]_ , \new_[1664]_ , \new_[1665]_ ,
    \new_[1666]_ , \new_[1667]_ , \new_[1668]_ , \new_[1669]_ ,
    \new_[1670]_ , \new_[1671]_ , \new_[1672]_ , \new_[1673]_ ,
    \new_[1674]_ , \new_[1675]_ , \new_[1676]_ , \new_[1677]_ ,
    \new_[1678]_ , \new_[1679]_ , \new_[1680]_ , \new_[1681]_ ,
    \new_[1682]_ , \new_[1683]_ , \new_[1684]_ , \new_[1685]_ ,
    \new_[1686]_ , \new_[1687]_ , \new_[1688]_ , \new_[1689]_ ,
    \new_[1690]_ , \new_[1691]_ , \new_[1692]_ , \new_[1693]_ ,
    \new_[1694]_ , \new_[1695]_ , \new_[1696]_ , \new_[1697]_ ,
    \new_[1698]_ , \new_[1699]_ , \new_[1700]_ , \new_[1701]_ ,
    \new_[1702]_ , \new_[1703]_ , \new_[1704]_ , \new_[1705]_ ,
    \new_[1706]_ , \new_[1707]_ , \new_[1708]_ , \new_[1709]_ ,
    \new_[1710]_ , \new_[1711]_ , \new_[1712]_ , \new_[1713]_ ,
    \new_[1714]_ , \new_[1715]_ , \new_[1716]_ , \new_[1717]_ ,
    \new_[1718]_ , \new_[1719]_ , \new_[1720]_ , \new_[1721]_ ,
    \new_[1722]_ , \new_[1723]_ , \new_[1724]_ , \new_[1725]_ ,
    \new_[1726]_ , \new_[1727]_ , \new_[1728]_ , \new_[1729]_ ,
    \new_[1730]_ , \new_[1731]_ , \new_[1732]_ , \new_[1733]_ ,
    \new_[1734]_ , \new_[1735]_ , \new_[1736]_ , \new_[1737]_ ,
    \new_[1738]_ , \new_[1753]_ , \new_[1754]_ , \new_[1755]_ ,
    \new_[1756]_ , \new_[1758]_ , \new_[1759]_ , \new_[1760]_ ,
    \new_[1761]_ , \new_[1762]_ , \new_[1763]_ , \new_[1764]_ ,
    \new_[1765]_ , \new_[1766]_ , \new_[1767]_ , \new_[1768]_ ,
    \new_[1769]_ , \new_[1770]_ , \new_[1771]_ , \new_[1772]_ ,
    \new_[1773]_ , \new_[1774]_ , \new_[1775]_ , \new_[1776]_ ,
    \new_[1777]_ , \new_[1778]_ , \new_[1779]_ , \new_[1780]_ ,
    \new_[1781]_ , \new_[1782]_ , \new_[1783]_ , \new_[1784]_ ,
    \new_[1785]_ , \new_[1786]_ , \new_[1787]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1791]_ , \new_[1793]_ ,
    \new_[1794]_ , \new_[1795]_ , \new_[1796]_ , \new_[1797]_ ,
    \new_[1798]_ , \new_[1799]_ , \new_[1800]_ , \new_[1801]_ ,
    \new_[1802]_ , \new_[1803]_ , \new_[1804]_ , \new_[1807]_ ,
    \new_[1808]_ , \new_[1836]_ , \new_[1842]_ , \new_[1851]_ ,
    \new_[1852]_ , \new_[1853]_ , \new_[1854]_ , \new_[1855]_ ,
    \new_[1856]_ , \new_[1857]_ , \new_[1858]_ , \new_[1859]_ ,
    \new_[1860]_ , \new_[1861]_ , \new_[1862]_ , \new_[1863]_ ,
    \new_[1864]_ , \new_[1865]_ , \new_[1866]_ , \new_[1867]_ ,
    \new_[1868]_ , \new_[1869]_ , \new_[1870]_ , \new_[1871]_ ,
    \new_[1872]_ , \new_[1873]_ , \new_[1874]_ , \new_[1875]_ ,
    \new_[1876]_ , \new_[1877]_ , \new_[1878]_ , \new_[1879]_ ,
    \new_[1880]_ , \new_[1881]_ , \new_[1882]_ , \new_[1883]_ ,
    \new_[1884]_ , \new_[1885]_ , \new_[1886]_ , \new_[1887]_ ,
    \new_[1888]_ , \new_[1889]_ , \new_[1890]_ , \new_[1891]_ ,
    \new_[1892]_ , \new_[1893]_ , \new_[1894]_ , \new_[1895]_ ,
    \new_[1896]_ , \new_[1897]_ , \new_[1898]_ , \new_[1899]_ ,
    \new_[1900]_ , \new_[1901]_ , \new_[1902]_ , \new_[1903]_ ,
    \new_[1904]_ , \new_[1905]_ , \new_[1906]_ , \new_[1907]_ ,
    \new_[1908]_ , \new_[1909]_ , \new_[1910]_ , \new_[1911]_ ,
    \new_[1912]_ , \new_[1915]_ , \new_[1924]_ , \new_[1931]_ ,
    \new_[1939]_ , \new_[1941]_ , \new_[1942]_ , \new_[1943]_ ,
    \new_[1944]_ , \new_[1945]_ , \new_[1946]_ , \new_[1947]_ ,
    \new_[1948]_ , \new_[1949]_ , \new_[1950]_ , \new_[1951]_ ,
    \new_[1952]_ , \new_[1953]_ , \new_[1954]_ , \new_[1955]_ ,
    \new_[1956]_ , \new_[1957]_ , \new_[1958]_ , \new_[1960]_ ,
    \new_[1961]_ , \new_[1962]_ , \new_[1963]_ , \new_[1964]_ ,
    \new_[1965]_ , \new_[1966]_ , \new_[1967]_ , \new_[1968]_ ,
    \new_[1969]_ , \new_[1970]_ , \new_[1971]_ , \new_[1972]_ ,
    \new_[1973]_ , \new_[1974]_ , \new_[1975]_ , \new_[1976]_ ,
    \new_[1977]_ , \new_[1983]_ , \new_[1984]_ , \new_[1995]_ ,
    \new_[1999]_ , \new_[2012]_ , \new_[2022]_ , \new_[2023]_ ,
    \new_[2024]_ , \new_[2025]_ , \new_[2028]_ , \new_[2029]_ ,
    \new_[2030]_ , \new_[2031]_ , \new_[2032]_ , \new_[2033]_ ,
    \new_[2034]_ , \new_[2035]_ , \new_[2036]_ , \new_[2037]_ ,
    \new_[2038]_ , \new_[2060]_ , \new_[2061]_ , \new_[2062]_ ,
    \new_[2063]_ , \new_[2064]_ , \new_[2065]_ , \new_[2066]_ ,
    \new_[2067]_ , \new_[2068]_ , \new_[2069]_ , \new_[2070]_ ,
    \new_[2071]_ , \new_[2072]_ , \new_[2073]_ , \new_[2074]_ ,
    \new_[2075]_ , \new_[2076]_ , \new_[2077]_ , \new_[2078]_ ,
    \new_[2079]_ , \new_[2080]_ , \new_[2081]_ , \new_[2082]_ ,
    \new_[2083]_ , \new_[2084]_ , \new_[2085]_ , \new_[2086]_ ,
    \new_[2087]_ , \new_[2088]_ , \new_[2089]_ , \new_[2090]_ ,
    \new_[2091]_ , \new_[2092]_ , \new_[2093]_ , \new_[2094]_ ,
    \new_[2095]_ , \new_[2096]_ , \new_[2097]_ , \new_[2098]_ ,
    \new_[2099]_ , \new_[2100]_ , \new_[2101]_ , \new_[2102]_ ,
    \new_[2103]_ , \new_[2104]_ , \new_[2105]_ , \new_[2106]_ ,
    \new_[2107]_ , \new_[2108]_ , \new_[2109]_ , \new_[2110]_ ,
    \new_[2111]_ , \new_[2112]_ , \new_[2113]_ , \new_[2114]_ ,
    \new_[2115]_ , \new_[2116]_ , \new_[2117]_ , \new_[2118]_ ,
    \new_[2119]_ , \new_[2120]_ , \new_[2121]_ , \new_[2122]_ ,
    \new_[2123]_ , \new_[2124]_ , \new_[2125]_ , \new_[2126]_ ,
    \new_[2127]_ , \new_[2128]_ , \new_[2129]_ , \new_[2130]_ ,
    \new_[2131]_ , \new_[2132]_ , \new_[2133]_ , \new_[2134]_ ,
    \new_[2135]_ , \new_[2136]_ , \new_[2137]_ , \new_[2138]_ ,
    \new_[2139]_ , \new_[2140]_ , \new_[2141]_ , \new_[2155]_ ,
    \new_[2157]_ , \new_[2158]_ , \new_[2159]_ , \new_[2160]_ ,
    \new_[2161]_ , \new_[2162]_ , \new_[2163]_ , \new_[2164]_ ,
    \new_[2165]_ , \new_[2166]_ , \new_[2167]_ , \new_[2168]_ ,
    \new_[2171]_ , \new_[2172]_ , \new_[2173]_ , \new_[2174]_ ,
    \new_[2175]_ , \new_[2176]_ , \new_[2177]_ , \new_[2178]_ ,
    \new_[2179]_ , \new_[2180]_ , \new_[2181]_ , \new_[2182]_ ,
    \new_[2183]_ , \new_[2184]_ , \new_[2185]_ , \new_[2186]_ ,
    \new_[2187]_ , \new_[2188]_ , \new_[2189]_ , \new_[2190]_ ,
    \new_[2191]_ , \new_[2192]_ , \new_[2193]_ , \new_[2194]_ ,
    \new_[2195]_ , \new_[2196]_ , \new_[2197]_ , \new_[2198]_ ,
    \new_[2199]_ , \new_[2200]_ , \new_[2201]_ , \new_[2202]_ ,
    \new_[2203]_ , \new_[2204]_ , \new_[2205]_ , \new_[2206]_ ,
    \new_[2207]_ , \new_[2208]_ , \new_[2209]_ , \new_[2210]_ ,
    \new_[2211]_ , \new_[2212]_ , \new_[2213]_ , \new_[2214]_ ,
    \new_[2215]_ , \new_[2216]_ , \new_[2217]_ , \new_[2218]_ ,
    \new_[2219]_ , \new_[2220]_ , \new_[2221]_ , \new_[2222]_ ,
    \new_[2223]_ , \new_[2224]_ , \new_[2225]_ , \new_[2226]_ ,
    \new_[2227]_ , \new_[2238]_ , \new_[2239]_ , \new_[2240]_ ,
    \new_[2241]_ , \new_[2242]_ , \new_[2243]_ , \new_[2244]_ ,
    \new_[2245]_ , \new_[2246]_ , \new_[2247]_ , \new_[2248]_ ,
    \new_[2249]_ , \new_[2250]_ , \new_[2251]_ , \new_[2266]_ ,
    \new_[2267]_ , \new_[2268]_ , \new_[2269]_ , \new_[2270]_ ,
    \new_[2271]_ , \new_[2272]_ , \new_[2273]_ , \new_[2274]_ ,
    \new_[2275]_ , \new_[2276]_ , \new_[2277]_ , \new_[2278]_ ,
    \new_[2279]_ , \new_[2280]_ , \new_[2281]_ , \new_[2282]_ ,
    \new_[2283]_ , \new_[2284]_ , \new_[2285]_ , \new_[2286]_ ,
    \new_[2287]_ , \new_[2288]_ , \new_[2289]_ , \new_[2290]_ ,
    \new_[2291]_ , \new_[2292]_ , \new_[2293]_ , \new_[2294]_ ,
    \new_[2295]_ , \new_[2296]_ , \new_[2297]_ , \new_[2298]_ ,
    \new_[2299]_ , \new_[2300]_ , \new_[2301]_ , \new_[2302]_ ,
    \new_[2303]_ , \new_[2304]_ , \new_[2305]_ , \new_[2306]_ ,
    \new_[2307]_ , \new_[2308]_ , \new_[2309]_ , \new_[2310]_ ,
    \new_[2311]_ , \new_[2312]_ , \new_[2313]_ , \new_[2314]_ ,
    \new_[2315]_ , \new_[2316]_ , \new_[2317]_ , \new_[2318]_ ,
    \new_[2319]_ , \new_[2320]_ , \new_[2321]_ , \new_[2322]_ ,
    \new_[2323]_ , \new_[2324]_ , \new_[2325]_ , \new_[2326]_ ,
    \new_[2327]_ , \new_[2328]_ , \new_[2329]_ , \new_[2330]_ ,
    \new_[2331]_ , \new_[2332]_ , \new_[2333]_ , \new_[2334]_ ,
    \new_[2347]_ , \new_[2348]_ , \new_[2353]_ , \new_[2354]_ ,
    \new_[2355]_ , \new_[2356]_ , \new_[2357]_ , \new_[2358]_ ,
    \new_[2359]_ , \new_[2360]_ , \new_[2361]_ , \new_[2362]_ ,
    \new_[2363]_ , \new_[2364]_ , \new_[2365]_ , \new_[2366]_ ,
    \new_[2367]_ , \new_[2368]_ , \new_[2369]_ , \new_[2370]_ ,
    \new_[2371]_ , \new_[2372]_ , \new_[2373]_ , \new_[2374]_ ,
    \new_[2375]_ , \new_[2376]_ , \new_[2377]_ , \new_[2378]_ ,
    \new_[2379]_ , \new_[2380]_ , \new_[2381]_ , \new_[2382]_ ,
    \new_[2383]_ , \new_[2384]_ , \new_[2385]_ , \new_[2386]_ ,
    \new_[2387]_ , \new_[2389]_ , \new_[2390]_ , \new_[2391]_ ,
    \new_[2392]_ , \new_[2393]_ , \new_[2394]_ , \new_[2395]_ ,
    \new_[2396]_ , \new_[2397]_ , \new_[2399]_ , \new_[2400]_ ,
    \new_[2401]_ , \new_[2402]_ , \new_[2403]_ , \new_[2404]_ ,
    \new_[2405]_ , \new_[2406]_ , \new_[2407]_ , \new_[2408]_ ,
    \new_[2409]_ , \new_[2410]_ , \new_[2411]_ , \new_[2412]_ ,
    \new_[2413]_ , \new_[2414]_ , \new_[2415]_ , \new_[2416]_ ,
    \new_[2417]_ , \new_[2418]_ , \new_[2420]_ , \new_[2421]_ ,
    \new_[2422]_ , \new_[2423]_ , \new_[2424]_ , \new_[2425]_ ,
    \new_[2426]_ , \new_[2427]_ , \new_[2428]_ , \new_[2429]_ ,
    \new_[2430]_ , \new_[2431]_ , \new_[2432]_ , \new_[2433]_ ,
    \new_[2434]_ , \new_[2435]_ , \new_[2436]_ , \new_[2438]_ ,
    \new_[2439]_ , \new_[2440]_ , \new_[2441]_ , \new_[2442]_ ,
    \new_[2443]_ , \new_[2444]_ , \new_[2445]_ , \new_[2446]_ ,
    \new_[2447]_ , \new_[2448]_ , \new_[2449]_ , \new_[2450]_ ,
    \new_[2451]_ , \new_[2452]_ , \new_[2453]_ , \new_[2454]_ ,
    \new_[2455]_ , \new_[2456]_ , \new_[2457]_ , \new_[2458]_ ,
    \new_[2459]_ , \new_[2460]_ , \new_[2461]_ , \new_[2462]_ ,
    \new_[2463]_ , \new_[2464]_ , \new_[2465]_ , \new_[2466]_ ,
    \new_[2467]_ , \new_[2468]_ , \new_[2469]_ , \new_[2470]_ ,
    \new_[2471]_ , \new_[2472]_ , \new_[2473]_ , \new_[2474]_ ,
    \new_[2475]_ , \new_[2476]_ , \new_[2477]_ , \new_[2478]_ ,
    \new_[2479]_ , \new_[2480]_ , \new_[2481]_ , \new_[2482]_ ,
    \new_[2483]_ , \new_[2484]_ , \new_[2485]_ , \new_[2486]_ ,
    \new_[2487]_ , \new_[2488]_ , \new_[2489]_ , \new_[2490]_ ,
    \new_[2491]_ , \new_[2492]_ , \new_[2493]_ , \new_[2494]_ ,
    \new_[2495]_ , \new_[2496]_ , \new_[2497]_ , \new_[2498]_ ,
    \new_[2499]_ , \new_[2500]_ , \new_[2501]_ , \new_[2502]_ ,
    \new_[2503]_ , \new_[2504]_ , \new_[2505]_ , \new_[2506]_ ,
    \new_[2507]_ , \new_[2508]_ , \new_[2509]_ , \new_[2510]_ ,
    \new_[2511]_ , \new_[2512]_ , \new_[2513]_ , \new_[2514]_ ,
    \new_[2515]_ , \new_[2516]_ , \new_[2517]_ , \new_[2518]_ ,
    \new_[2519]_ , \new_[2520]_ , \new_[2521]_ , \new_[2522]_ ,
    \new_[2523]_ , \new_[2524]_ , \new_[2525]_ , \new_[2526]_ ,
    \new_[2527]_ , \new_[2528]_ , \new_[2529]_ , \new_[2530]_ ,
    \new_[2531]_ , \new_[2532]_ , \new_[2533]_ , \new_[2534]_ ,
    \new_[2535]_ , \new_[2536]_ , \new_[2537]_ , \new_[2538]_ ,
    \new_[2539]_ , \new_[2540]_ , \new_[2541]_ , \new_[2542]_ ,
    \new_[2543]_ , \new_[2544]_ , \new_[2545]_ , \new_[2546]_ ,
    \new_[2547]_ , \new_[2548]_ , \new_[2549]_ , \new_[2550]_ ,
    \new_[2551]_ , \new_[2552]_ , \new_[2553]_ , \new_[2554]_ ,
    \new_[2555]_ , \new_[2556]_ , \new_[2557]_ , \new_[2558]_ ,
    \new_[2559]_ , \new_[2560]_ , \new_[2561]_ , \new_[2562]_ ,
    \new_[2563]_ , \new_[2564]_ , \new_[2565]_ , \new_[2566]_ ,
    \new_[2567]_ , \new_[2568]_ , \new_[2569]_ , \new_[2571]_ ,
    \new_[2572]_ , \new_[2573]_ , \new_[2574]_ , \new_[2575]_ ,
    \new_[2576]_ , \new_[2577]_ , \new_[2578]_ , \new_[2579]_ ,
    \new_[2580]_ , \new_[2581]_ , \new_[2582]_ , \new_[2583]_ ,
    \new_[2584]_ , \new_[2585]_ , \new_[2586]_ , \new_[2587]_ ,
    \new_[2588]_ , \new_[2589]_ , \new_[2590]_ , \new_[2591]_ ,
    \new_[2592]_ , \new_[2593]_ , \new_[2594]_ , \new_[2595]_ ,
    \new_[2596]_ , \new_[2597]_ , \new_[2598]_ , \new_[2599]_ ,
    \new_[2600]_ , \new_[2601]_ , \new_[2602]_ , \new_[2603]_ ,
    \new_[2604]_ , \new_[2605]_ , \new_[2606]_ , \new_[2607]_ ,
    \new_[2608]_ , \new_[2609]_ , \new_[2610]_ , \new_[2611]_ ,
    \new_[2612]_ , \new_[2613]_ , \new_[2614]_ , \new_[2615]_ ,
    \new_[2616]_ , \new_[2617]_ , \new_[2618]_ , \new_[2619]_ ,
    \new_[2620]_ , \new_[2621]_ , \new_[2622]_ , \new_[2623]_ ,
    \new_[2624]_ , \new_[2625]_ , \new_[2626]_ , \new_[2627]_ ,
    \new_[2628]_ , \new_[2629]_ , \new_[2630]_ , \new_[2631]_ ,
    \new_[2632]_ , \new_[2633]_ , \new_[2634]_ , \new_[2635]_ ,
    \new_[2636]_ , \new_[2637]_ , \new_[2638]_ , \new_[2639]_ ,
    \new_[2640]_ , \new_[2641]_ , \new_[2642]_ , \new_[2643]_ ,
    \new_[2644]_ , \new_[2645]_ , \new_[2646]_ , \new_[2647]_ ,
    \new_[2648]_ , \new_[2649]_ , \new_[2650]_ , \new_[2651]_ ,
    \new_[2652]_ , \new_[2653]_ , \new_[2654]_ , \new_[2655]_ ,
    \new_[2656]_ , \new_[2657]_ , \new_[2658]_ , \new_[2659]_ ,
    \new_[2661]_ , \new_[2662]_ , \new_[2663]_ , \new_[2664]_ ,
    \new_[2665]_ , \new_[2666]_ , \new_[2667]_ , \new_[2668]_ ,
    \new_[2669]_ , \new_[2670]_ , \new_[2671]_ , \new_[2672]_ ,
    \new_[2673]_ , \new_[2674]_ , \new_[2675]_ , \new_[2676]_ ,
    \new_[2677]_ , \new_[2678]_ , \new_[2679]_ , \new_[2680]_ ,
    \new_[2681]_ , \new_[2683]_ , \new_[2692]_ , \new_[2694]_ ,
    \new_[2697]_ , \new_[2698]_ , \new_[2699]_ , \new_[2700]_ ,
    \new_[2701]_ , \new_[2702]_ , \new_[2703]_ , \new_[2704]_ ,
    \new_[2705]_ , \new_[2706]_ , \new_[2707]_ , \new_[2708]_ ,
    \new_[2709]_ , \new_[2710]_ , \new_[2711]_ , \new_[2712]_ ,
    \new_[2713]_ , \new_[2714]_ , \new_[2715]_ , \new_[2716]_ ,
    \new_[2718]_ , \new_[2724]_ , \new_[2725]_ , \new_[2726]_ ,
    \new_[2727]_ , \new_[2728]_ , \new_[2729]_ , \new_[2730]_ ,
    \new_[2741]_ , \new_[2742]_ , \new_[2745]_ , \new_[2746]_ ,
    \new_[2747]_ , \new_[2748]_ , \new_[2749]_ , \new_[2750]_ ,
    \new_[2751]_ , \new_[2754]_ , \new_[2755]_ , \new_[2756]_ ,
    \new_[2757]_ , \new_[2758]_ , \new_[2759]_ , \new_[2760]_ ,
    \new_[2761]_ , \new_[2762]_ , \new_[2763]_ , \new_[2764]_ ,
    \new_[2765]_ , \new_[2766]_ , \new_[2767]_ , \new_[2768]_ ,
    \new_[2769]_ , \new_[2770]_ , \new_[2771]_ , \new_[2772]_ ,
    \new_[2773]_ , \new_[2774]_ , \new_[2775]_ , \new_[2776]_ ,
    \new_[2777]_ , \new_[2778]_ , \new_[2779]_ , \new_[2780]_ ,
    \new_[2781]_ , \new_[2782]_ , \new_[2783]_ , \new_[2784]_ ,
    \new_[2785]_ , \new_[2786]_ , \new_[2787]_ , \new_[2788]_ ,
    \new_[2789]_ , \new_[2790]_ , \new_[2791]_ , \new_[2792]_ ,
    \new_[2793]_ , \new_[2794]_ , \new_[2795]_ , \new_[2796]_ ,
    \new_[2797]_ , \new_[2798]_ , \new_[2799]_ , \new_[2800]_ ,
    \new_[2801]_ , \new_[2802]_ , \new_[2803]_ , \new_[2804]_ ,
    \new_[2805]_ , \new_[2806]_ , \new_[2807]_ , \new_[2808]_ ,
    \new_[2809]_ , \new_[2810]_ , \new_[2811]_ , \new_[2812]_ ,
    \new_[2813]_ , \new_[2814]_ , \new_[2815]_ , \new_[2816]_ ,
    \new_[2817]_ , \new_[2818]_ , \new_[2819]_ , \new_[2820]_ ,
    \new_[2821]_ , \new_[2822]_ , \new_[2823]_ , \new_[2824]_ ,
    \new_[2825]_ , \new_[2826]_ , \new_[2827]_ , \new_[2828]_ ,
    \new_[2829]_ , \new_[2830]_ , \new_[2831]_ , \new_[2832]_ ,
    \new_[2833]_ , \new_[2834]_ , \new_[2835]_ , \new_[2836]_ ,
    \new_[2837]_ , \new_[2838]_ , \new_[2839]_ , \new_[2840]_ ,
    \new_[2841]_ , \new_[2842]_ , \new_[2846]_ , \new_[2847]_ ,
    \new_[2848]_ , \new_[2849]_ , \new_[2850]_ , \new_[2851]_ ,
    \new_[2852]_ , \new_[2853]_ , \new_[2854]_ , \new_[2855]_ ,
    \new_[2856]_ , \new_[2857]_ , \new_[2858]_ , \new_[2859]_ ,
    \new_[2860]_ , \new_[2861]_ , \new_[2862]_ , \new_[2863]_ ,
    \new_[2864]_ , \new_[2865]_ , \new_[2866]_ , \new_[2867]_ ,
    \new_[2868]_ , \new_[2869]_ , \new_[2870]_ , \new_[2871]_ ,
    \new_[2872]_ , \new_[2873]_ , \new_[2874]_ , \new_[2875]_ ,
    \new_[2876]_ , \new_[2877]_ , \new_[2878]_ , \new_[2879]_ ,
    \new_[2880]_ , \new_[2881]_ , \new_[2882]_ , \new_[2883]_ ,
    \new_[2884]_ , \new_[2885]_ , \new_[2886]_ , \new_[2887]_ ,
    \new_[2888]_ , \new_[2889]_ , \new_[2890]_ , \new_[2891]_ ,
    \new_[2892]_ , \new_[2893]_ , \new_[2894]_ , \new_[2895]_ ,
    \new_[2896]_ , \new_[2897]_ , \new_[2898]_ , \new_[2899]_ ,
    \new_[2900]_ , \new_[2901]_ , \new_[2902]_ , \new_[2903]_ ,
    \new_[2904]_ , \new_[2905]_ , \new_[2906]_ , \new_[2907]_ ,
    \new_[2908]_ , \new_[2909]_ , \new_[2910]_ , \new_[2911]_ ,
    \new_[2912]_ , \new_[2913]_ , \new_[2914]_ , \new_[2916]_ ,
    \new_[2917]_ , \new_[2918]_ , \new_[2919]_ , \new_[2920]_ ,
    \new_[2921]_ , \new_[2922]_ , \new_[2923]_ , \new_[2924]_ ,
    \new_[2925]_ , \new_[2926]_ , \new_[2927]_ , \new_[2928]_ ,
    \new_[2929]_ , \new_[2930]_ , \new_[2931]_ , \new_[2932]_ ,
    \new_[2933]_ , \new_[2936]_ , \new_[2937]_ , \new_[2938]_ ,
    \new_[2939]_ , \new_[2940]_ , \new_[2944]_ , \new_[2945]_ ,
    \new_[2946]_ , \new_[2947]_ , \new_[2948]_ , \new_[2949]_ ,
    \new_[2950]_ , \new_[2951]_ , \new_[2952]_ , \new_[2953]_ ,
    \new_[2955]_ , \new_[2956]_ , \new_[2957]_ , \new_[2959]_ ,
    \new_[2960]_ , \new_[2961]_ , \new_[2962]_ , \new_[2963]_ ,
    \new_[2964]_ , \new_[2965]_ , \new_[2966]_ , \new_[2967]_ ,
    \new_[2968]_ , \new_[2969]_ , \new_[2970]_ , \new_[2971]_ ,
    \new_[2972]_ , \new_[2973]_ , \new_[2974]_ , \new_[2975]_ ,
    \new_[2976]_ , \new_[2977]_ , \new_[2978]_ , \new_[2979]_ ,
    \new_[2980]_ , \new_[2981]_ , \new_[2982]_ , \new_[2983]_ ,
    \new_[2984]_ , \new_[2985]_ , \new_[2986]_ , \new_[2987]_ ,
    \new_[2988]_ , \new_[2989]_ , \new_[2990]_ , \new_[2991]_ ,
    \new_[2992]_ , \new_[2993]_ , \new_[2994]_ , \new_[2995]_ ,
    \new_[2996]_ , \new_[2997]_ , \new_[2998]_ , \new_[2999]_ ,
    \new_[3000]_ , \new_[3001]_ , \new_[3002]_ , \new_[3003]_ ,
    \new_[3004]_ , \new_[3005]_ , \new_[3006]_ , \new_[3007]_ ,
    \new_[3008]_ , \new_[3009]_ , \new_[3010]_ , \new_[3011]_ ,
    \new_[3012]_ , \new_[3015]_ , \new_[3016]_ , \new_[3017]_ ,
    \new_[3018]_ , \new_[3019]_ , \new_[3020]_ , \new_[3021]_ ,
    \new_[3022]_ , \new_[3023]_ , \new_[3024]_ , \new_[3025]_ ,
    \new_[3026]_ , \new_[3027]_ , \new_[3028]_ , \new_[3029]_ ,
    \new_[3030]_ , \new_[3031]_ , \new_[3032]_ , \new_[3033]_ ,
    \new_[3036]_ , \new_[3038]_ , \new_[3039]_ , \new_[3041]_ ,
    \new_[3042]_ , \new_[3047]_ , \new_[3049]_ , \new_[3050]_ ,
    \new_[3051]_ , \new_[3052]_ , \new_[3053]_ , \new_[3054]_ ,
    \new_[3055]_ , \new_[3056]_ , \new_[3057]_ , \new_[3066]_ ,
    \new_[3067]_ , \new_[3068]_ , \new_[3069]_ , \new_[3070]_ ,
    \new_[3071]_ , \new_[3072]_ , \new_[3073]_ , \new_[3074]_ ,
    \new_[3075]_ , \new_[3076]_ , \new_[3077]_ , \new_[3078]_ ,
    \new_[3079]_ , \new_[3080]_ , \new_[3081]_ , \new_[3082]_ ,
    \new_[3083]_ , \new_[3084]_ , \new_[3085]_ , \new_[3086]_ ,
    \new_[3087]_ , \new_[3088]_ , \new_[3089]_ , \new_[3090]_ ,
    \new_[3091]_ , \new_[3092]_ , \new_[3093]_ , \new_[3094]_ ,
    \new_[3095]_ , \new_[3098]_ , \new_[3099]_ , \new_[3100]_ ,
    \new_[3101]_ , \new_[3102]_ , \new_[3103]_ , \new_[3105]_ ,
    \new_[3128]_ , \new_[3129]_ , \new_[3130]_ , \new_[3131]_ ,
    \new_[3132]_ , \new_[3156]_ , \new_[3157]_ , \new_[3158]_ ,
    \new_[3159]_ , \new_[3160]_ , \new_[3161]_ , \new_[3162]_ ,
    \new_[3163]_ , \new_[3164]_ , \new_[3165]_ , \new_[3166]_ ,
    \new_[3167]_ , \new_[3168]_ , \new_[3169]_ , \new_[3170]_ ,
    \new_[3171]_ , \new_[3172]_ , \new_[3173]_ , \new_[3174]_ ,
    \new_[3175]_ , \new_[3176]_ , \new_[3177]_ , \new_[3178]_ ,
    \new_[3179]_ , \new_[3180]_ , \new_[3181]_ , \new_[3182]_ ,
    \new_[3183]_ , \new_[3184]_ , \new_[3185]_ , \new_[3186]_ ,
    \new_[3187]_ , \new_[3188]_ , \new_[3189]_ , \new_[3190]_ ,
    \new_[3191]_ , \new_[3192]_ , \new_[3193]_ , \new_[3194]_ ,
    \new_[3195]_ , \new_[3197]_ , \new_[3198]_ , \new_[3199]_ ,
    \new_[3201]_ , \new_[3202]_ , \new_[3203]_ , \new_[3204]_ ,
    \new_[3205]_ , \new_[3206]_ , \new_[3207]_ , \new_[3208]_ ,
    \new_[3209]_ , \new_[3210]_ , \new_[3211]_ , \new_[3212]_ ,
    \new_[3213]_ , \new_[3214]_ , \new_[3215]_ , \new_[3216]_ ,
    \new_[3217]_ , \new_[3218]_ , \new_[3219]_ , \new_[3220]_ ,
    \new_[3221]_ , \new_[3222]_ , \new_[3223]_ , \new_[3224]_ ,
    \new_[3225]_ , \new_[3226]_ , \new_[3227]_ , \new_[3228]_ ,
    \new_[3230]_ , \new_[3231]_ , \new_[3232]_ , \new_[3233]_ ,
    \new_[3234]_ , \new_[3235]_ , \new_[3236]_ , \new_[3237]_ ,
    \new_[3238]_ , \new_[3239]_ , \new_[3240]_ , \new_[3241]_ ,
    \new_[3242]_ , \new_[3243]_ , \new_[3244]_ , \new_[3245]_ ,
    \new_[3246]_ , \new_[3247]_ , \new_[3248]_ , \new_[3249]_ ,
    \new_[3250]_ , \new_[3251]_ , \new_[3252]_ , \new_[3253]_ ,
    \new_[3254]_ , \new_[3255]_ , \new_[3256]_ , \new_[3257]_ ,
    \new_[3259]_ , \new_[3261]_ , \new_[3262]_ , \new_[3263]_ ,
    \new_[3264]_ , \new_[3265]_ , \new_[3266]_ , \new_[3267]_ ,
    \new_[3268]_ , \new_[3269]_ , \new_[3270]_ , \new_[3271]_ ,
    \new_[3272]_ , \new_[3273]_ , \new_[3274]_ , \new_[3275]_ ,
    \new_[3276]_ , \new_[3278]_ , \new_[3279]_ , \new_[3280]_ ,
    \new_[3282]_ , \new_[3284]_ , \new_[3285]_ , \new_[3286]_ ,
    \new_[3287]_ , \new_[3288]_ , \new_[3290]_ , \new_[3291]_ ,
    \new_[3292]_ , \new_[3293]_ , \new_[3294]_ , \new_[3295]_ ,
    \new_[3296]_ , \new_[3297]_ , \new_[3298]_ , \new_[3299]_ ,
    \new_[3300]_ , \new_[3301]_ , \new_[3302]_ , \new_[3303]_ ,
    \new_[3304]_ , \new_[3305]_ , \new_[3306]_ , \new_[3307]_ ,
    \new_[3308]_ , \new_[3309]_ , \new_[3311]_ , \new_[3313]_ ,
    \new_[3315]_ , \new_[3316]_ , \new_[3317]_ , \new_[3318]_ ,
    \new_[3320]_ , \new_[3321]_ , \new_[3322]_ , \new_[3323]_ ,
    \new_[3324]_ , \new_[3325]_ , \new_[3327]_ , \new_[3328]_ ,
    \new_[3329]_ , \new_[3330]_ , \new_[3331]_ , \new_[3332]_ ,
    \new_[3333]_ , \new_[3334]_ , \new_[3338]_ , \new_[3339]_ ,
    \new_[3340]_ , \new_[3343]_ , \new_[3344]_ , \new_[3345]_ ,
    \new_[3346]_ , \new_[3347]_ , \new_[3348]_ , \new_[3349]_ ,
    \new_[3350]_ , \new_[3354]_ , \new_[3355]_ , \new_[3356]_ ,
    \new_[3357]_ , \new_[3358]_ , \new_[3359]_ , \new_[3360]_ ,
    \new_[3361]_ , \new_[3362]_ , \new_[3363]_ , \new_[3364]_ ,
    \new_[3365]_ , \new_[3366]_ , \new_[3367]_ , \new_[3398]_ ,
    \new_[3401]_ , \new_[3412]_ , \new_[3413]_ , \new_[3414]_ ,
    \new_[3417]_ , \new_[3420]_ , \new_[3421]_ , \new_[3426]_ ,
    \new_[3427]_ , \new_[3428]_ , \new_[3429]_ , \new_[3430]_ ,
    \new_[3431]_ , \new_[3432]_ , \new_[3433]_ , \new_[3434]_ ,
    \new_[3436]_ , \new_[3437]_ , \new_[3438]_ , \new_[3439]_ ,
    \new_[3440]_ , \new_[3441]_ , \new_[3442]_ , \new_[3443]_ ,
    \new_[3444]_ , \new_[3445]_ , \new_[3446]_ , \new_[3447]_ ,
    \new_[3448]_ , \new_[3449]_ , \new_[3450]_ , \new_[3451]_ ,
    \new_[3452]_ , \new_[3453]_ , \new_[3454]_ , \new_[3455]_ ,
    \new_[3456]_ , \new_[3457]_ , \new_[3458]_ , \new_[3459]_ ,
    \new_[3460]_ , \new_[3461]_ , \new_[3462]_ , \new_[3463]_ ,
    \new_[3465]_ , \new_[3467]_ , \new_[3468]_ , \new_[3470]_ ,
    \new_[3471]_ , \new_[3472]_ , \new_[3473]_ , \new_[3475]_ ,
    \new_[3476]_ , \new_[3478]_ , \new_[3484]_ , \new_[3497]_ ,
    \new_[3502]_ , \new_[3503]_ , \new_[3504]_ , \new_[3505]_ ,
    \new_[3508]_ , \new_[3510]_ , \new_[3511]_ , \new_[3512]_ ,
    \new_[3513]_ , \new_[3515]_ , \new_[3516]_ , \new_[3517]_ ,
    \new_[3518]_ , \new_[3519]_ , \new_[3520]_ , \new_[3521]_ ,
    \new_[3522]_ , \new_[3523]_ , \new_[3524]_ , \new_[3525]_ ,
    \new_[3526]_ , \new_[3527]_ , \new_[3528]_ , \new_[3529]_ ,
    \new_[3534]_ , \new_[3535]_ , \new_[3536]_ , \new_[3537]_ ,
    \new_[3538]_ , \new_[3539]_ , \new_[3540]_ , \new_[3541]_ ,
    \new_[3542]_ , \new_[3543]_ , \new_[3544]_ , \new_[3545]_ ,
    \new_[3546]_ , \new_[3547]_ , \new_[3548]_ , \new_[3549]_ ,
    \new_[3550]_ , \new_[3551]_ , \new_[3552]_ , \new_[3553]_ ,
    \new_[3554]_ , \new_[3555]_ , \new_[3556]_ , \new_[3557]_ ,
    \new_[3558]_ , \new_[3559]_ , \new_[3560]_ , \new_[3561]_ ,
    \new_[3562]_ , \new_[3563]_ , \new_[3564]_ , \new_[3565]_ ,
    \new_[3566]_ , \new_[3567]_ , \new_[3568]_ , \new_[3569]_ ,
    \new_[3570]_ , \new_[3571]_ , \new_[3572]_ , \new_[3573]_ ,
    \new_[3574]_ , \new_[3575]_ , \new_[3576]_ , \new_[3577]_ ,
    \new_[3578]_ , \new_[3579]_ , \new_[3580]_ , \new_[3581]_ ,
    \new_[3582]_ , \new_[3583]_ , \new_[3584]_ , \new_[3585]_ ,
    \new_[3586]_ , \new_[3588]_ , \new_[3589]_ , \new_[3590]_ ,
    \new_[3591]_ , \new_[3592]_ , \new_[3593]_ , \new_[3594]_ ,
    \new_[3595]_ , \new_[3596]_ , \new_[3597]_ , \new_[3598]_ ,
    \new_[3599]_ , \new_[3600]_ , \new_[3601]_ , \new_[3602]_ ,
    \new_[3603]_ , \new_[3604]_ , \new_[3605]_ , \new_[3606]_ ,
    \new_[3607]_ , \new_[3608]_ , \new_[3609]_ , \new_[3610]_ ,
    \new_[3611]_ , \new_[3612]_ , \new_[3613]_ , \new_[3614]_ ,
    \new_[3615]_ , \new_[3616]_ , \new_[3617]_ , \new_[3618]_ ,
    \new_[3619]_ , \new_[3620]_ , \new_[3621]_ , \new_[3622]_ ,
    \new_[3624]_ , \new_[3625]_ , \new_[3626]_ , \new_[3627]_ ,
    \new_[3628]_ , \new_[3629]_ , \new_[3630]_ , \new_[3631]_ ,
    \new_[3632]_ , \new_[3633]_ , \new_[3634]_ , \new_[3635]_ ,
    \new_[3636]_ , \new_[3637]_ , \new_[3638]_ , \new_[3639]_ ,
    \new_[3640]_ , \new_[3641]_ , \new_[3642]_ , \new_[3643]_ ,
    \new_[3644]_ , \new_[3645]_ , \new_[3646]_ , \new_[3647]_ ,
    \new_[3648]_ , \new_[3649]_ , \new_[3650]_ , \new_[3651]_ ,
    \new_[3652]_ , \new_[3653]_ , \new_[3654]_ , \new_[3655]_ ,
    \new_[3656]_ , \new_[3657]_ , \new_[3658]_ , \new_[3659]_ ,
    \new_[3660]_ , \new_[3661]_ , \new_[3662]_ , \new_[3663]_ ,
    \new_[3664]_ , \new_[3665]_ , \new_[3666]_ , \new_[3667]_ ,
    \new_[3668]_ , \new_[3669]_ , \new_[3670]_ , \new_[3671]_ ,
    \new_[3672]_ , \new_[3678]_ , \new_[3682]_ , \new_[3690]_ ,
    \new_[3704]_ , \new_[3705]_ , \new_[3706]_ , \new_[3707]_ ,
    \new_[3709]_ , \new_[3710]_ , \new_[3711]_ , \new_[3712]_ ,
    \new_[3713]_ , \new_[3714]_ , \new_[3715]_ , \new_[3716]_ ,
    \new_[3717]_ , \new_[3718]_ , \new_[3719]_ , \new_[3722]_ ,
    \new_[3723]_ , \new_[3724]_ , \new_[3725]_ , \new_[3726]_ ,
    \new_[3727]_ , \new_[3728]_ , \new_[3729]_ , \new_[3730]_ ,
    \new_[3731]_ , \new_[3732]_ , \new_[3733]_ , \new_[3734]_ ,
    \new_[3735]_ , \new_[3736]_ , \new_[3737]_ , \new_[3738]_ ,
    \new_[3739]_ , \new_[3740]_ , \new_[3741]_ , \new_[3742]_ ,
    \new_[3743]_ , \new_[3744]_ , \new_[3745]_ , \new_[3746]_ ,
    \new_[3747]_ , \new_[3748]_ , \new_[3749]_ , \new_[3750]_ ,
    \new_[3751]_ , \new_[3752]_ , \new_[3753]_ , \new_[3754]_ ,
    \new_[3756]_ , \new_[3761]_ , \new_[3763]_ , \new_[3765]_ ,
    \new_[3768]_ , \new_[3770]_ , \new_[3771]_ , \new_[3772]_ ,
    \new_[3773]_ , \new_[3774]_ , \new_[3775]_ , \new_[3776]_ ,
    \new_[3777]_ , \new_[3779]_ , \new_[3781]_ , \new_[3784]_ ,
    \new_[3786]_ , \new_[3787]_ , \new_[3788]_ , \new_[3789]_ ,
    \new_[3790]_ , \new_[3791]_ , \new_[3792]_ , \new_[3793]_ ,
    \new_[3794]_ , \new_[3796]_ , \new_[3797]_ , \new_[3798]_ ,
    \new_[3799]_ , \new_[3803]_ , \new_[3804]_ , \new_[3805]_ ,
    \new_[3806]_ , \new_[3807]_ , \new_[3808]_ , \new_[3810]_ ,
    \new_[3812]_ , \new_[3814]_ , \new_[3817]_ , \new_[3819]_ ,
    \new_[3820]_ , \new_[3822]_ , \new_[3823]_ , \new_[3824]_ ,
    \new_[3825]_ , \new_[3826]_ , \new_[3827]_ , \new_[3828]_ ,
    \new_[3835]_ , \new_[3836]_ , \new_[3837]_ , \new_[3838]_ ,
    \new_[3839]_ , \new_[3840]_ , \new_[3841]_ , \new_[3842]_ ,
    \new_[3843]_ , \new_[3844]_ , \new_[3845]_ , \new_[3846]_ ,
    \new_[3847]_ , \new_[3848]_ , \new_[3850]_ , \new_[3851]_ ,
    \new_[3853]_ , \new_[3854]_ , \new_[3856]_ , \new_[3857]_ ,
    \new_[3858]_ , \new_[3859]_ , \new_[3860]_ , \new_[3861]_ ,
    \new_[3862]_ , \new_[3863]_ , \new_[3864]_ , \new_[3865]_ ,
    \new_[3866]_ , \new_[3867]_ , \new_[3868]_ , \new_[3869]_ ,
    \new_[3870]_ , \new_[3871]_ , \new_[3872]_ , \new_[3874]_ ,
    \new_[3875]_ , \new_[3876]_ , \new_[3877]_ , \new_[3878]_ ,
    \new_[3879]_ , \new_[3880]_ , \new_[3881]_ , \new_[3882]_ ,
    \new_[3883]_ , \new_[3884]_ , \new_[3885]_ , \new_[3886]_ ,
    \new_[3887]_ , \new_[3888]_ , \new_[3889]_ , \new_[3890]_ ,
    \new_[3891]_ , \new_[3892]_ , \new_[3893]_ , \new_[3894]_ ,
    \new_[3895]_ , \new_[3896]_ , \new_[3897]_ , \new_[3898]_ ,
    \new_[3899]_ , \new_[3900]_ , \new_[3901]_ , \new_[3902]_ ,
    \new_[3903]_ , \new_[3904]_ , \new_[3905]_ , \new_[3906]_ ,
    \new_[3907]_ , \new_[3908]_ , \new_[3909]_ , \new_[3910]_ ,
    \new_[3911]_ , \new_[3912]_ , \new_[3913]_ , \new_[3914]_ ,
    \new_[3915]_ , \new_[3916]_ , \new_[3917]_ , \new_[3918]_ ,
    \new_[3919]_ , \new_[3920]_ , \new_[3921]_ , \new_[3922]_ ,
    \new_[3923]_ , \new_[3924]_ , \new_[3925]_ , \new_[3926]_ ,
    \new_[3927]_ , \new_[3928]_ , \new_[3929]_ , \new_[3930]_ ,
    \new_[3931]_ , \new_[3932]_ , \new_[3933]_ , \new_[3934]_ ,
    \new_[3935]_ , \new_[3936]_ , \new_[3937]_ , \new_[3938]_ ,
    \new_[3939]_ , \new_[3940]_ , \new_[3941]_ , \new_[3942]_ ,
    \new_[3943]_ , \new_[3944]_ , \new_[3945]_ , \new_[3946]_ ,
    \new_[3947]_ , \new_[3948]_ , \new_[3949]_ , \new_[3950]_ ,
    \new_[3951]_ , \new_[3952]_ , \new_[3953]_ , \new_[3954]_ ,
    \new_[3955]_ , \new_[3956]_ , \new_[3957]_ , \new_[3958]_ ,
    \new_[3959]_ , \new_[3960]_ , \new_[3961]_ , \new_[3962]_ ,
    \new_[3963]_ , \new_[3964]_ , \new_[3965]_ , \new_[3966]_ ,
    \new_[3967]_ , \new_[3968]_ , \new_[3969]_ , \new_[3970]_ ,
    \new_[3971]_ , \new_[3972]_ , \new_[3973]_ , \new_[3974]_ ,
    \new_[3975]_ , \new_[3976]_ , \new_[3977]_ , \new_[3978]_ ,
    \new_[3979]_ , \new_[3980]_ , \new_[3981]_ , \new_[3982]_ ,
    \new_[3983]_ , \new_[3984]_ , \new_[3985]_ , \new_[3986]_ ,
    \new_[3987]_ , \new_[3988]_ , \new_[3989]_ , \new_[3990]_ ,
    \new_[3991]_ , \new_[3992]_ , \new_[3993]_ , \new_[3994]_ ,
    \new_[3995]_ , \new_[3996]_ , \new_[3997]_ , \new_[3998]_ ,
    \new_[3999]_ , \new_[4000]_ , \new_[4001]_ , \new_[4002]_ ,
    \new_[4003]_ , \new_[4004]_ , \new_[4005]_ , \new_[4006]_ ,
    \new_[4007]_ , \new_[4008]_ , \new_[4009]_ , \new_[4010]_ ,
    \new_[4011]_ , \new_[4012]_ , \new_[4013]_ , \new_[4014]_ ,
    \new_[4015]_ , \new_[4016]_ , \new_[4017]_ , \new_[4018]_ ,
    \new_[4019]_ , \new_[4020]_ , \new_[4021]_ , \new_[4022]_ ,
    \new_[4023]_ , \new_[4024]_ , \new_[4025]_ , \new_[4026]_ ,
    \new_[4027]_ , \new_[4028]_ , \new_[4029]_ , \new_[4030]_ ,
    \new_[4031]_ , \new_[4032]_ , \new_[4033]_ , \new_[4034]_ ,
    \new_[4035]_ , \new_[4036]_ , \new_[4037]_ , \new_[4038]_ ,
    \new_[4039]_ , \new_[4040]_ , \new_[4041]_ , \new_[4042]_ ,
    \new_[4043]_ , \new_[4045]_ , \new_[4046]_ , \new_[4047]_ ,
    \new_[4048]_ , \new_[4049]_ , \new_[4050]_ , \new_[4051]_ ,
    \new_[4052]_ , \new_[4053]_ , \new_[4054]_ , \new_[4055]_ ,
    \new_[4056]_ , \new_[4057]_ , \new_[4058]_ , \new_[4059]_ ,
    \new_[4060]_ , \new_[4061]_ , \new_[4062]_ , \new_[4063]_ ,
    \new_[4064]_ , \new_[4065]_ , \new_[4066]_ , \new_[4067]_ ,
    \new_[4068]_ , \new_[4069]_ , \new_[4070]_ , \new_[4071]_ ,
    \new_[4072]_ , \new_[4073]_ , \new_[4074]_ , \new_[4075]_ ,
    \new_[4076]_ , \new_[4077]_ , \new_[4078]_ , \new_[4079]_ ,
    \new_[4080]_ , \new_[4081]_ , \new_[4082]_ , \new_[4083]_ ,
    \new_[4084]_ , \new_[4085]_ , \new_[4086]_ , \new_[4087]_ ,
    \new_[4088]_ , \new_[4089]_ , \new_[4090]_ , \new_[4091]_ ,
    \new_[4092]_ , \new_[4093]_ , \new_[4094]_ , \new_[4095]_ ,
    \new_[4096]_ , \new_[4097]_ , \new_[4098]_ , \new_[4099]_ ,
    \new_[4100]_ , \new_[4101]_ , \new_[4102]_ , \new_[4103]_ ,
    \new_[4104]_ , \new_[4105]_ , \new_[4106]_ , \new_[4107]_ ,
    \new_[4108]_ , \new_[4109]_ , \new_[4110]_ , \new_[4111]_ ,
    \new_[4112]_ , \new_[4113]_ , \new_[4114]_ , \new_[4115]_ ,
    \new_[4116]_ , \new_[4117]_ , \new_[4118]_ , \new_[4119]_ ,
    \new_[4120]_ , \new_[4121]_ , \new_[4122]_ , \new_[4123]_ ,
    \new_[4124]_ , \new_[4125]_ , \new_[4126]_ , \new_[4127]_ ,
    \new_[4128]_ , \new_[4129]_ , \new_[4130]_ , \new_[4131]_ ,
    \new_[4132]_ , \new_[4133]_ , \new_[4134]_ , \new_[4135]_ ,
    \new_[4136]_ , \new_[4137]_ , \new_[4138]_ , \new_[4139]_ ,
    \new_[4140]_ , \new_[4141]_ , \new_[4142]_ , \new_[4143]_ ,
    \new_[4144]_ , \new_[4145]_ , \new_[4146]_ , \new_[4147]_ ,
    \new_[4148]_ , \new_[4149]_ , \new_[4150]_ , \new_[4151]_ ,
    \new_[4152]_ , \new_[4153]_ , \new_[4154]_ , \new_[4155]_ ,
    \new_[4156]_ , \new_[4157]_ , \new_[4158]_ , \new_[4159]_ ,
    \new_[4160]_ , \new_[4161]_ , \new_[4162]_ , \new_[4163]_ ,
    \new_[4164]_ , \new_[4165]_ , \new_[4166]_ , \new_[4167]_ ,
    \new_[4168]_ , \new_[4169]_ , \new_[4170]_ , \new_[4171]_ ,
    \new_[4172]_ , \new_[4173]_ , \new_[4174]_ , \new_[4175]_ ,
    \new_[4176]_ , \new_[4177]_ , \new_[4178]_ , \new_[4179]_ ,
    \new_[4180]_ , \new_[4181]_ , \new_[4182]_ , \new_[4183]_ ,
    \new_[4184]_ , \new_[4185]_ , \new_[4186]_ , \new_[4187]_ ,
    \new_[4188]_ , \new_[4189]_ , \new_[4190]_ , \new_[4191]_ ,
    \new_[4192]_ , \new_[4193]_ , \new_[4194]_ , \new_[4195]_ ,
    \new_[4196]_ , \new_[4197]_ , \new_[4198]_ , \new_[4199]_ ,
    \new_[4200]_ , \new_[4201]_ , \new_[4202]_ , \new_[4203]_ ,
    \new_[4204]_ , \new_[4206]_ , \new_[4207]_ , \new_[4208]_ ,
    \new_[4209]_ , \new_[4210]_ , \new_[4211]_ , \new_[4212]_ ,
    \new_[4213]_ , \new_[4214]_ , \new_[4215]_ , \new_[4216]_ ,
    \new_[4217]_ , \new_[4218]_ , \new_[4219]_ , \new_[4220]_ ,
    \new_[4221]_ , \new_[4222]_ , \new_[4223]_ , \new_[4224]_ ,
    \new_[4225]_ , \new_[4226]_ , \new_[4227]_ , \new_[4228]_ ,
    \new_[4229]_ , \new_[4230]_ , \new_[4231]_ , \new_[4232]_ ,
    \new_[4233]_ , \new_[4234]_ , \new_[4235]_ , \new_[4236]_ ,
    \new_[4237]_ , \new_[4238]_ , \new_[4239]_ , \new_[4240]_ ,
    \new_[4241]_ , \new_[4242]_ , \new_[4243]_ , \new_[4244]_ ,
    \new_[4245]_ , \new_[4246]_ , \new_[4247]_ , \new_[4248]_ ,
    \new_[4249]_ , \new_[4250]_ , \new_[4251]_ , \new_[4252]_ ,
    \new_[4253]_ , \new_[4254]_ , \new_[4255]_ , \new_[4256]_ ,
    \new_[4257]_ , \new_[4258]_ , \new_[4259]_ , \new_[4260]_ ,
    \new_[4261]_ , \new_[4263]_ , \new_[4264]_ , \new_[4265]_ ,
    \new_[4266]_ , \new_[4267]_ , \new_[4268]_ , \new_[4269]_ ,
    \new_[4270]_ , \new_[4271]_ , \new_[4272]_ , \new_[4273]_ ,
    \new_[4274]_ , \new_[4277]_ , \new_[4278]_ , \new_[4279]_ ,
    \new_[4280]_ , \new_[4281]_ , \new_[4282]_ , \new_[4283]_ ,
    \new_[4284]_ , \new_[4285]_ , \new_[4286]_ , \new_[4288]_ ,
    \new_[4289]_ , \new_[4290]_ , \new_[4291]_ , \new_[4292]_ ,
    \new_[4293]_ , \new_[4294]_ , \new_[4295]_ , \new_[4296]_ ,
    \new_[4298]_ , \new_[4299]_ , \new_[4300]_ , \new_[4301]_ ,
    \new_[4302]_ , \new_[4303]_ , \new_[4304]_ , \new_[4305]_ ,
    \new_[4306]_ , \new_[4307]_ , \new_[4308]_ , \new_[4309]_ ,
    \new_[4310]_ , \new_[4311]_ , \new_[4312]_ , \new_[4313]_ ,
    \new_[4314]_ , \new_[4315]_ , \new_[4316]_ , \new_[4317]_ ,
    \new_[4318]_ , \new_[4319]_ , \new_[4320]_ , \new_[4321]_ ,
    \new_[4322]_ , \new_[4323]_ , \new_[4324]_ , \new_[4325]_ ,
    \new_[4326]_ , \new_[4327]_ , \new_[4328]_ , \new_[4329]_ ,
    \new_[4330]_ , \new_[4331]_ , \new_[4332]_ , \new_[4333]_ ,
    \new_[4334]_ , \new_[4335]_ , \new_[4336]_ , \new_[4337]_ ,
    \new_[4338]_ , \new_[4339]_ , \new_[4340]_ , \new_[4341]_ ,
    \new_[4342]_ , \new_[4343]_ , \new_[4344]_ , \new_[4345]_ ,
    \new_[4346]_ , \new_[4347]_ , \new_[4348]_ , \new_[4349]_ ,
    \new_[4350]_ , \new_[4351]_ , \new_[4352]_ , \new_[4353]_ ,
    \new_[4354]_ , \new_[4355]_ , \new_[4356]_ , \new_[4357]_ ,
    \new_[4358]_ , \new_[4359]_ , \new_[4360]_ , \new_[4361]_ ,
    \new_[4362]_ , \new_[4363]_ , \new_[4364]_ , \new_[4365]_ ,
    \new_[4366]_ , \new_[4367]_ , \new_[4368]_ , \new_[4369]_ ,
    \new_[4370]_ , \new_[4371]_ , \new_[4372]_ , \new_[4373]_ ,
    \new_[4374]_ , \new_[4375]_ , \new_[4377]_ , \new_[4378]_ ,
    \new_[4379]_ , \new_[4380]_ , \new_[4381]_ , \new_[4382]_ ,
    \new_[4383]_ , \new_[4384]_ , \new_[4385]_ , \new_[4386]_ ,
    \new_[4387]_ , \new_[4388]_ , \new_[4389]_ , \new_[4390]_ ,
    \new_[4391]_ , \new_[4392]_ , \new_[4393]_ , \new_[4394]_ ,
    \new_[4395]_ , \new_[4396]_ , \new_[4397]_ , \new_[4398]_ ,
    \new_[4399]_ , \new_[4400]_ , \new_[4401]_ , \new_[4402]_ ,
    \new_[4403]_ , \new_[4404]_ , \new_[4405]_ , \new_[4406]_ ,
    \new_[4407]_ , \new_[4408]_ , \new_[4409]_ , \new_[4410]_ ,
    \new_[4411]_ , \new_[4412]_ , \new_[4413]_ , \new_[4414]_ ,
    \new_[4415]_ , \new_[4416]_ , \new_[4417]_ , \new_[4418]_ ,
    \new_[4419]_ , \new_[4420]_ , \new_[4421]_ , \new_[4422]_ ,
    \new_[4423]_ , \new_[4424]_ , \new_[4425]_ , \new_[4426]_ ,
    \new_[4427]_ , \new_[4428]_ , \new_[4429]_ , \new_[4430]_ ,
    \new_[4431]_ , \new_[4432]_ , \new_[4433]_ , \new_[4434]_ ,
    \new_[4435]_ , \new_[4436]_ , \new_[4437]_ , \new_[4438]_ ,
    \new_[4439]_ , \new_[4440]_ , \new_[4441]_ , \new_[4442]_ ,
    \new_[4443]_ , \new_[4444]_ , \new_[4445]_ , \new_[4446]_ ,
    \new_[4447]_ , \new_[4448]_ , n866, n871, n876, n881, n886, n891, n896,
    n901, n906, n911, n916, n921, n926, n931, n936, n941, n946, n951, n956,
    n961, n966, n971, n976, n981, n986, n991, n996, n1001, n1006, n1011,
    n1016, n1021, n1026, n1031, n1036, n1041, n1046, n1051, n1056, n1061,
    n1066, n1071, n1076, n1081, n1086, n1091, n1096, n1101, n1106, n1111,
    n1116, n1121, n1126, n1131, n1136, n1141, n1146, n1151, n1156, n1161,
    n1166, n1171, n1176, n1181, n1186, n1191, n1196, n1201, n1206, n1211,
    n1216, n1221, n1226, n1231, n1236, n1241, n1246, n1251, n1256, n1261,
    n1266, n1271, n1276, n1281, n1286, n1291, n1296, n1301, n1306, n1311,
    n1316, n1321, n1326, n1331, n1336, n1341, n1346, n1351, n1356, n1361,
    n1366, n1371, n1376, n1381, n1386, n1391, n1396, n1401, n1406, n1411,
    n1416, n1421, n1426, n1431, n1436, n1441, n1446, n1451, n1456, n1461,
    n1466, n1471, n1476, n1481, n1486, n1491, n1496, n1501, n1506, n1511,
    n1516, n1521, n1526, n1531, n1536, n1541, n1546, n1551, n1556, n1561,
    n1566, n1571, n1576, n1581, n1586, n1591, n1596, n1601, n1606, n1611,
    n1616, n1621, n1626, n1631, n1636, n1641, n1646, n1651, n1656, n1661,
    n1666, n1671, n1676, n1681, n1686, n1691, n1696, n1701, n1706, n1711,
    n1716, n1721, n1726, n1731, n1736, n1741, n1746, n1751, n1756, n1761,
    n1766, n1771, n1776, n1781, n1786, n1791, n1796, n1801, n1806, n1811,
    n1816, n1821, n1826, n1831, n1836, n1841, n1846, n1851, n1856, n1861,
    n1866, n1871, n1876, n1881, n1886, n1891, n1896, n1901, n1906, n1911,
    n1916, n1921, n1926, n1931, n1936, n1941, n1946, n1951, n1956, n1961,
    n1966, n1971, n1976, n1981, n1986, n1991, n1996, n2001, n2006, n2011,
    n2016, n2021, n2026, n2031, n2036, n2041, n2046, n2051, n2056, n2061,
    n2066, n2071, n2076, n2081, n2086, n2091, n2096, n2101, n2106, n2111,
    n2116, n2121, n2126, n2131, n2136, n2141, n2146, n2151, n2156, n2161,
    n2166, n2171, n2176, n2181, n2186, n2191, n2196, n2201, n2206, n2211,
    n2216, n2221, n2226, n2231, n2236, n2241, n2246, n2251, n2256, n2261,
    n2266, n2271, n2276, n2281, n2286, n2291, n2296, n2301, n2306, n2311,
    n2316, n2321, n2326, n2331, n2336, n2341, n2346, n2351, n2356, n2361,
    n2366, n2371, n2376, n2381, n2386, n2391, n2396, n2401, n2406, n2411,
    n2416, n2421, n2426, n2431, n2436, n2441, n2446, n2451, n2456, n2461,
    n2466, n2471, n2476, n2481, n2486, n2491, n2496, n2501, n2506, n2511,
    n2516, n2521, n2526, n2531, n2536, n2541, n2546, n2551, n2556, n2561,
    n2566, n2571, n2576, n2581, n2586, n2591, n2596, n2601, n2606, n2611,
    n2616, n2621, n2626, n2631, n2636, n2641, n2646, n2651, n2656, n2661,
    n2666, n2671, n2676, n2681, n2686, n2691, n2696, n2701, n2706, n2711,
    n2716, n2721, n2726, n2731, n2736, n2741, n2746, n2751, n2756, n2761,
    n2766, n2771, n2776, n2781, n2786, n2791, n2796, n2801, n2806, n2811,
    n2816, n2821, n2826, n2831, n2836, n2841, n2846, n2851, n2856, n2861,
    n2866, n2871, n2876, n2881, n2886, n2891, n2896, n2901, n2906, n2911,
    n2916, n2921, n2926, n2931, n2936, n2941, n2946, n2951, n2956, n2961,
    n2966, n2971, n2976, n2981, n2986, n2991, n2996, n3001, n3006, n3011,
    n3016, n3021, n3026, n3031, n3036, n3041, n3046, n3051, n3056, n3061,
    n3066, n3071, n3076, n3081, n3086, n3091, n3096, n3101, n3106, n3111,
    n3116, n3121, n3126, n3131, n3136, n3141, n3146, n3151, n3156, n3161,
    n3166, n3171, n3176, n3181, n3186, n3191, n3196, n3201, n3206, n3211,
    n3216, n3221, n3226, n3231, n3236, n3241, n3246, n3251, n3256, n3261,
    n3266, n3271, n3276, n3281, n3286, n3291, n3296, n3301, n3306, n3311,
    n3316, n3321, n3326, n3331, n3336, n3341, n3346, n3351, n3356, n3361,
    n3366, n3371, n3376, n3381, n3386, n3391, n3396, n3401, n3406, n3411,
    n3416, n3421, n3426, n3431, n3436, n3441, n3446, n3451, n3456, n3461,
    n3466, n3471, n3476, n3481, n3486, n3491, n3496, n3501, n3506, n3511,
    n3516, n3521, n3526, n3531, n3536, n3541, n3546, n3551, n3556, n3561,
    n3566, n3571, n3576, n3581, n3586, n3591, n3596, n3601, n3606, n3611,
    n3616, n3621, n3626, n3631, n3636, n3641, n3646, n3651, n3656, n3661,
    n3666, n3671, n3676;
  assign wb0_stb_o = wb1_stb_i ? \new_[3574]_  : \new_[1001]_ ;
  assign wb1_stb_o = wb0_stb_i ? \new_[3592]_  : \new_[1025]_ ;
  assign wb0_cyc_o = wb1_cyc_i ? \new_[3574]_  : \new_[1030]_ ;
  assign wb1_cyc_o = wb0_cyc_i ? \new_[3592]_  : \new_[1058]_ ;
  assign \new_[1001]_  = u3_u0_mast_stb_reg;
  assign \wb0_addr_o[3]  = \wb1_addr_i[3]  ? \new_[3574]_  : \new_[1060]_ ;
  assign \wb0_addr_o[2]  = \wb1_addr_i[2]  ? \new_[3574]_  : \new_[1061]_ ;
  assign \wb0_addr_o[27]  = \wb1_addr_i[27]  ? \new_[3574]_  : \new_[1091]_ ;
  assign \wb0_addr_o[26]  = \wb1_addr_i[26]  ? \new_[3574]_  : \new_[1092]_ ;
  assign \wb0_addr_o[25]  = \wb1_addr_i[25]  ? \new_[3574]_  : \new_[1070]_ ;
  assign \wb0_addr_o[24]  = \wb1_addr_i[24]  ? \new_[3574]_  : \new_[1093]_ ;
  assign \wb0_addr_o[23]  = \wb1_addr_i[23]  ? \new_[3574]_  : \new_[1067]_ ;
  assign \wb0_addr_o[22]  = \wb1_addr_i[22]  ? \new_[3574]_  : \new_[1068]_ ;
  assign \wb0_addr_o[21]  = \wb1_addr_i[21]  ? \new_[3574]_  : \new_[1069]_ ;
  assign \wb0_addr_o[20]  = \wb1_addr_i[20]  ? \new_[3574]_  : \new_[1071]_ ;
  assign \wb0_addr_o[19]  = \wb1_addr_i[19]  ? \new_[3574]_  : \new_[1072]_ ;
  assign \wb0_addr_o[18]  = \wb1_addr_i[18]  ? \new_[3659]_  : \new_[1073]_ ;
  assign \wb0_addr_o[15]  = \wb1_addr_i[15]  ? \new_[3659]_  : \new_[1075]_ ;
  assign \wb0_addr_o[14]  = \wb1_addr_i[14]  ? \new_[3574]_  : \new_[1076]_ ;
  assign \wb0_addr_o[13]  = \wb1_addr_i[13]  ? \new_[3659]_  : \new_[1077]_ ;
  assign \wb0_addr_o[12]  = \wb1_addr_i[12]  ? \new_[3659]_  : \new_[1078]_ ;
  assign \wb0_addr_o[11]  = \wb1_addr_i[11]  ? \new_[3574]_  : \new_[1079]_ ;
  assign \wb0_addr_o[10]  = \wb1_addr_i[10]  ? \new_[3659]_  : \new_[1080]_ ;
  assign \wb0_addr_o[9]  = \wb1_addr_i[9]  ? \new_[3659]_  : \new_[1081]_ ;
  assign \wb0_addr_o[16]  = \wb1_addr_i[16]  ? \new_[3659]_  : \new_[1074]_ ;
  assign \wb0_addr_o[4]  = \wb1_addr_i[4]  ? \new_[3574]_  : \new_[1084]_ ;
  assign \wb0_addr_o[6]  = \wb1_addr_i[6]  ? \new_[3574]_  : \new_[1082]_ ;
  assign \wb0_addr_o[5]  = \wb1_addr_i[5]  ? \new_[3659]_  : \new_[1083]_ ;
  assign \new_[1025]_  = u4_u0_mast_stb_reg;
  assign \wb0_addr_o[28]  = \wb1_addr_i[28]  ? \new_[3574]_  : \new_[1090]_ ;
  assign \wb0_addr_o[29]  = \wb1_addr_i[29]  ? \new_[3659]_  : \new_[1089]_ ;
  assign \wb0_addr_o[31]  = \wb1_addr_i[31]  ? \new_[3574]_  : \new_[1123]_ ;
  assign \wb0_addr_o[30]  = \wb1_addr_i[30]  ? \new_[3574]_  : \new_[1124]_ ;
  assign \new_[1030]_  = u3_u0_mast_cyc_reg;
  assign \wb0_addr_o[17]  = \wb1_addr_i[17]  ? \new_[3659]_  : \new_[1094]_ ;
  assign \wb0_addr_o[8]  = \wb1_addr_i[8]  ? \new_[3659]_  : \new_[1096]_ ;
  assign \wb0_addr_o[7]  = \wb1_addr_i[7]  ? \new_[3659]_  : \new_[1095]_ ;
  assign \wb1_addr_o[27]  = \wb0_addr_i[27]  ? \new_[3592]_  : \new_[1100]_ ;
  assign \wb1_addr_o[26]  = \wb0_addr_i[26]  ? \new_[3607]_  : \new_[1101]_ ;
  assign \wb1_addr_o[25]  = \wb0_addr_i[25]  ? \new_[3607]_  : \new_[1102]_ ;
  assign \wb1_addr_o[24]  = \wb0_addr_i[24]  ? \new_[3607]_  : \new_[1103]_ ;
  assign \wb1_addr_o[23]  = \wb0_addr_i[23]  ? \new_[3606]_  : \new_[1105]_ ;
  assign \wb1_addr_o[22]  = \wb0_addr_i[22]  ? \new_[3592]_  : \new_[1104]_ ;
  assign \wb1_addr_o[21]  = \wb0_addr_i[21]  ? \new_[3592]_  : \new_[1106]_ ;
  assign \wb1_addr_o[20]  = \wb0_addr_i[20]  ? \new_[3592]_  : \new_[1107]_ ;
  assign \wb1_addr_o[19]  = \wb0_addr_i[19]  ? \new_[3592]_  : \new_[1108]_ ;
  assign \wb1_addr_o[18]  = \wb0_addr_i[18]  ? \new_[3592]_  : \new_[1109]_ ;
  assign \wb1_addr_o[16]  = \wb0_addr_i[16]  ? \new_[3592]_  : \new_[1110]_ ;
  assign \wb1_addr_o[15]  = \wb0_addr_i[15]  ? \new_[3606]_  : \new_[1111]_ ;
  assign \wb1_addr_o[14]  = \wb0_addr_i[14]  ? \new_[3592]_  : \new_[1114]_ ;
  assign \wb1_addr_o[13]  = \wb0_addr_i[13]  ? \new_[3607]_  : \new_[1112]_ ;
  assign \wb1_addr_o[12]  = \wb0_addr_i[12]  ? \new_[3607]_  : \new_[1113]_ ;
  assign \wb1_addr_o[11]  = \wb0_addr_i[11]  ? \new_[3607]_  : \new_[1115]_ ;
  assign \wb1_addr_o[9]  = \wb0_addr_i[9]  ? \new_[3592]_  : \new_[1117]_ ;
  assign \wb1_addr_o[6]  = \wb0_addr_i[6]  ? \new_[3607]_  : \new_[1118]_ ;
  assign \wb1_addr_o[5]  = \wb0_addr_i[5]  ? \new_[3592]_  : \new_[1119]_ ;
  assign \wb1_addr_o[4]  = \wb0_addr_i[4]  ? \new_[3592]_  : \new_[1120]_ ;
  assign n866 = \new_[1157]_  & n876;
  assign \wb1_addr_o[29]  = \wb0_addr_i[29]  ? \new_[3592]_  : \new_[1098]_ ;
  assign \wb1_addr_o[28]  = \wb0_addr_i[28]  ? \new_[3606]_  : \new_[1099]_ ;
  assign \wb1_addr_o[10]  = \wb0_addr_i[10]  ? \new_[3592]_  : \new_[1116]_ ;
  assign \new_[1058]_  = u4_u0_mast_cyc_reg;
  assign n871 = ~\new_[1200]_  & ~\new_[1097]_ ;
  assign \new_[1060]_  = \\u2_mast0_adr_reg[3] ;
  assign \new_[1061]_  = \\u2_mast0_adr_reg[2] ;
  assign \wb1_addr_o[30]  = \wb0_addr_i[30]  ? \new_[3606]_  : \new_[1149]_ ;
  assign \wb1_addr_o[31]  = \wb0_addr_i[31]  ? \new_[3606]_  : \new_[1148]_ ;
  assign \wb1_addr_o[17]  = \wb0_addr_i[17]  ? \new_[3592]_  : \new_[1150]_ ;
  assign \wb1_addr_o[7]  = \wb0_addr_i[7]  ? \new_[3592]_  : \new_[1152]_ ;
  assign \wb1_addr_o[8]  = \wb0_addr_i[8]  ? \new_[3607]_  : \new_[1151]_ ;
  assign \new_[1067]_  = \\u2_mast0_adr_reg[23] ;
  assign \new_[1068]_  = \\u2_mast0_adr_reg[22] ;
  assign \new_[1069]_  = \\u2_mast0_adr_reg[21] ;
  assign \new_[1070]_  = \\u2_mast0_adr_reg[25] ;
  assign \new_[1071]_  = \\u2_mast0_adr_reg[20] ;
  assign \new_[1072]_  = \\u2_mast0_adr_reg[19] ;
  assign \new_[1073]_  = \\u2_mast0_adr_reg[18] ;
  assign \new_[1074]_  = \\u2_mast0_adr_reg[16] ;
  assign \new_[1075]_  = \\u2_mast0_adr_reg[15] ;
  assign \new_[1076]_  = \\u2_mast0_adr_reg[14] ;
  assign \new_[1077]_  = \\u2_mast0_adr_reg[13] ;
  assign \new_[1078]_  = \\u2_mast0_adr_reg[12] ;
  assign \new_[1079]_  = \\u2_mast0_adr_reg[11] ;
  assign \new_[1080]_  = \\u2_mast0_adr_reg[10] ;
  assign \new_[1081]_  = \\u2_mast0_adr_reg[9] ;
  assign \new_[1082]_  = \\u2_mast0_adr_reg[6] ;
  assign \new_[1083]_  = \\u2_mast0_adr_reg[5] ;
  assign \new_[1084]_  = \\u2_mast0_adr_reg[4] ;
  assign n876 = ~\new_[1195]_  | ~\new_[4200]_  | ~\new_[1165]_ ;
  assign n881 = ~\new_[1097]_ ;
  assign \wb1_addr_o[3]  = \wb0_addr_i[3]  ? \new_[3592]_  : \new_[1167]_ ;
  assign \wb1_addr_o[2]  = \wb0_addr_i[2]  ? \new_[3592]_  : \new_[1168]_ ;
  assign \new_[1089]_  = \\u2_mast0_adr_reg[29] ;
  assign \new_[1090]_  = \\u2_mast0_adr_reg[28] ;
  assign \new_[1091]_  = \\u2_mast0_adr_reg[27] ;
  assign \new_[1092]_  = \\u2_mast0_adr_reg[26] ;
  assign \new_[1093]_  = \\u2_mast0_adr_reg[24] ;
  assign \new_[1094]_  = \\u2_mast0_adr_reg[17] ;
  assign \new_[1095]_  = \\u2_mast0_adr_reg[7] ;
  assign \new_[1096]_  = \\u2_mast0_adr_reg[8] ;
  assign \new_[1097]_  = ~\new_[1166]_  & (~\new_[1255]_  | ~\new_[2541]_ );
  assign \new_[1098]_  = \\u2_mast1_adr_reg[29] ;
  assign \new_[1099]_  = \\u2_mast1_adr_reg[28] ;
  assign \new_[1100]_  = \\u2_mast1_adr_reg[27] ;
  assign \new_[1101]_  = \\u2_mast1_adr_reg[26] ;
  assign \new_[1102]_  = \\u2_mast1_adr_reg[25] ;
  assign \new_[1103]_  = \\u2_mast1_adr_reg[24] ;
  assign \new_[1104]_  = \\u2_mast1_adr_reg[22] ;
  assign \new_[1105]_  = \\u2_mast1_adr_reg[23] ;
  assign \new_[1106]_  = \\u2_mast1_adr_reg[21] ;
  assign \new_[1107]_  = \\u2_mast1_adr_reg[20] ;
  assign \new_[1108]_  = \\u2_mast1_adr_reg[19] ;
  assign \new_[1109]_  = \\u2_mast1_adr_reg[18] ;
  assign \new_[1110]_  = \\u2_mast1_adr_reg[16] ;
  assign \new_[1111]_  = \\u2_mast1_adr_reg[15] ;
  assign \new_[1112]_  = \\u2_mast1_adr_reg[13] ;
  assign \new_[1113]_  = \\u2_mast1_adr_reg[12] ;
  assign \new_[1114]_  = \\u2_mast1_adr_reg[14] ;
  assign \new_[1115]_  = \\u2_mast1_adr_reg[11] ;
  assign \new_[1116]_  = \\u2_mast1_adr_reg[10] ;
  assign \new_[1117]_  = \\u2_mast1_adr_reg[9] ;
  assign \new_[1118]_  = \\u2_mast1_adr_reg[6] ;
  assign \new_[1119]_  = \\u2_mast1_adr_reg[5] ;
  assign \new_[1120]_  = \\u2_mast1_adr_reg[4] ;
  assign n891 = ~\new_[1159]_  | ~\new_[1333]_ ;
  assign n886 = ~\new_[1162]_  | ~\new_[1332]_ ;
  assign \new_[1123]_  = \\u2_mast0_adr_reg[31] ;
  assign \new_[1124]_  = \\u2_mast0_adr_reg[30] ;
  assign n951 = ~\new_[4203]_  & ~\new_[1203]_ ;
  assign n956 = ~\new_[4203]_  & ~\new_[1201]_ ;
  assign n946 = ~\new_[4203]_  & ~\new_[1204]_ ;
  assign n941 = ~\new_[4204]_  & ~\new_[1205]_ ;
  assign n936 = ~\new_[4204]_  & ~\new_[1206]_ ;
  assign n931 = ~\new_[4203]_  & ~\new_[1207]_ ;
  assign n926 = ~\new_[4203]_  & ~\new_[1209]_ ;
  assign n916 = ~\new_[4203]_  & ~\new_[1211]_ ;
  assign n921 = ~\new_[4204]_  & ~\new_[1210]_ ;
  assign n906 = ~\new_[4204]_  & ~\new_[1212]_ ;
  assign n901 = ~\new_[4204]_  & ~\new_[1213]_ ;
  assign n896 = ~\new_[4203]_  & ~\new_[1214]_ ;
  assign n1006 = ~\new_[4204]_  & ~\new_[1215]_ ;
  assign n911 = ~\new_[4204]_  & ~\new_[1216]_ ;
  assign n1001 = ~\new_[4203]_  & ~\new_[1217]_ ;
  assign n996 = ~\new_[4203]_  & ~\new_[1218]_ ;
  assign n991 = ~\new_[4204]_  & ~\new_[1219]_ ;
  assign n986 = ~\new_[4203]_  & ~\new_[1220]_ ;
  assign n961 = ~\new_[4204]_  & ~\new_[1202]_ ;
  assign n981 = ~\new_[4204]_  & ~\new_[1189]_ ;
  assign n971 = ~\new_[4204]_  & ~\new_[1191]_ ;
  assign n976 = ~\new_[4203]_  & ~\new_[1190]_ ;
  assign n966 = ~\new_[4204]_  & ~\new_[1194]_ ;
  assign \new_[1148]_  = \\u2_mast1_adr_reg[31] ;
  assign \new_[1149]_  = \\u2_mast1_adr_reg[30] ;
  assign \new_[1150]_  = \\u2_mast1_adr_reg[17] ;
  assign \new_[1151]_  = \\u2_mast1_adr_reg[8] ;
  assign \new_[1152]_  = \\u2_mast1_adr_reg[7] ;
  assign n1136 = ~\new_[1189]_ ;
  assign n1131 = ~\new_[1190]_ ;
  assign n1126 = ~\new_[1191]_ ;
  assign n1121 = ~\new_[1194]_ ;
  assign \new_[1157]_  = ~\new_[1226]_  | ~\new_[1726]_ ;
  assign n1011 = ~\new_[4202]_  & ~\new_[1256]_ ;
  assign \new_[1159]_  = ~\new_[4200]_  | ~n1181;
  assign n1146 = ~\new_[4202]_  & ~\new_[1258]_ ;
  assign n1141 = ~\new_[4202]_  & ~\new_[1222]_ ;
  assign \new_[1162]_  = ~\new_[4200]_  | ~n1176;
  assign n1016 = ~\new_[4203]_  & ~\new_[1224]_ ;
  assign n1021 = ~\new_[4202]_  & ~\new_[1225]_ ;
  assign \new_[1165]_  = ~\new_[1255]_  | ~\new_[2508]_ ;
  assign \new_[1166]_  = ~\new_[1253]_  & ~\new_[1320]_ ;
  assign \new_[1167]_  = \\u2_mast1_adr_reg[3] ;
  assign \new_[1168]_  = \\u2_mast1_adr_reg[2] ;
  assign n1111 = ~\new_[1201]_ ;
  assign n1116 = ~\new_[1202]_ ;
  assign n1101 = ~\new_[1203]_ ;
  assign n1096 = ~\new_[1204]_ ;
  assign n1106 = ~\new_[1205]_ ;
  assign n1091 = ~\new_[1206]_ ;
  assign n1086 = ~\new_[1207]_ ;
  assign n1081 = ~\new_[1209]_ ;
  assign n1076 = ~\new_[1210]_ ;
  assign n1071 = ~\new_[1211]_ ;
  assign n1066 = ~\new_[1212]_ ;
  assign n1056 = ~\new_[1213]_ ;
  assign n1061 = ~\new_[1214]_ ;
  assign n1051 = ~\new_[1215]_ ;
  assign n1046 = ~\new_[1216]_ ;
  assign n1041 = ~\new_[1217]_ ;
  assign n1036 = ~\new_[1218]_ ;
  assign n1031 = ~\new_[1219]_ ;
  assign n1026 = ~\new_[1220]_ ;
  assign n1151 = ~\new_[1222]_ ;
  assign \new_[1189]_  = ~\new_[1278]_  & (~\new_[1324]_  | ~\new_[1239]_ );
  assign \new_[1190]_  = ~\new_[1279]_  & (~\new_[1325]_  | ~\new_[1240]_ );
  assign \new_[1191]_  = ~\new_[1280]_  & (~\new_[1324]_  | ~\new_[1241]_ );
  assign n1171 = ~\new_[1224]_ ;
  assign n1166 = ~\new_[1225]_ ;
  assign \new_[1194]_  = ~\new_[1281]_  & (~\new_[1324]_  | ~\new_[1244]_ );
  assign \new_[1195]_  = ~\new_[2568]_  | ~n1361 | ~\new_[1317]_ ;
  assign \new_[1196]_  = \\u2_state_reg[1] ;
  assign \new_[1197]_  = \\u2_state_reg[3] ;
  assign \new_[1198]_  = ~u2_chunk_dec_reg;
  assign \new_[1199]_  = ~u2_tsz_dec_reg;
  assign \new_[1200]_  = \new_[1282]_  & \new_[1729]_ ;
  assign \new_[1201]_  = ~\new_[1260]_  & (~\new_[1324]_  | ~\new_[1246]_ );
  assign \new_[1202]_  = ~\new_[1259]_  & (~\new_[1325]_  | ~\new_[1245]_ );
  assign \new_[1203]_  = ~\new_[1261]_  & (~\new_[1325]_  | ~\new_[1247]_ );
  assign \new_[1204]_  = ~\new_[1262]_  & (~\new_[1324]_  | ~\new_[1248]_ );
  assign \new_[1205]_  = ~\new_[1263]_  & (~\new_[1325]_  | ~\new_[1287]_ );
  assign \new_[1206]_  = ~\new_[1264]_  & (~\new_[1325]_  | ~\new_[1249]_ );
  assign \new_[1207]_  = ~\new_[1265]_  & (~\new_[1324]_  | ~\new_[1250]_ );
  assign n1161 = ~\new_[1256]_ ;
  assign \new_[1209]_  = ~\new_[1266]_  & (~\new_[1324]_  | ~\new_[1238]_ );
  assign \new_[1210]_  = ~\new_[1267]_  & (~\new_[1325]_  | ~\new_[1236]_ );
  assign \new_[1211]_  = ~\new_[1268]_  & (~\new_[1325]_  | ~\new_[1233]_ );
  assign \new_[1212]_  = ~\new_[1269]_  & (~\new_[1325]_  | ~\new_[1232]_ );
  assign \new_[1213]_  = ~\new_[1270]_  & (~\new_[1325]_  | ~\new_[1231]_ );
  assign \new_[1214]_  = ~\new_[1271]_  & (~\new_[1325]_  | ~\new_[1237]_ );
  assign \new_[1215]_  = ~\new_[1272]_  & (~\new_[1324]_  | ~\new_[1285]_ );
  assign \new_[1216]_  = ~\new_[1273]_  & (~\new_[1324]_  | ~\new_[1229]_ );
  assign \new_[1217]_  = ~\new_[1274]_  & (~\new_[1324]_  | ~\new_[3959]_ );
  assign \new_[1218]_  = ~\new_[1275]_  & (~\new_[1324]_  | ~\new_[1234]_ );
  assign \new_[1219]_  = ~\new_[1276]_  & (~\new_[1325]_  | ~\new_[1284]_ );
  assign \new_[1220]_  = ~\new_[1277]_  & (~\new_[1325]_  | ~\new_[1228]_ );
  assign n1156 = ~\new_[1258]_ ;
  assign \new_[1222]_  = \new_[1415]_  ? \new_[1326]_  : \new_[1235]_ ;
  assign n1176 = ~\new_[1292]_  | (~\new_[1326]_  & ~\new_[1592]_ );
  assign \new_[1224]_  = \new_[1385]_  ? \new_[1326]_  : \new_[1242]_ ;
  assign \new_[1225]_  = \new_[1386]_  ? \new_[1326]_  : \new_[1243]_ ;
  assign \new_[1226]_  = ~\new_[1291]_  & ~\new_[4201]_ ;
  assign \new_[1227]_  = ~\\u2_adr1_cnt_reg[28] ;
  assign \new_[1228]_  = \\u2_adr1_cnt_reg[27] ;
  assign \new_[1229]_  = \\u2_adr1_cnt_reg[23] ;
  assign \new_[1230]_  = ~\\u2_adr1_cnt_reg[24] ;
  assign \new_[1231]_  = \\u2_adr1_cnt_reg[20] ;
  assign \new_[1232]_  = \\u2_adr1_cnt_reg[19] ;
  assign \new_[1233]_  = \\u2_adr1_cnt_reg[18] ;
  assign \new_[1234]_  = \\u2_adr1_cnt_reg[25] ;
  assign \new_[1235]_  = ~\\u2_adr1_cnt_reg[29] ;
  assign \new_[1236]_  = \\u2_adr1_cnt_reg[17] ;
  assign \new_[1237]_  = \\u2_adr1_cnt_reg[21] ;
  assign \new_[1238]_  = \\u2_adr1_cnt_reg[16] ;
  assign \new_[1239]_  = \\u2_adr1_cnt_reg[2] ;
  assign \new_[1240]_  = \\u2_adr1_cnt_reg[3] ;
  assign \new_[1241]_  = \\u2_adr1_cnt_reg[4] ;
  assign \new_[1242]_  = ~\\u2_adr1_cnt_reg[5] ;
  assign \new_[1243]_  = ~\\u2_adr1_cnt_reg[6] ;
  assign \new_[1244]_  = \\u2_adr1_cnt_reg[7] ;
  assign \new_[1245]_  = \\u2_adr1_cnt_reg[8] ;
  assign \new_[1246]_  = \\u2_adr1_cnt_reg[9] ;
  assign \new_[1247]_  = \\u2_adr1_cnt_reg[10] ;
  assign \new_[1248]_  = \\u2_adr1_cnt_reg[11] ;
  assign \new_[1249]_  = \\u2_adr1_cnt_reg[13] ;
  assign \new_[1250]_  = \\u2_adr1_cnt_reg[14] ;
  assign \new_[1251]_  = ~\\u2_adr1_cnt_reg[15] ;
  assign \new_[1252]_  = u2_read_r_reg;
  assign \new_[1253]_  = ~\new_[1317]_  | ~\new_[2586]_ ;
  assign wb0_we_o = wb1_we_i ? \new_[3574]_  : \new_[1329]_ ;
  assign \new_[1255]_  = ~\new_[1318]_  | ~\new_[1319]_ ;
  assign \new_[1256]_  = \new_[1416]_  ? \new_[1326]_  : \new_[1251]_ ;
  assign n1181 = \new_[3973]_  ? \new_[1326]_  : \new_[3997]_ ;
  assign \new_[1258]_  = \new_[1369]_  ? \new_[1324]_  : \new_[1227]_ ;
  assign \new_[1259]_  = \new_[1327]_  & \new_[1387]_ ;
  assign \new_[1260]_  = \new_[1327]_  & \new_[1345]_ ;
  assign \new_[1261]_  = \new_[1327]_  & \new_[1376]_ ;
  assign \new_[1262]_  = \new_[1327]_  & \new_[1377]_ ;
  assign \new_[1263]_  = \new_[1327]_  & \new_[1378]_ ;
  assign \new_[1264]_  = \new_[1327]_  & \new_[1379]_ ;
  assign \new_[1265]_  = \new_[1327]_  & \new_[1406]_ ;
  assign \new_[1266]_  = \new_[1327]_  & \new_[1339]_ ;
  assign \new_[1267]_  = \new_[1327]_  & \new_[1380]_ ;
  assign \new_[1268]_  = \new_[1327]_  & \new_[1375]_ ;
  assign \new_[1269]_  = \new_[1327]_  & \new_[1414]_ ;
  assign \new_[1270]_  = ~\new_[1326]_  & ~\new_[1374]_ ;
  assign \new_[1271]_  = \new_[1327]_  & \new_[1381]_ ;
  assign \new_[1272]_  = \new_[1327]_  & \new_[1413]_ ;
  assign \new_[1273]_  = \new_[1327]_  & \new_[1372]_ ;
  assign \new_[1274]_  = \new_[1327]_  & \new_[1371]_ ;
  assign \new_[1275]_  = \new_[1327]_  & \new_[1382]_ ;
  assign \new_[1276]_  = \new_[1327]_  & \new_[1373]_ ;
  assign \new_[1277]_  = \new_[1327]_  & \new_[1370]_ ;
  assign \new_[1278]_  = \new_[1327]_  & \new_[1383]_ ;
  assign \new_[1279]_  = \new_[1327]_  & \new_[1384]_ ;
  assign \new_[1280]_  = \new_[1327]_  & \new_[1389]_ ;
  assign \new_[1281]_  = \new_[1327]_  & \new_[1388]_ ;
  assign \new_[1282]_  = ~\new_[1327]_  | ~\new_[2541]_ ;
  assign n1186 = ~\new_[2168]_  | ~\new_[1348]_  | ~\new_[3017]_  | ~\new_[3103]_ ;
  assign \new_[1284]_  = \\u2_adr1_cnt_reg[26] ;
  assign \new_[1285]_  = \\u2_adr1_cnt_reg[22] ;
  assign n3471 = ~\\u2_adr1_cnt_reg[0] ;
  assign \new_[1287]_  = \\u2_adr1_cnt_reg[12] ;
  assign \new_[1288]_  = ~\\u2_adr1_cnt_reg[1] ;
  assign n1191 = ~\new_[3019]_  | ~\new_[1331]_ ;
  assign n1201 = ~\new_[1324]_  & ~\new_[1252]_ ;
  assign \new_[1291]_  = ~\new_[1337]_  & ~\new_[2541]_ ;
  assign \new_[1292]_  = ~\new_[1337]_  | ~\new_[4066]_ ;
  assign n1221 = ~\new_[1958]_  | (~\new_[1367]_  & ~\new_[4308]_ );
  assign n1251 = ~\new_[1952]_  | (~\new_[1365]_  & ~\new_[4288]_ );
  assign n1256 = ~\new_[1942]_  | (~\new_[1366]_  & ~\new_[4288]_ );
  assign n1216 = ~\new_[1957]_  | (~\new_[1368]_  & ~\new_[4288]_ );
  assign n1266 = ~\new_[1860]_  | (~\new_[1351]_  & ~\new_[2245]_ );
  assign n1271 = ~\new_[1861]_  | (~\new_[1352]_  & ~\new_[4288]_ );
  assign n1276 = ~\new_[1862]_  | (~\new_[1354]_  & ~\new_[2243]_ );
  assign n1281 = ~\new_[1863]_  | (~\new_[1355]_  & ~\new_[4288]_ );
  assign n1286 = ~\new_[1864]_  | (~\new_[1356]_  & ~\new_[2245]_ );
  assign n1291 = ~\new_[1865]_  | (~\new_[1357]_  & ~\new_[4288]_ );
  assign n1296 = ~\new_[1866]_  | (~\new_[1358]_  & ~\new_[4288]_ );
  assign n1301 = ~\new_[1867]_  | (~\new_[1359]_  & ~\new_[4288]_ );
  assign n1306 = ~\new_[1945]_  | (~\new_[1360]_  & ~\new_[2243]_ );
  assign n1311 = ~\new_[1946]_  | (~\new_[1361]_  & ~\new_[4288]_ );
  assign n1316 = ~\new_[1948]_  | (~\new_[1362]_  & ~\new_[4288]_ );
  assign n1321 = ~\new_[1949]_  | (~\new_[1363]_  & ~\new_[2245]_ );
  assign n1326 = ~\new_[1950]_  | (~\new_[1364]_  & ~\new_[4288]_ );
  assign n1206 = ~\new_[1858]_  | (~\new_[1404]_  & ~\new_[4288]_ );
  assign n1211 = ~\new_[1857]_  | (~\new_[1349]_  & ~\new_[2246]_ );
  assign n1226 = ~\new_[1955]_  | (~\new_[1403]_  & ~\new_[4288]_ );
  assign n1236 = ~\new_[1953]_  | (~\new_[1346]_  & ~\new_[4288]_ );
  assign n1261 = ~\new_[1951]_  | ~\new_[1343]_ ;
  assign n1246 = ~\new_[1859]_  | (~\new_[1353]_  & ~\new_[2245]_ );
  assign n1231 = ~\new_[1954]_  | (~\new_[1344]_  & ~\new_[4288]_ );
  assign \new_[1317]_  = u2_write_hold_r_reg;
  assign \new_[1318]_  = ~\new_[1562]_  | ~n1361;
  assign \new_[1319]_  = ~\new_[1350]_  | ~\new_[1588]_ ;
  assign \new_[1320]_  = ~n1361;
  assign n1346 = ~\new_[1334]_ ;
  assign n1351 = ~\new_[1947]_  | (~\new_[1411]_  & ~\new_[2243]_ );
  assign n1356 = ~\new_[1335]_ ;
  assign \new_[1324]_  = ~n1331;
  assign \new_[1325]_  = \new_[1337]_ ;
  assign \new_[1326]_  = ~\new_[1338]_ ;
  assign \new_[1327]_  = ~\new_[1337]_ ;
  assign n1341 = ~\new_[1956]_  | (~\new_[1434]_  & ~\new_[2244]_ );
  assign \new_[1329]_  = u3_u0_mast_we_r_reg;
  assign n1336 = ~\new_[1856]_  | (~\new_[1412]_  & ~\new_[4288]_ );
  assign \new_[1331]_  = ~\new_[1347]_  & ~\new_[2061]_ ;
  assign \new_[1332]_  = ~\new_[4202]_  | ~\new_[1560]_  | ~\new_[2862]_ ;
  assign \new_[1333]_  = ~\new_[1560]_  | ~\new_[2821]_  | ~\new_[4202]_ ;
  assign \new_[1334]_  = (~\new_[1443]_  | ~\new_[2186]_ ) & (~\new_[4093]_  | ~\new_[2064]_ );
  assign \new_[1335]_  = (~\new_[1445]_  | ~\new_[2186]_ ) & (~\new_[3976]_  | ~\new_[2064]_ );
  assign n1331 = \new_[1350]_ ;
  assign \new_[1337]_  = ~\new_[1350]_ ;
  assign \new_[1338]_  = \new_[1350]_ ;
  assign \new_[1339]_  = \\u2_adr0_cnt_reg[16] ;
  assign \new_[1340]_  = ~\\u0_u0_int_src_r_reg[2] ;
  assign dma_ack_o = \\u1_ack_o_reg[0] ;
  assign \new_[1342]_  = u1_next_start_reg;
  assign \new_[1343]_  = ~\new_[1407]_  | ~\new_[2186]_ ;
  assign \new_[1344]_  = ~\new_[1439]_  & (~\new_[4293]_  | ~\new_[1232]_ );
  assign \new_[1345]_  = \\u2_adr0_cnt_reg[9] ;
  assign \new_[1346]_  = ~\new_[1444]_  & (~\new_[1493]_  | ~\new_[1233]_ );
  assign \new_[1347]_  = ~\new_[3222]_  & (~\new_[1492]_  | ~\new_[2428]_ );
  assign \new_[1348]_  = ~\new_[1405]_ ;
  assign \new_[1349]_  = ~\new_[1447]_  & (~\new_[4293]_  | ~\new_[1228]_ );
  assign \new_[1350]_  = ~\new_[4377]_ ;
  assign \new_[1351]_  = ~\new_[1448]_  & (~\new_[4293]_  | ~\new_[1239]_ );
  assign \new_[1352]_  = ~\new_[1449]_  & (~\new_[4293]_  | ~\new_[1240]_ );
  assign \new_[1353]_  = ~\new_[1462]_  & (~\new_[1493]_  | ~\new_[3987]_ );
  assign \new_[1354]_  = ~\new_[1450]_  & (~\new_[4293]_  | ~\new_[1241]_ );
  assign \new_[1355]_  = ~\new_[1451]_  & (~\new_[1518]_  | ~\new_[4154]_ );
  assign \new_[1356]_  = ~\new_[1452]_  & (~\new_[1518]_  | ~\new_[3989]_ );
  assign \new_[1357]_  = ~\new_[1453]_  & (~\new_[1518]_  | ~\new_[1244]_ );
  assign \new_[1358]_  = ~\new_[1454]_  & (~\new_[1518]_  | ~\new_[1245]_ );
  assign \new_[1359]_  = ~\new_[1455]_  & (~\new_[4293]_  | ~\new_[1246]_ );
  assign \new_[1360]_  = ~\new_[1456]_  & (~\new_[1518]_  | ~\new_[1247]_ );
  assign \new_[1361]_  = ~\new_[1458]_  & (~\new_[1517]_  | ~\new_[1248]_ );
  assign \new_[1362]_  = ~\new_[1459]_  & (~\new_[1517]_  | ~\new_[1249]_ );
  assign \new_[1363]_  = ~\new_[1460]_  & (~\new_[1517]_  | ~\new_[1250]_ );
  assign \new_[1364]_  = ~\new_[1461]_  & (~\new_[1517]_  | ~\new_[4080]_ );
  assign \new_[1365]_  = ~\new_[1464]_  & (~\new_[1517]_  | ~\new_[1236]_ );
  assign \new_[1366]_  = ~\new_[1465]_  & (~\new_[4293]_  | ~\new_[1237]_ );
  assign \new_[1367]_  = ~\new_[1471]_  & (~\new_[1493]_  | ~\new_[3959]_ );
  assign \new_[1368]_  = ~\new_[1470]_  & (~\new_[4293]_  | ~\new_[1229]_ );
  assign \new_[1369]_  = ~\\u2_adr0_cnt_reg[28] ;
  assign \new_[1370]_  = \\u2_adr0_cnt_reg[27] ;
  assign \new_[1371]_  = \\u2_adr0_cnt_reg[24] ;
  assign \new_[1372]_  = \\u2_adr0_cnt_reg[23] ;
  assign \new_[1373]_  = \\u2_adr0_cnt_reg[26] ;
  assign \new_[1374]_  = ~\\u2_adr0_cnt_reg[20] ;
  assign \new_[1375]_  = \\u2_adr0_cnt_reg[18] ;
  assign \new_[1376]_  = \\u2_adr0_cnt_reg[10] ;
  assign \new_[1377]_  = \\u2_adr0_cnt_reg[11] ;
  assign \new_[1378]_  = \\u2_adr0_cnt_reg[12] ;
  assign \new_[1379]_  = \\u2_adr0_cnt_reg[13] ;
  assign \new_[1380]_  = \\u2_adr0_cnt_reg[17] ;
  assign \new_[1381]_  = \\u2_adr0_cnt_reg[21] ;
  assign \new_[1382]_  = \\u2_adr0_cnt_reg[25] ;
  assign \new_[1383]_  = \\u2_adr0_cnt_reg[2] ;
  assign \new_[1384]_  = \\u2_adr0_cnt_reg[3] ;
  assign \new_[1385]_  = ~\\u2_adr0_cnt_reg[5] ;
  assign \new_[1386]_  = ~\\u2_adr0_cnt_reg[6] ;
  assign \new_[1387]_  = \\u2_adr0_cnt_reg[8] ;
  assign \new_[1388]_  = \\u2_adr0_cnt_reg[7] ;
  assign \new_[1389]_  = \\u2_adr0_cnt_reg[4] ;
  assign \new_[1390]_  = ~\\u0_u0_ch_csr_r_reg[0] ;
  assign \wb0s_data_o[11]  = \wb1m_data_i[11]  ? \new_[3659]_  : \new_[1504]_ ;
  assign \wb0s_data_o[10]  = \wb1m_data_i[10]  ? \new_[3659]_  : \new_[1505]_ ;
  assign \wb0s_data_o[9]  = \wb1m_data_i[9]  ? \new_[3659]_  : \new_[1506]_ ;
  assign \wb0s_data_o[8]  = \wb1m_data_i[8]  ? \new_[3574]_  : \new_[1508]_ ;
  assign \wb0s_data_o[7]  = \wb1m_data_i[7]  ? \new_[3574]_  : \new_[1509]_ ;
  assign \wb0s_data_o[6]  = \wb1m_data_i[6]  ? \new_[3659]_  : \new_[1510]_ ;
  assign \wb0s_data_o[5]  = \wb1m_data_i[5]  ? \new_[3659]_  : \new_[1511]_ ;
  assign \wb0s_data_o[4]  = \wb1m_data_i[4]  ? \new_[3659]_  : \new_[1512]_ ;
  assign \wb0s_data_o[3]  = \wb1m_data_i[3]  ? \new_[3659]_  : \new_[1500]_ ;
  assign \wb0s_data_o[2]  = \wb1m_data_i[2]  ? \new_[3659]_  : \new_[1501]_ ;
  assign \wb0s_data_o[1]  = \wb1m_data_i[1]  ? \new_[3574]_  : \new_[1502]_ ;
  assign \wb0s_data_o[0]  = \wb1m_data_i[0]  ? \new_[3659]_  : \new_[1503]_ ;
  assign \new_[1403]_  = ~\new_[1436]_  & (~\new_[1493]_  | ~\new_[1231]_ );
  assign \new_[1404]_  = ~\new_[1437]_  & (~\new_[4293]_  | ~\new_[3994]_ );
  assign \new_[1405]_  = ~\new_[1975]_  | (~\new_[2371]_  & ~\new_[1516]_ );
  assign \new_[1406]_  = \\u2_adr0_cnt_reg[14] ;
  assign \new_[1407]_  = ~\new_[1495]_  | (~\new_[1587]_  & ~\new_[1518]_ );
  assign n1386 = ~\new_[4206]_  & ~\new_[1490]_ ;
  assign n1381 = ~\new_[1440]_ ;
  assign n1376 = ~\new_[1491]_  | ~\new_[2792]_ ;
  assign \new_[1411]_  = ~\new_[1494]_  & (~\new_[4293]_  | ~\new_[1287]_ );
  assign \new_[1412]_  = ~\new_[1496]_  & (~\new_[4293]_  | ~\new_[1284]_ );
  assign \new_[1413]_  = \\u2_adr0_cnt_reg[22] ;
  assign \new_[1414]_  = \\u2_adr0_cnt_reg[19] ;
  assign \new_[1415]_  = ~\\u2_adr0_cnt_reg[29] ;
  assign \new_[1416]_  = ~\\u2_adr0_cnt_reg[15] ;
  assign \new_[1417]_  = u0_u0_ch_done_reg;
  assign \wb0s_data_o[30]  = ~\new_[3441]_  | (~\new_[2089]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[29]  = ~\new_[3446]_  | (~\new_[2090]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[28]  = ~\new_[3449]_  | (~\new_[2091]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[27]  = ~\new_[3476]_  | (~\new_[2093]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[26]  = ~\new_[3502]_  | (~\new_[2074]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[25]  = ~\new_[3450]_  | (~\new_[2075]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[24]  = ~\new_[3440]_  | (~\new_[2076]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[23]  = ~\new_[3438]_  | (~\new_[2077]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[22]  = ~\new_[3448]_  | (~\new_[2078]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[21]  = ~\new_[3447]_  | (~\new_[2079]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[19]  = ~\new_[3511]_  | (~\new_[2081]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[18]  = ~\new_[3512]_  | (~\new_[2082]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[17]  = ~\new_[3505]_  | (~\new_[2083]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[14]  = ~\new_[3442]_  | (~\new_[2086]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[16]  = ~\new_[3443]_  | (~\new_[2084]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[15]  = ~\new_[3439]_  | (~\new_[2085]_  & ~\new_[1551]_ );
  assign \new_[1434]_  = ~\new_[1507]_  & (~\new_[1517]_  | ~\new_[1285]_ );
  assign n1371 = ~\new_[1899]_  | ~\new_[1488]_ ;
  assign \new_[1436]_  = ~\new_[1598]_  & ~\new_[1519]_ ;
  assign \new_[1437]_  = ~\new_[1519]_  & (~\new_[1605]_  | ~\new_[1609]_ );
  assign n1411 = ~\new_[1906]_  | (~\new_[1543]_  & ~\new_[4288]_ );
  assign \new_[1439]_  = ~\new_[1519]_  & (~\new_[1713]_  | ~\new_[1681]_ );
  assign \new_[1440]_  = ~\new_[2604]_  | ~\new_[4210]_  | ~\new_[2670]_  | ~n1536;
  assign n1396 = ~\new_[1911]_  | (~\new_[1548]_  & ~\new_[4288]_ );
  assign n1426 = ~\new_[1901]_  | (~\new_[1549]_  & ~\new_[4288]_ );
  assign \new_[1443]_  = \new_[3749]_  ? \new_[4293]_  : \new_[3997]_ ;
  assign \new_[1444]_  = ~\new_[1601]_  & ~\new_[1519]_ ;
  assign \new_[1445]_  = \new_[3590]_  ? \new_[4293]_  : \new_[4066]_ ;
  assign n1501 = ~\new_[2797]_  | ~\new_[1521]_ ;
  assign \new_[1447]_  = ~\new_[1519]_  & (~\new_[1707]_  | ~\new_[1608]_ );
  assign \new_[1448]_  = ~\new_[1519]_  & (~\new_[1685]_  | ~\new_[4355]_ );
  assign \new_[1449]_  = ~\new_[1519]_  & (~\new_[1686]_  | ~\new_[1610]_ );
  assign \new_[1450]_  = ~\new_[1519]_  & (~\new_[1687]_  | ~\new_[1611]_ );
  assign \new_[1451]_  = ~\new_[1519]_  & (~\new_[1688]_  | ~\new_[1612]_ );
  assign \new_[1452]_  = ~\new_[1519]_  & (~\new_[1689]_  | ~\new_[1613]_ );
  assign \new_[1453]_  = ~\new_[1519]_  & (~\new_[1690]_  | ~\new_[1614]_ );
  assign \new_[1454]_  = ~\new_[1519]_  & (~\new_[1637]_  | ~\new_[1615]_ );
  assign \new_[1455]_  = ~\new_[1519]_  & (~\new_[1638]_  | ~\new_[1616]_ );
  assign \new_[1456]_  = ~\new_[1519]_  & (~\new_[1715]_  | ~\new_[1635]_ );
  assign n1421 = ~\new_[1903]_  | (~\new_[1547]_  & ~\new_[2246]_ );
  assign \new_[1458]_  = ~\new_[1519]_  & (~\new_[1716]_  | ~\new_[1675]_ );
  assign \new_[1459]_  = ~\new_[1519]_  & (~\new_[1645]_  | ~\new_[1677]_ );
  assign \new_[1460]_  = ~\new_[1519]_  & (~\new_[1717]_  | ~\new_[1678]_ );
  assign \new_[1461]_  = ~\new_[1519]_  & (~\new_[1718]_  | ~\new_[1679]_ );
  assign \new_[1462]_  = ~\new_[1640]_  & ~\new_[1519]_ ;
  assign n1401 = ~\new_[1910]_  | (~\new_[1523]_  & ~\new_[4288]_ );
  assign \new_[1464]_  = ~\new_[1519]_  & (~\new_[1596]_  | ~\new_[1680]_ );
  assign \new_[1465]_  = ~\new_[1519]_  & (~\new_[1656]_  | ~\new_[1682]_ );
  assign \wb0s_data_o[31]  = ~\new_[3445]_  | (~\new_[2092]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[20]  = ~\new_[3421]_  | (~\new_[2080]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[12]  = ~\new_[3444]_  | (~\new_[2088]_  & ~\new_[1551]_ );
  assign \wb0s_data_o[13]  = ~\new_[3503]_  | (~\new_[2087]_  & ~\new_[1551]_ );
  assign \new_[1470]_  = ~\new_[1519]_  & (~\new_[1723]_  | ~\new_[1684]_ );
  assign \new_[1471]_  = ~\new_[1651]_  & ~\new_[1519]_ ;
  assign n1431 = ~\new_[1851]_  | (~\new_[1524]_  & ~\new_[4288]_ );
  assign n1436 = ~\new_[1881]_  | (~\new_[1525]_  & ~\new_[4308]_ );
  assign n1441 = ~\new_[1896]_  | (~\new_[1526]_  & ~\new_[4288]_ );
  assign n1451 = ~\new_[1900]_  | (~\new_[1528]_  & ~\new_[4288]_ );
  assign n1456 = ~\new_[1904]_  | (~\new_[1529]_  & ~\new_[4288]_ );
  assign n1461 = ~\new_[1908]_  | (~\new_[1530]_  & ~\new_[4288]_ );
  assign n1416 = ~\new_[1909]_  | (~\new_[1537]_  & ~\new_[2243]_ );
  assign n1466 = ~\new_[1912]_  | (~\new_[1531]_  & ~\new_[4288]_ );
  assign n1471 = ~\new_[1915]_  | (~\new_[1533]_  & ~\new_[2244]_ );
  assign n1496 = ~\new_[1924]_  | (~\new_[1535]_  & ~\new_[2246]_ );
  assign n1476 = ~\new_[1931]_  | (~\new_[1536]_  & ~\new_[2246]_ );
  assign n1481 = ~\new_[1939]_  | (~\new_[1538]_  & ~\new_[2244]_ );
  assign n1491 = ~\new_[1941]_  | (~\new_[1539]_  & ~\new_[2244]_ );
  assign n1486 = ~\new_[1943]_  | (~\new_[1540]_  & ~\new_[4288]_ );
  assign n1391 = ~\new_[1944]_  | (~\new_[1541]_  & ~\new_[4288]_ );
  assign n1406 = ~\new_[1907]_  | (~\new_[1542]_  & ~\new_[4308]_ );
  assign \new_[1488]_  = ~\new_[1527]_  | ~\new_[2186]_ ;
  assign n1511 = ~\new_[1905]_  | (~\new_[1556]_  & ~\new_[4288]_ );
  assign \new_[1490]_  = ~u2_next_ch_reg;
  assign \new_[1491]_  = ~n1536 | ~\new_[2514]_ ;
  assign \new_[1492]_  = ~\new_[1532]_  & (~\new_[2368]_  | ~\new_[3907]_ );
  assign \new_[1493]_  = ~\new_[4296]_  | ~\new_[4186]_ ;
  assign \new_[1494]_  = ~\new_[4293]_  & (~\new_[1663]_  | ~\new_[1676]_ );
  assign \new_[1495]_  = ~\new_[4293]_  | ~\new_[1238]_ ;
  assign \new_[1496]_  = ~\new_[4293]_  & (~\new_[1647]_  | ~\new_[1665]_ );
  assign n1521 = ~\new_[1522]_ ;
  assign \new_[1498]_  = ~\\u0_u0_int_src_r_reg[1] ;
  assign \new_[1499]_  = \\u2_state_reg[0] ;
  assign \new_[1500]_  = \new_[2358]_  ? \new_[1551]_  : \new_[1701]_ ;
  assign \new_[1501]_  = \new_[2359]_  ? \new_[1551]_  : \new_[1659]_ ;
  assign \new_[1502]_  = \new_[2360]_  ? \new_[1551]_  : \new_[1700]_ ;
  assign \new_[1503]_  = \new_[2361]_  ? \new_[1551]_  : \new_[1693]_ ;
  assign \new_[1504]_  = \new_[2362]_  ? \new_[1551]_  : \new_[1699]_ ;
  assign \new_[1505]_  = \new_[2363]_  ? \new_[1551]_  : \new_[1698]_ ;
  assign \new_[1506]_  = \new_[2364]_  ? \new_[1551]_  : \new_[1702]_ ;
  assign \new_[1507]_  = ~\new_[4293]_  & (~\new_[1654]_  | ~\new_[1683]_ );
  assign \new_[1508]_  = \new_[2365]_  ? \new_[1551]_  : \new_[1657]_ ;
  assign \new_[1509]_  = \new_[2366]_  ? \new_[1551]_  : \new_[1697]_ ;
  assign \new_[1510]_  = \new_[2367]_  ? \new_[1551]_  : \new_[1696]_ ;
  assign \new_[1511]_  = \new_[2369]_  ? \new_[1551]_  : \new_[1695]_ ;
  assign \new_[1512]_  = \new_[2370]_  ? \new_[1551]_  : \new_[1694]_ ;
  assign n1516 = ~\new_[1902]_  | (~\new_[1550]_  & ~\new_[4288]_ );
  assign n1506 = ~\new_[1897]_  | (~\new_[1552]_  & ~\new_[4308]_ );
  assign n1526 = ~\new_[1898]_  | (~\new_[1554]_  & ~\new_[4288]_ );
  assign \new_[1516]_  = ~\new_[1553]_  & (~\new_[2368]_  | ~\new_[3909]_ );
  assign \new_[1517]_  = ~\new_[4296]_ ;
  assign \new_[1518]_  = ~\new_[4296]_ ;
  assign \new_[1519]_  = ~\new_[4296]_ ;
  assign \new_[1520]_  = ~\new_[4251]_  | ~\new_[2849]_ ;
  assign \new_[1521]_  = ~\new_[3966]_  | ~\new_[2873]_  | ~\new_[1580]_ ;
  assign \new_[1522]_  = (~\new_[1559]_  | ~\new_[2186]_ ) & (~\new_[3981]_  | ~\new_[2064]_ );
  assign \new_[1523]_  = ~\new_[1561]_  & (~\new_[2038]_  | ~\new_[1370]_ );
  assign \new_[1524]_  = ~\new_[1563]_  & (~\new_[2035]_  | ~\new_[1376]_ );
  assign \new_[1525]_  = ~\new_[1564]_  & (~\new_[2035]_  | ~\new_[1377]_ );
  assign \new_[1526]_  = ~\new_[1565]_  & (~\new_[2035]_  | ~\new_[1378]_ );
  assign \new_[1527]_  = ~\new_[1855]_  | (~\new_[1586]_  & ~\new_[2038]_ );
  assign \new_[1528]_  = ~\new_[1567]_  & (~\new_[2035]_  | ~\new_[1380]_ );
  assign \new_[1529]_  = ~\new_[1568]_  & (~\new_[2035]_  | ~\new_[1381]_ );
  assign \new_[1530]_  = ~\new_[1569]_  & (~\new_[2038]_  | ~\new_[1382]_ );
  assign \new_[1531]_  = ~\new_[1570]_  & (~\new_[2035]_  | ~\new_[1383]_ );
  assign \new_[1532]_  = ~\new_[2368]_  & ~\new_[1562]_ ;
  assign \new_[1533]_  = ~\new_[1571]_  & (~\new_[2035]_  | ~\new_[1384]_ );
  assign n1536 = ~\new_[1562]_  & ~\new_[4242]_ ;
  assign \new_[1535]_  = ~\new_[1572]_  & (~\new_[2035]_  | ~\new_[1389]_ );
  assign \new_[1536]_  = ~\new_[1573]_  & (~\new_[2035]_  | ~\new_[4082]_ );
  assign \new_[1537]_  = ~\new_[1578]_  & (~\new_[2035]_  | ~\new_[1373]_ );
  assign \new_[1538]_  = ~\new_[1574]_  & (~\new_[2035]_  | ~\new_[4185]_ );
  assign \new_[1539]_  = ~\new_[1575]_  & (~\new_[2035]_  | ~\new_[1388]_ );
  assign \new_[1540]_  = ~\new_[1576]_  & (~\new_[2035]_  | ~\new_[1387]_ );
  assign \new_[1541]_  = ~\new_[1577]_  & (~\new_[2035]_  | ~\new_[1345]_ );
  assign \new_[1542]_  = ~\new_[1566]_  & (~\new_[2035]_  | ~\new_[1371]_ );
  assign \new_[1543]_  = ~\new_[1579]_  & (~\new_[2035]_  | ~\new_[1372]_ );
  assign n1546 = ~\new_[1584]_  | ~\new_[1854]_  | ~\new_[3211]_ ;
  assign n1531 = ~\new_[1580]_  | ~\new_[4173]_ ;
  assign n1541 = ~\new_[2791]_  | ~\new_[1580]_ ;
  assign \new_[1547]_  = ~\new_[1581]_  & (~\new_[2035]_  | ~\new_[3935]_ );
  assign \new_[1548]_  = ~\new_[1557]_  & (~\new_[2035]_  | ~\new_[4011]_ );
  assign \new_[1549]_  = ~\new_[1558]_  & (~\new_[2035]_  | ~\new_[1375]_ );
  assign \new_[1550]_  = ~\new_[1585]_  & (~\new_[2035]_  | ~\new_[1414]_ );
  assign \new_[1551]_  = ~\new_[1560]_ ;
  assign \new_[1552]_  = ~\new_[1589]_  & (~\new_[2035]_  | ~\new_[1406]_ );
  assign \new_[1553]_  = ~\new_[2425]_  & ~\new_[1588]_ ;
  assign \new_[1554]_  = ~\new_[1590]_  & (~\new_[2035]_  | ~\new_[4070]_ );
  assign \new_[1555]_  = \\u2_state_reg[9] ;
  assign \new_[1556]_  = ~\new_[1593]_  & (~\new_[2035]_  | ~\new_[1413]_ );
  assign \new_[1557]_  = ~\new_[2035]_  & (~\new_[1606]_  | ~\new_[1626]_ );
  assign \new_[1558]_  = ~\new_[2035]_  & (~\new_[1661]_  | ~\new_[1621]_ );
  assign \new_[1559]_  = \new_[2171]_  ? \new_[1600]_  : \new_[3992]_ ;
  assign \new_[1560]_  = ~\new_[1583]_ ;
  assign \new_[1561]_  = ~\new_[2037]_  & (~\new_[1714]_  | ~\new_[1625]_ );
  assign \new_[1562]_  = ~\new_[1588]_ ;
  assign \new_[1563]_  = ~\new_[2035]_  & (~\new_[1703]_  | ~\new_[1617]_ );
  assign \new_[1564]_  = ~\new_[2037]_  & (~\new_[1704]_  | ~\new_[1618]_ );
  assign \new_[1565]_  = ~\new_[2035]_  & (~\new_[1603]_  | ~\new_[1666]_ );
  assign \new_[1566]_  = ~\new_[2023]_  & (~\new_[1722]_  | ~\new_[1623]_ );
  assign \new_[1567]_  = ~\new_[2036]_  & (~\new_[1655]_  | ~\new_[1620]_ );
  assign \new_[1568]_  = ~\new_[2036]_  & (~\new_[1597]_  | ~\new_[1671]_ );
  assign \new_[1569]_  = ~\new_[2035]_  & (~\new_[1649]_  | ~\new_[1624]_ );
  assign \new_[1570]_  = ~\new_[2035]_  & (~\new_[1708]_  | ~\new_[1627]_ );
  assign \new_[1571]_  = ~\new_[2037]_  & (~\new_[1709]_  | ~\new_[1628]_ );
  assign \new_[1572]_  = ~\new_[2035]_  & (~\new_[1710]_  | ~\new_[1629]_ );
  assign \new_[1573]_  = ~\new_[2038]_  & (~\new_[1711]_  | ~\new_[1630]_ );
  assign \new_[1574]_  = ~\new_[2037]_  & (~\new_[1641]_  | ~\new_[1631]_ );
  assign \new_[1575]_  = ~\new_[2036]_  & (~\new_[1642]_  | ~\new_[1632]_ );
  assign \new_[1576]_  = ~\new_[2023]_  & (~\new_[1643]_  | ~\new_[1633]_ );
  assign \new_[1577]_  = ~\new_[2023]_  & (~\new_[1644]_  | ~\new_[1634]_ );
  assign \new_[1578]_  = ~\new_[2035]_  & (~\new_[1650]_  | ~\new_[1674]_ );
  assign \new_[1579]_  = ~\new_[2036]_  & (~\new_[1652]_  | ~\new_[1673]_ );
  assign \new_[1580]_  = (~\new_[2407]_  | ~\new_[1599]_ ) & (~\new_[3950]_  | ~\new_[3728]_ );
  assign \new_[1581]_  = ~\new_[2035]_  & (~\new_[1658]_  | ~\new_[1622]_ );
  assign n1551 = ~\new_[3022]_  | (~\new_[1660]_  & ~\new_[3234]_ );
  assign \new_[1583]_  = ~\new_[3254]_  | (~\new_[1660]_  & ~\new_[4242]_ );
  assign \new_[1584]_  = ~\new_[3179]_  & (~\new_[1660]_  | ~\new_[3182]_ );
  assign \new_[1585]_  = ~\new_[2023]_  & (~\new_[1712]_  | ~\new_[1670]_ );
  assign \new_[1586]_  = ~\new_[1619]_  & (~\new_[2631]_  | ~\new_[4186]_ );
  assign \new_[1587]_  = ~\new_[1636]_  & (~\new_[4191]_  | ~\new_[2647]_ );
  assign \new_[1588]_  = ~\new_[1602]_  | ~\new_[2518]_ ;
  assign \new_[1589]_  = ~\new_[2035]_  & (~\new_[1705]_  | ~\new_[1668]_ );
  assign \new_[1590]_  = ~\new_[2035]_  & (~\new_[1706]_  | ~\new_[1669]_ );
  assign n3466 = ~\\u2_adr0_cnt_reg[0] ;
  assign \new_[1592]_  = ~\\u2_adr0_cnt_reg[1] ;
  assign \new_[1593]_  = ~\new_[2035]_  & (~\new_[1653]_  | ~\new_[1672]_ );
  assign \wb0m_data_o[10]  = \wb1s_data_i[10]  ? \new_[3606]_  : \new_[1664]_ ;
  assign wb1_we_o = wb0_we_i ? \new_[3592]_  : \new_[1662]_ ;
  assign \new_[1596]_  = ~\new_[4186]_  | ~\new_[2561]_ ;
  assign \new_[1597]_  = ~\new_[4198]_  | ~\new_[2396]_ ;
  assign \new_[1598]_  = ~\new_[4188]_  | ~\new_[2198]_ ;
  assign \new_[1599]_  = ~\new_[3837]_  & (~\new_[1738]_  | ~\new_[2416]_ );
  assign \new_[1600]_  = ~\new_[4306]_  | ~\new_[4186]_ ;
  assign \new_[1601]_  = ~\new_[4188]_  | ~\new_[2515]_ ;
  assign \new_[1602]_  = ~n2861 | ~\new_[1724]_ ;
  assign \new_[1603]_  = ~\new_[4198]_  | ~\new_[2756]_ ;
  assign \new_[1604]_  = \new_[1725]_  & \new_[2514]_ ;
  assign \new_[1605]_  = ~\new_[4186]_  | ~\new_[1785]_ ;
  assign \new_[1606]_  = ~\new_[4186]_  | ~\new_[1730]_ ;
  assign \new_[1607]_  = ~\new_[4195]_  | ~\new_[1234]_ ;
  assign \new_[1608]_  = ~\new_[4190]_  | ~\new_[1228]_ ;
  assign \new_[1609]_  = ~\new_[4194]_  | ~\new_[3994]_ ;
  assign \new_[1610]_  = ~\new_[4194]_  | ~\new_[1240]_ ;
  assign \new_[1611]_  = ~\new_[4194]_  | ~\new_[1241]_ ;
  assign \new_[1612]_  = ~\new_[4195]_  | ~\new_[4154]_ ;
  assign \new_[1613]_  = ~\new_[4189]_  | ~\new_[3989]_ ;
  assign \new_[1614]_  = ~\new_[4195]_  | ~\new_[1244]_ ;
  assign \new_[1615]_  = ~\new_[4194]_  | ~\new_[1245]_ ;
  assign \new_[1616]_  = ~\new_[4194]_  | ~\new_[1246]_ ;
  assign \new_[1617]_  = ~\new_[4195]_  | ~\new_[1376]_ ;
  assign \new_[1618]_  = ~\new_[4194]_  | ~\new_[1377]_ ;
  assign \new_[1619]_  = ~\new_[4191]_  & ~\new_[4139]_ ;
  assign \new_[1620]_  = ~\new_[4195]_  | ~\new_[1380]_ ;
  assign \new_[1621]_  = ~\new_[4194]_  | ~\new_[1375]_ ;
  assign \new_[1622]_  = ~\new_[4189]_  | ~\new_[3935]_ ;
  assign \new_[1623]_  = ~\new_[4194]_  | ~\new_[1371]_ ;
  assign \new_[1624]_  = ~\new_[4195]_  | ~\new_[1382]_ ;
  assign \new_[1625]_  = ~\new_[4195]_  | ~\new_[1370]_ ;
  assign \new_[1626]_  = ~\new_[4194]_  | ~\new_[4011]_ ;
  assign \new_[1627]_  = ~\new_[4195]_  | ~\new_[1383]_ ;
  assign \new_[1628]_  = ~\new_[4190]_  | ~\new_[1384]_ ;
  assign \new_[1629]_  = ~\new_[4190]_  | ~\new_[1389]_ ;
  assign \new_[1630]_  = ~\new_[4190]_  | ~\new_[4082]_ ;
  assign \new_[1631]_  = ~\new_[4189]_  | ~\new_[4185]_ ;
  assign \new_[1632]_  = ~\new_[4194]_  | ~\new_[1388]_ ;
  assign \new_[1633]_  = ~\new_[4195]_  | ~\new_[1387]_ ;
  assign \new_[1634]_  = ~\new_[4195]_  | ~\new_[1345]_ ;
  assign \new_[1635]_  = ~\new_[4189]_  | ~\new_[1247]_ ;
  assign \new_[1636]_  = ~\new_[4191]_  & ~\new_[4068]_ ;
  assign \new_[1637]_  = ~\new_[4186]_  | ~\new_[2847]_ ;
  assign \new_[1638]_  = ~\new_[4186]_  | ~\new_[3290]_ ;
  assign \new_[1639]_  = ~\new_[4186]_  | ~\new_[3023]_ ;
  assign \new_[1640]_  = ~\new_[4191]_  | ~\new_[2381]_ ;
  assign \new_[1641]_  = ~\new_[4197]_  | ~\new_[3285]_ ;
  assign \new_[1642]_  = ~\new_[4197]_  | ~\new_[2923]_ ;
  assign \new_[1643]_  = ~\new_[4186]_  | ~\new_[2848]_ ;
  assign \new_[1644]_  = ~\new_[4198]_  | ~\new_[3291]_ ;
  assign \new_[1645]_  = ~\new_[4186]_  | ~\new_[3024]_ ;
  assign n1556 = ~\new_[1719]_ ;
  assign \new_[1647]_  = ~\new_[4186]_  | ~\new_[1971]_ ;
  assign n1561 = ~\new_[1720]_ ;
  assign \new_[1649]_  = ~\new_[4186]_  | ~\new_[2199]_ ;
  assign \new_[1650]_  = ~\new_[4197]_  | ~\new_[1836]_ ;
  assign \new_[1651]_  = ~\new_[4191]_  | ~\new_[1972]_ ;
  assign \new_[1652]_  = ~\new_[4198]_  | ~\new_[2022]_ ;
  assign \new_[1653]_  = ~\new_[4186]_  | ~\new_[2025]_ ;
  assign \new_[1654]_  = ~\new_[4197]_  | ~\new_[2096]_ ;
  assign \new_[1655]_  = ~\new_[4198]_  | ~\new_[2421]_ ;
  assign \new_[1656]_  = ~\new_[4198]_  | ~\new_[2519]_ ;
  assign \new_[1657]_  = \\u2_tsz_cnt_reg[8] ;
  assign \new_[1658]_  = ~\new_[4197]_  | ~\new_[2140]_ ;
  assign \new_[1659]_  = \\u2_tsz_cnt_reg[2] ;
  assign \new_[1660]_  = \new_[4253]_ ;
  assign \new_[1661]_  = ~\new_[4198]_  | ~\new_[2433]_ ;
  assign \new_[1662]_  = u4_u0_mast_we_r_reg;
  assign \new_[1663]_  = ~\new_[4186]_  | ~\new_[2757]_ ;
  assign \new_[1664]_  = \\u0_wb_rf_dout_reg[10] ;
  assign \new_[1665]_  = ~\new_[4187]_  | ~\new_[1284]_ ;
  assign \new_[1666]_  = ~\new_[4187]_  | ~\new_[1378]_ ;
  assign \new_[1667]_  = ~\new_[4195]_  | ~\new_[1379]_ ;
  assign \new_[1668]_  = ~\new_[4194]_  | ~\new_[1406]_ ;
  assign \new_[1669]_  = ~\new_[4195]_  | ~\new_[4070]_ ;
  assign \new_[1670]_  = ~\new_[4187]_  | ~\new_[1414]_ ;
  assign \new_[1671]_  = ~\new_[4195]_  | ~\new_[1381]_ ;
  assign \new_[1672]_  = ~\new_[4195]_  | ~\new_[1413]_ ;
  assign \new_[1673]_  = ~\new_[4195]_  | ~\new_[1372]_ ;
  assign \new_[1674]_  = ~\new_[4194]_  | ~\new_[1373]_ ;
  assign \new_[1675]_  = ~\new_[4187]_  | ~\new_[1248]_ ;
  assign \new_[1676]_  = ~\new_[4194]_  | ~\new_[1287]_ ;
  assign \new_[1677]_  = ~\new_[4192]_  | ~\new_[1249]_ ;
  assign \new_[1678]_  = ~\new_[4194]_  | ~\new_[1250]_ ;
  assign \new_[1679]_  = ~\new_[4195]_  | ~\new_[4080]_ ;
  assign \new_[1680]_  = ~\new_[4187]_  | ~\new_[1236]_ ;
  assign \new_[1681]_  = ~\new_[4187]_  | ~\new_[1232]_ ;
  assign \new_[1682]_  = ~\new_[4187]_  | ~\new_[1237]_ ;
  assign \new_[1683]_  = ~\new_[4194]_  | ~\new_[1285]_ ;
  assign \new_[1684]_  = ~\new_[4187]_  | ~\new_[1229]_ ;
  assign \new_[1685]_  = ~\new_[4197]_  | ~\new_[3413]_ ;
  assign \new_[1686]_  = ~\new_[4198]_  | ~\new_[3271]_ ;
  assign \new_[1687]_  = ~\new_[4197]_  | ~\new_[3091]_ ;
  assign \new_[1688]_  = ~\new_[4186]_  | ~\new_[3401]_ ;
  assign \new_[1689]_  = ~\new_[4197]_  | ~\new_[3284]_ ;
  assign \new_[1690]_  = ~\new_[4198]_  | ~\new_[2922]_ ;
  assign \new_[1691]_  = \\u2_state_reg[10] ;
  assign \new_[1692]_  = \\u2_state_reg[4] ;
  assign \new_[1693]_  = \\u2_tsz_cnt_reg[0] ;
  assign \new_[1694]_  = \\u2_tsz_cnt_reg[4] ;
  assign \new_[1695]_  = \\u2_tsz_cnt_reg[5] ;
  assign \new_[1696]_  = \\u2_tsz_cnt_reg[6] ;
  assign \new_[1697]_  = \\u2_tsz_cnt_reg[7] ;
  assign \new_[1698]_  = \\u2_tsz_cnt_reg[10] ;
  assign \new_[1699]_  = \\u2_tsz_cnt_reg[11] ;
  assign \new_[1700]_  = \\u2_tsz_cnt_reg[1] ;
  assign \new_[1701]_  = \\u2_tsz_cnt_reg[3] ;
  assign \new_[1702]_  = \\u2_tsz_cnt_reg[9] ;
  assign \new_[1703]_  = ~\new_[4198]_  | ~\new_[3099]_ ;
  assign \new_[1704]_  = ~\new_[4197]_  | ~\new_[2754]_ ;
  assign \new_[1705]_  = ~\new_[4186]_  | ~\new_[2839]_ ;
  assign \new_[1706]_  = ~\new_[4186]_  | ~\new_[2671]_ ;
  assign \new_[1707]_  = ~\new_[4197]_  | ~\new_[1966]_ ;
  assign \new_[1708]_  = ~\new_[4198]_  | ~\new_[3420]_ ;
  assign \new_[1709]_  = ~\new_[4197]_  | ~\new_[3278]_ ;
  assign \new_[1710]_  = ~\new_[4197]_  | ~\new_[3092]_ ;
  assign \new_[1711]_  = ~\new_[4197]_  | ~\new_[3338]_ ;
  assign \new_[1712]_  = ~\new_[4198]_  | ~\new_[2357]_ ;
  assign \new_[1713]_  = ~\new_[4198]_  | ~\new_[2400]_ ;
  assign \new_[1714]_  = ~\new_[4186]_  | ~\new_[1808]_ ;
  assign \new_[1715]_  = ~\new_[4197]_  | ~\new_[3098]_ ;
  assign \new_[1716]_  = ~\new_[4198]_  | ~\new_[2755]_ ;
  assign \new_[1717]_  = ~\new_[4197]_  | ~\new_[2840]_ ;
  assign \new_[1718]_  = ~\new_[4186]_  | ~\new_[2672]_ ;
  assign \new_[1719]_  = (~\new_[1790]_  | ~\new_[2186]_ ) & (~\new_[3961]_  | ~\new_[2064]_ );
  assign \new_[1720]_  = (~\new_[1791]_  | ~\new_[2186]_ ) & (~\new_[4032]_  | ~\new_[2064]_ );
  assign \new_[1721]_  = ~\new_[4198]_  | ~\new_[2395]_ ;
  assign \new_[1722]_  = ~\new_[4197]_  | ~\new_[1842]_ ;
  assign \new_[1723]_  = ~\new_[4198]_  | ~\new_[2095]_ ;
  assign \new_[1724]_  = ~u2_chunk_0_reg;
  assign \new_[1725]_  = u2_write_r_reg;
  assign \new_[1726]_  = ~n1366;
  assign \new_[1727]_  = \\u2_state_reg[2] ;
  assign \new_[1728]_  = ~\\u0_u0_ch_tot_sz_r_reg[0] ;
  assign \new_[1729]_  = ~n1576;
  assign \new_[1730]_  = ~\new_[1807]_  | (~\new_[1970]_  & ~\new_[4011]_ );
  assign \new_[1731]_  = ~\\u0_u0_ch_adr1_r_reg[25] ;
  assign \new_[1732]_  = ~\\u0_u0_ch_adr0_r_reg[17] ;
  assign \new_[1733]_  = ~\\u0_u0_ch_adr0_r_reg[13] ;
  assign \new_[1734]_  = ~\\u0_u0_ch_adr1_r_reg[29] ;
  assign \new_[1735]_  = ~\\u0_u0_ch_adr1_r_reg[21] ;
  assign \new_[1736]_  = ~\\u0_u0_ch_adr1_r_reg[13] ;
  assign \new_[1737]_  = ~\\u0_u0_ch_adr1_r_reg[17] ;
  assign \new_[1738]_  = ~\new_[4217]_  | ~n2861;
  assign n1586 = ~\new_[1974]_  | ~\new_[3016]_  | ~\new_[2850]_ ;
  assign n1591 = ~\new_[2846]_  | (~\new_[1983]_  & ~\new_[3100]_ );
  assign n1621 = ~\new_[1868]_  | (~\new_[2919]_  & ~\new_[2242]_ );
  assign n1626 = ~\new_[1869]_  | (~\new_[2762]_  & ~\new_[4308]_ );
  assign n1631 = ~\new_[1870]_  | (~\new_[3437]_  & ~\new_[2242]_ );
  assign n1636 = ~\new_[1872]_  | (~\new_[3330]_  & ~\new_[4308]_ );
  assign n1641 = ~\new_[1875]_  | (~\new_[3031]_  & ~\new_[4308]_ );
  assign n1606 = ~\new_[1873]_  | (~\new_[3057]_  & ~\new_[2242]_ );
  assign n1611 = ~\new_[1852]_  | (~\new_[2953]_  & ~\new_[2242]_ );
  assign n1616 = ~\new_[1874]_  | (~\new_[2918]_  & ~\new_[2242]_ );
  assign n1596 = ~\new_[1793]_ ;
  assign n1601 = ~\new_[1794]_ ;
  assign n1566 = ~\new_[1795]_ ;
  assign n1366 = ~\new_[1961]_  & ~\new_[2586]_ ;
  assign \new_[1753]_  = ~\\u0_u0_ch_tot_sz_r_reg[1] ;
  assign \new_[1754]_  = ~\\u0_u0_ch_adr1_r_reg[10] ;
  assign \new_[1755]_  = ~\\u0_u0_ch_adr1_r_reg[11] ;
  assign \new_[1756]_  = ~\\u0_u0_ch_adr1_r_reg[12] ;
  assign n1576 = ~\new_[1961]_  & ~\new_[2568]_ ;
  assign \new_[1758]_  = ~\\u0_u0_ch_adr1_r_reg[14] ;
  assign \new_[1759]_  = ~\\u0_u0_ch_adr1_r_reg[15] ;
  assign \new_[1760]_  = ~\\u0_u0_ch_adr1_r_reg[16] ;
  assign \new_[1761]_  = ~\\u0_u0_ch_adr1_r_reg[18] ;
  assign \new_[1762]_  = ~\\u0_u0_ch_adr1_r_reg[19] ;
  assign \new_[1763]_  = ~\\u0_u0_ch_adr1_r_reg[20] ;
  assign \new_[1764]_  = ~\\u0_u0_ch_adr1_r_reg[22] ;
  assign \new_[1765]_  = ~\\u0_u0_ch_adr1_r_reg[23] ;
  assign \new_[1766]_  = ~\\u0_u0_ch_adr1_r_reg[24] ;
  assign \new_[1767]_  = ~\\u0_u0_ch_adr1_r_reg[26] ;
  assign \new_[1768]_  = ~\\u0_u0_ch_adr1_r_reg[27] ;
  assign \new_[1769]_  = ~\\u0_u0_ch_adr1_r_reg[28] ;
  assign \new_[1770]_  = ~\\u0_u0_ch_adr0_r_reg[10] ;
  assign \new_[1771]_  = ~\\u0_u0_ch_adr0_r_reg[11] ;
  assign \new_[1772]_  = ~\\u0_u0_ch_adr0_r_reg[12] ;
  assign \new_[1773]_  = ~\\u0_u0_ch_adr0_r_reg[14] ;
  assign \new_[1774]_  = ~\\u0_u0_ch_adr0_r_reg[15] ;
  assign \new_[1775]_  = ~\\u0_u0_ch_adr0_r_reg[16] ;
  assign \new_[1776]_  = ~\\u0_u0_ch_adr0_r_reg[18] ;
  assign \new_[1777]_  = ~\\u0_u0_ch_adr0_r_reg[19] ;
  assign \new_[1778]_  = ~\\u0_u0_ch_adr0_r_reg[20] ;
  assign \new_[1779]_  = ~\\u0_u0_ch_adr0_r_reg[22] ;
  assign \new_[1780]_  = ~\\u0_u0_ch_adr0_r_reg[23] ;
  assign \new_[1781]_  = ~\\u0_u0_ch_adr0_r_reg[24] ;
  assign \new_[1782]_  = ~\\u0_u0_ch_adr0_r_reg[26] ;
  assign \new_[1783]_  = ~\\u0_u0_ch_adr0_r_reg[27] ;
  assign \new_[1784]_  = ~\\u0_u0_ch_adr0_r_reg[28] ;
  assign \new_[1785]_  = ~\new_[1964]_  | (~\new_[1995]_  & ~\new_[3994]_ );
  assign \new_[1786]_  = ~\\u0_u0_ch_adr0_r_reg[21] ;
  assign \new_[1787]_  = ~\\u0_u0_ch_adr0_r_reg[29] ;
  assign \new_[1788]_  = ~\\u0_u0_ch_adr0_r_reg[25] ;
  assign \new_[1789]_  = ~\\u0_u0_ch_tot_sz_r_reg[9] ;
  assign \new_[1790]_  = \new_[3742]_  ? \new_[4307]_  : \new_[3973]_ ;
  assign \new_[1791]_  = \new_[3583]_  ? \new_[4307]_  : \new_[4069]_ ;
  assign n1656 = ~\new_[2067]_  | ~\new_[3018]_  | ~\new_[2066]_ ;
  assign \new_[1793]_  = ~\new_[2062]_  & (~\new_[4047]_  | ~\new_[2064]_ );
  assign \new_[1794]_  = ~\new_[2065]_  & (~\new_[3996]_  | ~\new_[2064]_ );
  assign \new_[1795]_  = ~\new_[2060]_  & (~\new_[4112]_  | ~\new_[2064]_ );
  assign \new_[1796]_  = ~\\u0_u0_ch_tot_sz_r_reg[5] ;
  assign \new_[1797]_  = ~\\u0_u0_ch_tot_sz_r_reg[10] ;
  assign \new_[1798]_  = ~\\u0_u0_ch_tot_sz_r_reg[11] ;
  assign \new_[1799]_  = ~\\u0_u0_ch_tot_sz_r_reg[2] ;
  assign \new_[1800]_  = ~\\u0_u0_ch_tot_sz_r_reg[3] ;
  assign \new_[1801]_  = ~\\u0_u0_ch_tot_sz_r_reg[4] ;
  assign \new_[1802]_  = ~\\u0_u0_ch_tot_sz_r_reg[6] ;
  assign \new_[1803]_  = ~\\u0_u0_ch_tot_sz_r_reg[7] ;
  assign \new_[1804]_  = ~\\u0_u0_ch_tot_sz_r_reg[8] ;
  assign n1661 = ~\new_[1984]_  | (~\new_[2883]_  & ~\new_[3882]_ );
  assign n1646 = ~\new_[1963]_ ;
  assign \new_[1807]_  = ~\new_[1970]_  | ~\new_[4011]_ ;
  assign \new_[1808]_  = ~\new_[1969]_  | (~\new_[2094]_  & ~\new_[1370]_ );
  assign n1781 = \new_[3931]_  ? \new_[4272]_  : \new_[2117]_ ;
  assign n1786 = \new_[3938]_  ? \new_[4272]_  : \new_[2118]_ ;
  assign n1791 = \new_[3923]_  ? \new_[4272]_  : \new_[2119]_ ;
  assign n1676 = \new_[3936]_  ? \new_[4272]_  : \new_[2120]_ ;
  assign n1796 = \new_[3946]_  ? \new_[4272]_  : \new_[2121]_ ;
  assign n1801 = \new_[3932]_  ? \new_[4272]_  : \new_[2122]_ ;
  assign n1806 = \new_[3884]_  ? \new_[4272]_  : \new_[2123]_ ;
  assign n1671 = \new_[3899]_  ? \new_[4272]_  : \new_[2124]_ ;
  assign n1811 = \new_[3906]_  ? \new_[4272]_  : \new_[2125]_ ;
  assign n1816 = \new_[3927]_  ? \new_[4272]_  : \new_[2126]_ ;
  assign n1821 = \new_[3952]_  ? \new_[4272]_  : \new_[2127]_ ;
  assign n1856 = \new_[3925]_  ? \new_[4272]_  : \new_[2128]_ ;
  assign n1826 = \new_[3896]_  ? \new_[4272]_  : \new_[2129]_ ;
  assign n1831 = \new_[3928]_  ? \new_[4272]_  : \new_[2130]_ ;
  assign n1836 = \new_[3912]_  ? \new_[4272]_  : \new_[2131]_ ;
  assign n1866 = \new_[3929]_  ? \new_[4272]_  : \new_[2132]_ ;
  assign n1841 = \new_[3915]_  ? \new_[4272]_  : \new_[2133]_ ;
  assign n1846 = \new_[3913]_  ? \new_[4272]_  : \new_[2134]_ ;
  assign n1851 = \new_[3910]_  ? \new_[4272]_  : \new_[2135]_ ;
  assign n1861 = \new_[3903]_  ? \new_[4272]_  : \new_[2136]_ ;
  assign n1706 = \new_[3931]_  ? \new_[2939]_  : \new_[2097]_ ;
  assign n1711 = \new_[3938]_  ? \new_[2939]_  : \new_[2098]_ ;
  assign n1716 = \new_[3923]_  ? \new_[2750]_  : \new_[2100]_ ;
  assign n1691 = \new_[3936]_  ? \new_[2939]_  : \new_[2101]_ ;
  assign n1721 = \new_[3946]_  ? \new_[2939]_  : \new_[2102]_ ;
  assign n1726 = \new_[3932]_  ? \new_[2939]_  : \new_[2103]_ ;
  assign n1731 = \new_[3884]_  ? \new_[2750]_  : \new_[2104]_ ;
  assign \new_[1836]_  = \new_[1373]_  ^ \new_[2138]_ ;
  assign n1696 = \new_[3899]_  ? \new_[2939]_  : \new_[2099]_ ;
  assign n1736 = \new_[3906]_  ? \new_[2750]_  : \new_[2105]_ ;
  assign n1741 = \new_[3927]_  ? \new_[2939]_  : \new_[2106]_ ;
  assign n1746 = \new_[3952]_  ? \new_[2939]_  : \new_[2107]_ ;
  assign n1686 = \new_[3925]_  ? \new_[2750]_  : \new_[2108]_ ;
  assign \new_[1842]_  = \new_[1371]_  ^ \new_[2137]_ ;
  assign n1751 = \new_[3896]_  ? \new_[2750]_  : \new_[2109]_ ;
  assign n1756 = \new_[3928]_  ? \new_[2750]_  : \new_[2110]_ ;
  assign n1761 = \new_[3912]_  ? \new_[2750]_  : \new_[2111]_ ;
  assign n1666 = \new_[3929]_  ? \new_[2750]_  : \new_[2112]_ ;
  assign n1766 = \new_[3915]_  ? \new_[2750]_  : \new_[2113]_ ;
  assign n1771 = \new_[3913]_  ? \new_[2750]_  : \new_[2114]_ ;
  assign n1776 = \new_[3910]_  ? \new_[2750]_  : \new_[2115]_ ;
  assign n1681 = \new_[3903]_  ? \new_[2750]_  : \new_[2116]_ ;
  assign \new_[1851]_  = ~\new_[4059]_  | ~\new_[2063]_ ;
  assign \new_[1852]_  = ~\new_[4104]_  | ~\new_[2064]_ ;
  assign \new_[1853]_  = ~\\u0_u0_ch_csr_r_reg[4] ;
  assign \new_[1854]_  = ~\new_[2931]_  & (~\new_[2167]_  | ~\new_[3472]_ );
  assign \new_[1855]_  = ~\new_[4307]_  | ~\new_[1339]_ ;
  assign \new_[1856]_  = ~\new_[4179]_  | ~\new_[2064]_ ;
  assign \new_[1857]_  = ~\new_[4148]_  | ~\new_[2064]_ ;
  assign \new_[1858]_  = ~\new_[4060]_  | ~\new_[2064]_ ;
  assign \new_[1859]_  = ~\new_[4037]_  | ~\new_[2064]_ ;
  assign \new_[1860]_  = ~\new_[4020]_  | ~\new_[2063]_ ;
  assign \new_[1861]_  = ~\new_[4162]_  | ~\new_[2063]_ ;
  assign \new_[1862]_  = ~\new_[4050]_  | ~\new_[2063]_ ;
  assign \new_[1863]_  = ~\new_[4001]_  | ~\new_[2063]_ ;
  assign \new_[1864]_  = ~\new_[4153]_  | ~\new_[2063]_ ;
  assign \new_[1865]_  = ~\new_[4087]_  | ~\new_[2064]_ ;
  assign \new_[1866]_  = ~\new_[4285]_  | ~\new_[2063]_ ;
  assign \new_[1867]_  = ~\new_[3967]_  | ~\new_[2064]_ ;
  assign \new_[1868]_  = ~\new_[4281]_  | ~\new_[2064]_ ;
  assign \new_[1869]_  = ~\new_[4088]_  | ~\new_[2063]_ ;
  assign \new_[1870]_  = ~\new_[4014]_  | ~\new_[2064]_ ;
  assign \new_[1871]_  = ~u0_u0_ch_err_reg;
  assign \new_[1872]_  = ~\new_[3998]_  | ~\new_[2064]_ ;
  assign \new_[1873]_  = ~\new_[4021]_  | ~\new_[2063]_ ;
  assign \new_[1874]_  = ~\new_[4012]_  | ~\new_[2064]_ ;
  assign \new_[1875]_  = ~\new_[2063]_  | ~\new_[4101]_ ;
  assign \new_[1876]_  = \\u0_u0_ch_csr_r_reg[1] ;
  assign \new_[1877]_  = \\u0_u0_ch_csr_r_reg[2] ;
  assign \new_[1878]_  = ~\\u0_u0_ch_csr_r_reg[3] ;
  assign \new_[1879]_  = ~\\u0_u0_ch_adr1_r_reg[0] ;
  assign \new_[1880]_  = ~\\u0_u0_ch_adr1_r_reg[1] ;
  assign \new_[1881]_  = ~\new_[4177]_  | ~\new_[2063]_ ;
  assign \new_[1882]_  = ~\\u0_u0_ch_adr1_r_reg[3] ;
  assign \new_[1883]_  = ~\\u0_u0_ch_adr1_r_reg[4] ;
  assign \new_[1884]_  = ~\\u0_u0_ch_adr1_r_reg[5] ;
  assign \new_[1885]_  = ~\\u0_u0_ch_adr1_r_reg[7] ;
  assign \new_[1886]_  = ~\\u0_u0_ch_adr1_r_reg[8] ;
  assign \new_[1887]_  = ~\\u0_u0_ch_adr1_r_reg[9] ;
  assign \new_[1888]_  = ~\\u0_u0_ch_adr0_r_reg[9] ;
  assign \new_[1889]_  = ~\\u0_u0_ch_adr0_r_reg[0] ;
  assign \new_[1890]_  = ~\\u0_u0_ch_adr0_r_reg[1] ;
  assign \new_[1891]_  = ~\\u0_u0_ch_adr0_r_reg[3] ;
  assign \new_[1892]_  = ~\\u0_u0_ch_adr0_r_reg[4] ;
  assign \new_[1893]_  = ~\\u0_u0_ch_adr0_r_reg[5] ;
  assign \new_[1894]_  = ~\\u0_u0_ch_adr0_r_reg[7] ;
  assign \new_[1895]_  = ~\\u0_u0_int_src_r_reg[0] ;
  assign \new_[1896]_  = ~\new_[4058]_  | ~\new_[2064]_ ;
  assign \new_[1897]_  = ~\new_[4176]_  | ~\new_[2064]_ ;
  assign \new_[1898]_  = ~\new_[4096]_  | ~\new_[2063]_ ;
  assign \new_[1899]_  = ~\new_[4075]_  | ~\new_[2063]_ ;
  assign \new_[1900]_  = ~\new_[4159]_  | ~\new_[2064]_ ;
  assign \new_[1901]_  = ~\new_[4005]_  | ~\new_[2064]_ ;
  assign \new_[1902]_  = ~\new_[4098]_  | ~\new_[2064]_ ;
  assign \new_[1903]_  = ~\new_[4164]_  | ~\new_[2064]_ ;
  assign \new_[1904]_  = ~\new_[4092]_  | ~\new_[2064]_ ;
  assign \new_[1905]_  = ~\new_[4120]_  | ~\new_[2064]_ ;
  assign \new_[1906]_  = ~\new_[4090]_  | ~\new_[2064]_ ;
  assign \new_[1907]_  = ~\new_[4119]_  | ~\new_[2063]_ ;
  assign \new_[1908]_  = ~\new_[3995]_  | ~\new_[2063]_ ;
  assign \new_[1909]_  = ~\new_[3988]_  | ~\new_[2064]_ ;
  assign \new_[1910]_  = ~\new_[3990]_  | ~\new_[2064]_ ;
  assign \new_[1911]_  = ~\new_[3978]_  | ~\new_[2063]_ ;
  assign \new_[1912]_  = ~\new_[4121]_  | ~\new_[2064]_ ;
  assign \wb0m_data_o[26]  = \wb1s_data_i[26]  ? \new_[3606]_  : \new_[2157]_ ;
  assign \wb0m_data_o[25]  = \wb1s_data_i[25]  ? \new_[3606]_  : \new_[2158]_ ;
  assign \new_[1915]_  = ~\new_[4045]_  | ~\new_[2064]_ ;
  assign \wb0m_data_o[24]  = \wb1s_data_i[24]  ? \new_[3606]_  : \new_[2159]_ ;
  assign \wb0m_data_o[23]  = \wb1s_data_i[23]  ? \new_[3606]_  : \new_[2160]_ ;
  assign \wb0m_data_o[22]  = \wb1s_data_i[22]  ? \new_[3592]_  : \new_[2172]_ ;
  assign \wb0m_data_o[21]  = \wb1s_data_i[21]  ? \new_[3607]_  : \new_[2173]_ ;
  assign \wb0m_data_o[20]  = \wb1s_data_i[20]  ? \new_[3607]_  : \new_[2174]_ ;
  assign \wb0m_data_o[19]  = \wb1s_data_i[19]  ? \new_[3606]_  : \new_[2175]_ ;
  assign \wb0m_data_o[18]  = \wb1s_data_i[18]  ? \new_[3592]_  : \new_[2176]_ ;
  assign \wb0m_data_o[17]  = \wb1s_data_i[17]  ? \new_[3592]_  : \new_[2177]_ ;
  assign \new_[1924]_  = ~\new_[4043]_  | ~\new_[2064]_ ;
  assign \wb0m_data_o[16]  = \wb1s_data_i[16]  ? \new_[3607]_  : \new_[2178]_ ;
  assign \wb0m_data_o[15]  = \wb1s_data_i[15]  ? \new_[3592]_  : \new_[2179]_ ;
  assign \wb0m_data_o[14]  = \wb1s_data_i[14]  ? \new_[3606]_  : \new_[2161]_ ;
  assign \wb0m_data_o[13]  = \wb1s_data_i[13]  ? \new_[3607]_  : \new_[2162]_ ;
  assign \wb0m_data_o[12]  = \wb1s_data_i[12]  ? \new_[3607]_  : \new_[2163]_ ;
  assign \wb0m_data_o[11]  = \wb1s_data_i[11]  ? \new_[3607]_  : \new_[2180]_ ;
  assign \new_[1931]_  = ~\new_[3984]_  | ~\new_[2064]_ ;
  assign \wb0m_data_o[8]  = \wb1s_data_i[8]  ? \new_[3592]_  : \new_[2181]_ ;
  assign \wb0m_data_o[7]  = \wb1s_data_i[7]  ? \new_[3606]_  : \new_[2182]_ ;
  assign \wb0m_data_o[6]  = \wb1s_data_i[6]  ? \new_[3606]_  : \new_[2183]_ ;
  assign \wb0m_data_o[5]  = \wb1s_data_i[5]  ? \new_[3592]_  : \new_[2184]_ ;
  assign \wb0m_data_o[4]  = \wb1s_data_i[4]  ? \new_[3607]_  : \new_[2185]_ ;
  assign \wb0m_data_o[3]  = \wb1s_data_i[3]  ? \new_[3606]_  : \new_[2164]_ ;
  assign \wb0m_data_o[2]  = \wb1s_data_i[2]  ? \new_[3607]_  : \new_[2165]_ ;
  assign \new_[1939]_  = ~\new_[4180]_  | ~\new_[2064]_ ;
  assign \wb0m_data_o[0]  = \wb1s_data_i[0]  ? \new_[3592]_  : \new_[2166]_ ;
  assign \new_[1941]_  = ~\new_[4100]_  | ~\new_[2064]_ ;
  assign \new_[1942]_  = ~\new_[4160]_  | ~\new_[2063]_ ;
  assign \new_[1943]_  = ~\new_[3975]_  | ~\new_[2064]_ ;
  assign \new_[1944]_  = ~\new_[4083]_  | ~\new_[2063]_ ;
  assign \new_[1945]_  = ~\new_[4165]_  | ~\new_[2063]_ ;
  assign \new_[1946]_  = ~\new_[4169]_  | ~\new_[2063]_ ;
  assign \new_[1947]_  = ~\new_[4052]_  | ~\new_[2064]_ ;
  assign \new_[1948]_  = ~\new_[4056]_  | ~\new_[2064]_ ;
  assign \new_[1949]_  = ~\new_[4064]_  | ~\new_[2064]_ ;
  assign \new_[1950]_  = ~\new_[4026]_  | ~\new_[2064]_ ;
  assign \new_[1951]_  = ~\new_[4138]_  | ~\new_[2063]_ ;
  assign \new_[1952]_  = ~\new_[4129]_  | ~\new_[2064]_ ;
  assign \new_[1953]_  = ~\new_[4063]_  | ~\new_[2064]_ ;
  assign \new_[1954]_  = ~\new_[4030]_  | ~\new_[2063]_ ;
  assign \new_[1955]_  = ~\new_[4142]_  | ~\new_[2064]_ ;
  assign \new_[1956]_  = ~\new_[4182]_  | ~\new_[2064]_ ;
  assign \new_[1957]_  = ~\new_[4145]_  | ~\new_[2063]_ ;
  assign \new_[1958]_  = ~\new_[4034]_  | ~\new_[2063]_ ;
  assign n1701 = \new_[3897]_  ? \new_[2883]_  : \new_[2073]_ ;
  assign \new_[1960]_  = ~\\u0_u0_ch_adr0_r_reg[6] ;
  assign \new_[1961]_  = ~n1651;
  assign \new_[1962]_  = ~\\u0_u0_ch_adr0_r_reg[2] ;
  assign \new_[1963]_  = ~\new_[2376]_  | ~\new_[2375]_  | ~\new_[2012]_  | ~\new_[2374]_ ;
  assign \new_[1964]_  = ~\new_[1995]_  | ~\new_[3994]_ ;
  assign \new_[1965]_  = ~\\u0_u0_ch_adr0_r_reg[8] ;
  assign \new_[1966]_  = ~\new_[2070]_  | (~\new_[2197]_  & ~\new_[1228]_ );
  assign \new_[1967]_  = ~\\u0_u0_ch_adr1_r_reg[6] ;
  assign \new_[1968]_  = ~\\u0_u0_ch_adr1_r_reg[2] ;
  assign \new_[1969]_  = ~\new_[2094]_  | ~\new_[1370]_ ;
  assign \new_[1970]_  = ~\new_[1373]_  | ~\new_[1370]_  | ~\new_[2137]_  | ~\new_[3851]_ ;
  assign \new_[1971]_  = \new_[1284]_  ^ \new_[2224]_ ;
  assign \new_[1972]_  = \new_[3959]_  ^ \new_[2225]_ ;
  assign \new_[1973]_  = \\u2_chunk_cnt_reg[8] ;
  assign \new_[1974]_  = \new_[2155]_  | \new_[3286]_ ;
  assign \new_[1975]_  = \new_[2139]_  | \new_[3100]_ ;
  assign \new_[1976]_  = \\u2_chunk_cnt_reg[7] ;
  assign \new_[1977]_  = \\u2_chunk_cnt_reg[6] ;
  assign \wb0m_data_o[30]  = \wb1s_data_i[30]  ? \new_[3607]_  : \new_[2238]_ ;
  assign \wb0m_data_o[29]  = \wb1s_data_i[29]  ? \new_[3607]_  : \new_[2239]_ ;
  assign \wb0m_data_o[28]  = \wb1s_data_i[28]  ? \new_[3606]_  : \new_[2240]_ ;
  assign \wb0m_data_o[27]  = \wb1s_data_i[27]  ? \new_[3607]_  : \new_[2241]_ ;
  assign \wb0m_data_o[9]  = \wb1s_data_i[9]  ? \new_[3607]_  : \new_[2226]_ ;
  assign \new_[1983]_  = ~\new_[2227]_  & (~\new_[2391]_  | ~\new_[3894]_ );
  assign \new_[1984]_  = ~\new_[2072]_  | ~\new_[2883]_ ;
  assign n1881 = ~\new_[2187]_  | (~\new_[2871]_  & ~\new_[2196]_ );
  assign n1886 = ~\new_[2188]_  | (~\new_[2872]_  & ~\new_[2196]_ );
  assign n1891 = ~\new_[2189]_  | (~\new_[2874]_  & ~\new_[2196]_ );
  assign n1896 = ~\new_[2190]_  | (~\new_[2823]_  & ~\new_[2196]_ );
  assign n1901 = ~\new_[2191]_  | (~\new_[2876]_  & ~\new_[2196]_ );
  assign n1876 = ~\new_[2192]_  | (~\new_[2828]_  & ~\new_[2196]_ );
  assign n1906 = ~\new_[2193]_  | (~\new_[2829]_  & ~\new_[2196]_ );
  assign n1911 = ~\new_[2194]_  | (~\new_[2830]_  & ~\new_[2196]_ );
  assign n1916 = ~\new_[2195]_  | (~\new_[2877]_  & ~\new_[2196]_ );
  assign n1871 = ~\new_[2071]_  | (~\new_[2869]_  & ~\new_[2196]_ );
  assign \new_[1995]_  = ~\new_[1284]_  | ~\new_[1228]_  | ~\new_[2225]_  | ~\new_[3803]_ ;
  assign n1931 = \new_[3897]_  ? \new_[2873]_  : \new_[2286]_ ;
  assign n1936 = \new_[3859]_  ? \new_[2873]_  : \new_[2287]_ ;
  assign n1941 = \new_[3845]_  ? \new_[2873]_  : \new_[2288]_ ;
  assign \new_[1999]_  = \\u1_ch_sel_r_reg[2] ;
  assign n1921 = \new_[3844]_  ? \new_[2873]_  : \new_[2289]_ ;
  assign n1946 = ~\new_[2203]_  | (~\new_[2947]_  & ~\new_[2406]_ );
  assign n2046 = ~\new_[2202]_  | (~\new_[2868]_  & ~\new_[2406]_ );
  assign n1951 = ~\new_[2205]_  | (~\new_[2864]_  & ~\new_[2406]_ );
  assign n1956 = ~\new_[2204]_  | (~\new_[2824]_  & ~\new_[2406]_ );
  assign n1961 = ~\new_[2206]_  | (~\new_[2825]_  & ~\new_[2406]_ );
  assign n1966 = ~\new_[2207]_  | (~\new_[2870]_  & ~\new_[2406]_ );
  assign n2041 = ~\new_[2208]_  | (~\new_[2879]_  & ~\new_[2406]_ );
  assign n1971 = ~\new_[2211]_  | (~\new_[2886]_  & ~\new_[2406]_ );
  assign n1976 = ~\new_[2210]_  | (~\new_[2881]_  & ~\new_[2406]_ );
  assign n1981 = ~\new_[2209]_  | (~\new_[2826]_  & ~\new_[2406]_ );
  assign n1986 = ~\new_[2212]_  | (~\new_[2946]_  & ~\new_[4270]_ );
  assign \new_[2012]_  = ~\new_[2201]_  & ~\new_[2200]_ ;
  assign n1991 = ~\new_[2214]_  | (~\new_[2880]_  & ~\new_[4270]_ );
  assign n1996 = ~\new_[2215]_  | (~\new_[2884]_  & ~\new_[4270]_ );
  assign n2031 = ~\new_[2216]_  | (~\new_[2888]_  & ~\new_[4270]_ );
  assign n2001 = ~\new_[2213]_  | (~\new_[2889]_  & ~\new_[4270]_ );
  assign n2006 = ~\new_[2217]_  | (~\new_[2890]_  & ~\new_[4270]_ );
  assign n2011 = ~\new_[2218]_  | (~\new_[2891]_  & ~\new_[4270]_ );
  assign n2026 = ~\new_[2219]_  | (~\new_[2892]_  & ~\new_[4270]_ );
  assign n2016 = ~\new_[2220]_  | (~\new_[2893]_  & ~\new_[4270]_ );
  assign n2036 = ~\new_[2221]_  | (~\new_[2896]_  & ~\new_[4270]_ );
  assign \new_[2022]_  = \new_[1372]_  ^ \new_[2330]_ ;
  assign \new_[2023]_  = ~\new_[4306]_ ;
  assign \new_[2024]_  = ~\new_[2569]_  & ~\new_[2222]_ ;
  assign \new_[2025]_  = \new_[1413]_  ^ \new_[2331]_ ;
  assign n1926 = ~\new_[2769]_  | ~\new_[2223]_ ;
  assign n2021 = ~\new_[2790]_  | ~\new_[2223]_ ;
  assign \new_[2028]_  = \\u1_ch_sel_r_reg[1] ;
  assign \new_[2029]_  = \\u1_ch_sel_r_reg[3] ;
  assign \new_[2030]_  = \\u1_ch_sel_r_reg[4] ;
  assign \new_[2031]_  = \\u2_chunk_cnt_reg[1] ;
  assign \new_[2032]_  = \\u2_chunk_cnt_reg[3] ;
  assign \new_[2033]_  = \\u2_chunk_cnt_reg[4] ;
  assign \new_[2034]_  = \\u2_chunk_cnt_reg[0] ;
  assign \new_[2035]_  = ~\new_[4306]_ ;
  assign \new_[2036]_  = ~\new_[4306]_ ;
  assign \new_[2037]_  = ~\new_[4306]_ ;
  assign \new_[2038]_  = ~\new_[4306]_ ;
  assign \wb0m_data_o[1]  = \wb1s_data_i[1]  ? \new_[3607]_  : \new_[2248]_ ;
  assign \wb1s_data_o[31]  = \wb0m_data_i[31]  ? \new_[3607]_  : \new_[2284]_ ;
  assign \wb1s_data_o[30]  = \wb0m_data_i[30]  ? \new_[3607]_  : \new_[2281]_ ;
  assign \wb1s_data_o[29]  = \wb0m_data_i[29]  ? \new_[3606]_  : \new_[2282]_ ;
  assign \wb1s_data_o[28]  = \wb0m_data_i[28]  ? \new_[3606]_  : \new_[2283]_ ;
  assign \wb1s_data_o[27]  = \wb0m_data_i[27]  ? \new_[3606]_  : \new_[2285]_ ;
  assign \wb1s_data_o[26]  = \wb0m_data_i[26]  ? \new_[3592]_  : \new_[2266]_ ;
  assign \wb1s_data_o[25]  = \wb0m_data_i[25]  ? \new_[3606]_  : \new_[2267]_ ;
  assign \wb1s_data_o[24]  = \wb0m_data_i[24]  ? \new_[3606]_  : \new_[2268]_ ;
  assign \wb1s_data_o[23]  = \wb0m_data_i[23]  ? \new_[3606]_  : \new_[2269]_ ;
  assign \wb1s_data_o[22]  = \wb0m_data_i[22]  ? \new_[3606]_  : \new_[2270]_ ;
  assign \wb1s_data_o[21]  = \wb0m_data_i[21]  ? \new_[3606]_  : \new_[2271]_ ;
  assign \wb1s_data_o[20]  = \wb0m_data_i[20]  ? \new_[3606]_  : \new_[2272]_ ;
  assign \wb1s_data_o[19]  = \wb0m_data_i[19]  ? \new_[3606]_  : \new_[2273]_ ;
  assign \wb1s_data_o[18]  = \wb0m_data_i[18]  ? \new_[3607]_  : \new_[2274]_ ;
  assign \wb1s_data_o[17]  = \wb0m_data_i[17]  ? \new_[3607]_  : \new_[2275]_ ;
  assign \wb1s_data_o[16]  = \wb0m_data_i[16]  ? \new_[3607]_  : \new_[2276]_ ;
  assign \wb1s_data_o[15]  = \wb0m_data_i[15]  ? \new_[3606]_  : \new_[2277]_ ;
  assign \wb1s_data_o[14]  = \wb0m_data_i[14]  ? \new_[3607]_  : \new_[2278]_ ;
  assign \wb1s_data_o[13]  = \wb0m_data_i[13]  ? \new_[3606]_  : \new_[2279]_ ;
  assign \wb1s_data_o[12]  = \wb0m_data_i[12]  ? \new_[3606]_  : \new_[2280]_ ;
  assign \new_[2060]_  = ~\new_[2247]_  & (~\new_[3734]_  | ~\new_[3194]_ );
  assign \new_[2061]_  = ~\new_[3131]_  & (~\new_[2249]_  | ~\new_[2428]_ );
  assign \new_[2062]_  = ~\new_[3657]_  & ~\new_[2247]_ ;
  assign \new_[2063]_  = ~\new_[4265]_ ;
  assign \new_[2064]_  = ~\new_[4267]_ ;
  assign \new_[2065]_  = ~\new_[2247]_  & (~\new_[3736]_  | ~\new_[3324]_ );
  assign \new_[2066]_  = ~\new_[3889]_  | ~\new_[3130]_  | ~\new_[2251]_ ;
  assign \new_[2067]_  = ~\new_[3224]_  | ~\new_[2428]_  | ~\new_[2250]_ ;
  assign \new_[2068]_  = \\u2_chunk_cnt_reg[5] ;
  assign \new_[2069]_  = \\u2_chunk_cnt_reg[2] ;
  assign \new_[2070]_  = ~\new_[2197]_  | ~\new_[1228]_ ;
  assign \new_[2071]_  = ~\new_[2788]_  & (~\new_[2789]_  | ~\new_[2355]_ );
  assign \new_[2072]_  = \new_[3066]_  ? \new_[2355]_  : \new_[4047]_ ;
  assign \new_[2073]_  = \new_[3067]_  ? \new_[2355]_  : \new_[4014]_ ;
  assign \new_[2074]_  = ~\new_[2266]_  | ~\new_[3659]_ ;
  assign \new_[2075]_  = ~\new_[2267]_  | ~\new_[3659]_ ;
  assign \new_[2076]_  = ~\new_[2268]_  | ~\new_[3659]_ ;
  assign \new_[2077]_  = ~\new_[2269]_  | ~\new_[3659]_ ;
  assign \new_[2078]_  = ~\new_[2270]_  | ~\new_[3659]_ ;
  assign \new_[2079]_  = ~\new_[2271]_  | ~\new_[3659]_ ;
  assign \new_[2080]_  = ~\new_[2272]_  | ~\new_[3659]_ ;
  assign \new_[2081]_  = ~\new_[2273]_  | ~\new_[3659]_ ;
  assign \new_[2082]_  = ~\new_[2274]_  | ~\new_[3659]_ ;
  assign \new_[2083]_  = ~\new_[2275]_  | ~\new_[3659]_ ;
  assign \new_[2084]_  = ~\new_[2276]_  | ~\new_[3659]_ ;
  assign \new_[2085]_  = ~\new_[2277]_  | ~\new_[3659]_ ;
  assign \new_[2086]_  = ~\new_[2278]_  | ~\new_[3659]_ ;
  assign \new_[2087]_  = ~\new_[2279]_  | ~\new_[3659]_ ;
  assign \new_[2088]_  = ~\new_[2280]_  | ~\new_[3659]_ ;
  assign \new_[2089]_  = ~\new_[2281]_  | ~\new_[3659]_ ;
  assign \new_[2090]_  = ~\new_[2282]_  | ~\new_[3659]_ ;
  assign \new_[2091]_  = ~\new_[2283]_  | ~\new_[3659]_ ;
  assign \new_[2092]_  = ~\new_[2284]_  | ~\new_[3659]_ ;
  assign \new_[2093]_  = ~\new_[2285]_  | ~\new_[3659]_ ;
  assign \new_[2094]_  = ~\new_[1382]_  | ~\new_[1373]_  | ~\new_[2330]_  | ~\new_[3836]_ ;
  assign \new_[2095]_  = \new_[1229]_  ^ \new_[2379]_ ;
  assign \new_[2096]_  = \new_[1285]_  ^ \new_[2377]_ ;
  assign \new_[2097]_  = ~\new_[2290]_  | (~\new_[3053]_  & ~\new_[2431]_ );
  assign \new_[2098]_  = ~\new_[2293]_  | (~\new_[2965]_  & ~\new_[2431]_ );
  assign \new_[2099]_  = ~\new_[2294]_  | (~\new_[2969]_  & ~\new_[2431]_ );
  assign \new_[2100]_  = ~\new_[2322]_  | (~\new_[2949]_  & ~\new_[2431]_ );
  assign \new_[2101]_  = ~\new_[2291]_  | (~\new_[2962]_  & ~\new_[2431]_ );
  assign \new_[2102]_  = ~\new_[2292]_  | (~\new_[2950]_  & ~\new_[2431]_ );
  assign \new_[2103]_  = ~\new_[2307]_  | (~\new_[3054]_  & ~\new_[2431]_ );
  assign \new_[2104]_  = ~\new_[2329]_  | (~\new_[3055]_  & ~\new_[2431]_ );
  assign \new_[2105]_  = ~\new_[2295]_  | (~\new_[2951]_  & ~\new_[2431]_ );
  assign \new_[2106]_  = ~\new_[2296]_  | (~\new_[2961]_  & ~\new_[2431]_ );
  assign \new_[2107]_  = ~\new_[2297]_  | (~\new_[2866]_  & ~\new_[2431]_ );
  assign \new_[2108]_  = ~\new_[2298]_  | (~\new_[2955]_  & ~\new_[2431]_ );
  assign \new_[2109]_  = ~\new_[2299]_  | (~\new_[2956]_  & ~\new_[2431]_ );
  assign \new_[2110]_  = ~\new_[2300]_  | (~\new_[2957]_  & ~\new_[2431]_ );
  assign \new_[2111]_  = ~\new_[2301]_  | (~\new_[2959]_  & ~\new_[2431]_ );
  assign \new_[2112]_  = ~\new_[2302]_  | (~\new_[2952]_  & ~\new_[2431]_ );
  assign \new_[2113]_  = ~\new_[2303]_  | (~\new_[2867]_  & ~\new_[2431]_ );
  assign \new_[2114]_  = ~\new_[2304]_  | (~\new_[2982]_  & ~\new_[2431]_ );
  assign \new_[2115]_  = ~\new_[2305]_  | (~\new_[2960]_  & ~\new_[2431]_ );
  assign \new_[2116]_  = ~\new_[2306]_  | (~\new_[2966]_  & ~\new_[2431]_ );
  assign \new_[2117]_  = ~\new_[2308]_  | (~\new_[2967]_  & ~\new_[2413]_ );
  assign \new_[2118]_  = ~\new_[2309]_  | (~\new_[2968]_  & ~\new_[2414]_ );
  assign \new_[2119]_  = ~\new_[2310]_  | (~\new_[2875]_  & ~\new_[2413]_ );
  assign \new_[2120]_  = ~\new_[2311]_  | (~\new_[2983]_  & ~\new_[2412]_ );
  assign \new_[2121]_  = ~\new_[2312]_  | (~\new_[2970]_  & ~\new_[2412]_ );
  assign \new_[2122]_  = ~\new_[2313]_  | (~\new_[2971]_  & ~\new_[2412]_ );
  assign \new_[2123]_  = ~\new_[2314]_  | (~\new_[2972]_  & ~\new_[2414]_ );
  assign \new_[2124]_  = ~\new_[2315]_  | (~\new_[2973]_  & ~\new_[2412]_ );
  assign \new_[2125]_  = ~\new_[2316]_  | (~\new_[2974]_  & ~\new_[2413]_ );
  assign \new_[2126]_  = ~\new_[2317]_  | (~\new_[2975]_  & ~\new_[2413]_ );
  assign \new_[2127]_  = ~\new_[2318]_  | (~\new_[2885]_  & ~\new_[2413]_ );
  assign \new_[2128]_  = ~\new_[2319]_  | (~\new_[2976]_  & ~\new_[2413]_ );
  assign \new_[2129]_  = ~\new_[2320]_  | (~\new_[2977]_  & ~\new_[2413]_ );
  assign \new_[2130]_  = ~\new_[2321]_  | (~\new_[2978]_  & ~\new_[2414]_ );
  assign \new_[2131]_  = ~\new_[2323]_  | (~\new_[2979]_  & ~\new_[2414]_ );
  assign \new_[2132]_  = ~\new_[2324]_  | (~\new_[2980]_  & ~\new_[2413]_ );
  assign \new_[2133]_  = ~\new_[2325]_  | (~\new_[2887]_  & ~\new_[2413]_ );
  assign \new_[2134]_  = ~\new_[2326]_  | (~\new_[2963]_  & ~\new_[2413]_ );
  assign \new_[2135]_  = ~\new_[2327]_  | (~\new_[2981]_  & ~\new_[2413]_ );
  assign \new_[2136]_  = ~\new_[2328]_  | (~\new_[2964]_  & ~\new_[2413]_ );
  assign \new_[2137]_  = ~\new_[2332]_  & ~\new_[3812]_ ;
  assign \new_[2138]_  = \new_[3791]_  & \new_[2331]_ ;
  assign \new_[2139]_  = ~\new_[2334]_  | ~\new_[2333]_ ;
  assign \new_[2140]_  = \new_[3935]_  ^ \new_[2348]_ ;
  assign \new_[2141]_  = \\u1_ch_sel_r_reg[0] ;
  assign \wb0m_data_o[31]  = \wb1s_data_i[31]  ? \new_[3592]_  : \new_[2347]_ ;
  assign \wb1s_data_o[11]  = \wb0m_data_i[11]  ? \new_[3592]_  : \new_[2362]_ ;
  assign \wb1s_data_o[10]  = \wb0m_data_i[10]  ? \new_[3606]_  : \new_[2363]_ ;
  assign \wb1s_data_o[9]  = \wb0m_data_i[9]  ? \new_[3607]_  : \new_[2364]_ ;
  assign \wb1s_data_o[8]  = \wb0m_data_i[8]  ? \new_[3592]_  : \new_[2365]_ ;
  assign \wb1s_data_o[7]  = \wb0m_data_i[7]  ? \new_[3592]_  : \new_[2366]_ ;
  assign \wb1s_data_o[6]  = \wb0m_data_i[6]  ? \new_[3607]_  : \new_[2367]_ ;
  assign \wb1s_data_o[5]  = \wb0m_data_i[5]  ? \new_[3592]_  : \new_[2369]_ ;
  assign \wb1s_data_o[4]  = \wb0m_data_i[4]  ? \new_[3592]_  : \new_[2370]_ ;
  assign \wb1s_data_o[3]  = \wb0m_data_i[3]  ? \new_[3607]_  : \new_[2358]_ ;
  assign \wb1s_data_o[2]  = \wb0m_data_i[2]  ? \new_[3606]_  : \new_[2359]_ ;
  assign \wb1s_data_o[1]  = \wb0m_data_i[1]  ? \new_[3606]_  : \new_[2360]_ ;
  assign \wb1s_data_o[0]  = \wb0m_data_i[0]  ? \new_[3607]_  : \new_[2361]_ ;
  assign \new_[2155]_  = ~\new_[2832]_  & (~\new_[2391]_  | ~\new_[3911]_ );
  assign n2051 = ~\new_[2380]_  | (~\new_[2394]_  & ~\new_[2375]_ );
  assign \new_[2157]_  = \\u0_wb_rf_dout_reg[26] ;
  assign \new_[2158]_  = \\u0_wb_rf_dout_reg[25] ;
  assign \new_[2159]_  = \\u0_wb_rf_dout_reg[24] ;
  assign \new_[2160]_  = \\u0_wb_rf_dout_reg[23] ;
  assign \new_[2161]_  = \\u0_wb_rf_dout_reg[14] ;
  assign \new_[2162]_  = \\u0_wb_rf_dout_reg[13] ;
  assign \new_[2163]_  = \\u0_wb_rf_dout_reg[12] ;
  assign \new_[2164]_  = \\u0_wb_rf_dout_reg[3] ;
  assign \new_[2165]_  = \\u0_wb_rf_dout_reg[2] ;
  assign \new_[2166]_  = \\u0_wb_rf_dout_reg[0] ;
  assign \new_[2167]_  = ~\new_[2417]_  & ~\new_[3286]_ ;
  assign \new_[2168]_  = ~\new_[3909]_  | ~\new_[3224]_  | ~\new_[2353]_ ;
  assign n2061 = ~\new_[2386]_  | (~\new_[2394]_  & ~\new_[2374]_ );
  assign n2056 = ~\new_[2387]_  | (~\new_[2394]_  & ~\new_[2376]_ );
  assign \new_[2171]_  = \new_[3992]_  ^ \new_[2354]_ ;
  assign \new_[2172]_  = \\u0_wb_rf_dout_reg[22] ;
  assign \new_[2173]_  = \\u0_wb_rf_dout_reg[21] ;
  assign \new_[2174]_  = \\u0_wb_rf_dout_reg[20] ;
  assign \new_[2175]_  = \\u0_wb_rf_dout_reg[19] ;
  assign \new_[2176]_  = \\u0_wb_rf_dout_reg[18] ;
  assign \new_[2177]_  = \\u0_wb_rf_dout_reg[17] ;
  assign \new_[2178]_  = \\u0_wb_rf_dout_reg[16] ;
  assign \new_[2179]_  = \\u0_wb_rf_dout_reg[15] ;
  assign \new_[2180]_  = \\u0_wb_rf_dout_reg[11] ;
  assign \new_[2181]_  = \\u0_wb_rf_dout_reg[8] ;
  assign \new_[2182]_  = \\u0_wb_rf_dout_reg[7] ;
  assign \new_[2183]_  = \\u0_wb_rf_dout_reg[6] ;
  assign \new_[2184]_  = \\u0_wb_rf_dout_reg[5] ;
  assign \new_[2185]_  = \\u0_wb_rf_dout_reg[4] ;
  assign \new_[2186]_  = ~\new_[2247]_ ;
  assign \new_[2187]_  = ~\new_[2770]_  & (~\new_[2771]_  | ~\new_[2355]_ );
  assign \new_[2188]_  = ~\new_[2772]_  & (~\new_[2773]_  | ~\new_[2355]_ );
  assign \new_[2189]_  = ~\new_[2774]_  & (~\new_[2775]_  | ~\new_[2355]_ );
  assign \new_[2190]_  = ~\new_[2776]_  & (~\new_[2777]_  | ~\new_[2355]_ );
  assign \new_[2191]_  = ~\new_[2778]_  & (~\new_[2779]_  | ~\new_[2355]_ );
  assign \new_[2192]_  = ~\new_[2780]_  & (~\new_[2781]_  | ~\new_[2355]_ );
  assign \new_[2193]_  = ~\new_[2782]_  & (~\new_[2783]_  | ~\new_[2355]_ );
  assign \new_[2194]_  = ~\new_[2784]_  & (~\new_[2785]_  | ~\new_[2355]_ );
  assign \new_[2195]_  = ~\new_[2786]_  & (~\new_[2787]_  | ~\new_[2355]_ );
  assign \new_[2196]_  = ~\new_[2356]_  | ~\new_[2883]_ ;
  assign \new_[2197]_  = ~\new_[1234]_  | ~\new_[1284]_  | ~\new_[2379]_  | ~\new_[3850]_ ;
  assign \new_[2198]_  = \new_[1231]_  ^ \new_[2392]_ ;
  assign \new_[2199]_  = \new_[1382]_  ^ \new_[2399]_ ;
  assign \new_[2200]_  = ~\new_[2393]_  | ~\new_[2409]_  | ~\new_[2408]_ ;
  assign \new_[2201]_  = ~\new_[2411]_  | ~\new_[2410]_  | ~\new_[2415]_ ;
  assign \new_[2202]_  = ~\new_[2704]_  & (~\new_[2708]_  | ~\new_[2431]_ );
  assign \new_[2203]_  = ~\new_[2702]_  & (~\new_[2703]_  | ~\new_[2431]_ );
  assign \new_[2204]_  = ~\new_[2727]_  & (~\new_[2709]_  | ~\new_[2431]_ );
  assign \new_[2205]_  = ~\new_[2705]_  & (~\new_[2706]_  | ~\new_[2431]_ );
  assign \new_[2206]_  = ~\new_[2714]_  & (~\new_[2710]_  | ~\new_[2431]_ );
  assign \new_[2207]_  = ~\new_[2711]_  & (~\new_[2707]_  | ~\new_[2431]_ );
  assign \new_[2208]_  = ~\new_[2712]_  & (~\new_[2713]_  | ~\new_[2431]_ );
  assign \new_[2209]_  = ~\new_[2715]_  & (~\new_[2716]_  | ~\new_[2431]_ );
  assign \new_[2210]_  = ~\new_[2725]_  & (~\new_[2724]_  | ~\new_[2431]_ );
  assign \new_[2211]_  = ~\new_[2728]_  & (~\new_[2726]_  | ~\new_[2431]_ );
  assign \new_[2212]_  = ~\new_[2763]_  & (~\new_[2764]_  | ~\new_[2412]_ );
  assign \new_[2213]_  = ~\new_[2765]_  & (~\new_[2802]_  | ~\new_[2412]_ );
  assign \new_[2214]_  = ~\new_[2795]_  & (~\new_[2796]_  | ~\new_[2412]_ );
  assign \new_[2215]_  = ~\new_[2798]_  & (~\new_[2799]_  | ~\new_[2412]_ );
  assign \new_[2216]_  = ~\new_[2800]_  & (~\new_[2801]_  | ~\new_[2412]_ );
  assign \new_[2217]_  = ~\new_[2803]_  & (~\new_[2804]_  | ~\new_[2412]_ );
  assign \new_[2218]_  = ~\new_[2805]_  & (~\new_[2806]_  | ~\new_[2414]_ );
  assign \new_[2219]_  = ~\new_[2807]_  & (~\new_[2808]_  | ~\new_[2414]_ );
  assign \new_[2220]_  = ~\new_[2809]_  & (~\new_[2810]_  | ~\new_[2412]_ );
  assign \new_[2221]_  = ~\new_[2811]_  & (~\new_[2812]_  | ~\new_[2412]_ );
  assign \new_[2222]_  = ~u0_u0_ch_busy_reg;
  assign \new_[2223]_  = ~\new_[2507]_  | ~\new_[2514]_ ;
  assign \new_[2224]_  = \new_[3730]_  & \new_[2377]_ ;
  assign \new_[2225]_  = ~\new_[2378]_  & ~\new_[3881]_ ;
  assign \new_[2226]_  = \\u0_wb_rf_dout_reg[9] ;
  assign \new_[2227]_  = ~\new_[2333]_ ;
  assign n2101 = ~\new_[2389]_  | (~\new_[2394]_  & ~\new_[2410]_ );
  assign n2086 = ~\new_[2382]_  | (~\new_[2394]_  & ~\new_[2415]_ );
  assign n2111 = ~\new_[2383]_  | (~\new_[2394]_  & ~\new_[2411]_ );
  assign n2091 = ~\new_[2384]_  | (~\new_[2394]_  & ~\new_[2409]_ );
  assign n2096 = ~\new_[2390]_  | (~\new_[2394]_  & ~\new_[2408]_ );
  assign n2106 = ~\new_[2385]_  | (~\new_[2394]_  & ~\new_[2393]_ );
  assign n2071 = \new_[2648]_  ? \new_[2394]_  : \new_[2028]_ ;
  assign n2066 = \new_[4053]_  ? \new_[2394]_  : \new_[1999]_ ;
  assign n2076 = \new_[2635]_  ? \new_[2394]_  : \new_[2029]_ ;
  assign n2081 = \new_[2641]_  ? \new_[2394]_  : \new_[2030]_ ;
  assign \new_[2238]_  = \\u0_wb_rf_dout_reg[30] ;
  assign \new_[2239]_  = \\u0_wb_rf_dout_reg[29] ;
  assign \new_[2240]_  = \\u0_wb_rf_dout_reg[28] ;
  assign \new_[2241]_  = \\u0_wb_rf_dout_reg[27] ;
  assign \new_[2242]_  = ~\new_[4290]_ ;
  assign \new_[2243]_  = ~\new_[4290]_ ;
  assign \new_[2244]_  = ~\new_[4290]_ ;
  assign \new_[2245]_  = ~\new_[4290]_ ;
  assign \new_[2246]_  = ~\new_[4290]_ ;
  assign \new_[2247]_  = ~\new_[4290]_ ;
  assign \new_[2248]_  = \\u0_wb_rf_dout_reg[1] ;
  assign \new_[2249]_  = \new_[2402]_  | \new_[4242]_ ;
  assign \new_[2250]_  = \new_[2402]_  | \new_[3889]_ ;
  assign \new_[2251]_  = ~\new_[2403]_  & ~\new_[2507]_ ;
  assign n2211 = ~\new_[2448]_  | ~\new_[4286]_  | ~\new_[2447]_  | ~\new_[2526]_ ;
  assign n2206 = ~\new_[2456]_  | ~\new_[4286]_  | ~\new_[2455]_  | ~\new_[2527]_ ;
  assign n2201 = ~\new_[2458]_  | ~\new_[4286]_  | ~\new_[2528]_  | ~\new_[2457]_ ;
  assign n2196 = ~\new_[4286]_  | ~\new_[2461]_  | ~\new_[2459]_  | ~\new_[2460]_ ;
  assign n2191 = ~\new_[4286]_  | ~\new_[2464]_  | ~\new_[2462]_  | ~\new_[2463]_ ;
  assign n2186 = ~\new_[4286]_  | ~\new_[2467]_  | ~\new_[2465]_  | ~\new_[2466]_ ;
  assign n2181 = ~\new_[4286]_  | ~\new_[2471]_  | ~\new_[2469]_  | ~\new_[2470]_ ;
  assign n2176 = ~\new_[4286]_  | ~\new_[2474]_  | ~\new_[2472]_  | ~\new_[2473]_ ;
  assign n2171 = ~\new_[4286]_  | ~\new_[2477]_  | ~\new_[2475]_  | ~\new_[2476]_ ;
  assign n2236 = ~\new_[2495]_  | ~\new_[4286]_  | ~\new_[2534]_  | ~\new_[2494]_ ;
  assign n2231 = ~\new_[2497]_  | ~\new_[4286]_  | ~\new_[2535]_  | ~\new_[2496]_ ;
  assign n2226 = ~\new_[2499]_  | ~\new_[4286]_  | ~\new_[2536]_  | ~\new_[2498]_ ;
  assign n2221 = ~\new_[2501]_  | ~\new_[4286]_  | ~\new_[2537]_  | ~\new_[2500]_ ;
  assign n2216 = ~\new_[2503]_  | ~\new_[4286]_  | ~\new_[2502]_  | ~\new_[2538]_ ;
  assign \new_[2266]_  = \new_[3555]_  ? \new_[2566]_  : \new_[3294]_ ;
  assign \new_[2267]_  = \new_[3557]_  ? \new_[2566]_  : \new_[3263]_ ;
  assign \new_[2268]_  = \new_[3560]_  ? \new_[2430]_  : \new_[3276]_ ;
  assign \new_[2269]_  = \new_[3518]_  ? \new_[2566]_  : \new_[3275]_ ;
  assign \new_[2270]_  = \new_[3522]_  ? \new_[2566]_  : \new_[3248]_ ;
  assign \new_[2271]_  = \new_[3558]_  ? \new_[2566]_  : \new_[3279]_ ;
  assign \new_[2272]_  = \new_[3519]_  ? \new_[2429]_  : \new_[3262]_ ;
  assign \new_[2273]_  = \new_[3572]_  ? \new_[2429]_  : \new_[3227]_ ;
  assign \new_[2274]_  = \new_[3568]_  ? \new_[2429]_  : \new_[3250]_ ;
  assign \new_[2275]_  = \new_[3562]_  ? \new_[2430]_  : \new_[3269]_ ;
  assign \new_[2276]_  = \new_[3521]_  ? \new_[2566]_  : \new_[3295]_ ;
  assign \new_[2277]_  = \new_[3575]_  ? \new_[2566]_  : \new_[3259]_ ;
  assign \new_[2278]_  = \new_[3564]_  ? \new_[2566]_  : \new_[3264]_ ;
  assign \new_[2279]_  = \new_[3547]_  ? \new_[2566]_  : \new_[3267]_ ;
  assign \new_[2280]_  = \new_[3525]_  ? \new_[2566]_  : \new_[3255]_ ;
  assign \new_[2281]_  = \new_[3576]_  ? \new_[2566]_  : \new_[3235]_ ;
  assign \new_[2282]_  = \new_[3569]_  ? \new_[2566]_  : \new_[3228]_ ;
  assign \new_[2283]_  = \new_[3566]_  ? \new_[2430]_  : \new_[3226]_ ;
  assign \new_[2284]_  = \new_[3563]_  ? \new_[2430]_  : \new_[3272]_ ;
  assign \new_[2285]_  = \new_[3553]_  ? \new_[2429]_  : \new_[3274]_ ;
  assign \new_[2286]_  = \new_[1876]_  ? \new_[2432]_  : \new_[3295]_ ;
  assign \new_[2287]_  = \new_[1877]_  ? \new_[2432]_  : \new_[3269]_ ;
  assign \new_[2288]_  = \new_[4130]_  ? \new_[2432]_  : \new_[3250]_ ;
  assign \new_[2289]_  = \new_[4175]_  ? \new_[2432]_  : \new_[3227]_ ;
  assign \new_[2290]_  = ~\new_[2431]_  | ~\new_[4165]_ ;
  assign \new_[2291]_  = ~\new_[2431]_  | ~\new_[4056]_ ;
  assign \new_[2292]_  = ~\new_[2431]_  | ~\new_[4064]_ ;
  assign \new_[2293]_  = ~\new_[2431]_  | ~\new_[4169]_ ;
  assign \new_[2294]_  = ~\new_[2431]_  | ~\new_[4129]_ ;
  assign \new_[2295]_  = ~\new_[2431]_  | ~\new_[4063]_ ;
  assign \new_[2296]_  = ~\new_[2431]_  | ~\new_[4030]_ ;
  assign \new_[2297]_  = ~\new_[2431]_  | ~\new_[4142]_ ;
  assign \new_[2298]_  = ~\new_[2431]_  | ~\new_[4160]_ ;
  assign \new_[2299]_  = ~\new_[2431]_  | ~\new_[4182]_ ;
  assign \new_[2300]_  = ~\new_[2431]_  | ~\new_[4145]_ ;
  assign \new_[2301]_  = ~\new_[2431]_  | ~\new_[4034]_ ;
  assign \new_[2302]_  = ~\new_[2431]_  | ~\new_[4061]_ ;
  assign \new_[2303]_  = ~\new_[2431]_  | ~\new_[4179]_ ;
  assign \new_[2304]_  = ~\new_[2431]_  | ~\new_[4148]_ ;
  assign \new_[2305]_  = ~\new_[2431]_  | ~\new_[4060]_ ;
  assign \new_[2306]_  = ~\new_[2431]_  | ~\new_[4037]_ ;
  assign \new_[2307]_  = ~\new_[2431]_  | ~\new_[4026]_ ;
  assign \new_[2308]_  = ~\new_[2414]_  | ~\new_[4059]_ ;
  assign \new_[2309]_  = ~\new_[2414]_  | ~\new_[4177]_ ;
  assign \new_[2310]_  = ~\new_[2414]_  | ~\new_[4058]_ ;
  assign \new_[2311]_  = ~\new_[2414]_  | ~\new_[4057]_ ;
  assign \new_[2312]_  = ~\new_[2414]_  | ~\new_[4176]_ ;
  assign \new_[2313]_  = ~\new_[2414]_  | ~\new_[4096]_ ;
  assign \new_[2314]_  = ~\new_[2414]_  | ~\new_[4075]_ ;
  assign \new_[2315]_  = ~\new_[2414]_  | ~\new_[4159]_ ;
  assign \new_[2316]_  = ~\new_[2414]_  | ~\new_[4005]_ ;
  assign \new_[2317]_  = ~\new_[2414]_  | ~\new_[4098]_ ;
  assign \new_[2318]_  = ~\new_[2414]_  | ~\new_[4164]_ ;
  assign \new_[2319]_  = ~\new_[2414]_  | ~\new_[4092]_ ;
  assign \new_[2320]_  = ~\new_[2414]_  | ~\new_[4120]_ ;
  assign \new_[2321]_  = ~\new_[2414]_  | ~\new_[4090]_ ;
  assign \new_[2322]_  = ~\new_[2431]_  | ~\new_[4052]_ ;
  assign \new_[2323]_  = ~\new_[2414]_  | ~\new_[4119]_ ;
  assign \new_[2324]_  = ~\new_[2414]_  | ~\new_[3995]_ ;
  assign \new_[2325]_  = ~\new_[2414]_  | ~\new_[3988]_ ;
  assign \new_[2326]_  = ~\new_[2414]_  | ~\new_[3990]_ ;
  assign \new_[2327]_  = ~\new_[2414]_  | ~\new_[3978]_ ;
  assign \new_[2328]_  = ~\new_[2414]_  | ~\new_[3981]_ ;
  assign \new_[2329]_  = ~\new_[2431]_  | ~\new_[4138]_ ;
  assign \new_[2330]_  = ~\new_[3784]_  & ~\new_[2404]_ ;
  assign \new_[2331]_  = ~\new_[3812]_  & ~\new_[2404]_ ;
  assign \new_[2332]_  = \new_[2404]_  | \new_[3942]_ ;
  assign \new_[2333]_  = ~\new_[2417]_  | ~\new_[2567]_ ;
  assign \new_[2334]_  = \new_[2417]_  | \new_[3909]_ ;
  assign n2116 = \new_[3887]_  ? \new_[2418]_  : \new_[2141]_ ;
  assign n2151 = ~\new_[2449]_  | ~\new_[4286]_  | ~\new_[2450]_  | ~\new_[2576]_ ;
  assign n2146 = ~\new_[2451]_  | ~\new_[4286]_  | ~\new_[2452]_  | ~\new_[2550]_ ;
  assign n2141 = ~\new_[2453]_  | ~\new_[4286]_  | ~\new_[2454]_  | ~\new_[2557]_ ;
  assign n2136 = ~\new_[2478]_  | ~\new_[4286]_  | ~\new_[2479]_  | ~\new_[2559]_ ;
  assign n2131 = ~\new_[2480]_  | ~\new_[4286]_  | ~\new_[2481]_  | ~\new_[2558]_ ;
  assign n2126 = ~\new_[2482]_  | ~\new_[4286]_  | ~\new_[2483]_  | ~\new_[2556]_ ;
  assign n2121 = ~\new_[2484]_  | ~\new_[4286]_  | ~\new_[2485]_  | ~\new_[2555]_ ;
  assign n2161 = ~\new_[2489]_  | ~\new_[2553]_  | ~\new_[2490]_  | ~\new_[2539]_ ;
  assign n2156 = ~\new_[2492]_  | ~\new_[2551]_  | ~\new_[2493]_  | ~\new_[2540]_ ;
  assign n2166 = ~\new_[2446]_  | ~\new_[2579]_  | ~\new_[2554]_  | ~\new_[2444]_ ;
  assign n2241 = \new_[3317]_  & \new_[2514]_ ;
  assign \new_[2347]_  = \\u0_wb_rf_dout_reg[31] ;
  assign \new_[2348]_  = ~\new_[2404]_ ;
  assign n2266 = ~\new_[4286]_  | ~\new_[2529]_  | ~\new_[2486]_ ;
  assign n2261 = ~\new_[4286]_  | ~\new_[2530]_  | ~\new_[2487]_ ;
  assign n2256 = ~\new_[4286]_  | ~\new_[2531]_  | ~\new_[2488]_ ;
  assign n2251 = ~\new_[4286]_  | ~\new_[2532]_  | ~\new_[2491]_ ;
  assign \new_[2353]_  = ~\new_[2507]_  & ~\new_[2424]_ ;
  assign \new_[2354]_  = ~\new_[2420]_  & ~\new_[3797]_ ;
  assign \new_[2355]_  = \new_[2397]_ ;
  assign \new_[2356]_  = ~\new_[2397]_ ;
  assign \new_[2357]_  = \new_[1414]_  ^ \new_[2435]_ ;
  assign \new_[2358]_  = \new_[3529]_  ? \new_[2566]_  : \new_[3245]_ ;
  assign \new_[2359]_  = \new_[3559]_  ? \new_[2509]_  : \new_[3270]_ ;
  assign \new_[2360]_  = \new_[3554]_  ? \new_[2509]_  : \new_[3230]_ ;
  assign \new_[2361]_  = \new_[3561]_  ? \new_[2566]_  : \new_[3256]_ ;
  assign \new_[2362]_  = \new_[3524]_  ? \new_[2566]_  : \new_[3268]_ ;
  assign \new_[2363]_  = \new_[3567]_  ? \new_[2510]_  : \new_[3253]_ ;
  assign \new_[2364]_  = \new_[3571]_  ? \new_[2510]_  : \new_[3266]_ ;
  assign \new_[2365]_  = \new_[3565]_  ? \new_[2509]_  : \new_[3233]_ ;
  assign \new_[2366]_  = \new_[3528]_  ? \new_[2566]_  : \new_[3282]_ ;
  assign \new_[2367]_  = \new_[3570]_  ? \new_[2510]_  : \new_[3273]_ ;
  assign \new_[2368]_  = ~\new_[2403]_ ;
  assign \new_[2369]_  = \new_[3523]_  ? \new_[2510]_  : \new_[3287]_ ;
  assign \new_[2370]_  = \new_[3552]_  ? \new_[2509]_  : \new_[3225]_ ;
  assign \new_[2371]_  = ~\new_[3130]_  | ~\new_[2428]_ ;
  assign \new_[2372]_  = \new_[3745]_  & \new_[2428]_ ;
  assign \new_[2373]_  = \new_[2428]_  & \new_[3744]_ ;
  assign \new_[2374]_  = ~\new_[4085]_  | ~\new_[2514]_ ;
  assign \new_[2375]_  = ~\new_[4081]_  | ~\new_[2514]_ ;
  assign \new_[2376]_  = ~\new_[4108]_  | ~\new_[2514]_ ;
  assign \new_[2377]_  = ~\new_[3881]_  & ~\new_[2426]_ ;
  assign \new_[2378]_  = \new_[2426]_  | \new_[3955]_ ;
  assign \new_[2379]_  = ~\new_[3776]_  & ~\new_[2426]_ ;
  assign \new_[2380]_  = ~\new_[2418]_  | ~\new_[2865]_ ;
  assign \new_[2381]_  = \new_[3987]_  ^ \new_[2438]_ ;
  assign \new_[2382]_  = ~\new_[3582]_  | ~\new_[2418]_ ;
  assign \new_[2383]_  = ~\new_[3288]_  | ~\new_[2418]_ ;
  assign \new_[2384]_  = ~\new_[3292]_  | ~\new_[2418]_ ;
  assign \new_[2385]_  = ~\new_[3102]_  | ~\new_[2418]_ ;
  assign \new_[2386]_  = ~\new_[2418]_  | ~\new_[3210]_ ;
  assign \new_[2387]_  = ~\new_[2418]_  | ~\new_[3198]_ ;
  assign n2246 = ~\new_[2524]_  | ~\new_[2599]_  | ~\new_[2505]_  | ~\new_[2504]_ ;
  assign \new_[2389]_  = ~\new_[2418]_  | ~\new_[3656]_ ;
  assign \new_[2390]_  = ~\new_[2418]_  | ~\new_[3197]_ ;
  assign \new_[2391]_  = ~\new_[2417]_ ;
  assign \new_[2392]_  = ~\new_[2426]_ ;
  assign \new_[2393]_  = ~\new_[4062]_  | ~\new_[2514]_ ;
  assign \new_[2394]_  = ~\new_[2517]_ ;
  assign \new_[2395]_  = \new_[1234]_  ^ \new_[2520]_ ;
  assign \new_[2396]_  = \new_[1381]_  ^ \new_[2522]_ ;
  assign \new_[2397]_  = \new_[2443]_  & \new_[2445]_ ;
  assign n2271 = ~\new_[2506]_  | ~\new_[2468]_ ;
  assign \new_[2399]_  = ~\new_[2441]_  & ~\new_[3671]_ ;
  assign \new_[2400]_  = \new_[1232]_  ^ \new_[2516]_ ;
  assign \new_[2401]_  = ~\new_[2548]_  | ~\new_[2572]_  | ~\new_[2615]_ ;
  assign \new_[2402]_  = \new_[2424]_ ;
  assign \new_[2403]_  = ~\new_[2425]_ ;
  assign \new_[2404]_  = ~\new_[2435]_  | ~\new_[1414]_ ;
  assign \new_[2405]_  = ~\new_[2596]_  | ~\new_[2512]_  | ~\new_[2595]_ ;
  assign \new_[2406]_  = ~\new_[2511]_  | ~\new_[2939]_ ;
  assign \new_[2407]_  = \new_[2514]_  & \new_[3907]_ ;
  assign \new_[2408]_  = ~\new_[2642]_  | ~\new_[2514]_ ;
  assign \new_[2409]_  = ~\new_[2637]_  | ~\new_[2514]_ ;
  assign \new_[2410]_  = ~\new_[4015]_  | ~\new_[2514]_ ;
  assign \new_[2411]_  = ~\new_[2640]_  | ~\new_[2514]_ ;
  assign \new_[2412]_  = \new_[2414]_ ;
  assign \new_[2413]_  = \new_[2414]_ ;
  assign \new_[2414]_  = ~\new_[4271]_ ;
  assign \new_[2415]_  = ~\new_[2639]_  | ~\new_[2514]_ ;
  assign \new_[2416]_  = ~u2_tsz_cnt_is_0_r_reg;
  assign \new_[2417]_  = ~\new_[2434]_ ;
  assign \new_[2418]_  = \new_[2436]_ ;
  assign n2276 = ~\new_[2533]_  | ~\new_[4286]_ ;
  assign \new_[2420]_  = ~\new_[1382]_  | ~\new_[2522]_  | ~\new_[3825]_ ;
  assign \new_[2421]_  = \new_[1380]_  ^ \new_[2630]_ ;
  assign \new_[2422]_  = ~\new_[2593]_  | (~\new_[2552]_  & ~\new_[4367]_ );
  assign \new_[2423]_  = ~\new_[2571]_  | (~\new_[2549]_  & ~\new_[4366]_ );
  assign \new_[2424]_  = ~\new_[2523]_  | ~\new_[2564]_ ;
  assign \new_[2425]_  = ~\new_[2442]_ ;
  assign \new_[2426]_  = ~\new_[2516]_  | ~\new_[1232]_ ;
  assign \new_[2427]_  = ~\new_[2588]_  | ~\new_[2547]_ ;
  assign \new_[2428]_  = ~\new_[2507]_ ;
  assign \new_[2429]_  = ~\new_[2541]_ ;
  assign \new_[2430]_  = ~\new_[2541]_ ;
  assign \new_[2431]_  = ~\new_[2511]_ ;
  assign \new_[2432]_  = ~\new_[2654]_  & (~\new_[3320]_  | ~\new_[3087]_ );
  assign \new_[2433]_  = \new_[1375]_  ^ \new_[2562]_ ;
  assign \new_[2434]_  = ~\new_[2542]_  | ~\new_[2517]_ ;
  assign \new_[2435]_  = \new_[2562]_  & \new_[1375]_ ;
  assign \new_[2436]_  = ~\new_[2517]_ ;
  assign n2281 = ~\new_[2518]_ ;
  assign \new_[2438]_  = ~\new_[2560]_  & ~\new_[3827]_ ;
  assign \new_[2439]_  = ~\new_[2521]_ ;
  assign \new_[2440]_  = ~\new_[2563]_  & (~\new_[2683]_  | ~\new_[4322]_ );
  assign \new_[2441]_  = ~\new_[2630]_  | ~\new_[3825]_ ;
  assign \new_[2442]_  = ~\new_[2565]_  | ~\new_[2583]_ ;
  assign \new_[2443]_  = ~\new_[4209]_  | ~\new_[3471]_  | ~\new_[2514]_ ;
  assign \new_[2444]_  = (~\new_[2619]_  | ~\new_[2745]_ ) & (~\new_[4280]_  | ~\new_[4047]_ );
  assign \new_[2445]_  = ~\new_[3359]_  | ~\new_[2514]_  | ~\new_[3781]_  | ~\new_[4229]_ ;
  assign \new_[2446]_  = (~\new_[2591]_  | ~\new_[3966]_ ) & (~\new_[2928]_  | ~\new_[2592]_ );
  assign \new_[2447]_  = (~\new_[2591]_  | ~\new_[1417]_ ) & (~\new_[4167]_  | ~\new_[2592]_ );
  assign \new_[2448]_  = (~\new_[4280]_  | ~\new_[4088]_ ) & (~\new_[4374]_  | ~\new_[3967]_ );
  assign \new_[2449]_  = (~\new_[2591]_  | ~\new_[4073]_ ) & (~\new_[4284]_  | ~\new_[4165]_ );
  assign \new_[2450]_  = (~\new_[4019]_  | ~\new_[2592]_ ) & (~\new_[4031]_  | ~\new_[2653]_ );
  assign \new_[2451]_  = (~\new_[2591]_  | ~\new_[2609]_ ) & (~\new_[4284]_  | ~\new_[4169]_ );
  assign \new_[2452]_  = (~\new_[4172]_  | ~\new_[2592]_ ) & (~\new_[3968]_  | ~\new_[2653]_ );
  assign \new_[2453]_  = (~\new_[2591]_  | ~\new_[4127]_ ) & (~\new_[4284]_  | ~\new_[4052]_ );
  assign \new_[2454]_  = (~\new_[4107]_  | ~\new_[2592]_ ) & (~\new_[4181]_  | ~\new_[2653]_ );
  assign \new_[2455]_  = (~\new_[2591]_  | ~\new_[4076]_ ) & (~\new_[3972]_  | ~\new_[2592]_ );
  assign \new_[2456]_  = (~\new_[4280]_  | ~\new_[2633]_ ) & (~\new_[4284]_  | ~\new_[4056]_ );
  assign \new_[2457]_  = (~\new_[2591]_  | ~\new_[4016]_ ) & (~\new_[4113]_  | ~\new_[2592]_ );
  assign \new_[2458]_  = (~\new_[4280]_  | ~\new_[4015]_ ) & (~\new_[4284]_  | ~\new_[4064]_ );
  assign \new_[2459]_  = (~\new_[4132]_  | ~\new_[2592]_ ) & (~\new_[3964]_  | ~\new_[2653]_ );
  assign \new_[2460]_  = (~\new_[4280]_  | ~\new_[2639]_ ) & (~\new_[4284]_  | ~\new_[4026]_ );
  assign \new_[2461]_  = (~\new_[2591]_  | ~\new_[2601]_ ) & (~\new_[2620]_  | ~\new_[4096]_ );
  assign \new_[2462]_  = (~\new_[4168]_  | ~\new_[2592]_ ) & (~\new_[4033]_  | ~\new_[2653]_ );
  assign \new_[2463]_  = (~\new_[4280]_  | ~\new_[2640]_ ) & (~\new_[4284]_  | ~\new_[4138]_ );
  assign \new_[2464]_  = (~\new_[2591]_  | ~\new_[2610]_ ) & (~\new_[2620]_  | ~\new_[4075]_ );
  assign \new_[2465]_  = (~\new_[4174]_  | ~\new_[2592]_ ) & (~\new_[4183]_  | ~\new_[2653]_ );
  assign \new_[2466]_  = (~\new_[4280]_  | ~\new_[2637]_ ) & (~\new_[4284]_  | ~\new_[4129]_ );
  assign \new_[2467]_  = (~\new_[2591]_  | ~\new_[2600]_ ) & (~\new_[2620]_  | ~\new_[4159]_ );
  assign \new_[2468]_  = (~\new_[4084]_  | ~\new_[2592]_ ) & (~\new_[4146]_  | ~\new_[2653]_ );
  assign \new_[2469]_  = (~\new_[4141]_  | ~\new_[2592]_ ) & (~\new_[4126]_  | ~\new_[2653]_ );
  assign \new_[2470]_  = (~\new_[4280]_  | ~\new_[2642]_ ) & (~\new_[4284]_  | ~\new_[4063]_ );
  assign \new_[2471]_  = (~\new_[2591]_  | ~\new_[4055]_ ) & (~\new_[2620]_  | ~\new_[4005]_ );
  assign \new_[2472]_  = (~\new_[3974]_  | ~\new_[2592]_ ) & (~\new_[4178]_  | ~\new_[2653]_ );
  assign \new_[2473]_  = (~\new_[4280]_  | ~\new_[4062]_ ) & (~\new_[4284]_  | ~\new_[4030]_ );
  assign \new_[2474]_  = (~\new_[2591]_  | ~\new_[4072]_ ) & (~\new_[2620]_  | ~\new_[4098]_ );
  assign \new_[2475]_  = (~\new_[4002]_  | ~\new_[2592]_ ) & (~\new_[4051]_  | ~\new_[2653]_ );
  assign \new_[2476]_  = (~\new_[4280]_  | ~\new_[4085]_ ) & (~\new_[4284]_  | ~\new_[4142]_ );
  assign \new_[2477]_  = (~\new_[2591]_  | ~\new_[4184]_ ) & (~\new_[2620]_  | ~\new_[4164]_ );
  assign \new_[2478]_  = (~\new_[4280]_  | ~\new_[4108]_ ) & (~\new_[4284]_  | ~\new_[4160]_ );
  assign \new_[2479]_  = (~\new_[4097]_  | ~\new_[2592]_ ) & (~\new_[4035]_  | ~\new_[2653]_ );
  assign \new_[2480]_  = (~\new_[4280]_  | ~\new_[4081]_ ) & (~\new_[4284]_  | ~\new_[4182]_ );
  assign \new_[2481]_  = (~\new_[3985]_  | ~\new_[2592]_ ) & (~\new_[4155]_  | ~\new_[2653]_ );
  assign \new_[2482]_  = (~\new_[4280]_  | ~\new_[4000]_ ) & (~\new_[4284]_  | ~\new_[4145]_ );
  assign \new_[2483]_  = (~\new_[4102]_  | ~\new_[2592]_ ) & (~\new_[4036]_  | ~\new_[2653]_ );
  assign \new_[2484]_  = (~\new_[4280]_  | ~\new_[4017]_ ) & (~\new_[4284]_  | ~\new_[4034]_ );
  assign \new_[2485]_  = (~\new_[4109]_  | ~\new_[2592]_ ) & (~\new_[4150]_  | ~\new_[2653]_ );
  assign \new_[2486]_  = (~\new_[4106]_  | ~\new_[2592]_ ) & (~\new_[4149]_  | ~\new_[2653]_ );
  assign \new_[2487]_  = (~\new_[4118]_  | ~\new_[2592]_ ) & (~\new_[4008]_  | ~\new_[2653]_ );
  assign \new_[2488]_  = (~\new_[4123]_  | ~\new_[2592]_ ) & (~\new_[4038]_  | ~\new_[2653]_ );
  assign \new_[2489]_  = (~\new_[4115]_  | ~\new_[2592]_ ) & (~\new_[4040]_  | ~\new_[2653]_ );
  assign \new_[2490]_  = (~\new_[4280]_  | ~\new_[4266]_ ) & (~\new_[4284]_  | ~\new_[4093]_ );
  assign \new_[2491]_  = (~\new_[4116]_  | ~\new_[2592]_ ) & (~\new_[4039]_  | ~\new_[2653]_ );
  assign \new_[2492]_  = (~\new_[3993]_  | ~\new_[2592]_ ) & (~\new_[3957]_  | ~\new_[2653]_ );
  assign \new_[2493]_  = (~\new_[4280]_  | ~\new_[3998]_ ) & (~\new_[4284]_  | ~\new_[3976]_ );
  assign \new_[2494]_  = (~\new_[2591]_  | ~\new_[4175]_ ) & (~\new_[4006]_  | ~\new_[2592]_ );
  assign \new_[2495]_  = (~\new_[4280]_  | ~\new_[3996]_ ) & (~\new_[4284]_  | ~\new_[4020]_ );
  assign \new_[2496]_  = (~\new_[2591]_  | ~\new_[2604]_ ) & (~\new_[4105]_  | ~\new_[2592]_ );
  assign \new_[2497]_  = (~\new_[4280]_  | ~\new_[4021]_ ) & (~\new_[4374]_  | ~\new_[4162]_ );
  assign \new_[2498]_  = (~\new_[2591]_  | ~\new_[2611]_ ) & (~\new_[4049]_  | ~\new_[2592]_ );
  assign \new_[2499]_  = (~\new_[4280]_  | ~\new_[4104]_ ) & (~\new_[4284]_  | ~\new_[4050]_ );
  assign \new_[2500]_  = (~\new_[2591]_  | ~\new_[2603]_ ) & (~\new_[4140]_  | ~\new_[2592]_ );
  assign \new_[2501]_  = (~\new_[4280]_  | ~\new_[4012]_ ) & (~\new_[4284]_  | ~\new_[4001]_ );
  assign \new_[2502]_  = (~\new_[2591]_  | ~\new_[2612]_ ) & (~\new_[4099]_  | ~\new_[2592]_ );
  assign \new_[2503]_  = (~\new_[4280]_  | ~\new_[4112]_ ) & (~\new_[4284]_  | ~\new_[4153]_ );
  assign \new_[2504]_  = (~\new_[2592]_  | ~\new_[3980]_ ) & (~\new_[2653]_  | ~\new_[4095]_ );
  assign \new_[2505]_  = (~\new_[4280]_  | ~\new_[4101]_ ) & (~\new_[4284]_  | ~\new_[4087]_ );
  assign \new_[2506]_  = (~\new_[4280]_  | ~\new_[4014]_ ) & (~\new_[2591]_  | ~\new_[1876]_ );
  assign \new_[2507]_  = u2_dma_abort_r_reg;
  assign \new_[2508]_  = ~\new_[2541]_ ;
  assign \new_[2509]_  = ~\new_[2541]_ ;
  assign \new_[2510]_  = ~\new_[2541]_ ;
  assign \new_[2511]_  = ~\new_[2543]_ ;
  assign \new_[2512]_  = ~\new_[2574]_  | ~\new_[4367]_ ;
  assign \new_[2513]_  = ~\new_[2623]_  | ~\new_[4363]_ ;
  assign \new_[2514]_  = ~\new_[2654]_ ;
  assign \new_[2515]_  = \new_[1233]_  ^ \new_[2580]_ ;
  assign \new_[2516]_  = \new_[2580]_  & \new_[1233]_ ;
  assign \new_[2517]_  = ~\new_[4158]_  | (~\new_[2629]_  & ~\new_[2546]_ );
  assign \new_[2518]_  = \new_[2632]_  | \new_[3774]_  | \new_[3786]_  | \new_[3653]_ ;
  assign \new_[2519]_  = \new_[1237]_  ^ \new_[2605]_ ;
  assign \new_[2520]_  = ~\new_[2581]_  & ~\new_[3799]_ ;
  assign \new_[2521]_  = ~\new_[2618]_  | ~\new_[2616]_  | ~\new_[2614]_ ;
  assign \new_[2522]_  = ~\new_[3671]_  & ~\new_[2584]_ ;
  assign \new_[2523]_  = ~wb1_ack_i | ~\new_[2585]_ ;
  assign \new_[2524]_  = ~\new_[2589]_  & (~\new_[2620]_  | ~\new_[4100]_ );
  assign \new_[2525]_  = ~\new_[2587]_  & (~\new_[2692]_  | ~\new_[2665]_ );
  assign \new_[2526]_  = (~\new_[3963]_  | ~\new_[2653]_ ) & (~\new_[2620]_  | ~\new_[4083]_ );
  assign \new_[2527]_  = (~\new_[4166]_  | ~\new_[2653]_ ) & (~\new_[2620]_  | ~\new_[4057]_ );
  assign \new_[2528]_  = (~\new_[4144]_  | ~\new_[2653]_ ) & (~\new_[2620]_  | ~\new_[4176]_ );
  assign \new_[2529]_  = (~\new_[4284]_  | ~\new_[4061]_ ) & (~\new_[2620]_  | ~\new_[3995]_ );
  assign \new_[2530]_  = (~\new_[4284]_  | ~\new_[4179]_ ) & (~\new_[2620]_  | ~\new_[3988]_ );
  assign \new_[2531]_  = (~\new_[4284]_  | ~\new_[4148]_ ) & (~\new_[2620]_  | ~\new_[3990]_ );
  assign \new_[2532]_  = (~\new_[4284]_  | ~\new_[4060]_ ) & (~\new_[2620]_  | ~\new_[3978]_ );
  assign \new_[2533]_  = (~\new_[4284]_  | ~\new_[4037]_ ) & (~\new_[2620]_  | ~\new_[3981]_ );
  assign \new_[2534]_  = (~\new_[4151]_  | ~\new_[2653]_ ) & (~\new_[2620]_  | ~\new_[4121]_ );
  assign \new_[2535]_  = (~\new_[4042]_  | ~\new_[2653]_ ) & (~\new_[2620]_  | ~\new_[4045]_ );
  assign \new_[2536]_  = (~\new_[4041]_  | ~\new_[2653]_ ) & (~\new_[2620]_  | ~\new_[4043]_ );
  assign \new_[2537]_  = (~\new_[4094]_  | ~\new_[2653]_ ) & (~\new_[2620]_  | ~\new_[3984]_ );
  assign \new_[2538]_  = (~\new_[4152]_  | ~\new_[2653]_ ) & (~\new_[2620]_  | ~\new_[4180]_ );
  assign \new_[2539]_  = ~\new_[2591]_  | ~\new_[1877]_ ;
  assign \new_[2540]_  = ~\new_[2591]_  | ~\new_[4130]_ ;
  assign \new_[2541]_  = ~\new_[2566]_ ;
  assign \new_[2542]_  = ~\new_[4073]_  | ~\new_[2514]_ ;
  assign \new_[2543]_  = ~\new_[3128]_  | ~\new_[2514]_ ;
  assign \new_[2544]_  = ~\new_[4364]_  | ~\new_[2697]_  | ~\new_[3636]_ ;
  assign \new_[2545]_  = ~\new_[2655]_  | ~\new_[2594]_ ;
  assign \new_[2546]_  = u1_de_start_r_reg;
  assign \new_[2547]_  = ~\new_[3633]_  | ~\new_[2751]_  | ~\new_[4364]_ ;
  assign \new_[2548]_  = ~\new_[2855]_  | ~\new_[3635]_  | ~\new_[2626]_ ;
  assign \new_[2549]_  = ~\new_[2621]_  & (~\new_[3718]_  | ~\new_[2667]_ );
  assign \new_[2550]_  = ~\new_[2620]_  | ~\new_[4177]_ ;
  assign \new_[2551]_  = ~\new_[2620]_  | ~\new_[4032]_ ;
  assign \new_[2552]_  = ~\new_[2622]_  & (~\new_[2667]_  | ~\new_[3629]_ );
  assign \new_[2553]_  = ~\new_[2620]_  | ~\new_[3961]_ ;
  assign \new_[2554]_  = ~\new_[2746]_  | ~\new_[2624]_  | ~\new_[2859]_ ;
  assign \new_[2555]_  = ~\new_[2620]_  | ~\new_[4119]_ ;
  assign \new_[2556]_  = ~\new_[2620]_  | ~\new_[4090]_ ;
  assign \new_[2557]_  = ~\new_[2620]_  | ~\new_[4058]_ ;
  assign \new_[2558]_  = ~\new_[2620]_  | ~\new_[4120]_ ;
  assign \new_[2559]_  = ~\new_[2620]_  | ~\new_[4092]_ ;
  assign \new_[2560]_  = ~\new_[1234]_  | ~\new_[2605]_  | ~\new_[3750]_ ;
  assign \new_[2561]_  = \new_[1236]_  ^ \new_[2646]_ ;
  assign \new_[2562]_  = \new_[2630]_  & \new_[1380]_ ;
  assign \new_[2563]_  = ~\new_[2834]_  & (~\new_[2659]_  | ~\new_[2656]_ );
  assign \new_[2564]_  = ~wb0_ack_i | ~\new_[2607]_ ;
  assign \new_[2565]_  = ~\new_[2613]_  | ~wb0_ack_i;
  assign \new_[2566]_  = ~\new_[2585]_ ;
  assign \new_[2567]_  = ~\new_[4013]_  & ~\new_[2654]_ ;
  assign \new_[2568]_  = ~\new_[2586]_ ;
  assign \new_[2569]_  = ~\new_[2591]_ ;
  assign n2286 = ~\new_[3872]_  | ~\new_[2625]_ ;
  assign \new_[2571]_  = ~\new_[2742]_  | ~\new_[4327]_ ;
  assign \new_[2572]_  = ~\new_[2694]_  | ~\new_[2628]_ ;
  assign \new_[2573]_  = ~\new_[2680]_  | ~\new_[2678]_ ;
  assign \new_[2574]_  = ~\new_[2680]_  | ~\new_[2679]_ ;
  assign \new_[2575]_  = \new_[2612]_  & \new_[2514]_ ;
  assign \new_[2576]_  = ~\new_[2620]_  | ~\new_[4059]_ ;
  assign \new_[2577]_  = \new_[1252]_  & \new_[2514]_ ;
  assign \new_[2578]_  = \\u2_state_reg[5] ;
  assign \new_[2579]_  = ~\new_[2833]_  | ~\new_[2653]_ ;
  assign \new_[2580]_  = \new_[2646]_  & \new_[1236]_ ;
  assign \new_[2581]_  = ~\new_[2646]_  | ~\new_[3750]_ ;
  assign \new_[2582]_  = ~\new_[2657]_  | ~\new_[2658]_ ;
  assign \new_[2583]_  = ~\new_[4311]_  | ~wb1_ack_i;
  assign \new_[2584]_  = ~\new_[2630]_ ;
  assign \new_[2585]_  = ~\new_[2607]_ ;
  assign \new_[2586]_  = ~\new_[2613]_ ;
  assign \new_[2587]_  = ~\new_[4386]_  & ~\new_[2835]_  & ~\new_[3719]_ ;
  assign \new_[2588]_  = ~\new_[3717]_  | ~\new_[2697]_  | ~\new_[4349]_ ;
  assign \new_[2589]_  = ~\new_[2617]_ ;
  assign \new_[2590]_  = ~\new_[2741]_  | ~\new_[2668]_ ;
  assign \new_[2591]_  = \new_[2661]_  & \new_[2859]_ ;
  assign \new_[2592]_  = ~\new_[2859]_  & ~\new_[2746]_  & ~\new_[3199]_  & ~\new_[2916]_ ;
  assign \new_[2593]_  = ~\new_[2669]_  | ~\new_[2663]_ ;
  assign \new_[2594]_  = ~\new_[2729]_  | ~\new_[4366]_ ;
  assign \new_[2595]_  = ~\new_[2664]_  | ~\new_[4367]_ ;
  assign \new_[2596]_  = ~\new_[2751]_  | ~\new_[2666]_ ;
  assign \new_[2597]_  = ~\new_[4349]_  | ~\new_[2751]_  | ~\new_[3626]_ ;
  assign \new_[2598]_  = ~\new_[2628]_ ;
  assign \new_[2599]_  = ~\new_[2916]_  | ~\new_[3056]_  | ~\new_[2677]_ ;
  assign \new_[2600]_  = \\u0_u0_ch_csr_r3_reg[2] ;
  assign \new_[2601]_  = \\u0_u0_ch_csr_r3_reg[0] ;
  assign \new_[2602]_  = ~u0_u0_rest_en_reg;
  assign \new_[2603]_  = \\u0_u0_ch_csr_r_reg[7] ;
  assign \new_[2604]_  = \\u0_u0_ch_csr_r_reg[5] ;
  assign \new_[2605]_  = ~\new_[3799]_  & ~\new_[2673]_ ;
  assign \new_[2606]_  = ~\\u0_u0_ch_csr_r2_reg[2] ;
  assign \new_[2607]_  = ~\new_[1877]_  | ~\new_[4211]_  | ~\new_[2834]_ ;
  assign \new_[2608]_  = ~\\u0_u0_ch_csr_r2_reg[1] ;
  assign \new_[2609]_  = \\u0_u0_ch_csr_r2_reg[0] ;
  assign \new_[2610]_  = \\u0_u0_ch_csr_r3_reg[1] ;
  assign \new_[2611]_  = \\u0_u0_ch_csr_r_reg[6] ;
  assign \new_[2612]_  = \\u0_u0_ch_csr_r_reg[8] ;
  assign \new_[2613]_  = ~\new_[4311]_ ;
  assign \new_[2614]_  = ~\new_[4211]_  | ~\new_[4368]_  | ~\new_[3625]_ ;
  assign \new_[2615]_  = ~\new_[3727]_  | ~\new_[2674]_ ;
  assign \new_[2616]_  = ~\new_[3624]_  | ~\new_[2835]_  | ~\new_[2729]_ ;
  assign \new_[2617]_  = ~\new_[2916]_  | ~\new_[3056]_  | ~\new_[2701]_ ;
  assign \new_[2618]_  = ~\new_[2815]_  | ~\new_[2681]_  | ~\new_[2819]_ ;
  assign \new_[2619]_  = \new_[2677]_  & \new_[3911]_ ;
  assign \new_[2620]_  = \new_[2677]_  & \new_[2936]_ ;
  assign \new_[2621]_  = ~\new_[3632]_  & ~\new_[2678]_ ;
  assign \new_[2622]_  = ~\new_[2678]_  & ~\new_[3672]_ ;
  assign \new_[2623]_  = ~\new_[2697]_  | ~\new_[4349]_ ;
  assign \new_[2624]_  = \new_[2718]_  | \new_[2676]_ ;
  assign \new_[2625]_  = ~u0_u0_ch_stop_reg;
  assign \new_[2626]_  = ~\new_[2837]_  & ~\new_[4328]_ ;
  assign \new_[2627]_  = ~\new_[2663]_ ;
  assign \new_[2628]_  = ~\new_[2856]_  & ~\new_[4328]_ ;
  assign \new_[2629]_  = ~\new_[4210]_  | ~\new_[2670]_  | ~\new_[3594]_ ;
  assign \new_[2630]_  = \new_[2758]_  & \new_[1339]_ ;
  assign \new_[2631]_  = \new_[2758]_  ^ \new_[1339]_ ;
  assign \new_[2632]_  = ~\new_[3999]_  & ~\new_[4343]_ ;
  assign \new_[2633]_  = u0_u0_ch_sz_inf_reg;
  assign \new_[2634]_  = \\u1_u1_state_reg[2] ;
  assign \new_[2635]_  = \\u1_u1_state_reg[3] ;
  assign \new_[2636]_  = ~\\u0_u0_ch_chk_sz_r_reg[5] ;
  assign \new_[2637]_  = \\u0_u0_ch_chk_sz_r_reg[3] ;
  assign \new_[2638]_  = ~\\u0_u0_ch_chk_sz_r_reg[7] ;
  assign \new_[2639]_  = \\u0_u0_ch_chk_sz_r_reg[1] ;
  assign \new_[2640]_  = \\u0_u0_ch_chk_sz_r_reg[2] ;
  assign \new_[2641]_  = \\u1_u1_state_reg[4] ;
  assign \new_[2642]_  = \\u0_u0_ch_chk_sz_r_reg[4] ;
  assign \new_[2643]_  = ~\\u0_u0_ch_chk_sz_r_reg[6] ;
  assign \new_[2644]_  = ~\\u0_u0_ch_chk_sz_r_reg[0] ;
  assign \new_[2645]_  = \\u1_u1_state_reg[0] ;
  assign \new_[2646]_  = ~\new_[2673]_ ;
  assign \new_[2647]_  = \new_[2759]_  ^ \new_[1238]_ ;
  assign \new_[2648]_  = \\u1_u1_state_reg[1] ;
  assign \new_[2649]_  = u4_u1_rf_ack_reg;
  assign \new_[2650]_  = ~\\u0_u0_ch_chk_sz_r_reg[10] ;
  assign \new_[2651]_  = ~\\u0_u0_ch_chk_sz_r_reg[8] ;
  assign \new_[2652]_  = ~\\u0_u0_ch_chk_sz_r_reg[9] ;
  assign \new_[2653]_  = \new_[2933]_  & \new_[2701]_ ;
  assign \new_[2654]_  = ~\new_[2674]_ ;
  assign \new_[2655]_  = ~\new_[2697]_  | ~\new_[4210]_ ;
  assign \new_[2656]_  = ~\new_[3630]_  | ~\new_[2730]_ ;
  assign \new_[2657]_  = ~\new_[4243]_  | ~\new_[3722]_ ;
  assign \new_[2658]_  = ~\new_[2730]_  | ~\new_[3640]_ ;
  assign \new_[2659]_  = ~\new_[3682]_  | ~\new_[4243]_ ;
  assign n2296 = ~\new_[2675]_ ;
  assign \new_[2661]_  = ~\new_[2746]_  & ~\new_[2852]_ ;
  assign \new_[2662]_  = ~\new_[2746]_  & ~\new_[2793]_ ;
  assign \new_[2663]_  = ~\new_[2857]_  & ~\new_[4325]_ ;
  assign \new_[2664]_  = ~\new_[2678]_ ;
  assign \new_[2665]_  = ~\new_[2749]_  & ~\new_[4383]_ ;
  assign \new_[2666]_  = ~\new_[2679]_ ;
  assign \new_[2667]_  = ~\new_[2680]_ ;
  assign \new_[2668]_  = ~\new_[4244]_  & ~\new_[2749]_ ;
  assign \new_[2669]_  = ~\new_[2748]_  | ~\new_[2747]_ ;
  assign \new_[2670]_  = ~\new_[2697]_ ;
  assign \new_[2671]_  = \\u2_u0_out_r_reg[15] ;
  assign \new_[2672]_  = \\u2_u1_out_r_reg[15] ;
  assign \new_[2673]_  = ~\new_[2759]_  | ~\new_[1238]_ ;
  assign \new_[2674]_  = ~\new_[4343]_ ;
  assign \new_[2675]_  = ~\new_[2820]_  & (~\new_[3610]_  | ~\new_[3212]_ );
  assign \new_[2676]_  = ~\new_[3431]_  & ~\new_[2793]_ ;
  assign \new_[2677]_  = ~\new_[2938]_  & ~\new_[2794]_ ;
  assign \new_[2678]_  = ~\new_[4385]_  | ~\new_[2815]_ ;
  assign \new_[2679]_  = ~\new_[4387]_  | ~\new_[4207]_  | ~\new_[2913]_  | ~\new_[2838]_ ;
  assign \new_[2680]_  = ~\new_[2817]_  | ~\new_[2816]_ ;
  assign \new_[2681]_  = \new_[3627]_  ? \new_[2836]_  : \new_[3628]_ ;
  assign n2326 = \new_[4076]_  ? \new_[2827]_  : \new_[3936]_ ;
  assign \new_[2683]_  = ~\new_[2813]_  | (~\new_[4368]_  & ~\new_[3690]_ );
  assign n2336 = \new_[2609]_  ? \new_[2827]_  : \new_[3938]_ ;
  assign n2306 = \new_[2601]_  ? \new_[2827]_  : \new_[3932]_ ;
  assign n2341 = \new_[2610]_  ? \new_[2827]_  : \new_[3884]_ ;
  assign n2301 = \new_[2600]_  ? \new_[2827]_  : \new_[3899]_ ;
  assign n2321 = ~\new_[2766]_  | (~\new_[2873]_  & ~\new_[3895]_ );
  assign n2346 = ~\new_[2767]_  | (~\new_[2873]_  & ~\new_[3904]_ );
  assign n2316 = (~\new_[2873]_  & ~\new_[3886]_ ) | (~\new_[2827]_  & ~\new_[4013]_ );
  assign n2331 = \new_[4127]_  ? \new_[2827]_  : \new_[3923]_ ;
  assign \new_[2692]_  = ~\new_[2814]_  | (~\new_[2837]_  & ~\new_[3654]_ );
  assign n2311 = \new_[4016]_  ? \new_[2827]_  : \new_[3946]_ ;
  assign \new_[2694]_  = \new_[3639]_  ? \new_[2837]_  : \new_[3637]_ ;
  assign n2351 = ~\new_[2768]_  | (~\new_[2873]_  & ~\new_[3920]_ );
  assign n2356 = ~\new_[2873]_  & ~\new_[3926]_ ;
  assign \new_[2697]_  = ~\new_[2751]_ ;
  assign \new_[2698]_  = \\u2_state_reg[8] ;
  assign \new_[2699]_  = \\u2_state_reg[7] ;
  assign \new_[2700]_  = \\u2_state_reg[6] ;
  assign \new_[2701]_  = ~\new_[2938]_  & ~\new_[2853]_ ;
  assign \new_[2702]_  = ~\new_[2939]_  & ~\new_[3919]_ ;
  assign \new_[2703]_  = \new_[2939]_  & \new_[4093]_ ;
  assign \new_[2704]_  = ~\new_[2939]_  & ~\new_[3875]_ ;
  assign \new_[2705]_  = ~\new_[2939]_  & ~\new_[3930]_ ;
  assign \new_[2706]_  = \new_[2939]_  & \new_[3976]_ ;
  assign \new_[2707]_  = \new_[2939]_  & \new_[4001]_ ;
  assign \new_[2708]_  = \new_[2939]_  & \new_[4020]_ ;
  assign \new_[2709]_  = \new_[2939]_  & \new_[4162]_ ;
  assign \new_[2710]_  = \new_[2939]_  & \new_[4050]_ ;
  assign \new_[2711]_  = ~\new_[2939]_  & ~\new_[3886]_ ;
  assign \new_[2712]_  = ~\new_[2939]_  & ~\new_[3920]_ ;
  assign \new_[2713]_  = \new_[2939]_  & \new_[4153]_ ;
  assign \new_[2714]_  = ~\new_[2939]_  & ~\new_[3904]_ ;
  assign \new_[2715]_  = ~\new_[2939]_  & ~\new_[3934]_ ;
  assign \new_[2716]_  = \new_[2939]_  & \new_[3967]_ ;
  assign n2431 = ~\new_[2760]_ ;
  assign \new_[2718]_  = ~\new_[3430]_  & ~\new_[2852]_ ;
  assign n2421 = \new_[2991]_  | \new_[3068]_  | \new_[2985]_  | \new_[2995]_ ;
  assign n2426 = \new_[2986]_  | \new_[2996]_  | \new_[2992]_  | \new_[3069]_ ;
  assign n2366 = \new_[2993]_  | \new_[3070]_  | \new_[2987]_  | \new_[2997]_ ;
  assign n2371 = \new_[2988]_  | \new_[2998]_  | \new_[2994]_  | \new_[3071]_ ;
  assign n2401 = \new_[2990]_  | \new_[3072]_  | \new_[2989]_  | \new_[2999]_ ;
  assign \new_[2724]_  = \new_[2939]_  & \new_[4285]_ ;
  assign \new_[2725]_  = ~\new_[2939]_  & ~\new_[3943]_ ;
  assign \new_[2726]_  = \new_[2939]_  & \new_[4087]_ ;
  assign \new_[2727]_  = ~\new_[2939]_  & ~\new_[3895]_ ;
  assign \new_[2728]_  = ~\new_[2939]_  & ~\new_[3926]_ ;
  assign \new_[2729]_  = ~\new_[4244]_  & ~\new_[4325]_ ;
  assign \new_[2730]_  = ~\new_[4350]_  & ~\new_[2857]_ ;
  assign n2416 = \new_[3946]_  ? \new_[2883]_  : \new_[4015]_ ;
  assign n2386 = \new_[3925]_  ? \new_[2883]_  : \new_[4108]_ ;
  assign n2391 = \new_[3932]_  ? \new_[2883]_  : \new_[2639]_ ;
  assign n2396 = \new_[3884]_  ? \new_[2883]_  : \new_[2640]_ ;
  assign n2381 = \new_[3899]_  ? \new_[2883]_  : \new_[2637]_ ;
  assign n2376 = \new_[3927]_  ? \new_[2883]_  : \new_[4062]_ ;
  assign n2411 = \new_[3952]_  ? \new_[2883]_  : \new_[4085]_ ;
  assign n2441 = \new_[3896]_  ? \new_[2883]_  : \new_[4081]_ ;
  assign n2446 = \new_[3928]_  ? \new_[2883]_  : \new_[4000]_ ;
  assign n2361 = \new_[3936]_  ? \new_[2883]_  : \new_[2633]_ ;
  assign \new_[2741]_  = \new_[3641]_  ? \new_[4368]_  : \new_[3715]_ ;
  assign \new_[2742]_  = \new_[3714]_  ? \new_[4368]_  : \new_[3634]_ ;
  assign n2436 = \new_[3912]_  ? \new_[2883]_  : \new_[4017]_ ;
  assign n2406 = \new_[3906]_  ? \new_[2883]_  : \new_[2642]_ ;
  assign \new_[2745]_  = ~\new_[2793]_ ;
  assign \new_[2746]_  = ~\new_[2794]_ ;
  assign \new_[2747]_  = ~\new_[2835]_  | ~\new_[3678]_ ;
  assign \new_[2748]_  = ~\new_[2837]_  | ~\new_[3712]_ ;
  assign \new_[2749]_  = ~\new_[2818]_ ;
  assign \new_[2750]_  = ~\new_[2822]_ ;
  assign \new_[2751]_  = ~\new_[2837]_ ;
  assign n2451 = \new_[1416]_  ^ \new_[3003]_ ;
  assign n2456 = \new_[1251]_  ^ \new_[3002]_ ;
  assign \new_[2754]_  = \\u2_u0_out_r_reg[11] ;
  assign \new_[2755]_  = \\u2_u1_out_r_reg[11] ;
  assign \new_[2756]_  = \\u2_u0_out_r_reg[12] ;
  assign \new_[2757]_  = \\u2_u1_out_r_reg[12] ;
  assign \new_[2758]_  = \\u2_u0_out_r_reg[16] ;
  assign \new_[2759]_  = \\u2_u1_out_r_reg[16] ;
  assign \new_[2760]_  = ~wb1_cyc_i | ~\new_[2937]_  | ~wb1_stb_i;
  assign \new_[2761]_  = ~\new_[4351]_  | ~\new_[4345]_ ;
  assign \new_[2762]_  = ~\new_[2940]_  & (~\new_[3848]_  | ~\new_[1699]_ );
  assign \new_[2763]_  = ~\new_[4272]_  & ~\new_[3934]_ ;
  assign \new_[2764]_  = \new_[4272]_  & \new_[4083]_ ;
  assign \new_[2765]_  = ~\new_[4272]_  & ~\new_[3895]_ ;
  assign \new_[2766]_  = ~\new_[2873]_  | ~\new_[2604]_ ;
  assign \new_[2767]_  = ~\new_[2873]_  | ~\new_[2611]_ ;
  assign \new_[2768]_  = ~\new_[2873]_  | ~\new_[2612]_ ;
  assign \new_[2769]_  = ~\new_[2944]_  | ~\new_[4073]_ ;
  assign \new_[2770]_  = ~\new_[2883]_  & ~\new_[3943]_ ;
  assign \new_[2771]_  = \new_[2883]_  & \new_[4281]_ ;
  assign \new_[2772]_  = ~\new_[2883]_  & ~\new_[3934]_ ;
  assign \new_[2773]_  = \new_[2883]_  & \new_[4088]_ ;
  assign \new_[2774]_  = ~\new_[2883]_  & ~\new_[3919]_ ;
  assign \new_[2775]_  = \new_[2883]_  & \new_[4266]_ ;
  assign \new_[2776]_  = ~\new_[2883]_  & ~\new_[3930]_ ;
  assign \new_[2777]_  = \new_[2883]_  & \new_[3998]_ ;
  assign \new_[2778]_  = ~\new_[2883]_  & ~\new_[3875]_ ;
  assign \new_[2779]_  = \new_[2883]_  & \new_[3996]_ ;
  assign \new_[2780]_  = ~\new_[2883]_  & ~\new_[3895]_ ;
  assign \new_[2781]_  = \new_[2883]_  & \new_[4021]_ ;
  assign \new_[2782]_  = ~\new_[2883]_  & ~\new_[3904]_ ;
  assign \new_[2783]_  = \new_[2883]_  & \new_[4104]_ ;
  assign \new_[2784]_  = ~\new_[2883]_  & ~\new_[3886]_ ;
  assign \new_[2785]_  = \new_[2883]_  & \new_[4012]_ ;
  assign \new_[2786]_  = ~\new_[2883]_  & ~\new_[3920]_ ;
  assign \new_[2787]_  = \new_[2883]_  & \new_[4112]_ ;
  assign \new_[2788]_  = ~\new_[2883]_  & ~\new_[3926]_ ;
  assign \new_[2789]_  = \new_[2883]_  & \new_[4101]_ ;
  assign \new_[2790]_  = ~\new_[2944]_  | ~\new_[4055]_ ;
  assign \new_[2791]_  = ~\new_[2944]_  | ~\new_[4072]_ ;
  assign \new_[2792]_  = ~\new_[2944]_  | ~\new_[4184]_ ;
  assign \new_[2793]_  = \new_[3199]_  | \new_[3084]_ ;
  assign \new_[2794]_  = ~\new_[2853]_ ;
  assign \new_[2795]_  = ~\new_[4272]_  & ~\new_[3919]_ ;
  assign \new_[2796]_  = \new_[4272]_  & \new_[3961]_ ;
  assign \new_[2797]_  = \new_[2873]_  | \new_[3882]_ ;
  assign \new_[2798]_  = ~\new_[4272]_  & ~\new_[3930]_ ;
  assign \new_[2799]_  = \new_[4272]_  & \new_[4032]_ ;
  assign \new_[2800]_  = ~\new_[4272]_  & ~\new_[3875]_ ;
  assign \new_[2801]_  = \new_[4272]_  & \new_[4121]_ ;
  assign \new_[2802]_  = \new_[4272]_  & \new_[4045]_ ;
  assign \new_[2803]_  = ~\new_[4272]_  & ~\new_[3904]_ ;
  assign \new_[2804]_  = \new_[4272]_  & \new_[4043]_ ;
  assign \new_[2805]_  = ~\new_[4272]_  & ~\new_[3886]_ ;
  assign \new_[2806]_  = \new_[4272]_  & \new_[3984]_ ;
  assign \new_[2807]_  = ~\new_[4272]_  & ~\new_[3920]_ ;
  assign \new_[2808]_  = \new_[4272]_  & \new_[4180]_ ;
  assign \new_[2809]_  = ~\new_[4272]_  & ~\new_[3926]_ ;
  assign \new_[2810]_  = \new_[4272]_  & \new_[4100]_ ;
  assign \new_[2811]_  = ~\new_[4272]_  & ~\new_[3943]_ ;
  assign \new_[2812]_  = \new_[4272]_  & \new_[3975]_ ;
  assign \new_[2813]_  = ~\new_[2900]_  | ~\new_[3716]_ ;
  assign \new_[2814]_  = ~\new_[2900]_  | ~\new_[3631]_ ;
  assign \new_[2815]_  = ~\new_[2856]_ ;
  assign \new_[2816]_  = ~\new_[2856]_ ;
  assign \new_[2817]_  = ~\new_[2857]_ ;
  assign \new_[2818]_  = ~\new_[2858]_ ;
  assign \new_[2819]_  = ~\new_[4244]_ ;
  assign \new_[2820]_  = ~\new_[2917]_  | (~\new_[3550]_  & ~\new_[3244]_ );
  assign \new_[2821]_  = ~\new_[3192]_  | ~\new_[3085]_  | ~\new_[3088]_  | ~\new_[3191]_ ;
  assign \new_[2822]_  = ~\new_[2939]_ ;
  assign \new_[2823]_  = ~\new_[3077]_  & (~\new_[3307]_  | ~\new_[1701]_ );
  assign \new_[2824]_  = ~\new_[3079]_  & (~\new_[3307]_  | ~\new_[1240]_ );
  assign \new_[2825]_  = ~\new_[3080]_  & (~\new_[3307]_  | ~\new_[1241]_ );
  assign \new_[2826]_  = ~\new_[3074]_  & (~\new_[3307]_  | ~\new_[1246]_ );
  assign \new_[2827]_  = ~\new_[2873]_ ;
  assign \new_[2828]_  = ~\new_[3079]_  & (~\new_[3307]_  | ~\new_[1695]_ );
  assign \new_[2829]_  = ~\new_[3080]_  & (~\new_[3307]_  | ~\new_[1696]_ );
  assign \new_[2830]_  = ~\new_[3081]_  & (~\new_[3307]_  | ~\new_[1697]_ );
  assign \new_[2831]_  = ~\\u0_int_maska_r_reg[11] ;
  assign \new_[2832]_  = \\u0_csr_r_reg[0] ;
  assign \new_[2833]_  = \\u0_int_maska_r_reg[0] ;
  assign \new_[2834]_  = ~\new_[4368]_ ;
  assign \new_[2835]_  = ~\new_[2900]_ ;
  assign \new_[2836]_  = ~\new_[2912]_ ;
  assign \new_[2837]_  = ~\new_[2912]_ ;
  assign \new_[2838]_  = ~\new_[2914]_ ;
  assign \new_[2839]_  = \\u2_u0_out_r_reg[14] ;
  assign \new_[2840]_  = \\u2_u1_out_r_reg[14] ;
  assign \new_[2841]_  = ~\\u0_int_maska_r_reg[10] ;
  assign \new_[2842]_  = ~\\u0_int_maska_r_reg[5] ;
  assign n2466 = \new_[3025]_  | \new_[3101]_ ;
  assign n2461 = ~\new_[3021]_  | (~\new_[3578]_  & ~\new_[3132]_ );
  assign n2471 = ~\new_[3020]_  | (~\new_[3611]_  & ~\new_[3193]_ );
  assign \new_[2846]_  = ~\new_[3894]_  | ~\new_[3015]_  | ~\new_[4065]_ ;
  assign \new_[2847]_  = \\u2_u1_out_r_reg[8] ;
  assign \new_[2848]_  = \\u2_u0_out_r_reg[8] ;
  assign \new_[2849]_  = \new_[3189]_  | \new_[4255]_  | \new_[3364]_  | \new_[4259]_ ;
  assign \new_[2850]_  = ~\new_[3911]_  | ~\new_[3029]_  | ~\new_[2832]_ ;
  assign \new_[2851]_  = ~\\u0_int_maska_r_reg[6] ;
  assign \new_[2852]_  = ~\new_[2933]_ ;
  assign \new_[2853]_  = ~\new_[3246]_  & ~\new_[2984]_ ;
  assign \new_[2854]_  = ~\\u0_int_maska_r_reg[7] ;
  assign \new_[2855]_  = ~\new_[4350]_ ;
  assign \new_[2856]_  = ~\new_[4207]_  | ~\new_[4315]_ ;
  assign \new_[2857]_  = ~\new_[3000]_  | ~\new_[4353]_ ;
  assign \new_[2858]_  = ~\new_[4388]_  | ~\new_[4348]_ ;
  assign \new_[2859]_  = \new_[2938]_ ;
  assign \new_[2860]_  = ~\\u0_int_maska_r_reg[8] ;
  assign \new_[2861]_  = ~\\u0_int_maska_r_reg[9] ;
  assign \new_[2862]_  = ~\new_[3085]_  | (~\new_[3094]_  & ~\new_[3826]_ );
  assign \new_[2863]_  = ~\\u0_int_maska_r_reg[2] ;
  assign \new_[2864]_  = ~\new_[3077]_  & (~\new_[3307]_  | ~\new_[4066]_ );
  assign \new_[2865]_  = ~\new_[3775]_  | (~\new_[3195]_  & ~\new_[3880]_ );
  assign \new_[2866]_  = ~\new_[3168]_  & (~\new_[3307]_  | ~\new_[1231]_ );
  assign \new_[2867]_  = ~\new_[3174]_  & (~\new_[3307]_  | ~\new_[1284]_ );
  assign \new_[2868]_  = ~\new_[3078]_  & (~\new_[3307]_  | ~\new_[1239]_ );
  assign \new_[2869]_  = ~\new_[3075]_  & (~\new_[3307]_  | ~\new_[1702]_ );
  assign \new_[2870]_  = ~\new_[3081]_  & (~\new_[3307]_  | ~\new_[4154]_ );
  assign \new_[2871]_  = ~\new_[3073]_  & (~\new_[3307]_  | ~\new_[1698]_ );
  assign \new_[2872]_  = ~\new_[3074]_  & (~\new_[3307]_  | ~\new_[1699]_ );
  assign \new_[2873]_  = ~\new_[3743]_  | ~\new_[4273]_  | ~\new_[3725]_ ;
  assign \new_[2874]_  = ~\new_[3076]_  & (~\new_[3307]_  | ~\new_[1659]_ );
  assign \new_[2875]_  = ~\new_[3178]_  & (~\new_[3307]_  | ~\new_[1378]_ );
  assign \new_[2876]_  = ~\new_[3078]_  & (~\new_[3307]_  | ~\new_[1694]_ );
  assign \new_[2877]_  = ~\new_[3082]_  & (~\new_[3307]_  | ~\new_[1657]_ );
  assign \new_[2878]_  = ~\\u0_int_maska_r_reg[4] ;
  assign \new_[2879]_  = ~\new_[3082]_  & (~\new_[3307]_  | ~\new_[3989]_ );
  assign \new_[2880]_  = ~\new_[3076]_  & (~\new_[3307]_  | ~\new_[3973]_ );
  assign \new_[2881]_  = ~\new_[3073]_  & (~\new_[3307]_  | ~\new_[1245]_ );
  assign \new_[2882]_  = ~\\u0_int_maska_r_reg[3] ;
  assign \new_[2883]_  = ~\new_[3470]_  | ~\new_[4273]_ ;
  assign \new_[2884]_  = ~\new_[3077]_  & (~\new_[3307]_  | ~\new_[4069]_ );
  assign \new_[2885]_  = ~\new_[3168]_  & (~\new_[3307]_  | ~\new_[3935]_ );
  assign \new_[2886]_  = ~\new_[3075]_  & (~\new_[3307]_  | ~\new_[1244]_ );
  assign \new_[2887]_  = ~\new_[3174]_  & (~\new_[3307]_  | ~\new_[1373]_ );
  assign \new_[2888]_  = ~\new_[3078]_  & (~\new_[3307]_  | ~\new_[1383]_ );
  assign \new_[2889]_  = ~\new_[3079]_  & (~\new_[3307]_  | ~\new_[1384]_ );
  assign \new_[2890]_  = ~\new_[3080]_  & (~\new_[3307]_  | ~\new_[1389]_ );
  assign \new_[2891]_  = ~\new_[3081]_  & (~\new_[3307]_  | ~\new_[4082]_ );
  assign \new_[2892]_  = ~\new_[3082]_  & (~\new_[3307]_  | ~\new_[4185]_ );
  assign \new_[2893]_  = ~\new_[3075]_  & (~\new_[3307]_  | ~\new_[1388]_ );
  assign \new_[2894]_  = ~\\u0_int_maska_r_reg[29] ;
  assign \new_[2895]_  = ~\\u0_int_maska_r_reg[26] ;
  assign \new_[2896]_  = ~\new_[3073]_  & (~\new_[3307]_  | ~\new_[1387]_ );
  assign \new_[2897]_  = ~\\u0_int_maska_r_reg[27] ;
  assign \new_[2898]_  = ~\\u0_int_maska_r_reg[28] ;
  assign \new_[2899]_  = ~\\u0_int_maska_r_reg[19] ;
  assign \new_[2900]_  = \new_[4369]_ ;
  assign \new_[2901]_  = ~\\u0_int_maska_r_reg[22] ;
  assign \new_[2902]_  = ~\\u0_int_maska_r_reg[24] ;
  assign \new_[2903]_  = ~\\u0_int_maska_r_reg[23] ;
  assign \new_[2904]_  = ~\\u0_int_maska_r_reg[1] ;
  assign \new_[2905]_  = ~\\u0_int_maska_r_reg[20] ;
  assign \new_[2906]_  = ~\\u0_int_maska_r_reg[16] ;
  assign \new_[2907]_  = ~\\u0_int_maska_r_reg[17] ;
  assign \new_[2908]_  = ~\\u0_int_maska_r_reg[15] ;
  assign \new_[2909]_  = ~\\u0_int_maska_r_reg[12] ;
  assign \new_[2910]_  = ~\\u0_int_maska_r_reg[13] ;
  assign \new_[2911]_  = ~\\u0_int_maska_r_reg[14] ;
  assign \new_[2912]_  = ~\new_[4369]_ ;
  assign \new_[2913]_  = ~\new_[3000]_ ;
  assign \new_[2914]_  = ~\new_[4245]_ ;
  assign n2476 = \new_[1377]_  ^ \new_[3209]_ ;
  assign \new_[2916]_  = ~\new_[3001]_ ;
  assign \new_[2917]_  = ~\new_[3090]_  | ~\new_[3610]_ ;
  assign \new_[2918]_  = ~\new_[3093]_  & (~\new_[3848]_  | ~\new_[1697]_ );
  assign \new_[2919]_  = ~\new_[3095]_  & (~\new_[3848]_  | ~\new_[1698]_ );
  assign \new_[2920]_  = ~\\u0_int_maskb_r_reg[6] ;
  assign \new_[2921]_  = ~\\u0_int_maskb_r_reg[9] ;
  assign \new_[2922]_  = \\u2_u1_out_r_reg[7] ;
  assign \new_[2923]_  = \\u2_u0_out_r_reg[7] ;
  assign \new_[2924]_  = ~\\u0_int_maska_r_reg[18] ;
  assign \new_[2925]_  = ~\\u0_int_maska_r_reg[21] ;
  assign \new_[2926]_  = ~\\u0_int_maska_r_reg[25] ;
  assign \new_[2927]_  = ~\\u0_int_maska_r_reg[30] ;
  assign \new_[2928]_  = \\u0_int_maskb_r_reg[0] ;
  assign \new_[2929]_  = ~\\u0_int_maskb_r_reg[7] ;
  assign \new_[2930]_  = ~\\u0_int_maskb_r_reg[8] ;
  assign \new_[2931]_  = ~\new_[3105]_  & (~\new_[2832]_  | ~\new_[4077]_ );
  assign \new_[2932]_  = ~\\u0_int_maskb_r_reg[5] ;
  assign \new_[2933]_  = ~\new_[3056]_  & ~\new_[3084]_ ;
  assign n2486 = \new_[1378]_  ^ \new_[3157]_ ;
  assign n2491 = \new_[1287]_  ^ \new_[3158]_ ;
  assign \new_[2936]_  = \new_[3199]_  & \new_[3084]_ ;
  assign \new_[2937]_  = ~\new_[2649]_  & (~\new_[3156]_  | ~\new_[4086]_ );
  assign \new_[2938]_  = ~\new_[3180]_  | ~\new_[3201]_  | ~\new_[3190]_ ;
  assign \new_[2939]_  = ~\new_[3846]_  | ~\new_[3743]_  | ~\new_[4273]_  | ~\new_[3861]_ ;
  assign \new_[2940]_  = ~\new_[3089]_  & ~\new_[3848]_ ;
  assign n2481 = \new_[1248]_  ^ \new_[3208]_ ;
  assign n2496 = ~\new_[3049]_ ;
  assign n2501 = ~\new_[3050]_ ;
  assign \new_[2944]_  = ~\new_[3202]_  | ~\new_[3083]_  | ~\new_[3743]_ ;
  assign \new_[2945]_  = ~\\u0_int_maskb_r_reg[11] ;
  assign \new_[2946]_  = ~\new_[3074]_  & (~\new_[3307]_  | ~\new_[1345]_ );
  assign \new_[2947]_  = ~\new_[3076]_  & (~\new_[3307]_  | ~\new_[3997]_ );
  assign \new_[2948]_  = ~\\u0_int_maskb_r_reg[10] ;
  assign \new_[2949]_  = ~\new_[3178]_  & (~\new_[3307]_  | ~\new_[1287]_ );
  assign \new_[2950]_  = ~\new_[3162]_  & (~\new_[3307]_  | ~\new_[1250]_ );
  assign \new_[2951]_  = ~\new_[3166]_  & (~\new_[3307]_  | ~\new_[1233]_ );
  assign \new_[2952]_  = ~\new_[3173]_  & (~\new_[3307]_  | ~\new_[1234]_ );
  assign \new_[2953]_  = ~\new_[3205]_  & (~\new_[3848]_  | ~\new_[1696]_ );
  assign n2546 = ~\new_[3183]_  | (~\new_[3322]_  & ~\new_[1387]_ );
  assign \new_[2955]_  = ~\new_[3169]_  & (~\new_[3307]_  | ~\new_[1237]_ );
  assign \new_[2956]_  = ~\new_[3170]_  & (~\new_[3307]_  | ~\new_[1285]_ );
  assign \new_[2957]_  = ~\new_[3171]_  & (~\new_[3307]_  | ~\new_[1229]_ );
  assign n2541 = ~\new_[3185]_  | (~\new_[3321]_  & ~\new_[1245]_ );
  assign \new_[2959]_  = ~\new_[3172]_  & (~\new_[3307]_  | ~\new_[3959]_ );
  assign \new_[2960]_  = ~\new_[3176]_  & (~\new_[3307]_  | ~\new_[3994]_ );
  assign \new_[2961]_  = ~\new_[3167]_  & (~\new_[3307]_  | ~\new_[1232]_ );
  assign \new_[2962]_  = ~\new_[3161]_  & (~\new_[3307]_  | ~\new_[1249]_ );
  assign \new_[2963]_  = ~\new_[3175]_  & (~\new_[3307]_  | ~\new_[1370]_ );
  assign \new_[2964]_  = ~\new_[3177]_  & (~\new_[3307]_  | ~\new_[3992]_ );
  assign \new_[2965]_  = ~\new_[3159]_  & (~\new_[3307]_  | ~\new_[1248]_ );
  assign \new_[2966]_  = ~\new_[3177]_  & (~\new_[3307]_  | ~\new_[3987]_ );
  assign \new_[2967]_  = ~\new_[3160]_  & (~\new_[3307]_  | ~\new_[1376]_ );
  assign \new_[2968]_  = ~\new_[3159]_  & (~\new_[3307]_  | ~\new_[1377]_ );
  assign \new_[2969]_  = ~\new_[3165]_  & (~\new_[3307]_  | ~\new_[1236]_ );
  assign \new_[2970]_  = ~\new_[3162]_  & (~\new_[3307]_  | ~\new_[1406]_ );
  assign \new_[2971]_  = ~\new_[3163]_  & (~\new_[3307]_  | ~\new_[4070]_ );
  assign \new_[2972]_  = ~\new_[3164]_  & (~\new_[3307]_  | ~\new_[1339]_ );
  assign \new_[2973]_  = ~\new_[3165]_  & (~\new_[3307]_  | ~\new_[1380]_ );
  assign \new_[2974]_  = ~\new_[3166]_  & (~\new_[3307]_  | ~\new_[1375]_ );
  assign \new_[2975]_  = ~\new_[3167]_  & (~\new_[3307]_  | ~\new_[1414]_ );
  assign \new_[2976]_  = ~\new_[3169]_  & (~\new_[3307]_  | ~\new_[1381]_ );
  assign \new_[2977]_  = ~\new_[3170]_  & (~\new_[3307]_  | ~\new_[1413]_ );
  assign \new_[2978]_  = ~\new_[3171]_  & (~\new_[3307]_  | ~\new_[1372]_ );
  assign \new_[2979]_  = ~\new_[3172]_  & (~\new_[3307]_  | ~\new_[1371]_ );
  assign \new_[2980]_  = ~\new_[3173]_  & (~\new_[3307]_  | ~\new_[1382]_ );
  assign \new_[2981]_  = ~\new_[3176]_  & (~\new_[3307]_  | ~\new_[4011]_ );
  assign \new_[2982]_  = ~\new_[3175]_  & (~\new_[3307]_  | ~\new_[1228]_ );
  assign \new_[2983]_  = ~\new_[3161]_  & (~\new_[3307]_  | ~\new_[1379]_ );
  assign \new_[2984]_  = ~\new_[3186]_  | ~\new_[3187]_ ;
  assign \new_[2985]_  = ~\new_[3347]_  & (~\new_[3252]_  | ~\new_[3308]_ );
  assign \new_[2986]_  = ~\new_[3348]_  & (~\new_[3252]_  | ~\new_[3308]_ );
  assign \new_[2987]_  = ~\new_[3346]_  & (~\new_[3252]_  | ~\new_[3308]_ );
  assign \new_[2988]_  = ~\new_[3344]_  & (~\new_[3252]_  | ~\new_[3308]_ );
  assign \new_[2989]_  = ~\new_[3343]_  & (~\new_[3252]_  | ~\new_[3308]_ );
  assign \new_[2990]_  = ~\new_[3343]_  & (~\new_[3249]_  | ~\new_[3306]_ );
  assign \new_[2991]_  = ~\new_[3347]_  & (~\new_[3249]_  | ~\new_[3306]_ );
  assign \new_[2992]_  = ~\new_[3348]_  & (~\new_[3249]_  | ~\new_[3306]_ );
  assign \new_[2993]_  = ~\new_[3346]_  & (~\new_[3249]_  | ~\new_[3306]_ );
  assign \new_[2994]_  = ~\new_[3344]_  & (~\new_[3249]_  | ~\new_[3306]_ );
  assign \new_[2995]_  = ~\new_[3347]_  & (~\new_[3247]_  | ~\new_[3356]_ );
  assign \new_[2996]_  = ~\new_[3348]_  & (~\new_[3247]_  | ~\new_[3356]_ );
  assign \new_[2997]_  = ~\new_[3346]_  & (~\new_[3247]_  | ~\new_[3356]_ );
  assign \new_[2998]_  = ~\new_[3344]_  & (~\new_[3247]_  | ~\new_[3356]_ );
  assign \new_[2999]_  = ~\new_[3343]_  & (~\new_[3247]_  | ~\new_[3356]_ );
  assign \new_[3000]_  = ~\new_[4352]_ ;
  assign \new_[3001]_  = ~\new_[3084]_ ;
  assign \new_[3002]_  = ~\new_[1250]_  | ~\new_[1249]_  | ~\new_[3208]_  | ~\new_[3870]_ ;
  assign \new_[3003]_  = ~\new_[1406]_  | ~\new_[1379]_  | ~\new_[3209]_  | ~\new_[3956]_ ;
  assign \new_[3004]_  = ~\\u0_int_maskb_r_reg[14] ;
  assign \new_[3005]_  = ~\\u0_int_maskb_r_reg[17] ;
  assign \new_[3006]_  = ~\\u0_int_maskb_r_reg[20] ;
  assign \new_[3007]_  = ~\\u0_int_maskb_r_reg[22] ;
  assign \new_[3008]_  = ~\\u0_int_maskb_r_reg[2] ;
  assign \new_[3009]_  = ~\\u0_int_maskb_r_reg[12] ;
  assign \new_[3010]_  = ~\\u0_int_maskb_r_reg[18] ;
  assign \new_[3011]_  = ~\\u0_int_maskb_r_reg[19] ;
  assign \new_[3012]_  = ~\\u0_int_maskb_r_reg[15] ;
  assign n2521 = ~\new_[3206]_  | (~\new_[3331]_  & ~\new_[1406]_ );
  assign n2526 = ~\new_[3207]_  | (~\new_[3332]_  & ~\new_[1250]_ );
  assign \new_[3015]_  = \new_[3188]_  | \new_[3212]_ ;
  assign \new_[3016]_  = ~\new_[3911]_  | ~\new_[3212]_  | ~\new_[4065]_ ;
  assign \new_[3017]_  = ~\new_[3909]_  | ~\new_[3212]_  | ~\new_[4065]_ ;
  assign \new_[3018]_  = ~\new_[3889]_  | ~\new_[3212]_  | ~\new_[4065]_ ;
  assign \new_[3019]_  = ~\new_[3907]_  | ~\new_[3212]_  | ~\new_[4065]_ ;
  assign \new_[3020]_  = ~\new_[3937]_  | ~\new_[3212]_  | ~\new_[4065]_ ;
  assign \new_[3021]_  = ~\new_[3883]_  | ~\new_[3212]_  | ~\new_[4065]_ ;
  assign \new_[3022]_  = ~\new_[3890]_  | ~\new_[3212]_  | ~\new_[4065]_ ;
  assign \new_[3023]_  = \\u2_u0_out_r_reg[13] ;
  assign \new_[3024]_  = \\u2_u1_out_r_reg[13] ;
  assign \new_[3025]_  = ~\new_[3132]_  & ~\new_[3704]_ ;
  assign \new_[3026]_  = ~\\u0_int_maskb_r_reg[24] ;
  assign \new_[3027]_  = ~\\u0_int_maskb_r_reg[30] ;
  assign \new_[3028]_  = ~\\u0_int_maskb_r_reg[3] ;
  assign \new_[3029]_  = ~\new_[3105]_ ;
  assign \new_[3030]_  = ~\\u0_int_maskb_r_reg[4] ;
  assign \new_[3031]_  = ~\new_[3223]_  & (~\new_[3848]_  | ~\new_[1702]_ );
  assign \new_[3032]_  = ~\\u0_int_maskb_r_reg[25] ;
  assign \new_[3033]_  = ~\\u0_int_maskb_r_reg[28] ;
  assign n2516 = ~\new_[3213]_  | (~\new_[3301]_  & ~\new_[3882]_ );
  assign n2531 = ~\new_[3214]_  | (~\new_[3301]_  & ~\new_[3943]_ );
  assign \new_[3036]_  = ~\\u0_int_maskb_r_reg[29] ;
  assign n2506 = ~\new_[3215]_  | (~\new_[3301]_  & ~\new_[3934]_ );
  assign \new_[3038]_  = ~\\u0_int_maskb_r_reg[26] ;
  assign \new_[3039]_  = ~\\u0_int_maskb_r_reg[27] ;
  assign n2561 = ~\new_[3219]_  | (~\new_[3301]_  & ~\new_[3920]_ );
  assign \new_[3041]_  = ~\\u0_int_maskb_r_reg[23] ;
  assign \new_[3042]_  = ~\\u0_int_maskb_r_reg[1] ;
  assign n2536 = ~\new_[3216]_  | (~\new_[3301]_  & ~\new_[3895]_ );
  assign n2551 = ~\new_[3217]_  | (~\new_[3301]_  & ~\new_[3904]_ );
  assign n2556 = ~\new_[3218]_  | (~\new_[3301]_  & ~\new_[3886]_ );
  assign n2566 = ~\new_[3220]_  | (~\new_[3301]_  & ~\new_[3926]_ );
  assign \new_[3047]_  = ~\\u0_int_maskb_r_reg[21] ;
  assign n2511 = ~\new_[3221]_  | (~\new_[3300]_  & ~\new_[3882]_ );
  assign \new_[3049]_  = ~\new_[4070]_  | ~\new_[1379]_  | ~\new_[3181]_  | ~\new_[1406]_ ;
  assign \new_[3050]_  = ~\new_[4080]_  | ~\new_[1249]_  | ~\new_[3184]_  | ~\new_[1250]_ ;
  assign \new_[3051]_  = ~\\u0_int_maskb_r_reg[16] ;
  assign \new_[3052]_  = ~\\u0_int_maskb_r_reg[13] ;
  assign \new_[3053]_  = ~\new_[3160]_  & (~\new_[3307]_  | ~\new_[1247]_ );
  assign \new_[3054]_  = ~\new_[3163]_  & (~\new_[3307]_  | ~\new_[4080]_ );
  assign \new_[3055]_  = ~\new_[3164]_  & (~\new_[3307]_  | ~\new_[1238]_ );
  assign \new_[3056]_  = ~\new_[3199]_ ;
  assign \new_[3057]_  = ~\new_[3232]_  & (~\new_[3848]_  | ~\new_[1695]_ );
  assign n2726 = ~\new_[3237]_  | (~\new_[3354]_  & ~\new_[3934]_ );
  assign n2731 = ~\new_[3236]_  | (~\new_[3354]_  & ~\new_[3943]_ );
  assign n2706 = ~\new_[3238]_  | (~\new_[3354]_  & ~\new_[3882]_ );
  assign n2721 = ~\new_[3239]_  | (~\new_[3354]_  & ~\new_[3895]_ );
  assign n2666 = ~\new_[3240]_  | (~\new_[3354]_  & ~\new_[3904]_ );
  assign n2711 = ~\new_[3241]_  | (~\new_[3354]_  & ~\new_[3886]_ );
  assign n2716 = ~\new_[3242]_  | (~\new_[3354]_  & ~\new_[3920]_ );
  assign n2671 = ~\new_[3243]_  | (~\new_[3354]_  & ~\new_[3926]_ );
  assign \new_[3066]_  = \new_[3256]_  ? \new_[3307]_  : \new_[1693]_ ;
  assign \new_[3067]_  = \new_[3230]_  ? \new_[3307]_  : \new_[1700]_ ;
  assign \new_[3068]_  = ~\new_[3347]_  & (~\new_[3309]_  | ~\new_[3316]_ );
  assign \new_[3069]_  = ~\new_[3348]_  & (~\new_[3309]_  | ~\new_[3316]_ );
  assign \new_[3070]_  = ~\new_[3346]_  & (~\new_[3309]_  | ~\new_[3316]_ );
  assign \new_[3071]_  = ~\new_[3344]_  & (~\new_[3309]_  | ~\new_[3316]_ );
  assign \new_[3072]_  = ~\new_[3343]_  & (~\new_[3309]_  | ~\new_[3316]_ );
  assign \new_[3073]_  = ~\new_[3307]_  & ~\new_[3960]_ ;
  assign \new_[3074]_  = ~\new_[3307]_  & ~\new_[4103]_ ;
  assign \new_[3075]_  = ~\new_[3307]_  & ~\new_[3962]_ ;
  assign \new_[3076]_  = ~\new_[3307]_  & ~\new_[3979]_ ;
  assign \new_[3077]_  = ~\new_[3307]_  & ~\new_[4025]_ ;
  assign \new_[3078]_  = ~\new_[3307]_  & ~\new_[3970]_ ;
  assign \new_[3079]_  = ~\new_[3307]_  & ~\new_[4029]_ ;
  assign \new_[3080]_  = ~\new_[3307]_  & ~\new_[4124]_ ;
  assign \new_[3081]_  = ~\new_[3307]_  & ~\new_[4131]_ ;
  assign \new_[3082]_  = ~\new_[3307]_  & ~\new_[4027]_ ;
  assign \new_[3083]_  = ~\new_[3180]_ ;
  assign \new_[3084]_  = ~\new_[3725]_  & ~\new_[3251]_ ;
  assign \new_[3085]_  = ~\new_[3534]_  | ~\new_[3879]_  | ~\new_[3257]_  | ~\new_[4199]_ ;
  assign \new_[3086]_  = u2_chunk_cnt_is_0_r_reg;
  assign \new_[3087]_  = ~\new_[3365]_  | ~\new_[3894]_  | ~\new_[3724]_  | ~\new_[3781]_ ;
  assign \new_[3088]_  = ~\new_[3826]_  | ~\new_[3261]_  | ~n3126;
  assign \new_[3089]_  = \new_[1699]_  ^ \new_[3323]_ ;
  assign \new_[3090]_  = ~\new_[3193]_ ;
  assign \new_[3091]_  = \\u2_u1_out_r_reg[4] ;
  assign \new_[3092]_  = \\u2_u0_out_r_reg[4] ;
  assign \new_[3093]_  = ~\new_[3265]_  & ~\new_[3848]_ ;
  assign \new_[3094]_  = ~\new_[3261]_  & ~n3126;
  assign \new_[3095]_  = ~\new_[3280]_  & ~\new_[3848]_ ;
  assign n2681 = \new_[1388]_  ^ \new_[3328]_ ;
  assign n2676 = \new_[1244]_  ^ \new_[3329]_ ;
  assign \new_[3098]_  = \\u2_u1_out_r_reg[10] ;
  assign \new_[3099]_  = \\u2_u0_out_r_reg[10] ;
  assign \new_[3100]_  = \new_[3286]_  | \new_[2832]_ ;
  assign \new_[3101]_  = (~\new_[3615]_  & ~\new_[3318]_ ) | (~\new_[3333]_  & ~\new_[3704]_ );
  assign \new_[3102]_  = ~\new_[3771]_  | (~\new_[3304]_  & ~\new_[3880]_ );
  assign \new_[3103]_  = ~\new_[3883]_  | ~\new_[3293]_  | ~\new_[3854]_ ;
  assign n2646 = \new_[3936]_  ? \new_[3301]_  : \new_[4166]_ ;
  assign \new_[3105]_  = ~\new_[3838]_  | ~\new_[3293]_  | ~\new_[3911]_ ;
  assign n2651 = \new_[3931]_  ? \new_[3301]_  : \new_[4031]_ ;
  assign n2656 = \new_[3938]_  ? \new_[3301]_  : \new_[3968]_ ;
  assign n2661 = \new_[3923]_  ? \new_[3301]_  : \new_[4181]_ ;
  assign n2636 = \new_[3946]_  ? \new_[3301]_  : \new_[4144]_ ;
  assign n2641 = \new_[3932]_  ? \new_[3301]_  : \new_[3964]_ ;
  assign n2686 = \new_[3884]_  ? \new_[3301]_  : \new_[4033]_ ;
  assign n2606 = \new_[3899]_  ? \new_[3301]_  : \new_[4183]_ ;
  assign n2626 = \new_[3897]_  ? \new_[3301]_  : \new_[4146]_ ;
  assign n2691 = \new_[3927]_  ? \new_[3301]_  : \new_[4178]_ ;
  assign n2616 = \new_[3896]_  ? \new_[3301]_  : \new_[4155]_ ;
  assign n2696 = \new_[3928]_  ? \new_[3301]_  : \new_[4036]_ ;
  assign n2591 = \new_[3912]_  ? \new_[3301]_  : \new_[4150]_ ;
  assign n2596 = \new_[3929]_  ? \new_[3301]_  : \new_[4149]_ ;
  assign n2601 = \new_[3915]_  ? \new_[3301]_  : \new_[4008]_ ;
  assign n2586 = \new_[3913]_  ? \new_[3301]_  : \new_[4038]_ ;
  assign n2571 = \new_[3859]_  ? \new_[3301]_  : \new_[4040]_ ;
  assign n2701 = \new_[3910]_  ? \new_[3301]_  : \new_[4039]_ ;
  assign n2581 = \new_[3845]_  ? \new_[3301]_  : \new_[3957]_ ;
  assign n2576 = \new_[3844]_  ? \new_[3301]_  : \new_[4151]_ ;
  assign n2621 = \new_[3925]_  ? \new_[3301]_  : \new_[4035]_ ;
  assign n2611 = \new_[3952]_  ? \new_[3301]_  : \new_[4051]_ ;
  assign n2631 = \new_[3906]_  ? \new_[3301]_  : \new_[4126]_ ;
  assign \new_[3128]_  = \new_[3303]_  ? \new_[3879]_  : \new_[3471]_ ;
  assign \new_[3129]_  = \new_[3303]_  ? \new_[3937]_  : \new_[3471]_ ;
  assign \new_[3130]_  = ~\new_[3222]_ ;
  assign \new_[3131]_  = ~\new_[3224]_ ;
  assign \new_[3132]_  = ~\new_[3879]_  | ~\new_[3297]_  | ~\new_[3658]_ ;
  assign n2781 = ~\new_[3299]_  | (~\new_[3434]_  & ~\new_[1379]_ );
  assign n2786 = ~\new_[3296]_  | (~\new_[3433]_  & ~\new_[1249]_ );
  assign n2736 = \new_[3923]_  ? \new_[3354]_  : \new_[4107]_ ;
  assign n2746 = \new_[3906]_  ? \new_[3354]_  : \new_[4141]_ ;
  assign n2761 = \new_[3931]_  ? \new_[3354]_  : \new_[4019]_ ;
  assign n2851 = \new_[3946]_  ? \new_[3354]_  : \new_[4113]_ ;
  assign n2766 = \new_[3884]_  ? \new_[3354]_  : \new_[4168]_ ;
  assign n2771 = \new_[3899]_  ? \new_[3354]_  : \new_[4174]_ ;
  assign n2846 = \new_[3927]_  ? \new_[3354]_  : \new_[3974]_ ;
  assign n2751 = \new_[3952]_  ? \new_[3354]_  : \new_[4002]_ ;
  assign n2836 = \new_[3925]_  ? \new_[3354]_  : \new_[4097]_ ;
  assign n2811 = \new_[3928]_  ? \new_[3354]_  : \new_[4102]_ ;
  assign n2826 = \new_[3912]_  ? \new_[3354]_  : \new_[4109]_ ;
  assign n2831 = \new_[3929]_  ? \new_[3354]_  : \new_[4106]_ ;
  assign n2816 = \new_[3915]_  ? \new_[3354]_  : \new_[4118]_ ;
  assign n2821 = \new_[3913]_  ? \new_[3354]_  : \new_[4123]_ ;
  assign n2796 = \new_[3910]_  ? \new_[3354]_  : \new_[4116]_ ;
  assign n2801 = \new_[3845]_  ? \new_[3354]_  : \new_[3993]_ ;
  assign n2806 = \new_[3844]_  ? \new_[3354]_  : \new_[4006]_ ;
  assign n2841 = \new_[3897]_  ? \new_[3354]_  : \new_[4084]_ ;
  assign n2741 = \new_[3932]_  ? \new_[3354]_  : \new_[4132]_ ;
  assign n2776 = \new_[3936]_  ? \new_[3354]_  : \new_[3972]_ ;
  assign n2856 = \new_[3938]_  ? \new_[3354]_  : \new_[4172]_ ;
  assign \new_[3156]_  = ~u4_u1_slv_we_reg;
  assign \new_[3157]_  = ~\new_[3322]_  & ~\new_[3733]_ ;
  assign \new_[3158]_  = ~\new_[3321]_  & ~\new_[3731]_ ;
  assign \new_[3159]_  = ~\new_[3307]_  & ~\new_[4054]_ ;
  assign \new_[3160]_  = ~\new_[3307]_  & ~\new_[3969]_ ;
  assign \new_[3161]_  = ~\new_[3307]_  & ~\new_[4009]_ ;
  assign \new_[3162]_  = ~\new_[3307]_  & ~\new_[4157]_ ;
  assign \new_[3163]_  = ~\new_[3307]_  & ~\new_[3977]_ ;
  assign \new_[3164]_  = ~\new_[3307]_  & ~\new_[3983]_ ;
  assign \new_[3165]_  = ~\new_[3307]_  & ~\new_[4170]_ ;
  assign \new_[3166]_  = ~\new_[3307]_  & ~\new_[4028]_ ;
  assign \new_[3167]_  = ~\new_[3307]_  & ~\new_[4137]_ ;
  assign \new_[3168]_  = ~\new_[3307]_  & ~\new_[4111]_ ;
  assign \new_[3169]_  = ~\new_[3307]_  & ~\new_[4024]_ ;
  assign \new_[3170]_  = ~\new_[3307]_  & ~\new_[4136]_ ;
  assign \new_[3171]_  = ~\new_[3307]_  & ~\new_[4135]_ ;
  assign \new_[3172]_  = ~\new_[3307]_  & ~\new_[4003]_ ;
  assign \new_[3173]_  = ~\new_[3307]_  & ~\new_[4079]_ ;
  assign \new_[3174]_  = ~\new_[3307]_  & ~\new_[4023]_ ;
  assign \new_[3175]_  = ~\new_[3307]_  & ~\new_[3965]_ ;
  assign \new_[3176]_  = ~\new_[3307]_  & ~\new_[3958]_ ;
  assign \new_[3177]_  = ~\new_[3307]_  & ~\new_[3971]_ ;
  assign \new_[3178]_  = ~\new_[3307]_  & ~\new_[4171]_ ;
  assign \new_[3179]_  = ~\new_[4077]_  & ~\new_[3318]_  & ~n3126;
  assign \new_[3180]_  = ~\new_[3725]_  | ~\new_[3311]_ ;
  assign \new_[3181]_  = ~\new_[3651]_  & ~\new_[3322]_ ;
  assign \new_[3182]_  = ~\new_[3234]_ ;
  assign \new_[3183]_  = ~\new_[3322]_  | ~\new_[1387]_ ;
  assign \new_[3184]_  = ~\new_[3652]_  & ~\new_[3321]_ ;
  assign \new_[3185]_  = ~\new_[3321]_  | ~\new_[1245]_ ;
  assign \new_[3186]_  = ~\new_[3861]_  | ~\new_[3311]_ ;
  assign \new_[3187]_  = ~\new_[3823]_  | ~\new_[3313]_ ;
  assign \new_[3188]_  = ~\new_[3244]_ ;
  assign \new_[3189]_  = (~\new_[3360]_  | ~\new_[3670]_ ) & (~\new_[3452]_  | ~\new_[4228]_ );
  assign \new_[3190]_  = ~\new_[3315]_  | ~\new_[3871]_ ;
  assign \new_[3191]_  = ~\new_[3455]_  | ~\new_[3398]_ ;
  assign \new_[3192]_  = \new_[3536]_  | \new_[3398]_ ;
  assign \new_[3193]_  = ~\new_[4209]_  | ~\new_[4242]_  | ~\new_[3468]_  | ~\new_[3398]_ ;
  assign \new_[3194]_  = \new_[3325]_  | \new_[3848]_ ;
  assign \new_[3195]_  = \new_[1973]_  ^ \new_[3345]_ ;
  assign n2756 = \new_[3859]_  ? \new_[3354]_  : \new_[4115]_ ;
  assign \new_[3197]_  = \new_[3414]_  ? \new_[3880]_  : \new_[2033]_ ;
  assign \new_[3198]_  = ~\new_[3773]_  | (~\new_[3412]_  & ~\new_[3880]_ );
  assign \new_[3199]_  = \new_[3350]_  ? \new_[3822]_  : \new_[3349]_ ;
  assign n2791 = \new_[3896]_  ? \new_[3354]_  : \new_[3985]_ ;
  assign \new_[3201]_  = ~\new_[3648]_  | ~\new_[3313]_ ;
  assign \new_[3202]_  = u3_u1_slv_re_reg;
  assign \new_[3203]_  = u4_u1_slv_re_reg;
  assign \new_[3204]_  = u3_u1_slv_we_reg;
  assign \new_[3205]_  = ~\new_[3327]_  & ~\new_[3848]_ ;
  assign \new_[3206]_  = ~\new_[3331]_  | ~\new_[1406]_ ;
  assign \new_[3207]_  = ~\new_[3332]_  | ~\new_[1250]_ ;
  assign \new_[3208]_  = \new_[3645]_  & \new_[3329]_ ;
  assign \new_[3209]_  = \new_[3644]_  & \new_[3328]_ ;
  assign \new_[3210]_  = ~\new_[3772]_  | (~\new_[3334]_  & ~\new_[3880]_ );
  assign \new_[3211]_  = \new_[3548]_  | \new_[3333]_ ;
  assign \new_[3212]_  = ~\new_[3333]_  | ~\new_[3318]_ ;
  assign \new_[3213]_  = ~\new_[3301]_  | ~\new_[2833]_ ;
  assign \new_[3214]_  = ~\new_[3301]_  | ~\new_[4143]_ ;
  assign \new_[3215]_  = ~\new_[3301]_  | ~\new_[3963]_ ;
  assign \new_[3216]_  = ~\new_[3301]_  | ~\new_[4042]_ ;
  assign \new_[3217]_  = ~\new_[3301]_  | ~\new_[4041]_ ;
  assign \new_[3218]_  = ~\new_[3301]_  | ~\new_[4094]_ ;
  assign \new_[3219]_  = ~\new_[3301]_  | ~\new_[4152]_ ;
  assign \new_[3220]_  = ~\new_[3301]_  | ~\new_[4095]_ ;
  assign \new_[3221]_  = ~\new_[3300]_  | ~\new_[2832]_ ;
  assign \new_[3222]_  = ~\new_[4077]_  | ~\new_[3298]_  | ~\new_[3745]_ ;
  assign \new_[3223]_  = ~\new_[3305]_  & ~\new_[3848]_ ;
  assign \new_[3224]_  = \new_[3605]_  & \new_[3298]_ ;
  assign \new_[3225]_  = \\u3_u0_mast_dout_reg[4] ;
  assign \new_[3226]_  = \\u3_u0_mast_dout_reg[28] ;
  assign \new_[3227]_  = \\u3_u0_mast_dout_reg[19] ;
  assign \new_[3228]_  = \\u3_u0_mast_dout_reg[29] ;
  assign inta_o = u0_inta_o_reg;
  assign \new_[3230]_  = \\u3_u0_mast_dout_reg[1] ;
  assign \new_[3231]_  = ~\new_[4319]_  | ~\new_[2635]_  | ~\new_[3543]_  | ~\new_[3551]_ ;
  assign \new_[3232]_  = ~\new_[3358]_  & ~\new_[3848]_ ;
  assign \new_[3233]_  = \\u3_u0_mast_dout_reg[8] ;
  assign \new_[3234]_  = ~\new_[3622]_  | ~\new_[3601]_  | ~\new_[3475]_ ;
  assign \new_[3235]_  = \\u3_u0_mast_dout_reg[30] ;
  assign \new_[3236]_  = ~\new_[3354]_  | ~\new_[3986]_ ;
  assign \new_[3237]_  = ~\new_[3354]_  | ~\new_[4167]_ ;
  assign \new_[3238]_  = ~\new_[3354]_  | ~\new_[2928]_ ;
  assign \new_[3239]_  = ~\new_[3354]_  | ~\new_[4105]_ ;
  assign \new_[3240]_  = ~\new_[3354]_  | ~\new_[4049]_ ;
  assign \new_[3241]_  = ~\new_[3354]_  | ~\new_[4140]_ ;
  assign \new_[3242]_  = ~\new_[3354]_  | ~\new_[4099]_ ;
  assign \new_[3243]_  = ~\new_[3354]_  | ~\new_[3980]_ ;
  assign \new_[3244]_  = ~\new_[3475]_  | ~\new_[3601]_  | ~\new_[3746]_ ;
  assign \new_[3245]_  = \\u3_u0_mast_dout_reg[3] ;
  assign \new_[3246]_  = ~\new_[3922]_  & ~\new_[3871]_  & ~\new_[3454]_ ;
  assign \new_[3247]_  = ~\new_[3361]_  & ~\new_[3366]_ ;
  assign \new_[3248]_  = \\u3_u0_mast_dout_reg[22] ;
  assign \new_[3249]_  = ~\new_[3456]_  & ~\new_[3363]_ ;
  assign \new_[3250]_  = \\u3_u0_mast_dout_reg[18] ;
  assign \new_[3251]_  = ~\new_[3311]_ ;
  assign \new_[3252]_  = ~\new_[3362]_  & ~\new_[3462]_ ;
  assign \new_[3253]_  = \\u3_u0_mast_dout_reg[10] ;
  assign \new_[3254]_  = ~\new_[3890]_  | ~\new_[3729]_  | ~\new_[3367]_  | ~\new_[3546]_ ;
  assign \new_[3255]_  = \\u3_u0_mast_dout_reg[12] ;
  assign \new_[3256]_  = \\u3_u0_mast_dout_reg[0] ;
  assign \new_[3257]_  = \new_[3365]_  & \new_[3398]_ ;
  assign n2866 = \new_[1241]_  ^ \new_[3513]_ ;
  assign \new_[3259]_  = \\u3_u0_mast_dout_reg[15] ;
  assign n2871 = \new_[1389]_  ^ \new_[3515]_ ;
  assign \new_[3261]_  = ~\new_[3398]_ ;
  assign \new_[3262]_  = \\u3_u0_mast_dout_reg[20] ;
  assign \new_[3263]_  = \\u3_u0_mast_dout_reg[25] ;
  assign \new_[3264]_  = \\u3_u0_mast_dout_reg[14] ;
  assign \new_[3265]_  = \new_[1697]_  ^ \new_[3497]_ ;
  assign \new_[3266]_  = \\u3_u0_mast_dout_reg[9] ;
  assign \new_[3267]_  = \\u3_u0_mast_dout_reg[13] ;
  assign \new_[3268]_  = \\u3_u0_mast_dout_reg[11] ;
  assign \new_[3269]_  = \\u3_u0_mast_dout_reg[17] ;
  assign \new_[3270]_  = \\u3_u0_mast_dout_reg[2] ;
  assign \new_[3271]_  = \\u2_u1_out_r_reg[3] ;
  assign \new_[3272]_  = \\u3_u0_mast_dout_reg[31] ;
  assign \new_[3273]_  = \\u3_u0_mast_dout_reg[6] ;
  assign \new_[3274]_  = \\u3_u0_mast_dout_reg[27] ;
  assign \new_[3275]_  = \\u3_u0_mast_dout_reg[23] ;
  assign \new_[3276]_  = \\u3_u0_mast_dout_reg[24] ;
  assign intb_o = u0_intb_o_reg;
  assign \new_[3278]_  = \\u2_u0_out_r_reg[3] ;
  assign \new_[3279]_  = \\u3_u0_mast_dout_reg[21] ;
  assign \new_[3280]_  = \new_[1698]_  ^ \new_[3508]_ ;
  assign n2881 = \new_[1376]_  ^ \new_[3426]_ ;
  assign \new_[3282]_  = \\u3_u0_mast_dout_reg[7] ;
  assign n2861 = \new_[3417]_  & \new_[3940]_ ;
  assign \new_[3284]_  = \\u2_u1_out_r_reg[6] ;
  assign \new_[3285]_  = \\u2_u0_out_r_reg[6] ;
  assign \new_[3286]_  = \new_[3909]_  | \new_[4077]_  | \new_[3340]_  | \new_[3889]_ ;
  assign \new_[3287]_  = \\u3_u0_mast_dout_reg[5] ;
  assign \new_[3288]_  = ~\new_[3768]_  | (~\new_[3436]_  & ~\new_[3880]_ );
  assign n2876 = \new_[1247]_  ^ \new_[3427]_ ;
  assign \new_[3290]_  = \\u2_u1_out_r_reg[9] ;
  assign \new_[3291]_  = \\u2_u0_out_r_reg[9] ;
  assign \new_[3292]_  = ~\new_[3796]_  | (~\new_[3510]_  & ~\new_[3880]_ );
  assign \new_[3293]_  = ~\new_[3339]_  & ~\new_[4255]_ ;
  assign \new_[3294]_  = \\u3_u0_mast_dout_reg[26] ;
  assign \new_[3295]_  = \\u3_u0_mast_dout_reg[16] ;
  assign \new_[3296]_  = ~\new_[3433]_  | ~\new_[1249]_ ;
  assign \new_[3297]_  = ~\new_[3339]_ ;
  assign \new_[3298]_  = ~\new_[3340]_ ;
  assign \new_[3299]_  = ~\new_[3434]_  | ~\new_[1379]_ ;
  assign \new_[3300]_  = ~\new_[3743]_  | ~\new_[3545]_  | ~\new_[3535]_ ;
  assign \new_[3301]_  = ~\new_[3822]_  | ~\new_[3545]_  | ~\new_[3535]_ ;
  assign \new_[3302]_  = ~\new_[2029]_  | ~\new_[4329]_ ;
  assign \new_[3303]_  = ~\new_[4242]_  & ~\new_[3868]_  & ~\new_[3432]_  & ~\new_[3894]_ ;
  assign \new_[3304]_  = ~\new_[3429]_  & (~\new_[3638]_  | ~\new_[2068]_ );
  assign \new_[3305]_  = \new_[1702]_  ^ \new_[3539]_ ;
  assign \new_[3306]_  = \new_[3459]_  & \new_[3461]_ ;
  assign \new_[3307]_  = ~\new_[3428]_ ;
  assign \new_[3308]_  = ~\new_[3463]_  & ~\new_[3540]_ ;
  assign \new_[3309]_  = ~\new_[3460]_  & ~\new_[3589]_ ;
  assign n2896 = \new_[3451]_  & \new_[3737]_ ;
  assign \new_[3311]_  = ~\new_[3349]_ ;
  assign n2891 = ~\new_[3453]_  & ~\new_[3792]_ ;
  assign \new_[3313]_  = ~\new_[3350]_ ;
  assign n2886 = ~\new_[3473]_  & ~\new_[3867]_ ;
  assign \new_[3315]_  = ~\new_[3908]_  & ~\new_[3454]_ ;
  assign \new_[3316]_  = ~\new_[3457]_  & (~\new_[3662]_  | ~\new_[3887]_ );
  assign \new_[3317]_  = ~\new_[3355]_ ;
  assign \new_[3318]_  = ~\new_[3705]_  | ~\new_[3937]_  | ~\new_[3465]_  | ~\new_[3601]_ ;
  assign n2901 = ~\new_[3357]_ ;
  assign \new_[3320]_  = ~\new_[3471]_  | ~\new_[4209]_ ;
  assign \new_[3321]_  = ~\new_[3916]_  | ~\new_[1244]_  | ~\new_[3513]_  | ~\new_[1241]_ ;
  assign \new_[3322]_  = ~\new_[3941]_  | ~\new_[1388]_  | ~\new_[3515]_  | ~\new_[1389]_ ;
  assign \new_[3323]_  = ~\new_[3892]_  | ~\new_[3949]_  | ~\new_[3520]_ ;
  assign \new_[3324]_  = \new_[3516]_  | \new_[3848]_ ;
  assign \new_[3325]_  = \new_[1657]_  ^ \new_[3556]_ ;
  assign wb1_ack_o = n3126 ? \new_[3659]_  : \new_[2649]_ ;
  assign \new_[3327]_  = \new_[1696]_  ^ \new_[3577]_ ;
  assign \new_[3328]_  = \new_[3504]_  & \new_[3941]_ ;
  assign \new_[3329]_  = \new_[3517]_  & \new_[3916]_ ;
  assign \new_[3330]_  = ~\new_[3484]_  & (~\new_[3848]_  | ~\new_[1701]_ );
  assign \new_[3331]_  = ~\new_[1378]_  | ~\new_[1379]_  | ~\new_[3426]_  | ~\new_[3954]_ ;
  assign \new_[3332]_  = ~\new_[1287]_  | ~\new_[1249]_  | ~\new_[3427]_  | ~\new_[3874]_ ;
  assign \new_[3333]_  = ~\new_[3706]_  | ~\new_[3854]_  | ~\new_[3467]_  | ~\new_[3526]_ ;
  assign \new_[3334]_  = \new_[1977]_  ^ \new_[3579]_ ;
  assign n3071 = \new_[1243]_  ^ \new_[3581]_ ;
  assign \wb1m_data_o[4]  = ~\new_[4125]_  & ~\new_[3659]_ ;
  assign \wb1m_data_o[13]  = \wb0s_data_i[13]  & \new_[3595]_ ;
  assign \new_[3338]_  = \\u2_u0_out_r_reg[5] ;
  assign \new_[3339]_  = ~\new_[3526]_  | ~\new_[3599]_ ;
  assign \new_[3340]_  = ~\new_[3526]_  | ~\new_[3601]_ ;
  assign n3091 = \new_[1345]_  ^ \new_[3588]_ ;
  assign n3086 = \new_[1246]_  ^ \new_[3608]_ ;
  assign \new_[3343]_  = ~\new_[3537]_  | ~\new_[2641]_ ;
  assign \new_[3344]_  = ~\new_[3537]_  | ~\new_[2635]_ ;
  assign \new_[3345]_  = ~\new_[3917]_  | ~\new_[3945]_  | ~\new_[3619]_ ;
  assign \new_[3346]_  = ~\new_[3537]_  | ~\new_[4053]_ ;
  assign \new_[3347]_  = ~\new_[3537]_  | ~\new_[3887]_ ;
  assign \new_[3348]_  = ~\new_[3537]_  | ~\new_[2648]_ ;
  assign \new_[3349]_  = ~\new_[4335]_  | ~\new_[3933]_ ;
  assign \new_[3350]_  = ~\new_[4335]_  | ~\new_[3847]_ ;
  assign n2926 = ~\new_[3430]_ ;
  assign \wb0_sel_o[1]  = \wb1_sel_i[1]  | \new_[3574]_ ;
  assign n3051 = ~\new_[3431]_ ;
  assign \new_[3354]_  = ~\new_[3908]_  | ~\new_[3204]_  | ~\new_[3538]_  | ~\new_[3823]_ ;
  assign \new_[3355]_  = ~\new_[4329]_ ;
  assign \new_[3356]_  = ~\new_[3541]_  & ~\new_[3544]_ ;
  assign \new_[3357]_  = ~wb0_we_i | ~\new_[4134]_  | ~\new_[3542]_  | ~wb0_stb_i;
  assign \new_[3358]_  = \new_[1695]_  ^ \new_[3593]_ ;
  assign \new_[3359]_  = ~\new_[3573]_  & ~\new_[3612]_ ;
  assign \new_[3360]_  = \new_[4228]_  & \new_[3862]_ ;
  assign \new_[3361]_  = ~\new_[3458]_ ;
  assign \new_[3362]_  = ~\new_[3887]_  & (~\new_[3600]_  | ~\new_[3602]_ );
  assign \new_[3363]_  = ~\new_[3887]_  & (~\new_[3738]_  | ~\new_[3603]_ );
  assign \new_[3364]_  = ~\new_[3546]_  | ~\new_[4077]_ ;
  assign \new_[3365]_  = \new_[3658]_  & \new_[3546]_ ;
  assign \new_[3366]_  = ~\new_[3887]_  & (~\new_[3740]_  | ~\new_[3604]_ );
  assign \new_[3367]_  = \new_[3549]_  & \new_[4199]_ ;
  assign n2916 = \new_[3227]_  ? n3126 : \wb0s_data_i[19] ;
  assign n2931 = \new_[3230]_  ? n3126 : \wb0s_data_i[1] ;
  assign n3096 = \new_[3294]_  ? n3126 : \wb0s_data_i[26] ;
  assign n2961 = \new_[3253]_  ? n3126 : \wb0s_data_i[10] ;
  assign n3016 = \new_[3270]_  ? n3126 : \wb0s_data_i[2] ;
  assign n2976 = \new_[3259]_  ? n3126 : \wb0s_data_i[15] ;
  assign n2991 = \new_[3264]_  ? n3126 : \wb0s_data_i[14] ;
  assign n3031 = \new_[3273]_  ? n3126 : \wb0s_data_i[6] ;
  assign n3011 = \new_[3269]_  ? n3126 : \wb0s_data_i[17] ;
  assign n2936 = \new_[3233]_  ? n3126 : \wb0s_data_i[8] ;
  assign n3001 = \new_[3267]_  ? n3126 : \wb0s_data_i[13] ;
  assign n3046 = \new_[3276]_  ? n3126 : \wb0s_data_i[24] ;
  assign n3006 = \new_[3268]_  ? n3126 : \wb0s_data_i[11] ;
  assign n2946 = \new_[3245]_  ? n3126 : \wb0s_data_i[3] ;
  assign n2996 = \new_[3266]_  ? n3126 : \wb0s_data_i[9] ;
  assign n3041 = \new_[3275]_  ? n3126 : \wb0s_data_i[23] ;
  assign n2941 = \new_[3235]_  ? n3126 : \wb0s_data_i[30] ;
  assign n2986 = \new_[3263]_  ? n3126 : \wb0s_data_i[25] ;
  assign n2951 = \new_[3248]_  ? n3126 : \wb0s_data_i[22] ;
  assign n2981 = \new_[3262]_  ? n3126 : \wb0s_data_i[20] ;
  assign n3026 = \new_[3272]_  ? n3126 : \wb0s_data_i[31] ;
  assign n2911 = \new_[3226]_  ? n3126 : \wb0s_data_i[28] ;
  assign n2971 = \new_[3256]_  ? n3126 : \wb0s_data_i[0] ;
  assign n2966 = \new_[3255]_  ? n3126 : \wb0s_data_i[12] ;
  assign n2956 = \new_[3250]_  ? n3126 : \wb0s_data_i[18] ;
  assign n3101 = \new_[3295]_  ? n3126 : \wb0s_data_i[16] ;
  assign n3066 = \new_[3282]_  ? n3126 : \wb0s_data_i[7] ;
  assign n3036 = \new_[3274]_  ? n3126 : \wb0s_data_i[27] ;
  assign n3061 = \new_[3279]_  ? n3126 : \wb0s_data_i[21] ;
  assign n2921 = \new_[3228]_  ? n3126 : \wb0s_data_i[29] ;
  assign \new_[3398]_  = ~\new_[3894]_  & ~\new_[3937]_ ;
  assign \wb1m_data_o[8]  = \wb0s_data_i[8]  & \new_[3595]_ ;
  assign n3076 = \new_[1386]_  ^ \new_[3580]_ ;
  assign \new_[3401]_  = \\u2_u1_out_r_reg[5] ;
  assign wb0_ack_o = \new_[3840]_  ? \new_[3607]_  : \new_[3478]_ ;
  assign \wb0_sel_o[3]  = \wb1_sel_i[3]  | \new_[3659]_ ;
  assign \wb0_sel_o[2]  = \wb1_sel_i[2]  | \new_[3574]_ ;
  assign \wb0_sel_o[0]  = \wb1_sel_i[0]  | \new_[3574]_ ;
  assign wb1_rty_o = ~\new_[4022]_  & ~\new_[3659]_ ;
  assign \wb1m_data_o[26]  = \wb0s_data_i[26]  & \new_[3595]_ ;
  assign \wb1m_data_o[18]  = \wb0s_data_i[18]  & \new_[3595]_ ;
  assign \wb1m_data_o[14]  = ~\new_[4048]_  & ~\new_[3659]_ ;
  assign \wb1m_data_o[12]  = \wb0s_data_i[12]  & \new_[3595]_ ;
  assign \wb1m_data_o[5]  = \wb0s_data_i[5]  & \new_[3595]_ ;
  assign \new_[3412]_  = \new_[1976]_  ^ \new_[3618]_ ;
  assign \new_[3413]_  = \\u2_u1_out_r_reg[2] ;
  assign \new_[3414]_  = \new_[2033]_  ^ \new_[3619]_ ;
  assign n3081 = \new_[3287]_  ? n3126 : \wb0s_data_i[5] ;
  assign n2906 = \new_[3225]_  ? n3126 : \wb0s_data_i[4] ;
  assign \new_[3417]_  = ~\new_[3527]_  & ~\new_[1977]_ ;
  assign n3021 = \new_[1240]_  ^ \new_[3585]_ ;
  assign n3056 = \new_[1384]_  ^ \new_[3617]_ ;
  assign \new_[3420]_  = \\u2_u0_out_r_reg[2] ;
  assign \new_[3421]_  = ~\wb1m_data_i[20]  | ~\new_[3616]_ ;
  assign \wb1m_data_o[6]  = \wb0s_data_i[6]  & \new_[3616]_ ;
  assign \wb0_addr_o[0]  = \wb1_addr_i[0]  & \new_[3616]_ ;
  assign \wb1m_data_o[28]  = \wb0s_data_i[28]  & \new_[3616]_ ;
  assign \wb1m_data_o[30]  = \wb0s_data_i[30]  & \new_[3616]_ ;
  assign \new_[3426]_  = ~\new_[3646]_  & ~\new_[3580]_ ;
  assign \new_[3427]_  = ~\new_[3643]_  & ~\new_[3581]_ ;
  assign \new_[3428]_  = \new_[3586]_  | \new_[3879]_ ;
  assign \new_[3429]_  = ~\new_[3527]_ ;
  assign \new_[3430]_  = ~\new_[2833]_  | ~\new_[3642]_  | ~\new_[3647]_ ;
  assign \new_[3431]_  = ~\new_[2928]_  | ~\new_[3642]_  | ~\new_[3647]_ ;
  assign \new_[3432]_  = ~\new_[4229]_  | ~\new_[3724]_  | ~\new_[3658]_ ;
  assign \new_[3433]_  = ~\new_[1247]_  | ~\new_[1246]_  | ~\new_[3608]_  | ~\new_[3870]_ ;
  assign \new_[3434]_  = ~\new_[1376]_  | ~\new_[1345]_  | ~\new_[3588]_  | ~\new_[3956]_ ;
  assign \wb1_addr_o[0]  = ~\new_[4128]_  & ~\new_[3592]_ ;
  assign \new_[3436]_  = \new_[3584]_  & \new_[3747]_ ;
  assign \new_[3437]_  = ~\new_[3613]_  & (~\new_[3848]_  | ~\new_[1700]_ );
  assign \new_[3438]_  = ~\wb1m_data_i[23]  | ~\new_[3616]_ ;
  assign \new_[3439]_  = ~\wb1m_data_i[15]  | ~\new_[3616]_ ;
  assign \new_[3440]_  = ~\wb1m_data_i[24]  | ~\new_[3616]_ ;
  assign \new_[3441]_  = ~\wb1m_data_i[30]  | ~\new_[3616]_ ;
  assign \new_[3442]_  = ~\wb1m_data_i[14]  | ~\new_[3616]_ ;
  assign \new_[3443]_  = ~\wb1m_data_i[16]  | ~\new_[3616]_ ;
  assign \new_[3444]_  = ~\wb1m_data_i[12]  | ~\new_[3616]_ ;
  assign \new_[3445]_  = ~\new_[3616]_  | ~\wb1m_data_i[31] ;
  assign \new_[3446]_  = ~\wb1m_data_i[29]  | ~\new_[3616]_ ;
  assign \new_[3447]_  = ~\wb1m_data_i[21]  | ~\new_[3616]_ ;
  assign \new_[3448]_  = ~\wb1m_data_i[22]  | ~\new_[3616]_ ;
  assign \new_[3449]_  = ~\wb1m_data_i[28]  | ~\new_[3616]_ ;
  assign \new_[3450]_  = ~\wb1m_data_i[25]  | ~\new_[3616]_ ;
  assign \new_[3451]_  = ~\new_[3203]_  & ~\new_[3591]_ ;
  assign \new_[3452]_  = ~\new_[3862]_  & ~\new_[3863]_ ;
  assign \new_[3453]_  = \new_[3202]_  | \new_[3614]_ ;
  assign \new_[3454]_  = ~\new_[4335]_ ;
  assign \new_[3455]_  = ~n3126 & ~\new_[3826]_ ;
  assign \new_[3456]_  = ~\new_[3596]_  | ~\new_[3609]_ ;
  assign \new_[3457]_  = \new_[3662]_  ? \new_[3887]_  : \new_[3655]_ ;
  assign \new_[3458]_  = (~\new_[3621]_  | ~\new_[3887]_ ) & (~\new_[3666]_  | ~\new_[3814]_ );
  assign \new_[3459]_  = (~\new_[3713]_  | ~\new_[3887]_ ) & (~\new_[3660]_  | ~\new_[3887]_ );
  assign \new_[3460]_  = \new_[3663]_  ? \new_[3887]_  : \new_[3668]_ ;
  assign \new_[3461]_  = ~\new_[3597]_  & (~\new_[3741]_  | ~\new_[3887]_ );
  assign \new_[3462]_  = \new_[3663]_  ? \new_[4046]_  : \new_[3668]_ ;
  assign \new_[3463]_  = ~\new_[4046]_  & (~\new_[3740]_  | ~\new_[3664]_ );
  assign \wb1_sel_o[3]  = \wb0_sel_i[3]  | \new_[3592]_ ;
  assign \new_[3465]_  = \new_[3599]_  & \new_[3862]_ ;
  assign \wb1_sel_o[1]  = \wb0_sel_i[1]  | \new_[3592]_ ;
  assign \new_[3467]_  = \new_[3599]_  & \new_[3890]_ ;
  assign \new_[3468]_  = \new_[3601]_  & \new_[3599]_ ;
  assign \wb1m_data_o[17]  = \wb0s_data_i[17]  & \new_[3616]_ ;
  assign \new_[3470]_  = \new_[3725]_  & \new_[3822]_ ;
  assign \new_[3471]_  = u2_mast0_drdy_r_reg;
  assign \new_[3472]_  = ~\new_[2832]_  & ~\new_[4077]_ ;
  assign \new_[3473]_  = \new_[3591]_  | \new_[2649]_ ;
  assign \wb1m_data_o[9]  = \wb0s_data_i[9]  & \new_[3616]_ ;
  assign \new_[3475]_  = \new_[3599]_  & \new_[3826]_ ;
  assign \new_[3476]_  = ~\wb1m_data_i[27]  | ~\new_[3616]_ ;
  assign \wb1m_data_o[15]  = \wb0s_data_i[15]  & \new_[3616]_ ;
  assign \new_[3478]_  = u3_u1_rf_ack_reg;
  assign \wb0_addr_o[1]  = \wb1_addr_i[1]  & \new_[3616]_ ;
  assign \wb1m_data_o[20]  = \wb0s_data_i[20]  & \new_[3616]_ ;
  assign \wb1m_data_o[11]  = \wb0s_data_i[11]  & \new_[3616]_ ;
  assign \wb1m_data_o[1]  = \wb0s_data_i[1]  & \new_[3616]_ ;
  assign wb1_err_o = wb0_err_i & \new_[3616]_ ;
  assign \new_[3484]_  = ~\new_[3848]_  & (~\new_[3711]_  | ~\new_[3709]_ );
  assign \wb1m_data_o[24]  = \wb0s_data_i[24]  & \new_[3616]_ ;
  assign \wb1m_data_o[22]  = \wb0s_data_i[22]  & \new_[3616]_ ;
  assign \wb1m_data_o[16]  = \wb0s_data_i[16]  & \new_[3616]_ ;
  assign \wb1m_data_o[10]  = \wb0s_data_i[10]  & \new_[3616]_ ;
  assign \wb1m_data_o[2]  = \wb0s_data_i[2]  & \new_[3616]_ ;
  assign \wb1m_data_o[25]  = \wb0s_data_i[25]  & \new_[3616]_ ;
  assign \wb1_sel_o[0]  = \wb0_sel_i[0]  | \new_[3592]_ ;
  assign \wb1m_data_o[23]  = \wb0s_data_i[23]  & \new_[3616]_ ;
  assign \wb1m_data_o[21]  = \wb0s_data_i[21]  & \new_[3616]_ ;
  assign \wb1m_data_o[29]  = \wb0s_data_i[29]  & \new_[3616]_ ;
  assign \wb1m_data_o[27]  = \wb0s_data_i[27]  & \new_[3616]_ ;
  assign \wb1m_data_o[31]  = \wb0s_data_i[31]  & \new_[3616]_ ;
  assign \new_[3497]_  = ~\new_[3520]_ ;
  assign \wb1_sel_o[2]  = \wb0_sel_i[2]  | \new_[3592]_ ;
  assign \wb1m_data_o[7]  = \wb0s_data_i[7]  & \new_[3616]_ ;
  assign \wb1_addr_o[1]  = ~\new_[4018]_  & ~\new_[3592]_ ;
  assign \wb1m_data_o[0]  = \wb0s_data_i[0]  & \new_[3616]_ ;
  assign \new_[3502]_  = ~\wb1m_data_i[26]  | ~\new_[3616]_ ;
  assign \new_[3503]_  = ~\wb1m_data_i[13]  | ~\new_[3616]_ ;
  assign \new_[3504]_  = \new_[3617]_  & \new_[3885]_ ;
  assign \new_[3505]_  = ~\wb1m_data_i[17]  | ~\new_[3616]_ ;
  assign \wb1m_data_o[3]  = \wb0s_data_i[3]  & \new_[3616]_ ;
  assign wb0_rty_o = ~\new_[4067]_  & ~\new_[3592]_ ;
  assign \new_[3508]_  = ~\new_[3953]_  | ~\new_[3598]_  | ~\new_[3947]_ ;
  assign wb0_err_o = ~\new_[4078]_  & ~\new_[3592]_ ;
  assign \new_[3510]_  = ~\new_[3619]_  & (~\new_[3747]_  | ~\new_[2032]_ );
  assign \new_[3511]_  = ~\wb1m_data_i[19]  | ~\new_[3616]_ ;
  assign \new_[3512]_  = ~\wb1m_data_i[18]  | ~\new_[3616]_ ;
  assign \new_[3513]_  = \new_[3585]_  & \new_[1240]_ ;
  assign \wb1m_data_o[19]  = \wb0s_data_i[19]  & \new_[3616]_ ;
  assign \new_[3515]_  = \new_[3617]_  & \new_[1384]_ ;
  assign \new_[3516]_  = \new_[1694]_  ^ \new_[3709]_ ;
  assign \new_[3517]_  = \new_[3585]_  & \new_[3914]_ ;
  assign \new_[3518]_  = \\u4_u0_mast_dout_reg[23] ;
  assign \new_[3519]_  = \\u4_u0_mast_dout_reg[20] ;
  assign \new_[3520]_  = ~\new_[3789]_  & ~\new_[3709]_ ;
  assign \new_[3521]_  = \\u4_u0_mast_dout_reg[16] ;
  assign \new_[3522]_  = \\u4_u0_mast_dout_reg[22] ;
  assign \new_[3523]_  = \\u4_u0_mast_dout_reg[5] ;
  assign \new_[3524]_  = \\u4_u0_mast_dout_reg[11] ;
  assign \new_[3525]_  = \\u4_u0_mast_dout_reg[12] ;
  assign \new_[3526]_  = ~\new_[3710]_  & ~\new_[3894]_ ;
  assign \new_[3527]_  = \new_[3638]_  | \new_[2068]_ ;
  assign \new_[3528]_  = \\u4_u0_mast_dout_reg[7] ;
  assign \new_[3529]_  = \\u4_u0_mast_dout_reg[3] ;
  assign n3106 = \new_[1385]_  ^ \new_[3726]_ ;
  assign n3111 = \new_[1242]_  ^ \new_[3748]_ ;
  assign n3121 = \new_[1383]_  ^ \new_[3756]_ ;
  assign n3116 = \new_[1239]_  ^ \new_[3754]_ ;
  assign \new_[3534]_  = \new_[3826]_  & \new_[4077]_ ;
  assign \new_[3535]_  = ~\new_[4340]_  & ~\new_[4010]_ ;
  assign \new_[3536]_  = \new_[4065]_  | \new_[3826]_ ;
  assign \new_[3537]_  = \new_[3707]_  | \new_[2609]_ ;
  assign \new_[3538]_  = ~\new_[4340]_  & ~\new_[3761]_ ;
  assign \new_[3539]_  = ~\new_[3892]_  | ~\new_[3650]_  | ~\new_[3869]_ ;
  assign \new_[3540]_  = ~\new_[3665]_  & (~\new_[3887]_  | ~\new_[4046]_ );
  assign \new_[3541]_  = ~\new_[3667]_  & (~\new_[3887]_  | ~\new_[4046]_ );
  assign \new_[3542]_  = ~\new_[3614]_ ;
  assign \new_[3543]_  = ~\new_[4215]_ ;
  assign \new_[3544]_  = ~\new_[3664]_  & ~\new_[3887]_ ;
  assign \new_[3545]_  = ~\new_[3761]_  & ~\new_[3669]_ ;
  assign \new_[3546]_  = \new_[4229]_  & \new_[4242]_ ;
  assign \new_[3547]_  = \\u4_u0_mast_dout_reg[13] ;
  assign \new_[3548]_  = ~n3126 & ~\new_[3868]_ ;
  assign \new_[3549]_  = ~\new_[3907]_  & ~\new_[3868]_ ;
  assign \new_[3550]_  = ~n3126 & ~\new_[4209]_ ;
  assign \new_[3551]_  = ~\new_[4227]_ ;
  assign \new_[3552]_  = \\u4_u0_mast_dout_reg[4] ;
  assign \new_[3553]_  = \\u4_u0_mast_dout_reg[27] ;
  assign \new_[3554]_  = \\u4_u0_mast_dout_reg[1] ;
  assign \new_[3555]_  = \\u4_u0_mast_dout_reg[26] ;
  assign \new_[3556]_  = \new_[3709]_  | \new_[3774]_ ;
  assign \new_[3557]_  = \\u4_u0_mast_dout_reg[25] ;
  assign \new_[3558]_  = \\u4_u0_mast_dout_reg[21] ;
  assign \new_[3559]_  = \\u4_u0_mast_dout_reg[2] ;
  assign \new_[3560]_  = \\u4_u0_mast_dout_reg[24] ;
  assign \new_[3561]_  = \\u4_u0_mast_dout_reg[0] ;
  assign \new_[3562]_  = \\u4_u0_mast_dout_reg[17] ;
  assign \new_[3563]_  = \\u4_u0_mast_dout_reg[31] ;
  assign \new_[3564]_  = \\u4_u0_mast_dout_reg[14] ;
  assign \new_[3565]_  = \\u4_u0_mast_dout_reg[8] ;
  assign \new_[3566]_  = \\u4_u0_mast_dout_reg[28] ;
  assign \new_[3567]_  = \\u4_u0_mast_dout_reg[10] ;
  assign \new_[3568]_  = \\u4_u0_mast_dout_reg[18] ;
  assign \new_[3569]_  = \\u4_u0_mast_dout_reg[29] ;
  assign \new_[3570]_  = \\u4_u0_mast_dout_reg[6] ;
  assign \new_[3571]_  = \\u4_u0_mast_dout_reg[9] ;
  assign \new_[3572]_  = \\u4_u0_mast_dout_reg[19] ;
  assign \new_[3573]_  = ~\new_[3746]_  & ~\new_[3622]_ ;
  assign \new_[3574]_  = ~\new_[3595]_ ;
  assign \new_[3575]_  = \\u4_u0_mast_dout_reg[15] ;
  assign \new_[3576]_  = \\u4_u0_mast_dout_reg[30] ;
  assign \new_[3577]_  = ~\new_[3598]_ ;
  assign \new_[3578]_  = ~n3126 & ~\new_[3883]_ ;
  assign \new_[3579]_  = ~\new_[3902]_  | ~\new_[3944]_  | ~\new_[3917]_ ;
  assign \new_[3580]_  = ~\new_[1383]_  | ~\new_[4082]_  | ~\new_[3756]_  | ~\new_[3885]_ ;
  assign \new_[3581]_  = ~\new_[1239]_  | ~\new_[4154]_  | ~\new_[3754]_  | ~\new_[3914]_ ;
  assign \new_[3582]_  = ~\new_[3794]_  | (~\new_[3763]_  & ~\new_[3880]_ );
  assign \new_[3583]_  = \\u2_u0_out_r_reg[1] ;
  assign \new_[3584]_  = ~\new_[3865]_  | ~\new_[2069]_ ;
  assign \new_[3585]_  = \new_[3754]_  & \new_[1239]_ ;
  assign \new_[3586]_  = ~\new_[3862]_  | ~\new_[3826]_ ;
  assign n3131 = ~\new_[3661]_ ;
  assign \new_[3588]_  = ~\new_[3726]_  & ~\new_[3798]_ ;
  assign \new_[3589]_  = ~\new_[3739]_  & (~\new_[3887]_  | ~\new_[4046]_ );
  assign \new_[3590]_  = \\u2_u1_out_r_reg[1] ;
  assign \new_[3591]_  = ~\new_[3732]_  | ~wb1_cyc_i;
  assign \new_[3592]_  = ~\new_[3649]_ ;
  assign \new_[3593]_  = ~\new_[3650]_ ;
  assign \new_[3594]_  = ~\new_[3707]_ ;
  assign \new_[3595]_  = ~\new_[3659]_ ;
  assign \new_[3596]_  = ~\new_[3887]_  | ~\new_[3806]_  | ~\new_[3805]_ ;
  assign \new_[3597]_  = \new_[3741]_  & \new_[4046]_ ;
  assign \new_[3598]_  = ~\new_[3753]_  & ~\new_[3820]_ ;
  assign \new_[3599]_  = ~\new_[3723]_  & ~\new_[3889]_ ;
  assign \new_[3600]_  = ~\new_[3713]_ ;
  assign \new_[3601]_  = ~\new_[3751]_  & ~\new_[4255]_ ;
  assign \new_[3602]_  = ~\new_[3660]_ ;
  assign \new_[3603]_  = ~\new_[3655]_ ;
  assign \new_[3604]_  = ~\new_[3621]_ ;
  assign \new_[3605]_  = \new_[3744]_  & \new_[4077]_ ;
  assign \new_[3606]_  = ~\new_[3649]_ ;
  assign \new_[3607]_  = ~\new_[3649]_ ;
  assign \new_[3608]_  = ~\new_[3748]_  & ~\new_[3765]_ ;
  assign \new_[3609]_  = \new_[3738]_  | \new_[4046]_ ;
  assign \new_[3610]_  = ~n3126 & ~\new_[4241]_ ;
  assign \new_[3611]_  = ~n3126 & ~\new_[3937]_ ;
  assign \new_[3612]_  = ~\new_[3807]_  | ~\new_[3826]_  | ~\new_[3808]_ ;
  assign \new_[3613]_  = ~\new_[3848]_  & (~\new_[3804]_  | ~\new_[3876]_ );
  assign \new_[3614]_  = ~\new_[3735]_  | ~wb0_cyc_i;
  assign \new_[3615]_  = ~n3126 & ~\new_[3879]_ ;
  assign \new_[3616]_  = ~\new_[3659]_ ;
  assign \new_[3617]_  = \new_[3756]_  & \new_[1383]_ ;
  assign \new_[3618]_  = \new_[3878]_  | \new_[1977]_  | \new_[3747]_  | \new_[2068]_ ;
  assign \new_[3619]_  = ~\new_[3747]_  & ~\new_[2032]_ ;
  assign \new_[3620]_  = ~\new_[3848]_  & (~\new_[3819]_  | ~\new_[3820]_ );
  assign \new_[3621]_  = \new_[3817]_  & \new_[3857]_ ;
  assign \new_[3622]_  = ~\new_[3894]_  & ~\new_[4242]_ ;
  assign n3291 = \new_[3576]_  ? wb1_ack_i : \wb1s_data_i[30] ;
  assign \new_[3624]_  = \\u1_ndr_r_reg[2] ;
  assign \new_[3625]_  = \\u1_ndr_r_reg[1] ;
  assign \new_[3626]_  = \\u1_ndr_r_reg[24] ;
  assign \new_[3627]_  = \\u1_ndr_r_reg[10] ;
  assign \new_[3628]_  = \\u1_ndr_r_reg[11] ;
  assign \new_[3629]_  = \\u1_ndr_r_reg[12] ;
  assign \new_[3630]_  = \\u1_ndr_r_reg[29] ;
  assign \new_[3631]_  = \\u1_ndr_r_reg[17] ;
  assign \new_[3632]_  = ~\\u1_ndr_r_reg[9] ;
  assign \new_[3633]_  = \\u1_ndr_r_reg[22] ;
  assign \new_[3634]_  = \\u1_ndr_r_reg[7] ;
  assign \new_[3635]_  = \\u1_ndr_r_reg[30] ;
  assign \new_[3636]_  = \\u1_ndr_r_reg[23] ;
  assign \new_[3637]_  = \\u1_ndr_r_reg[15] ;
  assign \new_[3638]_  = ~\new_[3787]_  | ~\new_[3902]_ ;
  assign \new_[3639]_  = \\u1_ndr_r_reg[14] ;
  assign \new_[3640]_  = \\u1_ndr_r_reg[28] ;
  assign \new_[3641]_  = \\u1_ndr_r_reg[18] ;
  assign \new_[3642]_  = ~\new_[4004]_  | ~\new_[3864]_  | ~\new_[3853]_ ;
  assign \new_[3643]_  = \new_[3777]_  | \new_[1243]_ ;
  assign \new_[3644]_  = \new_[3790]_  & \new_[1376]_ ;
  assign \new_[3645]_  = ~\new_[3777]_  & ~\new_[4114]_ ;
  assign \new_[3646]_  = ~\new_[3790]_  | ~\new_[4185]_ ;
  assign \new_[3647]_  = ~\new_[1895]_  | ~\new_[3864]_  | ~\new_[3853]_ ;
  assign \new_[3648]_  = ~\new_[3908]_  | (~\new_[3861]_  & ~\new_[3922]_ );
  assign \new_[3649]_  = \new_[3770]_  & wb0_cyc_i;
  assign \new_[3650]_  = \new_[3939]_  & \new_[3788]_ ;
  assign \new_[3651]_  = ~\new_[3824]_  | ~\new_[1378]_ ;
  assign \new_[3652]_  = ~\new_[3828]_  | ~\new_[1287]_ ;
  assign \new_[3653]_  = ~\new_[3788]_  | ~\new_[3953]_ ;
  assign \new_[3654]_  = ~\\u1_ndr_r_reg[16] ;
  assign \new_[3655]_  = \new_[3839]_  & \new_[3805]_ ;
  assign \new_[3656]_  = ~\new_[3793]_  | (~\new_[3880]_  & ~\new_[2034]_ );
  assign \new_[3657]_  = \new_[1693]_  ^ \new_[3848]_ ;
  assign \new_[3658]_  = \new_[3808]_  & \new_[4089]_ ;
  assign \new_[3659]_  = ~\new_[3835]_  | ~wb1_cyc_i;
  assign \new_[3660]_  = \new_[3814]_  & \new_[3858]_ ;
  assign \new_[3661]_  = ~wb0_cyc_i | ~\new_[4134]_  | ~\new_[3810]_  | ~wb0_stb_i;
  assign \new_[3662]_  = \new_[3856]_  & \new_[3806]_ ;
  assign \new_[3663]_  = \new_[3814]_  & \new_[3806]_ ;
  assign \new_[3664]_  = ~\new_[3806]_  | ~\new_[3857]_ ;
  assign \new_[3665]_  = ~\new_[3817]_  | ~\new_[3805]_ ;
  assign \new_[3666]_  = \new_[3817]_  & \new_[4046]_ ;
  assign \new_[3667]_  = ~\new_[3805]_  | ~\new_[3858]_ ;
  assign \new_[3668]_  = \new_[3856]_  & \new_[3817]_ ;
  assign \new_[3669]_  = ~\new_[3725]_ ;
  assign \new_[3670]_  = ~\new_[3826]_  & (~\new_[3937]_  | ~\new_[4209]_ );
  assign \new_[3671]_  = ~\new_[1414]_  | ~\new_[3935]_  | ~\new_[1380]_  | ~\new_[1375]_ ;
  assign \new_[3672]_  = ~\\u1_ndr_r_reg[8] ;
  assign n3181 = \new_[3547]_  ? \new_[3840]_  : \wb1s_data_i[13] ;
  assign n3246 = \new_[3565]_  ? \new_[3840]_  : \wb1s_data_i[8] ;
  assign n3186 = \new_[3552]_  ? \new_[3840]_  : \wb1s_data_i[4] ;
  assign n3261 = \new_[3568]_  ? \new_[3840]_  : \wb1s_data_i[18] ;
  assign n3161 = \new_[3524]_  ? \new_[3840]_  : \wb1s_data_i[11] ;
  assign \new_[3678]_  = \\u1_ndr_r_reg[4] ;
  assign n3151 = \new_[3522]_  ? \new_[3840]_  : \wb1s_data_i[22] ;
  assign n3281 = \new_[3572]_  ? wb1_ack_i : \wb1s_data_i[19] ;
  assign n3141 = \new_[3519]_  ? \new_[3840]_  : \wb1s_data_i[20] ;
  assign \new_[3682]_  = \\u1_ndr_r_reg[27] ;
  assign n3276 = \new_[3571]_  ? \new_[3840]_  : \wb1s_data_i[9] ;
  assign n3156 = \new_[3523]_  ? \new_[3840]_  : \wb1s_data_i[5] ;
  assign n3241 = \new_[3564]_  ? \new_[3840]_  : \wb1s_data_i[14] ;
  assign n3231 = \new_[3562]_  ? \new_[3840]_  : \wb1s_data_i[17] ;
  assign n3166 = \new_[3525]_  ? \new_[3840]_  : \wb1s_data_i[12] ;
  assign n3256 = \new_[3567]_  ? \new_[3840]_  : \wb1s_data_i[10] ;
  assign n3226 = \new_[3561]_  ? wb1_ack_i : \wb1s_data_i[0] ;
  assign \new_[3690]_  = ~\\u1_ndr_r_reg[20] ;
  assign n3146 = \new_[3521]_  ? \new_[3840]_  : \wb1s_data_i[16] ;
  assign n3196 = \new_[3554]_  ? \new_[3840]_  : \wb1s_data_i[1] ;
  assign n3286 = \new_[3575]_  ? \new_[3840]_  : \wb1s_data_i[15] ;
  assign n3251 = \new_[3566]_  ? \new_[3840]_  : \wb1s_data_i[28] ;
  assign n3266 = \new_[3569]_  ? \new_[3840]_  : \wb1s_data_i[29] ;
  assign n3271 = \new_[3570]_  ? \new_[3840]_  : \wb1s_data_i[6] ;
  assign n3206 = \new_[3557]_  ? \new_[3840]_  : \wb1s_data_i[25] ;
  assign n3236 = \new_[3563]_  ? \new_[3840]_  : \wb1s_data_i[31] ;
  assign n3176 = \new_[3529]_  ? wb1_ack_i : \wb1s_data_i[3] ;
  assign n3221 = \new_[3560]_  ? \new_[3840]_  : \wb1s_data_i[24] ;
  assign n3171 = \new_[3528]_  ? \new_[3840]_  : \wb1s_data_i[7] ;
  assign n3136 = \new_[3518]_  ? \new_[3840]_  : \wb1s_data_i[23] ;
  assign n3201 = \new_[3555]_  ? \new_[3840]_  : \wb1s_data_i[26] ;
  assign \new_[3704]_  = ~\new_[4065]_  | ~\new_[3879]_ ;
  assign \new_[3705]_  = ~\new_[4209]_  & ~\new_[3907]_ ;
  assign \new_[3706]_  = ~\new_[3879]_  & ~\new_[3883]_ ;
  assign \new_[3707]_  = ~\new_[3779]_  | ~\new_[3966]_ ;
  assign n3216 = \new_[3559]_  ? \new_[3840]_  : \wb1s_data_i[2] ;
  assign \new_[3709]_  = \new_[3820]_  | \new_[1701]_ ;
  assign \new_[3710]_  = ~\new_[3826]_  | ~\new_[4242]_ ;
  assign \new_[3711]_  = ~\new_[3820]_  | ~\new_[1701]_ ;
  assign \new_[3712]_  = \\u1_ndr_r_reg[5] ;
  assign \new_[3713]_  = \new_[3839]_  & \new_[3814]_ ;
  assign \new_[3714]_  = \\u1_ndr_r_reg[6] ;
  assign \new_[3715]_  = \\u1_ndr_r_reg[19] ;
  assign \new_[3716]_  = \\u1_ndr_r_reg[21] ;
  assign \new_[3717]_  = \\u1_ndr_r_reg[25] ;
  assign \new_[3718]_  = \\u1_ndr_r_reg[13] ;
  assign \new_[3719]_  = ~\\u1_ndr_r_reg[3] ;
  assign n3211 = \new_[3558]_  ? \new_[3840]_  : \wb1s_data_i[21] ;
  assign n3191 = \new_[3553]_  ? \new_[3840]_  : \wb1s_data_i[27] ;
  assign \new_[3722]_  = \\u1_ndr_r_reg[26] ;
  assign \new_[3723]_  = ~\new_[3842]_  | ~\new_[4077]_ ;
  assign \new_[3724]_  = ~\new_[3879]_  & ~\new_[3863]_ ;
  assign \new_[3725]_  = \new_[3861]_  & \new_[3908]_ ;
  assign \new_[3726]_  = ~\new_[1383]_  | ~\new_[3973]_  | ~\new_[3885]_  | ~\new_[4069]_ ;
  assign \new_[3727]_  = \\u1_ndr_r_reg[0] ;
  assign \new_[3728]_  = \\u1_ndnr_reg[0] ;
  assign \new_[3729]_  = ~\new_[4230]_ ;
  assign \new_[3730]_  = ~\new_[3955]_  & ~\new_[3860]_ ;
  assign \new_[3731]_  = ~\new_[3828]_ ;
  assign \new_[3732]_  = ~\new_[3835]_ ;
  assign \new_[3733]_  = ~\new_[3824]_ ;
  assign \new_[3734]_  = ~\new_[3848]_  | ~\new_[1657]_ ;
  assign \new_[3735]_  = ~\new_[3770]_ ;
  assign \new_[3736]_  = ~\new_[3848]_  | ~\new_[1694]_ ;
  assign \new_[3737]_  = ~\new_[3841]_  & ~\new_[2649]_ ;
  assign \new_[3738]_  = ~\new_[3839]_  | ~\new_[3857]_ ;
  assign \new_[3739]_  = ~\new_[3839]_  | ~\new_[3856]_ ;
  assign \new_[3740]_  = ~\new_[3857]_  | ~\new_[3858]_ ;
  assign \new_[3741]_  = \new_[3856]_  & \new_[3858]_ ;
  assign \new_[3742]_  = \\u2_u0_out_r_reg[0] ;
  assign \new_[3743]_  = ~\new_[3822]_ ;
  assign \new_[3744]_  = ~\new_[3889]_  & ~\new_[3842]_ ;
  assign \new_[3745]_  = \new_[3889]_  & \new_[3842]_ ;
  assign \new_[3746]_  = ~\new_[3862]_  & ~\new_[3907]_ ;
  assign \new_[3747]_  = \new_[3865]_  | \new_[2069]_ ;
  assign \new_[3748]_  = ~\new_[1239]_  | ~\new_[3997]_  | ~\new_[3914]_  | ~\new_[4066]_ ;
  assign \new_[3749]_  = \\u2_u1_out_r_reg[0] ;
  assign \new_[3750]_  = \new_[3877]_  & \new_[3850]_ ;
  assign \new_[3751]_  = ~\new_[3854]_  | ~\new_[4089]_ ;
  assign \new_[3752]_  = \\u1_req_r_reg[0] ;
  assign \new_[3753]_  = \new_[3843]_  | \new_[1701]_ ;
  assign \new_[3754]_  = \new_[4066]_  & \new_[3997]_ ;
  assign n3301 = \new_[4066]_  ^ \new_[3997]_ ;
  assign \new_[3756]_  = \new_[4069]_  & \new_[3973]_ ;
  assign n3296 = \new_[4069]_  ^ \new_[3973]_ ;
  assign n3386 = \new_[4431]_  & \new_[4401]_ ;
  assign n3331 = \new_[4437]_  & \new_[4407]_ ;
  assign n3311 = \new_[4448]_  & \new_[4418]_ ;
  assign \new_[3761]_  = \new_[3888]_  | \new_[3933]_ ;
  assign n3406 = \new_[4422]_  & \new_[4392]_ ;
  assign \new_[3763]_  = ~\new_[3902]_  & (~\new_[2034]_  | ~\new_[2031]_ );
  assign n3346 = \new_[4440]_  & \new_[4410]_ ;
  assign \new_[3765]_  = ~\new_[1245]_  | ~\new_[3916]_  | ~\new_[1244]_ ;
  assign n3416 = \new_[4444]_  & \new_[4414]_ ;
  assign n3366 = \new_[4426]_  & \new_[4396]_ ;
  assign \new_[3768]_  = ~\new_[3880]_  | ~\new_[2069]_ ;
  assign n3446 = \new_[4446]_  & \new_[4416]_ ;
  assign \new_[3770]_  = \wb0_addr_i[31]  | \wb0_addr_i[28]  | \wb0_addr_i[29]  | \wb0_addr_i[30] ;
  assign \new_[3771]_  = ~\new_[3880]_  | ~\new_[2068]_ ;
  assign \new_[3772]_  = ~\new_[3880]_  | ~\new_[1977]_ ;
  assign \new_[3773]_  = ~\new_[3880]_  | ~\new_[1976]_ ;
  assign \new_[3774]_  = ~\new_[3947]_  | ~\new_[3918]_ ;
  assign \new_[3775]_  = ~\new_[3880]_  | ~\new_[1973]_ ;
  assign \new_[3776]_  = ~\new_[3877]_  | ~\new_[1231]_ ;
  assign \new_[3777]_  = ~\new_[3924]_  | ~\new_[1244]_ ;
  assign n3316 = \new_[4425]_  & \new_[4395]_ ;
  assign \new_[3779]_  = ~\new_[2604]_  | (~\new_[4117]_  & ~dma_ack_o);
  assign n3356 = \new_[4442]_  & \new_[4412]_ ;
  assign \new_[3781]_  = ~\new_[4209]_  & ~\new_[3868]_ ;
  assign n3351 = \new_[4427]_  & \new_[4397]_ ;
  assign n3341 = \new_[4432]_  & \new_[4402]_ ;
  assign \new_[3784]_  = \new_[3900]_  | \new_[1374]_ ;
  assign n3321 = \new_[4439]_  & \new_[4409]_ ;
  assign \new_[3786]_  = ~\new_[3982]_  | ~\new_[4122]_  | ~\new_[4156]_ ;
  assign \new_[3787]_  = ~\new_[2069]_  & ~\new_[3878]_ ;
  assign \new_[3788]_  = ~\new_[3951]_  & ~\new_[1700]_ ;
  assign \new_[3789]_  = ~\new_[3869]_  | ~\new_[4147]_ ;
  assign \new_[3790]_  = \new_[3891]_  & \new_[1388]_ ;
  assign \new_[3791]_  = ~\new_[3942]_  & ~\new_[3901]_ ;
  assign \new_[3792]_  = ~\new_[3948]_  | ~wb0_stb_i;
  assign \new_[3793]_  = ~\new_[3880]_  | ~\new_[2034]_ ;
  assign \new_[3794]_  = ~\new_[3880]_  | ~\new_[2031]_ ;
  assign n3436 = \new_[4424]_  & \new_[4394]_ ;
  assign \new_[3796]_  = ~\new_[3880]_  | ~\new_[2032]_ ;
  assign \new_[3797]_  = ~\new_[4011]_  | ~\new_[1373]_  | ~\new_[1370]_ ;
  assign \new_[3798]_  = ~\new_[1387]_  | ~\new_[3941]_  | ~\new_[1388]_ ;
  assign \new_[3799]_  = ~\new_[1232]_  | ~\new_[1231]_  | ~\new_[1236]_  | ~\new_[1233]_ ;
  assign n3381 = \new_[4421]_  & \new_[4391]_ ;
  assign n3371 = \new_[4434]_  & \new_[4404]_ ;
  assign n3431 = \new_[4428]_  & \new_[4398]_ ;
  assign \new_[3803]_  = ~\new_[3860]_ ;
  assign \new_[3804]_  = ~\new_[1693]_  | ~\new_[1700]_ ;
  assign \new_[3805]_  = ~\new_[2635]_  & ~\new_[2641]_ ;
  assign \new_[3806]_  = ~\new_[2648]_  & ~\new_[4053]_ ;
  assign \new_[3807]_  = ~\new_[3879]_  & ~\new_[3883]_ ;
  assign \new_[3808]_  = ~\new_[1555]_  & ~\new_[3911]_ ;
  assign n3391 = \new_[4433]_  & \new_[4403]_ ;
  assign \new_[3810]_  = \new_[3204]_  | \new_[3202]_ ;
  assign n3306 = \new_[4447]_  & \new_[4417]_ ;
  assign \new_[3812]_  = ~\new_[3935]_  | ~\new_[1381]_ ;
  assign n3326 = \new_[4438]_  & \new_[4408]_ ;
  assign \new_[3814]_  = \new_[2635]_  & \new_[2641]_ ;
  assign n3441 = \new_[4436]_  & \new_[4406]_ ;
  assign n3376 = \new_[4435]_  & \new_[4405]_ ;
  assign \new_[3817]_  = \new_[2648]_  & \new_[4053]_ ;
  assign n3411 = \new_[4429]_  & \new_[4399]_ ;
  assign \new_[3819]_  = ~\new_[3876]_  | ~\new_[1659]_ ;
  assign \new_[3820]_  = \new_[3876]_  | \new_[1659]_ ;
  assign n3421 = \new_[4443]_  & \new_[4413]_ ;
  assign \new_[3822]_  = ~\new_[3922]_ ;
  assign \new_[3823]_  = \new_[3871]_  & \new_[3922]_ ;
  assign \new_[3824]_  = \new_[3891]_  & \new_[3954]_ ;
  assign \new_[3825]_  = ~\new_[3900]_  & ~\new_[3893]_ ;
  assign \new_[3826]_  = ~\new_[3863]_ ;
  assign \new_[3827]_  = ~\new_[3994]_  | ~\new_[1284]_  | ~\new_[1228]_ ;
  assign \new_[3828]_  = \new_[3924]_  & \new_[3874]_ ;
  assign n3426 = \new_[4430]_  & \new_[4400]_ ;
  assign n3336 = \new_[4420]_  & \new_[4390]_ ;
  assign n3361 = \new_[4419]_  & \new_[4389]_ ;
  assign n3451 = \new_[4423]_  & \new_[4393]_ ;
  assign n3396 = \new_[4441]_  & \new_[4411]_ ;
  assign n3401 = \new_[4445]_  & \new_[4415]_ ;
  assign \new_[3835]_  = \wb1_addr_i[31]  | \wb1_addr_i[28]  | \wb1_addr_i[29]  | \wb1_addr_i[30] ;
  assign \new_[3836]_  = ~\new_[3893]_ ;
  assign \new_[3837]_  = ~\new_[3950]_ ;
  assign \new_[3838]_  = ~\new_[3883]_ ;
  assign \new_[3839]_  = ~\new_[4161]_  & ~\new_[4053]_ ;
  assign \new_[3840]_  = ~\new_[3866]_ ;
  assign \new_[3841]_  = ~wb1_stb_i | ~\new_[4091]_ ;
  assign \new_[3842]_  = ~\new_[3909]_ ;
  assign \new_[3843]_  = ~\new_[3918]_ ;
  assign \new_[3844]_  = ~\new_[3875]_ ;
  assign \new_[3845]_  = ~\new_[3930]_ ;
  assign \new_[3846]_  = ~\new_[3908]_ ;
  assign \new_[3847]_  = ~\new_[3933]_ ;
  assign \new_[3848]_  = ~\new_[2416]_  | ~\new_[4163]_ ;
  assign n3461 = ~\new_[4074]_  & ~dma_req_i;
  assign \new_[3850]_  = \new_[1229]_  & \new_[3959]_ ;
  assign \new_[3851]_  = ~\new_[3901]_ ;
  assign n3456 = ~\new_[4074]_  & ~\new_[4007]_ ;
  assign \new_[3853]_  = ~\new_[2610]_  | ~\new_[4072]_ ;
  assign \new_[3854]_  = ~\new_[3911]_ ;
  assign n3476 = ~\new_[4007]_  & ~dma_ack_o;
  assign \new_[3856]_  = \new_[4110]_  & \new_[2641]_ ;
  assign \new_[3857]_  = ~\new_[4110]_  & ~\new_[2641]_ ;
  assign \new_[3858]_  = \new_[4161]_  & \new_[4053]_ ;
  assign \new_[3859]_  = ~\new_[3919]_ ;
  assign \new_[3860]_  = ~\new_[3959]_  | ~\new_[1234]_ ;
  assign \new_[3861]_  = ~\new_[3871]_ ;
  assign \new_[3862]_  = ~\new_[3894]_ ;
  assign \new_[3863]_  = ~\new_[4216]_  | ~\new_[4241]_ ;
  assign \new_[3864]_  = ~\new_[2600]_  | ~\new_[4184]_ ;
  assign \new_[3865]_  = ~\new_[3902]_ ;
  assign \new_[3866]_  = ~wb1_ack_i;
  assign \new_[3867]_  = ~wb1_stb_i | ~wb1_we_i;
  assign \new_[3868]_  = ~\new_[4077]_ ;
  assign \new_[3869]_  = ~\new_[1695]_  & ~\new_[1696]_ ;
  assign \new_[3870]_  = \new_[1248]_  & \new_[1287]_ ;
  assign \new_[3871]_  = \\u3_u1_slv_adr_reg[3] ;
  assign \new_[3872]_  = ~wb0_err_i & ~wb1_err_i;
  assign n3126 = ~\new_[4065]_ ;
  assign \new_[3874]_  = \new_[1247]_  & \new_[1248]_ ;
  assign \new_[3875]_  = ~\\u3_u1_slv_dout_reg[4] ;
  assign \new_[3876]_  = \new_[1693]_  | \new_[1700]_ ;
  assign \new_[3877]_  = \new_[1237]_  & \new_[1285]_ ;
  assign \new_[3878]_  = \new_[2033]_  | \new_[2032]_ ;
  assign \new_[3879]_  = ~\new_[4234]_ ;
  assign \new_[3880]_  = \new_[3086]_  | \new_[1198]_ ;
  assign \new_[3881]_  = ~\new_[1231]_  | ~\new_[1237]_ ;
  assign \new_[3882]_  = ~\\u3_u1_slv_dout_reg[0] ;
  assign \new_[3883]_  = ~\new_[4089]_ ;
  assign \new_[3884]_  = \\u3_u1_slv_dout_reg[18] ;
  assign \new_[3885]_  = \new_[1384]_  & \new_[1389]_ ;
  assign \new_[3886]_  = ~\\u3_u1_slv_dout_reg[7] ;
  assign \new_[3887]_  = ~\new_[4046]_ ;
  assign \new_[3888]_  = \\u3_u1_slv_adr_reg[6] ;
  assign \new_[3889]_  = ~\new_[4133]_ ;
  assign \new_[3890]_  = ~\new_[3991]_ ;
  assign \new_[3891]_  = \new_[1387]_  & \new_[1345]_ ;
  assign \new_[3892]_  = ~\new_[1697]_  & ~\new_[1657]_ ;
  assign \new_[3893]_  = ~\new_[1372]_  | ~\new_[1371]_ ;
  assign \new_[3894]_  = ~\new_[4235]_ ;
  assign \new_[3895]_  = ~\\u3_u1_slv_dout_reg[5] ;
  assign \new_[3896]_  = \\u3_u1_slv_dout_reg[24] ;
  assign \new_[3897]_  = \\u3_u1_slv_dout_reg[1] ;
  assign \new_[3898]_  = \\u3_u1_slv_adr_reg[8] ;
  assign \new_[3899]_  = \\u3_u1_slv_dout_reg[19] ;
  assign \new_[3900]_  = ~\new_[1381]_  | ~\new_[1413]_ ;
  assign \new_[3901]_  = ~\new_[1371]_  | ~\new_[1382]_ ;
  assign \new_[3902]_  = ~\new_[2034]_  & ~\new_[2031]_ ;
  assign \new_[3903]_  = \\u3_u1_slv_dout_reg[31] ;
  assign \new_[3904]_  = ~\\u3_u1_slv_dout_reg[6] ;
  assign \new_[3905]_  = \\u3_u1_slv_adr_reg[9] ;
  assign \new_[3906]_  = \\u3_u1_slv_dout_reg[20] ;
  assign \new_[3907]_  = ~\new_[4242]_ ;
  assign \new_[3908]_  = ~\\u3_u1_slv_adr_reg[4] ;
  assign \new_[3909]_  = ~\new_[4071]_ ;
  assign \new_[3910]_  = \\u3_u1_slv_dout_reg[30] ;
  assign \new_[3911]_  = ~\new_[4233]_ ;
  assign \new_[3912]_  = \\u3_u1_slv_dout_reg[26] ;
  assign \new_[3913]_  = \\u3_u1_slv_dout_reg[29] ;
  assign \new_[3914]_  = \new_[1240]_  & \new_[1241]_ ;
  assign \new_[3915]_  = \\u3_u1_slv_dout_reg[28] ;
  assign \new_[3916]_  = ~\new_[1242]_  & ~\new_[1243]_ ;
  assign \new_[3917]_  = ~\new_[2068]_  & ~\new_[2033]_ ;
  assign \new_[3918]_  = ~\new_[1694]_  & ~\new_[1695]_ ;
  assign \new_[3919]_  = ~\\u3_u1_slv_dout_reg[2] ;
  assign \new_[3920]_  = ~\\u3_u1_slv_dout_reg[8] ;
  assign \new_[3921]_  = \\u3_u1_slv_adr_reg[7] ;
  assign \new_[3922]_  = ~\\u3_u1_slv_adr_reg[2] ;
  assign \new_[3923]_  = \\u3_u1_slv_dout_reg[14] ;
  assign \new_[3924]_  = \new_[1245]_  & \new_[1246]_ ;
  assign \new_[3925]_  = \\u3_u1_slv_dout_reg[23] ;
  assign \new_[3926]_  = ~\\u3_u1_slv_dout_reg[9] ;
  assign \new_[3927]_  = \\u3_u1_slv_dout_reg[21] ;
  assign \new_[3928]_  = \\u3_u1_slv_dout_reg[25] ;
  assign \new_[3929]_  = \\u3_u1_slv_dout_reg[27] ;
  assign \new_[3930]_  = ~\\u3_u1_slv_dout_reg[3] ;
  assign \new_[3931]_  = \\u3_u1_slv_dout_reg[12] ;
  assign \new_[3932]_  = \\u3_u1_slv_dout_reg[17] ;
  assign \new_[3933]_  = \\u3_u1_slv_adr_reg[5] ;
  assign \new_[3934]_  = ~\\u3_u1_slv_dout_reg[11] ;
  assign \new_[3935]_  = ~\new_[1374]_ ;
  assign \new_[3936]_  = \\u3_u1_slv_dout_reg[15] ;
  assign \new_[3937]_  = ~\new_[4216]_ ;
  assign \new_[3938]_  = \\u3_u1_slv_dout_reg[13] ;
  assign \new_[3939]_  = ~\new_[1693]_  & ~\new_[1694]_ ;
  assign \new_[3940]_  = ~\new_[1976]_  & ~\new_[1973]_ ;
  assign \new_[3941]_  = ~\new_[1385]_  & ~\new_[1386]_ ;
  assign \new_[3942]_  = ~\new_[1413]_  | ~\new_[1372]_ ;
  assign \new_[3943]_  = ~\\u3_u1_slv_dout_reg[10] ;
  assign \new_[3944]_  = ~\new_[2069]_  & ~\new_[2032]_ ;
  assign \new_[3945]_  = ~\new_[1977]_  & ~\new_[1976]_ ;
  assign \new_[3946]_  = \\u3_u1_slv_dout_reg[16] ;
  assign \new_[3947]_  = ~\new_[1696]_  & ~\new_[1697]_ ;
  assign \new_[3948]_  = ~wb0_we_i & ~\new_[3478]_ ;
  assign \new_[3949]_  = ~\new_[1702]_  & ~\new_[1698]_ ;
  assign \new_[3950]_  = ~\new_[2611]_  & ~\new_[2603]_ ;
  assign \new_[3951]_  = \new_[1659]_  | \new_[1701]_ ;
  assign \new_[3952]_  = \\u3_u1_slv_dout_reg[22] ;
  assign \new_[3953]_  = ~\new_[1657]_  & ~\new_[1702]_ ;
  assign \new_[3954]_  = \new_[1376]_  & \new_[1377]_ ;
  assign \new_[3955]_  = ~\new_[1285]_  | ~\new_[1229]_ ;
  assign \new_[3956]_  = \new_[1377]_  & \new_[1378]_ ;
  assign \new_[3957]_  = ~\new_[2882]_ ;
  assign \new_[3958]_  = ~\new_[3235]_ ;
  assign \new_[3959]_  = ~\new_[1230]_ ;
  assign \new_[3960]_  = ~\new_[3253]_ ;
  assign \new_[3961]_  = ~\new_[1889]_ ;
  assign \new_[3962]_  = ~\new_[3266]_ ;
  assign \new_[3963]_  = ~\new_[2831]_ ;
  assign \new_[3964]_  = ~\new_[2907]_ ;
  assign \new_[3965]_  = ~\new_[3228]_ ;
  assign \new_[3966]_  = ~\new_[1390]_ ;
  assign \new_[3967]_  = ~\new_[1887]_ ;
  assign \new_[3968]_  = ~\new_[2910]_ ;
  assign \new_[3969]_  = ~\new_[3255]_ ;
  assign \new_[3970]_  = ~\new_[3225]_ ;
  assign \new_[3971]_  = ~\new_[3272]_ ;
  assign \new_[3972]_  = ~\new_[3012]_ ;
  assign \new_[3973]_  = ~n3466;
  assign \new_[3974]_  = ~\new_[3047]_ ;
  assign \new_[3975]_  = ~\new_[1965]_ ;
  assign \new_[3976]_  = ~\new_[1880]_ ;
  assign \new_[3977]_  = ~\new_[3269]_ ;
  assign \new_[3978]_  = ~\new_[1784]_ ;
  assign \new_[3979]_  = ~\new_[3270]_ ;
  assign \new_[3980]_  = ~\new_[2921]_ ;
  assign \new_[3981]_  = ~\new_[1787]_ ;
  assign \new_[3982]_  = ~\new_[1699]_ ;
  assign \new_[3983]_  = ~\new_[3250]_ ;
  assign \new_[3984]_  = ~\new_[1893]_ ;
  assign \new_[3985]_  = ~\new_[3026]_ ;
  assign \new_[3986]_  = ~\new_[2948]_ ;
  assign \new_[3987]_  = ~\new_[1235]_ ;
  assign \new_[3988]_  = ~\new_[1782]_ ;
  assign \new_[3989]_  = ~\new_[1243]_ ;
  assign \new_[3990]_  = ~\new_[1783]_ ;
  assign \new_[3991]_  = ~\new_[1555]_ ;
  assign \new_[3992]_  = ~\new_[1415]_ ;
  assign \new_[3993]_  = ~\new_[3028]_ ;
  assign \new_[3994]_  = ~\new_[1227]_ ;
  assign \new_[3995]_  = ~\new_[1788]_ ;
  assign \new_[3996]_  = ~\new_[1801]_ ;
  assign \new_[3997]_  = ~n3471;
  assign \new_[3998]_  = ~\new_[1800]_ ;
  assign \new_[3999]_  = ~\new_[2633]_ ;
  assign \new_[4000]_  = ~\new_[2652]_ ;
  assign \new_[4001]_  = ~\new_[1884]_ ;
  assign \new_[4002]_  = ~\new_[3007]_ ;
  assign \new_[4003]_  = ~\new_[3294]_ ;
  assign \new_[4004]_  = ~\new_[2601]_ ;
  assign \new_[4005]_  = ~\new_[1776]_ ;
  assign \new_[4006]_  = ~\new_[3030]_ ;
  assign \new_[4007]_  = ~dma_req_i;
  assign \new_[4008]_  = ~\new_[2898]_ ;
  assign \new_[4009]_  = ~\new_[3259]_ ;
  assign \new_[4010]_  = ~\new_[3204]_ ;
  assign \new_[4011]_  = ~\new_[1369]_ ;
  assign \new_[4012]_  = ~\new_[1803]_ ;
  assign \new_[4013]_  = ~\new_[2603]_ ;
  assign \new_[4014]_  = ~\new_[1753]_ ;
  assign \new_[4015]_  = ~\new_[2644]_ ;
  assign \new_[4016]_  = ~\new_[2602]_ ;
  assign \new_[4017]_  = ~\new_[2650]_ ;
  assign \new_[4018]_  = ~\wb0_addr_i[1] ;
  assign \new_[4019]_  = ~\new_[3009]_ ;
  assign \new_[4020]_  = ~\new_[1968]_ ;
  assign \new_[4021]_  = ~\new_[1796]_ ;
  assign \new_[4022]_  = ~wb0_rty_i;
  assign \new_[4023]_  = ~\new_[3226]_ ;
  assign \new_[4024]_  = ~\new_[3275]_ ;
  assign \new_[4025]_  = ~\new_[3245]_ ;
  assign \new_[4026]_  = ~\new_[1759]_ ;
  assign \new_[4027]_  = ~\new_[3233]_ ;
  assign \new_[4028]_  = ~\new_[3262]_ ;
  assign \new_[4029]_  = ~\new_[3287]_ ;
  assign \new_[4030]_  = ~\new_[1762]_ ;
  assign \new_[4031]_  = ~\new_[2909]_ ;
  assign \new_[4032]_  = ~\new_[1890]_ ;
  assign \new_[4033]_  = ~\new_[2924]_ ;
  assign \new_[4034]_  = ~\new_[1766]_ ;
  assign \new_[4035]_  = ~\new_[2903]_ ;
  assign \new_[4036]_  = ~\new_[2926]_ ;
  assign \new_[4037]_  = ~\new_[1734]_ ;
  assign \new_[4038]_  = ~\new_[2894]_ ;
  assign \new_[4039]_  = ~\new_[2927]_ ;
  assign \new_[4040]_  = ~\new_[2863]_ ;
  assign \new_[4041]_  = ~\new_[2851]_ ;
  assign \new_[4042]_  = ~\new_[2842]_ ;
  assign \new_[4043]_  = ~\new_[1892]_ ;
  assign \new_[4045]_  = ~\new_[1891]_ ;
  assign \new_[4046]_  = ~\new_[2645]_ ;
  assign \new_[4047]_  = ~\new_[1728]_ ;
  assign \new_[4048]_  = ~\wb0s_data_i[14] ;
  assign \new_[4049]_  = ~\new_[2920]_ ;
  assign \new_[4050]_  = ~\new_[1883]_ ;
  assign \new_[4051]_  = ~\new_[2901]_ ;
  assign \new_[4052]_  = ~\new_[1756]_ ;
  assign \new_[4053]_  = \new_[2634]_ ;
  assign \new_[4054]_  = ~\new_[3267]_ ;
  assign \new_[4055]_  = ~\new_[1895]_ ;
  assign \new_[4056]_  = ~\new_[1736]_ ;
  assign \new_[4057]_  = ~\new_[1733]_ ;
  assign \new_[4058]_  = ~\new_[1772]_ ;
  assign \new_[4059]_  = ~\new_[1770]_ ;
  assign \new_[4060]_  = ~\new_[1769]_ ;
  assign \new_[4061]_  = ~\new_[1731]_ ;
  assign \new_[4062]_  = ~\new_[2636]_ ;
  assign \new_[4063]_  = ~\new_[1761]_ ;
  assign \new_[4064]_  = ~\new_[1758]_ ;
  assign \new_[4065]_  = ~wb0_ack_i;
  assign \new_[4066]_  = ~\new_[1288]_ ;
  assign \new_[4067]_  = ~wb1_rty_i;
  assign \new_[4068]_  = ~\new_[1238]_ ;
  assign \new_[4069]_  = ~\new_[1592]_ ;
  assign \new_[4070]_  = ~\new_[1416]_ ;
  assign \new_[4071]_  = ~\new_[1196]_ ;
  assign \new_[4072]_  = ~\new_[1498]_ ;
  assign \new_[4073]_  = ~\new_[1871]_ ;
  assign \new_[4074]_  = ~dma_nd_i;
  assign \new_[4075]_  = ~\new_[1775]_ ;
  assign \new_[4076]_  = ~\new_[2606]_ ;
  assign \new_[4077]_  = ~\new_[1499]_ ;
  assign \new_[4078]_  = ~wb1_err_i;
  assign \new_[4079]_  = ~\new_[3274]_ ;
  assign \new_[4080]_  = ~\new_[1251]_ ;
  assign \new_[4081]_  = ~\new_[2651]_ ;
  assign \new_[4082]_  = ~\new_[1385]_ ;
  assign \new_[4083]_  = ~\new_[1888]_ ;
  assign \new_[4084]_  = ~\new_[3042]_ ;
  assign \new_[4085]_  = ~\new_[2643]_ ;
  assign \new_[4086]_  = ~\new_[3203]_ ;
  assign \new_[4087]_  = ~\new_[1885]_ ;
  assign \new_[4088]_  = ~\new_[1798]_ ;
  assign \new_[4089]_  = ~\new_[2698]_ ;
  assign \new_[4090]_  = ~\new_[1780]_ ;
  assign \new_[4091]_  = ~wb1_we_i;
  assign \new_[4092]_  = ~\new_[1786]_ ;
  assign \new_[4093]_  = ~\new_[1879]_ ;
  assign \new_[4094]_  = ~\new_[2854]_ ;
  assign \new_[4095]_  = ~\new_[2861]_ ;
  assign \new_[4096]_  = ~\new_[1774]_ ;
  assign \new_[4097]_  = ~\new_[3041]_ ;
  assign \new_[4098]_  = ~\new_[1777]_ ;
  assign \new_[4099]_  = ~\new_[2930]_ ;
  assign \new_[4100]_  = ~\new_[1894]_ ;
  assign \new_[4101]_  = ~\new_[1789]_ ;
  assign \new_[4102]_  = ~\new_[3032]_ ;
  assign \new_[4103]_  = ~\new_[3268]_ ;
  assign \new_[4104]_  = ~\new_[1802]_ ;
  assign \new_[4105]_  = ~\new_[2932]_ ;
  assign \new_[4106]_  = ~\new_[3039]_ ;
  assign \new_[4107]_  = ~\new_[3004]_ ;
  assign \new_[4108]_  = ~\new_[2638]_ ;
  assign \new_[4109]_  = ~\new_[3038]_ ;
  assign \new_[4110]_  = ~\new_[2635]_ ;
  assign \new_[4111]_  = ~\new_[3248]_ ;
  assign \new_[4112]_  = ~\new_[1804]_ ;
  assign \new_[4113]_  = ~\new_[3051]_ ;
  assign \new_[4114]_  = ~\new_[1247]_ ;
  assign \new_[4115]_  = ~\new_[3008]_ ;
  assign \new_[4116]_  = ~\new_[3027]_ ;
  assign \new_[4117]_  = ~\new_[3752]_ ;
  assign \new_[4118]_  = ~\new_[3033]_ ;
  assign \new_[4119]_  = ~\new_[1781]_ ;
  assign \new_[4120]_  = ~\new_[1779]_ ;
  assign \new_[4121]_  = ~\new_[1962]_ ;
  assign \new_[4122]_  = ~\new_[1693]_ ;
  assign \new_[4123]_  = ~\new_[3036]_ ;
  assign \new_[4124]_  = ~\new_[3273]_ ;
  assign \new_[4125]_  = ~\wb0s_data_i[4] ;
  assign \new_[4126]_  = ~\new_[2905]_ ;
  assign \new_[4127]_  = ~\new_[2608]_ ;
  assign \new_[4128]_  = ~\wb0_addr_i[0] ;
  assign \new_[4129]_  = ~\new_[1737]_ ;
  assign \new_[4130]_  = ~\new_[1878]_ ;
  assign \new_[4131]_  = ~\new_[3282]_ ;
  assign \new_[4132]_  = ~\new_[3005]_ ;
  assign \new_[4133]_  = ~\new_[1727]_ ;
  assign \new_[4134]_  = ~\new_[3478]_ ;
  assign \new_[4135]_  = ~\new_[3263]_ ;
  assign \new_[4136]_  = ~\new_[3276]_ ;
  assign \new_[4137]_  = ~\new_[3279]_ ;
  assign \new_[4138]_  = ~\new_[1760]_ ;
  assign \new_[4139]_  = ~\new_[1339]_ ;
  assign \new_[4140]_  = ~\new_[2929]_ ;
  assign \new_[4141]_  = ~\new_[3006]_ ;
  assign \new_[4142]_  = ~\new_[1763]_ ;
  assign \new_[4143]_  = ~\new_[2841]_ ;
  assign \new_[4144]_  = ~\new_[2906]_ ;
  assign \new_[4145]_  = ~\new_[1765]_ ;
  assign \new_[4146]_  = ~\new_[2904]_ ;
  assign \new_[4147]_  = ~\new_[1694]_ ;
  assign \new_[4148]_  = ~\new_[1768]_ ;
  assign \new_[4149]_  = ~\new_[2897]_ ;
  assign \new_[4150]_  = ~\new_[2895]_ ;
  assign \new_[4151]_  = ~\new_[2878]_ ;
  assign \new_[4152]_  = ~\new_[2860]_ ;
  assign \new_[4153]_  = ~\new_[1967]_ ;
  assign \new_[4154]_  = ~\new_[1242]_ ;
  assign \new_[4155]_  = ~\new_[2902]_ ;
  assign \new_[4156]_  = ~\new_[1698]_ ;
  assign \new_[4157]_  = ~\new_[3295]_ ;
  assign \new_[4158]_  = ~\new_[1342]_ ;
  assign \new_[4159]_  = ~\new_[1732]_ ;
  assign \new_[4160]_  = ~\new_[1735]_ ;
  assign \new_[4161]_  = ~\new_[2648]_ ;
  assign \new_[4162]_  = ~\new_[1882]_ ;
  assign \new_[4163]_  = ~\new_[1199]_ ;
  assign \new_[4164]_  = ~\new_[1778]_ ;
  assign \new_[4165]_  = ~\new_[1754]_ ;
  assign \new_[4166]_  = ~\new_[2908]_ ;
  assign \new_[4167]_  = ~\new_[2945]_ ;
  assign \new_[4168]_  = ~\new_[3010]_ ;
  assign \new_[4169]_  = ~\new_[1755]_ ;
  assign \new_[4170]_  = ~\new_[3227]_ ;
  assign \new_[4171]_  = ~\new_[3264]_ ;
  assign \new_[4172]_  = ~\new_[3052]_ ;
  assign \new_[4173]_  = ~\new_[1417]_ ;
  assign \new_[4174]_  = ~\new_[3011]_ ;
  assign \new_[4175]_  = ~\new_[1853]_ ;
  assign \new_[4176]_  = ~\new_[1773]_ ;
  assign \new_[4177]_  = ~\new_[1771]_ ;
  assign \new_[4178]_  = ~\new_[2925]_ ;
  assign \new_[4179]_  = ~\new_[1767]_ ;
  assign \new_[4180]_  = ~\new_[1960]_ ;
  assign \new_[4181]_  = ~\new_[2911]_ ;
  assign \new_[4182]_  = ~\new_[1764]_ ;
  assign \new_[4183]_  = ~\new_[2899]_ ;
  assign \new_[4184]_  = ~\new_[1340]_ ;
  assign \new_[4185]_  = ~\new_[1386]_ ;
  assign \new_[4186]_  = ~\new_[4193]_ ;
  assign \new_[4187]_  = \new_[4193]_ ;
  assign \new_[4188]_  = \new_[4191]_ ;
  assign \new_[4189]_  = ~\new_[4191]_ ;
  assign \new_[4190]_  = ~\new_[4191]_ ;
  assign \new_[4191]_  = ~\new_[4193]_ ;
  assign \new_[4192]_  = ~\new_[4191]_ ;
  assign \new_[4193]_  = ~\new_[4373]_ ;
  assign \new_[4194]_  = ~\new_[4356]_ ;
  assign \new_[4195]_  = ~\new_[4196]_ ;
  assign \new_[4196]_  = ~\new_[4357]_ ;
  assign \new_[4197]_  = \new_[4372]_ ;
  assign \new_[4198]_  = \new_[4373]_ ;
  assign \new_[4199]_  = ~\new_[4212]_ ;
  assign \new_[4200]_  = ~\new_[4201]_ ;
  assign \new_[4201]_  = \new_[1520]_ ;
  assign \new_[4202]_  = \new_[1520]_ ;
  assign \new_[4203]_  = \new_[1520]_ ;
  assign \new_[4204]_  = \new_[1520]_ ;
  assign n2291 = ~\new_[4206]_ ;
  assign \new_[4206]_  = \new_[2629]_ ;
  assign \new_[4207]_  = ~\new_[4348]_ ;
  assign \new_[4208]_  = ~\new_[4326]_ ;
  assign \new_[4209]_  = ~\new_[4241]_ ;
  assign \new_[4210]_  = \new_[4211]_ ;
  assign \new_[4211]_  = ~\new_[2761]_ ;
  assign \new_[4212]_  = ~\new_[4334]_  | ~\new_[4241]_ ;
  assign \new_[4213]_  = ~\new_[2648]_  | ~\new_[4319]_  | ~\new_[3551]_  | ~\new_[4237]_ ;
  assign \new_[4214]_  = ~\new_[2641]_  | ~\new_[4237]_  | ~\new_[4319]_ ;
  assign \new_[4215]_  = ~\new_[4237]_ ;
  assign \new_[4216]_  = \new_[4236]_ ;
  assign \new_[4217]_  = ~\new_[4225]_  | ~\new_[4222]_  | ~\new_[4218]_  | ~\new_[4221]_ ;
  assign \new_[4218]_  = ~\new_[4219]_ ;
  assign \new_[4219]_  = ~\new_[2597]_  | ~\new_[2440]_  | ~\new_[4220]_  | ~\new_[2439]_ ;
  assign \new_[4220]_  = ~\new_[2670]_  | ~\new_[2582]_ ;
  assign \new_[4221]_  = ~\new_[2422]_  & ~\new_[2427]_ ;
  assign \new_[4222]_  = ~\new_[4223]_  & ~\new_[4224]_ ;
  assign \new_[4223]_  = ~\new_[2544]_  | ~\new_[2590]_ ;
  assign \new_[4224]_  = ~\new_[2525]_ ;
  assign \new_[4225]_  = ~\new_[2401]_  & ~\new_[2423]_ ;
  assign \new_[4226]_  = ~\new_[4227]_ ;
  assign \new_[4227]_  = \new_[1555]_  | \new_[4230]_ ;
  assign \new_[4228]_  = \new_[4226]_ ;
  assign \new_[4229]_  = \new_[4319]_ ;
  assign \new_[4230]_  = ~\new_[4233]_  | ~\new_[4231]_  | ~\new_[4232]_ ;
  assign \new_[4231]_  = ~\new_[2698]_ ;
  assign \new_[4232]_  = ~\new_[2699]_ ;
  assign \new_[4233]_  = ~\new_[1691]_ ;
  assign \new_[4234]_  = \new_[4232]_ ;
  assign \new_[4235]_  = ~\new_[1692]_ ;
  assign \new_[4236]_  = ~\new_[2700]_ ;
  assign \new_[4237]_  = ~\new_[4238]_  & ~\new_[4331]_ ;
  assign \new_[4238]_  = ~\new_[4236]_  | ~\new_[4235]_ ;
  assign \new_[4239]_  = ~\new_[2578]_ ;
  assign \new_[4240]_  = ~\new_[1197]_ ;
  assign \new_[4241]_  = \new_[4239]_ ;
  assign \new_[4242]_  = \new_[4240]_ ;
  assign \new_[4243]_  = ~\new_[4350]_  & ~\new_[4244]_ ;
  assign \new_[4244]_  = ~\new_[4354]_  | ~\new_[4245]_ ;
  assign \new_[4245]_  = ~\new_[4353]_ ;
  assign \new_[4246]_  = ~\new_[2627]_  | ~\new_[4247]_  | ~\new_[2598]_ ;
  assign \new_[4247]_  = ~\new_[4349]_  | ~\new_[2751]_ ;
  assign \new_[4248]_  = ~\new_[4250]_  | ~\new_[2654]_  | ~\new_[4249]_ ;
  assign \new_[4249]_  = ~\new_[2665]_ ;
  assign \new_[4250]_  = ~\new_[2668]_ ;
  assign \new_[4251]_  = ~\new_[4252]_  | ~\new_[4256]_ ;
  assign \new_[4252]_  = ~\new_[4253]_  | ~\new_[4254]_ ;
  assign \new_[4253]_  = ~\new_[4217]_  | ~\new_[2567]_  | ~\new_[2575]_ ;
  assign \new_[4254]_  = ~\new_[4255]_ ;
  assign \new_[4255]_  = \new_[3890]_  | \new_[3879]_ ;
  assign \new_[4256]_  = \new_[4257]_  | \new_[4260]_ ;
  assign \new_[4257]_  = ~\new_[4258]_  & (~\new_[4255]_  | ~wb0_ack_i);
  assign \new_[4258]_  = ~\new_[4259]_ ;
  assign \new_[4259]_  = ~\new_[4242]_  | ~\new_[4234]_ ;
  assign \new_[4260]_  = ~\new_[4254]_  & ~\new_[4261]_ ;
  assign \new_[4261]_  = ~\new_[4258]_  | ~\new_[4065]_ ;
  assign n1571 = ~\new_[4264]_  | (~\new_[4308]_  & ~\new_[4263]_ );
  assign \new_[4263]_  = ~\new_[3620]_  & (~\new_[3848]_  | ~\new_[1659]_ );
  assign \new_[4264]_  = \new_[1799]_  | \new_[4265]_ ;
  assign \new_[4265]_  = ~\new_[4302]_  | ~\new_[2514]_ ;
  assign \new_[4266]_  = ~\new_[1799]_ ;
  assign \new_[4267]_  = ~\new_[4310]_  | ~\new_[2514]_ ;
  assign \new_[4268]_  = ~\new_[4269]_  | (~\new_[2751]_  & ~\new_[4386]_ );
  assign \new_[4269]_  = ~\new_[2573]_  | ~\new_[4366]_ ;
  assign \new_[4270]_  = ~\new_[4271]_  | ~\new_[4272]_ ;
  assign \new_[4271]_  = \new_[2514]_  & \new_[3129]_ ;
  assign \new_[4272]_  = ~\new_[4273]_  | ~\new_[4274]_ ;
  assign \new_[4273]_  = ~\new_[4010]_  & ~\new_[3251]_ ;
  assign \new_[4274]_  = \new_[3823]_  & \new_[3908]_ ;
  assign n1651 = ~\new_[4381]_ ;
  assign n1581 = ~\new_[4277]_  | ~\new_[4279]_  | ~\new_[4283]_  | ~\new_[4278]_ ;
  assign \new_[4277]_  = ~\new_[2024]_ ;
  assign \new_[4278]_  = (~\new_[3975]_  | ~\new_[2620]_ ) & (~\new_[2592]_  | ~\new_[3986]_ );
  assign \new_[4279]_  = ~\new_[4282]_  & (~\new_[4280]_  | ~\new_[4281]_ );
  assign \new_[4280]_  = \new_[2662]_  & \new_[2938]_ ;
  assign \new_[4281]_  = ~\new_[1797]_ ;
  assign \new_[4282]_  = ~\new_[2617]_  | ~\new_[2599]_ ;
  assign \new_[4283]_  = (~\new_[4143]_  | ~\new_[2653]_ ) & (~\new_[4284]_  | ~\new_[4285]_ );
  assign \new_[4284]_  = \new_[2936]_  & \new_[2701]_ ;
  assign \new_[4285]_  = ~\new_[1886]_ ;
  assign \new_[4286]_  = ~\new_[4282]_ ;
  assign n1241 = ~\new_[4295]_  | (~\new_[4288]_  & ~\new_[4291]_ );
  assign \new_[4288]_  = ~\new_[4289]_ ;
  assign \new_[4289]_  = \new_[4290]_ ;
  assign \new_[4290]_  = ~\new_[4302]_ ;
  assign \new_[4291]_  = (~\new_[4292]_  | ~\new_[4296]_ ) & (~\new_[4293]_  | ~\new_[1234]_ );
  assign \new_[4292]_  = ~\new_[1607]_  | ~\new_[1721]_ ;
  assign \new_[4293]_  = \new_[4294]_ ;
  assign \new_[4294]_  = ~\new_[4130]_  | ~\new_[2403]_  | ~\new_[1604]_ ;
  assign \new_[4295]_  = ~\new_[2063]_  | ~\new_[4061]_ ;
  assign \new_[4296]_  = ~\new_[4294]_ ;
  assign n1446 = ~\new_[4298]_  | ~\new_[4303]_ ;
  assign \new_[4298]_  = ~\new_[4299]_  | ~\new_[4300]_ ;
  assign \new_[4299]_  = ~\new_[1667]_  | ~\new_[1639]_ ;
  assign \new_[4300]_  = ~\new_[4301]_  & ~\new_[2035]_ ;
  assign \new_[4301]_  = \new_[4302]_ ;
  assign \new_[4302]_  = ~\new_[3838]_  | ~\new_[2436]_ ;
  assign \new_[4303]_  = (~\new_[4057]_  | ~\new_[2063]_ ) & (~\new_[4304]_  | ~\new_[2035]_ );
  assign \new_[4304]_  = ~\new_[4305]_  & ~\new_[4301]_ ;
  assign \new_[4305]_  = ~\new_[1379]_ ;
  assign \new_[4306]_  = ~\new_[4307]_ ;
  assign \new_[4307]_  = ~\new_[4175]_  | ~\new_[2402]_  | ~\new_[2577]_ ;
  assign \new_[4308]_  = ~\new_[4309]_ ;
  assign \new_[4309]_  = ~\new_[4301]_ ;
  assign \new_[4310]_  = ~\new_[3838]_  | ~\new_[2436]_ ;
  assign \new_[4311]_  = ~\new_[4312]_  & ~\new_[4343]_ ;
  assign \new_[4312]_  = ~\new_[1876]_ ;
  assign \new_[4313]_  = \new_[4227]_  | \new_[4214]_ ;
  assign \new_[4314]_  = ~\new_[4329]_  | ~\new_[2030]_ ;
  assign \new_[4315]_  = ~\new_[3302]_  | ~\new_[3231]_ ;
  assign \new_[4316]_  = ~\new_[4320]_  & (~\new_[2626]_  | ~\new_[2855]_ );
  assign \new_[4317]_  = ~\new_[4364]_  | ~\new_[2837]_ ;
  assign \new_[4318]_  = ~\new_[4329]_  | ~\new_[2028]_ ;
  assign \new_[4319]_  = ~\new_[4333]_ ;
  assign \new_[4320]_  = ~\new_[4324]_  | ~\new_[4321]_  | ~\new_[4323]_ ;
  assign \new_[4321]_  = ~\new_[4322]_ ;
  assign \new_[4322]_  = ~\new_[2857]_  & ~\new_[2749]_ ;
  assign \new_[4323]_  = ~\new_[2730]_  & ~\new_[4243]_ ;
  assign \new_[4324]_  = \new_[4325]_  | \new_[4326]_ ;
  assign \new_[4325]_  = ~\new_[4345]_ ;
  assign \new_[4326]_  = ~\new_[2914]_  | ~\new_[2913]_ ;
  assign \new_[4327]_  = ~\new_[4324]_ ;
  assign \new_[4328]_  = \new_[4326]_ ;
  assign \new_[4329]_  = ~\new_[4334]_  | ~\new_[4330]_  | ~\new_[4332]_ ;
  assign \new_[4330]_  = ~\new_[4331]_  & ~\new_[4230]_ ;
  assign \new_[4331]_  = ~\new_[1499]_  | ~\new_[4239]_  | ~\new_[4240]_ ;
  assign \new_[4332]_  = ~\new_[1555]_  & ~\new_[4333]_ ;
  assign \new_[4333]_  = ~\new_[4133]_  | ~\new_[4071]_ ;
  assign \new_[4334]_  = \new_[4235]_  & \new_[4236]_ ;
  assign \new_[4335]_  = ~\new_[4336]_ ;
  assign \new_[4336]_  = ~\new_[4339]_  | ~\new_[4337]_  | ~\new_[4338]_ ;
  assign \new_[4337]_  = ~\new_[3921]_  & ~\new_[3898]_ ;
  assign \new_[4338]_  = ~\new_[3905]_ ;
  assign \new_[4339]_  = ~\new_[3888]_ ;
  assign \new_[4340]_  = ~\new_[4338]_  | ~\new_[4337]_ ;
  assign \new_[4341]_  = ~\new_[2634]_  | ~\new_[4237]_  | ~\new_[4226]_  | ~\new_[4319]_ ;
  assign \new_[4342]_  = ~\new_[4329]_  | ~\new_[1999]_ ;
  assign \new_[4343]_  = ~\new_[4351]_  | ~\new_[4344]_  | ~\new_[4345]_ ;
  assign \new_[4344]_  = ~\new_[4369]_ ;
  assign \new_[4345]_  = ~\new_[4346]_  & ~\new_[4347]_ ;
  assign \new_[4346]_  = ~\new_[3231]_  | ~\new_[3302]_ ;
  assign \new_[4347]_  = ~\new_[4313]_  | ~\new_[4314]_ ;
  assign \new_[4348]_  = ~\new_[4314]_  | ~\new_[4313]_ ;
  assign \new_[4349]_  = ~\new_[4350]_  & ~\new_[4384]_ ;
  assign \new_[4350]_  = ~\new_[4315]_  | ~\new_[4348]_ ;
  assign \new_[4351]_  = ~\new_[4352]_  & ~\new_[4353]_ ;
  assign \new_[4352]_  = ~\new_[4318]_  | ~\new_[4213]_ ;
  assign \new_[4353]_  = ~\new_[4342]_  | ~\new_[4341]_ ;
  assign \new_[4354]_  = \new_[4352]_ ;
  assign \new_[4355]_  = ~\new_[4194]_  | ~\new_[1239]_ ;
  assign \new_[4356]_  = ~\new_[4357]_ ;
  assign \new_[4357]_  = ~\new_[4372]_ ;
  assign \new_[4358]_  = ~\new_[4362]_  | ~\new_[4361]_  | ~\new_[4359]_  | ~\new_[4360]_ ;
  assign \new_[4359]_  = ~\new_[2545]_  & ~\new_[4246]_ ;
  assign \new_[4360]_  = \new_[4316]_  & \new_[4317]_ ;
  assign \new_[4361]_  = ~\new_[2513]_  & ~\new_[4268]_ ;
  assign \new_[4362]_  = ~\new_[4248]_  & ~\new_[2405]_ ;
  assign \new_[4363]_  = ~\new_[4364]_  | ~\new_[4366]_ ;
  assign \new_[4364]_  = ~\new_[4365]_ ;
  assign \new_[4365]_  = ~\new_[4208]_  | ~\new_[2818]_ ;
  assign \new_[4366]_  = ~\new_[4367]_ ;
  assign \new_[4367]_  = \new_[4368]_ ;
  assign \new_[4368]_  = \new_[4369]_ ;
  assign \new_[4369]_  = ~\new_[4370]_  | ~\new_[4371]_ ;
  assign \new_[4370]_  = ~\new_[3317]_  | ~\new_[2141]_ ;
  assign \new_[4371]_  = ~\new_[2645]_  | ~\new_[3355]_ ;
  assign \new_[4372]_  = \new_[4358]_ ;
  assign \new_[4373]_  = \new_[4358]_ ;
  assign \new_[4374]_  = ~\new_[4375]_ ;
  assign \new_[4375]_  = ~\new_[4284]_ ;
  assign n1361 = ~\new_[4377]_  | ~\new_[4381]_ ;
  assign \new_[4377]_  = ~\new_[4378]_ ;
  assign \new_[4378]_  = ~\new_[4379]_  | ~\new_[4380]_ ;
  assign \new_[4379]_  = ~\new_[2353]_  | ~\new_[3744]_ ;
  assign \new_[4380]_  = ~\new_[1553]_  | ~\new_[2372]_ ;
  assign \new_[4381]_  = ~\new_[4382]_  & (~\new_[2251]_  | ~\new_[3745]_ );
  assign \new_[4382]_  = \new_[2402]_  & \new_[2373]_ ;
  assign \new_[4383]_  = ~\new_[4385]_ ;
  assign \new_[4384]_  = ~\new_[4385]_ ;
  assign \new_[4385]_  = \new_[4351]_ ;
  assign \new_[4386]_  = ~\new_[2729]_ ;
  assign \new_[4387]_  = ~\new_[4388]_ ;
  assign \new_[4388]_  = ~\new_[4315]_ ;
  assign \new_[4389]_  = 1'b0;
  assign \new_[4390]_  = 1'b0;
  assign \new_[4391]_  = 1'b0;
  assign \new_[4392]_  = 1'b0;
  assign \new_[4393]_  = 1'b0;
  assign \new_[4394]_  = 1'b0;
  assign \new_[4395]_  = 1'b0;
  assign \new_[4396]_  = 1'b0;
  assign \new_[4397]_  = 1'b0;
  assign \new_[4398]_  = 1'b0;
  assign \new_[4399]_  = 1'b0;
  assign \new_[4400]_  = 1'b0;
  assign \new_[4401]_  = 1'b0;
  assign \new_[4402]_  = 1'b0;
  assign \new_[4403]_  = 1'b0;
  assign \new_[4404]_  = 1'b0;
  assign \new_[4405]_  = 1'b0;
  assign \new_[4406]_  = 1'b0;
  assign \new_[4407]_  = 1'b0;
  assign \new_[4408]_  = 1'b0;
  assign \new_[4409]_  = 1'b0;
  assign \new_[4410]_  = 1'b0;
  assign \new_[4411]_  = 1'b0;
  assign \new_[4412]_  = 1'b0;
  assign \new_[4413]_  = 1'b0;
  assign \new_[4414]_  = 1'b0;
  assign \new_[4415]_  = 1'b0;
  assign \new_[4416]_  = 1'b0;
  assign \new_[4417]_  = 1'b0;
  assign \new_[4418]_  = 1'b0;
  assign \new_[4419]_  = 1'b0;
  assign \new_[4420]_  = 1'b0;
  assign \new_[4421]_  = 1'b0;
  assign \new_[4422]_  = 1'b0;
  assign \new_[4423]_  = 1'b0;
  assign \new_[4424]_  = 1'b0;
  assign \new_[4425]_  = 1'b0;
  assign \new_[4426]_  = 1'b0;
  assign \new_[4427]_  = 1'b0;
  assign \new_[4428]_  = 1'b0;
  assign \new_[4429]_  = 1'b0;
  assign \new_[4430]_  = 1'b0;
  assign \new_[4431]_  = 1'b0;
  assign \new_[4432]_  = 1'b0;
  assign \new_[4433]_  = 1'b0;
  assign \new_[4434]_  = 1'b0;
  assign \new_[4435]_  = 1'b0;
  assign \new_[4436]_  = 1'b0;
  assign \new_[4437]_  = 1'b0;
  assign \new_[4438]_  = 1'b0;
  assign \new_[4439]_  = 1'b0;
  assign \new_[4440]_  = 1'b0;
  assign \new_[4441]_  = 1'b0;
  assign \new_[4442]_  = 1'b0;
  assign \new_[4443]_  = 1'b0;
  assign \new_[4444]_  = 1'b0;
  assign \new_[4445]_  = 1'b0;
  assign \new_[4446]_  = 1'b0;
  assign \new_[4447]_  = 1'b0;
  assign \new_[4448]_  = 1'b0;
  assign n1196 = n1201;
  assign n3481 = \wb0_addr_i[3] ;
  assign n3486 = \wb0m_data_i[4] ;
  assign n3491 = \wb0m_data_i[0] ;
  assign n3496 = \wb0m_data_i[18] ;
  assign n3501 = \wb0m_data_i[7] ;
  assign n3506 = \wb0_addr_i[6] ;
  assign n3511 = \wb0m_data_i[5] ;
  assign n3516 = \wb0m_data_i[24] ;
  assign n3521 = \wb0m_data_i[1] ;
  assign n3526 = \wb0_addr_i[8] ;
  assign n3531 = \wb0m_data_i[19] ;
  assign n3536 = \wb0m_data_i[31] ;
  assign n3541 = \wb0m_data_i[6] ;
  assign n3546 = \wb0_addr_i[9] ;
  assign n3551 = \wb0m_data_i[20] ;
  assign n3556 = \wb0_addr_i[4] ;
  assign n3561 = \wb0m_data_i[30] ;
  assign n3566 = \wb0m_data_i[26] ;
  assign n3571 = \wb0m_data_i[29] ;
  assign n3576 = \wb0m_data_i[28] ;
  assign n3581 = \wb0m_data_i[2] ;
  assign n3586 = \wb0m_data_i[8] ;
  assign n3591 = \wb0_addr_i[7] ;
  assign n3596 = \wb0_addr_i[2] ;
  assign n3601 = \wb0m_data_i[14] ;
  assign n3606 = \wb0m_data_i[23] ;
  assign n3611 = \wb0m_data_i[9] ;
  assign n3616 = \wb0m_data_i[21] ;
  assign n3621 = \wb0m_data_i[25] ;
  assign n3626 = \wb0m_data_i[27] ;
  assign n3631 = \wb0m_data_i[3] ;
  assign n3636 = \wb0m_data_i[12] ;
  assign n3641 = \wb0m_data_i[17] ;
  assign n3646 = \wb0_addr_i[5] ;
  assign n3651 = \wb0m_data_i[11] ;
  assign n3656 = \wb0m_data_i[15] ;
  assign n3661 = \wb0m_data_i[13] ;
  assign n3666 = \wb0m_data_i[10] ;
  assign n3671 = \wb0m_data_i[16] ;
  assign n3676 = \wb0m_data_i[22] ;
  always @ (posedge clock) begin
    u3_u0_mast_stb_reg <= n866;
    u4_u0_mast_stb_reg <= n871;
    u3_u0_mast_cyc_reg <= n876;
    u4_u0_mast_cyc_reg <= n881;
    \\u2_mast0_adr_reg[3]  <= n886;
    \\u2_mast0_adr_reg[2]  <= n891;
    \\u2_mast0_adr_reg[23]  <= n896;
    \\u2_mast0_adr_reg[22]  <= n901;
    \\u2_mast0_adr_reg[21]  <= n906;
    \\u2_mast0_adr_reg[25]  <= n911;
    \\u2_mast0_adr_reg[20]  <= n916;
    \\u2_mast0_adr_reg[19]  <= n921;
    \\u2_mast0_adr_reg[18]  <= n926;
    \\u2_mast0_adr_reg[16]  <= n931;
    \\u2_mast0_adr_reg[15]  <= n936;
    \\u2_mast0_adr_reg[14]  <= n941;
    \\u2_mast0_adr_reg[13]  <= n946;
    \\u2_mast0_adr_reg[12]  <= n951;
    \\u2_mast0_adr_reg[11]  <= n956;
    \\u2_mast0_adr_reg[10]  <= n961;
    \\u2_mast0_adr_reg[9]  <= n966;
    \\u2_mast0_adr_reg[6]  <= n971;
    \\u2_mast0_adr_reg[5]  <= n976;
    \\u2_mast0_adr_reg[4]  <= n981;
    \\u2_mast0_adr_reg[29]  <= n986;
    \\u2_mast0_adr_reg[28]  <= n991;
    \\u2_mast0_adr_reg[27]  <= n996;
    \\u2_mast0_adr_reg[26]  <= n1001;
    \\u2_mast0_adr_reg[24]  <= n1006;
    \\u2_mast0_adr_reg[17]  <= n1011;
    \\u2_mast0_adr_reg[7]  <= n1016;
    \\u2_mast0_adr_reg[8]  <= n1021;
    \\u2_mast1_adr_reg[29]  <= n1026;
    \\u2_mast1_adr_reg[28]  <= n1031;
    \\u2_mast1_adr_reg[27]  <= n1036;
    \\u2_mast1_adr_reg[26]  <= n1041;
    \\u2_mast1_adr_reg[25]  <= n1046;
    \\u2_mast1_adr_reg[24]  <= n1051;
    \\u2_mast1_adr_reg[22]  <= n1056;
    \\u2_mast1_adr_reg[23]  <= n1061;
    \\u2_mast1_adr_reg[21]  <= n1066;
    \\u2_mast1_adr_reg[20]  <= n1071;
    \\u2_mast1_adr_reg[19]  <= n1076;
    \\u2_mast1_adr_reg[18]  <= n1081;
    \\u2_mast1_adr_reg[16]  <= n1086;
    \\u2_mast1_adr_reg[15]  <= n1091;
    \\u2_mast1_adr_reg[13]  <= n1096;
    \\u2_mast1_adr_reg[12]  <= n1101;
    \\u2_mast1_adr_reg[14]  <= n1106;
    \\u2_mast1_adr_reg[11]  <= n1111;
    \\u2_mast1_adr_reg[10]  <= n1116;
    \\u2_mast1_adr_reg[9]  <= n1121;
    \\u2_mast1_adr_reg[6]  <= n1126;
    \\u2_mast1_adr_reg[5]  <= n1131;
    \\u2_mast1_adr_reg[4]  <= n1136;
    \\u2_mast0_adr_reg[31]  <= n1141;
    \\u2_mast0_adr_reg[30]  <= n1146;
    \\u2_mast1_adr_reg[31]  <= n1151;
    \\u2_mast1_adr_reg[30]  <= n1156;
    \\u2_mast1_adr_reg[17]  <= n1161;
    \\u2_mast1_adr_reg[8]  <= n1166;
    \\u2_mast1_adr_reg[7]  <= n1171;
    \\u2_mast1_adr_reg[3]  <= n1176;
    \\u2_mast1_adr_reg[2]  <= n1181;
    \\u2_state_reg[1]  <= n1186;
    \\u2_state_reg[3]  <= n1191;
    u2_chunk_dec_reg <= n1196;
    u2_tsz_dec_reg <= n1201;
    \\u2_adr1_cnt_reg[28]  <= n1206;
    \\u2_adr1_cnt_reg[27]  <= n1211;
    \\u2_adr1_cnt_reg[23]  <= n1216;
    \\u2_adr1_cnt_reg[24]  <= n1221;
    \\u2_adr1_cnt_reg[20]  <= n1226;
    \\u2_adr1_cnt_reg[19]  <= n1231;
    \\u2_adr1_cnt_reg[18]  <= n1236;
    \\u2_adr1_cnt_reg[25]  <= n1241;
    \\u2_adr1_cnt_reg[29]  <= n1246;
    \\u2_adr1_cnt_reg[17]  <= n1251;
    \\u2_adr1_cnt_reg[21]  <= n1256;
    \\u2_adr1_cnt_reg[16]  <= n1261;
    \\u2_adr1_cnt_reg[2]  <= n1266;
    \\u2_adr1_cnt_reg[3]  <= n1271;
    \\u2_adr1_cnt_reg[4]  <= n1276;
    \\u2_adr1_cnt_reg[5]  <= n1281;
    \\u2_adr1_cnt_reg[6]  <= n1286;
    \\u2_adr1_cnt_reg[7]  <= n1291;
    \\u2_adr1_cnt_reg[8]  <= n1296;
    \\u2_adr1_cnt_reg[9]  <= n1301;
    \\u2_adr1_cnt_reg[10]  <= n1306;
    \\u2_adr1_cnt_reg[11]  <= n1311;
    \\u2_adr1_cnt_reg[13]  <= n1316;
    \\u2_adr1_cnt_reg[14]  <= n1321;
    \\u2_adr1_cnt_reg[15]  <= n1326;
    u2_read_r_reg <= n1331;
    \\u2_adr1_cnt_reg[26]  <= n1336;
    \\u2_adr1_cnt_reg[22]  <= n1341;
    \\u2_adr1_cnt_reg[0]  <= n1346;
    \\u2_adr1_cnt_reg[12]  <= n1351;
    \\u2_adr1_cnt_reg[1]  <= n1356;
    u2_write_hold_r_reg <= n1361;
    u3_u0_mast_we_r_reg <= n1366;
    \\u2_adr0_cnt_reg[16]  <= n1371;
    \\u0_u0_int_src_r_reg[2]  <= n1376;
    \\u1_ack_o_reg[0]  <= n1381;
    u1_next_start_reg <= n1386;
    \\u2_adr0_cnt_reg[9]  <= n1391;
    \\u2_adr0_cnt_reg[28]  <= n1396;
    \\u2_adr0_cnt_reg[27]  <= n1401;
    \\u2_adr0_cnt_reg[24]  <= n1406;
    \\u2_adr0_cnt_reg[23]  <= n1411;
    \\u2_adr0_cnt_reg[26]  <= n1416;
    \\u2_adr0_cnt_reg[20]  <= n1421;
    \\u2_adr0_cnt_reg[18]  <= n1426;
    \\u2_adr0_cnt_reg[10]  <= n1431;
    \\u2_adr0_cnt_reg[11]  <= n1436;
    \\u2_adr0_cnt_reg[12]  <= n1441;
    \\u2_adr0_cnt_reg[13]  <= n1446;
    \\u2_adr0_cnt_reg[17]  <= n1451;
    \\u2_adr0_cnt_reg[21]  <= n1456;
    \\u2_adr0_cnt_reg[25]  <= n1461;
    \\u2_adr0_cnt_reg[2]  <= n1466;
    \\u2_adr0_cnt_reg[3]  <= n1471;
    \\u2_adr0_cnt_reg[5]  <= n1476;
    \\u2_adr0_cnt_reg[6]  <= n1481;
    \\u2_adr0_cnt_reg[8]  <= n1486;
    \\u2_adr0_cnt_reg[7]  <= n1491;
    \\u2_adr0_cnt_reg[4]  <= n1496;
    \\u0_u0_ch_csr_r_reg[0]  <= n1501;
    \\u2_adr0_cnt_reg[14]  <= n1506;
    \\u2_adr0_cnt_reg[22]  <= n1511;
    \\u2_adr0_cnt_reg[19]  <= n1516;
    \\u2_adr0_cnt_reg[29]  <= n1521;
    \\u2_adr0_cnt_reg[15]  <= n1526;
    u0_u0_ch_done_reg <= n1531;
    u2_next_ch_reg <= n1536;
    \\u0_u0_int_src_r_reg[1]  <= n1541;
    \\u2_state_reg[0]  <= n1546;
    \\u2_state_reg[9]  <= n1551;
    \\u2_adr0_cnt_reg[0]  <= n1556;
    \\u2_adr0_cnt_reg[1]  <= n1561;
    \\u2_tsz_cnt_reg[8]  <= n1566;
    \\u2_tsz_cnt_reg[2]  <= n1571;
    u4_u0_mast_we_r_reg <= n1576;
    \\u0_wb_rf_dout_reg[10]  <= n1581;
    \\u2_state_reg[10]  <= n1586;
    \\u2_state_reg[4]  <= n1591;
    \\u2_tsz_cnt_reg[0]  <= n1596;
    \\u2_tsz_cnt_reg[4]  <= n1601;
    \\u2_tsz_cnt_reg[5]  <= n1606;
    \\u2_tsz_cnt_reg[6]  <= n1611;
    \\u2_tsz_cnt_reg[7]  <= n1616;
    \\u2_tsz_cnt_reg[10]  <= n1621;
    \\u2_tsz_cnt_reg[11]  <= n1626;
    \\u2_tsz_cnt_reg[1]  <= n1631;
    \\u2_tsz_cnt_reg[3]  <= n1636;
    \\u2_tsz_cnt_reg[9]  <= n1641;
    u2_chunk_0_reg <= n1646;
    u2_write_r_reg <= n1651;
    \\u2_state_reg[2]  <= n1656;
    \\u0_u0_ch_tot_sz_r_reg[0]  <= n1661;
    \\u0_u0_ch_adr1_r_reg[25]  <= n1666;
    \\u0_u0_ch_adr0_r_reg[17]  <= n1671;
    \\u0_u0_ch_adr0_r_reg[13]  <= n1676;
    \\u0_u0_ch_adr1_r_reg[29]  <= n1681;
    \\u0_u0_ch_adr1_r_reg[21]  <= n1686;
    \\u0_u0_ch_adr1_r_reg[13]  <= n1691;
    \\u0_u0_ch_adr1_r_reg[17]  <= n1696;
    \\u0_u0_ch_tot_sz_r_reg[1]  <= n1701;
    \\u0_u0_ch_adr1_r_reg[10]  <= n1706;
    \\u0_u0_ch_adr1_r_reg[11]  <= n1711;
    \\u0_u0_ch_adr1_r_reg[12]  <= n1716;
    \\u0_u0_ch_adr1_r_reg[14]  <= n1721;
    \\u0_u0_ch_adr1_r_reg[15]  <= n1726;
    \\u0_u0_ch_adr1_r_reg[16]  <= n1731;
    \\u0_u0_ch_adr1_r_reg[18]  <= n1736;
    \\u0_u0_ch_adr1_r_reg[19]  <= n1741;
    \\u0_u0_ch_adr1_r_reg[20]  <= n1746;
    \\u0_u0_ch_adr1_r_reg[22]  <= n1751;
    \\u0_u0_ch_adr1_r_reg[23]  <= n1756;
    \\u0_u0_ch_adr1_r_reg[24]  <= n1761;
    \\u0_u0_ch_adr1_r_reg[26]  <= n1766;
    \\u0_u0_ch_adr1_r_reg[27]  <= n1771;
    \\u0_u0_ch_adr1_r_reg[28]  <= n1776;
    \\u0_u0_ch_adr0_r_reg[10]  <= n1781;
    \\u0_u0_ch_adr0_r_reg[11]  <= n1786;
    \\u0_u0_ch_adr0_r_reg[12]  <= n1791;
    \\u0_u0_ch_adr0_r_reg[14]  <= n1796;
    \\u0_u0_ch_adr0_r_reg[15]  <= n1801;
    \\u0_u0_ch_adr0_r_reg[16]  <= n1806;
    \\u0_u0_ch_adr0_r_reg[18]  <= n1811;
    \\u0_u0_ch_adr0_r_reg[19]  <= n1816;
    \\u0_u0_ch_adr0_r_reg[20]  <= n1821;
    \\u0_u0_ch_adr0_r_reg[22]  <= n1826;
    \\u0_u0_ch_adr0_r_reg[23]  <= n1831;
    \\u0_u0_ch_adr0_r_reg[24]  <= n1836;
    \\u0_u0_ch_adr0_r_reg[26]  <= n1841;
    \\u0_u0_ch_adr0_r_reg[27]  <= n1846;
    \\u0_u0_ch_adr0_r_reg[28]  <= n1851;
    \\u0_u0_ch_adr0_r_reg[21]  <= n1856;
    \\u0_u0_ch_adr0_r_reg[29]  <= n1861;
    \\u0_u0_ch_adr0_r_reg[25]  <= n1866;
    \\u0_u0_ch_tot_sz_r_reg[9]  <= n1871;
    \\u0_u0_ch_tot_sz_r_reg[5]  <= n1876;
    \\u0_u0_ch_tot_sz_r_reg[10]  <= n1881;
    \\u0_u0_ch_tot_sz_r_reg[11]  <= n1886;
    \\u0_u0_ch_tot_sz_r_reg[2]  <= n1891;
    \\u0_u0_ch_tot_sz_r_reg[3]  <= n1896;
    \\u0_u0_ch_tot_sz_r_reg[4]  <= n1901;
    \\u0_u0_ch_tot_sz_r_reg[6]  <= n1906;
    \\u0_u0_ch_tot_sz_r_reg[7]  <= n1911;
    \\u0_u0_ch_tot_sz_r_reg[8]  <= n1916;
    \\u0_u0_ch_csr_r_reg[4]  <= n1921;
    u0_u0_ch_err_reg <= n1926;
    \\u0_u0_ch_csr_r_reg[1]  <= n1931;
    \\u0_u0_ch_csr_r_reg[2]  <= n1936;
    \\u0_u0_ch_csr_r_reg[3]  <= n1941;
    \\u0_u0_ch_adr1_r_reg[0]  <= n1946;
    \\u0_u0_ch_adr1_r_reg[1]  <= n1951;
    \\u0_u0_ch_adr1_r_reg[3]  <= n1956;
    \\u0_u0_ch_adr1_r_reg[4]  <= n1961;
    \\u0_u0_ch_adr1_r_reg[5]  <= n1966;
    \\u0_u0_ch_adr1_r_reg[7]  <= n1971;
    \\u0_u0_ch_adr1_r_reg[8]  <= n1976;
    \\u0_u0_ch_adr1_r_reg[9]  <= n1981;
    \\u0_u0_ch_adr0_r_reg[9]  <= n1986;
    \\u0_u0_ch_adr0_r_reg[0]  <= n1991;
    \\u0_u0_ch_adr0_r_reg[1]  <= n1996;
    \\u0_u0_ch_adr0_r_reg[3]  <= n2001;
    \\u0_u0_ch_adr0_r_reg[4]  <= n2006;
    \\u0_u0_ch_adr0_r_reg[5]  <= n2011;
    \\u0_u0_ch_adr0_r_reg[7]  <= n2016;
    \\u0_u0_int_src_r_reg[0]  <= n2021;
    \\u0_u0_ch_adr0_r_reg[6]  <= n2026;
    \\u0_u0_ch_adr0_r_reg[2]  <= n2031;
    \\u0_u0_ch_adr0_r_reg[8]  <= n2036;
    \\u0_u0_ch_adr1_r_reg[6]  <= n2041;
    \\u0_u0_ch_adr1_r_reg[2]  <= n2046;
    \\u2_chunk_cnt_reg[8]  <= n2051;
    \\u2_chunk_cnt_reg[7]  <= n2056;
    \\u2_chunk_cnt_reg[6]  <= n2061;
    \\u1_ch_sel_r_reg[2]  <= n2066;
    \\u1_ch_sel_r_reg[1]  <= n2071;
    \\u1_ch_sel_r_reg[3]  <= n2076;
    \\u1_ch_sel_r_reg[4]  <= n2081;
    \\u2_chunk_cnt_reg[1]  <= n2086;
    \\u2_chunk_cnt_reg[3]  <= n2091;
    \\u2_chunk_cnt_reg[4]  <= n2096;
    \\u2_chunk_cnt_reg[0]  <= n2101;
    \\u2_chunk_cnt_reg[5]  <= n2106;
    \\u2_chunk_cnt_reg[2]  <= n2111;
    \\u1_ch_sel_r_reg[0]  <= n2116;
    \\u0_wb_rf_dout_reg[26]  <= n2121;
    \\u0_wb_rf_dout_reg[25]  <= n2126;
    \\u0_wb_rf_dout_reg[24]  <= n2131;
    \\u0_wb_rf_dout_reg[23]  <= n2136;
    \\u0_wb_rf_dout_reg[14]  <= n2141;
    \\u0_wb_rf_dout_reg[13]  <= n2146;
    \\u0_wb_rf_dout_reg[12]  <= n2151;
    \\u0_wb_rf_dout_reg[3]  <= n2156;
    \\u0_wb_rf_dout_reg[2]  <= n2161;
    \\u0_wb_rf_dout_reg[0]  <= n2166;
    \\u0_wb_rf_dout_reg[22]  <= n2171;
    \\u0_wb_rf_dout_reg[21]  <= n2176;
    \\u0_wb_rf_dout_reg[20]  <= n2181;
    \\u0_wb_rf_dout_reg[19]  <= n2186;
    \\u0_wb_rf_dout_reg[18]  <= n2191;
    \\u0_wb_rf_dout_reg[17]  <= n2196;
    \\u0_wb_rf_dout_reg[16]  <= n2201;
    \\u0_wb_rf_dout_reg[15]  <= n2206;
    \\u0_wb_rf_dout_reg[11]  <= n2211;
    \\u0_wb_rf_dout_reg[8]  <= n2216;
    \\u0_wb_rf_dout_reg[7]  <= n2221;
    \\u0_wb_rf_dout_reg[6]  <= n2226;
    \\u0_wb_rf_dout_reg[5]  <= n2231;
    \\u0_wb_rf_dout_reg[4]  <= n2236;
    u0_u0_ch_busy_reg <= n2241;
    \\u0_wb_rf_dout_reg[9]  <= n2246;
    \\u0_wb_rf_dout_reg[30]  <= n2251;
    \\u0_wb_rf_dout_reg[29]  <= n2256;
    \\u0_wb_rf_dout_reg[28]  <= n2261;
    \\u0_wb_rf_dout_reg[27]  <= n2266;
    \\u0_wb_rf_dout_reg[1]  <= n2271;
    \\u0_wb_rf_dout_reg[31]  <= n2276;
    u2_tsz_cnt_is_0_r_reg <= n2281;
    u2_dma_abort_r_reg <= n2286;
    u1_de_start_r_reg <= n2291;
    \\u2_state_reg[5]  <= n2296;
    \\u0_u0_ch_csr_r3_reg[2]  <= n2301;
    \\u0_u0_ch_csr_r3_reg[0]  <= n2306;
    u0_u0_rest_en_reg <= n2311;
    \\u0_u0_ch_csr_r_reg[7]  <= n2316;
    \\u0_u0_ch_csr_r_reg[5]  <= n2321;
    \\u0_u0_ch_csr_r2_reg[2]  <= n2326;
    \\u0_u0_ch_csr_r2_reg[1]  <= n2331;
    \\u0_u0_ch_csr_r2_reg[0]  <= n2336;
    \\u0_u0_ch_csr_r3_reg[1]  <= n2341;
    \\u0_u0_ch_csr_r_reg[6]  <= n2346;
    \\u0_u0_ch_csr_r_reg[8]  <= n2351;
    u0_u0_ch_stop_reg <= n2356;
    u0_u0_ch_sz_inf_reg <= n2361;
    \\u1_u1_state_reg[2]  <= n2366;
    \\u1_u1_state_reg[3]  <= n2371;
    \\u0_u0_ch_chk_sz_r_reg[5]  <= n2376;
    \\u0_u0_ch_chk_sz_r_reg[3]  <= n2381;
    \\u0_u0_ch_chk_sz_r_reg[7]  <= n2386;
    \\u0_u0_ch_chk_sz_r_reg[1]  <= n2391;
    \\u0_u0_ch_chk_sz_r_reg[2]  <= n2396;
    \\u1_u1_state_reg[4]  <= n2401;
    \\u0_u0_ch_chk_sz_r_reg[4]  <= n2406;
    \\u0_u0_ch_chk_sz_r_reg[6]  <= n2411;
    \\u0_u0_ch_chk_sz_r_reg[0]  <= n2416;
    \\u1_u1_state_reg[0]  <= n2421;
    \\u1_u1_state_reg[1]  <= n2426;
    u4_u1_rf_ack_reg <= n2431;
    \\u0_u0_ch_chk_sz_r_reg[10]  <= n2436;
    \\u0_u0_ch_chk_sz_r_reg[8]  <= n2441;
    \\u0_u0_ch_chk_sz_r_reg[9]  <= n2446;
    \\u2_u0_out_r_reg[15]  <= n2451;
    \\u2_u1_out_r_reg[15]  <= n2456;
    \\u2_state_reg[8]  <= n2461;
    \\u2_state_reg[7]  <= n2466;
    \\u2_state_reg[6]  <= n2471;
    \\u2_u0_out_r_reg[11]  <= n2476;
    \\u2_u1_out_r_reg[11]  <= n2481;
    \\u2_u0_out_r_reg[12]  <= n2486;
    \\u2_u1_out_r_reg[12]  <= n2491;
    \\u2_u0_out_r_reg[16]  <= n2496;
    \\u2_u1_out_r_reg[16]  <= n2501;
    \\u0_int_maska_r_reg[11]  <= n2506;
    \\u0_csr_r_reg[0]  <= n2511;
    \\u0_int_maska_r_reg[0]  <= n2516;
    \\u2_u0_out_r_reg[14]  <= n2521;
    \\u2_u1_out_r_reg[14]  <= n2526;
    \\u0_int_maska_r_reg[10]  <= n2531;
    \\u0_int_maska_r_reg[5]  <= n2536;
    \\u2_u1_out_r_reg[8]  <= n2541;
    \\u2_u0_out_r_reg[8]  <= n2546;
    \\u0_int_maska_r_reg[6]  <= n2551;
    \\u0_int_maska_r_reg[7]  <= n2556;
    \\u0_int_maska_r_reg[8]  <= n2561;
    \\u0_int_maska_r_reg[9]  <= n2566;
    \\u0_int_maska_r_reg[2]  <= n2571;
    \\u0_int_maska_r_reg[4]  <= n2576;
    \\u0_int_maska_r_reg[3]  <= n2581;
    \\u0_int_maska_r_reg[29]  <= n2586;
    \\u0_int_maska_r_reg[26]  <= n2591;
    \\u0_int_maska_r_reg[27]  <= n2596;
    \\u0_int_maska_r_reg[28]  <= n2601;
    \\u0_int_maska_r_reg[19]  <= n2606;
    \\u0_int_maska_r_reg[22]  <= n2611;
    \\u0_int_maska_r_reg[24]  <= n2616;
    \\u0_int_maska_r_reg[23]  <= n2621;
    \\u0_int_maska_r_reg[1]  <= n2626;
    \\u0_int_maska_r_reg[20]  <= n2631;
    \\u0_int_maska_r_reg[16]  <= n2636;
    \\u0_int_maska_r_reg[17]  <= n2641;
    \\u0_int_maska_r_reg[15]  <= n2646;
    \\u0_int_maska_r_reg[12]  <= n2651;
    \\u0_int_maska_r_reg[13]  <= n2656;
    \\u0_int_maska_r_reg[14]  <= n2661;
    \\u0_int_maskb_r_reg[6]  <= n2666;
    \\u0_int_maskb_r_reg[9]  <= n2671;
    \\u2_u1_out_r_reg[7]  <= n2676;
    \\u2_u0_out_r_reg[7]  <= n2681;
    \\u0_int_maska_r_reg[18]  <= n2686;
    \\u0_int_maska_r_reg[21]  <= n2691;
    \\u0_int_maska_r_reg[25]  <= n2696;
    \\u0_int_maska_r_reg[30]  <= n2701;
    \\u0_int_maskb_r_reg[0]  <= n2706;
    \\u0_int_maskb_r_reg[7]  <= n2711;
    \\u0_int_maskb_r_reg[8]  <= n2716;
    \\u0_int_maskb_r_reg[5]  <= n2721;
    \\u0_int_maskb_r_reg[11]  <= n2726;
    \\u0_int_maskb_r_reg[10]  <= n2731;
    \\u0_int_maskb_r_reg[14]  <= n2736;
    \\u0_int_maskb_r_reg[17]  <= n2741;
    \\u0_int_maskb_r_reg[20]  <= n2746;
    \\u0_int_maskb_r_reg[22]  <= n2751;
    \\u0_int_maskb_r_reg[2]  <= n2756;
    \\u0_int_maskb_r_reg[12]  <= n2761;
    \\u0_int_maskb_r_reg[18]  <= n2766;
    \\u0_int_maskb_r_reg[19]  <= n2771;
    \\u0_int_maskb_r_reg[15]  <= n2776;
    \\u2_u0_out_r_reg[13]  <= n2781;
    \\u2_u1_out_r_reg[13]  <= n2786;
    \\u0_int_maskb_r_reg[24]  <= n2791;
    \\u0_int_maskb_r_reg[30]  <= n2796;
    \\u0_int_maskb_r_reg[3]  <= n2801;
    \\u0_int_maskb_r_reg[4]  <= n2806;
    \\u0_int_maskb_r_reg[25]  <= n2811;
    \\u0_int_maskb_r_reg[28]  <= n2816;
    \\u0_int_maskb_r_reg[29]  <= n2821;
    \\u0_int_maskb_r_reg[26]  <= n2826;
    \\u0_int_maskb_r_reg[27]  <= n2831;
    \\u0_int_maskb_r_reg[23]  <= n2836;
    \\u0_int_maskb_r_reg[1]  <= n2841;
    \\u0_int_maskb_r_reg[21]  <= n2846;
    \\u0_int_maskb_r_reg[16]  <= n2851;
    \\u0_int_maskb_r_reg[13]  <= n2856;
    u2_chunk_cnt_is_0_r_reg <= n2861;
    \\u2_u1_out_r_reg[4]  <= n2866;
    \\u2_u0_out_r_reg[4]  <= n2871;
    \\u2_u1_out_r_reg[10]  <= n2876;
    \\u2_u0_out_r_reg[10]  <= n2881;
    u4_u1_slv_we_reg <= n2886;
    u3_u1_slv_re_reg <= n2891;
    u4_u1_slv_re_reg <= n2896;
    u3_u1_slv_we_reg <= n2901;
    \\u3_u0_mast_dout_reg[4]  <= n2906;
    \\u3_u0_mast_dout_reg[28]  <= n2911;
    \\u3_u0_mast_dout_reg[19]  <= n2916;
    \\u3_u0_mast_dout_reg[29]  <= n2921;
    u0_inta_o_reg <= n2926;
    \\u3_u0_mast_dout_reg[1]  <= n2931;
    \\u3_u0_mast_dout_reg[8]  <= n2936;
    \\u3_u0_mast_dout_reg[30]  <= n2941;
    \\u3_u0_mast_dout_reg[3]  <= n2946;
    \\u3_u0_mast_dout_reg[22]  <= n2951;
    \\u3_u0_mast_dout_reg[18]  <= n2956;
    \\u3_u0_mast_dout_reg[10]  <= n2961;
    \\u3_u0_mast_dout_reg[12]  <= n2966;
    \\u3_u0_mast_dout_reg[0]  <= n2971;
    \\u3_u0_mast_dout_reg[15]  <= n2976;
    \\u3_u0_mast_dout_reg[20]  <= n2981;
    \\u3_u0_mast_dout_reg[25]  <= n2986;
    \\u3_u0_mast_dout_reg[14]  <= n2991;
    \\u3_u0_mast_dout_reg[9]  <= n2996;
    \\u3_u0_mast_dout_reg[13]  <= n3001;
    \\u3_u0_mast_dout_reg[11]  <= n3006;
    \\u3_u0_mast_dout_reg[17]  <= n3011;
    \\u3_u0_mast_dout_reg[2]  <= n3016;
    \\u2_u1_out_r_reg[3]  <= n3021;
    \\u3_u0_mast_dout_reg[31]  <= n3026;
    \\u3_u0_mast_dout_reg[6]  <= n3031;
    \\u3_u0_mast_dout_reg[27]  <= n3036;
    \\u3_u0_mast_dout_reg[23]  <= n3041;
    \\u3_u0_mast_dout_reg[24]  <= n3046;
    u0_intb_o_reg <= n3051;
    \\u2_u0_out_r_reg[3]  <= n3056;
    \\u3_u0_mast_dout_reg[21]  <= n3061;
    \\u3_u0_mast_dout_reg[7]  <= n3066;
    \\u2_u1_out_r_reg[6]  <= n3071;
    \\u2_u0_out_r_reg[6]  <= n3076;
    \\u3_u0_mast_dout_reg[5]  <= n3081;
    \\u2_u1_out_r_reg[9]  <= n3086;
    \\u2_u0_out_r_reg[9]  <= n3091;
    \\u3_u0_mast_dout_reg[26]  <= n3096;
    \\u3_u0_mast_dout_reg[16]  <= n3101;
    \\u2_u0_out_r_reg[5]  <= n3106;
    \\u2_u1_out_r_reg[5]  <= n3111;
    \\u2_u1_out_r_reg[2]  <= n3116;
    \\u2_u0_out_r_reg[2]  <= n3121;
    u2_mast0_drdy_r_reg <= n3126;
    u3_u1_rf_ack_reg <= n3131;
    \\u4_u0_mast_dout_reg[23]  <= n3136;
    \\u4_u0_mast_dout_reg[20]  <= n3141;
    \\u4_u0_mast_dout_reg[16]  <= n3146;
    \\u4_u0_mast_dout_reg[22]  <= n3151;
    \\u4_u0_mast_dout_reg[5]  <= n3156;
    \\u4_u0_mast_dout_reg[11]  <= n3161;
    \\u4_u0_mast_dout_reg[12]  <= n3166;
    \\u4_u0_mast_dout_reg[7]  <= n3171;
    \\u4_u0_mast_dout_reg[3]  <= n3176;
    \\u4_u0_mast_dout_reg[13]  <= n3181;
    \\u4_u0_mast_dout_reg[4]  <= n3186;
    \\u4_u0_mast_dout_reg[27]  <= n3191;
    \\u4_u0_mast_dout_reg[1]  <= n3196;
    \\u4_u0_mast_dout_reg[26]  <= n3201;
    \\u4_u0_mast_dout_reg[25]  <= n3206;
    \\u4_u0_mast_dout_reg[21]  <= n3211;
    \\u4_u0_mast_dout_reg[2]  <= n3216;
    \\u4_u0_mast_dout_reg[24]  <= n3221;
    \\u4_u0_mast_dout_reg[0]  <= n3226;
    \\u4_u0_mast_dout_reg[17]  <= n3231;
    \\u4_u0_mast_dout_reg[31]  <= n3236;
    \\u4_u0_mast_dout_reg[14]  <= n3241;
    \\u4_u0_mast_dout_reg[8]  <= n3246;
    \\u4_u0_mast_dout_reg[28]  <= n3251;
    \\u4_u0_mast_dout_reg[10]  <= n3256;
    \\u4_u0_mast_dout_reg[18]  <= n3261;
    \\u4_u0_mast_dout_reg[29]  <= n3266;
    \\u4_u0_mast_dout_reg[6]  <= n3271;
    \\u4_u0_mast_dout_reg[9]  <= n3276;
    \\u4_u0_mast_dout_reg[19]  <= n3281;
    \\u4_u0_mast_dout_reg[15]  <= n3286;
    \\u4_u0_mast_dout_reg[30]  <= n3291;
    \\u2_u0_out_r_reg[1]  <= n3296;
    \\u2_u1_out_r_reg[1]  <= n3301;
    \\u1_ndr_r_reg[2]  <= n3306;
    \\u1_ndr_r_reg[1]  <= n3311;
    \\u1_ndr_r_reg[24]  <= n3316;
    \\u1_ndr_r_reg[10]  <= n3321;
    \\u1_ndr_r_reg[11]  <= n3326;
    \\u1_ndr_r_reg[12]  <= n3331;
    \\u1_ndr_r_reg[29]  <= n3336;
    \\u1_ndr_r_reg[17]  <= n3341;
    \\u1_ndr_r_reg[9]  <= n3346;
    \\u1_ndr_r_reg[22]  <= n3351;
    \\u1_ndr_r_reg[7]  <= n3356;
    \\u1_ndr_r_reg[30]  <= n3361;
    \\u1_ndr_r_reg[23]  <= n3366;
    \\u1_ndr_r_reg[15]  <= n3371;
    \\u1_ndr_r_reg[14]  <= n3376;
    \\u1_ndr_r_reg[28]  <= n3381;
    \\u1_ndr_r_reg[18]  <= n3386;
    \\u1_ndr_r_reg[16]  <= n3391;
    \\u1_ndr_r_reg[8]  <= n3396;
    \\u1_ndr_r_reg[4]  <= n3401;
    \\u1_ndr_r_reg[27]  <= n3406;
    \\u1_ndr_r_reg[20]  <= n3411;
    \\u1_ndr_r_reg[5]  <= n3416;
    \\u1_ndr_r_reg[6]  <= n3421;
    \\u1_ndr_r_reg[19]  <= n3426;
    \\u1_ndr_r_reg[21]  <= n3431;
    \\u1_ndr_r_reg[25]  <= n3436;
    \\u1_ndr_r_reg[13]  <= n3441;
    \\u1_ndr_r_reg[3]  <= n3446;
    \\u1_ndr_r_reg[26]  <= n3451;
    \\u1_ndr_r_reg[0]  <= n3456;
    \\u1_ndnr_reg[0]  <= n3461;
    \\u2_u0_out_r_reg[0]  <= n3466;
    \\u2_u1_out_r_reg[0]  <= n3471;
    \\u1_req_r_reg[0]  <= n3476;
    \\u3_u1_slv_adr_reg[3]  <= n3481;
    \\u3_u1_slv_dout_reg[4]  <= n3486;
    \\u3_u1_slv_dout_reg[0]  <= n3491;
    \\u3_u1_slv_dout_reg[18]  <= n3496;
    \\u3_u1_slv_dout_reg[7]  <= n3501;
    \\u3_u1_slv_adr_reg[6]  <= n3506;
    \\u3_u1_slv_dout_reg[5]  <= n3511;
    \\u3_u1_slv_dout_reg[24]  <= n3516;
    \\u3_u1_slv_dout_reg[1]  <= n3521;
    \\u3_u1_slv_adr_reg[8]  <= n3526;
    \\u3_u1_slv_dout_reg[19]  <= n3531;
    \\u3_u1_slv_dout_reg[31]  <= n3536;
    \\u3_u1_slv_dout_reg[6]  <= n3541;
    \\u3_u1_slv_adr_reg[9]  <= n3546;
    \\u3_u1_slv_dout_reg[20]  <= n3551;
    \\u3_u1_slv_adr_reg[4]  <= n3556;
    \\u3_u1_slv_dout_reg[30]  <= n3561;
    \\u3_u1_slv_dout_reg[26]  <= n3566;
    \\u3_u1_slv_dout_reg[29]  <= n3571;
    \\u3_u1_slv_dout_reg[28]  <= n3576;
    \\u3_u1_slv_dout_reg[2]  <= n3581;
    \\u3_u1_slv_dout_reg[8]  <= n3586;
    \\u3_u1_slv_adr_reg[7]  <= n3591;
    \\u3_u1_slv_adr_reg[2]  <= n3596;
    \\u3_u1_slv_dout_reg[14]  <= n3601;
    \\u3_u1_slv_dout_reg[23]  <= n3606;
    \\u3_u1_slv_dout_reg[9]  <= n3611;
    \\u3_u1_slv_dout_reg[21]  <= n3616;
    \\u3_u1_slv_dout_reg[25]  <= n3621;
    \\u3_u1_slv_dout_reg[27]  <= n3626;
    \\u3_u1_slv_dout_reg[3]  <= n3631;
    \\u3_u1_slv_dout_reg[12]  <= n3636;
    \\u3_u1_slv_dout_reg[17]  <= n3641;
    \\u3_u1_slv_adr_reg[5]  <= n3646;
    \\u3_u1_slv_dout_reg[11]  <= n3651;
    \\u3_u1_slv_dout_reg[15]  <= n3656;
    \\u3_u1_slv_dout_reg[13]  <= n3661;
    \\u3_u1_slv_dout_reg[10]  <= n3666;
    \\u3_u1_slv_dout_reg[16]  <= n3671;
    \\u3_u1_slv_dout_reg[22]  <= n3676;
  end
  initial begin
    \\u2_state_reg[1]  <= 1'b0;
    \\u2_state_reg[3]  <= 1'b0;
    \\u0_u0_int_src_r_reg[2]  <= 1'b0;
    \\u0_u0_ch_csr_r_reg[0]  <= 1'b0;
    u0_u0_ch_done_reg <= 1'b0;
    \\u0_u0_int_src_r_reg[1]  <= 1'b0;
    \\u2_state_reg[0]  <= 1'b1;
    \\u2_state_reg[9]  <= 1'b0;
    \\u2_state_reg[10]  <= 1'b0;
    \\u2_state_reg[4]  <= 1'b0;
    \\u2_state_reg[2]  <= 1'b0;
    \\u0_u0_ch_csr_r_reg[4]  <= 1'b0;
    u0_u0_ch_err_reg <= 1'b0;
    \\u0_u0_ch_csr_r_reg[1]  <= 1'b0;
    \\u0_u0_ch_csr_r_reg[2]  <= 1'b0;
    \\u0_u0_ch_csr_r_reg[3]  <= 1'b0;
    \\u0_u0_int_src_r_reg[0]  <= 1'b0;
    \\u1_ch_sel_r_reg[2]  <= 1'b0;
    \\u1_ch_sel_r_reg[1]  <= 1'b0;
    \\u1_ch_sel_r_reg[3]  <= 1'b0;
    \\u1_ch_sel_r_reg[4]  <= 1'b0;
    \\u1_ch_sel_r_reg[0]  <= 1'b0;
    \\u2_state_reg[5]  <= 1'b0;
    \\u0_u0_ch_csr_r3_reg[2]  <= 1'b0;
    \\u0_u0_ch_csr_r3_reg[0]  <= 1'b0;
    u0_u0_rest_en_reg <= 1'b0;
    \\u0_u0_ch_csr_r_reg[7]  <= 1'b0;
    \\u0_u0_ch_csr_r_reg[5]  <= 1'b0;
    \\u0_u0_ch_csr_r2_reg[2]  <= 1'b0;
    \\u0_u0_ch_csr_r2_reg[1]  <= 1'b0;
    \\u0_u0_ch_csr_r2_reg[0]  <= 1'b0;
    \\u0_u0_ch_csr_r3_reg[1]  <= 1'b0;
    \\u0_u0_ch_csr_r_reg[6]  <= 1'b0;
    \\u0_u0_ch_csr_r_reg[8]  <= 1'b0;
    \\u1_u1_state_reg[2]  <= 1'b0;
    \\u1_u1_state_reg[3]  <= 1'b0;
    \\u1_u1_state_reg[4]  <= 1'b0;
    \\u1_u1_state_reg[0]  <= 1'b0;
    \\u1_u1_state_reg[1]  <= 1'b0;
    \\u2_state_reg[8]  <= 1'b0;
    \\u2_state_reg[7]  <= 1'b0;
    \\u2_state_reg[6]  <= 1'b0;
    \\u0_int_maska_r_reg[11]  <= 1'b0;
    \\u0_csr_r_reg[0]  <= 1'b0;
    \\u0_int_maska_r_reg[0]  <= 1'b0;
    \\u0_int_maska_r_reg[10]  <= 1'b0;
    \\u0_int_maska_r_reg[5]  <= 1'b0;
    \\u0_int_maska_r_reg[6]  <= 1'b0;
    \\u0_int_maska_r_reg[7]  <= 1'b0;
    \\u0_int_maska_r_reg[8]  <= 1'b0;
    \\u0_int_maska_r_reg[9]  <= 1'b0;
    \\u0_int_maska_r_reg[2]  <= 1'b0;
    \\u0_int_maska_r_reg[4]  <= 1'b0;
    \\u0_int_maska_r_reg[3]  <= 1'b0;
    \\u0_int_maska_r_reg[29]  <= 1'b0;
    \\u0_int_maska_r_reg[26]  <= 1'b0;
    \\u0_int_maska_r_reg[27]  <= 1'b0;
    \\u0_int_maska_r_reg[28]  <= 1'b0;
    \\u0_int_maska_r_reg[19]  <= 1'b0;
    \\u0_int_maska_r_reg[22]  <= 1'b0;
    \\u0_int_maska_r_reg[24]  <= 1'b0;
    \\u0_int_maska_r_reg[23]  <= 1'b0;
    \\u0_int_maska_r_reg[1]  <= 1'b0;
    \\u0_int_maska_r_reg[20]  <= 1'b0;
    \\u0_int_maska_r_reg[16]  <= 1'b0;
    \\u0_int_maska_r_reg[17]  <= 1'b0;
    \\u0_int_maska_r_reg[15]  <= 1'b0;
    \\u0_int_maska_r_reg[12]  <= 1'b0;
    \\u0_int_maska_r_reg[13]  <= 1'b0;
    \\u0_int_maska_r_reg[14]  <= 1'b0;
    \\u0_int_maskb_r_reg[6]  <= 1'b0;
    \\u0_int_maskb_r_reg[9]  <= 1'b0;
    \\u0_int_maska_r_reg[18]  <= 1'b0;
    \\u0_int_maska_r_reg[21]  <= 1'b0;
    \\u0_int_maska_r_reg[25]  <= 1'b0;
    \\u0_int_maska_r_reg[30]  <= 1'b0;
    \\u0_int_maskb_r_reg[0]  <= 1'b0;
    \\u0_int_maskb_r_reg[7]  <= 1'b0;
    \\u0_int_maskb_r_reg[8]  <= 1'b0;
    \\u0_int_maskb_r_reg[5]  <= 1'b0;
    \\u0_int_maskb_r_reg[11]  <= 1'b0;
    \\u0_int_maskb_r_reg[10]  <= 1'b0;
    \\u0_int_maskb_r_reg[14]  <= 1'b0;
    \\u0_int_maskb_r_reg[17]  <= 1'b0;
    \\u0_int_maskb_r_reg[20]  <= 1'b0;
    \\u0_int_maskb_r_reg[22]  <= 1'b0;
    \\u0_int_maskb_r_reg[2]  <= 1'b0;
    \\u0_int_maskb_r_reg[12]  <= 1'b0;
    \\u0_int_maskb_r_reg[18]  <= 1'b0;
    \\u0_int_maskb_r_reg[19]  <= 1'b0;
    \\u0_int_maskb_r_reg[15]  <= 1'b0;
    \\u0_int_maskb_r_reg[24]  <= 1'b0;
    \\u0_int_maskb_r_reg[30]  <= 1'b0;
    \\u0_int_maskb_r_reg[3]  <= 1'b0;
    \\u0_int_maskb_r_reg[4]  <= 1'b0;
    \\u0_int_maskb_r_reg[25]  <= 1'b0;
    \\u0_int_maskb_r_reg[28]  <= 1'b0;
    \\u0_int_maskb_r_reg[29]  <= 1'b0;
    \\u0_int_maskb_r_reg[26]  <= 1'b0;
    \\u0_int_maskb_r_reg[27]  <= 1'b0;
    \\u0_int_maskb_r_reg[23]  <= 1'b0;
    \\u0_int_maskb_r_reg[1]  <= 1'b0;
    \\u0_int_maskb_r_reg[21]  <= 1'b0;
    \\u0_int_maskb_r_reg[16]  <= 1'b0;
    \\u0_int_maskb_r_reg[13]  <= 1'b0;
  end
endmodule


