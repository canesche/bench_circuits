module top ( 
    i_89_, i_76_, i_63_, i_50_, i_75_, i_64_, i_78_, i_61_, i_99_, i_77_,
    i_62_, i_40_, i_120_, i_72_, i_67_, i_121_, i_71_, i_68_, i_122_,
    i_74_, i_65_, i_30_, i_123_, i_73_, i_66_, i_124_, i_94_, i_81_,
    i_125_, i_93_, i_82_, i_20_, i_126_, i_92_, i_83_, i_69_, i_9_, i_127_,
    i_91_, i_84_, i_128_, i_98_, i_85_, i_10_, i_7_, i_129_, i_97_, i_86_,
    i_79_, i_8_, i_96_, i_87_, i_5_, i_95_, i_88_, i_6_, i_27_, i_14_,
    i_3_, i_39_, i_28_, i_13_, i_4_, i_119_, i_108_, i_25_, i_12_, i_1_,
    i_118_, i_109_, i_26_, i_11_, i_2_, i_117_, i_106_, i_90_, i_49_,
    i_23_, i_18_, i_116_, i_107_, i_24_, i_17_, i_0_, i_115_, i_104_,
    i_21_, i_16_, i_114_, i_105_, i_80_, i_59_, i_22_, i_15_, i_113_,
    i_102_, i_58_, i_45_, i_32_, i_112_, i_103_, i_57_, i_46_, i_31_,
    i_111_, i_100_, i_70_, i_56_, i_47_, i_34_, i_110_, i_101_, i_55_,
    i_48_, i_33_, i_19_, i_54_, i_41_, i_36_, i_60_, i_53_, i_42_, i_35_,
    i_52_, i_43_, i_38_, i_29_, i_51_, i_44_, i_37_,
    o_0_  );
  input  i_89_, i_76_, i_63_, i_50_, i_75_, i_64_, i_78_, i_61_, i_99_,
    i_77_, i_62_, i_40_, i_120_, i_72_, i_67_, i_121_, i_71_, i_68_,
    i_122_, i_74_, i_65_, i_30_, i_123_, i_73_, i_66_, i_124_, i_94_,
    i_81_, i_125_, i_93_, i_82_, i_20_, i_126_, i_92_, i_83_, i_69_, i_9_,
    i_127_, i_91_, i_84_, i_128_, i_98_, i_85_, i_10_, i_7_, i_129_, i_97_,
    i_86_, i_79_, i_8_, i_96_, i_87_, i_5_, i_95_, i_88_, i_6_, i_27_,
    i_14_, i_3_, i_39_, i_28_, i_13_, i_4_, i_119_, i_108_, i_25_, i_12_,
    i_1_, i_118_, i_109_, i_26_, i_11_, i_2_, i_117_, i_106_, i_90_, i_49_,
    i_23_, i_18_, i_116_, i_107_, i_24_, i_17_, i_0_, i_115_, i_104_,
    i_21_, i_16_, i_114_, i_105_, i_80_, i_59_, i_22_, i_15_, i_113_,
    i_102_, i_58_, i_45_, i_32_, i_112_, i_103_, i_57_, i_46_, i_31_,
    i_111_, i_100_, i_70_, i_56_, i_47_, i_34_, i_110_, i_101_, i_55_,
    i_48_, i_33_, i_19_, i_54_, i_41_, i_36_, i_60_, i_53_, i_42_, i_35_,
    i_52_, i_43_, i_38_, i_29_, i_51_, i_44_, i_37_;
  output o_0_;
  wire new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_;
  assign new_n132_ = i_105_ & i_41_;
  assign new_n133_ = i_106_ & i_42_;
  assign new_n134_ = i_40_ & i_104_;
  assign new_n135_ = ~new_n132_ & ~new_n133_;
  assign new_n136_ = ~new_n134_ & new_n135_;
  assign new_n137_ = i_108_ & i_44_;
  assign new_n138_ = i_109_ & i_45_;
  assign new_n139_ = i_107_ & i_43_;
  assign new_n140_ = ~new_n137_ & ~new_n138_;
  assign new_n141_ = ~new_n139_ & new_n140_;
  assign new_n142_ = i_102_ & i_38_;
  assign new_n143_ = i_39_ & i_103_;
  assign new_n144_ = i_101_ & i_37_;
  assign new_n145_ = ~new_n142_ & ~new_n143_;
  assign new_n146_ = ~new_n144_ & new_n145_;
  assign new_n147_ = new_n136_ & new_n141_;
  assign new_n148_ = new_n146_ & new_n147_;
  assign new_n149_ = i_50_ & i_114_;
  assign new_n150_ = i_115_ & i_51_;
  assign new_n151_ = i_49_ & i_113_;
  assign new_n152_ = ~new_n149_ & ~new_n150_;
  assign new_n153_ = ~new_n151_ & new_n152_;
  assign new_n154_ = i_117_ & i_53_;
  assign new_n155_ = i_118_ & i_54_;
  assign new_n156_ = i_116_ & i_52_;
  assign new_n157_ = ~new_n154_ & ~new_n155_;
  assign new_n158_ = ~new_n156_ & new_n157_;
  assign new_n159_ = i_111_ & i_47_;
  assign new_n160_ = i_112_ & i_48_;
  assign new_n161_ = i_46_ & i_110_;
  assign new_n162_ = ~new_n159_ & ~new_n160_;
  assign new_n163_ = ~new_n161_ & new_n162_;
  assign new_n164_ = new_n153_ & new_n158_;
  assign new_n165_ = new_n163_ & new_n164_;
  assign new_n166_ = i_96_ & i_32_;
  assign new_n167_ = i_97_ & i_33_;
  assign new_n168_ = i_95_ & i_31_;
  assign new_n169_ = ~new_n166_ & ~new_n167_;
  assign new_n170_ = ~new_n168_ & new_n169_;
  assign new_n171_ = i_99_ & i_35_;
  assign new_n172_ = i_100_ & i_36_;
  assign new_n173_ = i_98_ & i_34_;
  assign new_n174_ = ~new_n171_ & ~new_n172_;
  assign new_n175_ = ~new_n173_ & new_n174_;
  assign new_n176_ = i_93_ & i_29_;
  assign new_n177_ = i_30_ & i_94_;
  assign new_n178_ = i_92_ & i_28_;
  assign new_n179_ = ~new_n176_ & ~new_n177_;
  assign new_n180_ = ~new_n178_ & new_n179_;
  assign new_n181_ = new_n170_ & new_n175_;
  assign new_n182_ = new_n180_ & new_n181_;
  assign new_n183_ = new_n148_ & new_n165_;
  assign new_n184_ = new_n182_ & new_n183_;
  assign new_n185_ = i_129_ & i_0_;
  assign new_n186_ = i_64_ & i_128_;
  assign new_n187_ = ~new_n185_ & ~new_n186_;
  assign new_n188_ = i_123_ & i_59_;
  assign new_n189_ = i_124_ & i_60_;
  assign new_n190_ = i_122_ & i_58_;
  assign new_n191_ = ~new_n188_ & ~new_n189_;
  assign new_n192_ = ~new_n190_ & new_n191_;
  assign new_n193_ = i_62_ & i_126_;
  assign new_n194_ = i_63_ & i_127_;
  assign new_n195_ = i_61_ & i_125_;
  assign new_n196_ = ~new_n193_ & ~new_n194_;
  assign new_n197_ = ~new_n195_ & new_n196_;
  assign new_n198_ = i_120_ & i_56_;
  assign new_n199_ = i_121_ & i_57_;
  assign new_n200_ = i_119_ & i_55_;
  assign new_n201_ = ~new_n198_ & ~new_n199_;
  assign new_n202_ = ~new_n200_ & new_n201_;
  assign new_n203_ = new_n192_ & new_n197_;
  assign new_n204_ = new_n202_ & new_n203_;
  assign new_n205_ = new_n187_ & new_n204_;
  assign new_n206_ = i_78_ & i_14_;
  assign new_n207_ = i_79_ & i_15_;
  assign new_n208_ = i_77_ & i_13_;
  assign new_n209_ = ~new_n206_ & ~new_n207_;
  assign new_n210_ = ~new_n208_ & new_n209_;
  assign new_n211_ = i_81_ & i_17_;
  assign new_n212_ = i_82_ & i_18_;
  assign new_n213_ = i_16_ & i_80_;
  assign new_n214_ = ~new_n211_ & ~new_n212_;
  assign new_n215_ = ~new_n213_ & new_n214_;
  assign new_n216_ = i_75_ & i_11_;
  assign new_n217_ = i_76_ & i_12_;
  assign new_n218_ = i_74_ & i_10_;
  assign new_n219_ = ~new_n216_ & ~new_n217_;
  assign new_n220_ = ~new_n218_ & new_n219_;
  assign new_n221_ = new_n210_ & new_n215_;
  assign new_n222_ = new_n220_ & new_n221_;
  assign new_n223_ = i_87_ & i_23_;
  assign new_n224_ = i_88_ & i_24_;
  assign new_n225_ = i_86_ & i_22_;
  assign new_n226_ = ~new_n223_ & ~new_n224_;
  assign new_n227_ = ~new_n225_ & new_n226_;
  assign new_n228_ = i_26_ & i_90_;
  assign new_n229_ = i_91_ & i_27_;
  assign new_n230_ = i_89_ & i_25_;
  assign new_n231_ = ~new_n228_ & ~new_n229_;
  assign new_n232_ = ~new_n230_ & new_n231_;
  assign new_n233_ = i_20_ & i_84_;
  assign new_n234_ = i_85_ & i_21_;
  assign new_n235_ = i_83_ & i_19_;
  assign new_n236_ = ~new_n233_ & ~new_n234_;
  assign new_n237_ = ~new_n235_ & new_n236_;
  assign new_n238_ = new_n227_ & new_n232_;
  assign new_n239_ = new_n237_ & new_n238_;
  assign new_n240_ = i_69_ & i_5_;
  assign new_n241_ = i_6_ & i_70_;
  assign new_n242_ = i_68_ & i_4_;
  assign new_n243_ = ~new_n240_ & ~new_n241_;
  assign new_n244_ = ~new_n242_ & new_n243_;
  assign new_n245_ = i_72_ & i_8_;
  assign new_n246_ = i_73_ & i_9_;
  assign new_n247_ = i_71_ & i_7_;
  assign new_n248_ = ~new_n245_ & ~new_n246_;
  assign new_n249_ = ~new_n247_ & new_n248_;
  assign new_n250_ = i_66_ & i_2_;
  assign new_n251_ = i_67_ & i_3_;
  assign new_n252_ = i_65_ & i_1_;
  assign new_n253_ = ~new_n250_ & ~new_n251_;
  assign new_n254_ = ~new_n252_ & new_n253_;
  assign new_n255_ = new_n244_ & new_n249_;
  assign new_n256_ = new_n254_ & new_n255_;
  assign new_n257_ = new_n222_ & new_n239_;
  assign new_n258_ = new_n256_ & new_n257_;
  assign new_n259_ = new_n184_ & new_n205_;
  assign o_0_ = ~new_n258_ | ~new_n259_;
endmodule

