module Min_Max9_4 ( clock, 
    \1 , 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12,
    40, 41, 42, 43, 44, 45, 46, 47, 48  );
  input  clock;
  input  \1 , 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12;
  output 40, 41, 42, 43, 44, 45, 46, 47, 48;
  reg 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29,
    30, 31, 32, 33, 34, 35, 36, 37, 38, 39;
  wire new_n103_, new_n104_1_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_1_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_1_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_1_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_1_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_1_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_1_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_1_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_1_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_1_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_1_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_1_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_1_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_1_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_1_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n435_,
    new_n436_, new_n438_, new_n439_, new_n441_, new_n442_, new_n444_,
    new_n445_, new_n447_, new_n448_, new_n450_, new_n451_, new_n453_,
    new_n454_, new_n456_, new_n457_, new_n459_, new_n460_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n516_, new_n517_, new_n519_, new_n520_,
    new_n522_, new_n523_, new_n525_, new_n526_, new_n528_, new_n529_,
    new_n531_, new_n532_, new_n534_, new_n535_, new_n537_, new_n538_,
    new_n540_, new_n541_, n44, n49, n54, n59, n64, n69, n74, n79, n84, n89,
    n94, n99, n104, n109, n114, n119, n124, n129, n134, n139, n144, n149,
    n154, n159, n164, n169, n174;
  assign new_n103_ = 12 & ~39;
  assign new_n104_1_ = ~12 & 39;
  assign new_n105_ = ~new_n103_ & ~new_n104_1_;
  assign new_n106_ = 11 & ~38;
  assign new_n107_ = ~11 & 38;
  assign new_n108_ = ~new_n106_ & ~new_n107_;
  assign new_n109_1_ = 10 & ~37;
  assign new_n110_ = ~10 & 37;
  assign new_n111_ = ~new_n109_1_ & ~new_n110_;
  assign new_n112_ = 9 & ~36;
  assign new_n113_ = ~9 & 36;
  assign new_n114_1_ = ~new_n112_ & ~new_n113_;
  assign new_n115_ = 8 & ~35;
  assign new_n116_ = ~8 & 35;
  assign new_n117_ = ~new_n115_ & ~new_n116_;
  assign new_n118_ = 7 & ~34;
  assign new_n119_1_ = ~7 & 34;
  assign new_n120_ = ~new_n118_ & ~new_n119_1_;
  assign new_n121_ = 6 & ~33;
  assign new_n122_ = ~6 & 33;
  assign new_n123_ = ~new_n121_ & ~new_n122_;
  assign new_n124_1_ = 5 & ~32;
  assign new_n125_ = ~5 & 32;
  assign new_n126_ = ~new_n124_1_ & ~new_n125_;
  assign new_n127_ = 4 & ~31;
  assign new_n128_ = ~4 & 31;
  assign new_n129_1_ = ~new_n127_ & ~new_n128_;
  assign new_n130_ = 4 & ~new_n129_1_;
  assign new_n131_ = new_n126_ & new_n130_;
  assign new_n132_ = 5 & ~new_n126_;
  assign new_n133_ = ~new_n131_ & ~new_n132_;
  assign new_n134_1_ = new_n123_ & ~new_n133_;
  assign new_n135_ = 6 & ~new_n123_;
  assign new_n136_ = ~new_n134_1_ & ~new_n135_;
  assign new_n137_ = new_n120_ & ~new_n136_;
  assign new_n138_ = 7 & ~new_n120_;
  assign new_n139_1_ = ~new_n137_ & ~new_n138_;
  assign new_n140_ = new_n117_ & ~new_n139_1_;
  assign new_n141_ = 8 & ~new_n117_;
  assign new_n142_ = ~new_n140_ & ~new_n141_;
  assign new_n143_ = new_n114_1_ & ~new_n142_;
  assign new_n144_1_ = 9 & ~new_n114_1_;
  assign new_n145_ = ~new_n143_ & ~new_n144_1_;
  assign new_n146_ = new_n111_ & ~new_n145_;
  assign new_n147_ = 10 & ~new_n111_;
  assign new_n148_ = ~new_n146_ & ~new_n147_;
  assign new_n149_1_ = new_n108_ & ~new_n148_;
  assign new_n150_ = 11 & ~new_n108_;
  assign new_n151_ = ~new_n149_1_ & ~new_n150_;
  assign new_n152_ = new_n105_ & ~new_n151_;
  assign new_n153_ = 12 & ~new_n105_;
  assign new_n154_1_ = ~new_n152_ & ~new_n153_;
  assign new_n155_ = 2 & ~3;
  assign new_n156_ = ~\1  & new_n155_;
  assign new_n157_ = ~new_n154_1_ & new_n156_;
  assign new_n158_ = 31 & ~new_n157_;
  assign new_n159_1_ = 4 & new_n157_;
  assign new_n160_ = ~new_n158_ & ~new_n159_1_;
  assign new_n161_ = new_n156_ & ~new_n160_;
  assign new_n162_ = 12 & ~30;
  assign new_n163_ = ~12 & 30;
  assign new_n164_1_ = ~new_n162_ & ~new_n163_;
  assign new_n165_ = 11 & ~29;
  assign new_n166_ = ~11 & 29;
  assign new_n167_ = ~new_n165_ & ~new_n166_;
  assign new_n168_ = 10 & ~28;
  assign new_n169_1_ = ~10 & 28;
  assign new_n170_ = ~new_n168_ & ~new_n169_1_;
  assign new_n171_ = 9 & ~27;
  assign new_n172_ = ~9 & 27;
  assign new_n173_ = ~new_n171_ & ~new_n172_;
  assign new_n174_1_ = 8 & ~26;
  assign new_n175_ = ~8 & 26;
  assign new_n176_ = ~new_n174_1_ & ~new_n175_;
  assign new_n177_ = 7 & ~25;
  assign new_n178_ = ~7 & 25;
  assign new_n179_ = ~new_n177_ & ~new_n178_;
  assign new_n180_ = 6 & ~24;
  assign new_n181_ = ~6 & 24;
  assign new_n182_ = ~new_n180_ & ~new_n181_;
  assign new_n183_ = 5 & ~23;
  assign new_n184_ = ~5 & 23;
  assign new_n185_ = ~new_n183_ & ~new_n184_;
  assign new_n186_ = 4 & ~22;
  assign new_n187_ = ~4 & 22;
  assign new_n188_ = ~new_n186_ & ~new_n187_;
  assign new_n189_ = 4 & ~new_n188_;
  assign new_n190_ = new_n185_ & new_n189_;
  assign new_n191_ = 5 & ~new_n185_;
  assign new_n192_ = ~new_n190_ & ~new_n191_;
  assign new_n193_ = new_n182_ & ~new_n192_;
  assign new_n194_ = 6 & ~new_n182_;
  assign new_n195_ = ~new_n193_ & ~new_n194_;
  assign new_n196_ = new_n179_ & ~new_n195_;
  assign new_n197_ = 7 & ~new_n179_;
  assign new_n198_ = ~new_n196_ & ~new_n197_;
  assign new_n199_ = new_n176_ & ~new_n198_;
  assign new_n200_ = 8 & ~new_n176_;
  assign new_n201_ = ~new_n199_ & ~new_n200_;
  assign new_n202_ = new_n173_ & ~new_n201_;
  assign new_n203_ = 9 & ~new_n173_;
  assign new_n204_ = ~new_n202_ & ~new_n203_;
  assign new_n205_ = new_n170_ & ~new_n204_;
  assign new_n206_ = 10 & ~new_n170_;
  assign new_n207_ = ~new_n205_ & ~new_n206_;
  assign new_n208_ = new_n167_ & ~new_n207_;
  assign new_n209_ = 11 & ~new_n167_;
  assign new_n210_ = ~new_n208_ & ~new_n209_;
  assign new_n211_ = new_n164_1_ & ~new_n210_;
  assign new_n212_ = 12 & ~new_n164_1_;
  assign new_n213_ = ~new_n211_ & ~new_n212_;
  assign new_n214_ = new_n156_ & ~new_n213_;
  assign new_n215_ = 22 & new_n214_;
  assign new_n216_ = 4 & ~new_n214_;
  assign new_n217_ = ~new_n215_ & ~new_n216_;
  assign new_n218_ = new_n156_ & ~new_n217_;
  assign new_n219_ = new_n161_ & new_n218_;
  assign new_n220_ = 32 & ~new_n157_;
  assign new_n221_ = 5 & new_n157_;
  assign new_n222_ = ~new_n220_ & ~new_n221_;
  assign new_n223_ = new_n156_ & ~new_n222_;
  assign new_n224_ = 23 & new_n214_;
  assign new_n225_ = 5 & ~new_n214_;
  assign new_n226_ = ~new_n224_ & ~new_n225_;
  assign new_n227_ = new_n156_ & ~new_n226_;
  assign new_n228_ = ~new_n223_ & ~new_n227_;
  assign new_n229_ = new_n223_ & new_n227_;
  assign new_n230_ = ~new_n228_ & ~new_n229_;
  assign new_n231_ = new_n219_ & ~new_n230_;
  assign new_n232_ = ~new_n223_ & new_n227_;
  assign new_n233_ = new_n223_ & ~new_n227_;
  assign new_n234_ = ~new_n232_ & ~new_n233_;
  assign new_n235_ = ~new_n219_ & ~new_n234_;
  assign new_n236_ = ~new_n231_ & ~new_n235_;
  assign new_n237_ = ~3 & ~new_n236_;
  assign new_n238_ = 3 & 4;
  assign new_n239_ = ~new_n237_ & ~new_n238_;
  assign new_n240_ = 2 & ~new_n239_;
  assign new_n241_ = ~2 & 13;
  assign new_n242_ = ~new_n240_ & ~new_n241_;
  assign 40 = ~\1  & ~new_n242_;
  assign new_n244_ = new_n219_ & ~new_n228_;
  assign new_n245_ = ~new_n229_ & ~new_n244_;
  assign new_n246_ = 33 & ~new_n157_;
  assign new_n247_ = 6 & new_n157_;
  assign new_n248_ = ~new_n246_ & ~new_n247_;
  assign new_n249_ = new_n156_ & ~new_n248_;
  assign new_n250_ = 24 & new_n214_;
  assign new_n251_ = 6 & ~new_n214_;
  assign new_n252_ = ~new_n250_ & ~new_n251_;
  assign new_n253_ = new_n156_ & ~new_n252_;
  assign new_n254_ = ~new_n249_ & ~new_n253_;
  assign new_n255_ = new_n249_ & new_n253_;
  assign new_n256_ = ~new_n254_ & ~new_n255_;
  assign new_n257_ = ~new_n245_ & ~new_n256_;
  assign new_n258_ = ~new_n249_ & new_n253_;
  assign new_n259_ = new_n249_ & ~new_n253_;
  assign new_n260_ = ~new_n258_ & ~new_n259_;
  assign new_n261_ = new_n245_ & ~new_n260_;
  assign new_n262_ = ~new_n257_ & ~new_n261_;
  assign new_n263_ = ~3 & ~new_n262_;
  assign new_n264_ = 3 & 5;
  assign new_n265_ = ~new_n263_ & ~new_n264_;
  assign new_n266_ = 2 & ~new_n265_;
  assign new_n267_ = ~2 & 14;
  assign new_n268_ = ~new_n266_ & ~new_n267_;
  assign 41 = ~\1  & ~new_n268_;
  assign new_n270_ = ~new_n245_ & ~new_n254_;
  assign new_n271_ = ~new_n255_ & ~new_n270_;
  assign new_n272_ = 34 & ~new_n157_;
  assign new_n273_ = 7 & new_n157_;
  assign new_n274_ = ~new_n272_ & ~new_n273_;
  assign new_n275_ = new_n156_ & ~new_n274_;
  assign new_n276_ = 25 & new_n214_;
  assign new_n277_ = 7 & ~new_n214_;
  assign new_n278_ = ~new_n276_ & ~new_n277_;
  assign new_n279_ = new_n156_ & ~new_n278_;
  assign new_n280_ = ~new_n275_ & ~new_n279_;
  assign new_n281_ = new_n275_ & new_n279_;
  assign new_n282_ = ~new_n280_ & ~new_n281_;
  assign new_n283_ = ~new_n271_ & ~new_n282_;
  assign new_n284_ = ~new_n275_ & new_n279_;
  assign new_n285_ = new_n275_ & ~new_n279_;
  assign new_n286_ = ~new_n284_ & ~new_n285_;
  assign new_n287_ = new_n271_ & ~new_n286_;
  assign new_n288_ = ~new_n283_ & ~new_n287_;
  assign new_n289_ = ~3 & ~new_n288_;
  assign new_n290_ = 3 & 6;
  assign new_n291_ = ~new_n289_ & ~new_n290_;
  assign new_n292_ = 2 & ~new_n291_;
  assign new_n293_ = ~2 & 15;
  assign new_n294_ = ~new_n292_ & ~new_n293_;
  assign 42 = ~\1  & ~new_n294_;
  assign new_n296_ = ~new_n271_ & ~new_n280_;
  assign new_n297_ = ~new_n281_ & ~new_n296_;
  assign new_n298_ = 35 & ~new_n157_;
  assign new_n299_ = 8 & new_n157_;
  assign new_n300_ = ~new_n298_ & ~new_n299_;
  assign new_n301_ = new_n156_ & ~new_n300_;
  assign new_n302_ = 26 & new_n214_;
  assign new_n303_ = 8 & ~new_n214_;
  assign new_n304_ = ~new_n302_ & ~new_n303_;
  assign new_n305_ = new_n156_ & ~new_n304_;
  assign new_n306_ = ~new_n301_ & ~new_n305_;
  assign new_n307_ = new_n301_ & new_n305_;
  assign new_n308_ = ~new_n306_ & ~new_n307_;
  assign new_n309_ = ~new_n297_ & ~new_n308_;
  assign new_n310_ = ~new_n301_ & new_n305_;
  assign new_n311_ = new_n301_ & ~new_n305_;
  assign new_n312_ = ~new_n310_ & ~new_n311_;
  assign new_n313_ = new_n297_ & ~new_n312_;
  assign new_n314_ = ~new_n309_ & ~new_n313_;
  assign new_n315_ = ~3 & ~new_n314_;
  assign new_n316_ = 3 & 7;
  assign new_n317_ = ~new_n315_ & ~new_n316_;
  assign new_n318_ = 2 & ~new_n317_;
  assign new_n319_ = ~2 & 16;
  assign new_n320_ = ~new_n318_ & ~new_n319_;
  assign 43 = ~\1  & ~new_n320_;
  assign new_n322_ = ~new_n297_ & ~new_n306_;
  assign new_n323_ = ~new_n307_ & ~new_n322_;
  assign new_n324_ = 36 & ~new_n157_;
  assign new_n325_ = 9 & new_n157_;
  assign new_n326_ = ~new_n324_ & ~new_n325_;
  assign new_n327_ = new_n156_ & ~new_n326_;
  assign new_n328_ = 27 & new_n214_;
  assign new_n329_ = 9 & ~new_n214_;
  assign new_n330_ = ~new_n328_ & ~new_n329_;
  assign new_n331_ = new_n156_ & ~new_n330_;
  assign new_n332_ = ~new_n327_ & ~new_n331_;
  assign new_n333_ = new_n327_ & new_n331_;
  assign new_n334_ = ~new_n332_ & ~new_n333_;
  assign new_n335_ = ~new_n323_ & ~new_n334_;
  assign new_n336_ = ~new_n327_ & new_n331_;
  assign new_n337_ = new_n327_ & ~new_n331_;
  assign new_n338_ = ~new_n336_ & ~new_n337_;
  assign new_n339_ = new_n323_ & ~new_n338_;
  assign new_n340_ = ~new_n335_ & ~new_n339_;
  assign new_n341_ = ~3 & ~new_n340_;
  assign new_n342_ = 3 & 8;
  assign new_n343_ = ~new_n341_ & ~new_n342_;
  assign new_n344_ = 2 & ~new_n343_;
  assign new_n345_ = ~2 & 17;
  assign new_n346_ = ~new_n344_ & ~new_n345_;
  assign 44 = ~\1  & ~new_n346_;
  assign new_n348_ = ~new_n323_ & ~new_n332_;
  assign new_n349_ = ~new_n333_ & ~new_n348_;
  assign new_n350_ = 37 & ~new_n157_;
  assign new_n351_ = 10 & new_n157_;
  assign new_n352_ = ~new_n350_ & ~new_n351_;
  assign new_n353_ = new_n156_ & ~new_n352_;
  assign new_n354_ = 28 & new_n214_;
  assign new_n355_ = 10 & ~new_n214_;
  assign new_n356_ = ~new_n354_ & ~new_n355_;
  assign new_n357_ = new_n156_ & ~new_n356_;
  assign new_n358_ = ~new_n353_ & ~new_n357_;
  assign new_n359_ = new_n353_ & new_n357_;
  assign new_n360_ = ~new_n358_ & ~new_n359_;
  assign new_n361_ = ~new_n349_ & ~new_n360_;
  assign new_n362_ = ~new_n353_ & new_n357_;
  assign new_n363_ = new_n353_ & ~new_n357_;
  assign new_n364_ = ~new_n362_ & ~new_n363_;
  assign new_n365_ = new_n349_ & ~new_n364_;
  assign new_n366_ = ~new_n361_ & ~new_n365_;
  assign new_n367_ = ~3 & ~new_n366_;
  assign new_n368_ = 3 & 9;
  assign new_n369_ = ~new_n367_ & ~new_n368_;
  assign new_n370_ = 2 & ~new_n369_;
  assign new_n371_ = ~2 & 18;
  assign new_n372_ = ~new_n370_ & ~new_n371_;
  assign 45 = ~\1  & ~new_n372_;
  assign new_n374_ = ~new_n349_ & ~new_n358_;
  assign new_n375_ = ~new_n359_ & ~new_n374_;
  assign new_n376_ = 38 & ~new_n157_;
  assign new_n377_ = 11 & new_n157_;
  assign new_n378_ = ~new_n376_ & ~new_n377_;
  assign new_n379_ = new_n156_ & ~new_n378_;
  assign new_n380_ = 29 & new_n214_;
  assign new_n381_ = 11 & ~new_n214_;
  assign new_n382_ = ~new_n380_ & ~new_n381_;
  assign new_n383_ = new_n156_ & ~new_n382_;
  assign new_n384_ = ~new_n379_ & ~new_n383_;
  assign new_n385_ = new_n379_ & new_n383_;
  assign new_n386_ = ~new_n384_ & ~new_n385_;
  assign new_n387_ = ~new_n375_ & ~new_n386_;
  assign new_n388_ = ~new_n379_ & new_n383_;
  assign new_n389_ = new_n379_ & ~new_n383_;
  assign new_n390_ = ~new_n388_ & ~new_n389_;
  assign new_n391_ = new_n375_ & ~new_n390_;
  assign new_n392_ = ~new_n387_ & ~new_n391_;
  assign new_n393_ = ~3 & ~new_n392_;
  assign new_n394_ = 3 & 10;
  assign new_n395_ = ~new_n393_ & ~new_n394_;
  assign new_n396_ = 2 & ~new_n395_;
  assign new_n397_ = ~2 & 19;
  assign new_n398_ = ~new_n396_ & ~new_n397_;
  assign 46 = ~\1  & ~new_n398_;
  assign new_n400_ = ~new_n375_ & ~new_n384_;
  assign new_n401_ = ~new_n385_ & ~new_n400_;
  assign new_n402_ = 39 & ~new_n157_;
  assign new_n403_ = 12 & new_n157_;
  assign new_n404_ = ~new_n402_ & ~new_n403_;
  assign new_n405_ = new_n156_ & ~new_n404_;
  assign new_n406_ = 30 & new_n214_;
  assign new_n407_ = 12 & ~new_n214_;
  assign new_n408_ = ~new_n406_ & ~new_n407_;
  assign new_n409_ = new_n156_ & ~new_n408_;
  assign new_n410_ = ~new_n405_ & ~new_n409_;
  assign new_n411_ = new_n405_ & new_n409_;
  assign new_n412_ = ~new_n410_ & ~new_n411_;
  assign new_n413_ = ~new_n401_ & ~new_n412_;
  assign new_n414_ = ~new_n405_ & new_n409_;
  assign new_n415_ = new_n405_ & ~new_n409_;
  assign new_n416_ = ~new_n414_ & ~new_n415_;
  assign new_n417_ = new_n401_ & ~new_n416_;
  assign new_n418_ = ~new_n413_ & ~new_n417_;
  assign new_n419_ = ~3 & ~new_n418_;
  assign new_n420_ = 3 & 11;
  assign new_n421_ = ~new_n419_ & ~new_n420_;
  assign new_n422_ = 2 & ~new_n421_;
  assign new_n423_ = ~2 & 20;
  assign new_n424_ = ~new_n422_ & ~new_n423_;
  assign 47 = ~\1  & ~new_n424_;
  assign new_n426_ = ~new_n401_ & ~new_n410_;
  assign new_n427_ = ~new_n411_ & ~new_n426_;
  assign new_n428_ = ~3 & ~new_n427_;
  assign new_n429_ = 3 & 12;
  assign new_n430_ = ~new_n428_ & ~new_n429_;
  assign new_n431_ = 2 & ~new_n430_;
  assign new_n432_ = ~2 & 21;
  assign new_n433_ = ~new_n431_ & ~new_n432_;
  assign 48 = ~\1  & ~new_n433_;
  assign new_n435_ = 2 & 4;
  assign new_n436_ = ~new_n241_ & ~new_n435_;
  assign n44 = ~\1  & ~new_n436_;
  assign new_n438_ = 2 & 5;
  assign new_n439_ = ~new_n267_ & ~new_n438_;
  assign n49 = ~\1  & ~new_n439_;
  assign new_n441_ = 2 & 6;
  assign new_n442_ = ~new_n293_ & ~new_n441_;
  assign n54 = ~\1  & ~new_n442_;
  assign new_n444_ = 2 & 7;
  assign new_n445_ = ~new_n319_ & ~new_n444_;
  assign n59 = ~\1  & ~new_n445_;
  assign new_n447_ = 2 & 8;
  assign new_n448_ = ~new_n345_ & ~new_n447_;
  assign n64 = ~\1  & ~new_n448_;
  assign new_n450_ = 2 & 9;
  assign new_n451_ = ~new_n371_ & ~new_n450_;
  assign n69 = ~\1  & ~new_n451_;
  assign new_n453_ = 2 & 10;
  assign new_n454_ = ~new_n397_ & ~new_n453_;
  assign n74 = ~\1  & ~new_n454_;
  assign new_n456_ = 2 & 11;
  assign new_n457_ = ~new_n423_ & ~new_n456_;
  assign n79 = ~\1  & ~new_n457_;
  assign new_n459_ = 2 & 12;
  assign new_n460_ = ~new_n432_ & ~new_n459_;
  assign n84 = ~\1  & ~new_n460_;
  assign new_n462_ = ~3 & new_n218_;
  assign new_n463_ = ~3 & ~new_n462_;
  assign new_n464_ = 2 & ~new_n463_;
  assign new_n465_ = 2 & ~new_n464_;
  assign new_n466_ = ~\1  & ~new_n465_;
  assign n89 = \1  | new_n466_;
  assign new_n468_ = ~3 & new_n227_;
  assign new_n469_ = ~3 & ~new_n468_;
  assign new_n470_ = 2 & ~new_n469_;
  assign new_n471_ = 2 & ~new_n470_;
  assign new_n472_ = ~\1  & ~new_n471_;
  assign n94 = \1  | new_n472_;
  assign new_n474_ = ~3 & new_n253_;
  assign new_n475_ = ~3 & ~new_n474_;
  assign new_n476_ = 2 & ~new_n475_;
  assign new_n477_ = 2 & ~new_n476_;
  assign new_n478_ = ~\1  & ~new_n477_;
  assign n99 = \1  | new_n478_;
  assign new_n480_ = ~3 & new_n279_;
  assign new_n481_ = ~3 & ~new_n480_;
  assign new_n482_ = 2 & ~new_n481_;
  assign new_n483_ = 2 & ~new_n482_;
  assign new_n484_ = ~\1  & ~new_n483_;
  assign n104 = \1  | new_n484_;
  assign new_n486_ = ~3 & new_n305_;
  assign new_n487_ = ~3 & ~new_n486_;
  assign new_n488_ = 2 & ~new_n487_;
  assign new_n489_ = 2 & ~new_n488_;
  assign new_n490_ = ~\1  & ~new_n489_;
  assign n109 = \1  | new_n490_;
  assign new_n492_ = ~3 & new_n331_;
  assign new_n493_ = ~3 & ~new_n492_;
  assign new_n494_ = 2 & ~new_n493_;
  assign new_n495_ = 2 & ~new_n494_;
  assign new_n496_ = ~\1  & ~new_n495_;
  assign n114 = \1  | new_n496_;
  assign new_n498_ = ~3 & new_n357_;
  assign new_n499_ = ~3 & ~new_n498_;
  assign new_n500_ = 2 & ~new_n499_;
  assign new_n501_ = 2 & ~new_n500_;
  assign new_n502_ = ~\1  & ~new_n501_;
  assign n119 = \1  | new_n502_;
  assign new_n504_ = ~3 & new_n383_;
  assign new_n505_ = ~3 & ~new_n504_;
  assign new_n506_ = 2 & ~new_n505_;
  assign new_n507_ = 2 & ~new_n506_;
  assign new_n508_ = ~\1  & ~new_n507_;
  assign n124 = \1  | new_n508_;
  assign new_n510_ = ~3 & new_n409_;
  assign new_n511_ = ~3 & ~new_n510_;
  assign new_n512_ = 2 & ~new_n511_;
  assign new_n513_ = 2 & ~new_n512_;
  assign new_n514_ = ~\1  & ~new_n513_;
  assign n129 = \1  | new_n514_;
  assign new_n516_ = ~3 & new_n161_;
  assign new_n517_ = 2 & new_n516_;
  assign n134 = ~\1  & new_n517_;
  assign new_n519_ = ~3 & new_n223_;
  assign new_n520_ = 2 & new_n519_;
  assign n139 = ~\1  & new_n520_;
  assign new_n522_ = ~3 & new_n249_;
  assign new_n523_ = 2 & new_n522_;
  assign n144 = ~\1  & new_n523_;
  assign new_n525_ = ~3 & new_n275_;
  assign new_n526_ = 2 & new_n525_;
  assign n149 = ~\1  & new_n526_;
  assign new_n528_ = ~3 & new_n301_;
  assign new_n529_ = 2 & new_n528_;
  assign n154 = ~\1  & new_n529_;
  assign new_n531_ = ~3 & new_n327_;
  assign new_n532_ = 2 & new_n531_;
  assign n159 = ~\1  & new_n532_;
  assign new_n534_ = ~3 & new_n353_;
  assign new_n535_ = 2 & new_n534_;
  assign n164 = ~\1  & new_n535_;
  assign new_n537_ = ~3 & new_n379_;
  assign new_n538_ = 2 & new_n537_;
  assign n169 = ~\1  & new_n538_;
  assign new_n540_ = ~3 & new_n405_;
  assign new_n541_ = 2 & new_n540_;
  assign n174 = ~\1  & new_n541_;
  always @ (posedge clock) begin
    13 <= n44;
    14 <= n49;
    15 <= n54;
    16 <= n59;
    17 <= n64;
    18 <= n69;
    19 <= n74;
    20 <= n79;
    21 <= n84;
    22 <= n89;
    23 <= n94;
    24 <= n99;
    25 <= n104;
    26 <= n109;
    27 <= n114;
    28 <= n119;
    29 <= n124;
    30 <= n129;
    31 <= n134;
    32 <= n139;
    33 <= n144;
    34 <= n149;
    35 <= n154;
    36 <= n159;
    37 <= n164;
    38 <= n169;
    39 <= n174;
  end
  initial begin
    22 <= 1'b1;
    23 <= 1'b1;
    24 <= 1'b1;
    25 <= 1'b1;
    26 <= 1'b1;
    27 <= 1'b1;
    28 <= 1'b1;
    29 <= 1'b1;
    30 <= 1'b1;
    31 <= 1'b0;
    32 <= 1'b0;
    33 <= 1'b0;
    34 <= 1'b0;
    35 <= 1'b0;
    36 <= 1'b0;
    37 <= 1'b0;
    38 <= 1'b0;
    39 <= 1'b0;
  end
endmodule

