module top ( clock, 
    pg1943, pg1249, pg3219, pg3229, pg3217, pg3228, pg3218, pg3227, pg2637,
    pg3222, pg3233, pg3212, pg3221, pg3234, pclk, pg3220, pg3215, pg3226,
    pg3216, pg3225, pg3230, pg3213, pg3224, pg3231, pg3214, pg3223, pg3232,
    pg51, pg563,
    pg8012, pg8023, pg8265, pg16297, pg8167, pg8266, pg8275, pg4090,
    pg7161, pg7194, pg8021, pg8175, pg8263, pg8274, pg7052, pg8264, pg8273,
    pg7390, pg8261, pg8272, pg8262, pg8271, pg16355, pg24734, pg6573,
    pg7084, pg7264, pg7334, pg8007, pg8106, pg8270, pg8251, pg8260, pg4590,
    pg6642, pg6750, pg7302, pg4450, pg6225, pg26135, pg4088, pg5472,
    pg6442, pg8030, pg16437, pg25435, pg5511, pg7014, pg16399, pg16496,
    pg27380, pg6313, pg5612, pg6231, pg26149, pg5437, pg5657, pg6979,
    pg25420, pg25442, pg3993, pg6911, pg6944, pg4323, pg6712, pg6837,
    pg7519, pg25489, pg5686, pg5738, pg6447, pg26104, pg4200, pg4321,
    pg5388, pg5555, pg7229, pg5549, pg5637, pg5648, pg5747, pg5629, pg6518,
    pg7425, pg5595, pg8082, pg5695, pg6368, pg6485, pg6782, pg7961, pg7357,
    pg5796, pg7909, pg7956, pg8096, pg8258, pg8269, pg6677, pg8087, pg8249,
    pg8267, pg6895, pg7487, pg8259, pg8268  );
  input  clock;
  input  pg1943, pg1249, pg3219, pg3229, pg3217, pg3228, pg3218, pg3227,
    pg2637, pg3222, pg3233, pg3212, pg3221, pg3234, pclk, pg3220, pg3215,
    pg3226, pg3216, pg3225, pg3230, pg3213, pg3224, pg3231, pg3214, pg3223,
    pg3232, pg51, pg563;
  output pg8012, pg8023, pg8265, pg16297, pg8167, pg8266, pg8275, pg4090,
    pg7161, pg7194, pg8021, pg8175, pg8263, pg8274, pg7052, pg8264, pg8273,
    pg7390, pg8261, pg8272, pg8262, pg8271, pg16355, pg24734, pg6573,
    pg7084, pg7264, pg7334, pg8007, pg8106, pg8270, pg8251, pg8260, pg4590,
    pg6642, pg6750, pg7302, pg4450, pg6225, pg26135, pg4088, pg5472,
    pg6442, pg8030, pg16437, pg25435, pg5511, pg7014, pg16399, pg16496,
    pg27380, pg6313, pg5612, pg6231, pg26149, pg5437, pg5657, pg6979,
    pg25420, pg25442, pg3993, pg6911, pg6944, pg4323, pg6712, pg6837,
    pg7519, pg25489, pg5686, pg5738, pg6447, pg26104, pg4200, pg4321,
    pg5388, pg5555, pg7229, pg5549, pg5637, pg5648, pg5747, pg5629, pg6518,
    pg7425, pg5595, pg8082, pg5695, pg6368, pg6485, pg6782, pg7961, pg7357,
    pg5796, pg7909, pg7956, pg8096, pg8258, pg8269, pg6677, pg8087, pg8249,
    pg8267, pg6895, pg7487, pg8259, pg8268;
  reg ng3097, ng3108, ng3185, ng3135, ng141, ng155, ng258, ng83, ng369,
    ng414, ng441, ng318, ng452, ng380, ng557, ng574, ng461, ng535, ng575,
    ng590, ng490, ng646, ng703, ng714, ng722, ng736, ng821, ng835, ng849,
    ng863, ng924, ng939, ng954, ng744, ng1085, ng1113, ng1000, ng1090,
    ng969, ng992, ng1053, ng1082, ng1255, ng1173, ng1151, ng1186, ng1267,
    ng1303, ng1211, ng1352, ng1392, ng1403, ng1411, ng1425, ng1527, ng1535,
    ng1552, ng1642, ng1453, ng1739, ng1798, ng1825, ng1700, ng1834, ng1890,
    ng1945, ng1858, ng1922, ng1959, ng1973, ng1991, ng1912, ng2033, ng2082,
    ng2090, ng2104, ng2237, ng2251, ng2312, ng2327, ng2342, ng2124, ng2436,
    ng2495, ng2523, ng2362, ng2426, ng2455, ng2631, ng2648, ng2536, ng2609,
    ng2649, ng2772, ng2786, ng2797, ng2805, ng3044, ng3098, ng3107, ng3088,
    ng3139, ng145, ng154, ng261, ng88, ng358, ng411, ng444, ng317, ng286,
    ng381, ng554, ng565, ng458, ng542, ng577, ng593, ng611, ng660, ng702,
    ng715, ng724, ng734, ng817, ng839, ng848, ng921, ng882, ng936, ng957,
    ng749, ng1075, ng1115, ng1001, ng1008, ng970, ng986, ng985, ng1083,
    ng1250, ng1174, ng1171, ng1244, ng1269, ng1306, ng1206, ng1365, ng1391,
    ng1404, ng1413, ng1423, ng1523, ng1539, ng1551, ng1585, ng1448, ng1750,
    ng1801, ng1822, ng1701, ng1833, ng1893, ng1954, ng1859, ng1915, ng1960,
    ng1970, ng1871, ng1911, ng2026, ng2078, ng2094, ng2103, ng2235, ng2247,
    ng2270, ng2324, ng2345, ng2129, ng2459, ng2492, ng2394, ng2363, ng2425,
    ng2456, ng2628, ng2639, ng2533, ng2616, ng2651, ng2727, ng2784, ng2793,
    ng2809, ng3043, ng3099, ng3158, ng3179, ng3110, ng164, ng178, ng264,
    ng74, ng343, ng408, ng448, ng450, ng285, ng382, ng513, ng572, ng455,
    ng543, ng580, ng584, ng608, ng672, ng705, ng712, ng723, ng738, ng820,
    ng836, ng844, ng885, ng900, ng912, ng753, ng1078, ng1119, ng1134,
    ng1010, ng1029, ng1055, ng1210, ng1175, ng1155, ng1234, ng1268, ng1291,
    ng1216, ng1315, ng1402, ng1416, ng1420, ng1525, ng1540, ng1554, ng1573,
    ng1444, ng1765, ng1792, ng1819, ng1703, ng1660, ng1903, ng1947, ng1839,
    ng1908, ng1958, ng1979, ng1874, ng1914, ng2020, ng2080, ng2113, ng2209,
    ng2239, ng2250, ng2306, ng2285, ng2348, ng2256, ng2444, ng2489, ng2395,
    ng2529, ng2457, ng2587, ng2646, ng2530, ng2617, ng2654, ng2720, ng2777,
    ng2795, ng2810, ng3046, ng3100, ng3155, ng3182, ng3120, ng162, ng174,
    ng222, ng79, ng346, ng391, ng319, ng451, ng284, ng383, ng510, ng573,
    ng488, ng544, ng579, ng587, ng605, ng666, ng701, ng710, ng719, ng739,
    ng822, ng837, ng846, ng888, ng942, ng915, ng758, ng1095, ng1116, ng999,
    ng1009, ng1036, ng1054, ng1081, ng1142, ng1152, ng1235, ng1264, ng1215,
    ng1217, ng1312, ng1406, ng1415, ng1424, ng1524, ng1538, ng1550, ng1555,
    ng1439, ng1742, ng1795, ng1816, ng1704, ng1835, ng1904, ng1946, ng1842,
    ng1852, ng1962, ng1976, ng1877, ng1913, ng2013, ng2079, ng2111, ng2205,
    ng2240, ng2252, ng2309, ng2282, ng2160, ng2120, ng2433, ng2486, ng2397,
    ng2528, ng2458, ng2584, ng2647, ng2563, ng2618, ng2653, ng2734, ng2776,
    ng2785, ng2808, ng3045, ng2900, ng3093, ng3104, ng3173, ng3123, ng195,
    ng255, ng270, ng52, ng388, ng298, ng367, ng570, ng487, ng529, ng659,
    ng721, ng737, ng856, ng876, ng1098, ng1125, ng1141, ng976, ng1145,
    ng1214, ng1263, ng1282, ng1183, ng1407, ng1418, ng1511, ng1531, ng1534,
    ng1545, ng1435, ng1757, ng1809, ng1693, ng1696, ng1783, ng1944, ng1870,
    ng1865, ng1929, ng1939, ng1966, ng1886, ng1917, ng2089, ng2100, ng2108,
    ng2207, ng2238, ng2255, ng2315, ng2294, ng2339, ng2142, ng2418, ng2483,
    ng2398, ng2355, ng2366, ng2439, ng2644, ng2562, ng2670, ng2571, ng2610,
    ng2812, ng3048, ng3094, ng3103, ng3176, ng3124, ng198, ng252, ng213,
    ng354, ng398, ng342, ng366, ng571, ng486, ng530, ng630, ng711, ng830,
    ng860, ng873, ng1101, ng1122, ng966, ng975, ng1148, ng1158, ng1270,
    ng1285, ng1180, ng1405, ng1414, ng1515, ng1530, ng1532, ng1541, ng1430,
    ng1754, ng1807, ng1828, ng1697, ng1785, ng1949, ng1948, ng1845, ng1928,
    ng1956, ng1965, ng1887, ng1916, ng2087, ng2096, ng2112, ng2206, ng2245,
    ng2254, ng2318, ng2291, ng2297, ng2147, ng2421, ng2466, ng2396, ng2354,
    ng2374, ng2432, ng2645, ng2561, ng2652, ng2580, ng2608, ng2813, ng3047,
    ng3095, ng3106, ng3167, ng3125, ng216, ng92, ng376, ng349, ng372,
    ng324, ng531, ng633, ng698, ng840, ng861, ng918, ng1002, ng1089, ng967,
    ng978, ng1164, ng1245, ng1272, ng1288, ng1193, ng1409, ng1417, ng1512,
    ng1526, ng1536, ng1544, ng1426, ng1769, ng1804, ng1830, ng1698, ng1832,
    ng1950, ng1868, ng1860, ng1924, ng1957, ng1967, ng2040, ng2081, ng2091,
    ng2099, ng2109, ng2117, ng2246, ng2261, ng2273, ng2288, ng2300, ng2133,
    ng2384, ng2463, ng2478, ng2357, ng2364, ng2428, ng2447, ng2399, ng2656,
    ng2676, ng2607, ng2811, ng3096, ng3105, ng3170, ng3126, ng219, ng273,
    ng56, ng368, ng379, ng397, ng532, ng640, ng653, ng847, ng859, ng879,
    ng1003, ng1091, ng968, ng977, ng1221, ng1262, ng1271, ng1300, ng1192,
    ng1410, ng1419, ng1513, ng1528, ng1537, ng1546, ng1735, ng1779, ng1808,
    ng1829, ng1699, ng1831, ng1951, ng1867, ng1861, ng1923, ng1955, ng1964,
    ng2052, ng2083, ng2092, ng2101, ng2110, ng2119, ng2244, ng2253, ng2276,
    ng2330, ng2303, ng2138, ng2429, ng2473, ng2479, ng2356, ng2365, ng2427,
    ng2454, ng2472, ng2657, ng2673, ng2568, ng3049, ng2888, ng130, ng144,
    ng158, ng172, ng192, ng207, ng449, ng322, ng279, ng290, ng357, ng578,
    ng599, ng506, ng537, ng700, ng838, ng852, ng866, ng894, ng909, ng1137,
    ng972, ng1044, ng1070, ng1209, ng1294, ng1223, ng1332, ng1389, ng1400,
    ng1560, ng1582, ng1597, ng1466, ng1666, ng1730, ng1753, ng1705, ng2217,
    ng2231, ng2248, ng2503, ng2387, ng2477, ng2359, ng2417, ng2443, ng2655,
    ng2691, ng2599, ng2704, ng2766, ng2783, ng2794, ng3050, ng3062, ng3073,
    ng3013, ng45, ng20, ng2896, ng131, ng146, ng156, ng168, ng231, ng204,
    ng427, ng323, ng454, ng291, ng353, ng582, ng596, ng507, ng536, ng707,
    ng831, ng850, ng862, ng897, ng951, ng1138, ng971, ng1051, ng1069,
    ng1252, ng1273, ng1224, ng1339, ng1387, ng1396, ng1561, ng1579, ng1600,
    ng1654, ng1667, ng1723, ng1760, ng1778, ng2221, ng2230, ng2264, ng2501,
    ng2522, ng2525, ng2358, ng2424, ng2442, ng2659, ng2688, ng2603, ng2615,
    ng2773, ng2782, ng2804, ng3051, ng3061, ng3074, ng3002, ng42, ng23,
    ng2892, ng129, ng149, ng153, ng170, ng234, ng249, ng428, ng312, ng453,
    ng299, ng365, ng484, ng549, ng520, ng541, ng720, ng826, ng857, ng865,
    ng767, ng1045, ng1139, ng974, ng1052, ng1196, ng1251, ng1276, ng1177,
    ng1227, ng1358, ng1384, ng1398, ng1529, ng1543, ng1559, ng1624, ng1636,
    ng1651, ng1784, ng1668, ng1732, ng1748, ng1777, ng2222, ng2233, ng2321,
    ng2504, ng2389, ng2526, ng2361, ng2380, ng2441, ng2559, ng2623, ng2660,
    ng2679, ng2581, ng2612, ng2774, ng2792, ng2803, ng3052, ng3064, ng3071,
    ng3006, ng39, ng11, ng1, ng2903, ng133, ng148, ng157, ng169, ng237,
    ng210, ng426, ng447, ng320, ng305, ng364, ng464, ng548, ng525, ng538,
    ng730, ng728, ng858, ng867, ng762, ng1056, ng1140, ng973, ng1074,
    ng1199, ng1260, ng1279, ng1297, ng1309, ng1346, ng1388, ng1397, ng1533,
    ng1542, ng1567, ng1621, ng1594, ng1648, ng1695, ng1669, ng1731, ng1749,
    ng1776, ng2220, ng2229, ng2333, ng2507, ng2388, ng2527, ng2360, ng2373,
    ng2440, ng2539, ng2622, ng2658, ng2694, ng2594, ng2611, ng2781, ng2790,
    ng2799, ng3053, ng3063, ng3072, ng2998, ng27, ng17, ng2817, ng3101,
    ng3164, ng134, ng151, ng159, ng176, ng179, ng240, ng225, ng65, ng373,
    ng429, ng314, ng404, ng283, ng350, ng387, ng524, ng568, ng480, ng465,
    ng558, ng585, ng620, ng679, ng704, ng718, ng729, ng732, ng853, ng834,
    ng845, ng927, ng906, ng776, ng1033, ng1048, ng1107, ng1135, ng1007,
    ng1037, ng1066, ng1240, ng1259, ng1165, ng1229, ng1266, ng1218, ng1345,
    ng1385, ng1393, ng1421, ng1514, ng1553, ng1615, ng1630, ng1609, ng1813,
    ng1662, ng1680, ng1746, ng1775, ng2224, ng2232, ng2156, ng2510, ng2391,
    ng2462, ng2598, ng2642, ng2555, ng2540, ng2632, ng2661, ng2685, ng2606,
    ng2746, ng2779, ng2787, ng2801, ng3054, ng3055, ng3066, ng3077, ng3028,
    ng3040, ng3083, ng2990, ng2933, ng3102, ng3161, ng132, ng147, ng163,
    ng175, ng177, ng201, ng228, ng70, ng423, ng432, ng313, ng402, ng282,
    ng287, ng394, ng523, ng489, ng479, ng468, ng499, ng586, ng617, ng686,
    ng706, ng716, ng725, ng733, ng823, ng832, ng841, ng930, ng903, ng771,
    ng1030, ng1071, ng1104, ng1136, ng1006, ng1038, ng1059, ng1243, ng1258,
    ng1253, ng1230, ng1265, ng1219, ng1316, ng1386, ng1395, ng1422, ng1516,
    ng1557, ng1612, ng1633, ng1606, ng1789, ng1663, ng1672, ng1747, ng1768,
    ng2225, ng2234, ng2258, ng2513, ng2390, ng2469, ng2597, ng2564, ng2554,
    ng2543, ng2574, ng2664, ng2682, ng2707, ng2740, ng2775, ng2791, ng2800,
    ng2802, ng3056, ng3065, ng3078, ng3018, ng2986, ng36, ng2991, ng2950,
    ng3191, ng185, ng142, ng150, ng160, ng171, ng186, ng246, ng267, ng361,
    ng420, ng435, ng316, ng321, ng281, ng288, ng352, ng395, ng569, ng566,
    ng478, ng471, ng576, ng583, ng614, ng493, ng534, ng692, ng709, ng713,
    ng727, ng731, ng819, ng829, ng843, ng864, ng933, ng948, ng960, ng1041,
    ng1060, ng1114, ng1128, ng1005, ng1039, ng1068, ng1084, ng1257, ng1254,
    ng1167, ng1261, ng1220, ng1319, ng1372, ng1394, ng1401, ng1412, ng1558,
    ng1576, ng1588, ng1603, ng1727, ng1664, ng1679, ng1738, ng1764, ng2448,
    ng2516, ng2393, ng2470, ng2643, ng2640, ng2553, ng2546, ng2650, ng2667,
    ng2604, ng2714, ng2753, ng2778, ng2788, ng2796, ng2806, ng3080, ng3057,
    ng3068, ng3075, ng3024, ng2987, ng2992, ng8, ng2883, ng3128, ng3147,
    ng143, ng152, ng161, ng173, ng189, ng243, ng61, ng384, ng417, ng438,
    ng315, ng403, ng280, ng289, ng351, ng396, ng564, ng567, ng477, ng528,
    ng559, ng581, ng602, ng496, ng533, ng699, ng708, ng717, ng726, ng735,
    ng818, ng833, ng842, ng851, ng891, ng945, ng780, ng740, ng1063, ng1110,
    ng1131, ng1004, ng1040, ng1067, ng1011, ng1256, ng1176, ng1166, ng1228,
    ng1222, ng1326, ng1378, ng1390, ng1399, ng1408, ng1556, ng1618, ng1591,
    ng1645, ng1457, ng1665, ng1686, ng1745, ng1763, ng2498, ng2519, ng2392,
    ng2471, ng2638, ng2641, ng2552, ng2602, ng2633, ng2565, ng2605, ng2733,
    ng2760, ng2780, ng2789, ng2798, ng2807, ng3079, ng3058, ng3067, ng3076,
    ng3010, ng48, ng26, ng2, ng809, ng2827, ng113, ng2200, ng3084, ng3059,
    ng3070, ng2867, ng789, ng2845, ng2857, ng3085, ng3060, ng3069, ng805,
    ng2830, ng117, ng2858, ng3086, ng2997, ng3032, ng2814, ng2870, ng785,
    ng2842, ng97, ng3087, ng2993, ng3036, ng2908, ng2935, ng2969, ng1481,
    ng3091, ng1570, ng1670, ng1734, ng2210, ng2227, ng30, ng5, ng2912,
    ng2934, ng2972, ng1486, ng3092, ng1627, ng1671, ng1733, ng2208, ng2223,
    ng33, ng14, ng2917, ng2941, ng2963, ng1491, ng1639, ng1761, ng1937,
    ng2218, ng2226, ng2524, ng2924, ng2938, ng2966, ng1496, ng1462, ng1762,
    ng1934, ng2219, ng2228, ng2502, ng2920, ng2947, ng2981, ng2861, ng793,
    ng2839, ng1724, ng1952, ng1836, ng2085, ng2093, ng2107, ng2118, ng2451,
    ng2984, ng2944, ng2874, ng2877, ng2824, ng121, ng1772, ng1953, ng1869,
    ng2086, ng2095, ng2105, ng2114, ng2257, ng2985, ng2956, ng2975, ng1471,
    ng101, ng2170, ng1810, ng1846, ng1938, ng2084, ng2098, ng2102, ng2116,
    ng2151, ng2930, ng2953, ng2978, ng1476, ng2854, ng2175, ng1694, ng1849,
    ng1880, ng2088, ng2097, ng2106, ng2115, ng2336, ng2929, ng2962, ng801,
    ng2833, ng105, ng2180, ng2165, ng1702, ng1963, ng1994, ng1997, ng1905,
    ng2010, ng2072, ng2279, ng2879, ng2959, ng2818, ng2873, ng2851, ng2185,
    ng2878, ng1661, ng1961, ng1982, ng2000, ng1900, ng2039, ng2066, ng2267,
    ng1506, ng2864, ng797, ng2836, ng109, ng2190, ng3210, ng1985, ng1910,
    ng1918, ng2059, ng2249, ng1501, ng813, ng2821, ng125, ng2848, ng2195,
    ng3211, ng1988, ng1909, ng1921, ng2046, ng2236;
  wire new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_1_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_1_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_1_, new_n4546_,
    new_n4547_, new_n4548_, new_n4549_, new_n4550_1_, new_n4551_,
    new_n4552_, new_n4553_, new_n4554_, new_n4555_1_, new_n4556_,
    new_n4557_, new_n4558_, new_n4559_, new_n4560_1_, new_n4561_,
    new_n4562_, new_n4563_, new_n4564_1_, new_n4565_, new_n4566_,
    new_n4567_, new_n4568_, new_n4569_1_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_1_, new_n4574_, new_n4575_, new_n4576_,
    new_n4577_1_, new_n4578_, new_n4579_, new_n4580_, new_n4581_1_,
    new_n4582_, new_n4583_, new_n4584_, new_n4585_1_, new_n4586_,
    new_n4587_, new_n4588_, new_n4589_, new_n4590_1_, new_n4591_,
    new_n4592_, new_n4593_, new_n4594_, new_n4595_1_, new_n4596_,
    new_n4597_, new_n4598_, new_n4599_1_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_1_, new_n4605_, new_n4606_,
    new_n4607_, new_n4608_, new_n4609_1_, new_n4610_, new_n4611_,
    new_n4612_, new_n4613_, new_n4614_1_, new_n4615_, new_n4616_,
    new_n4617_, new_n4618_, new_n4620_, new_n4621_, new_n4622_, new_n4623_,
    new_n4625_, new_n4627_, new_n4628_, new_n4629_1_, new_n4630_,
    new_n4631_, new_n4632_, new_n4633_, new_n4634_1_, new_n4635_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_1_, new_n4640_,
    new_n4641_, new_n4642_, new_n4643_, new_n4644_1_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4650_, new_n4651_, new_n4652_,
    new_n4653_, new_n4654_1_, new_n4655_, new_n4656_, new_n4657_1_,
    new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_1_,
    new_n4663_, new_n4664_, new_n4665_, new_n4666_1_, new_n4667_,
    new_n4668_, new_n4669_, new_n4670_, new_n4671_1_, new_n4672_,
    new_n4673_, new_n4674_, new_n4675_, new_n4676_1_, new_n4677_,
    new_n4678_, new_n4679_, new_n4681_1_, new_n4682_, new_n4683_,
    new_n4684_, new_n4686_1_, new_n4687_, new_n4688_, new_n4689_,
    new_n4691_1_, new_n4692_, new_n4693_, new_n4694_1_, new_n4695_,
    new_n4696_, new_n4697_, new_n4698_, new_n4699_1_, new_n4700_,
    new_n4701_, new_n4702_, new_n4703_, new_n4704_1_, new_n4705_,
    new_n4707_, new_n4708_1_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_1_, new_n4714_, new_n4715_, new_n4716_,
    new_n4717_, new_n4718_1_, new_n4719_, new_n4720_, new_n4721_,
    new_n4722_, new_n4723_1_, new_n4724_, new_n4725_, new_n4726_,
    new_n4727_, new_n4728_1_, new_n4729_, new_n4730_, new_n4731_,
    new_n4732_1_, new_n4733_, new_n4734_, new_n4735_, new_n4736_,
    new_n4737_1_, new_n4738_, new_n4739_, new_n4740_, new_n4742_1_,
    new_n4743_, new_n4744_, new_n4746_, new_n4747_1_, new_n4749_,
    new_n4750_, new_n4751_, new_n4752_1_, new_n4753_, new_n4754_,
    new_n4755_, new_n4757_1_, new_n4758_, new_n4759_, new_n4760_,
    new_n4762_1_, new_n4763_, new_n4764_, new_n4765_, new_n4767_1_,
    new_n4768_, new_n4770_, new_n4771_, new_n4773_, new_n4774_, new_n4775_,
    new_n4777_1_, new_n4778_, new_n4779_, new_n4781_, new_n4782_1_,
    new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_1_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_1_,
    new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_1_,
    new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_1_,
    new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_1_,
    new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_1_,
    new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_1_,
    new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_1_,
    new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_1_,
    new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_1_,
    new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_1_,
    new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_1_,
    new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_1_,
    new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_1_,
    new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_1_,
    new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_1_,
    new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_1_,
    new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_1_,
    new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_1_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_1_,
    new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_1_,
    new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_1_,
    new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_1_,
    new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_1_,
    new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_1_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_1_,
    new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_1_,
    new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_1_,
    new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_1_,
    new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_1_,
    new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_1_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_1_,
    new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_1_,
    new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_1_,
    new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_1_,
    new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_1_,
    new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_1_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_1_,
    new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_1_,
    new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_1_,
    new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_1_,
    new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_1_,
    new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_1_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_1_,
    new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_1_,
    new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_1_,
    new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_1_,
    new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_1_,
    new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_1_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_1_,
    new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_1_,
    new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_1_,
    new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_1_,
    new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_1_,
    new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_1_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_1_,
    new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_1_,
    new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_1_,
    new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_1_,
    new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_1_,
    new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_1_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_1_,
    new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_1_,
    new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_1_,
    new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_1_,
    new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_1_,
    new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_1_,
    new_n5118_, new_n5119_, new_n5120_, new_n5122_1_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_1_, new_n5128_,
    new_n5129_, new_n5130_, new_n5131_, new_n5132_1_, new_n5133_,
    new_n5135_, new_n5136_, new_n5137_1_, new_n5138_, new_n5139_,
    new_n5140_, new_n5141_, new_n5142_1_, new_n5143_, new_n5144_,
    new_n5145_, new_n5146_, new_n5147_1_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_, new_n5152_1_, new_n5153_, new_n5154_,
    new_n5155_, new_n5156_, new_n5157_1_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_1_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_1_, new_n5168_, new_n5169_, new_n5170_,
    new_n5171_, new_n5172_1_, new_n5174_, new_n5175_, new_n5176_,
    new_n5177_1_, new_n5178_, new_n5179_, new_n5180_, new_n5181_,
    new_n5182_1_, new_n5183_, new_n5184_, new_n5185_, new_n5186_,
    new_n5187_1_, new_n5188_, new_n5189_, new_n5190_, new_n5191_,
    new_n5192_1_, new_n5193_, new_n5194_, new_n5195_, new_n5196_,
    new_n5197_1_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_1_, new_n5203_, new_n5204_, new_n5205_, new_n5206_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_1_,
    new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_1_,
    new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_1_,
    new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_1_,
    new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_1_,
    new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_1_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5243_, new_n5244_,
    new_n5245_, new_n5246_, new_n5247_1_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_1_, new_n5253_, new_n5254_,
    new_n5255_, new_n5256_, new_n5257_1_, new_n5258_, new_n5259_,
    new_n5260_, new_n5261_, new_n5262_1_, new_n5263_, new_n5264_,
    new_n5265_, new_n5266_, new_n5267_1_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_1_, new_n5273_, new_n5274_,
    new_n5275_, new_n5277_1_, new_n5278_, new_n5280_, new_n5281_,
    new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_1_,
    new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_1_,
    new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_1_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_1_,
    new_n5303_, new_n5304_, new_n5305_1_, new_n5307_, new_n5308_,
    new_n5309_1_, new_n5310_, new_n5311_, new_n5312_, new_n5313_1_,
    new_n5314_, new_n5315_, new_n5316_1_, new_n5317_, new_n5318_,
    new_n5319_, new_n5320_, new_n5321_1_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_1_, new_n5327_, new_n5328_,
    new_n5329_, new_n5330_1_, new_n5331_, new_n5332_, new_n5333_,
    new_n5334_, new_n5335_1_, new_n5336_, new_n5337_, new_n5338_,
    new_n5339_, new_n5340_1_, new_n5341_, new_n5342_, new_n5344_,
    new_n5345_1_, new_n5346_, new_n5347_, new_n5348_, new_n5349_,
    new_n5350_1_, new_n5351_, new_n5352_, new_n5354_, new_n5355_1_,
    new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_1_,
    new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_1_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_1_, new_n5371_,
    new_n5372_, new_n5373_1_, new_n5374_, new_n5375_, new_n5376_,
    new_n5377_, new_n5378_1_, new_n5380_, new_n5381_, new_n5382_,
    new_n5383_1_, new_n5384_, new_n5385_, new_n5386_, new_n5387_,
    new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_1_,
    new_n5395_, new_n5396_, new_n5397_, new_n5399_, new_n5400_, new_n5401_,
    new_n5403_1_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_1_, new_n5409_, new_n5410_, new_n5411_, new_n5412_,
    new_n5413_1_, new_n5414_, new_n5415_, new_n5416_, new_n5417_,
    new_n5418_1_, new_n5419_, new_n5420_, new_n5421_, new_n5422_1_,
    new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_1_,
    new_n5428_, new_n5429_, new_n5430_, new_n5431_1_, new_n5432_,
    new_n5433_, new_n5434_, new_n5435_, new_n5436_1_, new_n5437_,
    new_n5438_, new_n5439_1_, new_n5440_, new_n5441_, new_n5442_,
    new_n5443_1_, new_n5444_, new_n5445_, new_n5446_, new_n5447_,
    new_n5448_1_, new_n5449_, new_n5450_, new_n5451_, new_n5452_,
    new_n5453_1_, new_n5454_, new_n5455_, new_n5456_, new_n5457_,
    new_n5458_1_, new_n5459_, new_n5460_, new_n5461_, new_n5462_,
    new_n5463_1_, new_n5464_, new_n5465_, new_n5466_, new_n5467_,
    new_n5468_1_, new_n5469_, new_n5470_, new_n5471_, new_n5472_,
    new_n5473_1_, new_n5474_, new_n5475_, new_n5476_, new_n5477_,
    new_n5478_1_, new_n5479_, new_n5480_, new_n5481_, new_n5482_,
    new_n5483_1_, new_n5484_, new_n5485_, new_n5486_, new_n5487_,
    new_n5488_1_, new_n5489_, new_n5490_, new_n5491_, new_n5492_,
    new_n5493_1_, new_n5494_, new_n5495_, new_n5496_, new_n5497_,
    new_n5498_1_, new_n5499_, new_n5500_, new_n5501_, new_n5502_,
    new_n5503_1_, new_n5504_, new_n5505_, new_n5506_, new_n5507_,
    new_n5508_1_, new_n5509_, new_n5510_, new_n5511_, new_n5512_,
    new_n5513_1_, new_n5514_, new_n5515_, new_n5517_1_, new_n5518_,
    new_n5519_, new_n5521_, new_n5522_1_, new_n5524_, new_n5525_,
    new_n5526_1_, new_n5527_, new_n5528_, new_n5529_, new_n5530_,
    new_n5532_, new_n5533_, new_n5534_, new_n5535_1_, new_n5536_,
    new_n5538_, new_n5539_, new_n5540_1_, new_n5542_, new_n5543_,
    new_n5544_, new_n5545_1_, new_n5546_, new_n5547_, new_n5548_,
    new_n5549_1_, new_n5550_, new_n5551_, new_n5552_, new_n5553_1_,
    new_n5554_, new_n5555_, new_n5556_1_, new_n5557_, new_n5558_,
    new_n5559_, new_n5560_, new_n5561_1_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_1_, new_n5567_, new_n5568_,
    new_n5569_, new_n5570_1_, new_n5571_, new_n5572_, new_n5573_,
    new_n5574_, new_n5575_1_, new_n5576_, new_n5577_, new_n5578_,
    new_n5579_, new_n5580_1_, new_n5581_, new_n5582_, new_n5583_,
    new_n5584_, new_n5585_1_, new_n5586_, new_n5587_, new_n5588_,
    new_n5589_, new_n5590_1_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_1_, new_n5596_, new_n5597_, new_n5598_,
    new_n5599_, new_n5600_1_, new_n5601_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_1_, new_n5606_, new_n5607_, new_n5608_,
    new_n5609_, new_n5610_1_, new_n5611_, new_n5612_, new_n5613_,
    new_n5614_, new_n5615_1_, new_n5616_, new_n5617_, new_n5618_,
    new_n5619_, new_n5620_1_, new_n5621_, new_n5622_, new_n5623_,
    new_n5624_, new_n5625_1_, new_n5626_, new_n5627_, new_n5628_,
    new_n5629_, new_n5630_1_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_1_, new_n5635_, new_n5636_, new_n5637_, new_n5638_,
    new_n5639_1_, new_n5640_, new_n5641_, new_n5642_, new_n5643_,
    new_n5644_1_, new_n5645_, new_n5646_, new_n5647_, new_n5648_,
    new_n5649_1_, new_n5650_, new_n5651_, new_n5652_, new_n5653_,
    new_n5654_1_, new_n5655_, new_n5656_, new_n5657_, new_n5658_,
    new_n5659_1_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_1_, new_n5665_, new_n5666_, new_n5667_, new_n5668_,
    new_n5669_1_, new_n5670_, new_n5671_, new_n5672_, new_n5673_,
    new_n5674_1_, new_n5675_, new_n5676_, new_n5677_, new_n5678_,
    new_n5679_1_, new_n5680_, new_n5681_, new_n5682_, new_n5683_,
    new_n5684_1_, new_n5685_, new_n5686_, new_n5687_, new_n5688_,
    new_n5689_1_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_1_, new_n5695_, new_n5696_, new_n5697_, new_n5698_,
    new_n5699_1_, new_n5700_, new_n5701_, new_n5702_, new_n5703_,
    new_n5704_1_, new_n5705_, new_n5706_, new_n5707_, new_n5708_,
    new_n5709_1_, new_n5710_, new_n5711_, new_n5712_, new_n5713_,
    new_n5714_1_, new_n5715_, new_n5716_, new_n5717_, new_n5718_,
    new_n5719_1_, new_n5720_, new_n5721_, new_n5722_, new_n5723_,
    new_n5724_1_, new_n5725_, new_n5726_, new_n5727_, new_n5728_,
    new_n5729_1_, new_n5730_, new_n5731_, new_n5732_, new_n5733_,
    new_n5734_1_, new_n5735_, new_n5736_, new_n5737_, new_n5738_1_,
    new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_1_,
    new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_1_,
    new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_1_,
    new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_1_,
    new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_1_,
    new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5768_1_,
    new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_1_,
    new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_1_,
    new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_1_,
    new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_1_,
    new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_1_,
    new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_1_,
    new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_1_,
    new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_1_,
    new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_1_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_1_,
    new_n5819_, new_n5820_, new_n5821_, new_n5822_, new_n5823_1_,
    new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_1_,
    new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_1_,
    new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_1_,
    new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_1_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_1_,
    new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_1_,
    new_n5854_, new_n5856_, new_n5857_, new_n5858_1_, new_n5859_,
    new_n5860_, new_n5861_, new_n5862_, new_n5863_1_, new_n5864_,
    new_n5865_, new_n5866_, new_n5867_, new_n5868_1_, new_n5869_,
    new_n5870_, new_n5871_, new_n5872_, new_n5873_1_, new_n5874_,
    new_n5875_, new_n5876_, new_n5877_, new_n5878_1_, new_n5879_,
    new_n5880_, new_n5882_, new_n5883_1_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_1_, new_n5889_, new_n5890_,
    new_n5891_, new_n5892_, new_n5893_1_, new_n5894_, new_n5895_,
    new_n5896_, new_n5897_, new_n5898_1_, new_n5899_, new_n5900_,
    new_n5901_, new_n5902_, new_n5903_1_, new_n5904_, new_n5905_,
    new_n5906_, new_n5907_, new_n5908_1_, new_n5909_, new_n5911_,
    new_n5912_, new_n5913_1_, new_n5914_, new_n5915_, new_n5916_,
    new_n5917_, new_n5918_1_, new_n5919_, new_n5920_, new_n5921_,
    new_n5923_1_, new_n5924_, new_n5925_, new_n5926_, new_n5927_,
    new_n5928_1_, new_n5929_, new_n5930_, new_n5931_, new_n5932_,
    new_n5933_1_, new_n5934_, new_n5935_, new_n5936_, new_n5937_,
    new_n5938_1_, new_n5939_, new_n5940_, new_n5941_, new_n5942_,
    new_n5943_1_, new_n5944_, new_n5945_, new_n5946_, new_n5947_,
    new_n5948_1_, new_n5949_, new_n5951_, new_n5952_, new_n5953_1_,
    new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_1_,
    new_n5959_, new_n5961_, new_n5962_1_, new_n5963_, new_n5964_,
    new_n5965_, new_n5966_, new_n5967_1_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_1_, new_n5973_, new_n5974_,
    new_n5975_, new_n5976_, new_n5977_1_, new_n5978_, new_n5979_,
    new_n5980_, new_n5981_, new_n5982_1_, new_n5983_, new_n5984_,
    new_n5985_, new_n5986_, new_n5987_1_, new_n5989_, new_n5990_,
    new_n5991_, new_n5992_1_, new_n5993_, new_n5994_, new_n5995_,
    new_n5996_, new_n5997_1_, new_n5998_, new_n5999_, new_n6000_,
    new_n6001_, new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6008_,
    new_n6009_, new_n6010_, new_n6011_, new_n6013_, new_n6014_, new_n6015_,
    new_n6016_, new_n6018_, new_n6019_, new_n6020_, new_n6021_,
    new_n6022_1_, new_n6023_, new_n6024_, new_n6026_, new_n6027_1_,
    new_n6029_, new_n6030_, new_n6031_, new_n6032_1_, new_n6033_,
    new_n6034_, new_n6035_, new_n6036_, new_n6037_1_, new_n6038_,
    new_n6039_, new_n6040_, new_n6041_, new_n6042_1_, new_n6043_,
    new_n6044_, new_n6045_, new_n6046_, new_n6047_1_, new_n6049_,
    new_n6050_, new_n6051_, new_n6052_1_, new_n6053_, new_n6054_,
    new_n6055_, new_n6056_, new_n6057_1_, new_n6058_, new_n6059_,
    new_n6060_, new_n6061_, new_n6062_1_, new_n6063_, new_n6064_,
    new_n6065_, new_n6066_, new_n6067_1_, new_n6068_, new_n6069_,
    new_n6070_, new_n6071_, new_n6072_1_, new_n6073_, new_n6074_,
    new_n6075_, new_n6076_, new_n6077_1_, new_n6078_, new_n6080_,
    new_n6081_, new_n6082_1_, new_n6083_, new_n6084_, new_n6085_,
    new_n6086_, new_n6087_1_, new_n6088_, new_n6089_, new_n6090_,
    new_n6091_, new_n6092_1_, new_n6093_, new_n6094_, new_n6095_,
    new_n6096_, new_n6097_1_, new_n6098_, new_n6099_, new_n6100_,
    new_n6101_, new_n6102_1_, new_n6103_, new_n6104_, new_n6105_,
    new_n6106_, new_n6107_1_, new_n6108_, new_n6109_, new_n6110_,
    new_n6111_, new_n6112_1_, new_n6113_, new_n6114_, new_n6115_,
    new_n6116_, new_n6117_1_, new_n6118_, new_n6119_, new_n6120_,
    new_n6121_, new_n6122_1_, new_n6123_, new_n6124_, new_n6125_,
    new_n6126_, new_n6127_1_, new_n6128_, new_n6129_, new_n6130_,
    new_n6131_, new_n6132_1_, new_n6133_, new_n6134_, new_n6135_,
    new_n6136_, new_n6137_1_, new_n6138_, new_n6139_, new_n6140_,
    new_n6141_, new_n6142_1_, new_n6143_, new_n6144_, new_n6145_,
    new_n6146_, new_n6147_1_, new_n6148_, new_n6149_, new_n6150_,
    new_n6151_, new_n6153_, new_n6154_, new_n6155_, new_n6156_,
    new_n6157_1_, new_n6158_, new_n6159_, new_n6160_, new_n6161_,
    new_n6162_1_, new_n6163_, new_n6164_, new_n6166_, new_n6167_1_,
    new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_1_,
    new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_1_,
    new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_1_,
    new_n6183_, new_n6184_, new_n6185_1_, new_n6186_, new_n6187_,
    new_n6188_, new_n6189_1_, new_n6190_, new_n6191_, new_n6192_,
    new_n6193_1_, new_n6194_, new_n6195_, new_n6196_, new_n6197_,
    new_n6198_1_, new_n6199_, new_n6200_, new_n6201_1_, new_n6202_,
    new_n6203_, new_n6204_, new_n6205_, new_n6206_1_, new_n6207_,
    new_n6208_, new_n6209_, new_n6210_, new_n6211_1_, new_n6212_,
    new_n6213_, new_n6214_1_, new_n6215_, new_n6216_, new_n6217_,
    new_n6218_, new_n6219_1_, new_n6220_, new_n6221_, new_n6222_,
    new_n6223_, new_n6224_1_, new_n6225_, new_n6226_, new_n6227_,
    new_n6228_, new_n6229_1_, new_n6230_, new_n6231_, new_n6232_,
    new_n6233_, new_n6234_1_, new_n6235_, new_n6236_, new_n6237_,
    new_n6238_, new_n6239_1_, new_n6241_, new_n6242_, new_n6243_,
    new_n6244_1_, new_n6245_, new_n6246_, new_n6247_, new_n6248_,
    new_n6249_1_, new_n6250_, new_n6251_, new_n6253_, new_n6254_1_,
    new_n6255_, new_n6256_, new_n6257_, new_n6259_1_, new_n6260_,
    new_n6261_, new_n6263_, new_n6264_1_, new_n6265_, new_n6267_,
    new_n6268_, new_n6269_1_, new_n6270_, new_n6272_, new_n6273_,
    new_n6275_, new_n6276_, new_n6278_, new_n6279_1_, new_n6280_,
    new_n6281_, new_n6282_, new_n6283_, new_n6285_, new_n6286_, new_n6287_,
    new_n6288_, new_n6289_1_, new_n6290_, new_n6291_, new_n6292_,
    new_n6293_, new_n6294_1_, new_n6295_, new_n6296_, new_n6297_,
    new_n6298_, new_n6299_1_, new_n6300_, new_n6301_, new_n6302_,
    new_n6303_, new_n6304_1_, new_n6305_, new_n6306_, new_n6307_,
    new_n6308_, new_n6309_1_, new_n6310_, new_n6311_, new_n6312_,
    new_n6313_, new_n6314_1_, new_n6315_, new_n6316_, new_n6317_,
    new_n6318_, new_n6319_1_, new_n6320_, new_n6321_, new_n6322_,
    new_n6323_1_, new_n6324_, new_n6325_, new_n6326_, new_n6327_,
    new_n6328_1_, new_n6329_, new_n6330_, new_n6331_1_, new_n6332_,
    new_n6333_, new_n6334_, new_n6335_, new_n6336_1_, new_n6337_,
    new_n6338_, new_n6339_1_, new_n6340_, new_n6341_, new_n6342_,
    new_n6343_, new_n6344_1_, new_n6345_, new_n6346_, new_n6347_,
    new_n6348_1_, new_n6349_, new_n6350_, new_n6351_, new_n6352_,
    new_n6353_1_, new_n6354_, new_n6355_, new_n6356_, new_n6357_,
    new_n6358_1_, new_n6359_, new_n6360_, new_n6361_, new_n6362_,
    new_n6363_1_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_1_, new_n6369_, new_n6370_, new_n6371_, new_n6372_,
    new_n6373_1_, new_n6374_, new_n6375_, new_n6376_, new_n6377_,
    new_n6378_1_, new_n6379_, new_n6380_, new_n6381_, new_n6382_,
    new_n6383_1_, new_n6384_, new_n6385_, new_n6386_, new_n6387_,
    new_n6388_1_, new_n6389_, new_n6390_, new_n6391_, new_n6392_,
    new_n6393_1_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_1_, new_n6399_, new_n6400_, new_n6401_, new_n6402_,
    new_n6403_1_, new_n6404_, new_n6405_, new_n6406_, new_n6407_,
    new_n6408_1_, new_n6409_, new_n6410_, new_n6411_, new_n6412_1_,
    new_n6413_, new_n6414_, new_n6415_, new_n6416_1_, new_n6417_,
    new_n6418_, new_n6419_, new_n6420_, new_n6421_1_, new_n6422_,
    new_n6423_, new_n6424_, new_n6425_1_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_1_, new_n6431_, new_n6432_,
    new_n6433_, new_n6434_, new_n6435_1_, new_n6436_, new_n6437_,
    new_n6438_, new_n6439_1_, new_n6440_, new_n6441_, new_n6442_,
    new_n6443_, new_n6444_1_, new_n6445_, new_n6446_, new_n6447_1_,
    new_n6448_, new_n6449_, new_n6450_, new_n6451_, new_n6452_1_,
    new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_1_,
    new_n6458_, new_n6459_, new_n6460_1_, new_n6461_, new_n6462_,
    new_n6463_, new_n6464_, new_n6465_1_, new_n6466_, new_n6467_,
    new_n6468_, new_n6469_, new_n6470_1_, new_n6471_, new_n6472_,
    new_n6473_, new_n6474_, new_n6475_1_, new_n6476_, new_n6477_,
    new_n6478_, new_n6479_, new_n6480_1_, new_n6481_, new_n6482_,
    new_n6483_, new_n6484_, new_n6485_1_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_1_, new_n6491_, new_n6492_,
    new_n6493_, new_n6494_, new_n6495_1_, new_n6496_, new_n6497_,
    new_n6498_, new_n6499_, new_n6500_1_, new_n6501_, new_n6502_,
    new_n6503_, new_n6504_, new_n6505_1_, new_n6506_, new_n6507_,
    new_n6508_, new_n6509_, new_n6510_1_, new_n6511_, new_n6512_,
    new_n6513_, new_n6514_, new_n6515_1_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_1_, new_n6521_, new_n6522_,
    new_n6523_, new_n6524_, new_n6525_1_, new_n6526_, new_n6527_,
    new_n6528_, new_n6529_, new_n6530_1_, new_n6531_, new_n6532_,
    new_n6533_, new_n6534_, new_n6535_1_, new_n6536_, new_n6537_,
    new_n6538_, new_n6539_, new_n6540_1_, new_n6541_, new_n6542_,
    new_n6543_, new_n6544_, new_n6545_1_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_1_, new_n6551_, new_n6552_,
    new_n6553_, new_n6554_, new_n6555_1_, new_n6556_, new_n6557_,
    new_n6558_, new_n6559_, new_n6560_1_, new_n6561_, new_n6562_,
    new_n6563_, new_n6564_, new_n6565_1_, new_n6566_, new_n6567_,
    new_n6568_, new_n6569_, new_n6570_1_, new_n6571_, new_n6572_,
    new_n6573_, new_n6574_, new_n6575_1_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_1_, new_n6581_, new_n6582_,
    new_n6583_, new_n6584_, new_n6585_1_, new_n6586_, new_n6587_,
    new_n6588_, new_n6589_, new_n6590_1_, new_n6591_, new_n6592_,
    new_n6593_, new_n6594_, new_n6595_1_, new_n6596_, new_n6597_,
    new_n6598_, new_n6599_, new_n6600_1_, new_n6601_, new_n6602_,
    new_n6603_, new_n6604_, new_n6605_1_, new_n6606_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_1_, new_n6611_, new_n6612_,
    new_n6613_, new_n6614_1_, new_n6615_, new_n6616_, new_n6617_,
    new_n6618_, new_n6619_1_, new_n6620_, new_n6621_, new_n6622_,
    new_n6623_, new_n6624_1_, new_n6626_, new_n6627_, new_n6628_,
    new_n6629_1_, new_n6630_, new_n6631_, new_n6633_1_, new_n6634_,
    new_n6635_, new_n6636_, new_n6637_, new_n6638_1_, new_n6639_,
    new_n6640_, new_n6641_, new_n6642_, new_n6643_1_, new_n6644_,
    new_n6645_, new_n6646_, new_n6647_, new_n6648_1_, new_n6649_,
    new_n6650_, new_n6651_, new_n6652_, new_n6653_1_, new_n6654_,
    new_n6655_, new_n6656_, new_n6657_1_, new_n6658_, new_n6659_,
    new_n6660_, new_n6662_1_, new_n6663_, new_n6664_, new_n6665_,
    new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_1_,
    new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_1_,
    new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_1_,
    new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_1_,
    new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_1_,
    new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_1_,
    new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_1_,
    new_n6702_, new_n6703_, new_n6704_, new_n6706_1_, new_n6707_,
    new_n6708_, new_n6709_, new_n6710_, new_n6711_1_, new_n6712_,
    new_n6713_, new_n6714_, new_n6715_1_, new_n6716_, new_n6717_,
    new_n6718_, new_n6719_, new_n6720_1_, new_n6721_, new_n6722_,
    new_n6723_, new_n6724_, new_n6725_1_, new_n6726_, new_n6727_,
    new_n6728_, new_n6729_, new_n6730_1_, new_n6731_, new_n6732_,
    new_n6733_, new_n6734_, new_n6735_1_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6741_, new_n6742_, new_n6743_, new_n6744_,
    new_n6745_1_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_1_, new_n6751_, new_n6752_, new_n6753_, new_n6754_,
    new_n6755_1_, new_n6756_, new_n6757_, new_n6758_, new_n6759_,
    new_n6760_1_, new_n6761_, new_n6762_, new_n6763_, new_n6764_,
    new_n6765_1_, new_n6766_, new_n6767_, new_n6768_, new_n6769_,
    new_n6770_1_, new_n6771_, new_n6772_, new_n6773_, new_n6775_1_,
    new_n6776_, new_n6778_, new_n6779_1_, new_n6781_, new_n6782_,
    new_n6783_1_, new_n6784_, new_n6785_, new_n6786_, new_n6787_,
    new_n6788_1_, new_n6789_, new_n6790_, new_n6791_, new_n6792_,
    new_n6793_1_, new_n6794_, new_n6795_, new_n6796_, new_n6797_,
    new_n6798_1_, new_n6799_, new_n6801_, new_n6802_, new_n6803_1_,
    new_n6804_, new_n6805_, new_n6806_, new_n6807_, new_n6808_1_,
    new_n6809_, new_n6810_, new_n6811_, new_n6812_, new_n6813_1_,
    new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_1_,
    new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_1_,
    new_n6824_, new_n6825_, new_n6827_, new_n6828_1_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_1_, new_n6834_,
    new_n6835_, new_n6837_, new_n6838_1_, new_n6839_, new_n6840_,
    new_n6841_, new_n6842_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_1_, new_n6849_, new_n6850_, new_n6851_, new_n6852_,
    new_n6853_1_, new_n6854_, new_n6855_, new_n6856_, new_n6857_,
    new_n6858_1_, new_n6859_, new_n6860_, new_n6861_, new_n6862_,
    new_n6863_1_, new_n6864_, new_n6865_, new_n6866_, new_n6867_,
    new_n6868_1_, new_n6869_, new_n6870_, new_n6871_, new_n6872_,
    new_n6873_1_, new_n6874_, new_n6875_, new_n6876_, new_n6877_1_,
    new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_1_,
    new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_1_,
    new_n6888_, new_n6889_, new_n6890_, new_n6891_, new_n6892_1_,
    new_n6893_, new_n6894_, new_n6895_, new_n6896_, new_n6897_1_,
    new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_1_,
    new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_1_,
    new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_1_,
    new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_1_,
    new_n6918_, new_n6919_, new_n6920_, new_n6921_, new_n6922_1_,
    new_n6923_, new_n6924_, new_n6925_, new_n6926_, new_n6927_1_,
    new_n6928_, new_n6929_, new_n6930_, new_n6931_1_, new_n6932_,
    new_n6933_, new_n6934_, new_n6935_, new_n6936_1_, new_n6937_,
    new_n6938_, new_n6939_, new_n6940_, new_n6941_1_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_1_, new_n6947_,
    new_n6948_, new_n6949_, new_n6950_, new_n6951_1_, new_n6952_,
    new_n6953_, new_n6954_, new_n6955_, new_n6956_1_, new_n6957_,
    new_n6958_, new_n6959_, new_n6960_, new_n6961_1_, new_n6962_,
    new_n6963_, new_n6964_, new_n6965_, new_n6966_1_, new_n6967_,
    new_n6968_, new_n6969_, new_n6970_, new_n6971_1_, new_n6972_,
    new_n6973_, new_n6974_, new_n6976_1_, new_n6977_, new_n6978_,
    new_n6979_, new_n6980_, new_n6981_1_, new_n6982_, new_n6983_,
    new_n6984_, new_n6985_, new_n6986_1_, new_n6987_, new_n6988_,
    new_n6989_, new_n6990_, new_n6991_1_, new_n6993_, new_n6994_,
    new_n6995_1_, new_n6996_, new_n6997_, new_n6998_, new_n6999_,
    new_n7001_, new_n7002_, new_n7003_, new_n7004_1_, new_n7005_,
    new_n7007_, new_n7008_, new_n7009_1_, new_n7011_, new_n7012_,
    new_n7013_, new_n7015_, new_n7016_, new_n7017_, new_n7018_,
    new_n7019_1_, new_n7020_, new_n7021_, new_n7023_, new_n7024_1_,
    new_n7026_, new_n7027_, new_n7028_, new_n7029_1_, new_n7030_,
    new_n7031_, new_n7032_, new_n7033_1_, new_n7034_, new_n7035_,
    new_n7036_, new_n7037_, new_n7038_1_, new_n7039_, new_n7040_,
    new_n7041_, new_n7042_, new_n7043_1_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_1_, new_n7049_, new_n7050_,
    new_n7051_, new_n7052_, new_n7053_1_, new_n7054_, new_n7055_,
    new_n7056_, new_n7057_, new_n7058_1_, new_n7059_, new_n7060_,
    new_n7061_, new_n7062_, new_n7063_1_, new_n7064_, new_n7065_,
    new_n7066_, new_n7067_, new_n7068_1_, new_n7069_, new_n7070_,
    new_n7071_, new_n7072_, new_n7073_1_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_1_, new_n7079_, new_n7080_,
    new_n7081_, new_n7082_1_, new_n7083_, new_n7084_, new_n7085_,
    new_n7086_, new_n7087_1_, new_n7088_, new_n7089_, new_n7090_,
    new_n7091_, new_n7092_1_, new_n7093_, new_n7094_, new_n7095_,
    new_n7096_, new_n7097_1_, new_n7098_, new_n7099_, new_n7100_,
    new_n7101_, new_n7102_1_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_1_, new_n7108_, new_n7109_, new_n7110_,
    new_n7111_, new_n7112_1_, new_n7113_, new_n7114_, new_n7115_,
    new_n7116_, new_n7117_1_, new_n7118_, new_n7119_, new_n7120_,
    new_n7121_, new_n7122_1_, new_n7123_, new_n7124_, new_n7125_,
    new_n7126_, new_n7127_1_, new_n7128_, new_n7129_, new_n7130_,
    new_n7131_1_, new_n7132_, new_n7133_, new_n7134_, new_n7135_,
    new_n7136_1_, new_n7137_, new_n7138_, new_n7139_, new_n7140_,
    new_n7141_1_, new_n7142_, new_n7143_, new_n7144_, new_n7145_1_,
    new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_1_,
    new_n7151_, new_n7152_, new_n7153_, new_n7154_, new_n7155_1_,
    new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_1_,
    new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_1_,
    new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_1_,
    new_n7171_, new_n7172_, new_n7173_, new_n7174_1_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_, new_n7179_1_, new_n7180_,
    new_n7181_, new_n7182_, new_n7183_1_, new_n7184_, new_n7185_,
    new_n7186_, new_n7187_, new_n7188_1_, new_n7189_, new_n7190_,
    new_n7191_, new_n7192_, new_n7193_1_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_1_, new_n7199_, new_n7200_,
    new_n7201_, new_n7202_, new_n7203_1_, new_n7204_, new_n7205_,
    new_n7206_, new_n7207_, new_n7208_1_, new_n7209_, new_n7210_,
    new_n7211_, new_n7212_, new_n7213_1_, new_n7214_, new_n7215_,
    new_n7216_, new_n7217_, new_n7218_1_, new_n7219_, new_n7220_,
    new_n7221_, new_n7222_, new_n7223_1_, new_n7224_, new_n7225_,
    new_n7226_, new_n7227_, new_n7228_1_, new_n7229_, new_n7230_,
    new_n7231_, new_n7232_, new_n7233_1_, new_n7234_, new_n7235_,
    new_n7236_, new_n7237_, new_n7238_1_, new_n7239_, new_n7240_,
    new_n7241_, new_n7242_, new_n7243_1_, new_n7244_, new_n7245_,
    new_n7246_, new_n7247_, new_n7248_1_, new_n7249_, new_n7250_,
    new_n7251_, new_n7252_, new_n7253_1_, new_n7254_, new_n7255_,
    new_n7256_, new_n7257_, new_n7258_1_, new_n7259_, new_n7260_,
    new_n7261_, new_n7262_1_, new_n7263_, new_n7264_, new_n7265_,
    new_n7266_, new_n7267_1_, new_n7268_, new_n7269_, new_n7270_,
    new_n7271_1_, new_n7272_, new_n7273_, new_n7274_, new_n7275_,
    new_n7276_1_, new_n7277_, new_n7278_, new_n7279_, new_n7280_,
    new_n7281_1_, new_n7282_, new_n7283_, new_n7284_, new_n7285_1_,
    new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_1_,
    new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_1_,
    new_n7296_, new_n7297_, new_n7298_, new_n7299_, new_n7300_1_,
    new_n7301_, new_n7302_, new_n7303_, new_n7304_1_, new_n7305_,
    new_n7306_, new_n7307_, new_n7308_, new_n7309_1_, new_n7310_,
    new_n7311_, new_n7312_, new_n7313_, new_n7314_1_, new_n7315_,
    new_n7316_, new_n7317_, new_n7318_, new_n7319_1_, new_n7320_,
    new_n7321_, new_n7322_, new_n7323_, new_n7324_1_, new_n7325_,
    new_n7326_, new_n7327_1_, new_n7328_, new_n7329_, new_n7330_,
    new_n7331_, new_n7332_1_, new_n7333_, new_n7334_, new_n7335_1_,
    new_n7336_, new_n7337_, new_n7338_, new_n7340_1_, new_n7341_,
    new_n7342_, new_n7343_, new_n7344_, new_n7345_1_, new_n7346_,
    new_n7347_, new_n7348_, new_n7349_, new_n7350_1_, new_n7351_,
    new_n7352_, new_n7353_, new_n7354_, new_n7355_1_, new_n7356_,
    new_n7357_, new_n7358_, new_n7359_, new_n7360_1_, new_n7361_,
    new_n7362_, new_n7363_, new_n7364_, new_n7366_, new_n7367_, new_n7368_,
    new_n7369_, new_n7370_1_, new_n7371_, new_n7372_, new_n7373_,
    new_n7374_, new_n7375_1_, new_n7376_, new_n7377_, new_n7378_,
    new_n7379_1_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_1_, new_n7385_, new_n7386_, new_n7387_1_, new_n7388_,
    new_n7389_, new_n7390_, new_n7391_, new_n7392_1_, new_n7393_,
    new_n7395_, new_n7396_1_, new_n7397_, new_n7398_, new_n7399_,
    new_n7400_, new_n7401_1_, new_n7402_, new_n7403_, new_n7404_,
    new_n7405_, new_n7407_, new_n7408_, new_n7409_, new_n7410_,
    new_n7411_1_, new_n7412_, new_n7413_, new_n7414_, new_n7415_,
    new_n7416_1_, new_n7417_, new_n7418_, new_n7419_, new_n7420_,
    new_n7421_1_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_1_, new_n7427_, new_n7428_, new_n7429_, new_n7430_,
    new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7441_, new_n7442_, new_n7443_, new_n7444_,
    new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_, new_n7450_,
    new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_, new_n7456_,
    new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_, new_n7462_,
    new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_, new_n7468_,
    new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_, new_n7474_,
    new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7480_, new_n7481_,
    new_n7482_, new_n7483_, new_n7484_, new_n7485_, new_n7486_, new_n7487_,
    new_n7488_, new_n7489_, new_n7490_, new_n7491_, new_n7492_, new_n7493_,
    new_n7494_, new_n7495_, new_n7496_, new_n7497_, new_n7498_, new_n7499_,
    new_n7500_, new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7505_,
    new_n7506_, new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_,
    new_n7512_, new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_,
    new_n7519_, new_n7520_, new_n7522_, new_n7523_, new_n7525_, new_n7526_,
    new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_,
    new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_,
    new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7545_,
    new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_,
    new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_,
    new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_,
    new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_,
    new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_,
    new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7582_,
    new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7588_, new_n7589_,
    new_n7590_, new_n7592_, new_n7593_, new_n7594_, new_n7596_, new_n7597_,
    new_n7598_, new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_,
    new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_,
    new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_,
    new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_,
    new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_,
    new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_,
    new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_,
    new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_,
    new_n7647_, new_n7648_, new_n7650_, new_n7651_, new_n7653_, new_n7654_,
    new_n7656_, new_n7657_, new_n7659_, new_n7660_, new_n7662_, new_n7663_,
    new_n7665_, new_n7666_, new_n7668_, new_n7669_, new_n7670_, new_n7672_,
    new_n7673_, new_n7674_, new_n7676_, new_n7677_, new_n7679_, new_n7680_,
    new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_,
    new_n7688_, new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_,
    new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_,
    new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_,
    new_n7706_, new_n7707_, new_n7709_, new_n7710_, new_n7712_, new_n7713_,
    new_n7715_, new_n7716_, new_n7717_, new_n7719_, new_n7720_, new_n7722_,
    new_n7723_, new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_,
    new_n7729_, new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7734_,
    new_n7735_, new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_,
    new_n7741_, new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_,
    new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_, new_n7752_,
    new_n7753_, new_n7754_, new_n7755_, new_n7756_, new_n7757_, new_n7758_,
    new_n7759_, new_n7760_, new_n7761_, new_n7762_, new_n7763_, new_n7764_,
    new_n7765_, new_n7766_, new_n7767_, new_n7768_, new_n7769_, new_n7770_,
    new_n7771_, new_n7772_, new_n7773_, new_n7774_, new_n7775_, new_n7776_,
    new_n7777_, new_n7778_, new_n7779_, new_n7780_, new_n7781_, new_n7782_,
    new_n7783_, new_n7784_, new_n7785_, new_n7786_, new_n7787_, new_n7788_,
    new_n7789_, new_n7790_, new_n7791_, new_n7792_, new_n7793_, new_n7794_,
    new_n7795_, new_n7796_, new_n7797_, new_n7798_, new_n7799_, new_n7800_,
    new_n7801_, new_n7802_, new_n7803_, new_n7804_, new_n7805_, new_n7806_,
    new_n7807_, new_n7808_, new_n7809_, new_n7810_, new_n7811_, new_n7812_,
    new_n7813_, new_n7814_, new_n7815_, new_n7816_, new_n7817_, new_n7818_,
    new_n7819_, new_n7820_, new_n7821_, new_n7822_, new_n7823_, new_n7824_,
    new_n7825_, new_n7826_, new_n7827_, new_n7828_, new_n7829_, new_n7830_,
    new_n7831_, new_n7832_, new_n7833_, new_n7834_, new_n7835_, new_n7836_,
    new_n7837_, new_n7838_, new_n7839_, new_n7840_, new_n7841_, new_n7842_,
    new_n7843_, new_n7844_, new_n7845_, new_n7846_, new_n7848_, new_n7849_,
    new_n7850_, new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_,
    new_n7856_, new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_,
    new_n7862_, new_n7863_, new_n7865_, new_n7866_, new_n7867_, new_n7868_,
    new_n7870_, new_n7871_, new_n7873_, new_n7874_, new_n7876_, new_n7877_,
    new_n7879_, new_n7880_, new_n7882_, new_n7883_, new_n7885_, new_n7886_,
    new_n7888_, new_n7889_, new_n7891_, new_n7892_, new_n7894_, new_n7895_,
    new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_,
    new_n7902_, new_n7903_, new_n7905_, new_n7906_, new_n7908_, new_n7909_,
    new_n7911_, new_n7912_, new_n7913_, new_n7915_, new_n7916_, new_n7917_,
    new_n7919_, new_n7920_, new_n7921_, new_n7923_, new_n7924_, new_n7926_,
    new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_, new_n7932_,
    new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_, new_n7938_,
    new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_, new_n7944_,
    new_n7945_, new_n7947_, new_n7948_, new_n7949_, new_n7950_, new_n7951_,
    new_n7952_, new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_,
    new_n7958_, new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_,
    new_n7964_, new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_,
    new_n7970_, new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_,
    new_n7976_, new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_,
    new_n7982_, new_n7983_, new_n7984_, new_n7985_, new_n7986_, new_n7987_,
    new_n7988_, new_n7989_, new_n7990_, new_n7991_, new_n7992_, new_n7993_,
    new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_, new_n7999_,
    new_n8001_, new_n8002_, new_n8004_, new_n8005_, new_n8007_, new_n8008_,
    new_n8009_, new_n8010_, new_n8012_, new_n8013_, new_n8014_, new_n8016_,
    new_n8017_, new_n8019_, new_n8020_, new_n8021_, new_n8022_, new_n8023_,
    new_n8025_, new_n8026_, new_n8027_, new_n8028_, new_n8030_, new_n8031_,
    new_n8032_, new_n8033_, new_n8035_, new_n8036_, new_n8038_, new_n8039_,
    new_n8041_, new_n8042_, new_n8044_, new_n8045_, new_n8046_, new_n8048_,
    new_n8049_, new_n8051_, new_n8052_, new_n8054_, new_n8055_, new_n8057_,
    new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_,
    new_n8064_, new_n8065_, new_n8067_, new_n8068_, new_n8069_, new_n8070_,
    new_n8072_, new_n8073_, new_n8074_, new_n8076_, new_n8077_, new_n8079_,
    new_n8080_, new_n8082_, new_n8083_, new_n8085_, new_n8086_, new_n8088_,
    new_n8089_, new_n8090_, new_n8092_, new_n8093_, new_n8095_, new_n8096_,
    new_n8097_, new_n8098_, new_n8099_, new_n8100_, new_n8101_, new_n8102_,
    new_n8104_, new_n8105_, new_n8106_, new_n8107_, new_n8109_, new_n8110_,
    new_n8112_, new_n8113_, new_n8115_, new_n8116_, new_n8118_, new_n8119_,
    new_n8121_, new_n8122_, new_n8123_, new_n8125_, new_n8126_, new_n8127_,
    new_n8128_, new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_,
    new_n8134_, new_n8136_, new_n8137_, new_n8139_, new_n8140_, new_n8142_,
    new_n8143_, new_n8144_, new_n8146_, new_n8147_, new_n8148_, new_n8149_,
    new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_, new_n8155_,
    new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_, new_n8161_,
    new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8167_, new_n8168_,
    new_n8170_, new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_,
    new_n8176_, new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_,
    new_n8182_, new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_,
    new_n8188_, new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_,
    new_n8194_, new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_,
    new_n8200_, new_n8201_, new_n8202_, new_n8204_, new_n8206_, new_n8207_,
    new_n8209_, new_n8210_, new_n8211_, new_n8213_, new_n8214_, new_n8215_,
    new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8221_, new_n8222_,
    new_n8224_, new_n8225_, new_n8227_, new_n8228_, new_n8229_, new_n8230_,
    new_n8231_, new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_,
    new_n8237_, new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_,
    new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_,
    new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_,
    new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_,
    new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_,
    new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_,
    new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_,
    new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_,
    new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_,
    new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_,
    new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_,
    new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_,
    new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_,
    new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_,
    new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_,
    new_n8327_, new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_,
    new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_,
    new_n8339_, new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_,
    new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_,
    new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8357_, new_n8358_,
    new_n8360_, new_n8361_, new_n8363_, new_n8364_, new_n8366_, new_n8367_,
    new_n8369_, new_n8370_, new_n8372_, new_n8373_, new_n8375_, new_n8376_,
    new_n8377_, new_n8378_, new_n8379_, new_n8381_, new_n8382_, new_n8383_,
    new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8389_,
    new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_, new_n8395_,
    new_n8396_, new_n8397_, new_n8398_, new_n8399_, new_n8401_, new_n8402_,
    new_n8404_, new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_,
    new_n8410_, new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_,
    new_n8417_, new_n8418_, new_n8420_, new_n8421_, new_n8422_, new_n8423_,
    new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_,
    new_n8431_, new_n8432_, new_n8434_, new_n8435_, new_n8436_, new_n8437_,
    new_n8438_, new_n8439_, new_n8440_, new_n8442_, new_n8443_, new_n8445_,
    new_n8446_, new_n8447_, new_n8448_, new_n8450_, new_n8451_, new_n8453_,
    new_n8454_, new_n8456_, new_n8457_, new_n8459_, new_n8460_, new_n8461_,
    new_n8462_, new_n8464_, new_n8465_, new_n8467_, new_n8468_, new_n8470_,
    new_n8471_, new_n8473_, new_n8474_, new_n8476_, new_n8477_, new_n8478_,
    new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_,
    new_n8485_, new_n8487_, new_n8488_, new_n8489_, new_n8490_, new_n8491_,
    new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_, new_n8498_,
    new_n8499_, new_n8500_, new_n8502_, new_n8503_, new_n8504_, new_n8506_,
    new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_,
    new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_,
    new_n8519_, new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_,
    new_n8525_, new_n8526_, new_n8527_, new_n8529_, new_n8530_, new_n8531_,
    new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_,
    new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_,
    new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_,
    new_n8550_, new_n8552_, new_n8553_, new_n8554_, new_n8556_, new_n8557_,
    new_n8559_, new_n8560_, new_n8562_, new_n8563_, new_n8564_, new_n8566_,
    new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_,
    new_n8573_, new_n8574_, new_n8575_, new_n8577_, new_n8578_, new_n8580_,
    new_n8581_, new_n8583_, new_n8584_, new_n8585_, new_n8586_, new_n8587_,
    new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_, new_n8593_,
    new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_, new_n8599_,
    new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_, new_n8605_,
    new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_, new_n8611_,
    new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_, new_n8617_,
    new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_, new_n8623_,
    new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_, new_n8629_,
    new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_, new_n8635_,
    new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_, new_n8641_,
    new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_, new_n8647_,
    new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_, new_n8653_,
    new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_, new_n8659_,
    new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_, new_n8665_,
    new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_, new_n8671_,
    new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_, new_n8677_,
    new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_, new_n8683_,
    new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_, new_n8689_,
    new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_, new_n8695_,
    new_n8697_, new_n8698_, new_n8700_, new_n8701_, new_n8703_, new_n8704_,
    new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_,
    new_n8712_, new_n8713_, new_n8714_, new_n8716_, new_n8717_, new_n8718_,
    new_n8719_, new_n8721_, new_n8722_, new_n8723_, new_n8724_, new_n8725_,
    new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_,
    new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_,
    new_n8738_, new_n8739_, new_n8741_, new_n8742_, new_n8743_, new_n8744_,
    new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_, new_n8750_,
    new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_, new_n8756_,
    new_n8757_, new_n8758_, new_n8759_, new_n8761_, new_n8762_, new_n8764_,
    new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_,
    new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8776_, new_n8777_,
    new_n8779_, new_n8780_, new_n8781_, new_n8783_, new_n8784_, new_n8785_,
    new_n8787_, new_n8788_, new_n8790_, new_n8791_, new_n8792_, new_n8794_,
    new_n8795_, new_n8797_, new_n8798_, new_n8800_, new_n8801_, new_n8803_,
    new_n8804_, new_n8806_, new_n8807_, new_n8809_, new_n8810_, new_n8812_,
    new_n8813_, new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_,
    new_n8819_, new_n8820_, new_n8822_, new_n8823_, new_n8825_, new_n8826_,
    new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_, new_n8833_,
    new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_, new_n8839_,
    new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_, new_n8845_,
    new_n8846_, new_n8848_, new_n8849_, new_n8851_, new_n8852_, new_n8853_,
    new_n8854_, new_n8856_, new_n8857_, new_n8859_, new_n8860_, new_n8861_,
    new_n8862_, new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_,
    new_n8869_, new_n8870_, new_n8871_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8878_, new_n8879_, new_n8881_, new_n8882_, new_n8884_,
    new_n8885_, new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_,
    new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_,
    new_n8898_, new_n8900_, new_n8901_, new_n8903_, new_n8905_, new_n8906_,
    new_n8908_, new_n8909_, new_n8911_, new_n8912_, new_n8914_, new_n8915_,
    new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8933_, new_n8934_,
    new_n8935_, new_n8937_, new_n8938_, new_n8939_, new_n8941_, new_n8942_,
    new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_, new_n8948_,
    new_n8950_, new_n8951_, new_n8953_, new_n8954_, new_n8956_, new_n8957_,
    new_n8959_, new_n8960_, new_n8961_, new_n8963_, new_n8964_, new_n8966_,
    new_n8967_, new_n8969_, new_n8970_, new_n8971_, new_n8972_, new_n8974_,
    new_n8975_, new_n8977_, new_n8978_, new_n8980_, new_n8981_, new_n8983_,
    new_n8984_, new_n8985_, new_n8987_, new_n8988_, new_n8990_, new_n8991_,
    new_n8993_, new_n8994_, new_n8996_, new_n8997_, new_n8999_, new_n9000_,
    new_n9002_, new_n9003_, new_n9005_, new_n9006_, new_n9007_, new_n9009_,
    new_n9010_, new_n9011_, new_n9012_, new_n9013_, new_n9014_, new_n9015_,
    new_n9016_, new_n9017_, new_n9018_, new_n9019_, new_n9020_, new_n9021_,
    new_n9022_, new_n9023_, new_n9024_, new_n9025_, new_n9026_, new_n9028_,
    new_n9029_, new_n9031_, new_n9032_, new_n9034_, new_n9035_, new_n9036_,
    new_n9038_, new_n9039_, new_n9041_, new_n9042_, new_n9044_, new_n9045_,
    new_n9046_, new_n9047_, new_n9049_, new_n9050_, new_n9051_, new_n9052_,
    new_n9053_, new_n9054_, new_n9055_, new_n9056_, new_n9057_, new_n9059_,
    new_n9060_, new_n9062_, new_n9063_, new_n9064_, new_n9066_, new_n9067_,
    new_n9068_, new_n9070_, new_n9071_, new_n9073_, new_n9074_, new_n9076_,
    new_n9077_, new_n9079_, new_n9080_, new_n9082_, new_n9083_, new_n9084_,
    new_n9085_, new_n9087_, new_n9088_, new_n9089_, new_n9091_, new_n9092_,
    new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_, new_n9099_,
    new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_, new_n9106_,
    new_n9107_, new_n9108_, new_n9110_, new_n9111_, new_n9113_, new_n9114_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_,
    new_n9128_, new_n9130_, new_n9131_, new_n9133_, new_n9134_, new_n9136_,
    new_n9137_, new_n9138_, new_n9140_, new_n9141_, new_n9143_, new_n9144_,
    new_n9145_, new_n9147_, new_n9148_, new_n9150_, new_n9151_, new_n9153_,
    new_n9154_, new_n9156_, new_n9157_, new_n9159_, new_n9160_, new_n9162_,
    new_n9163_, new_n9164_, new_n9166_, new_n9167_, new_n9168_, new_n9169_,
    new_n9171_, new_n9172_, new_n9173_, new_n9175_, new_n9176_, new_n9178_,
    new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_, new_n9184_,
    new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9190_, new_n9191_,
    new_n9193_, new_n9194_, new_n9196_, new_n9197_, new_n9198_, new_n9200_,
    new_n9201_, new_n9202_, new_n9203_, new_n9205_, new_n9206_, new_n9208_,
    new_n9209_, new_n9211_, new_n9212_, new_n9214_, new_n9215_, new_n9216_,
    new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_,
    new_n9223_, new_n9224_, new_n9225_, new_n9227_, new_n9228_, new_n9229_,
    new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_,
    new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_,
    new_n9242_, new_n9244_, new_n9245_, new_n9247_, new_n9248_, new_n9250_,
    new_n9251_, new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_,
    new_n9258_, new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9264_,
    new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_,
    new_n9271_, new_n9272_, new_n9273_, new_n9275_, new_n9276_, new_n9277_,
    new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_,
    new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_, new_n9290_,
    new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_,
    new_n9297_, new_n9299_, new_n9300_, new_n9302_, new_n9303_, new_n9304_,
    new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_, new_n9310_,
    new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_, new_n9316_,
    new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_, new_n9322_,
    new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_, new_n9328_,
    new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_, new_n9334_,
    new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_, new_n9340_,
    new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_,
    new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_,
    new_n9353_, new_n9354_, new_n9356_, new_n9357_, new_n9359_, new_n9360_,
    new_n9362_, new_n9363_, new_n9365_, new_n9366_, new_n9367_, new_n9369_,
    new_n9370_, new_n9371_, new_n9372_, new_n9373_, new_n9375_, new_n9376_,
    new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_,
    new_n9383_, new_n9385_, new_n9386_, new_n9388_, new_n9389_, new_n9390_,
    new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9397_,
    new_n9398_, new_n9400_, new_n9401_, new_n9402_, new_n9403_, new_n9404_,
    new_n9405_, new_n9406_, new_n9407_, new_n9408_, new_n9409_, new_n9410_,
    new_n9412_, new_n9413_, new_n9414_, new_n9416_, new_n9417_, new_n9418_,
    new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9425_,
    new_n9426_, new_n9428_, new_n9429_, new_n9431_, new_n9432_, new_n9434_,
    new_n9435_, new_n9437_, new_n9438_, new_n9440_, new_n9441_, new_n9443_,
    new_n9444_, new_n9445_, new_n9446_, new_n9448_, new_n9449_, new_n9451_,
    new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_, new_n9457_,
    new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_, new_n9464_,
    new_n9465_, new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_,
    new_n9471_, new_n9472_, new_n9473_, new_n9474_, new_n9475_, new_n9476_,
    new_n9478_, new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_,
    new_n9484_, new_n9485_, new_n9486_, new_n9487_, new_n9488_, new_n9489_,
    new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_,
    new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_,
    new_n9502_, new_n9503_, new_n9505_, new_n9506_, new_n9507_, new_n9508_,
    new_n9510_, new_n9511_, new_n9513_, new_n9514_, new_n9515_, new_n9516_,
    new_n9518_, new_n9519_, new_n9520_, new_n9521_, new_n9522_, new_n9523_,
    new_n9524_, new_n9526_, new_n9527_, new_n9529_, new_n9530_, new_n9532_,
    new_n9533_, new_n9535_, new_n9536_, new_n9538_, new_n9539_, new_n9541_,
    new_n9542_, new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_,
    new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_,
    new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_, new_n9561_,
    new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9567_, new_n9568_,
    new_n9569_, new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_,
    new_n9575_, new_n9576_, new_n9578_, new_n9579_, new_n9580_, new_n9582_,
    new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_,
    new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9594_, new_n9595_,
    new_n9597_, new_n9598_, new_n9599_, new_n9601_, new_n9602_, new_n9604_,
    new_n9605_, new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_,
    new_n9611_, new_n9612_, new_n9614_, new_n9615_, new_n9616_, new_n9617_,
    new_n9618_, new_n9619_, new_n9621_, new_n9622_, new_n9623_, new_n9624_,
    new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9630_, new_n9631_,
    new_n9632_, new_n9633_, new_n9635_, new_n9636_, new_n9637_, new_n9638_,
    new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_,
    new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9650_, new_n9651_,
    new_n9653_, new_n9654_, new_n9656_, new_n9657_, new_n9659_, new_n9660_,
    new_n9662_, new_n9663_, new_n9665_, new_n9666_, new_n9667_, new_n9668_,
    new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_, new_n9675_,
    new_n9676_, new_n9678_, new_n9679_, new_n9681_, new_n9682_, new_n9684_,
    new_n9685_, new_n9687_, new_n9688_, new_n9690_, new_n9691_, new_n9693_,
    new_n9694_, new_n9696_, new_n9697_, new_n9699_, new_n9700_, new_n9702_,
    new_n9703_, new_n9705_, new_n9706_, new_n9708_, new_n9709_, new_n9711_,
    new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_,
    new_n9719_, new_n9720_, new_n9722_, new_n9723_, new_n9725_, new_n9726_,
    new_n9728_, new_n9729_, new_n9730_, new_n9732_, new_n9733_, new_n9735_,
    new_n9736_, new_n9738_, new_n9739_, new_n9741_, new_n9742_, new_n9744_,
    new_n9745_, new_n9746_, new_n9747_, new_n9749_, new_n9750_, new_n9752_,
    new_n9753_, new_n9754_, new_n9756_, new_n9757_, new_n9758_, new_n9759_,
    new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_,
    new_n9766_, new_n9767_, new_n9769_, new_n9770_, new_n9772_, new_n9773_,
    new_n9774_, new_n9776_, new_n9777_, new_n9779_, new_n9780_, new_n9781_,
    new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_,
    new_n9788_, new_n9789_, new_n9791_, new_n9792_, new_n9794_, new_n9795_,
    new_n9797_, new_n9798_, new_n9800_, new_n9801_, new_n9802_, new_n9804_,
    new_n9805_, new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_,
    new_n9813_, new_n9814_, new_n9816_, new_n9817_, new_n9819_, new_n9820_,
    new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_, new_n9827_,
    new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9833_, new_n9834_,
    new_n9835_, new_n9837_, new_n9838_, new_n9840_, new_n9841_, new_n9842_,
    new_n9843_, new_n9844_, new_n9845_, new_n9846_, new_n9847_, new_n9849_,
    new_n9850_, new_n9851_, new_n9853_, new_n9854_, new_n9856_, new_n9857_,
    new_n9859_, new_n9860_, new_n9861_, new_n9863_, new_n9864_, new_n9865_,
    new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_, new_n9871_,
    new_n9872_, new_n9873_, new_n9874_, new_n9876_, new_n9877_, new_n9879_,
    new_n9880_, new_n9882_, new_n9883_, new_n9885_, new_n9886_, new_n9888_,
    new_n9889_, new_n9890_, new_n9892_, new_n9893_, new_n9894_, new_n9895_,
    new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_, new_n9901_,
    new_n9902_, new_n9904_, new_n9905_, new_n9906_, new_n9908_, new_n9909_,
    new_n9911_, new_n9912_, new_n9914_, new_n9915_, new_n9917_, new_n9918_,
    new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_,
    new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_,
    new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9950_,
    new_n9951_, new_n9953_, new_n9954_, new_n9956_, new_n9957_, new_n9959_,
    new_n9960_, new_n9962_, new_n9963_, new_n9965_, new_n9966_, new_n9968_,
    new_n9969_, new_n9971_, new_n9972_, new_n9974_, new_n9975_, new_n9977_,
    new_n9978_, new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9985_,
    new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_, new_n9991_,
    new_n9992_, new_n9994_, new_n9995_, new_n9997_, new_n9998_, new_n9999_,
    new_n10001_, new_n10002_, new_n10004_, new_n10005_, new_n10007_,
    new_n10008_, new_n10010_, new_n10011_, new_n10013_, new_n10014_,
    new_n10016_, new_n10017_, new_n10018_, new_n10019_, new_n10021_,
    new_n10022_, new_n10024_, new_n10025_, new_n10027_, new_n10028_,
    new_n10030_, new_n10031_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10038_, new_n10039_, new_n10041_, new_n10042_,
    new_n10043_, new_n10044_, new_n10045_, new_n10046_, new_n10047_,
    new_n10048_, new_n10049_, new_n10051_, new_n10052_, new_n10054_,
    new_n10055_, new_n10057_, new_n10058_, new_n10060_, new_n10061_,
    new_n10062_, new_n10064_, new_n10065_, new_n10067_, new_n10068_,
    new_n10069_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10083_, new_n10084_, new_n10086_,
    new_n10087_, new_n10088_, new_n10090_, new_n10091_, new_n10093_,
    new_n10094_, new_n10096_, new_n10097_, new_n10099_, new_n10100_,
    new_n10102_, new_n10103_, new_n10105_, new_n10106_, new_n10107_,
    new_n10109_, new_n10110_, new_n10111_, new_n10113_, new_n10114_,
    new_n10115_, new_n10117_, new_n10118_, new_n10120_, new_n10121_,
    new_n10123_, new_n10124_, new_n10126_, new_n10127_, new_n10129_,
    new_n10130_, new_n10132_, new_n10133_, new_n10135_, new_n10136_,
    new_n10138_, new_n10139_, new_n10141_, new_n10142_, new_n10144_,
    new_n10145_, new_n10147_, new_n10148_, new_n10150_, new_n10151_,
    new_n10153_, new_n10154_, new_n10156_, new_n10157_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10171_, new_n10172_, new_n10174_, new_n10175_, new_n10176_,
    new_n10178_, new_n10179_, new_n10180_, new_n10182_, new_n10183_,
    new_n10185_, new_n10186_, new_n10188_, new_n10189_, new_n10191_,
    new_n10192_, new_n10193_, new_n10194_, new_n10196_, new_n10197_,
    new_n10199_, new_n10200_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10207_, new_n10208_, new_n10210_, new_n10211_,
    new_n10213_, new_n10214_, new_n10216_, new_n10217_, new_n10219_,
    new_n10220_, new_n10221_, new_n10223_, new_n10224_, new_n10226_,
    new_n10227_, new_n10229_, new_n10230_, new_n10232_, new_n10233_,
    new_n10235_, new_n10236_, new_n10238_, new_n10239_, new_n10240_,
    new_n10242_, new_n10243_, new_n10245_, new_n10246_, new_n10248_,
    new_n10249_, new_n10251_, new_n10252_, new_n10254_, new_n10255_,
    new_n10257_, new_n10258_, new_n10260_, new_n10261_, new_n10262_,
    new_n10263_, new_n10264_, new_n10265_, new_n10266_, new_n10267_,
    new_n10268_, new_n10269_, new_n10270_, new_n10271_, new_n10272_,
    new_n10273_, new_n10274_, new_n10275_, new_n10276_, new_n10277_,
    new_n10278_, new_n10279_, new_n10280_, new_n10282_, new_n10283_,
    new_n10284_, new_n10286_, new_n10287_, new_n10289_, new_n10290_,
    new_n10292_, new_n10293_, new_n10295_, new_n10296_, new_n10298_,
    new_n10299_, new_n10300_, new_n10301_, new_n10302_, new_n10303_,
    new_n10304_, new_n10305_, new_n10306_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10318_, new_n10319_, new_n10320_,
    new_n10322_, new_n10323_, new_n10324_, new_n10325_, new_n10326_,
    new_n10327_, new_n10328_, new_n10329_, new_n10330_, new_n10331_,
    new_n10332_, new_n10334_, new_n10335_, new_n10337_, new_n10338_,
    new_n10339_, new_n10341_, new_n10342_, new_n10344_, new_n10345_,
    new_n10347_, new_n10348_, new_n10350_, new_n10351_, new_n10353_,
    new_n10354_, new_n10355_, new_n10356_, new_n10357_, new_n10358_,
    new_n10359_, new_n10360_, new_n10361_, new_n10363_, new_n10364_,
    new_n10366_, new_n10367_, new_n10369_, new_n10370_, new_n10371_,
    new_n10373_, new_n10374_, new_n10376_, new_n10377_, new_n10379_,
    new_n10380_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10394_, new_n10395_, new_n10396_,
    new_n10397_, new_n10398_, new_n10399_, new_n10400_, new_n10401_,
    new_n10402_, new_n10404_, new_n10405_, new_n10406_, new_n10408_,
    new_n10409_, new_n10411_, new_n10412_, new_n10414_, new_n10415_,
    new_n10417_, new_n10418_, new_n10419_, new_n10420_, new_n10421_,
    new_n10422_, new_n10423_, new_n10424_, new_n10425_, new_n10426_,
    new_n10427_, new_n10428_, new_n10430_, new_n10431_, new_n10432_,
    new_n10433_, new_n10434_, new_n10435_, new_n10436_, new_n10437_,
    new_n10438_, new_n10439_, new_n10440_, new_n10441_, new_n10442_,
    new_n10444_, new_n10445_, new_n10447_, new_n10448_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10588_, new_n10589_, new_n10591_, new_n10592_,
    new_n10593_, new_n10594_, new_n10595_, new_n10596_, new_n10597_,
    new_n10598_, new_n10600_, new_n10601_, new_n10603_, new_n10604_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10628_, new_n10629_, new_n10630_, new_n10631_,
    new_n10632_, new_n10633_, new_n10634_, new_n10635_, new_n10636_,
    new_n10637_, new_n10638_, new_n10639_, new_n10640_, new_n10641_,
    new_n10642_, new_n10643_, new_n10644_, new_n10645_, new_n10646_,
    new_n10647_, new_n10648_, new_n10649_, new_n10650_, new_n10651_,
    new_n10652_, new_n10653_, new_n10654_, new_n10655_, new_n10656_,
    new_n10657_, new_n10658_, new_n10659_, new_n10660_, new_n10661_,
    new_n10662_, new_n10663_, new_n10664_, new_n10665_, new_n10666_,
    new_n10667_, new_n10668_, new_n10669_, new_n10670_, new_n10671_,
    new_n10672_, new_n10673_, new_n10674_, new_n10675_, new_n10676_,
    new_n10677_, new_n10678_, new_n10679_, new_n10680_, new_n10681_,
    new_n10682_, new_n10683_, new_n10684_, new_n10685_, new_n10686_,
    new_n10687_, new_n10688_, new_n10689_, new_n10690_, new_n10691_,
    new_n10692_, new_n10693_, new_n10694_, new_n10695_, new_n10696_,
    new_n10697_, new_n10698_, new_n10699_, new_n10700_, new_n10701_,
    new_n10702_, new_n10703_, new_n10704_, new_n10705_, new_n10706_,
    new_n10707_, new_n10708_, new_n10709_, new_n10710_, new_n10711_,
    new_n10712_, new_n10713_, new_n10714_, new_n10715_, new_n10716_,
    new_n10717_, new_n10718_, new_n10719_, new_n10720_, new_n10721_,
    new_n10722_, new_n10723_, new_n10724_, new_n10725_, new_n10726_,
    new_n10727_, new_n10728_, new_n10729_, new_n10731_, new_n10732_,
    new_n10733_, new_n10734_, new_n10735_, new_n10736_, new_n10737_,
    new_n10738_, new_n10739_, new_n10740_, new_n10741_, new_n10742_,
    new_n10743_, new_n10744_, new_n10745_, new_n10746_, new_n10747_,
    new_n10748_, new_n10749_, new_n10750_, new_n10751_, new_n10752_,
    new_n10753_, new_n10754_, new_n10755_, new_n10756_, new_n10757_,
    new_n10758_, new_n10759_, new_n10760_, new_n10761_, new_n10762_,
    new_n10763_, new_n10764_, new_n10765_, new_n10766_, new_n10767_,
    new_n10768_, new_n10769_, new_n10770_, new_n10771_, new_n10772_,
    new_n10773_, new_n10774_, new_n10775_, new_n10776_, new_n10777_,
    new_n10779_, new_n10780_, new_n10781_, new_n10782_, new_n10783_,
    new_n10784_, new_n10785_, new_n10786_, new_n10787_, new_n10789_,
    new_n10790_, new_n10792_, new_n10793_, new_n10795_, new_n10796_,
    new_n10797_, new_n10799_, new_n10800_, new_n10802_, new_n10803_,
    new_n10805_, new_n10806_, new_n10808_, new_n10809_, new_n10810_,
    new_n10811_, new_n10812_, new_n10814_, new_n10815_, new_n10816_,
    new_n10817_, new_n10818_, new_n10819_, new_n10820_, new_n10821_,
    new_n10822_, new_n10823_, new_n10825_, new_n10826_, new_n10828_,
    new_n10829_, new_n10830_, new_n10831_, new_n10832_, new_n10833_,
    new_n10834_, new_n10835_, new_n10836_, new_n10837_, new_n10838_,
    new_n10839_, new_n10841_, new_n10842_, new_n10843_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10857_, new_n10858_, new_n10860_, new_n10861_, new_n10863_,
    new_n10864_, new_n10866_, new_n10867_, new_n10869_, new_n10870_,
    new_n10872_, new_n10873_, new_n10875_, new_n10876_, new_n10877_,
    new_n10878_, new_n10879_, new_n10880_, new_n10881_, new_n10882_,
    new_n10883_, new_n10884_, new_n10886_, new_n10887_, new_n10888_,
    new_n10890_, new_n10891_, new_n10893_, new_n10894_, new_n10895_,
    new_n10897_, new_n10898_, new_n10900_, new_n10901_, new_n10903_,
    new_n10904_, new_n10906_, new_n10907_, new_n10909_, new_n10910_,
    new_n10912_, new_n10913_, new_n10914_, new_n10915_, new_n10916_,
    new_n10917_, new_n10918_, new_n10919_, new_n10920_, new_n10921_,
    new_n10922_, new_n10923_, new_n10924_, new_n10925_, new_n10926_,
    new_n10927_, new_n10928_, new_n10929_, new_n10930_, new_n10931_,
    new_n10932_, new_n10934_, new_n10935_, new_n10937_, new_n10938_,
    new_n10940_, new_n10941_, new_n10943_, new_n10944_, new_n10945_,
    new_n10947_, new_n10948_, new_n10949_, new_n10951_, new_n10952_,
    new_n10953_, new_n10954_, new_n10955_, new_n10956_, new_n10957_,
    new_n10959_, new_n10960_, new_n10962_, new_n10963_, new_n10965_,
    new_n10966_, new_n10968_, new_n10969_, new_n10971_, new_n10972_,
    new_n10973_, new_n10974_, new_n10975_, new_n10976_, new_n10977_,
    new_n10978_, new_n10979_, new_n10980_, new_n10981_, new_n10982_,
    new_n10983_, new_n10984_, new_n10985_, new_n10986_, new_n10987_,
    new_n10988_, new_n10989_, new_n10990_, new_n10991_, new_n10992_,
    new_n10993_, new_n10994_, new_n10995_, new_n10996_, new_n10997_,
    new_n10998_, new_n10999_, new_n11000_, new_n11001_, new_n11002_,
    new_n11003_, new_n11004_, new_n11005_, new_n11006_, new_n11007_,
    new_n11008_, new_n11009_, new_n11010_, new_n11011_, new_n11012_,
    new_n11014_, new_n11015_, new_n11016_, new_n11017_, new_n11018_,
    new_n11019_, new_n11020_, new_n11021_, new_n11022_, new_n11023_,
    new_n11024_, new_n11025_, new_n11026_, new_n11027_, new_n11028_,
    new_n11029_, new_n11030_, new_n11031_, new_n11032_, new_n11033_,
    new_n11034_, new_n11035_, new_n11036_, new_n11037_, new_n11038_,
    new_n11039_, new_n11040_, new_n11041_, new_n11042_, new_n11043_,
    new_n11044_, new_n11045_, new_n11046_, new_n11047_, new_n11048_,
    new_n11049_, new_n11050_, new_n11051_, new_n11052_, new_n11053_,
    new_n11054_, new_n11055_, new_n11056_, new_n11057_, new_n11058_,
    new_n11059_, new_n11060_, new_n11061_, new_n11062_, new_n11063_,
    new_n11064_, new_n11065_, new_n11066_, new_n11067_, new_n11068_,
    new_n11069_, new_n11070_, new_n11071_, new_n11072_, new_n11073_,
    new_n11074_, new_n11075_, new_n11076_, new_n11077_, new_n11078_,
    new_n11079_, new_n11080_, new_n11081_, new_n11082_, new_n11083_,
    new_n11084_, new_n11085_, new_n11086_, new_n11087_, new_n11088_,
    new_n11089_, new_n11090_, new_n11091_, new_n11092_, new_n11093_,
    new_n11094_, new_n11095_, new_n11096_, new_n11097_, new_n11098_,
    new_n11099_, new_n11100_, new_n11101_, new_n11102_, new_n11103_,
    new_n11104_, new_n11105_, new_n11106_, new_n11107_, new_n11108_,
    new_n11109_, new_n11110_, new_n11111_, new_n11112_, new_n11113_,
    new_n11114_, new_n11115_, new_n11116_, new_n11117_, new_n11118_,
    new_n11119_, new_n11120_, new_n11121_, new_n11122_, new_n11123_,
    new_n11124_, new_n11125_, new_n11126_, new_n11127_, new_n11128_,
    new_n11129_, new_n11130_, new_n11131_, new_n11132_, new_n11133_,
    new_n11134_, new_n11135_, new_n11136_, new_n11137_, new_n11138_,
    new_n11139_, new_n11140_, new_n11141_, new_n11142_, new_n11143_,
    new_n11144_, new_n11145_, new_n11146_, new_n11147_, new_n11148_,
    new_n11149_, new_n11151_, new_n11152_, new_n11153_, new_n11154_,
    new_n11155_, new_n11156_, new_n11157_, new_n11158_, new_n11159_,
    new_n11160_, new_n11161_, new_n11162_, new_n11163_, new_n11164_,
    new_n11165_, new_n11167_, new_n11168_, new_n11169_, new_n11171_,
    new_n11172_, new_n11174_, new_n11175_, new_n11177_, new_n11178_,
    new_n11179_, new_n11181_, new_n11182_, new_n11184_, new_n11185_,
    new_n11187_, new_n11188_, new_n11190_, new_n11191_, new_n11193_,
    new_n11194_, new_n11196_, new_n11197_, new_n11199_, new_n11200_,
    new_n11201_, new_n11203_, new_n11204_, new_n11205_, new_n11206_,
    new_n11207_, new_n11208_, new_n11209_, new_n11210_, new_n11211_,
    new_n11212_, new_n11213_, new_n11214_, new_n11215_, new_n11217_,
    new_n11218_, new_n11220_, new_n11221_, new_n11222_, new_n11223_,
    new_n11225_, new_n11226_, new_n11228_, new_n11229_, new_n11231_,
    new_n11232_, new_n11234_, new_n11235_, new_n11236_, new_n11238_,
    new_n11239_, new_n11240_, new_n11241_, new_n11242_, new_n11243_,
    new_n11244_, new_n11245_, new_n11246_, new_n11248_, new_n11249_,
    new_n11251_, new_n11252_, new_n11254_, new_n11255_, new_n11257_,
    new_n11258_, new_n11259_, new_n11261_, new_n11262_, new_n11264_,
    new_n11265_, new_n11267_, new_n11268_, new_n11270_, new_n11271_,
    new_n11273_, new_n11274_, new_n11276_, new_n11277_, new_n11278_,
    new_n11279_, new_n11280_, new_n11281_, new_n11282_, new_n11283_,
    new_n11284_, new_n11285_, new_n11286_, new_n11288_, new_n11289_,
    new_n11290_, new_n11291_, new_n11292_, new_n11293_, new_n11294_,
    new_n11295_, new_n11296_, new_n11297_, new_n11299_, new_n11300_,
    new_n11302_, new_n11303_, new_n11305_, new_n11306_, new_n11308_,
    new_n11309_, new_n11311_, new_n11312_, new_n11314_, new_n11315_,
    new_n11316_, new_n11317_, new_n11318_, new_n11319_, new_n11320_,
    new_n11321_, new_n11322_, new_n11323_, new_n11324_, new_n11326_,
    new_n11327_, new_n11329_, new_n11330_, new_n11331_, new_n11332_,
    new_n11333_, new_n11334_, new_n11336_, new_n11337_, new_n11338_,
    new_n11339_, new_n11341_, new_n11342_, new_n11344_, new_n11345_,
    new_n11346_, new_n11347_, new_n11349_, new_n11350_, new_n11352_,
    new_n11353_, new_n11354_, new_n11355_, new_n11356_, new_n11357_,
    new_n11358_, new_n11359_, new_n11360_, new_n11361_, new_n11363_,
    new_n11364_, new_n11366_, new_n11367_, new_n11369_, new_n11370_,
    new_n11372_, new_n11373_, new_n11374_, new_n11376_, new_n11377_,
    new_n11378_, new_n11379_, new_n11380_, new_n11381_, new_n11382_,
    new_n11383_, new_n11384_, new_n11385_, new_n11386_, new_n11387_,
    new_n11388_, new_n11389_, new_n11390_, new_n11391_, new_n11393_,
    new_n11394_, new_n11395_, new_n11396_, new_n11397_, new_n11398_,
    new_n11399_, new_n11400_, new_n11401_, new_n11402_, new_n11403_,
    new_n11404_, new_n11405_, new_n11406_, new_n11407_, new_n11409_,
    new_n11410_, new_n11411_, new_n11412_, new_n11413_, new_n11414_,
    new_n11415_, new_n11416_, new_n11417_, new_n11418_, new_n11419_,
    new_n11420_, new_n11422_, new_n11423_, new_n11424_, new_n11426_,
    new_n11427_, new_n11429_, new_n11430_, new_n11432_, new_n11433_,
    new_n11434_, new_n11435_, new_n11436_, new_n11437_, new_n11438_,
    new_n11439_, new_n11440_, new_n11441_, new_n11442_, new_n11443_,
    new_n11444_, new_n11445_, new_n11446_, new_n11447_, new_n11448_,
    new_n11449_, new_n11450_, new_n11451_, new_n11452_, new_n11453_,
    new_n11454_, new_n11455_, new_n11456_, new_n11457_, new_n11458_,
    new_n11459_, new_n11460_, new_n11461_, new_n11462_, new_n11463_,
    new_n11465_, new_n11466_, new_n11467_, new_n11469_, new_n11470_,
    new_n11472_, new_n11473_, new_n11475_, new_n11476_, new_n11478_,
    new_n11479_, new_n11481_, new_n11482_, new_n11484_, new_n11485_,
    new_n11487_, new_n11488_, new_n11489_, new_n11491_, new_n11492_,
    new_n11493_, new_n11495_, new_n11496_, new_n11498_, new_n11499_,
    new_n11501_, new_n11502_, new_n11504_, new_n11505_, new_n11507_,
    new_n11508_, new_n11509_, new_n11511_, new_n11512_, new_n11514_,
    new_n11515_, new_n11517_, new_n11518_, new_n11519_, new_n11521_,
    new_n11522_, new_n11524_, new_n11525_, new_n11527_, new_n11528_,
    new_n11530_, new_n11531_, new_n11532_, new_n11534_, new_n11535_,
    new_n11537_, new_n11538_, new_n11540_, new_n11541_, new_n11543_,
    new_n11544_, new_n11546_, new_n11547_, new_n11549_, new_n11550_,
    new_n11552_, new_n11553_, new_n11555_, new_n11556_, new_n11558_,
    new_n11559_, new_n11561_, new_n11562_, new_n11564_, new_n11565_,
    new_n11567_, new_n11568_, new_n11570_, new_n11571_, new_n11573_,
    new_n11574_, new_n11576_, new_n11577_, new_n11578_, new_n11579_,
    new_n11580_, new_n11581_, new_n11582_, new_n11583_, new_n11584_,
    new_n11585_, new_n11586_, new_n11587_, new_n11588_, new_n11589_,
    new_n11590_, new_n11591_, new_n11592_, new_n11593_, new_n11594_,
    new_n11595_, new_n11596_, new_n11597_, new_n11598_, new_n11599_,
    new_n11600_, new_n11601_, new_n11602_, new_n11603_, new_n11604_,
    new_n11605_, new_n11606_, new_n11607_, new_n11608_, new_n11609_,
    new_n11610_, new_n11611_, new_n11612_, new_n11613_, new_n11614_,
    new_n11615_, new_n11616_, new_n11617_, new_n11618_, new_n11619_,
    new_n11620_, new_n11621_, new_n11622_, new_n11623_, new_n11624_,
    new_n11625_, new_n11626_, new_n11627_, new_n11628_, new_n11630_,
    new_n11631_, new_n11633_, new_n11634_, new_n11636_, new_n11637_,
    new_n11639_, new_n11640_, new_n11641_, new_n11642_, new_n11643_,
    new_n11644_, new_n11646_, new_n11647_, new_n11648_, new_n11649_,
    new_n11651_, new_n11652_, new_n11654_, new_n11655_, new_n11657_,
    new_n11658_, new_n11660_, new_n11661_, new_n11662_, new_n11663_,
    new_n11664_, new_n11665_, new_n11666_, new_n11667_, new_n11669_,
    new_n11670_, new_n11671_, new_n11672_, new_n11673_, new_n11674_,
    new_n11675_, new_n11676_, new_n11677_, new_n11678_, new_n11679_,
    new_n11680_, new_n11682_, new_n11683_, new_n11684_, new_n11685_,
    new_n11686_, new_n11687_, new_n11688_, new_n11689_, new_n11690_,
    new_n11691_, new_n11692_, new_n11693_, new_n11695_, new_n11696_,
    new_n11697_, new_n11698_, new_n11699_, new_n11701_, new_n11702_,
    new_n11704_, new_n11705_, new_n11708_, new_n11709_, new_n11711_,
    new_n11712_, new_n11714_, new_n11715_, new_n11717_, new_n11718_,
    new_n11720_, new_n11721_, new_n11723_, new_n11724_, new_n11726_,
    new_n11727_, new_n11729_, new_n11730_, new_n11731_, new_n11732_,
    new_n11733_, new_n11734_, new_n11735_, new_n11736_, new_n11737_,
    new_n11738_, new_n11739_, new_n11741_, new_n11742_, new_n11744_,
    new_n11745_, new_n11746_, new_n11748_, new_n11749_, new_n11751_,
    new_n11752_, new_n11753_, new_n11754_, new_n11755_, new_n11756_,
    new_n11757_, new_n11758_, new_n11759_, new_n11760_, new_n11761_,
    new_n11763_, new_n11764_, new_n11766_, new_n11767_, new_n11768_,
    new_n11770_, new_n11771_, new_n11773_, new_n11774_, new_n11776_,
    new_n11777_, new_n11778_, new_n11779_, new_n11781_, new_n11782_,
    new_n11784_, new_n11785_, new_n11786_, new_n11787_, new_n11788_,
    new_n11789_, new_n11790_, new_n11791_, new_n11792_, new_n11793_,
    new_n11795_, new_n11796_, new_n11797_, new_n11798_, new_n11800_,
    new_n11801_, new_n11803_, new_n11804_, new_n11806_, new_n11807_,
    new_n11808_, new_n11810_, new_n11811_, new_n11813_, new_n11814_,
    new_n11816_, new_n11817_, new_n11819_, new_n11820_, new_n11821_,
    new_n11822_, new_n11823_, new_n11824_, new_n11825_, new_n11826_,
    new_n11827_, new_n11828_, new_n11829_, new_n11831_, new_n11832_,
    new_n11834_, new_n11835_, new_n11836_, new_n11838_, new_n11839_,
    new_n11840_, new_n11841_, new_n11842_, new_n11843_, new_n11844_,
    new_n11845_, new_n11846_, new_n11847_, new_n11848_, new_n11849_,
    new_n11850_, new_n11851_, new_n11852_, new_n11853_, new_n11854_,
    new_n11855_, new_n11856_, new_n11858_, new_n11859_, new_n11861_,
    new_n11862_, new_n11863_, new_n11864_, new_n11865_, new_n11866_,
    new_n11867_, new_n11868_, new_n11869_, new_n11870_, new_n11871_,
    new_n11872_, new_n11873_, new_n11874_, new_n11875_, new_n11876_,
    new_n11877_, new_n11878_, new_n11879_, new_n11881_, new_n11882_,
    new_n11883_, new_n11885_, new_n11886_, new_n11887_, new_n11888_,
    new_n11889_, new_n11890_, new_n11891_, new_n11892_, new_n11893_,
    new_n11894_, new_n11895_, new_n11896_, new_n11897_, new_n11898_,
    new_n11899_, new_n11900_, new_n11901_, new_n11902_, new_n11903_,
    new_n11904_, new_n11905_, new_n11907_, new_n11909_, new_n11910_,
    new_n11912_, new_n11913_, new_n11914_, new_n11915_, new_n11917_,
    new_n11918_, new_n11920_, new_n11922_, new_n11923_, new_n11925_,
    new_n11926_, new_n11928_, new_n11929_, new_n11931_, new_n11932_,
    new_n11934_, new_n11935_, new_n11937_, new_n11938_, new_n11939_,
    new_n11940_, new_n11941_, new_n11942_, new_n11943_, new_n11944_,
    new_n11945_, new_n11946_, new_n11948_, new_n11949_, new_n11951_,
    new_n11952_, new_n11953_, new_n11954_, new_n11955_, new_n11956_,
    new_n11957_, new_n11958_, new_n11959_, new_n11960_, new_n11962_,
    new_n11963_, new_n11965_, new_n11966_, new_n11968_, new_n11969_,
    new_n11971_, new_n11972_, new_n11973_, new_n11975_, new_n11976_,
    new_n11978_, new_n11979_, new_n11980_, new_n11981_, new_n11982_,
    new_n11983_, new_n11984_, new_n11985_, new_n11986_, new_n11987_,
    new_n11988_, new_n11989_, new_n11990_, new_n11991_, new_n11992_,
    new_n11993_, new_n11994_, new_n11995_, new_n11996_, new_n11997_,
    new_n11998_, new_n11999_, new_n12000_, new_n12001_, new_n12002_,
    new_n12003_, new_n12005_, new_n12006_, new_n12008_, new_n12009_,
    new_n12011_, new_n12012_, new_n12013_, new_n12014_, new_n12016_,
    new_n12017_, new_n12018_, new_n12020_, new_n12021_, new_n12023_,
    new_n12024_, new_n12025_, new_n12027_, new_n12028_, new_n12030_,
    new_n12031_, new_n12033_, new_n12034_, new_n12037_, new_n12038_,
    new_n12039_, new_n12040_, new_n12041_, new_n12043_, new_n12044_,
    new_n12045_, new_n12046_, new_n12047_, new_n12048_, new_n12049_,
    new_n12050_, new_n12051_, new_n12052_, new_n12053_, new_n12054_,
    new_n12055_, new_n12056_, new_n12058_, new_n12059_, new_n12060_,
    new_n12061_, new_n12062_, new_n12063_, new_n12064_, new_n12065_,
    new_n12066_, new_n12067_, new_n12068_, new_n12069_, new_n12070_,
    new_n12071_, new_n12072_, new_n12073_, new_n12074_, new_n12075_,
    new_n12076_, new_n12077_, new_n12078_, new_n12080_, new_n12081_,
    new_n12082_, new_n12083_, new_n12084_, new_n12085_, new_n12086_,
    new_n12087_, new_n12088_, new_n12090_, new_n12091_, new_n12093_,
    new_n12094_, new_n12097_, new_n12098_, new_n12100_, new_n12101_,
    new_n12103_, new_n12104_, new_n12106_, new_n12107_, new_n12109_,
    new_n12110_, new_n12112_, new_n12113_, new_n12115_, new_n12116_,
    new_n12118_, new_n12119_, new_n12121_, new_n12122_, new_n12124_,
    new_n12125_, new_n12126_, new_n12128_, new_n12129_, new_n12130_,
    new_n12131_, new_n12132_, new_n12133_, new_n12134_, new_n12135_,
    new_n12136_, new_n12137_, new_n12138_, new_n12139_, new_n12140_,
    new_n12141_, new_n12142_, new_n12143_, new_n12144_, new_n12145_,
    new_n12146_, new_n12148_, new_n12149_, new_n12151_, new_n12152_,
    new_n12154_, new_n12155_, new_n12157_, new_n12158_, new_n12160_,
    new_n12161_, new_n12163_, new_n12164_, new_n12166_, new_n12167_,
    new_n12169_, new_n12170_, new_n12171_, new_n12172_, new_n12174_,
    new_n12175_, new_n12177_, new_n12178_, new_n12180_, new_n12181_,
    new_n12183_, new_n12184_, new_n12186_, new_n12187_, new_n12189_,
    new_n12190_, new_n12192_, new_n12193_, new_n12195_, new_n12196_,
    new_n12198_, new_n12199_, new_n12200_, new_n12202_, new_n12203_,
    new_n12205_, new_n12206_, new_n12207_, new_n12208_, new_n12209_,
    new_n12210_, new_n12211_, new_n12212_, new_n12213_, new_n12214_,
    new_n12215_, new_n12217_, new_n12218_, new_n12220_, new_n12221_,
    new_n12222_, new_n12224_, new_n12225_, new_n12227_, new_n12228_,
    new_n12230_, new_n12231_, new_n12233_, new_n12234_, new_n12236_,
    new_n12237_, new_n12239_, new_n12240_, new_n12242_, new_n12243_,
    new_n12245_, new_n12246_, new_n12248_, new_n12249_, new_n12251_,
    new_n12252_, new_n12254_, new_n12255_, new_n12257_, new_n12258_,
    new_n12260_, new_n12261_, new_n12263_, new_n12264_, new_n12266_,
    new_n12267_, new_n12269_, new_n12270_, new_n12271_, new_n12272_,
    new_n12273_, new_n12274_, new_n12275_, new_n12276_, new_n12278_,
    new_n12279_, new_n12281_, new_n12282_, new_n12284_, new_n12285_,
    new_n12287_, new_n12288_, new_n12290_, new_n12291_, new_n12293_,
    new_n12294_, new_n12295_, new_n12297_, new_n12298_, new_n12299_,
    new_n12301_, new_n12302_, new_n12304_, new_n12305_, new_n12307_,
    new_n12308_, new_n12310_, new_n12311_, new_n12313_, new_n12314_,
    new_n12315_, new_n12316_, new_n12317_, new_n12319_, new_n12320_,
    new_n12321_, new_n12322_, new_n12323_, new_n12324_, new_n12325_,
    new_n12326_, new_n12327_, new_n12328_, new_n12329_, new_n12330_,
    new_n12332_, new_n12333_, new_n12334_, new_n12335_, new_n12336_,
    new_n12337_, new_n12338_, new_n12339_, new_n12340_, new_n12341_,
    new_n12342_, new_n12343_, new_n12344_, new_n12345_, new_n12346_,
    new_n12347_, new_n12348_, new_n12349_, new_n12350_, new_n12351_,
    new_n12352_, new_n12354_, new_n12355_, new_n12356_, new_n12358_,
    new_n12359_, new_n12361_, new_n12362_, new_n12363_, new_n12366_,
    new_n12367_, new_n12369_, new_n12370_, new_n12372_, new_n12373_,
    new_n12375_, new_n12376_, new_n12378_, new_n12379_, new_n12381_,
    new_n12382_, new_n12384_, new_n12385_, new_n12387_, new_n12388_,
    new_n12390_, new_n12391_, new_n12393_, new_n12394_, new_n12396_,
    new_n12397_, new_n12399_, new_n12400_, new_n12401_, new_n12403_,
    new_n12404_, new_n12406_, new_n12407_, new_n12409_, new_n12410_,
    new_n12412_, new_n12413_, new_n12415_, new_n12416_, new_n12418_,
    new_n12419_, new_n12421_, new_n12422_, new_n12423_, new_n12424_,
    new_n12426_, new_n12427_, new_n12429_, new_n12430_, new_n12432_,
    new_n12433_, new_n12435_, new_n12436_, new_n12438_, new_n12439_,
    new_n12441_, new_n12442_, new_n12444_, new_n12445_, new_n12447_,
    new_n12448_, new_n12450_, new_n12451_, new_n12453_, new_n12454_,
    new_n12456_, new_n12457_, new_n12459_, new_n12460_, new_n12462_,
    new_n12463_, new_n12465_, new_n12466_, new_n12467_, new_n12469_,
    new_n12470_, new_n12472_, new_n12473_, new_n12475_, new_n12476_,
    new_n12478_, new_n12479_, new_n12481_, new_n12482_, new_n12483_,
    new_n12485_, new_n12486_, new_n12487_, new_n12488_, new_n12490_,
    new_n12491_, new_n12493_, new_n12494_, new_n12496_, new_n12497_,
    new_n12499_, new_n12500_, new_n12502_, new_n12503_, new_n12505_,
    new_n12506_, new_n12508_, new_n12509_, new_n12511_, new_n12512_,
    new_n12514_, new_n12515_, new_n12516_, new_n12517_, new_n12518_,
    new_n12519_, new_n12520_, new_n12521_, new_n12522_, new_n12523_,
    new_n12524_, new_n12525_, new_n12526_, new_n12527_, new_n12528_,
    new_n12529_, new_n12530_, new_n12531_, new_n12532_, new_n12533_,
    new_n12534_, new_n12535_, new_n12536_, new_n12537_, new_n12538_,
    new_n12539_, new_n12540_, new_n12541_, new_n12542_, new_n12543_,
    new_n12544_, new_n12545_, new_n12546_, new_n12547_, new_n12548_,
    new_n12549_, new_n12550_, new_n12551_, new_n12552_, new_n12553_,
    new_n12554_, new_n12555_, new_n12556_, new_n12557_, new_n12558_,
    new_n12559_, new_n12560_, new_n12561_, new_n12562_, new_n12563_,
    new_n12564_, new_n12565_, new_n12566_, new_n12568_, new_n12569_,
    new_n12571_, new_n12572_, new_n12574_, new_n12575_, new_n12577_,
    new_n12578_, new_n12580_, new_n12581_, new_n12583_, new_n12584_,
    new_n12586_, new_n12587_, new_n12589_, new_n12590_, new_n12591_,
    new_n12593_, new_n12594_, new_n12595_, new_n12597_, new_n12598_,
    new_n12600_, new_n12601_, new_n12603_, new_n12604_, new_n12606_,
    new_n12607_, new_n12610_, new_n12611_, new_n12612_, new_n12613_,
    new_n12614_, new_n12615_, new_n12616_, new_n12618_, new_n12619_,
    new_n12620_, new_n12621_, new_n12622_, new_n12623_, new_n12624_,
    new_n12625_, new_n12626_, new_n12627_, new_n12628_, new_n12629_,
    new_n12630_, new_n12631_, new_n12632_, new_n12633_, new_n12634_,
    new_n12635_, new_n12636_, new_n12637_, new_n12638_, new_n12640_,
    new_n12641_, new_n12642_, new_n12643_, new_n12644_, new_n12645_,
    new_n12646_, new_n12647_, new_n12648_, new_n12649_, new_n12650_,
    new_n12651_, new_n12652_, new_n12653_, new_n12655_, new_n12656_,
    new_n12657_, new_n12658_, new_n12659_, new_n12661_, new_n12662_,
    new_n12663_, new_n12664_, new_n12665_, new_n12666_, new_n12667_,
    new_n12668_, new_n12669_, new_n12670_, new_n12671_, new_n12672_,
    new_n12673_, new_n12674_, new_n12675_, new_n12676_, new_n12677_,
    new_n12678_, new_n12679_, new_n12680_, new_n12681_, new_n12682_,
    new_n12683_, new_n12684_, new_n12685_, new_n12686_, new_n12687_,
    new_n12688_, new_n12689_, new_n12690_, new_n12691_, new_n12693_,
    new_n12694_, new_n12696_, new_n12697_, new_n12698_, new_n12700_,
    new_n12701_, new_n12703_, new_n12704_, new_n12706_, new_n12707_,
    new_n12709_, new_n12710_, new_n12712_, new_n12713_, new_n12715_,
    new_n12716_, new_n12718_, new_n12719_, new_n12720_, new_n12722_,
    new_n12723_, new_n12725_, new_n12726_, new_n12728_, new_n12729_,
    new_n12731_, new_n12732_, new_n12734_, new_n12735_, new_n12737_,
    new_n12738_, new_n12740_, new_n12741_, new_n12743_, new_n12744_,
    new_n12746_, new_n12747_, new_n12749_, new_n12750_, new_n12752_,
    new_n12753_, new_n12755_, new_n12756_, new_n12758_, new_n12759_,
    new_n12761_, new_n12762_, new_n12764_, new_n12765_, new_n12767_,
    new_n12768_, new_n12770_, new_n12771_, new_n12773_, new_n12774_,
    new_n12776_, new_n12777_, new_n12779_, new_n12780_, new_n12782_,
    new_n12783_, new_n12784_, new_n12786_, new_n12787_, new_n12788_,
    new_n12789_, new_n12791_, new_n12792_, new_n12794_, new_n12795_,
    new_n12797_, new_n12798_, new_n12800_, new_n12801_, new_n12803_,
    new_n12804_, new_n12806_, new_n12807_, new_n12808_, new_n12810_,
    new_n12811_, new_n12812_, new_n12813_, new_n12815_, new_n12816_,
    new_n12818_, new_n12819_, new_n12821_, new_n12822_, new_n12824_,
    new_n12825_, new_n12827_, new_n12828_, new_n12830_, new_n12831_,
    new_n12833_, new_n12834_, new_n12836_, new_n12837_, new_n12838_,
    new_n12840_, new_n12841_, new_n12843_, new_n12844_, new_n12846_,
    new_n12847_, new_n12849_, new_n12850_, new_n12852_, new_n12853_,
    new_n12855_, new_n12857_, new_n12858_, new_n12859_, new_n12861_,
    new_n12862_, new_n12864_, new_n12865_, new_n12867_, new_n12868_,
    new_n12870_, new_n12871_, new_n12874_, new_n12875_, new_n12876_,
    new_n12877_, new_n12878_, new_n12880_, new_n12881_, new_n12882_,
    new_n12883_, new_n12884_, new_n12885_, new_n12886_, new_n12887_,
    new_n12888_, new_n12889_, new_n12890_, new_n12891_, new_n12893_,
    new_n12894_, new_n12895_, new_n12896_, new_n12897_, new_n12898_,
    new_n12899_, new_n12900_, new_n12901_, new_n12902_, new_n12903_,
    new_n12904_, new_n12906_, new_n12907_, new_n12908_, new_n12910_,
    new_n12911_, new_n12913_, new_n12914_, new_n12915_, new_n12917_,
    new_n12918_, new_n12920_, new_n12921_, new_n12923_, new_n12924_,
    new_n12926_, new_n12927_, new_n12929_, new_n12930_, new_n12931_,
    new_n12932_, new_n12933_, new_n12934_, new_n12935_, new_n12937_,
    new_n12938_, new_n12939_, new_n12940_, new_n12941_, new_n12942_,
    new_n12943_, new_n12944_, new_n12945_, new_n12946_, new_n12947_,
    new_n12948_, new_n12949_, new_n12950_, new_n12951_, new_n12952_,
    new_n12953_, new_n12954_, new_n12955_, new_n12956_, new_n12957_,
    new_n12958_, new_n12959_, new_n12960_, new_n12961_, new_n12962_,
    new_n12963_, new_n12964_, new_n12965_, new_n12966_, new_n12967_,
    new_n12968_, new_n12969_, new_n12970_, new_n12971_, new_n12972_,
    new_n12973_, new_n12974_, new_n12975_, new_n12976_, new_n12977_,
    new_n12978_, new_n12979_, new_n12980_, new_n12981_, new_n12982_,
    new_n12983_, new_n12984_, new_n12985_, new_n12986_, new_n12987_,
    new_n12988_, new_n12989_, new_n12990_, new_n12991_, new_n12992_,
    new_n12994_, new_n12995_, new_n12997_, new_n12998_, new_n13000_,
    new_n13001_, new_n13003_, new_n13004_, new_n13005_, new_n13006_,
    new_n13007_, new_n13008_, new_n13009_, new_n13011_, new_n13012_,
    new_n13013_, new_n13014_, new_n13015_, new_n13016_, new_n13017_,
    new_n13019_, new_n13020_, new_n13021_, new_n13022_, new_n13023_,
    new_n13024_, new_n13025_, new_n13026_, new_n13027_, new_n13028_,
    new_n13029_, new_n13030_, new_n13031_, new_n13032_, new_n13033_,
    new_n13034_, new_n13035_, new_n13036_, new_n13037_, new_n13038_,
    new_n13039_, new_n13040_, new_n13041_, new_n13042_, new_n13043_,
    new_n13044_, new_n13045_, new_n13046_, new_n13047_, new_n13048_,
    new_n13049_, new_n13050_, new_n13051_, new_n13052_, new_n13053_,
    new_n13055_, new_n13056_, new_n13057_, new_n13058_, new_n13059_,
    new_n13060_, new_n13061_, new_n13062_, new_n13063_, new_n13064_,
    new_n13065_, new_n13066_, new_n13067_, new_n13068_, new_n13069_,
    new_n13070_, new_n13071_, new_n13072_, new_n13073_, new_n13074_,
    new_n13075_, new_n13076_, new_n13077_, new_n13078_, new_n13079_,
    new_n13080_, new_n13081_, new_n13082_, new_n13083_, new_n13084_,
    new_n13085_, new_n13086_, new_n13087_, new_n13088_, new_n13090_,
    new_n13091_, new_n13093_, new_n13094_, new_n13095_, new_n13096_,
    new_n13097_, new_n13098_, new_n13099_, new_n13100_, new_n13101_,
    new_n13102_, new_n13103_, new_n13104_, new_n13105_, new_n13106_,
    new_n13107_, new_n13108_, new_n13109_, new_n13110_, new_n13111_,
    new_n13112_, new_n13113_, new_n13114_, new_n13115_, new_n13116_,
    new_n13117_, new_n13118_, new_n13119_, new_n13120_, new_n13121_,
    new_n13122_, new_n13123_, new_n13124_, new_n13125_, new_n13126_,
    new_n13127_, new_n13128_, new_n13129_, new_n13130_, new_n13131_,
    new_n13132_, new_n13133_, new_n13134_, new_n13136_, new_n13137_,
    new_n13138_, new_n13139_, new_n13140_, new_n13142_, new_n13143_,
    new_n13145_, new_n13146_, new_n13148_, new_n13149_, new_n13151_,
    new_n13152_, new_n13153_, new_n13154_, new_n13155_, new_n13157_,
    new_n13158_, new_n13159_, new_n13161_, new_n13162_, new_n13163_,
    new_n13164_, new_n13166_, new_n13167_, new_n13169_, new_n13170_,
    new_n13172_, new_n13173_, new_n13175_, new_n13176_, new_n13178_,
    new_n13179_, new_n13181_, new_n13182_, new_n13184_, new_n13185_,
    new_n13187_, new_n13188_, new_n13189_, new_n13190_, new_n13191_,
    new_n13192_, new_n13193_, new_n13194_, new_n13196_, new_n13197_,
    new_n13199_, new_n13200_, new_n13202_, new_n13203_, new_n13205_,
    new_n13206_, new_n13208_, new_n13209_, new_n13211_, new_n13212_,
    new_n13214_, new_n13215_, new_n13217_, new_n13218_, new_n13219_,
    new_n13220_, new_n13222_, new_n13223_, new_n13225_, new_n13226_,
    new_n13228_, new_n13229_, new_n13231_, new_n13232_, new_n13234_,
    new_n13235_, new_n13237_, new_n13238_, new_n13239_, new_n13241_,
    new_n13242_, new_n13243_, new_n13244_, new_n13246_, new_n13247_,
    new_n13249_, new_n13250_, new_n13251_, new_n13253_, new_n13255_,
    new_n13256_, new_n13258_, new_n13259_, new_n13261_, new_n13262_,
    new_n13263_, new_n13265_, new_n13266_, new_n13267_, new_n13268_,
    new_n13270_, new_n13271_, new_n13273_, new_n13274_, new_n13276_,
    new_n13277_, new_n13279_, new_n13280_, new_n13282_, new_n13283_,
    new_n13285_, new_n13286_, new_n13288_, new_n13289_, new_n13291_,
    new_n13292_, new_n13293_, new_n13295_, new_n13296_, new_n13298_,
    new_n13299_, new_n13300_, new_n13302_, new_n13303_, new_n13305_,
    new_n13306_, new_n13308_, new_n13309_, new_n13311_, new_n13312_,
    new_n13314_, new_n13315_, new_n13317_, new_n13318_, new_n13320_,
    new_n13321_, new_n13323_, new_n13324_, new_n13325_, new_n13326_,
    new_n13327_, new_n13328_, new_n13329_, new_n13330_, new_n13331_,
    new_n13332_, new_n13333_, new_n13334_, new_n13335_, new_n13336_,
    new_n13337_, new_n13338_, new_n13339_, new_n13340_, new_n13341_,
    new_n13342_, new_n13343_, new_n13344_, new_n13345_, new_n13346_,
    new_n13347_, new_n13348_, new_n13349_, new_n13350_, new_n13351_,
    new_n13352_, new_n13353_, new_n13354_, new_n13355_, new_n13356_,
    new_n13357_, new_n13358_, new_n13359_, new_n13360_, new_n13361_,
    new_n13362_, new_n13363_, new_n13364_, new_n13365_, new_n13366_,
    new_n13367_, new_n13368_, new_n13369_, new_n13370_, new_n13371_,
    new_n13372_, new_n13373_, new_n13374_, new_n13375_, new_n13376_,
    new_n13377_, new_n13378_, new_n13379_, new_n13380_, new_n13382_,
    new_n13383_, new_n13384_, new_n13386_, new_n13387_, new_n13389_,
    new_n13390_, new_n13392_, new_n13393_, new_n13395_, new_n13396_,
    new_n13398_, new_n13399_, new_n13400_, new_n13401_, new_n13403_,
    new_n13404_, new_n13406_, new_n13407_, new_n13409_, new_n13410_,
    new_n13412_, new_n13413_, new_n13415_, new_n13416_, new_n13417_,
    new_n13419_, new_n13420_, new_n13422_, new_n13423_, new_n13425_,
    new_n13426_, new_n13428_, new_n13429_, new_n13431_, new_n13432_,
    new_n13434_, new_n13435_, new_n13437_, new_n13438_, new_n13440_,
    new_n13441_, new_n13443_, new_n13444_, new_n13446_, new_n13447_,
    new_n13449_, new_n13450_, new_n13452_, new_n13453_, new_n13455_,
    new_n13456_, new_n13458_, new_n13459_, new_n13460_, new_n13462_,
    new_n13463_, new_n13465_, new_n13466_, new_n13467_, new_n13468_,
    new_n13469_, new_n13470_, new_n13471_, new_n13472_, new_n13473_,
    new_n13474_, new_n13476_, new_n13477_, new_n13479_, new_n13480_,
    new_n13482_, new_n13483_, new_n13484_, new_n13485_, new_n13486_,
    new_n13487_, new_n13488_, new_n13490_, new_n13491_, new_n13493_,
    new_n13495_, new_n13496_, new_n13498_, new_n13499_, new_n13501_,
    new_n13502_, new_n13504_, new_n13505_, new_n13507_, new_n13508_,
    new_n13510_, new_n13511_, new_n13513_, new_n13514_, new_n13516_,
    new_n13518_, new_n13519_, new_n13520_, new_n13522_, new_n13523_,
    new_n13525_, new_n13526_, new_n13528_, new_n13529_, new_n13531_,
    new_n13532_, new_n13534_, new_n13535_, new_n13537_, new_n13538_,
    new_n13540_, new_n13541_, new_n13543_, new_n13544_, new_n13546_,
    new_n13547_, new_n13548_, new_n13550_, new_n13551_, new_n13553_,
    new_n13554_, new_n13556_, new_n13557_, new_n13559_, new_n13560_,
    new_n13562_, new_n13563_, new_n13565_, new_n13566_, new_n13568_,
    new_n13569_, new_n13571_, new_n13572_, new_n13573_, new_n13575_,
    new_n13576_, n272, n277, n282, n287, n292, n297, n302, n307, n312,
    n317, n322, n327, n332, n337, n342, n347, n352, n357, n362, n367, n372,
    n377, n382, n387, n392, n397, n402, n407, n412, n417, n422, n427, n432,
    n437, n442, n447, n452, n457, n462, n467, n472, n477, n482, n487, n492,
    n497, n502, n507, n512, n517, n522, n527, n532, n537, n542, n547, n552,
    n557, n562, n567, n572, n577, n582, n587, n592, n597, n602, n607, n612,
    n617, n622, n627, n632, n637, n642, n647, n652, n657, n662, n667, n672,
    n677, n682, n687, n692, n697, n702, n707, n712, n717, n722, n727, n732,
    n737, n742, n747, n752, n757, n762, n767, n772, n777, n782, n787, n792,
    n797, n802, n807, n812, n817, n822, n826, n831, n835, n840, n844, n849,
    n854, n859, n864, n869, n874, n879, n884, n889, n894, n899, n904, n909,
    n914, n919, n924, n929, n934, n939, n944, n948, n953, n958, n962, n967,
    n971, n976, n981, n986, n991, n996, n1000, n1005, n1010, n1015, n1020,
    n1025, n1030, n1035, n1040, n1045, n1050, n1055, n1060, n1065, n1070,
    n1074, n1079, n1083, n1088, n1092, n1097, n1102, n1107, n1112, n1117,
    n1122, n1127, n1132, n1137, n1142, n1147, n1152, n1157, n1162, n1167,
    n1172, n1177, n1182, n1185, n1190, n1194, n1199, n1203, n1208, n1213,
    n1218, n1223, n1228, n1233, n1238, n1243, n1248, n1253, n1258, n1263,
    n1268, n1273, n1278, n1283, n1288, n1293, n1298, n1303, n1308, n1313,
    n1318, n1323, n1328, n1333, n1338, n1343, n1348, n1353, n1358, n1363,
    n1368, n1373, n1378, n1383, n1388, n1393, n1398, n1403, n1408, n1413,
    n1418, n1423, n1428, n1433, n1438, n1443, n1448, n1453, n1458, n1463,
    n1468, n1473, n1478, n1483, n1488, n1493, n1498, n1503, n1508, n1513,
    n1518, n1523, n1528, n1533, n1537, n1542, n1547, n1552, n1556, n1561,
    n1566, n1571, n1576, n1581, n1586, n1591, n1596, n1601, n1606, n1611,
    n1616, n1621, n1626, n1631, n1636, n1641, n1646, n1651, n1656, n1661,
    n1666, n1671, n1676, n1681, n1686, n1691, n1696, n1701, n1706, n1711,
    n1716, n1721, n1726, n1731, n1736, n1741, n1746, n1751, n1755, n1760,
    n1763, n1768, n1772, n1777, n1781, n1786, n1791, n1796, n1801, n1806,
    n1811, n1816, n1821, n1826, n1831, n1836, n1841, n1846, n1851, n1856,
    n1861, n1866, n1871, n1876, n1880, n1885, n1889, n1894, n1899, n1904,
    n1908, n1913, n1918, n1923, n1927, n1932, n1937, n1942, n1947, n1952,
    n1957, n1962, n1967, n1972, n1977, n1982, n1987, n1990, n1995, n1999,
    n2004, n2009, n2014, n2019, n2024, n2029, n2034, n2039, n2044, n2049,
    n2054, n2059, n2064, n2069, n2074, n2079, n2084, n2089, n2094, n2098,
    n2103, n2107, n2112, n2116, n2121, n2126, n2131, n2136, n2141, n2146,
    n2151, n2156, n2161, n2166, n2171, n2176, n2181, n2186, n2191, n2196,
    n2201, n2206, n2211, n2216, n2221, n2226, n2231, n2236, n2241, n2246,
    n2251, n2256, n2261, n2266, n2271, n2276, n2281, n2286, n2291, n2296,
    n2301, n2306, n2311, n2316, n2321, n2326, n2331, n2336, n2341, n2346,
    n2351, n2356, n2361, n2366, n2371, n2376, n2381, n2386, n2391, n2396,
    n2401, n2406, n2411, n2416, n2421, n2426, n2431, n2436, n2441, n2446,
    n2451, n2456, n2461, n2466, n2471, n2476, n2481, n2486, n2491, n2496,
    n2501, n2506, n2511, n2516, n2521, n2526, n2531, n2536, n2541, n2546,
    n2551, n2556, n2561, n2565, n2570, n2575, n2580, n2585, n2590, n2595,
    n2600, n2605, n2610, n2614, n2619, n2623, n2628, n2633, n2638, n2643,
    n2648, n2653, n2658, n2663, n2668, n2673, n2678, n2683, n2688, n2693,
    n2698, n2703, n2707, n2712, n2716, n2721, n2726, n2731, n2736, n2741,
    n2746, n2751, n2756, n2761, n2766, n2771, n2776, n2781, n2786, n2791,
    n2796, n2801, n2806, n2810, n2815, n2820, n2823, n2828, n2833, n2838,
    n2843, n2848, n2853, n2858, n2863, n2868, n2873, n2878, n2883, n2888,
    n2892, n2897, n2902, n2907, n2912, n2917, n2922, n2927, n2932, n2937,
    n2942, n2947, n2952, n2957, n2961, n2966, n2971, n2976, n2981, n2986,
    n2991, n2996, n3001, n3006, n3011, n3016, n3021, n3026, n3031, n3036,
    n3041, n3046, n3051, n3056, n3061, n3066, n3071, n3076, n3081, n3086,
    n3091, n3096, n3101, n3106, n3111, n3116, n3121, n3126, n3131, n3136,
    n3141, n3146, n3150, n3155, n3160, n3165, n3170, n3175, n3180, n3185,
    n3190, n3195, n3200, n3205, n3210, n3215, n3220, n3224, n3228, n3233,
    n3237, n3242, n3247, n3252, n3257, n3262, n3267, n3272, n3276, n3281,
    n3284, n3289, n3294, n3299, n3304, n3309, n3314, n3319, n3324, n3329,
    n3334, n3339, n3344, n3349, n3354, n3359, n3364, n3367, n3372, n3377,
    n3382, n3386, n3391, n3396, n3401, n3406, n3411, n3416, n3421, n3426,
    n3431, n3436, n3441, n3446, n3451, n3456, n3461, n3466, n3470, n3475,
    n3479, n3482, n3487, n3491, n3496, n3501, n3506, n3511, n3516, n3521,
    n3526, n3531, n3536, n3541, n3546, n3551, n3556, n3561, n3566, n3571,
    n3576, n3581, n3586, n3591, n3596, n3601, n3606, n3611, n3616, n3621,
    n3626, n3631, n3636, n3641, n3645, n3650, n3655, n3660, n3665, n3670,
    n3675, n3680, n3685, n3690, n3695, n3700, n3705, n3710, n3715, n3720,
    n3725, n3730, n3735, n3740, n3745, n3750, n3755, n3760, n3765, n3770,
    n3775, n3780, n3785, n3790, n3795, n3800, n3805, n3810, n3815, n3820,
    n3825, n3830, n3835, n3840, n3845, n3850, n3855, n3860, n3865, n3868,
    n3873, n3878, n3883, n3888, n3893, n3898, n3903, n3908, n3913, n3918,
    n3923, n3927, n3932, n3935, n3940, n3944, n3949, n3954, n3959, n3964,
    n3969, n3974, n3979, n3984, n3989, n3994, n3999, n4002, n4007, n4011,
    n4016, n4021, n4026, n4031, n4036, n4040, n4044, n4049, n4053, n4058,
    n4063, n4068, n4073, n4078, n4083, n4088, n4093, n4098, n4103, n4108,
    n4113, n4118, n4123, n4128, n4133, n4138, n4143, n4148, n4153, n4158,
    n4162, n4167, n4172, n4176, n4181, n4186, n4191, n4196, n4201, n4206,
    n4211, n4216, n4221, n4226, n4231, n4236, n4240, n4245, n4250, n4255,
    n4260, n4265, n4270, n4275, n4280, n4285, n4290, n4295, n4300, n4305,
    n4310, n4314, n4319, n4324, n4329, n4334, n4339, n4344, n4349, n4354,
    n4358, n4363, n4367, n4372, n4377, n4382, n4387, n4392, n4397, n4402,
    n4407, n4412, n4417, n4422, n4427, n4432, n4437, n4442, n4447, n4452,
    n4457, n4462, n4467, n4472, n4477, n4482, n4487, n4492, n4497, n4502,
    n4507, n4511, n4516, n4521, n4525, n4530, n4535, n4540, n4545, n4550,
    n4555, n4560, n4564, n4569, n4573, n4577, n4581, n4585, n4590, n4595,
    n4599, n4604, n4609, n4614, n4619, n4624, n4629, n4634, n4639, n4644,
    n4649, n4654, n4657, n4662, n4666, n4671, n4676, n4681, n4686, n4691,
    n4694, n4699, n4704, n4708, n4713, n4718, n4723, n4728, n4732, n4737,
    n4742, n4747, n4752, n4757, n4762, n4767, n4772, n4777, n4782, n4787,
    n4792, n4797, n4802, n4807, n4812, n4817, n4822, n4827, n4832, n4837,
    n4842, n4847, n4852, n4857, n4862, n4867, n4872, n4877, n4882, n4887,
    n4892, n4897, n4902, n4907, n4912, n4917, n4922, n4927, n4932, n4937,
    n4942, n4947, n4952, n4957, n4962, n4967, n4972, n4977, n4982, n4987,
    n4992, n4997, n5002, n5007, n5012, n5017, n5022, n5027, n5032, n5037,
    n5042, n5047, n5052, n5057, n5062, n5067, n5072, n5077, n5082, n5087,
    n5092, n5097, n5102, n5107, n5112, n5117, n5122, n5127, n5132, n5137,
    n5142, n5147, n5152, n5157, n5162, n5167, n5172, n5177, n5182, n5187,
    n5192, n5197, n5202, n5207, n5212, n5217, n5222, n5227, n5232, n5237,
    n5242, n5247, n5252, n5257, n5262, n5267, n5272, n5277, n5282, n5287,
    n5292, n5297, n5302, n5305, n5309, n5313, n5316, n5321, n5326, n5330,
    n5335, n5340, n5345, n5350, n5355, n5360, n5365, n5369, n5373, n5378,
    n5383, n5388, n5393, n5398, n5403, n5408, n5413, n5418, n5422, n5427,
    n5431, n5436, n5439, n5443, n5448, n5453, n5458, n5463, n5468, n5473,
    n5478, n5483, n5488, n5493, n5498, n5503, n5508, n5513, n5517, n5522,
    n5526, n5531, n5535, n5540, n5545, n5549, n5553, n5556, n5561, n5566,
    n5570, n5575, n5580, n5585, n5590, n5595, n5600, n5605, n5610, n5615,
    n5620, n5625, n5630, n5634, n5639, n5644, n5649, n5654, n5659, n5664,
    n5669, n5674, n5679, n5684, n5689, n5694, n5699, n5704, n5709, n5714,
    n5719, n5724, n5729, n5734, n5738, n5743, n5748, n5753, n5758, n5763,
    n5768, n5773, n5778, n5783, n5788, n5793, n5798, n5803, n5808, n5813,
    n5818, n5823, n5828, n5833, n5838, n5843, n5848, n5853, n5858, n5863,
    n5868, n5873, n5878, n5883, n5888, n5893, n5898, n5903, n5908, n5913,
    n5918, n5923, n5928, n5933, n5938, n5943, n5948, n5953, n5958, n5962,
    n5967, n5972, n5977, n5982, n5987, n5992, n5997, n6002, n6007, n6012,
    n6017, n6022, n6027, n6032, n6037, n6042, n6047, n6052, n6057, n6062,
    n6067, n6072, n6077, n6082, n6087, n6092, n6097, n6102, n6107, n6112,
    n6117, n6122, n6127, n6132, n6137, n6142, n6147, n6152, n6157, n6162,
    n6167, n6172, n6177, n6182, n6185, n6189, n6193, n6198, n6201, n6206,
    n6211, n6214, n6219, n6224, n6229, n6234, n6239, n6244, n6249, n6254,
    n6259, n6264, n6269, n6274, n6279, n6284, n6289, n6294, n6299, n6304,
    n6309, n6314, n6319, n6323, n6328, n6331, n6336, n6339, n6344, n6348,
    n6353, n6358, n6363, n6368, n6373, n6378, n6383, n6388, n6393, n6398,
    n6403, n6408, n6412, n6416, n6421, n6425, n6430, n6435, n6439, n6444,
    n6447, n6452, n6457, n6460, n6465, n6470, n6475, n6480, n6485, n6490,
    n6495, n6500, n6505, n6510, n6515, n6520, n6525, n6530, n6535, n6540,
    n6545, n6550, n6555, n6560, n6565, n6570, n6575, n6580, n6585, n6590,
    n6595, n6600, n6605, n6610, n6614, n6619, n6624, n6629, n6633, n6638,
    n6643, n6648, n6653, n6657, n6662, n6666, n6671, n6676, n6681, n6686,
    n6691, n6696, n6701, n6706, n6711, n6715, n6720, n6725, n6730, n6735,
    n6740, n6745, n6750, n6755, n6760, n6765, n6770, n6775, n6779, n6783,
    n6788, n6793, n6798, n6803, n6808, n6813, n6818, n6823, n6828, n6833,
    n6838, n6843, n6848, n6853, n6858, n6863, n6868, n6873, n6877, n6882,
    n6887, n6892, n6897, n6902, n6907, n6912, n6917, n6922, n6927, n6931,
    n6936, n6941, n6946, n6951, n6956, n6961, n6966, n6971, n6976, n6981,
    n6986, n6991, n6995, n7000, n7004, n7009, n7014, n7019, n7024, n7029,
    n7033, n7038, n7043, n7048, n7053, n7058, n7063, n7068, n7073, n7078,
    n7082, n7087, n7092, n7097, n7102, n7107, n7112, n7117, n7122, n7127,
    n7131, n7136, n7141, n7145, n7150, n7155, n7160, n7165, n7170, n7174,
    n7179, n7183, n7188, n7193, n7198, n7203, n7208, n7213, n7218, n7223,
    n7228, n7233, n7238, n7243, n7248, n7253, n7258, n7262, n7267, n7271,
    n7276, n7281, n7285, n7290, n7295, n7300, n7304, n7309, n7314, n7319,
    n7324, n7327, n7332, n7335, n7340, n7345, n7350, n7355, n7360, n7365,
    n7370, n7375, n7379, n7384, n7387, n7392, n7396, n7401, n7406, n7411,
    n7416, n7421, n7426;
  assign new_n4531_ = pg3233 & ~pg3230;
  assign new_n4532_ = ~ng3110 & ~ng3191;
  assign new_n4533_ = ~ng3124 & ~ng3126;
  assign new_n4534_ = new_n4532_ & new_n4533_;
  assign new_n4535_1_ = ng3135 & ng3120;
  assign new_n4536_ = ~ng3147 & new_n4535_1_;
  assign new_n4537_ = ~ng3139 & new_n4536_;
  assign new_n4538_ = new_n4534_ & new_n4537_;
  assign new_n4539_ = ~ng3123 & new_n4538_;
  assign new_n4540_1_ = new_n4531_ & new_n4539_;
  assign n2171 = new_n4531_ & ~new_n4540_1_;
  assign new_n4542_ = ng3110 & ~ng3191;
  assign new_n4543_ = ~ng3124 & new_n4542_;
  assign new_n4544_ = ~ng3126 & new_n4543_;
  assign new_n4545_1_ = ng3135 & ~ng3120;
  assign new_n4546_ = ~ng3147 & new_n4545_1_;
  assign new_n4547_ = ~ng3139 & new_n4546_;
  assign new_n4548_ = new_n4544_ & new_n4547_;
  assign new_n4549_ = ng3105 & new_n4548_;
  assign new_n4550_1_ = ng3139 & new_n4546_;
  assign new_n4551_ = new_n4544_ & new_n4550_1_;
  assign new_n4552_ = ng3106 & new_n4551_;
  assign new_n4553_ = ~ng3135 & ng3120;
  assign new_n4554_ = ng3147 & new_n4553_;
  assign new_n4555_1_ = ng3139 & new_n4554_;
  assign new_n4556_ = new_n4544_ & new_n4555_1_;
  assign new_n4557_ = ng3104 & new_n4556_;
  assign new_n4558_ = ~new_n4549_ & ~new_n4552_;
  assign new_n4559_ = ~new_n4557_ & new_n4558_;
  assign new_n4560_1_ = ~ng3135 & ~ng3120;
  assign new_n4561_ = ng3147 & new_n4560_1_;
  assign new_n4562_ = ng3139 & new_n4561_;
  assign new_n4563_ = new_n4544_ & new_n4562_;
  assign new_n4564_1_ = ng3102 & new_n4563_;
  assign new_n4565_ = ~ng3139 & new_n4554_;
  assign new_n4566_ = new_n4544_ & new_n4565_;
  assign new_n4567_ = ng3103 & new_n4566_;
  assign new_n4568_ = ~ng3139 & new_n4561_;
  assign new_n4569_1_ = new_n4544_ & new_n4568_;
  assign new_n4570_ = ng3101 & new_n4569_1_;
  assign new_n4571_ = ~new_n4564_1_ & ~new_n4567_;
  assign new_n4572_ = ~new_n4570_ & new_n4571_;
  assign new_n4573_1_ = ng3139 & new_n4536_;
  assign new_n4574_ = new_n4544_ & new_n4573_1_;
  assign new_n4575_ = ng3108 & new_n4574_;
  assign new_n4576_ = new_n4537_ & new_n4544_;
  assign new_n4577_1_ = ng3107 & new_n4576_;
  assign new_n4578_ = ~new_n4575_ & ~new_n4577_1_;
  assign new_n4579_ = new_n4559_ & new_n4572_;
  assign new_n4580_ = new_n4578_ & new_n4579_;
  assign new_n4581_1_ = ng3147 & new_n4535_1_;
  assign new_n4582_ = ~ng3139 & new_n4581_1_;
  assign new_n4583_ = new_n4534_ & new_n4582_;
  assign new_n4584_ = ng3147 & new_n4583_;
  assign new_n4585_1_ = ~ng3147 & new_n4560_1_;
  assign new_n4586_ = ~ng3139 & new_n4585_1_;
  assign new_n4587_ = new_n4544_ & new_n4586_;
  assign new_n4588_ = ng3097 & new_n4587_;
  assign new_n4589_ = ng3147 & new_n4545_1_;
  assign new_n4590_1_ = ~ng3139 & new_n4589_;
  assign new_n4591_ = new_n4534_ & new_n4590_1_;
  assign new_n4592_ = ng3147 & new_n4591_;
  assign new_n4593_ = ~new_n4584_ & ~new_n4588_;
  assign new_n4594_ = ~new_n4592_ & new_n4593_;
  assign new_n4595_1_ = new_n4534_ & new_n4568_;
  assign new_n4596_ = ng3147 & new_n4595_1_;
  assign new_n4597_ = ~ng3128 & new_n4538_;
  assign new_n4598_ = ~ng2991 & ~ng2992;
  assign new_n4599_1_ = new_n4534_ & new_n4586_;
  assign new_n4600_ = ~new_n4598_ & new_n4599_1_;
  assign new_n4601_ = ~new_n4596_ & ~new_n4597_;
  assign new_n4602_ = ~new_n4600_ & new_n4601_;
  assign new_n4603_ = ~ng3147 & new_n4553_;
  assign new_n4604_1_ = ~ng3139 & new_n4603_;
  assign new_n4605_ = new_n4544_ & new_n4604_1_;
  assign new_n4606_ = ng3099 & new_n4605_;
  assign new_n4607_ = ng3139 & new_n4603_;
  assign new_n4608_ = new_n4544_ & new_n4607_;
  assign new_n4609_1_ = ng3100 & new_n4608_;
  assign new_n4610_ = ng3139 & new_n4585_1_;
  assign new_n4611_ = new_n4544_ & new_n4610_;
  assign new_n4612_ = ng3098 & new_n4611_;
  assign new_n4613_ = ~new_n4606_ & ~new_n4609_1_;
  assign new_n4614_1_ = ~new_n4612_ & new_n4613_;
  assign new_n4615_ = new_n4580_ & new_n4594_;
  assign new_n4616_ = new_n4602_ & new_n4615_;
  assign new_n4617_ = new_n4614_1_ & new_n4616_;
  assign new_n4618_ = new_n4531_ & ~new_n4617_;
  assign n6112 = new_n4531_ & ~new_n4618_;
  assign new_n4620_ = ng3110 & new_n4595_1_;
  assign new_n4621_ = ~ng3125 & new_n4538_;
  assign new_n4622_ = ~new_n4620_ & ~new_n4621_;
  assign new_n4623_ = new_n4531_ & ~new_n4622_;
  assign n2873 = new_n4531_ & ~new_n4623_;
  assign new_n4625_ = ng3040 & ~ng2986;
  assign pg16496 = ~ng2987 | new_n4625_;
  assign new_n4627_ = ng3139 & new_n4591_;
  assign new_n4628_ = ng3139 & new_n4583_;
  assign new_n4629_1_ = ~ng185 & new_n4538_;
  assign new_n4630_ = ~new_n4627_ & ~new_n4628_;
  assign new_n4631_ = ~new_n4629_1_ & new_n4630_;
  assign new_n4632_ = new_n4534_ & new_n4550_1_;
  assign new_n4633_ = new_n4534_ & new_n4547_;
  assign new_n4634_1_ = ~new_n4599_1_ & ~new_n4632_;
  assign new_n4635_ = ~new_n4633_ & new_n4634_1_;
  assign new_n4636_ = ng3139 & new_n4589_;
  assign new_n4637_ = new_n4544_ & new_n4636_;
  assign new_n4638_ = ~ng185 & new_n4637_;
  assign new_n4639_1_ = ~ng2984 & ~ng2985;
  assign new_n4640_ = ng3120 & ~new_n4639_1_;
  assign new_n4641_ = ng3147 & ~new_n4598_;
  assign new_n4642_ = ~new_n4640_ & ~new_n4641_;
  assign new_n4643_ = new_n4544_ & new_n4590_1_;
  assign new_n4644_1_ = new_n4642_ & new_n4643_;
  assign new_n4645_ = ~new_n4638_ & ~new_n4644_1_;
  assign new_n4646_ = new_n4631_ & new_n4635_;
  assign new_n4647_ = new_n4645_ & new_n4646_;
  assign new_n4648_ = new_n4531_ & ~new_n4647_;
  assign n5659 = new_n4531_ & ~new_n4648_;
  assign new_n4650_ = ng3182 & new_n4551_;
  assign new_n4651_ = ng3185 & new_n4576_;
  assign new_n4652_ = ng3179 & new_n4548_;
  assign new_n4653_ = ~new_n4650_ & ~new_n4651_;
  assign new_n4654_1_ = ~new_n4652_ & new_n4653_;
  assign new_n4655_ = ng3173 & new_n4566_;
  assign new_n4656_ = ng3176 & new_n4556_;
  assign new_n4657_1_ = ng3170 & new_n4563_;
  assign new_n4658_ = ~new_n4655_ & ~new_n4656_;
  assign new_n4659_ = ~new_n4657_1_ & new_n4658_;
  assign new_n4660_ = ng3088 & new_n4574_;
  assign new_n4661_ = new_n4654_1_ & new_n4659_;
  assign new_n4662_1_ = ~new_n4660_ & new_n4661_;
  assign new_n4663_ = ng3155 & new_n4587_;
  assign new_n4664_ = ng3158 & new_n4611_;
  assign new_n4665_ = ng3135 & new_n4591_;
  assign new_n4666_1_ = ~new_n4663_ & ~new_n4664_;
  assign new_n4667_ = ~new_n4665_ & new_n4666_1_;
  assign new_n4668_ = ng3135 & new_n4538_;
  assign new_n4669_ = ng3135 & new_n4595_1_;
  assign new_n4670_ = ~new_n4668_ & ~new_n4669_;
  assign new_n4671_1_ = ng3164 & new_n4608_;
  assign new_n4672_ = ng3167 & new_n4569_1_;
  assign new_n4673_ = ng3161 & new_n4605_;
  assign new_n4674_ = ~new_n4671_1_ & ~new_n4672_;
  assign new_n4675_ = ~new_n4673_ & new_n4674_;
  assign new_n4676_1_ = new_n4662_1_ & new_n4667_;
  assign new_n4677_ = new_n4670_ & new_n4676_1_;
  assign new_n4678_ = new_n4675_ & new_n4677_;
  assign new_n4679_ = new_n4531_ & ~new_n4678_;
  assign pg26149 = ~new_n4531_ | new_n4679_;
  assign new_n4681_1_ = ng3126 & new_n4595_1_;
  assign new_n4682_ = ng3126 & new_n4538_;
  assign new_n4683_ = ~new_n4681_1_ & ~new_n4682_;
  assign new_n4684_ = new_n4531_ & ~new_n4683_;
  assign pg25420 = ~new_n4531_ | new_n4684_;
  assign new_n4686_1_ = ng3124 & new_n4595_1_;
  assign new_n4687_ = ng3124 & new_n4538_;
  assign new_n4688_ = ~new_n4686_1_ & ~new_n4687_;
  assign new_n4689_ = new_n4531_ & ~new_n4688_;
  assign pg25442 = ~new_n4531_ | new_n4689_;
  assign new_n4691_1_ = ~ng3120 & ~ng3147;
  assign new_n4692_ = ~ng3139 & new_n4691_1_;
  assign new_n4693_ = ~ng3097 & ng3139;
  assign new_n4694_1_ = ng3139 & ~new_n4693_;
  assign new_n4695_ = ng3120 & new_n4694_1_;
  assign new_n4696_ = ng3147 & ~new_n4695_;
  assign new_n4697_ = ~ng3139 & new_n4598_;
  assign new_n4698_ = ~ng3139 & ~new_n4697_;
  assign new_n4699_1_ = ng3120 & new_n4698_;
  assign new_n4700_ = ng3139 & new_n4639_1_;
  assign new_n4701_ = ~ng3120 & ~new_n4700_;
  assign new_n4702_ = ~new_n4699_1_ & ~new_n4701_;
  assign new_n4703_ = ~ng3147 & new_n4702_;
  assign new_n4704_1_ = ~new_n4696_ & ~new_n4703_;
  assign new_n4705_ = ~new_n4692_ & new_n4704_1_;
  assign pg25489 = new_n4692_ | new_n4705_;
  assign new_n4707_ = ng3093 & new_n4548_;
  assign new_n4708_1_ = ng3094 & new_n4551_;
  assign new_n4709_ = ng3092 & new_n4556_;
  assign new_n4710_ = ~new_n4707_ & ~new_n4708_1_;
  assign new_n4711_ = ~new_n4709_ & new_n4710_;
  assign new_n4712_ = ng3087 & new_n4563_;
  assign new_n4713_1_ = ng3091 & new_n4566_;
  assign new_n4714_ = ng3086 & new_n4569_1_;
  assign new_n4715_ = ~new_n4712_ & ~new_n4713_1_;
  assign new_n4716_ = ~new_n4714_ & new_n4715_;
  assign new_n4717_ = ng3096 & new_n4574_;
  assign new_n4718_1_ = ng3095 & new_n4576_;
  assign new_n4719_ = ~new_n4717_ & ~new_n4718_1_;
  assign new_n4720_ = new_n4711_ & new_n4716_;
  assign new_n4721_ = new_n4719_ & new_n4720_;
  assign new_n4722_ = ng3120 & new_n4583_;
  assign new_n4723_1_ = ng3210 & new_n4587_;
  assign new_n4724_ = ng3120 & new_n4591_;
  assign new_n4725_ = ~new_n4722_ & ~new_n4723_1_;
  assign new_n4726_ = ~new_n4724_ & new_n4725_;
  assign new_n4727_ = ng3120 & new_n4595_1_;
  assign new_n4728_1_ = ng3120 & new_n4538_;
  assign new_n4729_ = new_n4599_1_ & ~new_n4639_1_;
  assign new_n4730_ = ~new_n4727_ & ~new_n4728_1_;
  assign new_n4731_ = ~new_n4729_ & new_n4730_;
  assign new_n4732_1_ = ng3084 & new_n4605_;
  assign new_n4733_ = ng3085 & new_n4608_;
  assign new_n4734_ = ng3211 & new_n4611_;
  assign new_n4735_ = ~new_n4732_1_ & ~new_n4733_;
  assign new_n4736_ = ~new_n4734_ & new_n4735_;
  assign new_n4737_1_ = new_n4721_ & new_n4726_;
  assign new_n4738_ = new_n4731_ & new_n4737_1_;
  assign new_n4739_ = new_n4736_ & new_n4738_;
  assign new_n4740_ = new_n4531_ & ~new_n4739_;
  assign pg26104 = ~new_n4531_ | new_n4740_;
  assign new_n4742_1_ = ~ng544 & ng499;
  assign new_n4743_ = ng548 & ~ng1309;
  assign new_n4744_ = ~ng499 & ~new_n4743_;
  assign n4521 = ~new_n4742_1_ & ~new_n4744_;
  assign new_n4746_ = ng1309 & ~n4521;
  assign new_n4747_1_ = ~ng3097 & ~ng1309;
  assign n272 = ~new_n4746_ & ~new_n4747_1_;
  assign new_n4749_ = ~ng2618 & ng2574;
  assign new_n4750_ = ~ng1924 & ng1880;
  assign new_n4751_ = ng1186 & ~ng1230;
  assign new_n4752_1_ = ng1309 & n4521;
  assign new_n4753_ = ng1234 & ~ng1309;
  assign new_n4754_ = ~new_n4752_1_ & ~new_n4753_;
  assign new_n4755_ = ~ng1186 & new_n4754_;
  assign n1448 = ~new_n4751_ & ~new_n4755_;
  assign new_n4757_1_ = ng1309 & n1448;
  assign new_n4758_ = ng1928 & ~ng1309;
  assign new_n4759_ = ~new_n4757_1_ & ~new_n4758_;
  assign new_n4760_ = ~ng1880 & new_n4759_;
  assign n2721 = ~new_n4750_ & ~new_n4760_;
  assign new_n4762_1_ = ng1309 & n2721;
  assign new_n4763_ = ~ng1309 & ng2622;
  assign new_n4764_ = ~new_n4762_1_ & ~new_n4763_;
  assign new_n4765_ = ~ng2574 & new_n4764_;
  assign n4713 = ~new_n4749_ & ~new_n4765_;
  assign new_n4767_1_ = ng1315 & ~n4713;
  assign new_n4768_ = ~ng3108 & ~ng1315;
  assign n277 = ~new_n4767_1_ & ~new_n4768_;
  assign new_n4770_ = ng1312 & ~ng2574;
  assign new_n4771_ = ~ng3185 & ~ng1312;
  assign n282 = ~new_n4770_ & ~new_n4771_;
  assign new_n4773_ = ng853 & ng2257;
  assign new_n4774_ = ~ng141 & ~new_n4773_;
  assign new_n4775_ = ng105 & new_n4773_;
  assign n292 = ~new_n4774_ & ~new_n4775_;
  assign new_n4777_1_ = ng823 & ng2257;
  assign new_n4778_ = ~ng155 & ~new_n4777_1_;
  assign new_n4779_ = ng121 & new_n4777_1_;
  assign n297 = ~new_n4778_ & ~new_n4779_;
  assign new_n4781_ = ng823 & ~ng316;
  assign new_n4782_1_ = ~ng317 & ng853;
  assign new_n4783_ = ng826 & ~ng315;
  assign new_n4784_ = ~new_n4781_ & ~new_n4782_1_;
  assign new_n4785_ = ~new_n4783_ & new_n4784_;
  assign new_n4786_ = ~ng313 & ng823;
  assign new_n4787_1_ = ~ng314 & ng853;
  assign new_n4788_ = ~ng312 & ng826;
  assign new_n4789_ = ~new_n4786_ & ~new_n4787_1_;
  assign new_n4790_ = ~new_n4788_ & new_n4789_;
  assign new_n4791_ = ~ng319 & ng823;
  assign new_n4792_1_ = ~ng320 & ng853;
  assign new_n4793_ = ~ng318 & ng826;
  assign new_n4794_ = ~new_n4791_ & ~new_n4792_1_;
  assign new_n4795_ = ~new_n4793_ & new_n4794_;
  assign new_n4796_ = ~new_n4785_ & new_n4790_;
  assign new_n4797_1_ = new_n4795_ & new_n4796_;
  assign new_n4798_ = new_n4785_ & new_n4790_;
  assign new_n4799_ = new_n4795_ & new_n4798_;
  assign new_n4800_ = ~new_n4797_1_ & ~new_n4799_;
  assign new_n4801_ = ng198 & ng823;
  assign new_n4802_1_ = ng853 & ng201;
  assign new_n4803_ = ng195 & ng826;
  assign new_n4804_ = ~new_n4801_ & ~new_n4802_1_;
  assign new_n4805_ = ~new_n4803_ & new_n4804_;
  assign new_n4806_ = ng823 & ng243;
  assign new_n4807_1_ = ng853 & ng246;
  assign new_n4808_ = ng826 & ng240;
  assign new_n4809_ = ~new_n4806_ & ~new_n4807_1_;
  assign new_n4810_ = ~new_n4808_ & new_n4809_;
  assign new_n4811_ = ng234 & ng823;
  assign new_n4812_1_ = ng237 & ng853;
  assign new_n4813_ = ng231 & ng826;
  assign new_n4814_ = ~new_n4811_ & ~new_n4812_1_;
  assign new_n4815_ = ~new_n4813_ & new_n4814_;
  assign new_n4816_ = ~new_n4805_ & ~new_n4810_;
  assign new_n4817_1_ = ~new_n4815_ & new_n4816_;
  assign new_n4818_ = ng270 & ng823;
  assign new_n4819_ = ng273 & ng853;
  assign new_n4820_ = ng826 & ng267;
  assign new_n4821_ = ~new_n4818_ & ~new_n4819_;
  assign new_n4822_1_ = ~new_n4820_ & new_n4821_;
  assign new_n4823_ = ng261 & ng823;
  assign new_n4824_ = ng264 & ng853;
  assign new_n4825_ = ng258 & ng826;
  assign new_n4826_ = ~new_n4823_ & ~new_n4824_;
  assign new_n4827_1_ = ~new_n4825_ & new_n4826_;
  assign new_n4828_ = ng207 & ng823;
  assign new_n4829_ = ng210 & ng853;
  assign new_n4830_ = ng204 & ng826;
  assign new_n4831_ = ~new_n4828_ & ~new_n4829_;
  assign new_n4832_1_ = ~new_n4830_ & new_n4831_;
  assign new_n4833_ = ng252 & ng823;
  assign new_n4834_ = ng255 & ng853;
  assign new_n4835_ = ng249 & ng826;
  assign new_n4836_ = ~new_n4833_ & ~new_n4834_;
  assign new_n4837_1_ = ~new_n4835_ & new_n4836_;
  assign new_n4838_ = ng823 & ng189;
  assign new_n4839_ = ng192 & ng853;
  assign new_n4840_ = ng826 & ng186;
  assign new_n4841_ = ~new_n4838_ & ~new_n4839_;
  assign new_n4842_1_ = ~new_n4840_ & new_n4841_;
  assign new_n4843_ = new_n4832_1_ & new_n4837_1_;
  assign new_n4844_ = new_n4842_1_ & new_n4843_;
  assign new_n4845_ = ng216 & ng823;
  assign new_n4846_ = ng219 & ng853;
  assign new_n4847_1_ = ng213 & ng826;
  assign new_n4848_ = ~new_n4845_ & ~new_n4846_;
  assign new_n4849_ = ~new_n4847_1_ & new_n4848_;
  assign new_n4850_ = new_n4827_1_ & new_n4844_;
  assign new_n4851_ = new_n4849_ & new_n4850_;
  assign new_n4852_1_ = ng225 & ng823;
  assign new_n4853_ = ng853 & ng228;
  assign new_n4854_ = ng222 & ng826;
  assign new_n4855_ = ~new_n4852_1_ & ~new_n4853_;
  assign new_n4856_ = ~new_n4854_ & new_n4855_;
  assign new_n4857_1_ = new_n4817_1_ & ~new_n4822_1_;
  assign new_n4858_ = new_n4851_ & new_n4857_1_;
  assign new_n4859_ = ~new_n4856_ & new_n4858_;
  assign new_n4860_ = new_n4797_1_ & new_n4859_;
  assign new_n4861_ = new_n4805_ & new_n4810_;
  assign new_n4862_1_ = new_n4815_ & new_n4861_;
  assign new_n4863_ = new_n4822_1_ & new_n4862_1_;
  assign new_n4864_ = new_n4851_ & new_n4863_;
  assign new_n4865_ = new_n4856_ & new_n4864_;
  assign new_n4866_ = ~new_n4797_1_ & new_n4865_;
  assign new_n4867_1_ = ~new_n4860_ & ~new_n4866_;
  assign new_n4868_ = ~new_n4800_ & ~new_n4867_1_;
  assign new_n4869_ = ~ng170 & ng823;
  assign new_n4870_ = ~ng168 & ng853;
  assign new_n4871_ = ng826 & ~ng169;
  assign new_n4872_1_ = ~new_n4869_ & ~new_n4870_;
  assign new_n4873_ = ~new_n4871_ & new_n4872_1_;
  assign new_n4874_ = ng101 & ~new_n4815_;
  assign new_n4875_ = ng101 & ~new_n4874_;
  assign new_n4876_ = ~new_n4815_ & ~new_n4874_;
  assign new_n4877_1_ = ~new_n4875_ & ~new_n4876_;
  assign new_n4878_ = ng125 & ~new_n4827_1_;
  assign new_n4879_ = ng125 & ~new_n4878_;
  assign new_n4880_ = ~new_n4827_1_ & ~new_n4878_;
  assign new_n4881_ = ~new_n4879_ & ~new_n4880_;
  assign new_n4882_1_ = new_n4877_1_ & new_n4881_;
  assign new_n4883_ = ng109 & ~new_n4810_;
  assign new_n4884_ = ng109 & ~new_n4883_;
  assign new_n4885_ = ~new_n4810_ & ~new_n4883_;
  assign new_n4886_ = ~new_n4884_ & ~new_n4885_;
  assign new_n4887_1_ = ng823 & ~ng173;
  assign new_n4888_ = ng853 & ~ng171;
  assign new_n4889_ = ~ng172 & ng826;
  assign new_n4890_ = ~new_n4887_1_ & ~new_n4888_;
  assign new_n4891_ = ~new_n4889_ & new_n4890_;
  assign new_n4892_1_ = ~new_n4822_1_ & ~new_n4891_;
  assign new_n4893_ = ~new_n4891_ & ~new_n4892_1_;
  assign new_n4894_ = ~new_n4822_1_ & ~new_n4892_1_;
  assign new_n4895_ = ~new_n4893_ & ~new_n4894_;
  assign new_n4896_ = new_n4886_ & new_n4895_;
  assign new_n4897_1_ = ng117 & ~new_n4837_1_;
  assign new_n4898_ = ng117 & ~new_n4897_1_;
  assign new_n4899_ = ~new_n4837_1_ & ~new_n4897_1_;
  assign new_n4900_ = ~new_n4898_ & ~new_n4899_;
  assign new_n4901_ = ~new_n4882_1_ & ~new_n4896_;
  assign new_n4902_1_ = ~new_n4900_ & new_n4901_;
  assign new_n4903_ = new_n4881_ & new_n4900_;
  assign new_n4904_ = new_n4877_1_ & new_n4886_;
  assign new_n4905_ = ~new_n4903_ & ~new_n4904_;
  assign new_n4906_ = ~new_n4895_ & new_n4905_;
  assign new_n4907_1_ = new_n4881_ & new_n4895_;
  assign new_n4908_ = new_n4886_ & new_n4900_;
  assign new_n4909_ = ~new_n4907_1_ & ~new_n4908_;
  assign new_n4910_ = ~new_n4877_1_ & new_n4909_;
  assign new_n4911_ = ~new_n4902_1_ & ~new_n4906_;
  assign new_n4912_1_ = ~new_n4910_ & new_n4911_;
  assign new_n4913_ = ng2257 & ~new_n4873_;
  assign new_n4914_ = ~new_n4912_1_ & new_n4913_;
  assign new_n4915_ = ng97 & ~new_n4842_1_;
  assign new_n4916_ = ng97 & ~new_n4915_;
  assign new_n4917_1_ = ~new_n4842_1_ & ~new_n4915_;
  assign new_n4918_ = ~new_n4916_ & ~new_n4917_1_;
  assign new_n4919_ = ng121 & ~new_n4849_;
  assign new_n4920_ = ng121 & ~new_n4919_;
  assign new_n4921_ = ~new_n4849_ & ~new_n4919_;
  assign new_n4922_1_ = ~new_n4920_ & ~new_n4921_;
  assign new_n4923_ = new_n4918_ & new_n4922_1_;
  assign new_n4924_ = ng105 & ~new_n4805_;
  assign new_n4925_ = ng105 & ~new_n4924_;
  assign new_n4926_ = ~new_n4805_ & ~new_n4924_;
  assign new_n4927_1_ = ~new_n4925_ & ~new_n4926_;
  assign new_n4928_ = ~ng176 & ng823;
  assign new_n4929_ = ~ng174 & ng853;
  assign new_n4930_ = ng826 & ~ng175;
  assign new_n4931_ = ~new_n4928_ & ~new_n4929_;
  assign new_n4932_1_ = ~new_n4930_ & new_n4931_;
  assign new_n4933_ = ~new_n4856_ & ~new_n4932_1_;
  assign new_n4934_ = ~new_n4932_1_ & ~new_n4933_;
  assign new_n4935_ = ~new_n4856_ & ~new_n4933_;
  assign new_n4936_ = ~new_n4934_ & ~new_n4935_;
  assign new_n4937_1_ = new_n4927_1_ & new_n4936_;
  assign new_n4938_ = ng113 & ~new_n4832_1_;
  assign new_n4939_ = ng113 & ~new_n4938_;
  assign new_n4940_ = ~new_n4832_1_ & ~new_n4938_;
  assign new_n4941_ = ~new_n4939_ & ~new_n4940_;
  assign new_n4942_1_ = ~new_n4923_ & ~new_n4937_1_;
  assign new_n4943_ = ~new_n4941_ & new_n4942_1_;
  assign new_n4944_ = new_n4922_1_ & new_n4941_;
  assign new_n4945_ = new_n4918_ & new_n4927_1_;
  assign new_n4946_ = ~new_n4944_ & ~new_n4945_;
  assign new_n4947_1_ = ~new_n4936_ & new_n4946_;
  assign new_n4948_ = new_n4922_1_ & new_n4936_;
  assign new_n4949_ = new_n4927_1_ & new_n4941_;
  assign new_n4950_ = ~new_n4948_ & ~new_n4949_;
  assign new_n4951_ = ~new_n4918_ & new_n4950_;
  assign new_n4952_1_ = ~new_n4943_ & ~new_n4947_1_;
  assign new_n4953_ = ~new_n4951_ & new_n4952_1_;
  assign new_n4954_ = new_n4913_ & ~new_n4953_;
  assign new_n4955_ = ~new_n4914_ & ~new_n4954_;
  assign new_n4956_ = ~ng164 & ng823;
  assign new_n4957_1_ = ~ng162 & ng853;
  assign new_n4958_ = ng826 & ~ng163;
  assign new_n4959_ = ~new_n4956_ & ~new_n4957_1_;
  assign new_n4960_ = ~new_n4958_ & new_n4959_;
  assign new_n4961_ = ~new_n4891_ & ~new_n4960_;
  assign new_n4962_1_ = ~new_n4960_ & ~new_n4961_;
  assign new_n4963_ = ~new_n4891_ & ~new_n4961_;
  assign new_n4964_ = ~new_n4962_1_ & ~new_n4963_;
  assign new_n4965_ = ~ng155 & ng823;
  assign new_n4966_ = ~ng153 & ng853;
  assign new_n4967_1_ = ~ng154 & ng826;
  assign new_n4968_ = ~new_n4965_ & ~new_n4966_;
  assign new_n4969_ = ~new_n4967_1_ & new_n4968_;
  assign new_n4970_ = ng121 & ~new_n4969_;
  assign new_n4971_ = ~new_n4969_ & ~new_n4970_;
  assign new_n4972_1_ = ng121 & ~new_n4970_;
  assign new_n4973_ = ~new_n4971_ & ~new_n4972_1_;
  assign new_n4974_ = ~ng158 & ng823;
  assign new_n4975_ = ~ng156 & ng853;
  assign new_n4976_ = ng826 & ~ng157;
  assign new_n4977_1_ = ~new_n4974_ & ~new_n4975_;
  assign new_n4978_ = ~new_n4976_ & new_n4977_1_;
  assign new_n4979_ = ng125 & ~new_n4978_;
  assign new_n4980_ = ~new_n4978_ & ~new_n4979_;
  assign new_n4981_ = ng125 & ~new_n4979_;
  assign new_n4982_1_ = ~new_n4980_ & ~new_n4981_;
  assign new_n4983_ = ng823 & ~ng152;
  assign new_n4984_ = ng853 & ~ng150;
  assign new_n4985_ = ng826 & ~ng151;
  assign new_n4986_ = ~new_n4983_ & ~new_n4984_;
  assign new_n4987_1_ = ~new_n4985_ & new_n4986_;
  assign new_n4988_ = ng117 & ~new_n4987_1_;
  assign new_n4989_ = ~new_n4987_1_ & ~new_n4988_;
  assign new_n4990_ = ng117 & ~new_n4988_;
  assign new_n4991_ = ~new_n4989_ & ~new_n4990_;
  assign new_n4992_1_ = new_n4973_ & new_n4982_1_;
  assign new_n4993_ = new_n4991_ & new_n4992_1_;
  assign new_n4994_ = ng823 & ~ng161;
  assign new_n4995_ = ~ng159 & ng853;
  assign new_n4996_ = ng826 & ~ng160;
  assign new_n4997_1_ = ~new_n4994_ & ~new_n4995_;
  assign new_n4998_ = ~new_n4996_ & new_n4997_1_;
  assign new_n4999_ = ~new_n4932_1_ & ~new_n4998_;
  assign new_n5000_ = ~new_n4998_ & ~new_n4999_;
  assign new_n5001_ = ~new_n4932_1_ & ~new_n4999_;
  assign new_n5002_1_ = ~new_n5000_ & ~new_n5001_;
  assign new_n5003_ = new_n4964_ & new_n4993_;
  assign new_n5004_ = new_n5002_1_ & new_n5003_;
  assign new_n5005_ = ~ng149 & ng823;
  assign new_n5006_ = ng853 & ~ng147;
  assign new_n5007_1_ = ng826 & ~ng148;
  assign new_n5008_ = ~new_n5005_ & ~new_n5006_;
  assign new_n5009_ = ~new_n5007_1_ & new_n5008_;
  assign new_n5010_ = ng113 & ~new_n5009_;
  assign new_n5011_ = ~new_n5009_ & ~new_n5010_;
  assign new_n5012_1_ = ng113 & ~new_n5010_;
  assign new_n5013_ = ~new_n5011_ & ~new_n5012_1_;
  assign new_n5014_ = ~ng134 & ng823;
  assign new_n5015_ = ng853 & ~ng132;
  assign new_n5016_ = ng826 & ~ng133;
  assign new_n5017_1_ = ~new_n5014_ & ~new_n5015_;
  assign new_n5018_ = ~new_n5016_ & new_n5017_1_;
  assign new_n5019_ = ng101 & ~new_n5018_;
  assign new_n5020_ = ~new_n5018_ & ~new_n5019_;
  assign new_n5021_ = ng101 & ~new_n5019_;
  assign new_n5022_1_ = ~new_n5020_ & ~new_n5021_;
  assign new_n5023_ = ng823 & ~ng143;
  assign new_n5024_ = ~ng141 & ng853;
  assign new_n5025_ = ng826 & ~ng142;
  assign new_n5026_ = ~new_n5023_ & ~new_n5024_;
  assign new_n5027_1_ = ~new_n5025_ & new_n5026_;
  assign new_n5028_ = ng105 & ~new_n5027_1_;
  assign new_n5029_ = ~new_n5027_1_ & ~new_n5028_;
  assign new_n5030_ = ng105 & ~new_n5028_;
  assign new_n5031_ = ~new_n5029_ & ~new_n5030_;
  assign new_n5032_1_ = ~ng131 & ng823;
  assign new_n5033_ = ~ng129 & ng853;
  assign new_n5034_ = ~ng130 & ng826;
  assign new_n5035_ = ~new_n5032_1_ & ~new_n5033_;
  assign new_n5036_ = ~new_n5034_ & new_n5035_;
  assign new_n5037_1_ = ng97 & ~new_n5036_;
  assign new_n5038_ = ~new_n5036_ & ~new_n5037_1_;
  assign new_n5039_ = ng97 & ~new_n5037_1_;
  assign new_n5040_ = ~new_n5038_ & ~new_n5039_;
  assign new_n5041_ = new_n5022_1_ & new_n5031_;
  assign new_n5042_1_ = new_n5040_ & new_n5041_;
  assign new_n5043_ = ~ng146 & ng823;
  assign new_n5044_ = ~ng144 & ng853;
  assign new_n5045_ = ~ng145 & ng826;
  assign new_n5046_ = ~new_n5043_ & ~new_n5044_;
  assign new_n5047_1_ = ~new_n5045_ & new_n5046_;
  assign new_n5048_ = ng109 & ~new_n5047_1_;
  assign new_n5049_ = ~new_n5047_1_ & ~new_n5048_;
  assign new_n5050_ = ng109 & ~new_n5048_;
  assign new_n5051_ = ~new_n5049_ & ~new_n5050_;
  assign new_n5052_1_ = new_n5013_ & new_n5042_1_;
  assign new_n5053_ = new_n5051_ & new_n5052_1_;
  assign new_n5054_ = new_n5004_ & new_n5053_;
  assign new_n5055_ = ~new_n4873_ & new_n4955_;
  assign new_n5056_ = ng2257 & new_n5054_;
  assign new_n5057_1_ = new_n5055_ & new_n5056_;
  assign new_n5058_ = ~ng323 & ng823;
  assign new_n5059_ = ng853 & ~ng321;
  assign new_n5060_ = ~ng322 & ng826;
  assign new_n5061_ = ~new_n5058_ & ~new_n5059_;
  assign new_n5062_1_ = ~new_n5060_ & new_n5061_;
  assign new_n5063_ = new_n4785_ & ~new_n4790_;
  assign new_n5064_ = new_n4795_ & new_n5063_;
  assign new_n5065_ = new_n5057_1_ & ~new_n5062_1_;
  assign new_n5066_ = new_n5064_ & new_n5065_;
  assign new_n5067_1_ = new_n4913_ & new_n5054_;
  assign new_n5068_ = ~new_n4795_ & new_n5063_;
  assign new_n5069_ = ~new_n5062_1_ & new_n5067_1_;
  assign new_n5070_ = new_n5068_ & new_n5069_;
  assign new_n5071_ = ng2257 & new_n4873_;
  assign new_n5072_1_ = ~new_n4790_ & new_n5071_;
  assign new_n5073_ = ~new_n5066_ & ~new_n5070_;
  assign new_n5074_ = ~new_n5072_1_ & new_n5073_;
  assign new_n5075_ = ~ng404 & ng823;
  assign new_n5076_ = ng853 & ~ng402;
  assign new_n5077_1_ = ng826 & ~ng403;
  assign new_n5078_ = ~new_n5075_ & ~new_n5076_;
  assign new_n5079_ = ~new_n5077_1_ & new_n5078_;
  assign new_n5080_ = new_n5067_1_ & ~new_n5079_;
  assign new_n5081_ = new_n5074_ & ~new_n5080_;
  assign new_n5082_1_ = ~new_n4868_ & new_n5081_;
  assign new_n5083_ = new_n4868_ & new_n5081_;
  assign new_n5084_ = ng125 & ~new_n5083_;
  assign new_n5085_ = ~new_n5082_1_ & ~new_n5084_;
  assign new_n5086_ = new_n4797_1_ & ~new_n4849_;
  assign new_n5087_1_ = ~new_n4797_1_ & new_n4849_;
  assign new_n5088_ = ~new_n5086_ & ~new_n5087_1_;
  assign new_n5089_ = new_n4797_1_ & ~new_n4815_;
  assign new_n5090_ = ~new_n4797_1_ & new_n4815_;
  assign new_n5091_ = ~new_n5089_ & ~new_n5090_;
  assign new_n5092_1_ = new_n4797_1_ & new_n4842_1_;
  assign new_n5093_ = ~new_n4797_1_ & ~new_n4842_1_;
  assign new_n5094_ = ~new_n5092_1_ & ~new_n5093_;
  assign new_n5095_ = ~new_n4800_ & new_n5094_;
  assign new_n5096_ = ~new_n5091_ & new_n5095_;
  assign new_n5097_1_ = new_n4797_1_ & ~new_n4810_;
  assign new_n5098_ = ~new_n4797_1_ & new_n4810_;
  assign new_n5099_ = ~new_n5097_1_ & ~new_n5098_;
  assign new_n5100_ = new_n4797_1_ & ~new_n4805_;
  assign new_n5101_ = ~new_n4797_1_ & new_n4805_;
  assign new_n5102_1_ = ~new_n5100_ & ~new_n5101_;
  assign new_n5103_ = ~new_n5099_ & ~new_n5102_1_;
  assign new_n5104_ = new_n4797_1_ & ~new_n4837_1_;
  assign new_n5105_ = ~new_n4797_1_ & new_n4837_1_;
  assign new_n5106_ = ~new_n5104_ & ~new_n5105_;
  assign new_n5107_1_ = new_n4797_1_ & ~new_n4832_1_;
  assign new_n5108_ = ~new_n4797_1_ & new_n4832_1_;
  assign new_n5109_ = ~new_n5107_1_ & ~new_n5108_;
  assign new_n5110_ = ~new_n5106_ & ~new_n5109_;
  assign new_n5111_ = new_n5096_ & new_n5103_;
  assign new_n5112_1_ = new_n5110_ & new_n5111_;
  assign new_n5113_ = ~new_n5088_ & new_n5112_1_;
  assign new_n5114_ = new_n4827_1_ & new_n5113_;
  assign new_n5115_ = ~new_n4827_1_ & ~new_n5113_;
  assign new_n5116_ = ~new_n5114_ & ~new_n5115_;
  assign new_n5117_1_ = new_n5082_1_ & new_n5116_;
  assign new_n5118_ = ~new_n5085_ & ~new_n5117_1_;
  assign new_n5119_ = ng826 & ~new_n5118_;
  assign new_n5120_ = ~ng258 & ~ng826;
  assign n302 = ~new_n5119_ & ~new_n5120_;
  assign new_n5122_1_ = ~ng2892 & ~ng2903;
  assign new_n5123_ = ~ng2896 & new_n5122_1_;
  assign new_n5124_ = ~ng2908 & new_n5123_;
  assign new_n5125_ = ~ng2900 & new_n5124_;
  assign new_n5126_ = ng2257 & new_n5125_;
  assign new_n5127_1_ = ng853 & new_n5126_;
  assign new_n5128_ = ng853 & ~new_n5125_;
  assign new_n5129_ = ng92 & new_n5128_;
  assign new_n5130_ = ng88 & new_n5129_;
  assign new_n5131_ = ~ng83 & new_n5130_;
  assign new_n5132_1_ = ng83 & ~new_n5130_;
  assign new_n5133_ = ~new_n5131_ & ~new_n5132_1_;
  assign n307 = ~new_n5127_1_ & ~new_n5133_;
  assign new_n5135_ = ~new_n4799_ & new_n5125_;
  assign new_n5136_ = ~new_n4795_ & new_n4796_;
  assign new_n5137_1_ = ~new_n5135_ & ~new_n5136_;
  assign new_n5138_ = ng826 & new_n5137_1_;
  assign new_n5139_ = ~ng369 & ~new_n5138_;
  assign new_n5140_ = ~ng373 & ng823;
  assign new_n5141_ = ~ng376 & ng853;
  assign new_n5142_1_ = ng826 & ~ng384;
  assign new_n5143_ = ~new_n5140_ & ~new_n5141_;
  assign new_n5144_ = ~new_n5142_1_ & new_n5143_;
  assign new_n5145_ = ~ng343 & ng823;
  assign new_n5146_ = ~ng346 & ng853;
  assign new_n5147_1_ = ~ng354 & ng826;
  assign new_n5148_ = ~new_n5145_ & ~new_n5146_;
  assign new_n5149_ = ~new_n5147_1_ & new_n5148_;
  assign new_n5150_ = ~new_n5144_ & new_n5149_;
  assign new_n5151_ = ~pg3229 & new_n5150_;
  assign new_n5152_1_ = ~new_n5144_ & ~new_n5149_;
  assign new_n5153_ = pg3229 & new_n5152_1_;
  assign new_n5154_ = ~ng358 & ng823;
  assign new_n5155_ = ng853 & ~ng361;
  assign new_n5156_ = ~ng369 & ng826;
  assign new_n5157_1_ = ~new_n5154_ & ~new_n5155_;
  assign new_n5158_ = ~new_n5156_ & new_n5157_1_;
  assign new_n5159_ = new_n5144_ & ~new_n5158_;
  assign new_n5160_ = ~new_n5151_ & ~new_n5153_;
  assign new_n5161_ = ~new_n5159_ & new_n5160_;
  assign new_n5162_1_ = new_n5138_ & ~new_n5161_;
  assign n312 = ~new_n5139_ & ~new_n5162_1_;
  assign new_n5164_ = ng411 & ng823;
  assign new_n5165_ = ng414 & ng853;
  assign new_n5166_ = ng408 & ng826;
  assign new_n5167_1_ = ~new_n5164_ & ~new_n5165_;
  assign new_n5168_ = ~new_n5166_ & new_n5167_1_;
  assign new_n5169_ = ng823 & ng420;
  assign new_n5170_ = ng853 & ng423;
  assign new_n5171_ = ng826 & ng417;
  assign new_n5172_1_ = ~new_n5169_ & ~new_n5170_;
  assign n4167 = new_n5171_ | ~new_n5172_1_;
  assign new_n5174_ = ng117 & ng125;
  assign new_n5175_ = ng121 & new_n5174_;
  assign new_n5176_ = ng113 & new_n5175_;
  assign new_n5177_1_ = ng101 & ng109;
  assign new_n5178_ = ng105 & new_n5177_1_;
  assign new_n5179_ = ng97 & new_n5178_;
  assign new_n5180_ = new_n5176_ & new_n5179_;
  assign new_n5181_ = ~new_n4891_ & ~new_n4932_1_;
  assign new_n5182_1_ = new_n5180_ & new_n5181_;
  assign new_n5183_ = ~ng428 & ng823;
  assign new_n5184_ = ~ng426 & ng853;
  assign new_n5185_ = ~ng427 & ng826;
  assign new_n5186_ = ~new_n5183_ & ~new_n5184_;
  assign new_n5187_1_ = ~new_n5185_ & new_n5186_;
  assign new_n5188_ = ~new_n5182_1_ & new_n5187_1_;
  assign new_n5189_ = n4167 & new_n5188_;
  assign new_n5190_ = ~new_n5071_ & new_n5182_1_;
  assign new_n5191_ = new_n5187_1_ & new_n5190_;
  assign new_n5192_1_ = ~n4167 & new_n5191_;
  assign new_n5193_ = ~new_n5189_ & ~new_n5192_1_;
  assign new_n5194_ = ~new_n5168_ & new_n5193_;
  assign new_n5195_ = n4167 & new_n5182_1_;
  assign new_n5196_ = ~n4167 & ~new_n5190_;
  assign new_n5197_1_ = ~new_n5195_ & ~new_n5196_;
  assign new_n5198_ = new_n5168_ & new_n5197_1_;
  assign new_n5199_ = ~new_n5194_ & ~new_n5198_;
  assign new_n5200_ = ng2384 & ~new_n5199_;
  assign new_n5201_ = ~new_n5168_ & new_n5200_;
  assign new_n5202_1_ = ~new_n5168_ & ~new_n5201_;
  assign new_n5203_ = new_n5200_ & ~new_n5201_;
  assign new_n5204_ = ~new_n5202_1_ & ~new_n5203_;
  assign new_n5205_ = ng853 & new_n5204_;
  assign new_n5206_ = ~ng414 & ~ng853;
  assign n317 = ~new_n5205_ & ~new_n5206_;
  assign new_n5208_ = ng441 & ng823;
  assign new_n5209_ = ng444 & ng853;
  assign new_n5210_ = ng826 & ng438;
  assign new_n5211_ = ~new_n5208_ & ~new_n5209_;
  assign new_n5212_1_ = ~new_n5210_ & new_n5211_;
  assign new_n5213_ = ~ng449 & ng823;
  assign new_n5214_ = ~ng447 & ng853;
  assign new_n5215_ = ~ng448 & ng826;
  assign new_n5216_ = ~new_n5213_ & ~new_n5214_;
  assign new_n5217_1_ = ~new_n5215_ & new_n5216_;
  assign new_n5218_ = ng432 & ng823;
  assign new_n5219_ = ng853 & ng435;
  assign new_n5220_ = ng826 & ng429;
  assign new_n5221_ = ~new_n5218_ & ~new_n5219_;
  assign new_n5222_1_ = ~new_n5220_ & new_n5221_;
  assign new_n5223_ = ~ng179 & ng823;
  assign new_n5224_ = ng853 & ~ng177;
  assign new_n5225_ = ~ng178 & ng826;
  assign new_n5226_ = ~new_n5223_ & ~new_n5224_;
  assign new_n5227_1_ = ~new_n5225_ & new_n5226_;
  assign new_n5228_ = new_n5180_ & ~new_n5227_1_;
  assign new_n5229_ = new_n5212_1_ & ~new_n5222_1_;
  assign new_n5230_ = new_n5228_ & new_n5229_;
  assign new_n5231_ = ~new_n5212_1_ & new_n5222_1_;
  assign new_n5232_1_ = ~new_n5228_ & new_n5231_;
  assign new_n5233_ = ~new_n5230_ & ~new_n5232_1_;
  assign new_n5234_ = ng2384 & ~new_n5217_1_;
  assign new_n5235_ = ~new_n5233_ & new_n5234_;
  assign new_n5236_ = ~new_n5212_1_ & new_n5235_;
  assign new_n5237_1_ = ~new_n5212_1_ & ~new_n5236_;
  assign new_n5238_ = new_n5235_ & ~new_n5236_;
  assign new_n5239_ = ~new_n5237_1_ & ~new_n5238_;
  assign new_n5240_ = ng823 & new_n5239_;
  assign new_n5241_ = ~ng441 & ~ng823;
  assign n322 = ~new_n5240_ & ~new_n5241_;
  assign new_n5243_ = new_n4790_ & new_n4795_;
  assign new_n5244_ = new_n4795_ & ~new_n4954_;
  assign new_n5245_ = ng2384 & ~new_n4914_;
  assign new_n5246_ = new_n5244_ & new_n5245_;
  assign new_n5247_1_ = new_n4785_ & ~new_n5246_;
  assign new_n5248_ = new_n4877_1_ & new_n4908_;
  assign new_n5249_ = new_n4895_ & new_n5248_;
  assign new_n5250_ = new_n4881_ & new_n5249_;
  assign new_n5251_ = new_n4918_ & new_n4949_;
  assign new_n5252_1_ = new_n4936_ & new_n5251_;
  assign new_n5253_ = new_n4922_1_ & new_n5252_1_;
  assign new_n5254_ = new_n5250_ & new_n5253_;
  assign new_n5255_ = ng2257 & new_n5254_;
  assign new_n5256_ = ~new_n4873_ & new_n5255_;
  assign new_n5257_1_ = ~new_n5071_ & ~new_n5256_;
  assign new_n5258_ = new_n4795_ & ~new_n5257_1_;
  assign new_n5259_ = ~new_n4873_ & ~new_n5254_;
  assign new_n5260_ = ng2257 & new_n5259_;
  assign new_n5261_ = ~new_n4954_ & ~new_n5260_;
  assign new_n5262_1_ = ~new_n4914_ & new_n5261_;
  assign new_n5263_ = ~new_n4795_ & ~new_n5262_1_;
  assign new_n5264_ = ~new_n5258_ & ~new_n5263_;
  assign new_n5265_ = ~new_n4785_ & new_n5264_;
  assign new_n5266_ = ~new_n5247_1_ & ~new_n5265_;
  assign new_n5267_1_ = ~new_n4790_ & new_n5266_;
  assign new_n5268_ = ~new_n5243_ & ~new_n5267_1_;
  assign new_n5269_ = ~new_n4795_ & new_n5268_;
  assign new_n5270_ = ~new_n4795_ & ~new_n5269_;
  assign new_n5271_ = new_n5268_ & ~new_n5269_;
  assign new_n5272_1_ = ~new_n5270_ & ~new_n5271_;
  assign new_n5273_ = ~new_n5080_ & ~new_n5272_1_;
  assign new_n5274_ = ng826 & ~new_n5273_;
  assign new_n5275_ = ~ng318 & ~ng826;
  assign n327 = ~new_n5274_ & ~new_n5275_;
  assign new_n5277_1_ = ng554 & ng1315;
  assign new_n5278_ = ~ng557 & ~ng1315;
  assign n342 = ~new_n5277_1_ & ~new_n5278_;
  assign new_n5280_ = ng853 & ~new_n5136_;
  assign new_n5281_ = ~ng461 & ~ng853;
  assign n352 = ~new_n5280_ & ~new_n5281_;
  assign new_n5283_ = ng608 & ng1312;
  assign new_n5284_ = ng611 & ng1315;
  assign new_n5285_ = ng605 & ng1309;
  assign new_n5286_ = ~new_n5283_ & ~new_n5284_;
  assign new_n5287_1_ = ~new_n5285_ & new_n5286_;
  assign new_n5288_ = ng1312 & ng493;
  assign new_n5289_ = ng1315 & ng496;
  assign new_n5290_ = ng490 & ng1309;
  assign new_n5291_ = ~new_n5288_ & ~new_n5289_;
  assign new_n5292_1_ = ~new_n5290_ & new_n5291_;
  assign new_n5293_ = ~new_n5287_1_ & ~new_n5292_1_;
  assign new_n5294_ = ~ng3013 & ~ng3002;
  assign new_n5295_ = ~ng3006 & new_n5294_;
  assign new_n5296_ = ~ng3024 & new_n5295_;
  assign new_n5297_1_ = ~ng3010 & new_n5296_;
  assign new_n5298_ = ng1312 & ng617;
  assign new_n5299_ = ng1315 & ng620;
  assign new_n5300_ = ng1309 & ng614;
  assign new_n5301_ = ~new_n5298_ & ~new_n5299_;
  assign new_n5302_1_ = ~new_n5300_ & new_n5301_;
  assign new_n5303_ = ng510 & new_n5292_1_;
  assign new_n5304_ = ~new_n5302_1_ & new_n5303_;
  assign new_n5305_1_ = new_n5297_1_ & ~new_n5304_;
  assign n3888 = ~new_n5293_ & ~new_n5305_1_;
  assign new_n5307_ = ng1315 & n3888;
  assign new_n5308_ = ~ng575 & ~new_n5307_;
  assign new_n5309_1_ = ng1312 & ~ng586;
  assign new_n5310_ = ~ng584 & ng1315;
  assign new_n5311_ = ng1309 & ~ng585;
  assign new_n5312_ = ~new_n5309_1_ & ~new_n5310_;
  assign new_n5313_1_ = ~new_n5311_ & new_n5312_;
  assign new_n5314_ = ~ng580 & ng1312;
  assign new_n5315_ = ng1315 & ~ng578;
  assign new_n5316_1_ = ~ng579 & ng1309;
  assign new_n5317_ = ~new_n5314_ & ~new_n5315_;
  assign new_n5318_ = ~new_n5316_1_ & new_n5317_;
  assign new_n5319_ = ~ng577 & ng1312;
  assign new_n5320_ = ~ng575 & ng1315;
  assign new_n5321_1_ = ng1309 & ~ng576;
  assign new_n5322_ = ~new_n5319_ & ~new_n5320_;
  assign new_n5323_ = ~new_n5321_1_ & new_n5322_;
  assign new_n5324_ = pg3229 & ~new_n5323_;
  assign new_n5325_ = new_n5313_1_ & new_n5318_;
  assign new_n5326_1_ = new_n5324_ & new_n5325_;
  assign new_n5327_ = ng1312 & ~ng583;
  assign new_n5328_ = ng1315 & ~ng581;
  assign new_n5329_ = ~ng582 & ng1309;
  assign new_n5330_1_ = ~new_n5327_ & ~new_n5328_;
  assign new_n5331_ = ~new_n5329_ & new_n5330_1_;
  assign new_n5332_ = new_n5324_ & ~new_n5331_;
  assign new_n5333_ = ~new_n5326_1_ & ~new_n5332_;
  assign new_n5334_ = new_n5313_1_ & ~new_n5323_;
  assign new_n5335_1_ = ~pg3229 & new_n5334_;
  assign new_n5336_ = ~new_n5318_ & new_n5331_;
  assign new_n5337_ = ~pg3229 & new_n5336_;
  assign new_n5338_ = pg3229 & ~new_n5313_1_;
  assign new_n5339_ = ~new_n5335_1_ & ~new_n5337_;
  assign new_n5340_1_ = ~new_n5338_ & new_n5339_;
  assign new_n5341_ = new_n5333_ & new_n5340_1_;
  assign new_n5342_ = new_n5307_ & ~new_n5341_;
  assign n362 = ~new_n5308_ & ~new_n5342_;
  assign new_n5344_ = ng590 & ng1312;
  assign new_n5345_1_ = ng593 & ng1315;
  assign new_n5346_ = ng587 & ng1309;
  assign new_n5347_ = ~new_n5344_ & ~new_n5345_1_;
  assign new_n5348_ = ~new_n5346_ & new_n5347_;
  assign new_n5349_ = ng1312 & ng571;
  assign new_n5350_1_ = ng1315 & ng573;
  assign new_n5351_ = ng1309 & ng569;
  assign new_n5352_ = ~new_n5349_ & ~new_n5350_1_;
  assign n1308 = ~new_n5351_ & new_n5352_;
  assign new_n5354_ = ng524 & ~n1308;
  assign new_n5355_1_ = ng185 & new_n5354_;
  assign new_n5356_ = new_n5348_ & ~new_n5355_1_;
  assign new_n5357_ = ng3002 & ng2998;
  assign new_n5358_ = ~ng3006 & new_n5357_;
  assign new_n5359_ = ~ng2993 & new_n5358_;
  assign new_n5360_1_ = ~ng3010 & new_n5359_;
  assign new_n5361_ = ng3024 & new_n5360_1_;
  assign new_n5362_ = ng3013 & new_n5361_;
  assign new_n5363_ = ng3028 & ng3018;
  assign new_n5364_ = new_n5362_ & new_n5363_;
  assign new_n5365_1_ = ~ng3032 & new_n5364_;
  assign new_n5366_ = ~ng3036 & new_n5365_1_;
  assign new_n5367_ = ~new_n5356_ & ~new_n5366_;
  assign new_n5368_ = ng1312 & ~new_n5367_;
  assign new_n5369_1_ = ~ng590 & ~ng1312;
  assign n367 = ~new_n5368_ & ~new_n5369_1_;
  assign new_n5371_ = ng510 & new_n5302_1_;
  assign new_n5372_ = new_n5292_1_ & ~new_n5371_;
  assign new_n5373_1_ = ~new_n5292_1_ & new_n5372_;
  assign new_n5374_ = ~new_n5292_1_ & ~new_n5373_1_;
  assign new_n5375_ = new_n5372_ & ~new_n5373_1_;
  assign new_n5376_ = ~new_n5374_ & ~new_n5375_;
  assign new_n5377_ = ng1309 & ~new_n5376_;
  assign new_n5378_1_ = ~ng490 & ~ng1309;
  assign n372 = ~new_n5377_ & ~new_n5378_1_;
  assign new_n5380_ = ng1312 & ng630;
  assign new_n5381_ = ng1315 & ~ng659;
  assign new_n5382_ = ng640 & new_n5381_;
  assign new_n5383_1_ = ng633 & new_n5382_;
  assign new_n5384_ = ng653 & new_n5383_1_;
  assign new_n5385_ = ~ng646 & new_n5384_;
  assign new_n5386_ = ng646 & ~new_n5384_;
  assign new_n5387_ = ~new_n5385_ & ~new_n5386_;
  assign n377 = ~new_n5380_ & ~new_n5387_;
  assign new_n5389_ = ng525 & ng538;
  assign new_n5390_ = ~ng659 & new_n5389_;
  assign new_n5391_ = ng1312 & new_n5390_;
  assign new_n5392_ = ~ng703 & ~new_n5391_;
  assign new_n5393_1_ = ng633 & new_n5391_;
  assign n382 = ~new_n5392_ & ~new_n5393_1_;
  assign new_n5395_ = ng1309 & new_n5390_;
  assign new_n5396_ = ~ng714 & ~new_n5395_;
  assign new_n5397_ = ng672 & new_n5395_;
  assign n387 = ~new_n5396_ & ~new_n5397_;
  assign new_n5399_ = ng1315 & new_n5390_;
  assign new_n5400_ = ~ng722 & ~new_n5399_;
  assign new_n5401_ = ng686 & new_n5399_;
  assign n392 = ~new_n5400_ & ~new_n5401_;
  assign new_n5403_1_ = ~ng736 & ~new_n5391_;
  assign new_n5404_ = ng1312 & ~ng730;
  assign new_n5405_ = ng1315 & ~ng728;
  assign new_n5406_ = ng1309 & ~ng729;
  assign new_n5407_ = ~new_n5404_ & ~new_n5405_;
  assign new_n5408_1_ = ~new_n5406_ & new_n5407_;
  assign new_n5409_ = ~ng712 & ng1312;
  assign new_n5410_ = ng1315 & ~ng710;
  assign new_n5411_ = ~ng711 & ng1309;
  assign new_n5412_ = ~new_n5409_ & ~new_n5410_;
  assign new_n5413_1_ = ~new_n5411_ & new_n5412_;
  assign new_n5414_ = ~ng660 & ~new_n5413_1_;
  assign new_n5415_ = ~new_n5413_1_ & ~new_n5414_;
  assign new_n5416_ = ~ng660 & ~new_n5414_;
  assign new_n5417_ = ~new_n5415_ & ~new_n5416_;
  assign new_n5418_1_ = ~ng703 & ng1312;
  assign new_n5419_ = ng1315 & ~ng701;
  assign new_n5420_ = ~ng702 & ng1309;
  assign new_n5421_ = ~new_n5418_1_ & ~new_n5419_;
  assign new_n5422_1_ = ~new_n5420_ & new_n5421_;
  assign new_n5423_ = ~ng633 & ~new_n5422_1_;
  assign new_n5424_ = ~new_n5422_1_ & ~new_n5423_;
  assign new_n5425_ = ~ng633 & ~new_n5423_;
  assign new_n5426_ = ~new_n5424_ & ~new_n5425_;
  assign new_n5427_1_ = ng1312 & ~ng706;
  assign new_n5428_ = ng1315 & ~ng704;
  assign new_n5429_ = ~ng705 & ng1309;
  assign new_n5430_ = ~new_n5427_1_ & ~new_n5428_;
  assign new_n5431_1_ = ~new_n5429_ & new_n5430_;
  assign new_n5432_ = ~ng653 & ~new_n5431_1_;
  assign new_n5433_ = ~new_n5431_1_ & ~new_n5432_;
  assign new_n5434_ = ~ng653 & ~new_n5432_;
  assign new_n5435_ = ~new_n5433_ & ~new_n5434_;
  assign new_n5436_1_ = ng1312 & ~ng700;
  assign new_n5437_ = ng1315 & ~ng698;
  assign new_n5438_ = ng1309 & ~ng699;
  assign new_n5439_1_ = ~new_n5436_1_ & ~new_n5437_;
  assign new_n5440_ = ~new_n5438_ & new_n5439_1_;
  assign new_n5441_ = ~ng640 & ~new_n5440_;
  assign new_n5442_ = ~new_n5440_ & ~new_n5441_;
  assign new_n5443_1_ = ~ng640 & ~new_n5441_;
  assign new_n5444_ = ~new_n5442_ & ~new_n5443_1_;
  assign new_n5445_ = ~new_n5426_ & ~new_n5435_;
  assign new_n5446_ = ~new_n5444_ & new_n5445_;
  assign new_n5447_ = ng1312 & ~ng709;
  assign new_n5448_1_ = ng1315 & ~ng707;
  assign new_n5449_ = ng1309 & ~ng708;
  assign new_n5450_ = ~new_n5447_ & ~new_n5448_1_;
  assign new_n5451_ = ~new_n5449_ & new_n5450_;
  assign new_n5452_ = ~ng646 & ~new_n5451_;
  assign new_n5453_1_ = ~new_n5451_ & ~new_n5452_;
  assign new_n5454_ = ~ng646 & ~new_n5452_;
  assign new_n5455_ = ~new_n5453_1_ & ~new_n5454_;
  assign new_n5456_ = ~new_n5417_ & new_n5446_;
  assign new_n5457_ = ~new_n5455_ & new_n5456_;
  assign new_n5458_1_ = ng1312 & ~ng727;
  assign new_n5459_ = ng1315 & ~ng725;
  assign new_n5460_ = ng1309 & ~ng726;
  assign new_n5461_ = ~new_n5458_1_ & ~new_n5459_;
  assign new_n5462_ = ~new_n5460_ & new_n5461_;
  assign new_n5463_1_ = ~ng692 & ~new_n5462_;
  assign new_n5464_ = ~new_n5462_ & ~new_n5463_1_;
  assign new_n5465_ = ~ng692 & ~new_n5463_1_;
  assign new_n5466_ = ~new_n5464_ & ~new_n5465_;
  assign new_n5467_ = ng1312 & ~ng718;
  assign new_n5468_1_ = ng1315 & ~ng716;
  assign new_n5469_ = ng1309 & ~ng717;
  assign new_n5470_ = ~new_n5467_ & ~new_n5468_1_;
  assign new_n5471_ = ~new_n5469_ & new_n5470_;
  assign new_n5472_ = ~ng666 & ~new_n5471_;
  assign new_n5473_1_ = ~new_n5471_ & ~new_n5472_;
  assign new_n5474_ = ~ng666 & ~new_n5472_;
  assign new_n5475_ = ~new_n5473_1_ & ~new_n5474_;
  assign new_n5476_ = ng1312 & ~ng721;
  assign new_n5477_ = ng1315 & ~ng719;
  assign new_n5478_1_ = ~ng720 & ng1309;
  assign new_n5479_ = ~new_n5476_ & ~new_n5477_;
  assign new_n5480_ = ~new_n5478_1_ & new_n5479_;
  assign new_n5481_ = ~ng679 & ~new_n5480_;
  assign new_n5482_ = ~new_n5480_ & ~new_n5481_;
  assign new_n5483_1_ = ~ng679 & ~new_n5481_;
  assign new_n5484_ = ~new_n5482_ & ~new_n5483_1_;
  assign new_n5485_ = ~ng715 & ng1312;
  assign new_n5486_ = ng1315 & ~ng713;
  assign new_n5487_ = ~ng714 & ng1309;
  assign new_n5488_1_ = ~new_n5485_ & ~new_n5486_;
  assign new_n5489_ = ~new_n5487_ & new_n5488_1_;
  assign new_n5490_ = ~ng672 & ~new_n5489_;
  assign new_n5491_ = ~new_n5489_ & ~new_n5490_;
  assign new_n5492_ = ~ng672 & ~new_n5490_;
  assign new_n5493_1_ = ~new_n5491_ & ~new_n5492_;
  assign new_n5494_ = ~new_n5475_ & ~new_n5484_;
  assign new_n5495_ = ~new_n5493_1_ & new_n5494_;
  assign new_n5496_ = ~ng724 & ng1312;
  assign new_n5497_ = ~ng722 & ng1315;
  assign new_n5498_1_ = ~ng723 & ng1309;
  assign new_n5499_ = ~new_n5496_ & ~new_n5497_;
  assign new_n5500_ = ~new_n5498_1_ & new_n5499_;
  assign new_n5501_ = ~ng686 & ~new_n5500_;
  assign new_n5502_ = ~new_n5500_ & ~new_n5501_;
  assign new_n5503_1_ = ~ng686 & ~new_n5501_;
  assign new_n5504_ = ~new_n5502_ & ~new_n5503_1_;
  assign new_n5505_ = ~new_n5466_ & new_n5495_;
  assign new_n5506_ = ~new_n5504_ & new_n5505_;
  assign new_n5507_ = new_n5457_ & new_n5506_;
  assign new_n5508_1_ = ng1312 & ~ng733;
  assign new_n5509_ = ng1315 & ~ng731;
  assign new_n5510_ = ng1309 & ~ng732;
  assign new_n5511_ = ~new_n5508_1_ & ~new_n5509_;
  assign new_n5512_ = ~new_n5510_ & new_n5511_;
  assign new_n5513_1_ = new_n5408_1_ & ~new_n5507_;
  assign new_n5514_ = new_n5512_ & new_n5513_1_;
  assign new_n5515_ = new_n5391_ & ~new_n5514_;
  assign n397 = ~new_n5403_1_ & ~new_n5515_;
  assign new_n5517_1_ = ng826 & ng2257;
  assign new_n5518_ = ~ng821 & ~new_n5517_1_;
  assign new_n5519_ = ng789 & new_n5517_1_;
  assign n402 = ~new_n5518_ & ~new_n5519_;
  assign new_n5521_ = ~ng835 & ~new_n4773_;
  assign new_n5522_1_ = ng801 & new_n4773_;
  assign n407 = ~new_n5521_ & ~new_n5522_1_;
  assign new_n5524_ = ~ng849 & ~new_n4777_1_;
  assign new_n5525_ = ng823 & ~ng864;
  assign new_n5526_1_ = ~ng862 & ng853;
  assign new_n5527_ = ~ng863 & ng826;
  assign new_n5528_ = ~new_n5525_ & ~new_n5526_1_;
  assign new_n5529_ = ~new_n5527_ & new_n5528_;
  assign new_n5530_ = new_n4777_1_ & ~new_n5529_;
  assign n412 = ~new_n5524_ & ~new_n5530_;
  assign new_n5532_ = ~ng2917 & ~ng2920;
  assign new_n5533_ = ng2924 & new_n5532_;
  assign new_n5534_ = ~ng2912 & new_n5533_;
  assign new_n5535_1_ = ng2883 & new_n5125_;
  assign new_n5536_ = ~ng2888 & new_n5535_1_;
  assign n1621 = new_n5534_ & new_n5536_;
  assign new_n5538_ = ng826 & n1621;
  assign new_n5539_ = ~ng863 & ~new_n5538_;
  assign new_n5540_1_ = ng785 & new_n5538_;
  assign n417 = ~new_n5539_ & ~new_n5540_1_;
  assign new_n5542_ = ~ng1003 & ng823;
  assign new_n5543_ = ng853 & ~ng1004;
  assign new_n5544_ = ~ng1002 & ng826;
  assign new_n5545_1_ = ~new_n5542_ & ~new_n5543_;
  assign new_n5546_ = ~new_n5544_ & new_n5545_1_;
  assign new_n5547_ = ~ng1000 & ng823;
  assign new_n5548_ = ~ng1001 & ng853;
  assign new_n5549_1_ = ~ng999 & ng826;
  assign new_n5550_ = ~new_n5547_ & ~new_n5548_;
  assign new_n5551_ = ~new_n5549_1_ & new_n5550_;
  assign new_n5552_ = ng823 & ~ng1006;
  assign new_n5553_1_ = ng853 & ~ng1007;
  assign new_n5554_ = ng826 & ~ng1005;
  assign new_n5555_ = ~new_n5552_ & ~new_n5553_1_;
  assign new_n5556_1_ = ~new_n5554_ & new_n5555_;
  assign new_n5557_ = ~new_n5546_ & new_n5551_;
  assign new_n5558_ = new_n5556_1_ & new_n5557_;
  assign new_n5559_ = new_n5546_ & new_n5551_;
  assign new_n5560_ = new_n5556_1_ & new_n5559_;
  assign new_n5561_1_ = ~new_n5558_ & ~new_n5560_;
  assign new_n5562_ = ng885 & ng823;
  assign new_n5563_ = ng888 & ng853;
  assign new_n5564_ = ng882 & ng826;
  assign new_n5565_ = ~new_n5562_ & ~new_n5563_;
  assign new_n5566_1_ = ~new_n5564_ & new_n5565_;
  assign new_n5567_ = ng823 & ng930;
  assign new_n5568_ = ng853 & ng933;
  assign new_n5569_ = ng826 & ng927;
  assign new_n5570_1_ = ~new_n5567_ & ~new_n5568_;
  assign new_n5571_ = ~new_n5569_ & new_n5570_1_;
  assign new_n5572_ = ng921 & ng823;
  assign new_n5573_ = ng924 & ng853;
  assign new_n5574_ = ng918 & ng826;
  assign new_n5575_1_ = ~new_n5572_ & ~new_n5573_;
  assign new_n5576_ = ~new_n5574_ & new_n5575_1_;
  assign new_n5577_ = ~new_n5566_1_ & ~new_n5571_;
  assign new_n5578_ = ~new_n5576_ & new_n5577_;
  assign new_n5579_ = ng957 & ng823;
  assign new_n5580_1_ = ng853 & ng960;
  assign new_n5581_ = ng954 & ng826;
  assign new_n5582_ = ~new_n5579_ & ~new_n5580_1_;
  assign new_n5583_ = ~new_n5581_ & new_n5582_;
  assign new_n5584_ = ng823 & ng948;
  assign new_n5585_1_ = ng951 & ng853;
  assign new_n5586_ = ng826 & ng945;
  assign new_n5587_ = ~new_n5584_ & ~new_n5585_1_;
  assign new_n5588_ = ~new_n5586_ & new_n5587_;
  assign new_n5589_ = ng894 & ng823;
  assign new_n5590_1_ = ng897 & ng853;
  assign new_n5591_ = ng826 & ng891;
  assign new_n5592_ = ~new_n5589_ & ~new_n5590_1_;
  assign new_n5593_ = ~new_n5591_ & new_n5592_;
  assign new_n5594_ = ng939 & ng823;
  assign new_n5595_1_ = ng942 & ng853;
  assign new_n5596_ = ng936 & ng826;
  assign new_n5597_ = ~new_n5594_ & ~new_n5595_1_;
  assign new_n5598_ = ~new_n5596_ & new_n5597_;
  assign new_n5599_ = ng876 & ng823;
  assign new_n5600_1_ = ng879 & ng853;
  assign new_n5601_ = ng873 & ng826;
  assign new_n5602_ = ~new_n5599_ & ~new_n5600_1_;
  assign new_n5603_ = ~new_n5601_ & new_n5602_;
  assign new_n5604_ = new_n5593_ & new_n5598_;
  assign new_n5605_1_ = new_n5603_ & new_n5604_;
  assign new_n5606_ = ng823 & ng903;
  assign new_n5607_ = ng853 & ng906;
  assign new_n5608_ = ng900 & ng826;
  assign new_n5609_ = ~new_n5606_ & ~new_n5607_;
  assign new_n5610_1_ = ~new_n5608_ & new_n5609_;
  assign new_n5611_ = new_n5588_ & new_n5605_1_;
  assign new_n5612_ = new_n5610_1_ & new_n5611_;
  assign new_n5613_ = ng912 & ng823;
  assign new_n5614_ = ng915 & ng853;
  assign new_n5615_1_ = ng909 & ng826;
  assign new_n5616_ = ~new_n5613_ & ~new_n5614_;
  assign new_n5617_ = ~new_n5615_1_ & new_n5616_;
  assign new_n5618_ = new_n5578_ & ~new_n5583_;
  assign new_n5619_ = new_n5612_ & new_n5618_;
  assign new_n5620_1_ = ~new_n5617_ & new_n5619_;
  assign new_n5621_ = new_n5558_ & new_n5620_1_;
  assign new_n5622_ = new_n5566_1_ & new_n5571_;
  assign new_n5623_ = new_n5576_ & new_n5622_;
  assign new_n5624_ = new_n5583_ & new_n5623_;
  assign new_n5625_1_ = new_n5612_ & new_n5624_;
  assign new_n5626_ = new_n5617_ & new_n5625_1_;
  assign new_n5627_ = ~new_n5558_ & new_n5626_;
  assign new_n5628_ = ~new_n5621_ & ~new_n5627_;
  assign new_n5629_ = ~new_n5561_1_ & ~new_n5628_;
  assign new_n5630_1_ = ~ng858 & ng823;
  assign new_n5631_ = ~ng856 & ng853;
  assign new_n5632_ = ng826 & ~ng857;
  assign new_n5633_ = ~new_n5630_1_ & ~new_n5631_;
  assign new_n5634_1_ = ~new_n5632_ & new_n5633_;
  assign new_n5635_ = ng789 & ~new_n5576_;
  assign new_n5636_ = ng789 & ~new_n5635_;
  assign new_n5637_ = ~new_n5576_ & ~new_n5635_;
  assign new_n5638_ = ~new_n5636_ & ~new_n5637_;
  assign new_n5639_1_ = ng813 & ~new_n5588_;
  assign new_n5640_ = ng813 & ~new_n5639_1_;
  assign new_n5641_ = ~new_n5588_ & ~new_n5639_1_;
  assign new_n5642_ = ~new_n5640_ & ~new_n5641_;
  assign new_n5643_ = new_n5638_ & new_n5642_;
  assign new_n5644_1_ = ng797 & ~new_n5571_;
  assign new_n5645_ = ng797 & ~new_n5644_1_;
  assign new_n5646_ = ~new_n5571_ & ~new_n5644_1_;
  assign new_n5647_ = ~new_n5645_ & ~new_n5646_;
  assign new_n5648_ = ~ng861 & ng823;
  assign new_n5649_1_ = ~ng859 & ng853;
  assign new_n5650_ = ~ng860 & ng826;
  assign new_n5651_ = ~new_n5648_ & ~new_n5649_1_;
  assign new_n5652_ = ~new_n5650_ & new_n5651_;
  assign new_n5653_ = ~new_n5583_ & ~new_n5652_;
  assign new_n5654_1_ = ~new_n5652_ & ~new_n5653_;
  assign new_n5655_ = ~new_n5583_ & ~new_n5653_;
  assign new_n5656_ = ~new_n5654_1_ & ~new_n5655_;
  assign new_n5657_ = new_n5647_ & new_n5656_;
  assign new_n5658_ = ng805 & ~new_n5598_;
  assign new_n5659_1_ = ng805 & ~new_n5658_;
  assign new_n5660_ = ~new_n5598_ & ~new_n5658_;
  assign new_n5661_ = ~new_n5659_1_ & ~new_n5660_;
  assign new_n5662_ = ~new_n5643_ & ~new_n5657_;
  assign new_n5663_ = ~new_n5661_ & new_n5662_;
  assign new_n5664_1_ = new_n5642_ & new_n5661_;
  assign new_n5665_ = new_n5638_ & new_n5647_;
  assign new_n5666_ = ~new_n5664_1_ & ~new_n5665_;
  assign new_n5667_ = ~new_n5656_ & new_n5666_;
  assign new_n5668_ = new_n5642_ & new_n5656_;
  assign new_n5669_1_ = new_n5647_ & new_n5661_;
  assign new_n5670_ = ~new_n5668_ & ~new_n5669_1_;
  assign new_n5671_ = ~new_n5638_ & new_n5670_;
  assign new_n5672_ = ~new_n5663_ & ~new_n5667_;
  assign new_n5673_ = ~new_n5671_ & new_n5672_;
  assign new_n5674_1_ = ng2257 & ~new_n5634_1_;
  assign new_n5675_ = ~new_n5673_ & new_n5674_1_;
  assign new_n5676_ = ng785 & ~new_n5603_;
  assign new_n5677_ = ng785 & ~new_n5676_;
  assign new_n5678_ = ~new_n5603_ & ~new_n5676_;
  assign new_n5679_1_ = ~new_n5677_ & ~new_n5678_;
  assign new_n5680_ = ng809 & ~new_n5610_1_;
  assign new_n5681_ = ng809 & ~new_n5680_;
  assign new_n5682_ = ~new_n5610_1_ & ~new_n5680_;
  assign new_n5683_ = ~new_n5681_ & ~new_n5682_;
  assign new_n5684_1_ = new_n5679_1_ & new_n5683_;
  assign new_n5685_ = ng793 & ~new_n5566_1_;
  assign new_n5686_ = ng793 & ~new_n5685_;
  assign new_n5687_ = ~new_n5566_1_ & ~new_n5685_;
  assign new_n5688_ = ~new_n5686_ & ~new_n5687_;
  assign new_n5689_1_ = ~new_n5529_ & ~new_n5617_;
  assign new_n5690_ = ~new_n5529_ & ~new_n5689_1_;
  assign new_n5691_ = ~new_n5617_ & ~new_n5689_1_;
  assign new_n5692_ = ~new_n5690_ & ~new_n5691_;
  assign new_n5693_ = new_n5688_ & new_n5692_;
  assign new_n5694_1_ = ng801 & ~new_n5593_;
  assign new_n5695_ = ng801 & ~new_n5694_1_;
  assign new_n5696_ = ~new_n5593_ & ~new_n5694_1_;
  assign new_n5697_ = ~new_n5695_ & ~new_n5696_;
  assign new_n5698_ = ~new_n5684_1_ & ~new_n5693_;
  assign new_n5699_1_ = ~new_n5697_ & new_n5698_;
  assign new_n5700_ = new_n5683_ & new_n5697_;
  assign new_n5701_ = new_n5679_1_ & new_n5688_;
  assign new_n5702_ = ~new_n5700_ & ~new_n5701_;
  assign new_n5703_ = ~new_n5692_ & new_n5702_;
  assign new_n5704_1_ = new_n5683_ & new_n5692_;
  assign new_n5705_ = new_n5688_ & new_n5697_;
  assign new_n5706_ = ~new_n5704_1_ & ~new_n5705_;
  assign new_n5707_ = ~new_n5679_1_ & new_n5706_;
  assign new_n5708_ = ~new_n5699_1_ & ~new_n5703_;
  assign new_n5709_1_ = ~new_n5707_ & new_n5708_;
  assign new_n5710_ = new_n5674_1_ & ~new_n5709_1_;
  assign new_n5711_ = ~new_n5675_ & ~new_n5710_;
  assign new_n5712_ = ~ng852 & ng823;
  assign new_n5713_ = ~ng850 & ng853;
  assign new_n5714_1_ = ng826 & ~ng851;
  assign new_n5715_ = ~new_n5712_ & ~new_n5713_;
  assign new_n5716_ = ~new_n5714_1_ & new_n5715_;
  assign new_n5717_ = ~new_n5652_ & ~new_n5716_;
  assign new_n5718_ = ~new_n5716_ & ~new_n5717_;
  assign new_n5719_1_ = ~new_n5652_ & ~new_n5717_;
  assign new_n5720_ = ~new_n5718_ & ~new_n5719_1_;
  assign new_n5721_ = ng823 & ~ng843;
  assign new_n5722_ = ng853 & ~ng841;
  assign new_n5723_ = ng826 & ~ng842;
  assign new_n5724_1_ = ~new_n5721_ & ~new_n5722_;
  assign new_n5725_ = ~new_n5723_ & new_n5724_1_;
  assign new_n5726_ = ng809 & ~new_n5725_;
  assign new_n5727_ = ~new_n5725_ & ~new_n5726_;
  assign new_n5728_ = ng809 & ~new_n5726_;
  assign new_n5729_1_ = ~new_n5727_ & ~new_n5728_;
  assign new_n5730_ = ~ng846 & ng823;
  assign new_n5731_ = ~ng844 & ng853;
  assign new_n5732_ = ng826 & ~ng845;
  assign new_n5733_ = ~new_n5730_ & ~new_n5731_;
  assign new_n5734_1_ = ~new_n5732_ & new_n5733_;
  assign new_n5735_ = ng813 & ~new_n5734_1_;
  assign new_n5736_ = ~new_n5734_1_ & ~new_n5735_;
  assign new_n5737_ = ng813 & ~new_n5735_;
  assign new_n5738_1_ = ~new_n5736_ & ~new_n5737_;
  assign new_n5739_ = ~ng840 & ng823;
  assign new_n5740_ = ~ng838 & ng853;
  assign new_n5741_ = ~ng839 & ng826;
  assign new_n5742_ = ~new_n5739_ & ~new_n5740_;
  assign new_n5743_1_ = ~new_n5741_ & new_n5742_;
  assign new_n5744_ = ng805 & ~new_n5743_1_;
  assign new_n5745_ = ~new_n5743_1_ & ~new_n5744_;
  assign new_n5746_ = ng805 & ~new_n5744_;
  assign new_n5747_ = ~new_n5745_ & ~new_n5746_;
  assign new_n5748_1_ = new_n5729_1_ & new_n5738_1_;
  assign new_n5749_ = new_n5747_ & new_n5748_1_;
  assign new_n5750_ = ~ng849 & ng823;
  assign new_n5751_ = ~ng847 & ng853;
  assign new_n5752_ = ~ng848 & ng826;
  assign new_n5753_1_ = ~new_n5750_ & ~new_n5751_;
  assign new_n5754_ = ~new_n5752_ & new_n5753_1_;
  assign new_n5755_ = ~new_n5529_ & ~new_n5754_;
  assign new_n5756_ = ~new_n5754_ & ~new_n5755_;
  assign new_n5757_ = ~new_n5529_ & ~new_n5755_;
  assign new_n5758_1_ = ~new_n5756_ & ~new_n5757_;
  assign new_n5759_ = new_n5720_ & new_n5749_;
  assign new_n5760_ = new_n5758_1_ & new_n5759_;
  assign new_n5761_ = ~ng837 & ng823;
  assign new_n5762_ = ~ng835 & ng853;
  assign new_n5763_1_ = ~ng836 & ng826;
  assign new_n5764_ = ~new_n5761_ & ~new_n5762_;
  assign new_n5765_ = ~new_n5763_1_ & new_n5764_;
  assign new_n5766_ = ng801 & ~new_n5765_;
  assign new_n5767_ = ~new_n5765_ & ~new_n5766_;
  assign new_n5768_1_ = ng801 & ~new_n5766_;
  assign new_n5769_ = ~new_n5767_ & ~new_n5768_1_;
  assign new_n5770_ = ~ng822 & ng823;
  assign new_n5771_ = ~ng820 & ng853;
  assign new_n5772_ = ~ng821 & ng826;
  assign new_n5773_1_ = ~new_n5770_ & ~new_n5771_;
  assign new_n5774_ = ~new_n5772_ & new_n5773_1_;
  assign new_n5775_ = ng789 & ~new_n5774_;
  assign new_n5776_ = ~new_n5774_ & ~new_n5775_;
  assign new_n5777_ = ng789 & ~new_n5775_;
  assign new_n5778_1_ = ~new_n5776_ & ~new_n5777_;
  assign new_n5779_ = ~ng831 & ng823;
  assign new_n5780_ = ng853 & ~ng829;
  assign new_n5781_ = ~ng830 & ng826;
  assign new_n5782_ = ~new_n5779_ & ~new_n5780_;
  assign new_n5783_1_ = ~new_n5781_ & new_n5782_;
  assign new_n5784_ = ng793 & ~new_n5783_1_;
  assign new_n5785_ = ~new_n5783_1_ & ~new_n5784_;
  assign new_n5786_ = ng793 & ~new_n5784_;
  assign new_n5787_ = ~new_n5785_ & ~new_n5786_;
  assign new_n5788_1_ = ng823 & ~ng819;
  assign new_n5789_ = ~ng817 & ng853;
  assign new_n5790_ = ng826 & ~ng818;
  assign new_n5791_ = ~new_n5788_1_ & ~new_n5789_;
  assign new_n5792_ = ~new_n5790_ & new_n5791_;
  assign new_n5793_1_ = ng785 & ~new_n5792_;
  assign new_n5794_ = ~new_n5792_ & ~new_n5793_1_;
  assign new_n5795_ = ng785 & ~new_n5793_1_;
  assign new_n5796_ = ~new_n5794_ & ~new_n5795_;
  assign new_n5797_ = new_n5778_1_ & new_n5787_;
  assign new_n5798_1_ = new_n5796_ & new_n5797_;
  assign new_n5799_ = ~ng834 & ng823;
  assign new_n5800_ = ng853 & ~ng832;
  assign new_n5801_ = ng826 & ~ng833;
  assign new_n5802_ = ~new_n5799_ & ~new_n5800_;
  assign new_n5803_1_ = ~new_n5801_ & new_n5802_;
  assign new_n5804_ = ng797 & ~new_n5803_1_;
  assign new_n5805_ = ~new_n5803_1_ & ~new_n5804_;
  assign new_n5806_ = ng797 & ~new_n5804_;
  assign new_n5807_ = ~new_n5805_ & ~new_n5806_;
  assign new_n5808_1_ = new_n5769_ & new_n5798_1_;
  assign new_n5809_ = new_n5807_ & new_n5808_1_;
  assign new_n5810_ = new_n5760_ & new_n5809_;
  assign new_n5811_ = ~new_n5634_1_ & new_n5711_;
  assign new_n5812_ = ng2257 & new_n5810_;
  assign new_n5813_1_ = new_n5811_ & new_n5812_;
  assign new_n5814_ = ~ng1010 & ng823;
  assign new_n5815_ = ~ng1008 & ng853;
  assign new_n5816_ = ~ng1009 & ng826;
  assign new_n5817_ = ~new_n5814_ & ~new_n5815_;
  assign new_n5818_1_ = ~new_n5816_ & new_n5817_;
  assign new_n5819_ = new_n5546_ & ~new_n5551_;
  assign new_n5820_ = new_n5556_1_ & new_n5819_;
  assign new_n5821_ = new_n5813_1_ & ~new_n5818_1_;
  assign new_n5822_ = new_n5820_ & new_n5821_;
  assign new_n5823_1_ = new_n5674_1_ & new_n5810_;
  assign new_n5824_ = ~new_n5556_1_ & new_n5819_;
  assign new_n5825_ = ~new_n5818_1_ & new_n5823_1_;
  assign new_n5826_ = new_n5824_ & new_n5825_;
  assign new_n5827_ = ng2257 & new_n5634_1_;
  assign new_n5828_1_ = ~new_n5551_ & new_n5827_;
  assign new_n5829_ = ~new_n5822_ & ~new_n5826_;
  assign new_n5830_ = ~new_n5828_1_ & new_n5829_;
  assign new_n5831_ = ~ng1091 & ng823;
  assign new_n5832_ = ~ng1089 & ng853;
  assign new_n5833_1_ = ~ng1090 & ng826;
  assign new_n5834_ = ~new_n5831_ & ~new_n5832_;
  assign new_n5835_ = ~new_n5833_1_ & new_n5834_;
  assign new_n5836_ = new_n5823_1_ & ~new_n5835_;
  assign new_n5837_ = new_n5830_ & ~new_n5836_;
  assign new_n5838_1_ = ~new_n5629_ & new_n5837_;
  assign new_n5839_ = new_n5629_ & new_n5837_;
  assign new_n5840_ = ng789 & ~new_n5839_;
  assign new_n5841_ = ~new_n5558_ & new_n5839_;
  assign new_n5842_ = ~new_n5840_ & ~new_n5841_;
  assign new_n5843_1_ = ~new_n5838_1_ & new_n5842_;
  assign new_n5844_ = new_n5558_ & new_n5603_;
  assign new_n5845_ = ~new_n5558_ & ~new_n5603_;
  assign new_n5846_ = ~new_n5844_ & ~new_n5845_;
  assign new_n5847_ = ~new_n5561_1_ & new_n5846_;
  assign new_n5848_1_ = ~new_n5576_ & ~new_n5847_;
  assign new_n5849_ = new_n5576_ & new_n5847_;
  assign new_n5850_ = ~new_n5848_1_ & ~new_n5849_;
  assign new_n5851_ = new_n5838_1_ & new_n5850_;
  assign new_n5852_ = ~new_n5843_1_ & ~new_n5851_;
  assign new_n5853_1_ = ng853 & ~new_n5852_;
  assign new_n5854_ = ~ng924 & ~ng853;
  assign n422 = ~new_n5853_1_ & ~new_n5854_;
  assign new_n5856_ = ng805 & ~new_n5839_;
  assign new_n5857_ = ~new_n5838_1_ & ~new_n5856_;
  assign new_n5858_1_ = new_n5558_ & ~new_n5593_;
  assign new_n5859_ = ~new_n5558_ & new_n5593_;
  assign new_n5860_ = ~new_n5858_1_ & ~new_n5859_;
  assign new_n5861_ = new_n5558_ & ~new_n5576_;
  assign new_n5862_ = ~new_n5558_ & new_n5576_;
  assign new_n5863_1_ = ~new_n5861_ & ~new_n5862_;
  assign new_n5864_ = new_n5847_ & ~new_n5863_1_;
  assign new_n5865_ = new_n5558_ & ~new_n5571_;
  assign new_n5866_ = ~new_n5558_ & new_n5571_;
  assign new_n5867_ = ~new_n5865_ & ~new_n5866_;
  assign new_n5868_1_ = new_n5558_ & ~new_n5566_1_;
  assign new_n5869_ = ~new_n5558_ & new_n5566_1_;
  assign new_n5870_ = ~new_n5868_1_ & ~new_n5869_;
  assign new_n5871_ = ~new_n5867_ & ~new_n5870_;
  assign new_n5872_ = new_n5864_ & new_n5871_;
  assign new_n5873_1_ = ~new_n5860_ & new_n5872_;
  assign new_n5874_ = new_n5598_ & new_n5873_1_;
  assign new_n5875_ = ~new_n5598_ & ~new_n5873_1_;
  assign new_n5876_ = ~new_n5874_ & ~new_n5875_;
  assign new_n5877_ = new_n5838_1_ & new_n5876_;
  assign new_n5878_1_ = ~new_n5857_ & ~new_n5877_;
  assign new_n5879_ = ng823 & ~new_n5878_1_;
  assign new_n5880_ = ~ng939 & ~ng823;
  assign n427 = ~new_n5879_ & ~new_n5880_;
  assign new_n5882_ = ~new_n5652_ & ~new_n5839_;
  assign new_n5883_1_ = ~new_n5841_ & ~new_n5882_;
  assign new_n5884_ = ~new_n5838_1_ & new_n5883_1_;
  assign new_n5885_ = new_n5558_ & ~new_n5617_;
  assign new_n5886_ = ~new_n5558_ & new_n5617_;
  assign new_n5887_ = ~new_n5885_ & ~new_n5886_;
  assign new_n5888_1_ = new_n5558_ & ~new_n5598_;
  assign new_n5889_ = ~new_n5558_ & new_n5598_;
  assign new_n5890_ = ~new_n5888_1_ & ~new_n5889_;
  assign new_n5891_ = ~new_n5860_ & ~new_n5890_;
  assign new_n5892_ = new_n5558_ & ~new_n5588_;
  assign new_n5893_1_ = ~new_n5558_ & new_n5588_;
  assign new_n5894_ = ~new_n5892_ & ~new_n5893_1_;
  assign new_n5895_ = new_n5558_ & ~new_n5610_1_;
  assign new_n5896_ = ~new_n5558_ & new_n5610_1_;
  assign new_n5897_ = ~new_n5895_ & ~new_n5896_;
  assign new_n5898_1_ = ~new_n5894_ & ~new_n5897_;
  assign new_n5899_ = new_n5864_ & new_n5891_;
  assign new_n5900_ = new_n5871_ & new_n5898_1_;
  assign new_n5901_ = new_n5899_ & new_n5900_;
  assign new_n5902_ = ~new_n5887_ & new_n5901_;
  assign new_n5903_1_ = new_n5583_ & new_n5902_;
  assign new_n5904_ = ~new_n5583_ & ~new_n5902_;
  assign new_n5905_ = ~new_n5903_1_ & ~new_n5904_;
  assign new_n5906_ = new_n5838_1_ & new_n5905_;
  assign new_n5907_ = ~new_n5884_ & ~new_n5906_;
  assign new_n5908_1_ = ng826 & ~new_n5907_;
  assign new_n5909_ = ~ng954 & ~ng826;
  assign n432 = ~new_n5908_1_ & ~new_n5909_;
  assign new_n5911_ = ng780 & new_n5128_;
  assign new_n5912_ = ng776 & new_n5911_;
  assign new_n5913_1_ = ng771 & new_n5912_;
  assign new_n5914_ = ng767 & new_n5913_1_;
  assign new_n5915_ = ng762 & new_n5914_;
  assign new_n5916_ = ng758 & new_n5915_;
  assign new_n5917_ = ng753 & new_n5916_;
  assign new_n5918_1_ = ng749 & new_n5917_;
  assign new_n5919_ = ~ng744 & new_n5918_1_;
  assign new_n5920_ = ng744 & ~new_n5918_1_;
  assign new_n5921_ = ~new_n5919_ & ~new_n5920_;
  assign n437 = ~new_n5127_1_ & ~new_n5921_;
  assign new_n5923_1_ = new_n5125_ & ~new_n5560_;
  assign new_n5924_ = ~new_n5556_1_ & new_n5557_;
  assign new_n5925_ = ~new_n5923_1_ & ~new_n5924_;
  assign new_n5926_ = ng826 & new_n5925_;
  assign new_n5927_ = ~ng1085 & ~new_n5926_;
  assign new_n5928_1_ = ng823 & ~ng1030;
  assign new_n5929_ = ng853 & ~ng1033;
  assign new_n5930_ = ng826 & ~ng1041;
  assign new_n5931_ = ~new_n5928_1_ & ~new_n5929_;
  assign new_n5932_ = ~new_n5930_ & new_n5931_;
  assign new_n5933_1_ = ng823 & ~ng1060;
  assign new_n5934_ = ng853 & ~ng1063;
  assign new_n5935_ = ng826 & ~ng1071;
  assign new_n5936_ = ~new_n5933_1_ & ~new_n5934_;
  assign new_n5937_ = ~new_n5935_ & new_n5936_;
  assign new_n5938_1_ = ~ng1045 & ng823;
  assign new_n5939_ = ng853 & ~ng1048;
  assign new_n5940_ = ng826 & ~ng1056;
  assign new_n5941_ = ~new_n5938_1_ & ~new_n5939_;
  assign new_n5942_ = ~new_n5940_ & new_n5941_;
  assign new_n5943_1_ = new_n5937_ & new_n5942_;
  assign new_n5944_ = ~pg3229 & ~new_n5932_;
  assign new_n5945_ = new_n5943_1_ & new_n5944_;
  assign new_n5946_ = pg3229 & new_n5932_;
  assign new_n5947_ = new_n5943_1_ & new_n5946_;
  assign new_n5948_1_ = ~new_n5945_ & ~new_n5947_;
  assign new_n5949_ = new_n5926_ & ~new_n5948_1_;
  assign n442 = ~new_n5927_ & ~new_n5949_;
  assign new_n5951_ = ~ng1115 & ng823;
  assign new_n5952_ = ~ng1113 & ng853;
  assign new_n5953_1_ = ng826 & ~ng1114;
  assign new_n5954_ = ~new_n5951_ & ~new_n5952_;
  assign new_n5955_ = ~new_n5953_1_ & new_n5954_;
  assign new_n5956_ = ng1107 & ng823;
  assign new_n5957_ = ng853 & ng1110;
  assign new_n5958_1_ = ng826 & ng1104;
  assign new_n5959_ = ~new_n5956_ & ~new_n5957_;
  assign n953 = new_n5958_1_ | ~new_n5959_;
  assign new_n5961_ = ng805 & ng813;
  assign new_n5962_1_ = ng809 & new_n5961_;
  assign new_n5963_ = ng801 & new_n5962_1_;
  assign new_n5964_ = ng789 & ng797;
  assign new_n5965_ = ng793 & new_n5964_;
  assign new_n5966_ = ng785 & new_n5965_;
  assign new_n5967_1_ = new_n5963_ & new_n5966_;
  assign new_n5968_ = ~new_n5529_ & ~new_n5652_;
  assign new_n5969_ = new_n5967_1_ & new_n5968_;
  assign new_n5970_ = n953 & ~new_n5969_;
  assign new_n5971_ = ~new_n5827_ & new_n5969_;
  assign new_n5972_1_ = ~n953 & new_n5971_;
  assign new_n5973_ = ~new_n5970_ & ~new_n5972_1_;
  assign new_n5974_ = ng1098 & ng823;
  assign new_n5975_ = ng1101 & ng853;
  assign new_n5976_ = ng1095 & ng826;
  assign new_n5977_1_ = ~new_n5974_ & ~new_n5975_;
  assign new_n5978_ = ~new_n5976_ & new_n5977_1_;
  assign new_n5979_ = new_n5955_ & ~new_n5973_;
  assign new_n5980_ = ~new_n5978_ & new_n5979_;
  assign new_n5981_ = ng2384 & new_n5980_;
  assign new_n5982_1_ = ~new_n5973_ & new_n5978_;
  assign new_n5983_ = ng2384 & new_n5982_1_;
  assign new_n5984_ = ~new_n5981_ & ~new_n5983_;
  assign new_n5985_ = ng853 & ~new_n5984_;
  assign new_n5986_ = ~ng1113 & ~new_n5985_;
  assign new_n5987_1_ = new_n5981_ & new_n5985_;
  assign n447 = ~new_n5986_ & ~new_n5987_1_;
  assign new_n5989_ = ~new_n5546_ & new_n5556_1_;
  assign new_n5990_ = new_n5551_ & new_n5989_;
  assign new_n5991_ = new_n5546_ & ~new_n5556_1_;
  assign new_n5992_1_ = ~new_n5711_ & ~new_n5991_;
  assign new_n5993_ = ~new_n5551_ & ~new_n5992_1_;
  assign new_n5994_ = ~new_n5990_ & ~new_n5993_;
  assign new_n5995_ = ~new_n5551_ & new_n5994_;
  assign new_n5996_ = ~new_n5551_ & ~new_n5995_;
  assign new_n5997_1_ = new_n5994_ & ~new_n5995_;
  assign new_n5998_ = ~new_n5996_ & ~new_n5997_1_;
  assign new_n5999_ = ~new_n5836_ & new_n5998_;
  assign new_n6000_ = ng823 & ~new_n5999_;
  assign new_n6001_ = ~ng1000 & ~ng823;
  assign n452 = ~new_n6000_ & ~new_n6001_;
  assign new_n6003_ = ng2384 & ng826;
  assign new_n6004_ = ~ng1090 & ~new_n6003_;
  assign new_n6005_ = new_n5823_1_ & new_n5835_;
  assign new_n6006_ = new_n6003_ & new_n6005_;
  assign n457 = ~new_n6004_ & ~new_n6006_;
  assign new_n6008_ = ~ng986 & ng985;
  assign new_n6009_ = ng298 & ~ng299;
  assign new_n6010_ = ng305 & ~ng823;
  assign new_n6011_ = ng299 & ~new_n6010_;
  assign n4507 = ~new_n6009_ & ~new_n6011_;
  assign new_n6013_ = ng823 & n4507;
  assign new_n6014_ = ng992 & ~ng823;
  assign new_n6015_ = ~new_n6013_ & ~new_n6014_;
  assign new_n6016_ = ng986 & new_n6015_;
  assign n467 = ~new_n6008_ & ~new_n6016_;
  assign new_n6018_ = ng823 & ng1128;
  assign new_n6019_ = ng853 & ng1131;
  assign new_n6020_ = ng1125 & ng826;
  assign new_n6021_ = ~new_n6018_ & ~new_n6019_;
  assign new_n6022_1_ = ~new_n6020_ & new_n6021_;
  assign new_n6023_ = ng826 & new_n6022_1_;
  assign new_n6024_ = ~ng1173 & ~ng826;
  assign n487 = ~new_n6023_ & ~new_n6024_;
  assign new_n6026_ = ng853 & n953;
  assign new_n6027_1_ = ~ng1151 & ~ng853;
  assign n492 = ~new_n6026_ & ~new_n6027_1_;
  assign new_n6029_ = ng1312 & ng1294;
  assign new_n6030_ = ng1315 & ng1297;
  assign new_n6031_ = ng1291 & ng1309;
  assign new_n6032_1_ = ~new_n6029_ & ~new_n6030_;
  assign new_n6033_ = ~new_n6031_ & new_n6032_1_;
  assign new_n6034_ = ng1312 & ng1180;
  assign new_n6035_ = ng1315 & ng1183;
  assign new_n6036_ = ng1177 & ng1309;
  assign new_n6037_1_ = ~new_n6034_ & ~new_n6035_;
  assign new_n6038_ = ~new_n6036_ & new_n6037_1_;
  assign new_n6039_ = ~new_n6033_ & ~new_n6038_;
  assign new_n6040_ = ng1303 & ng1312;
  assign new_n6041_ = ng1306 & ng1315;
  assign new_n6042_1_ = ng1300 & ng1309;
  assign new_n6043_ = ~new_n6040_ & ~new_n6041_;
  assign new_n6044_ = ~new_n6042_1_ & new_n6043_;
  assign new_n6045_ = ng1196 & new_n6038_;
  assign new_n6046_ = ~new_n6044_ & new_n6045_;
  assign new_n6047_1_ = new_n5297_1_ & ~new_n6046_;
  assign n2976 = ~new_n6039_ & ~new_n6047_1_;
  assign new_n6049_ = ng1315 & n2976;
  assign new_n6050_ = ~ng1267 & ~new_n6049_;
  assign new_n6051_ = ng1312 & ~ng1263;
  assign new_n6052_1_ = ng1315 & ~ng1261;
  assign new_n6053_ = ~ng1262 & ng1309;
  assign new_n6054_ = ~new_n6051_ & ~new_n6052_1_;
  assign new_n6055_ = ~new_n6053_ & new_n6054_;
  assign new_n6056_ = ng1312 & ~ng1272;
  assign new_n6057_1_ = ng1315 & ~ng1270;
  assign new_n6058_ = ~ng1271 & ng1309;
  assign new_n6059_ = ~new_n6056_ & ~new_n6057_1_;
  assign new_n6060_ = ~new_n6058_ & new_n6059_;
  assign new_n6061_ = ng1312 & ~ng1266;
  assign new_n6062_1_ = ng1315 & ~ng1264;
  assign new_n6063_ = ng1309 & ~ng1265;
  assign new_n6064_ = ~new_n6061_ & ~new_n6062_1_;
  assign new_n6065_ = ~new_n6063_ & new_n6064_;
  assign new_n6066_ = new_n6060_ & new_n6065_;
  assign new_n6067_1_ = pg3229 & ~new_n6055_;
  assign new_n6068_ = new_n6066_ & new_n6067_1_;
  assign new_n6069_ = ~pg3229 & new_n6055_;
  assign new_n6070_ = new_n6066_ & new_n6069_;
  assign new_n6071_ = ~new_n6068_ & ~new_n6070_;
  assign new_n6072_1_ = ~new_n6055_ & ~new_n6065_;
  assign new_n6073_ = ~pg3229 & new_n6072_1_;
  assign new_n6074_ = new_n6055_ & ~new_n6065_;
  assign new_n6075_ = pg3229 & new_n6074_;
  assign new_n6076_ = ~new_n6073_ & ~new_n6075_;
  assign new_n6077_1_ = new_n6071_ & new_n6076_;
  assign new_n6078_ = new_n6049_ & ~new_n6077_1_;
  assign n502 = ~new_n6050_ & ~new_n6078_;
  assign new_n6080_ = ng1312 & ng1068;
  assign new_n6081_ = ng1315 & ng1070;
  assign new_n6082_1_ = ng1309 & ng1066;
  assign new_n6083_ = ~new_n6080_ & ~new_n6081_;
  assign new_n6084_ = ~new_n6082_1_ & new_n6083_;
  assign new_n6085_ = ng1053 & ng1312;
  assign new_n6086_ = ng1055 & ng1315;
  assign new_n6087_1_ = ng1051 & ng1309;
  assign new_n6088_ = ~new_n6085_ & ~new_n6086_;
  assign new_n6089_ = ~new_n6087_1_ & new_n6088_;
  assign new_n6090_ = ~new_n6065_ & ~new_n6084_;
  assign new_n6091_ = new_n6089_ & new_n6090_;
  assign new_n6092_1_ = new_n6055_ & new_n6091_;
  assign new_n6093_ = ~ng1269 & ng1312;
  assign new_n6094_ = ~ng1267 & ng1315;
  assign new_n6095_ = ~ng1268 & ng1309;
  assign new_n6096_ = ~new_n6093_ & ~new_n6094_;
  assign new_n6097_1_ = ~new_n6095_ & new_n6096_;
  assign new_n6098_ = ng1312 & ng1038;
  assign new_n6099_ = ng1315 & ng1040;
  assign new_n6100_ = ng1036 & ng1309;
  assign new_n6101_ = ~new_n6098_ & ~new_n6099_;
  assign new_n6102_1_ = ~new_n6100_ & new_n6101_;
  assign new_n6103_ = new_n6089_ & new_n6097_1_;
  assign new_n6104_ = new_n6102_1_ & new_n6103_;
  assign new_n6105_ = ~new_n6065_ & new_n6104_;
  assign new_n6106_ = ng1083 & ng1312;
  assign new_n6107_1_ = ng1315 & ng1011;
  assign new_n6108_ = ng1081 & ng1309;
  assign new_n6109_ = ~new_n6106_ & ~new_n6107_1_;
  assign new_n6110_ = ~new_n6108_ & new_n6109_;
  assign new_n6111_ = new_n6065_ & new_n6110_;
  assign new_n6112_1_ = new_n6097_1_ & new_n6111_;
  assign new_n6113_ = ~new_n6055_ & new_n6112_1_;
  assign new_n6114_ = ~new_n6092_1_ & ~new_n6105_;
  assign new_n6115_ = ~new_n6113_ & new_n6114_;
  assign new_n6116_ = new_n6089_ & ~new_n6097_1_;
  assign new_n6117_1_ = ~new_n6102_1_ & new_n6116_;
  assign new_n6118_ = new_n6055_ & new_n6117_1_;
  assign new_n6119_ = ~new_n6084_ & ~new_n6102_1_;
  assign new_n6120_ = ~new_n6089_ & new_n6119_;
  assign new_n6121_ = ~new_n6060_ & new_n6120_;
  assign new_n6122_1_ = ~new_n6065_ & new_n6084_;
  assign new_n6123_ = new_n6102_1_ & new_n6122_1_;
  assign new_n6124_ = ~new_n6055_ & new_n6123_;
  assign new_n6125_ = new_n6115_ & ~new_n6118_;
  assign new_n6126_ = ~new_n6121_ & ~new_n6124_;
  assign new_n6127_1_ = new_n6125_ & new_n6126_;
  assign new_n6128_ = new_n6055_ & new_n6066_;
  assign new_n6129_ = new_n6084_ & new_n6128_;
  assign new_n6130_ = ~new_n6102_1_ & new_n6129_;
  assign new_n6131_ = new_n6065_ & new_n6097_1_;
  assign new_n6132_1_ = new_n6055_ & new_n6131_;
  assign new_n6133_ = ~new_n6089_ & new_n6132_1_;
  assign new_n6134_ = ~new_n6110_ & new_n6133_;
  assign new_n6135_ = ~new_n6102_1_ & new_n6134_;
  assign new_n6136_ = ~new_n6097_1_ & new_n6102_1_;
  assign new_n6137_1_ = ~new_n6055_ & new_n6136_;
  assign new_n6138_ = ~new_n6110_ & new_n6137_1_;
  assign new_n6139_ = ~new_n6089_ & new_n6138_;
  assign new_n6140_ = ~new_n6055_ & new_n6066_;
  assign new_n6141_ = ~new_n6089_ & new_n6140_;
  assign new_n6142_1_ = ~new_n6084_ & new_n6141_;
  assign new_n6143_ = new_n6102_1_ & new_n6142_1_;
  assign new_n6144_ = ~new_n6130_ & ~new_n6135_;
  assign new_n6145_ = ~new_n6139_ & ~new_n6143_;
  assign new_n6146_ = new_n6144_ & new_n6145_;
  assign new_n6147_1_ = new_n6127_1_ & new_n6146_;
  assign new_n6148_ = ng1312 & ng1253;
  assign new_n6149_ = ng1315 & ng1176;
  assign new_n6150_ = ng1251 & ng1309;
  assign new_n6151_ = ~new_n6148_ & ~new_n6149_;
  assign n2276 = ~new_n6150_ & new_n6151_;
  assign new_n6153_ = ng185 & ~n2276;
  assign new_n6154_ = ng1228 & new_n6153_;
  assign new_n6155_ = ng1312 & ng1285;
  assign new_n6156_ = ng1315 & ng1288;
  assign new_n6157_1_ = ng1282 & ng1309;
  assign new_n6158_ = ~new_n6155_ & ~new_n6156_;
  assign new_n6159_ = ~new_n6157_1_ & new_n6158_;
  assign new_n6160_ = ~new_n6154_ & new_n6159_;
  assign new_n6161_ = ng1312 & ng1257;
  assign new_n6162_1_ = ng1315 & ng1259;
  assign new_n6163_ = ng1255 & ng1309;
  assign new_n6164_ = ~new_n6161_ & ~new_n6162_1_;
  assign n4577 = ~new_n6163_ & new_n6164_;
  assign new_n6166_ = ng1210 & ~n4577;
  assign new_n6167_1_ = ng185 & new_n6166_;
  assign new_n6168_ = ng1312 & ng1276;
  assign new_n6169_ = ng1315 & ng1279;
  assign new_n6170_ = ng1273 & ng1309;
  assign new_n6171_ = ~new_n6168_ & ~new_n6169_;
  assign new_n6172_1_ = ~new_n6170_ & new_n6171_;
  assign new_n6173_ = ~new_n6167_1_ & new_n6172_1_;
  assign new_n6174_ = new_n6147_1_ & ~new_n6160_;
  assign new_n6175_ = new_n6173_ & new_n6174_;
  assign new_n6176_ = ~new_n6097_1_ & ~new_n6102_1_;
  assign new_n6177_1_ = new_n6055_ & new_n6176_;
  assign new_n6178_ = ~new_n6084_ & new_n6177_1_;
  assign new_n6179_ = ~new_n6089_ & new_n6178_;
  assign new_n6180_ = new_n6097_1_ & ~new_n6102_1_;
  assign new_n6181_ = ~new_n6065_ & new_n6180_;
  assign new_n6182_1_ = ~new_n6110_ & new_n6181_;
  assign new_n6183_ = ~new_n6089_ & new_n6182_1_;
  assign new_n6184_ = new_n6065_ & new_n6089_;
  assign new_n6185_1_ = new_n6102_1_ & new_n6184_;
  assign new_n6186_ = ~new_n6055_ & new_n6185_1_;
  assign new_n6187_ = new_n6065_ & new_n6102_1_;
  assign new_n6188_ = new_n6055_ & new_n6187_;
  assign new_n6189_1_ = ~new_n6084_ & new_n6188_;
  assign new_n6190_ = ~new_n6089_ & new_n6189_1_;
  assign new_n6191_ = ~new_n6183_ & ~new_n6186_;
  assign new_n6192_ = ~new_n6190_ & new_n6191_;
  assign new_n6193_1_ = new_n6060_ & ~new_n6102_1_;
  assign new_n6194_ = ~new_n6055_ & new_n6193_1_;
  assign new_n6195_ = ~new_n6084_ & new_n6194_;
  assign new_n6196_ = new_n6089_ & new_n6195_;
  assign new_n6197_ = ~new_n6179_ & new_n6192_;
  assign new_n6198_1_ = ~new_n6196_ & new_n6197_;
  assign new_n6199_ = ~new_n6060_ & ~new_n6110_;
  assign new_n6200_ = new_n6102_1_ & new_n6199_;
  assign new_n6201_1_ = ~new_n6055_ & new_n6200_;
  assign new_n6202_ = new_n6084_ & ~new_n6102_1_;
  assign new_n6203_ = ~new_n6089_ & new_n6202_;
  assign new_n6204_ = ~new_n6065_ & new_n6203_;
  assign new_n6205_ = ~new_n6055_ & new_n6117_1_;
  assign new_n6206_1_ = new_n6097_1_ & new_n6102_1_;
  assign new_n6207_ = new_n6065_ & new_n6206_1_;
  assign new_n6208_ = new_n6084_ & new_n6207_;
  assign new_n6209_ = ~new_n6089_ & new_n6208_;
  assign new_n6210_ = ~new_n6204_ & ~new_n6205_;
  assign new_n6211_1_ = ~new_n6209_ & new_n6210_;
  assign new_n6212_ = new_n6060_ & new_n6110_;
  assign new_n6213_ = ~new_n6102_1_ & new_n6212_;
  assign new_n6214_1_ = new_n6055_ & new_n6213_;
  assign new_n6215_ = ~new_n6201_1_ & new_n6211_1_;
  assign new_n6216_ = ~new_n6214_1_ & new_n6215_;
  assign new_n6217_ = new_n6084_ & new_n6102_1_;
  assign new_n6218_ = ~new_n6060_ & new_n6217_;
  assign new_n6219_1_ = new_n6084_ & new_n6097_1_;
  assign new_n6220_ = ~new_n6102_1_ & new_n6219_1_;
  assign new_n6221_ = ~new_n6065_ & new_n6220_;
  assign new_n6222_ = ~new_n6097_1_ & new_n6110_;
  assign new_n6223_ = new_n6055_ & new_n6222_;
  assign new_n6224_1_ = ~new_n6084_ & ~new_n6097_1_;
  assign new_n6225_ = new_n6089_ & new_n6224_1_;
  assign new_n6226_ = ~new_n6055_ & new_n6225_;
  assign new_n6227_ = ~new_n6218_ & ~new_n6221_;
  assign new_n6228_ = ~new_n6223_ & ~new_n6226_;
  assign new_n6229_1_ = new_n6227_ & new_n6228_;
  assign new_n6230_ = new_n6198_1_ & new_n6216_;
  assign new_n6231_ = new_n6229_1_ & new_n6230_;
  assign new_n6232_ = new_n6160_ & ~new_n6231_;
  assign new_n6233_ = new_n6147_1_ & new_n6232_;
  assign new_n6234_1_ = ~new_n6175_ & ~new_n6233_;
  assign new_n6235_ = new_n5366_ & new_n6234_1_;
  assign new_n6236_ = ~new_n5366_ & new_n6044_;
  assign new_n6237_ = ~new_n6235_ & ~new_n6236_;
  assign new_n6238_ = ng1312 & ~new_n6237_;
  assign new_n6239_1_ = ~ng1303 & ~ng1312;
  assign n507 = ~new_n6238_ & ~new_n6239_1_;
  assign new_n6241_ = ng1312 & ng1316;
  assign new_n6242_ = ng1315 & ~ng1345;
  assign new_n6243_ = ng1326 & new_n6242_;
  assign new_n6244_1_ = ng1319 & new_n6243_;
  assign new_n6245_ = ng1339 & new_n6244_1_;
  assign new_n6246_ = ng1332 & new_n6245_;
  assign new_n6247_ = ng1346 & new_n6246_;
  assign new_n6248_ = ng1358 & new_n6247_;
  assign new_n6249_1_ = ng1352 & ~new_n6248_;
  assign new_n6250_ = ~ng1352 & new_n6248_;
  assign new_n6251_ = ~new_n6249_1_ & ~new_n6250_;
  assign n517 = ~new_n6241_ & ~new_n6251_;
  assign new_n6253_ = ng1211 & ng1224;
  assign new_n6254_1_ = ~ng1345 & new_n6253_;
  assign new_n6255_ = ng1312 & new_n6254_1_;
  assign new_n6256_ = ~ng1392 & ~new_n6255_;
  assign new_n6257_ = ng1339 & new_n6255_;
  assign n522 = ~new_n6256_ & ~new_n6257_;
  assign new_n6259_1_ = ng1309 & new_n6254_1_;
  assign new_n6260_ = ~ng1403 & ~new_n6259_1_;
  assign new_n6261_ = ng1352 & new_n6259_1_;
  assign n527 = ~new_n6260_ & ~new_n6261_;
  assign new_n6263_ = ng1315 & new_n6254_1_;
  assign new_n6264_1_ = ~ng1411 & ~new_n6263_;
  assign new_n6265_ = ng1378 & new_n6263_;
  assign n532 = ~new_n6264_1_ & ~new_n6265_;
  assign new_n6267_ = ~ng1316 & ~new_n6254_1_;
  assign new_n6268_ = ng1312 & ~new_n6267_;
  assign new_n6269_1_ = ~ng1425 & ~new_n6268_;
  assign new_n6270_ = ng1316 & new_n6268_;
  assign n537 = ~new_n6269_1_ & ~new_n6270_;
  assign new_n6272_ = ~ng1527 & ~new_n5517_1_;
  assign new_n6273_ = ng1486 & new_n5517_1_;
  assign n542 = ~new_n6272_ & ~new_n6273_;
  assign new_n6275_ = ~ng1535 & ~new_n4773_;
  assign new_n6276_ = ng1501 & new_n4773_;
  assign n547 = ~new_n6275_ & ~new_n6276_;
  assign new_n6278_ = ng823 & n1621;
  assign new_n6279_1_ = ~ng1552 & ~new_n6278_;
  assign new_n6280_ = ~ng1496 & ~ng1501;
  assign new_n6281_ = ng1506 & new_n6280_;
  assign new_n6282_ = ng1491 & new_n6281_;
  assign new_n6283_ = new_n6278_ & ~new_n6282_;
  assign n552 = ~new_n6279_1_ & ~new_n6283_;
  assign new_n6285_ = ~ng1697 & ng823;
  assign new_n6286_ = ~ng1698 & ng853;
  assign new_n6287_ = ~ng1696 & ng826;
  assign new_n6288_ = ~new_n6285_ & ~new_n6286_;
  assign new_n6289_1_ = ~new_n6287_ & new_n6288_;
  assign new_n6290_ = ng823 & ~ng1694;
  assign new_n6291_ = ~ng1695 & ng853;
  assign new_n6292_ = ~ng1693 & ng826;
  assign new_n6293_ = ~new_n6290_ & ~new_n6291_;
  assign new_n6294_1_ = ~new_n6292_ & new_n6293_;
  assign new_n6295_ = ~ng1700 & ng823;
  assign new_n6296_ = ~ng1701 & ng853;
  assign new_n6297_ = ~ng1699 & ng826;
  assign new_n6298_ = ~new_n6295_ & ~new_n6296_;
  assign new_n6299_1_ = ~new_n6297_ & new_n6298_;
  assign new_n6300_ = ~new_n6289_1_ & new_n6294_1_;
  assign new_n6301_ = new_n6299_1_ & new_n6300_;
  assign new_n6302_ = new_n6289_1_ & new_n6294_1_;
  assign new_n6303_ = new_n6299_1_ & new_n6302_;
  assign new_n6304_1_ = ~new_n6301_ & ~new_n6303_;
  assign new_n6305_ = ng1579 & ng823;
  assign new_n6306_ = ng1582 & ng853;
  assign new_n6307_ = ng826 & ng1576;
  assign new_n6308_ = ~new_n6305_ & ~new_n6306_;
  assign new_n6309_1_ = ~new_n6307_ & new_n6308_;
  assign new_n6310_ = ng1624 & ng823;
  assign new_n6311_ = ng853 & ng1627;
  assign new_n6312_ = ng826 & ng1621;
  assign new_n6313_ = ~new_n6310_ & ~new_n6311_;
  assign new_n6314_1_ = ~new_n6312_ & new_n6313_;
  assign new_n6315_ = ng1615 & ng823;
  assign new_n6316_ = ng853 & ng1618;
  assign new_n6317_ = ng826 & ng1612;
  assign new_n6318_ = ~new_n6315_ & ~new_n6316_;
  assign new_n6319_1_ = ~new_n6317_ & new_n6318_;
  assign new_n6320_ = ~new_n6309_1_ & ~new_n6314_1_;
  assign new_n6321_ = ~new_n6319_1_ & new_n6320_;
  assign new_n6322_ = ng1651 & ng823;
  assign new_n6323_1_ = ng1654 & ng853;
  assign new_n6324_ = ng826 & ng1648;
  assign new_n6325_ = ~new_n6322_ & ~new_n6323_1_;
  assign new_n6326_ = ~new_n6324_ & new_n6325_;
  assign new_n6327_ = ng1642 & ng823;
  assign new_n6328_1_ = ng853 & ng1645;
  assign new_n6329_ = ng826 & ng1639;
  assign new_n6330_ = ~new_n6327_ & ~new_n6328_1_;
  assign new_n6331_1_ = ~new_n6329_ & new_n6330_;
  assign new_n6332_ = ng823 & ng1588;
  assign new_n6333_ = ng853 & ng1591;
  assign new_n6334_ = ng1585 & ng826;
  assign new_n6335_ = ~new_n6332_ & ~new_n6333_;
  assign new_n6336_1_ = ~new_n6334_ & new_n6335_;
  assign new_n6337_ = ng823 & ng1633;
  assign new_n6338_ = ng1636 & ng853;
  assign new_n6339_1_ = ng826 & ng1630;
  assign new_n6340_ = ~new_n6337_ & ~new_n6338_;
  assign new_n6341_ = ~new_n6339_1_ & new_n6340_;
  assign new_n6342_ = ng823 & ng1570;
  assign new_n6343_ = ng1573 & ng853;
  assign new_n6344_1_ = ng826 & ng1567;
  assign new_n6345_ = ~new_n6342_ & ~new_n6343_;
  assign new_n6346_ = ~new_n6344_1_ & new_n6345_;
  assign new_n6347_ = new_n6336_1_ & new_n6341_;
  assign new_n6348_1_ = new_n6346_ & new_n6347_;
  assign new_n6349_ = ng1597 & ng823;
  assign new_n6350_ = ng1600 & ng853;
  assign new_n6351_ = ng826 & ng1594;
  assign new_n6352_ = ~new_n6349_ & ~new_n6350_;
  assign new_n6353_1_ = ~new_n6351_ & new_n6352_;
  assign new_n6354_ = new_n6331_1_ & new_n6348_1_;
  assign new_n6355_ = new_n6353_1_ & new_n6354_;
  assign new_n6356_ = ng823 & ng1606;
  assign new_n6357_ = ng853 & ng1609;
  assign new_n6358_1_ = ng826 & ng1603;
  assign new_n6359_ = ~new_n6356_ & ~new_n6357_;
  assign new_n6360_ = ~new_n6358_1_ & new_n6359_;
  assign new_n6361_ = new_n6321_ & ~new_n6326_;
  assign new_n6362_ = new_n6355_ & new_n6361_;
  assign new_n6363_1_ = ~new_n6360_ & new_n6362_;
  assign new_n6364_ = new_n6301_ & new_n6363_1_;
  assign new_n6365_ = new_n6309_1_ & new_n6314_1_;
  assign new_n6366_ = new_n6319_1_ & new_n6365_;
  assign new_n6367_ = new_n6326_ & new_n6366_;
  assign new_n6368_1_ = new_n6355_ & new_n6367_;
  assign new_n6369_ = new_n6360_ & new_n6368_1_;
  assign new_n6370_ = ~new_n6301_ & new_n6369_;
  assign new_n6371_ = ~new_n6364_ & ~new_n6370_;
  assign new_n6372_ = ~new_n6304_1_ & ~new_n6371_;
  assign new_n6373_1_ = ~ng1552 & ng823;
  assign new_n6374_ = ~ng1550 & ng853;
  assign new_n6375_ = ~ng1551 & ng826;
  assign new_n6376_ = ~new_n6373_1_ & ~new_n6374_;
  assign new_n6377_ = ~new_n6375_ & new_n6376_;
  assign new_n6378_1_ = ng1476 & ~new_n6319_1_;
  assign new_n6379_ = ng1476 & ~new_n6378_1_;
  assign new_n6380_ = ~new_n6319_1_ & ~new_n6378_1_;
  assign new_n6381_ = ~new_n6379_ & ~new_n6380_;
  assign new_n6382_ = ng1506 & ~new_n6331_1_;
  assign new_n6383_1_ = ng1506 & ~new_n6382_;
  assign new_n6384_ = ~new_n6331_1_ & ~new_n6382_;
  assign new_n6385_ = ~new_n6383_1_ & ~new_n6384_;
  assign new_n6386_ = new_n6381_ & new_n6385_;
  assign new_n6387_ = ng1486 & ~new_n6314_1_;
  assign new_n6388_1_ = ng1486 & ~new_n6387_;
  assign new_n6389_ = ~new_n6314_1_ & ~new_n6387_;
  assign new_n6390_ = ~new_n6388_1_ & ~new_n6389_;
  assign new_n6391_ = ~ng1555 & ng823;
  assign new_n6392_ = ng853 & ~ng1553;
  assign new_n6393_1_ = ~ng1554 & ng826;
  assign new_n6394_ = ~new_n6391_ & ~new_n6392_;
  assign new_n6395_ = ~new_n6393_1_ & new_n6394_;
  assign new_n6396_ = ~new_n6326_ & ~new_n6395_;
  assign new_n6397_ = ~new_n6395_ & ~new_n6396_;
  assign new_n6398_1_ = ~new_n6326_ & ~new_n6396_;
  assign new_n6399_ = ~new_n6397_ & ~new_n6398_1_;
  assign new_n6400_ = new_n6390_ & new_n6399_;
  assign new_n6401_ = ng1496 & ~new_n6341_;
  assign new_n6402_ = ng1496 & ~new_n6401_;
  assign new_n6403_1_ = ~new_n6341_ & ~new_n6401_;
  assign new_n6404_ = ~new_n6402_ & ~new_n6403_1_;
  assign new_n6405_ = ~new_n6386_ & ~new_n6400_;
  assign new_n6406_ = ~new_n6404_ & new_n6405_;
  assign new_n6407_ = new_n6385_ & new_n6404_;
  assign new_n6408_1_ = new_n6381_ & new_n6390_;
  assign new_n6409_ = ~new_n6407_ & ~new_n6408_1_;
  assign new_n6410_ = ~new_n6399_ & new_n6409_;
  assign new_n6411_ = new_n6385_ & new_n6399_;
  assign new_n6412_1_ = new_n6390_ & new_n6404_;
  assign new_n6413_ = ~new_n6411_ & ~new_n6412_1_;
  assign new_n6414_ = ~new_n6381_ & new_n6413_;
  assign new_n6415_ = ~new_n6406_ & ~new_n6410_;
  assign new_n6416_1_ = ~new_n6414_ & new_n6415_;
  assign new_n6417_ = ng2257 & ~new_n6377_;
  assign new_n6418_ = ~new_n6416_1_ & new_n6417_;
  assign new_n6419_ = ng1471 & ~new_n6346_;
  assign new_n6420_ = ng1471 & ~new_n6419_;
  assign new_n6421_1_ = ~new_n6346_ & ~new_n6419_;
  assign new_n6422_ = ~new_n6420_ & ~new_n6421_1_;
  assign new_n6423_ = ng1501 & ~new_n6353_1_;
  assign new_n6424_ = ng1501 & ~new_n6423_;
  assign new_n6425_1_ = ~new_n6353_1_ & ~new_n6423_;
  assign new_n6426_ = ~new_n6424_ & ~new_n6425_1_;
  assign new_n6427_ = new_n6422_ & new_n6426_;
  assign new_n6428_ = ng1481 & ~new_n6309_1_;
  assign new_n6429_ = ng1481 & ~new_n6428_;
  assign new_n6430_1_ = ~new_n6309_1_ & ~new_n6428_;
  assign new_n6431_ = ~new_n6429_ & ~new_n6430_1_;
  assign new_n6432_ = ng823 & ~ng1558;
  assign new_n6433_ = ng853 & ~ng1556;
  assign new_n6434_ = ng826 & ~ng1557;
  assign new_n6435_1_ = ~new_n6432_ & ~new_n6433_;
  assign new_n6436_ = ~new_n6434_ & new_n6435_1_;
  assign new_n6437_ = ~new_n6360_ & ~new_n6436_;
  assign new_n6438_ = ~new_n6436_ & ~new_n6437_;
  assign new_n6439_1_ = ~new_n6360_ & ~new_n6437_;
  assign new_n6440_ = ~new_n6438_ & ~new_n6439_1_;
  assign new_n6441_ = new_n6431_ & new_n6440_;
  assign new_n6442_ = ng1491 & ~new_n6336_1_;
  assign new_n6443_ = ng1491 & ~new_n6442_;
  assign new_n6444_1_ = ~new_n6336_1_ & ~new_n6442_;
  assign new_n6445_ = ~new_n6443_ & ~new_n6444_1_;
  assign new_n6446_ = ~new_n6427_ & ~new_n6441_;
  assign new_n6447_1_ = ~new_n6445_ & new_n6446_;
  assign new_n6448_ = new_n6426_ & new_n6445_;
  assign new_n6449_ = new_n6422_ & new_n6431_;
  assign new_n6450_ = ~new_n6448_ & ~new_n6449_;
  assign new_n6451_ = ~new_n6440_ & new_n6450_;
  assign new_n6452_1_ = new_n6426_ & new_n6440_;
  assign new_n6453_ = new_n6431_ & new_n6445_;
  assign new_n6454_ = ~new_n6452_1_ & ~new_n6453_;
  assign new_n6455_ = ~new_n6422_ & new_n6454_;
  assign new_n6456_ = ~new_n6447_1_ & ~new_n6451_;
  assign new_n6457_1_ = ~new_n6455_ & new_n6456_;
  assign new_n6458_ = new_n6417_ & ~new_n6457_1_;
  assign new_n6459_ = ~new_n6418_ & ~new_n6458_;
  assign new_n6460_1_ = ~ng1546 & ng823;
  assign new_n6461_ = ~ng1544 & ng853;
  assign new_n6462_ = ~ng1545 & ng826;
  assign new_n6463_ = ~new_n6460_1_ & ~new_n6461_;
  assign new_n6464_ = ~new_n6462_ & new_n6463_;
  assign new_n6465_1_ = ~new_n6395_ & ~new_n6464_;
  assign new_n6466_ = ~new_n6464_ & ~new_n6465_1_;
  assign new_n6467_ = ~new_n6395_ & ~new_n6465_1_;
  assign new_n6468_ = ~new_n6466_ & ~new_n6467_;
  assign new_n6469_ = ~ng1537 & ng823;
  assign new_n6470_1_ = ~ng1535 & ng853;
  assign new_n6471_ = ~ng1536 & ng826;
  assign new_n6472_ = ~new_n6469_ & ~new_n6470_1_;
  assign new_n6473_ = ~new_n6471_ & new_n6472_;
  assign new_n6474_ = ng1501 & ~new_n6473_;
  assign new_n6475_1_ = ~new_n6473_ & ~new_n6474_;
  assign new_n6476_ = ng1501 & ~new_n6474_;
  assign new_n6477_ = ~new_n6475_1_ & ~new_n6476_;
  assign new_n6478_ = ~ng1540 & ng823;
  assign new_n6479_ = ~ng1538 & ng853;
  assign new_n6480_1_ = ~ng1539 & ng826;
  assign new_n6481_ = ~new_n6478_ & ~new_n6479_;
  assign new_n6482_ = ~new_n6480_1_ & new_n6481_;
  assign new_n6483_ = ng1506 & ~new_n6482_;
  assign new_n6484_ = ~new_n6482_ & ~new_n6483_;
  assign new_n6485_1_ = ng1506 & ~new_n6483_;
  assign new_n6486_ = ~new_n6484_ & ~new_n6485_1_;
  assign new_n6487_ = ~ng1534 & ng823;
  assign new_n6488_ = ~ng1532 & ng853;
  assign new_n6489_ = ng826 & ~ng1533;
  assign new_n6490_1_ = ~new_n6487_ & ~new_n6488_;
  assign new_n6491_ = ~new_n6489_ & new_n6490_1_;
  assign new_n6492_ = ng1496 & ~new_n6491_;
  assign new_n6493_ = ~new_n6491_ & ~new_n6492_;
  assign new_n6494_ = ng1496 & ~new_n6492_;
  assign new_n6495_1_ = ~new_n6493_ & ~new_n6494_;
  assign new_n6496_ = new_n6477_ & new_n6486_;
  assign new_n6497_ = new_n6495_1_ & new_n6496_;
  assign new_n6498_ = ~ng1543 & ng823;
  assign new_n6499_ = ~ng1541 & ng853;
  assign new_n6500_1_ = ng826 & ~ng1542;
  assign new_n6501_ = ~new_n6498_ & ~new_n6499_;
  assign new_n6502_ = ~new_n6500_1_ & new_n6501_;
  assign new_n6503_ = ~new_n6436_ & ~new_n6502_;
  assign new_n6504_ = ~new_n6502_ & ~new_n6503_;
  assign new_n6505_1_ = ~new_n6436_ & ~new_n6503_;
  assign new_n6506_ = ~new_n6504_ & ~new_n6505_1_;
  assign new_n6507_ = new_n6468_ & new_n6497_;
  assign new_n6508_ = new_n6506_ & new_n6507_;
  assign new_n6509_ = ~ng1531 & ng823;
  assign new_n6510_1_ = ~ng1529 & ng853;
  assign new_n6511_ = ~ng1530 & ng826;
  assign new_n6512_ = ~new_n6509_ & ~new_n6510_1_;
  assign new_n6513_ = ~new_n6511_ & new_n6512_;
  assign new_n6514_ = ng1491 & ~new_n6513_;
  assign new_n6515_1_ = ~new_n6513_ & ~new_n6514_;
  assign new_n6516_ = ng1491 & ~new_n6514_;
  assign new_n6517_ = ~new_n6515_1_ & ~new_n6516_;
  assign new_n6518_ = ng823 & ~ng1516;
  assign new_n6519_ = ng853 & ~ng1514;
  assign new_n6520_1_ = ~ng1515 & ng826;
  assign new_n6521_ = ~new_n6518_ & ~new_n6519_;
  assign new_n6522_ = ~new_n6520_1_ & new_n6521_;
  assign new_n6523_ = ng1476 & ~new_n6522_;
  assign new_n6524_ = ~new_n6522_ & ~new_n6523_;
  assign new_n6525_1_ = ng1476 & ~new_n6523_;
  assign new_n6526_ = ~new_n6524_ & ~new_n6525_1_;
  assign new_n6527_ = ~ng1525 & ng823;
  assign new_n6528_ = ~ng1523 & ng853;
  assign new_n6529_ = ~ng1524 & ng826;
  assign new_n6530_1_ = ~new_n6527_ & ~new_n6528_;
  assign new_n6531_ = ~new_n6529_ & new_n6530_1_;
  assign new_n6532_ = ng1481 & ~new_n6531_;
  assign new_n6533_ = ~new_n6531_ & ~new_n6532_;
  assign new_n6534_ = ng1481 & ~new_n6532_;
  assign new_n6535_1_ = ~new_n6533_ & ~new_n6534_;
  assign new_n6536_ = ~ng1513 & ng823;
  assign new_n6537_ = ~ng1511 & ng853;
  assign new_n6538_ = ~ng1512 & ng826;
  assign new_n6539_ = ~new_n6536_ & ~new_n6537_;
  assign new_n6540_1_ = ~new_n6538_ & new_n6539_;
  assign new_n6541_ = ng1471 & ~new_n6540_1_;
  assign new_n6542_ = ~new_n6540_1_ & ~new_n6541_;
  assign new_n6543_ = ng1471 & ~new_n6541_;
  assign new_n6544_ = ~new_n6542_ & ~new_n6543_;
  assign new_n6545_1_ = new_n6526_ & new_n6535_1_;
  assign new_n6546_ = new_n6544_ & new_n6545_1_;
  assign new_n6547_ = ~ng1528 & ng823;
  assign new_n6548_ = ~ng1526 & ng853;
  assign new_n6549_ = ~ng1527 & ng826;
  assign new_n6550_1_ = ~new_n6547_ & ~new_n6548_;
  assign new_n6551_ = ~new_n6549_ & new_n6550_1_;
  assign new_n6552_ = ng1486 & ~new_n6551_;
  assign new_n6553_ = ~new_n6551_ & ~new_n6552_;
  assign new_n6554_ = ng1486 & ~new_n6552_;
  assign new_n6555_1_ = ~new_n6553_ & ~new_n6554_;
  assign new_n6556_ = new_n6517_ & new_n6546_;
  assign new_n6557_ = new_n6555_1_ & new_n6556_;
  assign new_n6558_ = new_n6508_ & new_n6557_;
  assign new_n6559_ = ~new_n6377_ & new_n6459_;
  assign new_n6560_1_ = ng2257 & new_n6558_;
  assign new_n6561_ = new_n6559_ & new_n6560_1_;
  assign new_n6562_ = ~ng1704 & ng823;
  assign new_n6563_ = ng853 & ~ng1702;
  assign new_n6564_ = ~ng1703 & ng826;
  assign new_n6565_1_ = ~new_n6562_ & ~new_n6563_;
  assign new_n6566_ = ~new_n6564_ & new_n6565_1_;
  assign new_n6567_ = new_n6289_1_ & ~new_n6294_1_;
  assign new_n6568_ = new_n6299_1_ & new_n6567_;
  assign new_n6569_ = new_n6561_ & ~new_n6566_;
  assign new_n6570_1_ = new_n6568_ & new_n6569_;
  assign new_n6571_ = new_n6417_ & new_n6558_;
  assign new_n6572_ = ~new_n6299_1_ & new_n6567_;
  assign new_n6573_ = ~new_n6566_ & new_n6571_;
  assign new_n6574_ = new_n6572_ & new_n6573_;
  assign new_n6575_1_ = ng2257 & new_n6377_;
  assign new_n6576_ = ~new_n6294_1_ & new_n6575_1_;
  assign new_n6577_ = ~new_n6570_1_ & ~new_n6574_;
  assign new_n6578_ = ~new_n6576_ & new_n6577_;
  assign new_n6579_ = ~ng1785 & ng823;
  assign new_n6580_1_ = ~ng1783 & ng853;
  assign new_n6581_ = ng826 & ~ng1784;
  assign new_n6582_ = ~new_n6579_ & ~new_n6580_1_;
  assign new_n6583_ = ~new_n6581_ & new_n6582_;
  assign new_n6584_ = new_n6571_ & ~new_n6583_;
  assign new_n6585_1_ = new_n6578_ & ~new_n6584_;
  assign new_n6586_ = ~new_n6372_ & new_n6585_1_;
  assign new_n6587_ = new_n6372_ & new_n6585_1_;
  assign new_n6588_ = ng1506 & ~new_n6587_;
  assign new_n6589_ = ~new_n6586_ & ~new_n6588_;
  assign new_n6590_1_ = new_n6301_ & ~new_n6353_1_;
  assign new_n6591_ = ~new_n6301_ & new_n6353_1_;
  assign new_n6592_ = ~new_n6590_1_ & ~new_n6591_;
  assign new_n6593_ = new_n6301_ & ~new_n6319_1_;
  assign new_n6594_ = ~new_n6301_ & new_n6319_1_;
  assign new_n6595_1_ = ~new_n6593_ & ~new_n6594_;
  assign new_n6596_ = new_n6301_ & new_n6346_;
  assign new_n6597_ = ~new_n6301_ & ~new_n6346_;
  assign new_n6598_ = ~new_n6596_ & ~new_n6597_;
  assign new_n6599_ = ~new_n6304_1_ & new_n6598_;
  assign new_n6600_1_ = ~new_n6595_1_ & new_n6599_;
  assign new_n6601_ = new_n6301_ & ~new_n6314_1_;
  assign new_n6602_ = ~new_n6301_ & new_n6314_1_;
  assign new_n6603_ = ~new_n6601_ & ~new_n6602_;
  assign new_n6604_ = new_n6301_ & ~new_n6309_1_;
  assign new_n6605_1_ = ~new_n6301_ & new_n6309_1_;
  assign new_n6606_ = ~new_n6604_ & ~new_n6605_1_;
  assign new_n6607_ = ~new_n6603_ & ~new_n6606_;
  assign new_n6608_ = new_n6301_ & ~new_n6341_;
  assign new_n6609_ = ~new_n6301_ & new_n6341_;
  assign new_n6610_1_ = ~new_n6608_ & ~new_n6609_;
  assign new_n6611_ = new_n6301_ & ~new_n6336_1_;
  assign new_n6612_ = ~new_n6301_ & new_n6336_1_;
  assign new_n6613_ = ~new_n6611_ & ~new_n6612_;
  assign new_n6614_1_ = ~new_n6610_1_ & ~new_n6613_;
  assign new_n6615_ = new_n6600_1_ & new_n6607_;
  assign new_n6616_ = new_n6614_1_ & new_n6615_;
  assign new_n6617_ = ~new_n6592_ & new_n6616_;
  assign new_n6618_ = new_n6331_1_ & new_n6617_;
  assign new_n6619_1_ = ~new_n6331_1_ & ~new_n6617_;
  assign new_n6620_ = ~new_n6618_ & ~new_n6619_1_;
  assign new_n6621_ = new_n6586_ & new_n6620_;
  assign new_n6622_ = ~new_n6589_ & ~new_n6621_;
  assign new_n6623_ = ng823 & ~new_n6622_;
  assign new_n6624_1_ = ~ng1642 & ~ng823;
  assign n557 = ~new_n6623_ & ~new_n6624_1_;
  assign new_n6626_ = ng1466 & new_n5128_;
  assign new_n6627_ = ng1462 & new_n6626_;
  assign new_n6628_ = ng1457 & new_n6627_;
  assign new_n6629_1_ = ng1453 & ~new_n6628_;
  assign new_n6630_ = ~ng1453 & new_n6628_;
  assign new_n6631_ = ~new_n6629_1_ & ~new_n6630_;
  assign n562 = ~new_n5127_1_ & ~new_n6631_;
  assign new_n6633_1_ = new_n5125_ & ~new_n6303_;
  assign new_n6634_ = ~new_n6299_1_ & new_n6300_;
  assign new_n6635_ = ~new_n6633_1_ & ~new_n6634_;
  assign new_n6636_ = ng823 & new_n6635_;
  assign new_n6637_ = ~ng1739 & ~new_n6636_;
  assign new_n6638_1_ = ~ng1754 & ng823;
  assign new_n6639_ = ~ng1757 & ng853;
  assign new_n6640_ = ~ng1765 & ng826;
  assign new_n6641_ = ~new_n6638_1_ & ~new_n6639_;
  assign new_n6642_ = ~new_n6640_ & new_n6641_;
  assign new_n6643_1_ = ng823 & ~ng1724;
  assign new_n6644_ = ng853 & ~ng1727;
  assign new_n6645_ = ~ng1735 & ng826;
  assign new_n6646_ = ~new_n6643_1_ & ~new_n6644_;
  assign new_n6647_ = ~new_n6645_ & new_n6646_;
  assign new_n6648_1_ = ~new_n6642_ & new_n6647_;
  assign new_n6649_ = ~pg3229 & new_n6648_1_;
  assign new_n6650_ = ~new_n6642_ & ~new_n6647_;
  assign new_n6651_ = pg3229 & new_n6650_;
  assign new_n6652_ = ~ng1739 & ng823;
  assign new_n6653_1_ = ~ng1742 & ng853;
  assign new_n6654_ = ~ng1750 & ng826;
  assign new_n6655_ = ~new_n6652_ & ~new_n6653_1_;
  assign new_n6656_ = ~new_n6654_ & new_n6655_;
  assign new_n6657_1_ = new_n6642_ & ~new_n6656_;
  assign new_n6658_ = ~new_n6649_ & ~new_n6651_;
  assign new_n6659_ = ~new_n6657_1_ & new_n6658_;
  assign new_n6660_ = new_n6636_ & ~new_n6659_;
  assign n567 = ~new_n6637_ & ~new_n6660_;
  assign new_n6662_1_ = ng1801 & ng823;
  assign new_n6663_ = ng1804 & ng853;
  assign new_n6664_ = ng1798 & ng826;
  assign new_n6665_ = ~new_n6662_1_ & ~new_n6663_;
  assign n5082 = new_n6664_ | ~new_n6665_;
  assign new_n6667_ = ng1792 & ng823;
  assign new_n6668_ = ng1795 & ng853;
  assign new_n6669_ = ng826 & ng1789;
  assign new_n6670_ = ~new_n6667_ & ~new_n6668_;
  assign new_n6671_1_ = ~new_n6669_ & new_n6670_;
  assign new_n6672_ = ng1496 & ng1506;
  assign new_n6673_ = ng1501 & new_n6672_;
  assign new_n6674_ = ng1491 & new_n6673_;
  assign new_n6675_ = ng1486 & ng1476;
  assign new_n6676_1_ = ng1481 & new_n6675_;
  assign new_n6677_ = ng1471 & new_n6676_1_;
  assign new_n6678_ = new_n6674_ & new_n6677_;
  assign new_n6679_ = ~new_n6395_ & ~new_n6436_;
  assign new_n6680_ = new_n6678_ & new_n6679_;
  assign new_n6681_1_ = ~ng1809 & ng823;
  assign new_n6682_ = ~ng1807 & ng853;
  assign new_n6683_ = ~ng1808 & ng826;
  assign new_n6684_ = ~new_n6681_1_ & ~new_n6682_;
  assign new_n6685_ = ~new_n6683_ & new_n6684_;
  assign new_n6686_1_ = ~new_n6680_ & ~new_n6685_;
  assign new_n6687_ = n5082 & ~new_n6686_1_;
  assign new_n6688_ = ~new_n6575_1_ & new_n6685_;
  assign new_n6689_ = new_n6680_ & ~new_n6688_;
  assign new_n6690_ = ~n5082 & ~new_n6689_;
  assign new_n6691_1_ = ~new_n6687_ & ~new_n6690_;
  assign new_n6692_ = ~new_n6671_1_ & new_n6691_1_;
  assign new_n6693_ = new_n6575_1_ & new_n6680_;
  assign new_n6694_ = ~n5082 & ~new_n6693_;
  assign new_n6695_ = ~n5082 & ~new_n6694_;
  assign new_n6696_1_ = new_n6671_1_ & new_n6695_;
  assign new_n6697_ = ~new_n6692_ & ~new_n6696_1_;
  assign new_n6698_ = ng2384 & ~new_n6697_;
  assign new_n6699_ = n5082 & new_n6698_;
  assign new_n6700_ = n5082 & ~new_n6699_;
  assign new_n6701_1_ = new_n6698_ & ~new_n6699_;
  assign new_n6702_ = ~new_n6700_ & ~new_n6701_1_;
  assign new_n6703_ = ng826 & new_n6702_;
  assign new_n6704_ = ~ng1798 & ~ng826;
  assign n572 = ~new_n6703_ & ~new_n6704_;
  assign new_n6706_1_ = ng1822 & ng823;
  assign new_n6707_ = ng1825 & ng853;
  assign new_n6708_ = ng1819 & ng826;
  assign new_n6709_ = ~new_n6706_1_ & ~new_n6707_;
  assign new_n6710_ = ~new_n6708_ & new_n6709_;
  assign new_n6711_1_ = ~ng1830 & ng823;
  assign new_n6712_ = ~ng1828 & ng853;
  assign new_n6713_ = ~ng1829 & ng826;
  assign new_n6714_ = ~new_n6711_1_ & ~new_n6712_;
  assign new_n6715_1_ = ~new_n6713_ & new_n6714_;
  assign new_n6716_ = ng1813 & ng823;
  assign new_n6717_ = ng1816 & ng853;
  assign new_n6718_ = ng826 & ng1810;
  assign new_n6719_ = ~new_n6716_ & ~new_n6717_;
  assign new_n6720_1_ = ~new_n6718_ & new_n6719_;
  assign new_n6721_ = ~ng1561 & ng823;
  assign new_n6722_ = ~ng1559 & ng853;
  assign new_n6723_ = ~ng1560 & ng826;
  assign new_n6724_ = ~new_n6721_ & ~new_n6722_;
  assign new_n6725_1_ = ~new_n6723_ & new_n6724_;
  assign new_n6726_ = new_n6678_ & ~new_n6725_1_;
  assign new_n6727_ = new_n6710_ & ~new_n6720_1_;
  assign new_n6728_ = new_n6726_ & new_n6727_;
  assign new_n6729_ = ~new_n6710_ & new_n6720_1_;
  assign new_n6730_1_ = ~new_n6726_ & new_n6729_;
  assign new_n6731_ = ~new_n6728_ & ~new_n6730_1_;
  assign new_n6732_ = ng2384 & ~new_n6715_1_;
  assign new_n6733_ = ~new_n6731_ & new_n6732_;
  assign new_n6734_ = ~new_n6710_ & new_n6733_;
  assign new_n6735_1_ = ~new_n6710_ & ~new_n6734_;
  assign new_n6736_ = new_n6733_ & ~new_n6734_;
  assign new_n6737_ = ~new_n6735_1_ & ~new_n6736_;
  assign new_n6738_ = ng853 & new_n6737_;
  assign new_n6739_ = ~ng1825 & ~ng853;
  assign n577 = ~new_n6738_ & ~new_n6739_;
  assign new_n6741_ = new_n6294_1_ & new_n6299_1_;
  assign new_n6742_ = new_n6299_1_ & ~new_n6458_;
  assign new_n6743_ = ng2384 & ~new_n6418_;
  assign new_n6744_ = new_n6742_ & new_n6743_;
  assign new_n6745_1_ = new_n6289_1_ & ~new_n6744_;
  assign new_n6746_ = new_n6381_ & new_n6412_1_;
  assign new_n6747_ = new_n6399_ & new_n6746_;
  assign new_n6748_ = new_n6385_ & new_n6747_;
  assign new_n6749_ = new_n6422_ & new_n6453_;
  assign new_n6750_1_ = new_n6440_ & new_n6749_;
  assign new_n6751_ = new_n6426_ & new_n6750_1_;
  assign new_n6752_ = new_n6748_ & new_n6751_;
  assign new_n6753_ = ng2257 & new_n6752_;
  assign new_n6754_ = ~new_n6377_ & new_n6753_;
  assign new_n6755_1_ = ~new_n6575_1_ & ~new_n6754_;
  assign new_n6756_ = new_n6299_1_ & ~new_n6755_1_;
  assign new_n6757_ = ~new_n6377_ & ~new_n6752_;
  assign new_n6758_ = ng2257 & new_n6757_;
  assign new_n6759_ = ~new_n6458_ & ~new_n6758_;
  assign new_n6760_1_ = ~new_n6418_ & new_n6759_;
  assign new_n6761_ = ~new_n6299_1_ & ~new_n6760_1_;
  assign new_n6762_ = ~new_n6756_ & ~new_n6761_;
  assign new_n6763_ = ~new_n6289_1_ & new_n6762_;
  assign new_n6764_ = ~new_n6745_1_ & ~new_n6763_;
  assign new_n6765_1_ = ~new_n6294_1_ & new_n6764_;
  assign new_n6766_ = ~new_n6741_ & ~new_n6765_1_;
  assign new_n6767_ = ~new_n6299_1_ & new_n6766_;
  assign new_n6768_ = ~new_n6299_1_ & ~new_n6767_;
  assign new_n6769_ = new_n6766_ & ~new_n6767_;
  assign new_n6770_1_ = ~new_n6768_ & ~new_n6769_;
  assign new_n6771_ = ~new_n6584_ & ~new_n6770_1_;
  assign new_n6772_ = ng823 & ~new_n6771_;
  assign new_n6773_ = ~ng1700 & ~ng823;
  assign n582 = ~new_n6772_ & ~new_n6773_;
  assign new_n6775_1_ = ng1315 & ~ng1937;
  assign new_n6776_ = ~ng1890 & ~ng1315;
  assign n592 = ~new_n6775_1_ & ~new_n6776_;
  assign new_n6778_ = ng826 & ~new_n6572_;
  assign new_n6779_1_ = ~ng1858 & ~ng826;
  assign n602 = ~new_n6778_ & ~new_n6779_1_;
  assign new_n6781_ = ng1312 & ng1988;
  assign new_n6782_ = ng1991 & ng1315;
  assign new_n6783_1_ = ng1309 & ng1985;
  assign new_n6784_ = ~new_n6781_ & ~new_n6782_;
  assign new_n6785_ = ~new_n6783_1_ & new_n6784_;
  assign new_n6786_ = ng1874 & ng1312;
  assign new_n6787_ = ng1315 & ng1877;
  assign new_n6788_1_ = ng1871 & ng1309;
  assign new_n6789_ = ~new_n6786_ & ~new_n6787_;
  assign new_n6790_ = ~new_n6788_1_ & new_n6789_;
  assign new_n6791_ = ~new_n6785_ & ~new_n6790_;
  assign new_n6792_ = ng1312 & ng1997;
  assign new_n6793_1_ = ng1315 & ng2000;
  assign new_n6794_ = ng1309 & ng1994;
  assign new_n6795_ = ~new_n6792_ & ~new_n6793_1_;
  assign new_n6796_ = ~new_n6794_ & new_n6795_;
  assign new_n6797_ = ng1890 & new_n6790_;
  assign new_n6798_1_ = ~new_n6796_ & new_n6797_;
  assign new_n6799_ = new_n5297_1_ & ~new_n6798_1_;
  assign n2736 = ~new_n6791_ & ~new_n6799_;
  assign new_n6801_ = ng1309 & n2736;
  assign new_n6802_ = ~ng1959 & ~new_n6801_;
  assign new_n6803_1_ = ng1312 & ~ng1963;
  assign new_n6804_ = ng1315 & ~ng1961;
  assign new_n6805_ = ~ng1962 & ng1309;
  assign new_n6806_ = ~new_n6803_1_ & ~new_n6804_;
  assign new_n6807_ = ~new_n6805_ & new_n6806_;
  assign new_n6808_1_ = ng1312 & ~ng1957;
  assign new_n6809_ = ng1315 & ~ng1955;
  assign new_n6810_ = ~ng1956 & ng1309;
  assign new_n6811_ = ~new_n6808_1_ & ~new_n6809_;
  assign new_n6812_ = ~new_n6810_ & new_n6811_;
  assign new_n6813_1_ = ~new_n6807_ & new_n6812_;
  assign new_n6814_ = ~pg3229 & new_n6813_1_;
  assign new_n6815_ = ~new_n6807_ & ~new_n6812_;
  assign new_n6816_ = pg3229 & new_n6815_;
  assign new_n6817_ = ~ng1960 & ng1312;
  assign new_n6818_1_ = ng1315 & ~ng1958;
  assign new_n6819_ = ~ng1959 & ng1309;
  assign new_n6820_ = ~new_n6817_ & ~new_n6818_1_;
  assign new_n6821_ = ~new_n6819_ & new_n6820_;
  assign new_n6822_ = new_n6807_ & ~new_n6821_;
  assign new_n6823_1_ = ~new_n6814_ & ~new_n6816_;
  assign new_n6824_ = ~new_n6822_ & new_n6823_1_;
  assign new_n6825_ = new_n6801_ & ~new_n6824_;
  assign n612 = ~new_n6802_ & ~new_n6825_;
  assign new_n6827_ = ng1970 & ng1312;
  assign new_n6828_1_ = ng1973 & ng1315;
  assign new_n6829_ = ng1967 & ng1309;
  assign new_n6830_ = ~new_n6827_ & ~new_n6828_1_;
  assign new_n6831_ = ~new_n6829_ & new_n6830_;
  assign new_n6832_ = ng1312 & ng1951;
  assign new_n6833_1_ = ng1315 & ng1953;
  assign new_n6834_ = ng1949 & ng1309;
  assign new_n6835_ = ~new_n6832_ & ~new_n6833_1_;
  assign n1074 = ~new_n6834_ & new_n6835_;
  assign new_n6837_ = ng1904 & ~n1074;
  assign new_n6838_1_ = ng185 & new_n6837_;
  assign new_n6839_ = new_n6831_ & ~new_n6838_1_;
  assign new_n6840_ = ~new_n5366_ & ~new_n6839_;
  assign new_n6841_ = ng1315 & ~new_n6840_;
  assign new_n6842_ = ~ng1973 & ~ng1315;
  assign n617 = ~new_n6841_ & ~new_n6842_;
  assign new_n6844_ = ng1312 & ng1762;
  assign new_n6845_ = ng1315 & ng1764;
  assign new_n6846_ = ng1760 & ng1309;
  assign new_n6847_ = ~new_n6844_ & ~new_n6845_;
  assign new_n6848_1_ = ~new_n6846_ & new_n6847_;
  assign new_n6849_ = ng1312 & ng1747;
  assign new_n6850_ = ng1315 & ng1749;
  assign new_n6851_ = ng1309 & ng1745;
  assign new_n6852_ = ~new_n6849_ & ~new_n6850_;
  assign new_n6853_1_ = ~new_n6851_ & new_n6852_;
  assign new_n6854_ = ~new_n6821_ & ~new_n6848_1_;
  assign new_n6855_ = new_n6853_1_ & new_n6854_;
  assign new_n6856_ = new_n6812_ & new_n6855_;
  assign new_n6857_ = ng1312 & ng1732;
  assign new_n6858_1_ = ng1315 & ng1734;
  assign new_n6859_ = ng1730 & ng1309;
  assign new_n6860_ = ~new_n6857_ & ~new_n6858_1_;
  assign new_n6861_ = ~new_n6859_ & new_n6860_;
  assign new_n6862_ = new_n6807_ & new_n6853_1_;
  assign new_n6863_1_ = new_n6861_ & new_n6862_;
  assign new_n6864_ = ~new_n6821_ & new_n6863_1_;
  assign new_n6865_ = ng1312 & ng1777;
  assign new_n6866_ = ng1315 & ng1705;
  assign new_n6867_ = ng1309 & ng1775;
  assign new_n6868_1_ = ~new_n6865_ & ~new_n6866_;
  assign new_n6869_ = ~new_n6867_ & new_n6868_1_;
  assign new_n6870_ = new_n6821_ & new_n6869_;
  assign new_n6871_ = new_n6807_ & new_n6870_;
  assign new_n6872_ = ~new_n6812_ & new_n6871_;
  assign new_n6873_1_ = ~new_n6856_ & ~new_n6864_;
  assign new_n6874_ = ~new_n6872_ & new_n6873_1_;
  assign new_n6875_ = ~new_n6807_ & new_n6853_1_;
  assign new_n6876_ = ~new_n6861_ & new_n6875_;
  assign new_n6877_1_ = new_n6812_ & new_n6876_;
  assign new_n6878_ = ng1312 & ~ng1966;
  assign new_n6879_ = ng1315 & ~ng1964;
  assign new_n6880_ = ~ng1965 & ng1309;
  assign new_n6881_ = ~new_n6878_ & ~new_n6879_;
  assign new_n6882_1_ = ~new_n6880_ & new_n6881_;
  assign new_n6883_ = ~new_n6848_1_ & ~new_n6861_;
  assign new_n6884_ = ~new_n6853_1_ & new_n6883_;
  assign new_n6885_ = ~new_n6882_1_ & new_n6884_;
  assign new_n6886_ = ~new_n6821_ & new_n6848_1_;
  assign new_n6887_1_ = new_n6861_ & new_n6886_;
  assign new_n6888_ = ~new_n6812_ & new_n6887_1_;
  assign new_n6889_ = new_n6874_ & ~new_n6877_1_;
  assign new_n6890_ = ~new_n6885_ & ~new_n6888_;
  assign new_n6891_ = new_n6889_ & new_n6890_;
  assign new_n6892_1_ = new_n6821_ & new_n6882_1_;
  assign new_n6893_ = new_n6812_ & new_n6892_1_;
  assign new_n6894_ = new_n6848_1_ & new_n6893_;
  assign new_n6895_ = ~new_n6861_ & new_n6894_;
  assign new_n6896_ = new_n6807_ & new_n6821_;
  assign new_n6897_1_ = new_n6812_ & new_n6896_;
  assign new_n6898_ = ~new_n6853_1_ & new_n6897_1_;
  assign new_n6899_ = ~new_n6869_ & new_n6898_;
  assign new_n6900_ = ~new_n6861_ & new_n6899_;
  assign new_n6901_ = ~new_n6807_ & new_n6861_;
  assign new_n6902_1_ = ~new_n6812_ & new_n6901_;
  assign new_n6903_ = ~new_n6869_ & new_n6902_1_;
  assign new_n6904_ = ~new_n6853_1_ & new_n6903_;
  assign new_n6905_ = ~new_n6812_ & new_n6892_1_;
  assign new_n6906_ = ~new_n6853_1_ & new_n6905_;
  assign new_n6907_1_ = ~new_n6848_1_ & new_n6906_;
  assign new_n6908_ = new_n6861_ & new_n6907_1_;
  assign new_n6909_ = ~new_n6895_ & ~new_n6900_;
  assign new_n6910_ = ~new_n6904_ & ~new_n6908_;
  assign new_n6911_ = new_n6909_ & new_n6910_;
  assign new_n6912_1_ = new_n6891_ & new_n6911_;
  assign new_n6913_ = ~new_n6807_ & ~new_n6861_;
  assign new_n6914_ = new_n6812_ & new_n6913_;
  assign new_n6915_ = ~new_n6848_1_ & new_n6914_;
  assign new_n6916_ = ~new_n6853_1_ & new_n6915_;
  assign new_n6917_1_ = new_n6807_ & ~new_n6861_;
  assign new_n6918_ = ~new_n6821_ & new_n6917_1_;
  assign new_n6919_ = ~new_n6869_ & new_n6918_;
  assign new_n6920_ = ~new_n6853_1_ & new_n6919_;
  assign new_n6921_ = new_n6821_ & new_n6853_1_;
  assign new_n6922_1_ = new_n6861_ & new_n6921_;
  assign new_n6923_ = ~new_n6812_ & new_n6922_1_;
  assign new_n6924_ = new_n6821_ & new_n6861_;
  assign new_n6925_ = new_n6812_ & new_n6924_;
  assign new_n6926_ = ~new_n6848_1_ & new_n6925_;
  assign new_n6927_1_ = ~new_n6853_1_ & new_n6926_;
  assign new_n6928_ = ~new_n6920_ & ~new_n6923_;
  assign new_n6929_ = ~new_n6927_1_ & new_n6928_;
  assign new_n6930_ = ~new_n6861_ & new_n6882_1_;
  assign new_n6931_1_ = ~new_n6812_ & new_n6930_;
  assign new_n6932_ = ~new_n6848_1_ & new_n6931_1_;
  assign new_n6933_ = new_n6853_1_ & new_n6932_;
  assign new_n6934_ = ~new_n6916_ & new_n6929_;
  assign new_n6935_ = ~new_n6933_ & new_n6934_;
  assign new_n6936_1_ = ~new_n6869_ & ~new_n6882_1_;
  assign new_n6937_ = new_n6861_ & new_n6936_1_;
  assign new_n6938_ = ~new_n6812_ & new_n6937_;
  assign new_n6939_ = new_n6848_1_ & ~new_n6861_;
  assign new_n6940_ = ~new_n6853_1_ & new_n6939_;
  assign new_n6941_1_ = ~new_n6821_ & new_n6940_;
  assign new_n6942_ = ~new_n6812_ & new_n6876_;
  assign new_n6943_ = new_n6807_ & new_n6861_;
  assign new_n6944_ = new_n6821_ & new_n6943_;
  assign new_n6945_ = new_n6848_1_ & new_n6944_;
  assign new_n6946_1_ = ~new_n6853_1_ & new_n6945_;
  assign new_n6947_ = ~new_n6941_1_ & ~new_n6942_;
  assign new_n6948_ = ~new_n6946_1_ & new_n6947_;
  assign new_n6949_ = new_n6869_ & new_n6882_1_;
  assign new_n6950_ = ~new_n6861_ & new_n6949_;
  assign new_n6951_1_ = new_n6812_ & new_n6950_;
  assign new_n6952_ = ~new_n6938_ & new_n6948_;
  assign new_n6953_ = ~new_n6951_1_ & new_n6952_;
  assign new_n6954_ = new_n6848_1_ & new_n6861_;
  assign new_n6955_ = ~new_n6882_1_ & new_n6954_;
  assign new_n6956_1_ = new_n6807_ & new_n6848_1_;
  assign new_n6957_ = ~new_n6861_ & new_n6956_1_;
  assign new_n6958_ = ~new_n6821_ & new_n6957_;
  assign new_n6959_ = ~new_n6807_ & new_n6869_;
  assign new_n6960_ = new_n6812_ & new_n6959_;
  assign new_n6961_1_ = ~new_n6807_ & ~new_n6848_1_;
  assign new_n6962_ = new_n6853_1_ & new_n6961_1_;
  assign new_n6963_ = ~new_n6812_ & new_n6962_;
  assign new_n6964_ = ~new_n6955_ & ~new_n6958_;
  assign new_n6965_ = ~new_n6960_ & ~new_n6963_;
  assign new_n6966_1_ = new_n6964_ & new_n6965_;
  assign new_n6967_ = new_n6935_ & new_n6953_;
  assign new_n6968_ = new_n6966_1_ & new_n6967_;
  assign new_n6969_ = ~new_n6912_1_ & new_n6968_;
  assign new_n6970_ = new_n6839_ & new_n6969_;
  assign new_n6971_1_ = ng1947 & ng1312;
  assign new_n6972_ = ng1315 & ng1870;
  assign new_n6973_ = ng1945 & ng1309;
  assign new_n6974_ = ~new_n6971_1_ & ~new_n6972_;
  assign n1552 = ~new_n6973_ & new_n6974_;
  assign new_n6976_1_ = ng185 & ~n1552;
  assign new_n6977_ = ng1922 & new_n6976_1_;
  assign new_n6978_ = ng1979 & ng1312;
  assign new_n6979_ = ng1315 & ng1982;
  assign new_n6980_ = ng1976 & ng1309;
  assign new_n6981_1_ = ~new_n6978_ & ~new_n6979_;
  assign new_n6982_ = ~new_n6980_ & new_n6981_1_;
  assign new_n6983_ = ~new_n6977_ & new_n6982_;
  assign new_n6984_ = new_n6968_ & new_n6983_;
  assign new_n6985_ = ~new_n6839_ & new_n6984_;
  assign new_n6986_1_ = ~new_n6970_ & ~new_n6985_;
  assign new_n6987_ = new_n5366_ & new_n6986_1_;
  assign new_n6988_ = ~new_n5366_ & new_n6785_;
  assign new_n6989_ = ~new_n6987_ & ~new_n6988_;
  assign new_n6990_ = ng1315 & ~new_n6989_;
  assign new_n6991_1_ = ~ng1991 & ~ng1315;
  assign n622 = ~new_n6990_ & ~new_n6991_1_;
  assign new_n6993_ = ng1312 & ng2010;
  assign new_n6994_ = ng1315 & ~ng2039;
  assign new_n6995_1_ = ng2020 & new_n6994_;
  assign new_n6996_ = ng2013 & new_n6995_1_;
  assign new_n6997_ = ng2033 & ~new_n6996_;
  assign new_n6998_ = ~ng2033 & new_n6996_;
  assign new_n6999_ = ~new_n6997_ & ~new_n6998_;
  assign n632 = ~new_n6993_ & ~new_n6999_;
  assign new_n7001_ = ng1905 & ng1918;
  assign new_n7002_ = ~ng2039 & new_n7001_;
  assign new_n7003_ = ng1309 & new_n7002_;
  assign new_n7004_1_ = ~ng2082 & ~new_n7003_;
  assign new_n7005_ = ng2013 & new_n7003_;
  assign n637 = ~new_n7004_1_ & ~new_n7005_;
  assign new_n7007_ = ng1315 & new_n7002_;
  assign new_n7008_ = ~ng2090 & ~new_n7007_;
  assign new_n7009_1_ = ng2040 & new_n7007_;
  assign n642 = ~new_n7008_ & ~new_n7009_1_;
  assign new_n7011_ = ng1312 & new_n7002_;
  assign new_n7012_ = ~ng2104 & ~new_n7011_;
  assign new_n7013_ = ng2066 & new_n7011_;
  assign n647 = ~new_n7012_ & ~new_n7013_;
  assign new_n7015_ = ~ng2237 & ~new_n4777_1_;
  assign new_n7016_ = ~ng2252 & ng823;
  assign new_n7017_ = ~ng2250 & ng853;
  assign new_n7018_ = ~ng2251 & ng826;
  assign new_n7019_1_ = ~new_n7016_ & ~new_n7017_;
  assign new_n7020_ = ~new_n7018_ & new_n7019_1_;
  assign new_n7021_ = new_n4777_1_ & ~new_n7020_;
  assign n652 = ~new_n7015_ & ~new_n7021_;
  assign new_n7023_ = ~ng2251 & ~new_n5538_;
  assign new_n7024_1_ = ng2165 & new_n5538_;
  assign n657 = ~new_n7023_ & ~new_n7024_1_;
  assign new_n7026_ = ~ng2391 & ng823;
  assign new_n7027_ = ng853 & ~ng2392;
  assign new_n7028_ = ng826 & ~ng2390;
  assign new_n7029_1_ = ~new_n7026_ & ~new_n7027_;
  assign new_n7030_ = ~new_n7028_ & new_n7029_1_;
  assign new_n7031_ = ~ng2388 & ng823;
  assign new_n7032_ = ~ng2389 & ng853;
  assign new_n7033_1_ = ~ng2387 & ng826;
  assign new_n7034_ = ~new_n7031_ & ~new_n7032_;
  assign new_n7035_ = ~new_n7033_1_ & new_n7034_;
  assign new_n7036_ = ~ng2394 & ng823;
  assign new_n7037_ = ~ng2395 & ng853;
  assign new_n7038_1_ = ng826 & ~ng2393;
  assign new_n7039_ = ~new_n7036_ & ~new_n7037_;
  assign new_n7040_ = ~new_n7038_1_ & new_n7039_;
  assign new_n7041_ = ~new_n7030_ & new_n7035_;
  assign new_n7042_ = new_n7040_ & new_n7041_;
  assign new_n7043_1_ = new_n7030_ & new_n7035_;
  assign new_n7044_ = new_n7040_ & new_n7043_1_;
  assign new_n7045_ = ~new_n7042_ & ~new_n7044_;
  assign new_n7046_ = ng2273 & ng823;
  assign new_n7047_ = ng2276 & ng853;
  assign new_n7048_1_ = ng2270 & ng826;
  assign new_n7049_ = ~new_n7046_ & ~new_n7047_;
  assign new_n7050_ = ~new_n7048_1_ & new_n7049_;
  assign new_n7051_ = ng2318 & ng823;
  assign new_n7052_ = ng2321 & ng853;
  assign new_n7053_1_ = ng2315 & ng826;
  assign new_n7054_ = ~new_n7051_ & ~new_n7052_;
  assign new_n7055_ = ~new_n7053_1_ & new_n7054_;
  assign new_n7056_ = ng2309 & ng823;
  assign new_n7057_ = ng2312 & ng853;
  assign new_n7058_1_ = ng2306 & ng826;
  assign new_n7059_ = ~new_n7056_ & ~new_n7057_;
  assign new_n7060_ = ~new_n7058_1_ & new_n7059_;
  assign new_n7061_ = ~new_n7050_ & ~new_n7055_;
  assign new_n7062_ = ~new_n7060_ & new_n7061_;
  assign new_n7063_1_ = ng2345 & ng823;
  assign new_n7064_ = ng2348 & ng853;
  assign new_n7065_ = ng2342 & ng826;
  assign new_n7066_ = ~new_n7063_1_ & ~new_n7064_;
  assign new_n7067_ = ~new_n7065_ & new_n7066_;
  assign new_n7068_1_ = ng823 & ng2336;
  assign new_n7069_ = ng2339 & ng853;
  assign new_n7070_ = ng826 & ng2333;
  assign new_n7071_ = ~new_n7068_1_ & ~new_n7069_;
  assign new_n7072_ = ~new_n7070_ & new_n7071_;
  assign new_n7073_1_ = ng2282 & ng823;
  assign new_n7074_ = ng2285 & ng853;
  assign new_n7075_ = ng826 & ng2279;
  assign new_n7076_ = ~new_n7073_1_ & ~new_n7074_;
  assign new_n7077_ = ~new_n7075_ & new_n7076_;
  assign new_n7078_1_ = ng2327 & ng823;
  assign new_n7079_ = ng2330 & ng853;
  assign new_n7080_ = ng2324 & ng826;
  assign new_n7081_ = ~new_n7078_1_ & ~new_n7079_;
  assign new_n7082_1_ = ~new_n7080_ & new_n7081_;
  assign new_n7083_ = ng2264 & ng823;
  assign new_n7084_ = ng853 & ng2267;
  assign new_n7085_ = ng2261 & ng826;
  assign new_n7086_ = ~new_n7083_ & ~new_n7084_;
  assign new_n7087_1_ = ~new_n7085_ & new_n7086_;
  assign new_n7088_ = new_n7077_ & new_n7082_1_;
  assign new_n7089_ = new_n7087_1_ & new_n7088_;
  assign new_n7090_ = ng2291 & ng823;
  assign new_n7091_ = ng2294 & ng853;
  assign new_n7092_1_ = ng2288 & ng826;
  assign new_n7093_ = ~new_n7090_ & ~new_n7091_;
  assign new_n7094_ = ~new_n7092_1_ & new_n7093_;
  assign new_n7095_ = new_n7072_ & new_n7089_;
  assign new_n7096_ = new_n7094_ & new_n7095_;
  assign new_n7097_1_ = ng2300 & ng823;
  assign new_n7098_ = ng2303 & ng853;
  assign new_n7099_ = ng2297 & ng826;
  assign new_n7100_ = ~new_n7097_1_ & ~new_n7098_;
  assign new_n7101_ = ~new_n7099_ & new_n7100_;
  assign new_n7102_1_ = new_n7062_ & ~new_n7067_;
  assign new_n7103_ = new_n7096_ & new_n7102_1_;
  assign new_n7104_ = ~new_n7101_ & new_n7103_;
  assign new_n7105_ = new_n7042_ & new_n7104_;
  assign new_n7106_ = new_n7050_ & new_n7055_;
  assign new_n7107_1_ = new_n7060_ & new_n7106_;
  assign new_n7108_ = new_n7067_ & new_n7107_1_;
  assign new_n7109_ = new_n7096_ & new_n7108_;
  assign new_n7110_ = new_n7101_ & new_n7109_;
  assign new_n7111_ = ~new_n7042_ & new_n7110_;
  assign new_n7112_1_ = ~new_n7105_ & ~new_n7111_;
  assign new_n7113_ = ~new_n7045_ & ~new_n7112_1_;
  assign new_n7114_ = ~ng2246 & ng823;
  assign new_n7115_ = ~ng2244 & ng853;
  assign new_n7116_ = ~ng2245 & ng826;
  assign new_n7117_1_ = ~new_n7114_ & ~new_n7115_;
  assign new_n7118_ = ~new_n7116_ & new_n7117_1_;
  assign new_n7119_ = ng2170 & ~new_n7060_;
  assign new_n7120_ = ng2170 & ~new_n7119_;
  assign new_n7121_ = ~new_n7060_ & ~new_n7119_;
  assign new_n7122_1_ = ~new_n7120_ & ~new_n7121_;
  assign new_n7123_ = ng2200 & ~new_n7072_;
  assign new_n7124_ = ng2200 & ~new_n7123_;
  assign new_n7125_ = ~new_n7072_ & ~new_n7123_;
  assign new_n7126_ = ~new_n7124_ & ~new_n7125_;
  assign new_n7127_1_ = new_n7122_1_ & new_n7126_;
  assign new_n7128_ = ng2180 & ~new_n7055_;
  assign new_n7129_ = ng2180 & ~new_n7128_;
  assign new_n7130_ = ~new_n7055_ & ~new_n7128_;
  assign new_n7131_1_ = ~new_n7129_ & ~new_n7130_;
  assign new_n7132_ = ng823 & ~ng2249;
  assign new_n7133_ = ~ng2247 & ng853;
  assign new_n7134_ = ~ng2248 & ng826;
  assign new_n7135_ = ~new_n7132_ & ~new_n7133_;
  assign new_n7136_1_ = ~new_n7134_ & new_n7135_;
  assign new_n7137_ = ~new_n7067_ & ~new_n7136_1_;
  assign new_n7138_ = ~new_n7136_1_ & ~new_n7137_;
  assign new_n7139_ = ~new_n7067_ & ~new_n7137_;
  assign new_n7140_ = ~new_n7138_ & ~new_n7139_;
  assign new_n7141_1_ = new_n7131_1_ & new_n7140_;
  assign new_n7142_ = ng2190 & ~new_n7082_1_;
  assign new_n7143_ = ng2190 & ~new_n7142_;
  assign new_n7144_ = ~new_n7082_1_ & ~new_n7142_;
  assign new_n7145_1_ = ~new_n7143_ & ~new_n7144_;
  assign new_n7146_ = ~new_n7127_1_ & ~new_n7141_1_;
  assign new_n7147_ = ~new_n7145_1_ & new_n7146_;
  assign new_n7148_ = new_n7126_ & new_n7145_1_;
  assign new_n7149_ = new_n7122_1_ & new_n7131_1_;
  assign new_n7150_1_ = ~new_n7148_ & ~new_n7149_;
  assign new_n7151_ = ~new_n7140_ & new_n7150_1_;
  assign new_n7152_ = new_n7126_ & new_n7140_;
  assign new_n7153_ = new_n7131_1_ & new_n7145_1_;
  assign new_n7154_ = ~new_n7152_ & ~new_n7153_;
  assign new_n7155_1_ = ~new_n7122_1_ & new_n7154_;
  assign new_n7156_ = ~new_n7147_ & ~new_n7151_;
  assign new_n7157_ = ~new_n7155_1_ & new_n7156_;
  assign new_n7158_ = ng2257 & ~new_n7118_;
  assign new_n7159_ = ~new_n7157_ & new_n7158_;
  assign new_n7160_1_ = ng2165 & ~new_n7087_1_;
  assign new_n7161_ = ng2165 & ~new_n7160_1_;
  assign new_n7162_ = ~new_n7087_1_ & ~new_n7160_1_;
  assign new_n7163_ = ~new_n7161_ & ~new_n7162_;
  assign new_n7164_ = ng2195 & ~new_n7094_;
  assign new_n7165_1_ = ng2195 & ~new_n7164_;
  assign new_n7166_ = ~new_n7094_ & ~new_n7164_;
  assign new_n7167_ = ~new_n7165_1_ & ~new_n7166_;
  assign new_n7168_ = new_n7163_ & new_n7167_;
  assign new_n7169_ = ng2175 & ~new_n7050_;
  assign new_n7170_1_ = ng2175 & ~new_n7169_;
  assign new_n7171_ = ~new_n7050_ & ~new_n7169_;
  assign new_n7172_ = ~new_n7170_1_ & ~new_n7171_;
  assign new_n7173_ = ~new_n7020_ & ~new_n7101_;
  assign new_n7174_1_ = ~new_n7020_ & ~new_n7173_;
  assign new_n7175_ = ~new_n7101_ & ~new_n7173_;
  assign new_n7176_ = ~new_n7174_1_ & ~new_n7175_;
  assign new_n7177_ = new_n7172_ & new_n7176_;
  assign new_n7178_ = ng2185 & ~new_n7077_;
  assign new_n7179_1_ = ng2185 & ~new_n7178_;
  assign new_n7180_ = ~new_n7077_ & ~new_n7178_;
  assign new_n7181_ = ~new_n7179_1_ & ~new_n7180_;
  assign new_n7182_ = ~new_n7168_ & ~new_n7177_;
  assign new_n7183_1_ = ~new_n7181_ & new_n7182_;
  assign new_n7184_ = new_n7167_ & new_n7181_;
  assign new_n7185_ = new_n7163_ & new_n7172_;
  assign new_n7186_ = ~new_n7184_ & ~new_n7185_;
  assign new_n7187_ = ~new_n7176_ & new_n7186_;
  assign new_n7188_1_ = new_n7167_ & new_n7176_;
  assign new_n7189_ = new_n7172_ & new_n7181_;
  assign new_n7190_ = ~new_n7188_1_ & ~new_n7189_;
  assign new_n7191_ = ~new_n7163_ & new_n7190_;
  assign new_n7192_ = ~new_n7183_1_ & ~new_n7187_;
  assign new_n7193_1_ = ~new_n7191_ & new_n7192_;
  assign new_n7194_ = new_n7158_ & ~new_n7193_1_;
  assign new_n7195_ = ~new_n7159_ & ~new_n7194_;
  assign new_n7196_ = ~ng2240 & ng823;
  assign new_n7197_ = ~ng2238 & ng853;
  assign new_n7198_1_ = ~ng2239 & ng826;
  assign new_n7199_ = ~new_n7196_ & ~new_n7197_;
  assign new_n7200_ = ~new_n7198_1_ & new_n7199_;
  assign new_n7201_ = ~new_n7136_1_ & ~new_n7200_;
  assign new_n7202_ = ~new_n7200_ & ~new_n7201_;
  assign new_n7203_1_ = ~new_n7136_1_ & ~new_n7201_;
  assign new_n7204_ = ~new_n7202_ & ~new_n7203_1_;
  assign new_n7205_ = ~ng2231 & ng823;
  assign new_n7206_ = ~ng2229 & ng853;
  assign new_n7207_ = ~ng2230 & ng826;
  assign new_n7208_1_ = ~new_n7205_ & ~new_n7206_;
  assign new_n7209_ = ~new_n7207_ & new_n7208_1_;
  assign new_n7210_ = ng2195 & ~new_n7209_;
  assign new_n7211_ = ~new_n7209_ & ~new_n7210_;
  assign new_n7212_ = ng2195 & ~new_n7210_;
  assign new_n7213_1_ = ~new_n7211_ & ~new_n7212_;
  assign new_n7214_ = ng823 & ~ng2234;
  assign new_n7215_ = ng853 & ~ng2232;
  assign new_n7216_ = ng826 & ~ng2233;
  assign new_n7217_ = ~new_n7214_ & ~new_n7215_;
  assign new_n7218_1_ = ~new_n7216_ & new_n7217_;
  assign new_n7219_ = ng2200 & ~new_n7218_1_;
  assign new_n7220_ = ~new_n7218_1_ & ~new_n7219_;
  assign new_n7221_ = ng2200 & ~new_n7219_;
  assign new_n7222_ = ~new_n7220_ & ~new_n7221_;
  assign new_n7223_1_ = ng823 & ~ng2228;
  assign new_n7224_ = ng853 & ~ng2226;
  assign new_n7225_ = ng826 & ~ng2227;
  assign new_n7226_ = ~new_n7223_1_ & ~new_n7224_;
  assign new_n7227_ = ~new_n7225_ & new_n7226_;
  assign new_n7228_1_ = ng2190 & ~new_n7227_;
  assign new_n7229_ = ~new_n7227_ & ~new_n7228_1_;
  assign new_n7230_ = ng2190 & ~new_n7228_1_;
  assign new_n7231_ = ~new_n7229_ & ~new_n7230_;
  assign new_n7232_ = new_n7213_1_ & new_n7222_;
  assign new_n7233_1_ = new_n7231_ & new_n7232_;
  assign new_n7234_ = ~ng2237 & ng823;
  assign new_n7235_ = ~ng2235 & ng853;
  assign new_n7236_ = ng826 & ~ng2236;
  assign new_n7237_ = ~new_n7234_ & ~new_n7235_;
  assign new_n7238_1_ = ~new_n7236_ & new_n7237_;
  assign new_n7239_ = ~new_n7020_ & ~new_n7238_1_;
  assign new_n7240_ = ~new_n7238_1_ & ~new_n7239_;
  assign new_n7241_ = ~new_n7020_ & ~new_n7239_;
  assign new_n7242_ = ~new_n7240_ & ~new_n7241_;
  assign new_n7243_1_ = new_n7204_ & new_n7233_1_;
  assign new_n7244_ = new_n7242_ & new_n7243_1_;
  assign new_n7245_ = ng823 & ~ng2225;
  assign new_n7246_ = ng853 & ~ng2223;
  assign new_n7247_ = ng826 & ~ng2224;
  assign new_n7248_1_ = ~new_n7245_ & ~new_n7246_;
  assign new_n7249_ = ~new_n7247_ & new_n7248_1_;
  assign new_n7250_ = ng2185 & ~new_n7249_;
  assign new_n7251_ = ~new_n7249_ & ~new_n7250_;
  assign new_n7252_ = ng2185 & ~new_n7250_;
  assign new_n7253_1_ = ~new_n7251_ & ~new_n7252_;
  assign new_n7254_ = ng823 & ~ng2210;
  assign new_n7255_ = ng853 & ~ng2208;
  assign new_n7256_ = ~ng2209 & ng826;
  assign new_n7257_ = ~new_n7254_ & ~new_n7255_;
  assign new_n7258_1_ = ~new_n7256_ & new_n7257_;
  assign new_n7259_ = ng2170 & ~new_n7258_1_;
  assign new_n7260_ = ~new_n7258_1_ & ~new_n7259_;
  assign new_n7261_ = ng2170 & ~new_n7259_;
  assign new_n7262_1_ = ~new_n7260_ & ~new_n7261_;
  assign new_n7263_ = ng823 & ~ng2219;
  assign new_n7264_ = ~ng2217 & ng853;
  assign new_n7265_ = ng826 & ~ng2218;
  assign new_n7266_ = ~new_n7263_ & ~new_n7264_;
  assign new_n7267_1_ = ~new_n7265_ & new_n7266_;
  assign new_n7268_ = ng2175 & ~new_n7267_1_;
  assign new_n7269_ = ~new_n7267_1_ & ~new_n7268_;
  assign new_n7270_ = ng2175 & ~new_n7268_;
  assign new_n7271_1_ = ~new_n7269_ & ~new_n7270_;
  assign new_n7272_ = ~ng2207 & ng823;
  assign new_n7273_ = ~ng2205 & ng853;
  assign new_n7274_ = ~ng2206 & ng826;
  assign new_n7275_ = ~new_n7272_ & ~new_n7273_;
  assign new_n7276_1_ = ~new_n7274_ & new_n7275_;
  assign new_n7277_ = ng2165 & ~new_n7276_1_;
  assign new_n7278_ = ~new_n7276_1_ & ~new_n7277_;
  assign new_n7279_ = ng2165 & ~new_n7277_;
  assign new_n7280_ = ~new_n7278_ & ~new_n7279_;
  assign new_n7281_1_ = new_n7262_1_ & new_n7271_1_;
  assign new_n7282_ = new_n7280_ & new_n7281_1_;
  assign new_n7283_ = ~ng2222 & ng823;
  assign new_n7284_ = ~ng2220 & ng853;
  assign new_n7285_1_ = ~ng2221 & ng826;
  assign new_n7286_ = ~new_n7283_ & ~new_n7284_;
  assign new_n7287_ = ~new_n7285_1_ & new_n7286_;
  assign new_n7288_ = ng2180 & ~new_n7287_;
  assign new_n7289_ = ~new_n7287_ & ~new_n7288_;
  assign new_n7290_1_ = ng2180 & ~new_n7288_;
  assign new_n7291_ = ~new_n7289_ & ~new_n7290_1_;
  assign new_n7292_ = new_n7253_1_ & new_n7282_;
  assign new_n7293_ = new_n7291_ & new_n7292_;
  assign new_n7294_ = new_n7244_ & new_n7293_;
  assign new_n7295_1_ = ~new_n7118_ & new_n7195_;
  assign new_n7296_ = ng2257 & new_n7294_;
  assign new_n7297_ = new_n7295_1_ & new_n7296_;
  assign new_n7298_ = ~ng2398 & ng823;
  assign new_n7299_ = ~ng2396 & ng853;
  assign new_n7300_1_ = ~ng2397 & ng826;
  assign new_n7301_ = ~new_n7298_ & ~new_n7299_;
  assign new_n7302_ = ~new_n7300_1_ & new_n7301_;
  assign new_n7303_ = new_n7030_ & ~new_n7035_;
  assign new_n7304_1_ = new_n7040_ & new_n7303_;
  assign new_n7305_ = new_n7297_ & ~new_n7302_;
  assign new_n7306_ = new_n7304_1_ & new_n7305_;
  assign new_n7307_ = new_n7158_ & new_n7294_;
  assign new_n7308_ = ~new_n7040_ & new_n7303_;
  assign new_n7309_1_ = ~new_n7302_ & new_n7307_;
  assign new_n7310_ = new_n7308_ & new_n7309_1_;
  assign new_n7311_ = ng2257 & new_n7118_;
  assign new_n7312_ = ~new_n7035_ & new_n7311_;
  assign new_n7313_ = ~new_n7306_ & ~new_n7310_;
  assign new_n7314_1_ = ~new_n7312_ & new_n7313_;
  assign new_n7315_ = ~ng2479 & ng823;
  assign new_n7316_ = ~ng2477 & ng853;
  assign new_n7317_ = ~ng2478 & ng826;
  assign new_n7318_ = ~new_n7315_ & ~new_n7316_;
  assign new_n7319_1_ = ~new_n7317_ & new_n7318_;
  assign new_n7320_ = new_n7307_ & ~new_n7319_1_;
  assign new_n7321_ = new_n7314_1_ & ~new_n7320_;
  assign new_n7322_ = ~new_n7113_ & new_n7321_;
  assign new_n7323_ = new_n7113_ & new_n7321_;
  assign new_n7324_1_ = ng2170 & ~new_n7323_;
  assign new_n7325_ = ~new_n7042_ & new_n7323_;
  assign new_n7326_ = ~new_n7324_1_ & ~new_n7325_;
  assign new_n7327_1_ = ~new_n7322_ & new_n7326_;
  assign new_n7328_ = new_n7042_ & new_n7087_1_;
  assign new_n7329_ = ~new_n7042_ & ~new_n7087_1_;
  assign new_n7330_ = ~new_n7328_ & ~new_n7329_;
  assign new_n7331_ = ~new_n7045_ & new_n7330_;
  assign new_n7332_1_ = ~new_n7060_ & ~new_n7331_;
  assign new_n7333_ = new_n7060_ & new_n7331_;
  assign new_n7334_ = ~new_n7332_1_ & ~new_n7333_;
  assign new_n7335_1_ = new_n7322_ & new_n7334_;
  assign new_n7336_ = ~new_n7327_1_ & ~new_n7335_1_;
  assign new_n7337_ = ng853 & ~new_n7336_;
  assign new_n7338_ = ~ng2312 & ~ng853;
  assign n662 = ~new_n7337_ & ~new_n7338_;
  assign new_n7340_1_ = ng2190 & ~new_n7323_;
  assign new_n7341_ = ~new_n7322_ & ~new_n7340_1_;
  assign new_n7342_ = new_n7042_ & ~new_n7077_;
  assign new_n7343_ = ~new_n7042_ & new_n7077_;
  assign new_n7344_ = ~new_n7342_ & ~new_n7343_;
  assign new_n7345_1_ = new_n7042_ & ~new_n7060_;
  assign new_n7346_ = ~new_n7042_ & new_n7060_;
  assign new_n7347_ = ~new_n7345_1_ & ~new_n7346_;
  assign new_n7348_ = new_n7331_ & ~new_n7347_;
  assign new_n7349_ = new_n7042_ & ~new_n7055_;
  assign new_n7350_1_ = ~new_n7042_ & new_n7055_;
  assign new_n7351_ = ~new_n7349_ & ~new_n7350_1_;
  assign new_n7352_ = new_n7042_ & ~new_n7050_;
  assign new_n7353_ = ~new_n7042_ & new_n7050_;
  assign new_n7354_ = ~new_n7352_ & ~new_n7353_;
  assign new_n7355_1_ = ~new_n7351_ & ~new_n7354_;
  assign new_n7356_ = new_n7348_ & new_n7355_1_;
  assign new_n7357_ = ~new_n7344_ & new_n7356_;
  assign new_n7358_ = new_n7082_1_ & new_n7357_;
  assign new_n7359_ = ~new_n7082_1_ & ~new_n7357_;
  assign new_n7360_1_ = ~new_n7358_ & ~new_n7359_;
  assign new_n7361_ = new_n7322_ & new_n7360_1_;
  assign new_n7362_ = ~new_n7341_ & ~new_n7361_;
  assign new_n7363_ = ng823 & ~new_n7362_;
  assign new_n7364_ = ~ng2327 & ~ng823;
  assign n667 = ~new_n7363_ & ~new_n7364_;
  assign new_n7366_ = ~new_n7136_1_ & ~new_n7323_;
  assign new_n7367_ = ~new_n7325_ & ~new_n7366_;
  assign new_n7368_ = ~new_n7322_ & new_n7367_;
  assign new_n7369_ = new_n7042_ & ~new_n7101_;
  assign new_n7370_1_ = ~new_n7042_ & new_n7101_;
  assign new_n7371_ = ~new_n7369_ & ~new_n7370_1_;
  assign new_n7372_ = new_n7042_ & ~new_n7082_1_;
  assign new_n7373_ = ~new_n7042_ & new_n7082_1_;
  assign new_n7374_ = ~new_n7372_ & ~new_n7373_;
  assign new_n7375_1_ = ~new_n7344_ & ~new_n7374_;
  assign new_n7376_ = new_n7042_ & ~new_n7072_;
  assign new_n7377_ = ~new_n7042_ & new_n7072_;
  assign new_n7378_ = ~new_n7376_ & ~new_n7377_;
  assign new_n7379_1_ = new_n7042_ & ~new_n7094_;
  assign new_n7380_ = ~new_n7042_ & new_n7094_;
  assign new_n7381_ = ~new_n7379_1_ & ~new_n7380_;
  assign new_n7382_ = ~new_n7378_ & ~new_n7381_;
  assign new_n7383_ = new_n7348_ & new_n7375_1_;
  assign new_n7384_1_ = new_n7355_1_ & new_n7382_;
  assign new_n7385_ = new_n7383_ & new_n7384_1_;
  assign new_n7386_ = ~new_n7371_ & new_n7385_;
  assign new_n7387_1_ = new_n7067_ & new_n7386_;
  assign new_n7388_ = ~new_n7067_ & ~new_n7386_;
  assign new_n7389_ = ~new_n7387_1_ & ~new_n7388_;
  assign new_n7390_ = new_n7322_ & new_n7389_;
  assign new_n7391_ = ~new_n7368_ & ~new_n7390_;
  assign new_n7392_1_ = ng826 & ~new_n7391_;
  assign new_n7393_ = ~ng2342 & ~ng826;
  assign n672 = ~new_n7392_1_ & ~new_n7393_;
  assign new_n7395_ = ng2160 & new_n5128_;
  assign new_n7396_1_ = ng2156 & new_n7395_;
  assign new_n7397_ = ng2151 & new_n7396_1_;
  assign new_n7398_ = ng2147 & new_n7397_;
  assign new_n7399_ = ng2142 & new_n7398_;
  assign new_n7400_ = ng2138 & new_n7399_;
  assign new_n7401_1_ = ng2133 & new_n7400_;
  assign new_n7402_ = ng2129 & new_n7401_1_;
  assign new_n7403_ = ~ng2124 & new_n7402_;
  assign new_n7404_ = ng2124 & ~new_n7402_;
  assign new_n7405_ = ~new_n7403_ & ~new_n7404_;
  assign n677 = ~new_n5127_1_ & ~new_n7405_;
  assign new_n7407_ = new_n5125_ & ~new_n7044_;
  assign new_n7408_ = ~new_n7040_ & new_n7041_;
  assign new_n7409_ = ~new_n7407_ & ~new_n7408_;
  assign new_n7410_ = ng853 & new_n7409_;
  assign new_n7411_1_ = ~ng2436 & ~new_n7410_;
  assign new_n7412_ = ng823 & ~ng2448;
  assign new_n7413_ = ng853 & ~ng2451;
  assign new_n7414_ = ~ng2459 & ng826;
  assign new_n7415_ = ~new_n7412_ & ~new_n7413_;
  assign new_n7416_1_ = ~new_n7414_ & new_n7415_;
  assign new_n7417_ = ~ng2418 & ng823;
  assign new_n7418_ = ~ng2421 & ng853;
  assign new_n7419_ = ~ng2429 & ng826;
  assign new_n7420_ = ~new_n7417_ & ~new_n7418_;
  assign new_n7421_1_ = ~new_n7419_ & new_n7420_;
  assign new_n7422_ = ~new_n7416_1_ & new_n7421_1_;
  assign new_n7423_ = ~pg3229 & new_n7422_;
  assign new_n7424_ = ~new_n7416_1_ & ~new_n7421_1_;
  assign new_n7425_ = pg3229 & new_n7424_;
  assign new_n7426_1_ = ~ng2433 & ng823;
  assign new_n7427_ = ~ng2436 & ng853;
  assign new_n7428_ = ~ng2444 & ng826;
  assign new_n7429_ = ~new_n7426_1_ & ~new_n7427_;
  assign new_n7430_ = ~new_n7428_ & new_n7429_;
  assign new_n7431_ = new_n7416_1_ & ~new_n7430_;
  assign new_n7432_ = ~new_n7423_ & ~new_n7425_;
  assign new_n7433_ = ~new_n7431_ & new_n7432_;
  assign new_n7434_ = new_n7410_ & ~new_n7433_;
  assign n682 = ~new_n7411_1_ & ~new_n7434_;
  assign new_n7436_ = ng2495 & ng823;
  assign new_n7437_ = ng853 & ng2498;
  assign new_n7438_ = ng2492 & ng826;
  assign new_n7439_ = ~new_n7436_ & ~new_n7437_;
  assign n2815 = new_n7438_ | ~new_n7439_;
  assign new_n7441_ = ng2486 & ng823;
  assign new_n7442_ = ng2489 & ng853;
  assign new_n7443_ = ng2483 & ng826;
  assign new_n7444_ = ~new_n7441_ & ~new_n7442_;
  assign new_n7445_ = ~new_n7443_ & new_n7444_;
  assign new_n7446_ = ng2200 & ng2190;
  assign new_n7447_ = ng2195 & new_n7446_;
  assign new_n7448_ = ng2185 & new_n7447_;
  assign new_n7449_ = ng2170 & ng2180;
  assign new_n7450_ = ng2175 & new_n7449_;
  assign new_n7451_ = ng2165 & new_n7450_;
  assign new_n7452_ = new_n7448_ & new_n7451_;
  assign new_n7453_ = ~new_n7020_ & ~new_n7136_1_;
  assign new_n7454_ = new_n7452_ & new_n7453_;
  assign new_n7455_ = ~ng2503 & ng823;
  assign new_n7456_ = ~ng2501 & ng853;
  assign new_n7457_ = ng826 & ~ng2502;
  assign new_n7458_ = ~new_n7455_ & ~new_n7456_;
  assign new_n7459_ = ~new_n7457_ & new_n7458_;
  assign new_n7460_ = ~new_n7454_ & ~new_n7459_;
  assign new_n7461_ = n2815 & ~new_n7460_;
  assign new_n7462_ = ~new_n7311_ & new_n7459_;
  assign new_n7463_ = new_n7454_ & ~new_n7462_;
  assign new_n7464_ = ~n2815 & ~new_n7463_;
  assign new_n7465_ = ~new_n7461_ & ~new_n7464_;
  assign new_n7466_ = ~new_n7445_ & new_n7465_;
  assign new_n7467_ = new_n7311_ & new_n7454_;
  assign new_n7468_ = ~n2815 & ~new_n7467_;
  assign new_n7469_ = ~n2815 & ~new_n7468_;
  assign new_n7470_ = new_n7445_ & new_n7469_;
  assign new_n7471_ = ~new_n7466_ & ~new_n7470_;
  assign new_n7472_ = ng2384 & ~new_n7471_;
  assign new_n7473_ = n2815 & new_n7472_;
  assign new_n7474_ = n2815 & ~new_n7473_;
  assign new_n7475_ = new_n7472_ & ~new_n7473_;
  assign new_n7476_ = ~new_n7474_ & ~new_n7475_;
  assign new_n7477_ = ng823 & new_n7476_;
  assign new_n7478_ = ~ng2495 & ~ng823;
  assign n687 = ~new_n7477_ & ~new_n7478_;
  assign new_n7480_ = ng823 & ~ng2524;
  assign new_n7481_ = ~ng2522 & ng853;
  assign new_n7482_ = ~ng2523 & ng826;
  assign new_n7483_ = ~new_n7480_ & ~new_n7481_;
  assign new_n7484_ = ~new_n7482_ & new_n7483_;
  assign new_n7485_ = ng823 & ng2516;
  assign new_n7486_ = ng853 & ng2519;
  assign new_n7487_ = ng826 & ng2513;
  assign new_n7488_ = ~new_n7485_ & ~new_n7486_;
  assign new_n7489_ = ~new_n7487_ & new_n7488_;
  assign new_n7490_ = ng2507 & ng823;
  assign new_n7491_ = ng853 & ng2510;
  assign new_n7492_ = ng826 & ng2504;
  assign new_n7493_ = ~new_n7490_ & ~new_n7491_;
  assign new_n7494_ = ~new_n7492_ & new_n7493_;
  assign new_n7495_ = ~ng2255 & ng823;
  assign new_n7496_ = ~ng2253 & ng853;
  assign new_n7497_ = ~ng2254 & ng826;
  assign new_n7498_ = ~new_n7495_ & ~new_n7496_;
  assign new_n7499_ = ~new_n7497_ & new_n7498_;
  assign new_n7500_ = new_n7452_ & ~new_n7499_;
  assign new_n7501_ = new_n7489_ & ~new_n7494_;
  assign new_n7502_ = new_n7500_ & new_n7501_;
  assign new_n7503_ = ~new_n7489_ & new_n7494_;
  assign new_n7504_ = ~new_n7500_ & new_n7503_;
  assign new_n7505_ = ~new_n7502_ & ~new_n7504_;
  assign new_n7506_ = new_n7484_ & ~new_n7505_;
  assign new_n7507_ = ng2384 & new_n7506_;
  assign new_n7508_ = ~new_n7489_ & ~new_n7494_;
  assign new_n7509_ = ~new_n7500_ & new_n7508_;
  assign new_n7510_ = new_n7489_ & new_n7494_;
  assign new_n7511_ = new_n7500_ & new_n7510_;
  assign new_n7512_ = ~new_n7509_ & ~new_n7511_;
  assign new_n7513_ = ng2384 & ~new_n7512_;
  assign new_n7514_ = ~new_n7507_ & ~new_n7513_;
  assign new_n7515_ = ng826 & ~new_n7514_;
  assign new_n7516_ = ~ng2523 & ~new_n7515_;
  assign new_n7517_ = new_n7507_ & new_n7515_;
  assign n692 = ~new_n7516_ & ~new_n7517_;
  assign new_n7519_ = ng2628 & ng1315;
  assign new_n7520_ = ~ng2631 & ~ng1315;
  assign n712 = ~new_n7519_ & ~new_n7520_;
  assign new_n7522_ = ng853 & ~new_n7408_;
  assign new_n7523_ = ~ng2536 & ~ng853;
  assign n722 = ~new_n7522_ & ~new_n7523_;
  assign new_n7525_ = ng1312 & ng2682;
  assign new_n7526_ = ng1315 & ng2685;
  assign new_n7527_ = ng2679 & ng1309;
  assign new_n7528_ = ~new_n7525_ & ~new_n7526_;
  assign new_n7529_ = ~new_n7527_ & new_n7528_;
  assign new_n7530_ = ng1312 & ng2568;
  assign new_n7531_ = ng1315 & ng2571;
  assign new_n7532_ = ng1309 & ng2565;
  assign new_n7533_ = ~new_n7530_ & ~new_n7531_;
  assign new_n7534_ = ~new_n7532_ & new_n7533_;
  assign new_n7535_ = ~new_n7529_ & ~new_n7534_;
  assign new_n7536_ = ng1312 & ng2691;
  assign new_n7537_ = ng1315 & ng2694;
  assign new_n7538_ = ng2688 & ng1309;
  assign new_n7539_ = ~new_n7536_ & ~new_n7537_;
  assign new_n7540_ = ~new_n7538_ & new_n7539_;
  assign new_n7541_ = ng2584 & new_n7534_;
  assign new_n7542_ = ~new_n7540_ & new_n7541_;
  assign new_n7543_ = new_n5297_1_ & ~new_n7542_;
  assign n4397 = ~new_n7535_ & ~new_n7543_;
  assign new_n7545_ = ng1315 & n4397;
  assign new_n7546_ = ~ng2649 & ~new_n7545_;
  assign new_n7547_ = ng1312 & ~ng2660;
  assign new_n7548_ = ng1315 & ~ng2658;
  assign new_n7549_ = ~ng2659 & ng1309;
  assign new_n7550_ = ~new_n7547_ & ~new_n7548_;
  assign new_n7551_ = ~new_n7549_ & new_n7550_;
  assign new_n7552_ = ~ng2654 & ng1312;
  assign new_n7553_ = ng1315 & ~ng2652;
  assign new_n7554_ = ~ng2653 & ng1309;
  assign new_n7555_ = ~new_n7552_ & ~new_n7553_;
  assign new_n7556_ = ~new_n7554_ & new_n7555_;
  assign new_n7557_ = ~ng2651 & ng1312;
  assign new_n7558_ = ~ng2649 & ng1315;
  assign new_n7559_ = ng1309 & ~ng2650;
  assign new_n7560_ = ~new_n7557_ & ~new_n7558_;
  assign new_n7561_ = ~new_n7559_ & new_n7560_;
  assign new_n7562_ = pg3229 & ~new_n7561_;
  assign new_n7563_ = new_n7551_ & new_n7556_;
  assign new_n7564_ = new_n7562_ & new_n7563_;
  assign new_n7565_ = ng1312 & ~ng2657;
  assign new_n7566_ = ng1315 & ~ng2655;
  assign new_n7567_ = ~ng2656 & ng1309;
  assign new_n7568_ = ~new_n7565_ & ~new_n7566_;
  assign new_n7569_ = ~new_n7567_ & new_n7568_;
  assign new_n7570_ = new_n7562_ & ~new_n7569_;
  assign new_n7571_ = ~new_n7564_ & ~new_n7570_;
  assign new_n7572_ = new_n7551_ & ~new_n7561_;
  assign new_n7573_ = ~pg3229 & new_n7572_;
  assign new_n7574_ = ~new_n7556_ & new_n7569_;
  assign new_n7575_ = ~pg3229 & new_n7574_;
  assign new_n7576_ = pg3229 & ~new_n7551_;
  assign new_n7577_ = ~new_n7573_ & ~new_n7575_;
  assign new_n7578_ = ~new_n7576_ & new_n7577_;
  assign new_n7579_ = new_n7571_ & new_n7578_;
  assign new_n7580_ = new_n7545_ & ~new_n7579_;
  assign n732 = ~new_n7546_ & ~new_n7580_;
  assign new_n7582_ = ng2599 & ng2612;
  assign new_n7583_ = ~ng2733 & new_n7582_;
  assign new_n7584_ = ng1315 & new_n7583_;
  assign new_n7585_ = ~ng2772 & ~new_n7584_;
  assign new_n7586_ = ng2714 & new_n7584_;
  assign n737 = ~new_n7585_ & ~new_n7586_;
  assign new_n7588_ = ng1312 & new_n7583_;
  assign new_n7589_ = ~ng2786 & ~new_n7588_;
  assign new_n7590_ = ng2734 & new_n7588_;
  assign n742 = ~new_n7589_ & ~new_n7590_;
  assign new_n7592_ = ng1309 & new_n7583_;
  assign new_n7593_ = ~ng2797 & ~new_n7592_;
  assign new_n7594_ = ng2760 & new_n7592_;
  assign n747 = ~new_n7593_ & ~new_n7594_;
  assign new_n7596_ = ng1315 & ng2704;
  assign new_n7597_ = ~ng2805 & ~new_n7596_;
  assign new_n7598_ = ~new_n7529_ & new_n7596_;
  assign n752 = ~new_n7597_ & ~new_n7598_;
  assign new_n7600_ = ~ng557 & ng510;
  assign new_n7601_ = ~ng557 & ~ng510;
  assign new_n7602_ = ng525 & new_n7601_;
  assign new_n7603_ = ~new_n7600_ & ~new_n7602_;
  assign new_n7604_ = ng557 & ~ng510;
  assign new_n7605_ = ~new_n7602_ & ~new_n7604_;
  assign new_n7606_ = ng1309 & ~ng499;
  assign new_n7607_ = ~ng559 & ~n4521;
  assign new_n7608_ = ~pg563 & ~new_n7606_;
  assign new_n7609_ = new_n7607_ & new_n7608_;
  assign new_n7610_ = ~ng530 & new_n7609_;
  assign new_n7611_ = ~new_n7605_ & new_n7610_;
  assign new_n7612_ = new_n5471_ & new_n5480_;
  assign new_n7613_ = new_n5489_ & new_n7612_;
  assign new_n7614_ = ~new_n5462_ & new_n7613_;
  assign new_n7615_ = ~new_n5500_ & new_n7614_;
  assign new_n7616_ = ~ng739 & ng1312;
  assign new_n7617_ = ng1315 & ~ng737;
  assign new_n7618_ = ~ng738 & ng1309;
  assign new_n7619_ = ~new_n7616_ & ~new_n7617_;
  assign new_n7620_ = ~new_n7618_ & new_n7619_;
  assign new_n7621_ = ~new_n5422_1_ & ~new_n5431_1_;
  assign new_n7622_ = new_n5440_ & new_n7621_;
  assign new_n7623_ = new_n5413_1_ & new_n7622_;
  assign new_n7624_ = ~new_n5451_ & new_n7623_;
  assign new_n7625_ = new_n7615_ & ~new_n7620_;
  assign new_n7626_ = ~new_n5512_ & new_n7624_;
  assign new_n7627_ = new_n7625_ & new_n7626_;
  assign new_n7628_ = ~new_n5471_ & ~new_n7627_;
  assign new_n7629_ = ~new_n5302_1_ & ~new_n7628_;
  assign new_n7630_ = ~new_n7628_ & ~new_n7629_;
  assign new_n7631_ = ~new_n5302_1_ & ~new_n7629_;
  assign new_n7632_ = ~new_n7630_ & ~new_n7631_;
  assign new_n7633_ = new_n7609_ & ~new_n7632_;
  assign new_n7634_ = ng499 & new_n7633_;
  assign new_n7635_ = new_n7605_ & new_n7634_;
  assign new_n7636_ = ~new_n7611_ & ~new_n7635_;
  assign new_n7637_ = ~new_n7603_ & new_n7636_;
  assign new_n7638_ = new_n7603_ & ~new_n7605_;
  assign new_n7639_ = ~ng736 & ng1312;
  assign new_n7640_ = ~ng734 & ng1315;
  assign new_n7641_ = ng1309 & ~ng735;
  assign new_n7642_ = ~new_n7639_ & ~new_n7640_;
  assign new_n7643_ = ~new_n7641_ & new_n7642_;
  assign new_n7644_ = ~new_n7627_ & new_n7643_;
  assign new_n7645_ = ng499 & ~new_n7644_;
  assign new_n7646_ = new_n7609_ & ~new_n7645_;
  assign new_n7647_ = new_n7638_ & ~new_n7646_;
  assign new_n7648_ = new_n7603_ & new_n7647_;
  assign n757 = new_n7637_ | new_n7648_;
  assign new_n7650_ = ng1312 & ~n4521;
  assign new_n7651_ = ~ng3098 & ~ng1312;
  assign n762 = ~new_n7650_ & ~new_n7651_;
  assign new_n7653_ = ng1312 & ~n4713;
  assign new_n7654_ = ~ng3107 & ~ng1312;
  assign n767 = ~new_n7653_ & ~new_n7654_;
  assign new_n7656_ = ng1315 & ~ng2574;
  assign new_n7657_ = ~ng3088 & ~ng1315;
  assign n772 = ~new_n7656_ & ~new_n7657_;
  assign new_n7659_ = ~ng145 & ~new_n5517_1_;
  assign new_n7660_ = ng109 & new_n5517_1_;
  assign n782 = ~new_n7659_ & ~new_n7660_;
  assign new_n7662_ = ~ng154 & ~new_n5517_1_;
  assign new_n7663_ = ng121 & new_n5517_1_;
  assign n787 = ~new_n7662_ & ~new_n7663_;
  assign new_n7665_ = ng823 & ~new_n5118_;
  assign new_n7666_ = ~ng261 & ~ng823;
  assign n792 = ~new_n7665_ & ~new_n7666_;
  assign new_n7668_ = ng88 & ~new_n5129_;
  assign new_n7669_ = ~ng88 & new_n5129_;
  assign new_n7670_ = ~new_n7668_ & ~new_n7669_;
  assign n797 = ~new_n5127_1_ & ~new_n7670_;
  assign new_n7672_ = ng823 & new_n5137_1_;
  assign new_n7673_ = ~ng358 & ~new_n7672_;
  assign new_n7674_ = ~new_n5161_ & new_n7672_;
  assign n802 = ~new_n7673_ & ~new_n7674_;
  assign new_n7676_ = ng823 & new_n5204_;
  assign new_n7677_ = ~ng411 & ~ng823;
  assign n807 = ~new_n7676_ & ~new_n7677_;
  assign new_n7679_ = ng853 & new_n5239_;
  assign new_n7680_ = ~ng444 & ~ng853;
  assign n812 = ~new_n7679_ & ~new_n7680_;
  assign new_n7682_ = new_n4785_ & new_n4795_;
  assign new_n7683_ = new_n4790_ & ~new_n7682_;
  assign new_n7684_ = new_n5065_ & new_n5260_;
  assign new_n7685_ = new_n5257_1_ & ~new_n7684_;
  assign new_n7686_ = ~new_n4914_ & new_n7685_;
  assign new_n7687_ = new_n4795_ & new_n7686_;
  assign new_n7688_ = ~new_n5069_ & ~new_n5071_;
  assign new_n7689_ = ~new_n4795_ & new_n7688_;
  assign new_n7690_ = ~new_n7687_ & ~new_n7689_;
  assign new_n7691_ = new_n4785_ & new_n7690_;
  assign new_n7692_ = ~new_n4914_ & new_n5260_;
  assign new_n7693_ = ~new_n4954_ & ~new_n7692_;
  assign new_n7694_ = new_n4795_ & new_n7693_;
  assign new_n7695_ = ~new_n4795_ & ~new_n4954_;
  assign new_n7696_ = ~new_n7694_ & ~new_n7695_;
  assign new_n7697_ = ~new_n4785_ & new_n7696_;
  assign new_n7698_ = ~new_n7691_ & ~new_n7697_;
  assign new_n7699_ = ~new_n4790_ & new_n7698_;
  assign new_n7700_ = ~new_n7683_ & ~new_n7699_;
  assign new_n7701_ = ~new_n4785_ & new_n7700_;
  assign new_n7702_ = ~new_n4785_ & ~new_n7701_;
  assign new_n7703_ = new_n7700_ & ~new_n7701_;
  assign new_n7704_ = ~new_n7702_ & ~new_n7703_;
  assign new_n7705_ = ~new_n5080_ & new_n7704_;
  assign new_n7706_ = ng853 & ~new_n7705_;
  assign new_n7707_ = ~ng317 & ~ng853;
  assign n817 = ~new_n7706_ & ~new_n7707_;
  assign new_n7709_ = ng1315 & new_n5366_;
  assign new_n7710_ = ~ng554 & ~ng1315;
  assign n831 = ~new_n7709_ & ~new_n7710_;
  assign new_n7712_ = ng823 & ~new_n5136_;
  assign new_n7713_ = ~ng458 & ~ng823;
  assign n840 = ~new_n7712_ & ~new_n7713_;
  assign new_n7715_ = ng1312 & n3888;
  assign new_n7716_ = ~ng577 & ~new_n7715_;
  assign new_n7717_ = ~new_n5341_ & new_n7715_;
  assign n849 = ~new_n7716_ & ~new_n7717_;
  assign new_n7719_ = ng1315 & ~new_n5367_;
  assign new_n7720_ = ~ng593 & ~ng1315;
  assign n854 = ~new_n7719_ & ~new_n7720_;
  assign new_n7722_ = ng381 & ng1312;
  assign new_n7723_ = ng1315 & ng383;
  assign new_n7724_ = ng379 & ng1309;
  assign new_n7725_ = ~new_n7722_ & ~new_n7723_;
  assign new_n7726_ = ~new_n7724_ & new_n7725_;
  assign new_n7727_ = ng1312 & ng366;
  assign new_n7728_ = ng1315 & ng368;
  assign new_n7729_ = ng364 & ng1309;
  assign new_n7730_ = ~new_n7727_ & ~new_n7728_;
  assign new_n7731_ = ~new_n7729_ & new_n7730_;
  assign new_n7732_ = ~new_n5318_ & ~new_n7726_;
  assign new_n7733_ = new_n7731_ & new_n7732_;
  assign new_n7734_ = new_n5323_ & new_n7733_;
  assign new_n7735_ = ng1312 & ng351;
  assign new_n7736_ = ng1315 & ng353;
  assign new_n7737_ = ng349 & ng1309;
  assign new_n7738_ = ~new_n7735_ & ~new_n7736_;
  assign new_n7739_ = ~new_n7737_ & new_n7738_;
  assign new_n7740_ = new_n5331_ & new_n7731_;
  assign new_n7741_ = new_n7739_ & new_n7740_;
  assign new_n7742_ = ~new_n5318_ & new_n7741_;
  assign new_n7743_ = ng1312 & ng396;
  assign new_n7744_ = ng1315 & ng324;
  assign new_n7745_ = ng1309 & ng394;
  assign new_n7746_ = ~new_n7743_ & ~new_n7744_;
  assign new_n7747_ = ~new_n7745_ & new_n7746_;
  assign new_n7748_ = new_n5318_ & new_n7747_;
  assign new_n7749_ = new_n5331_ & new_n7748_;
  assign new_n7750_ = ~new_n5323_ & new_n7749_;
  assign new_n7751_ = ~new_n7734_ & ~new_n7742_;
  assign new_n7752_ = ~new_n7750_ & new_n7751_;
  assign new_n7753_ = ~new_n5331_ & new_n7731_;
  assign new_n7754_ = ~new_n7739_ & new_n7753_;
  assign new_n7755_ = new_n5323_ & new_n7754_;
  assign new_n7756_ = ~new_n7726_ & ~new_n7739_;
  assign new_n7757_ = ~new_n7731_ & new_n7756_;
  assign new_n7758_ = ~new_n5313_1_ & new_n7757_;
  assign new_n7759_ = ~new_n5318_ & new_n7726_;
  assign new_n7760_ = new_n7739_ & new_n7759_;
  assign new_n7761_ = ~new_n5323_ & new_n7760_;
  assign new_n7762_ = new_n7752_ & ~new_n7755_;
  assign new_n7763_ = ~new_n7758_ & ~new_n7761_;
  assign new_n7764_ = new_n7762_ & new_n7763_;
  assign new_n7765_ = new_n5323_ & new_n5325_;
  assign new_n7766_ = new_n7726_ & new_n7765_;
  assign new_n7767_ = ~new_n7739_ & new_n7766_;
  assign new_n7768_ = new_n5318_ & new_n5331_;
  assign new_n7769_ = new_n5323_ & new_n7768_;
  assign new_n7770_ = ~new_n7731_ & new_n7769_;
  assign new_n7771_ = ~new_n7747_ & new_n7770_;
  assign new_n7772_ = ~new_n7739_ & new_n7771_;
  assign new_n7773_ = ~new_n5331_ & new_n7739_;
  assign new_n7774_ = ~new_n5323_ & new_n7773_;
  assign new_n7775_ = ~new_n7747_ & new_n7774_;
  assign new_n7776_ = ~new_n7731_ & new_n7775_;
  assign new_n7777_ = ~new_n5323_ & new_n5325_;
  assign new_n7778_ = ~new_n7731_ & new_n7777_;
  assign new_n7779_ = ~new_n7726_ & new_n7778_;
  assign new_n7780_ = new_n7739_ & new_n7779_;
  assign new_n7781_ = ~new_n7767_ & ~new_n7772_;
  assign new_n7782_ = ~new_n7776_ & ~new_n7780_;
  assign new_n7783_ = new_n7781_ & new_n7782_;
  assign new_n7784_ = new_n7764_ & new_n7783_;
  assign new_n7785_ = ~new_n5331_ & ~new_n7739_;
  assign new_n7786_ = new_n5323_ & new_n7785_;
  assign new_n7787_ = ~new_n7726_ & new_n7786_;
  assign new_n7788_ = ~new_n7731_ & new_n7787_;
  assign new_n7789_ = new_n5331_ & ~new_n7739_;
  assign new_n7790_ = ~new_n5318_ & new_n7789_;
  assign new_n7791_ = ~new_n7747_ & new_n7790_;
  assign new_n7792_ = ~new_n7731_ & new_n7791_;
  assign new_n7793_ = new_n5318_ & new_n7731_;
  assign new_n7794_ = new_n7739_ & new_n7793_;
  assign new_n7795_ = ~new_n5323_ & new_n7794_;
  assign new_n7796_ = new_n5318_ & new_n7739_;
  assign new_n7797_ = new_n5323_ & new_n7796_;
  assign new_n7798_ = ~new_n7726_ & new_n7797_;
  assign new_n7799_ = ~new_n7731_ & new_n7798_;
  assign new_n7800_ = ~new_n7792_ & ~new_n7795_;
  assign new_n7801_ = ~new_n7799_ & new_n7800_;
  assign new_n7802_ = new_n5313_1_ & ~new_n7739_;
  assign new_n7803_ = ~new_n5323_ & new_n7802_;
  assign new_n7804_ = ~new_n7726_ & new_n7803_;
  assign new_n7805_ = new_n7731_ & new_n7804_;
  assign new_n7806_ = ~new_n7788_ & new_n7801_;
  assign new_n7807_ = ~new_n7805_ & new_n7806_;
  assign new_n7808_ = ~new_n5313_1_ & ~new_n7747_;
  assign new_n7809_ = new_n7739_ & new_n7808_;
  assign new_n7810_ = ~new_n5323_ & new_n7809_;
  assign new_n7811_ = new_n7726_ & ~new_n7739_;
  assign new_n7812_ = ~new_n7731_ & new_n7811_;
  assign new_n7813_ = ~new_n5318_ & new_n7812_;
  assign new_n7814_ = ~new_n5323_ & new_n7754_;
  assign new_n7815_ = new_n5331_ & new_n7739_;
  assign new_n7816_ = new_n5318_ & new_n7815_;
  assign new_n7817_ = new_n7726_ & new_n7816_;
  assign new_n7818_ = ~new_n7731_ & new_n7817_;
  assign new_n7819_ = ~new_n7813_ & ~new_n7814_;
  assign new_n7820_ = ~new_n7818_ & new_n7819_;
  assign new_n7821_ = new_n5313_1_ & new_n7747_;
  assign new_n7822_ = ~new_n7739_ & new_n7821_;
  assign new_n7823_ = new_n5323_ & new_n7822_;
  assign new_n7824_ = ~new_n7810_ & new_n7820_;
  assign new_n7825_ = ~new_n7823_ & new_n7824_;
  assign new_n7826_ = new_n7726_ & new_n7739_;
  assign new_n7827_ = ~new_n5313_1_ & new_n7826_;
  assign new_n7828_ = new_n5331_ & new_n7726_;
  assign new_n7829_ = ~new_n7739_ & new_n7828_;
  assign new_n7830_ = ~new_n5318_ & new_n7829_;
  assign new_n7831_ = ~new_n5331_ & new_n7747_;
  assign new_n7832_ = new_n5323_ & new_n7831_;
  assign new_n7833_ = ~new_n5331_ & ~new_n7726_;
  assign new_n7834_ = new_n7731_ & new_n7833_;
  assign new_n7835_ = ~new_n5323_ & new_n7834_;
  assign new_n7836_ = ~new_n7827_ & ~new_n7830_;
  assign new_n7837_ = ~new_n7832_ & ~new_n7835_;
  assign new_n7838_ = new_n7836_ & new_n7837_;
  assign new_n7839_ = new_n7807_ & new_n7825_;
  assign new_n7840_ = new_n7838_ & new_n7839_;
  assign new_n7841_ = ~new_n7784_ & new_n7840_;
  assign new_n7842_ = new_n5356_ & new_n7841_;
  assign new_n7843_ = ng1312 & ng567;
  assign new_n7844_ = ng1315 & ng489;
  assign new_n7845_ = ng565 & ng1309;
  assign new_n7846_ = ~new_n7843_ & ~new_n7844_;
  assign n6211 = ~new_n7845_ & new_n7846_;
  assign new_n7848_ = ng185 & ~n6211;
  assign new_n7849_ = ng542 & new_n7848_;
  assign new_n7850_ = ng1312 & ng599;
  assign new_n7851_ = ng1315 & ng602;
  assign new_n7852_ = ng596 & ng1309;
  assign new_n7853_ = ~new_n7850_ & ~new_n7851_;
  assign new_n7854_ = ~new_n7852_ & new_n7853_;
  assign new_n7855_ = ~new_n7849_ & new_n7854_;
  assign new_n7856_ = new_n7840_ & new_n7855_;
  assign new_n7857_ = ~new_n5356_ & new_n7856_;
  assign new_n7858_ = ~new_n7842_ & ~new_n7857_;
  assign new_n7859_ = new_n5366_ & new_n7858_;
  assign new_n7860_ = new_n5287_1_ & ~new_n5366_;
  assign new_n7861_ = ~new_n7859_ & ~new_n7860_;
  assign new_n7862_ = ng1315 & ~new_n7861_;
  assign new_n7863_ = ~ng611 & ~ng1315;
  assign n859 = ~new_n7862_ & ~new_n7863_;
  assign new_n7865_ = ng646 & new_n5384_;
  assign new_n7866_ = ng660 & ~new_n7865_;
  assign new_n7867_ = ~ng660 & new_n7865_;
  assign new_n7868_ = ~new_n7866_ & ~new_n7867_;
  assign n864 = ~new_n5380_ & ~new_n7868_;
  assign new_n7870_ = ~ng702 & ~new_n5395_;
  assign new_n7871_ = ng633 & new_n5395_;
  assign n869 = ~new_n7870_ & ~new_n7871_;
  assign new_n7873_ = ~ng715 & ~new_n5391_;
  assign new_n7874_ = ng672 & new_n5391_;
  assign n874 = ~new_n7873_ & ~new_n7874_;
  assign new_n7876_ = ~ng724 & ~new_n5391_;
  assign new_n7877_ = ng686 & new_n5391_;
  assign n879 = ~new_n7876_ & ~new_n7877_;
  assign new_n7879_ = ~ng734 & ~new_n5399_;
  assign new_n7880_ = new_n5399_ & ~new_n5514_;
  assign n884 = ~new_n7879_ & ~new_n7880_;
  assign new_n7882_ = ~ng817 & ~new_n4773_;
  assign new_n7883_ = ng785 & new_n4773_;
  assign n889 = ~new_n7882_ & ~new_n7883_;
  assign new_n7885_ = ~ng839 & ~new_n5517_1_;
  assign new_n7886_ = ng805 & new_n5517_1_;
  assign n894 = ~new_n7885_ & ~new_n7886_;
  assign new_n7888_ = ~ng848 & ~new_n5517_1_;
  assign new_n7889_ = new_n5517_1_ & ~new_n5529_;
  assign n899 = ~new_n7888_ & ~new_n7889_;
  assign new_n7891_ = ng823 & ~new_n5852_;
  assign new_n7892_ = ~ng921 & ~ng823;
  assign n904 = ~new_n7891_ & ~new_n7892_;
  assign new_n7894_ = ng793 & ~new_n5839_;
  assign new_n7895_ = ~new_n5841_ & ~new_n7894_;
  assign new_n7896_ = ~new_n5838_1_ & new_n7895_;
  assign new_n7897_ = ~new_n5566_1_ & ~new_n5864_;
  assign new_n7898_ = new_n5566_1_ & new_n5864_;
  assign new_n7899_ = ~new_n7897_ & ~new_n7898_;
  assign new_n7900_ = new_n5838_1_ & new_n7899_;
  assign new_n7901_ = ~new_n7896_ & ~new_n7900_;
  assign new_n7902_ = ng826 & ~new_n7901_;
  assign new_n7903_ = ~ng882 & ~ng826;
  assign n909 = ~new_n7902_ & ~new_n7903_;
  assign new_n7905_ = ng826 & ~new_n5878_1_;
  assign new_n7906_ = ~ng936 & ~ng826;
  assign n914 = ~new_n7905_ & ~new_n7906_;
  assign new_n7908_ = ng823 & ~new_n5907_;
  assign new_n7909_ = ~ng957 & ~ng823;
  assign n919 = ~new_n7908_ & ~new_n7909_;
  assign new_n7911_ = ng749 & ~new_n5917_;
  assign new_n7912_ = ~ng749 & new_n5917_;
  assign new_n7913_ = ~new_n7911_ & ~new_n7912_;
  assign n924 = ~new_n5127_1_ & ~new_n7913_;
  assign new_n7915_ = ng823 & new_n5925_;
  assign new_n7916_ = ~ng1075 & ~new_n7915_;
  assign new_n7917_ = ~new_n5948_1_ & new_n7915_;
  assign n929 = ~new_n7916_ & ~new_n7917_;
  assign new_n7919_ = ng823 & ~new_n5984_;
  assign new_n7920_ = ~ng1115 & ~new_n7919_;
  assign new_n7921_ = new_n5981_ & new_n7919_;
  assign n934 = ~new_n7920_ & ~new_n7921_;
  assign new_n7923_ = ng853 & ~new_n5999_;
  assign new_n7924_ = ~ng1001 & ~ng853;
  assign n939 = ~new_n7923_ & ~new_n7924_;
  assign new_n7926_ = ~ng2384 & new_n5824_;
  assign new_n7927_ = new_n5638_ & new_n5669_1_;
  assign new_n7928_ = new_n5656_ & new_n7927_;
  assign new_n7929_ = new_n5642_ & new_n7928_;
  assign new_n7930_ = new_n5679_1_ & new_n5705_;
  assign new_n7931_ = new_n5692_ & new_n7930_;
  assign new_n7932_ = new_n5683_ & new_n7931_;
  assign new_n7933_ = new_n7929_ & new_n7932_;
  assign new_n7934_ = ~new_n5634_1_ & ~new_n7933_;
  assign new_n7935_ = ng2257 & new_n7934_;
  assign new_n7936_ = ~new_n5824_ & ~new_n7935_;
  assign new_n7937_ = ~new_n7926_ & ~new_n7936_;
  assign new_n7938_ = ng853 & new_n7937_;
  assign new_n7939_ = ~ng1008 & ~new_n7938_;
  assign new_n7940_ = ~new_n5556_1_ & new_n5823_1_;
  assign new_n7941_ = new_n5546_ & new_n7940_;
  assign new_n7942_ = new_n5556_1_ & new_n5813_1_;
  assign new_n7943_ = ~new_n7941_ & ~new_n7942_;
  assign new_n7944_ = ~new_n5551_ & ~new_n7943_;
  assign new_n7945_ = new_n7938_ & new_n7944_;
  assign n944 = ~new_n7939_ & ~new_n7945_;
  assign new_n7947_ = ng740 & new_n5583_;
  assign new_n7948_ = new_n5583_ & ~new_n7947_;
  assign new_n7949_ = ng740 & ~new_n7947_;
  assign new_n7950_ = ~new_n7948_ & ~new_n7949_;
  assign new_n7951_ = ng753 & new_n5610_1_;
  assign new_n7952_ = new_n5610_1_ & ~new_n7951_;
  assign new_n7953_ = ng753 & ~new_n7951_;
  assign new_n7954_ = ~new_n7952_ & ~new_n7953_;
  assign new_n7955_ = ng749 & new_n5588_;
  assign new_n7956_ = new_n5588_ & ~new_n7955_;
  assign new_n7957_ = ng749 & ~new_n7955_;
  assign new_n7958_ = ~new_n7956_ & ~new_n7957_;
  assign new_n7959_ = ng758 & new_n5598_;
  assign new_n7960_ = new_n5598_ & ~new_n7959_;
  assign new_n7961_ = ng758 & ~new_n7959_;
  assign new_n7962_ = ~new_n7960_ & ~new_n7961_;
  assign new_n7963_ = ~new_n7954_ & ~new_n7958_;
  assign new_n7964_ = ~new_n7962_ & new_n7963_;
  assign new_n7965_ = ng744 & new_n5617_;
  assign new_n7966_ = new_n5617_ & ~new_n7965_;
  assign new_n7967_ = ng744 & ~new_n7965_;
  assign new_n7968_ = ~new_n7966_ & ~new_n7967_;
  assign new_n7969_ = ~new_n7950_ & new_n7964_;
  assign new_n7970_ = ~new_n7968_ & new_n7969_;
  assign new_n7971_ = ng762 & new_n5593_;
  assign new_n7972_ = new_n5593_ & ~new_n7971_;
  assign new_n7973_ = ng762 & ~new_n7971_;
  assign new_n7974_ = ~new_n7972_ & ~new_n7973_;
  assign new_n7975_ = ng776 & new_n5576_;
  assign new_n7976_ = new_n5576_ & ~new_n7975_;
  assign new_n7977_ = ng776 & ~new_n7975_;
  assign new_n7978_ = ~new_n7976_ & ~new_n7977_;
  assign new_n7979_ = ng771 & new_n5566_1_;
  assign new_n7980_ = new_n5566_1_ & ~new_n7979_;
  assign new_n7981_ = ng771 & ~new_n7979_;
  assign new_n7982_ = ~new_n7980_ & ~new_n7981_;
  assign new_n7983_ = ng780 & new_n5603_;
  assign new_n7984_ = new_n5603_ & ~new_n7983_;
  assign new_n7985_ = ng780 & ~new_n7983_;
  assign new_n7986_ = ~new_n7984_ & ~new_n7985_;
  assign new_n7987_ = ~new_n7978_ & ~new_n7982_;
  assign new_n7988_ = ~new_n7986_ & new_n7987_;
  assign new_n7989_ = ng767 & new_n5571_;
  assign new_n7990_ = new_n5571_ & ~new_n7989_;
  assign new_n7991_ = ng767 & ~new_n7989_;
  assign new_n7992_ = ~new_n7990_ & ~new_n7991_;
  assign new_n7993_ = ~new_n7974_ & new_n7988_;
  assign new_n7994_ = ~new_n7992_ & new_n7993_;
  assign new_n7995_ = ~new_n5924_ & new_n7970_;
  assign new_n7996_ = new_n7994_ & new_n7995_;
  assign new_n7997_ = ~new_n5125_ & new_n7996_;
  assign new_n7998_ = new_n5560_ & new_n5626_;
  assign new_n7999_ = ~new_n7997_ & ~new_n7998_;
  assign n958 = ~new_n5925_ | new_n7999_;
  assign new_n8001_ = ng823 & new_n6022_1_;
  assign new_n8002_ = ~ng1174 & ~ng823;
  assign n971 = ~new_n8001_ & ~new_n8002_;
  assign new_n8004_ = ng823 & n953;
  assign new_n8005_ = ~ng1171 & ~ng823;
  assign n976 = ~new_n8004_ & ~new_n8005_;
  assign new_n8007_ = ~ng1174 & ng1315;
  assign new_n8008_ = ~ng1175 & ng1309;
  assign new_n8009_ = ~ng1173 & ng1312;
  assign new_n8010_ = ~new_n8007_ & ~new_n8008_;
  assign n981 = ~new_n8009_ & new_n8010_;
  assign new_n8012_ = ng1312 & n2976;
  assign new_n8013_ = ~ng1269 & ~new_n8012_;
  assign new_n8014_ = ~new_n6077_1_ & new_n8012_;
  assign n986 = ~new_n8013_ & ~new_n8014_;
  assign new_n8016_ = ng1315 & ~new_n6237_;
  assign new_n8017_ = ~ng1306 & ~ng1315;
  assign n991 = ~new_n8016_ & ~new_n8017_;
  assign new_n8019_ = ~ng1193 & ng1192;
  assign new_n8020_ = ng506 & ~ng507;
  assign new_n8021_ = ~ng1312 & ng520;
  assign new_n8022_ = ~ng1312 & ~new_n8021_;
  assign new_n8023_ = ~ng506 & new_n8022_;
  assign n4186 = ~new_n8020_ & ~new_n8023_;
  assign new_n8025_ = ng1312 & n4186;
  assign new_n8026_ = ng1206 & ~ng1312;
  assign new_n8027_ = ~new_n8025_ & ~new_n8026_;
  assign new_n8028_ = ~ng1192 & new_n8027_;
  assign n996 = ~new_n8019_ & ~new_n8028_;
  assign new_n8030_ = ng1352 & new_n6248_;
  assign new_n8031_ = ~ng1365 & new_n8030_;
  assign new_n8032_ = ng1365 & ~new_n8030_;
  assign new_n8033_ = ~new_n8031_ & ~new_n8032_;
  assign n1000 = ~new_n6241_ & ~new_n8033_;
  assign new_n8035_ = ~ng1391 & ~new_n6259_1_;
  assign new_n8036_ = ng1339 & new_n6259_1_;
  assign n1005 = ~new_n8035_ & ~new_n8036_;
  assign new_n8038_ = ~ng1404 & ~new_n6255_;
  assign new_n8039_ = ng1352 & new_n6255_;
  assign n1010 = ~new_n8038_ & ~new_n8039_;
  assign new_n8041_ = ~ng1413 & ~new_n6255_;
  assign new_n8042_ = ng1378 & new_n6255_;
  assign n1015 = ~new_n8041_ & ~new_n8042_;
  assign new_n8044_ = ng1315 & ~new_n6267_;
  assign new_n8045_ = ~ng1423 & ~new_n8044_;
  assign new_n8046_ = ng1316 & new_n8044_;
  assign n1020 = ~new_n8045_ & ~new_n8046_;
  assign new_n8048_ = ~ng1523 & ~new_n4773_;
  assign new_n8049_ = ng1481 & new_n4773_;
  assign n1025 = ~new_n8048_ & ~new_n8049_;
  assign new_n8051_ = ~ng1539 & ~new_n5517_1_;
  assign new_n8052_ = ng1506 & new_n5517_1_;
  assign n1030 = ~new_n8051_ & ~new_n8052_;
  assign new_n8054_ = ~ng1551 & ~new_n5538_;
  assign new_n8055_ = new_n5538_ & ~new_n6282_;
  assign n1035 = ~new_n8054_ & ~new_n8055_;
  assign new_n8057_ = ng1491 & ~new_n6587_;
  assign new_n8058_ = ~new_n6586_ & ~new_n8057_;
  assign new_n8059_ = ~new_n6336_1_ & ~new_n6615_;
  assign new_n8060_ = new_n6336_1_ & new_n6615_;
  assign new_n8061_ = ~new_n8059_ & ~new_n8060_;
  assign new_n8062_ = new_n6586_ & new_n8061_;
  assign new_n8063_ = ~new_n8058_ & ~new_n8062_;
  assign new_n8064_ = ng826 & ~new_n8063_;
  assign new_n8065_ = ~ng1585 & ~ng826;
  assign n1040 = ~new_n8064_ & ~new_n8065_;
  assign new_n8067_ = ng1453 & new_n6628_;
  assign new_n8068_ = ~ng1448 & new_n8067_;
  assign new_n8069_ = ng1448 & ~new_n8067_;
  assign new_n8070_ = ~new_n8068_ & ~new_n8069_;
  assign n1045 = ~new_n5127_1_ & ~new_n8070_;
  assign new_n8072_ = ng826 & new_n6635_;
  assign new_n8073_ = ~ng1750 & ~new_n8072_;
  assign new_n8074_ = ~new_n6659_ & new_n8072_;
  assign n1050 = ~new_n8073_ & ~new_n8074_;
  assign new_n8076_ = ng823 & new_n6702_;
  assign new_n8077_ = ~ng1801 & ~ng823;
  assign n1055 = ~new_n8076_ & ~new_n8077_;
  assign new_n8079_ = ng823 & new_n6737_;
  assign new_n8080_ = ~ng1822 & ~ng823;
  assign n1060 = ~new_n8079_ & ~new_n8080_;
  assign new_n8082_ = ng853 & ~new_n6771_;
  assign new_n8083_ = ~ng1701 & ~ng853;
  assign n1065 = ~new_n8082_ & ~new_n8083_;
  assign new_n8085_ = ng823 & ~new_n6572_;
  assign new_n8086_ = ~ng1859 & ~ng823;
  assign n1083 = ~new_n8085_ & ~new_n8086_;
  assign new_n8088_ = ng1312 & n2736;
  assign new_n8089_ = ~ng1960 & ~new_n8088_;
  assign new_n8090_ = ~new_n6824_ & new_n8088_;
  assign n1092 = ~new_n8089_ & ~new_n8090_;
  assign new_n8092_ = ng1312 & ~new_n6840_;
  assign new_n8093_ = ~ng1970 & ~ng1312;
  assign n1097 = ~new_n8092_ & ~new_n8093_;
  assign new_n8095_ = ng1890 & new_n6796_;
  assign new_n8096_ = new_n6790_ & ~new_n8095_;
  assign new_n8097_ = ~new_n6790_ & new_n8096_;
  assign new_n8098_ = ~new_n6790_ & ~new_n8097_;
  assign new_n8099_ = new_n8096_ & ~new_n8097_;
  assign new_n8100_ = ~new_n8098_ & ~new_n8099_;
  assign new_n8101_ = ng1309 & ~new_n8100_;
  assign new_n8102_ = ~ng1871 & ~ng1309;
  assign n1102 = ~new_n8101_ & ~new_n8102_;
  assign new_n8104_ = ng2033 & new_n6996_;
  assign new_n8105_ = ~ng2026 & new_n8104_;
  assign new_n8106_ = ng2026 & ~new_n8104_;
  assign new_n8107_ = ~new_n8105_ & ~new_n8106_;
  assign n1112 = ~new_n6993_ & ~new_n8107_;
  assign new_n8109_ = ~ng2078 & ~new_n7007_;
  assign new_n8110_ = ng2020 & new_n7007_;
  assign n1117 = ~new_n8109_ & ~new_n8110_;
  assign new_n8112_ = ~ng2094 & ~new_n7003_;
  assign new_n8113_ = ng2052 & new_n7003_;
  assign n1122 = ~new_n8112_ & ~new_n8113_;
  assign new_n8115_ = ~ng2103 & ~new_n7003_;
  assign new_n8116_ = ng2066 & new_n7003_;
  assign n1127 = ~new_n8115_ & ~new_n8116_;
  assign new_n8118_ = ~ng2235 & ~new_n4773_;
  assign new_n8119_ = new_n4773_ & ~new_n7020_;
  assign n1132 = ~new_n8118_ & ~new_n8119_;
  assign new_n8121_ = ng853 & n1621;
  assign new_n8122_ = ~ng2247 & ~new_n8121_;
  assign new_n8123_ = ng2170 & new_n8121_;
  assign n1137 = ~new_n8122_ & ~new_n8123_;
  assign new_n8125_ = ng2175 & ~new_n7323_;
  assign new_n8126_ = ~new_n7325_ & ~new_n8125_;
  assign new_n8127_ = ~new_n7322_ & new_n8126_;
  assign new_n8128_ = ~new_n7050_ & ~new_n7348_;
  assign new_n8129_ = new_n7050_ & new_n7348_;
  assign new_n8130_ = ~new_n8128_ & ~new_n8129_;
  assign new_n8131_ = new_n7322_ & new_n8130_;
  assign new_n8132_ = ~new_n8127_ & ~new_n8131_;
  assign new_n8133_ = ng826 & ~new_n8132_;
  assign new_n8134_ = ~ng2270 & ~ng826;
  assign n1142 = ~new_n8133_ & ~new_n8134_;
  assign new_n8136_ = ng826 & ~new_n7362_;
  assign new_n8137_ = ~ng2324 & ~ng826;
  assign n1147 = ~new_n8136_ & ~new_n8137_;
  assign new_n8139_ = ng823 & ~new_n7391_;
  assign new_n8140_ = ~ng2345 & ~ng823;
  assign n1152 = ~new_n8139_ & ~new_n8140_;
  assign new_n8142_ = ng2129 & ~new_n7401_1_;
  assign new_n8143_ = ~ng2129 & new_n7401_1_;
  assign new_n8144_ = ~new_n8142_ & ~new_n8143_;
  assign n1157 = ~new_n5127_1_ & ~new_n8144_;
  assign new_n8146_ = ng826 & new_n7409_;
  assign new_n8147_ = ~ng2459 & ~new_n8146_;
  assign new_n8148_ = ~ng2463 & ng823;
  assign new_n8149_ = ~ng2466 & ng853;
  assign new_n8150_ = ~ng2473 & ng826;
  assign new_n8151_ = ~new_n8148_ & ~new_n8149_;
  assign new_n8152_ = ~new_n8150_ & new_n8151_;
  assign new_n8153_ = new_n7430_ & new_n8152_;
  assign new_n8154_ = pg3229 & ~new_n7421_1_;
  assign new_n8155_ = new_n8153_ & new_n8154_;
  assign new_n8156_ = ~pg3229 & new_n7421_1_;
  assign new_n8157_ = new_n8153_ & new_n8156_;
  assign new_n8158_ = ~new_n8155_ & ~new_n8157_;
  assign new_n8159_ = ~new_n7421_1_ & ~new_n7430_;
  assign new_n8160_ = ~pg3229 & new_n8159_;
  assign new_n8161_ = new_n7421_1_ & ~new_n7430_;
  assign new_n8162_ = pg3229 & new_n8161_;
  assign new_n8163_ = ~new_n8160_ & ~new_n8162_;
  assign new_n8164_ = new_n8158_ & new_n8163_;
  assign new_n8165_ = new_n8146_ & ~new_n8164_;
  assign n1162 = ~new_n8147_ & ~new_n8165_;
  assign new_n8167_ = ng826 & new_n7476_;
  assign new_n8168_ = ~ng2492 & ~ng826;
  assign n1167 = ~new_n8167_ & ~new_n8168_;
  assign new_n8170_ = new_n7035_ & new_n7040_;
  assign new_n8171_ = new_n7040_ & ~new_n7194_;
  assign new_n8172_ = ng2384 & ~new_n7159_;
  assign new_n8173_ = new_n8171_ & new_n8172_;
  assign new_n8174_ = new_n7030_ & ~new_n8173_;
  assign new_n8175_ = new_n7122_1_ & new_n7153_;
  assign new_n8176_ = new_n7140_ & new_n8175_;
  assign new_n8177_ = new_n7126_ & new_n8176_;
  assign new_n8178_ = new_n7163_ & new_n7189_;
  assign new_n8179_ = new_n7176_ & new_n8178_;
  assign new_n8180_ = new_n7167_ & new_n8179_;
  assign new_n8181_ = new_n8177_ & new_n8180_;
  assign new_n8182_ = ng2257 & new_n8181_;
  assign new_n8183_ = ~new_n7118_ & new_n8182_;
  assign new_n8184_ = ~new_n7311_ & ~new_n8183_;
  assign new_n8185_ = new_n7040_ & ~new_n8184_;
  assign new_n8186_ = ~new_n7118_ & ~new_n8181_;
  assign new_n8187_ = ng2257 & new_n8186_;
  assign new_n8188_ = ~new_n7194_ & ~new_n8187_;
  assign new_n8189_ = ~new_n7159_ & new_n8188_;
  assign new_n8190_ = ~new_n7040_ & ~new_n8189_;
  assign new_n8191_ = ~new_n8185_ & ~new_n8190_;
  assign new_n8192_ = ~new_n7030_ & new_n8191_;
  assign new_n8193_ = ~new_n8174_ & ~new_n8192_;
  assign new_n8194_ = ~new_n7035_ & new_n8193_;
  assign new_n8195_ = ~new_n8170_ & ~new_n8194_;
  assign new_n8196_ = ~new_n7040_ & new_n8195_;
  assign new_n8197_ = ~new_n7040_ & ~new_n8196_;
  assign new_n8198_ = new_n8195_ & ~new_n8196_;
  assign new_n8199_ = ~new_n8197_ & ~new_n8198_;
  assign new_n8200_ = ~new_n7320_ & ~new_n8199_;
  assign new_n8201_ = ng823 & ~new_n8200_;
  assign new_n8202_ = ~ng2394 & ~ng823;
  assign n1172 = ~new_n8201_ & ~new_n8202_;
  assign new_n8204_ = ~ng2628 & ~ng1315;
  assign n1190 = ~new_n7709_ & ~new_n8204_;
  assign new_n8206_ = ng823 & ~new_n7408_;
  assign new_n8207_ = ~ng2533 & ~ng823;
  assign n1199 = ~new_n8206_ & ~new_n8207_;
  assign new_n8209_ = ng1312 & n4397;
  assign new_n8210_ = ~ng2651 & ~new_n8209_;
  assign new_n8211_ = ~new_n7579_ & new_n8209_;
  assign n1208 = ~new_n8210_ & ~new_n8211_;
  assign new_n8213_ = ng1312 & ng2704;
  assign new_n8214_ = ng1315 & ~ng2733;
  assign new_n8215_ = ng2714 & new_n8214_;
  assign new_n8216_ = ng2707 & new_n8215_;
  assign new_n8217_ = ng2727 & ~new_n8216_;
  assign new_n8218_ = ~ng2727 & new_n8216_;
  assign new_n8219_ = ~new_n8217_ & ~new_n8218_;
  assign n1213 = ~new_n8213_ & ~new_n8219_;
  assign new_n8221_ = ~ng2784 & ~new_n7584_;
  assign new_n8222_ = ng2734 & new_n7584_;
  assign n1218 = ~new_n8221_ & ~new_n8222_;
  assign new_n8224_ = ~ng2793 & ~new_n7584_;
  assign new_n8225_ = ng2753 & new_n7584_;
  assign n1223 = ~new_n8224_ & ~new_n8225_;
  assign new_n8227_ = ~ng2809 & ~new_n7592_;
  assign new_n8228_ = ng1312 & ~ng2804;
  assign new_n8229_ = ng1315 & ~ng2802;
  assign new_n8230_ = ~ng2803 & ng1309;
  assign new_n8231_ = ~new_n8228_ & ~new_n8229_;
  assign new_n8232_ = ~new_n8230_ & new_n8231_;
  assign new_n8233_ = ~ng2786 & ng1312;
  assign new_n8234_ = ~ng2784 & ng1315;
  assign new_n8235_ = ~ng2785 & ng1309;
  assign new_n8236_ = ~new_n8233_ & ~new_n8234_;
  assign new_n8237_ = ~new_n8235_ & new_n8236_;
  assign new_n8238_ = ~ng2734 & ~new_n8237_;
  assign new_n8239_ = ~new_n8237_ & ~new_n8238_;
  assign new_n8240_ = ~ng2734 & ~new_n8238_;
  assign new_n8241_ = ~new_n8239_ & ~new_n8240_;
  assign new_n8242_ = ~ng2777 & ng1312;
  assign new_n8243_ = ng1315 & ~ng2775;
  assign new_n8244_ = ~ng2776 & ng1309;
  assign new_n8245_ = ~new_n8242_ & ~new_n8243_;
  assign new_n8246_ = ~new_n8244_ & new_n8245_;
  assign new_n8247_ = ~ng2707 & ~new_n8246_;
  assign new_n8248_ = ~new_n8246_ & ~new_n8247_;
  assign new_n8249_ = ~ng2707 & ~new_n8247_;
  assign new_n8250_ = ~new_n8248_ & ~new_n8249_;
  assign new_n8251_ = ng1312 & ~ng2780;
  assign new_n8252_ = ng1315 & ~ng2778;
  assign new_n8253_ = ng1309 & ~ng2779;
  assign new_n8254_ = ~new_n8251_ & ~new_n8252_;
  assign new_n8255_ = ~new_n8253_ & new_n8254_;
  assign new_n8256_ = ~ng2727 & ~new_n8255_;
  assign new_n8257_ = ~new_n8255_ & ~new_n8256_;
  assign new_n8258_ = ~ng2727 & ~new_n8256_;
  assign new_n8259_ = ~new_n8257_ & ~new_n8258_;
  assign new_n8260_ = ng1312 & ~ng2774;
  assign new_n8261_ = ~ng2772 & ng1315;
  assign new_n8262_ = ~ng2773 & ng1309;
  assign new_n8263_ = ~new_n8260_ & ~new_n8261_;
  assign new_n8264_ = ~new_n8262_ & new_n8263_;
  assign new_n8265_ = ~ng2714 & ~new_n8264_;
  assign new_n8266_ = ~new_n8264_ & ~new_n8265_;
  assign new_n8267_ = ~ng2714 & ~new_n8265_;
  assign new_n8268_ = ~new_n8266_ & ~new_n8267_;
  assign new_n8269_ = ~new_n8250_ & ~new_n8259_;
  assign new_n8270_ = ~new_n8268_ & new_n8269_;
  assign new_n8271_ = ng1312 & ~ng2783;
  assign new_n8272_ = ng1315 & ~ng2781;
  assign new_n8273_ = ~ng2782 & ng1309;
  assign new_n8274_ = ~new_n8271_ & ~new_n8272_;
  assign new_n8275_ = ~new_n8273_ & new_n8274_;
  assign new_n8276_ = ~ng2720 & ~new_n8275_;
  assign new_n8277_ = ~new_n8275_ & ~new_n8276_;
  assign new_n8278_ = ~ng2720 & ~new_n8276_;
  assign new_n8279_ = ~new_n8277_ & ~new_n8278_;
  assign new_n8280_ = ~new_n8241_ & new_n8270_;
  assign new_n8281_ = ~new_n8279_ & new_n8280_;
  assign new_n8282_ = ng1312 & ~ng2801;
  assign new_n8283_ = ng1315 & ~ng2799;
  assign new_n8284_ = ng1309 & ~ng2800;
  assign new_n8285_ = ~new_n8282_ & ~new_n8283_;
  assign new_n8286_ = ~new_n8284_ & new_n8285_;
  assign new_n8287_ = ~ng2766 & ~new_n8286_;
  assign new_n8288_ = ~new_n8286_ & ~new_n8287_;
  assign new_n8289_ = ~ng2766 & ~new_n8287_;
  assign new_n8290_ = ~new_n8288_ & ~new_n8289_;
  assign new_n8291_ = ng1312 & ~ng2792;
  assign new_n8292_ = ng1315 & ~ng2790;
  assign new_n8293_ = ng1309 & ~ng2791;
  assign new_n8294_ = ~new_n8291_ & ~new_n8292_;
  assign new_n8295_ = ~new_n8293_ & new_n8294_;
  assign new_n8296_ = ~ng2740 & ~new_n8295_;
  assign new_n8297_ = ~new_n8295_ & ~new_n8296_;
  assign new_n8298_ = ~ng2740 & ~new_n8296_;
  assign new_n8299_ = ~new_n8297_ & ~new_n8298_;
  assign new_n8300_ = ~ng2795 & ng1312;
  assign new_n8301_ = ~ng2793 & ng1315;
  assign new_n8302_ = ~ng2794 & ng1309;
  assign new_n8303_ = ~new_n8300_ & ~new_n8301_;
  assign new_n8304_ = ~new_n8302_ & new_n8303_;
  assign new_n8305_ = ~ng2753 & ~new_n8304_;
  assign new_n8306_ = ~new_n8304_ & ~new_n8305_;
  assign new_n8307_ = ~ng2753 & ~new_n8305_;
  assign new_n8308_ = ~new_n8306_ & ~new_n8307_;
  assign new_n8309_ = ng1312 & ~ng2789;
  assign new_n8310_ = ng1315 & ~ng2787;
  assign new_n8311_ = ng1309 & ~ng2788;
  assign new_n8312_ = ~new_n8309_ & ~new_n8310_;
  assign new_n8313_ = ~new_n8311_ & new_n8312_;
  assign new_n8314_ = ~ng2746 & ~new_n8313_;
  assign new_n8315_ = ~new_n8313_ & ~new_n8314_;
  assign new_n8316_ = ~ng2746 & ~new_n8314_;
  assign new_n8317_ = ~new_n8315_ & ~new_n8316_;
  assign new_n8318_ = ~new_n8299_ & ~new_n8308_;
  assign new_n8319_ = ~new_n8317_ & new_n8318_;
  assign new_n8320_ = ng1312 & ~ng2798;
  assign new_n8321_ = ng1315 & ~ng2796;
  assign new_n8322_ = ~ng2797 & ng1309;
  assign new_n8323_ = ~new_n8320_ & ~new_n8321_;
  assign new_n8324_ = ~new_n8322_ & new_n8323_;
  assign new_n8325_ = ~ng2760 & ~new_n8324_;
  assign new_n8326_ = ~new_n8324_ & ~new_n8325_;
  assign new_n8327_ = ~ng2760 & ~new_n8325_;
  assign new_n8328_ = ~new_n8326_ & ~new_n8327_;
  assign new_n8329_ = ~new_n8290_ & new_n8319_;
  assign new_n8330_ = ~new_n8328_ & new_n8329_;
  assign new_n8331_ = new_n8281_ & new_n8330_;
  assign new_n8332_ = ng1312 & ~ng2807;
  assign new_n8333_ = ~ng2805 & ng1315;
  assign new_n8334_ = ng1309 & ~ng2806;
  assign new_n8335_ = ~new_n8332_ & ~new_n8333_;
  assign new_n8336_ = ~new_n8334_ & new_n8335_;
  assign new_n8337_ = new_n8232_ & ~new_n8331_;
  assign new_n8338_ = new_n8336_ & new_n8337_;
  assign new_n8339_ = new_n7592_ & ~new_n8338_;
  assign n1228 = ~new_n8227_ & ~new_n8339_;
  assign new_n8341_ = ~ng529 & new_n7609_;
  assign new_n8342_ = ~new_n7605_ & new_n8341_;
  assign new_n8343_ = ~new_n5480_ & ~new_n7627_;
  assign new_n8344_ = ~new_n5287_1_ & ~new_n8343_;
  assign new_n8345_ = ~new_n8343_ & ~new_n8344_;
  assign new_n8346_ = ~new_n5287_1_ & ~new_n8344_;
  assign new_n8347_ = ~new_n8345_ & ~new_n8346_;
  assign new_n8348_ = new_n7609_ & ~new_n8347_;
  assign new_n8349_ = ng499 & new_n8348_;
  assign new_n8350_ = new_n7605_ & new_n8349_;
  assign new_n8351_ = ~new_n8342_ & ~new_n8350_;
  assign new_n8352_ = ~new_n7603_ & new_n8351_;
  assign new_n8353_ = new_n7609_ & new_n7645_;
  assign new_n8354_ = new_n7638_ & ~new_n8353_;
  assign new_n8355_ = new_n7603_ & new_n8354_;
  assign n1233 = new_n8352_ | new_n8355_;
  assign new_n8357_ = ng1315 & ~n4521;
  assign new_n8358_ = ~ng3099 & ~ng1315;
  assign n1238 = ~new_n8357_ & ~new_n8358_;
  assign new_n8360_ = ng1312 & ~ng499;
  assign new_n8361_ = ~ng3158 & ~ng1312;
  assign n1243 = ~new_n8360_ & ~new_n8361_;
  assign new_n8363_ = ng1315 & ~ng1880;
  assign new_n8364_ = ~ng3179 & ~ng1315;
  assign n1248 = ~new_n8363_ & ~new_n8364_;
  assign new_n8366_ = ~ng164 & ~new_n4777_1_;
  assign new_n8367_ = new_n4777_1_ & ~new_n4891_;
  assign n1258 = ~new_n8366_ & ~new_n8367_;
  assign new_n8369_ = ~ng178 & ~new_n5538_;
  assign new_n8370_ = new_n5180_ & new_n5538_;
  assign n1263 = ~new_n8369_ & ~new_n8370_;
  assign new_n8372_ = ng853 & ~new_n5118_;
  assign new_n8373_ = ~ng264 & ~ng853;
  assign n1268 = ~new_n8372_ & ~new_n8373_;
  assign new_n8375_ = ng83 & new_n5130_;
  assign new_n8376_ = ng79 & new_n8375_;
  assign new_n8377_ = ~ng74 & new_n8376_;
  assign new_n8378_ = ng74 & ~new_n8376_;
  assign new_n8379_ = ~new_n8377_ & ~new_n8378_;
  assign n1273 = ~new_n5127_1_ & ~new_n8379_;
  assign new_n8381_ = ~ng343 & ~new_n7672_;
  assign new_n8382_ = ~ng388 & ng823;
  assign new_n8383_ = ~ng391 & ng853;
  assign new_n8384_ = ~ng398 & ng826;
  assign new_n8385_ = ~new_n8382_ & ~new_n8383_;
  assign new_n8386_ = ~new_n8384_ & new_n8385_;
  assign new_n8387_ = pg3229 & ~new_n5149_;
  assign new_n8388_ = new_n5158_ & new_n8386_;
  assign new_n8389_ = new_n8387_ & new_n8388_;
  assign new_n8390_ = ~new_n5144_ & new_n8387_;
  assign new_n8391_ = ~new_n8389_ & ~new_n8390_;
  assign new_n8392_ = ~new_n5149_ & new_n8386_;
  assign new_n8393_ = ~pg3229 & new_n8392_;
  assign new_n8394_ = ~pg3229 & new_n5159_;
  assign new_n8395_ = pg3229 & ~new_n8386_;
  assign new_n8396_ = ~new_n8393_ & ~new_n8394_;
  assign new_n8397_ = ~new_n8395_ & new_n8396_;
  assign new_n8398_ = new_n8391_ & new_n8397_;
  assign new_n8399_ = new_n7672_ & ~new_n8398_;
  assign n1278 = ~new_n8381_ & ~new_n8399_;
  assign new_n8401_ = ng826 & new_n5204_;
  assign new_n8402_ = ~ng408 & ~ng826;
  assign n1283 = ~new_n8401_ & ~new_n8402_;
  assign new_n8404_ = new_n5217_1_ & ~new_n5233_;
  assign new_n8405_ = ng2384 & new_n8404_;
  assign new_n8406_ = ~new_n5212_1_ & ~new_n5222_1_;
  assign new_n8407_ = ~new_n5228_ & new_n8406_;
  assign new_n8408_ = new_n5212_1_ & new_n5222_1_;
  assign new_n8409_ = new_n5228_ & new_n8408_;
  assign new_n8410_ = ~new_n8407_ & ~new_n8409_;
  assign new_n8411_ = ng2384 & ~new_n8410_;
  assign new_n8412_ = ~new_n8405_ & ~new_n8411_;
  assign new_n8413_ = ng826 & ~new_n8412_;
  assign new_n8414_ = ~ng448 & ~new_n8413_;
  assign new_n8415_ = new_n8405_ & new_n8413_;
  assign n1288 = ~new_n8414_ & ~new_n8415_;
  assign new_n8417_ = ng826 & ~new_n5136_;
  assign new_n8418_ = ~ng455 & ~ng826;
  assign n1318 = ~new_n8417_ & ~new_n8418_;
  assign new_n8420_ = ng1315 & ~ng478;
  assign new_n8421_ = ng1309 & ~ng479;
  assign new_n8422_ = ng1312 & ~ng477;
  assign new_n8423_ = ~new_n8420_ & ~new_n8421_;
  assign n1323 = ~new_n8422_ & new_n8423_;
  assign new_n8425_ = ~ng580 & ~new_n7715_;
  assign new_n8426_ = new_n5323_ & ~new_n5331_;
  assign new_n8427_ = ~pg3229 & new_n8426_;
  assign new_n8428_ = ~new_n5323_ & ~new_n5331_;
  assign new_n8429_ = pg3229 & new_n8428_;
  assign new_n8430_ = ~new_n8427_ & ~new_n8429_;
  assign new_n8431_ = ~new_n5336_ & new_n8430_;
  assign new_n8432_ = new_n7715_ & ~new_n8431_;
  assign n1328 = ~new_n8425_ & ~new_n8432_;
  assign new_n8434_ = ~ng584 & ~new_n5307_;
  assign new_n8435_ = ~pg3229 & ~new_n5323_;
  assign new_n8436_ = new_n7768_ & new_n8435_;
  assign new_n8437_ = pg3229 & new_n5323_;
  assign new_n8438_ = new_n7768_ & new_n8437_;
  assign new_n8439_ = ~new_n8436_ & ~new_n8438_;
  assign new_n8440_ = new_n5307_ & ~new_n8439_;
  assign n1333 = ~new_n8434_ & ~new_n8440_;
  assign new_n8442_ = ng1312 & ~new_n7861_;
  assign new_n8443_ = ~ng608 & ~ng1312;
  assign n1338 = ~new_n8442_ & ~new_n8443_;
  assign new_n8445_ = ng660 & new_n7865_;
  assign new_n8446_ = ~ng672 & new_n8445_;
  assign new_n8447_ = ng672 & ~new_n8445_;
  assign new_n8448_ = ~new_n8446_ & ~new_n8447_;
  assign n1343 = ~new_n5380_ & ~new_n8448_;
  assign new_n8450_ = ~ng705 & ~new_n5395_;
  assign new_n8451_ = ng653 & new_n5395_;
  assign n1348 = ~new_n8450_ & ~new_n8451_;
  assign new_n8453_ = ~ng712 & ~new_n5391_;
  assign new_n8454_ = ng660 & new_n5391_;
  assign n1353 = ~new_n8453_ & ~new_n8454_;
  assign new_n8456_ = ~ng723 & ~new_n5395_;
  assign new_n8457_ = ng686 & new_n5395_;
  assign n1358 = ~new_n8456_ & ~new_n8457_;
  assign new_n8459_ = ~ng630 & ~new_n5390_;
  assign new_n8460_ = ng1309 & ~new_n8459_;
  assign new_n8461_ = ~ng738 & ~new_n8460_;
  assign new_n8462_ = ng630 & new_n8460_;
  assign n1363 = ~new_n8461_ & ~new_n8462_;
  assign new_n8464_ = ~ng820 & ~new_n4773_;
  assign new_n8465_ = ng789 & new_n4773_;
  assign n1368 = ~new_n8464_ & ~new_n8465_;
  assign new_n8467_ = ~ng836 & ~new_n5517_1_;
  assign new_n8468_ = ng801 & new_n5517_1_;
  assign n1373 = ~new_n8467_ & ~new_n8468_;
  assign new_n8470_ = ~ng844 & ~new_n4773_;
  assign new_n8471_ = ng813 & new_n4773_;
  assign n1378 = ~new_n8470_ & ~new_n8471_;
  assign new_n8473_ = ng823 & ~new_n7901_;
  assign new_n8474_ = ~ng885 & ~ng823;
  assign n1383 = ~new_n8473_ & ~new_n8474_;
  assign new_n8476_ = ng809 & ~new_n5839_;
  assign new_n8477_ = ~new_n5838_1_ & ~new_n8476_;
  assign new_n8478_ = new_n5872_ & new_n5891_;
  assign new_n8479_ = ~new_n5610_1_ & ~new_n8478_;
  assign new_n8480_ = new_n5610_1_ & new_n8478_;
  assign new_n8481_ = ~new_n8479_ & ~new_n8480_;
  assign new_n8482_ = new_n5838_1_ & new_n8481_;
  assign new_n8483_ = ~new_n8477_ & ~new_n8482_;
  assign new_n8484_ = ng826 & ~new_n8483_;
  assign new_n8485_ = ~ng900 & ~ng826;
  assign n1388 = ~new_n8484_ & ~new_n8485_;
  assign new_n8487_ = ~new_n5529_ & ~new_n5839_;
  assign new_n8488_ = ~new_n5841_ & ~new_n8487_;
  assign new_n8489_ = ~new_n5838_1_ & new_n8488_;
  assign new_n8490_ = ~new_n5617_ & ~new_n5901_;
  assign new_n8491_ = new_n5617_ & new_n5901_;
  assign new_n8492_ = ~new_n8490_ & ~new_n8491_;
  assign new_n8493_ = new_n5838_1_ & new_n8492_;
  assign new_n8494_ = ~new_n8489_ & ~new_n8493_;
  assign new_n8495_ = ng823 & ~new_n8494_;
  assign new_n8496_ = ~ng912 & ~ng823;
  assign n1393 = ~new_n8495_ & ~new_n8496_;
  assign new_n8498_ = ~ng753 & new_n5916_;
  assign new_n8499_ = ng753 & ~new_n5916_;
  assign new_n8500_ = ~new_n8498_ & ~new_n8499_;
  assign n1398 = ~new_n5127_1_ & ~new_n8500_;
  assign new_n8502_ = ng853 & new_n5925_;
  assign new_n8503_ = ~ng1078 & ~new_n8502_;
  assign new_n8504_ = ~new_n5948_1_ & new_n8502_;
  assign n1403 = ~new_n8503_ & ~new_n8504_;
  assign new_n8506_ = ng1119 & ng823;
  assign new_n8507_ = ng1122 & ng853;
  assign new_n8508_ = ng1116 & ng826;
  assign new_n8509_ = ~new_n8506_ & ~new_n8507_;
  assign new_n8510_ = ~new_n8508_ & new_n8509_;
  assign new_n8511_ = ~ng867 & ng823;
  assign new_n8512_ = ~ng865 & ng853;
  assign new_n8513_ = ~ng866 & ng826;
  assign new_n8514_ = ~new_n8511_ & ~new_n8512_;
  assign new_n8515_ = ~new_n8513_ & new_n8514_;
  assign new_n8516_ = new_n5967_1_ & ~new_n8515_;
  assign new_n8517_ = ~new_n8510_ & new_n8516_;
  assign new_n8518_ = new_n8516_ & ~new_n8517_;
  assign new_n8519_ = ~new_n8510_ & ~new_n8517_;
  assign new_n8520_ = ~new_n8518_ & ~new_n8519_;
  assign new_n8521_ = ng2384 & ~new_n8520_;
  assign new_n8522_ = ~new_n8510_ & ~new_n8521_;
  assign new_n8523_ = ~new_n8510_ & ~new_n8522_;
  assign new_n8524_ = ~new_n8521_ & ~new_n8522_;
  assign new_n8525_ = ~new_n8523_ & ~new_n8524_;
  assign new_n8526_ = ng823 & ~new_n8525_;
  assign new_n8527_ = ~ng1119 & ~ng823;
  assign n1408 = ~new_n8526_ & ~new_n8527_;
  assign new_n8529_ = ng823 & ~ng1136;
  assign new_n8530_ = ~ng1134 & ng853;
  assign new_n8531_ = ng826 & ~ng1135;
  assign new_n8532_ = ~new_n8529_ & ~new_n8530_;
  assign new_n8533_ = ~new_n8531_ & new_n8532_;
  assign new_n8534_ = new_n6022_1_ & ~new_n8510_;
  assign new_n8535_ = new_n8516_ & new_n8534_;
  assign new_n8536_ = ~new_n6022_1_ & new_n8510_;
  assign new_n8537_ = ~new_n8516_ & new_n8536_;
  assign new_n8538_ = ~new_n8535_ & ~new_n8537_;
  assign new_n8539_ = new_n8533_ & ~new_n8538_;
  assign new_n8540_ = ng2384 & new_n8539_;
  assign new_n8541_ = ~new_n6022_1_ & ~new_n8510_;
  assign new_n8542_ = ~new_n8516_ & new_n8541_;
  assign new_n8543_ = new_n6022_1_ & new_n8510_;
  assign new_n8544_ = new_n8516_ & new_n8543_;
  assign new_n8545_ = ~new_n8542_ & ~new_n8544_;
  assign new_n8546_ = ng2384 & ~new_n8545_;
  assign new_n8547_ = ~new_n8540_ & ~new_n8546_;
  assign new_n8548_ = ng853 & ~new_n8547_;
  assign new_n8549_ = ~ng1134 & ~new_n8548_;
  assign new_n8550_ = new_n8540_ & new_n8548_;
  assign n1413 = ~new_n8549_ & ~new_n8550_;
  assign new_n8552_ = ng823 & new_n7937_;
  assign new_n8553_ = ~ng1010 & ~new_n8552_;
  assign new_n8554_ = new_n7944_ & new_n8552_;
  assign n1418 = ~new_n8553_ & ~new_n8554_;
  assign new_n8556_ = ng853 & new_n6022_1_;
  assign new_n8557_ = ~ng1175 & ~ng853;
  assign n1438 = ~new_n8556_ & ~new_n8557_;
  assign new_n8559_ = ng823 & ~new_n5560_;
  assign new_n8560_ = ~ng1155 & ~ng823;
  assign n1443 = ~new_n8559_ & ~new_n8560_;
  assign new_n8562_ = ng1309 & n2976;
  assign new_n8563_ = ~ng1268 & ~new_n8562_;
  assign new_n8564_ = ~new_n6077_1_ & new_n8562_;
  assign n1453 = ~new_n8563_ & ~new_n8564_;
  assign new_n8566_ = ~new_n6147_1_ & new_n6231_;
  assign new_n8567_ = new_n6173_ & new_n8566_;
  assign new_n8568_ = new_n6160_ & new_n6231_;
  assign new_n8569_ = ~new_n6173_ & new_n8568_;
  assign new_n8570_ = ~new_n8567_ & ~new_n8569_;
  assign new_n8571_ = new_n5366_ & new_n8570_;
  assign new_n8572_ = ~new_n5366_ & new_n6033_;
  assign new_n8573_ = ~new_n8571_ & ~new_n8572_;
  assign new_n8574_ = ng1309 & ~new_n8573_;
  assign new_n8575_ = ~ng1291 & ~ng1309;
  assign n1458 = ~new_n8574_ & ~new_n8575_;
  assign new_n8577_ = ~ng1402 & ~new_n6263_;
  assign new_n8578_ = ng1352 & new_n6263_;
  assign n1473 = ~new_n8577_ & ~new_n8578_;
  assign new_n8580_ = ~ng1416 & ~new_n6241_;
  assign new_n8581_ = ~new_n6044_ & new_n6241_;
  assign n1478 = ~new_n8580_ & ~new_n8581_;
  assign new_n8583_ = ~ng1420 & ~new_n6263_;
  assign new_n8584_ = ~ng1416 & ng1312;
  assign new_n8585_ = ng1315 & ~ng1414;
  assign new_n8586_ = ~ng1415 & ng1309;
  assign new_n8587_ = ~new_n8584_ & ~new_n8585_;
  assign new_n8588_ = ~new_n8586_ & new_n8587_;
  assign new_n8589_ = ng1312 & ~ng1398;
  assign new_n8590_ = ng1315 & ~ng1396;
  assign new_n8591_ = ng1309 & ~ng1397;
  assign new_n8592_ = ~new_n8589_ & ~new_n8590_;
  assign new_n8593_ = ~new_n8591_ & new_n8592_;
  assign new_n8594_ = ~ng1346 & ~new_n8593_;
  assign new_n8595_ = ~new_n8593_ & ~new_n8594_;
  assign new_n8596_ = ~ng1346 & ~new_n8594_;
  assign new_n8597_ = ~new_n8595_ & ~new_n8596_;
  assign new_n8598_ = ng1312 & ~ng1389;
  assign new_n8599_ = ng1315 & ~ng1387;
  assign new_n8600_ = ng1309 & ~ng1388;
  assign new_n8601_ = ~new_n8598_ & ~new_n8599_;
  assign new_n8602_ = ~new_n8600_ & new_n8601_;
  assign new_n8603_ = ~ng1319 & ~new_n8602_;
  assign new_n8604_ = ~new_n8602_ & ~new_n8603_;
  assign new_n8605_ = ~ng1319 & ~new_n8603_;
  assign new_n8606_ = ~new_n8604_ & ~new_n8605_;
  assign new_n8607_ = ~ng1392 & ng1312;
  assign new_n8608_ = ng1315 & ~ng1390;
  assign new_n8609_ = ~ng1391 & ng1309;
  assign new_n8610_ = ~new_n8607_ & ~new_n8608_;
  assign new_n8611_ = ~new_n8609_ & new_n8610_;
  assign new_n8612_ = ~ng1339 & ~new_n8611_;
  assign new_n8613_ = ~new_n8611_ & ~new_n8612_;
  assign new_n8614_ = ~ng1339 & ~new_n8612_;
  assign new_n8615_ = ~new_n8613_ & ~new_n8614_;
  assign new_n8616_ = ng1312 & ~ng1386;
  assign new_n8617_ = ng1315 & ~ng1384;
  assign new_n8618_ = ng1309 & ~ng1385;
  assign new_n8619_ = ~new_n8616_ & ~new_n8617_;
  assign new_n8620_ = ~new_n8618_ & new_n8619_;
  assign new_n8621_ = ~ng1326 & ~new_n8620_;
  assign new_n8622_ = ~new_n8620_ & ~new_n8621_;
  assign new_n8623_ = ~ng1326 & ~new_n8621_;
  assign new_n8624_ = ~new_n8622_ & ~new_n8623_;
  assign new_n8625_ = ~new_n8606_ & ~new_n8615_;
  assign new_n8626_ = ~new_n8624_ & new_n8625_;
  assign new_n8627_ = ng1312 & ~ng1395;
  assign new_n8628_ = ng1315 & ~ng1393;
  assign new_n8629_ = ng1309 & ~ng1394;
  assign new_n8630_ = ~new_n8627_ & ~new_n8628_;
  assign new_n8631_ = ~new_n8629_ & new_n8630_;
  assign new_n8632_ = ~ng1332 & ~new_n8631_;
  assign new_n8633_ = ~new_n8631_ & ~new_n8632_;
  assign new_n8634_ = ~ng1332 & ~new_n8632_;
  assign new_n8635_ = ~new_n8633_ & ~new_n8634_;
  assign new_n8636_ = ~new_n8597_ & new_n8626_;
  assign new_n8637_ = ~new_n8635_ & new_n8636_;
  assign new_n8638_ = ~ng1413 & ng1312;
  assign new_n8639_ = ~ng1411 & ng1315;
  assign new_n8640_ = ng1309 & ~ng1412;
  assign new_n8641_ = ~new_n8638_ & ~new_n8639_;
  assign new_n8642_ = ~new_n8640_ & new_n8641_;
  assign new_n8643_ = ~ng1378 & ~new_n8642_;
  assign new_n8644_ = ~new_n8642_ & ~new_n8643_;
  assign new_n8645_ = ~ng1378 & ~new_n8643_;
  assign new_n8646_ = ~new_n8644_ & ~new_n8645_;
  assign new_n8647_ = ~ng1404 & ng1312;
  assign new_n8648_ = ng1315 & ~ng1402;
  assign new_n8649_ = ~ng1403 & ng1309;
  assign new_n8650_ = ~new_n8647_ & ~new_n8648_;
  assign new_n8651_ = ~new_n8649_ & new_n8650_;
  assign new_n8652_ = ~ng1352 & ~new_n8651_;
  assign new_n8653_ = ~new_n8651_ & ~new_n8652_;
  assign new_n8654_ = ~ng1352 & ~new_n8652_;
  assign new_n8655_ = ~new_n8653_ & ~new_n8654_;
  assign new_n8656_ = ng1312 & ~ng1407;
  assign new_n8657_ = ng1315 & ~ng1405;
  assign new_n8658_ = ~ng1406 & ng1309;
  assign new_n8659_ = ~new_n8656_ & ~new_n8657_;
  assign new_n8660_ = ~new_n8658_ & new_n8659_;
  assign new_n8661_ = ~ng1365 & ~new_n8660_;
  assign new_n8662_ = ~new_n8660_ & ~new_n8661_;
  assign new_n8663_ = ~ng1365 & ~new_n8661_;
  assign new_n8664_ = ~new_n8662_ & ~new_n8663_;
  assign new_n8665_ = ng1312 & ~ng1401;
  assign new_n8666_ = ng1315 & ~ng1399;
  assign new_n8667_ = ~ng1400 & ng1309;
  assign new_n8668_ = ~new_n8665_ & ~new_n8666_;
  assign new_n8669_ = ~new_n8667_ & new_n8668_;
  assign new_n8670_ = ~ng1358 & ~new_n8669_;
  assign new_n8671_ = ~new_n8669_ & ~new_n8670_;
  assign new_n8672_ = ~ng1358 & ~new_n8670_;
  assign new_n8673_ = ~new_n8671_ & ~new_n8672_;
  assign new_n8674_ = ~new_n8655_ & ~new_n8664_;
  assign new_n8675_ = ~new_n8673_ & new_n8674_;
  assign new_n8676_ = ng1312 & ~ng1410;
  assign new_n8677_ = ng1315 & ~ng1408;
  assign new_n8678_ = ~ng1409 & ng1309;
  assign new_n8679_ = ~new_n8676_ & ~new_n8677_;
  assign new_n8680_ = ~new_n8678_ & new_n8679_;
  assign new_n8681_ = ~ng1372 & ~new_n8680_;
  assign new_n8682_ = ~new_n8680_ & ~new_n8681_;
  assign new_n8683_ = ~ng1372 & ~new_n8681_;
  assign new_n8684_ = ~new_n8682_ & ~new_n8683_;
  assign new_n8685_ = ~new_n8646_ & new_n8675_;
  assign new_n8686_ = ~new_n8684_ & new_n8685_;
  assign new_n8687_ = new_n8637_ & new_n8686_;
  assign new_n8688_ = ng1312 & ~ng1419;
  assign new_n8689_ = ng1315 & ~ng1417;
  assign new_n8690_ = ~ng1418 & ng1309;
  assign new_n8691_ = ~new_n8688_ & ~new_n8689_;
  assign new_n8692_ = ~new_n8690_ & new_n8691_;
  assign new_n8693_ = new_n8588_ & ~new_n8687_;
  assign new_n8694_ = new_n8692_ & new_n8693_;
  assign new_n8695_ = new_n6263_ & ~new_n8694_;
  assign n1483 = ~new_n8583_ & ~new_n8695_;
  assign new_n8697_ = ~ng1525 & ~new_n4777_1_;
  assign new_n8698_ = ng1481 & new_n4777_1_;
  assign n1488 = ~new_n8697_ & ~new_n8698_;
  assign new_n8700_ = ~ng1540 & ~new_n4777_1_;
  assign new_n8701_ = ng1506 & new_n4777_1_;
  assign n1493 = ~new_n8700_ & ~new_n8701_;
  assign new_n8703_ = ~ng1554 & ~new_n5538_;
  assign new_n8704_ = ng1476 & new_n5538_;
  assign n1498 = ~new_n8703_ & ~new_n8704_;
  assign new_n8706_ = ng1471 & ~new_n6587_;
  assign new_n8707_ = ~new_n6586_ & ~new_n8706_;
  assign new_n8708_ = ~new_n6304_1_ & new_n6346_;
  assign new_n8709_ = new_n6304_1_ & ~new_n6346_;
  assign new_n8710_ = ~new_n8708_ & ~new_n8709_;
  assign new_n8711_ = new_n6586_ & new_n8710_;
  assign new_n8712_ = ~new_n8707_ & ~new_n8711_;
  assign new_n8713_ = ng853 & ~new_n8712_;
  assign new_n8714_ = ~ng1573 & ~ng853;
  assign n1503 = ~new_n8713_ & ~new_n8714_;
  assign new_n8716_ = ng1448 & new_n8067_;
  assign new_n8717_ = ng1444 & ~new_n8716_;
  assign new_n8718_ = ~ng1444 & new_n8716_;
  assign new_n8719_ = ~new_n8717_ & ~new_n8718_;
  assign n1508 = ~new_n5127_1_ & ~new_n8719_;
  assign new_n8721_ = ~ng1765 & ~new_n8072_;
  assign new_n8722_ = ~ng1769 & ng823;
  assign new_n8723_ = ng853 & ~ng1772;
  assign new_n8724_ = ~ng1779 & ng826;
  assign new_n8725_ = ~new_n8722_ & ~new_n8723_;
  assign new_n8726_ = ~new_n8724_ & new_n8725_;
  assign new_n8727_ = new_n6656_ & new_n8726_;
  assign new_n8728_ = pg3229 & ~new_n6647_;
  assign new_n8729_ = new_n8727_ & new_n8728_;
  assign new_n8730_ = ~pg3229 & new_n6647_;
  assign new_n8731_ = new_n8727_ & new_n8730_;
  assign new_n8732_ = ~new_n8729_ & ~new_n8731_;
  assign new_n8733_ = ~new_n6647_ & ~new_n6656_;
  assign new_n8734_ = ~pg3229 & new_n8733_;
  assign new_n8735_ = new_n6647_ & ~new_n6656_;
  assign new_n8736_ = pg3229 & new_n8735_;
  assign new_n8737_ = ~new_n8734_ & ~new_n8736_;
  assign new_n8738_ = new_n8732_ & new_n8737_;
  assign new_n8739_ = new_n8072_ & ~new_n8738_;
  assign n1513 = ~new_n8721_ & ~new_n8739_;
  assign new_n8741_ = ~new_n6680_ & new_n6685_;
  assign new_n8742_ = n5082 & new_n8741_;
  assign new_n8743_ = ~new_n6575_1_ & new_n6680_;
  assign new_n8744_ = new_n6685_ & new_n8743_;
  assign new_n8745_ = ~n5082 & new_n8744_;
  assign new_n8746_ = ~new_n8742_ & ~new_n8745_;
  assign new_n8747_ = ~new_n6671_1_ & new_n8746_;
  assign new_n8748_ = n5082 & new_n6680_;
  assign new_n8749_ = ~n5082 & ~new_n8743_;
  assign new_n8750_ = ~new_n8748_ & ~new_n8749_;
  assign new_n8751_ = new_n6671_1_ & new_n8750_;
  assign new_n8752_ = ~new_n8747_ & ~new_n8751_;
  assign new_n8753_ = ng2384 & ~new_n8752_;
  assign new_n8754_ = ~new_n6671_1_ & new_n8753_;
  assign new_n8755_ = ~new_n6671_1_ & ~new_n8754_;
  assign new_n8756_ = new_n8753_ & ~new_n8754_;
  assign new_n8757_ = ~new_n8755_ & ~new_n8756_;
  assign new_n8758_ = ng823 & new_n8757_;
  assign new_n8759_ = ~ng1792 & ~ng823;
  assign n1518 = ~new_n8758_ & ~new_n8759_;
  assign new_n8761_ = ng826 & new_n6737_;
  assign new_n8762_ = ~ng1819 & ~ng826;
  assign n1523 = ~new_n8761_ & ~new_n8762_;
  assign new_n8764_ = ~ng2384 & new_n6572_;
  assign new_n8765_ = ~new_n6572_ & ~new_n6758_;
  assign new_n8766_ = ~new_n8764_ & ~new_n8765_;
  assign new_n8767_ = ng826 & new_n8766_;
  assign new_n8768_ = ~ng1703 & ~new_n8767_;
  assign new_n8769_ = ~new_n6299_1_ & new_n6571_;
  assign new_n8770_ = new_n6289_1_ & new_n8769_;
  assign new_n8771_ = new_n6299_1_ & new_n6561_;
  assign new_n8772_ = ~new_n8770_ & ~new_n8771_;
  assign new_n8773_ = ~new_n6294_1_ & ~new_n8772_;
  assign new_n8774_ = new_n8767_ & new_n8773_;
  assign n1528 = ~new_n8768_ & ~new_n8774_;
  assign new_n8776_ = ng823 & ~new_n6634_;
  assign new_n8777_ = ~ng1839 & ~ng823;
  assign n1547 = ~new_n8776_ & ~new_n8777_;
  assign new_n8779_ = ng1315 & n2736;
  assign new_n8780_ = ~ng1958 & ~new_n8779_;
  assign new_n8781_ = ~new_n6824_ & new_n8779_;
  assign n1556 = ~new_n8780_ & ~new_n8781_;
  assign new_n8783_ = ~new_n5366_ & ~new_n6983_;
  assign new_n8784_ = ng1312 & ~new_n8783_;
  assign new_n8785_ = ~ng1979 & ~ng1312;
  assign n1561 = ~new_n8784_ & ~new_n8785_;
  assign new_n8787_ = ng1312 & ~new_n8100_;
  assign new_n8788_ = ~ng1874 & ~ng1312;
  assign n1566 = ~new_n8787_ & ~new_n8788_;
  assign new_n8790_ = ng2020 & ~new_n6994_;
  assign new_n8791_ = ~ng2020 & new_n6994_;
  assign new_n8792_ = ~new_n8790_ & ~new_n8791_;
  assign n1576 = ~new_n6993_ & ~new_n8792_;
  assign new_n8794_ = ~ng2080 & ~new_n7011_;
  assign new_n8795_ = ng2020 & new_n7011_;
  assign n1581 = ~new_n8794_ & ~new_n8795_;
  assign new_n8797_ = ~ng2113 & ~new_n6993_;
  assign new_n8798_ = ~new_n6785_ & new_n6993_;
  assign n1586 = ~new_n8797_ & ~new_n8798_;
  assign new_n8800_ = ~ng2209 & ~new_n5517_1_;
  assign new_n8801_ = ng2170 & new_n5517_1_;
  assign n1591 = ~new_n8800_ & ~new_n8801_;
  assign new_n8803_ = ~ng2239 & ~new_n5517_1_;
  assign new_n8804_ = new_n5517_1_ & ~new_n7136_1_;
  assign n1596 = ~new_n8803_ & ~new_n8804_;
  assign new_n8806_ = ~ng2250 & ~new_n8121_;
  assign new_n8807_ = ng2165 & new_n8121_;
  assign n1601 = ~new_n8806_ & ~new_n8807_;
  assign new_n8809_ = ng826 & ~new_n7336_;
  assign new_n8810_ = ~ng2306 & ~ng826;
  assign n1606 = ~new_n8809_ & ~new_n8810_;
  assign new_n8812_ = ng2185 & ~new_n7323_;
  assign new_n8813_ = ~new_n7322_ & ~new_n8812_;
  assign new_n8814_ = ~new_n7077_ & ~new_n7356_;
  assign new_n8815_ = new_n7077_ & new_n7356_;
  assign new_n8816_ = ~new_n8814_ & ~new_n8815_;
  assign new_n8817_ = new_n7322_ & new_n8816_;
  assign new_n8818_ = ~new_n8813_ & ~new_n8817_;
  assign new_n8819_ = ng853 & ~new_n8818_;
  assign new_n8820_ = ~ng2285 & ~ng853;
  assign n1611 = ~new_n8819_ & ~new_n8820_;
  assign new_n8822_ = ng853 & ~new_n7391_;
  assign new_n8823_ = ~ng2348 & ~ng853;
  assign n1616 = ~new_n8822_ & ~new_n8823_;
  assign new_n8825_ = ~ng2444 & ~new_n8146_;
  assign new_n8826_ = ~new_n7433_ & new_n8146_;
  assign n1626 = ~new_n8825_ & ~new_n8826_;
  assign new_n8828_ = ~new_n7454_ & new_n7459_;
  assign new_n8829_ = n2815 & new_n8828_;
  assign new_n8830_ = ~new_n7311_ & new_n7454_;
  assign new_n8831_ = new_n7459_ & new_n8830_;
  assign new_n8832_ = ~n2815 & new_n8831_;
  assign new_n8833_ = ~new_n8829_ & ~new_n8832_;
  assign new_n8834_ = ~new_n7445_ & new_n8833_;
  assign new_n8835_ = n2815 & new_n7454_;
  assign new_n8836_ = ~n2815 & ~new_n8830_;
  assign new_n8837_ = ~new_n8835_ & ~new_n8836_;
  assign new_n8838_ = new_n7445_ & new_n8837_;
  assign new_n8839_ = ~new_n8834_ & ~new_n8838_;
  assign new_n8840_ = ng2384 & ~new_n8839_;
  assign new_n8841_ = ~new_n7445_ & new_n8840_;
  assign new_n8842_ = ~new_n7445_ & ~new_n8841_;
  assign new_n8843_ = new_n8840_ & ~new_n8841_;
  assign new_n8844_ = ~new_n8842_ & ~new_n8843_;
  assign new_n8845_ = ng853 & new_n8844_;
  assign new_n8846_ = ~ng2489 & ~ng853;
  assign n1631 = ~new_n8845_ & ~new_n8846_;
  assign new_n8848_ = ng853 & ~new_n8200_;
  assign new_n8849_ = ~ng2395 & ~ng853;
  assign n1636 = ~new_n8848_ & ~new_n8849_;
  assign new_n8851_ = ng1312 & ng2645;
  assign new_n8852_ = ng1315 & ng2647;
  assign new_n8853_ = ng1309 & ng2643;
  assign new_n8854_ = ~new_n8851_ & ~new_n8852_;
  assign n1651 = ~new_n8853_ & new_n8854_;
  assign new_n8856_ = ng826 & ~new_n7408_;
  assign new_n8857_ = ~ng2530 & ~ng826;
  assign n1661 = ~new_n8856_ & ~new_n8857_;
  assign new_n8859_ = ng1315 & ~ng2553;
  assign new_n8860_ = ng1309 & ~ng2554;
  assign new_n8861_ = ng1312 & ~ng2552;
  assign new_n8862_ = ~new_n8859_ & ~new_n8860_;
  assign n1666 = ~new_n8861_ & new_n8862_;
  assign new_n8864_ = ~ng2654 & ~new_n8209_;
  assign new_n8865_ = new_n7561_ & ~new_n7569_;
  assign new_n8866_ = ~pg3229 & new_n8865_;
  assign new_n8867_ = ~new_n7561_ & ~new_n7569_;
  assign new_n8868_ = pg3229 & new_n8867_;
  assign new_n8869_ = ~new_n8866_ & ~new_n8868_;
  assign new_n8870_ = ~new_n7574_ & new_n8869_;
  assign new_n8871_ = new_n8209_ & ~new_n8870_;
  assign n1671 = ~new_n8864_ & ~new_n8871_;
  assign new_n8873_ = ng2727 & new_n8216_;
  assign new_n8874_ = ~ng2720 & new_n8873_;
  assign new_n8875_ = ng2720 & ~new_n8873_;
  assign new_n8876_ = ~new_n8874_ & ~new_n8875_;
  assign n1676 = ~new_n8213_ & ~new_n8876_;
  assign new_n8878_ = ~ng2777 & ~new_n7588_;
  assign new_n8879_ = ng2707 & new_n7588_;
  assign n1681 = ~new_n8878_ & ~new_n8879_;
  assign new_n8881_ = ~ng2795 & ~new_n7588_;
  assign new_n8882_ = ng2753 & new_n7588_;
  assign n1686 = ~new_n8881_ & ~new_n8882_;
  assign new_n8884_ = ~ng2810 & ~new_n7588_;
  assign new_n8885_ = new_n7588_ & ~new_n8338_;
  assign n1691 = ~new_n8884_ & ~new_n8885_;
  assign new_n8887_ = ~ng532 & new_n7609_;
  assign new_n8888_ = ~new_n7605_ & new_n8887_;
  assign new_n8889_ = ~new_n5413_1_ & ~new_n7627_;
  assign new_n8890_ = ~new_n5302_1_ & ~new_n8889_;
  assign new_n8891_ = ~new_n8889_ & ~new_n8890_;
  assign new_n8892_ = ~new_n5302_1_ & ~new_n8890_;
  assign new_n8893_ = ~new_n8891_ & ~new_n8892_;
  assign new_n8894_ = new_n7609_ & ~new_n8893_;
  assign new_n8895_ = ng499 & new_n8894_;
  assign new_n8896_ = new_n7605_ & new_n8895_;
  assign new_n8897_ = ~new_n8888_ & ~new_n8896_;
  assign new_n8898_ = ~new_n7603_ & new_n8897_;
  assign n1696 = new_n8355_ | new_n8898_;
  assign new_n8900_ = ng1309 & ~n1448;
  assign new_n8901_ = ~ng3100 & ~ng1309;
  assign n1701 = ~new_n8900_ & ~new_n8901_;
  assign new_n8903_ = ~ng3155 & ~ng1309;
  assign n1706 = ~new_n7606_ & ~new_n8903_;
  assign new_n8905_ = ng1309 & ~ng2574;
  assign new_n8906_ = ~ng3182 & ~ng1309;
  assign n1711 = ~new_n8905_ & ~new_n8906_;
  assign new_n8908_ = ~ng162 & ~new_n4773_;
  assign new_n8909_ = new_n4773_ & ~new_n4891_;
  assign n1721 = ~new_n8908_ & ~new_n8909_;
  assign new_n8911_ = ~ng174 & ~new_n8121_;
  assign new_n8912_ = ng97 & new_n8121_;
  assign n1726 = ~new_n8911_ & ~new_n8912_;
  assign new_n8914_ = ~new_n4932_1_ & ~new_n5083_;
  assign new_n8915_ = ~new_n4797_1_ & new_n5083_;
  assign new_n8916_ = ~new_n8914_ & ~new_n8915_;
  assign new_n8917_ = ~new_n5082_1_ & new_n8916_;
  assign new_n8918_ = new_n4797_1_ & ~new_n4827_1_;
  assign new_n8919_ = ~new_n4797_1_ & new_n4827_1_;
  assign new_n8920_ = ~new_n8918_ & ~new_n8919_;
  assign new_n8921_ = ~new_n5088_ & ~new_n8920_;
  assign new_n8922_ = new_n5096_ & new_n5110_;
  assign new_n8923_ = new_n5103_ & new_n8921_;
  assign new_n8924_ = new_n8922_ & new_n8923_;
  assign new_n8925_ = ~new_n4856_ & ~new_n8924_;
  assign new_n8926_ = new_n4856_ & new_n8924_;
  assign new_n8927_ = ~new_n8925_ & ~new_n8926_;
  assign new_n8928_ = new_n5082_1_ & new_n8927_;
  assign new_n8929_ = ~new_n8917_ & ~new_n8928_;
  assign new_n8930_ = ng826 & ~new_n8929_;
  assign new_n8931_ = ~ng222 & ~ng826;
  assign n1731 = ~new_n8930_ & ~new_n8931_;
  assign new_n8933_ = ng79 & ~new_n8375_;
  assign new_n8934_ = ~ng79 & new_n8375_;
  assign new_n8935_ = ~new_n8933_ & ~new_n8934_;
  assign n1736 = ~new_n5127_1_ & ~new_n8935_;
  assign new_n8937_ = ng853 & new_n5137_1_;
  assign new_n8938_ = ~ng346 & ~new_n8937_;
  assign new_n8939_ = ~new_n8398_ & new_n8937_;
  assign n1741 = ~new_n8938_ & ~new_n8939_;
  assign new_n8941_ = ~ng391 & ~new_n8937_;
  assign new_n8942_ = new_n5144_ & new_n5158_;
  assign new_n8943_ = ~pg3229 & ~new_n5149_;
  assign new_n8944_ = new_n8942_ & new_n8943_;
  assign new_n8945_ = pg3229 & new_n5149_;
  assign new_n8946_ = new_n8942_ & new_n8945_;
  assign new_n8947_ = ~new_n8944_ & ~new_n8946_;
  assign new_n8948_ = new_n8937_ & ~new_n8947_;
  assign n1746 = ~new_n8941_ & ~new_n8948_;
  assign new_n8950_ = ng823 & ~new_n5273_;
  assign new_n8951_ = ~ng319 & ~ng823;
  assign n1751 = ~new_n8950_ & ~new_n8951_;
  assign new_n8953_ = ~ng557 & ng1315;
  assign new_n8954_ = ~ng1315 & ~ng510;
  assign n1768 = ~new_n8953_ & ~new_n8954_;
  assign new_n8956_ = ng853 & new_n5212_1_;
  assign new_n8957_ = ~ng488 & ~ng853;
  assign n1777 = ~new_n8956_ & ~new_n8957_;
  assign new_n8959_ = ng1309 & n3888;
  assign new_n8960_ = ~ng579 & ~new_n8959_;
  assign new_n8961_ = ~new_n8431_ & new_n8959_;
  assign n1786 = ~new_n8960_ & ~new_n8961_;
  assign new_n8963_ = ng1309 & ~new_n5367_;
  assign new_n8964_ = ~ng587 & ~ng1309;
  assign n1791 = ~new_n8963_ & ~new_n8964_;
  assign new_n8966_ = ng1309 & ~new_n7861_;
  assign new_n8967_ = ~ng605 & ~ng1309;
  assign n1796 = ~new_n8966_ & ~new_n8967_;
  assign new_n8969_ = ng672 & new_n8445_;
  assign new_n8970_ = ng666 & ~new_n8969_;
  assign new_n8971_ = ~ng666 & new_n8969_;
  assign new_n8972_ = ~new_n8970_ & ~new_n8971_;
  assign n1801 = ~new_n5380_ & ~new_n8972_;
  assign new_n8974_ = ~ng701 & ~new_n5399_;
  assign new_n8975_ = ng633 & new_n5399_;
  assign n1806 = ~new_n8974_ & ~new_n8975_;
  assign new_n8977_ = ~ng710 & ~new_n5399_;
  assign new_n8978_ = ng660 & new_n5399_;
  assign n1811 = ~new_n8977_ & ~new_n8978_;
  assign new_n8980_ = ~ng719 & ~new_n5399_;
  assign new_n8981_ = ng679 & new_n5399_;
  assign n1816 = ~new_n8980_ & ~new_n8981_;
  assign new_n8983_ = ng1312 & ~new_n8459_;
  assign new_n8984_ = ~ng739 & ~new_n8983_;
  assign new_n8985_ = ng630 & new_n8983_;
  assign n1821 = ~new_n8984_ & ~new_n8985_;
  assign new_n8987_ = ~ng822 & ~new_n4777_1_;
  assign new_n8988_ = ng789 & new_n4777_1_;
  assign n1826 = ~new_n8987_ & ~new_n8988_;
  assign new_n8990_ = ~ng837 & ~new_n4777_1_;
  assign new_n8991_ = ng801 & new_n4777_1_;
  assign n1831 = ~new_n8990_ & ~new_n8991_;
  assign new_n8993_ = ~ng846 & ~new_n4777_1_;
  assign new_n8994_ = ng813 & new_n4777_1_;
  assign n1836 = ~new_n8993_ & ~new_n8994_;
  assign new_n8996_ = ng853 & ~new_n7901_;
  assign new_n8997_ = ~ng888 & ~ng853;
  assign n1841 = ~new_n8996_ & ~new_n8997_;
  assign new_n8999_ = ng853 & ~new_n5878_1_;
  assign new_n9000_ = ~ng942 & ~ng853;
  assign n1846 = ~new_n8999_ & ~new_n9000_;
  assign new_n9002_ = ng853 & ~new_n8494_;
  assign new_n9003_ = ~ng915 & ~ng853;
  assign n1851 = ~new_n9002_ & ~new_n9003_;
  assign new_n9005_ = ng758 & ~new_n5915_;
  assign new_n9006_ = ~ng758 & new_n5915_;
  assign new_n9007_ = ~new_n9005_ & ~new_n9006_;
  assign n1856 = ~new_n5127_1_ & ~new_n9007_;
  assign new_n9009_ = new_n5955_ & ~new_n5969_;
  assign new_n9010_ = n953 & new_n9009_;
  assign new_n9011_ = new_n5955_ & new_n5971_;
  assign new_n9012_ = ~n953 & new_n9011_;
  assign new_n9013_ = ~new_n9010_ & ~new_n9012_;
  assign new_n9014_ = ~new_n5978_ & new_n9013_;
  assign new_n9015_ = n953 & new_n5969_;
  assign new_n9016_ = ~n953 & ~new_n5971_;
  assign new_n9017_ = ~new_n9015_ & ~new_n9016_;
  assign new_n9018_ = new_n5978_ & new_n9017_;
  assign new_n9019_ = ~new_n9014_ & ~new_n9018_;
  assign new_n9020_ = ng2384 & ~new_n9019_;
  assign new_n9021_ = ~new_n5978_ & new_n9020_;
  assign new_n9022_ = ~new_n5978_ & ~new_n9021_;
  assign new_n9023_ = new_n9020_ & ~new_n9021_;
  assign new_n9024_ = ~new_n9022_ & ~new_n9023_;
  assign new_n9025_ = ng826 & new_n9024_;
  assign new_n9026_ = ~ng1095 & ~ng826;
  assign n1861 = ~new_n9025_ & ~new_n9026_;
  assign new_n9028_ = ng826 & ~new_n8525_;
  assign new_n9029_ = ~ng1116 & ~ng826;
  assign n1866 = ~new_n9028_ & ~new_n9029_;
  assign new_n9031_ = ng826 & ~new_n5999_;
  assign new_n9032_ = ~ng999 & ~ng826;
  assign n1871 = ~new_n9031_ & ~new_n9032_;
  assign new_n9034_ = ng826 & new_n7937_;
  assign new_n9035_ = ~ng1009 & ~new_n9034_;
  assign new_n9036_ = new_n7944_ & new_n9034_;
  assign n1876 = ~new_n9035_ & ~new_n9036_;
  assign new_n9038_ = ng826 & ~new_n5924_;
  assign new_n9039_ = ~ng1142 & ~ng826;
  assign n1894 = ~new_n9038_ & ~new_n9039_;
  assign new_n9041_ = ng826 & ~new_n5560_;
  assign new_n9042_ = ~ng1152 & ~ng826;
  assign n1899 = ~new_n9041_ & ~new_n9042_;
  assign new_n9044_ = ~ng1171 & ng1315;
  assign new_n9045_ = ~ng1151 & ng1309;
  assign new_n9046_ = ng1312 & ~ng1167;
  assign new_n9047_ = ~new_n9044_ & ~new_n9045_;
  assign n1904 = ~new_n9046_ & new_n9047_;
  assign new_n9049_ = ~ng1264 & ~new_n6049_;
  assign new_n9050_ = new_n6055_ & ~new_n6097_1_;
  assign new_n9051_ = ~pg3229 & new_n9050_;
  assign new_n9052_ = ~new_n6055_ & ~new_n6097_1_;
  assign new_n9053_ = pg3229 & new_n9052_;
  assign new_n9054_ = ~new_n6065_ & new_n6097_1_;
  assign new_n9055_ = ~new_n9051_ & ~new_n9053_;
  assign new_n9056_ = ~new_n9054_ & new_n9055_;
  assign new_n9057_ = new_n6049_ & ~new_n9056_;
  assign n1908 = ~new_n9049_ & ~new_n9057_;
  assign new_n9059_ = ~ng1406 & ~new_n6259_1_;
  assign new_n9060_ = ng1365 & new_n6259_1_;
  assign n1927 = ~new_n9059_ & ~new_n9060_;
  assign new_n9062_ = ng1309 & ng1316;
  assign new_n9063_ = ~ng1415 & ~new_n9062_;
  assign new_n9064_ = ~new_n6044_ & new_n9062_;
  assign n1932 = ~new_n9063_ & ~new_n9064_;
  assign new_n9066_ = ng1309 & ~new_n6267_;
  assign new_n9067_ = ~ng1424 & ~new_n9066_;
  assign new_n9068_ = ng1316 & new_n9066_;
  assign n1937 = ~new_n9067_ & ~new_n9068_;
  assign new_n9070_ = ~ng1524 & ~new_n5517_1_;
  assign new_n9071_ = ng1481 & new_n5517_1_;
  assign n1942 = ~new_n9070_ & ~new_n9071_;
  assign new_n9073_ = ~ng1538 & ~new_n4773_;
  assign new_n9074_ = ng1506 & new_n4773_;
  assign n1947 = ~new_n9073_ & ~new_n9074_;
  assign new_n9076_ = ~ng1550 & ~new_n8121_;
  assign new_n9077_ = ~new_n6282_ & new_n8121_;
  assign n1952 = ~new_n9076_ & ~new_n9077_;
  assign new_n9079_ = ~ng1555 & ~new_n6278_;
  assign new_n9080_ = ng1476 & new_n6278_;
  assign n1957 = ~new_n9079_ & ~new_n9080_;
  assign new_n9082_ = ng1444 & new_n8716_;
  assign new_n9083_ = ~ng1439 & new_n9082_;
  assign new_n9084_ = ng1439 & ~new_n9082_;
  assign new_n9085_ = ~new_n9083_ & ~new_n9084_;
  assign n1962 = ~new_n5127_1_ & ~new_n9085_;
  assign new_n9087_ = ng853 & new_n6635_;
  assign new_n9088_ = ~ng1742 & ~new_n9087_;
  assign new_n9089_ = ~new_n6659_ & new_n9087_;
  assign n1967 = ~new_n9088_ & ~new_n9089_;
  assign new_n9091_ = ng853 & new_n8757_;
  assign new_n9092_ = ~ng1795 & ~ng853;
  assign n1972 = ~new_n9091_ & ~new_n9092_;
  assign new_n9094_ = ~new_n6720_1_ & new_n6726_;
  assign new_n9095_ = new_n6726_ & ~new_n9094_;
  assign new_n9096_ = ~new_n6720_1_ & ~new_n9094_;
  assign new_n9097_ = ~new_n9095_ & ~new_n9096_;
  assign new_n9098_ = ng2384 & ~new_n9097_;
  assign new_n9099_ = ~new_n6720_1_ & ~new_n9098_;
  assign new_n9100_ = ~new_n6720_1_ & ~new_n9099_;
  assign new_n9101_ = ~new_n9098_ & ~new_n9099_;
  assign new_n9102_ = ~new_n9100_ & ~new_n9101_;
  assign new_n9103_ = ng853 & ~new_n9102_;
  assign new_n9104_ = ~ng1816 & ~ng853;
  assign n1977 = ~new_n9103_ & ~new_n9104_;
  assign new_n9106_ = ng823 & new_n8766_;
  assign new_n9107_ = ~ng1704 & ~new_n9106_;
  assign new_n9108_ = new_n8773_ & new_n9106_;
  assign n1982 = ~new_n9107_ & ~new_n9108_;
  assign new_n9110_ = ng853 & ~new_n6634_;
  assign new_n9111_ = ~ng1842 & ~ng853;
  assign n1999 = ~new_n9110_ & ~new_n9111_;
  assign new_n9113_ = ng853 & ~new_n6303_;
  assign new_n9114_ = ~ng1852 & ~ng853;
  assign n2004 = ~new_n9113_ & ~new_n9114_;
  assign new_n9116_ = ~ng1962 & ~new_n6801_;
  assign new_n9117_ = pg3229 & ~new_n6812_;
  assign new_n9118_ = new_n6892_1_ & new_n9117_;
  assign new_n9119_ = ~pg3229 & new_n6812_;
  assign new_n9120_ = new_n6892_1_ & new_n9119_;
  assign new_n9121_ = ~new_n9118_ & ~new_n9120_;
  assign new_n9122_ = ~new_n6812_ & ~new_n6821_;
  assign new_n9123_ = ~pg3229 & new_n9122_;
  assign new_n9124_ = new_n6812_ & ~new_n6821_;
  assign new_n9125_ = pg3229 & new_n9124_;
  assign new_n9126_ = ~new_n9123_ & ~new_n9125_;
  assign new_n9127_ = new_n9121_ & new_n9126_;
  assign new_n9128_ = new_n6801_ & ~new_n9127_;
  assign n2009 = ~new_n9116_ & ~new_n9128_;
  assign new_n9130_ = ng1309 & ~new_n8783_;
  assign new_n9131_ = ~ng1976 & ~ng1309;
  assign n2014 = ~new_n9130_ & ~new_n9131_;
  assign new_n9133_ = ng1315 & ~new_n8100_;
  assign new_n9134_ = ~ng1315 & ~ng1877;
  assign n2019 = ~new_n9133_ & ~new_n9134_;
  assign new_n9136_ = ~ng2013 & new_n6995_1_;
  assign new_n9137_ = ng2013 & ~new_n6995_1_;
  assign new_n9138_ = ~new_n9136_ & ~new_n9137_;
  assign n2029 = ~new_n6993_ & ~new_n9138_;
  assign new_n9140_ = ~ng2079 & ~new_n7003_;
  assign new_n9141_ = ng2020 & new_n7003_;
  assign n2034 = ~new_n9140_ & ~new_n9141_;
  assign new_n9143_ = ng1315 & ng2010;
  assign new_n9144_ = ~ng2111 & ~new_n9143_;
  assign new_n9145_ = ~new_n6785_ & new_n9143_;
  assign n2039 = ~new_n9144_ & ~new_n9145_;
  assign new_n9147_ = ~ng2205 & ~new_n4773_;
  assign new_n9148_ = ng2165 & new_n4773_;
  assign n2044 = ~new_n9147_ & ~new_n9148_;
  assign new_n9150_ = ~ng2240 & ~new_n4777_1_;
  assign new_n9151_ = new_n4777_1_ & ~new_n7136_1_;
  assign n2049 = ~new_n9150_ & ~new_n9151_;
  assign new_n9153_ = ~ng2252 & ~new_n6278_;
  assign new_n9154_ = ng2165 & new_n6278_;
  assign n2054 = ~new_n9153_ & ~new_n9154_;
  assign new_n9156_ = ng823 & ~new_n7336_;
  assign new_n9157_ = ~ng2309 & ~ng823;
  assign n2059 = ~new_n9156_ & ~new_n9157_;
  assign new_n9159_ = ng823 & ~new_n8818_;
  assign new_n9160_ = ~ng2282 & ~ng823;
  assign n2064 = ~new_n9159_ & ~new_n9160_;
  assign new_n9162_ = ~ng2160 & new_n5128_;
  assign new_n9163_ = ng2160 & ~new_n5128_;
  assign new_n9164_ = ~new_n9162_ & ~new_n9163_;
  assign n2069 = ~new_n5127_1_ & ~new_n9164_;
  assign new_n9166_ = ng2124 & new_n7402_;
  assign new_n9167_ = ng2120 & ~new_n9166_;
  assign new_n9168_ = ~ng2120 & new_n9166_;
  assign new_n9169_ = ~new_n9167_ & ~new_n9168_;
  assign n2074 = ~new_n5127_1_ & ~new_n9169_;
  assign new_n9171_ = ng823 & new_n7409_;
  assign new_n9172_ = ~ng2433 & ~new_n9171_;
  assign new_n9173_ = ~new_n7433_ & new_n9171_;
  assign n2079 = ~new_n9172_ & ~new_n9173_;
  assign new_n9175_ = ng823 & new_n8844_;
  assign new_n9176_ = ~ng2486 & ~ng823;
  assign n2084 = ~new_n9175_ & ~new_n9176_;
  assign new_n9178_ = ~ng2384 & new_n7308_;
  assign new_n9179_ = ~new_n7308_ & ~new_n8187_;
  assign new_n9180_ = ~new_n9178_ & ~new_n9179_;
  assign new_n9181_ = ng826 & new_n9180_;
  assign new_n9182_ = ~ng2397 & ~new_n9181_;
  assign new_n9183_ = ~new_n7040_ & new_n7307_;
  assign new_n9184_ = new_n7030_ & new_n9183_;
  assign new_n9185_ = new_n7040_ & new_n7297_;
  assign new_n9186_ = ~new_n9184_ & ~new_n9185_;
  assign new_n9187_ = ~new_n7035_ & ~new_n9186_;
  assign new_n9188_ = new_n9181_ & new_n9187_;
  assign n2089 = ~new_n9182_ & ~new_n9188_;
  assign new_n9190_ = ~ng2631 & ng1315;
  assign new_n9191_ = ~ng1315 & ~ng2584;
  assign n2103 = ~new_n9190_ & ~new_n9191_;
  assign new_n9193_ = ng853 & new_n7489_;
  assign new_n9194_ = ~ng2563 & ~ng853;
  assign n2112 = ~new_n9193_ & ~new_n9194_;
  assign new_n9196_ = ng1309 & n4397;
  assign new_n9197_ = ~ng2653 & ~new_n9196_;
  assign new_n9198_ = ~new_n8870_ & new_n9196_;
  assign n2121 = ~new_n9197_ & ~new_n9198_;
  assign new_n9200_ = ng2720 & new_n8873_;
  assign new_n9201_ = ng2734 & ~new_n9200_;
  assign new_n9202_ = ~ng2734 & new_n9200_;
  assign new_n9203_ = ~new_n9201_ & ~new_n9202_;
  assign n2126 = ~new_n8213_ & ~new_n9203_;
  assign new_n9205_ = ~ng2776 & ~new_n7592_;
  assign new_n9206_ = ng2707 & new_n7592_;
  assign n2131 = ~new_n9205_ & ~new_n9206_;
  assign new_n9208_ = ~ng2785 & ~new_n7592_;
  assign new_n9209_ = ng2734 & new_n7592_;
  assign n2136 = ~new_n9208_ & ~new_n9209_;
  assign new_n9211_ = ~ng2808 & ~new_n7584_;
  assign new_n9212_ = new_n7584_ & ~new_n8338_;
  assign n2141 = ~new_n9211_ & ~new_n9212_;
  assign new_n9214_ = ~ng531 & new_n7609_;
  assign new_n9215_ = ~new_n7605_ & new_n9214_;
  assign new_n9216_ = ~new_n5489_ & ~new_n7627_;
  assign new_n9217_ = ~new_n5287_1_ & ~new_n9216_;
  assign new_n9218_ = ~new_n9216_ & ~new_n9217_;
  assign new_n9219_ = ~new_n5287_1_ & ~new_n9217_;
  assign new_n9220_ = ~new_n9218_ & ~new_n9219_;
  assign new_n9221_ = new_n7609_ & ~new_n9220_;
  assign new_n9222_ = ng499 & new_n9221_;
  assign new_n9223_ = new_n7605_ & new_n9222_;
  assign new_n9224_ = ~new_n9215_ & ~new_n9223_;
  assign new_n9225_ = ~new_n7603_ & new_n9224_;
  assign n2146 = new_n7648_ | new_n9225_;
  assign new_n9227_ = ng2903 & ng2908;
  assign new_n9228_ = ~ng2900 & new_n9227_;
  assign new_n9229_ = ng2892 & new_n9228_;
  assign new_n9230_ = ~ng2896 & ~ng2883;
  assign new_n9231_ = ng2888 & new_n9230_;
  assign new_n9232_ = ng2950 & new_n9231_;
  assign new_n9233_ = new_n9229_ & new_n9232_;
  assign new_n9234_ = ~ng2814 & ~new_n9233_;
  assign new_n9235_ = ng2950 & ng2883;
  assign new_n9236_ = ng2888 & new_n9235_;
  assign new_n9237_ = ng2896 & new_n9236_;
  assign new_n9238_ = ng2892 & new_n9237_;
  assign new_n9239_ = ng2903 & new_n9238_;
  assign new_n9240_ = ng2900 & ~new_n9239_;
  assign new_n9241_ = ~ng2900 & new_n9239_;
  assign new_n9242_ = ~new_n9240_ & ~new_n9241_;
  assign n2151 = new_n9234_ & ~new_n9242_;
  assign new_n9244_ = ng1315 & ~ng1939;
  assign new_n9245_ = ~ng1315 & ~ng3093;
  assign n2156 = ~new_n9244_ & ~new_n9245_;
  assign new_n9247_ = ng1312 & ~n2721;
  assign new_n9248_ = ~ng1312 & ~ng3104;
  assign n2161 = ~new_n9247_ & ~new_n9248_;
  assign new_n9250_ = ng1309 & ~ng1880;
  assign new_n9251_ = ~ng3173 & ~ng1309;
  assign n2166 = ~new_n9250_ & ~new_n9251_;
  assign new_n9253_ = ng105 & ~new_n5083_;
  assign new_n9254_ = ~new_n8915_ & ~new_n9253_;
  assign new_n9255_ = ~new_n5082_1_ & new_n9254_;
  assign new_n9256_ = ~new_n4805_ & ~new_n5096_;
  assign new_n9257_ = new_n4805_ & new_n5096_;
  assign new_n9258_ = ~new_n9256_ & ~new_n9257_;
  assign new_n9259_ = new_n5082_1_ & new_n9258_;
  assign new_n9260_ = ~new_n9255_ & ~new_n9259_;
  assign new_n9261_ = ng826 & ~new_n9260_;
  assign new_n9262_ = ~ng195 & ~ng826;
  assign n2176 = ~new_n9261_ & ~new_n9262_;
  assign new_n9264_ = ng117 & ~new_n5083_;
  assign new_n9265_ = ~new_n5082_1_ & ~new_n9264_;
  assign new_n9266_ = ~new_n5109_ & new_n5111_;
  assign new_n9267_ = new_n4837_1_ & new_n9266_;
  assign new_n9268_ = ~new_n4837_1_ & ~new_n9266_;
  assign new_n9269_ = ~new_n9267_ & ~new_n9268_;
  assign new_n9270_ = new_n5082_1_ & new_n9269_;
  assign new_n9271_ = ~new_n9265_ & ~new_n9270_;
  assign new_n9272_ = ng853 & ~new_n9271_;
  assign new_n9273_ = ~ng255 & ~ng853;
  assign n2181 = ~new_n9272_ & ~new_n9273_;
  assign new_n9275_ = ~new_n4891_ & ~new_n5083_;
  assign new_n9276_ = ~new_n8915_ & ~new_n9275_;
  assign new_n9277_ = ~new_n5082_1_ & new_n9276_;
  assign new_n9278_ = new_n4797_1_ & ~new_n4856_;
  assign new_n9279_ = ~new_n4797_1_ & new_n4856_;
  assign new_n9280_ = ~new_n9278_ & ~new_n9279_;
  assign new_n9281_ = new_n8924_ & ~new_n9280_;
  assign new_n9282_ = new_n4822_1_ & new_n9281_;
  assign new_n9283_ = ~new_n4822_1_ & ~new_n9281_;
  assign new_n9284_ = ~new_n9282_ & ~new_n9283_;
  assign new_n9285_ = new_n5082_1_ & new_n9284_;
  assign new_n9286_ = ~new_n9277_ & ~new_n9285_;
  assign new_n9287_ = ng823 & ~new_n9286_;
  assign new_n9288_ = ~ng270 & ~ng823;
  assign n2186 = ~new_n9287_ & ~new_n9288_;
  assign new_n9290_ = ng74 & new_n8376_;
  assign new_n9291_ = ng70 & new_n9290_;
  assign new_n9292_ = ng65 & new_n9291_;
  assign new_n9293_ = ng61 & new_n9292_;
  assign new_n9294_ = ng56 & new_n9293_;
  assign new_n9295_ = ng52 & ~new_n9294_;
  assign new_n9296_ = ~ng52 & new_n9294_;
  assign new_n9297_ = ~new_n9295_ & ~new_n9296_;
  assign n2191 = ~new_n5127_1_ & ~new_n9297_;
  assign new_n9299_ = ~ng388 & ~new_n7672_;
  assign new_n9300_ = new_n7672_ & ~new_n8947_;
  assign n2196 = ~new_n9299_ & ~new_n9300_;
  assign new_n9302_ = ng52 & new_n4822_1_;
  assign new_n9303_ = new_n4822_1_ & ~new_n9302_;
  assign new_n9304_ = ng52 & ~new_n9302_;
  assign new_n9305_ = ~new_n9303_ & ~new_n9304_;
  assign new_n9306_ = ng65 & new_n4849_;
  assign new_n9307_ = new_n4849_ & ~new_n9306_;
  assign new_n9308_ = ng65 & ~new_n9306_;
  assign new_n9309_ = ~new_n9307_ & ~new_n9308_;
  assign new_n9310_ = ng61 & new_n4827_1_;
  assign new_n9311_ = new_n4827_1_ & ~new_n9310_;
  assign new_n9312_ = ng61 & ~new_n9310_;
  assign new_n9313_ = ~new_n9311_ & ~new_n9312_;
  assign new_n9314_ = ng70 & new_n4837_1_;
  assign new_n9315_ = new_n4837_1_ & ~new_n9314_;
  assign new_n9316_ = ng70 & ~new_n9314_;
  assign new_n9317_ = ~new_n9315_ & ~new_n9316_;
  assign new_n9318_ = ~new_n9309_ & ~new_n9313_;
  assign new_n9319_ = ~new_n9317_ & new_n9318_;
  assign new_n9320_ = ng56 & new_n4856_;
  assign new_n9321_ = new_n4856_ & ~new_n9320_;
  assign new_n9322_ = ng56 & ~new_n9320_;
  assign new_n9323_ = ~new_n9321_ & ~new_n9322_;
  assign new_n9324_ = ~new_n9305_ & new_n9319_;
  assign new_n9325_ = ~new_n9323_ & new_n9324_;
  assign new_n9326_ = ng74 & new_n4832_1_;
  assign new_n9327_ = new_n4832_1_ & ~new_n9326_;
  assign new_n9328_ = ng74 & ~new_n9326_;
  assign new_n9329_ = ~new_n9327_ & ~new_n9328_;
  assign new_n9330_ = ng88 & new_n4815_;
  assign new_n9331_ = new_n4815_ & ~new_n9330_;
  assign new_n9332_ = ng88 & ~new_n9330_;
  assign new_n9333_ = ~new_n9331_ & ~new_n9332_;
  assign new_n9334_ = ng83 & new_n4805_;
  assign new_n9335_ = new_n4805_ & ~new_n9334_;
  assign new_n9336_ = ng83 & ~new_n9334_;
  assign new_n9337_ = ~new_n9335_ & ~new_n9336_;
  assign new_n9338_ = ng92 & new_n4842_1_;
  assign new_n9339_ = new_n4842_1_ & ~new_n9338_;
  assign new_n9340_ = ng92 & ~new_n9338_;
  assign new_n9341_ = ~new_n9339_ & ~new_n9340_;
  assign new_n9342_ = ~new_n9333_ & ~new_n9337_;
  assign new_n9343_ = ~new_n9341_ & new_n9342_;
  assign new_n9344_ = ng79 & new_n4810_;
  assign new_n9345_ = new_n4810_ & ~new_n9344_;
  assign new_n9346_ = ng79 & ~new_n9344_;
  assign new_n9347_ = ~new_n9345_ & ~new_n9346_;
  assign new_n9348_ = ~new_n9329_ & new_n9343_;
  assign new_n9349_ = ~new_n9347_ & new_n9348_;
  assign new_n9350_ = ~new_n5136_ & new_n9325_;
  assign new_n9351_ = new_n9349_ & new_n9350_;
  assign new_n9352_ = ~new_n5125_ & new_n9351_;
  assign new_n9353_ = new_n4799_ & new_n4865_;
  assign new_n9354_ = ~new_n9352_ & ~new_n9353_;
  assign n2201 = ~new_n5137_1_ | new_n9354_;
  assign new_n9356_ = ng823 & new_n5212_1_;
  assign new_n9357_ = ~ng487 & ~ng823;
  assign n2216 = ~new_n9356_ & ~new_n9357_;
  assign new_n9359_ = ng1315 & ~new_n5297_1_;
  assign new_n9360_ = ~ng1315 & ~ng659;
  assign n2226 = ~new_n9359_ & ~new_n9360_;
  assign new_n9362_ = ~ng721 & ~new_n5391_;
  assign new_n9363_ = ng679 & new_n5391_;
  assign n2231 = ~new_n9362_ & ~new_n9363_;
  assign new_n9365_ = ng1315 & ~new_n8459_;
  assign new_n9366_ = ~ng737 & ~new_n9365_;
  assign new_n9367_ = ng630 & new_n9365_;
  assign n2236 = ~new_n9366_ & ~new_n9367_;
  assign new_n9369_ = ~ng856 & ~new_n8121_;
  assign new_n9370_ = ~ng809 & ~ng805;
  assign new_n9371_ = ng813 & new_n9370_;
  assign new_n9372_ = ng801 & new_n9371_;
  assign new_n9373_ = new_n8121_ & ~new_n9372_;
  assign n2241 = ~new_n9369_ & ~new_n9373_;
  assign new_n9375_ = ng785 & ~new_n5839_;
  assign new_n9376_ = ~new_n5838_1_ & ~new_n9375_;
  assign new_n9377_ = ~new_n5561_1_ & new_n5603_;
  assign new_n9378_ = new_n5561_1_ & ~new_n5603_;
  assign new_n9379_ = ~new_n9377_ & ~new_n9378_;
  assign new_n9380_ = new_n5838_1_ & new_n9379_;
  assign new_n9381_ = ~new_n9376_ & ~new_n9380_;
  assign new_n9382_ = ng823 & ~new_n9381_;
  assign new_n9383_ = ~ng876 & ~ng823;
  assign n2246 = ~new_n9382_ & ~new_n9383_;
  assign new_n9385_ = ng823 & new_n9024_;
  assign new_n9386_ = ~ng1098 & ~ng823;
  assign n2251 = ~new_n9385_ & ~new_n9386_;
  assign new_n9388_ = ng2384 & ~new_n8533_;
  assign new_n9389_ = ~new_n8538_ & new_n9388_;
  assign new_n9390_ = ~new_n6022_1_ & new_n9389_;
  assign new_n9391_ = ~new_n6022_1_ & ~new_n9390_;
  assign new_n9392_ = new_n9389_ & ~new_n9390_;
  assign new_n9393_ = ~new_n9391_ & ~new_n9392_;
  assign new_n9394_ = ng826 & new_n9393_;
  assign new_n9395_ = ~ng1125 & ~ng826;
  assign n2256 = ~new_n9394_ & ~new_n9395_;
  assign new_n9397_ = ng823 & ~new_n5924_;
  assign new_n9398_ = ~ng1145 & ~ng823;
  assign n2271 = ~new_n9397_ & ~new_n9398_;
  assign new_n9400_ = ~ng1263 & ~new_n8012_;
  assign new_n9401_ = new_n6067_1_ & ~new_n6097_1_;
  assign new_n9402_ = ~new_n6068_ & ~new_n9401_;
  assign new_n9403_ = ~new_n6055_ & new_n6060_;
  assign new_n9404_ = ~pg3229 & new_n9403_;
  assign new_n9405_ = ~pg3229 & new_n9054_;
  assign new_n9406_ = pg3229 & ~new_n6060_;
  assign new_n9407_ = ~new_n9404_ & ~new_n9405_;
  assign new_n9408_ = ~new_n9406_ & new_n9407_;
  assign new_n9409_ = new_n9402_ & new_n9408_;
  assign new_n9410_ = new_n8012_ & ~new_n9409_;
  assign n2281 = ~new_n9400_ & ~new_n9410_;
  assign new_n9412_ = ~new_n5366_ & ~new_n6160_;
  assign new_n9413_ = ng1309 & ~new_n9412_;
  assign new_n9414_ = ~ng1282 & ~ng1309;
  assign n2286 = ~new_n9413_ & ~new_n9414_;
  assign new_n9416_ = ng1196 & new_n6044_;
  assign new_n9417_ = new_n6038_ & ~new_n9416_;
  assign new_n9418_ = ~new_n6038_ & new_n9417_;
  assign new_n9419_ = ~new_n6038_ & ~new_n9418_;
  assign new_n9420_ = new_n9417_ & ~new_n9418_;
  assign new_n9421_ = ~new_n9419_ & ~new_n9420_;
  assign new_n9422_ = ng1315 & ~new_n9421_;
  assign new_n9423_ = ~ng1315 & ~ng1183;
  assign n2291 = ~new_n9422_ & ~new_n9423_;
  assign new_n9425_ = ~ng1407 & ~new_n6255_;
  assign new_n9426_ = ng1365 & new_n6255_;
  assign n2296 = ~new_n9425_ & ~new_n9426_;
  assign new_n9428_ = ~ng1418 & ~new_n9062_;
  assign new_n9429_ = ~new_n6033_ & new_n9062_;
  assign n2301 = ~new_n9428_ & ~new_n9429_;
  assign new_n9431_ = ~ng1511 & ~new_n4773_;
  assign new_n9432_ = ng1471 & new_n4773_;
  assign n2306 = ~new_n9431_ & ~new_n9432_;
  assign new_n9434_ = ~ng1531 & ~new_n4777_1_;
  assign new_n9435_ = ng1491 & new_n4777_1_;
  assign n2311 = ~new_n9434_ & ~new_n9435_;
  assign new_n9437_ = ~ng1534 & ~new_n4777_1_;
  assign new_n9438_ = ng1496 & new_n4777_1_;
  assign n2316 = ~new_n9437_ & ~new_n9438_;
  assign new_n9440_ = ~ng1545 & ~new_n5517_1_;
  assign new_n9441_ = new_n5517_1_ & ~new_n6395_;
  assign n2321 = ~new_n9440_ & ~new_n9441_;
  assign new_n9443_ = ng1439 & new_n9082_;
  assign new_n9444_ = ng1435 & ~new_n9443_;
  assign new_n9445_ = ~ng1435 & new_n9443_;
  assign new_n9446_ = ~new_n9444_ & ~new_n9445_;
  assign n2326 = ~new_n5127_1_ & ~new_n9446_;
  assign new_n9448_ = ~ng1757 & ~new_n9087_;
  assign new_n9449_ = ~new_n8738_ & new_n9087_;
  assign n2331 = ~new_n9448_ & ~new_n9449_;
  assign new_n9451_ = n5082 & ~new_n6680_;
  assign new_n9452_ = ~n5082 & new_n8743_;
  assign new_n9453_ = ~new_n9451_ & ~new_n9452_;
  assign new_n9454_ = new_n6685_ & ~new_n9453_;
  assign new_n9455_ = ~new_n6671_1_ & new_n9454_;
  assign new_n9456_ = ng2384 & new_n9455_;
  assign new_n9457_ = new_n6671_1_ & ~new_n9453_;
  assign new_n9458_ = ng2384 & new_n9457_;
  assign new_n9459_ = ~new_n9456_ & ~new_n9458_;
  assign new_n9460_ = ng823 & ~new_n9459_;
  assign new_n9461_ = ~ng1809 & ~new_n9460_;
  assign new_n9462_ = new_n9456_ & new_n9460_;
  assign n2336 = ~new_n9461_ & ~new_n9462_;
  assign new_n9464_ = ~new_n6289_1_ & new_n6299_1_;
  assign new_n9465_ = new_n6294_1_ & new_n9464_;
  assign new_n9466_ = new_n6289_1_ & ~new_n6299_1_;
  assign new_n9467_ = ~new_n6459_ & ~new_n9466_;
  assign new_n9468_ = ~new_n6294_1_ & ~new_n9467_;
  assign new_n9469_ = ~new_n9465_ & ~new_n9468_;
  assign new_n9470_ = ~new_n6294_1_ & new_n9469_;
  assign new_n9471_ = ~new_n6294_1_ & ~new_n9470_;
  assign new_n9472_ = new_n9469_ & ~new_n9470_;
  assign new_n9473_ = ~new_n9471_ & ~new_n9472_;
  assign new_n9474_ = ~new_n6584_ & new_n9473_;
  assign new_n9475_ = ng826 & ~new_n9474_;
  assign new_n9476_ = ~ng1693 & ~ng826;
  assign n2341 = ~new_n9475_ & ~new_n9476_;
  assign new_n9478_ = new_n6289_1_ & new_n6299_1_;
  assign new_n9479_ = new_n6294_1_ & ~new_n9478_;
  assign new_n9480_ = new_n6569_ & new_n6758_;
  assign new_n9481_ = new_n6755_1_ & ~new_n9480_;
  assign new_n9482_ = ~new_n6418_ & new_n9481_;
  assign new_n9483_ = new_n6299_1_ & new_n9482_;
  assign new_n9484_ = ~new_n6573_ & ~new_n6575_1_;
  assign new_n9485_ = ~new_n6299_1_ & new_n9484_;
  assign new_n9486_ = ~new_n9483_ & ~new_n9485_;
  assign new_n9487_ = new_n6289_1_ & new_n9486_;
  assign new_n9488_ = ~new_n6418_ & new_n6758_;
  assign new_n9489_ = ~new_n6458_ & ~new_n9488_;
  assign new_n9490_ = new_n6299_1_ & new_n9489_;
  assign new_n9491_ = ~new_n6299_1_ & ~new_n6458_;
  assign new_n9492_ = ~new_n9490_ & ~new_n9491_;
  assign new_n9493_ = ~new_n6289_1_ & new_n9492_;
  assign new_n9494_ = ~new_n9487_ & ~new_n9493_;
  assign new_n9495_ = ~new_n6294_1_ & new_n9494_;
  assign new_n9496_ = ~new_n9479_ & ~new_n9495_;
  assign new_n9497_ = ~new_n6289_1_ & new_n9496_;
  assign new_n9498_ = ~new_n6289_1_ & ~new_n9497_;
  assign new_n9499_ = new_n9496_ & ~new_n9497_;
  assign new_n9500_ = ~new_n9498_ & ~new_n9499_;
  assign new_n9501_ = ~new_n6584_ & new_n9500_;
  assign new_n9502_ = ng826 & ~new_n9501_;
  assign new_n9503_ = ~ng1696 & ~ng826;
  assign n2346 = ~new_n9502_ & ~new_n9503_;
  assign new_n9505_ = ng2384 & ng853;
  assign new_n9506_ = ~ng1783 & ~new_n9505_;
  assign new_n9507_ = new_n6571_ & new_n6583_;
  assign new_n9508_ = new_n9505_ & new_n9507_;
  assign n2351 = ~new_n9506_ & ~new_n9508_;
  assign new_n9510_ = ng823 & n5082;
  assign new_n9511_ = ~ng1865 & ~ng823;
  assign n2366 = ~new_n9510_ & ~new_n9511_;
  assign new_n9513_ = ng1315 & ~ng1865;
  assign new_n9514_ = ~ng1845 & ng1309;
  assign new_n9515_ = ng1312 & ~ng1861;
  assign new_n9516_ = ~new_n9513_ & ~new_n9514_;
  assign n2371 = ~new_n9515_ & new_n9516_;
  assign new_n9518_ = ~ng1966 & ~new_n8088_;
  assign new_n9519_ = ~pg3229 & ~new_n6812_;
  assign new_n9520_ = new_n6896_ & new_n9519_;
  assign new_n9521_ = pg3229 & new_n6812_;
  assign new_n9522_ = new_n6896_ & new_n9521_;
  assign new_n9523_ = ~new_n9520_ & ~new_n9522_;
  assign new_n9524_ = new_n8088_ & ~new_n9523_;
  assign n2381 = ~new_n9518_ & ~new_n9524_;
  assign new_n9526_ = ~ng2089 & ~new_n7011_;
  assign new_n9527_ = ng2026 & new_n7011_;
  assign n2396 = ~new_n9526_ & ~new_n9527_;
  assign new_n9529_ = ~ng2100 & ~new_n7003_;
  assign new_n9530_ = ng2059 & new_n7003_;
  assign n2401 = ~new_n9529_ & ~new_n9530_;
  assign new_n9532_ = ~ng2108 & ~new_n9143_;
  assign new_n9533_ = ~new_n6796_ & new_n9143_;
  assign n2406 = ~new_n9532_ & ~new_n9533_;
  assign new_n9535_ = ~ng2207 & ~new_n4777_1_;
  assign new_n9536_ = ng2165 & new_n4777_1_;
  assign n2411 = ~new_n9535_ & ~new_n9536_;
  assign new_n9538_ = ~ng2238 & ~new_n4773_;
  assign new_n9539_ = new_n4773_ & ~new_n7136_1_;
  assign n2416 = ~new_n9538_ & ~new_n9539_;
  assign new_n9541_ = ~ng2255 & ~new_n6278_;
  assign new_n9542_ = new_n6278_ & new_n7452_;
  assign n2421 = ~new_n9541_ & ~new_n9542_;
  assign new_n9544_ = ng2180 & ~new_n7323_;
  assign new_n9545_ = ~new_n7325_ & ~new_n9544_;
  assign new_n9546_ = ~new_n7322_ & new_n9545_;
  assign new_n9547_ = new_n7348_ & ~new_n7354_;
  assign new_n9548_ = new_n7055_ & new_n9547_;
  assign new_n9549_ = ~new_n7055_ & ~new_n9547_;
  assign new_n9550_ = ~new_n9548_ & ~new_n9549_;
  assign new_n9551_ = new_n7322_ & new_n9550_;
  assign new_n9552_ = ~new_n9546_ & ~new_n9551_;
  assign new_n9553_ = ng826 & ~new_n9552_;
  assign new_n9554_ = ~ng2315 & ~ng826;
  assign n2426 = ~new_n9553_ & ~new_n9554_;
  assign new_n9556_ = ng2195 & ~new_n7323_;
  assign new_n9557_ = ~new_n7322_ & ~new_n9556_;
  assign new_n9558_ = new_n7356_ & new_n7375_1_;
  assign new_n9559_ = ~new_n7094_ & ~new_n9558_;
  assign new_n9560_ = new_n7094_ & new_n9558_;
  assign new_n9561_ = ~new_n9559_ & ~new_n9560_;
  assign new_n9562_ = new_n7322_ & new_n9561_;
  assign new_n9563_ = ~new_n9557_ & ~new_n9562_;
  assign new_n9564_ = ng853 & ~new_n9563_;
  assign new_n9565_ = ~ng2294 & ~ng853;
  assign n2431 = ~new_n9564_ & ~new_n9565_;
  assign new_n9567_ = ng2200 & ~new_n7323_;
  assign new_n9568_ = ~new_n7322_ & ~new_n9567_;
  assign new_n9569_ = ~new_n7381_ & new_n9558_;
  assign new_n9570_ = new_n7072_ & new_n9569_;
  assign new_n9571_ = ~new_n7072_ & ~new_n9569_;
  assign new_n9572_ = ~new_n9570_ & ~new_n9571_;
  assign new_n9573_ = new_n7322_ & new_n9572_;
  assign new_n9574_ = ~new_n9568_ & ~new_n9573_;
  assign new_n9575_ = ng853 & ~new_n9574_;
  assign new_n9576_ = ~ng2339 & ~ng853;
  assign n2436 = ~new_n9575_ & ~new_n9576_;
  assign new_n9578_ = ~ng2142 & new_n7398_;
  assign new_n9579_ = ng2142 & ~new_n7398_;
  assign new_n9580_ = ~new_n9578_ & ~new_n9579_;
  assign n2441 = ~new_n5127_1_ & ~new_n9580_;
  assign new_n9582_ = ~ng2418 & ~new_n9171_;
  assign new_n9583_ = ~new_n7416_1_ & new_n8154_;
  assign new_n9584_ = ~new_n8155_ & ~new_n9583_;
  assign new_n9585_ = ~new_n7421_1_ & new_n8152_;
  assign new_n9586_ = ~pg3229 & new_n9585_;
  assign new_n9587_ = ~pg3229 & new_n7431_;
  assign new_n9588_ = pg3229 & ~new_n8152_;
  assign new_n9589_ = ~new_n9586_ & ~new_n9587_;
  assign new_n9590_ = ~new_n9588_ & new_n9589_;
  assign new_n9591_ = new_n9584_ & new_n9590_;
  assign new_n9592_ = new_n9171_ & ~new_n9591_;
  assign n2446 = ~new_n9582_ & ~new_n9592_;
  assign new_n9594_ = ng826 & new_n8844_;
  assign new_n9595_ = ~ng2483 & ~ng826;
  assign n2451 = ~new_n9594_ & ~new_n9595_;
  assign new_n9597_ = ng823 & new_n9180_;
  assign new_n9598_ = ~ng2398 & ~new_n9597_;
  assign new_n9599_ = new_n9187_ & new_n9597_;
  assign n2456 = ~new_n9598_ & ~new_n9599_;
  assign new_n9601_ = ng823 & new_n7489_;
  assign new_n9602_ = ~ng2562 & ~ng823;
  assign n2481 = ~new_n9601_ & ~new_n9602_;
  assign new_n9604_ = ng1312 & ng2673;
  assign new_n9605_ = ng1315 & ng2676;
  assign new_n9606_ = ng2670 & ng1309;
  assign new_n9607_ = ~new_n9604_ & ~new_n9605_;
  assign new_n9608_ = ~new_n9606_ & new_n9607_;
  assign new_n9609_ = ng1312 & ng2641;
  assign new_n9610_ = ng1315 & ng2564;
  assign new_n9611_ = ng2639 & ng1309;
  assign new_n9612_ = ~new_n9609_ & ~new_n9610_;
  assign n6457 = ~new_n9611_ & new_n9612_;
  assign new_n9614_ = ng185 & ~n6457;
  assign new_n9615_ = ng2616 & new_n9614_;
  assign new_n9616_ = new_n9608_ & ~new_n9615_;
  assign new_n9617_ = ~new_n5366_ & ~new_n9616_;
  assign new_n9618_ = ng1309 & ~new_n9617_;
  assign new_n9619_ = ~ng2670 & ~ng1309;
  assign n2486 = ~new_n9618_ & ~new_n9619_;
  assign new_n9621_ = ng2584 & new_n7540_;
  assign new_n9622_ = new_n7534_ & ~new_n9621_;
  assign new_n9623_ = ~new_n7534_ & new_n9622_;
  assign new_n9624_ = ~new_n7534_ & ~new_n9623_;
  assign new_n9625_ = new_n9622_ & ~new_n9623_;
  assign new_n9626_ = ~new_n9624_ & ~new_n9625_;
  assign new_n9627_ = ng1315 & ~new_n9626_;
  assign new_n9628_ = ~ng1315 & ~ng2571;
  assign n2491 = ~new_n9627_ & ~new_n9628_;
  assign new_n9630_ = ~ng2704 & ~new_n7583_;
  assign new_n9631_ = ng1309 & ~new_n9630_;
  assign new_n9632_ = ~ng2812 & ~new_n9631_;
  assign new_n9633_ = ng2704 & new_n9631_;
  assign n2501 = ~new_n9632_ & ~new_n9633_;
  assign new_n9635_ = ~ng534 & new_n7609_;
  assign new_n9636_ = ~new_n7605_ & new_n9635_;
  assign new_n9637_ = ~new_n5431_1_ & ~new_n7627_;
  assign new_n9638_ = ~new_n5302_1_ & ~new_n9637_;
  assign new_n9639_ = ~new_n9637_ & ~new_n9638_;
  assign new_n9640_ = ~new_n5302_1_ & ~new_n9638_;
  assign new_n9641_ = ~new_n9639_ & ~new_n9640_;
  assign new_n9642_ = new_n7609_ & ~new_n9641_;
  assign new_n9643_ = ng499 & new_n9642_;
  assign new_n9644_ = new_n7605_ & new_n9643_;
  assign new_n9645_ = ~new_n9636_ & ~new_n9644_;
  assign new_n9646_ = ~new_n7603_ & new_n9645_;
  assign new_n9647_ = ~new_n7609_ & new_n7638_;
  assign new_n9648_ = new_n7603_ & new_n9647_;
  assign n2506 = new_n9646_ | new_n9648_;
  assign new_n9650_ = ng1309 & ~ng2633;
  assign new_n9651_ = ~ng3094 & ~ng1309;
  assign n2511 = ~new_n9650_ & ~new_n9651_;
  assign new_n9653_ = ng1309 & ~n2721;
  assign new_n9654_ = ~ng3103 & ~ng1309;
  assign n2516 = ~new_n9653_ & ~new_n9654_;
  assign new_n9656_ = ng1312 & ~ng1880;
  assign new_n9657_ = ~ng1312 & ~ng3176;
  assign n2521 = ~new_n9656_ & ~new_n9657_;
  assign new_n9659_ = ng823 & ~new_n9260_;
  assign new_n9660_ = ~ng198 & ~ng823;
  assign n2531 = ~new_n9659_ & ~new_n9660_;
  assign new_n9662_ = ng823 & ~new_n9271_;
  assign new_n9663_ = ~ng252 & ~ng823;
  assign n2536 = ~new_n9662_ & ~new_n9663_;
  assign new_n9665_ = ng121 & ~new_n5083_;
  assign new_n9666_ = ~new_n5082_1_ & ~new_n9665_;
  assign new_n9667_ = ~new_n4849_ & ~new_n5112_1_;
  assign new_n9668_ = new_n4849_ & new_n5112_1_;
  assign new_n9669_ = ~new_n9667_ & ~new_n9668_;
  assign new_n9670_ = new_n5082_1_ & new_n9669_;
  assign new_n9671_ = ~new_n9666_ & ~new_n9670_;
  assign new_n9672_ = ng826 & ~new_n9671_;
  assign new_n9673_ = ~ng213 & ~ng826;
  assign n2541 = ~new_n9672_ & ~new_n9673_;
  assign new_n9675_ = ~ng354 & ~new_n5138_;
  assign new_n9676_ = new_n5138_ & ~new_n8398_;
  assign n2546 = ~new_n9675_ & ~new_n9676_;
  assign new_n9678_ = ~ng398 & ~new_n5138_;
  assign new_n9679_ = new_n5138_ & ~new_n8947_;
  assign n2551 = ~new_n9678_ & ~new_n9679_;
  assign new_n9681_ = ng826 & new_n5212_1_;
  assign new_n9682_ = ~ng486 & ~ng826;
  assign n2570 = ~new_n9681_ & ~new_n9682_;
  assign new_n9684_ = ng1315 & ~ng510;
  assign new_n9685_ = ~ng1315 & ~ng630;
  assign n2580 = ~new_n9684_ & ~new_n9685_;
  assign new_n9687_ = ~ng711 & ~new_n5395_;
  assign new_n9688_ = ng660 & new_n5395_;
  assign n2585 = ~new_n9687_ & ~new_n9688_;
  assign new_n9690_ = ~ng830 & ~new_n5517_1_;
  assign new_n9691_ = ng793 & new_n5517_1_;
  assign n2590 = ~new_n9690_ & ~new_n9691_;
  assign new_n9693_ = ~ng860 & ~new_n5538_;
  assign new_n9694_ = ng789 & new_n5538_;
  assign n2595 = ~new_n9693_ & ~new_n9694_;
  assign new_n9696_ = ng826 & ~new_n9381_;
  assign new_n9697_ = ~ng873 & ~ng826;
  assign n2600 = ~new_n9696_ & ~new_n9697_;
  assign new_n9699_ = ng853 & new_n9024_;
  assign new_n9700_ = ~ng1101 & ~ng853;
  assign n2605 = ~new_n9699_ & ~new_n9700_;
  assign new_n9702_ = ng853 & ~new_n8525_;
  assign new_n9703_ = ~ng1122 & ~ng853;
  assign n2610 = ~new_n9702_ & ~new_n9703_;
  assign new_n9705_ = ng853 & ~new_n5924_;
  assign new_n9706_ = ~ng1148 & ~ng853;
  assign n2623 = ~new_n9705_ & ~new_n9706_;
  assign new_n9708_ = ng853 & ~new_n5560_;
  assign new_n9709_ = ~ng1158 & ~ng853;
  assign n2628 = ~new_n9708_ & ~new_n9709_;
  assign new_n9711_ = ~ng1270 & ~new_n6049_;
  assign new_n9712_ = ~pg3229 & ~new_n6055_;
  assign new_n9713_ = new_n6131_ & new_n9712_;
  assign new_n9714_ = pg3229 & new_n6055_;
  assign new_n9715_ = new_n6131_ & new_n9714_;
  assign new_n9716_ = ~new_n9713_ & ~new_n9715_;
  assign new_n9717_ = new_n6049_ & ~new_n9716_;
  assign n2633 = ~new_n9711_ & ~new_n9717_;
  assign new_n9719_ = ng1312 & ~new_n9412_;
  assign new_n9720_ = ~ng1312 & ~ng1285;
  assign n2638 = ~new_n9719_ & ~new_n9720_;
  assign new_n9722_ = ng1312 & ~new_n9421_;
  assign new_n9723_ = ~ng1312 & ~ng1180;
  assign n2643 = ~new_n9722_ & ~new_n9723_;
  assign new_n9725_ = ~ng1405 & ~new_n6263_;
  assign new_n9726_ = ng1365 & new_n6263_;
  assign n2648 = ~new_n9725_ & ~new_n9726_;
  assign new_n9728_ = ng1315 & ng1316;
  assign new_n9729_ = ~ng1414 & ~new_n9728_;
  assign new_n9730_ = ~new_n6044_ & new_n9728_;
  assign n2653 = ~new_n9729_ & ~new_n9730_;
  assign new_n9732_ = ~ng1515 & ~new_n5517_1_;
  assign new_n9733_ = ng1476 & new_n5517_1_;
  assign n2658 = ~new_n9732_ & ~new_n9733_;
  assign new_n9735_ = ~ng1530 & ~new_n5517_1_;
  assign new_n9736_ = ng1491 & new_n5517_1_;
  assign n2663 = ~new_n9735_ & ~new_n9736_;
  assign new_n9738_ = ~ng1532 & ~new_n4773_;
  assign new_n9739_ = ng1496 & new_n4773_;
  assign n2668 = ~new_n9738_ & ~new_n9739_;
  assign new_n9741_ = ~ng1541 & ~new_n4773_;
  assign new_n9742_ = new_n4773_ & ~new_n6436_;
  assign n2673 = ~new_n9741_ & ~new_n9742_;
  assign new_n9744_ = ng1435 & new_n9443_;
  assign new_n9745_ = ~ng1430 & new_n9744_;
  assign new_n9746_ = ng1430 & ~new_n9744_;
  assign new_n9747_ = ~new_n9745_ & ~new_n9746_;
  assign n2678 = ~new_n5127_1_ & ~new_n9747_;
  assign new_n9749_ = ~ng1754 & ~new_n6636_;
  assign new_n9750_ = new_n6636_ & ~new_n8738_;
  assign n2683 = ~new_n9749_ & ~new_n9750_;
  assign new_n9752_ = ng853 & ~new_n9459_;
  assign new_n9753_ = ~ng1807 & ~new_n9752_;
  assign new_n9754_ = new_n9456_ & new_n9752_;
  assign n2688 = ~new_n9753_ & ~new_n9754_;
  assign new_n9756_ = new_n6715_1_ & ~new_n6731_;
  assign new_n9757_ = ng2384 & new_n9756_;
  assign new_n9758_ = ~new_n6710_ & ~new_n6720_1_;
  assign new_n9759_ = ~new_n6726_ & new_n9758_;
  assign new_n9760_ = new_n6710_ & new_n6720_1_;
  assign new_n9761_ = new_n6726_ & new_n9760_;
  assign new_n9762_ = ~new_n9759_ & ~new_n9761_;
  assign new_n9763_ = ng2384 & ~new_n9762_;
  assign new_n9764_ = ~new_n9757_ & ~new_n9763_;
  assign new_n9765_ = ng853 & ~new_n9764_;
  assign new_n9766_ = ~ng1828 & ~new_n9765_;
  assign new_n9767_ = new_n9757_ & new_n9765_;
  assign n2693 = ~new_n9766_ & ~new_n9767_;
  assign new_n9769_ = ng823 & ~new_n9501_;
  assign new_n9770_ = ~ng1697 & ~ng823;
  assign n2698 = ~new_n9769_ & ~new_n9770_;
  assign new_n9772_ = ng2384 & ng823;
  assign new_n9773_ = ~ng1785 & ~new_n9772_;
  assign new_n9774_ = new_n9507_ & new_n9772_;
  assign n2703 = ~new_n9773_ & ~new_n9774_;
  assign new_n9776_ = ng853 & n5082;
  assign new_n9777_ = ~ng1845 & ~ng853;
  assign n2716 = ~new_n9776_ & ~new_n9777_;
  assign new_n9779_ = ~ng1956 & ~new_n6801_;
  assign new_n9780_ = ~new_n6807_ & new_n9117_;
  assign new_n9781_ = ~new_n9118_ & ~new_n9780_;
  assign new_n9782_ = ~new_n6812_ & new_n6882_1_;
  assign new_n9783_ = ~pg3229 & new_n9782_;
  assign new_n9784_ = ~pg3229 & new_n6822_;
  assign new_n9785_ = pg3229 & ~new_n6882_1_;
  assign new_n9786_ = ~new_n9783_ & ~new_n9784_;
  assign new_n9787_ = ~new_n9785_ & new_n9786_;
  assign new_n9788_ = new_n9781_ & new_n9787_;
  assign new_n9789_ = new_n6801_ & ~new_n9788_;
  assign n2726 = ~new_n9779_ & ~new_n9789_;
  assign new_n9791_ = ~ng1965 & ~new_n6801_;
  assign new_n9792_ = new_n6801_ & ~new_n9523_;
  assign n2731 = ~new_n9791_ & ~new_n9792_;
  assign new_n9794_ = ~ng2087 & ~new_n7007_;
  assign new_n9795_ = ng2026 & new_n7007_;
  assign n2746 = ~new_n9794_ & ~new_n9795_;
  assign new_n9797_ = ~ng2096 & ~new_n7007_;
  assign new_n9798_ = ng2046 & new_n7007_;
  assign n2751 = ~new_n9797_ & ~new_n9798_;
  assign new_n9800_ = ng1309 & ng2010;
  assign new_n9801_ = ~ng2112 & ~new_n9800_;
  assign new_n9802_ = ~new_n6785_ & new_n9800_;
  assign n2756 = ~new_n9801_ & ~new_n9802_;
  assign new_n9804_ = ~ng2206 & ~new_n5517_1_;
  assign new_n9805_ = ng2165 & new_n5517_1_;
  assign n2761 = ~new_n9804_ & ~new_n9805_;
  assign new_n9807_ = ~ng2245 & ~new_n5538_;
  assign new_n9808_ = ~ng2190 & ~ng2195;
  assign new_n9809_ = ng2200 & new_n9808_;
  assign new_n9810_ = ng2185 & new_n9809_;
  assign new_n9811_ = new_n5538_ & ~new_n9810_;
  assign n2766 = ~new_n9807_ & ~new_n9811_;
  assign new_n9813_ = ~ng2254 & ~new_n5538_;
  assign new_n9814_ = new_n5538_ & new_n7452_;
  assign n2771 = ~new_n9813_ & ~new_n9814_;
  assign new_n9816_ = ng823 & ~new_n9552_;
  assign new_n9817_ = ~ng2318 & ~ng823;
  assign n2776 = ~new_n9816_ & ~new_n9817_;
  assign new_n9819_ = ng823 & ~new_n9563_;
  assign new_n9820_ = ~ng2291 & ~ng823;
  assign n2781 = ~new_n9819_ & ~new_n9820_;
  assign new_n9822_ = ~new_n7020_ & ~new_n7323_;
  assign new_n9823_ = ~new_n7325_ & ~new_n9822_;
  assign new_n9824_ = ~new_n7322_ & new_n9823_;
  assign new_n9825_ = ~new_n7101_ & ~new_n7385_;
  assign new_n9826_ = new_n7101_ & new_n7385_;
  assign new_n9827_ = ~new_n9825_ & ~new_n9826_;
  assign new_n9828_ = new_n7322_ & new_n9827_;
  assign new_n9829_ = ~new_n9824_ & ~new_n9828_;
  assign new_n9830_ = ng826 & ~new_n9829_;
  assign new_n9831_ = ~ng2297 & ~ng826;
  assign n2786 = ~new_n9830_ & ~new_n9831_;
  assign new_n9833_ = ng2147 & ~new_n7397_;
  assign new_n9834_ = ~ng2147 & new_n7397_;
  assign new_n9835_ = ~new_n9833_ & ~new_n9834_;
  assign n2791 = ~new_n5127_1_ & ~new_n9835_;
  assign new_n9837_ = ~ng2421 & ~new_n7410_;
  assign new_n9838_ = new_n7410_ & ~new_n9591_;
  assign n2796 = ~new_n9837_ & ~new_n9838_;
  assign new_n9840_ = ~ng2466 & ~new_n7410_;
  assign new_n9841_ = new_n7416_1_ & new_n7430_;
  assign new_n9842_ = ~pg3229 & ~new_n7421_1_;
  assign new_n9843_ = new_n9841_ & new_n9842_;
  assign new_n9844_ = pg3229 & new_n7421_1_;
  assign new_n9845_ = new_n9841_ & new_n9844_;
  assign new_n9846_ = ~new_n9843_ & ~new_n9845_;
  assign new_n9847_ = new_n7410_ & ~new_n9846_;
  assign n2801 = ~new_n9840_ & ~new_n9847_;
  assign new_n9849_ = ng853 & new_n9180_;
  assign new_n9850_ = ~ng2396 & ~new_n9849_;
  assign new_n9851_ = new_n9187_ & new_n9849_;
  assign n2806 = ~new_n9850_ & ~new_n9851_;
  assign new_n9853_ = ng826 & new_n7489_;
  assign new_n9854_ = ~ng2561 & ~ng826;
  assign n2828 = ~new_n9853_ & ~new_n9854_;
  assign new_n9856_ = ~ng2652 & ~new_n7545_;
  assign new_n9857_ = new_n7545_ & ~new_n8870_;
  assign n2833 = ~new_n9856_ & ~new_n9857_;
  assign new_n9859_ = ng1312 & ~new_n9630_;
  assign new_n9860_ = ~ng2813 & ~new_n9859_;
  assign new_n9861_ = ng2704 & new_n9859_;
  assign n2848 = ~new_n9860_ & ~new_n9861_;
  assign new_n9863_ = ~ng533 & new_n7609_;
  assign new_n9864_ = ~new_n7605_ & new_n9863_;
  assign new_n9865_ = ~new_n5451_ & ~new_n7627_;
  assign new_n9866_ = ~new_n5287_1_ & ~new_n9865_;
  assign new_n9867_ = ~new_n9865_ & ~new_n9866_;
  assign new_n9868_ = ~new_n5287_1_ & ~new_n9866_;
  assign new_n9869_ = ~new_n9867_ & ~new_n9868_;
  assign new_n9870_ = new_n7609_ & ~new_n9869_;
  assign new_n9871_ = ng499 & new_n9870_;
  assign new_n9872_ = new_n7605_ & new_n9871_;
  assign new_n9873_ = ~new_n9864_ & ~new_n9872_;
  assign new_n9874_ = ~new_n7603_ & new_n9873_;
  assign n2853 = new_n9648_ | new_n9874_;
  assign new_n9876_ = ng1312 & ~ng2633;
  assign new_n9877_ = ~ng1312 & ~ng3095;
  assign n2858 = ~new_n9876_ & ~new_n9877_;
  assign new_n9879_ = ng1309 & ~n4713;
  assign new_n9880_ = ~ng3106 & ~ng1309;
  assign n2863 = ~new_n9879_ & ~new_n9880_;
  assign new_n9882_ = ~ng1186 & ng1312;
  assign new_n9883_ = ~ng1312 & ~ng3167;
  assign n2868 = ~new_n9882_ & ~new_n9883_;
  assign new_n9885_ = ng823 & ~new_n9671_;
  assign new_n9886_ = ~ng216 & ~ng823;
  assign n2878 = ~new_n9885_ & ~new_n9886_;
  assign new_n9888_ = ~ng92 & new_n5128_;
  assign new_n9889_ = ng92 & ~new_n5128_;
  assign new_n9890_ = ~new_n9888_ & ~new_n9889_;
  assign n2883 = ~new_n5127_1_ & ~new_n9890_;
  assign new_n9892_ = ~ng376 & ~new_n8937_;
  assign new_n9893_ = ~pg3229 & new_n5149_;
  assign new_n9894_ = new_n8388_ & new_n9893_;
  assign new_n9895_ = ~new_n8389_ & ~new_n9894_;
  assign new_n9896_ = ~new_n5149_ & ~new_n5158_;
  assign new_n9897_ = ~pg3229 & new_n9896_;
  assign new_n9898_ = new_n5149_ & ~new_n5158_;
  assign new_n9899_ = pg3229 & new_n9898_;
  assign new_n9900_ = ~new_n9897_ & ~new_n9899_;
  assign new_n9901_ = new_n9895_ & new_n9900_;
  assign new_n9902_ = new_n8937_ & ~new_n9901_;
  assign n2888 = ~new_n9892_ & ~new_n9902_;
  assign new_n9904_ = ~ng633 & new_n5382_;
  assign new_n9905_ = ng633 & ~new_n5382_;
  assign new_n9906_ = ~new_n9904_ & ~new_n9905_;
  assign n2912 = ~new_n5380_ & ~new_n9906_;
  assign new_n9908_ = ~ng698 & ~new_n5399_;
  assign new_n9909_ = ng640 & new_n5399_;
  assign n2917 = ~new_n9908_ & ~new_n9909_;
  assign new_n9911_ = ~ng840 & ~new_n4777_1_;
  assign new_n9912_ = ng805 & new_n4777_1_;
  assign n2922 = ~new_n9911_ & ~new_n9912_;
  assign new_n9914_ = ~ng861 & ~new_n6278_;
  assign new_n9915_ = ng789 & new_n6278_;
  assign n2927 = ~new_n9914_ & ~new_n9915_;
  assign new_n9917_ = ng826 & ~new_n5852_;
  assign new_n9918_ = ~ng918 & ~ng826;
  assign n2932 = ~new_n9917_ & ~new_n9918_;
  assign new_n9920_ = new_n5546_ & new_n5556_1_;
  assign new_n9921_ = new_n5551_ & ~new_n9920_;
  assign new_n9922_ = ng2257 & new_n7933_;
  assign new_n9923_ = ~new_n5634_1_ & new_n9922_;
  assign new_n9924_ = ~new_n5827_ & ~new_n9923_;
  assign new_n9925_ = new_n5821_ & new_n7935_;
  assign new_n9926_ = new_n9924_ & ~new_n9925_;
  assign new_n9927_ = ~new_n5675_ & new_n9926_;
  assign new_n9928_ = new_n5556_1_ & new_n9927_;
  assign new_n9929_ = ~new_n5825_ & ~new_n5827_;
  assign new_n9930_ = ~new_n5556_1_ & new_n9929_;
  assign new_n9931_ = ~new_n9928_ & ~new_n9930_;
  assign new_n9932_ = new_n5546_ & new_n9931_;
  assign new_n9933_ = ~new_n5675_ & new_n7935_;
  assign new_n9934_ = ~new_n5710_ & ~new_n9933_;
  assign new_n9935_ = new_n5556_1_ & new_n9934_;
  assign new_n9936_ = ~new_n5556_1_ & ~new_n5710_;
  assign new_n9937_ = ~new_n9935_ & ~new_n9936_;
  assign new_n9938_ = ~new_n5546_ & new_n9937_;
  assign new_n9939_ = ~new_n9932_ & ~new_n9938_;
  assign new_n9940_ = ~new_n5551_ & new_n9939_;
  assign new_n9941_ = ~new_n9921_ & ~new_n9940_;
  assign new_n9942_ = ~new_n5546_ & new_n9941_;
  assign new_n9943_ = ~new_n5546_ & ~new_n9942_;
  assign new_n9944_ = new_n9941_ & ~new_n9942_;
  assign new_n9945_ = ~new_n9943_ & ~new_n9944_;
  assign new_n9946_ = ~new_n5836_ & new_n9945_;
  assign new_n9947_ = ng826 & ~new_n9946_;
  assign new_n9948_ = ~ng1002 & ~ng826;
  assign n2937 = ~new_n9947_ & ~new_n9948_;
  assign new_n9950_ = ~ng1089 & ~new_n9505_;
  assign new_n9951_ = new_n6005_ & new_n9505_;
  assign n2942 = ~new_n9950_ & ~new_n9951_;
  assign new_n9953_ = ng826 & ~new_n5824_;
  assign new_n9954_ = ~ng1164 & ~ng826;
  assign n2957 = ~new_n9953_ & ~new_n9954_;
  assign new_n9956_ = ~ng1272 & ~new_n8012_;
  assign new_n9957_ = new_n8012_ & ~new_n9716_;
  assign n2966 = ~new_n9956_ & ~new_n9957_;
  assign new_n9959_ = ng1315 & ~new_n9412_;
  assign new_n9960_ = ~ng1315 & ~ng1288;
  assign n2971 = ~new_n9959_ & ~new_n9960_;
  assign new_n9962_ = ~ng1409 & ~new_n6259_1_;
  assign new_n9963_ = ng1372 & new_n6259_1_;
  assign n2981 = ~new_n9962_ & ~new_n9963_;
  assign new_n9965_ = ~ng1417 & ~new_n9728_;
  assign new_n9966_ = ~new_n6033_ & new_n9728_;
  assign n2986 = ~new_n9965_ & ~new_n9966_;
  assign new_n9968_ = ~ng1512 & ~new_n5517_1_;
  assign new_n9969_ = ng1471 & new_n5517_1_;
  assign n2991 = ~new_n9968_ & ~new_n9969_;
  assign new_n9971_ = ~ng1526 & ~new_n4773_;
  assign new_n9972_ = ng1486 & new_n4773_;
  assign n2996 = ~new_n9971_ & ~new_n9972_;
  assign new_n9974_ = ~ng1536 & ~new_n5517_1_;
  assign new_n9975_ = ng1501 & new_n5517_1_;
  assign n3001 = ~new_n9974_ & ~new_n9975_;
  assign new_n9977_ = ~ng1544 & ~new_n4773_;
  assign new_n9978_ = new_n4773_ & ~new_n6395_;
  assign n3006 = ~new_n9977_ & ~new_n9978_;
  assign new_n9980_ = ng1430 & new_n9744_;
  assign new_n9981_ = ng1426 & ~new_n9980_;
  assign new_n9982_ = ~ng1426 & new_n9980_;
  assign new_n9983_ = ~new_n9981_ & ~new_n9982_;
  assign n3011 = ~new_n5127_1_ & ~new_n9983_;
  assign new_n9985_ = ~ng1769 & ~new_n6636_;
  assign new_n9986_ = new_n6642_ & new_n6656_;
  assign new_n9987_ = ~pg3229 & ~new_n6647_;
  assign new_n9988_ = new_n9986_ & new_n9987_;
  assign new_n9989_ = pg3229 & new_n6647_;
  assign new_n9990_ = new_n9986_ & new_n9989_;
  assign new_n9991_ = ~new_n9988_ & ~new_n9990_;
  assign new_n9992_ = new_n6636_ & ~new_n9991_;
  assign n3016 = ~new_n9985_ & ~new_n9992_;
  assign new_n9994_ = ng853 & new_n6702_;
  assign new_n9995_ = ~ng1804 & ~ng853;
  assign n3021 = ~new_n9994_ & ~new_n9995_;
  assign new_n9997_ = ng823 & ~new_n9764_;
  assign new_n9998_ = ~ng1830 & ~new_n9997_;
  assign new_n9999_ = new_n9757_ & new_n9997_;
  assign n3026 = ~new_n9998_ & ~new_n9999_;
  assign new_n10001_ = ng853 & ~new_n9501_;
  assign new_n10002_ = ~ng1698 & ~ng853;
  assign n3031 = ~new_n10001_ & ~new_n10002_;
  assign new_n10004_ = ng823 & new_n6710_;
  assign new_n10005_ = ~ng1868 & ~ng823;
  assign n3046 = ~new_n10004_ & ~new_n10005_;
  assign new_n10007_ = ng853 & ~new_n6572_;
  assign new_n10008_ = ~ng1860 & ~ng853;
  assign n3051 = ~new_n10007_ & ~new_n10008_;
  assign new_n10010_ = ~ng1957 & ~new_n8088_;
  assign new_n10011_ = new_n8088_ & ~new_n9788_;
  assign n3061 = ~new_n10010_ & ~new_n10011_;
  assign new_n10013_ = ng1309 & ~new_n6840_;
  assign new_n10014_ = ~ng1967 & ~ng1309;
  assign n3066 = ~new_n10013_ & ~new_n10014_;
  assign new_n10016_ = ng2026 & new_n8104_;
  assign new_n10017_ = ng2040 & ~new_n10016_;
  assign new_n10018_ = ~ng2040 & new_n10016_;
  assign new_n10019_ = ~new_n10017_ & ~new_n10018_;
  assign n3071 = ~new_n6993_ & ~new_n10019_;
  assign new_n10021_ = ~ng2081 & ~new_n7007_;
  assign new_n10022_ = ng2013 & new_n7007_;
  assign n3076 = ~new_n10021_ & ~new_n10022_;
  assign new_n10024_ = ~ng2091 & ~new_n7003_;
  assign new_n10025_ = ng2040 & new_n7003_;
  assign n3081 = ~new_n10024_ & ~new_n10025_;
  assign new_n10027_ = ~ng2099 & ~new_n7007_;
  assign new_n10028_ = ng2059 & new_n7007_;
  assign n3086 = ~new_n10027_ & ~new_n10028_;
  assign new_n10030_ = ~ng2109 & ~new_n9800_;
  assign new_n10031_ = ~new_n6796_ & new_n9800_;
  assign n3091 = ~new_n10030_ & ~new_n10031_;
  assign new_n10033_ = ~ng2010 & ~new_n7002_;
  assign new_n10034_ = ng1315 & ~new_n10033_;
  assign new_n10035_ = ~ng2117 & ~new_n10034_;
  assign new_n10036_ = ng2010 & new_n10034_;
  assign n3096 = ~new_n10035_ & ~new_n10036_;
  assign new_n10038_ = ~ng2246 & ~new_n6278_;
  assign new_n10039_ = new_n6278_ & ~new_n9810_;
  assign n3101 = ~new_n10038_ & ~new_n10039_;
  assign new_n10041_ = ng2165 & ~new_n7323_;
  assign new_n10042_ = ~new_n7322_ & ~new_n10041_;
  assign new_n10043_ = ~new_n7045_ & new_n7087_1_;
  assign new_n10044_ = new_n7045_ & ~new_n7087_1_;
  assign new_n10045_ = ~new_n10043_ & ~new_n10044_;
  assign new_n10046_ = new_n7322_ & new_n10045_;
  assign new_n10047_ = ~new_n10042_ & ~new_n10046_;
  assign new_n10048_ = ng826 & ~new_n10047_;
  assign new_n10049_ = ~ng2261 & ~ng826;
  assign n3106 = ~new_n10048_ & ~new_n10049_;
  assign new_n10051_ = ng823 & ~new_n8132_;
  assign new_n10052_ = ~ng2273 & ~ng823;
  assign n3111 = ~new_n10051_ & ~new_n10052_;
  assign new_n10054_ = ng826 & ~new_n9563_;
  assign new_n10055_ = ~ng2288 & ~ng826;
  assign n3116 = ~new_n10054_ & ~new_n10055_;
  assign new_n10057_ = ng823 & ~new_n9829_;
  assign new_n10058_ = ~ng2300 & ~ng823;
  assign n3121 = ~new_n10057_ & ~new_n10058_;
  assign new_n10060_ = ~ng2133 & new_n7400_;
  assign new_n10061_ = ng2133 & ~new_n7400_;
  assign new_n10062_ = ~new_n10060_ & ~new_n10061_;
  assign n3126 = ~new_n5127_1_ & ~new_n10062_;
  assign new_n10064_ = ~ng2463 & ~new_n9171_;
  assign new_n10065_ = new_n9171_ & ~new_n9846_;
  assign n3136 = ~new_n10064_ & ~new_n10065_;
  assign new_n10067_ = ~ng2478 & ~new_n6003_;
  assign new_n10068_ = new_n7307_ & new_n7319_1_;
  assign new_n10069_ = new_n6003_ & new_n10068_;
  assign n3141 = ~new_n10067_ & ~new_n10069_;
  assign new_n10071_ = ~ng2656 & ~new_n9196_;
  assign new_n10072_ = ~pg3229 & new_n7561_;
  assign new_n10073_ = new_n7563_ & new_n10072_;
  assign new_n10074_ = ~new_n7564_ & ~new_n10073_;
  assign new_n10075_ = ~new_n7556_ & ~new_n7561_;
  assign new_n10076_ = ~pg3229 & new_n10075_;
  assign new_n10077_ = ~new_n7556_ & new_n7561_;
  assign new_n10078_ = pg3229 & new_n10077_;
  assign new_n10079_ = ~new_n10076_ & ~new_n10078_;
  assign new_n10080_ = new_n10074_ & new_n10079_;
  assign new_n10081_ = new_n9196_ & ~new_n10080_;
  assign n3170 = ~new_n10071_ & ~new_n10081_;
  assign new_n10083_ = ng1315 & ~new_n9617_;
  assign new_n10084_ = ~ng1315 & ~ng2676;
  assign n3175 = ~new_n10083_ & ~new_n10084_;
  assign new_n10086_ = ng1315 & ~new_n9630_;
  assign new_n10087_ = ~ng2811 & ~new_n10086_;
  assign new_n10088_ = ng2704 & new_n10086_;
  assign n3185 = ~new_n10087_ & ~new_n10088_;
  assign new_n10090_ = ng1315 & ~ng2633;
  assign new_n10091_ = ~ng1315 & ~ng3096;
  assign n3190 = ~new_n10090_ & ~new_n10091_;
  assign new_n10093_ = ng1315 & ~n2721;
  assign new_n10094_ = ~ng1315 & ~ng3105;
  assign n3195 = ~new_n10093_ & ~new_n10094_;
  assign new_n10096_ = ~ng1186 & ng1315;
  assign new_n10097_ = ~ng1315 & ~ng3170;
  assign n3200 = ~new_n10096_ & ~new_n10097_;
  assign new_n10099_ = ng853 & ~new_n9671_;
  assign new_n10100_ = ~ng219 & ~ng853;
  assign n3210 = ~new_n10099_ & ~new_n10100_;
  assign new_n10102_ = ng853 & ~new_n9286_;
  assign new_n10103_ = ~ng273 & ~ng853;
  assign n3215 = ~new_n10102_ & ~new_n10103_;
  assign new_n10105_ = ~ng56 & new_n9293_;
  assign new_n10106_ = ng56 & ~new_n9293_;
  assign new_n10107_ = ~new_n10105_ & ~new_n10106_;
  assign n3220 = ~new_n5127_1_ & ~new_n10107_;
  assign new_n10109_ = ng640 & ~new_n5381_;
  assign new_n10110_ = ~ng640 & new_n5381_;
  assign new_n10111_ = ~new_n10109_ & ~new_n10110_;
  assign n3242 = ~new_n5380_ & ~new_n10111_;
  assign new_n10113_ = ng653 & ~new_n5383_1_;
  assign new_n10114_ = ~ng653 & new_n5383_1_;
  assign new_n10115_ = ~new_n10113_ & ~new_n10114_;
  assign n3247 = ~new_n5380_ & ~new_n10115_;
  assign new_n10117_ = ~ng847 & ~new_n4773_;
  assign new_n10118_ = new_n4773_ & ~new_n5529_;
  assign n3252 = ~new_n10117_ & ~new_n10118_;
  assign new_n10120_ = ~ng859 & ~new_n8121_;
  assign new_n10121_ = ng789 & new_n8121_;
  assign n3257 = ~new_n10120_ & ~new_n10121_;
  assign new_n10123_ = ng853 & ~new_n9381_;
  assign new_n10124_ = ~ng879 & ~ng853;
  assign n3262 = ~new_n10123_ & ~new_n10124_;
  assign new_n10126_ = ng823 & ~new_n9946_;
  assign new_n10127_ = ~ng1003 & ~ng823;
  assign n3267 = ~new_n10126_ & ~new_n10127_;
  assign new_n10129_ = ~ng1091 & ~new_n9772_;
  assign new_n10130_ = new_n6005_ & new_n9772_;
  assign n3272 = ~new_n10129_ & ~new_n10130_;
  assign new_n10132_ = ~ng1262 & ~new_n8562_;
  assign new_n10133_ = new_n8562_ & ~new_n9409_;
  assign n3289 = ~new_n10132_ & ~new_n10133_;
  assign new_n10135_ = ~ng1271 & ~new_n8562_;
  assign new_n10136_ = new_n8562_ & ~new_n9716_;
  assign n3294 = ~new_n10135_ & ~new_n10136_;
  assign new_n10138_ = ng1309 & ~new_n6237_;
  assign new_n10139_ = ~ng1300 & ~ng1309;
  assign n3299 = ~new_n10138_ & ~new_n10139_;
  assign new_n10141_ = ~ng1410 & ~new_n6255_;
  assign new_n10142_ = ng1372 & new_n6255_;
  assign n3309 = ~new_n10141_ & ~new_n10142_;
  assign new_n10144_ = ~ng1419 & ~new_n6241_;
  assign new_n10145_ = ~new_n6033_ & new_n6241_;
  assign n3314 = ~new_n10144_ & ~new_n10145_;
  assign new_n10147_ = ~ng1513 & ~new_n4777_1_;
  assign new_n10148_ = ng1471 & new_n4777_1_;
  assign n3319 = ~new_n10147_ & ~new_n10148_;
  assign new_n10150_ = ~ng1528 & ~new_n4777_1_;
  assign new_n10151_ = ng1486 & new_n4777_1_;
  assign n3324 = ~new_n10150_ & ~new_n10151_;
  assign new_n10153_ = ~ng1537 & ~new_n4777_1_;
  assign new_n10154_ = ng1501 & new_n4777_1_;
  assign n3329 = ~new_n10153_ & ~new_n10154_;
  assign new_n10156_ = ~ng1546 & ~new_n4777_1_;
  assign new_n10157_ = new_n4777_1_ & ~new_n6395_;
  assign n3334 = ~new_n10156_ & ~new_n10157_;
  assign new_n10159_ = ~ng1735 & ~new_n8072_;
  assign new_n10160_ = ~new_n6642_ & new_n8728_;
  assign new_n10161_ = ~new_n8729_ & ~new_n10160_;
  assign new_n10162_ = ~new_n6647_ & new_n8726_;
  assign new_n10163_ = ~pg3229 & new_n10162_;
  assign new_n10164_ = ~pg3229 & new_n6657_1_;
  assign new_n10165_ = pg3229 & ~new_n8726_;
  assign new_n10166_ = ~new_n10163_ & ~new_n10164_;
  assign new_n10167_ = ~new_n10165_ & new_n10166_;
  assign new_n10168_ = new_n10161_ & new_n10167_;
  assign new_n10169_ = new_n8072_ & ~new_n10168_;
  assign n3339 = ~new_n10159_ & ~new_n10169_;
  assign new_n10171_ = ~ng1779 & ~new_n8072_;
  assign new_n10172_ = new_n8072_ & ~new_n9991_;
  assign n3344 = ~new_n10171_ & ~new_n10172_;
  assign new_n10174_ = ng826 & ~new_n9459_;
  assign new_n10175_ = ~ng1808 & ~new_n10174_;
  assign new_n10176_ = new_n9456_ & new_n10174_;
  assign n3349 = ~new_n10175_ & ~new_n10176_;
  assign new_n10178_ = ng826 & ~new_n9764_;
  assign new_n10179_ = ~ng1829 & ~new_n10178_;
  assign new_n10180_ = new_n9757_ & new_n10178_;
  assign n3354 = ~new_n10179_ & ~new_n10180_;
  assign new_n10182_ = ng826 & ~new_n6771_;
  assign new_n10183_ = ~ng1699 & ~ng826;
  assign n3359 = ~new_n10182_ & ~new_n10183_;
  assign new_n10185_ = ng826 & new_n6710_;
  assign new_n10186_ = ~ng1867 & ~ng826;
  assign n3372 = ~new_n10185_ & ~new_n10186_;
  assign new_n10188_ = ng826 & n5082;
  assign new_n10189_ = ~ng1861 & ~ng826;
  assign n3377 = ~new_n10188_ & ~new_n10189_;
  assign new_n10191_ = ~ng1859 & ng1315;
  assign new_n10192_ = ~ng1860 & ng1309;
  assign new_n10193_ = ~ng1858 & ng1312;
  assign new_n10194_ = ~new_n10191_ & ~new_n10192_;
  assign n3382 = ~new_n10193_ & new_n10194_;
  assign new_n10196_ = ~ng1955 & ~new_n8779_;
  assign new_n10197_ = new_n8779_ & ~new_n9788_;
  assign n3386 = ~new_n10196_ & ~new_n10197_;
  assign new_n10199_ = ~ng1964 & ~new_n8779_;
  assign new_n10200_ = new_n8779_ & ~new_n9523_;
  assign n3391 = ~new_n10199_ & ~new_n10200_;
  assign new_n10202_ = ng2040 & new_n10016_;
  assign new_n10203_ = ~ng2052 & new_n10202_;
  assign new_n10204_ = ng2052 & ~new_n10202_;
  assign new_n10205_ = ~new_n10203_ & ~new_n10204_;
  assign n3396 = ~new_n6993_ & ~new_n10205_;
  assign new_n10207_ = ~ng2083 & ~new_n7011_;
  assign new_n10208_ = ng2013 & new_n7011_;
  assign n3401 = ~new_n10207_ & ~new_n10208_;
  assign new_n10210_ = ~ng2092 & ~new_n7011_;
  assign new_n10211_ = ng2040 & new_n7011_;
  assign n3406 = ~new_n10210_ & ~new_n10211_;
  assign new_n10213_ = ~ng2101 & ~new_n7011_;
  assign new_n10214_ = ng2059 & new_n7011_;
  assign n3411 = ~new_n10213_ & ~new_n10214_;
  assign new_n10216_ = ~ng2110 & ~new_n6993_;
  assign new_n10217_ = ~new_n6796_ & new_n6993_;
  assign n3416 = ~new_n10216_ & ~new_n10217_;
  assign new_n10219_ = ng1312 & ~new_n10033_;
  assign new_n10220_ = ~ng2119 & ~new_n10219_;
  assign new_n10221_ = ng2010 & new_n10219_;
  assign n3421 = ~new_n10220_ & ~new_n10221_;
  assign new_n10223_ = ~ng2244 & ~new_n8121_;
  assign new_n10224_ = new_n8121_ & ~new_n9810_;
  assign n3426 = ~new_n10223_ & ~new_n10224_;
  assign new_n10226_ = ~ng2253 & ~new_n8121_;
  assign new_n10227_ = new_n7452_ & new_n8121_;
  assign n3431 = ~new_n10226_ & ~new_n10227_;
  assign new_n10229_ = ng853 & ~new_n8132_;
  assign new_n10230_ = ~ng2276 & ~ng853;
  assign n3436 = ~new_n10229_ & ~new_n10230_;
  assign new_n10232_ = ng853 & ~new_n7362_;
  assign new_n10233_ = ~ng2330 & ~ng853;
  assign n3441 = ~new_n10232_ & ~new_n10233_;
  assign new_n10235_ = ng853 & ~new_n9829_;
  assign new_n10236_ = ~ng2303 & ~ng853;
  assign n3446 = ~new_n10235_ & ~new_n10236_;
  assign new_n10238_ = ng2138 & ~new_n7399_;
  assign new_n10239_ = ~ng2138 & new_n7399_;
  assign new_n10240_ = ~new_n10238_ & ~new_n10239_;
  assign n3451 = ~new_n5127_1_ & ~new_n10240_;
  assign new_n10242_ = ~ng2429 & ~new_n8146_;
  assign new_n10243_ = new_n8146_ & ~new_n9591_;
  assign n3456 = ~new_n10242_ & ~new_n10243_;
  assign new_n10245_ = ~ng2473 & ~new_n8146_;
  assign new_n10246_ = new_n8146_ & ~new_n9846_;
  assign n3461 = ~new_n10245_ & ~new_n10246_;
  assign new_n10248_ = ~ng2479 & ~new_n9772_;
  assign new_n10249_ = new_n9772_ & new_n10068_;
  assign n3466 = ~new_n10248_ & ~new_n10249_;
  assign new_n10251_ = ~ng2657 & ~new_n8209_;
  assign new_n10252_ = new_n8209_ & ~new_n10080_;
  assign n3491 = ~new_n10251_ & ~new_n10252_;
  assign new_n10254_ = ng1312 & ~new_n9617_;
  assign new_n10255_ = ~ng1312 & ~ng2673;
  assign n3496 = ~new_n10254_ & ~new_n10255_;
  assign new_n10257_ = ng1312 & ~new_n9626_;
  assign new_n10258_ = ~ng1312 & ~ng2568;
  assign n3501 = ~new_n10257_ & ~new_n10258_;
  assign new_n10260_ = ~ng536 & new_n7609_;
  assign new_n10261_ = ~new_n7605_ & new_n10260_;
  assign new_n10262_ = ~new_n5422_1_ & ~new_n7627_;
  assign new_n10263_ = ~new_n5287_1_ & ~new_n10262_;
  assign new_n10264_ = ~new_n10262_ & ~new_n10263_;
  assign new_n10265_ = ~new_n5287_1_ & ~new_n10263_;
  assign new_n10266_ = ~new_n10264_ & ~new_n10265_;
  assign new_n10267_ = new_n7609_ & ~new_n10266_;
  assign new_n10268_ = ng499 & new_n10267_;
  assign new_n10269_ = new_n7605_ & new_n10268_;
  assign new_n10270_ = ~new_n10261_ & ~new_n10269_;
  assign new_n10271_ = ~new_n7603_ & new_n10270_;
  assign new_n10272_ = ~new_n5462_ & ~new_n7627_;
  assign new_n10273_ = ~new_n5287_1_ & ~new_n10272_;
  assign new_n10274_ = ~new_n10272_ & ~new_n10273_;
  assign new_n10275_ = ~new_n5287_1_ & ~new_n10273_;
  assign new_n10276_ = ~new_n10274_ & ~new_n10275_;
  assign new_n10277_ = new_n7609_ & ~new_n10276_;
  assign new_n10278_ = ng499 & new_n10277_;
  assign new_n10279_ = new_n7638_ & ~new_n10278_;
  assign new_n10280_ = new_n7603_ & new_n10279_;
  assign n3506 = new_n10271_ | new_n10280_;
  assign new_n10282_ = ng2888 & ~new_n9235_;
  assign new_n10283_ = ~ng2888 & new_n9235_;
  assign new_n10284_ = ~new_n10282_ & ~new_n10283_;
  assign n3511 = new_n9234_ & ~new_n10284_;
  assign new_n10286_ = ~ng130 & ~new_n5517_1_;
  assign new_n10287_ = ng97 & new_n5517_1_;
  assign n3516 = ~new_n10286_ & ~new_n10287_;
  assign new_n10289_ = ~ng144 & ~new_n4773_;
  assign new_n10290_ = ng109 & new_n4773_;
  assign n3521 = ~new_n10289_ & ~new_n10290_;
  assign new_n10292_ = ~ng158 & ~new_n4777_1_;
  assign new_n10293_ = ng125 & new_n4777_1_;
  assign n3526 = ~new_n10292_ & ~new_n10293_;
  assign new_n10295_ = ~ng172 & ~new_n5538_;
  assign new_n10296_ = ng101 & new_n5538_;
  assign n3531 = ~new_n10295_ & ~new_n10296_;
  assign new_n10298_ = ng97 & ~new_n5083_;
  assign new_n10299_ = ~new_n5082_1_ & ~new_n10298_;
  assign new_n10300_ = ~new_n4800_ & new_n4842_1_;
  assign new_n10301_ = new_n4800_ & ~new_n4842_1_;
  assign new_n10302_ = ~new_n10300_ & ~new_n10301_;
  assign new_n10303_ = new_n5082_1_ & new_n10302_;
  assign new_n10304_ = ~new_n10299_ & ~new_n10303_;
  assign new_n10305_ = ng853 & ~new_n10304_;
  assign new_n10306_ = ~ng192 & ~ng853;
  assign n3536 = ~new_n10305_ & ~new_n10306_;
  assign new_n10308_ = ng113 & ~new_n5083_;
  assign new_n10309_ = ~new_n5082_1_ & ~new_n10308_;
  assign new_n10310_ = ~new_n4832_1_ & ~new_n5111_;
  assign new_n10311_ = new_n4832_1_ & new_n5111_;
  assign new_n10312_ = ~new_n10310_ & ~new_n10311_;
  assign new_n10313_ = new_n5082_1_ & new_n10312_;
  assign new_n10314_ = ~new_n10309_ & ~new_n10313_;
  assign new_n10315_ = ng823 & ~new_n10314_;
  assign new_n10316_ = ~ng207 & ~ng823;
  assign n3541 = ~new_n10315_ & ~new_n10316_;
  assign new_n10318_ = ng823 & ~new_n8412_;
  assign new_n10319_ = ~ng449 & ~new_n10318_;
  assign new_n10320_ = new_n8405_ & new_n10318_;
  assign n3546 = ~new_n10319_ & ~new_n10320_;
  assign new_n10322_ = ~ng2384 & new_n5068_;
  assign new_n10323_ = ~new_n5068_ & ~new_n5260_;
  assign new_n10324_ = ~new_n10322_ & ~new_n10323_;
  assign new_n10325_ = ng826 & new_n10324_;
  assign new_n10326_ = ~ng322 & ~new_n10325_;
  assign new_n10327_ = ~new_n4795_ & new_n5067_1_;
  assign new_n10328_ = new_n4785_ & new_n10327_;
  assign new_n10329_ = new_n4795_ & new_n5057_1_;
  assign new_n10330_ = ~new_n10328_ & ~new_n10329_;
  assign new_n10331_ = ~new_n4790_ & ~new_n10330_;
  assign new_n10332_ = new_n10325_ & new_n10331_;
  assign n3551 = ~new_n10326_ & ~new_n10332_;
  assign new_n10334_ = ~ng578 & ~new_n5307_;
  assign new_n10335_ = new_n5307_ & ~new_n8431_;
  assign n3571 = ~new_n10334_ & ~new_n10335_;
  assign new_n10337_ = ~new_n5366_ & ~new_n7855_;
  assign new_n10338_ = ng1312 & ~new_n10337_;
  assign new_n10339_ = ~ng1312 & ~ng599;
  assign n3576 = ~new_n10338_ & ~new_n10339_;
  assign new_n10341_ = ~ng700 & ~new_n5391_;
  assign new_n10342_ = ng640 & new_n5391_;
  assign n3591 = ~new_n10341_ & ~new_n10342_;
  assign new_n10344_ = ~ng838 & ~new_n4773_;
  assign new_n10345_ = ng805 & new_n4773_;
  assign n3596 = ~new_n10344_ & ~new_n10345_;
  assign new_n10347_ = ~ng852 & ~new_n4777_1_;
  assign new_n10348_ = new_n4777_1_ & ~new_n5652_;
  assign n3601 = ~new_n10347_ & ~new_n10348_;
  assign new_n10350_ = ~ng866 & ~new_n5538_;
  assign new_n10351_ = new_n5538_ & new_n5967_1_;
  assign n3606 = ~new_n10350_ & ~new_n10351_;
  assign new_n10353_ = ng801 & ~new_n5839_;
  assign new_n10354_ = ~new_n5838_1_ & ~new_n10353_;
  assign new_n10355_ = ~new_n5593_ & ~new_n5872_;
  assign new_n10356_ = new_n5593_ & new_n5872_;
  assign new_n10357_ = ~new_n10355_ & ~new_n10356_;
  assign new_n10358_ = new_n5838_1_ & new_n10357_;
  assign new_n10359_ = ~new_n10354_ & ~new_n10358_;
  assign new_n10360_ = ng823 & ~new_n10359_;
  assign new_n10361_ = ~ng894 & ~ng823;
  assign n3611 = ~new_n10360_ & ~new_n10361_;
  assign new_n10363_ = ng826 & ~new_n8494_;
  assign new_n10364_ = ~ng909 & ~ng826;
  assign n3616 = ~new_n10363_ & ~new_n10364_;
  assign new_n10366_ = ng1312 & ~new_n8573_;
  assign new_n10367_ = ~ng1312 & ~ng1294;
  assign n3645 = ~new_n10366_ & ~new_n10367_;
  assign new_n10369_ = ~ng1332 & new_n6245_;
  assign new_n10370_ = ng1332 & ~new_n6245_;
  assign new_n10371_ = ~new_n10369_ & ~new_n10370_;
  assign n3655 = ~new_n6241_ & ~new_n10371_;
  assign new_n10373_ = ~ng1389 & ~new_n6255_;
  assign new_n10374_ = ng1319 & new_n6255_;
  assign n3660 = ~new_n10373_ & ~new_n10374_;
  assign new_n10376_ = ~ng1400 & ~new_n6259_1_;
  assign new_n10377_ = ng1358 & new_n6259_1_;
  assign n3665 = ~new_n10376_ & ~new_n10377_;
  assign new_n10379_ = ~ng1560 & ~new_n5538_;
  assign new_n10380_ = new_n5538_ & new_n6678_;
  assign n3670 = ~new_n10379_ & ~new_n10380_;
  assign new_n10382_ = ng1481 & ~new_n6587_;
  assign new_n10383_ = ~new_n6301_ & new_n6587_;
  assign new_n10384_ = ~new_n10382_ & ~new_n10383_;
  assign new_n10385_ = ~new_n6586_ & new_n10384_;
  assign new_n10386_ = ~new_n6309_1_ & ~new_n6600_1_;
  assign new_n10387_ = new_n6309_1_ & new_n6600_1_;
  assign new_n10388_ = ~new_n10386_ & ~new_n10387_;
  assign new_n10389_ = new_n6586_ & new_n10388_;
  assign new_n10390_ = ~new_n10385_ & ~new_n10389_;
  assign new_n10391_ = ng853 & ~new_n10390_;
  assign new_n10392_ = ~ng1582 & ~ng853;
  assign n3675 = ~new_n10391_ & ~new_n10392_;
  assign new_n10394_ = ng1501 & ~new_n6587_;
  assign new_n10395_ = ~new_n6586_ & ~new_n10394_;
  assign new_n10396_ = ~new_n6353_1_ & ~new_n6616_;
  assign new_n10397_ = new_n6353_1_ & new_n6616_;
  assign new_n10398_ = ~new_n10396_ & ~new_n10397_;
  assign new_n10399_ = new_n6586_ & new_n10398_;
  assign new_n10400_ = ~new_n10395_ & ~new_n10399_;
  assign new_n10401_ = ng823 & ~new_n10400_;
  assign new_n10402_ = ~ng1597 & ~ng823;
  assign n3680 = ~new_n10401_ & ~new_n10402_;
  assign new_n10404_ = ~ng1466 & new_n5128_;
  assign new_n10405_ = ng1466 & ~new_n5128_;
  assign new_n10406_ = ~new_n10404_ & ~new_n10405_;
  assign n3685 = ~new_n5127_1_ & ~new_n10406_;
  assign new_n10408_ = ~ng2217 & ~new_n4773_;
  assign new_n10409_ = ng2175 & new_n4773_;
  assign n3710 = ~new_n10408_ & ~new_n10409_;
  assign new_n10411_ = ~ng2231 & ~new_n4777_1_;
  assign new_n10412_ = ng2195 & new_n4777_1_;
  assign n3715 = ~new_n10411_ & ~new_n10412_;
  assign new_n10414_ = ~ng2248 & ~new_n5538_;
  assign new_n10415_ = ng2170 & new_n5538_;
  assign n3720 = ~new_n10414_ & ~new_n10415_;
  assign new_n10417_ = n2815 & ~new_n7454_;
  assign new_n10418_ = ~n2815 & new_n8830_;
  assign new_n10419_ = ~new_n10417_ & ~new_n10418_;
  assign new_n10420_ = new_n7459_ & ~new_n10419_;
  assign new_n10421_ = ~new_n7445_ & new_n10420_;
  assign new_n10422_ = ng2384 & new_n10421_;
  assign new_n10423_ = new_n7445_ & ~new_n10419_;
  assign new_n10424_ = ng2384 & new_n10423_;
  assign new_n10425_ = ~new_n10422_ & ~new_n10424_;
  assign new_n10426_ = ng823 & ~new_n10425_;
  assign new_n10427_ = ~ng2503 & ~new_n10426_;
  assign new_n10428_ = new_n10422_ & new_n10426_;
  assign n3725 = ~new_n10427_ & ~new_n10428_;
  assign new_n10430_ = ~new_n7030_ & new_n7040_;
  assign new_n10431_ = new_n7035_ & new_n10430_;
  assign new_n10432_ = new_n7030_ & ~new_n7040_;
  assign new_n10433_ = ~new_n7195_ & ~new_n10432_;
  assign new_n10434_ = ~new_n7035_ & ~new_n10433_;
  assign new_n10435_ = ~new_n10431_ & ~new_n10434_;
  assign new_n10436_ = ~new_n7035_ & new_n10435_;
  assign new_n10437_ = ~new_n7035_ & ~new_n10436_;
  assign new_n10438_ = new_n10435_ & ~new_n10436_;
  assign new_n10439_ = ~new_n10437_ & ~new_n10438_;
  assign new_n10440_ = ~new_n7320_ & new_n10439_;
  assign new_n10441_ = ng826 & ~new_n10440_;
  assign new_n10442_ = ~ng2387 & ~ng826;
  assign n3730 = ~new_n10441_ & ~new_n10442_;
  assign new_n10444_ = ~ng2477 & ~new_n9505_;
  assign new_n10445_ = new_n9505_ & new_n10068_;
  assign n3735 = ~new_n10444_ & ~new_n10445_;
  assign new_n10447_ = ~ng2655 & ~new_n7545_;
  assign new_n10448_ = new_n7545_ & ~new_n10080_;
  assign n3755 = ~new_n10447_ & ~new_n10448_;
  assign new_n10450_ = ng2456 & ng1312;
  assign new_n10451_ = ng1315 & ng2458;
  assign new_n10452_ = ng2454 & ng1309;
  assign new_n10453_ = ~new_n10450_ & ~new_n10451_;
  assign new_n10454_ = ~new_n10452_ & new_n10453_;
  assign new_n10455_ = ng1312 & ng2441;
  assign new_n10456_ = ng1315 & ng2443;
  assign new_n10457_ = ng2439 & ng1309;
  assign new_n10458_ = ~new_n10455_ & ~new_n10456_;
  assign new_n10459_ = ~new_n10457_ & new_n10458_;
  assign new_n10460_ = ~new_n7556_ & ~new_n10454_;
  assign new_n10461_ = new_n10459_ & new_n10460_;
  assign new_n10462_ = new_n7561_ & new_n10461_;
  assign new_n10463_ = ng2426 & ng1312;
  assign new_n10464_ = ng1315 & ng2428;
  assign new_n10465_ = ng2424 & ng1309;
  assign new_n10466_ = ~new_n10463_ & ~new_n10464_;
  assign new_n10467_ = ~new_n10465_ & new_n10466_;
  assign new_n10468_ = new_n7569_ & new_n10459_;
  assign new_n10469_ = new_n10467_ & new_n10468_;
  assign new_n10470_ = ~new_n7556_ & new_n10469_;
  assign new_n10471_ = ng1312 & ng2471;
  assign new_n10472_ = ng1315 & ng2399;
  assign new_n10473_ = ng1309 & ng2469;
  assign new_n10474_ = ~new_n10471_ & ~new_n10472_;
  assign new_n10475_ = ~new_n10473_ & new_n10474_;
  assign new_n10476_ = new_n7556_ & new_n10475_;
  assign new_n10477_ = new_n7569_ & new_n10476_;
  assign new_n10478_ = ~new_n7561_ & new_n10477_;
  assign new_n10479_ = ~new_n10462_ & ~new_n10470_;
  assign new_n10480_ = ~new_n10478_ & new_n10479_;
  assign new_n10481_ = ~new_n7569_ & new_n10459_;
  assign new_n10482_ = ~new_n10467_ & new_n10481_;
  assign new_n10483_ = new_n7561_ & new_n10482_;
  assign new_n10484_ = ~new_n10454_ & ~new_n10467_;
  assign new_n10485_ = ~new_n10459_ & new_n10484_;
  assign new_n10486_ = ~new_n7551_ & new_n10485_;
  assign new_n10487_ = ~new_n7556_ & new_n10454_;
  assign new_n10488_ = new_n10467_ & new_n10487_;
  assign new_n10489_ = ~new_n7561_ & new_n10488_;
  assign new_n10490_ = new_n10480_ & ~new_n10483_;
  assign new_n10491_ = ~new_n10486_ & ~new_n10489_;
  assign new_n10492_ = new_n10490_ & new_n10491_;
  assign new_n10493_ = new_n7561_ & new_n7563_;
  assign new_n10494_ = new_n10454_ & new_n10493_;
  assign new_n10495_ = ~new_n10467_ & new_n10494_;
  assign new_n10496_ = new_n7556_ & new_n7569_;
  assign new_n10497_ = new_n7561_ & new_n10496_;
  assign new_n10498_ = ~new_n10459_ & new_n10497_;
  assign new_n10499_ = ~new_n10475_ & new_n10498_;
  assign new_n10500_ = ~new_n10467_ & new_n10499_;
  assign new_n10501_ = ~new_n7569_ & new_n10467_;
  assign new_n10502_ = ~new_n7561_ & new_n10501_;
  assign new_n10503_ = ~new_n10475_ & new_n10502_;
  assign new_n10504_ = ~new_n10459_ & new_n10503_;
  assign new_n10505_ = ~new_n7561_ & new_n7563_;
  assign new_n10506_ = ~new_n10459_ & new_n10505_;
  assign new_n10507_ = ~new_n10454_ & new_n10506_;
  assign new_n10508_ = new_n10467_ & new_n10507_;
  assign new_n10509_ = ~new_n10495_ & ~new_n10500_;
  assign new_n10510_ = ~new_n10504_ & ~new_n10508_;
  assign new_n10511_ = new_n10509_ & new_n10510_;
  assign new_n10512_ = new_n10492_ & new_n10511_;
  assign new_n10513_ = ng2598 & ~n1651;
  assign new_n10514_ = ng185 & new_n10513_;
  assign new_n10515_ = ng1312 & ng2664;
  assign new_n10516_ = ng1315 & ng2667;
  assign new_n10517_ = ng1309 & ng2661;
  assign new_n10518_ = ~new_n10515_ & ~new_n10516_;
  assign new_n10519_ = ~new_n10517_ & new_n10518_;
  assign new_n10520_ = ~new_n10514_ & new_n10519_;
  assign new_n10521_ = ~new_n9616_ & new_n10512_;
  assign new_n10522_ = new_n10520_ & new_n10521_;
  assign new_n10523_ = ~new_n7569_ & ~new_n10467_;
  assign new_n10524_ = new_n7561_ & new_n10523_;
  assign new_n10525_ = ~new_n10454_ & new_n10524_;
  assign new_n10526_ = ~new_n10459_ & new_n10525_;
  assign new_n10527_ = new_n7569_ & ~new_n10467_;
  assign new_n10528_ = ~new_n7556_ & new_n10527_;
  assign new_n10529_ = ~new_n10475_ & new_n10528_;
  assign new_n10530_ = ~new_n10459_ & new_n10529_;
  assign new_n10531_ = new_n7556_ & new_n10459_;
  assign new_n10532_ = new_n10467_ & new_n10531_;
  assign new_n10533_ = ~new_n7561_ & new_n10532_;
  assign new_n10534_ = new_n7556_ & new_n10467_;
  assign new_n10535_ = new_n7561_ & new_n10534_;
  assign new_n10536_ = ~new_n10454_ & new_n10535_;
  assign new_n10537_ = ~new_n10459_ & new_n10536_;
  assign new_n10538_ = ~new_n10530_ & ~new_n10533_;
  assign new_n10539_ = ~new_n10537_ & new_n10538_;
  assign new_n10540_ = new_n7551_ & ~new_n10467_;
  assign new_n10541_ = ~new_n7561_ & new_n10540_;
  assign new_n10542_ = ~new_n10454_ & new_n10541_;
  assign new_n10543_ = new_n10459_ & new_n10542_;
  assign new_n10544_ = ~new_n10526_ & new_n10539_;
  assign new_n10545_ = ~new_n10543_ & new_n10544_;
  assign new_n10546_ = ~new_n7551_ & ~new_n10475_;
  assign new_n10547_ = new_n10467_ & new_n10546_;
  assign new_n10548_ = ~new_n7561_ & new_n10547_;
  assign new_n10549_ = new_n10454_ & ~new_n10467_;
  assign new_n10550_ = ~new_n10459_ & new_n10549_;
  assign new_n10551_ = ~new_n7556_ & new_n10550_;
  assign new_n10552_ = ~new_n7561_ & new_n10482_;
  assign new_n10553_ = new_n7569_ & new_n10467_;
  assign new_n10554_ = new_n7556_ & new_n10553_;
  assign new_n10555_ = new_n10454_ & new_n10554_;
  assign new_n10556_ = ~new_n10459_ & new_n10555_;
  assign new_n10557_ = ~new_n10551_ & ~new_n10552_;
  assign new_n10558_ = ~new_n10556_ & new_n10557_;
  assign new_n10559_ = new_n7551_ & new_n10475_;
  assign new_n10560_ = ~new_n10467_ & new_n10559_;
  assign new_n10561_ = new_n7561_ & new_n10560_;
  assign new_n10562_ = ~new_n10548_ & new_n10558_;
  assign new_n10563_ = ~new_n10561_ & new_n10562_;
  assign new_n10564_ = new_n10454_ & new_n10467_;
  assign new_n10565_ = ~new_n7551_ & new_n10564_;
  assign new_n10566_ = new_n7569_ & new_n10454_;
  assign new_n10567_ = ~new_n10467_ & new_n10566_;
  assign new_n10568_ = ~new_n7556_ & new_n10567_;
  assign new_n10569_ = ~new_n7569_ & new_n10475_;
  assign new_n10570_ = new_n7561_ & new_n10569_;
  assign new_n10571_ = ~new_n7569_ & ~new_n10454_;
  assign new_n10572_ = new_n10459_ & new_n10571_;
  assign new_n10573_ = ~new_n7561_ & new_n10572_;
  assign new_n10574_ = ~new_n10565_ & ~new_n10568_;
  assign new_n10575_ = ~new_n10570_ & ~new_n10573_;
  assign new_n10576_ = new_n10574_ & new_n10575_;
  assign new_n10577_ = new_n10545_ & new_n10563_;
  assign new_n10578_ = new_n10576_ & new_n10577_;
  assign new_n10579_ = new_n9616_ & ~new_n10578_;
  assign new_n10580_ = new_n10512_ & new_n10579_;
  assign new_n10581_ = ~new_n10522_ & ~new_n10580_;
  assign new_n10582_ = new_n5366_ & new_n10581_;
  assign new_n10583_ = ~new_n5366_ & new_n7540_;
  assign new_n10584_ = ~new_n10582_ & ~new_n10583_;
  assign new_n10585_ = ng1312 & ~new_n10584_;
  assign new_n10586_ = ~ng1312 & ~ng2691;
  assign n3760 = ~new_n10585_ & ~new_n10586_;
  assign new_n10588_ = ng1315 & ~ng2584;
  assign new_n10589_ = ~ng1315 & ~ng2704;
  assign n3770 = ~new_n10588_ & ~new_n10589_;
  assign new_n10591_ = ng2734 & new_n9200_;
  assign new_n10592_ = ng2746 & new_n10591_;
  assign new_n10593_ = ng2740 & new_n10592_;
  assign new_n10594_ = ng2753 & new_n10593_;
  assign new_n10595_ = ng2760 & new_n10594_;
  assign new_n10596_ = ~ng2766 & new_n10595_;
  assign new_n10597_ = ng2766 & ~new_n10595_;
  assign new_n10598_ = ~new_n10596_ & ~new_n10597_;
  assign n3775 = ~new_n8213_ & ~new_n10598_;
  assign new_n10600_ = ~ng2783 & ~new_n7588_;
  assign new_n10601_ = ng2720 & new_n7588_;
  assign n3780 = ~new_n10600_ & ~new_n10601_;
  assign new_n10603_ = ~ng2794 & ~new_n7592_;
  assign new_n10604_ = ng2753 & new_n7592_;
  assign n3785 = ~new_n10603_ & ~new_n10604_;
  assign new_n10606_ = ~ng537 & new_n7609_;
  assign new_n10607_ = ~new_n7605_ & new_n10606_;
  assign new_n10608_ = ~new_n5440_ & ~new_n7627_;
  assign new_n10609_ = ~new_n5302_1_ & ~new_n10608_;
  assign new_n10610_ = ~new_n10608_ & ~new_n10609_;
  assign new_n10611_ = ~new_n5302_1_ & ~new_n10609_;
  assign new_n10612_ = ~new_n10610_ & ~new_n10611_;
  assign new_n10613_ = new_n7609_ & ~new_n10612_;
  assign new_n10614_ = ng499 & new_n10613_;
  assign new_n10615_ = new_n7605_ & new_n10614_;
  assign new_n10616_ = ~new_n10607_ & ~new_n10615_;
  assign new_n10617_ = ~new_n7603_ & new_n10616_;
  assign new_n10618_ = ~new_n5500_ & ~new_n7627_;
  assign new_n10619_ = ~new_n5302_1_ & ~new_n10618_;
  assign new_n10620_ = ~new_n10618_ & ~new_n10619_;
  assign new_n10621_ = ~new_n5302_1_ & ~new_n10619_;
  assign new_n10622_ = ~new_n10620_ & ~new_n10621_;
  assign new_n10623_ = new_n7609_ & ~new_n10622_;
  assign new_n10624_ = ng499 & new_n10623_;
  assign new_n10625_ = new_n7638_ & ~new_n10624_;
  assign new_n10626_ = new_n7603_ & new_n10625_;
  assign n3790 = new_n10617_ | new_n10626_;
  assign new_n10628_ = ng1890 & ~ng1937;
  assign new_n10629_ = ~ng1890 & ~ng1937;
  assign new_n10630_ = ng1905 & new_n10629_;
  assign new_n10631_ = ~new_n10628_ & ~new_n10630_;
  assign new_n10632_ = ~ng1890 & ng1937;
  assign new_n10633_ = ~new_n10630_ & ~new_n10632_;
  assign new_n10634_ = ~ng1939 & ~n2721;
  assign new_n10635_ = ~pg1943 & new_n10634_;
  assign new_n10636_ = ~ng1909 & new_n10635_;
  assign new_n10637_ = ~new_n10633_ & new_n10636_;
  assign new_n10638_ = ng1312 & ~ng2101;
  assign new_n10639_ = ng1315 & ~ng2099;
  assign new_n10640_ = ~ng2100 & ng1309;
  assign new_n10641_ = ~new_n10638_ & ~new_n10639_;
  assign new_n10642_ = ~new_n10640_ & new_n10641_;
  assign new_n10643_ = ng1312 & ~ng2107;
  assign new_n10644_ = ng1315 & ~ng2105;
  assign new_n10645_ = ng1309 & ~ng2106;
  assign new_n10646_ = ~new_n10643_ & ~new_n10644_;
  assign new_n10647_ = ~new_n10645_ & new_n10646_;
  assign new_n10648_ = ng1312 & ~ng2098;
  assign new_n10649_ = ng1315 & ~ng2096;
  assign new_n10650_ = ng1309 & ~ng2097;
  assign new_n10651_ = ~new_n10648_ & ~new_n10649_;
  assign new_n10652_ = ~new_n10650_ & new_n10651_;
  assign new_n10653_ = ng1312 & ~ng2095;
  assign new_n10654_ = ng1315 & ~ng2093;
  assign new_n10655_ = ~ng2094 & ng1309;
  assign new_n10656_ = ~new_n10653_ & ~new_n10654_;
  assign new_n10657_ = ~new_n10655_ & new_n10656_;
  assign new_n10658_ = new_n10642_ & new_n10652_;
  assign new_n10659_ = new_n10657_ & new_n10658_;
  assign new_n10660_ = ~ng2104 & ng1312;
  assign new_n10661_ = ng1315 & ~ng2102;
  assign new_n10662_ = ~ng2103 & ng1309;
  assign new_n10663_ = ~new_n10660_ & ~new_n10661_;
  assign new_n10664_ = ~new_n10662_ & new_n10663_;
  assign new_n10665_ = ~new_n10647_ & new_n10659_;
  assign new_n10666_ = ~new_n10664_ & new_n10665_;
  assign new_n10667_ = ng1312 & ~ng2119;
  assign new_n10668_ = ng1315 & ~ng2117;
  assign new_n10669_ = ng1309 & ~ng2118;
  assign new_n10670_ = ~new_n10667_ & ~new_n10668_;
  assign new_n10671_ = ~new_n10669_ & new_n10670_;
  assign new_n10672_ = ng1312 & ~ng2092;
  assign new_n10673_ = ~ng2090 & ng1315;
  assign new_n10674_ = ~ng2091 & ng1309;
  assign new_n10675_ = ~new_n10672_ & ~new_n10673_;
  assign new_n10676_ = ~new_n10674_ & new_n10675_;
  assign new_n10677_ = ng1312 & ~ng2083;
  assign new_n10678_ = ng1315 & ~ng2081;
  assign new_n10679_ = ~ng2082 & ng1309;
  assign new_n10680_ = ~new_n10677_ & ~new_n10678_;
  assign new_n10681_ = ~new_n10679_ & new_n10680_;
  assign new_n10682_ = ng1312 & ~ng2086;
  assign new_n10683_ = ng1315 & ~ng2084;
  assign new_n10684_ = ng1309 & ~ng2085;
  assign new_n10685_ = ~new_n10682_ & ~new_n10683_;
  assign new_n10686_ = ~new_n10684_ & new_n10685_;
  assign new_n10687_ = ~ng2080 & ng1312;
  assign new_n10688_ = ~ng2078 & ng1315;
  assign new_n10689_ = ~ng2079 & ng1309;
  assign new_n10690_ = ~new_n10687_ & ~new_n10688_;
  assign new_n10691_ = ~new_n10689_ & new_n10690_;
  assign new_n10692_ = ~new_n10681_ & ~new_n10686_;
  assign new_n10693_ = new_n10691_ & new_n10692_;
  assign new_n10694_ = ng1312 & ~ng2089;
  assign new_n10695_ = ng1315 & ~ng2087;
  assign new_n10696_ = ng1309 & ~ng2088;
  assign new_n10697_ = ~new_n10694_ & ~new_n10695_;
  assign new_n10698_ = ~new_n10696_ & new_n10697_;
  assign new_n10699_ = new_n10676_ & new_n10693_;
  assign new_n10700_ = ~new_n10698_ & new_n10699_;
  assign new_n10701_ = ~ng2113 & ng1312;
  assign new_n10702_ = ng1315 & ~ng2111;
  assign new_n10703_ = ~ng2112 & ng1309;
  assign new_n10704_ = ~new_n10701_ & ~new_n10702_;
  assign new_n10705_ = ~new_n10703_ & new_n10704_;
  assign new_n10706_ = new_n10666_ & ~new_n10671_;
  assign new_n10707_ = new_n10700_ & ~new_n10705_;
  assign new_n10708_ = new_n10706_ & new_n10707_;
  assign new_n10709_ = ~new_n10642_ & ~new_n10708_;
  assign new_n10710_ = ~new_n6785_ & ~new_n10709_;
  assign new_n10711_ = ~new_n10709_ & ~new_n10710_;
  assign new_n10712_ = ~new_n6785_ & ~new_n10710_;
  assign new_n10713_ = ~new_n10711_ & ~new_n10712_;
  assign new_n10714_ = new_n10635_ & ~new_n10713_;
  assign new_n10715_ = ng1880 & new_n10714_;
  assign new_n10716_ = new_n10633_ & new_n10715_;
  assign new_n10717_ = ~new_n10637_ & ~new_n10716_;
  assign new_n10718_ = ~new_n10631_ & new_n10717_;
  assign new_n10719_ = new_n10631_ & ~new_n10633_;
  assign new_n10720_ = ng1312 & ~ng2116;
  assign new_n10721_ = ng1315 & ~ng2114;
  assign new_n10722_ = ng1309 & ~ng2115;
  assign new_n10723_ = ~new_n10720_ & ~new_n10721_;
  assign new_n10724_ = ~new_n10722_ & new_n10723_;
  assign new_n10725_ = ~new_n10708_ & new_n10724_;
  assign new_n10726_ = ng1880 & ~new_n10725_;
  assign new_n10727_ = new_n10635_ & new_n10726_;
  assign new_n10728_ = new_n10719_ & ~new_n10727_;
  assign new_n10729_ = new_n10631_ & new_n10728_;
  assign n3795 = new_n10718_ | new_n10729_;
  assign new_n10731_ = ~ng2631 & ng2584;
  assign new_n10732_ = ~ng2631 & ~ng2584;
  assign new_n10733_ = ng2599 & new_n10732_;
  assign new_n10734_ = ~new_n10731_ & ~new_n10733_;
  assign new_n10735_ = ng2631 & ~ng2584;
  assign new_n10736_ = ~new_n10733_ & ~new_n10735_;
  assign new_n10737_ = ~ng2633 & ~n4713;
  assign new_n10738_ = ~pg2637 & new_n10737_;
  assign new_n10739_ = ~ng2605 & new_n10738_;
  assign new_n10740_ = ~new_n10736_ & new_n10739_;
  assign new_n10741_ = new_n8295_ & new_n8304_;
  assign new_n10742_ = new_n8313_ & new_n10741_;
  assign new_n10743_ = ~new_n8286_ & new_n10742_;
  assign new_n10744_ = ~new_n8324_ & new_n10743_;
  assign new_n10745_ = ng1312 & ~ng2813;
  assign new_n10746_ = ng1315 & ~ng2811;
  assign new_n10747_ = ~ng2812 & ng1309;
  assign new_n10748_ = ~new_n10745_ & ~new_n10746_;
  assign new_n10749_ = ~new_n10747_ & new_n10748_;
  assign new_n10750_ = ~new_n8246_ & ~new_n8255_;
  assign new_n10751_ = new_n8264_ & new_n10750_;
  assign new_n10752_ = new_n8237_ & new_n10751_;
  assign new_n10753_ = ~new_n8275_ & new_n10752_;
  assign new_n10754_ = new_n10744_ & ~new_n10749_;
  assign new_n10755_ = ~new_n8336_ & new_n10753_;
  assign new_n10756_ = new_n10754_ & new_n10755_;
  assign new_n10757_ = ~new_n8313_ & ~new_n10756_;
  assign new_n10758_ = ~new_n7529_ & ~new_n10757_;
  assign new_n10759_ = ~new_n10757_ & ~new_n10758_;
  assign new_n10760_ = ~new_n7529_ & ~new_n10758_;
  assign new_n10761_ = ~new_n10759_ & ~new_n10760_;
  assign new_n10762_ = new_n10738_ & ~new_n10761_;
  assign new_n10763_ = ng2574 & new_n10762_;
  assign new_n10764_ = new_n10736_ & new_n10763_;
  assign new_n10765_ = ~new_n10740_ & ~new_n10764_;
  assign new_n10766_ = ~new_n10734_ & new_n10765_;
  assign new_n10767_ = new_n10734_ & ~new_n10736_;
  assign new_n10768_ = ~ng2810 & ng1312;
  assign new_n10769_ = ng1315 & ~ng2808;
  assign new_n10770_ = ~ng2809 & ng1309;
  assign new_n10771_ = ~new_n10768_ & ~new_n10769_;
  assign new_n10772_ = ~new_n10770_ & new_n10771_;
  assign new_n10773_ = ~new_n10756_ & new_n10772_;
  assign new_n10774_ = ng2574 & ~new_n10773_;
  assign new_n10775_ = new_n10738_ & ~new_n10774_;
  assign new_n10776_ = new_n10767_ & ~new_n10775_;
  assign new_n10777_ = new_n10734_ & new_n10776_;
  assign n3800 = new_n10766_ | new_n10777_;
  assign new_n10779_ = ng3080 & new_n5362_;
  assign new_n10780_ = ~pg3234 & ~new_n10779_;
  assign new_n10781_ = ng3080 & ng2993;
  assign new_n10782_ = ng2998 & new_n10781_;
  assign new_n10783_ = ng3006 & new_n10782_;
  assign new_n10784_ = ng3002 & new_n10783_;
  assign new_n10785_ = ~ng3013 & new_n10784_;
  assign new_n10786_ = ng3013 & ~new_n10784_;
  assign new_n10787_ = ~new_n10785_ & ~new_n10786_;
  assign n3805 = new_n10780_ & ~new_n10787_;
  assign new_n10789_ = ~ng3063 & ng2987;
  assign new_n10790_ = ~ng3044 & ~ng2987;
  assign n3810 = ~new_n10789_ & ~new_n10790_;
  assign new_n10792_ = ~ng3072 & ng2987;
  assign new_n10793_ = ~ng3053 & ~ng2987;
  assign n3815 = ~new_n10792_ & ~new_n10793_;
  assign new_n10795_ = ~ng2896 & new_n9236_;
  assign new_n10796_ = ng2896 & ~new_n9236_;
  assign new_n10797_ = ~new_n10795_ & ~new_n10796_;
  assign n3820 = new_n9234_ & ~new_n10797_;
  assign new_n10799_ = ~ng131 & ~new_n4777_1_;
  assign new_n10800_ = ng97 & new_n4777_1_;
  assign n3825 = ~new_n10799_ & ~new_n10800_;
  assign new_n10802_ = ~ng146 & ~new_n4777_1_;
  assign new_n10803_ = ng109 & new_n4777_1_;
  assign n3830 = ~new_n10802_ & ~new_n10803_;
  assign new_n10805_ = ~ng156 & ~new_n4773_;
  assign new_n10806_ = ng125 & new_n4773_;
  assign n3835 = ~new_n10805_ & ~new_n10806_;
  assign new_n10808_ = ~ng168 & ~new_n8121_;
  assign new_n10809_ = ~ng117 & ~ng121;
  assign new_n10810_ = ng125 & new_n10809_;
  assign new_n10811_ = ng113 & new_n10810_;
  assign new_n10812_ = new_n8121_ & ~new_n10811_;
  assign n3840 = ~new_n10808_ & ~new_n10812_;
  assign new_n10814_ = ng101 & ~new_n5083_;
  assign new_n10815_ = ~new_n8915_ & ~new_n10814_;
  assign new_n10816_ = ~new_n5082_1_ & new_n10815_;
  assign new_n10817_ = ~new_n4815_ & ~new_n5095_;
  assign new_n10818_ = new_n4815_ & new_n5095_;
  assign new_n10819_ = ~new_n10817_ & ~new_n10818_;
  assign new_n10820_ = new_n5082_1_ & new_n10819_;
  assign new_n10821_ = ~new_n10816_ & ~new_n10820_;
  assign new_n10822_ = ng826 & ~new_n10821_;
  assign new_n10823_ = ~ng231 & ~ng826;
  assign n3845 = ~new_n10822_ & ~new_n10823_;
  assign new_n10825_ = ng826 & ~new_n10314_;
  assign new_n10826_ = ~ng204 & ~ng826;
  assign n3850 = ~new_n10825_ & ~new_n10826_;
  assign new_n10828_ = n4167 & ~new_n5182_1_;
  assign new_n10829_ = ~n4167 & new_n5190_;
  assign new_n10830_ = ~new_n10828_ & ~new_n10829_;
  assign new_n10831_ = new_n5187_1_ & ~new_n10830_;
  assign new_n10832_ = ~new_n5168_ & new_n10831_;
  assign new_n10833_ = ng2384 & new_n10832_;
  assign new_n10834_ = new_n5168_ & ~new_n10830_;
  assign new_n10835_ = ng2384 & new_n10834_;
  assign new_n10836_ = ~new_n10833_ & ~new_n10835_;
  assign new_n10837_ = ng826 & ~new_n10836_;
  assign new_n10838_ = ~ng427 & ~new_n10837_;
  assign new_n10839_ = new_n10833_ & new_n10837_;
  assign n3855 = ~new_n10838_ & ~new_n10839_;
  assign new_n10841_ = ng823 & new_n10324_;
  assign new_n10842_ = ~ng323 & ~new_n10841_;
  assign new_n10843_ = new_n10331_ & new_n10841_;
  assign n3860 = ~new_n10842_ & ~new_n10843_;
  assign new_n10845_ = ~ng582 & ~new_n8959_;
  assign new_n10846_ = ~pg3229 & new_n5323_;
  assign new_n10847_ = new_n5325_ & new_n10846_;
  assign new_n10848_ = ~new_n5326_1_ & ~new_n10847_;
  assign new_n10849_ = ~new_n5318_ & ~new_n5323_;
  assign new_n10850_ = ~pg3229 & new_n10849_;
  assign new_n10851_ = ~new_n5318_ & new_n5323_;
  assign new_n10852_ = pg3229 & new_n10851_;
  assign new_n10853_ = ~new_n10850_ & ~new_n10852_;
  assign new_n10854_ = new_n10848_ & new_n10853_;
  assign new_n10855_ = new_n8959_ & ~new_n10854_;
  assign n3878 = ~new_n10845_ & ~new_n10855_;
  assign new_n10857_ = ng1309 & ~new_n10337_;
  assign new_n10858_ = ~ng596 & ~ng1309;
  assign n3883 = ~new_n10857_ & ~new_n10858_;
  assign new_n10860_ = ~ng707 & ~new_n5399_;
  assign new_n10861_ = ng646 & new_n5399_;
  assign n3898 = ~new_n10860_ & ~new_n10861_;
  assign new_n10863_ = ~ng831 & ~new_n4777_1_;
  assign new_n10864_ = ng793 & new_n4777_1_;
  assign n3903 = ~new_n10863_ & ~new_n10864_;
  assign new_n10866_ = ~ng850 & ~new_n4773_;
  assign new_n10867_ = new_n4773_ & ~new_n5652_;
  assign n3908 = ~new_n10866_ & ~new_n10867_;
  assign new_n10869_ = ~ng862 & ~new_n8121_;
  assign new_n10870_ = ng785 & new_n8121_;
  assign n3913 = ~new_n10869_ & ~new_n10870_;
  assign new_n10872_ = ng853 & ~new_n10359_;
  assign new_n10873_ = ~ng897 & ~ng853;
  assign n3918 = ~new_n10872_ & ~new_n10873_;
  assign new_n10875_ = ng813 & ~new_n5839_;
  assign new_n10876_ = ~new_n5838_1_ & ~new_n10875_;
  assign new_n10877_ = ~new_n5897_ & new_n8478_;
  assign new_n10878_ = new_n5588_ & new_n10877_;
  assign new_n10879_ = ~new_n5588_ & ~new_n10877_;
  assign new_n10880_ = ~new_n10878_ & ~new_n10879_;
  assign new_n10881_ = new_n5838_1_ & new_n10880_;
  assign new_n10882_ = ~new_n10876_ & ~new_n10881_;
  assign new_n10883_ = ng853 & ~new_n10882_;
  assign new_n10884_ = ~ng951 & ~ng853;
  assign n3923 = ~new_n10883_ & ~new_n10884_;
  assign new_n10886_ = ~new_n5366_ & ~new_n6173_;
  assign new_n10887_ = ng1309 & ~new_n10886_;
  assign new_n10888_ = ~ng1273 & ~ng1309;
  assign n3949 = ~new_n10887_ & ~new_n10888_;
  assign new_n10890_ = ~pg3229 & ~ng992;
  assign new_n10891_ = pg3229 & ng978;
  assign n3954 = ~new_n10890_ & ~new_n10891_;
  assign new_n10893_ = ng1339 & ~new_n6244_1_;
  assign new_n10894_ = ~ng1339 & new_n6244_1_;
  assign new_n10895_ = ~new_n10893_ & ~new_n10894_;
  assign n3959 = ~new_n6241_ & ~new_n10895_;
  assign new_n10897_ = ~ng1387 & ~new_n6263_;
  assign new_n10898_ = ng1319 & new_n6263_;
  assign n3964 = ~new_n10897_ & ~new_n10898_;
  assign new_n10900_ = ~ng1396 & ~new_n6263_;
  assign new_n10901_ = ng1346 & new_n6263_;
  assign n3969 = ~new_n10900_ & ~new_n10901_;
  assign new_n10903_ = ~ng1561 & ~new_n6278_;
  assign new_n10904_ = new_n6278_ & new_n6678_;
  assign n3974 = ~new_n10903_ & ~new_n10904_;
  assign new_n10906_ = ng823 & ~new_n10390_;
  assign new_n10907_ = ~ng1579 & ~ng823;
  assign n3979 = ~new_n10906_ & ~new_n10907_;
  assign new_n10909_ = ng853 & ~new_n10400_;
  assign new_n10910_ = ~ng1600 & ~ng853;
  assign n3984 = ~new_n10909_ & ~new_n10910_;
  assign new_n10912_ = ~new_n6395_ & ~new_n6587_;
  assign new_n10913_ = ~new_n10383_ & ~new_n10912_;
  assign new_n10914_ = ~new_n6586_ & new_n10913_;
  assign new_n10915_ = new_n6301_ & ~new_n6360_;
  assign new_n10916_ = ~new_n6301_ & new_n6360_;
  assign new_n10917_ = ~new_n10915_ & ~new_n10916_;
  assign new_n10918_ = new_n6301_ & ~new_n6331_1_;
  assign new_n10919_ = ~new_n6301_ & new_n6331_1_;
  assign new_n10920_ = ~new_n10918_ & ~new_n10919_;
  assign new_n10921_ = ~new_n6592_ & ~new_n10920_;
  assign new_n10922_ = new_n6600_1_ & new_n6614_1_;
  assign new_n10923_ = new_n6607_ & new_n10921_;
  assign new_n10924_ = new_n10922_ & new_n10923_;
  assign new_n10925_ = ~new_n10917_ & new_n10924_;
  assign new_n10926_ = new_n6326_ & new_n10925_;
  assign new_n10927_ = ~new_n6326_ & ~new_n10925_;
  assign new_n10928_ = ~new_n10926_ & ~new_n10927_;
  assign new_n10929_ = new_n6586_ & new_n10928_;
  assign new_n10930_ = ~new_n10914_ & ~new_n10929_;
  assign new_n10931_ = ng853 & ~new_n10930_;
  assign new_n10932_ = ~ng1654 & ~ng853;
  assign n3989 = ~new_n10931_ & ~new_n10932_;
  assign new_n10934_ = ~ng2221 & ~new_n5517_1_;
  assign new_n10935_ = ng2180 & new_n5517_1_;
  assign n4011 = ~new_n10934_ & ~new_n10935_;
  assign new_n10937_ = ~ng2230 & ~new_n5517_1_;
  assign new_n10938_ = ng2195 & new_n5517_1_;
  assign n4016 = ~new_n10937_ & ~new_n10938_;
  assign new_n10940_ = ng823 & ~new_n10047_;
  assign new_n10941_ = ~ng2264 & ~ng823;
  assign n4021 = ~new_n10940_ & ~new_n10941_;
  assign new_n10943_ = ng853 & ~new_n10425_;
  assign new_n10944_ = ~ng2501 & ~new_n10943_;
  assign new_n10945_ = new_n10422_ & new_n10943_;
  assign n4026 = ~new_n10944_ & ~new_n10945_;
  assign new_n10947_ = ng853 & ~new_n7514_;
  assign new_n10948_ = ~ng2522 & ~new_n10947_;
  assign new_n10949_ = new_n7507_ & new_n10947_;
  assign n4031 = ~new_n10948_ & ~new_n10949_;
  assign new_n10951_ = ~ng2659 & ~new_n9196_;
  assign new_n10952_ = ~pg3229 & ~new_n7561_;
  assign new_n10953_ = new_n10496_ & new_n10952_;
  assign new_n10954_ = pg3229 & new_n7561_;
  assign new_n10955_ = new_n10496_ & new_n10954_;
  assign new_n10956_ = ~new_n10953_ & ~new_n10955_;
  assign new_n10957_ = new_n9196_ & ~new_n10956_;
  assign n4053 = ~new_n10951_ & ~new_n10957_;
  assign new_n10959_ = ng1309 & ~new_n10584_;
  assign new_n10960_ = ~ng2688 & ~ng1309;
  assign n4058 = ~new_n10959_ & ~new_n10960_;
  assign new_n10962_ = ~ng2773 & ~new_n7592_;
  assign new_n10963_ = ng2714 & new_n7592_;
  assign n4073 = ~new_n10962_ & ~new_n10963_;
  assign new_n10965_ = ~ng2782 & ~new_n7592_;
  assign new_n10966_ = ng2720 & new_n7592_;
  assign n4078 = ~new_n10965_ & ~new_n10966_;
  assign new_n10968_ = ~ng2804 & ~new_n8213_;
  assign new_n10969_ = ~new_n7540_ & new_n8213_;
  assign n4083 = ~new_n10968_ & ~new_n10969_;
  assign new_n10971_ = new_n10278_ & new_n10624_;
  assign new_n10972_ = new_n10278_ & ~new_n10971_;
  assign new_n10973_ = new_n10624_ & ~new_n10971_;
  assign new_n10974_ = ~new_n10972_ & ~new_n10973_;
  assign new_n10975_ = ng557 & ~new_n10974_;
  assign new_n10976_ = new_n7634_ & new_n8349_;
  assign new_n10977_ = new_n8349_ & ~new_n10976_;
  assign new_n10978_ = new_n7634_ & ~new_n10976_;
  assign new_n10979_ = ~new_n10977_ & ~new_n10978_;
  assign new_n10980_ = new_n8895_ & new_n9222_;
  assign new_n10981_ = new_n9222_ & ~new_n10980_;
  assign new_n10982_ = new_n8895_ & ~new_n10980_;
  assign new_n10983_ = ~new_n10981_ & ~new_n10982_;
  assign new_n10984_ = ~new_n10979_ & ~new_n10983_;
  assign new_n10985_ = ~new_n10979_ & ~new_n10984_;
  assign new_n10986_ = ~new_n10983_ & ~new_n10984_;
  assign new_n10987_ = ~new_n10985_ & ~new_n10986_;
  assign new_n10988_ = new_n9643_ & new_n9871_;
  assign new_n10989_ = new_n9871_ & ~new_n10988_;
  assign new_n10990_ = new_n9643_ & ~new_n10988_;
  assign new_n10991_ = ~new_n10989_ & ~new_n10990_;
  assign new_n10992_ = new_n10268_ & new_n10614_;
  assign new_n10993_ = new_n10268_ & ~new_n10992_;
  assign new_n10994_ = new_n10614_ & ~new_n10992_;
  assign new_n10995_ = ~new_n10993_ & ~new_n10994_;
  assign new_n10996_ = ~new_n10991_ & ~new_n10995_;
  assign new_n10997_ = ~new_n10991_ & ~new_n10996_;
  assign new_n10998_ = ~new_n10995_ & ~new_n10996_;
  assign new_n10999_ = ~new_n10997_ & ~new_n10998_;
  assign new_n11000_ = ~new_n10987_ & ~new_n10999_;
  assign new_n11001_ = ~new_n10987_ & ~new_n11000_;
  assign new_n11002_ = ~new_n10999_ & ~new_n11000_;
  assign new_n11003_ = ~new_n11001_ & ~new_n11002_;
  assign new_n11004_ = ng510 & ~new_n11003_;
  assign new_n11005_ = ~pg3229 & ~ng541;
  assign new_n11006_ = pg3229 & ~ng538;
  assign new_n11007_ = ~new_n11005_ & ~new_n11006_;
  assign new_n11008_ = new_n7609_ & new_n11007_;
  assign new_n11009_ = ~new_n7603_ & ~new_n7605_;
  assign new_n11010_ = new_n11008_ & new_n11009_;
  assign new_n11011_ = new_n7601_ & new_n11010_;
  assign new_n11012_ = ~new_n10975_ & ~new_n11004_;
  assign n4088 = new_n11011_ | ~new_n11012_;
  assign new_n11014_ = ~ng1245 & ~n1448;
  assign new_n11015_ = ~pg1249 & new_n11014_;
  assign new_n11016_ = new_n8651_ & new_n8660_;
  assign new_n11017_ = new_n8669_ & new_n11016_;
  assign new_n11018_ = ~new_n8642_ & new_n11017_;
  assign new_n11019_ = ~new_n8680_ & new_n11018_;
  assign new_n11020_ = ~ng1425 & ng1312;
  assign new_n11021_ = ~ng1423 & ng1315;
  assign new_n11022_ = ~ng1424 & ng1309;
  assign new_n11023_ = ~new_n11020_ & ~new_n11021_;
  assign new_n11024_ = ~new_n11022_ & new_n11023_;
  assign new_n11025_ = ~new_n8602_ & ~new_n8611_;
  assign new_n11026_ = new_n8620_ & new_n11025_;
  assign new_n11027_ = new_n8593_ & new_n11026_;
  assign new_n11028_ = ~new_n8631_ & new_n11027_;
  assign new_n11029_ = new_n11019_ & ~new_n11024_;
  assign new_n11030_ = ~new_n8692_ & new_n11028_;
  assign new_n11031_ = new_n11029_ & new_n11030_;
  assign new_n11032_ = ~new_n8642_ & ~new_n11031_;
  assign new_n11033_ = ~new_n6033_ & ~new_n11032_;
  assign new_n11034_ = ~new_n11032_ & ~new_n11033_;
  assign new_n11035_ = ~new_n6033_ & ~new_n11033_;
  assign new_n11036_ = ~new_n11034_ & ~new_n11035_;
  assign new_n11037_ = new_n11015_ & ~new_n11036_;
  assign new_n11038_ = ng1186 & new_n11037_;
  assign new_n11039_ = ~new_n8680_ & ~new_n11031_;
  assign new_n11040_ = ~new_n6044_ & ~new_n11039_;
  assign new_n11041_ = ~new_n11039_ & ~new_n11040_;
  assign new_n11042_ = ~new_n6044_ & ~new_n11040_;
  assign new_n11043_ = ~new_n11041_ & ~new_n11042_;
  assign new_n11044_ = new_n11015_ & ~new_n11043_;
  assign new_n11045_ = ng1186 & new_n11044_;
  assign new_n11046_ = new_n11038_ & new_n11045_;
  assign new_n11047_ = new_n11038_ & ~new_n11046_;
  assign new_n11048_ = new_n11045_ & ~new_n11046_;
  assign new_n11049_ = ~new_n11047_ & ~new_n11048_;
  assign new_n11050_ = ng1243 & ~new_n11049_;
  assign new_n11051_ = ~new_n8660_ & ~new_n11031_;
  assign new_n11052_ = ~new_n6033_ & ~new_n11051_;
  assign new_n11053_ = ~new_n11051_ & ~new_n11052_;
  assign new_n11054_ = ~new_n6033_ & ~new_n11052_;
  assign new_n11055_ = ~new_n11053_ & ~new_n11054_;
  assign new_n11056_ = new_n11015_ & ~new_n11055_;
  assign new_n11057_ = ng1186 & new_n11056_;
  assign new_n11058_ = ~new_n8651_ & ~new_n11031_;
  assign new_n11059_ = ~new_n6044_ & ~new_n11058_;
  assign new_n11060_ = ~new_n11058_ & ~new_n11059_;
  assign new_n11061_ = ~new_n6044_ & ~new_n11059_;
  assign new_n11062_ = ~new_n11060_ & ~new_n11061_;
  assign new_n11063_ = new_n11015_ & ~new_n11062_;
  assign new_n11064_ = ng1186 & new_n11063_;
  assign new_n11065_ = new_n11057_ & new_n11064_;
  assign new_n11066_ = new_n11057_ & ~new_n11065_;
  assign new_n11067_ = new_n11064_ & ~new_n11065_;
  assign new_n11068_ = ~new_n11066_ & ~new_n11067_;
  assign new_n11069_ = ~new_n8669_ & ~new_n11031_;
  assign new_n11070_ = ~new_n6033_ & ~new_n11069_;
  assign new_n11071_ = ~new_n11069_ & ~new_n11070_;
  assign new_n11072_ = ~new_n6033_ & ~new_n11070_;
  assign new_n11073_ = ~new_n11071_ & ~new_n11072_;
  assign new_n11074_ = new_n11015_ & ~new_n11073_;
  assign new_n11075_ = ng1186 & new_n11074_;
  assign new_n11076_ = ~new_n8593_ & ~new_n11031_;
  assign new_n11077_ = ~new_n6044_ & ~new_n11076_;
  assign new_n11078_ = ~new_n11076_ & ~new_n11077_;
  assign new_n11079_ = ~new_n6044_ & ~new_n11077_;
  assign new_n11080_ = ~new_n11078_ & ~new_n11079_;
  assign new_n11081_ = new_n11015_ & ~new_n11080_;
  assign new_n11082_ = ng1186 & new_n11081_;
  assign new_n11083_ = new_n11075_ & new_n11082_;
  assign new_n11084_ = new_n11075_ & ~new_n11083_;
  assign new_n11085_ = new_n11082_ & ~new_n11083_;
  assign new_n11086_ = ~new_n11084_ & ~new_n11085_;
  assign new_n11087_ = ~new_n11068_ & ~new_n11086_;
  assign new_n11088_ = ~new_n11068_ & ~new_n11087_;
  assign new_n11089_ = ~new_n11086_ & ~new_n11087_;
  assign new_n11090_ = ~new_n11088_ & ~new_n11089_;
  assign new_n11091_ = ~new_n8631_ & ~new_n11031_;
  assign new_n11092_ = ~new_n6033_ & ~new_n11091_;
  assign new_n11093_ = ~new_n11091_ & ~new_n11092_;
  assign new_n11094_ = ~new_n6033_ & ~new_n11092_;
  assign new_n11095_ = ~new_n11093_ & ~new_n11094_;
  assign new_n11096_ = new_n11015_ & ~new_n11095_;
  assign new_n11097_ = ng1186 & new_n11096_;
  assign new_n11098_ = ~new_n8611_ & ~new_n11031_;
  assign new_n11099_ = ~new_n6044_ & ~new_n11098_;
  assign new_n11100_ = ~new_n11098_ & ~new_n11099_;
  assign new_n11101_ = ~new_n6044_ & ~new_n11099_;
  assign new_n11102_ = ~new_n11100_ & ~new_n11101_;
  assign new_n11103_ = new_n11015_ & ~new_n11102_;
  assign new_n11104_ = ng1186 & new_n11103_;
  assign new_n11105_ = new_n11097_ & new_n11104_;
  assign new_n11106_ = new_n11097_ & ~new_n11105_;
  assign new_n11107_ = new_n11104_ & ~new_n11105_;
  assign new_n11108_ = ~new_n11106_ & ~new_n11107_;
  assign new_n11109_ = ~new_n8602_ & ~new_n11031_;
  assign new_n11110_ = ~new_n6033_ & ~new_n11109_;
  assign new_n11111_ = ~new_n11109_ & ~new_n11110_;
  assign new_n11112_ = ~new_n6033_ & ~new_n11110_;
  assign new_n11113_ = ~new_n11111_ & ~new_n11112_;
  assign new_n11114_ = new_n11015_ & ~new_n11113_;
  assign new_n11115_ = ng1186 & new_n11114_;
  assign new_n11116_ = ~new_n8620_ & ~new_n11031_;
  assign new_n11117_ = ~new_n6044_ & ~new_n11116_;
  assign new_n11118_ = ~new_n11116_ & ~new_n11117_;
  assign new_n11119_ = ~new_n6044_ & ~new_n11117_;
  assign new_n11120_ = ~new_n11118_ & ~new_n11119_;
  assign new_n11121_ = new_n11015_ & ~new_n11120_;
  assign new_n11122_ = ng1186 & new_n11121_;
  assign new_n11123_ = new_n11115_ & new_n11122_;
  assign new_n11124_ = new_n11115_ & ~new_n11123_;
  assign new_n11125_ = new_n11122_ & ~new_n11123_;
  assign new_n11126_ = ~new_n11124_ & ~new_n11125_;
  assign new_n11127_ = ~new_n11108_ & ~new_n11126_;
  assign new_n11128_ = ~new_n11108_ & ~new_n11127_;
  assign new_n11129_ = ~new_n11126_ & ~new_n11127_;
  assign new_n11130_ = ~new_n11128_ & ~new_n11129_;
  assign new_n11131_ = ~new_n11090_ & ~new_n11130_;
  assign new_n11132_ = ~new_n11090_ & ~new_n11131_;
  assign new_n11133_ = ~new_n11130_ & ~new_n11131_;
  assign new_n11134_ = ~new_n11132_ & ~new_n11133_;
  assign new_n11135_ = ng1196 & ~new_n11134_;
  assign new_n11136_ = ~ng1196 & ~ng1243;
  assign new_n11137_ = ng1211 & new_n11136_;
  assign new_n11138_ = ~ng1196 & ng1243;
  assign new_n11139_ = ~new_n11137_ & ~new_n11138_;
  assign new_n11140_ = ng1196 & ~ng1243;
  assign new_n11141_ = ~new_n11137_ & ~new_n11140_;
  assign new_n11142_ = ~pg3229 & ~ng1227;
  assign new_n11143_ = pg3229 & ~ng1224;
  assign new_n11144_ = ~new_n11142_ & ~new_n11143_;
  assign new_n11145_ = new_n11015_ & new_n11144_;
  assign new_n11146_ = ~new_n11139_ & ~new_n11141_;
  assign new_n11147_ = new_n11145_ & new_n11146_;
  assign new_n11148_ = new_n11136_ & new_n11147_;
  assign new_n11149_ = ~new_n11050_ & ~new_n11135_;
  assign n4093 = new_n11148_ | ~new_n11149_;
  assign new_n11151_ = ~ng2606 & new_n10738_;
  assign new_n11152_ = ~new_n10736_ & new_n11151_;
  assign new_n11153_ = ~new_n8237_ & ~new_n10756_;
  assign new_n11154_ = ~new_n7540_ & ~new_n11153_;
  assign new_n11155_ = ~new_n11153_ & ~new_n11154_;
  assign new_n11156_ = ~new_n7540_ & ~new_n11154_;
  assign new_n11157_ = ~new_n11155_ & ~new_n11156_;
  assign new_n11158_ = new_n10738_ & ~new_n11157_;
  assign new_n11159_ = ng2574 & new_n11158_;
  assign new_n11160_ = new_n10736_ & new_n11159_;
  assign new_n11161_ = ~new_n11152_ & ~new_n11160_;
  assign new_n11162_ = ~new_n10734_ & new_n11161_;
  assign new_n11163_ = new_n10738_ & new_n10774_;
  assign new_n11164_ = new_n10767_ & ~new_n11163_;
  assign new_n11165_ = new_n10734_ & new_n11164_;
  assign n4098 = new_n11162_ | new_n11165_;
  assign new_n11167_ = ng3002 & ~new_n10783_;
  assign new_n11168_ = ~ng3002 & new_n10783_;
  assign new_n11169_ = ~new_n11167_ & ~new_n11168_;
  assign n4103 = new_n10780_ & ~new_n11169_;
  assign new_n11171_ = ~ng3064 & ng2987;
  assign new_n11172_ = ~ng3045 & ~ng2987;
  assign n4108 = ~new_n11171_ & ~new_n11172_;
  assign new_n11174_ = ~ng3071 & ng2987;
  assign new_n11175_ = ~ng3052 & ~ng2987;
  assign n4113 = ~new_n11174_ & ~new_n11175_;
  assign new_n11177_ = ng2892 & ~new_n9237_;
  assign new_n11178_ = ~ng2892 & new_n9237_;
  assign new_n11179_ = ~new_n11177_ & ~new_n11178_;
  assign n4118 = new_n9234_ & ~new_n11179_;
  assign new_n11181_ = ~ng129 & ~new_n4773_;
  assign new_n11182_ = ng97 & new_n4773_;
  assign n4123 = ~new_n11181_ & ~new_n11182_;
  assign new_n11184_ = ~ng149 & ~new_n4777_1_;
  assign new_n11185_ = ng113 & new_n4777_1_;
  assign n4128 = ~new_n11184_ & ~new_n11185_;
  assign new_n11187_ = ~ng153 & ~new_n4773_;
  assign new_n11188_ = ng121 & new_n4773_;
  assign n4133 = ~new_n11187_ & ~new_n11188_;
  assign new_n11190_ = ~ng170 & ~new_n6278_;
  assign new_n11191_ = new_n6278_ & ~new_n10811_;
  assign n4138 = ~new_n11190_ & ~new_n11191_;
  assign new_n11193_ = ng823 & ~new_n10821_;
  assign new_n11194_ = ~ng234 & ~ng823;
  assign n4143 = ~new_n11193_ & ~new_n11194_;
  assign new_n11196_ = ng826 & ~new_n9271_;
  assign new_n11197_ = ~ng249 & ~ng826;
  assign n4148 = ~new_n11196_ & ~new_n11197_;
  assign new_n11199_ = ng823 & ~new_n10836_;
  assign new_n11200_ = ~ng428 & ~new_n11199_;
  assign new_n11201_ = new_n10833_ & new_n11199_;
  assign n4153 = ~new_n11200_ & ~new_n11201_;
  assign new_n11203_ = ~new_n4785_ & new_n4795_;
  assign new_n11204_ = new_n4790_ & new_n11203_;
  assign new_n11205_ = new_n4785_ & ~new_n4795_;
  assign new_n11206_ = ~new_n4955_ & ~new_n11205_;
  assign new_n11207_ = ~new_n4790_ & ~new_n11206_;
  assign new_n11208_ = ~new_n11204_ & ~new_n11207_;
  assign new_n11209_ = ~new_n4790_ & new_n11208_;
  assign new_n11210_ = ~new_n4790_ & ~new_n11209_;
  assign new_n11211_ = new_n11208_ & ~new_n11209_;
  assign new_n11212_ = ~new_n11210_ & ~new_n11211_;
  assign new_n11213_ = ~new_n5080_ & new_n11212_;
  assign new_n11214_ = ng826 & ~new_n11213_;
  assign new_n11215_ = ~ng312 & ~ng826;
  assign n4158 = ~new_n11214_ & ~new_n11215_;
  assign new_n11217_ = ng823 & n4167;
  assign new_n11218_ = ~ng484 & ~ng823;
  assign n4176 = ~new_n11217_ & ~new_n11218_;
  assign new_n11220_ = ng1315 & ~ng484;
  assign new_n11221_ = ~ng464 & ng1309;
  assign new_n11222_ = ng1312 & ~ng480;
  assign new_n11223_ = ~new_n11220_ & ~new_n11221_;
  assign n4181 = ~new_n11222_ & new_n11223_;
  assign new_n11225_ = ~ng720 & ~new_n5395_;
  assign new_n11226_ = ng679 & new_n5395_;
  assign n4196 = ~new_n11225_ & ~new_n11226_;
  assign new_n11228_ = ~ng857 & ~new_n5538_;
  assign new_n11229_ = new_n5538_ & ~new_n9372_;
  assign n4206 = ~new_n11228_ & ~new_n11229_;
  assign new_n11231_ = ~ng865 & ~new_n8121_;
  assign new_n11232_ = new_n5967_1_ & new_n8121_;
  assign n4211 = ~new_n11231_ & ~new_n11232_;
  assign new_n11234_ = ng767 & ~new_n5913_1_;
  assign new_n11235_ = ~ng767 & new_n5913_1_;
  assign new_n11236_ = ~new_n11234_ & ~new_n11235_;
  assign n4216 = ~new_n5127_1_ & ~new_n11236_;
  assign new_n11238_ = ~ng1045 & ~new_n7915_;
  assign new_n11239_ = new_n5932_ & ~new_n5937_;
  assign new_n11240_ = ~pg3229 & new_n11239_;
  assign new_n11241_ = ~new_n5932_ & ~new_n5937_;
  assign new_n11242_ = pg3229 & new_n11241_;
  assign new_n11243_ = new_n5937_ & ~new_n5942_;
  assign new_n11244_ = ~new_n11240_ & ~new_n11242_;
  assign new_n11245_ = ~new_n11243_ & new_n11244_;
  assign new_n11246_ = new_n7915_ & ~new_n11245_;
  assign n4221 = ~new_n11238_ & ~new_n11246_;
  assign new_n11248_ = ng1315 & ~ng1243;
  assign new_n11249_ = ~ng1315 & ~ng1196;
  assign n4240 = ~new_n11248_ & ~new_n11249_;
  assign new_n11251_ = ng1312 & ~new_n10886_;
  assign new_n11252_ = ~ng1312 & ~ng1276;
  assign n4250 = ~new_n11251_ & ~new_n11252_;
  assign new_n11254_ = ng1309 & ~new_n9421_;
  assign new_n11255_ = ~ng1177 & ~ng1309;
  assign n4255 = ~new_n11254_ & ~new_n11255_;
  assign new_n11257_ = ~ng1358 & new_n6247_;
  assign new_n11258_ = ng1358 & ~new_n6247_;
  assign new_n11259_ = ~new_n11257_ & ~new_n11258_;
  assign n4265 = ~new_n6241_ & ~new_n11259_;
  assign new_n11261_ = ~ng1384 & ~new_n6263_;
  assign new_n11262_ = ng1326 & new_n6263_;
  assign n4270 = ~new_n11261_ & ~new_n11262_;
  assign new_n11264_ = ~ng1398 & ~new_n6255_;
  assign new_n11265_ = ng1346 & new_n6255_;
  assign n4275 = ~new_n11264_ & ~new_n11265_;
  assign new_n11267_ = ~ng1529 & ~new_n4773_;
  assign new_n11268_ = ng1491 & new_n4773_;
  assign n4280 = ~new_n11267_ & ~new_n11268_;
  assign new_n11270_ = ~ng1543 & ~new_n4777_1_;
  assign new_n11271_ = new_n4777_1_ & ~new_n6436_;
  assign n4285 = ~new_n11270_ & ~new_n11271_;
  assign new_n11273_ = ~ng1559 & ~new_n8121_;
  assign new_n11274_ = new_n6678_ & new_n8121_;
  assign n4290 = ~new_n11273_ & ~new_n11274_;
  assign new_n11276_ = ng1486 & ~new_n6587_;
  assign new_n11277_ = ~new_n10383_ & ~new_n11276_;
  assign new_n11278_ = ~new_n6586_ & new_n11277_;
  assign new_n11279_ = new_n6600_1_ & ~new_n6606_;
  assign new_n11280_ = new_n6314_1_ & new_n11279_;
  assign new_n11281_ = ~new_n6314_1_ & ~new_n11279_;
  assign new_n11282_ = ~new_n11280_ & ~new_n11281_;
  assign new_n11283_ = new_n6586_ & new_n11282_;
  assign new_n11284_ = ~new_n11278_ & ~new_n11283_;
  assign new_n11285_ = ng823 & ~new_n11284_;
  assign new_n11286_ = ~ng1624 & ~ng823;
  assign n4295 = ~new_n11285_ & ~new_n11286_;
  assign new_n11288_ = ng1496 & ~new_n6587_;
  assign new_n11289_ = ~new_n6586_ & ~new_n11288_;
  assign new_n11290_ = ~new_n6613_ & new_n6615_;
  assign new_n11291_ = new_n6341_ & new_n11290_;
  assign new_n11292_ = ~new_n6341_ & ~new_n11290_;
  assign new_n11293_ = ~new_n11291_ & ~new_n11292_;
  assign new_n11294_ = new_n6586_ & new_n11293_;
  assign new_n11295_ = ~new_n11289_ & ~new_n11294_;
  assign new_n11296_ = ng853 & ~new_n11295_;
  assign new_n11297_ = ~ng1636 & ~ng853;
  assign n4300 = ~new_n11296_ & ~new_n11297_;
  assign new_n11299_ = ng823 & ~new_n10930_;
  assign new_n11300_ = ~ng1651 & ~ng823;
  assign n4305 = ~new_n11299_ & ~new_n11300_;
  assign new_n11302_ = ~ng1784 & ~new_n6003_;
  assign new_n11303_ = new_n6003_ & new_n9507_;
  assign n4310 = ~new_n11302_ & ~new_n11303_;
  assign new_n11305_ = ~ng2222 & ~new_n4777_1_;
  assign new_n11306_ = ng2180 & new_n4777_1_;
  assign n4334 = ~new_n11305_ & ~new_n11306_;
  assign new_n11308_ = ~ng2233 & ~new_n5517_1_;
  assign new_n11309_ = ng2200 & new_n5517_1_;
  assign n4339 = ~new_n11308_ & ~new_n11309_;
  assign new_n11311_ = ng853 & ~new_n9552_;
  assign new_n11312_ = ~ng2321 & ~ng853;
  assign n4344 = ~new_n11311_ & ~new_n11312_;
  assign new_n11314_ = ~new_n7494_ & new_n7500_;
  assign new_n11315_ = new_n7500_ & ~new_n11314_;
  assign new_n11316_ = ~new_n7494_ & ~new_n11314_;
  assign new_n11317_ = ~new_n11315_ & ~new_n11316_;
  assign new_n11318_ = ng2384 & ~new_n11317_;
  assign new_n11319_ = ~new_n7494_ & ~new_n11318_;
  assign new_n11320_ = ~new_n7494_ & ~new_n11319_;
  assign new_n11321_ = ~new_n11318_ & ~new_n11319_;
  assign new_n11322_ = ~new_n11320_ & ~new_n11321_;
  assign new_n11323_ = ng826 & ~new_n11322_;
  assign new_n11324_ = ~ng826 & ~ng2504;
  assign n4349 = ~new_n11323_ & ~new_n11324_;
  assign new_n11326_ = ng853 & ~new_n10440_;
  assign new_n11327_ = ~ng2389 & ~ng853;
  assign n4354 = ~new_n11326_ & ~new_n11327_;
  assign new_n11329_ = ~ng2374 & ng2373;
  assign new_n11330_ = ~ng1680 & ng1679;
  assign new_n11331_ = ng823 & n467;
  assign new_n11332_ = ~ng823 & ng1686;
  assign new_n11333_ = ~new_n11331_ & ~new_n11332_;
  assign new_n11334_ = ng1680 & new_n11333_;
  assign n6412 = ~new_n11330_ & ~new_n11334_;
  assign new_n11336_ = ng823 & n6412;
  assign new_n11337_ = ng2380 & ~ng823;
  assign new_n11338_ = ~new_n11336_ & ~new_n11337_;
  assign new_n11339_ = ng2374 & new_n11338_;
  assign n4367 = ~new_n11329_ & ~new_n11339_;
  assign new_n11341_ = ng823 & n2815;
  assign new_n11342_ = ~ng2559 & ~ng823;
  assign n4377 = ~new_n11341_ & ~new_n11342_;
  assign new_n11344_ = ng1315 & ~ng2559;
  assign new_n11345_ = ng1309 & ~ng2539;
  assign new_n11346_ = ng1312 & ~ng2555;
  assign new_n11347_ = ~new_n11344_ & ~new_n11345_;
  assign n4382 = ~new_n11346_ & new_n11347_;
  assign new_n11349_ = ~ng2660 & ~new_n8209_;
  assign new_n11350_ = new_n8209_ & ~new_n10956_;
  assign n4387 = ~new_n11349_ & ~new_n11350_;
  assign new_n11352_ = ~new_n10512_ & new_n10578_;
  assign new_n11353_ = new_n10520_ & new_n11352_;
  assign new_n11354_ = new_n9616_ & new_n10578_;
  assign new_n11355_ = ~new_n10520_ & new_n11354_;
  assign new_n11356_ = ~new_n11353_ & ~new_n11355_;
  assign new_n11357_ = new_n5366_ & new_n11356_;
  assign new_n11358_ = ~new_n5366_ & new_n7529_;
  assign new_n11359_ = ~new_n11357_ & ~new_n11358_;
  assign new_n11360_ = ng1309 & ~new_n11359_;
  assign new_n11361_ = ~ng2679 & ~ng1309;
  assign n4392 = ~new_n11360_ & ~new_n11361_;
  assign new_n11363_ = ~pg3229 & ~ng2380;
  assign new_n11364_ = pg3229 & ng2366;
  assign n4402 = ~new_n11363_ & ~new_n11364_;
  assign new_n11366_ = ~ng2774 & ~new_n7588_;
  assign new_n11367_ = ng2714 & new_n7588_;
  assign n4407 = ~new_n11366_ & ~new_n11367_;
  assign new_n11369_ = ~ng2792 & ~new_n7588_;
  assign new_n11370_ = ng2740 & new_n7588_;
  assign n4412 = ~new_n11369_ & ~new_n11370_;
  assign new_n11372_ = ng2704 & ng1309;
  assign new_n11373_ = ~ng2803 & ~new_n11372_;
  assign new_n11374_ = ~new_n7540_ & new_n11372_;
  assign n4417 = ~new_n11373_ & ~new_n11374_;
  assign new_n11376_ = ~ng1215 & new_n11015_;
  assign new_n11377_ = ~new_n11139_ & new_n11376_;
  assign new_n11378_ = new_n11057_ & new_n11139_;
  assign new_n11379_ = ~new_n11377_ & ~new_n11378_;
  assign new_n11380_ = ~new_n11141_ & new_n11379_;
  assign new_n11381_ = ~new_n11139_ & new_n11141_;
  assign new_n11382_ = ng1312 & ~ng1422;
  assign new_n11383_ = ng1315 & ~ng1420;
  assign new_n11384_ = ng1309 & ~ng1421;
  assign new_n11385_ = ~new_n11382_ & ~new_n11383_;
  assign new_n11386_ = ~new_n11384_ & new_n11385_;
  assign new_n11387_ = ~new_n11031_ & new_n11386_;
  assign new_n11388_ = ng1186 & ~new_n11387_;
  assign new_n11389_ = new_n11015_ & new_n11388_;
  assign new_n11390_ = new_n11381_ & ~new_n11389_;
  assign new_n11391_ = new_n11141_ & new_n11390_;
  assign n4422 = new_n11380_ | new_n11391_;
  assign new_n11393_ = ~ng1911 & new_n10635_;
  assign new_n11394_ = ~new_n10633_ & new_n11393_;
  assign new_n11395_ = ~new_n10657_ & ~new_n10708_;
  assign new_n11396_ = ~new_n6785_ & ~new_n11395_;
  assign new_n11397_ = ~new_n11395_ & ~new_n11396_;
  assign new_n11398_ = ~new_n6785_ & ~new_n11396_;
  assign new_n11399_ = ~new_n11397_ & ~new_n11398_;
  assign new_n11400_ = new_n10635_ & ~new_n11399_;
  assign new_n11401_ = ng1880 & new_n11400_;
  assign new_n11402_ = new_n10633_ & new_n11401_;
  assign new_n11403_ = ~new_n11394_ & ~new_n11402_;
  assign new_n11404_ = ~new_n10631_ & new_n11403_;
  assign new_n11405_ = new_n10635_ & ~new_n10726_;
  assign new_n11406_ = new_n10719_ & ~new_n11405_;
  assign new_n11407_ = new_n10631_ & new_n11406_;
  assign n4427 = new_n11404_ | new_n11407_;
  assign new_n11409_ = ~ng2603 & new_n10738_;
  assign new_n11410_ = ~new_n10736_ & new_n11409_;
  assign new_n11411_ = ~new_n8304_ & ~new_n10756_;
  assign new_n11412_ = ~new_n7529_ & ~new_n11411_;
  assign new_n11413_ = ~new_n11411_ & ~new_n11412_;
  assign new_n11414_ = ~new_n7529_ & ~new_n11412_;
  assign new_n11415_ = ~new_n11413_ & ~new_n11414_;
  assign new_n11416_ = new_n10738_ & ~new_n11415_;
  assign new_n11417_ = ng2574 & new_n11416_;
  assign new_n11418_ = new_n10736_ & new_n11417_;
  assign new_n11419_ = ~new_n11410_ & ~new_n11418_;
  assign new_n11420_ = ~new_n10734_ & new_n11419_;
  assign n4432 = new_n11165_ | new_n11420_;
  assign new_n11422_ = ~ng3006 & new_n10782_;
  assign new_n11423_ = ng3006 & ~new_n10782_;
  assign new_n11424_ = ~new_n11422_ & ~new_n11423_;
  assign n4437 = new_n10780_ & ~new_n11424_;
  assign new_n11426_ = ~ng3065 & ng2987;
  assign new_n11427_ = ~ng3046 & ~ng2987;
  assign n4442 = ~new_n11426_ & ~new_n11427_;
  assign new_n11429_ = ~ng3074 & ng2987;
  assign new_n11430_ = ~ng3056 & ~ng2987;
  assign n4447 = ~new_n11429_ & ~new_n11430_;
  assign new_n11432_ = ~pg3231 & ng3120;
  assign new_n11433_ = ~ng20 & ~ng23;
  assign new_n11434_ = ~ng23 & ~new_n11433_;
  assign new_n11435_ = ~ng20 & ~new_n11433_;
  assign new_n11436_ = ~new_n11434_ & ~new_n11435_;
  assign new_n11437_ = ~ng11 & ~ng17;
  assign new_n11438_ = ~ng17 & ~new_n11437_;
  assign new_n11439_ = ~ng11 & ~new_n11437_;
  assign new_n11440_ = ~new_n11438_ & ~new_n11439_;
  assign new_n11441_ = ~new_n11436_ & ~new_n11440_;
  assign new_n11442_ = ~new_n11436_ & ~new_n11441_;
  assign new_n11443_ = ~new_n11440_ & ~new_n11441_;
  assign new_n11444_ = ~new_n11442_ & ~new_n11443_;
  assign new_n11445_ = ~ng5 & ~ng14;
  assign new_n11446_ = ~ng14 & ~new_n11445_;
  assign new_n11447_ = ~ng5 & ~new_n11445_;
  assign new_n11448_ = ~new_n11446_ & ~new_n11447_;
  assign new_n11449_ = ~ng8 & ~ng2;
  assign new_n11450_ = ~ng8 & ~new_n11449_;
  assign new_n11451_ = ~ng2 & ~new_n11449_;
  assign new_n11452_ = ~new_n11450_ & ~new_n11451_;
  assign new_n11453_ = ~new_n11448_ & ~new_n11452_;
  assign new_n11454_ = ~new_n11448_ & ~new_n11453_;
  assign new_n11455_ = ~new_n11452_ & ~new_n11453_;
  assign new_n11456_ = ~new_n11454_ & ~new_n11455_;
  assign new_n11457_ = ~new_n11444_ & ~new_n11456_;
  assign new_n11458_ = ~new_n11444_ & ~new_n11457_;
  assign new_n11459_ = ~new_n11456_ & ~new_n11457_;
  assign new_n11460_ = ~new_n11458_ & ~new_n11459_;
  assign new_n11461_ = new_n11432_ & ~new_n11460_;
  assign new_n11462_ = new_n11432_ & ~new_n11461_;
  assign new_n11463_ = ~new_n11460_ & ~new_n11461_;
  assign n4452 = new_n11462_ | new_n11463_;
  assign new_n11465_ = ~ng2903 & new_n9238_;
  assign new_n11466_ = ng2903 & ~new_n9238_;
  assign new_n11467_ = ~new_n11465_ & ~new_n11466_;
  assign n4457 = new_n9234_ & ~new_n11467_;
  assign new_n11469_ = ~ng133 & ~new_n5517_1_;
  assign new_n11470_ = ng101 & new_n5517_1_;
  assign n4462 = ~new_n11469_ & ~new_n11470_;
  assign new_n11472_ = ~ng148 & ~new_n5517_1_;
  assign new_n11473_ = ng113 & new_n5517_1_;
  assign n4467 = ~new_n11472_ & ~new_n11473_;
  assign new_n11475_ = ~ng157 & ~new_n5517_1_;
  assign new_n11476_ = ng125 & new_n5517_1_;
  assign n4472 = ~new_n11475_ & ~new_n11476_;
  assign new_n11478_ = ~ng169 & ~new_n5538_;
  assign new_n11479_ = new_n5538_ & ~new_n10811_;
  assign n4477 = ~new_n11478_ & ~new_n11479_;
  assign new_n11481_ = ng853 & ~new_n10821_;
  assign new_n11482_ = ~ng237 & ~ng853;
  assign n4482 = ~new_n11481_ & ~new_n11482_;
  assign new_n11484_ = ng853 & ~new_n10314_;
  assign new_n11485_ = ~ng210 & ~ng853;
  assign n4487 = ~new_n11484_ & ~new_n11485_;
  assign new_n11487_ = ng853 & ~new_n10836_;
  assign new_n11488_ = ~ng426 & ~new_n11487_;
  assign new_n11489_ = new_n10833_ & new_n11487_;
  assign n4492 = ~new_n11488_ & ~new_n11489_;
  assign new_n11491_ = ng853 & ~new_n8412_;
  assign new_n11492_ = ~ng447 & ~new_n11491_;
  assign new_n11493_ = new_n8405_ & new_n11491_;
  assign n4497 = ~new_n11492_ & ~new_n11493_;
  assign new_n11495_ = ng853 & ~new_n5273_;
  assign new_n11496_ = ~ng320 & ~ng853;
  assign n4502 = ~new_n11495_ & ~new_n11496_;
  assign new_n11498_ = ng853 & n4167;
  assign new_n11499_ = ~ng464 & ~ng853;
  assign n4516 = ~new_n11498_ & ~new_n11499_;
  assign new_n11501_ = ~pg3229 & ~ng305;
  assign new_n11502_ = pg3229 & ng291;
  assign n4530 = ~new_n11501_ & ~new_n11502_;
  assign new_n11504_ = ~ng730 & ~new_n5380_;
  assign new_n11505_ = ~new_n5302_1_ & new_n5380_;
  assign n4535 = ~new_n11504_ & ~new_n11505_;
  assign new_n11507_ = ng1315 & ng630;
  assign new_n11508_ = ~ng728 & ~new_n11507_;
  assign new_n11509_ = ~new_n5302_1_ & new_n11507_;
  assign n4540 = ~new_n11508_ & ~new_n11509_;
  assign new_n11511_ = ~ng858 & ~new_n6278_;
  assign new_n11512_ = new_n6278_ & ~new_n9372_;
  assign n4545 = ~new_n11511_ & ~new_n11512_;
  assign new_n11514_ = ~ng867 & ~new_n6278_;
  assign new_n11515_ = new_n5967_1_ & new_n6278_;
  assign n4550 = ~new_n11514_ & ~new_n11515_;
  assign new_n11517_ = ~ng762 & new_n5914_;
  assign new_n11518_ = ng762 & ~new_n5914_;
  assign new_n11519_ = ~new_n11517_ & ~new_n11518_;
  assign n4555 = ~new_n5127_1_ & ~new_n11519_;
  assign new_n11521_ = ~ng1056 & ~new_n5926_;
  assign new_n11522_ = new_n5926_ & ~new_n11245_;
  assign n4560 = ~new_n11521_ & ~new_n11522_;
  assign new_n11524_ = ng1315 & ~new_n10886_;
  assign new_n11525_ = ~ng1315 & ~ng1279;
  assign n4585 = ~new_n11524_ & ~new_n11525_;
  assign new_n11527_ = ng1315 & ~new_n8573_;
  assign new_n11528_ = ~ng1315 & ~ng1297;
  assign n4590 = ~new_n11527_ & ~new_n11528_;
  assign new_n11530_ = ng1346 & ~new_n6246_;
  assign new_n11531_ = ~ng1346 & new_n6246_;
  assign new_n11532_ = ~new_n11530_ & ~new_n11531_;
  assign n4599 = ~new_n6241_ & ~new_n11532_;
  assign new_n11534_ = ~ng1388 & ~new_n6259_1_;
  assign new_n11535_ = ng1319 & new_n6259_1_;
  assign n4604 = ~new_n11534_ & ~new_n11535_;
  assign new_n11537_ = ~ng1397 & ~new_n6259_1_;
  assign new_n11538_ = ng1346 & new_n6259_1_;
  assign n4609 = ~new_n11537_ & ~new_n11538_;
  assign new_n11540_ = ~ng1533 & ~new_n5517_1_;
  assign new_n11541_ = ng1496 & new_n5517_1_;
  assign n4614 = ~new_n11540_ & ~new_n11541_;
  assign new_n11543_ = ~ng1542 & ~new_n5517_1_;
  assign new_n11544_ = new_n5517_1_ & ~new_n6436_;
  assign n4619 = ~new_n11543_ & ~new_n11544_;
  assign new_n11546_ = ng826 & ~new_n8712_;
  assign new_n11547_ = ~ng826 & ~ng1567;
  assign n4624 = ~new_n11546_ & ~new_n11547_;
  assign new_n11549_ = ng826 & ~new_n11284_;
  assign new_n11550_ = ~ng826 & ~ng1621;
  assign n4629 = ~new_n11549_ & ~new_n11550_;
  assign new_n11552_ = ng826 & ~new_n10400_;
  assign new_n11553_ = ~ng826 & ~ng1594;
  assign n4634 = ~new_n11552_ & ~new_n11553_;
  assign new_n11555_ = ng826 & ~new_n10930_;
  assign new_n11556_ = ~ng826 & ~ng1648;
  assign n4639 = ~new_n11555_ & ~new_n11556_;
  assign new_n11558_ = ng853 & ~new_n9474_;
  assign new_n11559_ = ~ng1695 & ~ng853;
  assign n4644 = ~new_n11558_ & ~new_n11559_;
  assign new_n11561_ = ~ng2220 & ~new_n4773_;
  assign new_n11562_ = ng2180 & new_n4773_;
  assign n4666 = ~new_n11561_ & ~new_n11562_;
  assign new_n11564_ = ~ng2229 & ~new_n4773_;
  assign new_n11565_ = ng2195 & new_n4773_;
  assign n4671 = ~new_n11564_ & ~new_n11565_;
  assign new_n11567_ = ng826 & ~new_n9574_;
  assign new_n11568_ = ~ng826 & ~ng2333;
  assign n4676 = ~new_n11567_ & ~new_n11568_;
  assign new_n11570_ = ng823 & ~new_n11322_;
  assign new_n11571_ = ~ng2507 & ~ng823;
  assign n4681 = ~new_n11570_ & ~new_n11571_;
  assign new_n11573_ = ng823 & ~new_n10440_;
  assign new_n11574_ = ~ng2388 & ~ng823;
  assign n4686 = ~new_n11573_ & ~new_n11574_;
  assign new_n11576_ = ng2120 & new_n7067_;
  assign new_n11577_ = new_n7067_ & ~new_n11576_;
  assign new_n11578_ = ng2120 & ~new_n11576_;
  assign new_n11579_ = ~new_n11577_ & ~new_n11578_;
  assign new_n11580_ = ng2133 & new_n7094_;
  assign new_n11581_ = new_n7094_ & ~new_n11580_;
  assign new_n11582_ = ng2133 & ~new_n11580_;
  assign new_n11583_ = ~new_n11581_ & ~new_n11582_;
  assign new_n11584_ = ng2129 & new_n7072_;
  assign new_n11585_ = new_n7072_ & ~new_n11584_;
  assign new_n11586_ = ng2129 & ~new_n11584_;
  assign new_n11587_ = ~new_n11585_ & ~new_n11586_;
  assign new_n11588_ = ng2138 & new_n7082_1_;
  assign new_n11589_ = new_n7082_1_ & ~new_n11588_;
  assign new_n11590_ = ng2138 & ~new_n11588_;
  assign new_n11591_ = ~new_n11589_ & ~new_n11590_;
  assign new_n11592_ = ~new_n11583_ & ~new_n11587_;
  assign new_n11593_ = ~new_n11591_ & new_n11592_;
  assign new_n11594_ = ng2124 & new_n7101_;
  assign new_n11595_ = new_n7101_ & ~new_n11594_;
  assign new_n11596_ = ng2124 & ~new_n11594_;
  assign new_n11597_ = ~new_n11595_ & ~new_n11596_;
  assign new_n11598_ = ~new_n11579_ & new_n11593_;
  assign new_n11599_ = ~new_n11597_ & new_n11598_;
  assign new_n11600_ = ng2142 & new_n7077_;
  assign new_n11601_ = new_n7077_ & ~new_n11600_;
  assign new_n11602_ = ng2142 & ~new_n11600_;
  assign new_n11603_ = ~new_n11601_ & ~new_n11602_;
  assign new_n11604_ = ng2156 & new_n7060_;
  assign new_n11605_ = new_n7060_ & ~new_n11604_;
  assign new_n11606_ = ng2156 & ~new_n11604_;
  assign new_n11607_ = ~new_n11605_ & ~new_n11606_;
  assign new_n11608_ = ng2151 & new_n7050_;
  assign new_n11609_ = new_n7050_ & ~new_n11608_;
  assign new_n11610_ = ng2151 & ~new_n11608_;
  assign new_n11611_ = ~new_n11609_ & ~new_n11610_;
  assign new_n11612_ = ng2160 & new_n7087_1_;
  assign new_n11613_ = new_n7087_1_ & ~new_n11612_;
  assign new_n11614_ = ng2160 & ~new_n11612_;
  assign new_n11615_ = ~new_n11613_ & ~new_n11614_;
  assign new_n11616_ = ~new_n11607_ & ~new_n11611_;
  assign new_n11617_ = ~new_n11615_ & new_n11616_;
  assign new_n11618_ = ng2147 & new_n7055_;
  assign new_n11619_ = new_n7055_ & ~new_n11618_;
  assign new_n11620_ = ng2147 & ~new_n11618_;
  assign new_n11621_ = ~new_n11619_ & ~new_n11620_;
  assign new_n11622_ = ~new_n11603_ & new_n11617_;
  assign new_n11623_ = ~new_n11621_ & new_n11622_;
  assign new_n11624_ = ~new_n7408_ & new_n11599_;
  assign new_n11625_ = new_n11623_ & new_n11624_;
  assign new_n11626_ = ~new_n5125_ & new_n11625_;
  assign new_n11627_ = new_n7044_ & new_n7110_;
  assign new_n11628_ = ~new_n11626_ & ~new_n11627_;
  assign n4699 = ~new_n7409_ | new_n11628_;
  assign new_n11630_ = ng853 & n2815;
  assign new_n11631_ = ~ng2539 & ~ng853;
  assign n4708 = ~new_n11630_ & ~new_n11631_;
  assign new_n11633_ = ~ng2658 & ~new_n7545_;
  assign new_n11634_ = new_n7545_ & ~new_n10956_;
  assign n4718 = ~new_n11633_ & ~new_n11634_;
  assign new_n11636_ = ng1315 & ~new_n10584_;
  assign new_n11637_ = ~ng1315 & ~ng2694;
  assign n4723 = ~new_n11636_ & ~new_n11637_;
  assign new_n11639_ = ng2580 & ~ng2581;
  assign new_n11640_ = ng1886 & ~ng1887;
  assign new_n11641_ = ng1312 & n996;
  assign new_n11642_ = ~ng1312 & ng1900;
  assign new_n11643_ = ~new_n11641_ & ~new_n11642_;
  assign new_n11644_ = ~ng1886 & new_n11643_;
  assign n7300 = ~new_n11640_ & ~new_n11644_;
  assign new_n11646_ = ng1312 & n7300;
  assign new_n11647_ = ~ng1312 & ng2594;
  assign new_n11648_ = ~new_n11646_ & ~new_n11647_;
  assign new_n11649_ = ~ng2580 & new_n11648_;
  assign n4728 = ~new_n11639_ & ~new_n11649_;
  assign new_n11651_ = ~ng2781 & ~new_n7584_;
  assign new_n11652_ = ng2720 & new_n7584_;
  assign n4737 = ~new_n11651_ & ~new_n11652_;
  assign new_n11654_ = ~ng2790 & ~new_n7584_;
  assign new_n11655_ = ng2740 & new_n7584_;
  assign n4742 = ~new_n11654_ & ~new_n11655_;
  assign new_n11657_ = ~ng2799 & ~new_n7584_;
  assign new_n11658_ = ng2766 & new_n7584_;
  assign n4747 = ~new_n11657_ & ~new_n11658_;
  assign new_n11660_ = ~ng1216 & new_n11015_;
  assign new_n11661_ = ~new_n11139_ & new_n11660_;
  assign new_n11662_ = new_n11064_ & new_n11139_;
  assign new_n11663_ = ~new_n11661_ & ~new_n11662_;
  assign new_n11664_ = ~new_n11141_ & new_n11663_;
  assign new_n11665_ = new_n11015_ & ~new_n11388_;
  assign new_n11666_ = new_n11381_ & ~new_n11665_;
  assign new_n11667_ = new_n11141_ & new_n11666_;
  assign n4752 = new_n11664_ | new_n11667_;
  assign new_n11669_ = ~ng1910 & new_n10635_;
  assign new_n11670_ = ~new_n10633_ & new_n11669_;
  assign new_n11671_ = ~new_n10652_ & ~new_n10708_;
  assign new_n11672_ = ~new_n6796_ & ~new_n11671_;
  assign new_n11673_ = ~new_n11671_ & ~new_n11672_;
  assign new_n11674_ = ~new_n6796_ & ~new_n11672_;
  assign new_n11675_ = ~new_n11673_ & ~new_n11674_;
  assign new_n11676_ = new_n10635_ & ~new_n11675_;
  assign new_n11677_ = ng1880 & new_n11676_;
  assign new_n11678_ = new_n10633_ & new_n11677_;
  assign new_n11679_ = ~new_n11670_ & ~new_n11678_;
  assign new_n11680_ = ~new_n10631_ & new_n11679_;
  assign n4757 = new_n11407_ | new_n11680_;
  assign new_n11682_ = ~ng2604 & new_n10738_;
  assign new_n11683_ = ~new_n10736_ & new_n11682_;
  assign new_n11684_ = ~new_n8295_ & ~new_n10756_;
  assign new_n11685_ = ~new_n7540_ & ~new_n11684_;
  assign new_n11686_ = ~new_n11684_ & ~new_n11685_;
  assign new_n11687_ = ~new_n7540_ & ~new_n11685_;
  assign new_n11688_ = ~new_n11686_ & ~new_n11687_;
  assign new_n11689_ = new_n10738_ & ~new_n11688_;
  assign new_n11690_ = ng2574 & new_n11689_;
  assign new_n11691_ = new_n10736_ & new_n11690_;
  assign new_n11692_ = ~new_n11683_ & ~new_n11691_;
  assign new_n11693_ = ~new_n10734_ & new_n11692_;
  assign n4762 = new_n10777_ | new_n11693_;
  assign new_n11695_ = ~pg3234 & ~new_n10780_;
  assign new_n11696_ = ng2998 & ~new_n10781_;
  assign new_n11697_ = ~ng2998 & new_n10781_;
  assign new_n11698_ = ~new_n11696_ & ~new_n11697_;
  assign new_n11699_ = new_n10780_ & new_n11698_;
  assign n4767 = ~new_n11695_ & ~new_n11699_;
  assign new_n11701_ = ~ng3066 & ng2987;
  assign new_n11702_ = ~ng3047 & ~ng2987;
  assign n4772 = ~new_n11701_ & ~new_n11702_;
  assign new_n11704_ = ~ng3073 & ng2987;
  assign new_n11705_ = ~ng3055 & ~ng2987;
  assign n4777 = ~new_n11704_ & ~new_n11705_;
  assign n4782 = ~pg51 & ng2950;
  assign new_n11708_ = ng1312 & ~n1448;
  assign new_n11709_ = ~ng1312 & ~ng3101;
  assign n4787 = ~new_n11708_ & ~new_n11709_;
  assign new_n11711_ = ~ng1186 & ng1309;
  assign new_n11712_ = ~ng1309 & ~ng3164;
  assign n4792 = ~new_n11711_ & ~new_n11712_;
  assign new_n11714_ = ~ng134 & ~new_n4777_1_;
  assign new_n11715_ = ng101 & new_n4777_1_;
  assign n4797 = ~new_n11714_ & ~new_n11715_;
  assign new_n11717_ = ~ng151 & ~new_n5517_1_;
  assign new_n11718_ = ng117 & new_n5517_1_;
  assign n4802 = ~new_n11717_ & ~new_n11718_;
  assign new_n11720_ = ~ng159 & ~new_n4773_;
  assign new_n11721_ = new_n4773_ & ~new_n4932_1_;
  assign n4807 = ~new_n11720_ & ~new_n11721_;
  assign new_n11723_ = ~ng176 & ~new_n6278_;
  assign new_n11724_ = ng97 & new_n6278_;
  assign n4812 = ~new_n11723_ & ~new_n11724_;
  assign new_n11726_ = ~ng179 & ~new_n6278_;
  assign new_n11727_ = new_n5180_ & new_n6278_;
  assign n4817 = ~new_n11726_ & ~new_n11727_;
  assign new_n11729_ = ng109 & ~new_n5083_;
  assign new_n11730_ = ~new_n8915_ & ~new_n11729_;
  assign new_n11731_ = ~new_n5082_1_ & new_n11730_;
  assign new_n11732_ = new_n5096_ & ~new_n5102_1_;
  assign new_n11733_ = new_n4810_ & new_n11732_;
  assign new_n11734_ = ~new_n4810_ & ~new_n11732_;
  assign new_n11735_ = ~new_n11733_ & ~new_n11734_;
  assign new_n11736_ = new_n5082_1_ & new_n11735_;
  assign new_n11737_ = ~new_n11731_ & ~new_n11736_;
  assign new_n11738_ = ng826 & ~new_n11737_;
  assign new_n11739_ = ~ng826 & ~ng240;
  assign n4822 = ~new_n11738_ & ~new_n11739_;
  assign new_n11741_ = ng823 & ~new_n8929_;
  assign new_n11742_ = ~ng225 & ~ng823;
  assign n4827 = ~new_n11741_ & ~new_n11742_;
  assign new_n11744_ = ~ng65 & new_n9291_;
  assign new_n11745_ = ng65 & ~new_n9291_;
  assign new_n11746_ = ~new_n11744_ & ~new_n11745_;
  assign n4832 = ~new_n5127_1_ & ~new_n11746_;
  assign new_n11748_ = ~ng373 & ~new_n7672_;
  assign new_n11749_ = new_n7672_ & ~new_n9901_;
  assign n4837 = ~new_n11748_ & ~new_n11749_;
  assign new_n11751_ = ~new_n5222_1_ & new_n5228_;
  assign new_n11752_ = new_n5228_ & ~new_n11751_;
  assign new_n11753_ = ~new_n5222_1_ & ~new_n11751_;
  assign new_n11754_ = ~new_n11752_ & ~new_n11753_;
  assign new_n11755_ = ng2384 & ~new_n11754_;
  assign new_n11756_ = ~new_n5222_1_ & ~new_n11755_;
  assign new_n11757_ = ~new_n5222_1_ & ~new_n11756_;
  assign new_n11758_ = ~new_n11755_ & ~new_n11756_;
  assign new_n11759_ = ~new_n11757_ & ~new_n11758_;
  assign new_n11760_ = ng826 & ~new_n11759_;
  assign new_n11761_ = ~ng826 & ~ng429;
  assign n4842 = ~new_n11760_ & ~new_n11761_;
  assign new_n11763_ = ng853 & ~new_n11213_;
  assign new_n11764_ = ~ng314 & ~ng853;
  assign n4847 = ~new_n11763_ & ~new_n11764_;
  assign new_n11766_ = ~ng404 & ~new_n9772_;
  assign new_n11767_ = new_n5067_1_ & new_n5079_;
  assign new_n11768_ = new_n9772_ & new_n11767_;
  assign n4852 = ~new_n11766_ & ~new_n11768_;
  assign new_n11770_ = ng826 & n4167;
  assign new_n11771_ = ~ng826 & ~ng480;
  assign n4882 = ~new_n11770_ & ~new_n11771_;
  assign new_n11773_ = ng826 & ~new_n4799_;
  assign new_n11774_ = ~ng826 & ~ng465;
  assign n4887 = ~new_n11773_ & ~new_n11774_;
  assign new_n11776_ = ng1315 & ~ng487;
  assign new_n11777_ = ~ng488 & ng1309;
  assign new_n11778_ = ng1312 & ~ng486;
  assign new_n11779_ = ~new_n11776_ & ~new_n11777_;
  assign n4892 = ~new_n11778_ & new_n11779_;
  assign new_n11781_ = ~ng585 & ~new_n8959_;
  assign new_n11782_ = ~new_n8439_ & new_n8959_;
  assign n4897 = ~new_n11781_ & ~new_n11782_;
  assign new_n11784_ = new_n7784_ & ~new_n7855_;
  assign new_n11785_ = new_n5356_ & new_n11784_;
  assign new_n11786_ = ~new_n7840_ & new_n7855_;
  assign new_n11787_ = new_n7784_ & new_n11786_;
  assign new_n11788_ = ~new_n11785_ & ~new_n11787_;
  assign new_n11789_ = new_n5366_ & new_n11788_;
  assign new_n11790_ = new_n5302_1_ & ~new_n5366_;
  assign new_n11791_ = ~new_n11789_ & ~new_n11790_;
  assign new_n11792_ = ng1315 & ~new_n11791_;
  assign new_n11793_ = ~ng1315 & ~ng620;
  assign n4902 = ~new_n11792_ & ~new_n11793_;
  assign new_n11795_ = ng666 & new_n8969_;
  assign new_n11796_ = ~ng679 & new_n11795_;
  assign new_n11797_ = ng679 & ~new_n11795_;
  assign new_n11798_ = ~new_n11796_ & ~new_n11797_;
  assign n4907 = ~new_n5380_ & ~new_n11798_;
  assign new_n11800_ = ~ng704 & ~new_n5399_;
  assign new_n11801_ = ng653 & new_n5399_;
  assign n4912 = ~new_n11800_ & ~new_n11801_;
  assign new_n11803_ = ~ng718 & ~new_n5391_;
  assign new_n11804_ = ng666 & new_n5391_;
  assign n4917 = ~new_n11803_ & ~new_n11804_;
  assign new_n11806_ = ng630 & ng1309;
  assign new_n11807_ = ~ng729 & ~new_n11806_;
  assign new_n11808_ = ~new_n5302_1_ & new_n11806_;
  assign n4922 = ~new_n11807_ & ~new_n11808_;
  assign new_n11810_ = ~ng732 & ~new_n11806_;
  assign new_n11811_ = ~new_n5287_1_ & new_n11806_;
  assign n4927 = ~new_n11810_ & ~new_n11811_;
  assign new_n11813_ = ~ng834 & ~new_n4777_1_;
  assign new_n11814_ = ng797 & new_n4777_1_;
  assign n4937 = ~new_n11813_ & ~new_n11814_;
  assign new_n11816_ = ~ng845 & ~new_n5517_1_;
  assign new_n11817_ = ng813 & new_n5517_1_;
  assign n4942 = ~new_n11816_ & ~new_n11817_;
  assign new_n11819_ = ng797 & ~new_n5839_;
  assign new_n11820_ = ~new_n5841_ & ~new_n11819_;
  assign new_n11821_ = ~new_n5838_1_ & new_n11820_;
  assign new_n11822_ = new_n5864_ & ~new_n5870_;
  assign new_n11823_ = new_n5571_ & new_n11822_;
  assign new_n11824_ = ~new_n5571_ & ~new_n11822_;
  assign new_n11825_ = ~new_n11823_ & ~new_n11824_;
  assign new_n11826_ = new_n5838_1_ & new_n11825_;
  assign new_n11827_ = ~new_n11821_ & ~new_n11826_;
  assign new_n11828_ = ng826 & ~new_n11827_;
  assign new_n11829_ = ~ng826 & ~ng927;
  assign n4947 = ~new_n11828_ & ~new_n11829_;
  assign new_n11831_ = ng853 & ~new_n8483_;
  assign new_n11832_ = ~ng853 & ~ng906;
  assign n4952 = ~new_n11831_ & ~new_n11832_;
  assign new_n11834_ = ng776 & ~new_n5911_;
  assign new_n11835_ = ~ng776 & new_n5911_;
  assign new_n11836_ = ~new_n11834_ & ~new_n11835_;
  assign n4957 = ~new_n5127_1_ & ~new_n11836_;
  assign new_n11838_ = ~ng1033 & ~new_n8502_;
  assign new_n11839_ = ~ng1075 & ng823;
  assign new_n11840_ = ~ng1078 & ng853;
  assign new_n11841_ = ~ng1085 & ng826;
  assign new_n11842_ = ~new_n11839_ & ~new_n11840_;
  assign new_n11843_ = ~new_n11841_ & new_n11842_;
  assign new_n11844_ = pg3229 & ~new_n5932_;
  assign new_n11845_ = new_n5942_ & new_n11843_;
  assign new_n11846_ = new_n11844_ & new_n11845_;
  assign new_n11847_ = ~new_n5937_ & new_n11844_;
  assign new_n11848_ = ~new_n11846_ & ~new_n11847_;
  assign new_n11849_ = ~new_n5932_ & new_n11843_;
  assign new_n11850_ = ~pg3229 & new_n11849_;
  assign new_n11851_ = ~pg3229 & new_n11243_;
  assign new_n11852_ = pg3229 & ~new_n11843_;
  assign new_n11853_ = ~new_n11850_ & ~new_n11851_;
  assign new_n11854_ = ~new_n11852_ & new_n11853_;
  assign new_n11855_ = new_n11848_ & new_n11854_;
  assign new_n11856_ = new_n8502_ & ~new_n11855_;
  assign n4962 = ~new_n11838_ & ~new_n11856_;
  assign new_n11858_ = ~ng1048 & ~new_n8502_;
  assign new_n11859_ = new_n8502_ & ~new_n11245_;
  assign n4967 = ~new_n11858_ & ~new_n11859_;
  assign new_n11861_ = ~new_n5955_ & ~new_n5969_;
  assign new_n11862_ = n953 & ~new_n11861_;
  assign new_n11863_ = ~new_n5827_ & new_n5955_;
  assign new_n11864_ = new_n5969_ & ~new_n11863_;
  assign new_n11865_ = ~n953 & ~new_n11864_;
  assign new_n11866_ = ~new_n11862_ & ~new_n11865_;
  assign new_n11867_ = ~new_n5978_ & new_n11866_;
  assign new_n11868_ = new_n5827_ & new_n5969_;
  assign new_n11869_ = ~n953 & ~new_n11868_;
  assign new_n11870_ = ~n953 & ~new_n11869_;
  assign new_n11871_ = new_n5978_ & new_n11870_;
  assign new_n11872_ = ~new_n11867_ & ~new_n11871_;
  assign new_n11873_ = ng2384 & ~new_n11872_;
  assign new_n11874_ = n953 & new_n11873_;
  assign new_n11875_ = n953 & ~new_n11874_;
  assign new_n11876_ = new_n11873_ & ~new_n11874_;
  assign new_n11877_ = ~new_n11875_ & ~new_n11876_;
  assign new_n11878_ = ng823 & new_n11877_;
  assign new_n11879_ = ~ng1107 & ~ng823;
  assign n4972 = ~new_n11878_ & ~new_n11879_;
  assign new_n11881_ = ng826 & ~new_n8547_;
  assign new_n11882_ = ~ng1135 & ~new_n11881_;
  assign new_n11883_ = new_n8540_ & new_n11881_;
  assign n4977 = ~new_n11882_ & ~new_n11883_;
  assign new_n11885_ = new_n5551_ & new_n5556_1_;
  assign new_n11886_ = new_n5556_1_ & ~new_n5710_;
  assign new_n11887_ = ng2384 & ~new_n5675_;
  assign new_n11888_ = new_n11886_ & new_n11887_;
  assign new_n11889_ = new_n5546_ & ~new_n11888_;
  assign new_n11890_ = new_n5556_1_ & ~new_n9924_;
  assign new_n11891_ = ~new_n5710_ & ~new_n7935_;
  assign new_n11892_ = ~new_n5675_ & new_n11891_;
  assign new_n11893_ = ~new_n5556_1_ & ~new_n11892_;
  assign new_n11894_ = ~new_n11890_ & ~new_n11893_;
  assign new_n11895_ = ~new_n5546_ & new_n11894_;
  assign new_n11896_ = ~new_n11889_ & ~new_n11895_;
  assign new_n11897_ = ~new_n5551_ & new_n11896_;
  assign new_n11898_ = ~new_n11885_ & ~new_n11897_;
  assign new_n11899_ = ~new_n5556_1_ & new_n11898_;
  assign new_n11900_ = ~new_n5556_1_ & ~new_n11899_;
  assign new_n11901_ = new_n11898_ & ~new_n11899_;
  assign new_n11902_ = ~new_n11900_ & ~new_n11901_;
  assign new_n11903_ = ~new_n5836_ & ~new_n11902_;
  assign new_n11904_ = ng853 & ~new_n11903_;
  assign new_n11905_ = ~ng853 & ~ng1007;
  assign n4982 = ~new_n11904_ & ~new_n11905_;
  assign new_n11907_ = ~ng1315 & ~ng1240;
  assign n4997 = ~new_n7709_ & ~new_n11907_;
  assign new_n11909_ = ng823 & ~new_n5824_;
  assign new_n11910_ = ~ng1165 & ~ng823;
  assign n5007 = ~new_n11909_ & ~new_n11910_;
  assign new_n11912_ = ng1315 & ~ng1165;
  assign new_n11913_ = ng1309 & ~ng1166;
  assign new_n11914_ = ng1312 & ~ng1164;
  assign new_n11915_ = ~new_n11912_ & ~new_n11913_;
  assign n5012 = ~new_n11914_ & new_n11915_;
  assign new_n11917_ = ~ng1266 & ~new_n8012_;
  assign new_n11918_ = new_n8012_ & ~new_n9056_;
  assign n5017 = ~new_n11917_ & ~new_n11918_;
  assign new_n11920_ = ~ng1315 & ~ng1345;
  assign n5027 = ~new_n9359_ & ~new_n11920_;
  assign new_n11922_ = ~ng1385 & ~new_n6259_1_;
  assign new_n11923_ = ng1326 & new_n6259_1_;
  assign n5032 = ~new_n11922_ & ~new_n11923_;
  assign new_n11925_ = ~ng1393 & ~new_n6263_;
  assign new_n11926_ = ng1332 & new_n6263_;
  assign n5037 = ~new_n11925_ & ~new_n11926_;
  assign new_n11928_ = ~ng1421 & ~new_n6259_1_;
  assign new_n11929_ = new_n6259_1_ & ~new_n8694_;
  assign n5042 = ~new_n11928_ & ~new_n11929_;
  assign new_n11931_ = ~ng1514 & ~new_n4773_;
  assign new_n11932_ = ng1476 & new_n4773_;
  assign n5047 = ~new_n11931_ & ~new_n11932_;
  assign new_n11934_ = ~ng1553 & ~new_n8121_;
  assign new_n11935_ = ng1476 & new_n8121_;
  assign n5052 = ~new_n11934_ & ~new_n11935_;
  assign new_n11937_ = ng1476 & ~new_n6587_;
  assign new_n11938_ = ~new_n10383_ & ~new_n11937_;
  assign new_n11939_ = ~new_n6586_ & new_n11938_;
  assign new_n11940_ = ~new_n6319_1_ & ~new_n6599_;
  assign new_n11941_ = new_n6319_1_ & new_n6599_;
  assign new_n11942_ = ~new_n11940_ & ~new_n11941_;
  assign new_n11943_ = new_n6586_ & new_n11942_;
  assign new_n11944_ = ~new_n11939_ & ~new_n11943_;
  assign new_n11945_ = ng823 & ~new_n11944_;
  assign new_n11946_ = ~ng1615 & ~ng823;
  assign n5057 = ~new_n11945_ & ~new_n11946_;
  assign new_n11948_ = ng826 & ~new_n11295_;
  assign new_n11949_ = ~ng826 & ~ng1630;
  assign n5062 = ~new_n11948_ & ~new_n11949_;
  assign new_n11951_ = ~new_n6436_ & ~new_n6587_;
  assign new_n11952_ = ~new_n10383_ & ~new_n11951_;
  assign new_n11953_ = ~new_n6586_ & new_n11952_;
  assign new_n11954_ = ~new_n6360_ & ~new_n10924_;
  assign new_n11955_ = new_n6360_ & new_n10924_;
  assign new_n11956_ = ~new_n11954_ & ~new_n11955_;
  assign new_n11957_ = new_n6586_ & new_n11956_;
  assign new_n11958_ = ~new_n11953_ & ~new_n11957_;
  assign new_n11959_ = ng853 & ~new_n11958_;
  assign new_n11960_ = ~ng853 & ~ng1609;
  assign n5067 = ~new_n11959_ & ~new_n11960_;
  assign new_n11962_ = ng823 & ~new_n9102_;
  assign new_n11963_ = ~ng1813 & ~ng823;
  assign n5072 = ~new_n11962_ & ~new_n11963_;
  assign new_n11965_ = ~ng2224 & ~new_n5517_1_;
  assign new_n11966_ = ng2185 & new_n5517_1_;
  assign n5097 = ~new_n11965_ & ~new_n11966_;
  assign new_n11968_ = ~ng2232 & ~new_n4773_;
  assign new_n11969_ = ng2200 & new_n4773_;
  assign n5102 = ~new_n11968_ & ~new_n11969_;
  assign new_n11971_ = ng2156 & ~new_n7395_;
  assign new_n11972_ = ~ng2156 & new_n7395_;
  assign new_n11973_ = ~new_n11971_ & ~new_n11972_;
  assign n5107 = ~new_n5127_1_ & ~new_n11973_;
  assign new_n11975_ = ng853 & ~new_n11322_;
  assign new_n11976_ = ~ng853 & ~ng2510;
  assign n5112 = ~new_n11975_ & ~new_n11976_;
  assign new_n11978_ = new_n7030_ & new_n7040_;
  assign new_n11979_ = new_n7035_ & ~new_n11978_;
  assign new_n11980_ = new_n7305_ & new_n8187_;
  assign new_n11981_ = new_n8184_ & ~new_n11980_;
  assign new_n11982_ = ~new_n7159_ & new_n11981_;
  assign new_n11983_ = new_n7040_ & new_n11982_;
  assign new_n11984_ = ~new_n7309_1_ & ~new_n7311_;
  assign new_n11985_ = ~new_n7040_ & new_n11984_;
  assign new_n11986_ = ~new_n11983_ & ~new_n11985_;
  assign new_n11987_ = new_n7030_ & new_n11986_;
  assign new_n11988_ = ~new_n7159_ & new_n8187_;
  assign new_n11989_ = ~new_n7194_ & ~new_n11988_;
  assign new_n11990_ = new_n7040_ & new_n11989_;
  assign new_n11991_ = ~new_n7040_ & ~new_n7194_;
  assign new_n11992_ = ~new_n11990_ & ~new_n11991_;
  assign new_n11993_ = ~new_n7030_ & new_n11992_;
  assign new_n11994_ = ~new_n11987_ & ~new_n11993_;
  assign new_n11995_ = ~new_n7035_ & new_n11994_;
  assign new_n11996_ = ~new_n11979_ & ~new_n11995_;
  assign new_n11997_ = ~new_n7030_ & new_n11996_;
  assign new_n11998_ = ~new_n7030_ & ~new_n11997_;
  assign new_n11999_ = new_n11996_ & ~new_n11997_;
  assign new_n12000_ = ~new_n11998_ & ~new_n11999_;
  assign new_n12001_ = ~new_n7320_ & new_n12000_;
  assign new_n12002_ = ng823 & ~new_n12001_;
  assign new_n12003_ = ~ng2391 & ~ng823;
  assign n5117 = ~new_n12002_ & ~new_n12003_;
  assign new_n12005_ = ng826 & n2815;
  assign new_n12006_ = ~ng826 & ~ng2555;
  assign n5137 = ~new_n12005_ & ~new_n12006_;
  assign new_n12008_ = ng826 & ~new_n7044_;
  assign new_n12009_ = ~ng826 & ~ng2540;
  assign n5142 = ~new_n12008_ & ~new_n12009_;
  assign new_n12011_ = ng1315 & ~ng2562;
  assign new_n12012_ = ~ng2563 & ng1309;
  assign new_n12013_ = ng1312 & ~ng2561;
  assign new_n12014_ = ~new_n12011_ & ~new_n12012_;
  assign n5147 = ~new_n12013_ & new_n12014_;
  assign new_n12016_ = ~new_n5366_ & ~new_n10520_;
  assign new_n12017_ = ng1309 & ~new_n12016_;
  assign new_n12018_ = ~ng1309 & ~ng2661;
  assign n5152 = ~new_n12017_ & ~new_n12018_;
  assign new_n12020_ = ng1315 & ~new_n11359_;
  assign new_n12021_ = ~ng1315 & ~ng2685;
  assign n5157 = ~new_n12020_ & ~new_n12021_;
  assign new_n12023_ = ~ng2746 & new_n10591_;
  assign new_n12024_ = ng2746 & ~new_n10591_;
  assign new_n12025_ = ~new_n12023_ & ~new_n12024_;
  assign n5167 = ~new_n8213_ & ~new_n12025_;
  assign new_n12027_ = ~ng2779 & ~new_n7592_;
  assign new_n12028_ = ng2727 & new_n7592_;
  assign n5172 = ~new_n12027_ & ~new_n12028_;
  assign new_n12030_ = ~ng2787 & ~new_n7584_;
  assign new_n12031_ = ng2746 & new_n7584_;
  assign n5177 = ~new_n12030_ & ~new_n12031_;
  assign new_n12033_ = ~ng2801 & ~new_n7588_;
  assign new_n12034_ = ng2766 & new_n7588_;
  assign n5182 = ~new_n12033_ & ~new_n12034_;
  assign n5187 = ~pg3234 & ng3080;
  assign new_n12037_ = ~ng1217 & new_n11015_;
  assign new_n12038_ = ~new_n11139_ & new_n12037_;
  assign new_n12039_ = new_n11075_ & new_n11139_;
  assign new_n12040_ = ~new_n12038_ & ~new_n12039_;
  assign new_n12041_ = ~new_n11141_ & new_n12040_;
  assign n5192 = new_n11667_ | new_n12041_;
  assign new_n12043_ = ~ng1913 & new_n10635_;
  assign new_n12044_ = ~new_n10633_ & new_n12043_;
  assign new_n12045_ = ~new_n10698_ & ~new_n10708_;
  assign new_n12046_ = ~new_n6785_ & ~new_n12045_;
  assign new_n12047_ = ~new_n12045_ & ~new_n12046_;
  assign new_n12048_ = ~new_n6785_ & ~new_n12046_;
  assign new_n12049_ = ~new_n12047_ & ~new_n12048_;
  assign new_n12050_ = new_n10635_ & ~new_n12049_;
  assign new_n12051_ = ng1880 & new_n12050_;
  assign new_n12052_ = new_n10633_ & new_n12051_;
  assign new_n12053_ = ~new_n12044_ & ~new_n12052_;
  assign new_n12054_ = ~new_n10631_ & new_n12053_;
  assign new_n12055_ = ~new_n10635_ & new_n10719_;
  assign new_n12056_ = new_n10631_ & new_n12055_;
  assign n5197 = new_n12054_ | new_n12056_;
  assign new_n12058_ = ~ng2610 & new_n10738_;
  assign new_n12059_ = ~new_n10736_ & new_n12058_;
  assign new_n12060_ = ~new_n8246_ & ~new_n10756_;
  assign new_n12061_ = ~new_n7529_ & ~new_n12060_;
  assign new_n12062_ = ~new_n12060_ & ~new_n12061_;
  assign new_n12063_ = ~new_n7529_ & ~new_n12061_;
  assign new_n12064_ = ~new_n12062_ & ~new_n12063_;
  assign new_n12065_ = new_n10738_ & ~new_n12064_;
  assign new_n12066_ = ng2574 & new_n12065_;
  assign new_n12067_ = new_n10736_ & new_n12066_;
  assign new_n12068_ = ~new_n12059_ & ~new_n12067_;
  assign new_n12069_ = ~new_n10734_ & new_n12068_;
  assign new_n12070_ = ~new_n8286_ & ~new_n10756_;
  assign new_n12071_ = ~new_n7529_ & ~new_n12070_;
  assign new_n12072_ = ~new_n12070_ & ~new_n12071_;
  assign new_n12073_ = ~new_n7529_ & ~new_n12071_;
  assign new_n12074_ = ~new_n12072_ & ~new_n12073_;
  assign new_n12075_ = new_n10738_ & ~new_n12074_;
  assign new_n12076_ = ng2574 & new_n12075_;
  assign new_n12077_ = new_n10767_ & ~new_n12076_;
  assign new_n12078_ = new_n10734_ & new_n12077_;
  assign n5202 = new_n12069_ | new_n12078_;
  assign new_n12080_ = ~ng3028 & ng3018;
  assign new_n12081_ = new_n10779_ & new_n12080_;
  assign new_n12082_ = ng3032 & new_n12081_;
  assign new_n12083_ = ~ng3036 & new_n12082_;
  assign new_n12084_ = ~pg3234 & ~new_n12083_;
  assign new_n12085_ = ng3018 & new_n10779_;
  assign new_n12086_ = ng3028 & ~new_n12085_;
  assign new_n12087_ = ~ng3028 & new_n12085_;
  assign new_n12088_ = ~new_n12086_ & ~new_n12087_;
  assign n5207 = new_n12084_ & ~new_n12088_;
  assign new_n12090_ = ng2987 & ~ng3070;
  assign new_n12091_ = ~ng3051 & ~ng2987;
  assign n5217 = ~new_n12090_ & ~new_n12091_;
  assign new_n12093_ = ng2987 & ~ng2997;
  assign new_n12094_ = ~ng3061 & ~ng2987;
  assign n5222 = ~new_n12093_ & ~new_n12094_;
  assign n5227 = ~pg51 & ng2817;
  assign new_n12097_ = ng1315 & ~n1448;
  assign new_n12098_ = ~ng1315 & ~ng3102;
  assign n5232 = ~new_n12097_ & ~new_n12098_;
  assign new_n12100_ = ng1315 & ~ng499;
  assign new_n12101_ = ~ng1315 & ~ng3161;
  assign n5237 = ~new_n12100_ & ~new_n12101_;
  assign new_n12103_ = ~ng132 & ~new_n4773_;
  assign new_n12104_ = ng101 & new_n4773_;
  assign n5242 = ~new_n12103_ & ~new_n12104_;
  assign new_n12106_ = ~ng147 & ~new_n4773_;
  assign new_n12107_ = ng113 & new_n4773_;
  assign n5247 = ~new_n12106_ & ~new_n12107_;
  assign new_n12109_ = ~ng163 & ~new_n5517_1_;
  assign new_n12110_ = ~new_n4891_ & new_n5517_1_;
  assign n5252 = ~new_n12109_ & ~new_n12110_;
  assign new_n12112_ = ~ng175 & ~new_n5538_;
  assign new_n12113_ = ng97 & new_n5538_;
  assign n5257 = ~new_n12112_ & ~new_n12113_;
  assign new_n12115_ = ~ng177 & ~new_n8121_;
  assign new_n12116_ = new_n5180_ & new_n8121_;
  assign n5262 = ~new_n12115_ & ~new_n12116_;
  assign new_n12118_ = ng853 & ~new_n9260_;
  assign new_n12119_ = ~ng853 & ~ng201;
  assign n5267 = ~new_n12118_ & ~new_n12119_;
  assign new_n12121_ = ng853 & ~new_n8929_;
  assign new_n12122_ = ~ng853 & ~ng228;
  assign n5272 = ~new_n12121_ & ~new_n12122_;
  assign new_n12124_ = ng70 & ~new_n9290_;
  assign new_n12125_ = ~ng70 & new_n9290_;
  assign new_n12126_ = ~new_n12124_ & ~new_n12125_;
  assign n5277 = ~new_n5127_1_ & ~new_n12126_;
  assign new_n12128_ = ~new_n5182_1_ & ~new_n5187_1_;
  assign new_n12129_ = n4167 & ~new_n12128_;
  assign new_n12130_ = ~new_n5071_ & new_n5187_1_;
  assign new_n12131_ = new_n5182_1_ & ~new_n12130_;
  assign new_n12132_ = ~n4167 & ~new_n12131_;
  assign new_n12133_ = ~new_n12129_ & ~new_n12132_;
  assign new_n12134_ = ~new_n5168_ & new_n12133_;
  assign new_n12135_ = new_n5071_ & new_n5182_1_;
  assign new_n12136_ = ~n4167 & ~new_n12135_;
  assign new_n12137_ = ~n4167 & ~new_n12136_;
  assign new_n12138_ = new_n5168_ & new_n12137_;
  assign new_n12139_ = ~new_n12134_ & ~new_n12138_;
  assign new_n12140_ = ng2384 & ~new_n12139_;
  assign new_n12141_ = n4167 & new_n12140_;
  assign new_n12142_ = n4167 & ~new_n12141_;
  assign new_n12143_ = new_n12140_ & ~new_n12141_;
  assign new_n12144_ = ~new_n12142_ & ~new_n12143_;
  assign new_n12145_ = ng853 & new_n12144_;
  assign new_n12146_ = ~ng853 & ~ng423;
  assign n5282 = ~new_n12145_ & ~new_n12146_;
  assign new_n12148_ = ng823 & ~new_n11759_;
  assign new_n12149_ = ~ng432 & ~ng823;
  assign n5287 = ~new_n12148_ & ~new_n12149_;
  assign new_n12151_ = ng823 & ~new_n11213_;
  assign new_n12152_ = ~ng313 & ~ng823;
  assign n5292 = ~new_n12151_ & ~new_n12152_;
  assign new_n12154_ = ~ng402 & ~new_n9505_;
  assign new_n12155_ = new_n9505_ & new_n11767_;
  assign n5297 = ~new_n12154_ & ~new_n12155_;
  assign new_n12157_ = ng853 & ~new_n5068_;
  assign new_n12158_ = ~ng853 & ~ng479;
  assign n5321 = ~new_n12157_ & ~new_n12158_;
  assign new_n12160_ = ng823 & ~new_n4799_;
  assign new_n12161_ = ~ng468 & ~ng823;
  assign n5326 = ~new_n12160_ & ~new_n12161_;
  assign new_n12163_ = ~ng586 & ~new_n7715_;
  assign new_n12164_ = new_n7715_ & ~new_n8439_;
  assign n5335 = ~new_n12163_ & ~new_n12164_;
  assign new_n12166_ = ng1312 & ~new_n11791_;
  assign new_n12167_ = ~ng1312 & ~ng617;
  assign n5340 = ~new_n12166_ & ~new_n12167_;
  assign new_n12169_ = ng679 & new_n11795_;
  assign new_n12170_ = ng686 & ~new_n12169_;
  assign new_n12171_ = ~ng686 & new_n12169_;
  assign new_n12172_ = ~new_n12170_ & ~new_n12171_;
  assign n5345 = ~new_n5380_ & ~new_n12172_;
  assign new_n12174_ = ~ng706 & ~new_n5391_;
  assign new_n12175_ = ng653 & new_n5391_;
  assign n5350 = ~new_n12174_ & ~new_n12175_;
  assign new_n12177_ = ~ng716 & ~new_n5399_;
  assign new_n12178_ = ng666 & new_n5399_;
  assign n5355 = ~new_n12177_ & ~new_n12178_;
  assign new_n12180_ = ~ng725 & ~new_n5399_;
  assign new_n12181_ = ng692 & new_n5399_;
  assign n5360 = ~new_n12180_ & ~new_n12181_;
  assign new_n12183_ = ~ng733 & ~new_n5380_;
  assign new_n12184_ = ~new_n5287_1_ & new_n5380_;
  assign n5365 = ~new_n12183_ & ~new_n12184_;
  assign new_n12186_ = ~ng832 & ~new_n4773_;
  assign new_n12187_ = ng797 & new_n4773_;
  assign n5373 = ~new_n12186_ & ~new_n12187_;
  assign new_n12189_ = ~ng841 & ~new_n4773_;
  assign new_n12190_ = ng809 & new_n4773_;
  assign n5378 = ~new_n12189_ & ~new_n12190_;
  assign new_n12192_ = ng823 & ~new_n11827_;
  assign new_n12193_ = ~ng823 & ~ng930;
  assign n5383 = ~new_n12192_ & ~new_n12193_;
  assign new_n12195_ = ng823 & ~new_n8483_;
  assign new_n12196_ = ~ng823 & ~ng903;
  assign n5388 = ~new_n12195_ & ~new_n12196_;
  assign new_n12198_ = ~ng771 & new_n5912_;
  assign new_n12199_ = ng771 & ~new_n5912_;
  assign new_n12200_ = ~new_n12198_ & ~new_n12199_;
  assign n5393 = ~new_n5127_1_ & ~new_n12200_;
  assign new_n12202_ = ~ng1030 & ~new_n7915_;
  assign new_n12203_ = new_n7915_ & ~new_n11855_;
  assign n5398 = ~new_n12202_ & ~new_n12203_;
  assign new_n12205_ = ~ng1071 & ~new_n5926_;
  assign new_n12206_ = ~pg3229 & new_n5932_;
  assign new_n12207_ = new_n11845_ & new_n12206_;
  assign new_n12208_ = ~new_n11846_ & ~new_n12207_;
  assign new_n12209_ = ~new_n5932_ & ~new_n5942_;
  assign new_n12210_ = ~pg3229 & new_n12209_;
  assign new_n12211_ = new_n5932_ & ~new_n5942_;
  assign new_n12212_ = pg3229 & new_n12211_;
  assign new_n12213_ = ~new_n12210_ & ~new_n12212_;
  assign new_n12214_ = new_n12208_ & new_n12213_;
  assign new_n12215_ = new_n5926_ & ~new_n12214_;
  assign n5403 = ~new_n12205_ & ~new_n12215_;
  assign new_n12217_ = ng826 & new_n11877_;
  assign new_n12218_ = ~ng826 & ~ng1104;
  assign n5408 = ~new_n12217_ & ~new_n12218_;
  assign new_n12220_ = ng823 & ~new_n8547_;
  assign new_n12221_ = ~ng1136 & ~new_n12220_;
  assign new_n12222_ = new_n8540_ & new_n12220_;
  assign n5413 = ~new_n12221_ & ~new_n12222_;
  assign new_n12224_ = ng823 & ~new_n11903_;
  assign new_n12225_ = ~ng823 & ~ng1006;
  assign n5418 = ~new_n12224_ & ~new_n12225_;
  assign new_n12227_ = ng1315 & ng1240;
  assign new_n12228_ = ~ng1315 & ~ng1243;
  assign n5431 = ~new_n12227_ & ~new_n12228_;
  assign new_n12230_ = ~ng1265 & ~new_n8562_;
  assign new_n12231_ = new_n8562_ & ~new_n9056_;
  assign n5448 = ~new_n12230_ & ~new_n12231_;
  assign new_n12233_ = ng1315 & ~ng1196;
  assign new_n12234_ = ~ng1315 & ~ng1316;
  assign n5458 = ~new_n12233_ & ~new_n12234_;
  assign new_n12236_ = ~ng1386 & ~new_n6255_;
  assign new_n12237_ = ng1326 & new_n6255_;
  assign n5463 = ~new_n12236_ & ~new_n12237_;
  assign new_n12239_ = ~ng1395 & ~new_n6255_;
  assign new_n12240_ = ng1332 & new_n6255_;
  assign n5468 = ~new_n12239_ & ~new_n12240_;
  assign new_n12242_ = ~ng1422 & ~new_n6255_;
  assign new_n12243_ = new_n6255_ & ~new_n8694_;
  assign n5473 = ~new_n12242_ & ~new_n12243_;
  assign new_n12245_ = ~ng1516 & ~new_n4777_1_;
  assign new_n12246_ = ng1476 & new_n4777_1_;
  assign n5478 = ~new_n12245_ & ~new_n12246_;
  assign new_n12248_ = ~ng1557 & ~new_n5538_;
  assign new_n12249_ = ng1471 & new_n5538_;
  assign n5483 = ~new_n12248_ & ~new_n12249_;
  assign new_n12251_ = ng826 & ~new_n11944_;
  assign new_n12252_ = ~ng826 & ~ng1612;
  assign n5488 = ~new_n12251_ & ~new_n12252_;
  assign new_n12254_ = ng823 & ~new_n11295_;
  assign new_n12255_ = ~ng823 & ~ng1633;
  assign n5493 = ~new_n12254_ & ~new_n12255_;
  assign new_n12257_ = ng823 & ~new_n11958_;
  assign new_n12258_ = ~ng823 & ~ng1606;
  assign n5498 = ~new_n12257_ & ~new_n12258_;
  assign new_n12260_ = ng826 & new_n8757_;
  assign new_n12261_ = ~ng826 & ~ng1789;
  assign n5503 = ~new_n12260_ & ~new_n12261_;
  assign new_n12263_ = ~ng2225 & ~new_n4777_1_;
  assign new_n12264_ = ng2185 & new_n4777_1_;
  assign n5526 = ~new_n12263_ & ~new_n12264_;
  assign new_n12266_ = ~ng2234 & ~new_n4777_1_;
  assign new_n12267_ = ng2200 & new_n4777_1_;
  assign n5531 = ~new_n12266_ & ~new_n12267_;
  assign new_n12269_ = ng2384 & ~new_n7484_;
  assign new_n12270_ = ~new_n7505_ & new_n12269_;
  assign new_n12271_ = ~new_n7489_ & new_n12270_;
  assign new_n12272_ = ~new_n7489_ & ~new_n12271_;
  assign new_n12273_ = new_n12270_ & ~new_n12271_;
  assign new_n12274_ = ~new_n12272_ & ~new_n12273_;
  assign new_n12275_ = ng826 & new_n12274_;
  assign new_n12276_ = ~ng826 & ~ng2513;
  assign n5540 = ~new_n12275_ & ~new_n12276_;
  assign new_n12278_ = ng826 & ~new_n12001_;
  assign new_n12279_ = ~ng826 & ~ng2390;
  assign n5545 = ~new_n12278_ & ~new_n12279_;
  assign new_n12281_ = ng853 & ~new_n7308_;
  assign new_n12282_ = ~ng853 & ~ng2554;
  assign n5561 = ~new_n12281_ & ~new_n12282_;
  assign new_n12284_ = ng823 & ~new_n7044_;
  assign new_n12285_ = ~ng823 & ~ng2543;
  assign n5566 = ~new_n12284_ & ~new_n12285_;
  assign new_n12287_ = ng1312 & ~new_n12016_;
  assign new_n12288_ = ~ng1312 & ~ng2664;
  assign n5575 = ~new_n12287_ & ~new_n12288_;
  assign new_n12290_ = ng1312 & ~new_n11359_;
  assign new_n12291_ = ~ng1312 & ~ng2682;
  assign n5580 = ~new_n12290_ & ~new_n12291_;
  assign new_n12293_ = ~ng2707 & new_n8215_;
  assign new_n12294_ = ng2707 & ~new_n8215_;
  assign new_n12295_ = ~new_n12293_ & ~new_n12294_;
  assign n5585 = ~new_n8213_ & ~new_n12295_;
  assign new_n12297_ = ng2740 & ~new_n10592_;
  assign new_n12298_ = ~ng2740 & new_n10592_;
  assign new_n12299_ = ~new_n12297_ & ~new_n12298_;
  assign n5590 = ~new_n8213_ & ~new_n12299_;
  assign new_n12301_ = ~ng2775 & ~new_n7584_;
  assign new_n12302_ = ng2707 & new_n7584_;
  assign n5595 = ~new_n12301_ & ~new_n12302_;
  assign new_n12304_ = ~ng2791 & ~new_n7592_;
  assign new_n12305_ = ng2740 & new_n7592_;
  assign n5600 = ~new_n12304_ & ~new_n12305_;
  assign new_n12307_ = ~ng2800 & ~new_n7592_;
  assign new_n12308_ = ng2766 & new_n7592_;
  assign n5605 = ~new_n12307_ & ~new_n12308_;
  assign new_n12310_ = ~ng2802 & ~new_n7596_;
  assign new_n12311_ = ~new_n7540_ & new_n7596_;
  assign n5610 = ~new_n12310_ & ~new_n12311_;
  assign new_n12313_ = ~ng1218 & new_n11015_;
  assign new_n12314_ = ~new_n11139_ & new_n12313_;
  assign new_n12315_ = new_n11082_ & new_n11139_;
  assign new_n12316_ = ~new_n12314_ & ~new_n12315_;
  assign new_n12317_ = ~new_n11141_ & new_n12316_;
  assign n5615 = new_n11391_ | new_n12317_;
  assign new_n12319_ = ~ng1912 & new_n10635_;
  assign new_n12320_ = ~new_n10633_ & new_n12319_;
  assign new_n12321_ = ~new_n10676_ & ~new_n10708_;
  assign new_n12322_ = ~new_n6796_ & ~new_n12321_;
  assign new_n12323_ = ~new_n12321_ & ~new_n12322_;
  assign new_n12324_ = ~new_n6796_ & ~new_n12322_;
  assign new_n12325_ = ~new_n12323_ & ~new_n12324_;
  assign new_n12326_ = new_n10635_ & ~new_n12325_;
  assign new_n12327_ = ng1880 & new_n12326_;
  assign new_n12328_ = new_n10633_ & new_n12327_;
  assign new_n12329_ = ~new_n12320_ & ~new_n12328_;
  assign new_n12330_ = ~new_n10631_ & new_n12329_;
  assign n5620 = new_n10729_ | new_n12330_;
  assign new_n12332_ = ~ng2611 & new_n10738_;
  assign new_n12333_ = ~new_n10736_ & new_n12332_;
  assign new_n12334_ = ~new_n8264_ & ~new_n10756_;
  assign new_n12335_ = ~new_n7540_ & ~new_n12334_;
  assign new_n12336_ = ~new_n12334_ & ~new_n12335_;
  assign new_n12337_ = ~new_n7540_ & ~new_n12335_;
  assign new_n12338_ = ~new_n12336_ & ~new_n12337_;
  assign new_n12339_ = new_n10738_ & ~new_n12338_;
  assign new_n12340_ = ng2574 & new_n12339_;
  assign new_n12341_ = new_n10736_ & new_n12340_;
  assign new_n12342_ = ~new_n12333_ & ~new_n12341_;
  assign new_n12343_ = ~new_n10734_ & new_n12342_;
  assign new_n12344_ = ~new_n8324_ & ~new_n10756_;
  assign new_n12345_ = ~new_n7540_ & ~new_n12344_;
  assign new_n12346_ = ~new_n12344_ & ~new_n12345_;
  assign new_n12347_ = ~new_n7540_ & ~new_n12345_;
  assign new_n12348_ = ~new_n12346_ & ~new_n12347_;
  assign new_n12349_ = new_n10738_ & ~new_n12348_;
  assign new_n12350_ = ng2574 & new_n12349_;
  assign new_n12351_ = new_n10767_ & ~new_n12350_;
  assign new_n12352_ = new_n10734_ & new_n12351_;
  assign n5625 = new_n12343_ | new_n12352_;
  assign new_n12354_ = ~ng3018 & new_n10779_;
  assign new_n12355_ = ng3018 & ~new_n10779_;
  assign new_n12356_ = ~new_n12354_ & ~new_n12355_;
  assign n5630 = ~new_n12084_ | ~new_n12356_;
  assign new_n12358_ = ng2987 & ~ng3069;
  assign new_n12359_ = ~ng3050 & ~ng2987;
  assign n5639 = ~new_n12358_ & ~new_n12359_;
  assign new_n12361_ = ~ng2990 & ~new_n11460_;
  assign new_n12362_ = ~new_n11460_ & ~new_n12361_;
  assign new_n12363_ = ~ng2990 & ~new_n12361_;
  assign n5644 = ~new_n12362_ & ~new_n12363_;
  assign n5649 = pg51 | ng2933;
  assign new_n12366_ = ~ng142 & ~new_n5517_1_;
  assign new_n12367_ = ng105 & new_n5517_1_;
  assign n5664 = ~new_n12366_ & ~new_n12367_;
  assign new_n12369_ = ~ng150 & ~new_n4773_;
  assign new_n12370_ = ng117 & new_n4773_;
  assign n5669 = ~new_n12369_ & ~new_n12370_;
  assign new_n12372_ = ~ng160 & ~new_n5517_1_;
  assign new_n12373_ = ~new_n4932_1_ & new_n5517_1_;
  assign n5674 = ~new_n12372_ & ~new_n12373_;
  assign new_n12375_ = ~ng171 & ~new_n8121_;
  assign new_n12376_ = ng101 & new_n8121_;
  assign n5679 = ~new_n12375_ & ~new_n12376_;
  assign new_n12378_ = ng826 & ~new_n10304_;
  assign new_n12379_ = ~ng826 & ~ng186;
  assign n5684 = ~new_n12378_ & ~new_n12379_;
  assign new_n12381_ = ng853 & ~new_n11737_;
  assign new_n12382_ = ~ng853 & ~ng246;
  assign n5689 = ~new_n12381_ & ~new_n12382_;
  assign new_n12384_ = ng826 & ~new_n9286_;
  assign new_n12385_ = ~ng826 & ~ng267;
  assign n5694 = ~new_n12384_ & ~new_n12385_;
  assign new_n12387_ = ~ng361 & ~new_n8937_;
  assign new_n12388_ = ~new_n5161_ & new_n8937_;
  assign n5699 = ~new_n12387_ & ~new_n12388_;
  assign new_n12390_ = ng823 & new_n12144_;
  assign new_n12391_ = ~ng823 & ~ng420;
  assign n5704 = ~new_n12390_ & ~new_n12391_;
  assign new_n12393_ = ng853 & ~new_n11759_;
  assign new_n12394_ = ~ng853 & ~ng435;
  assign n5709 = ~new_n12393_ & ~new_n12394_;
  assign new_n12396_ = ng823 & ~new_n7705_;
  assign new_n12397_ = ~ng823 & ~ng316;
  assign n5714 = ~new_n12396_ & ~new_n12397_;
  assign new_n12399_ = ng853 & new_n10324_;
  assign new_n12400_ = ~ng321 & ~new_n12399_;
  assign new_n12401_ = new_n10331_ & new_n12399_;
  assign n5719 = ~new_n12400_ & ~new_n12401_;
  assign new_n12403_ = ng823 & ~new_n5068_;
  assign new_n12404_ = ~ng823 & ~ng478;
  assign n5753 = ~new_n12403_ & ~new_n12404_;
  assign new_n12406_ = ng853 & ~new_n4799_;
  assign new_n12407_ = ~ng853 & ~ng471;
  assign n5758 = ~new_n12406_ & ~new_n12407_;
  assign new_n12409_ = ~ng576 & ~new_n8959_;
  assign new_n12410_ = ~new_n5341_ & new_n8959_;
  assign n5763 = ~new_n12409_ & ~new_n12410_;
  assign new_n12412_ = ~ng583 & ~new_n7715_;
  assign new_n12413_ = new_n7715_ & ~new_n10854_;
  assign n5768 = ~new_n12412_ & ~new_n12413_;
  assign new_n12415_ = ng1309 & ~new_n11791_;
  assign new_n12416_ = ~ng1309 & ~ng614;
  assign n5773 = ~new_n12415_ & ~new_n12416_;
  assign new_n12418_ = ng1312 & ~new_n5376_;
  assign new_n12419_ = ~ng1312 & ~ng493;
  assign n5778 = ~new_n12418_ & ~new_n12419_;
  assign new_n12421_ = ng686 & new_n12169_;
  assign new_n12422_ = ~ng692 & new_n12421_;
  assign new_n12423_ = ng692 & ~new_n12421_;
  assign new_n12424_ = ~new_n12422_ & ~new_n12423_;
  assign n5788 = ~new_n5380_ & ~new_n12424_;
  assign new_n12426_ = ~ng709 & ~new_n5391_;
  assign new_n12427_ = ng646 & new_n5391_;
  assign n5793 = ~new_n12426_ & ~new_n12427_;
  assign new_n12429_ = ~ng713 & ~new_n5399_;
  assign new_n12430_ = ng672 & new_n5399_;
  assign n5798 = ~new_n12429_ & ~new_n12430_;
  assign new_n12432_ = ~ng727 & ~new_n5391_;
  assign new_n12433_ = ng692 & new_n5391_;
  assign n5803 = ~new_n12432_ & ~new_n12433_;
  assign new_n12435_ = ~ng731 & ~new_n11507_;
  assign new_n12436_ = ~new_n5287_1_ & new_n11507_;
  assign n5808 = ~new_n12435_ & ~new_n12436_;
  assign new_n12438_ = ~ng819 & ~new_n4777_1_;
  assign new_n12439_ = ng785 & new_n4777_1_;
  assign n5813 = ~new_n12438_ & ~new_n12439_;
  assign new_n12441_ = ~ng829 & ~new_n4773_;
  assign new_n12442_ = ng793 & new_n4773_;
  assign n5818 = ~new_n12441_ & ~new_n12442_;
  assign new_n12444_ = ~ng843 & ~new_n4777_1_;
  assign new_n12445_ = ng809 & new_n4777_1_;
  assign n5823 = ~new_n12444_ & ~new_n12445_;
  assign new_n12447_ = ~ng864 & ~new_n6278_;
  assign new_n12448_ = ng785 & new_n6278_;
  assign n5828 = ~new_n12447_ & ~new_n12448_;
  assign new_n12450_ = ng853 & ~new_n11827_;
  assign new_n12451_ = ~ng853 & ~ng933;
  assign n5833 = ~new_n12450_ & ~new_n12451_;
  assign new_n12453_ = ng823 & ~new_n10882_;
  assign new_n12454_ = ~ng823 & ~ng948;
  assign n5838 = ~new_n12453_ & ~new_n12454_;
  assign new_n12456_ = ng853 & ~new_n5907_;
  assign new_n12457_ = ~ng853 & ~ng960;
  assign n5843 = ~new_n12456_ & ~new_n12457_;
  assign new_n12459_ = ~ng1041 & ~new_n5926_;
  assign new_n12460_ = new_n5926_ & ~new_n11855_;
  assign n5848 = ~new_n12459_ & ~new_n12460_;
  assign new_n12462_ = ~ng1060 & ~new_n7915_;
  assign new_n12463_ = new_n7915_ & ~new_n12214_;
  assign n5853 = ~new_n12462_ & ~new_n12463_;
  assign new_n12465_ = ng826 & ~new_n5984_;
  assign new_n12466_ = ~ng1114 & ~new_n12465_;
  assign new_n12467_ = new_n5981_ & new_n12465_;
  assign n5858 = ~new_n12466_ & ~new_n12467_;
  assign new_n12469_ = ng823 & new_n9393_;
  assign new_n12470_ = ~ng823 & ~ng1128;
  assign n5863 = ~new_n12469_ & ~new_n12470_;
  assign new_n12472_ = ng826 & ~new_n11903_;
  assign new_n12473_ = ~ng826 & ~ng1005;
  assign n5868 = ~new_n12472_ & ~new_n12473_;
  assign new_n12475_ = ng826 & n953;
  assign new_n12476_ = ~ng826 & ~ng1167;
  assign n5898 = ~new_n12475_ & ~new_n12476_;
  assign new_n12478_ = ~ng1261 & ~new_n6049_;
  assign new_n12479_ = new_n6049_ & ~new_n9409_;
  assign n5903 = ~new_n12478_ & ~new_n12479_;
  assign new_n12481_ = ~ng1319 & new_n6243_;
  assign new_n12482_ = ng1319 & ~new_n6243_;
  assign new_n12483_ = ~new_n12481_ & ~new_n12482_;
  assign n5913 = ~new_n6241_ & ~new_n12483_;
  assign new_n12485_ = ng1365 & new_n8030_;
  assign new_n12486_ = ng1372 & ~new_n12485_;
  assign new_n12487_ = ~ng1372 & new_n12485_;
  assign new_n12488_ = ~new_n12486_ & ~new_n12487_;
  assign n5918 = ~new_n6241_ & ~new_n12488_;
  assign new_n12490_ = ~ng1394 & ~new_n6259_1_;
  assign new_n12491_ = ng1332 & new_n6259_1_;
  assign n5923 = ~new_n12490_ & ~new_n12491_;
  assign new_n12493_ = ~ng1401 & ~new_n6255_;
  assign new_n12494_ = ng1358 & new_n6255_;
  assign n5928 = ~new_n12493_ & ~new_n12494_;
  assign new_n12496_ = ~ng1412 & ~new_n6259_1_;
  assign new_n12497_ = ng1378 & new_n6259_1_;
  assign n5933 = ~new_n12496_ & ~new_n12497_;
  assign new_n12499_ = ~ng1558 & ~new_n6278_;
  assign new_n12500_ = ng1471 & new_n6278_;
  assign n5938 = ~new_n12499_ & ~new_n12500_;
  assign new_n12502_ = ng826 & ~new_n10390_;
  assign new_n12503_ = ~ng826 & ~ng1576;
  assign n5943 = ~new_n12502_ & ~new_n12503_;
  assign new_n12505_ = ng823 & ~new_n8063_;
  assign new_n12506_ = ~ng823 & ~ng1588;
  assign n5948 = ~new_n12505_ & ~new_n12506_;
  assign new_n12508_ = ng826 & ~new_n11958_;
  assign new_n12509_ = ~ng826 & ~ng1603;
  assign n5953 = ~new_n12508_ & ~new_n12509_;
  assign new_n12511_ = ~ng1727 & ~new_n9087_;
  assign new_n12512_ = new_n9087_ & ~new_n10168_;
  assign n5958 = ~new_n12511_ & ~new_n12512_;
  assign new_n12514_ = ng1426 & new_n6326_;
  assign new_n12515_ = new_n6326_ & ~new_n12514_;
  assign new_n12516_ = ng1426 & ~new_n12514_;
  assign new_n12517_ = ~new_n12515_ & ~new_n12516_;
  assign new_n12518_ = ng1439 & new_n6353_1_;
  assign new_n12519_ = new_n6353_1_ & ~new_n12518_;
  assign new_n12520_ = ng1439 & ~new_n12518_;
  assign new_n12521_ = ~new_n12519_ & ~new_n12520_;
  assign new_n12522_ = ng1435 & new_n6331_1_;
  assign new_n12523_ = new_n6331_1_ & ~new_n12522_;
  assign new_n12524_ = ng1435 & ~new_n12522_;
  assign new_n12525_ = ~new_n12523_ & ~new_n12524_;
  assign new_n12526_ = ng1444 & new_n6341_;
  assign new_n12527_ = new_n6341_ & ~new_n12526_;
  assign new_n12528_ = ng1444 & ~new_n12526_;
  assign new_n12529_ = ~new_n12527_ & ~new_n12528_;
  assign new_n12530_ = ~new_n12521_ & ~new_n12525_;
  assign new_n12531_ = ~new_n12529_ & new_n12530_;
  assign new_n12532_ = ng1430 & new_n6360_;
  assign new_n12533_ = new_n6360_ & ~new_n12532_;
  assign new_n12534_ = ng1430 & ~new_n12532_;
  assign new_n12535_ = ~new_n12533_ & ~new_n12534_;
  assign new_n12536_ = ~new_n12517_ & new_n12531_;
  assign new_n12537_ = ~new_n12535_ & new_n12536_;
  assign new_n12538_ = ng1448 & new_n6336_1_;
  assign new_n12539_ = new_n6336_1_ & ~new_n12538_;
  assign new_n12540_ = ng1448 & ~new_n12538_;
  assign new_n12541_ = ~new_n12539_ & ~new_n12540_;
  assign new_n12542_ = ng1462 & new_n6319_1_;
  assign new_n12543_ = new_n6319_1_ & ~new_n12542_;
  assign new_n12544_ = ng1462 & ~new_n12542_;
  assign new_n12545_ = ~new_n12543_ & ~new_n12544_;
  assign new_n12546_ = ng1457 & new_n6309_1_;
  assign new_n12547_ = new_n6309_1_ & ~new_n12546_;
  assign new_n12548_ = ng1457 & ~new_n12546_;
  assign new_n12549_ = ~new_n12547_ & ~new_n12548_;
  assign new_n12550_ = ng1466 & new_n6346_;
  assign new_n12551_ = new_n6346_ & ~new_n12550_;
  assign new_n12552_ = ng1466 & ~new_n12550_;
  assign new_n12553_ = ~new_n12551_ & ~new_n12552_;
  assign new_n12554_ = ~new_n12545_ & ~new_n12549_;
  assign new_n12555_ = ~new_n12553_ & new_n12554_;
  assign new_n12556_ = ng1453 & new_n6314_1_;
  assign new_n12557_ = new_n6314_1_ & ~new_n12556_;
  assign new_n12558_ = ng1453 & ~new_n12556_;
  assign new_n12559_ = ~new_n12557_ & ~new_n12558_;
  assign new_n12560_ = ~new_n12541_ & new_n12555_;
  assign new_n12561_ = ~new_n12559_ & new_n12560_;
  assign new_n12562_ = ~new_n6634_ & new_n12537_;
  assign new_n12563_ = new_n12561_ & new_n12562_;
  assign new_n12564_ = ~new_n5125_ & new_n12563_;
  assign new_n12565_ = new_n6303_ & new_n6369_;
  assign new_n12566_ = ~new_n12564_ & ~new_n12565_;
  assign n5967 = ~new_n6635_ | new_n12566_;
  assign new_n12568_ = ~ng2448 & ~new_n9171_;
  assign new_n12569_ = ~new_n8164_ & new_n9171_;
  assign n5982 = ~new_n12568_ & ~new_n12569_;
  assign new_n12571_ = ng823 & new_n12274_;
  assign new_n12572_ = ~ng823 & ~ng2516;
  assign n5987 = ~new_n12571_ & ~new_n12572_;
  assign new_n12574_ = ng826 & ~new_n8200_;
  assign new_n12575_ = ~ng826 & ~ng2393;
  assign n5992 = ~new_n12574_ & ~new_n12575_;
  assign new_n12577_ = ng823 & ~new_n7308_;
  assign new_n12578_ = ~ng823 & ~ng2553;
  assign n6012 = ~new_n12577_ & ~new_n12578_;
  assign new_n12580_ = ng853 & ~new_n7044_;
  assign new_n12581_ = ~ng853 & ~ng2546;
  assign n6017 = ~new_n12580_ & ~new_n12581_;
  assign new_n12583_ = ~ng2650 & ~new_n9196_;
  assign new_n12584_ = ~new_n7579_ & new_n9196_;
  assign n6022 = ~new_n12583_ & ~new_n12584_;
  assign new_n12586_ = ng1315 & ~new_n12016_;
  assign new_n12587_ = ~ng1315 & ~ng2667;
  assign n6027 = ~new_n12586_ & ~new_n12587_;
  assign new_n12589_ = ng2714 & ~new_n8214_;
  assign new_n12590_ = ~ng2714 & new_n8214_;
  assign new_n12591_ = ~new_n12589_ & ~new_n12590_;
  assign n6037 = ~new_n8213_ & ~new_n12591_;
  assign new_n12593_ = ~ng2753 & new_n10593_;
  assign new_n12594_ = ng2753 & ~new_n10593_;
  assign new_n12595_ = ~new_n12593_ & ~new_n12594_;
  assign n6042 = ~new_n8213_ & ~new_n12595_;
  assign new_n12597_ = ~ng2778 & ~new_n7584_;
  assign new_n12598_ = ng2727 & new_n7584_;
  assign n6047 = ~new_n12597_ & ~new_n12598_;
  assign new_n12600_ = ~ng2788 & ~new_n7592_;
  assign new_n12601_ = ng2746 & new_n7592_;
  assign n6052 = ~new_n12600_ & ~new_n12601_;
  assign new_n12603_ = ~ng2796 & ~new_n7584_;
  assign new_n12604_ = ng2760 & new_n7584_;
  assign n6057 = ~new_n12603_ & ~new_n12604_;
  assign new_n12606_ = ~ng2806 & ~new_n11372_;
  assign new_n12607_ = ~new_n7529_ & new_n11372_;
  assign n6062 = ~new_n12606_ & ~new_n12607_;
  assign n6067 = pg3234 | ng3079;
  assign new_n12610_ = ~ng1219 & new_n11015_;
  assign new_n12611_ = ~new_n11139_ & new_n12610_;
  assign new_n12612_ = new_n11097_ & new_n11139_;
  assign new_n12613_ = ~new_n12611_ & ~new_n12612_;
  assign new_n12614_ = ~new_n11141_ & new_n12613_;
  assign new_n12615_ = ~new_n11015_ & new_n11381_;
  assign new_n12616_ = new_n11141_ & new_n12615_;
  assign n6072 = new_n12614_ | new_n12616_;
  assign new_n12618_ = ~ng1916 & new_n10635_;
  assign new_n12619_ = ~new_n10633_ & new_n12618_;
  assign new_n12620_ = ~new_n10681_ & ~new_n10708_;
  assign new_n12621_ = ~new_n6785_ & ~new_n12620_;
  assign new_n12622_ = ~new_n12620_ & ~new_n12621_;
  assign new_n12623_ = ~new_n6785_ & ~new_n12621_;
  assign new_n12624_ = ~new_n12622_ & ~new_n12623_;
  assign new_n12625_ = new_n10635_ & ~new_n12624_;
  assign new_n12626_ = ng1880 & new_n12625_;
  assign new_n12627_ = new_n10633_ & new_n12626_;
  assign new_n12628_ = ~new_n12619_ & ~new_n12627_;
  assign new_n12629_ = ~new_n10631_ & new_n12628_;
  assign new_n12630_ = ~new_n10647_ & ~new_n10708_;
  assign new_n12631_ = ~new_n6785_ & ~new_n12630_;
  assign new_n12632_ = ~new_n12630_ & ~new_n12631_;
  assign new_n12633_ = ~new_n6785_ & ~new_n12631_;
  assign new_n12634_ = ~new_n12632_ & ~new_n12633_;
  assign new_n12635_ = new_n10635_ & ~new_n12634_;
  assign new_n12636_ = ng1880 & new_n12635_;
  assign new_n12637_ = new_n10719_ & ~new_n12636_;
  assign new_n12638_ = new_n10631_ & new_n12637_;
  assign n6077 = new_n12629_ | new_n12638_;
  assign new_n12640_ = ~ng2607 & new_n10738_;
  assign new_n12641_ = ~new_n10736_ & new_n12640_;
  assign new_n12642_ = ~new_n8275_ & ~new_n10756_;
  assign new_n12643_ = ~new_n7529_ & ~new_n12642_;
  assign new_n12644_ = ~new_n12642_ & ~new_n12643_;
  assign new_n12645_ = ~new_n7529_ & ~new_n12643_;
  assign new_n12646_ = ~new_n12644_ & ~new_n12645_;
  assign new_n12647_ = new_n10738_ & ~new_n12646_;
  assign new_n12648_ = ng2574 & new_n12647_;
  assign new_n12649_ = new_n10736_ & new_n12648_;
  assign new_n12650_ = ~new_n12641_ & ~new_n12649_;
  assign new_n12651_ = ~new_n10734_ & new_n12650_;
  assign new_n12652_ = ~new_n10738_ & new_n10767_;
  assign new_n12653_ = new_n10734_ & new_n12652_;
  assign n6082 = new_n12651_ | new_n12653_;
  assign new_n12655_ = ng3013 & new_n10784_;
  assign new_n12656_ = ng3010 & new_n12655_;
  assign new_n12657_ = ~ng3024 & new_n12656_;
  assign new_n12658_ = ng3024 & ~new_n12656_;
  assign new_n12659_ = ~new_n12657_ & ~new_n12658_;
  assign n6087 = new_n10780_ & ~new_n12659_;
  assign new_n12661_ = ~ng45 & ~ng48;
  assign new_n12662_ = ~ng48 & ~new_n12661_;
  assign new_n12663_ = ~ng45 & ~new_n12661_;
  assign new_n12664_ = ~new_n12662_ & ~new_n12663_;
  assign new_n12665_ = ~ng42 & ~ng39;
  assign new_n12666_ = ~ng42 & ~new_n12665_;
  assign new_n12667_ = ~ng39 & ~new_n12665_;
  assign new_n12668_ = ~new_n12666_ & ~new_n12667_;
  assign new_n12669_ = ~new_n12664_ & ~new_n12668_;
  assign new_n12670_ = ~new_n12664_ & ~new_n12669_;
  assign new_n12671_ = ~new_n12668_ & ~new_n12669_;
  assign new_n12672_ = ~new_n12670_ & ~new_n12671_;
  assign new_n12673_ = ~ng27 & ~ng30;
  assign new_n12674_ = ~ng27 & ~new_n12673_;
  assign new_n12675_ = ~ng30 & ~new_n12673_;
  assign new_n12676_ = ~new_n12674_ & ~new_n12675_;
  assign new_n12677_ = ~ng36 & ~ng33;
  assign new_n12678_ = ~ng33 & ~new_n12677_;
  assign new_n12679_ = ~ng36 & ~new_n12677_;
  assign new_n12680_ = ~new_n12678_ & ~new_n12679_;
  assign new_n12681_ = ~new_n12676_ & ~new_n12680_;
  assign new_n12682_ = ~new_n12676_ & ~new_n12681_;
  assign new_n12683_ = ~new_n12680_ & ~new_n12681_;
  assign new_n12684_ = ~new_n12682_ & ~new_n12683_;
  assign new_n12685_ = ~new_n12672_ & ~new_n12684_;
  assign new_n12686_ = ~new_n12672_ & ~new_n12685_;
  assign new_n12687_ = ~new_n12684_ & ~new_n12685_;
  assign new_n12688_ = ~new_n12686_ & ~new_n12687_;
  assign new_n12689_ = ~ng3083 & ~new_n12688_;
  assign new_n12690_ = ~new_n12688_ & ~new_n12689_;
  assign new_n12691_ = ~ng3083 & ~new_n12689_;
  assign n6097 = ~new_n12690_ & ~new_n12691_;
  assign new_n12693_ = ~ng3077 & ng2987;
  assign new_n12694_ = ~ng2987 & ~ng3059;
  assign n6102 = ~new_n12693_ & ~new_n12694_;
  assign new_n12696_ = ng2950 & ~ng2883;
  assign new_n12697_ = ~ng2950 & ng2883;
  assign new_n12698_ = ~new_n12696_ & ~new_n12697_;
  assign n6107 = ~new_n9234_ | ~new_n12698_;
  assign new_n12700_ = ~ng143 & ~new_n4777_1_;
  assign new_n12701_ = ng105 & new_n4777_1_;
  assign n6122 = ~new_n12700_ & ~new_n12701_;
  assign new_n12703_ = ~ng152 & ~new_n4777_1_;
  assign new_n12704_ = ng117 & new_n4777_1_;
  assign n6127 = ~new_n12703_ & ~new_n12704_;
  assign new_n12706_ = ~ng161 & ~new_n4777_1_;
  assign new_n12707_ = new_n4777_1_ & ~new_n4932_1_;
  assign n6132 = ~new_n12706_ & ~new_n12707_;
  assign new_n12709_ = ~ng173 & ~new_n6278_;
  assign new_n12710_ = ng101 & new_n6278_;
  assign n6137 = ~new_n12709_ & ~new_n12710_;
  assign new_n12712_ = ng823 & ~new_n10304_;
  assign new_n12713_ = ~ng823 & ~ng189;
  assign n6142 = ~new_n12712_ & ~new_n12713_;
  assign new_n12715_ = ng823 & ~new_n11737_;
  assign new_n12716_ = ~ng823 & ~ng243;
  assign n6147 = ~new_n12715_ & ~new_n12716_;
  assign new_n12718_ = ng61 & ~new_n9292_;
  assign new_n12719_ = ~ng61 & new_n9292_;
  assign new_n12720_ = ~new_n12718_ & ~new_n12719_;
  assign n6152 = ~new_n5127_1_ & ~new_n12720_;
  assign new_n12722_ = ~ng384 & ~new_n5138_;
  assign new_n12723_ = new_n5138_ & ~new_n9901_;
  assign n6157 = ~new_n12722_ & ~new_n12723_;
  assign new_n12725_ = ng826 & new_n12144_;
  assign new_n12726_ = ~ng826 & ~ng417;
  assign n6162 = ~new_n12725_ & ~new_n12726_;
  assign new_n12728_ = ng826 & new_n5239_;
  assign new_n12729_ = ~ng826 & ~ng438;
  assign n6167 = ~new_n12728_ & ~new_n12729_;
  assign new_n12731_ = ng826 & ~new_n7705_;
  assign new_n12732_ = ~ng826 & ~ng315;
  assign n6172 = ~new_n12731_ & ~new_n12732_;
  assign new_n12734_ = ~ng403 & ~new_n6003_;
  assign new_n12735_ = new_n6003_ & new_n11767_;
  assign n6177 = ~new_n12734_ & ~new_n12735_;
  assign new_n12737_ = ng826 & ~new_n5068_;
  assign new_n12738_ = ~ng826 & ~ng477;
  assign n6206 = ~new_n12737_ & ~new_n12738_;
  assign new_n12740_ = ~ng581 & ~new_n5307_;
  assign new_n12741_ = new_n5307_ & ~new_n10854_;
  assign n6219 = ~new_n12740_ & ~new_n12741_;
  assign new_n12743_ = ng1315 & ~new_n10337_;
  assign new_n12744_ = ~ng1315 & ~ng602;
  assign n6224 = ~new_n12743_ & ~new_n12744_;
  assign new_n12746_ = ng1315 & ~new_n5376_;
  assign new_n12747_ = ~ng1315 & ~ng496;
  assign n6229 = ~new_n12746_ & ~new_n12747_;
  assign new_n12749_ = ~ng699 & ~new_n5395_;
  assign new_n12750_ = ng640 & new_n5395_;
  assign n6239 = ~new_n12749_ & ~new_n12750_;
  assign new_n12752_ = ~ng708 & ~new_n5395_;
  assign new_n12753_ = ng646 & new_n5395_;
  assign n6244 = ~new_n12752_ & ~new_n12753_;
  assign new_n12755_ = ~ng717 & ~new_n5395_;
  assign new_n12756_ = ng666 & new_n5395_;
  assign n6249 = ~new_n12755_ & ~new_n12756_;
  assign new_n12758_ = ~ng726 & ~new_n5395_;
  assign new_n12759_ = ng692 & new_n5395_;
  assign n6254 = ~new_n12758_ & ~new_n12759_;
  assign new_n12761_ = ~ng735 & ~new_n5395_;
  assign new_n12762_ = new_n5395_ & ~new_n5514_;
  assign n6259 = ~new_n12761_ & ~new_n12762_;
  assign new_n12764_ = ~ng818 & ~new_n5517_1_;
  assign new_n12765_ = ng785 & new_n5517_1_;
  assign n6264 = ~new_n12764_ & ~new_n12765_;
  assign new_n12767_ = ~ng833 & ~new_n5517_1_;
  assign new_n12768_ = ng797 & new_n5517_1_;
  assign n6269 = ~new_n12767_ & ~new_n12768_;
  assign new_n12770_ = ~ng842 & ~new_n5517_1_;
  assign new_n12771_ = ng809 & new_n5517_1_;
  assign n6274 = ~new_n12770_ & ~new_n12771_;
  assign new_n12773_ = ~ng851 & ~new_n5517_1_;
  assign new_n12774_ = new_n5517_1_ & ~new_n5652_;
  assign n6279 = ~new_n12773_ & ~new_n12774_;
  assign new_n12776_ = ng826 & ~new_n10359_;
  assign new_n12777_ = ~ng826 & ~ng891;
  assign n6284 = ~new_n12776_ & ~new_n12777_;
  assign new_n12779_ = ng826 & ~new_n10882_;
  assign new_n12780_ = ~ng826 & ~ng945;
  assign n6289 = ~new_n12779_ & ~new_n12780_;
  assign new_n12782_ = ~ng780 & new_n5128_;
  assign new_n12783_ = ng780 & ~new_n5128_;
  assign new_n12784_ = ~new_n12782_ & ~new_n12783_;
  assign n6294 = ~new_n5127_1_ & ~new_n12784_;
  assign new_n12786_ = ng744 & new_n5918_1_;
  assign new_n12787_ = ng740 & ~new_n12786_;
  assign new_n12788_ = ~ng740 & new_n12786_;
  assign new_n12789_ = ~new_n12787_ & ~new_n12788_;
  assign n6299 = ~new_n5127_1_ & ~new_n12789_;
  assign new_n12791_ = ~ng1063 & ~new_n8502_;
  assign new_n12792_ = new_n8502_ & ~new_n12214_;
  assign n6304 = ~new_n12791_ & ~new_n12792_;
  assign new_n12794_ = ng853 & new_n11877_;
  assign new_n12795_ = ~ng853 & ~ng1110;
  assign n6309 = ~new_n12794_ & ~new_n12795_;
  assign new_n12797_ = ng853 & new_n9393_;
  assign new_n12798_ = ~ng853 & ~ng1131;
  assign n6314 = ~new_n12797_ & ~new_n12798_;
  assign new_n12800_ = ng853 & ~new_n9946_;
  assign new_n12801_ = ~ng853 & ~ng1004;
  assign n6319 = ~new_n12800_ & ~new_n12801_;
  assign new_n12803_ = ng853 & ~new_n5824_;
  assign new_n12804_ = ~ng853 & ~ng1166;
  assign n6344 = ~new_n12803_ & ~new_n12804_;
  assign new_n12806_ = ng1326 & ~new_n6242_;
  assign new_n12807_ = ~ng1326 & new_n6242_;
  assign new_n12808_ = ~new_n12806_ & ~new_n12807_;
  assign n6358 = ~new_n6241_ & ~new_n12808_;
  assign new_n12810_ = ng1372 & new_n12485_;
  assign new_n12811_ = ~ng1378 & new_n12810_;
  assign new_n12812_ = ng1378 & ~new_n12810_;
  assign new_n12813_ = ~new_n12811_ & ~new_n12812_;
  assign n6363 = ~new_n6241_ & ~new_n12813_;
  assign new_n12815_ = ~ng1390 & ~new_n6263_;
  assign new_n12816_ = ng1339 & new_n6263_;
  assign n6368 = ~new_n12815_ & ~new_n12816_;
  assign new_n12818_ = ~ng1399 & ~new_n6263_;
  assign new_n12819_ = ng1358 & new_n6263_;
  assign n6373 = ~new_n12818_ & ~new_n12819_;
  assign new_n12821_ = ~ng1408 & ~new_n6263_;
  assign new_n12822_ = ng1372 & new_n6263_;
  assign n6378 = ~new_n12821_ & ~new_n12822_;
  assign new_n12824_ = ~ng1556 & ~new_n8121_;
  assign new_n12825_ = ng1471 & new_n8121_;
  assign n6383 = ~new_n12824_ & ~new_n12825_;
  assign new_n12827_ = ng853 & ~new_n11944_;
  assign new_n12828_ = ~ng853 & ~ng1618;
  assign n6388 = ~new_n12827_ & ~new_n12828_;
  assign new_n12830_ = ng853 & ~new_n8063_;
  assign new_n12831_ = ~ng853 & ~ng1591;
  assign n6393 = ~new_n12830_ & ~new_n12831_;
  assign new_n12833_ = ng853 & ~new_n6622_;
  assign new_n12834_ = ~ng853 & ~ng1645;
  assign n6398 = ~new_n12833_ & ~new_n12834_;
  assign new_n12836_ = ~ng1457 & new_n6627_;
  assign new_n12837_ = ng1457 & ~new_n6627_;
  assign new_n12838_ = ~new_n12836_ & ~new_n12837_;
  assign n6403 = ~new_n5127_1_ & ~new_n12838_;
  assign new_n12840_ = ng853 & new_n7476_;
  assign new_n12841_ = ~ng853 & ~ng2498;
  assign n6425 = ~new_n12840_ & ~new_n12841_;
  assign new_n12843_ = ng853 & new_n12274_;
  assign new_n12844_ = ~ng853 & ~ng2519;
  assign n6430 = ~new_n12843_ & ~new_n12844_;
  assign new_n12846_ = ng853 & ~new_n12001_;
  assign new_n12847_ = ~ng853 & ~ng2392;
  assign n6435 = ~new_n12846_ & ~new_n12847_;
  assign new_n12849_ = ng826 & ~new_n7308_;
  assign new_n12850_ = ~ng826 & ~ng2552;
  assign n6452 = ~new_n12849_ & ~new_n12850_;
  assign new_n12852_ = ng1309 & ~new_n9626_;
  assign new_n12853_ = ~ng1309 & ~ng2565;
  assign n6465 = ~new_n12852_ & ~new_n12853_;
  assign new_n12855_ = ~ng1315 & ~ng2733;
  assign n6475 = ~new_n9359_ & ~new_n12855_;
  assign new_n12857_ = ng2760 & ~new_n10594_;
  assign new_n12858_ = ~ng2760 & new_n10594_;
  assign new_n12859_ = ~new_n12857_ & ~new_n12858_;
  assign n6480 = ~new_n8213_ & ~new_n12859_;
  assign new_n12861_ = ~ng2780 & ~new_n7588_;
  assign new_n12862_ = ng2727 & new_n7588_;
  assign n6485 = ~new_n12861_ & ~new_n12862_;
  assign new_n12864_ = ~ng2789 & ~new_n7588_;
  assign new_n12865_ = ng2746 & new_n7588_;
  assign n6490 = ~new_n12864_ & ~new_n12865_;
  assign new_n12867_ = ~ng2798 & ~new_n7588_;
  assign new_n12868_ = ng2760 & new_n7588_;
  assign n6495 = ~new_n12867_ & ~new_n12868_;
  assign new_n12870_ = ~ng2807 & ~new_n8213_;
  assign new_n12871_ = ~new_n7529_ & new_n8213_;
  assign n6500 = ~new_n12870_ & ~new_n12871_;
  assign n6505 = ~pg3234 & ng3054;
  assign new_n12874_ = ~ng1220 & new_n11015_;
  assign new_n12875_ = ~new_n11139_ & new_n12874_;
  assign new_n12876_ = new_n11104_ & new_n11139_;
  assign new_n12877_ = ~new_n12875_ & ~new_n12876_;
  assign new_n12878_ = ~new_n11141_ & new_n12877_;
  assign n6510 = new_n12616_ | new_n12878_;
  assign new_n12880_ = ~ng1914 & new_n10635_;
  assign new_n12881_ = ~new_n10633_ & new_n12880_;
  assign new_n12882_ = ~new_n10686_ & ~new_n10708_;
  assign new_n12883_ = ~new_n6796_ & ~new_n12882_;
  assign new_n12884_ = ~new_n12882_ & ~new_n12883_;
  assign new_n12885_ = ~new_n6796_ & ~new_n12883_;
  assign new_n12886_ = ~new_n12884_ & ~new_n12885_;
  assign new_n12887_ = new_n10635_ & ~new_n12886_;
  assign new_n12888_ = ng1880 & new_n12887_;
  assign new_n12889_ = new_n10633_ & new_n12888_;
  assign new_n12890_ = ~new_n12881_ & ~new_n12889_;
  assign new_n12891_ = ~new_n10631_ & new_n12890_;
  assign n6515 = new_n12056_ | new_n12891_;
  assign new_n12893_ = ~ng2608 & new_n10738_;
  assign new_n12894_ = ~new_n10736_ & new_n12893_;
  assign new_n12895_ = ~new_n8255_ & ~new_n10756_;
  assign new_n12896_ = ~new_n7540_ & ~new_n12895_;
  assign new_n12897_ = ~new_n12895_ & ~new_n12896_;
  assign new_n12898_ = ~new_n7540_ & ~new_n12896_;
  assign new_n12899_ = ~new_n12897_ & ~new_n12898_;
  assign new_n12900_ = new_n10738_ & ~new_n12899_;
  assign new_n12901_ = ng2574 & new_n12900_;
  assign new_n12902_ = new_n10736_ & new_n12901_;
  assign new_n12903_ = ~new_n12894_ & ~new_n12902_;
  assign new_n12904_ = ~new_n10734_ & new_n12903_;
  assign n6520 = new_n12653_ | new_n12904_;
  assign new_n12906_ = ng3010 & ~new_n12655_;
  assign new_n12907_ = ~ng3010 & new_n12655_;
  assign new_n12908_ = ~new_n12906_ & ~new_n12907_;
  assign n6525 = new_n10780_ & ~new_n12908_;
  assign new_n12910_ = ~ng3062 & ng2987;
  assign new_n12911_ = ~ng3043 & ~ng2987;
  assign n6530 = ~new_n12910_ & ~new_n12911_;
  assign new_n12913_ = new_n11432_ & ~new_n12688_;
  assign new_n12914_ = new_n11432_ & ~new_n12913_;
  assign new_n12915_ = ~new_n12688_ & ~new_n12913_;
  assign n6535 = new_n12914_ | new_n12915_;
  assign new_n12917_ = ~ng3078 & ng2987;
  assign new_n12918_ = ~ng2987 & ~ng3060;
  assign n6540 = ~new_n12917_ & ~new_n12918_;
  assign new_n12920_ = ~ng2963 & ~ng2879;
  assign new_n12921_ = ~ng2827 & ng2879;
  assign n6550 = ~new_n12920_ & ~new_n12921_;
  assign new_n12923_ = ~ng2874 & ng2879;
  assign new_n12924_ = ~ng2200 & ~ng2879;
  assign n6560 = ~new_n12923_ & ~new_n12924_;
  assign new_n12926_ = ng1315 & ~ng559;
  assign new_n12927_ = ~ng1315 & ~ng3084;
  assign n6565 = ~new_n12926_ & ~new_n12927_;
  assign new_n12929_ = ~ng1222 & new_n11015_;
  assign new_n12930_ = ~new_n11139_ & new_n12929_;
  assign new_n12931_ = new_n11115_ & new_n11139_;
  assign new_n12932_ = ~new_n12930_ & ~new_n12931_;
  assign new_n12933_ = ~new_n11141_ & new_n12932_;
  assign new_n12934_ = ~new_n11038_ & new_n11381_;
  assign new_n12935_ = new_n11141_ & new_n12934_;
  assign n6570 = new_n12933_ | new_n12935_;
  assign new_n12937_ = ~new_n10664_ & ~new_n10708_;
  assign new_n12938_ = ~new_n6796_ & ~new_n12937_;
  assign new_n12939_ = ~new_n12937_ & ~new_n12938_;
  assign new_n12940_ = ~new_n6796_ & ~new_n12938_;
  assign new_n12941_ = ~new_n12939_ & ~new_n12940_;
  assign new_n12942_ = new_n10635_ & ~new_n12941_;
  assign new_n12943_ = ng1880 & new_n12942_;
  assign new_n12944_ = new_n12636_ & new_n12943_;
  assign new_n12945_ = new_n12636_ & ~new_n12944_;
  assign new_n12946_ = new_n12943_ & ~new_n12944_;
  assign new_n12947_ = ~new_n12945_ & ~new_n12946_;
  assign new_n12948_ = ng1937 & ~new_n12947_;
  assign new_n12949_ = new_n10715_ & new_n11677_;
  assign new_n12950_ = new_n10715_ & ~new_n12949_;
  assign new_n12951_ = new_n11677_ & ~new_n12949_;
  assign new_n12952_ = ~new_n12950_ & ~new_n12951_;
  assign new_n12953_ = new_n11401_ & new_n12327_;
  assign new_n12954_ = new_n11401_ & ~new_n12953_;
  assign new_n12955_ = new_n12327_ & ~new_n12953_;
  assign new_n12956_ = ~new_n12954_ & ~new_n12955_;
  assign new_n12957_ = ~new_n12952_ & ~new_n12956_;
  assign new_n12958_ = ~new_n12952_ & ~new_n12957_;
  assign new_n12959_ = ~new_n12956_ & ~new_n12957_;
  assign new_n12960_ = ~new_n12958_ & ~new_n12959_;
  assign new_n12961_ = new_n12051_ & new_n12888_;
  assign new_n12962_ = new_n12051_ & ~new_n12961_;
  assign new_n12963_ = new_n12888_ & ~new_n12961_;
  assign new_n12964_ = ~new_n12962_ & ~new_n12963_;
  assign new_n12965_ = ~new_n10691_ & ~new_n10708_;
  assign new_n12966_ = ~new_n6796_ & ~new_n12965_;
  assign new_n12967_ = ~new_n12965_ & ~new_n12966_;
  assign new_n12968_ = ~new_n6796_ & ~new_n12966_;
  assign new_n12969_ = ~new_n12967_ & ~new_n12968_;
  assign new_n12970_ = new_n10635_ & ~new_n12969_;
  assign new_n12971_ = ng1880 & new_n12970_;
  assign new_n12972_ = new_n12626_ & new_n12971_;
  assign new_n12973_ = new_n12626_ & ~new_n12972_;
  assign new_n12974_ = new_n12971_ & ~new_n12972_;
  assign new_n12975_ = ~new_n12973_ & ~new_n12974_;
  assign new_n12976_ = ~new_n12964_ & ~new_n12975_;
  assign new_n12977_ = ~new_n12964_ & ~new_n12976_;
  assign new_n12978_ = ~new_n12975_ & ~new_n12976_;
  assign new_n12979_ = ~new_n12977_ & ~new_n12978_;
  assign new_n12980_ = ~new_n12960_ & ~new_n12979_;
  assign new_n12981_ = ~new_n12960_ & ~new_n12980_;
  assign new_n12982_ = ~new_n12979_ & ~new_n12980_;
  assign new_n12983_ = ~new_n12981_ & ~new_n12982_;
  assign new_n12984_ = ng1890 & ~new_n12983_;
  assign new_n12985_ = ~pg3229 & ~ng1921;
  assign new_n12986_ = pg3229 & ~ng1918;
  assign new_n12987_ = ~new_n12985_ & ~new_n12986_;
  assign new_n12988_ = new_n10635_ & new_n12987_;
  assign new_n12989_ = ~new_n10631_ & ~new_n10633_;
  assign new_n12990_ = new_n12988_ & new_n12989_;
  assign new_n12991_ = new_n10629_ & new_n12990_;
  assign new_n12992_ = ~new_n12948_ & ~new_n12984_;
  assign n6575 = new_n12991_ | ~new_n12992_;
  assign new_n12994_ = ~ng2978 & ~ng2879;
  assign new_n12995_ = ~ng2867 & ng2879;
  assign n6580 = ~new_n12994_ & ~new_n12995_;
  assign new_n12997_ = ~ng2944 & ~ng2879;
  assign new_n12998_ = ~ng2845 & ng2879;
  assign n6590 = ~new_n12997_ & ~new_n12998_;
  assign new_n13000_ = ~ng1245 & ng1309;
  assign new_n13001_ = ~ng1309 & ~ng3085;
  assign n6600 = ~new_n13000_ & ~new_n13001_;
  assign new_n13003_ = ~ng1223 & new_n11015_;
  assign new_n13004_ = ~new_n11139_ & new_n13003_;
  assign new_n13005_ = new_n11122_ & new_n11139_;
  assign new_n13006_ = ~new_n13004_ & ~new_n13005_;
  assign new_n13007_ = ~new_n11141_ & new_n13006_;
  assign new_n13008_ = ~new_n11045_ & new_n11381_;
  assign new_n13009_ = new_n11141_ & new_n13008_;
  assign n6605 = new_n13007_ | new_n13009_;
  assign new_n13011_ = ~ng1917 & new_n10635_;
  assign new_n13012_ = ~new_n10633_ & new_n13011_;
  assign new_n13013_ = new_n10633_ & new_n12971_;
  assign new_n13014_ = ~new_n13012_ & ~new_n13013_;
  assign new_n13015_ = ~new_n10631_ & new_n13014_;
  assign new_n13016_ = new_n10719_ & ~new_n12943_;
  assign new_n13017_ = new_n10631_ & new_n13016_;
  assign n6610 = new_n13015_ | new_n13017_;
  assign new_n13019_ = ~pg3231 & ng3139;
  assign new_n13020_ = ng2981 & ng2874;
  assign new_n13021_ = ng2874 & ~new_n13020_;
  assign new_n13022_ = ng2981 & ~new_n13020_;
  assign new_n13023_ = ~new_n13021_ & ~new_n13022_;
  assign new_n13024_ = ng2975 & ng2978;
  assign new_n13025_ = ng2978 & ~new_n13024_;
  assign new_n13026_ = ng2975 & ~new_n13024_;
  assign new_n13027_ = ~new_n13025_ & ~new_n13026_;
  assign new_n13028_ = ~new_n13023_ & ~new_n13027_;
  assign new_n13029_ = ~new_n13023_ & ~new_n13028_;
  assign new_n13030_ = ~new_n13027_ & ~new_n13028_;
  assign new_n13031_ = ~new_n13029_ & ~new_n13030_;
  assign new_n13032_ = ng2969 & ng2972;
  assign new_n13033_ = ng2972 & ~new_n13032_;
  assign new_n13034_ = ng2969 & ~new_n13032_;
  assign new_n13035_ = ~new_n13033_ & ~new_n13034_;
  assign new_n13036_ = ng2963 & ng2966;
  assign new_n13037_ = ng2966 & ~new_n13036_;
  assign new_n13038_ = ng2963 & ~new_n13036_;
  assign new_n13039_ = ~new_n13037_ & ~new_n13038_;
  assign new_n13040_ = ~new_n13035_ & ~new_n13039_;
  assign new_n13041_ = ~new_n13035_ & ~new_n13040_;
  assign new_n13042_ = ~new_n13039_ & ~new_n13040_;
  assign new_n13043_ = ~new_n13041_ & ~new_n13042_;
  assign new_n13044_ = ~new_n13031_ & ~new_n13043_;
  assign new_n13045_ = ~new_n13031_ & ~new_n13044_;
  assign new_n13046_ = ~new_n13043_ & ~new_n13044_;
  assign new_n13047_ = ~new_n13045_ & ~new_n13046_;
  assign new_n13048_ = new_n13019_ & ~new_n13047_;
  assign new_n13049_ = new_n13019_ & ~new_n13048_;
  assign new_n13050_ = ~new_n13047_ & ~new_n13048_;
  assign new_n13051_ = ~new_n13049_ & ~new_n13050_;
  assign new_n13052_ = ~ng2879 & ~new_n13051_;
  assign new_n13053_ = ~ng2830 & ng2879;
  assign n6619 = ~new_n13052_ & ~new_n13053_;
  assign new_n13055_ = ng2956 & ng2959;
  assign new_n13056_ = ng2959 & ~new_n13055_;
  assign new_n13057_ = ng2956 & ~new_n13055_;
  assign new_n13058_ = ~new_n13056_ & ~new_n13057_;
  assign new_n13059_ = ng2947 & ng2953;
  assign new_n13060_ = ng2953 & ~new_n13059_;
  assign new_n13061_ = ng2947 & ~new_n13059_;
  assign new_n13062_ = ~new_n13060_ & ~new_n13061_;
  assign new_n13063_ = ~new_n13058_ & ~new_n13062_;
  assign new_n13064_ = ~new_n13058_ & ~new_n13063_;
  assign new_n13065_ = ~new_n13062_ & ~new_n13063_;
  assign new_n13066_ = ~new_n13064_ & ~new_n13065_;
  assign new_n13067_ = ng2941 & ng2944;
  assign new_n13068_ = ng2944 & ~new_n13067_;
  assign new_n13069_ = ng2941 & ~new_n13067_;
  assign new_n13070_ = ~new_n13068_ & ~new_n13069_;
  assign new_n13071_ = ng2935 & ng2938;
  assign new_n13072_ = ng2938 & ~new_n13071_;
  assign new_n13073_ = ng2935 & ~new_n13071_;
  assign new_n13074_ = ~new_n13072_ & ~new_n13073_;
  assign new_n13075_ = ~new_n13070_ & ~new_n13074_;
  assign new_n13076_ = ~new_n13070_ & ~new_n13075_;
  assign new_n13077_ = ~new_n13074_ & ~new_n13075_;
  assign new_n13078_ = ~new_n13076_ & ~new_n13077_;
  assign new_n13079_ = ~new_n13066_ & ~new_n13078_;
  assign new_n13080_ = ~new_n13066_ & ~new_n13079_;
  assign new_n13081_ = ~new_n13078_ & ~new_n13079_;
  assign new_n13082_ = ~new_n13080_ & ~new_n13081_;
  assign new_n13083_ = new_n13019_ & ~new_n13082_;
  assign new_n13084_ = new_n13019_ & ~new_n13083_;
  assign new_n13085_ = ~new_n13082_ & ~new_n13083_;
  assign new_n13086_ = ~new_n13084_ & ~new_n13085_;
  assign new_n13087_ = ~ng2879 & ~new_n13086_;
  assign new_n13088_ = ~ng2858 & ng2879;
  assign n6629 = ~new_n13087_ & ~new_n13088_;
  assign new_n13090_ = ng1312 & ~ng1245;
  assign new_n13091_ = ~ng1312 & ~ng3086;
  assign n6633 = ~new_n13090_ & ~new_n13091_;
  assign new_n13093_ = new_n12076_ & new_n12350_;
  assign new_n13094_ = new_n12076_ & ~new_n13093_;
  assign new_n13095_ = new_n12350_ & ~new_n13093_;
  assign new_n13096_ = ~new_n13094_ & ~new_n13095_;
  assign new_n13097_ = ng2631 & ~new_n13096_;
  assign new_n13098_ = new_n11417_ & new_n11690_;
  assign new_n13099_ = new_n11417_ & ~new_n13098_;
  assign new_n13100_ = new_n11690_ & ~new_n13098_;
  assign new_n13101_ = ~new_n13099_ & ~new_n13100_;
  assign new_n13102_ = new_n10763_ & new_n11159_;
  assign new_n13103_ = new_n10763_ & ~new_n13102_;
  assign new_n13104_ = new_n11159_ & ~new_n13102_;
  assign new_n13105_ = ~new_n13103_ & ~new_n13104_;
  assign new_n13106_ = ~new_n13101_ & ~new_n13105_;
  assign new_n13107_ = ~new_n13101_ & ~new_n13106_;
  assign new_n13108_ = ~new_n13105_ & ~new_n13106_;
  assign new_n13109_ = ~new_n13107_ & ~new_n13108_;
  assign new_n13110_ = new_n12648_ & new_n12901_;
  assign new_n13111_ = new_n12648_ & ~new_n13110_;
  assign new_n13112_ = new_n12901_ & ~new_n13110_;
  assign new_n13113_ = ~new_n13111_ & ~new_n13112_;
  assign new_n13114_ = new_n12066_ & new_n12340_;
  assign new_n13115_ = new_n12066_ & ~new_n13114_;
  assign new_n13116_ = new_n12340_ & ~new_n13114_;
  assign new_n13117_ = ~new_n13115_ & ~new_n13116_;
  assign new_n13118_ = ~new_n13113_ & ~new_n13117_;
  assign new_n13119_ = ~new_n13113_ & ~new_n13118_;
  assign new_n13120_ = ~new_n13117_ & ~new_n13118_;
  assign new_n13121_ = ~new_n13119_ & ~new_n13120_;
  assign new_n13122_ = ~new_n13109_ & ~new_n13121_;
  assign new_n13123_ = ~new_n13109_ & ~new_n13122_;
  assign new_n13124_ = ~new_n13121_ & ~new_n13122_;
  assign new_n13125_ = ~new_n13123_ & ~new_n13124_;
  assign new_n13126_ = ng2584 & ~new_n13125_;
  assign new_n13127_ = ~pg3229 & ~ng2615;
  assign new_n13128_ = pg3229 & ~ng2612;
  assign new_n13129_ = ~new_n13127_ & ~new_n13128_;
  assign new_n13130_ = new_n10738_ & new_n13129_;
  assign new_n13131_ = ~new_n10734_ & ~new_n10736_;
  assign new_n13132_ = new_n13130_ & new_n13131_;
  assign new_n13133_ = new_n10732_ & new_n13132_;
  assign new_n13134_ = ~new_n13097_ & ~new_n13126_;
  assign n6638 = new_n13133_ | ~new_n13134_;
  assign new_n13136_ = ng3028 & new_n12085_;
  assign new_n13137_ = ng3036 & new_n13136_;
  assign new_n13138_ = ng3032 & ~new_n13137_;
  assign new_n13139_ = ~ng3032 & new_n13137_;
  assign new_n13140_ = ~new_n13138_ & ~new_n13139_;
  assign n6643 = new_n12084_ & ~new_n13140_;
  assign new_n13142_ = ~ng2975 & ~ng2879;
  assign new_n13143_ = ~ng2870 & ng2879;
  assign n6653 = ~new_n13142_ & ~new_n13143_;
  assign new_n13145_ = ~ng2947 & ~ng2879;
  assign new_n13146_ = ~ng2842 & ng2879;
  assign n6662 = ~new_n13145_ & ~new_n13146_;
  assign new_n13148_ = ng1315 & ~ng1245;
  assign new_n13149_ = ~ng1315 & ~ng3087;
  assign n6671 = ~new_n13148_ & ~new_n13149_;
  assign new_n13151_ = ng3080 & ~ng2993;
  assign new_n13152_ = ~ng3080 & ng2993;
  assign new_n13153_ = ~new_n13151_ & ~new_n13152_;
  assign new_n13154_ = new_n10780_ & new_n13153_;
  assign new_n13155_ = pg3234 & ~new_n10780_;
  assign n6676 = ~new_n13154_ & ~new_n13155_;
  assign new_n13157_ = ~ng3036 & new_n13136_;
  assign new_n13158_ = ng3036 & ~new_n13136_;
  assign new_n13159_ = ~new_n13157_ & ~new_n13158_;
  assign n6681 = new_n12084_ & ~new_n13159_;
  assign new_n13161_ = ng2900 & new_n9239_;
  assign new_n13162_ = ~ng2908 & new_n13161_;
  assign new_n13163_ = ng2908 & ~new_n13161_;
  assign new_n13164_ = ~new_n13162_ & ~new_n13163_;
  assign n6686 = new_n9234_ & ~new_n13164_;
  assign new_n13166_ = ~ng2941 & ng2879;
  assign new_n13167_ = ~ng1481 & ~ng2879;
  assign n6701 = ~new_n13166_ & ~new_n13167_;
  assign new_n13169_ = ~ng1939 & ng1309;
  assign new_n13170_ = ~ng1309 & ~ng3091;
  assign n6706 = ~new_n13169_ & ~new_n13170_;
  assign new_n13172_ = ng823 & ~new_n8712_;
  assign new_n13173_ = ~ng823 & ~ng1570;
  assign n6711 = ~new_n13172_ & ~new_n13173_;
  assign new_n13175_ = ~ng2210 & ~new_n4777_1_;
  assign new_n13176_ = ng2170 & new_n4777_1_;
  assign n6725 = ~new_n13175_ & ~new_n13176_;
  assign new_n13178_ = ~ng2227 & ~new_n5517_1_;
  assign new_n13179_ = ng2190 & new_n5517_1_;
  assign n6730 = ~new_n13178_ & ~new_n13179_;
  assign new_n13181_ = ng2987 & ~ng3067;
  assign new_n13182_ = ~ng3048 & ~ng2987;
  assign n6735 = ~new_n13181_ & ~new_n13182_;
  assign new_n13184_ = ng2987 & ~ng3076;
  assign new_n13185_ = ~ng2987 & ~ng3058;
  assign n6740 = ~new_n13184_ & ~new_n13185_;
  assign new_n13187_ = ng2912 & ~ng2917;
  assign new_n13188_ = new_n9233_ & new_n13187_;
  assign new_n13189_ = ng2920 & new_n13188_;
  assign new_n13190_ = ~ng2924 & new_n13189_;
  assign new_n13191_ = ~ng2814 & ~new_n13190_;
  assign new_n13192_ = ~ng2912 & new_n9233_;
  assign new_n13193_ = ng2912 & ~new_n9233_;
  assign new_n13194_ = ~new_n13192_ & ~new_n13193_;
  assign n6745 = ~new_n13191_ | ~new_n13194_;
  assign new_n13196_ = ~ng2944 & ng2879;
  assign new_n13197_ = ~ng1486 & ~ng2879;
  assign n6760 = ~new_n13196_ & ~new_n13197_;
  assign new_n13199_ = ng1312 & ~ng1939;
  assign new_n13200_ = ~ng1312 & ~ng3092;
  assign n6765 = ~new_n13199_ & ~new_n13200_;
  assign new_n13202_ = ng853 & ~new_n11284_;
  assign new_n13203_ = ~ng853 & ~ng1627;
  assign n6770 = ~new_n13202_ & ~new_n13203_;
  assign new_n13205_ = ~ng2208 & ~new_n4773_;
  assign new_n13206_ = ng2170 & new_n4773_;
  assign n6783 = ~new_n13205_ & ~new_n13206_;
  assign new_n13208_ = ~ng2223 & ~new_n4773_;
  assign new_n13209_ = ng2185 & new_n4773_;
  assign n6788 = ~new_n13208_ & ~new_n13209_;
  assign new_n13211_ = ~ng3068 & ng2987;
  assign new_n13212_ = ~ng3049 & ~ng2987;
  assign n6793 = ~new_n13211_ & ~new_n13212_;
  assign new_n13214_ = ~ng3075 & ng2987;
  assign new_n13215_ = ~ng3057 & ~ng2987;
  assign n6798 = ~new_n13214_ & ~new_n13215_;
  assign new_n13217_ = ng2912 & new_n9233_;
  assign new_n13218_ = ng2917 & ~new_n13217_;
  assign new_n13219_ = ~ng2917 & new_n13217_;
  assign new_n13220_ = ~new_n13218_ & ~new_n13219_;
  assign n6803 = new_n13191_ & ~new_n13220_;
  assign new_n13222_ = ~ng2947 & ng2879;
  assign new_n13223_ = ~ng1491 & ~ng2879;
  assign n6818 = ~new_n13222_ & ~new_n13223_;
  assign new_n13225_ = ng826 & ~new_n6622_;
  assign new_n13226_ = ~ng826 & ~ng1639;
  assign n6823 = ~new_n13225_ & ~new_n13226_;
  assign new_n13228_ = ng1315 & ng1934;
  assign new_n13229_ = ~ng1315 & ~ng1937;
  assign n6833 = ~new_n13228_ & ~new_n13229_;
  assign new_n13231_ = ~ng2218 & ~new_n5517_1_;
  assign new_n13232_ = ng2175 & new_n5517_1_;
  assign n6838 = ~new_n13231_ & ~new_n13232_;
  assign new_n13234_ = ~ng2226 & ~new_n4773_;
  assign new_n13235_ = ng2190 & new_n4773_;
  assign n6843 = ~new_n13234_ & ~new_n13235_;
  assign new_n13237_ = ng823 & ~new_n7514_;
  assign new_n13238_ = ~ng2524 & ~new_n13237_;
  assign new_n13239_ = new_n7507_ & new_n13237_;
  assign n6848 = ~new_n13238_ & ~new_n13239_;
  assign new_n13241_ = ng2917 & new_n13217_;
  assign new_n13242_ = ~ng2924 & new_n13241_;
  assign new_n13243_ = ng2924 & ~new_n13241_;
  assign new_n13244_ = ~new_n13242_ & ~new_n13243_;
  assign n6853 = new_n13191_ & ~new_n13244_;
  assign new_n13246_ = ~ng2953 & ng2879;
  assign new_n13247_ = ~ng1496 & ~ng2879;
  assign n6868 = ~new_n13246_ & ~new_n13247_;
  assign new_n13249_ = ng1462 & ~new_n6626_;
  assign new_n13250_ = ~ng1462 & new_n6626_;
  assign new_n13251_ = ~new_n13249_ & ~new_n13250_;
  assign n6873 = ~new_n5127_1_ & ~new_n13251_;
  assign new_n13253_ = ~ng1315 & ~ng1934;
  assign n6882 = ~new_n7709_ & ~new_n13253_;
  assign new_n13255_ = ~ng2219 & ~new_n4777_1_;
  assign new_n13256_ = ng2175 & new_n4777_1_;
  assign n6887 = ~new_n13255_ & ~new_n13256_;
  assign new_n13258_ = ~ng2228 & ~new_n4777_1_;
  assign new_n13259_ = ng2190 & new_n4777_1_;
  assign n6892 = ~new_n13258_ & ~new_n13259_;
  assign new_n13261_ = ng826 & ~new_n10425_;
  assign new_n13262_ = ~ng2502 & ~new_n13261_;
  assign new_n13263_ = new_n10422_ & new_n13261_;
  assign n6897 = ~new_n13262_ & ~new_n13263_;
  assign new_n13265_ = ng2924 & new_n13241_;
  assign new_n13266_ = ng2920 & ~new_n13265_;
  assign new_n13267_ = ~ng2920 & new_n13265_;
  assign new_n13268_ = ~new_n13266_ & ~new_n13267_;
  assign n6902 = new_n13191_ & ~new_n13268_;
  assign new_n13270_ = ~ng2874 & ~ng2879;
  assign new_n13271_ = ~ng2861 & ng2879;
  assign n6917 = ~new_n13270_ & ~new_n13271_;
  assign new_n13273_ = ~ng2953 & ~ng2879;
  assign new_n13274_ = ~ng2839 & ng2879;
  assign n6927 = ~new_n13273_ & ~new_n13274_;
  assign new_n13276_ = ~ng1724 & ~new_n6636_;
  assign new_n13277_ = new_n6636_ & ~new_n10168_;
  assign n6931 = ~new_n13276_ & ~new_n13277_;
  assign new_n13279_ = ng826 & ~new_n6634_;
  assign new_n13280_ = ~ng826 & ~ng1836;
  assign n6941 = ~new_n13279_ & ~new_n13280_;
  assign new_n13282_ = ~ng2085 & ~new_n7003_;
  assign new_n13283_ = ng2033 & new_n7003_;
  assign n6946 = ~new_n13282_ & ~new_n13283_;
  assign new_n13285_ = ~ng2093 & ~new_n7007_;
  assign new_n13286_ = ng2052 & new_n7007_;
  assign n6951 = ~new_n13285_ & ~new_n13286_;
  assign new_n13288_ = ~ng2107 & ~new_n7011_;
  assign new_n13289_ = ng2072 & new_n7011_;
  assign n6956 = ~new_n13288_ & ~new_n13289_;
  assign new_n13291_ = ng1309 & ~new_n10033_;
  assign new_n13292_ = ~ng2118 & ~new_n13291_;
  assign new_n13293_ = ng2010 & new_n13291_;
  assign n6961 = ~new_n13292_ & ~new_n13293_;
  assign new_n13295_ = ~ng2451 & ~new_n7410_;
  assign new_n13296_ = new_n7410_ & ~new_n8164_;
  assign n6966 = ~new_n13295_ & ~new_n13296_;
  assign new_n13298_ = ng2934 & ~new_n13082_;
  assign new_n13299_ = ~new_n13082_ & ~new_n13298_;
  assign new_n13300_ = ng2934 & ~new_n13298_;
  assign n6971 = new_n13299_ | new_n13300_;
  assign new_n13302_ = ng2879 & ~new_n13086_;
  assign new_n13303_ = ~ng2877 & ~ng2879;
  assign n6986 = ~new_n13302_ & ~new_n13303_;
  assign new_n13305_ = ~ng2966 & ~ng2879;
  assign new_n13306_ = ~ng2824 & ng2879;
  assign n6991 = ~new_n13305_ & ~new_n13306_;
  assign new_n13308_ = ~ng1772 & ~new_n9087_;
  assign new_n13309_ = new_n9087_ & ~new_n9991_;
  assign n7000 = ~new_n13308_ & ~new_n13309_;
  assign new_n13311_ = ng853 & new_n6710_;
  assign new_n13312_ = ~ng853 & ~ng1869;
  assign n7009 = ~new_n13311_ & ~new_n13312_;
  assign new_n13314_ = ~ng2086 & ~new_n7011_;
  assign new_n13315_ = ng2033 & new_n7011_;
  assign n7014 = ~new_n13314_ & ~new_n13315_;
  assign new_n13317_ = ~ng2095 & ~new_n7011_;
  assign new_n13318_ = ng2052 & new_n7011_;
  assign n7019 = ~new_n13317_ & ~new_n13318_;
  assign new_n13320_ = ~ng2105 & ~new_n7007_;
  assign new_n13321_ = ng2072 & new_n7007_;
  assign n7024 = ~new_n13320_ & ~new_n13321_;
  assign new_n13323_ = ~ng2114 & ~new_n7007_;
  assign new_n13324_ = ng1312 & ~ng2110;
  assign new_n13325_ = ng1315 & ~ng2108;
  assign new_n13326_ = ~ng2109 & ng1309;
  assign new_n13327_ = ~new_n13324_ & ~new_n13325_;
  assign new_n13328_ = ~new_n13326_ & new_n13327_;
  assign new_n13329_ = ~ng2040 & ~new_n10676_;
  assign new_n13330_ = ~new_n10676_ & ~new_n13329_;
  assign new_n13331_ = ~ng2040 & ~new_n13329_;
  assign new_n13332_ = ~new_n13330_ & ~new_n13331_;
  assign new_n13333_ = ~ng2013 & ~new_n10681_;
  assign new_n13334_ = ~new_n10681_ & ~new_n13333_;
  assign new_n13335_ = ~ng2013 & ~new_n13333_;
  assign new_n13336_ = ~new_n13334_ & ~new_n13335_;
  assign new_n13337_ = ~ng2033 & ~new_n10686_;
  assign new_n13338_ = ~new_n10686_ & ~new_n13337_;
  assign new_n13339_ = ~ng2033 & ~new_n13337_;
  assign new_n13340_ = ~new_n13338_ & ~new_n13339_;
  assign new_n13341_ = ~ng2020 & ~new_n10691_;
  assign new_n13342_ = ~new_n10691_ & ~new_n13341_;
  assign new_n13343_ = ~ng2020 & ~new_n13341_;
  assign new_n13344_ = ~new_n13342_ & ~new_n13343_;
  assign new_n13345_ = ~new_n13336_ & ~new_n13340_;
  assign new_n13346_ = ~new_n13344_ & new_n13345_;
  assign new_n13347_ = ~ng2026 & ~new_n10698_;
  assign new_n13348_ = ~new_n10698_ & ~new_n13347_;
  assign new_n13349_ = ~ng2026 & ~new_n13347_;
  assign new_n13350_ = ~new_n13348_ & ~new_n13349_;
  assign new_n13351_ = ~new_n13332_ & new_n13346_;
  assign new_n13352_ = ~new_n13350_ & new_n13351_;
  assign new_n13353_ = ~ng2072 & ~new_n10647_;
  assign new_n13354_ = ~new_n10647_ & ~new_n13353_;
  assign new_n13355_ = ~ng2072 & ~new_n13353_;
  assign new_n13356_ = ~new_n13354_ & ~new_n13355_;
  assign new_n13357_ = ~ng2046 & ~new_n10652_;
  assign new_n13358_ = ~new_n10652_ & ~new_n13357_;
  assign new_n13359_ = ~ng2046 & ~new_n13357_;
  assign new_n13360_ = ~new_n13358_ & ~new_n13359_;
  assign new_n13361_ = ~ng2059 & ~new_n10642_;
  assign new_n13362_ = ~new_n10642_ & ~new_n13361_;
  assign new_n13363_ = ~ng2059 & ~new_n13361_;
  assign new_n13364_ = ~new_n13362_ & ~new_n13363_;
  assign new_n13365_ = ~ng2052 & ~new_n10657_;
  assign new_n13366_ = ~new_n10657_ & ~new_n13365_;
  assign new_n13367_ = ~ng2052 & ~new_n13365_;
  assign new_n13368_ = ~new_n13366_ & ~new_n13367_;
  assign new_n13369_ = ~new_n13360_ & ~new_n13364_;
  assign new_n13370_ = ~new_n13368_ & new_n13369_;
  assign new_n13371_ = ~ng2066 & ~new_n10664_;
  assign new_n13372_ = ~new_n10664_ & ~new_n13371_;
  assign new_n13373_ = ~ng2066 & ~new_n13371_;
  assign new_n13374_ = ~new_n13372_ & ~new_n13373_;
  assign new_n13375_ = ~new_n13356_ & new_n13370_;
  assign new_n13376_ = ~new_n13374_ & new_n13375_;
  assign new_n13377_ = new_n13352_ & new_n13376_;
  assign new_n13378_ = new_n13328_ & ~new_n13377_;
  assign new_n13379_ = new_n10705_ & new_n13378_;
  assign new_n13380_ = new_n7007_ & ~new_n13379_;
  assign n7029 = ~new_n13323_ & ~new_n13380_;
  assign new_n13382_ = ng2962 & ~new_n13047_;
  assign new_n13383_ = ~new_n13047_ & ~new_n13382_;
  assign new_n13384_ = ng2962 & ~new_n13382_;
  assign n7038 = new_n13383_ | new_n13384_;
  assign new_n13386_ = ~ng2935 & ng2879;
  assign new_n13387_ = ~ng1471 & ~ng2879;
  assign n7053 = ~new_n13386_ & ~new_n13387_;
  assign new_n13389_ = ~ng2966 & ng2879;
  assign new_n13390_ = ~ng2170 & ~ng2879;
  assign n7063 = ~new_n13389_ & ~new_n13390_;
  assign new_n13392_ = ng826 & ~new_n9102_;
  assign new_n13393_ = ~ng826 & ~ng1810;
  assign n7068 = ~new_n13392_ & ~new_n13393_;
  assign new_n13395_ = ng826 & ~new_n6303_;
  assign new_n13396_ = ~ng826 & ~ng1846;
  assign n7073 = ~new_n13395_ & ~new_n13396_;
  assign new_n13398_ = ng1315 & ~ng1868;
  assign new_n13399_ = ng1309 & ~ng1869;
  assign new_n13400_ = ng1312 & ~ng1867;
  assign new_n13401_ = ~new_n13398_ & ~new_n13399_;
  assign n7078 = ~new_n13400_ & new_n13401_;
  assign new_n13403_ = ~ng2084 & ~new_n7007_;
  assign new_n13404_ = ng2033 & new_n7007_;
  assign n7082 = ~new_n13403_ & ~new_n13404_;
  assign new_n13406_ = ~ng2098 & ~new_n7011_;
  assign new_n13407_ = ng2046 & new_n7011_;
  assign n7087 = ~new_n13406_ & ~new_n13407_;
  assign new_n13409_ = ~ng2102 & ~new_n7007_;
  assign new_n13410_ = ng2066 & new_n7007_;
  assign n7092 = ~new_n13409_ & ~new_n13410_;
  assign new_n13412_ = ~ng2116 & ~new_n7011_;
  assign new_n13413_ = new_n7011_ & ~new_n13379_;
  assign n7097 = ~new_n13412_ & ~new_n13413_;
  assign new_n13415_ = ~ng2151 & new_n7396_1_;
  assign new_n13416_ = ng2151 & ~new_n7396_1_;
  assign new_n13417_ = ~new_n13415_ & ~new_n13416_;
  assign n7102 = ~new_n5127_1_ & ~new_n13417_;
  assign new_n13419_ = ~ng2938 & ng2879;
  assign new_n13420_ = ~ng1476 & ~ng2879;
  assign n7122 = ~new_n13419_ & ~new_n13420_;
  assign new_n13422_ = ~ng2935 & ~ng2879;
  assign new_n13423_ = ~ng2854 & ng2879;
  assign n7127 = ~new_n13422_ & ~new_n13423_;
  assign new_n13425_ = ~ng2969 & ng2879;
  assign new_n13426_ = ~ng2175 & ~ng2879;
  assign n7131 = ~new_n13425_ & ~new_n13426_;
  assign new_n13428_ = ng823 & ~new_n9474_;
  assign new_n13429_ = ~ng823 & ~ng1694;
  assign n7136 = ~new_n13428_ & ~new_n13429_;
  assign new_n13431_ = ng823 & ~new_n6303_;
  assign new_n13432_ = ~ng823 & ~ng1849;
  assign n7141 = ~new_n13431_ & ~new_n13432_;
  assign new_n13434_ = ~ng2088 & ~new_n7003_;
  assign new_n13435_ = ng2026 & new_n7003_;
  assign n7150 = ~new_n13434_ & ~new_n13435_;
  assign new_n13437_ = ~ng2097 & ~new_n7003_;
  assign new_n13438_ = ng2046 & new_n7003_;
  assign n7155 = ~new_n13437_ & ~new_n13438_;
  assign new_n13440_ = ~ng2106 & ~new_n7003_;
  assign new_n13441_ = ng2072 & new_n7003_;
  assign n7160 = ~new_n13440_ & ~new_n13441_;
  assign new_n13443_ = ~ng2115 & ~new_n7003_;
  assign new_n13444_ = new_n7003_ & ~new_n13379_;
  assign n7165 = ~new_n13443_ & ~new_n13444_;
  assign new_n13446_ = ng823 & ~new_n9574_;
  assign new_n13447_ = ~ng823 & ~ng2336;
  assign n7170 = ~new_n13446_ & ~new_n13447_;
  assign new_n13449_ = ~ng2879 & ~ng2959;
  assign new_n13450_ = ~ng2833 & ng2879;
  assign n7188 = ~new_n13449_ & ~new_n13450_;
  assign new_n13452_ = ~ng2972 & ng2879;
  assign new_n13453_ = ~ng2180 & ~ng2879;
  assign n7198 = ~new_n13452_ & ~new_n13453_;
  assign new_n13455_ = ~ng2963 & ng2879;
  assign new_n13456_ = ~ng2165 & ~ng2879;
  assign n7203 = ~new_n13455_ & ~new_n13456_;
  assign new_n13458_ = ng853 & new_n8766_;
  assign new_n13459_ = ~ng1702 & ~new_n13458_;
  assign new_n13460_ = new_n8773_ & new_n13458_;
  assign n7208 = ~new_n13459_ & ~new_n13460_;
  assign new_n13462_ = ~ng1963 & ~new_n8088_;
  assign new_n13463_ = new_n8088_ & ~new_n9127_;
  assign n7213 = ~new_n13462_ & ~new_n13463_;
  assign new_n13465_ = new_n6912_1_ & ~new_n6983_;
  assign new_n13466_ = new_n6839_ & new_n13465_;
  assign new_n13467_ = ~new_n6968_ & new_n6983_;
  assign new_n13468_ = new_n6912_1_ & new_n13467_;
  assign new_n13469_ = ~new_n13466_ & ~new_n13468_;
  assign new_n13470_ = new_n5366_ & new_n13469_;
  assign new_n13471_ = ~new_n5366_ & new_n6796_;
  assign new_n13472_ = ~new_n13470_ & ~new_n13471_;
  assign new_n13473_ = ng1309 & ~new_n13472_;
  assign new_n13474_ = ~ng1309 & ~ng1994;
  assign n7218 = ~new_n13473_ & ~new_n13474_;
  assign new_n13476_ = ng1312 & ~new_n13472_;
  assign new_n13477_ = ~ng1312 & ~ng1997;
  assign n7223 = ~new_n13476_ & ~new_n13477_;
  assign new_n13479_ = ~ng1890 & ng1315;
  assign new_n13480_ = ~ng1315 & ~ng2010;
  assign n7233 = ~new_n13479_ & ~new_n13480_;
  assign new_n13482_ = ng2052 & new_n10202_;
  assign new_n13483_ = ng2046 & new_n13482_;
  assign new_n13484_ = ng2059 & new_n13483_;
  assign new_n13485_ = ng2066 & new_n13484_;
  assign new_n13486_ = ~ng2072 & new_n13485_;
  assign new_n13487_ = ng2072 & ~new_n13485_;
  assign new_n13488_ = ~new_n13486_ & ~new_n13487_;
  assign n7238 = ~new_n6993_ & ~new_n13488_;
  assign new_n13490_ = ng826 & ~new_n8818_;
  assign new_n13491_ = ~ng826 & ~ng2279;
  assign n7243 = ~new_n13490_ & ~new_n13491_;
  assign new_n13493_ = ng2930 & ~ng2929;
  assign n7248 = ~ng2879 | new_n13493_;
  assign new_n13495_ = ~ng2972 & ~ng2879;
  assign new_n13496_ = ng2879 & ~ng2818;
  assign n7258 = ~new_n13495_ & ~new_n13496_;
  assign new_n13498_ = ~ng2938 & ~ng2879;
  assign new_n13499_ = ng2879 & ~ng2851;
  assign n7267 = ~new_n13498_ & ~new_n13499_;
  assign new_n13501_ = ~ng2975 & ng2879;
  assign new_n13502_ = ~ng2879 & ~ng2185;
  assign n7271 = ~new_n13501_ & ~new_n13502_;
  assign new_n13504_ = ng2879 & ~new_n13051_;
  assign new_n13505_ = ~ng2879 & ~ng2878;
  assign n7276 = ~new_n13504_ & ~new_n13505_;
  assign new_n13507_ = ~ng1961 & ~new_n8779_;
  assign new_n13508_ = new_n8779_ & ~new_n9127_;
  assign n7285 = ~new_n13507_ & ~new_n13508_;
  assign new_n13510_ = ng1315 & ~new_n8783_;
  assign new_n13511_ = ~ng1315 & ~ng1982;
  assign n7290 = ~new_n13510_ & ~new_n13511_;
  assign new_n13513_ = ng1315 & ~new_n13472_;
  assign new_n13514_ = ~ng1315 & ~ng2000;
  assign n7295 = ~new_n13513_ & ~new_n13514_;
  assign new_n13516_ = ~ng1315 & ~ng2039;
  assign n7304 = ~new_n9359_ & ~new_n13516_;
  assign new_n13518_ = ng2066 & ~new_n13484_;
  assign new_n13519_ = ~ng2066 & new_n13484_;
  assign new_n13520_ = ~new_n13518_ & ~new_n13519_;
  assign n7309 = ~new_n6993_ & ~new_n13520_;
  assign new_n13522_ = ng853 & ~new_n10047_;
  assign new_n13523_ = ~ng853 & ~ng2267;
  assign n7314 = ~new_n13522_ & ~new_n13523_;
  assign new_n13525_ = ng2879 & ~ng2959;
  assign new_n13526_ = ~ng2879 & ~ng1506;
  assign n7319 = ~new_n13525_ & ~new_n13526_;
  assign new_n13528_ = ~ng2981 & ~ng2879;
  assign new_n13529_ = ng2879 & ~ng2864;
  assign n7324 = ~new_n13528_ & ~new_n13529_;
  assign new_n13531_ = ~ng2956 & ~ng2879;
  assign new_n13532_ = ng2879 & ~ng2836;
  assign n7332 = ~new_n13531_ & ~new_n13532_;
  assign new_n13534_ = ~ng2978 & ng2879;
  assign new_n13535_ = ~ng2879 & ~ng2190;
  assign n7340 = ~new_n13534_ & ~new_n13535_;
  assign new_n13537_ = ng1309 & ~ng559;
  assign new_n13538_ = ~ng1309 & ~ng3210;
  assign n7345 = ~new_n13537_ & ~new_n13538_;
  assign new_n13540_ = ng1309 & ~new_n6989_;
  assign new_n13541_ = ~ng1309 & ~ng1985;
  assign n7350 = ~new_n13540_ & ~new_n13541_;
  assign new_n13543_ = ~pg3229 & ~ng1686;
  assign new_n13544_ = pg3229 & ng1672;
  assign n7360 = ~new_n13543_ & ~new_n13544_;
  assign new_n13546_ = ~ng2059 & new_n13483_;
  assign new_n13547_ = ng2059 & ~new_n13483_;
  assign new_n13548_ = ~new_n13546_ & ~new_n13547_;
  assign n7365 = ~new_n6993_ & ~new_n13548_;
  assign new_n13550_ = ~ng2249 & ~new_n6278_;
  assign new_n13551_ = ng2170 & new_n6278_;
  assign n7370 = ~new_n13550_ & ~new_n13551_;
  assign new_n13553_ = ~ng2956 & ng2879;
  assign new_n13554_ = ~ng2879 & ~ng1501;
  assign n7375 = ~new_n13553_ & ~new_n13554_;
  assign new_n13556_ = ~ng2969 & ~ng2879;
  assign new_n13557_ = ng2879 & ~ng2821;
  assign n7384 = ~new_n13556_ & ~new_n13557_;
  assign new_n13559_ = ~ng2941 & ~ng2879;
  assign new_n13560_ = ng2879 & ~ng2848;
  assign n7392 = ~new_n13559_ & ~new_n13560_;
  assign new_n13562_ = ~ng2981 & ng2879;
  assign new_n13563_ = ~ng2879 & ~ng2195;
  assign n7396 = ~new_n13562_ & ~new_n13563_;
  assign new_n13565_ = ng1312 & ~ng559;
  assign new_n13566_ = ~ng1312 & ~ng3211;
  assign n7401 = ~new_n13565_ & ~new_n13566_;
  assign new_n13568_ = ng1312 & ~new_n6989_;
  assign new_n13569_ = ~ng1312 & ~ng1988;
  assign n7406 = ~new_n13568_ & ~new_n13569_;
  assign new_n13571_ = ng2046 & ~new_n13482_;
  assign new_n13572_ = ~ng2046 & new_n13482_;
  assign new_n13573_ = ~new_n13571_ & ~new_n13572_;
  assign n7421 = ~new_n6993_ & ~new_n13573_;
  assign new_n13575_ = ~ng2236 & ~new_n5517_1_;
  assign new_n13576_ = new_n5517_1_ & ~new_n7020_;
  assign n7426 = ~new_n13575_ & ~new_n13576_;
  assign pg24734 = ~n2171;
  assign pg26135 = ~n6112;
  assign pg25435 = ~n2873;
  assign pg27380 = ~n5659;
  assign n332 = ~ng121;
  assign n462 = ~ng797;
  assign n627 = ~ng1662;
  assign n822 = ~ng101;
  assign n1070 = ~ng1501;
  assign n1107 = ~ng1660;
  assign n1177 = ~ng2165;
  assign n1293 = ~ng125;
  assign n1463 = ~ng1140;
  assign n1571 = ~ng1666;
  assign n1641 = ~ng2190;
  assign n1760 = ~ng105;
  assign n1913 = ~ng1138;
  assign n1918 = ~ng966;
  assign n1987 = ~ng1496;
  assign n2024 = ~ng1664;
  assign n2221 = ~ng451;
  assign n2261 = ~ng805;
  assign n2391 = ~ng1670;
  assign n2461 = ~ng2185;
  assign n2496 = ~ng2362;
  assign n2575 = ~ng453;
  assign n2619 = ~ng785;
  assign n2741 = ~ng1668;
  assign n2843 = ~ng2360;
  assign n2907 = ~ng279;
  assign n2947 = ~ng801;
  assign n3146 = ~ng2180;
  assign n3180 = ~ng2358;
  assign n3237 = ~ng281;
  assign n3364 = ~ng1506;
  assign n3586 = ~ng289;
  assign n3621 = ~ng813;
  assign n3650 = ~ng976;
  assign n3740 = ~ng2175;
  assign n3865 = ~ng117;
  assign n3893 = ~ng287;
  assign n3932 = ~ng793;
  assign n3994 = ~ng1476;
  assign n4036 = ~ng2200;
  assign n4063 = ~ng2526;
  assign n4068 = ~ng2366;
  assign n4191 = ~ng291;
  assign n4226 = ~ng809;
  assign n4260 = ~ng978;
  assign n4363 = ~ng2170;
  assign n4569 = ~ng789;
  assign n4649 = ~ng1471;
  assign n4691 = ~ng2195;
  assign n4732 = ~ng2364;
  assign n5022 = ~ng968;
  assign n5162 = ~ng2356;
  assign n5302 = ~ng109;
  assign n5453 = ~ng970;
  assign n5508 = ~ng1486;
  assign n5729 = ~ng97;
  assign n5783 = ~ng285;
  assign n5908 = ~ng972;
  assign n6032 = ~ng2528;
  assign n6182 = ~ng113;
  assign n6234 = ~ng283;
  assign n6353 = ~ng974;
  assign n6408 = ~ng1481;
  assign n6470 = ~ng2354;
  assign n7281 = ~ng1491;
  assign n7355 = ~ng1834;
  assign n7411 = ~ng1832;
  assign n7416 = ~ng1672;
  assign pg8012 = ng826;
  assign pg8023 = ng2842;
  assign pg8265 = ng20;
  assign pg16297 = ng520;
  assign pg8167 = ng823;
  assign pg8266 = ng23;
  assign pg8275 = ng48;
  assign pg4090 = ng2864;
  assign pg7161 = ng1312;
  assign pg7194 = ng1312;
  assign pg8021 = ng2930;
  assign pg8175 = ng2845;
  assign pg8263 = ng14;
  assign pg8274 = ng45;
  assign pg7052 = ng1309;
  assign pg8264 = ng17;
  assign pg8273 = ng42;
  assign pg7390 = ng1312;
  assign pg8261 = ng8;
  assign pg8272 = ng39;
  assign pg8262 = ng11;
  assign pg8271 = ng36;
  assign pg16355 = ng1206;
  assign pg6573 = ng826;
  assign pg7084 = ng823;
  assign pg7264 = ng823;
  assign pg7334 = ng2827;
  assign pg8007 = ng823;
  assign pg8106 = ng1309;
  assign pg8270 = ng33;
  assign pg8251 = ng2861;
  assign pg8260 = ng5;
  assign pg4590 = ng2870;
  assign pg6642 = ng1312;
  assign pg6750 = ng1309;
  assign pg7302 = ng1309;
  assign pg4450 = ng2854;
  assign pg6225 = ng2818;
  assign pg4088 = ng2836;
  assign pg5472 = ng826;
  assign pg6442 = ng2821;
  assign pg8030 = ng1312;
  assign pg16437 = ng2594;
  assign pg5511 = ng826;
  assign pg7014 = ng823;
  assign pg16399 = ng1900;
  assign pg6313 = ng823;
  assign pg5612 = ng2258;
  assign pg6231 = ng826;
  assign pg5437 = ng826;
  assign pg5657 = ng1309;
  assign pg6979 = ng1309;
  assign pg3993 = ng2848;
  assign pg6911 = ng1312;
  assign pg6944 = ng1312;
  assign pg4323 = ng2867;
  assign pg6712 = ng823;
  assign pg6837 = ng826;
  assign pg7519 = ng2830;
  assign pg5686 = ng1312;
  assign pg5738 = ng1312;
  assign pg6447 = ng823;
  assign pg4200 = ng2851;
  assign pg4321 = ng2839;
  assign pg5388 = ng3040;
  assign pg5555 = ng826;
  assign pg7229 = ng1309;
  assign pg5549 = ng2258;
  assign pg5637 = ng2258;
  assign pg5648 = ng1312;
  assign pg5747 = ng1309;
  assign pg5629 = ng1309;
  assign pg6518 = ng823;
  assign pg7425 = ng1309;
  assign pg5595 = ng2258;
  assign pg8082 = ng823;
  assign pg5695 = ng1309;
  assign pg6368 = ng826;
  assign pg6485 = ng1309;
  assign pg6782 = ng823;
  assign pg7961 = ng826;
  assign pg7357 = ng1312;
  assign pg5796 = ng1312;
  assign pg7909 = ng826;
  assign pg7956 = ng823;
  assign pg8096 = ng2858;
  assign pg8258 = ng1;
  assign pg8269 = ng30;
  assign pg6677 = ng1309;
  assign pg8087 = ng826;
  assign pg8249 = ng2833;
  assign pg8267 = ng26;
  assign pg6895 = ng2824;
  assign pg7487 = ng1312;
  assign pg8259 = ng2;
  assign pg8268 = ng27;
  assign n287 = pg26149;
  assign n337 = ng373;
  assign n347 = ng465;
  assign n357 = ng528;
  assign n472 = ng1052;
  assign n477 = ng1075;
  assign n482 = ng1250;
  assign n497 = ng1235;
  assign n512 = ng1206;
  assign n587 = ng1833;
  assign n597 = ng1954;
  assign n607 = ng1915;
  assign n697 = ng2361;
  assign n702 = ng2425;
  assign n707 = ng2448;
  assign n717 = ng2540;
  assign n727 = ng2602;
  assign n777 = pg27380;
  assign n826 = ng380;
  assign n835 = ng574;
  assign n844 = ng535;
  assign n948 = ng969;
  assign n962 = ng1082;
  assign n967 = ng1142;
  assign n1079 = ng1846;
  assign n1088 = ng1908;
  assign n1182 = ng2418;
  assign n1185 = ng2455;
  assign n1194 = ng2648;
  assign n1203 = ng2609;
  assign n1253 = pg25435;
  assign n1298 = ng284;
  assign n1303 = ng376;
  assign n1313 = ng461;
  assign n1423 = ng1041;
  assign n1428 = ng1054;
  assign n1433 = ng1209;
  assign n1468 = ng1312;
  assign n1533 = ng1835;
  assign n1537 = ng1893;
  assign n1542 = ng1946;
  assign n1646 = ng2451;
  assign n1656 = ng2536;
  assign n1716 = pg26104;
  assign n1755 = ng450;
  assign n1763 = ng382;
  assign n1772 = ng572;
  assign n1781 = ng543;
  assign n1880 = ng1029;
  assign n1885 = ng1048;
  assign n1889 = ng1074;
  assign n1923 = ng1309;
  assign n1990 = ng1903;
  assign n1995 = ng1849;
  assign n2094 = ng2527;
  assign n2098 = ng2457;
  assign n2107 = ng2646;
  assign n2116 = ng2617;
  assign n2206 = ng361;
  assign n2211 = ng458;
  assign n2266 = ng975;
  assign n2356 = ng1836;
  assign n2361 = ng1948;
  assign n2376 = ng1938;
  assign n2386 = ng1880;
  assign n2466 = ng2365;
  assign n2471 = ng2432;
  assign n2476 = ng2533;
  assign n2526 = pg25442;
  assign n2556 = ng354;
  assign n2561 = ng365;
  assign n2565 = ng570;
  assign n2614 = ng1141;
  assign n2707 = ng1944;
  assign n2712 = ng1852;
  assign n2810 = ng2529;
  assign n2820 = ng2444;
  assign n2823 = ng2644;
  assign n2838 = ng2574;
  assign n2892 = ng342;
  assign n2897 = ng384;
  assign n2902 = ng397;
  assign n2952 = ng977;
  assign n2961 = ng1244;
  assign n3036 = ng1831;
  assign n3041 = ng1839;
  assign n3056 = ng1923;
  assign n3131 = ng2258;
  assign n3150 = ng2363;
  assign n3155 = ng2427;
  assign n3160 = ng2459;
  assign n3165 = ng2472;
  assign n3205 = pg25420;
  assign n3224 = ng367;
  assign n3228 = ng372;
  assign n3233 = ng391;
  assign n3276 = ng967;
  assign n3281 = ng2873;
  assign n3284 = ng1214;
  assign n3304 = ng1186;
  assign n3367 = ng1950;
  assign n3470 = ng2355;
  assign n3475 = ng2878;
  assign n3479 = ng2421;
  assign n3482 = ng2447;
  assign n3487 = ng2466;
  assign n3556 = ng454;
  assign n3561 = ng2857;
  assign n3566 = ng369;
  assign n3581 = ng499;
  assign n3626 = ng971;
  assign n3631 = ng1056;
  assign n3636 = ng1069;
  assign n3641 = ng1199;
  assign n3690 = ng1665;
  assign n3695 = ng1723;
  assign n3700 = ng1765;
  assign n3705 = ng1778;
  assign n3745 = ng2429;
  assign n3750 = ng2442;
  assign n3765 = ng2594;
  assign n3868 = ng290;
  assign n3873 = ng352;
  assign n3927 = ng1137;
  assign n3935 = ng1044;
  assign n3940 = ng1063;
  assign n3944 = ng1155;
  assign n3999 = ng1735;
  assign n4002 = ng1753;
  assign n4007 = ng1772;
  assign n4040 = ng2357;
  assign n4044 = ng2417;
  assign n4049 = ng2436;
  assign n4162 = ng452;
  assign n4172 = ng358;
  assign n4201 = ng2950;
  assign n4231 = ng973;
  assign n4236 = ng1045;
  assign n4245 = ng1260;
  assign n4314 = ng1667;
  assign n4319 = ng1731;
  assign n4324 = ng1742;
  assign n4329 = ng1776;
  assign n4358 = ng2525;
  assign n4372 = ng2440;
  assign n4511 = ng357;
  assign n4525 = ng520;
  assign n4564 = ng1139;
  assign n4573 = ng1085;
  assign n4581 = ng1152;
  assign n4595 = ng3080;
  assign n4654 = ng1724;
  assign n4657 = ng1748;
  assign n4662 = ng1769;
  assign n4694 = ng2359;
  assign n4704 = ng2433;
  assign n4857 = ng282;
  assign n4862 = ng343;
  assign n4867 = ng398;
  assign n4872 = ng523;
  assign n4877 = ng471;
  assign n4932 = ng823;
  assign n4987 = ng1030;
  assign n4992 = ng1059;
  assign n5002 = ng1258;
  assign n5077 = ng1661;
  assign n5087 = ng1739;
  assign n5092 = ng1768;
  assign n5122 = ng2473;
  assign n5127 = ng2597;
  assign n5132 = ng2546;
  assign n5212 = pg3234;
  assign n5305 = ng286;
  assign n5309 = ng387;
  assign n5313 = ng513;
  assign n5316 = ng568;
  assign n5330 = ng549;
  assign n5369 = ng826;
  assign n5422 = ng1037;
  assign n5427 = ng1071;
  assign n5436 = ng1148;
  assign n5439 = ng1252;
  assign n5443 = ng1229;
  assign n5513 = ng1671;
  assign n5517 = ng1746;
  assign n5522 = ng1779;
  assign n5535 = ng2256;
  assign n5549 = ng2462;
  assign n5553 = ng2587;
  assign n5556 = ng2642;
  assign n5570 = ng2623;
  assign n5634 = ng3040;
  assign n5654 = pg24734;
  assign n5724 = ng280;
  assign n5734 = ng346;
  assign n5738 = ng388;
  assign n5743 = ng564;
  assign n5748 = ng468;
  assign n5873 = ng1033;
  assign n5878 = ng1067;
  assign n5883 = ng1078;
  assign n5888 = ng1256;
  assign n5893 = ng1158;
  assign n5962 = ng1663;
  assign n5972 = ng1750;
  assign n5977 = ng1763;
  assign n5997 = ng2463;
  assign n6002 = ng2638;
  assign n6007 = ng2543;
  assign n6092 = pg16496;
  assign n6117 = pg26135;
  assign n6185 = ng288;
  assign n6189 = ng350;
  assign n6193 = ng395;
  assign n6198 = ng455;
  assign n6201 = ng566;
  assign n6214 = ng558;
  assign n6323 = ng1039;
  assign n6328 = ng1060;
  assign n6331 = ng1084;
  assign n6336 = ng1145;
  assign n6339 = ng1254;
  assign n6348 = ng1221;
  assign n6416 = ng1738;
  assign n6421 = ng1757;
  assign n6439 = ng2470;
  assign n6444 = ng2530;
  assign n6447 = ng2640;
  assign n6460 = ng2632;
  assign n6545 = ng2864;
  assign n6555 = ng2842;
  assign n6585 = ng2824;
  assign n6595 = ng2858;
  assign n6614 = ng2867;
  assign n6624 = ng2839;
  assign n6648 = pg51;
  assign n6657 = ng2827;
  assign n6666 = ng2854;
  assign n6691 = pg3228;
  assign n6696 = pg3218;
  assign n6715 = ng1669;
  assign n6720 = ng1733;
  assign n6750 = pg3212;
  assign n6755 = pg3217;
  assign n6775 = ng2877;
  assign n6779 = ng1727;
  assign n6808 = pg3226;
  assign n6813 = pg3220;
  assign n6828 = ng1754;
  assign n6858 = pg3227;
  assign n6863 = pg3219;
  assign n6877 = ng1761;
  assign n6907 = pg3224;
  assign n6912 = pg3214;
  assign n6922 = ng2821;
  assign n6936 = ng1842;
  assign n6976 = pg3225;
  assign n6981 = pg3213;
  assign n6995 = ng2836;
  assign n7004 = ng1952;
  assign n7033 = ng2258;
  assign n7043 = pg3222;
  assign n7048 = pg3216;
  assign n7058 = ng2851;
  assign n7107 = pg51;
  assign n7112 = pg3223;
  assign n7117 = pg3215;
  assign n7145 = ng1929;
  assign n7174 = ng2930;
  assign n7179 = pg3232;
  assign n7183 = ng2870;
  assign n7193 = ng2848;
  assign n7228 = ng1900;
  assign n7253 = pg3221;
  assign n7262 = ng2830;
  assign n7327 = ng2818;
  assign n7335 = ng2845;
  assign n7379 = ng2861;
  assign n7387 = ng2833;
  always @ (posedge clock) begin
    ng3097 <= n272;
    ng3108 <= n277;
    ng3185 <= n282;
    ng3135 <= n287;
    ng141 <= n292;
    ng155 <= n297;
    ng258 <= n302;
    ng83 <= n307;
    ng369 <= n312;
    ng414 <= n317;
    ng441 <= n322;
    ng318 <= n327;
    ng452 <= n332;
    ng380 <= n337;
    ng557 <= n342;
    ng574 <= n347;
    ng461 <= n352;
    ng535 <= n357;
    ng575 <= n362;
    ng590 <= n367;
    ng490 <= n372;
    ng646 <= n377;
    ng703 <= n382;
    ng714 <= n387;
    ng722 <= n392;
    ng736 <= n397;
    ng821 <= n402;
    ng835 <= n407;
    ng849 <= n412;
    ng863 <= n417;
    ng924 <= n422;
    ng939 <= n427;
    ng954 <= n432;
    ng744 <= n437;
    ng1085 <= n442;
    ng1113 <= n447;
    ng1000 <= n452;
    ng1090 <= n457;
    ng969 <= n462;
    ng992 <= n467;
    ng1053 <= n472;
    ng1082 <= n477;
    ng1255 <= n482;
    ng1173 <= n487;
    ng1151 <= n492;
    ng1186 <= n497;
    ng1267 <= n502;
    ng1303 <= n507;
    ng1211 <= n512;
    ng1352 <= n517;
    ng1392 <= n522;
    ng1403 <= n527;
    ng1411 <= n532;
    ng1425 <= n537;
    ng1527 <= n542;
    ng1535 <= n547;
    ng1552 <= n552;
    ng1642 <= n557;
    ng1453 <= n562;
    ng1739 <= n567;
    ng1798 <= n572;
    ng1825 <= n577;
    ng1700 <= n582;
    ng1834 <= n587;
    ng1890 <= n592;
    ng1945 <= n597;
    ng1858 <= n602;
    ng1922 <= n607;
    ng1959 <= n612;
    ng1973 <= n617;
    ng1991 <= n622;
    ng1912 <= n627;
    ng2033 <= n632;
    ng2082 <= n637;
    ng2090 <= n642;
    ng2104 <= n647;
    ng2237 <= n652;
    ng2251 <= n657;
    ng2312 <= n662;
    ng2327 <= n667;
    ng2342 <= n672;
    ng2124 <= n677;
    ng2436 <= n682;
    ng2495 <= n687;
    ng2523 <= n692;
    ng2362 <= n697;
    ng2426 <= n702;
    ng2455 <= n707;
    ng2631 <= n712;
    ng2648 <= n717;
    ng2536 <= n722;
    ng2609 <= n727;
    ng2649 <= n732;
    ng2772 <= n737;
    ng2786 <= n742;
    ng2797 <= n747;
    ng2805 <= n752;
    ng3044 <= n757;
    ng3098 <= n762;
    ng3107 <= n767;
    ng3088 <= n772;
    ng3139 <= n777;
    ng145 <= n782;
    ng154 <= n787;
    ng261 <= n792;
    ng88 <= n797;
    ng358 <= n802;
    ng411 <= n807;
    ng444 <= n812;
    ng317 <= n817;
    ng286 <= n822;
    ng381 <= n826;
    ng554 <= n831;
    ng565 <= n835;
    ng458 <= n840;
    ng542 <= n844;
    ng577 <= n849;
    ng593 <= n854;
    ng611 <= n859;
    ng660 <= n864;
    ng702 <= n869;
    ng715 <= n874;
    ng724 <= n879;
    ng734 <= n884;
    ng817 <= n889;
    ng839 <= n894;
    ng848 <= n899;
    ng921 <= n904;
    ng882 <= n909;
    ng936 <= n914;
    ng957 <= n919;
    ng749 <= n924;
    ng1075 <= n929;
    ng1115 <= n934;
    ng1001 <= n939;
    ng1008 <= n944;
    ng970 <= n948;
    ng986 <= n953;
    ng985 <= n958;
    ng1083 <= n962;
    ng1250 <= n967;
    ng1174 <= n971;
    ng1171 <= n976;
    ng1244 <= n981;
    ng1269 <= n986;
    ng1306 <= n991;
    ng1206 <= n996;
    ng1365 <= n1000;
    ng1391 <= n1005;
    ng1404 <= n1010;
    ng1413 <= n1015;
    ng1423 <= n1020;
    ng1523 <= n1025;
    ng1539 <= n1030;
    ng1551 <= n1035;
    ng1585 <= n1040;
    ng1448 <= n1045;
    ng1750 <= n1050;
    ng1801 <= n1055;
    ng1822 <= n1060;
    ng1701 <= n1065;
    ng1833 <= n1070;
    ng1893 <= n1074;
    ng1954 <= n1079;
    ng1859 <= n1083;
    ng1915 <= n1088;
    ng1960 <= n1092;
    ng1970 <= n1097;
    ng1871 <= n1102;
    ng1911 <= n1107;
    ng2026 <= n1112;
    ng2078 <= n1117;
    ng2094 <= n1122;
    ng2103 <= n1127;
    ng2235 <= n1132;
    ng2247 <= n1137;
    ng2270 <= n1142;
    ng2324 <= n1147;
    ng2345 <= n1152;
    ng2129 <= n1157;
    ng2459 <= n1162;
    ng2492 <= n1167;
    ng2394 <= n1172;
    ng2363 <= n1177;
    ng2425 <= n1182;
    ng2456 <= n1185;
    ng2628 <= n1190;
    ng2639 <= n1194;
    ng2533 <= n1199;
    ng2616 <= n1203;
    ng2651 <= n1208;
    ng2727 <= n1213;
    ng2784 <= n1218;
    ng2793 <= n1223;
    ng2809 <= n1228;
    ng3043 <= n1233;
    ng3099 <= n1238;
    ng3158 <= n1243;
    ng3179 <= n1248;
    ng3110 <= n1253;
    ng164 <= n1258;
    ng178 <= n1263;
    ng264 <= n1268;
    ng74 <= n1273;
    ng343 <= n1278;
    ng408 <= n1283;
    ng448 <= n1288;
    ng450 <= n1293;
    ng285 <= n1298;
    ng382 <= n1303;
    ng513 <= n1308;
    ng572 <= n1313;
    ng455 <= n1318;
    ng543 <= n1323;
    ng580 <= n1328;
    ng584 <= n1333;
    ng608 <= n1338;
    ng672 <= n1343;
    ng705 <= n1348;
    ng712 <= n1353;
    ng723 <= n1358;
    ng738 <= n1363;
    ng820 <= n1368;
    ng836 <= n1373;
    ng844 <= n1378;
    ng885 <= n1383;
    ng900 <= n1388;
    ng912 <= n1393;
    ng753 <= n1398;
    ng1078 <= n1403;
    ng1119 <= n1408;
    ng1134 <= n1413;
    ng1010 <= n1418;
    ng1029 <= n1423;
    ng1055 <= n1428;
    ng1210 <= n1433;
    ng1175 <= n1438;
    ng1155 <= n1443;
    ng1234 <= n1448;
    ng1268 <= n1453;
    ng1291 <= n1458;
    ng1216 <= n1463;
    ng1315 <= n1468;
    ng1402 <= n1473;
    ng1416 <= n1478;
    ng1420 <= n1483;
    ng1525 <= n1488;
    ng1540 <= n1493;
    ng1554 <= n1498;
    ng1573 <= n1503;
    ng1444 <= n1508;
    ng1765 <= n1513;
    ng1792 <= n1518;
    ng1819 <= n1523;
    ng1703 <= n1528;
    ng1660 <= n1533;
    ng1903 <= n1537;
    ng1947 <= n1542;
    ng1839 <= n1547;
    ng1908 <= n1552;
    ng1958 <= n1556;
    ng1979 <= n1561;
    ng1874 <= n1566;
    ng1914 <= n1571;
    ng2020 <= n1576;
    ng2080 <= n1581;
    ng2113 <= n1586;
    ng2209 <= n1591;
    ng2239 <= n1596;
    ng2250 <= n1601;
    ng2306 <= n1606;
    ng2285 <= n1611;
    ng2348 <= n1616;
    ng2256 <= n1621;
    ng2444 <= n1626;
    ng2489 <= n1631;
    ng2395 <= n1636;
    ng2529 <= n1641;
    ng2457 <= n1646;
    ng2587 <= n1651;
    ng2646 <= n1656;
    ng2530 <= n1661;
    ng2617 <= n1666;
    ng2654 <= n1671;
    ng2720 <= n1676;
    ng2777 <= n1681;
    ng2795 <= n1686;
    ng2810 <= n1691;
    ng3046 <= n1696;
    ng3100 <= n1701;
    ng3155 <= n1706;
    ng3182 <= n1711;
    ng3120 <= n1716;
    ng162 <= n1721;
    ng174 <= n1726;
    ng222 <= n1731;
    ng79 <= n1736;
    ng346 <= n1741;
    ng391 <= n1746;
    ng319 <= n1751;
    ng451 <= n1755;
    ng284 <= n1760;
    ng383 <= n1763;
    ng510 <= n1768;
    ng573 <= n1772;
    ng488 <= n1777;
    ng544 <= n1781;
    ng579 <= n1786;
    ng587 <= n1791;
    ng605 <= n1796;
    ng666 <= n1801;
    ng701 <= n1806;
    ng710 <= n1811;
    ng719 <= n1816;
    ng739 <= n1821;
    ng822 <= n1826;
    ng837 <= n1831;
    ng846 <= n1836;
    ng888 <= n1841;
    ng942 <= n1846;
    ng915 <= n1851;
    ng758 <= n1856;
    ng1095 <= n1861;
    ng1116 <= n1866;
    ng999 <= n1871;
    ng1009 <= n1876;
    ng1036 <= n1880;
    ng1054 <= n1885;
    ng1081 <= n1889;
    ng1142 <= n1894;
    ng1152 <= n1899;
    ng1235 <= n1904;
    ng1264 <= n1908;
    ng1215 <= n1913;
    ng1217 <= n1918;
    ng1312 <= n1923;
    ng1406 <= n1927;
    ng1415 <= n1932;
    ng1424 <= n1937;
    ng1524 <= n1942;
    ng1538 <= n1947;
    ng1550 <= n1952;
    ng1555 <= n1957;
    ng1439 <= n1962;
    ng1742 <= n1967;
    ng1795 <= n1972;
    ng1816 <= n1977;
    ng1704 <= n1982;
    ng1835 <= n1987;
    ng1904 <= n1990;
    ng1946 <= n1995;
    ng1842 <= n1999;
    ng1852 <= n2004;
    ng1962 <= n2009;
    ng1976 <= n2014;
    ng1877 <= n2019;
    ng1913 <= n2024;
    ng2013 <= n2029;
    ng2079 <= n2034;
    ng2111 <= n2039;
    ng2205 <= n2044;
    ng2240 <= n2049;
    ng2252 <= n2054;
    ng2309 <= n2059;
    ng2282 <= n2064;
    ng2160 <= n2069;
    ng2120 <= n2074;
    ng2433 <= n2079;
    ng2486 <= n2084;
    ng2397 <= n2089;
    ng2528 <= n2094;
    ng2458 <= n2098;
    ng2584 <= n2103;
    ng2647 <= n2107;
    ng2563 <= n2112;
    ng2618 <= n2116;
    ng2653 <= n2121;
    ng2734 <= n2126;
    ng2776 <= n2131;
    ng2785 <= n2136;
    ng2808 <= n2141;
    ng3045 <= n2146;
    ng2900 <= n2151;
    ng3093 <= n2156;
    ng3104 <= n2161;
    ng3173 <= n2166;
    ng3123 <= n2171;
    ng195 <= n2176;
    ng255 <= n2181;
    ng270 <= n2186;
    ng52 <= n2191;
    ng388 <= n2196;
    ng298 <= n2201;
    ng367 <= n2206;
    ng570 <= n2211;
    ng487 <= n2216;
    ng529 <= n2221;
    ng659 <= n2226;
    ng721 <= n2231;
    ng737 <= n2236;
    ng856 <= n2241;
    ng876 <= n2246;
    ng1098 <= n2251;
    ng1125 <= n2256;
    ng1141 <= n2261;
    ng976 <= n2266;
    ng1145 <= n2271;
    ng1214 <= n2276;
    ng1263 <= n2281;
    ng1282 <= n2286;
    ng1183 <= n2291;
    ng1407 <= n2296;
    ng1418 <= n2301;
    ng1511 <= n2306;
    ng1531 <= n2311;
    ng1534 <= n2316;
    ng1545 <= n2321;
    ng1435 <= n2326;
    ng1757 <= n2331;
    ng1809 <= n2336;
    ng1693 <= n2341;
    ng1696 <= n2346;
    ng1783 <= n2351;
    ng1944 <= n2356;
    ng1870 <= n2361;
    ng1865 <= n2366;
    ng1929 <= n2371;
    ng1939 <= n2376;
    ng1966 <= n2381;
    ng1886 <= n2386;
    ng1917 <= n2391;
    ng2089 <= n2396;
    ng2100 <= n2401;
    ng2108 <= n2406;
    ng2207 <= n2411;
    ng2238 <= n2416;
    ng2255 <= n2421;
    ng2315 <= n2426;
    ng2294 <= n2431;
    ng2339 <= n2436;
    ng2142 <= n2441;
    ng2418 <= n2446;
    ng2483 <= n2451;
    ng2398 <= n2456;
    ng2355 <= n2461;
    ng2366 <= n2466;
    ng2439 <= n2471;
    ng2644 <= n2476;
    ng2562 <= n2481;
    ng2670 <= n2486;
    ng2571 <= n2491;
    ng2610 <= n2496;
    ng2812 <= n2501;
    ng3048 <= n2506;
    ng3094 <= n2511;
    ng3103 <= n2516;
    ng3176 <= n2521;
    ng3124 <= n2526;
    ng198 <= n2531;
    ng252 <= n2536;
    ng213 <= n2541;
    ng354 <= n2546;
    ng398 <= n2551;
    ng342 <= n2556;
    ng366 <= n2561;
    ng571 <= n2565;
    ng486 <= n2570;
    ng530 <= n2575;
    ng630 <= n2580;
    ng711 <= n2585;
    ng830 <= n2590;
    ng860 <= n2595;
    ng873 <= n2600;
    ng1101 <= n2605;
    ng1122 <= n2610;
    ng966 <= n2614;
    ng975 <= n2619;
    ng1148 <= n2623;
    ng1158 <= n2628;
    ng1270 <= n2633;
    ng1285 <= n2638;
    ng1180 <= n2643;
    ng1405 <= n2648;
    ng1414 <= n2653;
    ng1515 <= n2658;
    ng1530 <= n2663;
    ng1532 <= n2668;
    ng1541 <= n2673;
    ng1430 <= n2678;
    ng1754 <= n2683;
    ng1807 <= n2688;
    ng1828 <= n2693;
    ng1697 <= n2698;
    ng1785 <= n2703;
    ng1949 <= n2707;
    ng1948 <= n2712;
    ng1845 <= n2716;
    ng1928 <= n2721;
    ng1956 <= n2726;
    ng1965 <= n2731;
    ng1887 <= n2736;
    ng1916 <= n2741;
    ng2087 <= n2746;
    ng2096 <= n2751;
    ng2112 <= n2756;
    ng2206 <= n2761;
    ng2245 <= n2766;
    ng2254 <= n2771;
    ng2318 <= n2776;
    ng2291 <= n2781;
    ng2297 <= n2786;
    ng2147 <= n2791;
    ng2421 <= n2796;
    ng2466 <= n2801;
    ng2396 <= n2806;
    ng2354 <= n2810;
    ng2374 <= n2815;
    ng2432 <= n2820;
    ng2645 <= n2823;
    ng2561 <= n2828;
    ng2652 <= n2833;
    ng2580 <= n2838;
    ng2608 <= n2843;
    ng2813 <= n2848;
    ng3047 <= n2853;
    ng3095 <= n2858;
    ng3106 <= n2863;
    ng3167 <= n2868;
    ng3125 <= n2873;
    ng216 <= n2878;
    ng92 <= n2883;
    ng376 <= n2888;
    ng349 <= n2892;
    ng372 <= n2897;
    ng324 <= n2902;
    ng531 <= n2907;
    ng633 <= n2912;
    ng698 <= n2917;
    ng840 <= n2922;
    ng861 <= n2927;
    ng918 <= n2932;
    ng1002 <= n2937;
    ng1089 <= n2942;
    ng967 <= n2947;
    ng978 <= n2952;
    ng1164 <= n2957;
    ng1245 <= n2961;
    ng1272 <= n2966;
    ng1288 <= n2971;
    ng1193 <= n2976;
    ng1409 <= n2981;
    ng1417 <= n2986;
    ng1512 <= n2991;
    ng1526 <= n2996;
    ng1536 <= n3001;
    ng1544 <= n3006;
    ng1426 <= n3011;
    ng1769 <= n3016;
    ng1804 <= n3021;
    ng1830 <= n3026;
    ng1698 <= n3031;
    ng1832 <= n3036;
    ng1950 <= n3041;
    ng1868 <= n3046;
    ng1860 <= n3051;
    ng1924 <= n3056;
    ng1957 <= n3061;
    ng1967 <= n3066;
    ng2040 <= n3071;
    ng2081 <= n3076;
    ng2091 <= n3081;
    ng2099 <= n3086;
    ng2109 <= n3091;
    ng2117 <= n3096;
    ng2246 <= n3101;
    ng2261 <= n3106;
    ng2273 <= n3111;
    ng2288 <= n3116;
    ng2300 <= n3121;
    ng2133 <= n3126;
    ng2384 <= n3131;
    ng2463 <= n3136;
    ng2478 <= n3141;
    ng2357 <= n3146;
    ng2364 <= n3150;
    ng2428 <= n3155;
    ng2447 <= n3160;
    ng2399 <= n3165;
    ng2656 <= n3170;
    ng2676 <= n3175;
    ng2607 <= n3180;
    ng2811 <= n3185;
    ng3096 <= n3190;
    ng3105 <= n3195;
    ng3170 <= n3200;
    ng3126 <= n3205;
    ng219 <= n3210;
    ng273 <= n3215;
    ng56 <= n3220;
    ng368 <= n3224;
    ng379 <= n3228;
    ng397 <= n3233;
    ng532 <= n3237;
    ng640 <= n3242;
    ng653 <= n3247;
    ng847 <= n3252;
    ng859 <= n3257;
    ng879 <= n3262;
    ng1003 <= n3267;
    ng1091 <= n3272;
    ng968 <= n3276;
    ng977 <= n3281;
    ng1221 <= n3284;
    ng1262 <= n3289;
    ng1271 <= n3294;
    ng1300 <= n3299;
    ng1192 <= n3304;
    ng1410 <= n3309;
    ng1419 <= n3314;
    ng1513 <= n3319;
    ng1528 <= n3324;
    ng1537 <= n3329;
    ng1546 <= n3334;
    ng1735 <= n3339;
    ng1779 <= n3344;
    ng1808 <= n3349;
    ng1829 <= n3354;
    ng1699 <= n3359;
    ng1831 <= n3364;
    ng1951 <= n3367;
    ng1867 <= n3372;
    ng1861 <= n3377;
    ng1923 <= n3382;
    ng1955 <= n3386;
    ng1964 <= n3391;
    ng2052 <= n3396;
    ng2083 <= n3401;
    ng2092 <= n3406;
    ng2101 <= n3411;
    ng2110 <= n3416;
    ng2119 <= n3421;
    ng2244 <= n3426;
    ng2253 <= n3431;
    ng2276 <= n3436;
    ng2330 <= n3441;
    ng2303 <= n3446;
    ng2138 <= n3451;
    ng2429 <= n3456;
    ng2473 <= n3461;
    ng2479 <= n3466;
    ng2356 <= n3470;
    ng2365 <= n3475;
    ng2427 <= n3479;
    ng2454 <= n3482;
    ng2472 <= n3487;
    ng2657 <= n3491;
    ng2673 <= n3496;
    ng2568 <= n3501;
    ng3049 <= n3506;
    ng2888 <= n3511;
    ng130 <= n3516;
    ng144 <= n3521;
    ng158 <= n3526;
    ng172 <= n3531;
    ng192 <= n3536;
    ng207 <= n3541;
    ng449 <= n3546;
    ng322 <= n3551;
    ng279 <= n3556;
    ng290 <= n3561;
    ng357 <= n3566;
    ng578 <= n3571;
    ng599 <= n3576;
    ng506 <= n3581;
    ng537 <= n3586;
    ng700 <= n3591;
    ng838 <= n3596;
    ng852 <= n3601;
    ng866 <= n3606;
    ng894 <= n3611;
    ng909 <= n3616;
    ng1137 <= n3621;
    ng972 <= n3626;
    ng1044 <= n3631;
    ng1070 <= n3636;
    ng1209 <= n3641;
    ng1294 <= n3645;
    ng1223 <= n3650;
    ng1332 <= n3655;
    ng1389 <= n3660;
    ng1400 <= n3665;
    ng1560 <= n3670;
    ng1582 <= n3675;
    ng1597 <= n3680;
    ng1466 <= n3685;
    ng1666 <= n3690;
    ng1730 <= n3695;
    ng1753 <= n3700;
    ng1705 <= n3705;
    ng2217 <= n3710;
    ng2231 <= n3715;
    ng2248 <= n3720;
    ng2503 <= n3725;
    ng2387 <= n3730;
    ng2477 <= n3735;
    ng2359 <= n3740;
    ng2417 <= n3745;
    ng2443 <= n3750;
    ng2655 <= n3755;
    ng2691 <= n3760;
    ng2599 <= n3765;
    ng2704 <= n3770;
    ng2766 <= n3775;
    ng2783 <= n3780;
    ng2794 <= n3785;
    ng3050 <= n3790;
    ng3062 <= n3795;
    ng3073 <= n3800;
    ng3013 <= n3805;
    ng45 <= n3810;
    ng20 <= n3815;
    ng2896 <= n3820;
    ng131 <= n3825;
    ng146 <= n3830;
    ng156 <= n3835;
    ng168 <= n3840;
    ng231 <= n3845;
    ng204 <= n3850;
    ng427 <= n3855;
    ng323 <= n3860;
    ng454 <= n3865;
    ng291 <= n3868;
    ng353 <= n3873;
    ng582 <= n3878;
    ng596 <= n3883;
    ng507 <= n3888;
    ng536 <= n3893;
    ng707 <= n3898;
    ng831 <= n3903;
    ng850 <= n3908;
    ng862 <= n3913;
    ng897 <= n3918;
    ng951 <= n3923;
    ng1138 <= n3927;
    ng971 <= n3932;
    ng1051 <= n3935;
    ng1069 <= n3940;
    ng1252 <= n3944;
    ng1273 <= n3949;
    ng1224 <= n3954;
    ng1339 <= n3959;
    ng1387 <= n3964;
    ng1396 <= n3969;
    ng1561 <= n3974;
    ng1579 <= n3979;
    ng1600 <= n3984;
    ng1654 <= n3989;
    ng1667 <= n3994;
    ng1723 <= n3999;
    ng1760 <= n4002;
    ng1778 <= n4007;
    ng2221 <= n4011;
    ng2230 <= n4016;
    ng2264 <= n4021;
    ng2501 <= n4026;
    ng2522 <= n4031;
    ng2525 <= n4036;
    ng2358 <= n4040;
    ng2424 <= n4044;
    ng2442 <= n4049;
    ng2659 <= n4053;
    ng2688 <= n4058;
    ng2603 <= n4063;
    ng2615 <= n4068;
    ng2773 <= n4073;
    ng2782 <= n4078;
    ng2804 <= n4083;
    ng3051 <= n4088;
    ng3061 <= n4093;
    ng3074 <= n4098;
    ng3002 <= n4103;
    ng42 <= n4108;
    ng23 <= n4113;
    ng2892 <= n4118;
    ng129 <= n4123;
    ng149 <= n4128;
    ng153 <= n4133;
    ng170 <= n4138;
    ng234 <= n4143;
    ng249 <= n4148;
    ng428 <= n4153;
    ng312 <= n4158;
    ng453 <= n4162;
    ng299 <= n4167;
    ng365 <= n4172;
    ng484 <= n4176;
    ng549 <= n4181;
    ng520 <= n4186;
    ng541 <= n4191;
    ng720 <= n4196;
    ng826 <= n4201;
    ng857 <= n4206;
    ng865 <= n4211;
    ng767 <= n4216;
    ng1045 <= n4221;
    ng1139 <= n4226;
    ng974 <= n4231;
    ng1052 <= n4236;
    ng1196 <= n4240;
    ng1251 <= n4245;
    ng1276 <= n4250;
    ng1177 <= n4255;
    ng1227 <= n4260;
    ng1358 <= n4265;
    ng1384 <= n4270;
    ng1398 <= n4275;
    ng1529 <= n4280;
    ng1543 <= n4285;
    ng1559 <= n4290;
    ng1624 <= n4295;
    ng1636 <= n4300;
    ng1651 <= n4305;
    ng1784 <= n4310;
    ng1668 <= n4314;
    ng1732 <= n4319;
    ng1748 <= n4324;
    ng1777 <= n4329;
    ng2222 <= n4334;
    ng2233 <= n4339;
    ng2321 <= n4344;
    ng2504 <= n4349;
    ng2389 <= n4354;
    ng2526 <= n4358;
    ng2361 <= n4363;
    ng2380 <= n4367;
    ng2441 <= n4372;
    ng2559 <= n4377;
    ng2623 <= n4382;
    ng2660 <= n4387;
    ng2679 <= n4392;
    ng2581 <= n4397;
    ng2612 <= n4402;
    ng2774 <= n4407;
    ng2792 <= n4412;
    ng2803 <= n4417;
    ng3052 <= n4422;
    ng3064 <= n4427;
    ng3071 <= n4432;
    ng3006 <= n4437;
    ng39 <= n4442;
    ng11 <= n4447;
    ng1 <= n4452;
    ng2903 <= n4457;
    ng133 <= n4462;
    ng148 <= n4467;
    ng157 <= n4472;
    ng169 <= n4477;
    ng237 <= n4482;
    ng210 <= n4487;
    ng426 <= n4492;
    ng447 <= n4497;
    ng320 <= n4502;
    ng305 <= n4507;
    ng364 <= n4511;
    ng464 <= n4516;
    ng548 <= n4521;
    ng525 <= n4525;
    ng538 <= n4530;
    ng730 <= n4535;
    ng728 <= n4540;
    ng858 <= n4545;
    ng867 <= n4550;
    ng762 <= n4555;
    ng1056 <= n4560;
    ng1140 <= n4564;
    ng973 <= n4569;
    ng1074 <= n4573;
    ng1199 <= n4577;
    ng1260 <= n4581;
    ng1279 <= n4585;
    ng1297 <= n4590;
    ng1309 <= n4595;
    ng1346 <= n4599;
    ng1388 <= n4604;
    ng1397 <= n4609;
    ng1533 <= n4614;
    ng1542 <= n4619;
    ng1567 <= n4624;
    ng1621 <= n4629;
    ng1594 <= n4634;
    ng1648 <= n4639;
    ng1695 <= n4644;
    ng1669 <= n4649;
    ng1731 <= n4654;
    ng1749 <= n4657;
    ng1776 <= n4662;
    ng2220 <= n4666;
    ng2229 <= n4671;
    ng2333 <= n4676;
    ng2507 <= n4681;
    ng2388 <= n4686;
    ng2527 <= n4691;
    ng2360 <= n4694;
    ng2373 <= n4699;
    ng2440 <= n4704;
    ng2539 <= n4708;
    ng2622 <= n4713;
    ng2658 <= n4718;
    ng2694 <= n4723;
    ng2594 <= n4728;
    ng2611 <= n4732;
    ng2781 <= n4737;
    ng2790 <= n4742;
    ng2799 <= n4747;
    ng3053 <= n4752;
    ng3063 <= n4757;
    ng3072 <= n4762;
    ng2998 <= n4767;
    ng27 <= n4772;
    ng17 <= n4777;
    ng2817 <= n4782;
    ng3101 <= n4787;
    ng3164 <= n4792;
    ng134 <= n4797;
    ng151 <= n4802;
    ng159 <= n4807;
    ng176 <= n4812;
    ng179 <= n4817;
    ng240 <= n4822;
    ng225 <= n4827;
    ng65 <= n4832;
    ng373 <= n4837;
    ng429 <= n4842;
    ng314 <= n4847;
    ng404 <= n4852;
    ng283 <= n4857;
    ng350 <= n4862;
    ng387 <= n4867;
    ng524 <= n4872;
    ng568 <= n4877;
    ng480 <= n4882;
    ng465 <= n4887;
    ng558 <= n4892;
    ng585 <= n4897;
    ng620 <= n4902;
    ng679 <= n4907;
    ng704 <= n4912;
    ng718 <= n4917;
    ng729 <= n4922;
    ng732 <= n4927;
    ng853 <= n4932;
    ng834 <= n4937;
    ng845 <= n4942;
    ng927 <= n4947;
    ng906 <= n4952;
    ng776 <= n4957;
    ng1033 <= n4962;
    ng1048 <= n4967;
    ng1107 <= n4972;
    ng1135 <= n4977;
    ng1007 <= n4982;
    ng1037 <= n4987;
    ng1066 <= n4992;
    ng1240 <= n4997;
    ng1259 <= n5002;
    ng1165 <= n5007;
    ng1229 <= n5012;
    ng1266 <= n5017;
    ng1218 <= n5022;
    ng1345 <= n5027;
    ng1385 <= n5032;
    ng1393 <= n5037;
    ng1421 <= n5042;
    ng1514 <= n5047;
    ng1553 <= n5052;
    ng1615 <= n5057;
    ng1630 <= n5062;
    ng1609 <= n5067;
    ng1813 <= n5072;
    ng1662 <= n5077;
    ng1680 <= n5082;
    ng1746 <= n5087;
    ng1775 <= n5092;
    ng2224 <= n5097;
    ng2232 <= n5102;
    ng2156 <= n5107;
    ng2510 <= n5112;
    ng2391 <= n5117;
    ng2462 <= n5122;
    ng2598 <= n5127;
    ng2642 <= n5132;
    ng2555 <= n5137;
    ng2540 <= n5142;
    ng2632 <= n5147;
    ng2661 <= n5152;
    ng2685 <= n5157;
    ng2606 <= n5162;
    ng2746 <= n5167;
    ng2779 <= n5172;
    ng2787 <= n5177;
    ng2801 <= n5182;
    ng3054 <= n5187;
    ng3055 <= n5192;
    ng3066 <= n5197;
    ng3077 <= n5202;
    ng3028 <= n5207;
    ng3040 <= n5212;
    ng3083 <= n5217;
    ng2990 <= n5222;
    ng2933 <= n5227;
    ng3102 <= n5232;
    ng3161 <= n5237;
    ng132 <= n5242;
    ng147 <= n5247;
    ng163 <= n5252;
    ng175 <= n5257;
    ng177 <= n5262;
    ng201 <= n5267;
    ng228 <= n5272;
    ng70 <= n5277;
    ng423 <= n5282;
    ng432 <= n5287;
    ng313 <= n5292;
    ng402 <= n5297;
    ng282 <= n5302;
    ng287 <= n5305;
    ng394 <= n5309;
    ng523 <= n5313;
    ng489 <= n5316;
    ng479 <= n5321;
    ng468 <= n5326;
    ng499 <= n5330;
    ng586 <= n5335;
    ng617 <= n5340;
    ng686 <= n5345;
    ng706 <= n5350;
    ng716 <= n5355;
    ng725 <= n5360;
    ng733 <= n5365;
    ng823 <= n5369;
    ng832 <= n5373;
    ng841 <= n5378;
    ng930 <= n5383;
    ng903 <= n5388;
    ng771 <= n5393;
    ng1030 <= n5398;
    ng1071 <= n5403;
    ng1104 <= n5408;
    ng1136 <= n5413;
    ng1006 <= n5418;
    ng1038 <= n5422;
    ng1059 <= n5427;
    ng1243 <= n5431;
    ng1258 <= n5436;
    ng1253 <= n5439;
    ng1230 <= n5443;
    ng1265 <= n5448;
    ng1219 <= n5453;
    ng1316 <= n5458;
    ng1386 <= n5463;
    ng1395 <= n5468;
    ng1422 <= n5473;
    ng1516 <= n5478;
    ng1557 <= n5483;
    ng1612 <= n5488;
    ng1633 <= n5493;
    ng1606 <= n5498;
    ng1789 <= n5503;
    ng1663 <= n5508;
    ng1672 <= n5513;
    ng1747 <= n5517;
    ng1768 <= n5522;
    ng2225 <= n5526;
    ng2234 <= n5531;
    ng2258 <= n5535;
    ng2513 <= n5540;
    ng2390 <= n5545;
    ng2469 <= n5549;
    ng2597 <= n5553;
    ng2564 <= n5556;
    ng2554 <= n5561;
    ng2543 <= n5566;
    ng2574 <= n5570;
    ng2664 <= n5575;
    ng2682 <= n5580;
    ng2707 <= n5585;
    ng2740 <= n5590;
    ng2775 <= n5595;
    ng2791 <= n5600;
    ng2800 <= n5605;
    ng2802 <= n5610;
    ng3056 <= n5615;
    ng3065 <= n5620;
    ng3078 <= n5625;
    ng3018 <= n5630;
    ng2986 <= n5634;
    ng36 <= n5639;
    ng2991 <= n5644;
    ng2950 <= n5649;
    ng3191 <= n5654;
    ng185 <= n5659;
    ng142 <= n5664;
    ng150 <= n5669;
    ng160 <= n5674;
    ng171 <= n5679;
    ng186 <= n5684;
    ng246 <= n5689;
    ng267 <= n5694;
    ng361 <= n5699;
    ng420 <= n5704;
    ng435 <= n5709;
    ng316 <= n5714;
    ng321 <= n5719;
    ng281 <= n5724;
    ng288 <= n5729;
    ng352 <= n5734;
    ng395 <= n5738;
    ng569 <= n5743;
    ng566 <= n5748;
    ng478 <= n5753;
    ng471 <= n5758;
    ng576 <= n5763;
    ng583 <= n5768;
    ng614 <= n5773;
    ng493 <= n5778;
    ng534 <= n5783;
    ng692 <= n5788;
    ng709 <= n5793;
    ng713 <= n5798;
    ng727 <= n5803;
    ng731 <= n5808;
    ng819 <= n5813;
    ng829 <= n5818;
    ng843 <= n5823;
    ng864 <= n5828;
    ng933 <= n5833;
    ng948 <= n5838;
    ng960 <= n5843;
    ng1041 <= n5848;
    ng1060 <= n5853;
    ng1114 <= n5858;
    ng1128 <= n5863;
    ng1005 <= n5868;
    ng1039 <= n5873;
    ng1068 <= n5878;
    ng1084 <= n5883;
    ng1257 <= n5888;
    ng1254 <= n5893;
    ng1167 <= n5898;
    ng1261 <= n5903;
    ng1220 <= n5908;
    ng1319 <= n5913;
    ng1372 <= n5918;
    ng1394 <= n5923;
    ng1401 <= n5928;
    ng1412 <= n5933;
    ng1558 <= n5938;
    ng1576 <= n5943;
    ng1588 <= n5948;
    ng1603 <= n5953;
    ng1727 <= n5958;
    ng1664 <= n5962;
    ng1679 <= n5967;
    ng1738 <= n5972;
    ng1764 <= n5977;
    ng2448 <= n5982;
    ng2516 <= n5987;
    ng2393 <= n5992;
    ng2470 <= n5997;
    ng2643 <= n6002;
    ng2640 <= n6007;
    ng2553 <= n6012;
    ng2546 <= n6017;
    ng2650 <= n6022;
    ng2667 <= n6027;
    ng2604 <= n6032;
    ng2714 <= n6037;
    ng2753 <= n6042;
    ng2778 <= n6047;
    ng2788 <= n6052;
    ng2796 <= n6057;
    ng2806 <= n6062;
    ng3080 <= n6067;
    ng3057 <= n6072;
    ng3068 <= n6077;
    ng3075 <= n6082;
    ng3024 <= n6087;
    ng2987 <= n6092;
    ng2992 <= n6097;
    ng8 <= n6102;
    ng2883 <= n6107;
    ng3128 <= n6112;
    ng3147 <= n6117;
    ng143 <= n6122;
    ng152 <= n6127;
    ng161 <= n6132;
    ng173 <= n6137;
    ng189 <= n6142;
    ng243 <= n6147;
    ng61 <= n6152;
    ng384 <= n6157;
    ng417 <= n6162;
    ng438 <= n6167;
    ng315 <= n6172;
    ng403 <= n6177;
    ng280 <= n6182;
    ng289 <= n6185;
    ng351 <= n6189;
    ng396 <= n6193;
    ng564 <= n6198;
    ng567 <= n6201;
    ng477 <= n6206;
    ng528 <= n6211;
    ng559 <= n6214;
    ng581 <= n6219;
    ng602 <= n6224;
    ng496 <= n6229;
    ng533 <= n6234;
    ng699 <= n6239;
    ng708 <= n6244;
    ng717 <= n6249;
    ng726 <= n6254;
    ng735 <= n6259;
    ng818 <= n6264;
    ng833 <= n6269;
    ng842 <= n6274;
    ng851 <= n6279;
    ng891 <= n6284;
    ng945 <= n6289;
    ng780 <= n6294;
    ng740 <= n6299;
    ng1063 <= n6304;
    ng1110 <= n6309;
    ng1131 <= n6314;
    ng1004 <= n6319;
    ng1040 <= n6323;
    ng1067 <= n6328;
    ng1011 <= n6331;
    ng1256 <= n6336;
    ng1176 <= n6339;
    ng1166 <= n6344;
    ng1228 <= n6348;
    ng1222 <= n6353;
    ng1326 <= n6358;
    ng1378 <= n6363;
    ng1390 <= n6368;
    ng1399 <= n6373;
    ng1408 <= n6378;
    ng1556 <= n6383;
    ng1618 <= n6388;
    ng1591 <= n6393;
    ng1645 <= n6398;
    ng1457 <= n6403;
    ng1665 <= n6408;
    ng1686 <= n6412;
    ng1745 <= n6416;
    ng1763 <= n6421;
    ng2498 <= n6425;
    ng2519 <= n6430;
    ng2392 <= n6435;
    ng2471 <= n6439;
    ng2638 <= n6444;
    ng2641 <= n6447;
    ng2552 <= n6452;
    ng2602 <= n6457;
    ng2633 <= n6460;
    ng2565 <= n6465;
    ng2605 <= n6470;
    ng2733 <= n6475;
    ng2760 <= n6480;
    ng2780 <= n6485;
    ng2789 <= n6490;
    ng2798 <= n6495;
    ng2807 <= n6500;
    ng3079 <= n6505;
    ng3058 <= n6510;
    ng3067 <= n6515;
    ng3076 <= n6520;
    ng3010 <= n6525;
    ng48 <= n6530;
    ng26 <= n6535;
    ng2 <= n6540;
    ng809 <= n6545;
    ng2827 <= n6550;
    ng113 <= n6555;
    ng2200 <= n6560;
    ng3084 <= n6565;
    ng3059 <= n6570;
    ng3070 <= n6575;
    ng2867 <= n6580;
    ng789 <= n6585;
    ng2845 <= n6590;
    ng2857 <= n6595;
    ng3085 <= n6600;
    ng3060 <= n6605;
    ng3069 <= n6610;
    ng805 <= n6614;
    ng2830 <= n6619;
    ng117 <= n6624;
    ng2858 <= n6629;
    ng3086 <= n6633;
    ng2997 <= n6638;
    ng3032 <= n6643;
    ng2814 <= n6648;
    ng2870 <= n6653;
    ng785 <= n6657;
    ng2842 <= n6662;
    ng97 <= n6666;
    ng3087 <= n6671;
    ng2993 <= n6676;
    ng3036 <= n6681;
    ng2908 <= n6686;
    ng2935 <= n6691;
    ng2969 <= n6696;
    ng1481 <= n6701;
    ng3091 <= n6706;
    ng1570 <= n6711;
    ng1670 <= n6715;
    ng1734 <= n6720;
    ng2210 <= n6725;
    ng2227 <= n6730;
    ng30 <= n6735;
    ng5 <= n6740;
    ng2912 <= n6745;
    ng2934 <= n6750;
    ng2972 <= n6755;
    ng1486 <= n6760;
    ng3092 <= n6765;
    ng1627 <= n6770;
    ng1671 <= n6775;
    ng1733 <= n6779;
    ng2208 <= n6783;
    ng2223 <= n6788;
    ng33 <= n6793;
    ng14 <= n6798;
    ng2917 <= n6803;
    ng2941 <= n6808;
    ng2963 <= n6813;
    ng1491 <= n6818;
    ng1639 <= n6823;
    ng1761 <= n6828;
    ng1937 <= n6833;
    ng2218 <= n6838;
    ng2226 <= n6843;
    ng2524 <= n6848;
    ng2924 <= n6853;
    ng2938 <= n6858;
    ng2966 <= n6863;
    ng1496 <= n6868;
    ng1462 <= n6873;
    ng1762 <= n6877;
    ng1934 <= n6882;
    ng2219 <= n6887;
    ng2228 <= n6892;
    ng2502 <= n6897;
    ng2920 <= n6902;
    ng2947 <= n6907;
    ng2981 <= n6912;
    ng2861 <= n6917;
    ng793 <= n6922;
    ng2839 <= n6927;
    ng1724 <= n6931;
    ng1952 <= n6936;
    ng1836 <= n6941;
    ng2085 <= n6946;
    ng2093 <= n6951;
    ng2107 <= n6956;
    ng2118 <= n6961;
    ng2451 <= n6966;
    ng2984 <= n6971;
    ng2944 <= n6976;
    ng2874 <= n6981;
    ng2877 <= n6986;
    ng2824 <= n6991;
    ng121 <= n6995;
    ng1772 <= n7000;
    ng1953 <= n7004;
    ng1869 <= n7009;
    ng2086 <= n7014;
    ng2095 <= n7019;
    ng2105 <= n7024;
    ng2114 <= n7029;
    ng2257 <= n7033;
    ng2985 <= n7038;
    ng2956 <= n7043;
    ng2975 <= n7048;
    ng1471 <= n7053;
    ng101 <= n7058;
    ng2170 <= n7063;
    ng1810 <= n7068;
    ng1846 <= n7073;
    ng1938 <= n7078;
    ng2084 <= n7082;
    ng2098 <= n7087;
    ng2102 <= n7092;
    ng2116 <= n7097;
    ng2151 <= n7102;
    ng2930 <= n7107;
    ng2953 <= n7112;
    ng2978 <= n7117;
    ng1476 <= n7122;
    ng2854 <= n7127;
    ng2175 <= n7131;
    ng1694 <= n7136;
    ng1849 <= n7141;
    ng1880 <= n7145;
    ng2088 <= n7150;
    ng2097 <= n7155;
    ng2106 <= n7160;
    ng2115 <= n7165;
    ng2336 <= n7170;
    ng2929 <= n7174;
    ng2962 <= n7179;
    ng801 <= n7183;
    ng2833 <= n7188;
    ng105 <= n7193;
    ng2180 <= n7198;
    ng2165 <= n7203;
    ng1702 <= n7208;
    ng1963 <= n7213;
    ng1994 <= n7218;
    ng1997 <= n7223;
    ng1905 <= n7228;
    ng2010 <= n7233;
    ng2072 <= n7238;
    ng2279 <= n7243;
    ng2879 <= n7248;
    ng2959 <= n7253;
    ng2818 <= n7258;
    ng2873 <= n7262;
    ng2851 <= n7267;
    ng2185 <= n7271;
    ng2878 <= n7276;
    ng1661 <= n7281;
    ng1961 <= n7285;
    ng1982 <= n7290;
    ng2000 <= n7295;
    ng1900 <= n7300;
    ng2039 <= n7304;
    ng2066 <= n7309;
    ng2267 <= n7314;
    ng1506 <= n7319;
    ng2864 <= n7324;
    ng797 <= n7327;
    ng2836 <= n7332;
    ng109 <= n7335;
    ng2190 <= n7340;
    ng3210 <= n7345;
    ng1985 <= n7350;
    ng1910 <= n7355;
    ng1918 <= n7360;
    ng2059 <= n7365;
    ng2249 <= n7370;
    ng1501 <= n7375;
    ng813 <= n7379;
    ng2821 <= n7384;
    ng125 <= n7387;
    ng2848 <= n7392;
    ng2195 <= n7396;
    ng3211 <= n7401;
    ng1988 <= n7406;
    ng1909 <= n7411;
    ng1921 <= n7416;
    ng2046 <= n7421;
    ng2236 <= n7426;
  end
endmodule

