// Benchmark "top" written by ABC on Thu Oct  8 22:51:56 2020

module top ( 
    \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
    \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
    \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
    \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
    \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
    \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
    \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
    \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
    \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
    \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
    \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
    \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
    \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
    \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
    \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
    \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
    \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
    \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
    \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
    \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
    \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
    \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
    \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
    \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
    \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
    \priority[100] , \priority[101] , \priority[102] , \priority[103] ,
    \priority[104] , \priority[105] , \priority[106] , \priority[107] ,
    \priority[108] , \priority[109] , \priority[110] , \priority[111] ,
    \priority[112] , \priority[113] , \priority[114] , \priority[115] ,
    \priority[116] , \priority[117] , \priority[118] , \priority[119] ,
    \priority[120] , \priority[121] , \priority[122] , \priority[123] ,
    \priority[124] , \priority[125] , \priority[126] , \priority[127] ,
    \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] , \req[6] ,
    \req[7] , \req[8] , \req[9] , \req[10] , \req[11] , \req[12] ,
    \req[13] , \req[14] , \req[15] , \req[16] , \req[17] , \req[18] ,
    \req[19] , \req[20] , \req[21] , \req[22] , \req[23] , \req[24] ,
    \req[25] , \req[26] , \req[27] , \req[28] , \req[29] , \req[30] ,
    \req[31] , \req[32] , \req[33] , \req[34] , \req[35] , \req[36] ,
    \req[37] , \req[38] , \req[39] , \req[40] , \req[41] , \req[42] ,
    \req[43] , \req[44] , \req[45] , \req[46] , \req[47] , \req[48] ,
    \req[49] , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
    \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60] ,
    \req[61] , \req[62] , \req[63] , \req[64] , \req[65] , \req[66] ,
    \req[67] , \req[68] , \req[69] , \req[70] , \req[71] , \req[72] ,
    \req[73] , \req[74] , \req[75] , \req[76] , \req[77] , \req[78] ,
    \req[79] , \req[80] , \req[81] , \req[82] , \req[83] , \req[84] ,
    \req[85] , \req[86] , \req[87] , \req[88] , \req[89] , \req[90] ,
    \req[91] , \req[92] , \req[93] , \req[94] , \req[95] , \req[96] ,
    \req[97] , \req[98] , \req[99] , \req[100] , \req[101] , \req[102] ,
    \req[103] , \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
    \req[109] , \req[110] , \req[111] , \req[112] , \req[113] , \req[114] ,
    \req[115] , \req[116] , \req[117] , \req[118] , \req[119] , \req[120] ,
    \req[121] , \req[122] , \req[123] , \req[124] , \req[125] , \req[126] ,
    \req[127] ,
    \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] , \grant[5] ,
    \grant[6] , \grant[7] , \grant[8] , \grant[9] , \grant[10] ,
    \grant[11] , \grant[12] , \grant[13] , \grant[14] , \grant[15] ,
    \grant[16] , \grant[17] , \grant[18] , \grant[19] , \grant[20] ,
    \grant[21] , \grant[22] , \grant[23] , \grant[24] , \grant[25] ,
    \grant[26] , \grant[27] , \grant[28] , \grant[29] , \grant[30] ,
    \grant[31] , \grant[32] , \grant[33] , \grant[34] , \grant[35] ,
    \grant[36] , \grant[37] , \grant[38] , \grant[39] , \grant[40] ,
    \grant[41] , \grant[42] , \grant[43] , \grant[44] , \grant[45] ,
    \grant[46] , \grant[47] , \grant[48] , \grant[49] , \grant[50] ,
    \grant[51] , \grant[52] , \grant[53] , \grant[54] , \grant[55] ,
    \grant[56] , \grant[57] , \grant[58] , \grant[59] , \grant[60] ,
    \grant[61] , \grant[62] , \grant[63] , \grant[64] , \grant[65] ,
    \grant[66] , \grant[67] , \grant[68] , \grant[69] , \grant[70] ,
    \grant[71] , \grant[72] , \grant[73] , \grant[74] , \grant[75] ,
    \grant[76] , \grant[77] , \grant[78] , \grant[79] , \grant[80] ,
    \grant[81] , \grant[82] , \grant[83] , \grant[84] , \grant[85] ,
    \grant[86] , \grant[87] , \grant[88] , \grant[89] , \grant[90] ,
    \grant[91] , \grant[92] , \grant[93] , \grant[94] , \grant[95] ,
    \grant[96] , \grant[97] , \grant[98] , \grant[99] , \grant[100] ,
    \grant[101] , \grant[102] , \grant[103] , \grant[104] , \grant[105] ,
    \grant[106] , \grant[107] , \grant[108] , \grant[109] , \grant[110] ,
    \grant[111] , \grant[112] , \grant[113] , \grant[114] , \grant[115] ,
    \grant[116] , \grant[117] , \grant[118] , \grant[119] , \grant[120] ,
    \grant[121] , \grant[122] , \grant[123] , \grant[124] , \grant[125] ,
    \grant[126] , \grant[127] , anyGrant  );
  input  \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
    \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
    \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
    \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
    \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
    \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
    \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
    \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
    \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
    \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
    \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
    \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
    \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
    \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
    \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
    \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
    \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
    \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
    \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
    \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
    \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
    \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
    \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
    \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
    \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
    \priority[100] , \priority[101] , \priority[102] , \priority[103] ,
    \priority[104] , \priority[105] , \priority[106] , \priority[107] ,
    \priority[108] , \priority[109] , \priority[110] , \priority[111] ,
    \priority[112] , \priority[113] , \priority[114] , \priority[115] ,
    \priority[116] , \priority[117] , \priority[118] , \priority[119] ,
    \priority[120] , \priority[121] , \priority[122] , \priority[123] ,
    \priority[124] , \priority[125] , \priority[126] , \priority[127] ,
    \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] , \req[6] ,
    \req[7] , \req[8] , \req[9] , \req[10] , \req[11] , \req[12] ,
    \req[13] , \req[14] , \req[15] , \req[16] , \req[17] , \req[18] ,
    \req[19] , \req[20] , \req[21] , \req[22] , \req[23] , \req[24] ,
    \req[25] , \req[26] , \req[27] , \req[28] , \req[29] , \req[30] ,
    \req[31] , \req[32] , \req[33] , \req[34] , \req[35] , \req[36] ,
    \req[37] , \req[38] , \req[39] , \req[40] , \req[41] , \req[42] ,
    \req[43] , \req[44] , \req[45] , \req[46] , \req[47] , \req[48] ,
    \req[49] , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
    \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60] ,
    \req[61] , \req[62] , \req[63] , \req[64] , \req[65] , \req[66] ,
    \req[67] , \req[68] , \req[69] , \req[70] , \req[71] , \req[72] ,
    \req[73] , \req[74] , \req[75] , \req[76] , \req[77] , \req[78] ,
    \req[79] , \req[80] , \req[81] , \req[82] , \req[83] , \req[84] ,
    \req[85] , \req[86] , \req[87] , \req[88] , \req[89] , \req[90] ,
    \req[91] , \req[92] , \req[93] , \req[94] , \req[95] , \req[96] ,
    \req[97] , \req[98] , \req[99] , \req[100] , \req[101] , \req[102] ,
    \req[103] , \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
    \req[109] , \req[110] , \req[111] , \req[112] , \req[113] , \req[114] ,
    \req[115] , \req[116] , \req[117] , \req[118] , \req[119] , \req[120] ,
    \req[121] , \req[122] , \req[123] , \req[124] , \req[125] , \req[126] ,
    \req[127] ;
  output \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] ,
    \grant[5] , \grant[6] , \grant[7] , \grant[8] , \grant[9] ,
    \grant[10] , \grant[11] , \grant[12] , \grant[13] , \grant[14] ,
    \grant[15] , \grant[16] , \grant[17] , \grant[18] , \grant[19] ,
    \grant[20] , \grant[21] , \grant[22] , \grant[23] , \grant[24] ,
    \grant[25] , \grant[26] , \grant[27] , \grant[28] , \grant[29] ,
    \grant[30] , \grant[31] , \grant[32] , \grant[33] , \grant[34] ,
    \grant[35] , \grant[36] , \grant[37] , \grant[38] , \grant[39] ,
    \grant[40] , \grant[41] , \grant[42] , \grant[43] , \grant[44] ,
    \grant[45] , \grant[46] , \grant[47] , \grant[48] , \grant[49] ,
    \grant[50] , \grant[51] , \grant[52] , \grant[53] , \grant[54] ,
    \grant[55] , \grant[56] , \grant[57] , \grant[58] , \grant[59] ,
    \grant[60] , \grant[61] , \grant[62] , \grant[63] , \grant[64] ,
    \grant[65] , \grant[66] , \grant[67] , \grant[68] , \grant[69] ,
    \grant[70] , \grant[71] , \grant[72] , \grant[73] , \grant[74] ,
    \grant[75] , \grant[76] , \grant[77] , \grant[78] , \grant[79] ,
    \grant[80] , \grant[81] , \grant[82] , \grant[83] , \grant[84] ,
    \grant[85] , \grant[86] , \grant[87] , \grant[88] , \grant[89] ,
    \grant[90] , \grant[91] , \grant[92] , \grant[93] , \grant[94] ,
    \grant[95] , \grant[96] , \grant[97] , \grant[98] , \grant[99] ,
    \grant[100] , \grant[101] , \grant[102] , \grant[103] , \grant[104] ,
    \grant[105] , \grant[106] , \grant[107] , \grant[108] , \grant[109] ,
    \grant[110] , \grant[111] , \grant[112] , \grant[113] , \grant[114] ,
    \grant[115] , \grant[116] , \grant[117] , \grant[118] , \grant[119] ,
    \grant[120] , \grant[121] , \grant[122] , \grant[123] , \grant[124] ,
    \grant[125] , \grant[126] , \grant[127] , anyGrant;
  wire new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1489_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_,
    new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_,
    new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_,
    new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_,
    new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_,
    new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_,
    new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_,
    new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_,
    new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_,
    new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_,
    new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_,
    new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_,
    new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_,
    new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_,
    new_n1839_, new_n1840_, new_n1842_, new_n1843_, new_n1844_, new_n1845_,
    new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_,
    new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_,
    new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_,
    new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_,
    new_n1924_, new_n1925_, new_n1926_, new_n1928_, new_n1929_, new_n1930_,
    new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_,
    new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_,
    new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_,
    new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_,
    new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_,
    new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_,
    new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_,
    new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_,
    new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_,
    new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2014_, new_n2015_,
    new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_,
    new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_,
    new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_,
    new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_,
    new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_,
    new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_,
    new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_,
    new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_,
    new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_,
    new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_,
    new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_,
    new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_,
    new_n2355_, new_n2356_, new_n2358_, new_n2359_, new_n2360_, new_n2361_,
    new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_,
    new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_,
    new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_,
    new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_,
    new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_,
    new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_,
    new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_,
    new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_,
    new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_,
    new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_,
    new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_,
    new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_,
    new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_,
    new_n2440_, new_n2441_, new_n2442_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_,
    new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_,
    new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_,
    new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_,
    new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_,
    new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_,
    new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_,
    new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_,
    new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_,
    new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_,
    new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_,
    new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_,
    new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_,
    new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_,
    new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_,
    new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_,
    new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_,
    new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_,
    new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_,
    new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_,
    new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_,
    new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_,
    new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_,
    new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_,
    new_n2871_, new_n2872_, new_n2874_, new_n2875_, new_n2876_, new_n2877_,
    new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_,
    new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_,
    new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_,
    new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_,
    new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_,
    new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_,
    new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_,
    new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_,
    new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_,
    new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_,
    new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_,
    new_n2956_, new_n2957_, new_n2958_, new_n2960_, new_n2961_, new_n2962_,
    new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_,
    new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_,
    new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_,
    new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_,
    new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_,
    new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_,
    new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_,
    new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_,
    new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_,
    new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_,
    new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_,
    new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_,
    new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_,
    new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3132_,
    new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_,
    new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_,
    new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_,
    new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_,
    new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_,
    new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_,
    new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_,
    new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_,
    new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_,
    new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_,
    new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_,
    new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_,
    new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_,
    new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_,
    new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_,
    new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_,
    new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_,
    new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_,
    new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_,
    new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_,
    new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_,
    new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_,
    new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_,
    new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_,
    new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_,
    new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_,
    new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_,
    new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_,
    new_n3302_, new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_,
    new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_,
    new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_,
    new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_,
    new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_,
    new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_,
    new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_,
    new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_,
    new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_,
    new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_,
    new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_,
    new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_,
    new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_,
    new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_,
    new_n3387_, new_n3388_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_,
    new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_,
    new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_,
    new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_,
    new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_,
    new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_,
    new_n3472_, new_n3473_, new_n3474_, new_n3476_, new_n3477_, new_n3478_,
    new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_,
    new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_,
    new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_,
    new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_,
    new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_,
    new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_,
    new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_,
    new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_,
    new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_,
    new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_,
    new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_,
    new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_,
    new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_,
    new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3648_,
    new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_,
    new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_,
    new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_,
    new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_,
    new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_,
    new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_,
    new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_,
    new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_,
    new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_,
    new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_,
    new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_,
    new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_,
    new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_,
    new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_,
    new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_,
    new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_,
    new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_,
    new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_,
    new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_,
    new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_,
    new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_,
    new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_,
    new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_,
    new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_,
    new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_,
    new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_,
    new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_,
    new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_,
    new_n3818_, new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_,
    new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_,
    new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_,
    new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_,
    new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_,
    new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_,
    new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_,
    new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_,
    new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_,
    new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_,
    new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_,
    new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_,
    new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_,
    new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_,
    new_n3903_, new_n3904_, new_n3906_, new_n3907_, new_n3908_, new_n3909_,
    new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_,
    new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_,
    new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_,
    new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_,
    new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_,
    new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_,
    new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_,
    new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_,
    new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_,
    new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_,
    new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_,
    new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_,
    new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_,
    new_n3988_, new_n3989_, new_n3990_, new_n3992_, new_n3993_, new_n3994_,
    new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_,
    new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_,
    new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_,
    new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_,
    new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_,
    new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_,
    new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_,
    new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_,
    new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_,
    new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_,
    new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_,
    new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_,
    new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_,
    new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_,
    new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4164_,
    new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_,
    new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_,
    new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_,
    new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_,
    new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_,
    new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_,
    new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_, new_n4255_,
    new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_, new_n4261_,
    new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_, new_n4267_,
    new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_, new_n4273_,
    new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_, new_n4279_,
    new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_,
    new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_,
    new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_, new_n4297_,
    new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4336_, new_n4337_, new_n4338_, new_n4339_, new_n4340_,
    new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_,
    new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_,
    new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_, new_n4358_,
    new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_, new_n4364_,
    new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_, new_n4370_,
    new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_, new_n4376_,
    new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_, new_n4382_,
    new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_, new_n4388_,
    new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_, new_n4394_,
    new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_, new_n4400_,
    new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_, new_n4406_,
    new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_, new_n4412_,
    new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_, new_n4418_,
    new_n4419_, new_n4420_, new_n4422_, new_n4423_, new_n4424_, new_n4425_,
    new_n4426_, new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_,
    new_n4432_, new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_,
    new_n4438_, new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_,
    new_n4444_, new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4449_,
    new_n4450_, new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_,
    new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_,
    new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_,
    new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_,
    new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_,
    new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_,
    new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_, new_n4491_,
    new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_, new_n4497_,
    new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_, new_n4503_,
    new_n4504_, new_n4505_, new_n4506_, new_n4508_, new_n4509_, new_n4510_,
    new_n4511_, new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_,
    new_n4517_, new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_,
    new_n4523_, new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_,
    new_n4529_, new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_,
    new_n4535_, new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_,
    new_n4541_, new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_,
    new_n4547_, new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_,
    new_n4553_, new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_,
    new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_,
    new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_,
    new_n4571_, new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_,
    new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_,
    new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_,
    new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_,
    new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_,
    new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_,
    new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_,
    new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_,
    new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_,
    new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_,
    new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_,
    new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_,
    new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_,
    new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4680_,
    new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_,
    new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_,
    new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_,
    new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_,
    new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_,
    new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_,
    new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_,
    new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_,
    new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_,
    new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_,
    new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_,
    new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_,
    new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_,
    new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_,
    new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_,
    new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_,
    new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_,
    new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_,
    new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_,
    new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_,
    new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_,
    new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_,
    new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_,
    new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_,
    new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_,
    new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_,
    new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_,
    new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_,
    new_n4850_, new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_,
    new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_,
    new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_,
    new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_,
    new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_,
    new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_,
    new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_,
    new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_,
    new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_,
    new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_,
    new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_,
    new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_,
    new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_,
    new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_,
    new_n4935_, new_n4936_, new_n4938_, new_n4939_, new_n4940_, new_n4941_,
    new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_,
    new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_,
    new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_,
    new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_,
    new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_,
    new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_,
    new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_,
    new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_,
    new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_,
    new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_,
    new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_,
    new_n5020_, new_n5021_, new_n5022_, new_n5024_, new_n5025_, new_n5026_,
    new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_,
    new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_,
    new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_,
    new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_,
    new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_,
    new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_,
    new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_,
    new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_,
    new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_,
    new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_,
    new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_,
    new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_,
    new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_,
    new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5196_,
    new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_,
    new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_,
    new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_,
    new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_,
    new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_,
    new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_,
    new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_,
    new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_,
    new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_,
    new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_,
    new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_,
    new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_,
    new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_,
    new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_,
    new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_,
    new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_,
    new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_,
    new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5368_, new_n5369_, new_n5370_, new_n5371_, new_n5372_,
    new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_, new_n5378_,
    new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_,
    new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_,
    new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_,
    new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_,
    new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_,
    new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_, new_n5414_,
    new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_, new_n5420_,
    new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_,
    new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_,
    new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_,
    new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_,
    new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_,
    new_n5451_, new_n5452_, new_n5454_, new_n5455_, new_n5456_, new_n5457_,
    new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_,
    new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_,
    new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_,
    new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_,
    new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_,
    new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_,
    new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_,
    new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_,
    new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_,
    new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_,
    new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_,
    new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_,
    new_n5530_, new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_,
    new_n5536_, new_n5537_, new_n5538_, new_n5540_, new_n5541_, new_n5542_,
    new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_,
    new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_,
    new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_,
    new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_,
    new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_,
    new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_,
    new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_,
    new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_,
    new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_,
    new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_,
    new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_,
    new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_,
    new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_,
    new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5626_, new_n5627_,
    new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_,
    new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_,
    new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_,
    new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_,
    new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5712_,
    new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_,
    new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_,
    new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_,
    new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_,
    new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_,
    new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_,
    new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_,
    new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_,
    new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_,
    new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_,
    new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_,
    new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_,
    new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_,
    new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_,
    new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_,
    new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_,
    new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_,
    new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_,
    new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_,
    new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_,
    new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_,
    new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_,
    new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5850_, new_n5851_,
    new_n5852_, new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_,
    new_n5858_, new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_,
    new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_,
    new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_,
    new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_,
    new_n5882_, new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_,
    new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_,
    new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_,
    new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_,
    new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_,
    new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_,
    new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_,
    new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_,
    new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_,
    new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_,
    new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_,
    new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_,
    new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_,
    new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_,
    new_n5967_, new_n5968_, new_n5970_, new_n5971_, new_n5972_, new_n5973_,
    new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_, new_n5979_,
    new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_, new_n5985_,
    new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_, new_n5991_,
    new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_, new_n5997_,
    new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_, new_n6003_,
    new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_, new_n6009_,
    new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_, new_n6015_,
    new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_,
    new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_,
    new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_, new_n6033_,
    new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_,
    new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_, new_n6045_,
    new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_,
    new_n6052_, new_n6053_, new_n6054_, new_n6056_, new_n6057_, new_n6058_,
    new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_,
    new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_,
    new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_,
    new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_,
    new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_,
    new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_,
    new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_,
    new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_,
    new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_,
    new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_,
    new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_,
    new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_,
    new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_,
    new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6142_, new_n6143_,
    new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_,
    new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_,
    new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_,
    new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_,
    new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_,
    new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_,
    new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_,
    new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_,
    new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_,
    new_n6198_, new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_,
    new_n6204_, new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_,
    new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_,
    new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_,
    new_n6222_, new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6228_,
    new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_,
    new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_,
    new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_,
    new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_,
    new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_,
    new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_,
    new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_,
    new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_,
    new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_,
    new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_,
    new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_,
    new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_,
    new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_,
    new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_,
    new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_, new_n6319_,
    new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_, new_n6325_,
    new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_, new_n6331_,
    new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_, new_n6337_,
    new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_, new_n6343_,
    new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_,
    new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_,
    new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_,
    new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6400_, new_n6401_, new_n6402_, new_n6403_, new_n6404_,
    new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_, new_n6410_,
    new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_, new_n6416_,
    new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_, new_n6422_,
    new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_, new_n6428_,
    new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_, new_n6434_,
    new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_, new_n6440_,
    new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_, new_n6446_,
    new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_, new_n6452_,
    new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_, new_n6458_,
    new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_, new_n6464_,
    new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_, new_n6470_,
    new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_, new_n6476_,
    new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_, new_n6482_,
    new_n6483_, new_n6484_, new_n6486_, new_n6487_, new_n6488_, new_n6489_,
    new_n6490_, new_n6491_, new_n6492_, new_n6493_, new_n6494_, new_n6495_,
    new_n6496_, new_n6497_, new_n6498_, new_n6499_, new_n6500_, new_n6501_,
    new_n6502_, new_n6503_, new_n6504_, new_n6505_, new_n6506_, new_n6507_,
    new_n6508_, new_n6509_, new_n6510_, new_n6511_, new_n6512_, new_n6513_,
    new_n6514_, new_n6515_, new_n6516_, new_n6517_, new_n6518_, new_n6519_,
    new_n6520_, new_n6521_, new_n6522_, new_n6523_, new_n6524_, new_n6525_,
    new_n6526_, new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_,
    new_n6532_, new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_,
    new_n6538_, new_n6539_, new_n6540_, new_n6541_, new_n6542_, new_n6543_,
    new_n6544_, new_n6545_, new_n6546_, new_n6547_, new_n6548_, new_n6549_,
    new_n6550_, new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n6555_,
    new_n6556_, new_n6557_, new_n6558_, new_n6559_, new_n6560_, new_n6561_,
    new_n6562_, new_n6563_, new_n6564_, new_n6565_, new_n6566_, new_n6567_,
    new_n6568_, new_n6569_, new_n6570_, new_n6572_, new_n6573_, new_n6574_,
    new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_,
    new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_,
    new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_,
    new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_,
    new_n6599_, new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_,
    new_n6605_, new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_,
    new_n6611_, new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_,
    new_n6617_, new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_,
    new_n6623_, new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_,
    new_n6629_, new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_,
    new_n6635_, new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_,
    new_n6641_, new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_,
    new_n6647_, new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_,
    new_n6653_, new_n6654_, new_n6655_, new_n6656_, new_n6658_, new_n6659_,
    new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_,
    new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_,
    new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_,
    new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_,
    new_n6684_, new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_,
    new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_,
    new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_,
    new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_,
    new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_,
    new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_,
    new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_,
    new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6744_,
    new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_,
    new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_,
    new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_,
    new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_,
    new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_,
    new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_,
    new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_,
    new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_,
    new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_,
    new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_,
    new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_,
    new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_,
    new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_,
    new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_,
    new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_,
    new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_,
    new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_,
    new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_,
    new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_,
    new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_,
    new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_,
    new_n6914_, new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6920_,
    new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_,
    new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_,
    new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_,
    new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_,
    new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6950_,
    new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_, new_n6956_,
    new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_, new_n6962_,
    new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_, new_n6968_,
    new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_, new_n6974_,
    new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_, new_n6980_,
    new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_, new_n6986_,
    new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_, new_n6992_,
    new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_, new_n6998_,
    new_n6999_, new_n7000_, new_n7002_, new_n7003_, new_n7004_, new_n7005_,
    new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_, new_n7011_,
    new_n7012_, new_n7013_, new_n7014_, new_n7015_, new_n7016_, new_n7017_,
    new_n7018_, new_n7019_, new_n7020_, new_n7021_, new_n7022_, new_n7023_,
    new_n7024_, new_n7025_, new_n7026_, new_n7027_, new_n7028_, new_n7029_,
    new_n7030_, new_n7031_, new_n7032_, new_n7033_, new_n7034_, new_n7035_,
    new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7040_, new_n7041_,
    new_n7042_, new_n7043_, new_n7044_, new_n7045_, new_n7046_, new_n7047_,
    new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_, new_n7053_,
    new_n7054_, new_n7055_, new_n7056_, new_n7057_, new_n7058_, new_n7059_,
    new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_, new_n7065_,
    new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_, new_n7071_,
    new_n7072_, new_n7073_, new_n7074_, new_n7075_, new_n7076_, new_n7077_,
    new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_,
    new_n7084_, new_n7085_, new_n7086_, new_n7088_, new_n7089_, new_n7090_,
    new_n7091_, new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_,
    new_n7097_, new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_,
    new_n7103_, new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_,
    new_n7109_, new_n7110_, new_n7111_, new_n7112_, new_n7113_, new_n7114_,
    new_n7115_, new_n7116_, new_n7117_, new_n7118_, new_n7119_, new_n7120_,
    new_n7121_, new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_,
    new_n7127_, new_n7128_, new_n7129_, new_n7130_, new_n7131_, new_n7132_,
    new_n7133_, new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_,
    new_n7139_, new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_,
    new_n7145_, new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_,
    new_n7151_, new_n7152_, new_n7153_, new_n7154_, new_n7155_, new_n7156_,
    new_n7157_, new_n7158_, new_n7159_, new_n7160_, new_n7161_, new_n7162_,
    new_n7163_, new_n7164_, new_n7165_, new_n7166_, new_n7167_, new_n7168_,
    new_n7169_, new_n7170_, new_n7171_, new_n7172_, new_n7174_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_,
    new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_,
    new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_,
    new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_,
    new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_,
    new_n7206_, new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_,
    new_n7212_, new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_,
    new_n7218_, new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_,
    new_n7224_, new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_,
    new_n7230_, new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_,
    new_n7236_, new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_,
    new_n7242_, new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_,
    new_n7248_, new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_,
    new_n7254_, new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7260_,
    new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_,
    new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_,
    new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_,
    new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_,
    new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_,
    new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_,
    new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_,
    new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_,
    new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_,
    new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_,
    new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_,
    new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_,
    new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_,
    new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_,
    new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_,
    new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_,
    new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_,
    new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_,
    new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_,
    new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_,
    new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_,
    new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_,
    new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_,
    new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_,
    new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_,
    new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_,
    new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_,
    new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_,
    new_n7430_, new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_,
    new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_,
    new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_,
    new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_,
    new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_,
    new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_,
    new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_,
    new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_,
    new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_,
    new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_,
    new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_,
    new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_,
    new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_,
    new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_,
    new_n7515_, new_n7516_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_,
    new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_,
    new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_,
    new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_,
    new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_,
    new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_,
    new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_,
    new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_,
    new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_,
    new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_,
    new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_,
    new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_,
    new_n7600_, new_n7601_, new_n7602_, new_n7604_, new_n7605_, new_n7606_,
    new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_,
    new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_,
    new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_,
    new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_,
    new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_,
    new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_,
    new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_,
    new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_,
    new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_,
    new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_,
    new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_,
    new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_,
    new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_,
    new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7690_, new_n7691_,
    new_n7692_, new_n7693_, new_n7694_, new_n7695_, new_n7696_, new_n7697_,
    new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_, new_n7703_,
    new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_, new_n7709_,
    new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_, new_n7715_,
    new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_, new_n7721_,
    new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_, new_n7727_,
    new_n7728_, new_n7729_, new_n7730_, new_n7731_, new_n7732_, new_n7733_,
    new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_, new_n7739_,
    new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7744_, new_n7745_,
    new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_,
    new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_, new_n7757_,
    new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_, new_n7763_,
    new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_, new_n7769_,
    new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_, new_n7776_,
    new_n7777_, new_n7778_, new_n7779_, new_n7780_, new_n7781_, new_n7782_,
    new_n7783_, new_n7784_, new_n7785_, new_n7786_, new_n7787_, new_n7788_,
    new_n7789_, new_n7790_, new_n7791_, new_n7792_, new_n7793_, new_n7794_,
    new_n7795_, new_n7796_, new_n7797_, new_n7798_, new_n7799_, new_n7800_,
    new_n7801_, new_n7802_, new_n7803_, new_n7804_, new_n7805_, new_n7806_,
    new_n7807_, new_n7808_, new_n7809_, new_n7810_, new_n7811_, new_n7812_,
    new_n7813_, new_n7814_, new_n7815_, new_n7816_, new_n7817_, new_n7818_,
    new_n7819_, new_n7820_, new_n7821_, new_n7822_, new_n7823_, new_n7824_,
    new_n7825_, new_n7826_, new_n7827_, new_n7828_, new_n7829_, new_n7830_,
    new_n7831_, new_n7832_, new_n7833_, new_n7834_, new_n7835_, new_n7836_,
    new_n7837_, new_n7838_, new_n7839_, new_n7840_, new_n7841_, new_n7842_,
    new_n7843_, new_n7844_, new_n7845_, new_n7846_, new_n7847_, new_n7848_,
    new_n7849_, new_n7850_, new_n7851_, new_n7852_, new_n7853_, new_n7854_,
    new_n7855_, new_n7856_, new_n7857_, new_n7858_, new_n7859_, new_n7860_,
    new_n7862_, new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_,
    new_n7868_, new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_,
    new_n7874_, new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_,
    new_n7880_, new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_,
    new_n7886_, new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_,
    new_n7892_, new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_,
    new_n7898_, new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_,
    new_n7904_, new_n7905_, new_n7906_, new_n7907_, new_n7908_, new_n7909_,
    new_n7910_, new_n7911_, new_n7912_, new_n7913_, new_n7914_, new_n7915_,
    new_n7916_, new_n7917_, new_n7918_, new_n7919_, new_n7920_, new_n7921_,
    new_n7922_, new_n7923_, new_n7924_, new_n7925_, new_n7926_, new_n7927_,
    new_n7928_, new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_,
    new_n7934_, new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_,
    new_n7940_, new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_,
    new_n7946_, new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_,
    new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_,
    new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_,
    new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_,
    new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_,
    new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_,
    new_n7983_, new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_,
    new_n7989_, new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_,
    new_n7995_, new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_,
    new_n8001_, new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_,
    new_n8007_, new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_,
    new_n8013_, new_n8014_, new_n8015_, new_n8016_, new_n8017_, new_n8018_,
    new_n8019_, new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_,
    new_n8025_, new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8030_,
    new_n8031_, new_n8032_, new_n8034_, new_n8035_, new_n8036_, new_n8037_,
    new_n8038_, new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_,
    new_n8044_, new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_,
    new_n8050_, new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_,
    new_n8056_, new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_,
    new_n8062_, new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_,
    new_n8068_, new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_,
    new_n8074_, new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_,
    new_n8080_, new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_,
    new_n8086_, new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_,
    new_n8092_, new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_,
    new_n8098_, new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_,
    new_n8104_, new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_,
    new_n8110_, new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_,
    new_n8116_, new_n8117_, new_n8118_, new_n8120_, new_n8121_, new_n8122_,
    new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_,
    new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_,
    new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_,
    new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_,
    new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_,
    new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_,
    new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_,
    new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_,
    new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_,
    new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_,
    new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_,
    new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_,
    new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_,
    new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8206_, new_n8207_,
    new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_,
    new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8292_,
    new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_,
    new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_,
    new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_,
    new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_,
    new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_,
    new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_, new_n8328_,
    new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_, new_n8334_,
    new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_,
    new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_, new_n8346_,
    new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_, new_n8352_,
    new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_,
    new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_,
    new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_, new_n8370_,
    new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_, new_n8376_,
    new_n8378_, new_n8379_, new_n8380_, new_n8381_, new_n8382_, new_n8383_,
    new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8389_,
    new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_, new_n8395_,
    new_n8396_, new_n8397_, new_n8398_, new_n8399_, new_n8400_, new_n8401_,
    new_n8402_, new_n8403_, new_n8404_, new_n8405_, new_n8406_, new_n8407_,
    new_n8408_, new_n8409_, new_n8410_, new_n8411_, new_n8412_, new_n8413_,
    new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_, new_n8419_,
    new_n8420_, new_n8421_, new_n8422_, new_n8423_, new_n8424_, new_n8425_,
    new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_, new_n8431_,
    new_n8432_, new_n8433_, new_n8434_, new_n8435_, new_n8436_, new_n8437_,
    new_n8438_, new_n8439_, new_n8440_, new_n8441_, new_n8442_, new_n8443_,
    new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8448_, new_n8449_,
    new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_, new_n8455_,
    new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_, new_n8461_,
    new_n8462_, new_n8464_, new_n8465_, new_n8466_, new_n8467_, new_n8468_,
    new_n8469_, new_n8470_, new_n8471_, new_n8472_, new_n8473_, new_n8474_,
    new_n8475_, new_n8476_, new_n8477_, new_n8478_, new_n8479_, new_n8480_,
    new_n8481_, new_n8482_, new_n8483_, new_n8484_, new_n8485_, new_n8486_,
    new_n8487_, new_n8488_, new_n8489_, new_n8490_, new_n8491_, new_n8492_,
    new_n8493_, new_n8494_, new_n8495_, new_n8496_, new_n8497_, new_n8498_,
    new_n8499_, new_n8500_, new_n8501_, new_n8502_, new_n8503_, new_n8504_,
    new_n8505_, new_n8506_, new_n8507_, new_n8508_, new_n8509_, new_n8510_,
    new_n8511_, new_n8512_, new_n8513_, new_n8514_, new_n8515_, new_n8516_,
    new_n8517_, new_n8518_, new_n8519_, new_n8520_, new_n8521_, new_n8522_,
    new_n8523_, new_n8524_, new_n8525_, new_n8526_, new_n8527_, new_n8528_,
    new_n8529_, new_n8530_, new_n8531_, new_n8532_, new_n8533_, new_n8534_,
    new_n8535_, new_n8536_, new_n8537_, new_n8538_, new_n8539_, new_n8540_,
    new_n8541_, new_n8542_, new_n8543_, new_n8544_, new_n8545_, new_n8546_,
    new_n8547_, new_n8548_, new_n8550_, new_n8551_, new_n8552_, new_n8553_,
    new_n8554_, new_n8555_, new_n8556_, new_n8557_, new_n8558_, new_n8559_,
    new_n8560_, new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_,
    new_n8566_, new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_,
    new_n8572_, new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_,
    new_n8578_, new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_,
    new_n8584_, new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_,
    new_n8590_, new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_,
    new_n8596_, new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_,
    new_n8602_, new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_,
    new_n8608_, new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_,
    new_n8614_, new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_,
    new_n8620_, new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_,
    new_n8626_, new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_,
    new_n8632_, new_n8633_, new_n8634_, new_n8636_, new_n8637_, new_n8638_,
    new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_,
    new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_,
    new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_,
    new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_,
    new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_,
    new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_,
    new_n8675_, new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_,
    new_n8681_, new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_,
    new_n8687_, new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_,
    new_n8693_, new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_,
    new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_,
    new_n8705_, new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_,
    new_n8711_, new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_,
    new_n8717_, new_n8718_, new_n8719_, new_n8720_, new_n8722_, new_n8723_,
    new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_,
    new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_,
    new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_,
    new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_,
    new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_,
    new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_,
    new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_,
    new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_,
    new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_,
    new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_,
    new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_,
    new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_,
    new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_,
    new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8808_,
    new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_,
    new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_,
    new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_,
    new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_,
    new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_,
    new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_,
    new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_,
    new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_,
    new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_,
    new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_,
    new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_,
    new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_,
    new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_,
    new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_,
    new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_, new_n8899_,
    new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_,
    new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8980_, new_n8981_, new_n8982_, new_n8983_, new_n8984_,
    new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_, new_n8990_,
    new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_, new_n8996_,
    new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_, new_n9002_,
    new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_, new_n9008_,
    new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_, new_n9014_,
    new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_, new_n9020_,
    new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_, new_n9026_,
    new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_, new_n9032_,
    new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_, new_n9038_,
    new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_, new_n9044_,
    new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_, new_n9050_,
    new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_, new_n9056_,
    new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_,
    new_n9063_, new_n9064_, new_n9066_, new_n9067_, new_n9068_, new_n9069_,
    new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_, new_n9075_,
    new_n9076_, new_n9077_, new_n9078_, new_n9079_, new_n9080_, new_n9081_,
    new_n9082_, new_n9083_, new_n9084_, new_n9085_, new_n9086_, new_n9087_,
    new_n9088_, new_n9089_, new_n9090_, new_n9091_, new_n9092_, new_n9093_,
    new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_, new_n9099_,
    new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_, new_n9105_,
    new_n9106_, new_n9107_, new_n9108_, new_n9109_, new_n9110_, new_n9111_,
    new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_, new_n9117_,
    new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_, new_n9123_,
    new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_, new_n9129_,
    new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_, new_n9135_,
    new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_, new_n9141_,
    new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9147_,
    new_n9148_, new_n9149_, new_n9150_, new_n9152_, new_n9153_, new_n9154_,
    new_n9155_, new_n9156_, new_n9157_, new_n9158_, new_n9159_, new_n9160_,
    new_n9161_, new_n9162_, new_n9163_, new_n9164_, new_n9165_, new_n9166_,
    new_n9167_, new_n9168_, new_n9169_, new_n9170_, new_n9171_, new_n9172_,
    new_n9173_, new_n9174_, new_n9175_, new_n9176_, new_n9177_, new_n9178_,
    new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_, new_n9184_,
    new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_, new_n9190_,
    new_n9191_, new_n9192_, new_n9193_, new_n9194_, new_n9195_, new_n9196_,
    new_n9197_, new_n9198_, new_n9199_, new_n9200_, new_n9201_, new_n9202_,
    new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_, new_n9208_,
    new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_, new_n9214_,
    new_n9215_, new_n9216_, new_n9217_, new_n9218_, new_n9219_, new_n9220_,
    new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_, new_n9226_,
    new_n9227_, new_n9228_, new_n9229_, new_n9230_, new_n9231_, new_n9232_,
    new_n9233_, new_n9234_, new_n9235_, new_n9236_, new_n9238_, new_n9239_,
    new_n9240_, new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_,
    new_n9246_, new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_,
    new_n9252_, new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_,
    new_n9258_, new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_,
    new_n9264_, new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_,
    new_n9270_, new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_,
    new_n9276_, new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_,
    new_n9282_, new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_,
    new_n9288_, new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_,
    new_n9294_, new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_,
    new_n9300_, new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_,
    new_n9306_, new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_,
    new_n9312_, new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_,
    new_n9318_, new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9324_,
    new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_,
    new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_,
    new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_,
    new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_,
    new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_,
    new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_,
    new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_,
    new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_,
    new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_,
    new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_,
    new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_,
    new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_,
    new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_,
    new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_,
    new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_, new_n9415_,
    new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_, new_n9421_,
    new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_, new_n9427_,
    new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_, new_n9433_,
    new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_, new_n9439_,
    new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_, new_n9445_,
    new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_, new_n9451_,
    new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_, new_n9457_,
    new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_, new_n9463_,
    new_n9464_, new_n9465_, new_n9466_, new_n9467_, new_n9468_, new_n9469_,
    new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_, new_n9475_,
    new_n9476_, new_n9477_, new_n9478_, new_n9479_, new_n9480_, new_n9481_,
    new_n9482_, new_n9483_, new_n9484_, new_n9485_, new_n9486_, new_n9487_,
    new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_, new_n9493_,
    new_n9494_, new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_,
    new_n9501_, new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_,
    new_n9507_, new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_,
    new_n9513_, new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_,
    new_n9519_, new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_,
    new_n9525_, new_n9526_, new_n9527_, new_n9528_, new_n9529_, new_n9530_,
    new_n9531_, new_n9532_, new_n9533_, new_n9534_, new_n9535_, new_n9536_,
    new_n9537_, new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9542_,
    new_n9543_, new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_,
    new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_,
    new_n9555_, new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_,
    new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_,
    new_n9567_, new_n9568_, new_n9569_, new_n9570_, new_n9571_, new_n9572_,
    new_n9573_, new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_,
    new_n9579_, new_n9580_, new_n9582_, new_n9583_, new_n9584_, new_n9585_,
    new_n9586_, new_n9587_, new_n9588_, new_n9589_, new_n9590_, new_n9591_,
    new_n9592_, new_n9593_, new_n9594_, new_n9595_, new_n9596_, new_n9597_,
    new_n9598_, new_n9599_, new_n9600_, new_n9601_, new_n9602_, new_n9603_,
    new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_, new_n9609_,
    new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_, new_n9615_,
    new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9621_,
    new_n9622_, new_n9623_, new_n9624_, new_n9625_, new_n9626_, new_n9627_,
    new_n9628_, new_n9629_, new_n9630_, new_n9631_, new_n9632_, new_n9633_,
    new_n9634_, new_n9635_, new_n9636_, new_n9637_, new_n9638_, new_n9639_,
    new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_,
    new_n9646_, new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_,
    new_n9652_, new_n9653_, new_n9654_, new_n9655_, new_n9656_, new_n9657_,
    new_n9658_, new_n9659_, new_n9660_, new_n9661_, new_n9662_, new_n9663_,
    new_n9664_, new_n9665_, new_n9666_, new_n9668_, new_n9669_, new_n9670_,
    new_n9671_, new_n9672_, new_n9673_, new_n9674_, new_n9675_, new_n9676_,
    new_n9677_, new_n9678_, new_n9679_, new_n9680_, new_n9681_, new_n9682_,
    new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_, new_n9688_,
    new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_, new_n9694_,
    new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_, new_n9700_,
    new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_, new_n9706_,
    new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_, new_n9712_,
    new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_, new_n9718_,
    new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_, new_n9724_,
    new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_, new_n9730_,
    new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_, new_n9736_,
    new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_, new_n9742_,
    new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_, new_n9748_,
    new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9754_, new_n9755_,
    new_n9756_, new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_,
    new_n9762_, new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_,
    new_n9768_, new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9773_,
    new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9778_, new_n9779_,
    new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9784_, new_n9785_,
    new_n9786_, new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_,
    new_n9792_, new_n9793_, new_n9794_, new_n9795_, new_n9796_, new_n9797_,
    new_n9798_, new_n9799_, new_n9800_, new_n9801_, new_n9802_, new_n9803_,
    new_n9804_, new_n9805_, new_n9806_, new_n9807_, new_n9808_, new_n9809_,
    new_n9810_, new_n9811_, new_n9812_, new_n9813_, new_n9814_, new_n9815_,
    new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_, new_n9821_,
    new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_, new_n9827_,
    new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_, new_n9833_,
    new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_, new_n9840_,
    new_n9841_, new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_,
    new_n9847_, new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_,
    new_n9853_, new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_,
    new_n9859_, new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_,
    new_n9865_, new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_,
    new_n9871_, new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_,
    new_n9877_, new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_,
    new_n9883_, new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_,
    new_n9889_, new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_,
    new_n9895_, new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_,
    new_n9901_, new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_,
    new_n9907_, new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_,
    new_n9913_, new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_,
    new_n9919_, new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_,
    new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_,
    new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9949_,
    new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_, new_n9955_,
    new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_, new_n9961_,
    new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_, new_n9967_,
    new_n9968_, new_n9969_, new_n9970_, new_n9971_, new_n9972_, new_n9973_,
    new_n9974_, new_n9975_, new_n9976_, new_n9977_, new_n9978_, new_n9979_,
    new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9984_, new_n9985_,
    new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_, new_n9991_,
    new_n9992_, new_n9993_, new_n9994_, new_n9995_, new_n9996_, new_n9997_,
    new_n9998_, new_n9999_, new_n10000_, new_n10001_, new_n10002_,
    new_n10003_, new_n10004_, new_n10005_, new_n10006_, new_n10007_,
    new_n10008_, new_n10009_, new_n10010_, new_n10012_, new_n10013_,
    new_n10014_, new_n10015_, new_n10016_, new_n10017_, new_n10018_,
    new_n10019_, new_n10020_, new_n10021_, new_n10022_, new_n10023_,
    new_n10024_, new_n10025_, new_n10026_, new_n10027_, new_n10028_,
    new_n10029_, new_n10030_, new_n10031_, new_n10032_, new_n10033_,
    new_n10034_, new_n10035_, new_n10036_, new_n10037_, new_n10038_,
    new_n10039_, new_n10040_, new_n10041_, new_n10042_, new_n10043_,
    new_n10044_, new_n10045_, new_n10046_, new_n10047_, new_n10048_,
    new_n10049_, new_n10050_, new_n10051_, new_n10052_, new_n10053_,
    new_n10054_, new_n10055_, new_n10056_, new_n10057_, new_n10058_,
    new_n10059_, new_n10060_, new_n10061_, new_n10062_, new_n10063_,
    new_n10064_, new_n10065_, new_n10066_, new_n10067_, new_n10068_,
    new_n10069_, new_n10070_, new_n10071_, new_n10072_, new_n10073_,
    new_n10074_, new_n10075_, new_n10076_, new_n10077_, new_n10078_,
    new_n10079_, new_n10080_, new_n10081_, new_n10082_, new_n10083_,
    new_n10084_, new_n10085_, new_n10086_, new_n10087_, new_n10088_,
    new_n10089_, new_n10090_, new_n10091_, new_n10092_, new_n10093_,
    new_n10094_, new_n10095_, new_n10096_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10191_, new_n10192_, new_n10193_, new_n10194_, new_n10195_,
    new_n10196_, new_n10197_, new_n10198_, new_n10199_, new_n10200_,
    new_n10201_, new_n10202_, new_n10203_, new_n10204_, new_n10205_,
    new_n10206_, new_n10207_, new_n10208_, new_n10209_, new_n10210_,
    new_n10211_, new_n10212_, new_n10213_, new_n10214_, new_n10215_,
    new_n10216_, new_n10217_, new_n10218_, new_n10219_, new_n10220_,
    new_n10221_, new_n10222_, new_n10223_, new_n10224_, new_n10225_,
    new_n10226_, new_n10227_, new_n10228_, new_n10229_, new_n10230_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10241_, new_n10242_, new_n10243_, new_n10244_, new_n10245_,
    new_n10246_, new_n10247_, new_n10248_, new_n10249_, new_n10250_,
    new_n10251_, new_n10252_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10257_, new_n10258_, new_n10259_, new_n10260_,
    new_n10261_, new_n10262_, new_n10263_, new_n10264_, new_n10265_,
    new_n10266_, new_n10267_, new_n10268_, new_n10270_, new_n10271_,
    new_n10272_, new_n10273_, new_n10274_, new_n10275_, new_n10276_,
    new_n10277_, new_n10278_, new_n10279_, new_n10280_, new_n10281_,
    new_n10282_, new_n10283_, new_n10284_, new_n10285_, new_n10286_,
    new_n10287_, new_n10288_, new_n10289_, new_n10290_, new_n10291_,
    new_n10292_, new_n10293_, new_n10294_, new_n10295_, new_n10296_,
    new_n10297_, new_n10298_, new_n10299_, new_n10300_, new_n10301_,
    new_n10302_, new_n10303_, new_n10304_, new_n10305_, new_n10306_,
    new_n10307_, new_n10308_, new_n10309_, new_n10310_, new_n10311_,
    new_n10312_, new_n10313_, new_n10314_, new_n10315_, new_n10316_,
    new_n10317_, new_n10318_, new_n10319_, new_n10320_, new_n10321_,
    new_n10322_, new_n10323_, new_n10324_, new_n10325_, new_n10326_,
    new_n10327_, new_n10328_, new_n10329_, new_n10330_, new_n10331_,
    new_n10332_, new_n10333_, new_n10334_, new_n10335_, new_n10336_,
    new_n10337_, new_n10338_, new_n10339_, new_n10340_, new_n10341_,
    new_n10342_, new_n10343_, new_n10344_, new_n10345_, new_n10346_,
    new_n10347_, new_n10348_, new_n10349_, new_n10350_, new_n10351_,
    new_n10352_, new_n10353_, new_n10354_, new_n10356_, new_n10357_,
    new_n10358_, new_n10359_, new_n10360_, new_n10361_, new_n10362_,
    new_n10363_, new_n10364_, new_n10365_, new_n10366_, new_n10367_,
    new_n10368_, new_n10369_, new_n10370_, new_n10371_, new_n10372_,
    new_n10373_, new_n10374_, new_n10375_, new_n10376_, new_n10377_,
    new_n10378_, new_n10379_, new_n10380_, new_n10381_, new_n10382_,
    new_n10383_, new_n10384_, new_n10385_, new_n10386_, new_n10387_,
    new_n10388_, new_n10389_, new_n10390_, new_n10391_, new_n10392_,
    new_n10393_, new_n10394_, new_n10395_, new_n10396_, new_n10397_,
    new_n10398_, new_n10399_, new_n10400_, new_n10401_, new_n10402_,
    new_n10403_, new_n10404_, new_n10405_, new_n10406_, new_n10407_,
    new_n10408_, new_n10409_, new_n10410_, new_n10411_, new_n10412_,
    new_n10413_, new_n10414_, new_n10415_, new_n10416_, new_n10417_,
    new_n10418_, new_n10419_, new_n10420_, new_n10421_, new_n10422_,
    new_n10423_, new_n10424_, new_n10425_, new_n10426_, new_n10427_,
    new_n10428_, new_n10429_, new_n10430_, new_n10431_, new_n10432_,
    new_n10433_, new_n10434_, new_n10435_, new_n10436_, new_n10437_,
    new_n10438_, new_n10439_, new_n10440_, new_n10442_, new_n10443_,
    new_n10444_, new_n10445_, new_n10446_, new_n10447_, new_n10448_,
    new_n10449_, new_n10450_, new_n10451_, new_n10452_, new_n10453_,
    new_n10454_, new_n10455_, new_n10456_, new_n10457_, new_n10458_,
    new_n10459_, new_n10460_, new_n10461_, new_n10462_, new_n10463_,
    new_n10464_, new_n10465_, new_n10466_, new_n10467_, new_n10468_,
    new_n10469_, new_n10470_, new_n10471_, new_n10472_, new_n10473_,
    new_n10474_, new_n10475_, new_n10476_, new_n10477_, new_n10478_,
    new_n10479_, new_n10480_, new_n10481_, new_n10482_, new_n10483_,
    new_n10484_, new_n10485_, new_n10486_, new_n10487_, new_n10488_,
    new_n10489_, new_n10490_, new_n10491_, new_n10492_, new_n10493_,
    new_n10494_, new_n10495_, new_n10496_, new_n10497_, new_n10498_,
    new_n10499_, new_n10500_, new_n10501_, new_n10502_, new_n10503_,
    new_n10504_, new_n10505_, new_n10506_, new_n10507_, new_n10508_,
    new_n10509_, new_n10510_, new_n10511_, new_n10512_, new_n10513_,
    new_n10514_, new_n10515_, new_n10516_, new_n10517_, new_n10518_,
    new_n10519_, new_n10520_, new_n10521_, new_n10522_, new_n10523_,
    new_n10524_, new_n10525_, new_n10526_, new_n10528_, new_n10529_,
    new_n10530_, new_n10531_, new_n10532_, new_n10533_, new_n10534_,
    new_n10535_, new_n10536_, new_n10537_, new_n10538_, new_n10539_,
    new_n10540_, new_n10541_, new_n10542_, new_n10543_, new_n10544_,
    new_n10545_, new_n10546_, new_n10547_, new_n10548_, new_n10549_,
    new_n10550_, new_n10551_, new_n10552_, new_n10553_, new_n10554_,
    new_n10555_, new_n10556_, new_n10557_, new_n10558_, new_n10559_,
    new_n10560_, new_n10561_, new_n10562_, new_n10563_, new_n10564_,
    new_n10565_, new_n10566_, new_n10567_, new_n10568_, new_n10569_,
    new_n10570_, new_n10571_, new_n10572_, new_n10573_, new_n10574_,
    new_n10575_, new_n10576_, new_n10577_, new_n10578_, new_n10579_,
    new_n10580_, new_n10581_, new_n10582_, new_n10583_, new_n10584_,
    new_n10585_, new_n10586_, new_n10587_, new_n10588_, new_n10589_,
    new_n10590_, new_n10591_, new_n10592_, new_n10593_, new_n10594_,
    new_n10595_, new_n10596_, new_n10597_, new_n10598_, new_n10599_,
    new_n10600_, new_n10601_, new_n10602_, new_n10603_, new_n10604_,
    new_n10605_, new_n10606_, new_n10607_, new_n10608_, new_n10609_,
    new_n10610_, new_n10611_, new_n10612_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10700_, new_n10701_,
    new_n10702_, new_n10703_, new_n10704_, new_n10705_, new_n10706_,
    new_n10707_, new_n10708_, new_n10709_, new_n10710_, new_n10711_,
    new_n10712_, new_n10713_, new_n10714_, new_n10715_, new_n10716_,
    new_n10717_, new_n10718_, new_n10719_, new_n10720_, new_n10721_,
    new_n10722_, new_n10723_, new_n10724_, new_n10725_, new_n10726_,
    new_n10727_, new_n10728_, new_n10729_, new_n10730_, new_n10731_,
    new_n10732_, new_n10733_, new_n10734_, new_n10735_, new_n10736_,
    new_n10737_, new_n10738_, new_n10739_, new_n10740_, new_n10741_,
    new_n10742_, new_n10743_, new_n10744_, new_n10745_, new_n10746_,
    new_n10747_, new_n10748_, new_n10749_, new_n10750_, new_n10751_,
    new_n10752_, new_n10753_, new_n10754_, new_n10755_, new_n10756_,
    new_n10757_, new_n10758_, new_n10759_, new_n10760_, new_n10761_,
    new_n10762_, new_n10763_, new_n10764_, new_n10765_, new_n10766_,
    new_n10767_, new_n10768_, new_n10769_, new_n10770_, new_n10771_,
    new_n10772_, new_n10773_, new_n10774_, new_n10775_, new_n10776_,
    new_n10777_, new_n10778_, new_n10779_, new_n10780_, new_n10781_,
    new_n10782_, new_n10783_, new_n10784_, new_n10786_, new_n10787_,
    new_n10788_, new_n10789_, new_n10790_, new_n10791_, new_n10792_,
    new_n10793_, new_n10794_, new_n10795_, new_n10796_, new_n10797_,
    new_n10798_, new_n10799_, new_n10800_, new_n10801_, new_n10802_,
    new_n10803_, new_n10804_, new_n10805_, new_n10806_, new_n10807_,
    new_n10808_, new_n10809_, new_n10810_, new_n10811_, new_n10812_,
    new_n10813_, new_n10814_, new_n10815_, new_n10816_, new_n10817_,
    new_n10818_, new_n10819_, new_n10820_, new_n10821_, new_n10822_,
    new_n10823_, new_n10824_, new_n10825_, new_n10826_, new_n10827_,
    new_n10828_, new_n10829_, new_n10830_, new_n10831_, new_n10832_,
    new_n10833_, new_n10834_, new_n10835_, new_n10836_, new_n10837_,
    new_n10838_, new_n10839_, new_n10840_, new_n10841_, new_n10842_,
    new_n10843_, new_n10844_, new_n10845_, new_n10846_, new_n10847_,
    new_n10848_, new_n10849_, new_n10850_, new_n10851_, new_n10852_,
    new_n10853_, new_n10854_, new_n10855_, new_n10856_, new_n10857_,
    new_n10858_, new_n10859_, new_n10860_, new_n10861_, new_n10862_,
    new_n10863_, new_n10864_, new_n10865_, new_n10866_, new_n10867_,
    new_n10868_, new_n10869_, new_n10870_, new_n10872_, new_n10873_,
    new_n10874_, new_n10875_, new_n10876_, new_n10877_, new_n10878_,
    new_n10879_, new_n10880_, new_n10881_, new_n10882_, new_n10883_,
    new_n10884_, new_n10885_, new_n10886_, new_n10887_, new_n10888_,
    new_n10889_, new_n10890_, new_n10891_, new_n10892_, new_n10893_,
    new_n10894_, new_n10895_, new_n10896_, new_n10897_, new_n10898_,
    new_n10899_, new_n10900_, new_n10901_, new_n10902_, new_n10903_,
    new_n10904_, new_n10905_, new_n10906_, new_n10907_, new_n10908_,
    new_n10909_, new_n10910_, new_n10911_, new_n10912_, new_n10913_,
    new_n10914_, new_n10915_, new_n10916_, new_n10917_, new_n10918_,
    new_n10919_, new_n10920_, new_n10921_, new_n10922_, new_n10923_,
    new_n10924_, new_n10925_, new_n10926_, new_n10927_, new_n10928_,
    new_n10929_, new_n10930_, new_n10931_, new_n10932_, new_n10933_,
    new_n10934_, new_n10935_, new_n10936_, new_n10937_, new_n10938_,
    new_n10939_, new_n10940_, new_n10941_, new_n10942_, new_n10943_,
    new_n10944_, new_n10945_, new_n10946_, new_n10947_, new_n10948_,
    new_n10949_, new_n10950_, new_n10951_, new_n10952_, new_n10953_,
    new_n10954_, new_n10955_, new_n10956_, new_n10958_, new_n10959_,
    new_n10960_, new_n10961_, new_n10962_, new_n10963_, new_n10964_,
    new_n10965_, new_n10966_, new_n10967_, new_n10968_, new_n10969_,
    new_n10970_, new_n10971_, new_n10972_, new_n10973_, new_n10974_,
    new_n10975_, new_n10976_, new_n10977_, new_n10978_, new_n10979_,
    new_n10980_, new_n10981_, new_n10982_, new_n10983_, new_n10984_,
    new_n10985_, new_n10986_, new_n10987_, new_n10988_, new_n10989_,
    new_n10990_, new_n10991_, new_n10992_, new_n10993_, new_n10994_,
    new_n10995_, new_n10996_, new_n10997_, new_n10998_, new_n10999_,
    new_n11000_, new_n11001_, new_n11002_, new_n11003_, new_n11004_,
    new_n11005_, new_n11006_, new_n11007_, new_n11008_, new_n11009_,
    new_n11010_, new_n11011_, new_n11012_, new_n11013_, new_n11014_,
    new_n11015_, new_n11016_, new_n11017_, new_n11018_, new_n11019_,
    new_n11020_, new_n11021_, new_n11022_, new_n11023_, new_n11024_,
    new_n11025_, new_n11026_, new_n11027_, new_n11028_, new_n11029_,
    new_n11030_, new_n11031_, new_n11032_, new_n11033_, new_n11034_,
    new_n11035_, new_n11036_, new_n11037_, new_n11038_, new_n11039_,
    new_n11040_, new_n11041_, new_n11042_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11072_, new_n11073_, new_n11074_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11094_, new_n11095_,
    new_n11096_, new_n11097_, new_n11098_, new_n11099_, new_n11100_,
    new_n11101_, new_n11102_, new_n11103_, new_n11104_, new_n11105_,
    new_n11106_, new_n11107_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11113_, new_n11114_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11130_, new_n11131_,
    new_n11132_, new_n11133_, new_n11134_, new_n11135_, new_n11136_,
    new_n11137_, new_n11138_, new_n11139_, new_n11140_, new_n11141_,
    new_n11142_, new_n11143_, new_n11144_, new_n11145_, new_n11146_,
    new_n11147_, new_n11148_, new_n11149_, new_n11150_, new_n11151_,
    new_n11152_, new_n11153_, new_n11154_, new_n11155_, new_n11156_,
    new_n11157_, new_n11158_, new_n11159_, new_n11160_, new_n11161_,
    new_n11162_, new_n11163_, new_n11164_, new_n11165_, new_n11166_,
    new_n11167_, new_n11168_, new_n11169_, new_n11170_, new_n11171_,
    new_n11172_, new_n11173_, new_n11174_, new_n11175_, new_n11176_,
    new_n11177_, new_n11178_, new_n11179_, new_n11180_, new_n11181_,
    new_n11182_, new_n11183_, new_n11184_, new_n11185_, new_n11186_,
    new_n11187_, new_n11188_, new_n11189_, new_n11190_, new_n11191_,
    new_n11192_, new_n11193_, new_n11194_, new_n11195_, new_n11196_,
    new_n11197_, new_n11198_, new_n11199_, new_n11200_, new_n11201_,
    new_n11202_, new_n11203_, new_n11204_, new_n11205_, new_n11206_,
    new_n11207_, new_n11208_, new_n11209_, new_n11210_, new_n11211_,
    new_n11212_, new_n11213_, new_n11214_, new_n11216_, new_n11217_,
    new_n11218_, new_n11219_, new_n11220_, new_n11221_, new_n11222_,
    new_n11223_, new_n11224_, new_n11225_, new_n11226_, new_n11227_,
    new_n11228_, new_n11229_, new_n11230_, new_n11231_, new_n11232_,
    new_n11233_, new_n11234_, new_n11235_, new_n11236_, new_n11237_,
    new_n11238_, new_n11239_, new_n11240_, new_n11241_, new_n11242_,
    new_n11243_, new_n11244_, new_n11245_, new_n11246_, new_n11247_,
    new_n11248_, new_n11249_, new_n11250_, new_n11251_, new_n11252_,
    new_n11253_, new_n11254_, new_n11255_, new_n11256_, new_n11257_,
    new_n11258_, new_n11259_, new_n11260_, new_n11261_, new_n11262_,
    new_n11263_, new_n11264_, new_n11265_, new_n11266_, new_n11267_,
    new_n11268_, new_n11269_, new_n11270_, new_n11271_, new_n11272_,
    new_n11273_, new_n11274_, new_n11275_, new_n11276_, new_n11277_,
    new_n11278_, new_n11279_, new_n11280_, new_n11281_, new_n11282_,
    new_n11283_, new_n11284_, new_n11285_, new_n11286_, new_n11287_,
    new_n11288_, new_n11289_, new_n11290_, new_n11291_, new_n11292_,
    new_n11293_, new_n11294_, new_n11295_, new_n11296_, new_n11297_,
    new_n11298_, new_n11299_, new_n11300_, new_n11302_, new_n11303_,
    new_n11304_, new_n11305_, new_n11306_, new_n11307_, new_n11308_,
    new_n11309_, new_n11310_, new_n11311_, new_n11312_, new_n11313_,
    new_n11314_, new_n11315_, new_n11316_, new_n11317_, new_n11318_,
    new_n11319_, new_n11320_, new_n11321_, new_n11322_, new_n11323_,
    new_n11324_, new_n11325_, new_n11326_, new_n11327_, new_n11328_,
    new_n11329_, new_n11330_, new_n11331_, new_n11332_, new_n11333_,
    new_n11334_, new_n11335_, new_n11336_, new_n11337_, new_n11338_,
    new_n11339_, new_n11340_, new_n11341_, new_n11342_, new_n11343_,
    new_n11344_, new_n11345_, new_n11346_, new_n11347_, new_n11348_,
    new_n11349_, new_n11350_, new_n11351_, new_n11352_, new_n11353_,
    new_n11354_, new_n11355_, new_n11356_, new_n11357_, new_n11358_,
    new_n11359_, new_n11360_, new_n11361_, new_n11362_, new_n11363_,
    new_n11364_, new_n11365_, new_n11366_, new_n11367_, new_n11368_,
    new_n11369_, new_n11370_, new_n11371_, new_n11372_, new_n11373_,
    new_n11374_, new_n11375_, new_n11376_, new_n11377_, new_n11378_,
    new_n11379_, new_n11380_, new_n11381_, new_n11382_, new_n11383_,
    new_n11384_, new_n11385_, new_n11386_, new_n11388_, new_n11389_,
    new_n11390_, new_n11391_, new_n11392_, new_n11393_, new_n11394_,
    new_n11395_, new_n11396_, new_n11397_, new_n11398_, new_n11399_,
    new_n11400_, new_n11401_, new_n11402_, new_n11403_, new_n11404_,
    new_n11405_, new_n11406_, new_n11407_, new_n11408_, new_n11409_,
    new_n11410_, new_n11411_, new_n11412_, new_n11413_, new_n11414_,
    new_n11415_, new_n11416_, new_n11417_, new_n11418_, new_n11419_,
    new_n11420_, new_n11421_, new_n11422_, new_n11423_, new_n11424_,
    new_n11425_, new_n11426_, new_n11427_, new_n11428_, new_n11429_,
    new_n11430_, new_n11431_, new_n11432_, new_n11433_, new_n11434_,
    new_n11435_, new_n11436_, new_n11437_, new_n11438_, new_n11439_,
    new_n11440_, new_n11441_, new_n11442_, new_n11443_, new_n11444_,
    new_n11445_, new_n11446_, new_n11447_, new_n11448_, new_n11449_,
    new_n11450_, new_n11451_, new_n11452_, new_n11453_, new_n11454_,
    new_n11455_, new_n11456_, new_n11457_, new_n11458_, new_n11459_,
    new_n11460_, new_n11461_, new_n11462_, new_n11463_, new_n11464_,
    new_n11465_, new_n11466_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11472_, new_n11474_, new_n11475_,
    new_n11476_, new_n11477_, new_n11478_, new_n11479_, new_n11480_,
    new_n11481_, new_n11482_, new_n11483_, new_n11484_, new_n11485_,
    new_n11486_, new_n11487_, new_n11488_, new_n11489_, new_n11490_,
    new_n11491_, new_n11492_, new_n11493_, new_n11494_, new_n11495_,
    new_n11496_, new_n11497_, new_n11498_, new_n11499_, new_n11500_,
    new_n11501_, new_n11502_, new_n11503_, new_n11504_, new_n11505_,
    new_n11506_, new_n11507_, new_n11508_, new_n11509_, new_n11510_,
    new_n11511_, new_n11512_, new_n11513_, new_n11514_, new_n11515_,
    new_n11516_, new_n11517_, new_n11518_, new_n11519_, new_n11520_,
    new_n11521_, new_n11522_, new_n11523_, new_n11524_, new_n11525_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11560_, new_n11561_,
    new_n11562_, new_n11563_, new_n11564_, new_n11565_, new_n11566_,
    new_n11567_, new_n11568_, new_n11569_, new_n11570_, new_n11571_,
    new_n11572_, new_n11573_, new_n11574_, new_n11575_, new_n11576_,
    new_n11577_, new_n11578_, new_n11579_, new_n11580_, new_n11581_,
    new_n11582_, new_n11583_, new_n11584_, new_n11585_, new_n11586_,
    new_n11587_, new_n11588_, new_n11589_, new_n11590_, new_n11591_,
    new_n11592_, new_n11593_, new_n11594_, new_n11595_, new_n11596_,
    new_n11597_, new_n11598_, new_n11599_, new_n11600_, new_n11601_,
    new_n11602_, new_n11603_, new_n11604_, new_n11605_, new_n11606_,
    new_n11607_, new_n11608_, new_n11609_, new_n11610_, new_n11611_,
    new_n11612_, new_n11613_, new_n11614_, new_n11615_, new_n11616_,
    new_n11617_, new_n11618_, new_n11619_, new_n11620_, new_n11621_,
    new_n11622_, new_n11623_, new_n11624_, new_n11625_, new_n11626_,
    new_n11627_, new_n11628_, new_n11629_, new_n11630_, new_n11631_,
    new_n11632_, new_n11633_, new_n11634_, new_n11635_, new_n11636_,
    new_n11637_, new_n11638_, new_n11639_, new_n11640_, new_n11641_,
    new_n11642_, new_n11643_, new_n11644_, new_n11646_, new_n11647_,
    new_n11648_, new_n11649_, new_n11650_, new_n11651_, new_n11652_,
    new_n11653_, new_n11654_, new_n11655_, new_n11656_, new_n11657_,
    new_n11658_, new_n11659_, new_n11660_, new_n11661_, new_n11662_,
    new_n11663_, new_n11664_, new_n11665_, new_n11666_, new_n11667_,
    new_n11668_, new_n11669_, new_n11670_, new_n11671_, new_n11672_,
    new_n11673_, new_n11674_, new_n11675_, new_n11676_, new_n11677_,
    new_n11678_, new_n11679_, new_n11680_, new_n11681_, new_n11682_,
    new_n11683_, new_n11684_, new_n11685_, new_n11686_, new_n11687_,
    new_n11688_, new_n11689_, new_n11690_, new_n11691_, new_n11692_,
    new_n11693_, new_n11694_, new_n11695_, new_n11696_, new_n11697_,
    new_n11698_, new_n11699_, new_n11700_, new_n11701_, new_n11702_,
    new_n11703_, new_n11704_, new_n11705_, new_n11706_, new_n11707_,
    new_n11708_, new_n11709_, new_n11710_, new_n11711_, new_n11712_,
    new_n11713_, new_n11714_, new_n11715_, new_n11716_, new_n11717_,
    new_n11718_, new_n11719_, new_n11720_, new_n11721_, new_n11722_,
    new_n11723_, new_n11724_, new_n11725_, new_n11726_, new_n11727_,
    new_n11728_, new_n11729_, new_n11730_, new_n11732_, new_n11733_,
    new_n11734_, new_n11735_, new_n11736_, new_n11737_, new_n11738_,
    new_n11739_, new_n11740_, new_n11741_, new_n11742_, new_n11743_,
    new_n11744_, new_n11745_, new_n11746_, new_n11747_, new_n11748_,
    new_n11749_, new_n11750_, new_n11751_, new_n11752_, new_n11753_,
    new_n11754_, new_n11755_, new_n11756_, new_n11757_, new_n11758_,
    new_n11759_, new_n11760_, new_n11761_, new_n11762_, new_n11763_,
    new_n11764_, new_n11765_, new_n11766_, new_n11767_, new_n11768_,
    new_n11769_, new_n11770_, new_n11771_, new_n11772_, new_n11773_,
    new_n11774_, new_n11775_, new_n11776_, new_n11777_, new_n11778_,
    new_n11779_, new_n11780_, new_n11781_, new_n11782_, new_n11783_,
    new_n11784_, new_n11785_, new_n11786_, new_n11787_, new_n11788_,
    new_n11789_, new_n11790_, new_n11791_, new_n11792_, new_n11793_,
    new_n11794_, new_n11795_, new_n11796_, new_n11797_, new_n11798_,
    new_n11799_, new_n11800_, new_n11801_, new_n11802_, new_n11803_,
    new_n11804_, new_n11805_, new_n11806_, new_n11807_, new_n11808_,
    new_n11809_, new_n11810_, new_n11811_, new_n11812_, new_n11813_,
    new_n11814_, new_n11815_, new_n11816_, new_n11818_, new_n11819_,
    new_n11820_, new_n11821_, new_n11822_, new_n11823_, new_n11824_,
    new_n11825_, new_n11826_, new_n11827_, new_n11828_, new_n11829_,
    new_n11830_, new_n11831_, new_n11832_, new_n11833_, new_n11834_,
    new_n11835_, new_n11836_, new_n11837_, new_n11838_, new_n11839_,
    new_n11840_, new_n11841_, new_n11842_, new_n11843_, new_n11844_,
    new_n11845_, new_n11846_, new_n11847_, new_n11848_, new_n11849_,
    new_n11850_, new_n11851_, new_n11852_, new_n11853_, new_n11854_,
    new_n11855_, new_n11856_, new_n11857_, new_n11858_, new_n11859_,
    new_n11860_, new_n11861_, new_n11862_, new_n11863_, new_n11864_,
    new_n11865_, new_n11866_, new_n11867_, new_n11868_, new_n11869_,
    new_n11870_, new_n11871_, new_n11872_, new_n11873_, new_n11874_,
    new_n11875_, new_n11876_, new_n11877_, new_n11878_, new_n11879_,
    new_n11880_, new_n11881_, new_n11882_, new_n11883_, new_n11884_,
    new_n11885_, new_n11886_, new_n11887_, new_n11888_, new_n11889_,
    new_n11890_, new_n11891_, new_n11892_, new_n11893_, new_n11894_,
    new_n11895_, new_n11896_, new_n11897_, new_n11898_, new_n11899_,
    new_n11900_, new_n11901_, new_n11902_, new_n11904_, new_n11905_,
    new_n11906_, new_n11907_, new_n11908_, new_n11909_, new_n11910_,
    new_n11911_, new_n11912_, new_n11913_, new_n11914_, new_n11915_,
    new_n11916_, new_n11917_, new_n11918_, new_n11919_, new_n11920_,
    new_n11921_, new_n11922_, new_n11923_, new_n11924_, new_n11925_,
    new_n11926_, new_n11927_, new_n11928_, new_n11929_, new_n11930_,
    new_n11931_, new_n11932_, new_n11933_, new_n11934_, new_n11935_,
    new_n11936_, new_n11937_, new_n11938_, new_n11939_, new_n11940_,
    new_n11941_, new_n11942_, new_n11943_, new_n11944_, new_n11945_,
    new_n11946_, new_n11947_, new_n11948_, new_n11949_, new_n11950_,
    new_n11951_, new_n11952_, new_n11953_, new_n11954_, new_n11955_,
    new_n11956_, new_n11957_, new_n11958_, new_n11959_, new_n11960_,
    new_n11961_, new_n11962_, new_n11963_, new_n11964_, new_n11965_,
    new_n11966_, new_n11967_, new_n11968_, new_n11969_, new_n11970_,
    new_n11971_, new_n11972_, new_n11973_, new_n11974_, new_n11975_,
    new_n11976_, new_n11977_, new_n11978_, new_n11979_, new_n11980_,
    new_n11981_, new_n11982_, new_n11983_, new_n11984_, new_n11985_,
    new_n11986_, new_n11987_, new_n11988_, new_n11990_, new_n11991_,
    new_n11992_, new_n11993_, new_n11994_, new_n11995_, new_n11996_,
    new_n11997_, new_n11998_, new_n11999_, new_n12000_, new_n12001_,
    new_n12002_, new_n12003_, new_n12004_, new_n12005_, new_n12006_,
    new_n12007_, new_n12008_, new_n12009_, new_n12010_, new_n12011_,
    new_n12012_, new_n12013_, new_n12014_, new_n12015_, new_n12016_,
    new_n12017_, new_n12018_, new_n12019_, new_n12020_, new_n12021_,
    new_n12022_, new_n12023_, new_n12024_, new_n12025_, new_n12026_,
    new_n12027_, new_n12028_, new_n12029_, new_n12030_, new_n12031_,
    new_n12032_, new_n12033_, new_n12034_, new_n12035_, new_n12036_,
    new_n12037_, new_n12038_, new_n12039_, new_n12040_, new_n12041_,
    new_n12042_, new_n12043_, new_n12044_, new_n12045_, new_n12046_,
    new_n12047_, new_n12048_, new_n12049_, new_n12050_, new_n12051_,
    new_n12052_, new_n12053_, new_n12054_, new_n12055_, new_n12056_,
    new_n12057_, new_n12058_, new_n12059_, new_n12060_, new_n12061_,
    new_n12062_, new_n12063_, new_n12064_, new_n12065_, new_n12066_,
    new_n12067_, new_n12068_, new_n12069_, new_n12070_, new_n12071_,
    new_n12072_, new_n12073_, new_n12074_, new_n12076_, new_n12077_,
    new_n12078_, new_n12079_, new_n12080_, new_n12081_, new_n12082_,
    new_n12083_, new_n12084_, new_n12085_, new_n12086_, new_n12087_,
    new_n12088_, new_n12089_, new_n12090_, new_n12091_, new_n12092_,
    new_n12093_, new_n12094_, new_n12095_, new_n12096_, new_n12097_,
    new_n12098_, new_n12099_, new_n12100_, new_n12101_, new_n12102_,
    new_n12103_, new_n12104_, new_n12105_, new_n12106_, new_n12107_,
    new_n12108_, new_n12109_, new_n12110_, new_n12111_, new_n12112_,
    new_n12113_, new_n12114_, new_n12115_, new_n12116_, new_n12117_,
    new_n12118_, new_n12119_, new_n12120_, new_n12121_, new_n12122_,
    new_n12123_, new_n12124_, new_n12125_, new_n12126_, new_n12127_,
    new_n12128_, new_n12129_, new_n12130_, new_n12131_, new_n12132_,
    new_n12133_, new_n12134_, new_n12135_, new_n12136_, new_n12137_,
    new_n12138_, new_n12139_, new_n12140_, new_n12141_, new_n12142_,
    new_n12143_, new_n12144_, new_n12145_, new_n12146_, new_n12147_,
    new_n12148_, new_n12149_, new_n12150_, new_n12151_, new_n12152_,
    new_n12153_, new_n12154_, new_n12155_, new_n12156_, new_n12157_,
    new_n12158_, new_n12159_, new_n12160_, new_n12162_, new_n12163_,
    new_n12164_, new_n12165_, new_n12166_, new_n12167_, new_n12168_,
    new_n12169_, new_n12170_, new_n12171_, new_n12172_, new_n12173_,
    new_n12174_, new_n12175_, new_n12176_, new_n12177_, new_n12178_,
    new_n12179_, new_n12180_, new_n12181_, new_n12182_, new_n12183_,
    new_n12184_, new_n12185_, new_n12186_, new_n12187_, new_n12188_,
    new_n12189_, new_n12190_, new_n12191_, new_n12192_, new_n12193_,
    new_n12194_, new_n12195_, new_n12196_, new_n12197_, new_n12198_,
    new_n12199_, new_n12200_, new_n12201_, new_n12202_, new_n12203_,
    new_n12204_, new_n12205_, new_n12206_, new_n12207_, new_n12208_,
    new_n12209_, new_n12210_, new_n12211_, new_n12212_, new_n12213_,
    new_n12214_, new_n12215_, new_n12216_, new_n12217_, new_n12218_,
    new_n12219_, new_n12220_, new_n12221_, new_n12222_, new_n12223_;
  assign new_n386_ = \priority[1]  & ~\req[1] ;
  assign new_n387_ = ~\priority[2]  & ~new_n386_;
  assign new_n388_ = ~\req[2]  & ~\req[3] ;
  assign new_n389_ = ~new_n387_ & new_n388_;
  assign new_n390_ = \priority[3]  & ~\req[3] ;
  assign new_n391_ = ~\priority[4]  & ~new_n390_;
  assign new_n392_ = ~\priority[5]  & new_n391_;
  assign new_n393_ = ~new_n389_ & new_n392_;
  assign new_n394_ = ~\priority[5]  & \req[4] ;
  assign new_n395_ = ~\req[5]  & ~\req[6] ;
  assign new_n396_ = ~new_n394_ & new_n395_;
  assign new_n397_ = ~new_n393_ & new_n396_;
  assign new_n398_ = \priority[6]  & ~\req[6] ;
  assign new_n399_ = ~\priority[7]  & ~new_n398_;
  assign new_n400_ = ~\priority[8]  & new_n399_;
  assign new_n401_ = ~new_n397_ & new_n400_;
  assign new_n402_ = ~\priority[8]  & \req[7] ;
  assign new_n403_ = ~\req[8]  & ~\req[9] ;
  assign new_n404_ = ~new_n402_ & new_n403_;
  assign new_n405_ = ~new_n401_ & new_n404_;
  assign new_n406_ = \priority[9]  & ~\req[9] ;
  assign new_n407_ = ~\priority[10]  & ~new_n406_;
  assign new_n408_ = ~\priority[11]  & new_n407_;
  assign new_n409_ = ~new_n405_ & new_n408_;
  assign new_n410_ = ~\priority[11]  & \req[10] ;
  assign new_n411_ = ~\req[11]  & ~\req[12] ;
  assign new_n412_ = ~new_n410_ & new_n411_;
  assign new_n413_ = ~new_n409_ & new_n412_;
  assign new_n414_ = \priority[12]  & ~\req[12] ;
  assign new_n415_ = ~\priority[13]  & ~new_n414_;
  assign new_n416_ = ~\priority[14]  & new_n415_;
  assign new_n417_ = ~new_n413_ & new_n416_;
  assign new_n418_ = ~\priority[14]  & \req[13] ;
  assign new_n419_ = ~\req[14]  & ~\req[15] ;
  assign new_n420_ = ~new_n418_ & new_n419_;
  assign new_n421_ = ~new_n417_ & new_n420_;
  assign new_n422_ = \priority[15]  & ~\req[15] ;
  assign new_n423_ = ~\priority[16]  & ~new_n422_;
  assign new_n424_ = ~\priority[17]  & new_n423_;
  assign new_n425_ = ~new_n421_ & new_n424_;
  assign new_n426_ = ~\priority[17]  & \req[16] ;
  assign new_n427_ = ~\req[17]  & ~\req[18] ;
  assign new_n428_ = ~new_n426_ & new_n427_;
  assign new_n429_ = ~new_n425_ & new_n428_;
  assign new_n430_ = \priority[18]  & ~\req[18] ;
  assign new_n431_ = ~\priority[19]  & ~new_n430_;
  assign new_n432_ = ~\priority[20]  & new_n431_;
  assign new_n433_ = ~new_n429_ & new_n432_;
  assign new_n434_ = ~\priority[20]  & \req[19] ;
  assign new_n435_ = ~\req[20]  & ~\req[21] ;
  assign new_n436_ = ~new_n434_ & new_n435_;
  assign new_n437_ = ~new_n433_ & new_n436_;
  assign new_n438_ = \priority[21]  & ~\req[21] ;
  assign new_n439_ = ~\priority[22]  & ~new_n438_;
  assign new_n440_ = ~\priority[23]  & new_n439_;
  assign new_n441_ = ~new_n437_ & new_n440_;
  assign new_n442_ = ~\priority[23]  & \req[22] ;
  assign new_n443_ = ~\req[23]  & ~\req[24] ;
  assign new_n444_ = ~new_n442_ & new_n443_;
  assign new_n445_ = ~new_n441_ & new_n444_;
  assign new_n446_ = \priority[24]  & ~\req[24] ;
  assign new_n447_ = ~\priority[25]  & ~new_n446_;
  assign new_n448_ = ~\priority[26]  & new_n447_;
  assign new_n449_ = ~new_n445_ & new_n448_;
  assign new_n450_ = ~\priority[26]  & \req[25] ;
  assign new_n451_ = ~\req[26]  & ~\req[27] ;
  assign new_n452_ = ~new_n450_ & new_n451_;
  assign new_n453_ = ~new_n449_ & new_n452_;
  assign new_n454_ = \priority[27]  & ~\req[27] ;
  assign new_n455_ = ~\priority[28]  & ~new_n454_;
  assign new_n456_ = ~\priority[29]  & new_n455_;
  assign new_n457_ = ~new_n453_ & new_n456_;
  assign new_n458_ = ~\priority[29]  & \req[28] ;
  assign new_n459_ = ~\req[29]  & ~\req[30] ;
  assign new_n460_ = ~new_n458_ & new_n459_;
  assign new_n461_ = ~new_n457_ & new_n460_;
  assign new_n462_ = \priority[30]  & ~\req[30] ;
  assign new_n463_ = ~\priority[31]  & ~new_n462_;
  assign new_n464_ = ~\priority[32]  & new_n463_;
  assign new_n465_ = ~new_n461_ & new_n464_;
  assign new_n466_ = ~\priority[32]  & \req[31] ;
  assign new_n467_ = ~\req[32]  & ~\req[33] ;
  assign new_n468_ = ~new_n466_ & new_n467_;
  assign new_n469_ = ~new_n465_ & new_n468_;
  assign new_n470_ = \priority[33]  & ~\req[33] ;
  assign new_n471_ = ~\priority[34]  & ~new_n470_;
  assign new_n472_ = ~\priority[35]  & new_n471_;
  assign new_n473_ = ~new_n469_ & new_n472_;
  assign new_n474_ = ~\priority[35]  & \req[34] ;
  assign new_n475_ = ~\req[35]  & ~\req[36] ;
  assign new_n476_ = ~new_n474_ & new_n475_;
  assign new_n477_ = ~new_n473_ & new_n476_;
  assign new_n478_ = \priority[36]  & ~\req[36] ;
  assign new_n479_ = ~\priority[37]  & ~new_n478_;
  assign new_n480_ = ~\priority[38]  & new_n479_;
  assign new_n481_ = ~new_n477_ & new_n480_;
  assign new_n482_ = ~\priority[38]  & \req[37] ;
  assign new_n483_ = ~\req[38]  & ~\req[39] ;
  assign new_n484_ = ~new_n482_ & new_n483_;
  assign new_n485_ = ~new_n481_ & new_n484_;
  assign new_n486_ = \priority[39]  & ~\req[39] ;
  assign new_n487_ = ~\priority[40]  & ~new_n486_;
  assign new_n488_ = ~\priority[41]  & new_n487_;
  assign new_n489_ = ~new_n485_ & new_n488_;
  assign new_n490_ = ~\priority[41]  & \req[40] ;
  assign new_n491_ = ~\req[41]  & ~\req[42] ;
  assign new_n492_ = ~new_n490_ & new_n491_;
  assign new_n493_ = ~new_n489_ & new_n492_;
  assign new_n494_ = \priority[42]  & ~\req[42] ;
  assign new_n495_ = ~\priority[43]  & ~new_n494_;
  assign new_n496_ = ~\priority[44]  & new_n495_;
  assign new_n497_ = ~new_n493_ & new_n496_;
  assign new_n498_ = ~\priority[44]  & \req[43] ;
  assign new_n499_ = ~\req[44]  & ~\req[45] ;
  assign new_n500_ = ~new_n498_ & new_n499_;
  assign new_n501_ = ~new_n497_ & new_n500_;
  assign new_n502_ = \priority[45]  & ~\req[45] ;
  assign new_n503_ = ~\priority[46]  & ~new_n502_;
  assign new_n504_ = ~\priority[47]  & new_n503_;
  assign new_n505_ = ~new_n501_ & new_n504_;
  assign new_n506_ = ~\priority[47]  & \req[46] ;
  assign new_n507_ = ~\req[47]  & ~\req[48] ;
  assign new_n508_ = ~new_n506_ & new_n507_;
  assign new_n509_ = ~new_n505_ & new_n508_;
  assign new_n510_ = \priority[48]  & ~\req[48] ;
  assign new_n511_ = ~\priority[49]  & ~new_n510_;
  assign new_n512_ = ~\priority[50]  & new_n511_;
  assign new_n513_ = ~new_n509_ & new_n512_;
  assign new_n514_ = ~\priority[50]  & \req[49] ;
  assign new_n515_ = ~\req[50]  & ~\req[51] ;
  assign new_n516_ = ~new_n514_ & new_n515_;
  assign new_n517_ = ~new_n513_ & new_n516_;
  assign new_n518_ = \priority[51]  & ~\req[51] ;
  assign new_n519_ = ~\priority[52]  & ~new_n518_;
  assign new_n520_ = ~\priority[53]  & new_n519_;
  assign new_n521_ = ~new_n517_ & new_n520_;
  assign new_n522_ = ~\priority[53]  & \req[52] ;
  assign new_n523_ = ~\req[53]  & ~\req[54] ;
  assign new_n524_ = ~new_n522_ & new_n523_;
  assign new_n525_ = ~new_n521_ & new_n524_;
  assign new_n526_ = \priority[54]  & ~\req[54] ;
  assign new_n527_ = ~\priority[55]  & ~new_n526_;
  assign new_n528_ = ~\priority[56]  & new_n527_;
  assign new_n529_ = ~new_n525_ & new_n528_;
  assign new_n530_ = ~\priority[56]  & \req[55] ;
  assign new_n531_ = ~\req[56]  & ~\req[57] ;
  assign new_n532_ = ~new_n530_ & new_n531_;
  assign new_n533_ = ~new_n529_ & new_n532_;
  assign new_n534_ = \priority[57]  & ~\req[57] ;
  assign new_n535_ = ~\priority[58]  & ~new_n534_;
  assign new_n536_ = ~\priority[59]  & new_n535_;
  assign new_n537_ = ~new_n533_ & new_n536_;
  assign new_n538_ = ~\priority[59]  & \req[58] ;
  assign new_n539_ = ~\req[59]  & ~\req[60] ;
  assign new_n540_ = ~new_n538_ & new_n539_;
  assign new_n541_ = ~new_n537_ & new_n540_;
  assign new_n542_ = \priority[60]  & ~\req[60] ;
  assign new_n543_ = ~\priority[61]  & ~new_n542_;
  assign new_n544_ = ~\priority[62]  & new_n543_;
  assign new_n545_ = ~new_n541_ & new_n544_;
  assign new_n546_ = ~\priority[62]  & \req[61] ;
  assign new_n547_ = ~\req[62]  & ~\req[63] ;
  assign new_n548_ = ~new_n546_ & new_n547_;
  assign new_n549_ = ~new_n545_ & new_n548_;
  assign new_n550_ = \priority[63]  & ~\req[63] ;
  assign new_n551_ = ~\priority[64]  & ~new_n550_;
  assign new_n552_ = ~\priority[65]  & new_n551_;
  assign new_n553_ = ~new_n549_ & new_n552_;
  assign new_n554_ = ~\priority[65]  & \req[64] ;
  assign new_n555_ = ~\req[65]  & ~\req[66] ;
  assign new_n556_ = ~new_n554_ & new_n555_;
  assign new_n557_ = ~new_n553_ & new_n556_;
  assign new_n558_ = \priority[66]  & ~\req[66] ;
  assign new_n559_ = ~\priority[67]  & ~new_n558_;
  assign new_n560_ = ~\priority[68]  & new_n559_;
  assign new_n561_ = ~new_n557_ & new_n560_;
  assign new_n562_ = ~\priority[68]  & \req[67] ;
  assign new_n563_ = ~\req[68]  & ~\req[69] ;
  assign new_n564_ = ~new_n562_ & new_n563_;
  assign new_n565_ = ~new_n561_ & new_n564_;
  assign new_n566_ = \priority[69]  & ~\req[69] ;
  assign new_n567_ = ~\priority[70]  & ~new_n566_;
  assign new_n568_ = ~\priority[71]  & new_n567_;
  assign new_n569_ = ~new_n565_ & new_n568_;
  assign new_n570_ = ~\priority[71]  & \req[70] ;
  assign new_n571_ = ~\req[71]  & ~\req[72] ;
  assign new_n572_ = ~new_n570_ & new_n571_;
  assign new_n573_ = ~new_n569_ & new_n572_;
  assign new_n574_ = \priority[72]  & ~\req[72] ;
  assign new_n575_ = ~\priority[73]  & ~new_n574_;
  assign new_n576_ = ~\priority[74]  & new_n575_;
  assign new_n577_ = ~new_n573_ & new_n576_;
  assign new_n578_ = ~\priority[74]  & \req[73] ;
  assign new_n579_ = ~\req[74]  & ~\req[75] ;
  assign new_n580_ = ~new_n578_ & new_n579_;
  assign new_n581_ = ~new_n577_ & new_n580_;
  assign new_n582_ = \priority[75]  & ~\req[75] ;
  assign new_n583_ = ~\priority[76]  & ~new_n582_;
  assign new_n584_ = ~\priority[77]  & new_n583_;
  assign new_n585_ = ~new_n581_ & new_n584_;
  assign new_n586_ = ~\priority[77]  & \req[76] ;
  assign new_n587_ = ~\req[77]  & ~\req[78] ;
  assign new_n588_ = ~new_n586_ & new_n587_;
  assign new_n589_ = ~new_n585_ & new_n588_;
  assign new_n590_ = \priority[78]  & ~\req[78] ;
  assign new_n591_ = ~\priority[79]  & ~new_n590_;
  assign new_n592_ = ~\priority[80]  & new_n591_;
  assign new_n593_ = ~new_n589_ & new_n592_;
  assign new_n594_ = ~\priority[80]  & \req[79] ;
  assign new_n595_ = ~\req[80]  & ~\req[81] ;
  assign new_n596_ = ~new_n594_ & new_n595_;
  assign new_n597_ = ~new_n593_ & new_n596_;
  assign new_n598_ = \priority[81]  & ~\req[81] ;
  assign new_n599_ = ~\priority[82]  & ~new_n598_;
  assign new_n600_ = ~\priority[83]  & new_n599_;
  assign new_n601_ = ~new_n597_ & new_n600_;
  assign new_n602_ = ~\priority[83]  & \req[82] ;
  assign new_n603_ = ~\req[83]  & ~\req[84] ;
  assign new_n604_ = ~new_n602_ & new_n603_;
  assign new_n605_ = ~new_n601_ & new_n604_;
  assign new_n606_ = \priority[84]  & ~\req[84] ;
  assign new_n607_ = ~\priority[85]  & ~new_n606_;
  assign new_n608_ = ~\priority[86]  & new_n607_;
  assign new_n609_ = ~new_n605_ & new_n608_;
  assign new_n610_ = ~\priority[86]  & \req[85] ;
  assign new_n611_ = ~\req[86]  & ~\req[87] ;
  assign new_n612_ = ~new_n610_ & new_n611_;
  assign new_n613_ = ~new_n609_ & new_n612_;
  assign new_n614_ = \priority[87]  & ~\req[87] ;
  assign new_n615_ = ~\priority[88]  & ~new_n614_;
  assign new_n616_ = ~\priority[89]  & new_n615_;
  assign new_n617_ = ~new_n613_ & new_n616_;
  assign new_n618_ = ~\priority[89]  & \req[88] ;
  assign new_n619_ = ~\req[89]  & ~\req[90] ;
  assign new_n620_ = ~new_n618_ & new_n619_;
  assign new_n621_ = ~new_n617_ & new_n620_;
  assign new_n622_ = \priority[90]  & ~\req[90] ;
  assign new_n623_ = ~\priority[91]  & ~new_n622_;
  assign new_n624_ = ~\priority[92]  & new_n623_;
  assign new_n625_ = ~new_n621_ & new_n624_;
  assign new_n626_ = ~\priority[92]  & \req[91] ;
  assign new_n627_ = ~\req[92]  & ~\req[93] ;
  assign new_n628_ = ~new_n626_ & new_n627_;
  assign new_n629_ = ~new_n625_ & new_n628_;
  assign new_n630_ = \priority[93]  & ~\req[93] ;
  assign new_n631_ = ~\priority[94]  & ~new_n630_;
  assign new_n632_ = ~\priority[95]  & new_n631_;
  assign new_n633_ = ~new_n629_ & new_n632_;
  assign new_n634_ = ~\priority[95]  & \req[94] ;
  assign new_n635_ = ~\req[95]  & ~\req[96] ;
  assign new_n636_ = ~new_n634_ & new_n635_;
  assign new_n637_ = ~new_n633_ & new_n636_;
  assign new_n638_ = \priority[96]  & ~\req[96] ;
  assign new_n639_ = ~\priority[97]  & ~new_n638_;
  assign new_n640_ = ~\priority[98]  & new_n639_;
  assign new_n641_ = ~new_n637_ & new_n640_;
  assign new_n642_ = ~\priority[98]  & \req[97] ;
  assign new_n643_ = ~\req[98]  & ~\req[99] ;
  assign new_n644_ = ~new_n642_ & new_n643_;
  assign new_n645_ = ~new_n641_ & new_n644_;
  assign new_n646_ = \priority[99]  & ~\req[99] ;
  assign new_n647_ = ~\priority[100]  & ~new_n646_;
  assign new_n648_ = ~\priority[101]  & new_n647_;
  assign new_n649_ = ~new_n645_ & new_n648_;
  assign new_n650_ = ~\priority[101]  & \req[100] ;
  assign new_n651_ = ~\req[101]  & ~\req[102] ;
  assign new_n652_ = ~new_n650_ & new_n651_;
  assign new_n653_ = ~new_n649_ & new_n652_;
  assign new_n654_ = \priority[102]  & ~\req[102] ;
  assign new_n655_ = ~\priority[103]  & ~new_n654_;
  assign new_n656_ = ~\priority[104]  & new_n655_;
  assign new_n657_ = ~new_n653_ & new_n656_;
  assign new_n658_ = ~\priority[104]  & \req[103] ;
  assign new_n659_ = ~\req[104]  & ~\req[105] ;
  assign new_n660_ = ~new_n658_ & new_n659_;
  assign new_n661_ = ~new_n657_ & new_n660_;
  assign new_n662_ = \priority[105]  & ~\req[105] ;
  assign new_n663_ = ~\priority[106]  & ~new_n662_;
  assign new_n664_ = ~\priority[107]  & new_n663_;
  assign new_n665_ = ~new_n661_ & new_n664_;
  assign new_n666_ = ~\priority[107]  & \req[106] ;
  assign new_n667_ = ~\req[107]  & ~\req[108] ;
  assign new_n668_ = ~new_n666_ & new_n667_;
  assign new_n669_ = ~new_n665_ & new_n668_;
  assign new_n670_ = \priority[108]  & ~\req[108] ;
  assign new_n671_ = ~\priority[109]  & ~new_n670_;
  assign new_n672_ = ~\priority[110]  & new_n671_;
  assign new_n673_ = ~new_n669_ & new_n672_;
  assign new_n674_ = ~\priority[110]  & \req[109] ;
  assign new_n675_ = ~\req[110]  & ~\req[111] ;
  assign new_n676_ = ~new_n674_ & new_n675_;
  assign new_n677_ = ~new_n673_ & new_n676_;
  assign new_n678_ = \priority[111]  & ~\req[111] ;
  assign new_n679_ = ~\priority[112]  & ~new_n678_;
  assign new_n680_ = ~\priority[113]  & new_n679_;
  assign new_n681_ = ~new_n677_ & new_n680_;
  assign new_n682_ = ~\priority[113]  & \req[112] ;
  assign new_n683_ = ~\req[113]  & ~\req[114] ;
  assign new_n684_ = ~new_n682_ & new_n683_;
  assign new_n685_ = ~new_n681_ & new_n684_;
  assign new_n686_ = \priority[114]  & ~\req[114] ;
  assign new_n687_ = ~\priority[115]  & ~new_n686_;
  assign new_n688_ = ~\priority[116]  & new_n687_;
  assign new_n689_ = ~new_n685_ & new_n688_;
  assign new_n690_ = ~\priority[116]  & \req[115] ;
  assign new_n691_ = ~\req[116]  & ~\req[117] ;
  assign new_n692_ = ~new_n690_ & new_n691_;
  assign new_n693_ = ~new_n689_ & new_n692_;
  assign new_n694_ = \priority[117]  & ~\req[117] ;
  assign new_n695_ = ~\priority[118]  & ~new_n694_;
  assign new_n696_ = ~\priority[119]  & new_n695_;
  assign new_n697_ = ~new_n693_ & new_n696_;
  assign new_n698_ = ~\priority[119]  & \req[118] ;
  assign new_n699_ = ~\req[119]  & ~\req[120] ;
  assign new_n700_ = ~new_n698_ & new_n699_;
  assign new_n701_ = ~new_n697_ & new_n700_;
  assign new_n702_ = \priority[120]  & ~\req[120] ;
  assign new_n703_ = ~\priority[121]  & ~new_n702_;
  assign new_n704_ = ~\priority[122]  & new_n703_;
  assign new_n705_ = ~new_n701_ & new_n704_;
  assign new_n706_ = ~\priority[122]  & \req[121] ;
  assign new_n707_ = ~\req[122]  & ~\req[123] ;
  assign new_n708_ = ~new_n706_ & new_n707_;
  assign new_n709_ = ~new_n705_ & new_n708_;
  assign new_n710_ = \priority[123]  & ~\req[123] ;
  assign new_n711_ = ~\priority[124]  & ~new_n710_;
  assign new_n712_ = ~\priority[125]  & new_n711_;
  assign new_n713_ = ~new_n709_ & new_n712_;
  assign new_n714_ = ~\priority[125]  & \req[124] ;
  assign new_n715_ = ~\req[125]  & ~\req[126] ;
  assign new_n716_ = ~new_n714_ & new_n715_;
  assign new_n717_ = ~new_n713_ & new_n716_;
  assign new_n718_ = \priority[126]  & ~\req[126] ;
  assign new_n719_ = ~\priority[127]  & ~new_n718_;
  assign new_n720_ = ~\priority[0]  & new_n719_;
  assign new_n721_ = ~new_n717_ & new_n720_;
  assign new_n722_ = ~\priority[0]  & \req[127] ;
  assign new_n723_ = \req[0]  & ~new_n722_;
  assign \grant[0]  = ~new_n721_ & new_n723_;
  assign new_n725_ = \priority[2]  & ~\req[2] ;
  assign new_n726_ = ~\priority[3]  & ~new_n725_;
  assign new_n727_ = ~\req[3]  & ~\req[4] ;
  assign new_n728_ = ~new_n726_ & new_n727_;
  assign new_n729_ = \priority[4]  & ~\req[4] ;
  assign new_n730_ = ~\priority[5]  & ~new_n729_;
  assign new_n731_ = ~\priority[6]  & new_n730_;
  assign new_n732_ = ~new_n728_ & new_n731_;
  assign new_n733_ = ~\priority[6]  & \req[5] ;
  assign new_n734_ = ~\req[6]  & ~\req[7] ;
  assign new_n735_ = ~new_n733_ & new_n734_;
  assign new_n736_ = ~new_n732_ & new_n735_;
  assign new_n737_ = \priority[7]  & ~\req[7] ;
  assign new_n738_ = ~\priority[8]  & ~new_n737_;
  assign new_n739_ = ~\priority[9]  & new_n738_;
  assign new_n740_ = ~new_n736_ & new_n739_;
  assign new_n741_ = ~\priority[9]  & \req[8] ;
  assign new_n742_ = ~\req[9]  & ~\req[10] ;
  assign new_n743_ = ~new_n741_ & new_n742_;
  assign new_n744_ = ~new_n740_ & new_n743_;
  assign new_n745_ = \priority[10]  & ~\req[10] ;
  assign new_n746_ = ~\priority[11]  & ~new_n745_;
  assign new_n747_ = ~\priority[12]  & new_n746_;
  assign new_n748_ = ~new_n744_ & new_n747_;
  assign new_n749_ = ~\priority[12]  & \req[11] ;
  assign new_n750_ = ~\req[12]  & ~\req[13] ;
  assign new_n751_ = ~new_n749_ & new_n750_;
  assign new_n752_ = ~new_n748_ & new_n751_;
  assign new_n753_ = \priority[13]  & ~\req[13] ;
  assign new_n754_ = ~\priority[14]  & ~new_n753_;
  assign new_n755_ = ~\priority[15]  & new_n754_;
  assign new_n756_ = ~new_n752_ & new_n755_;
  assign new_n757_ = ~\priority[15]  & \req[14] ;
  assign new_n758_ = ~\req[15]  & ~\req[16] ;
  assign new_n759_ = ~new_n757_ & new_n758_;
  assign new_n760_ = ~new_n756_ & new_n759_;
  assign new_n761_ = \priority[16]  & ~\req[16] ;
  assign new_n762_ = ~\priority[17]  & ~new_n761_;
  assign new_n763_ = ~\priority[18]  & new_n762_;
  assign new_n764_ = ~new_n760_ & new_n763_;
  assign new_n765_ = ~\priority[18]  & \req[17] ;
  assign new_n766_ = ~\req[18]  & ~\req[19] ;
  assign new_n767_ = ~new_n765_ & new_n766_;
  assign new_n768_ = ~new_n764_ & new_n767_;
  assign new_n769_ = \priority[19]  & ~\req[19] ;
  assign new_n770_ = ~\priority[20]  & ~new_n769_;
  assign new_n771_ = ~\priority[21]  & new_n770_;
  assign new_n772_ = ~new_n768_ & new_n771_;
  assign new_n773_ = ~\priority[21]  & \req[20] ;
  assign new_n774_ = ~\req[21]  & ~\req[22] ;
  assign new_n775_ = ~new_n773_ & new_n774_;
  assign new_n776_ = ~new_n772_ & new_n775_;
  assign new_n777_ = \priority[22]  & ~\req[22] ;
  assign new_n778_ = ~\priority[23]  & ~new_n777_;
  assign new_n779_ = ~\priority[24]  & new_n778_;
  assign new_n780_ = ~new_n776_ & new_n779_;
  assign new_n781_ = ~\priority[24]  & \req[23] ;
  assign new_n782_ = ~\req[24]  & ~\req[25] ;
  assign new_n783_ = ~new_n781_ & new_n782_;
  assign new_n784_ = ~new_n780_ & new_n783_;
  assign new_n785_ = \priority[25]  & ~\req[25] ;
  assign new_n786_ = ~\priority[26]  & ~new_n785_;
  assign new_n787_ = ~\priority[27]  & new_n786_;
  assign new_n788_ = ~new_n784_ & new_n787_;
  assign new_n789_ = ~\priority[27]  & \req[26] ;
  assign new_n790_ = ~\req[27]  & ~\req[28] ;
  assign new_n791_ = ~new_n789_ & new_n790_;
  assign new_n792_ = ~new_n788_ & new_n791_;
  assign new_n793_ = \priority[28]  & ~\req[28] ;
  assign new_n794_ = ~\priority[29]  & ~new_n793_;
  assign new_n795_ = ~\priority[30]  & new_n794_;
  assign new_n796_ = ~new_n792_ & new_n795_;
  assign new_n797_ = ~\priority[30]  & \req[29] ;
  assign new_n798_ = ~\req[30]  & ~\req[31] ;
  assign new_n799_ = ~new_n797_ & new_n798_;
  assign new_n800_ = ~new_n796_ & new_n799_;
  assign new_n801_ = \priority[31]  & ~\req[31] ;
  assign new_n802_ = ~\priority[32]  & ~new_n801_;
  assign new_n803_ = ~\priority[33]  & new_n802_;
  assign new_n804_ = ~new_n800_ & new_n803_;
  assign new_n805_ = ~\priority[33]  & \req[32] ;
  assign new_n806_ = ~\req[33]  & ~\req[34] ;
  assign new_n807_ = ~new_n805_ & new_n806_;
  assign new_n808_ = ~new_n804_ & new_n807_;
  assign new_n809_ = \priority[34]  & ~\req[34] ;
  assign new_n810_ = ~\priority[35]  & ~new_n809_;
  assign new_n811_ = ~\priority[36]  & new_n810_;
  assign new_n812_ = ~new_n808_ & new_n811_;
  assign new_n813_ = ~\priority[36]  & \req[35] ;
  assign new_n814_ = ~\req[36]  & ~\req[37] ;
  assign new_n815_ = ~new_n813_ & new_n814_;
  assign new_n816_ = ~new_n812_ & new_n815_;
  assign new_n817_ = \priority[37]  & ~\req[37] ;
  assign new_n818_ = ~\priority[38]  & ~new_n817_;
  assign new_n819_ = ~\priority[39]  & new_n818_;
  assign new_n820_ = ~new_n816_ & new_n819_;
  assign new_n821_ = ~\priority[39]  & \req[38] ;
  assign new_n822_ = ~\req[39]  & ~\req[40] ;
  assign new_n823_ = ~new_n821_ & new_n822_;
  assign new_n824_ = ~new_n820_ & new_n823_;
  assign new_n825_ = \priority[40]  & ~\req[40] ;
  assign new_n826_ = ~\priority[41]  & ~new_n825_;
  assign new_n827_ = ~\priority[42]  & new_n826_;
  assign new_n828_ = ~new_n824_ & new_n827_;
  assign new_n829_ = ~\priority[42]  & \req[41] ;
  assign new_n830_ = ~\req[42]  & ~\req[43] ;
  assign new_n831_ = ~new_n829_ & new_n830_;
  assign new_n832_ = ~new_n828_ & new_n831_;
  assign new_n833_ = \priority[43]  & ~\req[43] ;
  assign new_n834_ = ~\priority[44]  & ~new_n833_;
  assign new_n835_ = ~\priority[45]  & new_n834_;
  assign new_n836_ = ~new_n832_ & new_n835_;
  assign new_n837_ = ~\priority[45]  & \req[44] ;
  assign new_n838_ = ~\req[45]  & ~\req[46] ;
  assign new_n839_ = ~new_n837_ & new_n838_;
  assign new_n840_ = ~new_n836_ & new_n839_;
  assign new_n841_ = \priority[46]  & ~\req[46] ;
  assign new_n842_ = ~\priority[47]  & ~new_n841_;
  assign new_n843_ = ~\priority[48]  & new_n842_;
  assign new_n844_ = ~new_n840_ & new_n843_;
  assign new_n845_ = ~\priority[48]  & \req[47] ;
  assign new_n846_ = ~\req[48]  & ~\req[49] ;
  assign new_n847_ = ~new_n845_ & new_n846_;
  assign new_n848_ = ~new_n844_ & new_n847_;
  assign new_n849_ = \priority[49]  & ~\req[49] ;
  assign new_n850_ = ~\priority[50]  & ~new_n849_;
  assign new_n851_ = ~\priority[51]  & new_n850_;
  assign new_n852_ = ~new_n848_ & new_n851_;
  assign new_n853_ = ~\priority[51]  & \req[50] ;
  assign new_n854_ = ~\req[51]  & ~\req[52] ;
  assign new_n855_ = ~new_n853_ & new_n854_;
  assign new_n856_ = ~new_n852_ & new_n855_;
  assign new_n857_ = \priority[52]  & ~\req[52] ;
  assign new_n858_ = ~\priority[53]  & ~new_n857_;
  assign new_n859_ = ~\priority[54]  & new_n858_;
  assign new_n860_ = ~new_n856_ & new_n859_;
  assign new_n861_ = ~\priority[54]  & \req[53] ;
  assign new_n862_ = ~\req[54]  & ~\req[55] ;
  assign new_n863_ = ~new_n861_ & new_n862_;
  assign new_n864_ = ~new_n860_ & new_n863_;
  assign new_n865_ = \priority[55]  & ~\req[55] ;
  assign new_n866_ = ~\priority[56]  & ~new_n865_;
  assign new_n867_ = ~\priority[57]  & new_n866_;
  assign new_n868_ = ~new_n864_ & new_n867_;
  assign new_n869_ = ~\priority[57]  & \req[56] ;
  assign new_n870_ = ~\req[57]  & ~\req[58] ;
  assign new_n871_ = ~new_n869_ & new_n870_;
  assign new_n872_ = ~new_n868_ & new_n871_;
  assign new_n873_ = \priority[58]  & ~\req[58] ;
  assign new_n874_ = ~\priority[59]  & ~new_n873_;
  assign new_n875_ = ~\priority[60]  & new_n874_;
  assign new_n876_ = ~new_n872_ & new_n875_;
  assign new_n877_ = ~\priority[60]  & \req[59] ;
  assign new_n878_ = ~\req[60]  & ~\req[61] ;
  assign new_n879_ = ~new_n877_ & new_n878_;
  assign new_n880_ = ~new_n876_ & new_n879_;
  assign new_n881_ = \priority[61]  & ~\req[61] ;
  assign new_n882_ = ~\priority[62]  & ~new_n881_;
  assign new_n883_ = ~\priority[63]  & new_n882_;
  assign new_n884_ = ~new_n880_ & new_n883_;
  assign new_n885_ = ~\priority[63]  & \req[62] ;
  assign new_n886_ = ~\req[63]  & ~\req[64] ;
  assign new_n887_ = ~new_n885_ & new_n886_;
  assign new_n888_ = ~new_n884_ & new_n887_;
  assign new_n889_ = \priority[64]  & ~\req[64] ;
  assign new_n890_ = ~\priority[65]  & ~new_n889_;
  assign new_n891_ = ~\priority[66]  & new_n890_;
  assign new_n892_ = ~new_n888_ & new_n891_;
  assign new_n893_ = ~\priority[66]  & \req[65] ;
  assign new_n894_ = ~\req[66]  & ~\req[67] ;
  assign new_n895_ = ~new_n893_ & new_n894_;
  assign new_n896_ = ~new_n892_ & new_n895_;
  assign new_n897_ = \priority[67]  & ~\req[67] ;
  assign new_n898_ = ~\priority[68]  & ~new_n897_;
  assign new_n899_ = ~\priority[69]  & new_n898_;
  assign new_n900_ = ~new_n896_ & new_n899_;
  assign new_n901_ = ~\priority[69]  & \req[68] ;
  assign new_n902_ = ~\req[69]  & ~\req[70] ;
  assign new_n903_ = ~new_n901_ & new_n902_;
  assign new_n904_ = ~new_n900_ & new_n903_;
  assign new_n905_ = \priority[70]  & ~\req[70] ;
  assign new_n906_ = ~\priority[71]  & ~new_n905_;
  assign new_n907_ = ~\priority[72]  & new_n906_;
  assign new_n908_ = ~new_n904_ & new_n907_;
  assign new_n909_ = ~\priority[72]  & \req[71] ;
  assign new_n910_ = ~\req[72]  & ~\req[73] ;
  assign new_n911_ = ~new_n909_ & new_n910_;
  assign new_n912_ = ~new_n908_ & new_n911_;
  assign new_n913_ = \priority[73]  & ~\req[73] ;
  assign new_n914_ = ~\priority[74]  & ~new_n913_;
  assign new_n915_ = ~\priority[75]  & new_n914_;
  assign new_n916_ = ~new_n912_ & new_n915_;
  assign new_n917_ = ~\priority[75]  & \req[74] ;
  assign new_n918_ = ~\req[75]  & ~\req[76] ;
  assign new_n919_ = ~new_n917_ & new_n918_;
  assign new_n920_ = ~new_n916_ & new_n919_;
  assign new_n921_ = \priority[76]  & ~\req[76] ;
  assign new_n922_ = ~\priority[77]  & ~new_n921_;
  assign new_n923_ = ~\priority[78]  & new_n922_;
  assign new_n924_ = ~new_n920_ & new_n923_;
  assign new_n925_ = ~\priority[78]  & \req[77] ;
  assign new_n926_ = ~\req[78]  & ~\req[79] ;
  assign new_n927_ = ~new_n925_ & new_n926_;
  assign new_n928_ = ~new_n924_ & new_n927_;
  assign new_n929_ = \priority[79]  & ~\req[79] ;
  assign new_n930_ = ~\priority[80]  & ~new_n929_;
  assign new_n931_ = ~\priority[81]  & new_n930_;
  assign new_n932_ = ~new_n928_ & new_n931_;
  assign new_n933_ = ~\priority[81]  & \req[80] ;
  assign new_n934_ = ~\req[81]  & ~\req[82] ;
  assign new_n935_ = ~new_n933_ & new_n934_;
  assign new_n936_ = ~new_n932_ & new_n935_;
  assign new_n937_ = \priority[82]  & ~\req[82] ;
  assign new_n938_ = ~\priority[83]  & ~new_n937_;
  assign new_n939_ = ~\priority[84]  & new_n938_;
  assign new_n940_ = ~new_n936_ & new_n939_;
  assign new_n941_ = ~\priority[84]  & \req[83] ;
  assign new_n942_ = ~\req[84]  & ~\req[85] ;
  assign new_n943_ = ~new_n941_ & new_n942_;
  assign new_n944_ = ~new_n940_ & new_n943_;
  assign new_n945_ = \priority[85]  & ~\req[85] ;
  assign new_n946_ = ~\priority[86]  & ~new_n945_;
  assign new_n947_ = ~\priority[87]  & new_n946_;
  assign new_n948_ = ~new_n944_ & new_n947_;
  assign new_n949_ = ~\priority[87]  & \req[86] ;
  assign new_n950_ = ~\req[87]  & ~\req[88] ;
  assign new_n951_ = ~new_n949_ & new_n950_;
  assign new_n952_ = ~new_n948_ & new_n951_;
  assign new_n953_ = \priority[88]  & ~\req[88] ;
  assign new_n954_ = ~\priority[89]  & ~new_n953_;
  assign new_n955_ = ~\priority[90]  & new_n954_;
  assign new_n956_ = ~new_n952_ & new_n955_;
  assign new_n957_ = ~\priority[90]  & \req[89] ;
  assign new_n958_ = ~\req[90]  & ~\req[91] ;
  assign new_n959_ = ~new_n957_ & new_n958_;
  assign new_n960_ = ~new_n956_ & new_n959_;
  assign new_n961_ = \priority[91]  & ~\req[91] ;
  assign new_n962_ = ~\priority[92]  & ~new_n961_;
  assign new_n963_ = ~\priority[93]  & new_n962_;
  assign new_n964_ = ~new_n960_ & new_n963_;
  assign new_n965_ = ~\priority[93]  & \req[92] ;
  assign new_n966_ = ~\req[93]  & ~\req[94] ;
  assign new_n967_ = ~new_n965_ & new_n966_;
  assign new_n968_ = ~new_n964_ & new_n967_;
  assign new_n969_ = \priority[94]  & ~\req[94] ;
  assign new_n970_ = ~\priority[95]  & ~new_n969_;
  assign new_n971_ = ~\priority[96]  & new_n970_;
  assign new_n972_ = ~new_n968_ & new_n971_;
  assign new_n973_ = ~\priority[96]  & \req[95] ;
  assign new_n974_ = ~\req[96]  & ~\req[97] ;
  assign new_n975_ = ~new_n973_ & new_n974_;
  assign new_n976_ = ~new_n972_ & new_n975_;
  assign new_n977_ = \priority[97]  & ~\req[97] ;
  assign new_n978_ = ~\priority[98]  & ~new_n977_;
  assign new_n979_ = ~\priority[99]  & new_n978_;
  assign new_n980_ = ~new_n976_ & new_n979_;
  assign new_n981_ = ~\priority[99]  & \req[98] ;
  assign new_n982_ = ~\req[99]  & ~\req[100] ;
  assign new_n983_ = ~new_n981_ & new_n982_;
  assign new_n984_ = ~new_n980_ & new_n983_;
  assign new_n985_ = \priority[100]  & ~\req[100] ;
  assign new_n986_ = ~\priority[101]  & ~new_n985_;
  assign new_n987_ = ~\priority[102]  & new_n986_;
  assign new_n988_ = ~new_n984_ & new_n987_;
  assign new_n989_ = ~\priority[102]  & \req[101] ;
  assign new_n990_ = ~\req[102]  & ~\req[103] ;
  assign new_n991_ = ~new_n989_ & new_n990_;
  assign new_n992_ = ~new_n988_ & new_n991_;
  assign new_n993_ = \priority[103]  & ~\req[103] ;
  assign new_n994_ = ~\priority[104]  & ~new_n993_;
  assign new_n995_ = ~\priority[105]  & new_n994_;
  assign new_n996_ = ~new_n992_ & new_n995_;
  assign new_n997_ = ~\priority[105]  & \req[104] ;
  assign new_n998_ = ~\req[105]  & ~\req[106] ;
  assign new_n999_ = ~new_n997_ & new_n998_;
  assign new_n1000_ = ~new_n996_ & new_n999_;
  assign new_n1001_ = \priority[106]  & ~\req[106] ;
  assign new_n1002_ = ~\priority[107]  & ~new_n1001_;
  assign new_n1003_ = ~\priority[108]  & new_n1002_;
  assign new_n1004_ = ~new_n1000_ & new_n1003_;
  assign new_n1005_ = ~\priority[108]  & \req[107] ;
  assign new_n1006_ = ~\req[108]  & ~\req[109] ;
  assign new_n1007_ = ~new_n1005_ & new_n1006_;
  assign new_n1008_ = ~new_n1004_ & new_n1007_;
  assign new_n1009_ = \priority[109]  & ~\req[109] ;
  assign new_n1010_ = ~\priority[110]  & ~new_n1009_;
  assign new_n1011_ = ~\priority[111]  & new_n1010_;
  assign new_n1012_ = ~new_n1008_ & new_n1011_;
  assign new_n1013_ = ~\priority[111]  & \req[110] ;
  assign new_n1014_ = ~\req[111]  & ~\req[112] ;
  assign new_n1015_ = ~new_n1013_ & new_n1014_;
  assign new_n1016_ = ~new_n1012_ & new_n1015_;
  assign new_n1017_ = \priority[112]  & ~\req[112] ;
  assign new_n1018_ = ~\priority[113]  & ~new_n1017_;
  assign new_n1019_ = ~\priority[114]  & new_n1018_;
  assign new_n1020_ = ~new_n1016_ & new_n1019_;
  assign new_n1021_ = ~\priority[114]  & \req[113] ;
  assign new_n1022_ = ~\req[114]  & ~\req[115] ;
  assign new_n1023_ = ~new_n1021_ & new_n1022_;
  assign new_n1024_ = ~new_n1020_ & new_n1023_;
  assign new_n1025_ = \priority[115]  & ~\req[115] ;
  assign new_n1026_ = ~\priority[116]  & ~new_n1025_;
  assign new_n1027_ = ~\priority[117]  & new_n1026_;
  assign new_n1028_ = ~new_n1024_ & new_n1027_;
  assign new_n1029_ = ~\priority[117]  & \req[116] ;
  assign new_n1030_ = ~\req[117]  & ~\req[118] ;
  assign new_n1031_ = ~new_n1029_ & new_n1030_;
  assign new_n1032_ = ~new_n1028_ & new_n1031_;
  assign new_n1033_ = \priority[118]  & ~\req[118] ;
  assign new_n1034_ = ~\priority[119]  & ~new_n1033_;
  assign new_n1035_ = ~\priority[120]  & new_n1034_;
  assign new_n1036_ = ~new_n1032_ & new_n1035_;
  assign new_n1037_ = ~\priority[120]  & \req[119] ;
  assign new_n1038_ = ~\req[120]  & ~\req[121] ;
  assign new_n1039_ = ~new_n1037_ & new_n1038_;
  assign new_n1040_ = ~new_n1036_ & new_n1039_;
  assign new_n1041_ = \priority[121]  & ~\req[121] ;
  assign new_n1042_ = ~\priority[122]  & ~new_n1041_;
  assign new_n1043_ = ~\priority[123]  & new_n1042_;
  assign new_n1044_ = ~new_n1040_ & new_n1043_;
  assign new_n1045_ = ~\priority[123]  & \req[122] ;
  assign new_n1046_ = ~\req[123]  & ~\req[124] ;
  assign new_n1047_ = ~new_n1045_ & new_n1046_;
  assign new_n1048_ = ~new_n1044_ & new_n1047_;
  assign new_n1049_ = \priority[124]  & ~\req[124] ;
  assign new_n1050_ = ~\priority[125]  & ~new_n1049_;
  assign new_n1051_ = ~\priority[126]  & new_n1050_;
  assign new_n1052_ = ~new_n1048_ & new_n1051_;
  assign new_n1053_ = ~\priority[126]  & \req[125] ;
  assign new_n1054_ = ~\req[126]  & ~\req[127] ;
  assign new_n1055_ = ~new_n1053_ & new_n1054_;
  assign new_n1056_ = ~new_n1052_ & new_n1055_;
  assign new_n1057_ = \priority[127]  & ~\req[127] ;
  assign new_n1058_ = ~\priority[0]  & ~new_n1057_;
  assign new_n1059_ = ~\priority[1]  & new_n1058_;
  assign new_n1060_ = ~new_n1056_ & new_n1059_;
  assign new_n1061_ = ~\priority[1]  & \req[0] ;
  assign new_n1062_ = \req[1]  & ~new_n1061_;
  assign \grant[1]  = ~new_n1060_ & new_n1062_;
  assign new_n1064_ = ~\req[4]  & ~\req[5] ;
  assign new_n1065_ = ~new_n391_ & new_n1064_;
  assign new_n1066_ = \priority[5]  & ~\req[5] ;
  assign new_n1067_ = ~\priority[6]  & ~new_n1066_;
  assign new_n1068_ = ~\priority[7]  & new_n1067_;
  assign new_n1069_ = ~new_n1065_ & new_n1068_;
  assign new_n1070_ = ~\priority[7]  & \req[6] ;
  assign new_n1071_ = ~\req[7]  & ~\req[8] ;
  assign new_n1072_ = ~new_n1070_ & new_n1071_;
  assign new_n1073_ = ~new_n1069_ & new_n1072_;
  assign new_n1074_ = \priority[8]  & ~\req[8] ;
  assign new_n1075_ = ~\priority[9]  & ~new_n1074_;
  assign new_n1076_ = ~\priority[10]  & new_n1075_;
  assign new_n1077_ = ~new_n1073_ & new_n1076_;
  assign new_n1078_ = ~\priority[10]  & \req[9] ;
  assign new_n1079_ = ~\req[10]  & ~\req[11] ;
  assign new_n1080_ = ~new_n1078_ & new_n1079_;
  assign new_n1081_ = ~new_n1077_ & new_n1080_;
  assign new_n1082_ = \priority[11]  & ~\req[11] ;
  assign new_n1083_ = ~\priority[12]  & ~new_n1082_;
  assign new_n1084_ = ~\priority[13]  & new_n1083_;
  assign new_n1085_ = ~new_n1081_ & new_n1084_;
  assign new_n1086_ = ~\priority[13]  & \req[12] ;
  assign new_n1087_ = ~\req[13]  & ~\req[14] ;
  assign new_n1088_ = ~new_n1086_ & new_n1087_;
  assign new_n1089_ = ~new_n1085_ & new_n1088_;
  assign new_n1090_ = \priority[14]  & ~\req[14] ;
  assign new_n1091_ = ~\priority[15]  & ~new_n1090_;
  assign new_n1092_ = ~\priority[16]  & new_n1091_;
  assign new_n1093_ = ~new_n1089_ & new_n1092_;
  assign new_n1094_ = ~\priority[16]  & \req[15] ;
  assign new_n1095_ = ~\req[16]  & ~\req[17] ;
  assign new_n1096_ = ~new_n1094_ & new_n1095_;
  assign new_n1097_ = ~new_n1093_ & new_n1096_;
  assign new_n1098_ = \priority[17]  & ~\req[17] ;
  assign new_n1099_ = ~\priority[18]  & ~new_n1098_;
  assign new_n1100_ = ~\priority[19]  & new_n1099_;
  assign new_n1101_ = ~new_n1097_ & new_n1100_;
  assign new_n1102_ = ~\priority[19]  & \req[18] ;
  assign new_n1103_ = ~\req[19]  & ~\req[20] ;
  assign new_n1104_ = ~new_n1102_ & new_n1103_;
  assign new_n1105_ = ~new_n1101_ & new_n1104_;
  assign new_n1106_ = \priority[20]  & ~\req[20] ;
  assign new_n1107_ = ~\priority[21]  & ~new_n1106_;
  assign new_n1108_ = ~\priority[22]  & new_n1107_;
  assign new_n1109_ = ~new_n1105_ & new_n1108_;
  assign new_n1110_ = ~\priority[22]  & \req[21] ;
  assign new_n1111_ = ~\req[22]  & ~\req[23] ;
  assign new_n1112_ = ~new_n1110_ & new_n1111_;
  assign new_n1113_ = ~new_n1109_ & new_n1112_;
  assign new_n1114_ = \priority[23]  & ~\req[23] ;
  assign new_n1115_ = ~\priority[24]  & ~new_n1114_;
  assign new_n1116_ = ~\priority[25]  & new_n1115_;
  assign new_n1117_ = ~new_n1113_ & new_n1116_;
  assign new_n1118_ = ~\priority[25]  & \req[24] ;
  assign new_n1119_ = ~\req[25]  & ~\req[26] ;
  assign new_n1120_ = ~new_n1118_ & new_n1119_;
  assign new_n1121_ = ~new_n1117_ & new_n1120_;
  assign new_n1122_ = \priority[26]  & ~\req[26] ;
  assign new_n1123_ = ~\priority[27]  & ~new_n1122_;
  assign new_n1124_ = ~\priority[28]  & new_n1123_;
  assign new_n1125_ = ~new_n1121_ & new_n1124_;
  assign new_n1126_ = ~\priority[28]  & \req[27] ;
  assign new_n1127_ = ~\req[28]  & ~\req[29] ;
  assign new_n1128_ = ~new_n1126_ & new_n1127_;
  assign new_n1129_ = ~new_n1125_ & new_n1128_;
  assign new_n1130_ = \priority[29]  & ~\req[29] ;
  assign new_n1131_ = ~\priority[30]  & ~new_n1130_;
  assign new_n1132_ = ~\priority[31]  & new_n1131_;
  assign new_n1133_ = ~new_n1129_ & new_n1132_;
  assign new_n1134_ = ~\priority[31]  & \req[30] ;
  assign new_n1135_ = ~\req[31]  & ~\req[32] ;
  assign new_n1136_ = ~new_n1134_ & new_n1135_;
  assign new_n1137_ = ~new_n1133_ & new_n1136_;
  assign new_n1138_ = \priority[32]  & ~\req[32] ;
  assign new_n1139_ = ~\priority[33]  & ~new_n1138_;
  assign new_n1140_ = ~\priority[34]  & new_n1139_;
  assign new_n1141_ = ~new_n1137_ & new_n1140_;
  assign new_n1142_ = ~\priority[34]  & \req[33] ;
  assign new_n1143_ = ~\req[34]  & ~\req[35] ;
  assign new_n1144_ = ~new_n1142_ & new_n1143_;
  assign new_n1145_ = ~new_n1141_ & new_n1144_;
  assign new_n1146_ = \priority[35]  & ~\req[35] ;
  assign new_n1147_ = ~\priority[36]  & ~new_n1146_;
  assign new_n1148_ = ~\priority[37]  & new_n1147_;
  assign new_n1149_ = ~new_n1145_ & new_n1148_;
  assign new_n1150_ = ~\priority[37]  & \req[36] ;
  assign new_n1151_ = ~\req[37]  & ~\req[38] ;
  assign new_n1152_ = ~new_n1150_ & new_n1151_;
  assign new_n1153_ = ~new_n1149_ & new_n1152_;
  assign new_n1154_ = \priority[38]  & ~\req[38] ;
  assign new_n1155_ = ~\priority[39]  & ~new_n1154_;
  assign new_n1156_ = ~\priority[40]  & new_n1155_;
  assign new_n1157_ = ~new_n1153_ & new_n1156_;
  assign new_n1158_ = ~\priority[40]  & \req[39] ;
  assign new_n1159_ = ~\req[40]  & ~\req[41] ;
  assign new_n1160_ = ~new_n1158_ & new_n1159_;
  assign new_n1161_ = ~new_n1157_ & new_n1160_;
  assign new_n1162_ = \priority[41]  & ~\req[41] ;
  assign new_n1163_ = ~\priority[42]  & ~new_n1162_;
  assign new_n1164_ = ~\priority[43]  & new_n1163_;
  assign new_n1165_ = ~new_n1161_ & new_n1164_;
  assign new_n1166_ = ~\priority[43]  & \req[42] ;
  assign new_n1167_ = ~\req[43]  & ~\req[44] ;
  assign new_n1168_ = ~new_n1166_ & new_n1167_;
  assign new_n1169_ = ~new_n1165_ & new_n1168_;
  assign new_n1170_ = \priority[44]  & ~\req[44] ;
  assign new_n1171_ = ~\priority[45]  & ~new_n1170_;
  assign new_n1172_ = ~\priority[46]  & new_n1171_;
  assign new_n1173_ = ~new_n1169_ & new_n1172_;
  assign new_n1174_ = ~\priority[46]  & \req[45] ;
  assign new_n1175_ = ~\req[46]  & ~\req[47] ;
  assign new_n1176_ = ~new_n1174_ & new_n1175_;
  assign new_n1177_ = ~new_n1173_ & new_n1176_;
  assign new_n1178_ = \priority[47]  & ~\req[47] ;
  assign new_n1179_ = ~\priority[48]  & ~new_n1178_;
  assign new_n1180_ = ~\priority[49]  & new_n1179_;
  assign new_n1181_ = ~new_n1177_ & new_n1180_;
  assign new_n1182_ = ~\priority[49]  & \req[48] ;
  assign new_n1183_ = ~\req[49]  & ~\req[50] ;
  assign new_n1184_ = ~new_n1182_ & new_n1183_;
  assign new_n1185_ = ~new_n1181_ & new_n1184_;
  assign new_n1186_ = \priority[50]  & ~\req[50] ;
  assign new_n1187_ = ~\priority[51]  & ~new_n1186_;
  assign new_n1188_ = ~\priority[52]  & new_n1187_;
  assign new_n1189_ = ~new_n1185_ & new_n1188_;
  assign new_n1190_ = ~\priority[52]  & \req[51] ;
  assign new_n1191_ = ~\req[52]  & ~\req[53] ;
  assign new_n1192_ = ~new_n1190_ & new_n1191_;
  assign new_n1193_ = ~new_n1189_ & new_n1192_;
  assign new_n1194_ = \priority[53]  & ~\req[53] ;
  assign new_n1195_ = ~\priority[54]  & ~new_n1194_;
  assign new_n1196_ = ~\priority[55]  & new_n1195_;
  assign new_n1197_ = ~new_n1193_ & new_n1196_;
  assign new_n1198_ = ~\priority[55]  & \req[54] ;
  assign new_n1199_ = ~\req[55]  & ~\req[56] ;
  assign new_n1200_ = ~new_n1198_ & new_n1199_;
  assign new_n1201_ = ~new_n1197_ & new_n1200_;
  assign new_n1202_ = \priority[56]  & ~\req[56] ;
  assign new_n1203_ = ~\priority[57]  & ~new_n1202_;
  assign new_n1204_ = ~\priority[58]  & new_n1203_;
  assign new_n1205_ = ~new_n1201_ & new_n1204_;
  assign new_n1206_ = ~\priority[58]  & \req[57] ;
  assign new_n1207_ = ~\req[58]  & ~\req[59] ;
  assign new_n1208_ = ~new_n1206_ & new_n1207_;
  assign new_n1209_ = ~new_n1205_ & new_n1208_;
  assign new_n1210_ = \priority[59]  & ~\req[59] ;
  assign new_n1211_ = ~\priority[60]  & ~new_n1210_;
  assign new_n1212_ = ~\priority[61]  & new_n1211_;
  assign new_n1213_ = ~new_n1209_ & new_n1212_;
  assign new_n1214_ = ~\priority[61]  & \req[60] ;
  assign new_n1215_ = ~\req[61]  & ~\req[62] ;
  assign new_n1216_ = ~new_n1214_ & new_n1215_;
  assign new_n1217_ = ~new_n1213_ & new_n1216_;
  assign new_n1218_ = \priority[62]  & ~\req[62] ;
  assign new_n1219_ = ~\priority[63]  & ~new_n1218_;
  assign new_n1220_ = ~\priority[64]  & new_n1219_;
  assign new_n1221_ = ~new_n1217_ & new_n1220_;
  assign new_n1222_ = ~\priority[64]  & \req[63] ;
  assign new_n1223_ = ~\req[64]  & ~\req[65] ;
  assign new_n1224_ = ~new_n1222_ & new_n1223_;
  assign new_n1225_ = ~new_n1221_ & new_n1224_;
  assign new_n1226_ = \priority[65]  & ~\req[65] ;
  assign new_n1227_ = ~\priority[66]  & ~new_n1226_;
  assign new_n1228_ = ~\priority[67]  & new_n1227_;
  assign new_n1229_ = ~new_n1225_ & new_n1228_;
  assign new_n1230_ = ~\priority[67]  & \req[66] ;
  assign new_n1231_ = ~\req[67]  & ~\req[68] ;
  assign new_n1232_ = ~new_n1230_ & new_n1231_;
  assign new_n1233_ = ~new_n1229_ & new_n1232_;
  assign new_n1234_ = \priority[68]  & ~\req[68] ;
  assign new_n1235_ = ~\priority[69]  & ~new_n1234_;
  assign new_n1236_ = ~\priority[70]  & new_n1235_;
  assign new_n1237_ = ~new_n1233_ & new_n1236_;
  assign new_n1238_ = ~\priority[70]  & \req[69] ;
  assign new_n1239_ = ~\req[70]  & ~\req[71] ;
  assign new_n1240_ = ~new_n1238_ & new_n1239_;
  assign new_n1241_ = ~new_n1237_ & new_n1240_;
  assign new_n1242_ = \priority[71]  & ~\req[71] ;
  assign new_n1243_ = ~\priority[72]  & ~new_n1242_;
  assign new_n1244_ = ~\priority[73]  & new_n1243_;
  assign new_n1245_ = ~new_n1241_ & new_n1244_;
  assign new_n1246_ = ~\priority[73]  & \req[72] ;
  assign new_n1247_ = ~\req[73]  & ~\req[74] ;
  assign new_n1248_ = ~new_n1246_ & new_n1247_;
  assign new_n1249_ = ~new_n1245_ & new_n1248_;
  assign new_n1250_ = \priority[74]  & ~\req[74] ;
  assign new_n1251_ = ~\priority[75]  & ~new_n1250_;
  assign new_n1252_ = ~\priority[76]  & new_n1251_;
  assign new_n1253_ = ~new_n1249_ & new_n1252_;
  assign new_n1254_ = ~\priority[76]  & \req[75] ;
  assign new_n1255_ = ~\req[76]  & ~\req[77] ;
  assign new_n1256_ = ~new_n1254_ & new_n1255_;
  assign new_n1257_ = ~new_n1253_ & new_n1256_;
  assign new_n1258_ = \priority[77]  & ~\req[77] ;
  assign new_n1259_ = ~\priority[78]  & ~new_n1258_;
  assign new_n1260_ = ~\priority[79]  & new_n1259_;
  assign new_n1261_ = ~new_n1257_ & new_n1260_;
  assign new_n1262_ = ~\priority[79]  & \req[78] ;
  assign new_n1263_ = ~\req[79]  & ~\req[80] ;
  assign new_n1264_ = ~new_n1262_ & new_n1263_;
  assign new_n1265_ = ~new_n1261_ & new_n1264_;
  assign new_n1266_ = \priority[80]  & ~\req[80] ;
  assign new_n1267_ = ~\priority[81]  & ~new_n1266_;
  assign new_n1268_ = ~\priority[82]  & new_n1267_;
  assign new_n1269_ = ~new_n1265_ & new_n1268_;
  assign new_n1270_ = ~\priority[82]  & \req[81] ;
  assign new_n1271_ = ~\req[82]  & ~\req[83] ;
  assign new_n1272_ = ~new_n1270_ & new_n1271_;
  assign new_n1273_ = ~new_n1269_ & new_n1272_;
  assign new_n1274_ = \priority[83]  & ~\req[83] ;
  assign new_n1275_ = ~\priority[84]  & ~new_n1274_;
  assign new_n1276_ = ~\priority[85]  & new_n1275_;
  assign new_n1277_ = ~new_n1273_ & new_n1276_;
  assign new_n1278_ = ~\priority[85]  & \req[84] ;
  assign new_n1279_ = ~\req[85]  & ~\req[86] ;
  assign new_n1280_ = ~new_n1278_ & new_n1279_;
  assign new_n1281_ = ~new_n1277_ & new_n1280_;
  assign new_n1282_ = \priority[86]  & ~\req[86] ;
  assign new_n1283_ = ~\priority[87]  & ~new_n1282_;
  assign new_n1284_ = ~\priority[88]  & new_n1283_;
  assign new_n1285_ = ~new_n1281_ & new_n1284_;
  assign new_n1286_ = ~\priority[88]  & \req[87] ;
  assign new_n1287_ = ~\req[88]  & ~\req[89] ;
  assign new_n1288_ = ~new_n1286_ & new_n1287_;
  assign new_n1289_ = ~new_n1285_ & new_n1288_;
  assign new_n1290_ = \priority[89]  & ~\req[89] ;
  assign new_n1291_ = ~\priority[90]  & ~new_n1290_;
  assign new_n1292_ = ~\priority[91]  & new_n1291_;
  assign new_n1293_ = ~new_n1289_ & new_n1292_;
  assign new_n1294_ = ~\priority[91]  & \req[90] ;
  assign new_n1295_ = ~\req[91]  & ~\req[92] ;
  assign new_n1296_ = ~new_n1294_ & new_n1295_;
  assign new_n1297_ = ~new_n1293_ & new_n1296_;
  assign new_n1298_ = \priority[92]  & ~\req[92] ;
  assign new_n1299_ = ~\priority[93]  & ~new_n1298_;
  assign new_n1300_ = ~\priority[94]  & new_n1299_;
  assign new_n1301_ = ~new_n1297_ & new_n1300_;
  assign new_n1302_ = ~\priority[94]  & \req[93] ;
  assign new_n1303_ = ~\req[94]  & ~\req[95] ;
  assign new_n1304_ = ~new_n1302_ & new_n1303_;
  assign new_n1305_ = ~new_n1301_ & new_n1304_;
  assign new_n1306_ = \priority[95]  & ~\req[95] ;
  assign new_n1307_ = ~\priority[96]  & ~new_n1306_;
  assign new_n1308_ = ~\priority[97]  & new_n1307_;
  assign new_n1309_ = ~new_n1305_ & new_n1308_;
  assign new_n1310_ = ~\priority[97]  & \req[96] ;
  assign new_n1311_ = ~\req[97]  & ~\req[98] ;
  assign new_n1312_ = ~new_n1310_ & new_n1311_;
  assign new_n1313_ = ~new_n1309_ & new_n1312_;
  assign new_n1314_ = \priority[98]  & ~\req[98] ;
  assign new_n1315_ = ~\priority[99]  & ~new_n1314_;
  assign new_n1316_ = ~\priority[100]  & new_n1315_;
  assign new_n1317_ = ~new_n1313_ & new_n1316_;
  assign new_n1318_ = ~\priority[100]  & \req[99] ;
  assign new_n1319_ = ~\req[100]  & ~\req[101] ;
  assign new_n1320_ = ~new_n1318_ & new_n1319_;
  assign new_n1321_ = ~new_n1317_ & new_n1320_;
  assign new_n1322_ = \priority[101]  & ~\req[101] ;
  assign new_n1323_ = ~\priority[102]  & ~new_n1322_;
  assign new_n1324_ = ~\priority[103]  & new_n1323_;
  assign new_n1325_ = ~new_n1321_ & new_n1324_;
  assign new_n1326_ = ~\priority[103]  & \req[102] ;
  assign new_n1327_ = ~\req[103]  & ~\req[104] ;
  assign new_n1328_ = ~new_n1326_ & new_n1327_;
  assign new_n1329_ = ~new_n1325_ & new_n1328_;
  assign new_n1330_ = \priority[104]  & ~\req[104] ;
  assign new_n1331_ = ~\priority[105]  & ~new_n1330_;
  assign new_n1332_ = ~\priority[106]  & new_n1331_;
  assign new_n1333_ = ~new_n1329_ & new_n1332_;
  assign new_n1334_ = ~\priority[106]  & \req[105] ;
  assign new_n1335_ = ~\req[106]  & ~\req[107] ;
  assign new_n1336_ = ~new_n1334_ & new_n1335_;
  assign new_n1337_ = ~new_n1333_ & new_n1336_;
  assign new_n1338_ = \priority[107]  & ~\req[107] ;
  assign new_n1339_ = ~\priority[108]  & ~new_n1338_;
  assign new_n1340_ = ~\priority[109]  & new_n1339_;
  assign new_n1341_ = ~new_n1337_ & new_n1340_;
  assign new_n1342_ = ~\priority[109]  & \req[108] ;
  assign new_n1343_ = ~\req[109]  & ~\req[110] ;
  assign new_n1344_ = ~new_n1342_ & new_n1343_;
  assign new_n1345_ = ~new_n1341_ & new_n1344_;
  assign new_n1346_ = \priority[110]  & ~\req[110] ;
  assign new_n1347_ = ~\priority[111]  & ~new_n1346_;
  assign new_n1348_ = ~\priority[112]  & new_n1347_;
  assign new_n1349_ = ~new_n1345_ & new_n1348_;
  assign new_n1350_ = ~\priority[112]  & \req[111] ;
  assign new_n1351_ = ~\req[112]  & ~\req[113] ;
  assign new_n1352_ = ~new_n1350_ & new_n1351_;
  assign new_n1353_ = ~new_n1349_ & new_n1352_;
  assign new_n1354_ = \priority[113]  & ~\req[113] ;
  assign new_n1355_ = ~\priority[114]  & ~new_n1354_;
  assign new_n1356_ = ~\priority[115]  & new_n1355_;
  assign new_n1357_ = ~new_n1353_ & new_n1356_;
  assign new_n1358_ = ~\priority[115]  & \req[114] ;
  assign new_n1359_ = ~\req[115]  & ~\req[116] ;
  assign new_n1360_ = ~new_n1358_ & new_n1359_;
  assign new_n1361_ = ~new_n1357_ & new_n1360_;
  assign new_n1362_ = \priority[116]  & ~\req[116] ;
  assign new_n1363_ = ~\priority[117]  & ~new_n1362_;
  assign new_n1364_ = ~\priority[118]  & new_n1363_;
  assign new_n1365_ = ~new_n1361_ & new_n1364_;
  assign new_n1366_ = ~\priority[118]  & \req[117] ;
  assign new_n1367_ = ~\req[118]  & ~\req[119] ;
  assign new_n1368_ = ~new_n1366_ & new_n1367_;
  assign new_n1369_ = ~new_n1365_ & new_n1368_;
  assign new_n1370_ = \priority[119]  & ~\req[119] ;
  assign new_n1371_ = ~\priority[120]  & ~new_n1370_;
  assign new_n1372_ = ~\priority[121]  & new_n1371_;
  assign new_n1373_ = ~new_n1369_ & new_n1372_;
  assign new_n1374_ = ~\priority[121]  & \req[120] ;
  assign new_n1375_ = ~\req[121]  & ~\req[122] ;
  assign new_n1376_ = ~new_n1374_ & new_n1375_;
  assign new_n1377_ = ~new_n1373_ & new_n1376_;
  assign new_n1378_ = \priority[122]  & ~\req[122] ;
  assign new_n1379_ = ~\priority[123]  & ~new_n1378_;
  assign new_n1380_ = ~\priority[124]  & new_n1379_;
  assign new_n1381_ = ~new_n1377_ & new_n1380_;
  assign new_n1382_ = ~\priority[124]  & \req[123] ;
  assign new_n1383_ = ~\req[124]  & ~\req[125] ;
  assign new_n1384_ = ~new_n1382_ & new_n1383_;
  assign new_n1385_ = ~new_n1381_ & new_n1384_;
  assign new_n1386_ = \priority[125]  & ~\req[125] ;
  assign new_n1387_ = ~\priority[126]  & ~new_n1386_;
  assign new_n1388_ = ~\priority[127]  & new_n1387_;
  assign new_n1389_ = ~new_n1385_ & new_n1388_;
  assign new_n1390_ = ~\priority[127]  & \req[126] ;
  assign new_n1391_ = ~\req[0]  & ~\req[127] ;
  assign new_n1392_ = ~new_n1390_ & new_n1391_;
  assign new_n1393_ = ~new_n1389_ & new_n1392_;
  assign new_n1394_ = \priority[0]  & ~\req[0] ;
  assign new_n1395_ = ~\priority[1]  & ~new_n1394_;
  assign new_n1396_ = ~\priority[2]  & new_n1395_;
  assign new_n1397_ = ~new_n1393_ & new_n1396_;
  assign new_n1398_ = ~\priority[2]  & \req[1] ;
  assign new_n1399_ = \req[2]  & ~new_n1398_;
  assign \grant[2]  = ~new_n1397_ & new_n1399_;
  assign new_n1401_ = new_n395_ & ~new_n730_;
  assign new_n1402_ = new_n400_ & ~new_n1401_;
  assign new_n1403_ = new_n404_ & ~new_n1402_;
  assign new_n1404_ = new_n408_ & ~new_n1403_;
  assign new_n1405_ = new_n412_ & ~new_n1404_;
  assign new_n1406_ = new_n416_ & ~new_n1405_;
  assign new_n1407_ = new_n420_ & ~new_n1406_;
  assign new_n1408_ = new_n424_ & ~new_n1407_;
  assign new_n1409_ = new_n428_ & ~new_n1408_;
  assign new_n1410_ = new_n432_ & ~new_n1409_;
  assign new_n1411_ = new_n436_ & ~new_n1410_;
  assign new_n1412_ = new_n440_ & ~new_n1411_;
  assign new_n1413_ = new_n444_ & ~new_n1412_;
  assign new_n1414_ = new_n448_ & ~new_n1413_;
  assign new_n1415_ = new_n452_ & ~new_n1414_;
  assign new_n1416_ = new_n456_ & ~new_n1415_;
  assign new_n1417_ = new_n460_ & ~new_n1416_;
  assign new_n1418_ = new_n464_ & ~new_n1417_;
  assign new_n1419_ = new_n468_ & ~new_n1418_;
  assign new_n1420_ = new_n472_ & ~new_n1419_;
  assign new_n1421_ = new_n476_ & ~new_n1420_;
  assign new_n1422_ = new_n480_ & ~new_n1421_;
  assign new_n1423_ = new_n484_ & ~new_n1422_;
  assign new_n1424_ = new_n488_ & ~new_n1423_;
  assign new_n1425_ = new_n492_ & ~new_n1424_;
  assign new_n1426_ = new_n496_ & ~new_n1425_;
  assign new_n1427_ = new_n500_ & ~new_n1426_;
  assign new_n1428_ = new_n504_ & ~new_n1427_;
  assign new_n1429_ = new_n508_ & ~new_n1428_;
  assign new_n1430_ = new_n512_ & ~new_n1429_;
  assign new_n1431_ = new_n516_ & ~new_n1430_;
  assign new_n1432_ = new_n520_ & ~new_n1431_;
  assign new_n1433_ = new_n524_ & ~new_n1432_;
  assign new_n1434_ = new_n528_ & ~new_n1433_;
  assign new_n1435_ = new_n532_ & ~new_n1434_;
  assign new_n1436_ = new_n536_ & ~new_n1435_;
  assign new_n1437_ = new_n540_ & ~new_n1436_;
  assign new_n1438_ = new_n544_ & ~new_n1437_;
  assign new_n1439_ = new_n548_ & ~new_n1438_;
  assign new_n1440_ = new_n552_ & ~new_n1439_;
  assign new_n1441_ = new_n556_ & ~new_n1440_;
  assign new_n1442_ = new_n560_ & ~new_n1441_;
  assign new_n1443_ = new_n564_ & ~new_n1442_;
  assign new_n1444_ = new_n568_ & ~new_n1443_;
  assign new_n1445_ = new_n572_ & ~new_n1444_;
  assign new_n1446_ = new_n576_ & ~new_n1445_;
  assign new_n1447_ = new_n580_ & ~new_n1446_;
  assign new_n1448_ = new_n584_ & ~new_n1447_;
  assign new_n1449_ = new_n588_ & ~new_n1448_;
  assign new_n1450_ = new_n592_ & ~new_n1449_;
  assign new_n1451_ = new_n596_ & ~new_n1450_;
  assign new_n1452_ = new_n600_ & ~new_n1451_;
  assign new_n1453_ = new_n604_ & ~new_n1452_;
  assign new_n1454_ = new_n608_ & ~new_n1453_;
  assign new_n1455_ = new_n612_ & ~new_n1454_;
  assign new_n1456_ = new_n616_ & ~new_n1455_;
  assign new_n1457_ = new_n620_ & ~new_n1456_;
  assign new_n1458_ = new_n624_ & ~new_n1457_;
  assign new_n1459_ = new_n628_ & ~new_n1458_;
  assign new_n1460_ = new_n632_ & ~new_n1459_;
  assign new_n1461_ = new_n636_ & ~new_n1460_;
  assign new_n1462_ = new_n640_ & ~new_n1461_;
  assign new_n1463_ = new_n644_ & ~new_n1462_;
  assign new_n1464_ = new_n648_ & ~new_n1463_;
  assign new_n1465_ = new_n652_ & ~new_n1464_;
  assign new_n1466_ = new_n656_ & ~new_n1465_;
  assign new_n1467_ = new_n660_ & ~new_n1466_;
  assign new_n1468_ = new_n664_ & ~new_n1467_;
  assign new_n1469_ = new_n668_ & ~new_n1468_;
  assign new_n1470_ = new_n672_ & ~new_n1469_;
  assign new_n1471_ = new_n676_ & ~new_n1470_;
  assign new_n1472_ = new_n680_ & ~new_n1471_;
  assign new_n1473_ = new_n684_ & ~new_n1472_;
  assign new_n1474_ = new_n688_ & ~new_n1473_;
  assign new_n1475_ = new_n692_ & ~new_n1474_;
  assign new_n1476_ = new_n696_ & ~new_n1475_;
  assign new_n1477_ = new_n700_ & ~new_n1476_;
  assign new_n1478_ = new_n704_ & ~new_n1477_;
  assign new_n1479_ = new_n708_ & ~new_n1478_;
  assign new_n1480_ = new_n712_ & ~new_n1479_;
  assign new_n1481_ = new_n716_ & ~new_n1480_;
  assign new_n1482_ = new_n720_ & ~new_n1481_;
  assign new_n1483_ = ~\req[0]  & ~\req[1] ;
  assign new_n1484_ = ~new_n722_ & new_n1483_;
  assign new_n1485_ = ~new_n1482_ & new_n1484_;
  assign new_n1486_ = ~\priority[3]  & new_n387_;
  assign new_n1487_ = ~new_n1485_ & new_n1486_;
  assign new_n1488_ = ~\priority[3]  & \req[2] ;
  assign new_n1489_ = \req[3]  & ~new_n1488_;
  assign \grant[3]  = ~new_n1487_ & new_n1489_;
  assign new_n1491_ = new_n734_ & ~new_n1067_;
  assign new_n1492_ = new_n739_ & ~new_n1491_;
  assign new_n1493_ = new_n743_ & ~new_n1492_;
  assign new_n1494_ = new_n747_ & ~new_n1493_;
  assign new_n1495_ = new_n751_ & ~new_n1494_;
  assign new_n1496_ = new_n755_ & ~new_n1495_;
  assign new_n1497_ = new_n759_ & ~new_n1496_;
  assign new_n1498_ = new_n763_ & ~new_n1497_;
  assign new_n1499_ = new_n767_ & ~new_n1498_;
  assign new_n1500_ = new_n771_ & ~new_n1499_;
  assign new_n1501_ = new_n775_ & ~new_n1500_;
  assign new_n1502_ = new_n779_ & ~new_n1501_;
  assign new_n1503_ = new_n783_ & ~new_n1502_;
  assign new_n1504_ = new_n787_ & ~new_n1503_;
  assign new_n1505_ = new_n791_ & ~new_n1504_;
  assign new_n1506_ = new_n795_ & ~new_n1505_;
  assign new_n1507_ = new_n799_ & ~new_n1506_;
  assign new_n1508_ = new_n803_ & ~new_n1507_;
  assign new_n1509_ = new_n807_ & ~new_n1508_;
  assign new_n1510_ = new_n811_ & ~new_n1509_;
  assign new_n1511_ = new_n815_ & ~new_n1510_;
  assign new_n1512_ = new_n819_ & ~new_n1511_;
  assign new_n1513_ = new_n823_ & ~new_n1512_;
  assign new_n1514_ = new_n827_ & ~new_n1513_;
  assign new_n1515_ = new_n831_ & ~new_n1514_;
  assign new_n1516_ = new_n835_ & ~new_n1515_;
  assign new_n1517_ = new_n839_ & ~new_n1516_;
  assign new_n1518_ = new_n843_ & ~new_n1517_;
  assign new_n1519_ = new_n847_ & ~new_n1518_;
  assign new_n1520_ = new_n851_ & ~new_n1519_;
  assign new_n1521_ = new_n855_ & ~new_n1520_;
  assign new_n1522_ = new_n859_ & ~new_n1521_;
  assign new_n1523_ = new_n863_ & ~new_n1522_;
  assign new_n1524_ = new_n867_ & ~new_n1523_;
  assign new_n1525_ = new_n871_ & ~new_n1524_;
  assign new_n1526_ = new_n875_ & ~new_n1525_;
  assign new_n1527_ = new_n879_ & ~new_n1526_;
  assign new_n1528_ = new_n883_ & ~new_n1527_;
  assign new_n1529_ = new_n887_ & ~new_n1528_;
  assign new_n1530_ = new_n891_ & ~new_n1529_;
  assign new_n1531_ = new_n895_ & ~new_n1530_;
  assign new_n1532_ = new_n899_ & ~new_n1531_;
  assign new_n1533_ = new_n903_ & ~new_n1532_;
  assign new_n1534_ = new_n907_ & ~new_n1533_;
  assign new_n1535_ = new_n911_ & ~new_n1534_;
  assign new_n1536_ = new_n915_ & ~new_n1535_;
  assign new_n1537_ = new_n919_ & ~new_n1536_;
  assign new_n1538_ = new_n923_ & ~new_n1537_;
  assign new_n1539_ = new_n927_ & ~new_n1538_;
  assign new_n1540_ = new_n931_ & ~new_n1539_;
  assign new_n1541_ = new_n935_ & ~new_n1540_;
  assign new_n1542_ = new_n939_ & ~new_n1541_;
  assign new_n1543_ = new_n943_ & ~new_n1542_;
  assign new_n1544_ = new_n947_ & ~new_n1543_;
  assign new_n1545_ = new_n951_ & ~new_n1544_;
  assign new_n1546_ = new_n955_ & ~new_n1545_;
  assign new_n1547_ = new_n959_ & ~new_n1546_;
  assign new_n1548_ = new_n963_ & ~new_n1547_;
  assign new_n1549_ = new_n967_ & ~new_n1548_;
  assign new_n1550_ = new_n971_ & ~new_n1549_;
  assign new_n1551_ = new_n975_ & ~new_n1550_;
  assign new_n1552_ = new_n979_ & ~new_n1551_;
  assign new_n1553_ = new_n983_ & ~new_n1552_;
  assign new_n1554_ = new_n987_ & ~new_n1553_;
  assign new_n1555_ = new_n991_ & ~new_n1554_;
  assign new_n1556_ = new_n995_ & ~new_n1555_;
  assign new_n1557_ = new_n999_ & ~new_n1556_;
  assign new_n1558_ = new_n1003_ & ~new_n1557_;
  assign new_n1559_ = new_n1007_ & ~new_n1558_;
  assign new_n1560_ = new_n1011_ & ~new_n1559_;
  assign new_n1561_ = new_n1015_ & ~new_n1560_;
  assign new_n1562_ = new_n1019_ & ~new_n1561_;
  assign new_n1563_ = new_n1023_ & ~new_n1562_;
  assign new_n1564_ = new_n1027_ & ~new_n1563_;
  assign new_n1565_ = new_n1031_ & ~new_n1564_;
  assign new_n1566_ = new_n1035_ & ~new_n1565_;
  assign new_n1567_ = new_n1039_ & ~new_n1566_;
  assign new_n1568_ = new_n1043_ & ~new_n1567_;
  assign new_n1569_ = new_n1047_ & ~new_n1568_;
  assign new_n1570_ = new_n1051_ & ~new_n1569_;
  assign new_n1571_ = new_n1055_ & ~new_n1570_;
  assign new_n1572_ = new_n1059_ & ~new_n1571_;
  assign new_n1573_ = ~\req[1]  & ~\req[2] ;
  assign new_n1574_ = ~new_n1061_ & new_n1573_;
  assign new_n1575_ = ~new_n1572_ & new_n1574_;
  assign new_n1576_ = ~\priority[4]  & new_n726_;
  assign new_n1577_ = ~new_n1575_ & new_n1576_;
  assign new_n1578_ = ~\priority[4]  & \req[3] ;
  assign new_n1579_ = \req[4]  & ~new_n1578_;
  assign \grant[4]  = ~new_n1577_ & new_n1579_;
  assign new_n1581_ = ~new_n399_ & new_n1071_;
  assign new_n1582_ = new_n1076_ & ~new_n1581_;
  assign new_n1583_ = new_n1080_ & ~new_n1582_;
  assign new_n1584_ = new_n1084_ & ~new_n1583_;
  assign new_n1585_ = new_n1088_ & ~new_n1584_;
  assign new_n1586_ = new_n1092_ & ~new_n1585_;
  assign new_n1587_ = new_n1096_ & ~new_n1586_;
  assign new_n1588_ = new_n1100_ & ~new_n1587_;
  assign new_n1589_ = new_n1104_ & ~new_n1588_;
  assign new_n1590_ = new_n1108_ & ~new_n1589_;
  assign new_n1591_ = new_n1112_ & ~new_n1590_;
  assign new_n1592_ = new_n1116_ & ~new_n1591_;
  assign new_n1593_ = new_n1120_ & ~new_n1592_;
  assign new_n1594_ = new_n1124_ & ~new_n1593_;
  assign new_n1595_ = new_n1128_ & ~new_n1594_;
  assign new_n1596_ = new_n1132_ & ~new_n1595_;
  assign new_n1597_ = new_n1136_ & ~new_n1596_;
  assign new_n1598_ = new_n1140_ & ~new_n1597_;
  assign new_n1599_ = new_n1144_ & ~new_n1598_;
  assign new_n1600_ = new_n1148_ & ~new_n1599_;
  assign new_n1601_ = new_n1152_ & ~new_n1600_;
  assign new_n1602_ = new_n1156_ & ~new_n1601_;
  assign new_n1603_ = new_n1160_ & ~new_n1602_;
  assign new_n1604_ = new_n1164_ & ~new_n1603_;
  assign new_n1605_ = new_n1168_ & ~new_n1604_;
  assign new_n1606_ = new_n1172_ & ~new_n1605_;
  assign new_n1607_ = new_n1176_ & ~new_n1606_;
  assign new_n1608_ = new_n1180_ & ~new_n1607_;
  assign new_n1609_ = new_n1184_ & ~new_n1608_;
  assign new_n1610_ = new_n1188_ & ~new_n1609_;
  assign new_n1611_ = new_n1192_ & ~new_n1610_;
  assign new_n1612_ = new_n1196_ & ~new_n1611_;
  assign new_n1613_ = new_n1200_ & ~new_n1612_;
  assign new_n1614_ = new_n1204_ & ~new_n1613_;
  assign new_n1615_ = new_n1208_ & ~new_n1614_;
  assign new_n1616_ = new_n1212_ & ~new_n1615_;
  assign new_n1617_ = new_n1216_ & ~new_n1616_;
  assign new_n1618_ = new_n1220_ & ~new_n1617_;
  assign new_n1619_ = new_n1224_ & ~new_n1618_;
  assign new_n1620_ = new_n1228_ & ~new_n1619_;
  assign new_n1621_ = new_n1232_ & ~new_n1620_;
  assign new_n1622_ = new_n1236_ & ~new_n1621_;
  assign new_n1623_ = new_n1240_ & ~new_n1622_;
  assign new_n1624_ = new_n1244_ & ~new_n1623_;
  assign new_n1625_ = new_n1248_ & ~new_n1624_;
  assign new_n1626_ = new_n1252_ & ~new_n1625_;
  assign new_n1627_ = new_n1256_ & ~new_n1626_;
  assign new_n1628_ = new_n1260_ & ~new_n1627_;
  assign new_n1629_ = new_n1264_ & ~new_n1628_;
  assign new_n1630_ = new_n1268_ & ~new_n1629_;
  assign new_n1631_ = new_n1272_ & ~new_n1630_;
  assign new_n1632_ = new_n1276_ & ~new_n1631_;
  assign new_n1633_ = new_n1280_ & ~new_n1632_;
  assign new_n1634_ = new_n1284_ & ~new_n1633_;
  assign new_n1635_ = new_n1288_ & ~new_n1634_;
  assign new_n1636_ = new_n1292_ & ~new_n1635_;
  assign new_n1637_ = new_n1296_ & ~new_n1636_;
  assign new_n1638_ = new_n1300_ & ~new_n1637_;
  assign new_n1639_ = new_n1304_ & ~new_n1638_;
  assign new_n1640_ = new_n1308_ & ~new_n1639_;
  assign new_n1641_ = new_n1312_ & ~new_n1640_;
  assign new_n1642_ = new_n1316_ & ~new_n1641_;
  assign new_n1643_ = new_n1320_ & ~new_n1642_;
  assign new_n1644_ = new_n1324_ & ~new_n1643_;
  assign new_n1645_ = new_n1328_ & ~new_n1644_;
  assign new_n1646_ = new_n1332_ & ~new_n1645_;
  assign new_n1647_ = new_n1336_ & ~new_n1646_;
  assign new_n1648_ = new_n1340_ & ~new_n1647_;
  assign new_n1649_ = new_n1344_ & ~new_n1648_;
  assign new_n1650_ = new_n1348_ & ~new_n1649_;
  assign new_n1651_ = new_n1352_ & ~new_n1650_;
  assign new_n1652_ = new_n1356_ & ~new_n1651_;
  assign new_n1653_ = new_n1360_ & ~new_n1652_;
  assign new_n1654_ = new_n1364_ & ~new_n1653_;
  assign new_n1655_ = new_n1368_ & ~new_n1654_;
  assign new_n1656_ = new_n1372_ & ~new_n1655_;
  assign new_n1657_ = new_n1376_ & ~new_n1656_;
  assign new_n1658_ = new_n1380_ & ~new_n1657_;
  assign new_n1659_ = new_n1384_ & ~new_n1658_;
  assign new_n1660_ = new_n1388_ & ~new_n1659_;
  assign new_n1661_ = new_n1392_ & ~new_n1660_;
  assign new_n1662_ = new_n1396_ & ~new_n1661_;
  assign new_n1663_ = new_n388_ & ~new_n1398_;
  assign new_n1664_ = ~new_n1662_ & new_n1663_;
  assign new_n1665_ = new_n392_ & ~new_n1664_;
  assign new_n1666_ = \req[5]  & ~new_n394_;
  assign \grant[5]  = ~new_n1665_ & new_n1666_;
  assign new_n1668_ = new_n403_ & ~new_n738_;
  assign new_n1669_ = new_n408_ & ~new_n1668_;
  assign new_n1670_ = new_n412_ & ~new_n1669_;
  assign new_n1671_ = new_n416_ & ~new_n1670_;
  assign new_n1672_ = new_n420_ & ~new_n1671_;
  assign new_n1673_ = new_n424_ & ~new_n1672_;
  assign new_n1674_ = new_n428_ & ~new_n1673_;
  assign new_n1675_ = new_n432_ & ~new_n1674_;
  assign new_n1676_ = new_n436_ & ~new_n1675_;
  assign new_n1677_ = new_n440_ & ~new_n1676_;
  assign new_n1678_ = new_n444_ & ~new_n1677_;
  assign new_n1679_ = new_n448_ & ~new_n1678_;
  assign new_n1680_ = new_n452_ & ~new_n1679_;
  assign new_n1681_ = new_n456_ & ~new_n1680_;
  assign new_n1682_ = new_n460_ & ~new_n1681_;
  assign new_n1683_ = new_n464_ & ~new_n1682_;
  assign new_n1684_ = new_n468_ & ~new_n1683_;
  assign new_n1685_ = new_n472_ & ~new_n1684_;
  assign new_n1686_ = new_n476_ & ~new_n1685_;
  assign new_n1687_ = new_n480_ & ~new_n1686_;
  assign new_n1688_ = new_n484_ & ~new_n1687_;
  assign new_n1689_ = new_n488_ & ~new_n1688_;
  assign new_n1690_ = new_n492_ & ~new_n1689_;
  assign new_n1691_ = new_n496_ & ~new_n1690_;
  assign new_n1692_ = new_n500_ & ~new_n1691_;
  assign new_n1693_ = new_n504_ & ~new_n1692_;
  assign new_n1694_ = new_n508_ & ~new_n1693_;
  assign new_n1695_ = new_n512_ & ~new_n1694_;
  assign new_n1696_ = new_n516_ & ~new_n1695_;
  assign new_n1697_ = new_n520_ & ~new_n1696_;
  assign new_n1698_ = new_n524_ & ~new_n1697_;
  assign new_n1699_ = new_n528_ & ~new_n1698_;
  assign new_n1700_ = new_n532_ & ~new_n1699_;
  assign new_n1701_ = new_n536_ & ~new_n1700_;
  assign new_n1702_ = new_n540_ & ~new_n1701_;
  assign new_n1703_ = new_n544_ & ~new_n1702_;
  assign new_n1704_ = new_n548_ & ~new_n1703_;
  assign new_n1705_ = new_n552_ & ~new_n1704_;
  assign new_n1706_ = new_n556_ & ~new_n1705_;
  assign new_n1707_ = new_n560_ & ~new_n1706_;
  assign new_n1708_ = new_n564_ & ~new_n1707_;
  assign new_n1709_ = new_n568_ & ~new_n1708_;
  assign new_n1710_ = new_n572_ & ~new_n1709_;
  assign new_n1711_ = new_n576_ & ~new_n1710_;
  assign new_n1712_ = new_n580_ & ~new_n1711_;
  assign new_n1713_ = new_n584_ & ~new_n1712_;
  assign new_n1714_ = new_n588_ & ~new_n1713_;
  assign new_n1715_ = new_n592_ & ~new_n1714_;
  assign new_n1716_ = new_n596_ & ~new_n1715_;
  assign new_n1717_ = new_n600_ & ~new_n1716_;
  assign new_n1718_ = new_n604_ & ~new_n1717_;
  assign new_n1719_ = new_n608_ & ~new_n1718_;
  assign new_n1720_ = new_n612_ & ~new_n1719_;
  assign new_n1721_ = new_n616_ & ~new_n1720_;
  assign new_n1722_ = new_n620_ & ~new_n1721_;
  assign new_n1723_ = new_n624_ & ~new_n1722_;
  assign new_n1724_ = new_n628_ & ~new_n1723_;
  assign new_n1725_ = new_n632_ & ~new_n1724_;
  assign new_n1726_ = new_n636_ & ~new_n1725_;
  assign new_n1727_ = new_n640_ & ~new_n1726_;
  assign new_n1728_ = new_n644_ & ~new_n1727_;
  assign new_n1729_ = new_n648_ & ~new_n1728_;
  assign new_n1730_ = new_n652_ & ~new_n1729_;
  assign new_n1731_ = new_n656_ & ~new_n1730_;
  assign new_n1732_ = new_n660_ & ~new_n1731_;
  assign new_n1733_ = new_n664_ & ~new_n1732_;
  assign new_n1734_ = new_n668_ & ~new_n1733_;
  assign new_n1735_ = new_n672_ & ~new_n1734_;
  assign new_n1736_ = new_n676_ & ~new_n1735_;
  assign new_n1737_ = new_n680_ & ~new_n1736_;
  assign new_n1738_ = new_n684_ & ~new_n1737_;
  assign new_n1739_ = new_n688_ & ~new_n1738_;
  assign new_n1740_ = new_n692_ & ~new_n1739_;
  assign new_n1741_ = new_n696_ & ~new_n1740_;
  assign new_n1742_ = new_n700_ & ~new_n1741_;
  assign new_n1743_ = new_n704_ & ~new_n1742_;
  assign new_n1744_ = new_n708_ & ~new_n1743_;
  assign new_n1745_ = new_n712_ & ~new_n1744_;
  assign new_n1746_ = new_n716_ & ~new_n1745_;
  assign new_n1747_ = new_n720_ & ~new_n1746_;
  assign new_n1748_ = new_n1484_ & ~new_n1747_;
  assign new_n1749_ = new_n1486_ & ~new_n1748_;
  assign new_n1750_ = new_n727_ & ~new_n1488_;
  assign new_n1751_ = ~new_n1749_ & new_n1750_;
  assign new_n1752_ = new_n731_ & ~new_n1751_;
  assign new_n1753_ = \req[6]  & ~new_n733_;
  assign \grant[6]  = ~new_n1752_ & new_n1753_;
  assign new_n1755_ = new_n742_ & ~new_n1075_;
  assign new_n1756_ = new_n747_ & ~new_n1755_;
  assign new_n1757_ = new_n751_ & ~new_n1756_;
  assign new_n1758_ = new_n755_ & ~new_n1757_;
  assign new_n1759_ = new_n759_ & ~new_n1758_;
  assign new_n1760_ = new_n763_ & ~new_n1759_;
  assign new_n1761_ = new_n767_ & ~new_n1760_;
  assign new_n1762_ = new_n771_ & ~new_n1761_;
  assign new_n1763_ = new_n775_ & ~new_n1762_;
  assign new_n1764_ = new_n779_ & ~new_n1763_;
  assign new_n1765_ = new_n783_ & ~new_n1764_;
  assign new_n1766_ = new_n787_ & ~new_n1765_;
  assign new_n1767_ = new_n791_ & ~new_n1766_;
  assign new_n1768_ = new_n795_ & ~new_n1767_;
  assign new_n1769_ = new_n799_ & ~new_n1768_;
  assign new_n1770_ = new_n803_ & ~new_n1769_;
  assign new_n1771_ = new_n807_ & ~new_n1770_;
  assign new_n1772_ = new_n811_ & ~new_n1771_;
  assign new_n1773_ = new_n815_ & ~new_n1772_;
  assign new_n1774_ = new_n819_ & ~new_n1773_;
  assign new_n1775_ = new_n823_ & ~new_n1774_;
  assign new_n1776_ = new_n827_ & ~new_n1775_;
  assign new_n1777_ = new_n831_ & ~new_n1776_;
  assign new_n1778_ = new_n835_ & ~new_n1777_;
  assign new_n1779_ = new_n839_ & ~new_n1778_;
  assign new_n1780_ = new_n843_ & ~new_n1779_;
  assign new_n1781_ = new_n847_ & ~new_n1780_;
  assign new_n1782_ = new_n851_ & ~new_n1781_;
  assign new_n1783_ = new_n855_ & ~new_n1782_;
  assign new_n1784_ = new_n859_ & ~new_n1783_;
  assign new_n1785_ = new_n863_ & ~new_n1784_;
  assign new_n1786_ = new_n867_ & ~new_n1785_;
  assign new_n1787_ = new_n871_ & ~new_n1786_;
  assign new_n1788_ = new_n875_ & ~new_n1787_;
  assign new_n1789_ = new_n879_ & ~new_n1788_;
  assign new_n1790_ = new_n883_ & ~new_n1789_;
  assign new_n1791_ = new_n887_ & ~new_n1790_;
  assign new_n1792_ = new_n891_ & ~new_n1791_;
  assign new_n1793_ = new_n895_ & ~new_n1792_;
  assign new_n1794_ = new_n899_ & ~new_n1793_;
  assign new_n1795_ = new_n903_ & ~new_n1794_;
  assign new_n1796_ = new_n907_ & ~new_n1795_;
  assign new_n1797_ = new_n911_ & ~new_n1796_;
  assign new_n1798_ = new_n915_ & ~new_n1797_;
  assign new_n1799_ = new_n919_ & ~new_n1798_;
  assign new_n1800_ = new_n923_ & ~new_n1799_;
  assign new_n1801_ = new_n927_ & ~new_n1800_;
  assign new_n1802_ = new_n931_ & ~new_n1801_;
  assign new_n1803_ = new_n935_ & ~new_n1802_;
  assign new_n1804_ = new_n939_ & ~new_n1803_;
  assign new_n1805_ = new_n943_ & ~new_n1804_;
  assign new_n1806_ = new_n947_ & ~new_n1805_;
  assign new_n1807_ = new_n951_ & ~new_n1806_;
  assign new_n1808_ = new_n955_ & ~new_n1807_;
  assign new_n1809_ = new_n959_ & ~new_n1808_;
  assign new_n1810_ = new_n963_ & ~new_n1809_;
  assign new_n1811_ = new_n967_ & ~new_n1810_;
  assign new_n1812_ = new_n971_ & ~new_n1811_;
  assign new_n1813_ = new_n975_ & ~new_n1812_;
  assign new_n1814_ = new_n979_ & ~new_n1813_;
  assign new_n1815_ = new_n983_ & ~new_n1814_;
  assign new_n1816_ = new_n987_ & ~new_n1815_;
  assign new_n1817_ = new_n991_ & ~new_n1816_;
  assign new_n1818_ = new_n995_ & ~new_n1817_;
  assign new_n1819_ = new_n999_ & ~new_n1818_;
  assign new_n1820_ = new_n1003_ & ~new_n1819_;
  assign new_n1821_ = new_n1007_ & ~new_n1820_;
  assign new_n1822_ = new_n1011_ & ~new_n1821_;
  assign new_n1823_ = new_n1015_ & ~new_n1822_;
  assign new_n1824_ = new_n1019_ & ~new_n1823_;
  assign new_n1825_ = new_n1023_ & ~new_n1824_;
  assign new_n1826_ = new_n1027_ & ~new_n1825_;
  assign new_n1827_ = new_n1031_ & ~new_n1826_;
  assign new_n1828_ = new_n1035_ & ~new_n1827_;
  assign new_n1829_ = new_n1039_ & ~new_n1828_;
  assign new_n1830_ = new_n1043_ & ~new_n1829_;
  assign new_n1831_ = new_n1047_ & ~new_n1830_;
  assign new_n1832_ = new_n1051_ & ~new_n1831_;
  assign new_n1833_ = new_n1055_ & ~new_n1832_;
  assign new_n1834_ = new_n1059_ & ~new_n1833_;
  assign new_n1835_ = new_n1574_ & ~new_n1834_;
  assign new_n1836_ = new_n1576_ & ~new_n1835_;
  assign new_n1837_ = new_n1064_ & ~new_n1578_;
  assign new_n1838_ = ~new_n1836_ & new_n1837_;
  assign new_n1839_ = new_n1068_ & ~new_n1838_;
  assign new_n1840_ = \req[7]  & ~new_n1070_;
  assign \grant[7]  = ~new_n1839_ & new_n1840_;
  assign new_n1842_ = ~new_n407_ & new_n1079_;
  assign new_n1843_ = new_n1084_ & ~new_n1842_;
  assign new_n1844_ = new_n1088_ & ~new_n1843_;
  assign new_n1845_ = new_n1092_ & ~new_n1844_;
  assign new_n1846_ = new_n1096_ & ~new_n1845_;
  assign new_n1847_ = new_n1100_ & ~new_n1846_;
  assign new_n1848_ = new_n1104_ & ~new_n1847_;
  assign new_n1849_ = new_n1108_ & ~new_n1848_;
  assign new_n1850_ = new_n1112_ & ~new_n1849_;
  assign new_n1851_ = new_n1116_ & ~new_n1850_;
  assign new_n1852_ = new_n1120_ & ~new_n1851_;
  assign new_n1853_ = new_n1124_ & ~new_n1852_;
  assign new_n1854_ = new_n1128_ & ~new_n1853_;
  assign new_n1855_ = new_n1132_ & ~new_n1854_;
  assign new_n1856_ = new_n1136_ & ~new_n1855_;
  assign new_n1857_ = new_n1140_ & ~new_n1856_;
  assign new_n1858_ = new_n1144_ & ~new_n1857_;
  assign new_n1859_ = new_n1148_ & ~new_n1858_;
  assign new_n1860_ = new_n1152_ & ~new_n1859_;
  assign new_n1861_ = new_n1156_ & ~new_n1860_;
  assign new_n1862_ = new_n1160_ & ~new_n1861_;
  assign new_n1863_ = new_n1164_ & ~new_n1862_;
  assign new_n1864_ = new_n1168_ & ~new_n1863_;
  assign new_n1865_ = new_n1172_ & ~new_n1864_;
  assign new_n1866_ = new_n1176_ & ~new_n1865_;
  assign new_n1867_ = new_n1180_ & ~new_n1866_;
  assign new_n1868_ = new_n1184_ & ~new_n1867_;
  assign new_n1869_ = new_n1188_ & ~new_n1868_;
  assign new_n1870_ = new_n1192_ & ~new_n1869_;
  assign new_n1871_ = new_n1196_ & ~new_n1870_;
  assign new_n1872_ = new_n1200_ & ~new_n1871_;
  assign new_n1873_ = new_n1204_ & ~new_n1872_;
  assign new_n1874_ = new_n1208_ & ~new_n1873_;
  assign new_n1875_ = new_n1212_ & ~new_n1874_;
  assign new_n1876_ = new_n1216_ & ~new_n1875_;
  assign new_n1877_ = new_n1220_ & ~new_n1876_;
  assign new_n1878_ = new_n1224_ & ~new_n1877_;
  assign new_n1879_ = new_n1228_ & ~new_n1878_;
  assign new_n1880_ = new_n1232_ & ~new_n1879_;
  assign new_n1881_ = new_n1236_ & ~new_n1880_;
  assign new_n1882_ = new_n1240_ & ~new_n1881_;
  assign new_n1883_ = new_n1244_ & ~new_n1882_;
  assign new_n1884_ = new_n1248_ & ~new_n1883_;
  assign new_n1885_ = new_n1252_ & ~new_n1884_;
  assign new_n1886_ = new_n1256_ & ~new_n1885_;
  assign new_n1887_ = new_n1260_ & ~new_n1886_;
  assign new_n1888_ = new_n1264_ & ~new_n1887_;
  assign new_n1889_ = new_n1268_ & ~new_n1888_;
  assign new_n1890_ = new_n1272_ & ~new_n1889_;
  assign new_n1891_ = new_n1276_ & ~new_n1890_;
  assign new_n1892_ = new_n1280_ & ~new_n1891_;
  assign new_n1893_ = new_n1284_ & ~new_n1892_;
  assign new_n1894_ = new_n1288_ & ~new_n1893_;
  assign new_n1895_ = new_n1292_ & ~new_n1894_;
  assign new_n1896_ = new_n1296_ & ~new_n1895_;
  assign new_n1897_ = new_n1300_ & ~new_n1896_;
  assign new_n1898_ = new_n1304_ & ~new_n1897_;
  assign new_n1899_ = new_n1308_ & ~new_n1898_;
  assign new_n1900_ = new_n1312_ & ~new_n1899_;
  assign new_n1901_ = new_n1316_ & ~new_n1900_;
  assign new_n1902_ = new_n1320_ & ~new_n1901_;
  assign new_n1903_ = new_n1324_ & ~new_n1902_;
  assign new_n1904_ = new_n1328_ & ~new_n1903_;
  assign new_n1905_ = new_n1332_ & ~new_n1904_;
  assign new_n1906_ = new_n1336_ & ~new_n1905_;
  assign new_n1907_ = new_n1340_ & ~new_n1906_;
  assign new_n1908_ = new_n1344_ & ~new_n1907_;
  assign new_n1909_ = new_n1348_ & ~new_n1908_;
  assign new_n1910_ = new_n1352_ & ~new_n1909_;
  assign new_n1911_ = new_n1356_ & ~new_n1910_;
  assign new_n1912_ = new_n1360_ & ~new_n1911_;
  assign new_n1913_ = new_n1364_ & ~new_n1912_;
  assign new_n1914_ = new_n1368_ & ~new_n1913_;
  assign new_n1915_ = new_n1372_ & ~new_n1914_;
  assign new_n1916_ = new_n1376_ & ~new_n1915_;
  assign new_n1917_ = new_n1380_ & ~new_n1916_;
  assign new_n1918_ = new_n1384_ & ~new_n1917_;
  assign new_n1919_ = new_n1388_ & ~new_n1918_;
  assign new_n1920_ = new_n1392_ & ~new_n1919_;
  assign new_n1921_ = new_n1396_ & ~new_n1920_;
  assign new_n1922_ = new_n1663_ & ~new_n1921_;
  assign new_n1923_ = new_n392_ & ~new_n1922_;
  assign new_n1924_ = new_n396_ & ~new_n1923_;
  assign new_n1925_ = new_n400_ & ~new_n1924_;
  assign new_n1926_ = \req[8]  & ~new_n402_;
  assign \grant[8]  = ~new_n1925_ & new_n1926_;
  assign new_n1928_ = new_n411_ & ~new_n746_;
  assign new_n1929_ = new_n416_ & ~new_n1928_;
  assign new_n1930_ = new_n420_ & ~new_n1929_;
  assign new_n1931_ = new_n424_ & ~new_n1930_;
  assign new_n1932_ = new_n428_ & ~new_n1931_;
  assign new_n1933_ = new_n432_ & ~new_n1932_;
  assign new_n1934_ = new_n436_ & ~new_n1933_;
  assign new_n1935_ = new_n440_ & ~new_n1934_;
  assign new_n1936_ = new_n444_ & ~new_n1935_;
  assign new_n1937_ = new_n448_ & ~new_n1936_;
  assign new_n1938_ = new_n452_ & ~new_n1937_;
  assign new_n1939_ = new_n456_ & ~new_n1938_;
  assign new_n1940_ = new_n460_ & ~new_n1939_;
  assign new_n1941_ = new_n464_ & ~new_n1940_;
  assign new_n1942_ = new_n468_ & ~new_n1941_;
  assign new_n1943_ = new_n472_ & ~new_n1942_;
  assign new_n1944_ = new_n476_ & ~new_n1943_;
  assign new_n1945_ = new_n480_ & ~new_n1944_;
  assign new_n1946_ = new_n484_ & ~new_n1945_;
  assign new_n1947_ = new_n488_ & ~new_n1946_;
  assign new_n1948_ = new_n492_ & ~new_n1947_;
  assign new_n1949_ = new_n496_ & ~new_n1948_;
  assign new_n1950_ = new_n500_ & ~new_n1949_;
  assign new_n1951_ = new_n504_ & ~new_n1950_;
  assign new_n1952_ = new_n508_ & ~new_n1951_;
  assign new_n1953_ = new_n512_ & ~new_n1952_;
  assign new_n1954_ = new_n516_ & ~new_n1953_;
  assign new_n1955_ = new_n520_ & ~new_n1954_;
  assign new_n1956_ = new_n524_ & ~new_n1955_;
  assign new_n1957_ = new_n528_ & ~new_n1956_;
  assign new_n1958_ = new_n532_ & ~new_n1957_;
  assign new_n1959_ = new_n536_ & ~new_n1958_;
  assign new_n1960_ = new_n540_ & ~new_n1959_;
  assign new_n1961_ = new_n544_ & ~new_n1960_;
  assign new_n1962_ = new_n548_ & ~new_n1961_;
  assign new_n1963_ = new_n552_ & ~new_n1962_;
  assign new_n1964_ = new_n556_ & ~new_n1963_;
  assign new_n1965_ = new_n560_ & ~new_n1964_;
  assign new_n1966_ = new_n564_ & ~new_n1965_;
  assign new_n1967_ = new_n568_ & ~new_n1966_;
  assign new_n1968_ = new_n572_ & ~new_n1967_;
  assign new_n1969_ = new_n576_ & ~new_n1968_;
  assign new_n1970_ = new_n580_ & ~new_n1969_;
  assign new_n1971_ = new_n584_ & ~new_n1970_;
  assign new_n1972_ = new_n588_ & ~new_n1971_;
  assign new_n1973_ = new_n592_ & ~new_n1972_;
  assign new_n1974_ = new_n596_ & ~new_n1973_;
  assign new_n1975_ = new_n600_ & ~new_n1974_;
  assign new_n1976_ = new_n604_ & ~new_n1975_;
  assign new_n1977_ = new_n608_ & ~new_n1976_;
  assign new_n1978_ = new_n612_ & ~new_n1977_;
  assign new_n1979_ = new_n616_ & ~new_n1978_;
  assign new_n1980_ = new_n620_ & ~new_n1979_;
  assign new_n1981_ = new_n624_ & ~new_n1980_;
  assign new_n1982_ = new_n628_ & ~new_n1981_;
  assign new_n1983_ = new_n632_ & ~new_n1982_;
  assign new_n1984_ = new_n636_ & ~new_n1983_;
  assign new_n1985_ = new_n640_ & ~new_n1984_;
  assign new_n1986_ = new_n644_ & ~new_n1985_;
  assign new_n1987_ = new_n648_ & ~new_n1986_;
  assign new_n1988_ = new_n652_ & ~new_n1987_;
  assign new_n1989_ = new_n656_ & ~new_n1988_;
  assign new_n1990_ = new_n660_ & ~new_n1989_;
  assign new_n1991_ = new_n664_ & ~new_n1990_;
  assign new_n1992_ = new_n668_ & ~new_n1991_;
  assign new_n1993_ = new_n672_ & ~new_n1992_;
  assign new_n1994_ = new_n676_ & ~new_n1993_;
  assign new_n1995_ = new_n680_ & ~new_n1994_;
  assign new_n1996_ = new_n684_ & ~new_n1995_;
  assign new_n1997_ = new_n688_ & ~new_n1996_;
  assign new_n1998_ = new_n692_ & ~new_n1997_;
  assign new_n1999_ = new_n696_ & ~new_n1998_;
  assign new_n2000_ = new_n700_ & ~new_n1999_;
  assign new_n2001_ = new_n704_ & ~new_n2000_;
  assign new_n2002_ = new_n708_ & ~new_n2001_;
  assign new_n2003_ = new_n712_ & ~new_n2002_;
  assign new_n2004_ = new_n716_ & ~new_n2003_;
  assign new_n2005_ = new_n720_ & ~new_n2004_;
  assign new_n2006_ = new_n1484_ & ~new_n2005_;
  assign new_n2007_ = new_n1486_ & ~new_n2006_;
  assign new_n2008_ = new_n1750_ & ~new_n2007_;
  assign new_n2009_ = new_n731_ & ~new_n2008_;
  assign new_n2010_ = new_n735_ & ~new_n2009_;
  assign new_n2011_ = new_n739_ & ~new_n2010_;
  assign new_n2012_ = \req[9]  & ~new_n741_;
  assign \grant[9]  = ~new_n2011_ & new_n2012_;
  assign new_n2014_ = new_n750_ & ~new_n1083_;
  assign new_n2015_ = new_n755_ & ~new_n2014_;
  assign new_n2016_ = new_n759_ & ~new_n2015_;
  assign new_n2017_ = new_n763_ & ~new_n2016_;
  assign new_n2018_ = new_n767_ & ~new_n2017_;
  assign new_n2019_ = new_n771_ & ~new_n2018_;
  assign new_n2020_ = new_n775_ & ~new_n2019_;
  assign new_n2021_ = new_n779_ & ~new_n2020_;
  assign new_n2022_ = new_n783_ & ~new_n2021_;
  assign new_n2023_ = new_n787_ & ~new_n2022_;
  assign new_n2024_ = new_n791_ & ~new_n2023_;
  assign new_n2025_ = new_n795_ & ~new_n2024_;
  assign new_n2026_ = new_n799_ & ~new_n2025_;
  assign new_n2027_ = new_n803_ & ~new_n2026_;
  assign new_n2028_ = new_n807_ & ~new_n2027_;
  assign new_n2029_ = new_n811_ & ~new_n2028_;
  assign new_n2030_ = new_n815_ & ~new_n2029_;
  assign new_n2031_ = new_n819_ & ~new_n2030_;
  assign new_n2032_ = new_n823_ & ~new_n2031_;
  assign new_n2033_ = new_n827_ & ~new_n2032_;
  assign new_n2034_ = new_n831_ & ~new_n2033_;
  assign new_n2035_ = new_n835_ & ~new_n2034_;
  assign new_n2036_ = new_n839_ & ~new_n2035_;
  assign new_n2037_ = new_n843_ & ~new_n2036_;
  assign new_n2038_ = new_n847_ & ~new_n2037_;
  assign new_n2039_ = new_n851_ & ~new_n2038_;
  assign new_n2040_ = new_n855_ & ~new_n2039_;
  assign new_n2041_ = new_n859_ & ~new_n2040_;
  assign new_n2042_ = new_n863_ & ~new_n2041_;
  assign new_n2043_ = new_n867_ & ~new_n2042_;
  assign new_n2044_ = new_n871_ & ~new_n2043_;
  assign new_n2045_ = new_n875_ & ~new_n2044_;
  assign new_n2046_ = new_n879_ & ~new_n2045_;
  assign new_n2047_ = new_n883_ & ~new_n2046_;
  assign new_n2048_ = new_n887_ & ~new_n2047_;
  assign new_n2049_ = new_n891_ & ~new_n2048_;
  assign new_n2050_ = new_n895_ & ~new_n2049_;
  assign new_n2051_ = new_n899_ & ~new_n2050_;
  assign new_n2052_ = new_n903_ & ~new_n2051_;
  assign new_n2053_ = new_n907_ & ~new_n2052_;
  assign new_n2054_ = new_n911_ & ~new_n2053_;
  assign new_n2055_ = new_n915_ & ~new_n2054_;
  assign new_n2056_ = new_n919_ & ~new_n2055_;
  assign new_n2057_ = new_n923_ & ~new_n2056_;
  assign new_n2058_ = new_n927_ & ~new_n2057_;
  assign new_n2059_ = new_n931_ & ~new_n2058_;
  assign new_n2060_ = new_n935_ & ~new_n2059_;
  assign new_n2061_ = new_n939_ & ~new_n2060_;
  assign new_n2062_ = new_n943_ & ~new_n2061_;
  assign new_n2063_ = new_n947_ & ~new_n2062_;
  assign new_n2064_ = new_n951_ & ~new_n2063_;
  assign new_n2065_ = new_n955_ & ~new_n2064_;
  assign new_n2066_ = new_n959_ & ~new_n2065_;
  assign new_n2067_ = new_n963_ & ~new_n2066_;
  assign new_n2068_ = new_n967_ & ~new_n2067_;
  assign new_n2069_ = new_n971_ & ~new_n2068_;
  assign new_n2070_ = new_n975_ & ~new_n2069_;
  assign new_n2071_ = new_n979_ & ~new_n2070_;
  assign new_n2072_ = new_n983_ & ~new_n2071_;
  assign new_n2073_ = new_n987_ & ~new_n2072_;
  assign new_n2074_ = new_n991_ & ~new_n2073_;
  assign new_n2075_ = new_n995_ & ~new_n2074_;
  assign new_n2076_ = new_n999_ & ~new_n2075_;
  assign new_n2077_ = new_n1003_ & ~new_n2076_;
  assign new_n2078_ = new_n1007_ & ~new_n2077_;
  assign new_n2079_ = new_n1011_ & ~new_n2078_;
  assign new_n2080_ = new_n1015_ & ~new_n2079_;
  assign new_n2081_ = new_n1019_ & ~new_n2080_;
  assign new_n2082_ = new_n1023_ & ~new_n2081_;
  assign new_n2083_ = new_n1027_ & ~new_n2082_;
  assign new_n2084_ = new_n1031_ & ~new_n2083_;
  assign new_n2085_ = new_n1035_ & ~new_n2084_;
  assign new_n2086_ = new_n1039_ & ~new_n2085_;
  assign new_n2087_ = new_n1043_ & ~new_n2086_;
  assign new_n2088_ = new_n1047_ & ~new_n2087_;
  assign new_n2089_ = new_n1051_ & ~new_n2088_;
  assign new_n2090_ = new_n1055_ & ~new_n2089_;
  assign new_n2091_ = new_n1059_ & ~new_n2090_;
  assign new_n2092_ = new_n1574_ & ~new_n2091_;
  assign new_n2093_ = new_n1576_ & ~new_n2092_;
  assign new_n2094_ = new_n1837_ & ~new_n2093_;
  assign new_n2095_ = new_n1068_ & ~new_n2094_;
  assign new_n2096_ = new_n1072_ & ~new_n2095_;
  assign new_n2097_ = new_n1076_ & ~new_n2096_;
  assign new_n2098_ = \req[10]  & ~new_n1078_;
  assign \grant[10]  = ~new_n2097_ & new_n2098_;
  assign new_n2100_ = ~new_n415_ & new_n1087_;
  assign new_n2101_ = new_n1092_ & ~new_n2100_;
  assign new_n2102_ = new_n1096_ & ~new_n2101_;
  assign new_n2103_ = new_n1100_ & ~new_n2102_;
  assign new_n2104_ = new_n1104_ & ~new_n2103_;
  assign new_n2105_ = new_n1108_ & ~new_n2104_;
  assign new_n2106_ = new_n1112_ & ~new_n2105_;
  assign new_n2107_ = new_n1116_ & ~new_n2106_;
  assign new_n2108_ = new_n1120_ & ~new_n2107_;
  assign new_n2109_ = new_n1124_ & ~new_n2108_;
  assign new_n2110_ = new_n1128_ & ~new_n2109_;
  assign new_n2111_ = new_n1132_ & ~new_n2110_;
  assign new_n2112_ = new_n1136_ & ~new_n2111_;
  assign new_n2113_ = new_n1140_ & ~new_n2112_;
  assign new_n2114_ = new_n1144_ & ~new_n2113_;
  assign new_n2115_ = new_n1148_ & ~new_n2114_;
  assign new_n2116_ = new_n1152_ & ~new_n2115_;
  assign new_n2117_ = new_n1156_ & ~new_n2116_;
  assign new_n2118_ = new_n1160_ & ~new_n2117_;
  assign new_n2119_ = new_n1164_ & ~new_n2118_;
  assign new_n2120_ = new_n1168_ & ~new_n2119_;
  assign new_n2121_ = new_n1172_ & ~new_n2120_;
  assign new_n2122_ = new_n1176_ & ~new_n2121_;
  assign new_n2123_ = new_n1180_ & ~new_n2122_;
  assign new_n2124_ = new_n1184_ & ~new_n2123_;
  assign new_n2125_ = new_n1188_ & ~new_n2124_;
  assign new_n2126_ = new_n1192_ & ~new_n2125_;
  assign new_n2127_ = new_n1196_ & ~new_n2126_;
  assign new_n2128_ = new_n1200_ & ~new_n2127_;
  assign new_n2129_ = new_n1204_ & ~new_n2128_;
  assign new_n2130_ = new_n1208_ & ~new_n2129_;
  assign new_n2131_ = new_n1212_ & ~new_n2130_;
  assign new_n2132_ = new_n1216_ & ~new_n2131_;
  assign new_n2133_ = new_n1220_ & ~new_n2132_;
  assign new_n2134_ = new_n1224_ & ~new_n2133_;
  assign new_n2135_ = new_n1228_ & ~new_n2134_;
  assign new_n2136_ = new_n1232_ & ~new_n2135_;
  assign new_n2137_ = new_n1236_ & ~new_n2136_;
  assign new_n2138_ = new_n1240_ & ~new_n2137_;
  assign new_n2139_ = new_n1244_ & ~new_n2138_;
  assign new_n2140_ = new_n1248_ & ~new_n2139_;
  assign new_n2141_ = new_n1252_ & ~new_n2140_;
  assign new_n2142_ = new_n1256_ & ~new_n2141_;
  assign new_n2143_ = new_n1260_ & ~new_n2142_;
  assign new_n2144_ = new_n1264_ & ~new_n2143_;
  assign new_n2145_ = new_n1268_ & ~new_n2144_;
  assign new_n2146_ = new_n1272_ & ~new_n2145_;
  assign new_n2147_ = new_n1276_ & ~new_n2146_;
  assign new_n2148_ = new_n1280_ & ~new_n2147_;
  assign new_n2149_ = new_n1284_ & ~new_n2148_;
  assign new_n2150_ = new_n1288_ & ~new_n2149_;
  assign new_n2151_ = new_n1292_ & ~new_n2150_;
  assign new_n2152_ = new_n1296_ & ~new_n2151_;
  assign new_n2153_ = new_n1300_ & ~new_n2152_;
  assign new_n2154_ = new_n1304_ & ~new_n2153_;
  assign new_n2155_ = new_n1308_ & ~new_n2154_;
  assign new_n2156_ = new_n1312_ & ~new_n2155_;
  assign new_n2157_ = new_n1316_ & ~new_n2156_;
  assign new_n2158_ = new_n1320_ & ~new_n2157_;
  assign new_n2159_ = new_n1324_ & ~new_n2158_;
  assign new_n2160_ = new_n1328_ & ~new_n2159_;
  assign new_n2161_ = new_n1332_ & ~new_n2160_;
  assign new_n2162_ = new_n1336_ & ~new_n2161_;
  assign new_n2163_ = new_n1340_ & ~new_n2162_;
  assign new_n2164_ = new_n1344_ & ~new_n2163_;
  assign new_n2165_ = new_n1348_ & ~new_n2164_;
  assign new_n2166_ = new_n1352_ & ~new_n2165_;
  assign new_n2167_ = new_n1356_ & ~new_n2166_;
  assign new_n2168_ = new_n1360_ & ~new_n2167_;
  assign new_n2169_ = new_n1364_ & ~new_n2168_;
  assign new_n2170_ = new_n1368_ & ~new_n2169_;
  assign new_n2171_ = new_n1372_ & ~new_n2170_;
  assign new_n2172_ = new_n1376_ & ~new_n2171_;
  assign new_n2173_ = new_n1380_ & ~new_n2172_;
  assign new_n2174_ = new_n1384_ & ~new_n2173_;
  assign new_n2175_ = new_n1388_ & ~new_n2174_;
  assign new_n2176_ = new_n1392_ & ~new_n2175_;
  assign new_n2177_ = new_n1396_ & ~new_n2176_;
  assign new_n2178_ = new_n1663_ & ~new_n2177_;
  assign new_n2179_ = new_n392_ & ~new_n2178_;
  assign new_n2180_ = new_n396_ & ~new_n2179_;
  assign new_n2181_ = new_n400_ & ~new_n2180_;
  assign new_n2182_ = new_n404_ & ~new_n2181_;
  assign new_n2183_ = new_n408_ & ~new_n2182_;
  assign new_n2184_ = \req[11]  & ~new_n410_;
  assign \grant[11]  = ~new_n2183_ & new_n2184_;
  assign new_n2186_ = new_n419_ & ~new_n754_;
  assign new_n2187_ = new_n424_ & ~new_n2186_;
  assign new_n2188_ = new_n428_ & ~new_n2187_;
  assign new_n2189_ = new_n432_ & ~new_n2188_;
  assign new_n2190_ = new_n436_ & ~new_n2189_;
  assign new_n2191_ = new_n440_ & ~new_n2190_;
  assign new_n2192_ = new_n444_ & ~new_n2191_;
  assign new_n2193_ = new_n448_ & ~new_n2192_;
  assign new_n2194_ = new_n452_ & ~new_n2193_;
  assign new_n2195_ = new_n456_ & ~new_n2194_;
  assign new_n2196_ = new_n460_ & ~new_n2195_;
  assign new_n2197_ = new_n464_ & ~new_n2196_;
  assign new_n2198_ = new_n468_ & ~new_n2197_;
  assign new_n2199_ = new_n472_ & ~new_n2198_;
  assign new_n2200_ = new_n476_ & ~new_n2199_;
  assign new_n2201_ = new_n480_ & ~new_n2200_;
  assign new_n2202_ = new_n484_ & ~new_n2201_;
  assign new_n2203_ = new_n488_ & ~new_n2202_;
  assign new_n2204_ = new_n492_ & ~new_n2203_;
  assign new_n2205_ = new_n496_ & ~new_n2204_;
  assign new_n2206_ = new_n500_ & ~new_n2205_;
  assign new_n2207_ = new_n504_ & ~new_n2206_;
  assign new_n2208_ = new_n508_ & ~new_n2207_;
  assign new_n2209_ = new_n512_ & ~new_n2208_;
  assign new_n2210_ = new_n516_ & ~new_n2209_;
  assign new_n2211_ = new_n520_ & ~new_n2210_;
  assign new_n2212_ = new_n524_ & ~new_n2211_;
  assign new_n2213_ = new_n528_ & ~new_n2212_;
  assign new_n2214_ = new_n532_ & ~new_n2213_;
  assign new_n2215_ = new_n536_ & ~new_n2214_;
  assign new_n2216_ = new_n540_ & ~new_n2215_;
  assign new_n2217_ = new_n544_ & ~new_n2216_;
  assign new_n2218_ = new_n548_ & ~new_n2217_;
  assign new_n2219_ = new_n552_ & ~new_n2218_;
  assign new_n2220_ = new_n556_ & ~new_n2219_;
  assign new_n2221_ = new_n560_ & ~new_n2220_;
  assign new_n2222_ = new_n564_ & ~new_n2221_;
  assign new_n2223_ = new_n568_ & ~new_n2222_;
  assign new_n2224_ = new_n572_ & ~new_n2223_;
  assign new_n2225_ = new_n576_ & ~new_n2224_;
  assign new_n2226_ = new_n580_ & ~new_n2225_;
  assign new_n2227_ = new_n584_ & ~new_n2226_;
  assign new_n2228_ = new_n588_ & ~new_n2227_;
  assign new_n2229_ = new_n592_ & ~new_n2228_;
  assign new_n2230_ = new_n596_ & ~new_n2229_;
  assign new_n2231_ = new_n600_ & ~new_n2230_;
  assign new_n2232_ = new_n604_ & ~new_n2231_;
  assign new_n2233_ = new_n608_ & ~new_n2232_;
  assign new_n2234_ = new_n612_ & ~new_n2233_;
  assign new_n2235_ = new_n616_ & ~new_n2234_;
  assign new_n2236_ = new_n620_ & ~new_n2235_;
  assign new_n2237_ = new_n624_ & ~new_n2236_;
  assign new_n2238_ = new_n628_ & ~new_n2237_;
  assign new_n2239_ = new_n632_ & ~new_n2238_;
  assign new_n2240_ = new_n636_ & ~new_n2239_;
  assign new_n2241_ = new_n640_ & ~new_n2240_;
  assign new_n2242_ = new_n644_ & ~new_n2241_;
  assign new_n2243_ = new_n648_ & ~new_n2242_;
  assign new_n2244_ = new_n652_ & ~new_n2243_;
  assign new_n2245_ = new_n656_ & ~new_n2244_;
  assign new_n2246_ = new_n660_ & ~new_n2245_;
  assign new_n2247_ = new_n664_ & ~new_n2246_;
  assign new_n2248_ = new_n668_ & ~new_n2247_;
  assign new_n2249_ = new_n672_ & ~new_n2248_;
  assign new_n2250_ = new_n676_ & ~new_n2249_;
  assign new_n2251_ = new_n680_ & ~new_n2250_;
  assign new_n2252_ = new_n684_ & ~new_n2251_;
  assign new_n2253_ = new_n688_ & ~new_n2252_;
  assign new_n2254_ = new_n692_ & ~new_n2253_;
  assign new_n2255_ = new_n696_ & ~new_n2254_;
  assign new_n2256_ = new_n700_ & ~new_n2255_;
  assign new_n2257_ = new_n704_ & ~new_n2256_;
  assign new_n2258_ = new_n708_ & ~new_n2257_;
  assign new_n2259_ = new_n712_ & ~new_n2258_;
  assign new_n2260_ = new_n716_ & ~new_n2259_;
  assign new_n2261_ = new_n720_ & ~new_n2260_;
  assign new_n2262_ = new_n1484_ & ~new_n2261_;
  assign new_n2263_ = new_n1486_ & ~new_n2262_;
  assign new_n2264_ = new_n1750_ & ~new_n2263_;
  assign new_n2265_ = new_n731_ & ~new_n2264_;
  assign new_n2266_ = new_n735_ & ~new_n2265_;
  assign new_n2267_ = new_n739_ & ~new_n2266_;
  assign new_n2268_ = new_n743_ & ~new_n2267_;
  assign new_n2269_ = new_n747_ & ~new_n2268_;
  assign new_n2270_ = \req[12]  & ~new_n749_;
  assign \grant[12]  = ~new_n2269_ & new_n2270_;
  assign new_n2272_ = new_n758_ & ~new_n1091_;
  assign new_n2273_ = new_n763_ & ~new_n2272_;
  assign new_n2274_ = new_n767_ & ~new_n2273_;
  assign new_n2275_ = new_n771_ & ~new_n2274_;
  assign new_n2276_ = new_n775_ & ~new_n2275_;
  assign new_n2277_ = new_n779_ & ~new_n2276_;
  assign new_n2278_ = new_n783_ & ~new_n2277_;
  assign new_n2279_ = new_n787_ & ~new_n2278_;
  assign new_n2280_ = new_n791_ & ~new_n2279_;
  assign new_n2281_ = new_n795_ & ~new_n2280_;
  assign new_n2282_ = new_n799_ & ~new_n2281_;
  assign new_n2283_ = new_n803_ & ~new_n2282_;
  assign new_n2284_ = new_n807_ & ~new_n2283_;
  assign new_n2285_ = new_n811_ & ~new_n2284_;
  assign new_n2286_ = new_n815_ & ~new_n2285_;
  assign new_n2287_ = new_n819_ & ~new_n2286_;
  assign new_n2288_ = new_n823_ & ~new_n2287_;
  assign new_n2289_ = new_n827_ & ~new_n2288_;
  assign new_n2290_ = new_n831_ & ~new_n2289_;
  assign new_n2291_ = new_n835_ & ~new_n2290_;
  assign new_n2292_ = new_n839_ & ~new_n2291_;
  assign new_n2293_ = new_n843_ & ~new_n2292_;
  assign new_n2294_ = new_n847_ & ~new_n2293_;
  assign new_n2295_ = new_n851_ & ~new_n2294_;
  assign new_n2296_ = new_n855_ & ~new_n2295_;
  assign new_n2297_ = new_n859_ & ~new_n2296_;
  assign new_n2298_ = new_n863_ & ~new_n2297_;
  assign new_n2299_ = new_n867_ & ~new_n2298_;
  assign new_n2300_ = new_n871_ & ~new_n2299_;
  assign new_n2301_ = new_n875_ & ~new_n2300_;
  assign new_n2302_ = new_n879_ & ~new_n2301_;
  assign new_n2303_ = new_n883_ & ~new_n2302_;
  assign new_n2304_ = new_n887_ & ~new_n2303_;
  assign new_n2305_ = new_n891_ & ~new_n2304_;
  assign new_n2306_ = new_n895_ & ~new_n2305_;
  assign new_n2307_ = new_n899_ & ~new_n2306_;
  assign new_n2308_ = new_n903_ & ~new_n2307_;
  assign new_n2309_ = new_n907_ & ~new_n2308_;
  assign new_n2310_ = new_n911_ & ~new_n2309_;
  assign new_n2311_ = new_n915_ & ~new_n2310_;
  assign new_n2312_ = new_n919_ & ~new_n2311_;
  assign new_n2313_ = new_n923_ & ~new_n2312_;
  assign new_n2314_ = new_n927_ & ~new_n2313_;
  assign new_n2315_ = new_n931_ & ~new_n2314_;
  assign new_n2316_ = new_n935_ & ~new_n2315_;
  assign new_n2317_ = new_n939_ & ~new_n2316_;
  assign new_n2318_ = new_n943_ & ~new_n2317_;
  assign new_n2319_ = new_n947_ & ~new_n2318_;
  assign new_n2320_ = new_n951_ & ~new_n2319_;
  assign new_n2321_ = new_n955_ & ~new_n2320_;
  assign new_n2322_ = new_n959_ & ~new_n2321_;
  assign new_n2323_ = new_n963_ & ~new_n2322_;
  assign new_n2324_ = new_n967_ & ~new_n2323_;
  assign new_n2325_ = new_n971_ & ~new_n2324_;
  assign new_n2326_ = new_n975_ & ~new_n2325_;
  assign new_n2327_ = new_n979_ & ~new_n2326_;
  assign new_n2328_ = new_n983_ & ~new_n2327_;
  assign new_n2329_ = new_n987_ & ~new_n2328_;
  assign new_n2330_ = new_n991_ & ~new_n2329_;
  assign new_n2331_ = new_n995_ & ~new_n2330_;
  assign new_n2332_ = new_n999_ & ~new_n2331_;
  assign new_n2333_ = new_n1003_ & ~new_n2332_;
  assign new_n2334_ = new_n1007_ & ~new_n2333_;
  assign new_n2335_ = new_n1011_ & ~new_n2334_;
  assign new_n2336_ = new_n1015_ & ~new_n2335_;
  assign new_n2337_ = new_n1019_ & ~new_n2336_;
  assign new_n2338_ = new_n1023_ & ~new_n2337_;
  assign new_n2339_ = new_n1027_ & ~new_n2338_;
  assign new_n2340_ = new_n1031_ & ~new_n2339_;
  assign new_n2341_ = new_n1035_ & ~new_n2340_;
  assign new_n2342_ = new_n1039_ & ~new_n2341_;
  assign new_n2343_ = new_n1043_ & ~new_n2342_;
  assign new_n2344_ = new_n1047_ & ~new_n2343_;
  assign new_n2345_ = new_n1051_ & ~new_n2344_;
  assign new_n2346_ = new_n1055_ & ~new_n2345_;
  assign new_n2347_ = new_n1059_ & ~new_n2346_;
  assign new_n2348_ = new_n1574_ & ~new_n2347_;
  assign new_n2349_ = new_n1576_ & ~new_n2348_;
  assign new_n2350_ = new_n1837_ & ~new_n2349_;
  assign new_n2351_ = new_n1068_ & ~new_n2350_;
  assign new_n2352_ = new_n1072_ & ~new_n2351_;
  assign new_n2353_ = new_n1076_ & ~new_n2352_;
  assign new_n2354_ = new_n1080_ & ~new_n2353_;
  assign new_n2355_ = new_n1084_ & ~new_n2354_;
  assign new_n2356_ = \req[13]  & ~new_n1086_;
  assign \grant[13]  = ~new_n2355_ & new_n2356_;
  assign new_n2358_ = ~new_n423_ & new_n1095_;
  assign new_n2359_ = new_n1100_ & ~new_n2358_;
  assign new_n2360_ = new_n1104_ & ~new_n2359_;
  assign new_n2361_ = new_n1108_ & ~new_n2360_;
  assign new_n2362_ = new_n1112_ & ~new_n2361_;
  assign new_n2363_ = new_n1116_ & ~new_n2362_;
  assign new_n2364_ = new_n1120_ & ~new_n2363_;
  assign new_n2365_ = new_n1124_ & ~new_n2364_;
  assign new_n2366_ = new_n1128_ & ~new_n2365_;
  assign new_n2367_ = new_n1132_ & ~new_n2366_;
  assign new_n2368_ = new_n1136_ & ~new_n2367_;
  assign new_n2369_ = new_n1140_ & ~new_n2368_;
  assign new_n2370_ = new_n1144_ & ~new_n2369_;
  assign new_n2371_ = new_n1148_ & ~new_n2370_;
  assign new_n2372_ = new_n1152_ & ~new_n2371_;
  assign new_n2373_ = new_n1156_ & ~new_n2372_;
  assign new_n2374_ = new_n1160_ & ~new_n2373_;
  assign new_n2375_ = new_n1164_ & ~new_n2374_;
  assign new_n2376_ = new_n1168_ & ~new_n2375_;
  assign new_n2377_ = new_n1172_ & ~new_n2376_;
  assign new_n2378_ = new_n1176_ & ~new_n2377_;
  assign new_n2379_ = new_n1180_ & ~new_n2378_;
  assign new_n2380_ = new_n1184_ & ~new_n2379_;
  assign new_n2381_ = new_n1188_ & ~new_n2380_;
  assign new_n2382_ = new_n1192_ & ~new_n2381_;
  assign new_n2383_ = new_n1196_ & ~new_n2382_;
  assign new_n2384_ = new_n1200_ & ~new_n2383_;
  assign new_n2385_ = new_n1204_ & ~new_n2384_;
  assign new_n2386_ = new_n1208_ & ~new_n2385_;
  assign new_n2387_ = new_n1212_ & ~new_n2386_;
  assign new_n2388_ = new_n1216_ & ~new_n2387_;
  assign new_n2389_ = new_n1220_ & ~new_n2388_;
  assign new_n2390_ = new_n1224_ & ~new_n2389_;
  assign new_n2391_ = new_n1228_ & ~new_n2390_;
  assign new_n2392_ = new_n1232_ & ~new_n2391_;
  assign new_n2393_ = new_n1236_ & ~new_n2392_;
  assign new_n2394_ = new_n1240_ & ~new_n2393_;
  assign new_n2395_ = new_n1244_ & ~new_n2394_;
  assign new_n2396_ = new_n1248_ & ~new_n2395_;
  assign new_n2397_ = new_n1252_ & ~new_n2396_;
  assign new_n2398_ = new_n1256_ & ~new_n2397_;
  assign new_n2399_ = new_n1260_ & ~new_n2398_;
  assign new_n2400_ = new_n1264_ & ~new_n2399_;
  assign new_n2401_ = new_n1268_ & ~new_n2400_;
  assign new_n2402_ = new_n1272_ & ~new_n2401_;
  assign new_n2403_ = new_n1276_ & ~new_n2402_;
  assign new_n2404_ = new_n1280_ & ~new_n2403_;
  assign new_n2405_ = new_n1284_ & ~new_n2404_;
  assign new_n2406_ = new_n1288_ & ~new_n2405_;
  assign new_n2407_ = new_n1292_ & ~new_n2406_;
  assign new_n2408_ = new_n1296_ & ~new_n2407_;
  assign new_n2409_ = new_n1300_ & ~new_n2408_;
  assign new_n2410_ = new_n1304_ & ~new_n2409_;
  assign new_n2411_ = new_n1308_ & ~new_n2410_;
  assign new_n2412_ = new_n1312_ & ~new_n2411_;
  assign new_n2413_ = new_n1316_ & ~new_n2412_;
  assign new_n2414_ = new_n1320_ & ~new_n2413_;
  assign new_n2415_ = new_n1324_ & ~new_n2414_;
  assign new_n2416_ = new_n1328_ & ~new_n2415_;
  assign new_n2417_ = new_n1332_ & ~new_n2416_;
  assign new_n2418_ = new_n1336_ & ~new_n2417_;
  assign new_n2419_ = new_n1340_ & ~new_n2418_;
  assign new_n2420_ = new_n1344_ & ~new_n2419_;
  assign new_n2421_ = new_n1348_ & ~new_n2420_;
  assign new_n2422_ = new_n1352_ & ~new_n2421_;
  assign new_n2423_ = new_n1356_ & ~new_n2422_;
  assign new_n2424_ = new_n1360_ & ~new_n2423_;
  assign new_n2425_ = new_n1364_ & ~new_n2424_;
  assign new_n2426_ = new_n1368_ & ~new_n2425_;
  assign new_n2427_ = new_n1372_ & ~new_n2426_;
  assign new_n2428_ = new_n1376_ & ~new_n2427_;
  assign new_n2429_ = new_n1380_ & ~new_n2428_;
  assign new_n2430_ = new_n1384_ & ~new_n2429_;
  assign new_n2431_ = new_n1388_ & ~new_n2430_;
  assign new_n2432_ = new_n1392_ & ~new_n2431_;
  assign new_n2433_ = new_n1396_ & ~new_n2432_;
  assign new_n2434_ = new_n1663_ & ~new_n2433_;
  assign new_n2435_ = new_n392_ & ~new_n2434_;
  assign new_n2436_ = new_n396_ & ~new_n2435_;
  assign new_n2437_ = new_n400_ & ~new_n2436_;
  assign new_n2438_ = new_n404_ & ~new_n2437_;
  assign new_n2439_ = new_n408_ & ~new_n2438_;
  assign new_n2440_ = new_n412_ & ~new_n2439_;
  assign new_n2441_ = new_n416_ & ~new_n2440_;
  assign new_n2442_ = \req[14]  & ~new_n418_;
  assign \grant[14]  = ~new_n2441_ & new_n2442_;
  assign new_n2444_ = new_n427_ & ~new_n762_;
  assign new_n2445_ = new_n432_ & ~new_n2444_;
  assign new_n2446_ = new_n436_ & ~new_n2445_;
  assign new_n2447_ = new_n440_ & ~new_n2446_;
  assign new_n2448_ = new_n444_ & ~new_n2447_;
  assign new_n2449_ = new_n448_ & ~new_n2448_;
  assign new_n2450_ = new_n452_ & ~new_n2449_;
  assign new_n2451_ = new_n456_ & ~new_n2450_;
  assign new_n2452_ = new_n460_ & ~new_n2451_;
  assign new_n2453_ = new_n464_ & ~new_n2452_;
  assign new_n2454_ = new_n468_ & ~new_n2453_;
  assign new_n2455_ = new_n472_ & ~new_n2454_;
  assign new_n2456_ = new_n476_ & ~new_n2455_;
  assign new_n2457_ = new_n480_ & ~new_n2456_;
  assign new_n2458_ = new_n484_ & ~new_n2457_;
  assign new_n2459_ = new_n488_ & ~new_n2458_;
  assign new_n2460_ = new_n492_ & ~new_n2459_;
  assign new_n2461_ = new_n496_ & ~new_n2460_;
  assign new_n2462_ = new_n500_ & ~new_n2461_;
  assign new_n2463_ = new_n504_ & ~new_n2462_;
  assign new_n2464_ = new_n508_ & ~new_n2463_;
  assign new_n2465_ = new_n512_ & ~new_n2464_;
  assign new_n2466_ = new_n516_ & ~new_n2465_;
  assign new_n2467_ = new_n520_ & ~new_n2466_;
  assign new_n2468_ = new_n524_ & ~new_n2467_;
  assign new_n2469_ = new_n528_ & ~new_n2468_;
  assign new_n2470_ = new_n532_ & ~new_n2469_;
  assign new_n2471_ = new_n536_ & ~new_n2470_;
  assign new_n2472_ = new_n540_ & ~new_n2471_;
  assign new_n2473_ = new_n544_ & ~new_n2472_;
  assign new_n2474_ = new_n548_ & ~new_n2473_;
  assign new_n2475_ = new_n552_ & ~new_n2474_;
  assign new_n2476_ = new_n556_ & ~new_n2475_;
  assign new_n2477_ = new_n560_ & ~new_n2476_;
  assign new_n2478_ = new_n564_ & ~new_n2477_;
  assign new_n2479_ = new_n568_ & ~new_n2478_;
  assign new_n2480_ = new_n572_ & ~new_n2479_;
  assign new_n2481_ = new_n576_ & ~new_n2480_;
  assign new_n2482_ = new_n580_ & ~new_n2481_;
  assign new_n2483_ = new_n584_ & ~new_n2482_;
  assign new_n2484_ = new_n588_ & ~new_n2483_;
  assign new_n2485_ = new_n592_ & ~new_n2484_;
  assign new_n2486_ = new_n596_ & ~new_n2485_;
  assign new_n2487_ = new_n600_ & ~new_n2486_;
  assign new_n2488_ = new_n604_ & ~new_n2487_;
  assign new_n2489_ = new_n608_ & ~new_n2488_;
  assign new_n2490_ = new_n612_ & ~new_n2489_;
  assign new_n2491_ = new_n616_ & ~new_n2490_;
  assign new_n2492_ = new_n620_ & ~new_n2491_;
  assign new_n2493_ = new_n624_ & ~new_n2492_;
  assign new_n2494_ = new_n628_ & ~new_n2493_;
  assign new_n2495_ = new_n632_ & ~new_n2494_;
  assign new_n2496_ = new_n636_ & ~new_n2495_;
  assign new_n2497_ = new_n640_ & ~new_n2496_;
  assign new_n2498_ = new_n644_ & ~new_n2497_;
  assign new_n2499_ = new_n648_ & ~new_n2498_;
  assign new_n2500_ = new_n652_ & ~new_n2499_;
  assign new_n2501_ = new_n656_ & ~new_n2500_;
  assign new_n2502_ = new_n660_ & ~new_n2501_;
  assign new_n2503_ = new_n664_ & ~new_n2502_;
  assign new_n2504_ = new_n668_ & ~new_n2503_;
  assign new_n2505_ = new_n672_ & ~new_n2504_;
  assign new_n2506_ = new_n676_ & ~new_n2505_;
  assign new_n2507_ = new_n680_ & ~new_n2506_;
  assign new_n2508_ = new_n684_ & ~new_n2507_;
  assign new_n2509_ = new_n688_ & ~new_n2508_;
  assign new_n2510_ = new_n692_ & ~new_n2509_;
  assign new_n2511_ = new_n696_ & ~new_n2510_;
  assign new_n2512_ = new_n700_ & ~new_n2511_;
  assign new_n2513_ = new_n704_ & ~new_n2512_;
  assign new_n2514_ = new_n708_ & ~new_n2513_;
  assign new_n2515_ = new_n712_ & ~new_n2514_;
  assign new_n2516_ = new_n716_ & ~new_n2515_;
  assign new_n2517_ = new_n720_ & ~new_n2516_;
  assign new_n2518_ = new_n1484_ & ~new_n2517_;
  assign new_n2519_ = new_n1486_ & ~new_n2518_;
  assign new_n2520_ = new_n1750_ & ~new_n2519_;
  assign new_n2521_ = new_n731_ & ~new_n2520_;
  assign new_n2522_ = new_n735_ & ~new_n2521_;
  assign new_n2523_ = new_n739_ & ~new_n2522_;
  assign new_n2524_ = new_n743_ & ~new_n2523_;
  assign new_n2525_ = new_n747_ & ~new_n2524_;
  assign new_n2526_ = new_n751_ & ~new_n2525_;
  assign new_n2527_ = new_n755_ & ~new_n2526_;
  assign new_n2528_ = \req[15]  & ~new_n757_;
  assign \grant[15]  = ~new_n2527_ & new_n2528_;
  assign new_n2530_ = new_n766_ & ~new_n1099_;
  assign new_n2531_ = new_n771_ & ~new_n2530_;
  assign new_n2532_ = new_n775_ & ~new_n2531_;
  assign new_n2533_ = new_n779_ & ~new_n2532_;
  assign new_n2534_ = new_n783_ & ~new_n2533_;
  assign new_n2535_ = new_n787_ & ~new_n2534_;
  assign new_n2536_ = new_n791_ & ~new_n2535_;
  assign new_n2537_ = new_n795_ & ~new_n2536_;
  assign new_n2538_ = new_n799_ & ~new_n2537_;
  assign new_n2539_ = new_n803_ & ~new_n2538_;
  assign new_n2540_ = new_n807_ & ~new_n2539_;
  assign new_n2541_ = new_n811_ & ~new_n2540_;
  assign new_n2542_ = new_n815_ & ~new_n2541_;
  assign new_n2543_ = new_n819_ & ~new_n2542_;
  assign new_n2544_ = new_n823_ & ~new_n2543_;
  assign new_n2545_ = new_n827_ & ~new_n2544_;
  assign new_n2546_ = new_n831_ & ~new_n2545_;
  assign new_n2547_ = new_n835_ & ~new_n2546_;
  assign new_n2548_ = new_n839_ & ~new_n2547_;
  assign new_n2549_ = new_n843_ & ~new_n2548_;
  assign new_n2550_ = new_n847_ & ~new_n2549_;
  assign new_n2551_ = new_n851_ & ~new_n2550_;
  assign new_n2552_ = new_n855_ & ~new_n2551_;
  assign new_n2553_ = new_n859_ & ~new_n2552_;
  assign new_n2554_ = new_n863_ & ~new_n2553_;
  assign new_n2555_ = new_n867_ & ~new_n2554_;
  assign new_n2556_ = new_n871_ & ~new_n2555_;
  assign new_n2557_ = new_n875_ & ~new_n2556_;
  assign new_n2558_ = new_n879_ & ~new_n2557_;
  assign new_n2559_ = new_n883_ & ~new_n2558_;
  assign new_n2560_ = new_n887_ & ~new_n2559_;
  assign new_n2561_ = new_n891_ & ~new_n2560_;
  assign new_n2562_ = new_n895_ & ~new_n2561_;
  assign new_n2563_ = new_n899_ & ~new_n2562_;
  assign new_n2564_ = new_n903_ & ~new_n2563_;
  assign new_n2565_ = new_n907_ & ~new_n2564_;
  assign new_n2566_ = new_n911_ & ~new_n2565_;
  assign new_n2567_ = new_n915_ & ~new_n2566_;
  assign new_n2568_ = new_n919_ & ~new_n2567_;
  assign new_n2569_ = new_n923_ & ~new_n2568_;
  assign new_n2570_ = new_n927_ & ~new_n2569_;
  assign new_n2571_ = new_n931_ & ~new_n2570_;
  assign new_n2572_ = new_n935_ & ~new_n2571_;
  assign new_n2573_ = new_n939_ & ~new_n2572_;
  assign new_n2574_ = new_n943_ & ~new_n2573_;
  assign new_n2575_ = new_n947_ & ~new_n2574_;
  assign new_n2576_ = new_n951_ & ~new_n2575_;
  assign new_n2577_ = new_n955_ & ~new_n2576_;
  assign new_n2578_ = new_n959_ & ~new_n2577_;
  assign new_n2579_ = new_n963_ & ~new_n2578_;
  assign new_n2580_ = new_n967_ & ~new_n2579_;
  assign new_n2581_ = new_n971_ & ~new_n2580_;
  assign new_n2582_ = new_n975_ & ~new_n2581_;
  assign new_n2583_ = new_n979_ & ~new_n2582_;
  assign new_n2584_ = new_n983_ & ~new_n2583_;
  assign new_n2585_ = new_n987_ & ~new_n2584_;
  assign new_n2586_ = new_n991_ & ~new_n2585_;
  assign new_n2587_ = new_n995_ & ~new_n2586_;
  assign new_n2588_ = new_n999_ & ~new_n2587_;
  assign new_n2589_ = new_n1003_ & ~new_n2588_;
  assign new_n2590_ = new_n1007_ & ~new_n2589_;
  assign new_n2591_ = new_n1011_ & ~new_n2590_;
  assign new_n2592_ = new_n1015_ & ~new_n2591_;
  assign new_n2593_ = new_n1019_ & ~new_n2592_;
  assign new_n2594_ = new_n1023_ & ~new_n2593_;
  assign new_n2595_ = new_n1027_ & ~new_n2594_;
  assign new_n2596_ = new_n1031_ & ~new_n2595_;
  assign new_n2597_ = new_n1035_ & ~new_n2596_;
  assign new_n2598_ = new_n1039_ & ~new_n2597_;
  assign new_n2599_ = new_n1043_ & ~new_n2598_;
  assign new_n2600_ = new_n1047_ & ~new_n2599_;
  assign new_n2601_ = new_n1051_ & ~new_n2600_;
  assign new_n2602_ = new_n1055_ & ~new_n2601_;
  assign new_n2603_ = new_n1059_ & ~new_n2602_;
  assign new_n2604_ = new_n1574_ & ~new_n2603_;
  assign new_n2605_ = new_n1576_ & ~new_n2604_;
  assign new_n2606_ = new_n1837_ & ~new_n2605_;
  assign new_n2607_ = new_n1068_ & ~new_n2606_;
  assign new_n2608_ = new_n1072_ & ~new_n2607_;
  assign new_n2609_ = new_n1076_ & ~new_n2608_;
  assign new_n2610_ = new_n1080_ & ~new_n2609_;
  assign new_n2611_ = new_n1084_ & ~new_n2610_;
  assign new_n2612_ = new_n1088_ & ~new_n2611_;
  assign new_n2613_ = new_n1092_ & ~new_n2612_;
  assign new_n2614_ = \req[16]  & ~new_n1094_;
  assign \grant[16]  = ~new_n2613_ & new_n2614_;
  assign new_n2616_ = ~new_n431_ & new_n1103_;
  assign new_n2617_ = new_n1108_ & ~new_n2616_;
  assign new_n2618_ = new_n1112_ & ~new_n2617_;
  assign new_n2619_ = new_n1116_ & ~new_n2618_;
  assign new_n2620_ = new_n1120_ & ~new_n2619_;
  assign new_n2621_ = new_n1124_ & ~new_n2620_;
  assign new_n2622_ = new_n1128_ & ~new_n2621_;
  assign new_n2623_ = new_n1132_ & ~new_n2622_;
  assign new_n2624_ = new_n1136_ & ~new_n2623_;
  assign new_n2625_ = new_n1140_ & ~new_n2624_;
  assign new_n2626_ = new_n1144_ & ~new_n2625_;
  assign new_n2627_ = new_n1148_ & ~new_n2626_;
  assign new_n2628_ = new_n1152_ & ~new_n2627_;
  assign new_n2629_ = new_n1156_ & ~new_n2628_;
  assign new_n2630_ = new_n1160_ & ~new_n2629_;
  assign new_n2631_ = new_n1164_ & ~new_n2630_;
  assign new_n2632_ = new_n1168_ & ~new_n2631_;
  assign new_n2633_ = new_n1172_ & ~new_n2632_;
  assign new_n2634_ = new_n1176_ & ~new_n2633_;
  assign new_n2635_ = new_n1180_ & ~new_n2634_;
  assign new_n2636_ = new_n1184_ & ~new_n2635_;
  assign new_n2637_ = new_n1188_ & ~new_n2636_;
  assign new_n2638_ = new_n1192_ & ~new_n2637_;
  assign new_n2639_ = new_n1196_ & ~new_n2638_;
  assign new_n2640_ = new_n1200_ & ~new_n2639_;
  assign new_n2641_ = new_n1204_ & ~new_n2640_;
  assign new_n2642_ = new_n1208_ & ~new_n2641_;
  assign new_n2643_ = new_n1212_ & ~new_n2642_;
  assign new_n2644_ = new_n1216_ & ~new_n2643_;
  assign new_n2645_ = new_n1220_ & ~new_n2644_;
  assign new_n2646_ = new_n1224_ & ~new_n2645_;
  assign new_n2647_ = new_n1228_ & ~new_n2646_;
  assign new_n2648_ = new_n1232_ & ~new_n2647_;
  assign new_n2649_ = new_n1236_ & ~new_n2648_;
  assign new_n2650_ = new_n1240_ & ~new_n2649_;
  assign new_n2651_ = new_n1244_ & ~new_n2650_;
  assign new_n2652_ = new_n1248_ & ~new_n2651_;
  assign new_n2653_ = new_n1252_ & ~new_n2652_;
  assign new_n2654_ = new_n1256_ & ~new_n2653_;
  assign new_n2655_ = new_n1260_ & ~new_n2654_;
  assign new_n2656_ = new_n1264_ & ~new_n2655_;
  assign new_n2657_ = new_n1268_ & ~new_n2656_;
  assign new_n2658_ = new_n1272_ & ~new_n2657_;
  assign new_n2659_ = new_n1276_ & ~new_n2658_;
  assign new_n2660_ = new_n1280_ & ~new_n2659_;
  assign new_n2661_ = new_n1284_ & ~new_n2660_;
  assign new_n2662_ = new_n1288_ & ~new_n2661_;
  assign new_n2663_ = new_n1292_ & ~new_n2662_;
  assign new_n2664_ = new_n1296_ & ~new_n2663_;
  assign new_n2665_ = new_n1300_ & ~new_n2664_;
  assign new_n2666_ = new_n1304_ & ~new_n2665_;
  assign new_n2667_ = new_n1308_ & ~new_n2666_;
  assign new_n2668_ = new_n1312_ & ~new_n2667_;
  assign new_n2669_ = new_n1316_ & ~new_n2668_;
  assign new_n2670_ = new_n1320_ & ~new_n2669_;
  assign new_n2671_ = new_n1324_ & ~new_n2670_;
  assign new_n2672_ = new_n1328_ & ~new_n2671_;
  assign new_n2673_ = new_n1332_ & ~new_n2672_;
  assign new_n2674_ = new_n1336_ & ~new_n2673_;
  assign new_n2675_ = new_n1340_ & ~new_n2674_;
  assign new_n2676_ = new_n1344_ & ~new_n2675_;
  assign new_n2677_ = new_n1348_ & ~new_n2676_;
  assign new_n2678_ = new_n1352_ & ~new_n2677_;
  assign new_n2679_ = new_n1356_ & ~new_n2678_;
  assign new_n2680_ = new_n1360_ & ~new_n2679_;
  assign new_n2681_ = new_n1364_ & ~new_n2680_;
  assign new_n2682_ = new_n1368_ & ~new_n2681_;
  assign new_n2683_ = new_n1372_ & ~new_n2682_;
  assign new_n2684_ = new_n1376_ & ~new_n2683_;
  assign new_n2685_ = new_n1380_ & ~new_n2684_;
  assign new_n2686_ = new_n1384_ & ~new_n2685_;
  assign new_n2687_ = new_n1388_ & ~new_n2686_;
  assign new_n2688_ = new_n1392_ & ~new_n2687_;
  assign new_n2689_ = new_n1396_ & ~new_n2688_;
  assign new_n2690_ = new_n1663_ & ~new_n2689_;
  assign new_n2691_ = new_n392_ & ~new_n2690_;
  assign new_n2692_ = new_n396_ & ~new_n2691_;
  assign new_n2693_ = new_n400_ & ~new_n2692_;
  assign new_n2694_ = new_n404_ & ~new_n2693_;
  assign new_n2695_ = new_n408_ & ~new_n2694_;
  assign new_n2696_ = new_n412_ & ~new_n2695_;
  assign new_n2697_ = new_n416_ & ~new_n2696_;
  assign new_n2698_ = new_n420_ & ~new_n2697_;
  assign new_n2699_ = new_n424_ & ~new_n2698_;
  assign new_n2700_ = \req[17]  & ~new_n426_;
  assign \grant[17]  = ~new_n2699_ & new_n2700_;
  assign new_n2702_ = new_n435_ & ~new_n770_;
  assign new_n2703_ = new_n440_ & ~new_n2702_;
  assign new_n2704_ = new_n444_ & ~new_n2703_;
  assign new_n2705_ = new_n448_ & ~new_n2704_;
  assign new_n2706_ = new_n452_ & ~new_n2705_;
  assign new_n2707_ = new_n456_ & ~new_n2706_;
  assign new_n2708_ = new_n460_ & ~new_n2707_;
  assign new_n2709_ = new_n464_ & ~new_n2708_;
  assign new_n2710_ = new_n468_ & ~new_n2709_;
  assign new_n2711_ = new_n472_ & ~new_n2710_;
  assign new_n2712_ = new_n476_ & ~new_n2711_;
  assign new_n2713_ = new_n480_ & ~new_n2712_;
  assign new_n2714_ = new_n484_ & ~new_n2713_;
  assign new_n2715_ = new_n488_ & ~new_n2714_;
  assign new_n2716_ = new_n492_ & ~new_n2715_;
  assign new_n2717_ = new_n496_ & ~new_n2716_;
  assign new_n2718_ = new_n500_ & ~new_n2717_;
  assign new_n2719_ = new_n504_ & ~new_n2718_;
  assign new_n2720_ = new_n508_ & ~new_n2719_;
  assign new_n2721_ = new_n512_ & ~new_n2720_;
  assign new_n2722_ = new_n516_ & ~new_n2721_;
  assign new_n2723_ = new_n520_ & ~new_n2722_;
  assign new_n2724_ = new_n524_ & ~new_n2723_;
  assign new_n2725_ = new_n528_ & ~new_n2724_;
  assign new_n2726_ = new_n532_ & ~new_n2725_;
  assign new_n2727_ = new_n536_ & ~new_n2726_;
  assign new_n2728_ = new_n540_ & ~new_n2727_;
  assign new_n2729_ = new_n544_ & ~new_n2728_;
  assign new_n2730_ = new_n548_ & ~new_n2729_;
  assign new_n2731_ = new_n552_ & ~new_n2730_;
  assign new_n2732_ = new_n556_ & ~new_n2731_;
  assign new_n2733_ = new_n560_ & ~new_n2732_;
  assign new_n2734_ = new_n564_ & ~new_n2733_;
  assign new_n2735_ = new_n568_ & ~new_n2734_;
  assign new_n2736_ = new_n572_ & ~new_n2735_;
  assign new_n2737_ = new_n576_ & ~new_n2736_;
  assign new_n2738_ = new_n580_ & ~new_n2737_;
  assign new_n2739_ = new_n584_ & ~new_n2738_;
  assign new_n2740_ = new_n588_ & ~new_n2739_;
  assign new_n2741_ = new_n592_ & ~new_n2740_;
  assign new_n2742_ = new_n596_ & ~new_n2741_;
  assign new_n2743_ = new_n600_ & ~new_n2742_;
  assign new_n2744_ = new_n604_ & ~new_n2743_;
  assign new_n2745_ = new_n608_ & ~new_n2744_;
  assign new_n2746_ = new_n612_ & ~new_n2745_;
  assign new_n2747_ = new_n616_ & ~new_n2746_;
  assign new_n2748_ = new_n620_ & ~new_n2747_;
  assign new_n2749_ = new_n624_ & ~new_n2748_;
  assign new_n2750_ = new_n628_ & ~new_n2749_;
  assign new_n2751_ = new_n632_ & ~new_n2750_;
  assign new_n2752_ = new_n636_ & ~new_n2751_;
  assign new_n2753_ = new_n640_ & ~new_n2752_;
  assign new_n2754_ = new_n644_ & ~new_n2753_;
  assign new_n2755_ = new_n648_ & ~new_n2754_;
  assign new_n2756_ = new_n652_ & ~new_n2755_;
  assign new_n2757_ = new_n656_ & ~new_n2756_;
  assign new_n2758_ = new_n660_ & ~new_n2757_;
  assign new_n2759_ = new_n664_ & ~new_n2758_;
  assign new_n2760_ = new_n668_ & ~new_n2759_;
  assign new_n2761_ = new_n672_ & ~new_n2760_;
  assign new_n2762_ = new_n676_ & ~new_n2761_;
  assign new_n2763_ = new_n680_ & ~new_n2762_;
  assign new_n2764_ = new_n684_ & ~new_n2763_;
  assign new_n2765_ = new_n688_ & ~new_n2764_;
  assign new_n2766_ = new_n692_ & ~new_n2765_;
  assign new_n2767_ = new_n696_ & ~new_n2766_;
  assign new_n2768_ = new_n700_ & ~new_n2767_;
  assign new_n2769_ = new_n704_ & ~new_n2768_;
  assign new_n2770_ = new_n708_ & ~new_n2769_;
  assign new_n2771_ = new_n712_ & ~new_n2770_;
  assign new_n2772_ = new_n716_ & ~new_n2771_;
  assign new_n2773_ = new_n720_ & ~new_n2772_;
  assign new_n2774_ = new_n1484_ & ~new_n2773_;
  assign new_n2775_ = new_n1486_ & ~new_n2774_;
  assign new_n2776_ = new_n1750_ & ~new_n2775_;
  assign new_n2777_ = new_n731_ & ~new_n2776_;
  assign new_n2778_ = new_n735_ & ~new_n2777_;
  assign new_n2779_ = new_n739_ & ~new_n2778_;
  assign new_n2780_ = new_n743_ & ~new_n2779_;
  assign new_n2781_ = new_n747_ & ~new_n2780_;
  assign new_n2782_ = new_n751_ & ~new_n2781_;
  assign new_n2783_ = new_n755_ & ~new_n2782_;
  assign new_n2784_ = new_n759_ & ~new_n2783_;
  assign new_n2785_ = new_n763_ & ~new_n2784_;
  assign new_n2786_ = \req[18]  & ~new_n765_;
  assign \grant[18]  = ~new_n2785_ & new_n2786_;
  assign new_n2788_ = new_n774_ & ~new_n1107_;
  assign new_n2789_ = new_n779_ & ~new_n2788_;
  assign new_n2790_ = new_n783_ & ~new_n2789_;
  assign new_n2791_ = new_n787_ & ~new_n2790_;
  assign new_n2792_ = new_n791_ & ~new_n2791_;
  assign new_n2793_ = new_n795_ & ~new_n2792_;
  assign new_n2794_ = new_n799_ & ~new_n2793_;
  assign new_n2795_ = new_n803_ & ~new_n2794_;
  assign new_n2796_ = new_n807_ & ~new_n2795_;
  assign new_n2797_ = new_n811_ & ~new_n2796_;
  assign new_n2798_ = new_n815_ & ~new_n2797_;
  assign new_n2799_ = new_n819_ & ~new_n2798_;
  assign new_n2800_ = new_n823_ & ~new_n2799_;
  assign new_n2801_ = new_n827_ & ~new_n2800_;
  assign new_n2802_ = new_n831_ & ~new_n2801_;
  assign new_n2803_ = new_n835_ & ~new_n2802_;
  assign new_n2804_ = new_n839_ & ~new_n2803_;
  assign new_n2805_ = new_n843_ & ~new_n2804_;
  assign new_n2806_ = new_n847_ & ~new_n2805_;
  assign new_n2807_ = new_n851_ & ~new_n2806_;
  assign new_n2808_ = new_n855_ & ~new_n2807_;
  assign new_n2809_ = new_n859_ & ~new_n2808_;
  assign new_n2810_ = new_n863_ & ~new_n2809_;
  assign new_n2811_ = new_n867_ & ~new_n2810_;
  assign new_n2812_ = new_n871_ & ~new_n2811_;
  assign new_n2813_ = new_n875_ & ~new_n2812_;
  assign new_n2814_ = new_n879_ & ~new_n2813_;
  assign new_n2815_ = new_n883_ & ~new_n2814_;
  assign new_n2816_ = new_n887_ & ~new_n2815_;
  assign new_n2817_ = new_n891_ & ~new_n2816_;
  assign new_n2818_ = new_n895_ & ~new_n2817_;
  assign new_n2819_ = new_n899_ & ~new_n2818_;
  assign new_n2820_ = new_n903_ & ~new_n2819_;
  assign new_n2821_ = new_n907_ & ~new_n2820_;
  assign new_n2822_ = new_n911_ & ~new_n2821_;
  assign new_n2823_ = new_n915_ & ~new_n2822_;
  assign new_n2824_ = new_n919_ & ~new_n2823_;
  assign new_n2825_ = new_n923_ & ~new_n2824_;
  assign new_n2826_ = new_n927_ & ~new_n2825_;
  assign new_n2827_ = new_n931_ & ~new_n2826_;
  assign new_n2828_ = new_n935_ & ~new_n2827_;
  assign new_n2829_ = new_n939_ & ~new_n2828_;
  assign new_n2830_ = new_n943_ & ~new_n2829_;
  assign new_n2831_ = new_n947_ & ~new_n2830_;
  assign new_n2832_ = new_n951_ & ~new_n2831_;
  assign new_n2833_ = new_n955_ & ~new_n2832_;
  assign new_n2834_ = new_n959_ & ~new_n2833_;
  assign new_n2835_ = new_n963_ & ~new_n2834_;
  assign new_n2836_ = new_n967_ & ~new_n2835_;
  assign new_n2837_ = new_n971_ & ~new_n2836_;
  assign new_n2838_ = new_n975_ & ~new_n2837_;
  assign new_n2839_ = new_n979_ & ~new_n2838_;
  assign new_n2840_ = new_n983_ & ~new_n2839_;
  assign new_n2841_ = new_n987_ & ~new_n2840_;
  assign new_n2842_ = new_n991_ & ~new_n2841_;
  assign new_n2843_ = new_n995_ & ~new_n2842_;
  assign new_n2844_ = new_n999_ & ~new_n2843_;
  assign new_n2845_ = new_n1003_ & ~new_n2844_;
  assign new_n2846_ = new_n1007_ & ~new_n2845_;
  assign new_n2847_ = new_n1011_ & ~new_n2846_;
  assign new_n2848_ = new_n1015_ & ~new_n2847_;
  assign new_n2849_ = new_n1019_ & ~new_n2848_;
  assign new_n2850_ = new_n1023_ & ~new_n2849_;
  assign new_n2851_ = new_n1027_ & ~new_n2850_;
  assign new_n2852_ = new_n1031_ & ~new_n2851_;
  assign new_n2853_ = new_n1035_ & ~new_n2852_;
  assign new_n2854_ = new_n1039_ & ~new_n2853_;
  assign new_n2855_ = new_n1043_ & ~new_n2854_;
  assign new_n2856_ = new_n1047_ & ~new_n2855_;
  assign new_n2857_ = new_n1051_ & ~new_n2856_;
  assign new_n2858_ = new_n1055_ & ~new_n2857_;
  assign new_n2859_ = new_n1059_ & ~new_n2858_;
  assign new_n2860_ = new_n1574_ & ~new_n2859_;
  assign new_n2861_ = new_n1576_ & ~new_n2860_;
  assign new_n2862_ = new_n1837_ & ~new_n2861_;
  assign new_n2863_ = new_n1068_ & ~new_n2862_;
  assign new_n2864_ = new_n1072_ & ~new_n2863_;
  assign new_n2865_ = new_n1076_ & ~new_n2864_;
  assign new_n2866_ = new_n1080_ & ~new_n2865_;
  assign new_n2867_ = new_n1084_ & ~new_n2866_;
  assign new_n2868_ = new_n1088_ & ~new_n2867_;
  assign new_n2869_ = new_n1092_ & ~new_n2868_;
  assign new_n2870_ = new_n1096_ & ~new_n2869_;
  assign new_n2871_ = new_n1100_ & ~new_n2870_;
  assign new_n2872_ = \req[19]  & ~new_n1102_;
  assign \grant[19]  = ~new_n2871_ & new_n2872_;
  assign new_n2874_ = ~new_n439_ & new_n1111_;
  assign new_n2875_ = new_n1116_ & ~new_n2874_;
  assign new_n2876_ = new_n1120_ & ~new_n2875_;
  assign new_n2877_ = new_n1124_ & ~new_n2876_;
  assign new_n2878_ = new_n1128_ & ~new_n2877_;
  assign new_n2879_ = new_n1132_ & ~new_n2878_;
  assign new_n2880_ = new_n1136_ & ~new_n2879_;
  assign new_n2881_ = new_n1140_ & ~new_n2880_;
  assign new_n2882_ = new_n1144_ & ~new_n2881_;
  assign new_n2883_ = new_n1148_ & ~new_n2882_;
  assign new_n2884_ = new_n1152_ & ~new_n2883_;
  assign new_n2885_ = new_n1156_ & ~new_n2884_;
  assign new_n2886_ = new_n1160_ & ~new_n2885_;
  assign new_n2887_ = new_n1164_ & ~new_n2886_;
  assign new_n2888_ = new_n1168_ & ~new_n2887_;
  assign new_n2889_ = new_n1172_ & ~new_n2888_;
  assign new_n2890_ = new_n1176_ & ~new_n2889_;
  assign new_n2891_ = new_n1180_ & ~new_n2890_;
  assign new_n2892_ = new_n1184_ & ~new_n2891_;
  assign new_n2893_ = new_n1188_ & ~new_n2892_;
  assign new_n2894_ = new_n1192_ & ~new_n2893_;
  assign new_n2895_ = new_n1196_ & ~new_n2894_;
  assign new_n2896_ = new_n1200_ & ~new_n2895_;
  assign new_n2897_ = new_n1204_ & ~new_n2896_;
  assign new_n2898_ = new_n1208_ & ~new_n2897_;
  assign new_n2899_ = new_n1212_ & ~new_n2898_;
  assign new_n2900_ = new_n1216_ & ~new_n2899_;
  assign new_n2901_ = new_n1220_ & ~new_n2900_;
  assign new_n2902_ = new_n1224_ & ~new_n2901_;
  assign new_n2903_ = new_n1228_ & ~new_n2902_;
  assign new_n2904_ = new_n1232_ & ~new_n2903_;
  assign new_n2905_ = new_n1236_ & ~new_n2904_;
  assign new_n2906_ = new_n1240_ & ~new_n2905_;
  assign new_n2907_ = new_n1244_ & ~new_n2906_;
  assign new_n2908_ = new_n1248_ & ~new_n2907_;
  assign new_n2909_ = new_n1252_ & ~new_n2908_;
  assign new_n2910_ = new_n1256_ & ~new_n2909_;
  assign new_n2911_ = new_n1260_ & ~new_n2910_;
  assign new_n2912_ = new_n1264_ & ~new_n2911_;
  assign new_n2913_ = new_n1268_ & ~new_n2912_;
  assign new_n2914_ = new_n1272_ & ~new_n2913_;
  assign new_n2915_ = new_n1276_ & ~new_n2914_;
  assign new_n2916_ = new_n1280_ & ~new_n2915_;
  assign new_n2917_ = new_n1284_ & ~new_n2916_;
  assign new_n2918_ = new_n1288_ & ~new_n2917_;
  assign new_n2919_ = new_n1292_ & ~new_n2918_;
  assign new_n2920_ = new_n1296_ & ~new_n2919_;
  assign new_n2921_ = new_n1300_ & ~new_n2920_;
  assign new_n2922_ = new_n1304_ & ~new_n2921_;
  assign new_n2923_ = new_n1308_ & ~new_n2922_;
  assign new_n2924_ = new_n1312_ & ~new_n2923_;
  assign new_n2925_ = new_n1316_ & ~new_n2924_;
  assign new_n2926_ = new_n1320_ & ~new_n2925_;
  assign new_n2927_ = new_n1324_ & ~new_n2926_;
  assign new_n2928_ = new_n1328_ & ~new_n2927_;
  assign new_n2929_ = new_n1332_ & ~new_n2928_;
  assign new_n2930_ = new_n1336_ & ~new_n2929_;
  assign new_n2931_ = new_n1340_ & ~new_n2930_;
  assign new_n2932_ = new_n1344_ & ~new_n2931_;
  assign new_n2933_ = new_n1348_ & ~new_n2932_;
  assign new_n2934_ = new_n1352_ & ~new_n2933_;
  assign new_n2935_ = new_n1356_ & ~new_n2934_;
  assign new_n2936_ = new_n1360_ & ~new_n2935_;
  assign new_n2937_ = new_n1364_ & ~new_n2936_;
  assign new_n2938_ = new_n1368_ & ~new_n2937_;
  assign new_n2939_ = new_n1372_ & ~new_n2938_;
  assign new_n2940_ = new_n1376_ & ~new_n2939_;
  assign new_n2941_ = new_n1380_ & ~new_n2940_;
  assign new_n2942_ = new_n1384_ & ~new_n2941_;
  assign new_n2943_ = new_n1388_ & ~new_n2942_;
  assign new_n2944_ = new_n1392_ & ~new_n2943_;
  assign new_n2945_ = new_n1396_ & ~new_n2944_;
  assign new_n2946_ = new_n1663_ & ~new_n2945_;
  assign new_n2947_ = new_n392_ & ~new_n2946_;
  assign new_n2948_ = new_n396_ & ~new_n2947_;
  assign new_n2949_ = new_n400_ & ~new_n2948_;
  assign new_n2950_ = new_n404_ & ~new_n2949_;
  assign new_n2951_ = new_n408_ & ~new_n2950_;
  assign new_n2952_ = new_n412_ & ~new_n2951_;
  assign new_n2953_ = new_n416_ & ~new_n2952_;
  assign new_n2954_ = new_n420_ & ~new_n2953_;
  assign new_n2955_ = new_n424_ & ~new_n2954_;
  assign new_n2956_ = new_n428_ & ~new_n2955_;
  assign new_n2957_ = new_n432_ & ~new_n2956_;
  assign new_n2958_ = \req[20]  & ~new_n434_;
  assign \grant[20]  = ~new_n2957_ & new_n2958_;
  assign new_n2960_ = new_n443_ & ~new_n778_;
  assign new_n2961_ = new_n448_ & ~new_n2960_;
  assign new_n2962_ = new_n452_ & ~new_n2961_;
  assign new_n2963_ = new_n456_ & ~new_n2962_;
  assign new_n2964_ = new_n460_ & ~new_n2963_;
  assign new_n2965_ = new_n464_ & ~new_n2964_;
  assign new_n2966_ = new_n468_ & ~new_n2965_;
  assign new_n2967_ = new_n472_ & ~new_n2966_;
  assign new_n2968_ = new_n476_ & ~new_n2967_;
  assign new_n2969_ = new_n480_ & ~new_n2968_;
  assign new_n2970_ = new_n484_ & ~new_n2969_;
  assign new_n2971_ = new_n488_ & ~new_n2970_;
  assign new_n2972_ = new_n492_ & ~new_n2971_;
  assign new_n2973_ = new_n496_ & ~new_n2972_;
  assign new_n2974_ = new_n500_ & ~new_n2973_;
  assign new_n2975_ = new_n504_ & ~new_n2974_;
  assign new_n2976_ = new_n508_ & ~new_n2975_;
  assign new_n2977_ = new_n512_ & ~new_n2976_;
  assign new_n2978_ = new_n516_ & ~new_n2977_;
  assign new_n2979_ = new_n520_ & ~new_n2978_;
  assign new_n2980_ = new_n524_ & ~new_n2979_;
  assign new_n2981_ = new_n528_ & ~new_n2980_;
  assign new_n2982_ = new_n532_ & ~new_n2981_;
  assign new_n2983_ = new_n536_ & ~new_n2982_;
  assign new_n2984_ = new_n540_ & ~new_n2983_;
  assign new_n2985_ = new_n544_ & ~new_n2984_;
  assign new_n2986_ = new_n548_ & ~new_n2985_;
  assign new_n2987_ = new_n552_ & ~new_n2986_;
  assign new_n2988_ = new_n556_ & ~new_n2987_;
  assign new_n2989_ = new_n560_ & ~new_n2988_;
  assign new_n2990_ = new_n564_ & ~new_n2989_;
  assign new_n2991_ = new_n568_ & ~new_n2990_;
  assign new_n2992_ = new_n572_ & ~new_n2991_;
  assign new_n2993_ = new_n576_ & ~new_n2992_;
  assign new_n2994_ = new_n580_ & ~new_n2993_;
  assign new_n2995_ = new_n584_ & ~new_n2994_;
  assign new_n2996_ = new_n588_ & ~new_n2995_;
  assign new_n2997_ = new_n592_ & ~new_n2996_;
  assign new_n2998_ = new_n596_ & ~new_n2997_;
  assign new_n2999_ = new_n600_ & ~new_n2998_;
  assign new_n3000_ = new_n604_ & ~new_n2999_;
  assign new_n3001_ = new_n608_ & ~new_n3000_;
  assign new_n3002_ = new_n612_ & ~new_n3001_;
  assign new_n3003_ = new_n616_ & ~new_n3002_;
  assign new_n3004_ = new_n620_ & ~new_n3003_;
  assign new_n3005_ = new_n624_ & ~new_n3004_;
  assign new_n3006_ = new_n628_ & ~new_n3005_;
  assign new_n3007_ = new_n632_ & ~new_n3006_;
  assign new_n3008_ = new_n636_ & ~new_n3007_;
  assign new_n3009_ = new_n640_ & ~new_n3008_;
  assign new_n3010_ = new_n644_ & ~new_n3009_;
  assign new_n3011_ = new_n648_ & ~new_n3010_;
  assign new_n3012_ = new_n652_ & ~new_n3011_;
  assign new_n3013_ = new_n656_ & ~new_n3012_;
  assign new_n3014_ = new_n660_ & ~new_n3013_;
  assign new_n3015_ = new_n664_ & ~new_n3014_;
  assign new_n3016_ = new_n668_ & ~new_n3015_;
  assign new_n3017_ = new_n672_ & ~new_n3016_;
  assign new_n3018_ = new_n676_ & ~new_n3017_;
  assign new_n3019_ = new_n680_ & ~new_n3018_;
  assign new_n3020_ = new_n684_ & ~new_n3019_;
  assign new_n3021_ = new_n688_ & ~new_n3020_;
  assign new_n3022_ = new_n692_ & ~new_n3021_;
  assign new_n3023_ = new_n696_ & ~new_n3022_;
  assign new_n3024_ = new_n700_ & ~new_n3023_;
  assign new_n3025_ = new_n704_ & ~new_n3024_;
  assign new_n3026_ = new_n708_ & ~new_n3025_;
  assign new_n3027_ = new_n712_ & ~new_n3026_;
  assign new_n3028_ = new_n716_ & ~new_n3027_;
  assign new_n3029_ = new_n720_ & ~new_n3028_;
  assign new_n3030_ = new_n1484_ & ~new_n3029_;
  assign new_n3031_ = new_n1486_ & ~new_n3030_;
  assign new_n3032_ = new_n1750_ & ~new_n3031_;
  assign new_n3033_ = new_n731_ & ~new_n3032_;
  assign new_n3034_ = new_n735_ & ~new_n3033_;
  assign new_n3035_ = new_n739_ & ~new_n3034_;
  assign new_n3036_ = new_n743_ & ~new_n3035_;
  assign new_n3037_ = new_n747_ & ~new_n3036_;
  assign new_n3038_ = new_n751_ & ~new_n3037_;
  assign new_n3039_ = new_n755_ & ~new_n3038_;
  assign new_n3040_ = new_n759_ & ~new_n3039_;
  assign new_n3041_ = new_n763_ & ~new_n3040_;
  assign new_n3042_ = new_n767_ & ~new_n3041_;
  assign new_n3043_ = new_n771_ & ~new_n3042_;
  assign new_n3044_ = \req[21]  & ~new_n773_;
  assign \grant[21]  = ~new_n3043_ & new_n3044_;
  assign new_n3046_ = new_n782_ & ~new_n1115_;
  assign new_n3047_ = new_n787_ & ~new_n3046_;
  assign new_n3048_ = new_n791_ & ~new_n3047_;
  assign new_n3049_ = new_n795_ & ~new_n3048_;
  assign new_n3050_ = new_n799_ & ~new_n3049_;
  assign new_n3051_ = new_n803_ & ~new_n3050_;
  assign new_n3052_ = new_n807_ & ~new_n3051_;
  assign new_n3053_ = new_n811_ & ~new_n3052_;
  assign new_n3054_ = new_n815_ & ~new_n3053_;
  assign new_n3055_ = new_n819_ & ~new_n3054_;
  assign new_n3056_ = new_n823_ & ~new_n3055_;
  assign new_n3057_ = new_n827_ & ~new_n3056_;
  assign new_n3058_ = new_n831_ & ~new_n3057_;
  assign new_n3059_ = new_n835_ & ~new_n3058_;
  assign new_n3060_ = new_n839_ & ~new_n3059_;
  assign new_n3061_ = new_n843_ & ~new_n3060_;
  assign new_n3062_ = new_n847_ & ~new_n3061_;
  assign new_n3063_ = new_n851_ & ~new_n3062_;
  assign new_n3064_ = new_n855_ & ~new_n3063_;
  assign new_n3065_ = new_n859_ & ~new_n3064_;
  assign new_n3066_ = new_n863_ & ~new_n3065_;
  assign new_n3067_ = new_n867_ & ~new_n3066_;
  assign new_n3068_ = new_n871_ & ~new_n3067_;
  assign new_n3069_ = new_n875_ & ~new_n3068_;
  assign new_n3070_ = new_n879_ & ~new_n3069_;
  assign new_n3071_ = new_n883_ & ~new_n3070_;
  assign new_n3072_ = new_n887_ & ~new_n3071_;
  assign new_n3073_ = new_n891_ & ~new_n3072_;
  assign new_n3074_ = new_n895_ & ~new_n3073_;
  assign new_n3075_ = new_n899_ & ~new_n3074_;
  assign new_n3076_ = new_n903_ & ~new_n3075_;
  assign new_n3077_ = new_n907_ & ~new_n3076_;
  assign new_n3078_ = new_n911_ & ~new_n3077_;
  assign new_n3079_ = new_n915_ & ~new_n3078_;
  assign new_n3080_ = new_n919_ & ~new_n3079_;
  assign new_n3081_ = new_n923_ & ~new_n3080_;
  assign new_n3082_ = new_n927_ & ~new_n3081_;
  assign new_n3083_ = new_n931_ & ~new_n3082_;
  assign new_n3084_ = new_n935_ & ~new_n3083_;
  assign new_n3085_ = new_n939_ & ~new_n3084_;
  assign new_n3086_ = new_n943_ & ~new_n3085_;
  assign new_n3087_ = new_n947_ & ~new_n3086_;
  assign new_n3088_ = new_n951_ & ~new_n3087_;
  assign new_n3089_ = new_n955_ & ~new_n3088_;
  assign new_n3090_ = new_n959_ & ~new_n3089_;
  assign new_n3091_ = new_n963_ & ~new_n3090_;
  assign new_n3092_ = new_n967_ & ~new_n3091_;
  assign new_n3093_ = new_n971_ & ~new_n3092_;
  assign new_n3094_ = new_n975_ & ~new_n3093_;
  assign new_n3095_ = new_n979_ & ~new_n3094_;
  assign new_n3096_ = new_n983_ & ~new_n3095_;
  assign new_n3097_ = new_n987_ & ~new_n3096_;
  assign new_n3098_ = new_n991_ & ~new_n3097_;
  assign new_n3099_ = new_n995_ & ~new_n3098_;
  assign new_n3100_ = new_n999_ & ~new_n3099_;
  assign new_n3101_ = new_n1003_ & ~new_n3100_;
  assign new_n3102_ = new_n1007_ & ~new_n3101_;
  assign new_n3103_ = new_n1011_ & ~new_n3102_;
  assign new_n3104_ = new_n1015_ & ~new_n3103_;
  assign new_n3105_ = new_n1019_ & ~new_n3104_;
  assign new_n3106_ = new_n1023_ & ~new_n3105_;
  assign new_n3107_ = new_n1027_ & ~new_n3106_;
  assign new_n3108_ = new_n1031_ & ~new_n3107_;
  assign new_n3109_ = new_n1035_ & ~new_n3108_;
  assign new_n3110_ = new_n1039_ & ~new_n3109_;
  assign new_n3111_ = new_n1043_ & ~new_n3110_;
  assign new_n3112_ = new_n1047_ & ~new_n3111_;
  assign new_n3113_ = new_n1051_ & ~new_n3112_;
  assign new_n3114_ = new_n1055_ & ~new_n3113_;
  assign new_n3115_ = new_n1059_ & ~new_n3114_;
  assign new_n3116_ = new_n1574_ & ~new_n3115_;
  assign new_n3117_ = new_n1576_ & ~new_n3116_;
  assign new_n3118_ = new_n1837_ & ~new_n3117_;
  assign new_n3119_ = new_n1068_ & ~new_n3118_;
  assign new_n3120_ = new_n1072_ & ~new_n3119_;
  assign new_n3121_ = new_n1076_ & ~new_n3120_;
  assign new_n3122_ = new_n1080_ & ~new_n3121_;
  assign new_n3123_ = new_n1084_ & ~new_n3122_;
  assign new_n3124_ = new_n1088_ & ~new_n3123_;
  assign new_n3125_ = new_n1092_ & ~new_n3124_;
  assign new_n3126_ = new_n1096_ & ~new_n3125_;
  assign new_n3127_ = new_n1100_ & ~new_n3126_;
  assign new_n3128_ = new_n1104_ & ~new_n3127_;
  assign new_n3129_ = new_n1108_ & ~new_n3128_;
  assign new_n3130_ = \req[22]  & ~new_n1110_;
  assign \grant[22]  = ~new_n3129_ & new_n3130_;
  assign new_n3132_ = ~new_n447_ & new_n1119_;
  assign new_n3133_ = new_n1124_ & ~new_n3132_;
  assign new_n3134_ = new_n1128_ & ~new_n3133_;
  assign new_n3135_ = new_n1132_ & ~new_n3134_;
  assign new_n3136_ = new_n1136_ & ~new_n3135_;
  assign new_n3137_ = new_n1140_ & ~new_n3136_;
  assign new_n3138_ = new_n1144_ & ~new_n3137_;
  assign new_n3139_ = new_n1148_ & ~new_n3138_;
  assign new_n3140_ = new_n1152_ & ~new_n3139_;
  assign new_n3141_ = new_n1156_ & ~new_n3140_;
  assign new_n3142_ = new_n1160_ & ~new_n3141_;
  assign new_n3143_ = new_n1164_ & ~new_n3142_;
  assign new_n3144_ = new_n1168_ & ~new_n3143_;
  assign new_n3145_ = new_n1172_ & ~new_n3144_;
  assign new_n3146_ = new_n1176_ & ~new_n3145_;
  assign new_n3147_ = new_n1180_ & ~new_n3146_;
  assign new_n3148_ = new_n1184_ & ~new_n3147_;
  assign new_n3149_ = new_n1188_ & ~new_n3148_;
  assign new_n3150_ = new_n1192_ & ~new_n3149_;
  assign new_n3151_ = new_n1196_ & ~new_n3150_;
  assign new_n3152_ = new_n1200_ & ~new_n3151_;
  assign new_n3153_ = new_n1204_ & ~new_n3152_;
  assign new_n3154_ = new_n1208_ & ~new_n3153_;
  assign new_n3155_ = new_n1212_ & ~new_n3154_;
  assign new_n3156_ = new_n1216_ & ~new_n3155_;
  assign new_n3157_ = new_n1220_ & ~new_n3156_;
  assign new_n3158_ = new_n1224_ & ~new_n3157_;
  assign new_n3159_ = new_n1228_ & ~new_n3158_;
  assign new_n3160_ = new_n1232_ & ~new_n3159_;
  assign new_n3161_ = new_n1236_ & ~new_n3160_;
  assign new_n3162_ = new_n1240_ & ~new_n3161_;
  assign new_n3163_ = new_n1244_ & ~new_n3162_;
  assign new_n3164_ = new_n1248_ & ~new_n3163_;
  assign new_n3165_ = new_n1252_ & ~new_n3164_;
  assign new_n3166_ = new_n1256_ & ~new_n3165_;
  assign new_n3167_ = new_n1260_ & ~new_n3166_;
  assign new_n3168_ = new_n1264_ & ~new_n3167_;
  assign new_n3169_ = new_n1268_ & ~new_n3168_;
  assign new_n3170_ = new_n1272_ & ~new_n3169_;
  assign new_n3171_ = new_n1276_ & ~new_n3170_;
  assign new_n3172_ = new_n1280_ & ~new_n3171_;
  assign new_n3173_ = new_n1284_ & ~new_n3172_;
  assign new_n3174_ = new_n1288_ & ~new_n3173_;
  assign new_n3175_ = new_n1292_ & ~new_n3174_;
  assign new_n3176_ = new_n1296_ & ~new_n3175_;
  assign new_n3177_ = new_n1300_ & ~new_n3176_;
  assign new_n3178_ = new_n1304_ & ~new_n3177_;
  assign new_n3179_ = new_n1308_ & ~new_n3178_;
  assign new_n3180_ = new_n1312_ & ~new_n3179_;
  assign new_n3181_ = new_n1316_ & ~new_n3180_;
  assign new_n3182_ = new_n1320_ & ~new_n3181_;
  assign new_n3183_ = new_n1324_ & ~new_n3182_;
  assign new_n3184_ = new_n1328_ & ~new_n3183_;
  assign new_n3185_ = new_n1332_ & ~new_n3184_;
  assign new_n3186_ = new_n1336_ & ~new_n3185_;
  assign new_n3187_ = new_n1340_ & ~new_n3186_;
  assign new_n3188_ = new_n1344_ & ~new_n3187_;
  assign new_n3189_ = new_n1348_ & ~new_n3188_;
  assign new_n3190_ = new_n1352_ & ~new_n3189_;
  assign new_n3191_ = new_n1356_ & ~new_n3190_;
  assign new_n3192_ = new_n1360_ & ~new_n3191_;
  assign new_n3193_ = new_n1364_ & ~new_n3192_;
  assign new_n3194_ = new_n1368_ & ~new_n3193_;
  assign new_n3195_ = new_n1372_ & ~new_n3194_;
  assign new_n3196_ = new_n1376_ & ~new_n3195_;
  assign new_n3197_ = new_n1380_ & ~new_n3196_;
  assign new_n3198_ = new_n1384_ & ~new_n3197_;
  assign new_n3199_ = new_n1388_ & ~new_n3198_;
  assign new_n3200_ = new_n1392_ & ~new_n3199_;
  assign new_n3201_ = new_n1396_ & ~new_n3200_;
  assign new_n3202_ = new_n1663_ & ~new_n3201_;
  assign new_n3203_ = new_n392_ & ~new_n3202_;
  assign new_n3204_ = new_n396_ & ~new_n3203_;
  assign new_n3205_ = new_n400_ & ~new_n3204_;
  assign new_n3206_ = new_n404_ & ~new_n3205_;
  assign new_n3207_ = new_n408_ & ~new_n3206_;
  assign new_n3208_ = new_n412_ & ~new_n3207_;
  assign new_n3209_ = new_n416_ & ~new_n3208_;
  assign new_n3210_ = new_n420_ & ~new_n3209_;
  assign new_n3211_ = new_n424_ & ~new_n3210_;
  assign new_n3212_ = new_n428_ & ~new_n3211_;
  assign new_n3213_ = new_n432_ & ~new_n3212_;
  assign new_n3214_ = new_n436_ & ~new_n3213_;
  assign new_n3215_ = new_n440_ & ~new_n3214_;
  assign new_n3216_ = \req[23]  & ~new_n442_;
  assign \grant[23]  = ~new_n3215_ & new_n3216_;
  assign new_n3218_ = new_n451_ & ~new_n786_;
  assign new_n3219_ = new_n456_ & ~new_n3218_;
  assign new_n3220_ = new_n460_ & ~new_n3219_;
  assign new_n3221_ = new_n464_ & ~new_n3220_;
  assign new_n3222_ = new_n468_ & ~new_n3221_;
  assign new_n3223_ = new_n472_ & ~new_n3222_;
  assign new_n3224_ = new_n476_ & ~new_n3223_;
  assign new_n3225_ = new_n480_ & ~new_n3224_;
  assign new_n3226_ = new_n484_ & ~new_n3225_;
  assign new_n3227_ = new_n488_ & ~new_n3226_;
  assign new_n3228_ = new_n492_ & ~new_n3227_;
  assign new_n3229_ = new_n496_ & ~new_n3228_;
  assign new_n3230_ = new_n500_ & ~new_n3229_;
  assign new_n3231_ = new_n504_ & ~new_n3230_;
  assign new_n3232_ = new_n508_ & ~new_n3231_;
  assign new_n3233_ = new_n512_ & ~new_n3232_;
  assign new_n3234_ = new_n516_ & ~new_n3233_;
  assign new_n3235_ = new_n520_ & ~new_n3234_;
  assign new_n3236_ = new_n524_ & ~new_n3235_;
  assign new_n3237_ = new_n528_ & ~new_n3236_;
  assign new_n3238_ = new_n532_ & ~new_n3237_;
  assign new_n3239_ = new_n536_ & ~new_n3238_;
  assign new_n3240_ = new_n540_ & ~new_n3239_;
  assign new_n3241_ = new_n544_ & ~new_n3240_;
  assign new_n3242_ = new_n548_ & ~new_n3241_;
  assign new_n3243_ = new_n552_ & ~new_n3242_;
  assign new_n3244_ = new_n556_ & ~new_n3243_;
  assign new_n3245_ = new_n560_ & ~new_n3244_;
  assign new_n3246_ = new_n564_ & ~new_n3245_;
  assign new_n3247_ = new_n568_ & ~new_n3246_;
  assign new_n3248_ = new_n572_ & ~new_n3247_;
  assign new_n3249_ = new_n576_ & ~new_n3248_;
  assign new_n3250_ = new_n580_ & ~new_n3249_;
  assign new_n3251_ = new_n584_ & ~new_n3250_;
  assign new_n3252_ = new_n588_ & ~new_n3251_;
  assign new_n3253_ = new_n592_ & ~new_n3252_;
  assign new_n3254_ = new_n596_ & ~new_n3253_;
  assign new_n3255_ = new_n600_ & ~new_n3254_;
  assign new_n3256_ = new_n604_ & ~new_n3255_;
  assign new_n3257_ = new_n608_ & ~new_n3256_;
  assign new_n3258_ = new_n612_ & ~new_n3257_;
  assign new_n3259_ = new_n616_ & ~new_n3258_;
  assign new_n3260_ = new_n620_ & ~new_n3259_;
  assign new_n3261_ = new_n624_ & ~new_n3260_;
  assign new_n3262_ = new_n628_ & ~new_n3261_;
  assign new_n3263_ = new_n632_ & ~new_n3262_;
  assign new_n3264_ = new_n636_ & ~new_n3263_;
  assign new_n3265_ = new_n640_ & ~new_n3264_;
  assign new_n3266_ = new_n644_ & ~new_n3265_;
  assign new_n3267_ = new_n648_ & ~new_n3266_;
  assign new_n3268_ = new_n652_ & ~new_n3267_;
  assign new_n3269_ = new_n656_ & ~new_n3268_;
  assign new_n3270_ = new_n660_ & ~new_n3269_;
  assign new_n3271_ = new_n664_ & ~new_n3270_;
  assign new_n3272_ = new_n668_ & ~new_n3271_;
  assign new_n3273_ = new_n672_ & ~new_n3272_;
  assign new_n3274_ = new_n676_ & ~new_n3273_;
  assign new_n3275_ = new_n680_ & ~new_n3274_;
  assign new_n3276_ = new_n684_ & ~new_n3275_;
  assign new_n3277_ = new_n688_ & ~new_n3276_;
  assign new_n3278_ = new_n692_ & ~new_n3277_;
  assign new_n3279_ = new_n696_ & ~new_n3278_;
  assign new_n3280_ = new_n700_ & ~new_n3279_;
  assign new_n3281_ = new_n704_ & ~new_n3280_;
  assign new_n3282_ = new_n708_ & ~new_n3281_;
  assign new_n3283_ = new_n712_ & ~new_n3282_;
  assign new_n3284_ = new_n716_ & ~new_n3283_;
  assign new_n3285_ = new_n720_ & ~new_n3284_;
  assign new_n3286_ = new_n1484_ & ~new_n3285_;
  assign new_n3287_ = new_n1486_ & ~new_n3286_;
  assign new_n3288_ = new_n1750_ & ~new_n3287_;
  assign new_n3289_ = new_n731_ & ~new_n3288_;
  assign new_n3290_ = new_n735_ & ~new_n3289_;
  assign new_n3291_ = new_n739_ & ~new_n3290_;
  assign new_n3292_ = new_n743_ & ~new_n3291_;
  assign new_n3293_ = new_n747_ & ~new_n3292_;
  assign new_n3294_ = new_n751_ & ~new_n3293_;
  assign new_n3295_ = new_n755_ & ~new_n3294_;
  assign new_n3296_ = new_n759_ & ~new_n3295_;
  assign new_n3297_ = new_n763_ & ~new_n3296_;
  assign new_n3298_ = new_n767_ & ~new_n3297_;
  assign new_n3299_ = new_n771_ & ~new_n3298_;
  assign new_n3300_ = new_n775_ & ~new_n3299_;
  assign new_n3301_ = new_n779_ & ~new_n3300_;
  assign new_n3302_ = \req[24]  & ~new_n781_;
  assign \grant[24]  = ~new_n3301_ & new_n3302_;
  assign new_n3304_ = new_n790_ & ~new_n1123_;
  assign new_n3305_ = new_n795_ & ~new_n3304_;
  assign new_n3306_ = new_n799_ & ~new_n3305_;
  assign new_n3307_ = new_n803_ & ~new_n3306_;
  assign new_n3308_ = new_n807_ & ~new_n3307_;
  assign new_n3309_ = new_n811_ & ~new_n3308_;
  assign new_n3310_ = new_n815_ & ~new_n3309_;
  assign new_n3311_ = new_n819_ & ~new_n3310_;
  assign new_n3312_ = new_n823_ & ~new_n3311_;
  assign new_n3313_ = new_n827_ & ~new_n3312_;
  assign new_n3314_ = new_n831_ & ~new_n3313_;
  assign new_n3315_ = new_n835_ & ~new_n3314_;
  assign new_n3316_ = new_n839_ & ~new_n3315_;
  assign new_n3317_ = new_n843_ & ~new_n3316_;
  assign new_n3318_ = new_n847_ & ~new_n3317_;
  assign new_n3319_ = new_n851_ & ~new_n3318_;
  assign new_n3320_ = new_n855_ & ~new_n3319_;
  assign new_n3321_ = new_n859_ & ~new_n3320_;
  assign new_n3322_ = new_n863_ & ~new_n3321_;
  assign new_n3323_ = new_n867_ & ~new_n3322_;
  assign new_n3324_ = new_n871_ & ~new_n3323_;
  assign new_n3325_ = new_n875_ & ~new_n3324_;
  assign new_n3326_ = new_n879_ & ~new_n3325_;
  assign new_n3327_ = new_n883_ & ~new_n3326_;
  assign new_n3328_ = new_n887_ & ~new_n3327_;
  assign new_n3329_ = new_n891_ & ~new_n3328_;
  assign new_n3330_ = new_n895_ & ~new_n3329_;
  assign new_n3331_ = new_n899_ & ~new_n3330_;
  assign new_n3332_ = new_n903_ & ~new_n3331_;
  assign new_n3333_ = new_n907_ & ~new_n3332_;
  assign new_n3334_ = new_n911_ & ~new_n3333_;
  assign new_n3335_ = new_n915_ & ~new_n3334_;
  assign new_n3336_ = new_n919_ & ~new_n3335_;
  assign new_n3337_ = new_n923_ & ~new_n3336_;
  assign new_n3338_ = new_n927_ & ~new_n3337_;
  assign new_n3339_ = new_n931_ & ~new_n3338_;
  assign new_n3340_ = new_n935_ & ~new_n3339_;
  assign new_n3341_ = new_n939_ & ~new_n3340_;
  assign new_n3342_ = new_n943_ & ~new_n3341_;
  assign new_n3343_ = new_n947_ & ~new_n3342_;
  assign new_n3344_ = new_n951_ & ~new_n3343_;
  assign new_n3345_ = new_n955_ & ~new_n3344_;
  assign new_n3346_ = new_n959_ & ~new_n3345_;
  assign new_n3347_ = new_n963_ & ~new_n3346_;
  assign new_n3348_ = new_n967_ & ~new_n3347_;
  assign new_n3349_ = new_n971_ & ~new_n3348_;
  assign new_n3350_ = new_n975_ & ~new_n3349_;
  assign new_n3351_ = new_n979_ & ~new_n3350_;
  assign new_n3352_ = new_n983_ & ~new_n3351_;
  assign new_n3353_ = new_n987_ & ~new_n3352_;
  assign new_n3354_ = new_n991_ & ~new_n3353_;
  assign new_n3355_ = new_n995_ & ~new_n3354_;
  assign new_n3356_ = new_n999_ & ~new_n3355_;
  assign new_n3357_ = new_n1003_ & ~new_n3356_;
  assign new_n3358_ = new_n1007_ & ~new_n3357_;
  assign new_n3359_ = new_n1011_ & ~new_n3358_;
  assign new_n3360_ = new_n1015_ & ~new_n3359_;
  assign new_n3361_ = new_n1019_ & ~new_n3360_;
  assign new_n3362_ = new_n1023_ & ~new_n3361_;
  assign new_n3363_ = new_n1027_ & ~new_n3362_;
  assign new_n3364_ = new_n1031_ & ~new_n3363_;
  assign new_n3365_ = new_n1035_ & ~new_n3364_;
  assign new_n3366_ = new_n1039_ & ~new_n3365_;
  assign new_n3367_ = new_n1043_ & ~new_n3366_;
  assign new_n3368_ = new_n1047_ & ~new_n3367_;
  assign new_n3369_ = new_n1051_ & ~new_n3368_;
  assign new_n3370_ = new_n1055_ & ~new_n3369_;
  assign new_n3371_ = new_n1059_ & ~new_n3370_;
  assign new_n3372_ = new_n1574_ & ~new_n3371_;
  assign new_n3373_ = new_n1576_ & ~new_n3372_;
  assign new_n3374_ = new_n1837_ & ~new_n3373_;
  assign new_n3375_ = new_n1068_ & ~new_n3374_;
  assign new_n3376_ = new_n1072_ & ~new_n3375_;
  assign new_n3377_ = new_n1076_ & ~new_n3376_;
  assign new_n3378_ = new_n1080_ & ~new_n3377_;
  assign new_n3379_ = new_n1084_ & ~new_n3378_;
  assign new_n3380_ = new_n1088_ & ~new_n3379_;
  assign new_n3381_ = new_n1092_ & ~new_n3380_;
  assign new_n3382_ = new_n1096_ & ~new_n3381_;
  assign new_n3383_ = new_n1100_ & ~new_n3382_;
  assign new_n3384_ = new_n1104_ & ~new_n3383_;
  assign new_n3385_ = new_n1108_ & ~new_n3384_;
  assign new_n3386_ = new_n1112_ & ~new_n3385_;
  assign new_n3387_ = new_n1116_ & ~new_n3386_;
  assign new_n3388_ = \req[25]  & ~new_n1118_;
  assign \grant[25]  = ~new_n3387_ & new_n3388_;
  assign new_n3390_ = ~new_n455_ & new_n1127_;
  assign new_n3391_ = new_n1132_ & ~new_n3390_;
  assign new_n3392_ = new_n1136_ & ~new_n3391_;
  assign new_n3393_ = new_n1140_ & ~new_n3392_;
  assign new_n3394_ = new_n1144_ & ~new_n3393_;
  assign new_n3395_ = new_n1148_ & ~new_n3394_;
  assign new_n3396_ = new_n1152_ & ~new_n3395_;
  assign new_n3397_ = new_n1156_ & ~new_n3396_;
  assign new_n3398_ = new_n1160_ & ~new_n3397_;
  assign new_n3399_ = new_n1164_ & ~new_n3398_;
  assign new_n3400_ = new_n1168_ & ~new_n3399_;
  assign new_n3401_ = new_n1172_ & ~new_n3400_;
  assign new_n3402_ = new_n1176_ & ~new_n3401_;
  assign new_n3403_ = new_n1180_ & ~new_n3402_;
  assign new_n3404_ = new_n1184_ & ~new_n3403_;
  assign new_n3405_ = new_n1188_ & ~new_n3404_;
  assign new_n3406_ = new_n1192_ & ~new_n3405_;
  assign new_n3407_ = new_n1196_ & ~new_n3406_;
  assign new_n3408_ = new_n1200_ & ~new_n3407_;
  assign new_n3409_ = new_n1204_ & ~new_n3408_;
  assign new_n3410_ = new_n1208_ & ~new_n3409_;
  assign new_n3411_ = new_n1212_ & ~new_n3410_;
  assign new_n3412_ = new_n1216_ & ~new_n3411_;
  assign new_n3413_ = new_n1220_ & ~new_n3412_;
  assign new_n3414_ = new_n1224_ & ~new_n3413_;
  assign new_n3415_ = new_n1228_ & ~new_n3414_;
  assign new_n3416_ = new_n1232_ & ~new_n3415_;
  assign new_n3417_ = new_n1236_ & ~new_n3416_;
  assign new_n3418_ = new_n1240_ & ~new_n3417_;
  assign new_n3419_ = new_n1244_ & ~new_n3418_;
  assign new_n3420_ = new_n1248_ & ~new_n3419_;
  assign new_n3421_ = new_n1252_ & ~new_n3420_;
  assign new_n3422_ = new_n1256_ & ~new_n3421_;
  assign new_n3423_ = new_n1260_ & ~new_n3422_;
  assign new_n3424_ = new_n1264_ & ~new_n3423_;
  assign new_n3425_ = new_n1268_ & ~new_n3424_;
  assign new_n3426_ = new_n1272_ & ~new_n3425_;
  assign new_n3427_ = new_n1276_ & ~new_n3426_;
  assign new_n3428_ = new_n1280_ & ~new_n3427_;
  assign new_n3429_ = new_n1284_ & ~new_n3428_;
  assign new_n3430_ = new_n1288_ & ~new_n3429_;
  assign new_n3431_ = new_n1292_ & ~new_n3430_;
  assign new_n3432_ = new_n1296_ & ~new_n3431_;
  assign new_n3433_ = new_n1300_ & ~new_n3432_;
  assign new_n3434_ = new_n1304_ & ~new_n3433_;
  assign new_n3435_ = new_n1308_ & ~new_n3434_;
  assign new_n3436_ = new_n1312_ & ~new_n3435_;
  assign new_n3437_ = new_n1316_ & ~new_n3436_;
  assign new_n3438_ = new_n1320_ & ~new_n3437_;
  assign new_n3439_ = new_n1324_ & ~new_n3438_;
  assign new_n3440_ = new_n1328_ & ~new_n3439_;
  assign new_n3441_ = new_n1332_ & ~new_n3440_;
  assign new_n3442_ = new_n1336_ & ~new_n3441_;
  assign new_n3443_ = new_n1340_ & ~new_n3442_;
  assign new_n3444_ = new_n1344_ & ~new_n3443_;
  assign new_n3445_ = new_n1348_ & ~new_n3444_;
  assign new_n3446_ = new_n1352_ & ~new_n3445_;
  assign new_n3447_ = new_n1356_ & ~new_n3446_;
  assign new_n3448_ = new_n1360_ & ~new_n3447_;
  assign new_n3449_ = new_n1364_ & ~new_n3448_;
  assign new_n3450_ = new_n1368_ & ~new_n3449_;
  assign new_n3451_ = new_n1372_ & ~new_n3450_;
  assign new_n3452_ = new_n1376_ & ~new_n3451_;
  assign new_n3453_ = new_n1380_ & ~new_n3452_;
  assign new_n3454_ = new_n1384_ & ~new_n3453_;
  assign new_n3455_ = new_n1388_ & ~new_n3454_;
  assign new_n3456_ = new_n1392_ & ~new_n3455_;
  assign new_n3457_ = new_n1396_ & ~new_n3456_;
  assign new_n3458_ = new_n1663_ & ~new_n3457_;
  assign new_n3459_ = new_n392_ & ~new_n3458_;
  assign new_n3460_ = new_n396_ & ~new_n3459_;
  assign new_n3461_ = new_n400_ & ~new_n3460_;
  assign new_n3462_ = new_n404_ & ~new_n3461_;
  assign new_n3463_ = new_n408_ & ~new_n3462_;
  assign new_n3464_ = new_n412_ & ~new_n3463_;
  assign new_n3465_ = new_n416_ & ~new_n3464_;
  assign new_n3466_ = new_n420_ & ~new_n3465_;
  assign new_n3467_ = new_n424_ & ~new_n3466_;
  assign new_n3468_ = new_n428_ & ~new_n3467_;
  assign new_n3469_ = new_n432_ & ~new_n3468_;
  assign new_n3470_ = new_n436_ & ~new_n3469_;
  assign new_n3471_ = new_n440_ & ~new_n3470_;
  assign new_n3472_ = new_n444_ & ~new_n3471_;
  assign new_n3473_ = new_n448_ & ~new_n3472_;
  assign new_n3474_ = \req[26]  & ~new_n450_;
  assign \grant[26]  = ~new_n3473_ & new_n3474_;
  assign new_n3476_ = new_n459_ & ~new_n794_;
  assign new_n3477_ = new_n464_ & ~new_n3476_;
  assign new_n3478_ = new_n468_ & ~new_n3477_;
  assign new_n3479_ = new_n472_ & ~new_n3478_;
  assign new_n3480_ = new_n476_ & ~new_n3479_;
  assign new_n3481_ = new_n480_ & ~new_n3480_;
  assign new_n3482_ = new_n484_ & ~new_n3481_;
  assign new_n3483_ = new_n488_ & ~new_n3482_;
  assign new_n3484_ = new_n492_ & ~new_n3483_;
  assign new_n3485_ = new_n496_ & ~new_n3484_;
  assign new_n3486_ = new_n500_ & ~new_n3485_;
  assign new_n3487_ = new_n504_ & ~new_n3486_;
  assign new_n3488_ = new_n508_ & ~new_n3487_;
  assign new_n3489_ = new_n512_ & ~new_n3488_;
  assign new_n3490_ = new_n516_ & ~new_n3489_;
  assign new_n3491_ = new_n520_ & ~new_n3490_;
  assign new_n3492_ = new_n524_ & ~new_n3491_;
  assign new_n3493_ = new_n528_ & ~new_n3492_;
  assign new_n3494_ = new_n532_ & ~new_n3493_;
  assign new_n3495_ = new_n536_ & ~new_n3494_;
  assign new_n3496_ = new_n540_ & ~new_n3495_;
  assign new_n3497_ = new_n544_ & ~new_n3496_;
  assign new_n3498_ = new_n548_ & ~new_n3497_;
  assign new_n3499_ = new_n552_ & ~new_n3498_;
  assign new_n3500_ = new_n556_ & ~new_n3499_;
  assign new_n3501_ = new_n560_ & ~new_n3500_;
  assign new_n3502_ = new_n564_ & ~new_n3501_;
  assign new_n3503_ = new_n568_ & ~new_n3502_;
  assign new_n3504_ = new_n572_ & ~new_n3503_;
  assign new_n3505_ = new_n576_ & ~new_n3504_;
  assign new_n3506_ = new_n580_ & ~new_n3505_;
  assign new_n3507_ = new_n584_ & ~new_n3506_;
  assign new_n3508_ = new_n588_ & ~new_n3507_;
  assign new_n3509_ = new_n592_ & ~new_n3508_;
  assign new_n3510_ = new_n596_ & ~new_n3509_;
  assign new_n3511_ = new_n600_ & ~new_n3510_;
  assign new_n3512_ = new_n604_ & ~new_n3511_;
  assign new_n3513_ = new_n608_ & ~new_n3512_;
  assign new_n3514_ = new_n612_ & ~new_n3513_;
  assign new_n3515_ = new_n616_ & ~new_n3514_;
  assign new_n3516_ = new_n620_ & ~new_n3515_;
  assign new_n3517_ = new_n624_ & ~new_n3516_;
  assign new_n3518_ = new_n628_ & ~new_n3517_;
  assign new_n3519_ = new_n632_ & ~new_n3518_;
  assign new_n3520_ = new_n636_ & ~new_n3519_;
  assign new_n3521_ = new_n640_ & ~new_n3520_;
  assign new_n3522_ = new_n644_ & ~new_n3521_;
  assign new_n3523_ = new_n648_ & ~new_n3522_;
  assign new_n3524_ = new_n652_ & ~new_n3523_;
  assign new_n3525_ = new_n656_ & ~new_n3524_;
  assign new_n3526_ = new_n660_ & ~new_n3525_;
  assign new_n3527_ = new_n664_ & ~new_n3526_;
  assign new_n3528_ = new_n668_ & ~new_n3527_;
  assign new_n3529_ = new_n672_ & ~new_n3528_;
  assign new_n3530_ = new_n676_ & ~new_n3529_;
  assign new_n3531_ = new_n680_ & ~new_n3530_;
  assign new_n3532_ = new_n684_ & ~new_n3531_;
  assign new_n3533_ = new_n688_ & ~new_n3532_;
  assign new_n3534_ = new_n692_ & ~new_n3533_;
  assign new_n3535_ = new_n696_ & ~new_n3534_;
  assign new_n3536_ = new_n700_ & ~new_n3535_;
  assign new_n3537_ = new_n704_ & ~new_n3536_;
  assign new_n3538_ = new_n708_ & ~new_n3537_;
  assign new_n3539_ = new_n712_ & ~new_n3538_;
  assign new_n3540_ = new_n716_ & ~new_n3539_;
  assign new_n3541_ = new_n720_ & ~new_n3540_;
  assign new_n3542_ = new_n1484_ & ~new_n3541_;
  assign new_n3543_ = new_n1486_ & ~new_n3542_;
  assign new_n3544_ = new_n1750_ & ~new_n3543_;
  assign new_n3545_ = new_n731_ & ~new_n3544_;
  assign new_n3546_ = new_n735_ & ~new_n3545_;
  assign new_n3547_ = new_n739_ & ~new_n3546_;
  assign new_n3548_ = new_n743_ & ~new_n3547_;
  assign new_n3549_ = new_n747_ & ~new_n3548_;
  assign new_n3550_ = new_n751_ & ~new_n3549_;
  assign new_n3551_ = new_n755_ & ~new_n3550_;
  assign new_n3552_ = new_n759_ & ~new_n3551_;
  assign new_n3553_ = new_n763_ & ~new_n3552_;
  assign new_n3554_ = new_n767_ & ~new_n3553_;
  assign new_n3555_ = new_n771_ & ~new_n3554_;
  assign new_n3556_ = new_n775_ & ~new_n3555_;
  assign new_n3557_ = new_n779_ & ~new_n3556_;
  assign new_n3558_ = new_n783_ & ~new_n3557_;
  assign new_n3559_ = new_n787_ & ~new_n3558_;
  assign new_n3560_ = \req[27]  & ~new_n789_;
  assign \grant[27]  = ~new_n3559_ & new_n3560_;
  assign new_n3562_ = new_n798_ & ~new_n1131_;
  assign new_n3563_ = new_n803_ & ~new_n3562_;
  assign new_n3564_ = new_n807_ & ~new_n3563_;
  assign new_n3565_ = new_n811_ & ~new_n3564_;
  assign new_n3566_ = new_n815_ & ~new_n3565_;
  assign new_n3567_ = new_n819_ & ~new_n3566_;
  assign new_n3568_ = new_n823_ & ~new_n3567_;
  assign new_n3569_ = new_n827_ & ~new_n3568_;
  assign new_n3570_ = new_n831_ & ~new_n3569_;
  assign new_n3571_ = new_n835_ & ~new_n3570_;
  assign new_n3572_ = new_n839_ & ~new_n3571_;
  assign new_n3573_ = new_n843_ & ~new_n3572_;
  assign new_n3574_ = new_n847_ & ~new_n3573_;
  assign new_n3575_ = new_n851_ & ~new_n3574_;
  assign new_n3576_ = new_n855_ & ~new_n3575_;
  assign new_n3577_ = new_n859_ & ~new_n3576_;
  assign new_n3578_ = new_n863_ & ~new_n3577_;
  assign new_n3579_ = new_n867_ & ~new_n3578_;
  assign new_n3580_ = new_n871_ & ~new_n3579_;
  assign new_n3581_ = new_n875_ & ~new_n3580_;
  assign new_n3582_ = new_n879_ & ~new_n3581_;
  assign new_n3583_ = new_n883_ & ~new_n3582_;
  assign new_n3584_ = new_n887_ & ~new_n3583_;
  assign new_n3585_ = new_n891_ & ~new_n3584_;
  assign new_n3586_ = new_n895_ & ~new_n3585_;
  assign new_n3587_ = new_n899_ & ~new_n3586_;
  assign new_n3588_ = new_n903_ & ~new_n3587_;
  assign new_n3589_ = new_n907_ & ~new_n3588_;
  assign new_n3590_ = new_n911_ & ~new_n3589_;
  assign new_n3591_ = new_n915_ & ~new_n3590_;
  assign new_n3592_ = new_n919_ & ~new_n3591_;
  assign new_n3593_ = new_n923_ & ~new_n3592_;
  assign new_n3594_ = new_n927_ & ~new_n3593_;
  assign new_n3595_ = new_n931_ & ~new_n3594_;
  assign new_n3596_ = new_n935_ & ~new_n3595_;
  assign new_n3597_ = new_n939_ & ~new_n3596_;
  assign new_n3598_ = new_n943_ & ~new_n3597_;
  assign new_n3599_ = new_n947_ & ~new_n3598_;
  assign new_n3600_ = new_n951_ & ~new_n3599_;
  assign new_n3601_ = new_n955_ & ~new_n3600_;
  assign new_n3602_ = new_n959_ & ~new_n3601_;
  assign new_n3603_ = new_n963_ & ~new_n3602_;
  assign new_n3604_ = new_n967_ & ~new_n3603_;
  assign new_n3605_ = new_n971_ & ~new_n3604_;
  assign new_n3606_ = new_n975_ & ~new_n3605_;
  assign new_n3607_ = new_n979_ & ~new_n3606_;
  assign new_n3608_ = new_n983_ & ~new_n3607_;
  assign new_n3609_ = new_n987_ & ~new_n3608_;
  assign new_n3610_ = new_n991_ & ~new_n3609_;
  assign new_n3611_ = new_n995_ & ~new_n3610_;
  assign new_n3612_ = new_n999_ & ~new_n3611_;
  assign new_n3613_ = new_n1003_ & ~new_n3612_;
  assign new_n3614_ = new_n1007_ & ~new_n3613_;
  assign new_n3615_ = new_n1011_ & ~new_n3614_;
  assign new_n3616_ = new_n1015_ & ~new_n3615_;
  assign new_n3617_ = new_n1019_ & ~new_n3616_;
  assign new_n3618_ = new_n1023_ & ~new_n3617_;
  assign new_n3619_ = new_n1027_ & ~new_n3618_;
  assign new_n3620_ = new_n1031_ & ~new_n3619_;
  assign new_n3621_ = new_n1035_ & ~new_n3620_;
  assign new_n3622_ = new_n1039_ & ~new_n3621_;
  assign new_n3623_ = new_n1043_ & ~new_n3622_;
  assign new_n3624_ = new_n1047_ & ~new_n3623_;
  assign new_n3625_ = new_n1051_ & ~new_n3624_;
  assign new_n3626_ = new_n1055_ & ~new_n3625_;
  assign new_n3627_ = new_n1059_ & ~new_n3626_;
  assign new_n3628_ = new_n1574_ & ~new_n3627_;
  assign new_n3629_ = new_n1576_ & ~new_n3628_;
  assign new_n3630_ = new_n1837_ & ~new_n3629_;
  assign new_n3631_ = new_n1068_ & ~new_n3630_;
  assign new_n3632_ = new_n1072_ & ~new_n3631_;
  assign new_n3633_ = new_n1076_ & ~new_n3632_;
  assign new_n3634_ = new_n1080_ & ~new_n3633_;
  assign new_n3635_ = new_n1084_ & ~new_n3634_;
  assign new_n3636_ = new_n1088_ & ~new_n3635_;
  assign new_n3637_ = new_n1092_ & ~new_n3636_;
  assign new_n3638_ = new_n1096_ & ~new_n3637_;
  assign new_n3639_ = new_n1100_ & ~new_n3638_;
  assign new_n3640_ = new_n1104_ & ~new_n3639_;
  assign new_n3641_ = new_n1108_ & ~new_n3640_;
  assign new_n3642_ = new_n1112_ & ~new_n3641_;
  assign new_n3643_ = new_n1116_ & ~new_n3642_;
  assign new_n3644_ = new_n1120_ & ~new_n3643_;
  assign new_n3645_ = new_n1124_ & ~new_n3644_;
  assign new_n3646_ = \req[28]  & ~new_n1126_;
  assign \grant[28]  = ~new_n3645_ & new_n3646_;
  assign new_n3648_ = ~new_n463_ & new_n1135_;
  assign new_n3649_ = new_n1140_ & ~new_n3648_;
  assign new_n3650_ = new_n1144_ & ~new_n3649_;
  assign new_n3651_ = new_n1148_ & ~new_n3650_;
  assign new_n3652_ = new_n1152_ & ~new_n3651_;
  assign new_n3653_ = new_n1156_ & ~new_n3652_;
  assign new_n3654_ = new_n1160_ & ~new_n3653_;
  assign new_n3655_ = new_n1164_ & ~new_n3654_;
  assign new_n3656_ = new_n1168_ & ~new_n3655_;
  assign new_n3657_ = new_n1172_ & ~new_n3656_;
  assign new_n3658_ = new_n1176_ & ~new_n3657_;
  assign new_n3659_ = new_n1180_ & ~new_n3658_;
  assign new_n3660_ = new_n1184_ & ~new_n3659_;
  assign new_n3661_ = new_n1188_ & ~new_n3660_;
  assign new_n3662_ = new_n1192_ & ~new_n3661_;
  assign new_n3663_ = new_n1196_ & ~new_n3662_;
  assign new_n3664_ = new_n1200_ & ~new_n3663_;
  assign new_n3665_ = new_n1204_ & ~new_n3664_;
  assign new_n3666_ = new_n1208_ & ~new_n3665_;
  assign new_n3667_ = new_n1212_ & ~new_n3666_;
  assign new_n3668_ = new_n1216_ & ~new_n3667_;
  assign new_n3669_ = new_n1220_ & ~new_n3668_;
  assign new_n3670_ = new_n1224_ & ~new_n3669_;
  assign new_n3671_ = new_n1228_ & ~new_n3670_;
  assign new_n3672_ = new_n1232_ & ~new_n3671_;
  assign new_n3673_ = new_n1236_ & ~new_n3672_;
  assign new_n3674_ = new_n1240_ & ~new_n3673_;
  assign new_n3675_ = new_n1244_ & ~new_n3674_;
  assign new_n3676_ = new_n1248_ & ~new_n3675_;
  assign new_n3677_ = new_n1252_ & ~new_n3676_;
  assign new_n3678_ = new_n1256_ & ~new_n3677_;
  assign new_n3679_ = new_n1260_ & ~new_n3678_;
  assign new_n3680_ = new_n1264_ & ~new_n3679_;
  assign new_n3681_ = new_n1268_ & ~new_n3680_;
  assign new_n3682_ = new_n1272_ & ~new_n3681_;
  assign new_n3683_ = new_n1276_ & ~new_n3682_;
  assign new_n3684_ = new_n1280_ & ~new_n3683_;
  assign new_n3685_ = new_n1284_ & ~new_n3684_;
  assign new_n3686_ = new_n1288_ & ~new_n3685_;
  assign new_n3687_ = new_n1292_ & ~new_n3686_;
  assign new_n3688_ = new_n1296_ & ~new_n3687_;
  assign new_n3689_ = new_n1300_ & ~new_n3688_;
  assign new_n3690_ = new_n1304_ & ~new_n3689_;
  assign new_n3691_ = new_n1308_ & ~new_n3690_;
  assign new_n3692_ = new_n1312_ & ~new_n3691_;
  assign new_n3693_ = new_n1316_ & ~new_n3692_;
  assign new_n3694_ = new_n1320_ & ~new_n3693_;
  assign new_n3695_ = new_n1324_ & ~new_n3694_;
  assign new_n3696_ = new_n1328_ & ~new_n3695_;
  assign new_n3697_ = new_n1332_ & ~new_n3696_;
  assign new_n3698_ = new_n1336_ & ~new_n3697_;
  assign new_n3699_ = new_n1340_ & ~new_n3698_;
  assign new_n3700_ = new_n1344_ & ~new_n3699_;
  assign new_n3701_ = new_n1348_ & ~new_n3700_;
  assign new_n3702_ = new_n1352_ & ~new_n3701_;
  assign new_n3703_ = new_n1356_ & ~new_n3702_;
  assign new_n3704_ = new_n1360_ & ~new_n3703_;
  assign new_n3705_ = new_n1364_ & ~new_n3704_;
  assign new_n3706_ = new_n1368_ & ~new_n3705_;
  assign new_n3707_ = new_n1372_ & ~new_n3706_;
  assign new_n3708_ = new_n1376_ & ~new_n3707_;
  assign new_n3709_ = new_n1380_ & ~new_n3708_;
  assign new_n3710_ = new_n1384_ & ~new_n3709_;
  assign new_n3711_ = new_n1388_ & ~new_n3710_;
  assign new_n3712_ = new_n1392_ & ~new_n3711_;
  assign new_n3713_ = new_n1396_ & ~new_n3712_;
  assign new_n3714_ = new_n1663_ & ~new_n3713_;
  assign new_n3715_ = new_n392_ & ~new_n3714_;
  assign new_n3716_ = new_n396_ & ~new_n3715_;
  assign new_n3717_ = new_n400_ & ~new_n3716_;
  assign new_n3718_ = new_n404_ & ~new_n3717_;
  assign new_n3719_ = new_n408_ & ~new_n3718_;
  assign new_n3720_ = new_n412_ & ~new_n3719_;
  assign new_n3721_ = new_n416_ & ~new_n3720_;
  assign new_n3722_ = new_n420_ & ~new_n3721_;
  assign new_n3723_ = new_n424_ & ~new_n3722_;
  assign new_n3724_ = new_n428_ & ~new_n3723_;
  assign new_n3725_ = new_n432_ & ~new_n3724_;
  assign new_n3726_ = new_n436_ & ~new_n3725_;
  assign new_n3727_ = new_n440_ & ~new_n3726_;
  assign new_n3728_ = new_n444_ & ~new_n3727_;
  assign new_n3729_ = new_n448_ & ~new_n3728_;
  assign new_n3730_ = new_n452_ & ~new_n3729_;
  assign new_n3731_ = new_n456_ & ~new_n3730_;
  assign new_n3732_ = \req[29]  & ~new_n458_;
  assign \grant[29]  = ~new_n3731_ & new_n3732_;
  assign new_n3734_ = new_n467_ & ~new_n802_;
  assign new_n3735_ = new_n472_ & ~new_n3734_;
  assign new_n3736_ = new_n476_ & ~new_n3735_;
  assign new_n3737_ = new_n480_ & ~new_n3736_;
  assign new_n3738_ = new_n484_ & ~new_n3737_;
  assign new_n3739_ = new_n488_ & ~new_n3738_;
  assign new_n3740_ = new_n492_ & ~new_n3739_;
  assign new_n3741_ = new_n496_ & ~new_n3740_;
  assign new_n3742_ = new_n500_ & ~new_n3741_;
  assign new_n3743_ = new_n504_ & ~new_n3742_;
  assign new_n3744_ = new_n508_ & ~new_n3743_;
  assign new_n3745_ = new_n512_ & ~new_n3744_;
  assign new_n3746_ = new_n516_ & ~new_n3745_;
  assign new_n3747_ = new_n520_ & ~new_n3746_;
  assign new_n3748_ = new_n524_ & ~new_n3747_;
  assign new_n3749_ = new_n528_ & ~new_n3748_;
  assign new_n3750_ = new_n532_ & ~new_n3749_;
  assign new_n3751_ = new_n536_ & ~new_n3750_;
  assign new_n3752_ = new_n540_ & ~new_n3751_;
  assign new_n3753_ = new_n544_ & ~new_n3752_;
  assign new_n3754_ = new_n548_ & ~new_n3753_;
  assign new_n3755_ = new_n552_ & ~new_n3754_;
  assign new_n3756_ = new_n556_ & ~new_n3755_;
  assign new_n3757_ = new_n560_ & ~new_n3756_;
  assign new_n3758_ = new_n564_ & ~new_n3757_;
  assign new_n3759_ = new_n568_ & ~new_n3758_;
  assign new_n3760_ = new_n572_ & ~new_n3759_;
  assign new_n3761_ = new_n576_ & ~new_n3760_;
  assign new_n3762_ = new_n580_ & ~new_n3761_;
  assign new_n3763_ = new_n584_ & ~new_n3762_;
  assign new_n3764_ = new_n588_ & ~new_n3763_;
  assign new_n3765_ = new_n592_ & ~new_n3764_;
  assign new_n3766_ = new_n596_ & ~new_n3765_;
  assign new_n3767_ = new_n600_ & ~new_n3766_;
  assign new_n3768_ = new_n604_ & ~new_n3767_;
  assign new_n3769_ = new_n608_ & ~new_n3768_;
  assign new_n3770_ = new_n612_ & ~new_n3769_;
  assign new_n3771_ = new_n616_ & ~new_n3770_;
  assign new_n3772_ = new_n620_ & ~new_n3771_;
  assign new_n3773_ = new_n624_ & ~new_n3772_;
  assign new_n3774_ = new_n628_ & ~new_n3773_;
  assign new_n3775_ = new_n632_ & ~new_n3774_;
  assign new_n3776_ = new_n636_ & ~new_n3775_;
  assign new_n3777_ = new_n640_ & ~new_n3776_;
  assign new_n3778_ = new_n644_ & ~new_n3777_;
  assign new_n3779_ = new_n648_ & ~new_n3778_;
  assign new_n3780_ = new_n652_ & ~new_n3779_;
  assign new_n3781_ = new_n656_ & ~new_n3780_;
  assign new_n3782_ = new_n660_ & ~new_n3781_;
  assign new_n3783_ = new_n664_ & ~new_n3782_;
  assign new_n3784_ = new_n668_ & ~new_n3783_;
  assign new_n3785_ = new_n672_ & ~new_n3784_;
  assign new_n3786_ = new_n676_ & ~new_n3785_;
  assign new_n3787_ = new_n680_ & ~new_n3786_;
  assign new_n3788_ = new_n684_ & ~new_n3787_;
  assign new_n3789_ = new_n688_ & ~new_n3788_;
  assign new_n3790_ = new_n692_ & ~new_n3789_;
  assign new_n3791_ = new_n696_ & ~new_n3790_;
  assign new_n3792_ = new_n700_ & ~new_n3791_;
  assign new_n3793_ = new_n704_ & ~new_n3792_;
  assign new_n3794_ = new_n708_ & ~new_n3793_;
  assign new_n3795_ = new_n712_ & ~new_n3794_;
  assign new_n3796_ = new_n716_ & ~new_n3795_;
  assign new_n3797_ = new_n720_ & ~new_n3796_;
  assign new_n3798_ = new_n1484_ & ~new_n3797_;
  assign new_n3799_ = new_n1486_ & ~new_n3798_;
  assign new_n3800_ = new_n1750_ & ~new_n3799_;
  assign new_n3801_ = new_n731_ & ~new_n3800_;
  assign new_n3802_ = new_n735_ & ~new_n3801_;
  assign new_n3803_ = new_n739_ & ~new_n3802_;
  assign new_n3804_ = new_n743_ & ~new_n3803_;
  assign new_n3805_ = new_n747_ & ~new_n3804_;
  assign new_n3806_ = new_n751_ & ~new_n3805_;
  assign new_n3807_ = new_n755_ & ~new_n3806_;
  assign new_n3808_ = new_n759_ & ~new_n3807_;
  assign new_n3809_ = new_n763_ & ~new_n3808_;
  assign new_n3810_ = new_n767_ & ~new_n3809_;
  assign new_n3811_ = new_n771_ & ~new_n3810_;
  assign new_n3812_ = new_n775_ & ~new_n3811_;
  assign new_n3813_ = new_n779_ & ~new_n3812_;
  assign new_n3814_ = new_n783_ & ~new_n3813_;
  assign new_n3815_ = new_n787_ & ~new_n3814_;
  assign new_n3816_ = new_n791_ & ~new_n3815_;
  assign new_n3817_ = new_n795_ & ~new_n3816_;
  assign new_n3818_ = \req[30]  & ~new_n797_;
  assign \grant[30]  = ~new_n3817_ & new_n3818_;
  assign new_n3820_ = new_n806_ & ~new_n1139_;
  assign new_n3821_ = new_n811_ & ~new_n3820_;
  assign new_n3822_ = new_n815_ & ~new_n3821_;
  assign new_n3823_ = new_n819_ & ~new_n3822_;
  assign new_n3824_ = new_n823_ & ~new_n3823_;
  assign new_n3825_ = new_n827_ & ~new_n3824_;
  assign new_n3826_ = new_n831_ & ~new_n3825_;
  assign new_n3827_ = new_n835_ & ~new_n3826_;
  assign new_n3828_ = new_n839_ & ~new_n3827_;
  assign new_n3829_ = new_n843_ & ~new_n3828_;
  assign new_n3830_ = new_n847_ & ~new_n3829_;
  assign new_n3831_ = new_n851_ & ~new_n3830_;
  assign new_n3832_ = new_n855_ & ~new_n3831_;
  assign new_n3833_ = new_n859_ & ~new_n3832_;
  assign new_n3834_ = new_n863_ & ~new_n3833_;
  assign new_n3835_ = new_n867_ & ~new_n3834_;
  assign new_n3836_ = new_n871_ & ~new_n3835_;
  assign new_n3837_ = new_n875_ & ~new_n3836_;
  assign new_n3838_ = new_n879_ & ~new_n3837_;
  assign new_n3839_ = new_n883_ & ~new_n3838_;
  assign new_n3840_ = new_n887_ & ~new_n3839_;
  assign new_n3841_ = new_n891_ & ~new_n3840_;
  assign new_n3842_ = new_n895_ & ~new_n3841_;
  assign new_n3843_ = new_n899_ & ~new_n3842_;
  assign new_n3844_ = new_n903_ & ~new_n3843_;
  assign new_n3845_ = new_n907_ & ~new_n3844_;
  assign new_n3846_ = new_n911_ & ~new_n3845_;
  assign new_n3847_ = new_n915_ & ~new_n3846_;
  assign new_n3848_ = new_n919_ & ~new_n3847_;
  assign new_n3849_ = new_n923_ & ~new_n3848_;
  assign new_n3850_ = new_n927_ & ~new_n3849_;
  assign new_n3851_ = new_n931_ & ~new_n3850_;
  assign new_n3852_ = new_n935_ & ~new_n3851_;
  assign new_n3853_ = new_n939_ & ~new_n3852_;
  assign new_n3854_ = new_n943_ & ~new_n3853_;
  assign new_n3855_ = new_n947_ & ~new_n3854_;
  assign new_n3856_ = new_n951_ & ~new_n3855_;
  assign new_n3857_ = new_n955_ & ~new_n3856_;
  assign new_n3858_ = new_n959_ & ~new_n3857_;
  assign new_n3859_ = new_n963_ & ~new_n3858_;
  assign new_n3860_ = new_n967_ & ~new_n3859_;
  assign new_n3861_ = new_n971_ & ~new_n3860_;
  assign new_n3862_ = new_n975_ & ~new_n3861_;
  assign new_n3863_ = new_n979_ & ~new_n3862_;
  assign new_n3864_ = new_n983_ & ~new_n3863_;
  assign new_n3865_ = new_n987_ & ~new_n3864_;
  assign new_n3866_ = new_n991_ & ~new_n3865_;
  assign new_n3867_ = new_n995_ & ~new_n3866_;
  assign new_n3868_ = new_n999_ & ~new_n3867_;
  assign new_n3869_ = new_n1003_ & ~new_n3868_;
  assign new_n3870_ = new_n1007_ & ~new_n3869_;
  assign new_n3871_ = new_n1011_ & ~new_n3870_;
  assign new_n3872_ = new_n1015_ & ~new_n3871_;
  assign new_n3873_ = new_n1019_ & ~new_n3872_;
  assign new_n3874_ = new_n1023_ & ~new_n3873_;
  assign new_n3875_ = new_n1027_ & ~new_n3874_;
  assign new_n3876_ = new_n1031_ & ~new_n3875_;
  assign new_n3877_ = new_n1035_ & ~new_n3876_;
  assign new_n3878_ = new_n1039_ & ~new_n3877_;
  assign new_n3879_ = new_n1043_ & ~new_n3878_;
  assign new_n3880_ = new_n1047_ & ~new_n3879_;
  assign new_n3881_ = new_n1051_ & ~new_n3880_;
  assign new_n3882_ = new_n1055_ & ~new_n3881_;
  assign new_n3883_ = new_n1059_ & ~new_n3882_;
  assign new_n3884_ = new_n1574_ & ~new_n3883_;
  assign new_n3885_ = new_n1576_ & ~new_n3884_;
  assign new_n3886_ = new_n1837_ & ~new_n3885_;
  assign new_n3887_ = new_n1068_ & ~new_n3886_;
  assign new_n3888_ = new_n1072_ & ~new_n3887_;
  assign new_n3889_ = new_n1076_ & ~new_n3888_;
  assign new_n3890_ = new_n1080_ & ~new_n3889_;
  assign new_n3891_ = new_n1084_ & ~new_n3890_;
  assign new_n3892_ = new_n1088_ & ~new_n3891_;
  assign new_n3893_ = new_n1092_ & ~new_n3892_;
  assign new_n3894_ = new_n1096_ & ~new_n3893_;
  assign new_n3895_ = new_n1100_ & ~new_n3894_;
  assign new_n3896_ = new_n1104_ & ~new_n3895_;
  assign new_n3897_ = new_n1108_ & ~new_n3896_;
  assign new_n3898_ = new_n1112_ & ~new_n3897_;
  assign new_n3899_ = new_n1116_ & ~new_n3898_;
  assign new_n3900_ = new_n1120_ & ~new_n3899_;
  assign new_n3901_ = new_n1124_ & ~new_n3900_;
  assign new_n3902_ = new_n1128_ & ~new_n3901_;
  assign new_n3903_ = new_n1132_ & ~new_n3902_;
  assign new_n3904_ = \req[31]  & ~new_n1134_;
  assign \grant[31]  = ~new_n3903_ & new_n3904_;
  assign new_n3906_ = ~new_n471_ & new_n1143_;
  assign new_n3907_ = new_n1148_ & ~new_n3906_;
  assign new_n3908_ = new_n1152_ & ~new_n3907_;
  assign new_n3909_ = new_n1156_ & ~new_n3908_;
  assign new_n3910_ = new_n1160_ & ~new_n3909_;
  assign new_n3911_ = new_n1164_ & ~new_n3910_;
  assign new_n3912_ = new_n1168_ & ~new_n3911_;
  assign new_n3913_ = new_n1172_ & ~new_n3912_;
  assign new_n3914_ = new_n1176_ & ~new_n3913_;
  assign new_n3915_ = new_n1180_ & ~new_n3914_;
  assign new_n3916_ = new_n1184_ & ~new_n3915_;
  assign new_n3917_ = new_n1188_ & ~new_n3916_;
  assign new_n3918_ = new_n1192_ & ~new_n3917_;
  assign new_n3919_ = new_n1196_ & ~new_n3918_;
  assign new_n3920_ = new_n1200_ & ~new_n3919_;
  assign new_n3921_ = new_n1204_ & ~new_n3920_;
  assign new_n3922_ = new_n1208_ & ~new_n3921_;
  assign new_n3923_ = new_n1212_ & ~new_n3922_;
  assign new_n3924_ = new_n1216_ & ~new_n3923_;
  assign new_n3925_ = new_n1220_ & ~new_n3924_;
  assign new_n3926_ = new_n1224_ & ~new_n3925_;
  assign new_n3927_ = new_n1228_ & ~new_n3926_;
  assign new_n3928_ = new_n1232_ & ~new_n3927_;
  assign new_n3929_ = new_n1236_ & ~new_n3928_;
  assign new_n3930_ = new_n1240_ & ~new_n3929_;
  assign new_n3931_ = new_n1244_ & ~new_n3930_;
  assign new_n3932_ = new_n1248_ & ~new_n3931_;
  assign new_n3933_ = new_n1252_ & ~new_n3932_;
  assign new_n3934_ = new_n1256_ & ~new_n3933_;
  assign new_n3935_ = new_n1260_ & ~new_n3934_;
  assign new_n3936_ = new_n1264_ & ~new_n3935_;
  assign new_n3937_ = new_n1268_ & ~new_n3936_;
  assign new_n3938_ = new_n1272_ & ~new_n3937_;
  assign new_n3939_ = new_n1276_ & ~new_n3938_;
  assign new_n3940_ = new_n1280_ & ~new_n3939_;
  assign new_n3941_ = new_n1284_ & ~new_n3940_;
  assign new_n3942_ = new_n1288_ & ~new_n3941_;
  assign new_n3943_ = new_n1292_ & ~new_n3942_;
  assign new_n3944_ = new_n1296_ & ~new_n3943_;
  assign new_n3945_ = new_n1300_ & ~new_n3944_;
  assign new_n3946_ = new_n1304_ & ~new_n3945_;
  assign new_n3947_ = new_n1308_ & ~new_n3946_;
  assign new_n3948_ = new_n1312_ & ~new_n3947_;
  assign new_n3949_ = new_n1316_ & ~new_n3948_;
  assign new_n3950_ = new_n1320_ & ~new_n3949_;
  assign new_n3951_ = new_n1324_ & ~new_n3950_;
  assign new_n3952_ = new_n1328_ & ~new_n3951_;
  assign new_n3953_ = new_n1332_ & ~new_n3952_;
  assign new_n3954_ = new_n1336_ & ~new_n3953_;
  assign new_n3955_ = new_n1340_ & ~new_n3954_;
  assign new_n3956_ = new_n1344_ & ~new_n3955_;
  assign new_n3957_ = new_n1348_ & ~new_n3956_;
  assign new_n3958_ = new_n1352_ & ~new_n3957_;
  assign new_n3959_ = new_n1356_ & ~new_n3958_;
  assign new_n3960_ = new_n1360_ & ~new_n3959_;
  assign new_n3961_ = new_n1364_ & ~new_n3960_;
  assign new_n3962_ = new_n1368_ & ~new_n3961_;
  assign new_n3963_ = new_n1372_ & ~new_n3962_;
  assign new_n3964_ = new_n1376_ & ~new_n3963_;
  assign new_n3965_ = new_n1380_ & ~new_n3964_;
  assign new_n3966_ = new_n1384_ & ~new_n3965_;
  assign new_n3967_ = new_n1388_ & ~new_n3966_;
  assign new_n3968_ = new_n1392_ & ~new_n3967_;
  assign new_n3969_ = new_n1396_ & ~new_n3968_;
  assign new_n3970_ = new_n1663_ & ~new_n3969_;
  assign new_n3971_ = new_n392_ & ~new_n3970_;
  assign new_n3972_ = new_n396_ & ~new_n3971_;
  assign new_n3973_ = new_n400_ & ~new_n3972_;
  assign new_n3974_ = new_n404_ & ~new_n3973_;
  assign new_n3975_ = new_n408_ & ~new_n3974_;
  assign new_n3976_ = new_n412_ & ~new_n3975_;
  assign new_n3977_ = new_n416_ & ~new_n3976_;
  assign new_n3978_ = new_n420_ & ~new_n3977_;
  assign new_n3979_ = new_n424_ & ~new_n3978_;
  assign new_n3980_ = new_n428_ & ~new_n3979_;
  assign new_n3981_ = new_n432_ & ~new_n3980_;
  assign new_n3982_ = new_n436_ & ~new_n3981_;
  assign new_n3983_ = new_n440_ & ~new_n3982_;
  assign new_n3984_ = new_n444_ & ~new_n3983_;
  assign new_n3985_ = new_n448_ & ~new_n3984_;
  assign new_n3986_ = new_n452_ & ~new_n3985_;
  assign new_n3987_ = new_n456_ & ~new_n3986_;
  assign new_n3988_ = new_n460_ & ~new_n3987_;
  assign new_n3989_ = new_n464_ & ~new_n3988_;
  assign new_n3990_ = \req[32]  & ~new_n466_;
  assign \grant[32]  = ~new_n3989_ & new_n3990_;
  assign new_n3992_ = new_n475_ & ~new_n810_;
  assign new_n3993_ = new_n480_ & ~new_n3992_;
  assign new_n3994_ = new_n484_ & ~new_n3993_;
  assign new_n3995_ = new_n488_ & ~new_n3994_;
  assign new_n3996_ = new_n492_ & ~new_n3995_;
  assign new_n3997_ = new_n496_ & ~new_n3996_;
  assign new_n3998_ = new_n500_ & ~new_n3997_;
  assign new_n3999_ = new_n504_ & ~new_n3998_;
  assign new_n4000_ = new_n508_ & ~new_n3999_;
  assign new_n4001_ = new_n512_ & ~new_n4000_;
  assign new_n4002_ = new_n516_ & ~new_n4001_;
  assign new_n4003_ = new_n520_ & ~new_n4002_;
  assign new_n4004_ = new_n524_ & ~new_n4003_;
  assign new_n4005_ = new_n528_ & ~new_n4004_;
  assign new_n4006_ = new_n532_ & ~new_n4005_;
  assign new_n4007_ = new_n536_ & ~new_n4006_;
  assign new_n4008_ = new_n540_ & ~new_n4007_;
  assign new_n4009_ = new_n544_ & ~new_n4008_;
  assign new_n4010_ = new_n548_ & ~new_n4009_;
  assign new_n4011_ = new_n552_ & ~new_n4010_;
  assign new_n4012_ = new_n556_ & ~new_n4011_;
  assign new_n4013_ = new_n560_ & ~new_n4012_;
  assign new_n4014_ = new_n564_ & ~new_n4013_;
  assign new_n4015_ = new_n568_ & ~new_n4014_;
  assign new_n4016_ = new_n572_ & ~new_n4015_;
  assign new_n4017_ = new_n576_ & ~new_n4016_;
  assign new_n4018_ = new_n580_ & ~new_n4017_;
  assign new_n4019_ = new_n584_ & ~new_n4018_;
  assign new_n4020_ = new_n588_ & ~new_n4019_;
  assign new_n4021_ = new_n592_ & ~new_n4020_;
  assign new_n4022_ = new_n596_ & ~new_n4021_;
  assign new_n4023_ = new_n600_ & ~new_n4022_;
  assign new_n4024_ = new_n604_ & ~new_n4023_;
  assign new_n4025_ = new_n608_ & ~new_n4024_;
  assign new_n4026_ = new_n612_ & ~new_n4025_;
  assign new_n4027_ = new_n616_ & ~new_n4026_;
  assign new_n4028_ = new_n620_ & ~new_n4027_;
  assign new_n4029_ = new_n624_ & ~new_n4028_;
  assign new_n4030_ = new_n628_ & ~new_n4029_;
  assign new_n4031_ = new_n632_ & ~new_n4030_;
  assign new_n4032_ = new_n636_ & ~new_n4031_;
  assign new_n4033_ = new_n640_ & ~new_n4032_;
  assign new_n4034_ = new_n644_ & ~new_n4033_;
  assign new_n4035_ = new_n648_ & ~new_n4034_;
  assign new_n4036_ = new_n652_ & ~new_n4035_;
  assign new_n4037_ = new_n656_ & ~new_n4036_;
  assign new_n4038_ = new_n660_ & ~new_n4037_;
  assign new_n4039_ = new_n664_ & ~new_n4038_;
  assign new_n4040_ = new_n668_ & ~new_n4039_;
  assign new_n4041_ = new_n672_ & ~new_n4040_;
  assign new_n4042_ = new_n676_ & ~new_n4041_;
  assign new_n4043_ = new_n680_ & ~new_n4042_;
  assign new_n4044_ = new_n684_ & ~new_n4043_;
  assign new_n4045_ = new_n688_ & ~new_n4044_;
  assign new_n4046_ = new_n692_ & ~new_n4045_;
  assign new_n4047_ = new_n696_ & ~new_n4046_;
  assign new_n4048_ = new_n700_ & ~new_n4047_;
  assign new_n4049_ = new_n704_ & ~new_n4048_;
  assign new_n4050_ = new_n708_ & ~new_n4049_;
  assign new_n4051_ = new_n712_ & ~new_n4050_;
  assign new_n4052_ = new_n716_ & ~new_n4051_;
  assign new_n4053_ = new_n720_ & ~new_n4052_;
  assign new_n4054_ = new_n1484_ & ~new_n4053_;
  assign new_n4055_ = new_n1486_ & ~new_n4054_;
  assign new_n4056_ = new_n1750_ & ~new_n4055_;
  assign new_n4057_ = new_n731_ & ~new_n4056_;
  assign new_n4058_ = new_n735_ & ~new_n4057_;
  assign new_n4059_ = new_n739_ & ~new_n4058_;
  assign new_n4060_ = new_n743_ & ~new_n4059_;
  assign new_n4061_ = new_n747_ & ~new_n4060_;
  assign new_n4062_ = new_n751_ & ~new_n4061_;
  assign new_n4063_ = new_n755_ & ~new_n4062_;
  assign new_n4064_ = new_n759_ & ~new_n4063_;
  assign new_n4065_ = new_n763_ & ~new_n4064_;
  assign new_n4066_ = new_n767_ & ~new_n4065_;
  assign new_n4067_ = new_n771_ & ~new_n4066_;
  assign new_n4068_ = new_n775_ & ~new_n4067_;
  assign new_n4069_ = new_n779_ & ~new_n4068_;
  assign new_n4070_ = new_n783_ & ~new_n4069_;
  assign new_n4071_ = new_n787_ & ~new_n4070_;
  assign new_n4072_ = new_n791_ & ~new_n4071_;
  assign new_n4073_ = new_n795_ & ~new_n4072_;
  assign new_n4074_ = new_n799_ & ~new_n4073_;
  assign new_n4075_ = new_n803_ & ~new_n4074_;
  assign new_n4076_ = \req[33]  & ~new_n805_;
  assign \grant[33]  = ~new_n4075_ & new_n4076_;
  assign new_n4078_ = new_n814_ & ~new_n1147_;
  assign new_n4079_ = new_n819_ & ~new_n4078_;
  assign new_n4080_ = new_n823_ & ~new_n4079_;
  assign new_n4081_ = new_n827_ & ~new_n4080_;
  assign new_n4082_ = new_n831_ & ~new_n4081_;
  assign new_n4083_ = new_n835_ & ~new_n4082_;
  assign new_n4084_ = new_n839_ & ~new_n4083_;
  assign new_n4085_ = new_n843_ & ~new_n4084_;
  assign new_n4086_ = new_n847_ & ~new_n4085_;
  assign new_n4087_ = new_n851_ & ~new_n4086_;
  assign new_n4088_ = new_n855_ & ~new_n4087_;
  assign new_n4089_ = new_n859_ & ~new_n4088_;
  assign new_n4090_ = new_n863_ & ~new_n4089_;
  assign new_n4091_ = new_n867_ & ~new_n4090_;
  assign new_n4092_ = new_n871_ & ~new_n4091_;
  assign new_n4093_ = new_n875_ & ~new_n4092_;
  assign new_n4094_ = new_n879_ & ~new_n4093_;
  assign new_n4095_ = new_n883_ & ~new_n4094_;
  assign new_n4096_ = new_n887_ & ~new_n4095_;
  assign new_n4097_ = new_n891_ & ~new_n4096_;
  assign new_n4098_ = new_n895_ & ~new_n4097_;
  assign new_n4099_ = new_n899_ & ~new_n4098_;
  assign new_n4100_ = new_n903_ & ~new_n4099_;
  assign new_n4101_ = new_n907_ & ~new_n4100_;
  assign new_n4102_ = new_n911_ & ~new_n4101_;
  assign new_n4103_ = new_n915_ & ~new_n4102_;
  assign new_n4104_ = new_n919_ & ~new_n4103_;
  assign new_n4105_ = new_n923_ & ~new_n4104_;
  assign new_n4106_ = new_n927_ & ~new_n4105_;
  assign new_n4107_ = new_n931_ & ~new_n4106_;
  assign new_n4108_ = new_n935_ & ~new_n4107_;
  assign new_n4109_ = new_n939_ & ~new_n4108_;
  assign new_n4110_ = new_n943_ & ~new_n4109_;
  assign new_n4111_ = new_n947_ & ~new_n4110_;
  assign new_n4112_ = new_n951_ & ~new_n4111_;
  assign new_n4113_ = new_n955_ & ~new_n4112_;
  assign new_n4114_ = new_n959_ & ~new_n4113_;
  assign new_n4115_ = new_n963_ & ~new_n4114_;
  assign new_n4116_ = new_n967_ & ~new_n4115_;
  assign new_n4117_ = new_n971_ & ~new_n4116_;
  assign new_n4118_ = new_n975_ & ~new_n4117_;
  assign new_n4119_ = new_n979_ & ~new_n4118_;
  assign new_n4120_ = new_n983_ & ~new_n4119_;
  assign new_n4121_ = new_n987_ & ~new_n4120_;
  assign new_n4122_ = new_n991_ & ~new_n4121_;
  assign new_n4123_ = new_n995_ & ~new_n4122_;
  assign new_n4124_ = new_n999_ & ~new_n4123_;
  assign new_n4125_ = new_n1003_ & ~new_n4124_;
  assign new_n4126_ = new_n1007_ & ~new_n4125_;
  assign new_n4127_ = new_n1011_ & ~new_n4126_;
  assign new_n4128_ = new_n1015_ & ~new_n4127_;
  assign new_n4129_ = new_n1019_ & ~new_n4128_;
  assign new_n4130_ = new_n1023_ & ~new_n4129_;
  assign new_n4131_ = new_n1027_ & ~new_n4130_;
  assign new_n4132_ = new_n1031_ & ~new_n4131_;
  assign new_n4133_ = new_n1035_ & ~new_n4132_;
  assign new_n4134_ = new_n1039_ & ~new_n4133_;
  assign new_n4135_ = new_n1043_ & ~new_n4134_;
  assign new_n4136_ = new_n1047_ & ~new_n4135_;
  assign new_n4137_ = new_n1051_ & ~new_n4136_;
  assign new_n4138_ = new_n1055_ & ~new_n4137_;
  assign new_n4139_ = new_n1059_ & ~new_n4138_;
  assign new_n4140_ = new_n1574_ & ~new_n4139_;
  assign new_n4141_ = new_n1576_ & ~new_n4140_;
  assign new_n4142_ = new_n1837_ & ~new_n4141_;
  assign new_n4143_ = new_n1068_ & ~new_n4142_;
  assign new_n4144_ = new_n1072_ & ~new_n4143_;
  assign new_n4145_ = new_n1076_ & ~new_n4144_;
  assign new_n4146_ = new_n1080_ & ~new_n4145_;
  assign new_n4147_ = new_n1084_ & ~new_n4146_;
  assign new_n4148_ = new_n1088_ & ~new_n4147_;
  assign new_n4149_ = new_n1092_ & ~new_n4148_;
  assign new_n4150_ = new_n1096_ & ~new_n4149_;
  assign new_n4151_ = new_n1100_ & ~new_n4150_;
  assign new_n4152_ = new_n1104_ & ~new_n4151_;
  assign new_n4153_ = new_n1108_ & ~new_n4152_;
  assign new_n4154_ = new_n1112_ & ~new_n4153_;
  assign new_n4155_ = new_n1116_ & ~new_n4154_;
  assign new_n4156_ = new_n1120_ & ~new_n4155_;
  assign new_n4157_ = new_n1124_ & ~new_n4156_;
  assign new_n4158_ = new_n1128_ & ~new_n4157_;
  assign new_n4159_ = new_n1132_ & ~new_n4158_;
  assign new_n4160_ = new_n1136_ & ~new_n4159_;
  assign new_n4161_ = new_n1140_ & ~new_n4160_;
  assign new_n4162_ = \req[34]  & ~new_n1142_;
  assign \grant[34]  = ~new_n4161_ & new_n4162_;
  assign new_n4164_ = ~new_n479_ & new_n1151_;
  assign new_n4165_ = new_n1156_ & ~new_n4164_;
  assign new_n4166_ = new_n1160_ & ~new_n4165_;
  assign new_n4167_ = new_n1164_ & ~new_n4166_;
  assign new_n4168_ = new_n1168_ & ~new_n4167_;
  assign new_n4169_ = new_n1172_ & ~new_n4168_;
  assign new_n4170_ = new_n1176_ & ~new_n4169_;
  assign new_n4171_ = new_n1180_ & ~new_n4170_;
  assign new_n4172_ = new_n1184_ & ~new_n4171_;
  assign new_n4173_ = new_n1188_ & ~new_n4172_;
  assign new_n4174_ = new_n1192_ & ~new_n4173_;
  assign new_n4175_ = new_n1196_ & ~new_n4174_;
  assign new_n4176_ = new_n1200_ & ~new_n4175_;
  assign new_n4177_ = new_n1204_ & ~new_n4176_;
  assign new_n4178_ = new_n1208_ & ~new_n4177_;
  assign new_n4179_ = new_n1212_ & ~new_n4178_;
  assign new_n4180_ = new_n1216_ & ~new_n4179_;
  assign new_n4181_ = new_n1220_ & ~new_n4180_;
  assign new_n4182_ = new_n1224_ & ~new_n4181_;
  assign new_n4183_ = new_n1228_ & ~new_n4182_;
  assign new_n4184_ = new_n1232_ & ~new_n4183_;
  assign new_n4185_ = new_n1236_ & ~new_n4184_;
  assign new_n4186_ = new_n1240_ & ~new_n4185_;
  assign new_n4187_ = new_n1244_ & ~new_n4186_;
  assign new_n4188_ = new_n1248_ & ~new_n4187_;
  assign new_n4189_ = new_n1252_ & ~new_n4188_;
  assign new_n4190_ = new_n1256_ & ~new_n4189_;
  assign new_n4191_ = new_n1260_ & ~new_n4190_;
  assign new_n4192_ = new_n1264_ & ~new_n4191_;
  assign new_n4193_ = new_n1268_ & ~new_n4192_;
  assign new_n4194_ = new_n1272_ & ~new_n4193_;
  assign new_n4195_ = new_n1276_ & ~new_n4194_;
  assign new_n4196_ = new_n1280_ & ~new_n4195_;
  assign new_n4197_ = new_n1284_ & ~new_n4196_;
  assign new_n4198_ = new_n1288_ & ~new_n4197_;
  assign new_n4199_ = new_n1292_ & ~new_n4198_;
  assign new_n4200_ = new_n1296_ & ~new_n4199_;
  assign new_n4201_ = new_n1300_ & ~new_n4200_;
  assign new_n4202_ = new_n1304_ & ~new_n4201_;
  assign new_n4203_ = new_n1308_ & ~new_n4202_;
  assign new_n4204_ = new_n1312_ & ~new_n4203_;
  assign new_n4205_ = new_n1316_ & ~new_n4204_;
  assign new_n4206_ = new_n1320_ & ~new_n4205_;
  assign new_n4207_ = new_n1324_ & ~new_n4206_;
  assign new_n4208_ = new_n1328_ & ~new_n4207_;
  assign new_n4209_ = new_n1332_ & ~new_n4208_;
  assign new_n4210_ = new_n1336_ & ~new_n4209_;
  assign new_n4211_ = new_n1340_ & ~new_n4210_;
  assign new_n4212_ = new_n1344_ & ~new_n4211_;
  assign new_n4213_ = new_n1348_ & ~new_n4212_;
  assign new_n4214_ = new_n1352_ & ~new_n4213_;
  assign new_n4215_ = new_n1356_ & ~new_n4214_;
  assign new_n4216_ = new_n1360_ & ~new_n4215_;
  assign new_n4217_ = new_n1364_ & ~new_n4216_;
  assign new_n4218_ = new_n1368_ & ~new_n4217_;
  assign new_n4219_ = new_n1372_ & ~new_n4218_;
  assign new_n4220_ = new_n1376_ & ~new_n4219_;
  assign new_n4221_ = new_n1380_ & ~new_n4220_;
  assign new_n4222_ = new_n1384_ & ~new_n4221_;
  assign new_n4223_ = new_n1388_ & ~new_n4222_;
  assign new_n4224_ = new_n1392_ & ~new_n4223_;
  assign new_n4225_ = new_n1396_ & ~new_n4224_;
  assign new_n4226_ = new_n1663_ & ~new_n4225_;
  assign new_n4227_ = new_n392_ & ~new_n4226_;
  assign new_n4228_ = new_n396_ & ~new_n4227_;
  assign new_n4229_ = new_n400_ & ~new_n4228_;
  assign new_n4230_ = new_n404_ & ~new_n4229_;
  assign new_n4231_ = new_n408_ & ~new_n4230_;
  assign new_n4232_ = new_n412_ & ~new_n4231_;
  assign new_n4233_ = new_n416_ & ~new_n4232_;
  assign new_n4234_ = new_n420_ & ~new_n4233_;
  assign new_n4235_ = new_n424_ & ~new_n4234_;
  assign new_n4236_ = new_n428_ & ~new_n4235_;
  assign new_n4237_ = new_n432_ & ~new_n4236_;
  assign new_n4238_ = new_n436_ & ~new_n4237_;
  assign new_n4239_ = new_n440_ & ~new_n4238_;
  assign new_n4240_ = new_n444_ & ~new_n4239_;
  assign new_n4241_ = new_n448_ & ~new_n4240_;
  assign new_n4242_ = new_n452_ & ~new_n4241_;
  assign new_n4243_ = new_n456_ & ~new_n4242_;
  assign new_n4244_ = new_n460_ & ~new_n4243_;
  assign new_n4245_ = new_n464_ & ~new_n4244_;
  assign new_n4246_ = new_n468_ & ~new_n4245_;
  assign new_n4247_ = new_n472_ & ~new_n4246_;
  assign new_n4248_ = \req[35]  & ~new_n474_;
  assign \grant[35]  = ~new_n4247_ & new_n4248_;
  assign new_n4250_ = new_n483_ & ~new_n818_;
  assign new_n4251_ = new_n488_ & ~new_n4250_;
  assign new_n4252_ = new_n492_ & ~new_n4251_;
  assign new_n4253_ = new_n496_ & ~new_n4252_;
  assign new_n4254_ = new_n500_ & ~new_n4253_;
  assign new_n4255_ = new_n504_ & ~new_n4254_;
  assign new_n4256_ = new_n508_ & ~new_n4255_;
  assign new_n4257_ = new_n512_ & ~new_n4256_;
  assign new_n4258_ = new_n516_ & ~new_n4257_;
  assign new_n4259_ = new_n520_ & ~new_n4258_;
  assign new_n4260_ = new_n524_ & ~new_n4259_;
  assign new_n4261_ = new_n528_ & ~new_n4260_;
  assign new_n4262_ = new_n532_ & ~new_n4261_;
  assign new_n4263_ = new_n536_ & ~new_n4262_;
  assign new_n4264_ = new_n540_ & ~new_n4263_;
  assign new_n4265_ = new_n544_ & ~new_n4264_;
  assign new_n4266_ = new_n548_ & ~new_n4265_;
  assign new_n4267_ = new_n552_ & ~new_n4266_;
  assign new_n4268_ = new_n556_ & ~new_n4267_;
  assign new_n4269_ = new_n560_ & ~new_n4268_;
  assign new_n4270_ = new_n564_ & ~new_n4269_;
  assign new_n4271_ = new_n568_ & ~new_n4270_;
  assign new_n4272_ = new_n572_ & ~new_n4271_;
  assign new_n4273_ = new_n576_ & ~new_n4272_;
  assign new_n4274_ = new_n580_ & ~new_n4273_;
  assign new_n4275_ = new_n584_ & ~new_n4274_;
  assign new_n4276_ = new_n588_ & ~new_n4275_;
  assign new_n4277_ = new_n592_ & ~new_n4276_;
  assign new_n4278_ = new_n596_ & ~new_n4277_;
  assign new_n4279_ = new_n600_ & ~new_n4278_;
  assign new_n4280_ = new_n604_ & ~new_n4279_;
  assign new_n4281_ = new_n608_ & ~new_n4280_;
  assign new_n4282_ = new_n612_ & ~new_n4281_;
  assign new_n4283_ = new_n616_ & ~new_n4282_;
  assign new_n4284_ = new_n620_ & ~new_n4283_;
  assign new_n4285_ = new_n624_ & ~new_n4284_;
  assign new_n4286_ = new_n628_ & ~new_n4285_;
  assign new_n4287_ = new_n632_ & ~new_n4286_;
  assign new_n4288_ = new_n636_ & ~new_n4287_;
  assign new_n4289_ = new_n640_ & ~new_n4288_;
  assign new_n4290_ = new_n644_ & ~new_n4289_;
  assign new_n4291_ = new_n648_ & ~new_n4290_;
  assign new_n4292_ = new_n652_ & ~new_n4291_;
  assign new_n4293_ = new_n656_ & ~new_n4292_;
  assign new_n4294_ = new_n660_ & ~new_n4293_;
  assign new_n4295_ = new_n664_ & ~new_n4294_;
  assign new_n4296_ = new_n668_ & ~new_n4295_;
  assign new_n4297_ = new_n672_ & ~new_n4296_;
  assign new_n4298_ = new_n676_ & ~new_n4297_;
  assign new_n4299_ = new_n680_ & ~new_n4298_;
  assign new_n4300_ = new_n684_ & ~new_n4299_;
  assign new_n4301_ = new_n688_ & ~new_n4300_;
  assign new_n4302_ = new_n692_ & ~new_n4301_;
  assign new_n4303_ = new_n696_ & ~new_n4302_;
  assign new_n4304_ = new_n700_ & ~new_n4303_;
  assign new_n4305_ = new_n704_ & ~new_n4304_;
  assign new_n4306_ = new_n708_ & ~new_n4305_;
  assign new_n4307_ = new_n712_ & ~new_n4306_;
  assign new_n4308_ = new_n716_ & ~new_n4307_;
  assign new_n4309_ = new_n720_ & ~new_n4308_;
  assign new_n4310_ = new_n1484_ & ~new_n4309_;
  assign new_n4311_ = new_n1486_ & ~new_n4310_;
  assign new_n4312_ = new_n1750_ & ~new_n4311_;
  assign new_n4313_ = new_n731_ & ~new_n4312_;
  assign new_n4314_ = new_n735_ & ~new_n4313_;
  assign new_n4315_ = new_n739_ & ~new_n4314_;
  assign new_n4316_ = new_n743_ & ~new_n4315_;
  assign new_n4317_ = new_n747_ & ~new_n4316_;
  assign new_n4318_ = new_n751_ & ~new_n4317_;
  assign new_n4319_ = new_n755_ & ~new_n4318_;
  assign new_n4320_ = new_n759_ & ~new_n4319_;
  assign new_n4321_ = new_n763_ & ~new_n4320_;
  assign new_n4322_ = new_n767_ & ~new_n4321_;
  assign new_n4323_ = new_n771_ & ~new_n4322_;
  assign new_n4324_ = new_n775_ & ~new_n4323_;
  assign new_n4325_ = new_n779_ & ~new_n4324_;
  assign new_n4326_ = new_n783_ & ~new_n4325_;
  assign new_n4327_ = new_n787_ & ~new_n4326_;
  assign new_n4328_ = new_n791_ & ~new_n4327_;
  assign new_n4329_ = new_n795_ & ~new_n4328_;
  assign new_n4330_ = new_n799_ & ~new_n4329_;
  assign new_n4331_ = new_n803_ & ~new_n4330_;
  assign new_n4332_ = new_n807_ & ~new_n4331_;
  assign new_n4333_ = new_n811_ & ~new_n4332_;
  assign new_n4334_ = \req[36]  & ~new_n813_;
  assign \grant[36]  = ~new_n4333_ & new_n4334_;
  assign new_n4336_ = new_n822_ & ~new_n1155_;
  assign new_n4337_ = new_n827_ & ~new_n4336_;
  assign new_n4338_ = new_n831_ & ~new_n4337_;
  assign new_n4339_ = new_n835_ & ~new_n4338_;
  assign new_n4340_ = new_n839_ & ~new_n4339_;
  assign new_n4341_ = new_n843_ & ~new_n4340_;
  assign new_n4342_ = new_n847_ & ~new_n4341_;
  assign new_n4343_ = new_n851_ & ~new_n4342_;
  assign new_n4344_ = new_n855_ & ~new_n4343_;
  assign new_n4345_ = new_n859_ & ~new_n4344_;
  assign new_n4346_ = new_n863_ & ~new_n4345_;
  assign new_n4347_ = new_n867_ & ~new_n4346_;
  assign new_n4348_ = new_n871_ & ~new_n4347_;
  assign new_n4349_ = new_n875_ & ~new_n4348_;
  assign new_n4350_ = new_n879_ & ~new_n4349_;
  assign new_n4351_ = new_n883_ & ~new_n4350_;
  assign new_n4352_ = new_n887_ & ~new_n4351_;
  assign new_n4353_ = new_n891_ & ~new_n4352_;
  assign new_n4354_ = new_n895_ & ~new_n4353_;
  assign new_n4355_ = new_n899_ & ~new_n4354_;
  assign new_n4356_ = new_n903_ & ~new_n4355_;
  assign new_n4357_ = new_n907_ & ~new_n4356_;
  assign new_n4358_ = new_n911_ & ~new_n4357_;
  assign new_n4359_ = new_n915_ & ~new_n4358_;
  assign new_n4360_ = new_n919_ & ~new_n4359_;
  assign new_n4361_ = new_n923_ & ~new_n4360_;
  assign new_n4362_ = new_n927_ & ~new_n4361_;
  assign new_n4363_ = new_n931_ & ~new_n4362_;
  assign new_n4364_ = new_n935_ & ~new_n4363_;
  assign new_n4365_ = new_n939_ & ~new_n4364_;
  assign new_n4366_ = new_n943_ & ~new_n4365_;
  assign new_n4367_ = new_n947_ & ~new_n4366_;
  assign new_n4368_ = new_n951_ & ~new_n4367_;
  assign new_n4369_ = new_n955_ & ~new_n4368_;
  assign new_n4370_ = new_n959_ & ~new_n4369_;
  assign new_n4371_ = new_n963_ & ~new_n4370_;
  assign new_n4372_ = new_n967_ & ~new_n4371_;
  assign new_n4373_ = new_n971_ & ~new_n4372_;
  assign new_n4374_ = new_n975_ & ~new_n4373_;
  assign new_n4375_ = new_n979_ & ~new_n4374_;
  assign new_n4376_ = new_n983_ & ~new_n4375_;
  assign new_n4377_ = new_n987_ & ~new_n4376_;
  assign new_n4378_ = new_n991_ & ~new_n4377_;
  assign new_n4379_ = new_n995_ & ~new_n4378_;
  assign new_n4380_ = new_n999_ & ~new_n4379_;
  assign new_n4381_ = new_n1003_ & ~new_n4380_;
  assign new_n4382_ = new_n1007_ & ~new_n4381_;
  assign new_n4383_ = new_n1011_ & ~new_n4382_;
  assign new_n4384_ = new_n1015_ & ~new_n4383_;
  assign new_n4385_ = new_n1019_ & ~new_n4384_;
  assign new_n4386_ = new_n1023_ & ~new_n4385_;
  assign new_n4387_ = new_n1027_ & ~new_n4386_;
  assign new_n4388_ = new_n1031_ & ~new_n4387_;
  assign new_n4389_ = new_n1035_ & ~new_n4388_;
  assign new_n4390_ = new_n1039_ & ~new_n4389_;
  assign new_n4391_ = new_n1043_ & ~new_n4390_;
  assign new_n4392_ = new_n1047_ & ~new_n4391_;
  assign new_n4393_ = new_n1051_ & ~new_n4392_;
  assign new_n4394_ = new_n1055_ & ~new_n4393_;
  assign new_n4395_ = new_n1059_ & ~new_n4394_;
  assign new_n4396_ = new_n1574_ & ~new_n4395_;
  assign new_n4397_ = new_n1576_ & ~new_n4396_;
  assign new_n4398_ = new_n1837_ & ~new_n4397_;
  assign new_n4399_ = new_n1068_ & ~new_n4398_;
  assign new_n4400_ = new_n1072_ & ~new_n4399_;
  assign new_n4401_ = new_n1076_ & ~new_n4400_;
  assign new_n4402_ = new_n1080_ & ~new_n4401_;
  assign new_n4403_ = new_n1084_ & ~new_n4402_;
  assign new_n4404_ = new_n1088_ & ~new_n4403_;
  assign new_n4405_ = new_n1092_ & ~new_n4404_;
  assign new_n4406_ = new_n1096_ & ~new_n4405_;
  assign new_n4407_ = new_n1100_ & ~new_n4406_;
  assign new_n4408_ = new_n1104_ & ~new_n4407_;
  assign new_n4409_ = new_n1108_ & ~new_n4408_;
  assign new_n4410_ = new_n1112_ & ~new_n4409_;
  assign new_n4411_ = new_n1116_ & ~new_n4410_;
  assign new_n4412_ = new_n1120_ & ~new_n4411_;
  assign new_n4413_ = new_n1124_ & ~new_n4412_;
  assign new_n4414_ = new_n1128_ & ~new_n4413_;
  assign new_n4415_ = new_n1132_ & ~new_n4414_;
  assign new_n4416_ = new_n1136_ & ~new_n4415_;
  assign new_n4417_ = new_n1140_ & ~new_n4416_;
  assign new_n4418_ = new_n1144_ & ~new_n4417_;
  assign new_n4419_ = new_n1148_ & ~new_n4418_;
  assign new_n4420_ = \req[37]  & ~new_n1150_;
  assign \grant[37]  = ~new_n4419_ & new_n4420_;
  assign new_n4422_ = ~new_n487_ & new_n1159_;
  assign new_n4423_ = new_n1164_ & ~new_n4422_;
  assign new_n4424_ = new_n1168_ & ~new_n4423_;
  assign new_n4425_ = new_n1172_ & ~new_n4424_;
  assign new_n4426_ = new_n1176_ & ~new_n4425_;
  assign new_n4427_ = new_n1180_ & ~new_n4426_;
  assign new_n4428_ = new_n1184_ & ~new_n4427_;
  assign new_n4429_ = new_n1188_ & ~new_n4428_;
  assign new_n4430_ = new_n1192_ & ~new_n4429_;
  assign new_n4431_ = new_n1196_ & ~new_n4430_;
  assign new_n4432_ = new_n1200_ & ~new_n4431_;
  assign new_n4433_ = new_n1204_ & ~new_n4432_;
  assign new_n4434_ = new_n1208_ & ~new_n4433_;
  assign new_n4435_ = new_n1212_ & ~new_n4434_;
  assign new_n4436_ = new_n1216_ & ~new_n4435_;
  assign new_n4437_ = new_n1220_ & ~new_n4436_;
  assign new_n4438_ = new_n1224_ & ~new_n4437_;
  assign new_n4439_ = new_n1228_ & ~new_n4438_;
  assign new_n4440_ = new_n1232_ & ~new_n4439_;
  assign new_n4441_ = new_n1236_ & ~new_n4440_;
  assign new_n4442_ = new_n1240_ & ~new_n4441_;
  assign new_n4443_ = new_n1244_ & ~new_n4442_;
  assign new_n4444_ = new_n1248_ & ~new_n4443_;
  assign new_n4445_ = new_n1252_ & ~new_n4444_;
  assign new_n4446_ = new_n1256_ & ~new_n4445_;
  assign new_n4447_ = new_n1260_ & ~new_n4446_;
  assign new_n4448_ = new_n1264_ & ~new_n4447_;
  assign new_n4449_ = new_n1268_ & ~new_n4448_;
  assign new_n4450_ = new_n1272_ & ~new_n4449_;
  assign new_n4451_ = new_n1276_ & ~new_n4450_;
  assign new_n4452_ = new_n1280_ & ~new_n4451_;
  assign new_n4453_ = new_n1284_ & ~new_n4452_;
  assign new_n4454_ = new_n1288_ & ~new_n4453_;
  assign new_n4455_ = new_n1292_ & ~new_n4454_;
  assign new_n4456_ = new_n1296_ & ~new_n4455_;
  assign new_n4457_ = new_n1300_ & ~new_n4456_;
  assign new_n4458_ = new_n1304_ & ~new_n4457_;
  assign new_n4459_ = new_n1308_ & ~new_n4458_;
  assign new_n4460_ = new_n1312_ & ~new_n4459_;
  assign new_n4461_ = new_n1316_ & ~new_n4460_;
  assign new_n4462_ = new_n1320_ & ~new_n4461_;
  assign new_n4463_ = new_n1324_ & ~new_n4462_;
  assign new_n4464_ = new_n1328_ & ~new_n4463_;
  assign new_n4465_ = new_n1332_ & ~new_n4464_;
  assign new_n4466_ = new_n1336_ & ~new_n4465_;
  assign new_n4467_ = new_n1340_ & ~new_n4466_;
  assign new_n4468_ = new_n1344_ & ~new_n4467_;
  assign new_n4469_ = new_n1348_ & ~new_n4468_;
  assign new_n4470_ = new_n1352_ & ~new_n4469_;
  assign new_n4471_ = new_n1356_ & ~new_n4470_;
  assign new_n4472_ = new_n1360_ & ~new_n4471_;
  assign new_n4473_ = new_n1364_ & ~new_n4472_;
  assign new_n4474_ = new_n1368_ & ~new_n4473_;
  assign new_n4475_ = new_n1372_ & ~new_n4474_;
  assign new_n4476_ = new_n1376_ & ~new_n4475_;
  assign new_n4477_ = new_n1380_ & ~new_n4476_;
  assign new_n4478_ = new_n1384_ & ~new_n4477_;
  assign new_n4479_ = new_n1388_ & ~new_n4478_;
  assign new_n4480_ = new_n1392_ & ~new_n4479_;
  assign new_n4481_ = new_n1396_ & ~new_n4480_;
  assign new_n4482_ = new_n1663_ & ~new_n4481_;
  assign new_n4483_ = new_n392_ & ~new_n4482_;
  assign new_n4484_ = new_n396_ & ~new_n4483_;
  assign new_n4485_ = new_n400_ & ~new_n4484_;
  assign new_n4486_ = new_n404_ & ~new_n4485_;
  assign new_n4487_ = new_n408_ & ~new_n4486_;
  assign new_n4488_ = new_n412_ & ~new_n4487_;
  assign new_n4489_ = new_n416_ & ~new_n4488_;
  assign new_n4490_ = new_n420_ & ~new_n4489_;
  assign new_n4491_ = new_n424_ & ~new_n4490_;
  assign new_n4492_ = new_n428_ & ~new_n4491_;
  assign new_n4493_ = new_n432_ & ~new_n4492_;
  assign new_n4494_ = new_n436_ & ~new_n4493_;
  assign new_n4495_ = new_n440_ & ~new_n4494_;
  assign new_n4496_ = new_n444_ & ~new_n4495_;
  assign new_n4497_ = new_n448_ & ~new_n4496_;
  assign new_n4498_ = new_n452_ & ~new_n4497_;
  assign new_n4499_ = new_n456_ & ~new_n4498_;
  assign new_n4500_ = new_n460_ & ~new_n4499_;
  assign new_n4501_ = new_n464_ & ~new_n4500_;
  assign new_n4502_ = new_n468_ & ~new_n4501_;
  assign new_n4503_ = new_n472_ & ~new_n4502_;
  assign new_n4504_ = new_n476_ & ~new_n4503_;
  assign new_n4505_ = new_n480_ & ~new_n4504_;
  assign new_n4506_ = \req[38]  & ~new_n482_;
  assign \grant[38]  = ~new_n4505_ & new_n4506_;
  assign new_n4508_ = new_n491_ & ~new_n826_;
  assign new_n4509_ = new_n496_ & ~new_n4508_;
  assign new_n4510_ = new_n500_ & ~new_n4509_;
  assign new_n4511_ = new_n504_ & ~new_n4510_;
  assign new_n4512_ = new_n508_ & ~new_n4511_;
  assign new_n4513_ = new_n512_ & ~new_n4512_;
  assign new_n4514_ = new_n516_ & ~new_n4513_;
  assign new_n4515_ = new_n520_ & ~new_n4514_;
  assign new_n4516_ = new_n524_ & ~new_n4515_;
  assign new_n4517_ = new_n528_ & ~new_n4516_;
  assign new_n4518_ = new_n532_ & ~new_n4517_;
  assign new_n4519_ = new_n536_ & ~new_n4518_;
  assign new_n4520_ = new_n540_ & ~new_n4519_;
  assign new_n4521_ = new_n544_ & ~new_n4520_;
  assign new_n4522_ = new_n548_ & ~new_n4521_;
  assign new_n4523_ = new_n552_ & ~new_n4522_;
  assign new_n4524_ = new_n556_ & ~new_n4523_;
  assign new_n4525_ = new_n560_ & ~new_n4524_;
  assign new_n4526_ = new_n564_ & ~new_n4525_;
  assign new_n4527_ = new_n568_ & ~new_n4526_;
  assign new_n4528_ = new_n572_ & ~new_n4527_;
  assign new_n4529_ = new_n576_ & ~new_n4528_;
  assign new_n4530_ = new_n580_ & ~new_n4529_;
  assign new_n4531_ = new_n584_ & ~new_n4530_;
  assign new_n4532_ = new_n588_ & ~new_n4531_;
  assign new_n4533_ = new_n592_ & ~new_n4532_;
  assign new_n4534_ = new_n596_ & ~new_n4533_;
  assign new_n4535_ = new_n600_ & ~new_n4534_;
  assign new_n4536_ = new_n604_ & ~new_n4535_;
  assign new_n4537_ = new_n608_ & ~new_n4536_;
  assign new_n4538_ = new_n612_ & ~new_n4537_;
  assign new_n4539_ = new_n616_ & ~new_n4538_;
  assign new_n4540_ = new_n620_ & ~new_n4539_;
  assign new_n4541_ = new_n624_ & ~new_n4540_;
  assign new_n4542_ = new_n628_ & ~new_n4541_;
  assign new_n4543_ = new_n632_ & ~new_n4542_;
  assign new_n4544_ = new_n636_ & ~new_n4543_;
  assign new_n4545_ = new_n640_ & ~new_n4544_;
  assign new_n4546_ = new_n644_ & ~new_n4545_;
  assign new_n4547_ = new_n648_ & ~new_n4546_;
  assign new_n4548_ = new_n652_ & ~new_n4547_;
  assign new_n4549_ = new_n656_ & ~new_n4548_;
  assign new_n4550_ = new_n660_ & ~new_n4549_;
  assign new_n4551_ = new_n664_ & ~new_n4550_;
  assign new_n4552_ = new_n668_ & ~new_n4551_;
  assign new_n4553_ = new_n672_ & ~new_n4552_;
  assign new_n4554_ = new_n676_ & ~new_n4553_;
  assign new_n4555_ = new_n680_ & ~new_n4554_;
  assign new_n4556_ = new_n684_ & ~new_n4555_;
  assign new_n4557_ = new_n688_ & ~new_n4556_;
  assign new_n4558_ = new_n692_ & ~new_n4557_;
  assign new_n4559_ = new_n696_ & ~new_n4558_;
  assign new_n4560_ = new_n700_ & ~new_n4559_;
  assign new_n4561_ = new_n704_ & ~new_n4560_;
  assign new_n4562_ = new_n708_ & ~new_n4561_;
  assign new_n4563_ = new_n712_ & ~new_n4562_;
  assign new_n4564_ = new_n716_ & ~new_n4563_;
  assign new_n4565_ = new_n720_ & ~new_n4564_;
  assign new_n4566_ = new_n1484_ & ~new_n4565_;
  assign new_n4567_ = new_n1486_ & ~new_n4566_;
  assign new_n4568_ = new_n1750_ & ~new_n4567_;
  assign new_n4569_ = new_n731_ & ~new_n4568_;
  assign new_n4570_ = new_n735_ & ~new_n4569_;
  assign new_n4571_ = new_n739_ & ~new_n4570_;
  assign new_n4572_ = new_n743_ & ~new_n4571_;
  assign new_n4573_ = new_n747_ & ~new_n4572_;
  assign new_n4574_ = new_n751_ & ~new_n4573_;
  assign new_n4575_ = new_n755_ & ~new_n4574_;
  assign new_n4576_ = new_n759_ & ~new_n4575_;
  assign new_n4577_ = new_n763_ & ~new_n4576_;
  assign new_n4578_ = new_n767_ & ~new_n4577_;
  assign new_n4579_ = new_n771_ & ~new_n4578_;
  assign new_n4580_ = new_n775_ & ~new_n4579_;
  assign new_n4581_ = new_n779_ & ~new_n4580_;
  assign new_n4582_ = new_n783_ & ~new_n4581_;
  assign new_n4583_ = new_n787_ & ~new_n4582_;
  assign new_n4584_ = new_n791_ & ~new_n4583_;
  assign new_n4585_ = new_n795_ & ~new_n4584_;
  assign new_n4586_ = new_n799_ & ~new_n4585_;
  assign new_n4587_ = new_n803_ & ~new_n4586_;
  assign new_n4588_ = new_n807_ & ~new_n4587_;
  assign new_n4589_ = new_n811_ & ~new_n4588_;
  assign new_n4590_ = new_n815_ & ~new_n4589_;
  assign new_n4591_ = new_n819_ & ~new_n4590_;
  assign new_n4592_ = \req[39]  & ~new_n821_;
  assign \grant[39]  = ~new_n4591_ & new_n4592_;
  assign new_n4594_ = new_n830_ & ~new_n1163_;
  assign new_n4595_ = new_n835_ & ~new_n4594_;
  assign new_n4596_ = new_n839_ & ~new_n4595_;
  assign new_n4597_ = new_n843_ & ~new_n4596_;
  assign new_n4598_ = new_n847_ & ~new_n4597_;
  assign new_n4599_ = new_n851_ & ~new_n4598_;
  assign new_n4600_ = new_n855_ & ~new_n4599_;
  assign new_n4601_ = new_n859_ & ~new_n4600_;
  assign new_n4602_ = new_n863_ & ~new_n4601_;
  assign new_n4603_ = new_n867_ & ~new_n4602_;
  assign new_n4604_ = new_n871_ & ~new_n4603_;
  assign new_n4605_ = new_n875_ & ~new_n4604_;
  assign new_n4606_ = new_n879_ & ~new_n4605_;
  assign new_n4607_ = new_n883_ & ~new_n4606_;
  assign new_n4608_ = new_n887_ & ~new_n4607_;
  assign new_n4609_ = new_n891_ & ~new_n4608_;
  assign new_n4610_ = new_n895_ & ~new_n4609_;
  assign new_n4611_ = new_n899_ & ~new_n4610_;
  assign new_n4612_ = new_n903_ & ~new_n4611_;
  assign new_n4613_ = new_n907_ & ~new_n4612_;
  assign new_n4614_ = new_n911_ & ~new_n4613_;
  assign new_n4615_ = new_n915_ & ~new_n4614_;
  assign new_n4616_ = new_n919_ & ~new_n4615_;
  assign new_n4617_ = new_n923_ & ~new_n4616_;
  assign new_n4618_ = new_n927_ & ~new_n4617_;
  assign new_n4619_ = new_n931_ & ~new_n4618_;
  assign new_n4620_ = new_n935_ & ~new_n4619_;
  assign new_n4621_ = new_n939_ & ~new_n4620_;
  assign new_n4622_ = new_n943_ & ~new_n4621_;
  assign new_n4623_ = new_n947_ & ~new_n4622_;
  assign new_n4624_ = new_n951_ & ~new_n4623_;
  assign new_n4625_ = new_n955_ & ~new_n4624_;
  assign new_n4626_ = new_n959_ & ~new_n4625_;
  assign new_n4627_ = new_n963_ & ~new_n4626_;
  assign new_n4628_ = new_n967_ & ~new_n4627_;
  assign new_n4629_ = new_n971_ & ~new_n4628_;
  assign new_n4630_ = new_n975_ & ~new_n4629_;
  assign new_n4631_ = new_n979_ & ~new_n4630_;
  assign new_n4632_ = new_n983_ & ~new_n4631_;
  assign new_n4633_ = new_n987_ & ~new_n4632_;
  assign new_n4634_ = new_n991_ & ~new_n4633_;
  assign new_n4635_ = new_n995_ & ~new_n4634_;
  assign new_n4636_ = new_n999_ & ~new_n4635_;
  assign new_n4637_ = new_n1003_ & ~new_n4636_;
  assign new_n4638_ = new_n1007_ & ~new_n4637_;
  assign new_n4639_ = new_n1011_ & ~new_n4638_;
  assign new_n4640_ = new_n1015_ & ~new_n4639_;
  assign new_n4641_ = new_n1019_ & ~new_n4640_;
  assign new_n4642_ = new_n1023_ & ~new_n4641_;
  assign new_n4643_ = new_n1027_ & ~new_n4642_;
  assign new_n4644_ = new_n1031_ & ~new_n4643_;
  assign new_n4645_ = new_n1035_ & ~new_n4644_;
  assign new_n4646_ = new_n1039_ & ~new_n4645_;
  assign new_n4647_ = new_n1043_ & ~new_n4646_;
  assign new_n4648_ = new_n1047_ & ~new_n4647_;
  assign new_n4649_ = new_n1051_ & ~new_n4648_;
  assign new_n4650_ = new_n1055_ & ~new_n4649_;
  assign new_n4651_ = new_n1059_ & ~new_n4650_;
  assign new_n4652_ = new_n1574_ & ~new_n4651_;
  assign new_n4653_ = new_n1576_ & ~new_n4652_;
  assign new_n4654_ = new_n1837_ & ~new_n4653_;
  assign new_n4655_ = new_n1068_ & ~new_n4654_;
  assign new_n4656_ = new_n1072_ & ~new_n4655_;
  assign new_n4657_ = new_n1076_ & ~new_n4656_;
  assign new_n4658_ = new_n1080_ & ~new_n4657_;
  assign new_n4659_ = new_n1084_ & ~new_n4658_;
  assign new_n4660_ = new_n1088_ & ~new_n4659_;
  assign new_n4661_ = new_n1092_ & ~new_n4660_;
  assign new_n4662_ = new_n1096_ & ~new_n4661_;
  assign new_n4663_ = new_n1100_ & ~new_n4662_;
  assign new_n4664_ = new_n1104_ & ~new_n4663_;
  assign new_n4665_ = new_n1108_ & ~new_n4664_;
  assign new_n4666_ = new_n1112_ & ~new_n4665_;
  assign new_n4667_ = new_n1116_ & ~new_n4666_;
  assign new_n4668_ = new_n1120_ & ~new_n4667_;
  assign new_n4669_ = new_n1124_ & ~new_n4668_;
  assign new_n4670_ = new_n1128_ & ~new_n4669_;
  assign new_n4671_ = new_n1132_ & ~new_n4670_;
  assign new_n4672_ = new_n1136_ & ~new_n4671_;
  assign new_n4673_ = new_n1140_ & ~new_n4672_;
  assign new_n4674_ = new_n1144_ & ~new_n4673_;
  assign new_n4675_ = new_n1148_ & ~new_n4674_;
  assign new_n4676_ = new_n1152_ & ~new_n4675_;
  assign new_n4677_ = new_n1156_ & ~new_n4676_;
  assign new_n4678_ = \req[40]  & ~new_n1158_;
  assign \grant[40]  = ~new_n4677_ & new_n4678_;
  assign new_n4680_ = ~new_n495_ & new_n1167_;
  assign new_n4681_ = new_n1172_ & ~new_n4680_;
  assign new_n4682_ = new_n1176_ & ~new_n4681_;
  assign new_n4683_ = new_n1180_ & ~new_n4682_;
  assign new_n4684_ = new_n1184_ & ~new_n4683_;
  assign new_n4685_ = new_n1188_ & ~new_n4684_;
  assign new_n4686_ = new_n1192_ & ~new_n4685_;
  assign new_n4687_ = new_n1196_ & ~new_n4686_;
  assign new_n4688_ = new_n1200_ & ~new_n4687_;
  assign new_n4689_ = new_n1204_ & ~new_n4688_;
  assign new_n4690_ = new_n1208_ & ~new_n4689_;
  assign new_n4691_ = new_n1212_ & ~new_n4690_;
  assign new_n4692_ = new_n1216_ & ~new_n4691_;
  assign new_n4693_ = new_n1220_ & ~new_n4692_;
  assign new_n4694_ = new_n1224_ & ~new_n4693_;
  assign new_n4695_ = new_n1228_ & ~new_n4694_;
  assign new_n4696_ = new_n1232_ & ~new_n4695_;
  assign new_n4697_ = new_n1236_ & ~new_n4696_;
  assign new_n4698_ = new_n1240_ & ~new_n4697_;
  assign new_n4699_ = new_n1244_ & ~new_n4698_;
  assign new_n4700_ = new_n1248_ & ~new_n4699_;
  assign new_n4701_ = new_n1252_ & ~new_n4700_;
  assign new_n4702_ = new_n1256_ & ~new_n4701_;
  assign new_n4703_ = new_n1260_ & ~new_n4702_;
  assign new_n4704_ = new_n1264_ & ~new_n4703_;
  assign new_n4705_ = new_n1268_ & ~new_n4704_;
  assign new_n4706_ = new_n1272_ & ~new_n4705_;
  assign new_n4707_ = new_n1276_ & ~new_n4706_;
  assign new_n4708_ = new_n1280_ & ~new_n4707_;
  assign new_n4709_ = new_n1284_ & ~new_n4708_;
  assign new_n4710_ = new_n1288_ & ~new_n4709_;
  assign new_n4711_ = new_n1292_ & ~new_n4710_;
  assign new_n4712_ = new_n1296_ & ~new_n4711_;
  assign new_n4713_ = new_n1300_ & ~new_n4712_;
  assign new_n4714_ = new_n1304_ & ~new_n4713_;
  assign new_n4715_ = new_n1308_ & ~new_n4714_;
  assign new_n4716_ = new_n1312_ & ~new_n4715_;
  assign new_n4717_ = new_n1316_ & ~new_n4716_;
  assign new_n4718_ = new_n1320_ & ~new_n4717_;
  assign new_n4719_ = new_n1324_ & ~new_n4718_;
  assign new_n4720_ = new_n1328_ & ~new_n4719_;
  assign new_n4721_ = new_n1332_ & ~new_n4720_;
  assign new_n4722_ = new_n1336_ & ~new_n4721_;
  assign new_n4723_ = new_n1340_ & ~new_n4722_;
  assign new_n4724_ = new_n1344_ & ~new_n4723_;
  assign new_n4725_ = new_n1348_ & ~new_n4724_;
  assign new_n4726_ = new_n1352_ & ~new_n4725_;
  assign new_n4727_ = new_n1356_ & ~new_n4726_;
  assign new_n4728_ = new_n1360_ & ~new_n4727_;
  assign new_n4729_ = new_n1364_ & ~new_n4728_;
  assign new_n4730_ = new_n1368_ & ~new_n4729_;
  assign new_n4731_ = new_n1372_ & ~new_n4730_;
  assign new_n4732_ = new_n1376_ & ~new_n4731_;
  assign new_n4733_ = new_n1380_ & ~new_n4732_;
  assign new_n4734_ = new_n1384_ & ~new_n4733_;
  assign new_n4735_ = new_n1388_ & ~new_n4734_;
  assign new_n4736_ = new_n1392_ & ~new_n4735_;
  assign new_n4737_ = new_n1396_ & ~new_n4736_;
  assign new_n4738_ = new_n1663_ & ~new_n4737_;
  assign new_n4739_ = new_n392_ & ~new_n4738_;
  assign new_n4740_ = new_n396_ & ~new_n4739_;
  assign new_n4741_ = new_n400_ & ~new_n4740_;
  assign new_n4742_ = new_n404_ & ~new_n4741_;
  assign new_n4743_ = new_n408_ & ~new_n4742_;
  assign new_n4744_ = new_n412_ & ~new_n4743_;
  assign new_n4745_ = new_n416_ & ~new_n4744_;
  assign new_n4746_ = new_n420_ & ~new_n4745_;
  assign new_n4747_ = new_n424_ & ~new_n4746_;
  assign new_n4748_ = new_n428_ & ~new_n4747_;
  assign new_n4749_ = new_n432_ & ~new_n4748_;
  assign new_n4750_ = new_n436_ & ~new_n4749_;
  assign new_n4751_ = new_n440_ & ~new_n4750_;
  assign new_n4752_ = new_n444_ & ~new_n4751_;
  assign new_n4753_ = new_n448_ & ~new_n4752_;
  assign new_n4754_ = new_n452_ & ~new_n4753_;
  assign new_n4755_ = new_n456_ & ~new_n4754_;
  assign new_n4756_ = new_n460_ & ~new_n4755_;
  assign new_n4757_ = new_n464_ & ~new_n4756_;
  assign new_n4758_ = new_n468_ & ~new_n4757_;
  assign new_n4759_ = new_n472_ & ~new_n4758_;
  assign new_n4760_ = new_n476_ & ~new_n4759_;
  assign new_n4761_ = new_n480_ & ~new_n4760_;
  assign new_n4762_ = new_n484_ & ~new_n4761_;
  assign new_n4763_ = new_n488_ & ~new_n4762_;
  assign new_n4764_ = \req[41]  & ~new_n490_;
  assign \grant[41]  = ~new_n4763_ & new_n4764_;
  assign new_n4766_ = new_n499_ & ~new_n834_;
  assign new_n4767_ = new_n504_ & ~new_n4766_;
  assign new_n4768_ = new_n508_ & ~new_n4767_;
  assign new_n4769_ = new_n512_ & ~new_n4768_;
  assign new_n4770_ = new_n516_ & ~new_n4769_;
  assign new_n4771_ = new_n520_ & ~new_n4770_;
  assign new_n4772_ = new_n524_ & ~new_n4771_;
  assign new_n4773_ = new_n528_ & ~new_n4772_;
  assign new_n4774_ = new_n532_ & ~new_n4773_;
  assign new_n4775_ = new_n536_ & ~new_n4774_;
  assign new_n4776_ = new_n540_ & ~new_n4775_;
  assign new_n4777_ = new_n544_ & ~new_n4776_;
  assign new_n4778_ = new_n548_ & ~new_n4777_;
  assign new_n4779_ = new_n552_ & ~new_n4778_;
  assign new_n4780_ = new_n556_ & ~new_n4779_;
  assign new_n4781_ = new_n560_ & ~new_n4780_;
  assign new_n4782_ = new_n564_ & ~new_n4781_;
  assign new_n4783_ = new_n568_ & ~new_n4782_;
  assign new_n4784_ = new_n572_ & ~new_n4783_;
  assign new_n4785_ = new_n576_ & ~new_n4784_;
  assign new_n4786_ = new_n580_ & ~new_n4785_;
  assign new_n4787_ = new_n584_ & ~new_n4786_;
  assign new_n4788_ = new_n588_ & ~new_n4787_;
  assign new_n4789_ = new_n592_ & ~new_n4788_;
  assign new_n4790_ = new_n596_ & ~new_n4789_;
  assign new_n4791_ = new_n600_ & ~new_n4790_;
  assign new_n4792_ = new_n604_ & ~new_n4791_;
  assign new_n4793_ = new_n608_ & ~new_n4792_;
  assign new_n4794_ = new_n612_ & ~new_n4793_;
  assign new_n4795_ = new_n616_ & ~new_n4794_;
  assign new_n4796_ = new_n620_ & ~new_n4795_;
  assign new_n4797_ = new_n624_ & ~new_n4796_;
  assign new_n4798_ = new_n628_ & ~new_n4797_;
  assign new_n4799_ = new_n632_ & ~new_n4798_;
  assign new_n4800_ = new_n636_ & ~new_n4799_;
  assign new_n4801_ = new_n640_ & ~new_n4800_;
  assign new_n4802_ = new_n644_ & ~new_n4801_;
  assign new_n4803_ = new_n648_ & ~new_n4802_;
  assign new_n4804_ = new_n652_ & ~new_n4803_;
  assign new_n4805_ = new_n656_ & ~new_n4804_;
  assign new_n4806_ = new_n660_ & ~new_n4805_;
  assign new_n4807_ = new_n664_ & ~new_n4806_;
  assign new_n4808_ = new_n668_ & ~new_n4807_;
  assign new_n4809_ = new_n672_ & ~new_n4808_;
  assign new_n4810_ = new_n676_ & ~new_n4809_;
  assign new_n4811_ = new_n680_ & ~new_n4810_;
  assign new_n4812_ = new_n684_ & ~new_n4811_;
  assign new_n4813_ = new_n688_ & ~new_n4812_;
  assign new_n4814_ = new_n692_ & ~new_n4813_;
  assign new_n4815_ = new_n696_ & ~new_n4814_;
  assign new_n4816_ = new_n700_ & ~new_n4815_;
  assign new_n4817_ = new_n704_ & ~new_n4816_;
  assign new_n4818_ = new_n708_ & ~new_n4817_;
  assign new_n4819_ = new_n712_ & ~new_n4818_;
  assign new_n4820_ = new_n716_ & ~new_n4819_;
  assign new_n4821_ = new_n720_ & ~new_n4820_;
  assign new_n4822_ = new_n1484_ & ~new_n4821_;
  assign new_n4823_ = new_n1486_ & ~new_n4822_;
  assign new_n4824_ = new_n1750_ & ~new_n4823_;
  assign new_n4825_ = new_n731_ & ~new_n4824_;
  assign new_n4826_ = new_n735_ & ~new_n4825_;
  assign new_n4827_ = new_n739_ & ~new_n4826_;
  assign new_n4828_ = new_n743_ & ~new_n4827_;
  assign new_n4829_ = new_n747_ & ~new_n4828_;
  assign new_n4830_ = new_n751_ & ~new_n4829_;
  assign new_n4831_ = new_n755_ & ~new_n4830_;
  assign new_n4832_ = new_n759_ & ~new_n4831_;
  assign new_n4833_ = new_n763_ & ~new_n4832_;
  assign new_n4834_ = new_n767_ & ~new_n4833_;
  assign new_n4835_ = new_n771_ & ~new_n4834_;
  assign new_n4836_ = new_n775_ & ~new_n4835_;
  assign new_n4837_ = new_n779_ & ~new_n4836_;
  assign new_n4838_ = new_n783_ & ~new_n4837_;
  assign new_n4839_ = new_n787_ & ~new_n4838_;
  assign new_n4840_ = new_n791_ & ~new_n4839_;
  assign new_n4841_ = new_n795_ & ~new_n4840_;
  assign new_n4842_ = new_n799_ & ~new_n4841_;
  assign new_n4843_ = new_n803_ & ~new_n4842_;
  assign new_n4844_ = new_n807_ & ~new_n4843_;
  assign new_n4845_ = new_n811_ & ~new_n4844_;
  assign new_n4846_ = new_n815_ & ~new_n4845_;
  assign new_n4847_ = new_n819_ & ~new_n4846_;
  assign new_n4848_ = new_n823_ & ~new_n4847_;
  assign new_n4849_ = new_n827_ & ~new_n4848_;
  assign new_n4850_ = \req[42]  & ~new_n829_;
  assign \grant[42]  = ~new_n4849_ & new_n4850_;
  assign new_n4852_ = new_n838_ & ~new_n1171_;
  assign new_n4853_ = new_n843_ & ~new_n4852_;
  assign new_n4854_ = new_n847_ & ~new_n4853_;
  assign new_n4855_ = new_n851_ & ~new_n4854_;
  assign new_n4856_ = new_n855_ & ~new_n4855_;
  assign new_n4857_ = new_n859_ & ~new_n4856_;
  assign new_n4858_ = new_n863_ & ~new_n4857_;
  assign new_n4859_ = new_n867_ & ~new_n4858_;
  assign new_n4860_ = new_n871_ & ~new_n4859_;
  assign new_n4861_ = new_n875_ & ~new_n4860_;
  assign new_n4862_ = new_n879_ & ~new_n4861_;
  assign new_n4863_ = new_n883_ & ~new_n4862_;
  assign new_n4864_ = new_n887_ & ~new_n4863_;
  assign new_n4865_ = new_n891_ & ~new_n4864_;
  assign new_n4866_ = new_n895_ & ~new_n4865_;
  assign new_n4867_ = new_n899_ & ~new_n4866_;
  assign new_n4868_ = new_n903_ & ~new_n4867_;
  assign new_n4869_ = new_n907_ & ~new_n4868_;
  assign new_n4870_ = new_n911_ & ~new_n4869_;
  assign new_n4871_ = new_n915_ & ~new_n4870_;
  assign new_n4872_ = new_n919_ & ~new_n4871_;
  assign new_n4873_ = new_n923_ & ~new_n4872_;
  assign new_n4874_ = new_n927_ & ~new_n4873_;
  assign new_n4875_ = new_n931_ & ~new_n4874_;
  assign new_n4876_ = new_n935_ & ~new_n4875_;
  assign new_n4877_ = new_n939_ & ~new_n4876_;
  assign new_n4878_ = new_n943_ & ~new_n4877_;
  assign new_n4879_ = new_n947_ & ~new_n4878_;
  assign new_n4880_ = new_n951_ & ~new_n4879_;
  assign new_n4881_ = new_n955_ & ~new_n4880_;
  assign new_n4882_ = new_n959_ & ~new_n4881_;
  assign new_n4883_ = new_n963_ & ~new_n4882_;
  assign new_n4884_ = new_n967_ & ~new_n4883_;
  assign new_n4885_ = new_n971_ & ~new_n4884_;
  assign new_n4886_ = new_n975_ & ~new_n4885_;
  assign new_n4887_ = new_n979_ & ~new_n4886_;
  assign new_n4888_ = new_n983_ & ~new_n4887_;
  assign new_n4889_ = new_n987_ & ~new_n4888_;
  assign new_n4890_ = new_n991_ & ~new_n4889_;
  assign new_n4891_ = new_n995_ & ~new_n4890_;
  assign new_n4892_ = new_n999_ & ~new_n4891_;
  assign new_n4893_ = new_n1003_ & ~new_n4892_;
  assign new_n4894_ = new_n1007_ & ~new_n4893_;
  assign new_n4895_ = new_n1011_ & ~new_n4894_;
  assign new_n4896_ = new_n1015_ & ~new_n4895_;
  assign new_n4897_ = new_n1019_ & ~new_n4896_;
  assign new_n4898_ = new_n1023_ & ~new_n4897_;
  assign new_n4899_ = new_n1027_ & ~new_n4898_;
  assign new_n4900_ = new_n1031_ & ~new_n4899_;
  assign new_n4901_ = new_n1035_ & ~new_n4900_;
  assign new_n4902_ = new_n1039_ & ~new_n4901_;
  assign new_n4903_ = new_n1043_ & ~new_n4902_;
  assign new_n4904_ = new_n1047_ & ~new_n4903_;
  assign new_n4905_ = new_n1051_ & ~new_n4904_;
  assign new_n4906_ = new_n1055_ & ~new_n4905_;
  assign new_n4907_ = new_n1059_ & ~new_n4906_;
  assign new_n4908_ = new_n1574_ & ~new_n4907_;
  assign new_n4909_ = new_n1576_ & ~new_n4908_;
  assign new_n4910_ = new_n1837_ & ~new_n4909_;
  assign new_n4911_ = new_n1068_ & ~new_n4910_;
  assign new_n4912_ = new_n1072_ & ~new_n4911_;
  assign new_n4913_ = new_n1076_ & ~new_n4912_;
  assign new_n4914_ = new_n1080_ & ~new_n4913_;
  assign new_n4915_ = new_n1084_ & ~new_n4914_;
  assign new_n4916_ = new_n1088_ & ~new_n4915_;
  assign new_n4917_ = new_n1092_ & ~new_n4916_;
  assign new_n4918_ = new_n1096_ & ~new_n4917_;
  assign new_n4919_ = new_n1100_ & ~new_n4918_;
  assign new_n4920_ = new_n1104_ & ~new_n4919_;
  assign new_n4921_ = new_n1108_ & ~new_n4920_;
  assign new_n4922_ = new_n1112_ & ~new_n4921_;
  assign new_n4923_ = new_n1116_ & ~new_n4922_;
  assign new_n4924_ = new_n1120_ & ~new_n4923_;
  assign new_n4925_ = new_n1124_ & ~new_n4924_;
  assign new_n4926_ = new_n1128_ & ~new_n4925_;
  assign new_n4927_ = new_n1132_ & ~new_n4926_;
  assign new_n4928_ = new_n1136_ & ~new_n4927_;
  assign new_n4929_ = new_n1140_ & ~new_n4928_;
  assign new_n4930_ = new_n1144_ & ~new_n4929_;
  assign new_n4931_ = new_n1148_ & ~new_n4930_;
  assign new_n4932_ = new_n1152_ & ~new_n4931_;
  assign new_n4933_ = new_n1156_ & ~new_n4932_;
  assign new_n4934_ = new_n1160_ & ~new_n4933_;
  assign new_n4935_ = new_n1164_ & ~new_n4934_;
  assign new_n4936_ = \req[43]  & ~new_n1166_;
  assign \grant[43]  = ~new_n4935_ & new_n4936_;
  assign new_n4938_ = ~new_n503_ & new_n1175_;
  assign new_n4939_ = new_n1180_ & ~new_n4938_;
  assign new_n4940_ = new_n1184_ & ~new_n4939_;
  assign new_n4941_ = new_n1188_ & ~new_n4940_;
  assign new_n4942_ = new_n1192_ & ~new_n4941_;
  assign new_n4943_ = new_n1196_ & ~new_n4942_;
  assign new_n4944_ = new_n1200_ & ~new_n4943_;
  assign new_n4945_ = new_n1204_ & ~new_n4944_;
  assign new_n4946_ = new_n1208_ & ~new_n4945_;
  assign new_n4947_ = new_n1212_ & ~new_n4946_;
  assign new_n4948_ = new_n1216_ & ~new_n4947_;
  assign new_n4949_ = new_n1220_ & ~new_n4948_;
  assign new_n4950_ = new_n1224_ & ~new_n4949_;
  assign new_n4951_ = new_n1228_ & ~new_n4950_;
  assign new_n4952_ = new_n1232_ & ~new_n4951_;
  assign new_n4953_ = new_n1236_ & ~new_n4952_;
  assign new_n4954_ = new_n1240_ & ~new_n4953_;
  assign new_n4955_ = new_n1244_ & ~new_n4954_;
  assign new_n4956_ = new_n1248_ & ~new_n4955_;
  assign new_n4957_ = new_n1252_ & ~new_n4956_;
  assign new_n4958_ = new_n1256_ & ~new_n4957_;
  assign new_n4959_ = new_n1260_ & ~new_n4958_;
  assign new_n4960_ = new_n1264_ & ~new_n4959_;
  assign new_n4961_ = new_n1268_ & ~new_n4960_;
  assign new_n4962_ = new_n1272_ & ~new_n4961_;
  assign new_n4963_ = new_n1276_ & ~new_n4962_;
  assign new_n4964_ = new_n1280_ & ~new_n4963_;
  assign new_n4965_ = new_n1284_ & ~new_n4964_;
  assign new_n4966_ = new_n1288_ & ~new_n4965_;
  assign new_n4967_ = new_n1292_ & ~new_n4966_;
  assign new_n4968_ = new_n1296_ & ~new_n4967_;
  assign new_n4969_ = new_n1300_ & ~new_n4968_;
  assign new_n4970_ = new_n1304_ & ~new_n4969_;
  assign new_n4971_ = new_n1308_ & ~new_n4970_;
  assign new_n4972_ = new_n1312_ & ~new_n4971_;
  assign new_n4973_ = new_n1316_ & ~new_n4972_;
  assign new_n4974_ = new_n1320_ & ~new_n4973_;
  assign new_n4975_ = new_n1324_ & ~new_n4974_;
  assign new_n4976_ = new_n1328_ & ~new_n4975_;
  assign new_n4977_ = new_n1332_ & ~new_n4976_;
  assign new_n4978_ = new_n1336_ & ~new_n4977_;
  assign new_n4979_ = new_n1340_ & ~new_n4978_;
  assign new_n4980_ = new_n1344_ & ~new_n4979_;
  assign new_n4981_ = new_n1348_ & ~new_n4980_;
  assign new_n4982_ = new_n1352_ & ~new_n4981_;
  assign new_n4983_ = new_n1356_ & ~new_n4982_;
  assign new_n4984_ = new_n1360_ & ~new_n4983_;
  assign new_n4985_ = new_n1364_ & ~new_n4984_;
  assign new_n4986_ = new_n1368_ & ~new_n4985_;
  assign new_n4987_ = new_n1372_ & ~new_n4986_;
  assign new_n4988_ = new_n1376_ & ~new_n4987_;
  assign new_n4989_ = new_n1380_ & ~new_n4988_;
  assign new_n4990_ = new_n1384_ & ~new_n4989_;
  assign new_n4991_ = new_n1388_ & ~new_n4990_;
  assign new_n4992_ = new_n1392_ & ~new_n4991_;
  assign new_n4993_ = new_n1396_ & ~new_n4992_;
  assign new_n4994_ = new_n1663_ & ~new_n4993_;
  assign new_n4995_ = new_n392_ & ~new_n4994_;
  assign new_n4996_ = new_n396_ & ~new_n4995_;
  assign new_n4997_ = new_n400_ & ~new_n4996_;
  assign new_n4998_ = new_n404_ & ~new_n4997_;
  assign new_n4999_ = new_n408_ & ~new_n4998_;
  assign new_n5000_ = new_n412_ & ~new_n4999_;
  assign new_n5001_ = new_n416_ & ~new_n5000_;
  assign new_n5002_ = new_n420_ & ~new_n5001_;
  assign new_n5003_ = new_n424_ & ~new_n5002_;
  assign new_n5004_ = new_n428_ & ~new_n5003_;
  assign new_n5005_ = new_n432_ & ~new_n5004_;
  assign new_n5006_ = new_n436_ & ~new_n5005_;
  assign new_n5007_ = new_n440_ & ~new_n5006_;
  assign new_n5008_ = new_n444_ & ~new_n5007_;
  assign new_n5009_ = new_n448_ & ~new_n5008_;
  assign new_n5010_ = new_n452_ & ~new_n5009_;
  assign new_n5011_ = new_n456_ & ~new_n5010_;
  assign new_n5012_ = new_n460_ & ~new_n5011_;
  assign new_n5013_ = new_n464_ & ~new_n5012_;
  assign new_n5014_ = new_n468_ & ~new_n5013_;
  assign new_n5015_ = new_n472_ & ~new_n5014_;
  assign new_n5016_ = new_n476_ & ~new_n5015_;
  assign new_n5017_ = new_n480_ & ~new_n5016_;
  assign new_n5018_ = new_n484_ & ~new_n5017_;
  assign new_n5019_ = new_n488_ & ~new_n5018_;
  assign new_n5020_ = new_n492_ & ~new_n5019_;
  assign new_n5021_ = new_n496_ & ~new_n5020_;
  assign new_n5022_ = \req[44]  & ~new_n498_;
  assign \grant[44]  = ~new_n5021_ & new_n5022_;
  assign new_n5024_ = new_n507_ & ~new_n842_;
  assign new_n5025_ = new_n512_ & ~new_n5024_;
  assign new_n5026_ = new_n516_ & ~new_n5025_;
  assign new_n5027_ = new_n520_ & ~new_n5026_;
  assign new_n5028_ = new_n524_ & ~new_n5027_;
  assign new_n5029_ = new_n528_ & ~new_n5028_;
  assign new_n5030_ = new_n532_ & ~new_n5029_;
  assign new_n5031_ = new_n536_ & ~new_n5030_;
  assign new_n5032_ = new_n540_ & ~new_n5031_;
  assign new_n5033_ = new_n544_ & ~new_n5032_;
  assign new_n5034_ = new_n548_ & ~new_n5033_;
  assign new_n5035_ = new_n552_ & ~new_n5034_;
  assign new_n5036_ = new_n556_ & ~new_n5035_;
  assign new_n5037_ = new_n560_ & ~new_n5036_;
  assign new_n5038_ = new_n564_ & ~new_n5037_;
  assign new_n5039_ = new_n568_ & ~new_n5038_;
  assign new_n5040_ = new_n572_ & ~new_n5039_;
  assign new_n5041_ = new_n576_ & ~new_n5040_;
  assign new_n5042_ = new_n580_ & ~new_n5041_;
  assign new_n5043_ = new_n584_ & ~new_n5042_;
  assign new_n5044_ = new_n588_ & ~new_n5043_;
  assign new_n5045_ = new_n592_ & ~new_n5044_;
  assign new_n5046_ = new_n596_ & ~new_n5045_;
  assign new_n5047_ = new_n600_ & ~new_n5046_;
  assign new_n5048_ = new_n604_ & ~new_n5047_;
  assign new_n5049_ = new_n608_ & ~new_n5048_;
  assign new_n5050_ = new_n612_ & ~new_n5049_;
  assign new_n5051_ = new_n616_ & ~new_n5050_;
  assign new_n5052_ = new_n620_ & ~new_n5051_;
  assign new_n5053_ = new_n624_ & ~new_n5052_;
  assign new_n5054_ = new_n628_ & ~new_n5053_;
  assign new_n5055_ = new_n632_ & ~new_n5054_;
  assign new_n5056_ = new_n636_ & ~new_n5055_;
  assign new_n5057_ = new_n640_ & ~new_n5056_;
  assign new_n5058_ = new_n644_ & ~new_n5057_;
  assign new_n5059_ = new_n648_ & ~new_n5058_;
  assign new_n5060_ = new_n652_ & ~new_n5059_;
  assign new_n5061_ = new_n656_ & ~new_n5060_;
  assign new_n5062_ = new_n660_ & ~new_n5061_;
  assign new_n5063_ = new_n664_ & ~new_n5062_;
  assign new_n5064_ = new_n668_ & ~new_n5063_;
  assign new_n5065_ = new_n672_ & ~new_n5064_;
  assign new_n5066_ = new_n676_ & ~new_n5065_;
  assign new_n5067_ = new_n680_ & ~new_n5066_;
  assign new_n5068_ = new_n684_ & ~new_n5067_;
  assign new_n5069_ = new_n688_ & ~new_n5068_;
  assign new_n5070_ = new_n692_ & ~new_n5069_;
  assign new_n5071_ = new_n696_ & ~new_n5070_;
  assign new_n5072_ = new_n700_ & ~new_n5071_;
  assign new_n5073_ = new_n704_ & ~new_n5072_;
  assign new_n5074_ = new_n708_ & ~new_n5073_;
  assign new_n5075_ = new_n712_ & ~new_n5074_;
  assign new_n5076_ = new_n716_ & ~new_n5075_;
  assign new_n5077_ = new_n720_ & ~new_n5076_;
  assign new_n5078_ = new_n1484_ & ~new_n5077_;
  assign new_n5079_ = new_n1486_ & ~new_n5078_;
  assign new_n5080_ = new_n1750_ & ~new_n5079_;
  assign new_n5081_ = new_n731_ & ~new_n5080_;
  assign new_n5082_ = new_n735_ & ~new_n5081_;
  assign new_n5083_ = new_n739_ & ~new_n5082_;
  assign new_n5084_ = new_n743_ & ~new_n5083_;
  assign new_n5085_ = new_n747_ & ~new_n5084_;
  assign new_n5086_ = new_n751_ & ~new_n5085_;
  assign new_n5087_ = new_n755_ & ~new_n5086_;
  assign new_n5088_ = new_n759_ & ~new_n5087_;
  assign new_n5089_ = new_n763_ & ~new_n5088_;
  assign new_n5090_ = new_n767_ & ~new_n5089_;
  assign new_n5091_ = new_n771_ & ~new_n5090_;
  assign new_n5092_ = new_n775_ & ~new_n5091_;
  assign new_n5093_ = new_n779_ & ~new_n5092_;
  assign new_n5094_ = new_n783_ & ~new_n5093_;
  assign new_n5095_ = new_n787_ & ~new_n5094_;
  assign new_n5096_ = new_n791_ & ~new_n5095_;
  assign new_n5097_ = new_n795_ & ~new_n5096_;
  assign new_n5098_ = new_n799_ & ~new_n5097_;
  assign new_n5099_ = new_n803_ & ~new_n5098_;
  assign new_n5100_ = new_n807_ & ~new_n5099_;
  assign new_n5101_ = new_n811_ & ~new_n5100_;
  assign new_n5102_ = new_n815_ & ~new_n5101_;
  assign new_n5103_ = new_n819_ & ~new_n5102_;
  assign new_n5104_ = new_n823_ & ~new_n5103_;
  assign new_n5105_ = new_n827_ & ~new_n5104_;
  assign new_n5106_ = new_n831_ & ~new_n5105_;
  assign new_n5107_ = new_n835_ & ~new_n5106_;
  assign new_n5108_ = \req[45]  & ~new_n837_;
  assign \grant[45]  = ~new_n5107_ & new_n5108_;
  assign new_n5110_ = new_n846_ & ~new_n1179_;
  assign new_n5111_ = new_n851_ & ~new_n5110_;
  assign new_n5112_ = new_n855_ & ~new_n5111_;
  assign new_n5113_ = new_n859_ & ~new_n5112_;
  assign new_n5114_ = new_n863_ & ~new_n5113_;
  assign new_n5115_ = new_n867_ & ~new_n5114_;
  assign new_n5116_ = new_n871_ & ~new_n5115_;
  assign new_n5117_ = new_n875_ & ~new_n5116_;
  assign new_n5118_ = new_n879_ & ~new_n5117_;
  assign new_n5119_ = new_n883_ & ~new_n5118_;
  assign new_n5120_ = new_n887_ & ~new_n5119_;
  assign new_n5121_ = new_n891_ & ~new_n5120_;
  assign new_n5122_ = new_n895_ & ~new_n5121_;
  assign new_n5123_ = new_n899_ & ~new_n5122_;
  assign new_n5124_ = new_n903_ & ~new_n5123_;
  assign new_n5125_ = new_n907_ & ~new_n5124_;
  assign new_n5126_ = new_n911_ & ~new_n5125_;
  assign new_n5127_ = new_n915_ & ~new_n5126_;
  assign new_n5128_ = new_n919_ & ~new_n5127_;
  assign new_n5129_ = new_n923_ & ~new_n5128_;
  assign new_n5130_ = new_n927_ & ~new_n5129_;
  assign new_n5131_ = new_n931_ & ~new_n5130_;
  assign new_n5132_ = new_n935_ & ~new_n5131_;
  assign new_n5133_ = new_n939_ & ~new_n5132_;
  assign new_n5134_ = new_n943_ & ~new_n5133_;
  assign new_n5135_ = new_n947_ & ~new_n5134_;
  assign new_n5136_ = new_n951_ & ~new_n5135_;
  assign new_n5137_ = new_n955_ & ~new_n5136_;
  assign new_n5138_ = new_n959_ & ~new_n5137_;
  assign new_n5139_ = new_n963_ & ~new_n5138_;
  assign new_n5140_ = new_n967_ & ~new_n5139_;
  assign new_n5141_ = new_n971_ & ~new_n5140_;
  assign new_n5142_ = new_n975_ & ~new_n5141_;
  assign new_n5143_ = new_n979_ & ~new_n5142_;
  assign new_n5144_ = new_n983_ & ~new_n5143_;
  assign new_n5145_ = new_n987_ & ~new_n5144_;
  assign new_n5146_ = new_n991_ & ~new_n5145_;
  assign new_n5147_ = new_n995_ & ~new_n5146_;
  assign new_n5148_ = new_n999_ & ~new_n5147_;
  assign new_n5149_ = new_n1003_ & ~new_n5148_;
  assign new_n5150_ = new_n1007_ & ~new_n5149_;
  assign new_n5151_ = new_n1011_ & ~new_n5150_;
  assign new_n5152_ = new_n1015_ & ~new_n5151_;
  assign new_n5153_ = new_n1019_ & ~new_n5152_;
  assign new_n5154_ = new_n1023_ & ~new_n5153_;
  assign new_n5155_ = new_n1027_ & ~new_n5154_;
  assign new_n5156_ = new_n1031_ & ~new_n5155_;
  assign new_n5157_ = new_n1035_ & ~new_n5156_;
  assign new_n5158_ = new_n1039_ & ~new_n5157_;
  assign new_n5159_ = new_n1043_ & ~new_n5158_;
  assign new_n5160_ = new_n1047_ & ~new_n5159_;
  assign new_n5161_ = new_n1051_ & ~new_n5160_;
  assign new_n5162_ = new_n1055_ & ~new_n5161_;
  assign new_n5163_ = new_n1059_ & ~new_n5162_;
  assign new_n5164_ = new_n1574_ & ~new_n5163_;
  assign new_n5165_ = new_n1576_ & ~new_n5164_;
  assign new_n5166_ = new_n1837_ & ~new_n5165_;
  assign new_n5167_ = new_n1068_ & ~new_n5166_;
  assign new_n5168_ = new_n1072_ & ~new_n5167_;
  assign new_n5169_ = new_n1076_ & ~new_n5168_;
  assign new_n5170_ = new_n1080_ & ~new_n5169_;
  assign new_n5171_ = new_n1084_ & ~new_n5170_;
  assign new_n5172_ = new_n1088_ & ~new_n5171_;
  assign new_n5173_ = new_n1092_ & ~new_n5172_;
  assign new_n5174_ = new_n1096_ & ~new_n5173_;
  assign new_n5175_ = new_n1100_ & ~new_n5174_;
  assign new_n5176_ = new_n1104_ & ~new_n5175_;
  assign new_n5177_ = new_n1108_ & ~new_n5176_;
  assign new_n5178_ = new_n1112_ & ~new_n5177_;
  assign new_n5179_ = new_n1116_ & ~new_n5178_;
  assign new_n5180_ = new_n1120_ & ~new_n5179_;
  assign new_n5181_ = new_n1124_ & ~new_n5180_;
  assign new_n5182_ = new_n1128_ & ~new_n5181_;
  assign new_n5183_ = new_n1132_ & ~new_n5182_;
  assign new_n5184_ = new_n1136_ & ~new_n5183_;
  assign new_n5185_ = new_n1140_ & ~new_n5184_;
  assign new_n5186_ = new_n1144_ & ~new_n5185_;
  assign new_n5187_ = new_n1148_ & ~new_n5186_;
  assign new_n5188_ = new_n1152_ & ~new_n5187_;
  assign new_n5189_ = new_n1156_ & ~new_n5188_;
  assign new_n5190_ = new_n1160_ & ~new_n5189_;
  assign new_n5191_ = new_n1164_ & ~new_n5190_;
  assign new_n5192_ = new_n1168_ & ~new_n5191_;
  assign new_n5193_ = new_n1172_ & ~new_n5192_;
  assign new_n5194_ = \req[46]  & ~new_n1174_;
  assign \grant[46]  = ~new_n5193_ & new_n5194_;
  assign new_n5196_ = ~new_n511_ & new_n1183_;
  assign new_n5197_ = new_n1188_ & ~new_n5196_;
  assign new_n5198_ = new_n1192_ & ~new_n5197_;
  assign new_n5199_ = new_n1196_ & ~new_n5198_;
  assign new_n5200_ = new_n1200_ & ~new_n5199_;
  assign new_n5201_ = new_n1204_ & ~new_n5200_;
  assign new_n5202_ = new_n1208_ & ~new_n5201_;
  assign new_n5203_ = new_n1212_ & ~new_n5202_;
  assign new_n5204_ = new_n1216_ & ~new_n5203_;
  assign new_n5205_ = new_n1220_ & ~new_n5204_;
  assign new_n5206_ = new_n1224_ & ~new_n5205_;
  assign new_n5207_ = new_n1228_ & ~new_n5206_;
  assign new_n5208_ = new_n1232_ & ~new_n5207_;
  assign new_n5209_ = new_n1236_ & ~new_n5208_;
  assign new_n5210_ = new_n1240_ & ~new_n5209_;
  assign new_n5211_ = new_n1244_ & ~new_n5210_;
  assign new_n5212_ = new_n1248_ & ~new_n5211_;
  assign new_n5213_ = new_n1252_ & ~new_n5212_;
  assign new_n5214_ = new_n1256_ & ~new_n5213_;
  assign new_n5215_ = new_n1260_ & ~new_n5214_;
  assign new_n5216_ = new_n1264_ & ~new_n5215_;
  assign new_n5217_ = new_n1268_ & ~new_n5216_;
  assign new_n5218_ = new_n1272_ & ~new_n5217_;
  assign new_n5219_ = new_n1276_ & ~new_n5218_;
  assign new_n5220_ = new_n1280_ & ~new_n5219_;
  assign new_n5221_ = new_n1284_ & ~new_n5220_;
  assign new_n5222_ = new_n1288_ & ~new_n5221_;
  assign new_n5223_ = new_n1292_ & ~new_n5222_;
  assign new_n5224_ = new_n1296_ & ~new_n5223_;
  assign new_n5225_ = new_n1300_ & ~new_n5224_;
  assign new_n5226_ = new_n1304_ & ~new_n5225_;
  assign new_n5227_ = new_n1308_ & ~new_n5226_;
  assign new_n5228_ = new_n1312_ & ~new_n5227_;
  assign new_n5229_ = new_n1316_ & ~new_n5228_;
  assign new_n5230_ = new_n1320_ & ~new_n5229_;
  assign new_n5231_ = new_n1324_ & ~new_n5230_;
  assign new_n5232_ = new_n1328_ & ~new_n5231_;
  assign new_n5233_ = new_n1332_ & ~new_n5232_;
  assign new_n5234_ = new_n1336_ & ~new_n5233_;
  assign new_n5235_ = new_n1340_ & ~new_n5234_;
  assign new_n5236_ = new_n1344_ & ~new_n5235_;
  assign new_n5237_ = new_n1348_ & ~new_n5236_;
  assign new_n5238_ = new_n1352_ & ~new_n5237_;
  assign new_n5239_ = new_n1356_ & ~new_n5238_;
  assign new_n5240_ = new_n1360_ & ~new_n5239_;
  assign new_n5241_ = new_n1364_ & ~new_n5240_;
  assign new_n5242_ = new_n1368_ & ~new_n5241_;
  assign new_n5243_ = new_n1372_ & ~new_n5242_;
  assign new_n5244_ = new_n1376_ & ~new_n5243_;
  assign new_n5245_ = new_n1380_ & ~new_n5244_;
  assign new_n5246_ = new_n1384_ & ~new_n5245_;
  assign new_n5247_ = new_n1388_ & ~new_n5246_;
  assign new_n5248_ = new_n1392_ & ~new_n5247_;
  assign new_n5249_ = new_n1396_ & ~new_n5248_;
  assign new_n5250_ = new_n1663_ & ~new_n5249_;
  assign new_n5251_ = new_n392_ & ~new_n5250_;
  assign new_n5252_ = new_n396_ & ~new_n5251_;
  assign new_n5253_ = new_n400_ & ~new_n5252_;
  assign new_n5254_ = new_n404_ & ~new_n5253_;
  assign new_n5255_ = new_n408_ & ~new_n5254_;
  assign new_n5256_ = new_n412_ & ~new_n5255_;
  assign new_n5257_ = new_n416_ & ~new_n5256_;
  assign new_n5258_ = new_n420_ & ~new_n5257_;
  assign new_n5259_ = new_n424_ & ~new_n5258_;
  assign new_n5260_ = new_n428_ & ~new_n5259_;
  assign new_n5261_ = new_n432_ & ~new_n5260_;
  assign new_n5262_ = new_n436_ & ~new_n5261_;
  assign new_n5263_ = new_n440_ & ~new_n5262_;
  assign new_n5264_ = new_n444_ & ~new_n5263_;
  assign new_n5265_ = new_n448_ & ~new_n5264_;
  assign new_n5266_ = new_n452_ & ~new_n5265_;
  assign new_n5267_ = new_n456_ & ~new_n5266_;
  assign new_n5268_ = new_n460_ & ~new_n5267_;
  assign new_n5269_ = new_n464_ & ~new_n5268_;
  assign new_n5270_ = new_n468_ & ~new_n5269_;
  assign new_n5271_ = new_n472_ & ~new_n5270_;
  assign new_n5272_ = new_n476_ & ~new_n5271_;
  assign new_n5273_ = new_n480_ & ~new_n5272_;
  assign new_n5274_ = new_n484_ & ~new_n5273_;
  assign new_n5275_ = new_n488_ & ~new_n5274_;
  assign new_n5276_ = new_n492_ & ~new_n5275_;
  assign new_n5277_ = new_n496_ & ~new_n5276_;
  assign new_n5278_ = new_n500_ & ~new_n5277_;
  assign new_n5279_ = new_n504_ & ~new_n5278_;
  assign new_n5280_ = \req[47]  & ~new_n506_;
  assign \grant[47]  = ~new_n5279_ & new_n5280_;
  assign new_n5282_ = new_n515_ & ~new_n850_;
  assign new_n5283_ = new_n520_ & ~new_n5282_;
  assign new_n5284_ = new_n524_ & ~new_n5283_;
  assign new_n5285_ = new_n528_ & ~new_n5284_;
  assign new_n5286_ = new_n532_ & ~new_n5285_;
  assign new_n5287_ = new_n536_ & ~new_n5286_;
  assign new_n5288_ = new_n540_ & ~new_n5287_;
  assign new_n5289_ = new_n544_ & ~new_n5288_;
  assign new_n5290_ = new_n548_ & ~new_n5289_;
  assign new_n5291_ = new_n552_ & ~new_n5290_;
  assign new_n5292_ = new_n556_ & ~new_n5291_;
  assign new_n5293_ = new_n560_ & ~new_n5292_;
  assign new_n5294_ = new_n564_ & ~new_n5293_;
  assign new_n5295_ = new_n568_ & ~new_n5294_;
  assign new_n5296_ = new_n572_ & ~new_n5295_;
  assign new_n5297_ = new_n576_ & ~new_n5296_;
  assign new_n5298_ = new_n580_ & ~new_n5297_;
  assign new_n5299_ = new_n584_ & ~new_n5298_;
  assign new_n5300_ = new_n588_ & ~new_n5299_;
  assign new_n5301_ = new_n592_ & ~new_n5300_;
  assign new_n5302_ = new_n596_ & ~new_n5301_;
  assign new_n5303_ = new_n600_ & ~new_n5302_;
  assign new_n5304_ = new_n604_ & ~new_n5303_;
  assign new_n5305_ = new_n608_ & ~new_n5304_;
  assign new_n5306_ = new_n612_ & ~new_n5305_;
  assign new_n5307_ = new_n616_ & ~new_n5306_;
  assign new_n5308_ = new_n620_ & ~new_n5307_;
  assign new_n5309_ = new_n624_ & ~new_n5308_;
  assign new_n5310_ = new_n628_ & ~new_n5309_;
  assign new_n5311_ = new_n632_ & ~new_n5310_;
  assign new_n5312_ = new_n636_ & ~new_n5311_;
  assign new_n5313_ = new_n640_ & ~new_n5312_;
  assign new_n5314_ = new_n644_ & ~new_n5313_;
  assign new_n5315_ = new_n648_ & ~new_n5314_;
  assign new_n5316_ = new_n652_ & ~new_n5315_;
  assign new_n5317_ = new_n656_ & ~new_n5316_;
  assign new_n5318_ = new_n660_ & ~new_n5317_;
  assign new_n5319_ = new_n664_ & ~new_n5318_;
  assign new_n5320_ = new_n668_ & ~new_n5319_;
  assign new_n5321_ = new_n672_ & ~new_n5320_;
  assign new_n5322_ = new_n676_ & ~new_n5321_;
  assign new_n5323_ = new_n680_ & ~new_n5322_;
  assign new_n5324_ = new_n684_ & ~new_n5323_;
  assign new_n5325_ = new_n688_ & ~new_n5324_;
  assign new_n5326_ = new_n692_ & ~new_n5325_;
  assign new_n5327_ = new_n696_ & ~new_n5326_;
  assign new_n5328_ = new_n700_ & ~new_n5327_;
  assign new_n5329_ = new_n704_ & ~new_n5328_;
  assign new_n5330_ = new_n708_ & ~new_n5329_;
  assign new_n5331_ = new_n712_ & ~new_n5330_;
  assign new_n5332_ = new_n716_ & ~new_n5331_;
  assign new_n5333_ = new_n720_ & ~new_n5332_;
  assign new_n5334_ = new_n1484_ & ~new_n5333_;
  assign new_n5335_ = new_n1486_ & ~new_n5334_;
  assign new_n5336_ = new_n1750_ & ~new_n5335_;
  assign new_n5337_ = new_n731_ & ~new_n5336_;
  assign new_n5338_ = new_n735_ & ~new_n5337_;
  assign new_n5339_ = new_n739_ & ~new_n5338_;
  assign new_n5340_ = new_n743_ & ~new_n5339_;
  assign new_n5341_ = new_n747_ & ~new_n5340_;
  assign new_n5342_ = new_n751_ & ~new_n5341_;
  assign new_n5343_ = new_n755_ & ~new_n5342_;
  assign new_n5344_ = new_n759_ & ~new_n5343_;
  assign new_n5345_ = new_n763_ & ~new_n5344_;
  assign new_n5346_ = new_n767_ & ~new_n5345_;
  assign new_n5347_ = new_n771_ & ~new_n5346_;
  assign new_n5348_ = new_n775_ & ~new_n5347_;
  assign new_n5349_ = new_n779_ & ~new_n5348_;
  assign new_n5350_ = new_n783_ & ~new_n5349_;
  assign new_n5351_ = new_n787_ & ~new_n5350_;
  assign new_n5352_ = new_n791_ & ~new_n5351_;
  assign new_n5353_ = new_n795_ & ~new_n5352_;
  assign new_n5354_ = new_n799_ & ~new_n5353_;
  assign new_n5355_ = new_n803_ & ~new_n5354_;
  assign new_n5356_ = new_n807_ & ~new_n5355_;
  assign new_n5357_ = new_n811_ & ~new_n5356_;
  assign new_n5358_ = new_n815_ & ~new_n5357_;
  assign new_n5359_ = new_n819_ & ~new_n5358_;
  assign new_n5360_ = new_n823_ & ~new_n5359_;
  assign new_n5361_ = new_n827_ & ~new_n5360_;
  assign new_n5362_ = new_n831_ & ~new_n5361_;
  assign new_n5363_ = new_n835_ & ~new_n5362_;
  assign new_n5364_ = new_n839_ & ~new_n5363_;
  assign new_n5365_ = new_n843_ & ~new_n5364_;
  assign new_n5366_ = \req[48]  & ~new_n845_;
  assign \grant[48]  = ~new_n5365_ & new_n5366_;
  assign new_n5368_ = new_n854_ & ~new_n1187_;
  assign new_n5369_ = new_n859_ & ~new_n5368_;
  assign new_n5370_ = new_n863_ & ~new_n5369_;
  assign new_n5371_ = new_n867_ & ~new_n5370_;
  assign new_n5372_ = new_n871_ & ~new_n5371_;
  assign new_n5373_ = new_n875_ & ~new_n5372_;
  assign new_n5374_ = new_n879_ & ~new_n5373_;
  assign new_n5375_ = new_n883_ & ~new_n5374_;
  assign new_n5376_ = new_n887_ & ~new_n5375_;
  assign new_n5377_ = new_n891_ & ~new_n5376_;
  assign new_n5378_ = new_n895_ & ~new_n5377_;
  assign new_n5379_ = new_n899_ & ~new_n5378_;
  assign new_n5380_ = new_n903_ & ~new_n5379_;
  assign new_n5381_ = new_n907_ & ~new_n5380_;
  assign new_n5382_ = new_n911_ & ~new_n5381_;
  assign new_n5383_ = new_n915_ & ~new_n5382_;
  assign new_n5384_ = new_n919_ & ~new_n5383_;
  assign new_n5385_ = new_n923_ & ~new_n5384_;
  assign new_n5386_ = new_n927_ & ~new_n5385_;
  assign new_n5387_ = new_n931_ & ~new_n5386_;
  assign new_n5388_ = new_n935_ & ~new_n5387_;
  assign new_n5389_ = new_n939_ & ~new_n5388_;
  assign new_n5390_ = new_n943_ & ~new_n5389_;
  assign new_n5391_ = new_n947_ & ~new_n5390_;
  assign new_n5392_ = new_n951_ & ~new_n5391_;
  assign new_n5393_ = new_n955_ & ~new_n5392_;
  assign new_n5394_ = new_n959_ & ~new_n5393_;
  assign new_n5395_ = new_n963_ & ~new_n5394_;
  assign new_n5396_ = new_n967_ & ~new_n5395_;
  assign new_n5397_ = new_n971_ & ~new_n5396_;
  assign new_n5398_ = new_n975_ & ~new_n5397_;
  assign new_n5399_ = new_n979_ & ~new_n5398_;
  assign new_n5400_ = new_n983_ & ~new_n5399_;
  assign new_n5401_ = new_n987_ & ~new_n5400_;
  assign new_n5402_ = new_n991_ & ~new_n5401_;
  assign new_n5403_ = new_n995_ & ~new_n5402_;
  assign new_n5404_ = new_n999_ & ~new_n5403_;
  assign new_n5405_ = new_n1003_ & ~new_n5404_;
  assign new_n5406_ = new_n1007_ & ~new_n5405_;
  assign new_n5407_ = new_n1011_ & ~new_n5406_;
  assign new_n5408_ = new_n1015_ & ~new_n5407_;
  assign new_n5409_ = new_n1019_ & ~new_n5408_;
  assign new_n5410_ = new_n1023_ & ~new_n5409_;
  assign new_n5411_ = new_n1027_ & ~new_n5410_;
  assign new_n5412_ = new_n1031_ & ~new_n5411_;
  assign new_n5413_ = new_n1035_ & ~new_n5412_;
  assign new_n5414_ = new_n1039_ & ~new_n5413_;
  assign new_n5415_ = new_n1043_ & ~new_n5414_;
  assign new_n5416_ = new_n1047_ & ~new_n5415_;
  assign new_n5417_ = new_n1051_ & ~new_n5416_;
  assign new_n5418_ = new_n1055_ & ~new_n5417_;
  assign new_n5419_ = new_n1059_ & ~new_n5418_;
  assign new_n5420_ = new_n1574_ & ~new_n5419_;
  assign new_n5421_ = new_n1576_ & ~new_n5420_;
  assign new_n5422_ = new_n1837_ & ~new_n5421_;
  assign new_n5423_ = new_n1068_ & ~new_n5422_;
  assign new_n5424_ = new_n1072_ & ~new_n5423_;
  assign new_n5425_ = new_n1076_ & ~new_n5424_;
  assign new_n5426_ = new_n1080_ & ~new_n5425_;
  assign new_n5427_ = new_n1084_ & ~new_n5426_;
  assign new_n5428_ = new_n1088_ & ~new_n5427_;
  assign new_n5429_ = new_n1092_ & ~new_n5428_;
  assign new_n5430_ = new_n1096_ & ~new_n5429_;
  assign new_n5431_ = new_n1100_ & ~new_n5430_;
  assign new_n5432_ = new_n1104_ & ~new_n5431_;
  assign new_n5433_ = new_n1108_ & ~new_n5432_;
  assign new_n5434_ = new_n1112_ & ~new_n5433_;
  assign new_n5435_ = new_n1116_ & ~new_n5434_;
  assign new_n5436_ = new_n1120_ & ~new_n5435_;
  assign new_n5437_ = new_n1124_ & ~new_n5436_;
  assign new_n5438_ = new_n1128_ & ~new_n5437_;
  assign new_n5439_ = new_n1132_ & ~new_n5438_;
  assign new_n5440_ = new_n1136_ & ~new_n5439_;
  assign new_n5441_ = new_n1140_ & ~new_n5440_;
  assign new_n5442_ = new_n1144_ & ~new_n5441_;
  assign new_n5443_ = new_n1148_ & ~new_n5442_;
  assign new_n5444_ = new_n1152_ & ~new_n5443_;
  assign new_n5445_ = new_n1156_ & ~new_n5444_;
  assign new_n5446_ = new_n1160_ & ~new_n5445_;
  assign new_n5447_ = new_n1164_ & ~new_n5446_;
  assign new_n5448_ = new_n1168_ & ~new_n5447_;
  assign new_n5449_ = new_n1172_ & ~new_n5448_;
  assign new_n5450_ = new_n1176_ & ~new_n5449_;
  assign new_n5451_ = new_n1180_ & ~new_n5450_;
  assign new_n5452_ = \req[49]  & ~new_n1182_;
  assign \grant[49]  = ~new_n5451_ & new_n5452_;
  assign new_n5454_ = ~new_n519_ & new_n1191_;
  assign new_n5455_ = new_n1196_ & ~new_n5454_;
  assign new_n5456_ = new_n1200_ & ~new_n5455_;
  assign new_n5457_ = new_n1204_ & ~new_n5456_;
  assign new_n5458_ = new_n1208_ & ~new_n5457_;
  assign new_n5459_ = new_n1212_ & ~new_n5458_;
  assign new_n5460_ = new_n1216_ & ~new_n5459_;
  assign new_n5461_ = new_n1220_ & ~new_n5460_;
  assign new_n5462_ = new_n1224_ & ~new_n5461_;
  assign new_n5463_ = new_n1228_ & ~new_n5462_;
  assign new_n5464_ = new_n1232_ & ~new_n5463_;
  assign new_n5465_ = new_n1236_ & ~new_n5464_;
  assign new_n5466_ = new_n1240_ & ~new_n5465_;
  assign new_n5467_ = new_n1244_ & ~new_n5466_;
  assign new_n5468_ = new_n1248_ & ~new_n5467_;
  assign new_n5469_ = new_n1252_ & ~new_n5468_;
  assign new_n5470_ = new_n1256_ & ~new_n5469_;
  assign new_n5471_ = new_n1260_ & ~new_n5470_;
  assign new_n5472_ = new_n1264_ & ~new_n5471_;
  assign new_n5473_ = new_n1268_ & ~new_n5472_;
  assign new_n5474_ = new_n1272_ & ~new_n5473_;
  assign new_n5475_ = new_n1276_ & ~new_n5474_;
  assign new_n5476_ = new_n1280_ & ~new_n5475_;
  assign new_n5477_ = new_n1284_ & ~new_n5476_;
  assign new_n5478_ = new_n1288_ & ~new_n5477_;
  assign new_n5479_ = new_n1292_ & ~new_n5478_;
  assign new_n5480_ = new_n1296_ & ~new_n5479_;
  assign new_n5481_ = new_n1300_ & ~new_n5480_;
  assign new_n5482_ = new_n1304_ & ~new_n5481_;
  assign new_n5483_ = new_n1308_ & ~new_n5482_;
  assign new_n5484_ = new_n1312_ & ~new_n5483_;
  assign new_n5485_ = new_n1316_ & ~new_n5484_;
  assign new_n5486_ = new_n1320_ & ~new_n5485_;
  assign new_n5487_ = new_n1324_ & ~new_n5486_;
  assign new_n5488_ = new_n1328_ & ~new_n5487_;
  assign new_n5489_ = new_n1332_ & ~new_n5488_;
  assign new_n5490_ = new_n1336_ & ~new_n5489_;
  assign new_n5491_ = new_n1340_ & ~new_n5490_;
  assign new_n5492_ = new_n1344_ & ~new_n5491_;
  assign new_n5493_ = new_n1348_ & ~new_n5492_;
  assign new_n5494_ = new_n1352_ & ~new_n5493_;
  assign new_n5495_ = new_n1356_ & ~new_n5494_;
  assign new_n5496_ = new_n1360_ & ~new_n5495_;
  assign new_n5497_ = new_n1364_ & ~new_n5496_;
  assign new_n5498_ = new_n1368_ & ~new_n5497_;
  assign new_n5499_ = new_n1372_ & ~new_n5498_;
  assign new_n5500_ = new_n1376_ & ~new_n5499_;
  assign new_n5501_ = new_n1380_ & ~new_n5500_;
  assign new_n5502_ = new_n1384_ & ~new_n5501_;
  assign new_n5503_ = new_n1388_ & ~new_n5502_;
  assign new_n5504_ = new_n1392_ & ~new_n5503_;
  assign new_n5505_ = new_n1396_ & ~new_n5504_;
  assign new_n5506_ = new_n1663_ & ~new_n5505_;
  assign new_n5507_ = new_n392_ & ~new_n5506_;
  assign new_n5508_ = new_n396_ & ~new_n5507_;
  assign new_n5509_ = new_n400_ & ~new_n5508_;
  assign new_n5510_ = new_n404_ & ~new_n5509_;
  assign new_n5511_ = new_n408_ & ~new_n5510_;
  assign new_n5512_ = new_n412_ & ~new_n5511_;
  assign new_n5513_ = new_n416_ & ~new_n5512_;
  assign new_n5514_ = new_n420_ & ~new_n5513_;
  assign new_n5515_ = new_n424_ & ~new_n5514_;
  assign new_n5516_ = new_n428_ & ~new_n5515_;
  assign new_n5517_ = new_n432_ & ~new_n5516_;
  assign new_n5518_ = new_n436_ & ~new_n5517_;
  assign new_n5519_ = new_n440_ & ~new_n5518_;
  assign new_n5520_ = new_n444_ & ~new_n5519_;
  assign new_n5521_ = new_n448_ & ~new_n5520_;
  assign new_n5522_ = new_n452_ & ~new_n5521_;
  assign new_n5523_ = new_n456_ & ~new_n5522_;
  assign new_n5524_ = new_n460_ & ~new_n5523_;
  assign new_n5525_ = new_n464_ & ~new_n5524_;
  assign new_n5526_ = new_n468_ & ~new_n5525_;
  assign new_n5527_ = new_n472_ & ~new_n5526_;
  assign new_n5528_ = new_n476_ & ~new_n5527_;
  assign new_n5529_ = new_n480_ & ~new_n5528_;
  assign new_n5530_ = new_n484_ & ~new_n5529_;
  assign new_n5531_ = new_n488_ & ~new_n5530_;
  assign new_n5532_ = new_n492_ & ~new_n5531_;
  assign new_n5533_ = new_n496_ & ~new_n5532_;
  assign new_n5534_ = new_n500_ & ~new_n5533_;
  assign new_n5535_ = new_n504_ & ~new_n5534_;
  assign new_n5536_ = new_n508_ & ~new_n5535_;
  assign new_n5537_ = new_n512_ & ~new_n5536_;
  assign new_n5538_ = \req[50]  & ~new_n514_;
  assign \grant[50]  = ~new_n5537_ & new_n5538_;
  assign new_n5540_ = new_n523_ & ~new_n858_;
  assign new_n5541_ = new_n528_ & ~new_n5540_;
  assign new_n5542_ = new_n532_ & ~new_n5541_;
  assign new_n5543_ = new_n536_ & ~new_n5542_;
  assign new_n5544_ = new_n540_ & ~new_n5543_;
  assign new_n5545_ = new_n544_ & ~new_n5544_;
  assign new_n5546_ = new_n548_ & ~new_n5545_;
  assign new_n5547_ = new_n552_ & ~new_n5546_;
  assign new_n5548_ = new_n556_ & ~new_n5547_;
  assign new_n5549_ = new_n560_ & ~new_n5548_;
  assign new_n5550_ = new_n564_ & ~new_n5549_;
  assign new_n5551_ = new_n568_ & ~new_n5550_;
  assign new_n5552_ = new_n572_ & ~new_n5551_;
  assign new_n5553_ = new_n576_ & ~new_n5552_;
  assign new_n5554_ = new_n580_ & ~new_n5553_;
  assign new_n5555_ = new_n584_ & ~new_n5554_;
  assign new_n5556_ = new_n588_ & ~new_n5555_;
  assign new_n5557_ = new_n592_ & ~new_n5556_;
  assign new_n5558_ = new_n596_ & ~new_n5557_;
  assign new_n5559_ = new_n600_ & ~new_n5558_;
  assign new_n5560_ = new_n604_ & ~new_n5559_;
  assign new_n5561_ = new_n608_ & ~new_n5560_;
  assign new_n5562_ = new_n612_ & ~new_n5561_;
  assign new_n5563_ = new_n616_ & ~new_n5562_;
  assign new_n5564_ = new_n620_ & ~new_n5563_;
  assign new_n5565_ = new_n624_ & ~new_n5564_;
  assign new_n5566_ = new_n628_ & ~new_n5565_;
  assign new_n5567_ = new_n632_ & ~new_n5566_;
  assign new_n5568_ = new_n636_ & ~new_n5567_;
  assign new_n5569_ = new_n640_ & ~new_n5568_;
  assign new_n5570_ = new_n644_ & ~new_n5569_;
  assign new_n5571_ = new_n648_ & ~new_n5570_;
  assign new_n5572_ = new_n652_ & ~new_n5571_;
  assign new_n5573_ = new_n656_ & ~new_n5572_;
  assign new_n5574_ = new_n660_ & ~new_n5573_;
  assign new_n5575_ = new_n664_ & ~new_n5574_;
  assign new_n5576_ = new_n668_ & ~new_n5575_;
  assign new_n5577_ = new_n672_ & ~new_n5576_;
  assign new_n5578_ = new_n676_ & ~new_n5577_;
  assign new_n5579_ = new_n680_ & ~new_n5578_;
  assign new_n5580_ = new_n684_ & ~new_n5579_;
  assign new_n5581_ = new_n688_ & ~new_n5580_;
  assign new_n5582_ = new_n692_ & ~new_n5581_;
  assign new_n5583_ = new_n696_ & ~new_n5582_;
  assign new_n5584_ = new_n700_ & ~new_n5583_;
  assign new_n5585_ = new_n704_ & ~new_n5584_;
  assign new_n5586_ = new_n708_ & ~new_n5585_;
  assign new_n5587_ = new_n712_ & ~new_n5586_;
  assign new_n5588_ = new_n716_ & ~new_n5587_;
  assign new_n5589_ = new_n720_ & ~new_n5588_;
  assign new_n5590_ = new_n1484_ & ~new_n5589_;
  assign new_n5591_ = new_n1486_ & ~new_n5590_;
  assign new_n5592_ = new_n1750_ & ~new_n5591_;
  assign new_n5593_ = new_n731_ & ~new_n5592_;
  assign new_n5594_ = new_n735_ & ~new_n5593_;
  assign new_n5595_ = new_n739_ & ~new_n5594_;
  assign new_n5596_ = new_n743_ & ~new_n5595_;
  assign new_n5597_ = new_n747_ & ~new_n5596_;
  assign new_n5598_ = new_n751_ & ~new_n5597_;
  assign new_n5599_ = new_n755_ & ~new_n5598_;
  assign new_n5600_ = new_n759_ & ~new_n5599_;
  assign new_n5601_ = new_n763_ & ~new_n5600_;
  assign new_n5602_ = new_n767_ & ~new_n5601_;
  assign new_n5603_ = new_n771_ & ~new_n5602_;
  assign new_n5604_ = new_n775_ & ~new_n5603_;
  assign new_n5605_ = new_n779_ & ~new_n5604_;
  assign new_n5606_ = new_n783_ & ~new_n5605_;
  assign new_n5607_ = new_n787_ & ~new_n5606_;
  assign new_n5608_ = new_n791_ & ~new_n5607_;
  assign new_n5609_ = new_n795_ & ~new_n5608_;
  assign new_n5610_ = new_n799_ & ~new_n5609_;
  assign new_n5611_ = new_n803_ & ~new_n5610_;
  assign new_n5612_ = new_n807_ & ~new_n5611_;
  assign new_n5613_ = new_n811_ & ~new_n5612_;
  assign new_n5614_ = new_n815_ & ~new_n5613_;
  assign new_n5615_ = new_n819_ & ~new_n5614_;
  assign new_n5616_ = new_n823_ & ~new_n5615_;
  assign new_n5617_ = new_n827_ & ~new_n5616_;
  assign new_n5618_ = new_n831_ & ~new_n5617_;
  assign new_n5619_ = new_n835_ & ~new_n5618_;
  assign new_n5620_ = new_n839_ & ~new_n5619_;
  assign new_n5621_ = new_n843_ & ~new_n5620_;
  assign new_n5622_ = new_n847_ & ~new_n5621_;
  assign new_n5623_ = new_n851_ & ~new_n5622_;
  assign new_n5624_ = \req[51]  & ~new_n853_;
  assign \grant[51]  = ~new_n5623_ & new_n5624_;
  assign new_n5626_ = new_n862_ & ~new_n1195_;
  assign new_n5627_ = new_n867_ & ~new_n5626_;
  assign new_n5628_ = new_n871_ & ~new_n5627_;
  assign new_n5629_ = new_n875_ & ~new_n5628_;
  assign new_n5630_ = new_n879_ & ~new_n5629_;
  assign new_n5631_ = new_n883_ & ~new_n5630_;
  assign new_n5632_ = new_n887_ & ~new_n5631_;
  assign new_n5633_ = new_n891_ & ~new_n5632_;
  assign new_n5634_ = new_n895_ & ~new_n5633_;
  assign new_n5635_ = new_n899_ & ~new_n5634_;
  assign new_n5636_ = new_n903_ & ~new_n5635_;
  assign new_n5637_ = new_n907_ & ~new_n5636_;
  assign new_n5638_ = new_n911_ & ~new_n5637_;
  assign new_n5639_ = new_n915_ & ~new_n5638_;
  assign new_n5640_ = new_n919_ & ~new_n5639_;
  assign new_n5641_ = new_n923_ & ~new_n5640_;
  assign new_n5642_ = new_n927_ & ~new_n5641_;
  assign new_n5643_ = new_n931_ & ~new_n5642_;
  assign new_n5644_ = new_n935_ & ~new_n5643_;
  assign new_n5645_ = new_n939_ & ~new_n5644_;
  assign new_n5646_ = new_n943_ & ~new_n5645_;
  assign new_n5647_ = new_n947_ & ~new_n5646_;
  assign new_n5648_ = new_n951_ & ~new_n5647_;
  assign new_n5649_ = new_n955_ & ~new_n5648_;
  assign new_n5650_ = new_n959_ & ~new_n5649_;
  assign new_n5651_ = new_n963_ & ~new_n5650_;
  assign new_n5652_ = new_n967_ & ~new_n5651_;
  assign new_n5653_ = new_n971_ & ~new_n5652_;
  assign new_n5654_ = new_n975_ & ~new_n5653_;
  assign new_n5655_ = new_n979_ & ~new_n5654_;
  assign new_n5656_ = new_n983_ & ~new_n5655_;
  assign new_n5657_ = new_n987_ & ~new_n5656_;
  assign new_n5658_ = new_n991_ & ~new_n5657_;
  assign new_n5659_ = new_n995_ & ~new_n5658_;
  assign new_n5660_ = new_n999_ & ~new_n5659_;
  assign new_n5661_ = new_n1003_ & ~new_n5660_;
  assign new_n5662_ = new_n1007_ & ~new_n5661_;
  assign new_n5663_ = new_n1011_ & ~new_n5662_;
  assign new_n5664_ = new_n1015_ & ~new_n5663_;
  assign new_n5665_ = new_n1019_ & ~new_n5664_;
  assign new_n5666_ = new_n1023_ & ~new_n5665_;
  assign new_n5667_ = new_n1027_ & ~new_n5666_;
  assign new_n5668_ = new_n1031_ & ~new_n5667_;
  assign new_n5669_ = new_n1035_ & ~new_n5668_;
  assign new_n5670_ = new_n1039_ & ~new_n5669_;
  assign new_n5671_ = new_n1043_ & ~new_n5670_;
  assign new_n5672_ = new_n1047_ & ~new_n5671_;
  assign new_n5673_ = new_n1051_ & ~new_n5672_;
  assign new_n5674_ = new_n1055_ & ~new_n5673_;
  assign new_n5675_ = new_n1059_ & ~new_n5674_;
  assign new_n5676_ = new_n1574_ & ~new_n5675_;
  assign new_n5677_ = new_n1576_ & ~new_n5676_;
  assign new_n5678_ = new_n1837_ & ~new_n5677_;
  assign new_n5679_ = new_n1068_ & ~new_n5678_;
  assign new_n5680_ = new_n1072_ & ~new_n5679_;
  assign new_n5681_ = new_n1076_ & ~new_n5680_;
  assign new_n5682_ = new_n1080_ & ~new_n5681_;
  assign new_n5683_ = new_n1084_ & ~new_n5682_;
  assign new_n5684_ = new_n1088_ & ~new_n5683_;
  assign new_n5685_ = new_n1092_ & ~new_n5684_;
  assign new_n5686_ = new_n1096_ & ~new_n5685_;
  assign new_n5687_ = new_n1100_ & ~new_n5686_;
  assign new_n5688_ = new_n1104_ & ~new_n5687_;
  assign new_n5689_ = new_n1108_ & ~new_n5688_;
  assign new_n5690_ = new_n1112_ & ~new_n5689_;
  assign new_n5691_ = new_n1116_ & ~new_n5690_;
  assign new_n5692_ = new_n1120_ & ~new_n5691_;
  assign new_n5693_ = new_n1124_ & ~new_n5692_;
  assign new_n5694_ = new_n1128_ & ~new_n5693_;
  assign new_n5695_ = new_n1132_ & ~new_n5694_;
  assign new_n5696_ = new_n1136_ & ~new_n5695_;
  assign new_n5697_ = new_n1140_ & ~new_n5696_;
  assign new_n5698_ = new_n1144_ & ~new_n5697_;
  assign new_n5699_ = new_n1148_ & ~new_n5698_;
  assign new_n5700_ = new_n1152_ & ~new_n5699_;
  assign new_n5701_ = new_n1156_ & ~new_n5700_;
  assign new_n5702_ = new_n1160_ & ~new_n5701_;
  assign new_n5703_ = new_n1164_ & ~new_n5702_;
  assign new_n5704_ = new_n1168_ & ~new_n5703_;
  assign new_n5705_ = new_n1172_ & ~new_n5704_;
  assign new_n5706_ = new_n1176_ & ~new_n5705_;
  assign new_n5707_ = new_n1180_ & ~new_n5706_;
  assign new_n5708_ = new_n1184_ & ~new_n5707_;
  assign new_n5709_ = new_n1188_ & ~new_n5708_;
  assign new_n5710_ = \req[52]  & ~new_n1190_;
  assign \grant[52]  = ~new_n5709_ & new_n5710_;
  assign new_n5712_ = ~new_n527_ & new_n1199_;
  assign new_n5713_ = new_n1204_ & ~new_n5712_;
  assign new_n5714_ = new_n1208_ & ~new_n5713_;
  assign new_n5715_ = new_n1212_ & ~new_n5714_;
  assign new_n5716_ = new_n1216_ & ~new_n5715_;
  assign new_n5717_ = new_n1220_ & ~new_n5716_;
  assign new_n5718_ = new_n1224_ & ~new_n5717_;
  assign new_n5719_ = new_n1228_ & ~new_n5718_;
  assign new_n5720_ = new_n1232_ & ~new_n5719_;
  assign new_n5721_ = new_n1236_ & ~new_n5720_;
  assign new_n5722_ = new_n1240_ & ~new_n5721_;
  assign new_n5723_ = new_n1244_ & ~new_n5722_;
  assign new_n5724_ = new_n1248_ & ~new_n5723_;
  assign new_n5725_ = new_n1252_ & ~new_n5724_;
  assign new_n5726_ = new_n1256_ & ~new_n5725_;
  assign new_n5727_ = new_n1260_ & ~new_n5726_;
  assign new_n5728_ = new_n1264_ & ~new_n5727_;
  assign new_n5729_ = new_n1268_ & ~new_n5728_;
  assign new_n5730_ = new_n1272_ & ~new_n5729_;
  assign new_n5731_ = new_n1276_ & ~new_n5730_;
  assign new_n5732_ = new_n1280_ & ~new_n5731_;
  assign new_n5733_ = new_n1284_ & ~new_n5732_;
  assign new_n5734_ = new_n1288_ & ~new_n5733_;
  assign new_n5735_ = new_n1292_ & ~new_n5734_;
  assign new_n5736_ = new_n1296_ & ~new_n5735_;
  assign new_n5737_ = new_n1300_ & ~new_n5736_;
  assign new_n5738_ = new_n1304_ & ~new_n5737_;
  assign new_n5739_ = new_n1308_ & ~new_n5738_;
  assign new_n5740_ = new_n1312_ & ~new_n5739_;
  assign new_n5741_ = new_n1316_ & ~new_n5740_;
  assign new_n5742_ = new_n1320_ & ~new_n5741_;
  assign new_n5743_ = new_n1324_ & ~new_n5742_;
  assign new_n5744_ = new_n1328_ & ~new_n5743_;
  assign new_n5745_ = new_n1332_ & ~new_n5744_;
  assign new_n5746_ = new_n1336_ & ~new_n5745_;
  assign new_n5747_ = new_n1340_ & ~new_n5746_;
  assign new_n5748_ = new_n1344_ & ~new_n5747_;
  assign new_n5749_ = new_n1348_ & ~new_n5748_;
  assign new_n5750_ = new_n1352_ & ~new_n5749_;
  assign new_n5751_ = new_n1356_ & ~new_n5750_;
  assign new_n5752_ = new_n1360_ & ~new_n5751_;
  assign new_n5753_ = new_n1364_ & ~new_n5752_;
  assign new_n5754_ = new_n1368_ & ~new_n5753_;
  assign new_n5755_ = new_n1372_ & ~new_n5754_;
  assign new_n5756_ = new_n1376_ & ~new_n5755_;
  assign new_n5757_ = new_n1380_ & ~new_n5756_;
  assign new_n5758_ = new_n1384_ & ~new_n5757_;
  assign new_n5759_ = new_n1388_ & ~new_n5758_;
  assign new_n5760_ = new_n1392_ & ~new_n5759_;
  assign new_n5761_ = new_n1396_ & ~new_n5760_;
  assign new_n5762_ = new_n1663_ & ~new_n5761_;
  assign new_n5763_ = new_n392_ & ~new_n5762_;
  assign new_n5764_ = new_n396_ & ~new_n5763_;
  assign new_n5765_ = new_n400_ & ~new_n5764_;
  assign new_n5766_ = new_n404_ & ~new_n5765_;
  assign new_n5767_ = new_n408_ & ~new_n5766_;
  assign new_n5768_ = new_n412_ & ~new_n5767_;
  assign new_n5769_ = new_n416_ & ~new_n5768_;
  assign new_n5770_ = new_n420_ & ~new_n5769_;
  assign new_n5771_ = new_n424_ & ~new_n5770_;
  assign new_n5772_ = new_n428_ & ~new_n5771_;
  assign new_n5773_ = new_n432_ & ~new_n5772_;
  assign new_n5774_ = new_n436_ & ~new_n5773_;
  assign new_n5775_ = new_n440_ & ~new_n5774_;
  assign new_n5776_ = new_n444_ & ~new_n5775_;
  assign new_n5777_ = new_n448_ & ~new_n5776_;
  assign new_n5778_ = new_n452_ & ~new_n5777_;
  assign new_n5779_ = new_n456_ & ~new_n5778_;
  assign new_n5780_ = new_n460_ & ~new_n5779_;
  assign new_n5781_ = new_n464_ & ~new_n5780_;
  assign new_n5782_ = new_n468_ & ~new_n5781_;
  assign new_n5783_ = new_n472_ & ~new_n5782_;
  assign new_n5784_ = new_n476_ & ~new_n5783_;
  assign new_n5785_ = new_n480_ & ~new_n5784_;
  assign new_n5786_ = new_n484_ & ~new_n5785_;
  assign new_n5787_ = new_n488_ & ~new_n5786_;
  assign new_n5788_ = new_n492_ & ~new_n5787_;
  assign new_n5789_ = new_n496_ & ~new_n5788_;
  assign new_n5790_ = new_n500_ & ~new_n5789_;
  assign new_n5791_ = new_n504_ & ~new_n5790_;
  assign new_n5792_ = new_n508_ & ~new_n5791_;
  assign new_n5793_ = new_n512_ & ~new_n5792_;
  assign new_n5794_ = new_n516_ & ~new_n5793_;
  assign new_n5795_ = new_n520_ & ~new_n5794_;
  assign new_n5796_ = \req[53]  & ~new_n522_;
  assign \grant[53]  = ~new_n5795_ & new_n5796_;
  assign new_n5798_ = new_n531_ & ~new_n866_;
  assign new_n5799_ = new_n536_ & ~new_n5798_;
  assign new_n5800_ = new_n540_ & ~new_n5799_;
  assign new_n5801_ = new_n544_ & ~new_n5800_;
  assign new_n5802_ = new_n548_ & ~new_n5801_;
  assign new_n5803_ = new_n552_ & ~new_n5802_;
  assign new_n5804_ = new_n556_ & ~new_n5803_;
  assign new_n5805_ = new_n560_ & ~new_n5804_;
  assign new_n5806_ = new_n564_ & ~new_n5805_;
  assign new_n5807_ = new_n568_ & ~new_n5806_;
  assign new_n5808_ = new_n572_ & ~new_n5807_;
  assign new_n5809_ = new_n576_ & ~new_n5808_;
  assign new_n5810_ = new_n580_ & ~new_n5809_;
  assign new_n5811_ = new_n584_ & ~new_n5810_;
  assign new_n5812_ = new_n588_ & ~new_n5811_;
  assign new_n5813_ = new_n592_ & ~new_n5812_;
  assign new_n5814_ = new_n596_ & ~new_n5813_;
  assign new_n5815_ = new_n600_ & ~new_n5814_;
  assign new_n5816_ = new_n604_ & ~new_n5815_;
  assign new_n5817_ = new_n608_ & ~new_n5816_;
  assign new_n5818_ = new_n612_ & ~new_n5817_;
  assign new_n5819_ = new_n616_ & ~new_n5818_;
  assign new_n5820_ = new_n620_ & ~new_n5819_;
  assign new_n5821_ = new_n624_ & ~new_n5820_;
  assign new_n5822_ = new_n628_ & ~new_n5821_;
  assign new_n5823_ = new_n632_ & ~new_n5822_;
  assign new_n5824_ = new_n636_ & ~new_n5823_;
  assign new_n5825_ = new_n640_ & ~new_n5824_;
  assign new_n5826_ = new_n644_ & ~new_n5825_;
  assign new_n5827_ = new_n648_ & ~new_n5826_;
  assign new_n5828_ = new_n652_ & ~new_n5827_;
  assign new_n5829_ = new_n656_ & ~new_n5828_;
  assign new_n5830_ = new_n660_ & ~new_n5829_;
  assign new_n5831_ = new_n664_ & ~new_n5830_;
  assign new_n5832_ = new_n668_ & ~new_n5831_;
  assign new_n5833_ = new_n672_ & ~new_n5832_;
  assign new_n5834_ = new_n676_ & ~new_n5833_;
  assign new_n5835_ = new_n680_ & ~new_n5834_;
  assign new_n5836_ = new_n684_ & ~new_n5835_;
  assign new_n5837_ = new_n688_ & ~new_n5836_;
  assign new_n5838_ = new_n692_ & ~new_n5837_;
  assign new_n5839_ = new_n696_ & ~new_n5838_;
  assign new_n5840_ = new_n700_ & ~new_n5839_;
  assign new_n5841_ = new_n704_ & ~new_n5840_;
  assign new_n5842_ = new_n708_ & ~new_n5841_;
  assign new_n5843_ = new_n712_ & ~new_n5842_;
  assign new_n5844_ = new_n716_ & ~new_n5843_;
  assign new_n5845_ = new_n720_ & ~new_n5844_;
  assign new_n5846_ = new_n1484_ & ~new_n5845_;
  assign new_n5847_ = new_n1486_ & ~new_n5846_;
  assign new_n5848_ = new_n1750_ & ~new_n5847_;
  assign new_n5849_ = new_n731_ & ~new_n5848_;
  assign new_n5850_ = new_n735_ & ~new_n5849_;
  assign new_n5851_ = new_n739_ & ~new_n5850_;
  assign new_n5852_ = new_n743_ & ~new_n5851_;
  assign new_n5853_ = new_n747_ & ~new_n5852_;
  assign new_n5854_ = new_n751_ & ~new_n5853_;
  assign new_n5855_ = new_n755_ & ~new_n5854_;
  assign new_n5856_ = new_n759_ & ~new_n5855_;
  assign new_n5857_ = new_n763_ & ~new_n5856_;
  assign new_n5858_ = new_n767_ & ~new_n5857_;
  assign new_n5859_ = new_n771_ & ~new_n5858_;
  assign new_n5860_ = new_n775_ & ~new_n5859_;
  assign new_n5861_ = new_n779_ & ~new_n5860_;
  assign new_n5862_ = new_n783_ & ~new_n5861_;
  assign new_n5863_ = new_n787_ & ~new_n5862_;
  assign new_n5864_ = new_n791_ & ~new_n5863_;
  assign new_n5865_ = new_n795_ & ~new_n5864_;
  assign new_n5866_ = new_n799_ & ~new_n5865_;
  assign new_n5867_ = new_n803_ & ~new_n5866_;
  assign new_n5868_ = new_n807_ & ~new_n5867_;
  assign new_n5869_ = new_n811_ & ~new_n5868_;
  assign new_n5870_ = new_n815_ & ~new_n5869_;
  assign new_n5871_ = new_n819_ & ~new_n5870_;
  assign new_n5872_ = new_n823_ & ~new_n5871_;
  assign new_n5873_ = new_n827_ & ~new_n5872_;
  assign new_n5874_ = new_n831_ & ~new_n5873_;
  assign new_n5875_ = new_n835_ & ~new_n5874_;
  assign new_n5876_ = new_n839_ & ~new_n5875_;
  assign new_n5877_ = new_n843_ & ~new_n5876_;
  assign new_n5878_ = new_n847_ & ~new_n5877_;
  assign new_n5879_ = new_n851_ & ~new_n5878_;
  assign new_n5880_ = new_n855_ & ~new_n5879_;
  assign new_n5881_ = new_n859_ & ~new_n5880_;
  assign new_n5882_ = \req[54]  & ~new_n861_;
  assign \grant[54]  = ~new_n5881_ & new_n5882_;
  assign new_n5884_ = new_n870_ & ~new_n1203_;
  assign new_n5885_ = new_n875_ & ~new_n5884_;
  assign new_n5886_ = new_n879_ & ~new_n5885_;
  assign new_n5887_ = new_n883_ & ~new_n5886_;
  assign new_n5888_ = new_n887_ & ~new_n5887_;
  assign new_n5889_ = new_n891_ & ~new_n5888_;
  assign new_n5890_ = new_n895_ & ~new_n5889_;
  assign new_n5891_ = new_n899_ & ~new_n5890_;
  assign new_n5892_ = new_n903_ & ~new_n5891_;
  assign new_n5893_ = new_n907_ & ~new_n5892_;
  assign new_n5894_ = new_n911_ & ~new_n5893_;
  assign new_n5895_ = new_n915_ & ~new_n5894_;
  assign new_n5896_ = new_n919_ & ~new_n5895_;
  assign new_n5897_ = new_n923_ & ~new_n5896_;
  assign new_n5898_ = new_n927_ & ~new_n5897_;
  assign new_n5899_ = new_n931_ & ~new_n5898_;
  assign new_n5900_ = new_n935_ & ~new_n5899_;
  assign new_n5901_ = new_n939_ & ~new_n5900_;
  assign new_n5902_ = new_n943_ & ~new_n5901_;
  assign new_n5903_ = new_n947_ & ~new_n5902_;
  assign new_n5904_ = new_n951_ & ~new_n5903_;
  assign new_n5905_ = new_n955_ & ~new_n5904_;
  assign new_n5906_ = new_n959_ & ~new_n5905_;
  assign new_n5907_ = new_n963_ & ~new_n5906_;
  assign new_n5908_ = new_n967_ & ~new_n5907_;
  assign new_n5909_ = new_n971_ & ~new_n5908_;
  assign new_n5910_ = new_n975_ & ~new_n5909_;
  assign new_n5911_ = new_n979_ & ~new_n5910_;
  assign new_n5912_ = new_n983_ & ~new_n5911_;
  assign new_n5913_ = new_n987_ & ~new_n5912_;
  assign new_n5914_ = new_n991_ & ~new_n5913_;
  assign new_n5915_ = new_n995_ & ~new_n5914_;
  assign new_n5916_ = new_n999_ & ~new_n5915_;
  assign new_n5917_ = new_n1003_ & ~new_n5916_;
  assign new_n5918_ = new_n1007_ & ~new_n5917_;
  assign new_n5919_ = new_n1011_ & ~new_n5918_;
  assign new_n5920_ = new_n1015_ & ~new_n5919_;
  assign new_n5921_ = new_n1019_ & ~new_n5920_;
  assign new_n5922_ = new_n1023_ & ~new_n5921_;
  assign new_n5923_ = new_n1027_ & ~new_n5922_;
  assign new_n5924_ = new_n1031_ & ~new_n5923_;
  assign new_n5925_ = new_n1035_ & ~new_n5924_;
  assign new_n5926_ = new_n1039_ & ~new_n5925_;
  assign new_n5927_ = new_n1043_ & ~new_n5926_;
  assign new_n5928_ = new_n1047_ & ~new_n5927_;
  assign new_n5929_ = new_n1051_ & ~new_n5928_;
  assign new_n5930_ = new_n1055_ & ~new_n5929_;
  assign new_n5931_ = new_n1059_ & ~new_n5930_;
  assign new_n5932_ = new_n1574_ & ~new_n5931_;
  assign new_n5933_ = new_n1576_ & ~new_n5932_;
  assign new_n5934_ = new_n1837_ & ~new_n5933_;
  assign new_n5935_ = new_n1068_ & ~new_n5934_;
  assign new_n5936_ = new_n1072_ & ~new_n5935_;
  assign new_n5937_ = new_n1076_ & ~new_n5936_;
  assign new_n5938_ = new_n1080_ & ~new_n5937_;
  assign new_n5939_ = new_n1084_ & ~new_n5938_;
  assign new_n5940_ = new_n1088_ & ~new_n5939_;
  assign new_n5941_ = new_n1092_ & ~new_n5940_;
  assign new_n5942_ = new_n1096_ & ~new_n5941_;
  assign new_n5943_ = new_n1100_ & ~new_n5942_;
  assign new_n5944_ = new_n1104_ & ~new_n5943_;
  assign new_n5945_ = new_n1108_ & ~new_n5944_;
  assign new_n5946_ = new_n1112_ & ~new_n5945_;
  assign new_n5947_ = new_n1116_ & ~new_n5946_;
  assign new_n5948_ = new_n1120_ & ~new_n5947_;
  assign new_n5949_ = new_n1124_ & ~new_n5948_;
  assign new_n5950_ = new_n1128_ & ~new_n5949_;
  assign new_n5951_ = new_n1132_ & ~new_n5950_;
  assign new_n5952_ = new_n1136_ & ~new_n5951_;
  assign new_n5953_ = new_n1140_ & ~new_n5952_;
  assign new_n5954_ = new_n1144_ & ~new_n5953_;
  assign new_n5955_ = new_n1148_ & ~new_n5954_;
  assign new_n5956_ = new_n1152_ & ~new_n5955_;
  assign new_n5957_ = new_n1156_ & ~new_n5956_;
  assign new_n5958_ = new_n1160_ & ~new_n5957_;
  assign new_n5959_ = new_n1164_ & ~new_n5958_;
  assign new_n5960_ = new_n1168_ & ~new_n5959_;
  assign new_n5961_ = new_n1172_ & ~new_n5960_;
  assign new_n5962_ = new_n1176_ & ~new_n5961_;
  assign new_n5963_ = new_n1180_ & ~new_n5962_;
  assign new_n5964_ = new_n1184_ & ~new_n5963_;
  assign new_n5965_ = new_n1188_ & ~new_n5964_;
  assign new_n5966_ = new_n1192_ & ~new_n5965_;
  assign new_n5967_ = new_n1196_ & ~new_n5966_;
  assign new_n5968_ = \req[55]  & ~new_n1198_;
  assign \grant[55]  = ~new_n5967_ & new_n5968_;
  assign new_n5970_ = ~new_n535_ & new_n1207_;
  assign new_n5971_ = new_n1212_ & ~new_n5970_;
  assign new_n5972_ = new_n1216_ & ~new_n5971_;
  assign new_n5973_ = new_n1220_ & ~new_n5972_;
  assign new_n5974_ = new_n1224_ & ~new_n5973_;
  assign new_n5975_ = new_n1228_ & ~new_n5974_;
  assign new_n5976_ = new_n1232_ & ~new_n5975_;
  assign new_n5977_ = new_n1236_ & ~new_n5976_;
  assign new_n5978_ = new_n1240_ & ~new_n5977_;
  assign new_n5979_ = new_n1244_ & ~new_n5978_;
  assign new_n5980_ = new_n1248_ & ~new_n5979_;
  assign new_n5981_ = new_n1252_ & ~new_n5980_;
  assign new_n5982_ = new_n1256_ & ~new_n5981_;
  assign new_n5983_ = new_n1260_ & ~new_n5982_;
  assign new_n5984_ = new_n1264_ & ~new_n5983_;
  assign new_n5985_ = new_n1268_ & ~new_n5984_;
  assign new_n5986_ = new_n1272_ & ~new_n5985_;
  assign new_n5987_ = new_n1276_ & ~new_n5986_;
  assign new_n5988_ = new_n1280_ & ~new_n5987_;
  assign new_n5989_ = new_n1284_ & ~new_n5988_;
  assign new_n5990_ = new_n1288_ & ~new_n5989_;
  assign new_n5991_ = new_n1292_ & ~new_n5990_;
  assign new_n5992_ = new_n1296_ & ~new_n5991_;
  assign new_n5993_ = new_n1300_ & ~new_n5992_;
  assign new_n5994_ = new_n1304_ & ~new_n5993_;
  assign new_n5995_ = new_n1308_ & ~new_n5994_;
  assign new_n5996_ = new_n1312_ & ~new_n5995_;
  assign new_n5997_ = new_n1316_ & ~new_n5996_;
  assign new_n5998_ = new_n1320_ & ~new_n5997_;
  assign new_n5999_ = new_n1324_ & ~new_n5998_;
  assign new_n6000_ = new_n1328_ & ~new_n5999_;
  assign new_n6001_ = new_n1332_ & ~new_n6000_;
  assign new_n6002_ = new_n1336_ & ~new_n6001_;
  assign new_n6003_ = new_n1340_ & ~new_n6002_;
  assign new_n6004_ = new_n1344_ & ~new_n6003_;
  assign new_n6005_ = new_n1348_ & ~new_n6004_;
  assign new_n6006_ = new_n1352_ & ~new_n6005_;
  assign new_n6007_ = new_n1356_ & ~new_n6006_;
  assign new_n6008_ = new_n1360_ & ~new_n6007_;
  assign new_n6009_ = new_n1364_ & ~new_n6008_;
  assign new_n6010_ = new_n1368_ & ~new_n6009_;
  assign new_n6011_ = new_n1372_ & ~new_n6010_;
  assign new_n6012_ = new_n1376_ & ~new_n6011_;
  assign new_n6013_ = new_n1380_ & ~new_n6012_;
  assign new_n6014_ = new_n1384_ & ~new_n6013_;
  assign new_n6015_ = new_n1388_ & ~new_n6014_;
  assign new_n6016_ = new_n1392_ & ~new_n6015_;
  assign new_n6017_ = new_n1396_ & ~new_n6016_;
  assign new_n6018_ = new_n1663_ & ~new_n6017_;
  assign new_n6019_ = new_n392_ & ~new_n6018_;
  assign new_n6020_ = new_n396_ & ~new_n6019_;
  assign new_n6021_ = new_n400_ & ~new_n6020_;
  assign new_n6022_ = new_n404_ & ~new_n6021_;
  assign new_n6023_ = new_n408_ & ~new_n6022_;
  assign new_n6024_ = new_n412_ & ~new_n6023_;
  assign new_n6025_ = new_n416_ & ~new_n6024_;
  assign new_n6026_ = new_n420_ & ~new_n6025_;
  assign new_n6027_ = new_n424_ & ~new_n6026_;
  assign new_n6028_ = new_n428_ & ~new_n6027_;
  assign new_n6029_ = new_n432_ & ~new_n6028_;
  assign new_n6030_ = new_n436_ & ~new_n6029_;
  assign new_n6031_ = new_n440_ & ~new_n6030_;
  assign new_n6032_ = new_n444_ & ~new_n6031_;
  assign new_n6033_ = new_n448_ & ~new_n6032_;
  assign new_n6034_ = new_n452_ & ~new_n6033_;
  assign new_n6035_ = new_n456_ & ~new_n6034_;
  assign new_n6036_ = new_n460_ & ~new_n6035_;
  assign new_n6037_ = new_n464_ & ~new_n6036_;
  assign new_n6038_ = new_n468_ & ~new_n6037_;
  assign new_n6039_ = new_n472_ & ~new_n6038_;
  assign new_n6040_ = new_n476_ & ~new_n6039_;
  assign new_n6041_ = new_n480_ & ~new_n6040_;
  assign new_n6042_ = new_n484_ & ~new_n6041_;
  assign new_n6043_ = new_n488_ & ~new_n6042_;
  assign new_n6044_ = new_n492_ & ~new_n6043_;
  assign new_n6045_ = new_n496_ & ~new_n6044_;
  assign new_n6046_ = new_n500_ & ~new_n6045_;
  assign new_n6047_ = new_n504_ & ~new_n6046_;
  assign new_n6048_ = new_n508_ & ~new_n6047_;
  assign new_n6049_ = new_n512_ & ~new_n6048_;
  assign new_n6050_ = new_n516_ & ~new_n6049_;
  assign new_n6051_ = new_n520_ & ~new_n6050_;
  assign new_n6052_ = new_n524_ & ~new_n6051_;
  assign new_n6053_ = new_n528_ & ~new_n6052_;
  assign new_n6054_ = \req[56]  & ~new_n530_;
  assign \grant[56]  = ~new_n6053_ & new_n6054_;
  assign new_n6056_ = new_n539_ & ~new_n874_;
  assign new_n6057_ = new_n544_ & ~new_n6056_;
  assign new_n6058_ = new_n548_ & ~new_n6057_;
  assign new_n6059_ = new_n552_ & ~new_n6058_;
  assign new_n6060_ = new_n556_ & ~new_n6059_;
  assign new_n6061_ = new_n560_ & ~new_n6060_;
  assign new_n6062_ = new_n564_ & ~new_n6061_;
  assign new_n6063_ = new_n568_ & ~new_n6062_;
  assign new_n6064_ = new_n572_ & ~new_n6063_;
  assign new_n6065_ = new_n576_ & ~new_n6064_;
  assign new_n6066_ = new_n580_ & ~new_n6065_;
  assign new_n6067_ = new_n584_ & ~new_n6066_;
  assign new_n6068_ = new_n588_ & ~new_n6067_;
  assign new_n6069_ = new_n592_ & ~new_n6068_;
  assign new_n6070_ = new_n596_ & ~new_n6069_;
  assign new_n6071_ = new_n600_ & ~new_n6070_;
  assign new_n6072_ = new_n604_ & ~new_n6071_;
  assign new_n6073_ = new_n608_ & ~new_n6072_;
  assign new_n6074_ = new_n612_ & ~new_n6073_;
  assign new_n6075_ = new_n616_ & ~new_n6074_;
  assign new_n6076_ = new_n620_ & ~new_n6075_;
  assign new_n6077_ = new_n624_ & ~new_n6076_;
  assign new_n6078_ = new_n628_ & ~new_n6077_;
  assign new_n6079_ = new_n632_ & ~new_n6078_;
  assign new_n6080_ = new_n636_ & ~new_n6079_;
  assign new_n6081_ = new_n640_ & ~new_n6080_;
  assign new_n6082_ = new_n644_ & ~new_n6081_;
  assign new_n6083_ = new_n648_ & ~new_n6082_;
  assign new_n6084_ = new_n652_ & ~new_n6083_;
  assign new_n6085_ = new_n656_ & ~new_n6084_;
  assign new_n6086_ = new_n660_ & ~new_n6085_;
  assign new_n6087_ = new_n664_ & ~new_n6086_;
  assign new_n6088_ = new_n668_ & ~new_n6087_;
  assign new_n6089_ = new_n672_ & ~new_n6088_;
  assign new_n6090_ = new_n676_ & ~new_n6089_;
  assign new_n6091_ = new_n680_ & ~new_n6090_;
  assign new_n6092_ = new_n684_ & ~new_n6091_;
  assign new_n6093_ = new_n688_ & ~new_n6092_;
  assign new_n6094_ = new_n692_ & ~new_n6093_;
  assign new_n6095_ = new_n696_ & ~new_n6094_;
  assign new_n6096_ = new_n700_ & ~new_n6095_;
  assign new_n6097_ = new_n704_ & ~new_n6096_;
  assign new_n6098_ = new_n708_ & ~new_n6097_;
  assign new_n6099_ = new_n712_ & ~new_n6098_;
  assign new_n6100_ = new_n716_ & ~new_n6099_;
  assign new_n6101_ = new_n720_ & ~new_n6100_;
  assign new_n6102_ = new_n1484_ & ~new_n6101_;
  assign new_n6103_ = new_n1486_ & ~new_n6102_;
  assign new_n6104_ = new_n1750_ & ~new_n6103_;
  assign new_n6105_ = new_n731_ & ~new_n6104_;
  assign new_n6106_ = new_n735_ & ~new_n6105_;
  assign new_n6107_ = new_n739_ & ~new_n6106_;
  assign new_n6108_ = new_n743_ & ~new_n6107_;
  assign new_n6109_ = new_n747_ & ~new_n6108_;
  assign new_n6110_ = new_n751_ & ~new_n6109_;
  assign new_n6111_ = new_n755_ & ~new_n6110_;
  assign new_n6112_ = new_n759_ & ~new_n6111_;
  assign new_n6113_ = new_n763_ & ~new_n6112_;
  assign new_n6114_ = new_n767_ & ~new_n6113_;
  assign new_n6115_ = new_n771_ & ~new_n6114_;
  assign new_n6116_ = new_n775_ & ~new_n6115_;
  assign new_n6117_ = new_n779_ & ~new_n6116_;
  assign new_n6118_ = new_n783_ & ~new_n6117_;
  assign new_n6119_ = new_n787_ & ~new_n6118_;
  assign new_n6120_ = new_n791_ & ~new_n6119_;
  assign new_n6121_ = new_n795_ & ~new_n6120_;
  assign new_n6122_ = new_n799_ & ~new_n6121_;
  assign new_n6123_ = new_n803_ & ~new_n6122_;
  assign new_n6124_ = new_n807_ & ~new_n6123_;
  assign new_n6125_ = new_n811_ & ~new_n6124_;
  assign new_n6126_ = new_n815_ & ~new_n6125_;
  assign new_n6127_ = new_n819_ & ~new_n6126_;
  assign new_n6128_ = new_n823_ & ~new_n6127_;
  assign new_n6129_ = new_n827_ & ~new_n6128_;
  assign new_n6130_ = new_n831_ & ~new_n6129_;
  assign new_n6131_ = new_n835_ & ~new_n6130_;
  assign new_n6132_ = new_n839_ & ~new_n6131_;
  assign new_n6133_ = new_n843_ & ~new_n6132_;
  assign new_n6134_ = new_n847_ & ~new_n6133_;
  assign new_n6135_ = new_n851_ & ~new_n6134_;
  assign new_n6136_ = new_n855_ & ~new_n6135_;
  assign new_n6137_ = new_n859_ & ~new_n6136_;
  assign new_n6138_ = new_n863_ & ~new_n6137_;
  assign new_n6139_ = new_n867_ & ~new_n6138_;
  assign new_n6140_ = \req[57]  & ~new_n869_;
  assign \grant[57]  = ~new_n6139_ & new_n6140_;
  assign new_n6142_ = new_n878_ & ~new_n1211_;
  assign new_n6143_ = new_n883_ & ~new_n6142_;
  assign new_n6144_ = new_n887_ & ~new_n6143_;
  assign new_n6145_ = new_n891_ & ~new_n6144_;
  assign new_n6146_ = new_n895_ & ~new_n6145_;
  assign new_n6147_ = new_n899_ & ~new_n6146_;
  assign new_n6148_ = new_n903_ & ~new_n6147_;
  assign new_n6149_ = new_n907_ & ~new_n6148_;
  assign new_n6150_ = new_n911_ & ~new_n6149_;
  assign new_n6151_ = new_n915_ & ~new_n6150_;
  assign new_n6152_ = new_n919_ & ~new_n6151_;
  assign new_n6153_ = new_n923_ & ~new_n6152_;
  assign new_n6154_ = new_n927_ & ~new_n6153_;
  assign new_n6155_ = new_n931_ & ~new_n6154_;
  assign new_n6156_ = new_n935_ & ~new_n6155_;
  assign new_n6157_ = new_n939_ & ~new_n6156_;
  assign new_n6158_ = new_n943_ & ~new_n6157_;
  assign new_n6159_ = new_n947_ & ~new_n6158_;
  assign new_n6160_ = new_n951_ & ~new_n6159_;
  assign new_n6161_ = new_n955_ & ~new_n6160_;
  assign new_n6162_ = new_n959_ & ~new_n6161_;
  assign new_n6163_ = new_n963_ & ~new_n6162_;
  assign new_n6164_ = new_n967_ & ~new_n6163_;
  assign new_n6165_ = new_n971_ & ~new_n6164_;
  assign new_n6166_ = new_n975_ & ~new_n6165_;
  assign new_n6167_ = new_n979_ & ~new_n6166_;
  assign new_n6168_ = new_n983_ & ~new_n6167_;
  assign new_n6169_ = new_n987_ & ~new_n6168_;
  assign new_n6170_ = new_n991_ & ~new_n6169_;
  assign new_n6171_ = new_n995_ & ~new_n6170_;
  assign new_n6172_ = new_n999_ & ~new_n6171_;
  assign new_n6173_ = new_n1003_ & ~new_n6172_;
  assign new_n6174_ = new_n1007_ & ~new_n6173_;
  assign new_n6175_ = new_n1011_ & ~new_n6174_;
  assign new_n6176_ = new_n1015_ & ~new_n6175_;
  assign new_n6177_ = new_n1019_ & ~new_n6176_;
  assign new_n6178_ = new_n1023_ & ~new_n6177_;
  assign new_n6179_ = new_n1027_ & ~new_n6178_;
  assign new_n6180_ = new_n1031_ & ~new_n6179_;
  assign new_n6181_ = new_n1035_ & ~new_n6180_;
  assign new_n6182_ = new_n1039_ & ~new_n6181_;
  assign new_n6183_ = new_n1043_ & ~new_n6182_;
  assign new_n6184_ = new_n1047_ & ~new_n6183_;
  assign new_n6185_ = new_n1051_ & ~new_n6184_;
  assign new_n6186_ = new_n1055_ & ~new_n6185_;
  assign new_n6187_ = new_n1059_ & ~new_n6186_;
  assign new_n6188_ = new_n1574_ & ~new_n6187_;
  assign new_n6189_ = new_n1576_ & ~new_n6188_;
  assign new_n6190_ = new_n1837_ & ~new_n6189_;
  assign new_n6191_ = new_n1068_ & ~new_n6190_;
  assign new_n6192_ = new_n1072_ & ~new_n6191_;
  assign new_n6193_ = new_n1076_ & ~new_n6192_;
  assign new_n6194_ = new_n1080_ & ~new_n6193_;
  assign new_n6195_ = new_n1084_ & ~new_n6194_;
  assign new_n6196_ = new_n1088_ & ~new_n6195_;
  assign new_n6197_ = new_n1092_ & ~new_n6196_;
  assign new_n6198_ = new_n1096_ & ~new_n6197_;
  assign new_n6199_ = new_n1100_ & ~new_n6198_;
  assign new_n6200_ = new_n1104_ & ~new_n6199_;
  assign new_n6201_ = new_n1108_ & ~new_n6200_;
  assign new_n6202_ = new_n1112_ & ~new_n6201_;
  assign new_n6203_ = new_n1116_ & ~new_n6202_;
  assign new_n6204_ = new_n1120_ & ~new_n6203_;
  assign new_n6205_ = new_n1124_ & ~new_n6204_;
  assign new_n6206_ = new_n1128_ & ~new_n6205_;
  assign new_n6207_ = new_n1132_ & ~new_n6206_;
  assign new_n6208_ = new_n1136_ & ~new_n6207_;
  assign new_n6209_ = new_n1140_ & ~new_n6208_;
  assign new_n6210_ = new_n1144_ & ~new_n6209_;
  assign new_n6211_ = new_n1148_ & ~new_n6210_;
  assign new_n6212_ = new_n1152_ & ~new_n6211_;
  assign new_n6213_ = new_n1156_ & ~new_n6212_;
  assign new_n6214_ = new_n1160_ & ~new_n6213_;
  assign new_n6215_ = new_n1164_ & ~new_n6214_;
  assign new_n6216_ = new_n1168_ & ~new_n6215_;
  assign new_n6217_ = new_n1172_ & ~new_n6216_;
  assign new_n6218_ = new_n1176_ & ~new_n6217_;
  assign new_n6219_ = new_n1180_ & ~new_n6218_;
  assign new_n6220_ = new_n1184_ & ~new_n6219_;
  assign new_n6221_ = new_n1188_ & ~new_n6220_;
  assign new_n6222_ = new_n1192_ & ~new_n6221_;
  assign new_n6223_ = new_n1196_ & ~new_n6222_;
  assign new_n6224_ = new_n1200_ & ~new_n6223_;
  assign new_n6225_ = new_n1204_ & ~new_n6224_;
  assign new_n6226_ = \req[58]  & ~new_n1206_;
  assign \grant[58]  = ~new_n6225_ & new_n6226_;
  assign new_n6228_ = ~new_n543_ & new_n1215_;
  assign new_n6229_ = new_n1220_ & ~new_n6228_;
  assign new_n6230_ = new_n1224_ & ~new_n6229_;
  assign new_n6231_ = new_n1228_ & ~new_n6230_;
  assign new_n6232_ = new_n1232_ & ~new_n6231_;
  assign new_n6233_ = new_n1236_ & ~new_n6232_;
  assign new_n6234_ = new_n1240_ & ~new_n6233_;
  assign new_n6235_ = new_n1244_ & ~new_n6234_;
  assign new_n6236_ = new_n1248_ & ~new_n6235_;
  assign new_n6237_ = new_n1252_ & ~new_n6236_;
  assign new_n6238_ = new_n1256_ & ~new_n6237_;
  assign new_n6239_ = new_n1260_ & ~new_n6238_;
  assign new_n6240_ = new_n1264_ & ~new_n6239_;
  assign new_n6241_ = new_n1268_ & ~new_n6240_;
  assign new_n6242_ = new_n1272_ & ~new_n6241_;
  assign new_n6243_ = new_n1276_ & ~new_n6242_;
  assign new_n6244_ = new_n1280_ & ~new_n6243_;
  assign new_n6245_ = new_n1284_ & ~new_n6244_;
  assign new_n6246_ = new_n1288_ & ~new_n6245_;
  assign new_n6247_ = new_n1292_ & ~new_n6246_;
  assign new_n6248_ = new_n1296_ & ~new_n6247_;
  assign new_n6249_ = new_n1300_ & ~new_n6248_;
  assign new_n6250_ = new_n1304_ & ~new_n6249_;
  assign new_n6251_ = new_n1308_ & ~new_n6250_;
  assign new_n6252_ = new_n1312_ & ~new_n6251_;
  assign new_n6253_ = new_n1316_ & ~new_n6252_;
  assign new_n6254_ = new_n1320_ & ~new_n6253_;
  assign new_n6255_ = new_n1324_ & ~new_n6254_;
  assign new_n6256_ = new_n1328_ & ~new_n6255_;
  assign new_n6257_ = new_n1332_ & ~new_n6256_;
  assign new_n6258_ = new_n1336_ & ~new_n6257_;
  assign new_n6259_ = new_n1340_ & ~new_n6258_;
  assign new_n6260_ = new_n1344_ & ~new_n6259_;
  assign new_n6261_ = new_n1348_ & ~new_n6260_;
  assign new_n6262_ = new_n1352_ & ~new_n6261_;
  assign new_n6263_ = new_n1356_ & ~new_n6262_;
  assign new_n6264_ = new_n1360_ & ~new_n6263_;
  assign new_n6265_ = new_n1364_ & ~new_n6264_;
  assign new_n6266_ = new_n1368_ & ~new_n6265_;
  assign new_n6267_ = new_n1372_ & ~new_n6266_;
  assign new_n6268_ = new_n1376_ & ~new_n6267_;
  assign new_n6269_ = new_n1380_ & ~new_n6268_;
  assign new_n6270_ = new_n1384_ & ~new_n6269_;
  assign new_n6271_ = new_n1388_ & ~new_n6270_;
  assign new_n6272_ = new_n1392_ & ~new_n6271_;
  assign new_n6273_ = new_n1396_ & ~new_n6272_;
  assign new_n6274_ = new_n1663_ & ~new_n6273_;
  assign new_n6275_ = new_n392_ & ~new_n6274_;
  assign new_n6276_ = new_n396_ & ~new_n6275_;
  assign new_n6277_ = new_n400_ & ~new_n6276_;
  assign new_n6278_ = new_n404_ & ~new_n6277_;
  assign new_n6279_ = new_n408_ & ~new_n6278_;
  assign new_n6280_ = new_n412_ & ~new_n6279_;
  assign new_n6281_ = new_n416_ & ~new_n6280_;
  assign new_n6282_ = new_n420_ & ~new_n6281_;
  assign new_n6283_ = new_n424_ & ~new_n6282_;
  assign new_n6284_ = new_n428_ & ~new_n6283_;
  assign new_n6285_ = new_n432_ & ~new_n6284_;
  assign new_n6286_ = new_n436_ & ~new_n6285_;
  assign new_n6287_ = new_n440_ & ~new_n6286_;
  assign new_n6288_ = new_n444_ & ~new_n6287_;
  assign new_n6289_ = new_n448_ & ~new_n6288_;
  assign new_n6290_ = new_n452_ & ~new_n6289_;
  assign new_n6291_ = new_n456_ & ~new_n6290_;
  assign new_n6292_ = new_n460_ & ~new_n6291_;
  assign new_n6293_ = new_n464_ & ~new_n6292_;
  assign new_n6294_ = new_n468_ & ~new_n6293_;
  assign new_n6295_ = new_n472_ & ~new_n6294_;
  assign new_n6296_ = new_n476_ & ~new_n6295_;
  assign new_n6297_ = new_n480_ & ~new_n6296_;
  assign new_n6298_ = new_n484_ & ~new_n6297_;
  assign new_n6299_ = new_n488_ & ~new_n6298_;
  assign new_n6300_ = new_n492_ & ~new_n6299_;
  assign new_n6301_ = new_n496_ & ~new_n6300_;
  assign new_n6302_ = new_n500_ & ~new_n6301_;
  assign new_n6303_ = new_n504_ & ~new_n6302_;
  assign new_n6304_ = new_n508_ & ~new_n6303_;
  assign new_n6305_ = new_n512_ & ~new_n6304_;
  assign new_n6306_ = new_n516_ & ~new_n6305_;
  assign new_n6307_ = new_n520_ & ~new_n6306_;
  assign new_n6308_ = new_n524_ & ~new_n6307_;
  assign new_n6309_ = new_n528_ & ~new_n6308_;
  assign new_n6310_ = new_n532_ & ~new_n6309_;
  assign new_n6311_ = new_n536_ & ~new_n6310_;
  assign new_n6312_ = \req[59]  & ~new_n538_;
  assign \grant[59]  = ~new_n6311_ & new_n6312_;
  assign new_n6314_ = new_n547_ & ~new_n882_;
  assign new_n6315_ = new_n552_ & ~new_n6314_;
  assign new_n6316_ = new_n556_ & ~new_n6315_;
  assign new_n6317_ = new_n560_ & ~new_n6316_;
  assign new_n6318_ = new_n564_ & ~new_n6317_;
  assign new_n6319_ = new_n568_ & ~new_n6318_;
  assign new_n6320_ = new_n572_ & ~new_n6319_;
  assign new_n6321_ = new_n576_ & ~new_n6320_;
  assign new_n6322_ = new_n580_ & ~new_n6321_;
  assign new_n6323_ = new_n584_ & ~new_n6322_;
  assign new_n6324_ = new_n588_ & ~new_n6323_;
  assign new_n6325_ = new_n592_ & ~new_n6324_;
  assign new_n6326_ = new_n596_ & ~new_n6325_;
  assign new_n6327_ = new_n600_ & ~new_n6326_;
  assign new_n6328_ = new_n604_ & ~new_n6327_;
  assign new_n6329_ = new_n608_ & ~new_n6328_;
  assign new_n6330_ = new_n612_ & ~new_n6329_;
  assign new_n6331_ = new_n616_ & ~new_n6330_;
  assign new_n6332_ = new_n620_ & ~new_n6331_;
  assign new_n6333_ = new_n624_ & ~new_n6332_;
  assign new_n6334_ = new_n628_ & ~new_n6333_;
  assign new_n6335_ = new_n632_ & ~new_n6334_;
  assign new_n6336_ = new_n636_ & ~new_n6335_;
  assign new_n6337_ = new_n640_ & ~new_n6336_;
  assign new_n6338_ = new_n644_ & ~new_n6337_;
  assign new_n6339_ = new_n648_ & ~new_n6338_;
  assign new_n6340_ = new_n652_ & ~new_n6339_;
  assign new_n6341_ = new_n656_ & ~new_n6340_;
  assign new_n6342_ = new_n660_ & ~new_n6341_;
  assign new_n6343_ = new_n664_ & ~new_n6342_;
  assign new_n6344_ = new_n668_ & ~new_n6343_;
  assign new_n6345_ = new_n672_ & ~new_n6344_;
  assign new_n6346_ = new_n676_ & ~new_n6345_;
  assign new_n6347_ = new_n680_ & ~new_n6346_;
  assign new_n6348_ = new_n684_ & ~new_n6347_;
  assign new_n6349_ = new_n688_ & ~new_n6348_;
  assign new_n6350_ = new_n692_ & ~new_n6349_;
  assign new_n6351_ = new_n696_ & ~new_n6350_;
  assign new_n6352_ = new_n700_ & ~new_n6351_;
  assign new_n6353_ = new_n704_ & ~new_n6352_;
  assign new_n6354_ = new_n708_ & ~new_n6353_;
  assign new_n6355_ = new_n712_ & ~new_n6354_;
  assign new_n6356_ = new_n716_ & ~new_n6355_;
  assign new_n6357_ = new_n720_ & ~new_n6356_;
  assign new_n6358_ = new_n1484_ & ~new_n6357_;
  assign new_n6359_ = new_n1486_ & ~new_n6358_;
  assign new_n6360_ = new_n1750_ & ~new_n6359_;
  assign new_n6361_ = new_n731_ & ~new_n6360_;
  assign new_n6362_ = new_n735_ & ~new_n6361_;
  assign new_n6363_ = new_n739_ & ~new_n6362_;
  assign new_n6364_ = new_n743_ & ~new_n6363_;
  assign new_n6365_ = new_n747_ & ~new_n6364_;
  assign new_n6366_ = new_n751_ & ~new_n6365_;
  assign new_n6367_ = new_n755_ & ~new_n6366_;
  assign new_n6368_ = new_n759_ & ~new_n6367_;
  assign new_n6369_ = new_n763_ & ~new_n6368_;
  assign new_n6370_ = new_n767_ & ~new_n6369_;
  assign new_n6371_ = new_n771_ & ~new_n6370_;
  assign new_n6372_ = new_n775_ & ~new_n6371_;
  assign new_n6373_ = new_n779_ & ~new_n6372_;
  assign new_n6374_ = new_n783_ & ~new_n6373_;
  assign new_n6375_ = new_n787_ & ~new_n6374_;
  assign new_n6376_ = new_n791_ & ~new_n6375_;
  assign new_n6377_ = new_n795_ & ~new_n6376_;
  assign new_n6378_ = new_n799_ & ~new_n6377_;
  assign new_n6379_ = new_n803_ & ~new_n6378_;
  assign new_n6380_ = new_n807_ & ~new_n6379_;
  assign new_n6381_ = new_n811_ & ~new_n6380_;
  assign new_n6382_ = new_n815_ & ~new_n6381_;
  assign new_n6383_ = new_n819_ & ~new_n6382_;
  assign new_n6384_ = new_n823_ & ~new_n6383_;
  assign new_n6385_ = new_n827_ & ~new_n6384_;
  assign new_n6386_ = new_n831_ & ~new_n6385_;
  assign new_n6387_ = new_n835_ & ~new_n6386_;
  assign new_n6388_ = new_n839_ & ~new_n6387_;
  assign new_n6389_ = new_n843_ & ~new_n6388_;
  assign new_n6390_ = new_n847_ & ~new_n6389_;
  assign new_n6391_ = new_n851_ & ~new_n6390_;
  assign new_n6392_ = new_n855_ & ~new_n6391_;
  assign new_n6393_ = new_n859_ & ~new_n6392_;
  assign new_n6394_ = new_n863_ & ~new_n6393_;
  assign new_n6395_ = new_n867_ & ~new_n6394_;
  assign new_n6396_ = new_n871_ & ~new_n6395_;
  assign new_n6397_ = new_n875_ & ~new_n6396_;
  assign new_n6398_ = \req[60]  & ~new_n877_;
  assign \grant[60]  = ~new_n6397_ & new_n6398_;
  assign new_n6400_ = new_n886_ & ~new_n1219_;
  assign new_n6401_ = new_n891_ & ~new_n6400_;
  assign new_n6402_ = new_n895_ & ~new_n6401_;
  assign new_n6403_ = new_n899_ & ~new_n6402_;
  assign new_n6404_ = new_n903_ & ~new_n6403_;
  assign new_n6405_ = new_n907_ & ~new_n6404_;
  assign new_n6406_ = new_n911_ & ~new_n6405_;
  assign new_n6407_ = new_n915_ & ~new_n6406_;
  assign new_n6408_ = new_n919_ & ~new_n6407_;
  assign new_n6409_ = new_n923_ & ~new_n6408_;
  assign new_n6410_ = new_n927_ & ~new_n6409_;
  assign new_n6411_ = new_n931_ & ~new_n6410_;
  assign new_n6412_ = new_n935_ & ~new_n6411_;
  assign new_n6413_ = new_n939_ & ~new_n6412_;
  assign new_n6414_ = new_n943_ & ~new_n6413_;
  assign new_n6415_ = new_n947_ & ~new_n6414_;
  assign new_n6416_ = new_n951_ & ~new_n6415_;
  assign new_n6417_ = new_n955_ & ~new_n6416_;
  assign new_n6418_ = new_n959_ & ~new_n6417_;
  assign new_n6419_ = new_n963_ & ~new_n6418_;
  assign new_n6420_ = new_n967_ & ~new_n6419_;
  assign new_n6421_ = new_n971_ & ~new_n6420_;
  assign new_n6422_ = new_n975_ & ~new_n6421_;
  assign new_n6423_ = new_n979_ & ~new_n6422_;
  assign new_n6424_ = new_n983_ & ~new_n6423_;
  assign new_n6425_ = new_n987_ & ~new_n6424_;
  assign new_n6426_ = new_n991_ & ~new_n6425_;
  assign new_n6427_ = new_n995_ & ~new_n6426_;
  assign new_n6428_ = new_n999_ & ~new_n6427_;
  assign new_n6429_ = new_n1003_ & ~new_n6428_;
  assign new_n6430_ = new_n1007_ & ~new_n6429_;
  assign new_n6431_ = new_n1011_ & ~new_n6430_;
  assign new_n6432_ = new_n1015_ & ~new_n6431_;
  assign new_n6433_ = new_n1019_ & ~new_n6432_;
  assign new_n6434_ = new_n1023_ & ~new_n6433_;
  assign new_n6435_ = new_n1027_ & ~new_n6434_;
  assign new_n6436_ = new_n1031_ & ~new_n6435_;
  assign new_n6437_ = new_n1035_ & ~new_n6436_;
  assign new_n6438_ = new_n1039_ & ~new_n6437_;
  assign new_n6439_ = new_n1043_ & ~new_n6438_;
  assign new_n6440_ = new_n1047_ & ~new_n6439_;
  assign new_n6441_ = new_n1051_ & ~new_n6440_;
  assign new_n6442_ = new_n1055_ & ~new_n6441_;
  assign new_n6443_ = new_n1059_ & ~new_n6442_;
  assign new_n6444_ = new_n1574_ & ~new_n6443_;
  assign new_n6445_ = new_n1576_ & ~new_n6444_;
  assign new_n6446_ = new_n1837_ & ~new_n6445_;
  assign new_n6447_ = new_n1068_ & ~new_n6446_;
  assign new_n6448_ = new_n1072_ & ~new_n6447_;
  assign new_n6449_ = new_n1076_ & ~new_n6448_;
  assign new_n6450_ = new_n1080_ & ~new_n6449_;
  assign new_n6451_ = new_n1084_ & ~new_n6450_;
  assign new_n6452_ = new_n1088_ & ~new_n6451_;
  assign new_n6453_ = new_n1092_ & ~new_n6452_;
  assign new_n6454_ = new_n1096_ & ~new_n6453_;
  assign new_n6455_ = new_n1100_ & ~new_n6454_;
  assign new_n6456_ = new_n1104_ & ~new_n6455_;
  assign new_n6457_ = new_n1108_ & ~new_n6456_;
  assign new_n6458_ = new_n1112_ & ~new_n6457_;
  assign new_n6459_ = new_n1116_ & ~new_n6458_;
  assign new_n6460_ = new_n1120_ & ~new_n6459_;
  assign new_n6461_ = new_n1124_ & ~new_n6460_;
  assign new_n6462_ = new_n1128_ & ~new_n6461_;
  assign new_n6463_ = new_n1132_ & ~new_n6462_;
  assign new_n6464_ = new_n1136_ & ~new_n6463_;
  assign new_n6465_ = new_n1140_ & ~new_n6464_;
  assign new_n6466_ = new_n1144_ & ~new_n6465_;
  assign new_n6467_ = new_n1148_ & ~new_n6466_;
  assign new_n6468_ = new_n1152_ & ~new_n6467_;
  assign new_n6469_ = new_n1156_ & ~new_n6468_;
  assign new_n6470_ = new_n1160_ & ~new_n6469_;
  assign new_n6471_ = new_n1164_ & ~new_n6470_;
  assign new_n6472_ = new_n1168_ & ~new_n6471_;
  assign new_n6473_ = new_n1172_ & ~new_n6472_;
  assign new_n6474_ = new_n1176_ & ~new_n6473_;
  assign new_n6475_ = new_n1180_ & ~new_n6474_;
  assign new_n6476_ = new_n1184_ & ~new_n6475_;
  assign new_n6477_ = new_n1188_ & ~new_n6476_;
  assign new_n6478_ = new_n1192_ & ~new_n6477_;
  assign new_n6479_ = new_n1196_ & ~new_n6478_;
  assign new_n6480_ = new_n1200_ & ~new_n6479_;
  assign new_n6481_ = new_n1204_ & ~new_n6480_;
  assign new_n6482_ = new_n1208_ & ~new_n6481_;
  assign new_n6483_ = new_n1212_ & ~new_n6482_;
  assign new_n6484_ = \req[61]  & ~new_n1214_;
  assign \grant[61]  = ~new_n6483_ & new_n6484_;
  assign new_n6486_ = ~new_n551_ & new_n1223_;
  assign new_n6487_ = new_n1228_ & ~new_n6486_;
  assign new_n6488_ = new_n1232_ & ~new_n6487_;
  assign new_n6489_ = new_n1236_ & ~new_n6488_;
  assign new_n6490_ = new_n1240_ & ~new_n6489_;
  assign new_n6491_ = new_n1244_ & ~new_n6490_;
  assign new_n6492_ = new_n1248_ & ~new_n6491_;
  assign new_n6493_ = new_n1252_ & ~new_n6492_;
  assign new_n6494_ = new_n1256_ & ~new_n6493_;
  assign new_n6495_ = new_n1260_ & ~new_n6494_;
  assign new_n6496_ = new_n1264_ & ~new_n6495_;
  assign new_n6497_ = new_n1268_ & ~new_n6496_;
  assign new_n6498_ = new_n1272_ & ~new_n6497_;
  assign new_n6499_ = new_n1276_ & ~new_n6498_;
  assign new_n6500_ = new_n1280_ & ~new_n6499_;
  assign new_n6501_ = new_n1284_ & ~new_n6500_;
  assign new_n6502_ = new_n1288_ & ~new_n6501_;
  assign new_n6503_ = new_n1292_ & ~new_n6502_;
  assign new_n6504_ = new_n1296_ & ~new_n6503_;
  assign new_n6505_ = new_n1300_ & ~new_n6504_;
  assign new_n6506_ = new_n1304_ & ~new_n6505_;
  assign new_n6507_ = new_n1308_ & ~new_n6506_;
  assign new_n6508_ = new_n1312_ & ~new_n6507_;
  assign new_n6509_ = new_n1316_ & ~new_n6508_;
  assign new_n6510_ = new_n1320_ & ~new_n6509_;
  assign new_n6511_ = new_n1324_ & ~new_n6510_;
  assign new_n6512_ = new_n1328_ & ~new_n6511_;
  assign new_n6513_ = new_n1332_ & ~new_n6512_;
  assign new_n6514_ = new_n1336_ & ~new_n6513_;
  assign new_n6515_ = new_n1340_ & ~new_n6514_;
  assign new_n6516_ = new_n1344_ & ~new_n6515_;
  assign new_n6517_ = new_n1348_ & ~new_n6516_;
  assign new_n6518_ = new_n1352_ & ~new_n6517_;
  assign new_n6519_ = new_n1356_ & ~new_n6518_;
  assign new_n6520_ = new_n1360_ & ~new_n6519_;
  assign new_n6521_ = new_n1364_ & ~new_n6520_;
  assign new_n6522_ = new_n1368_ & ~new_n6521_;
  assign new_n6523_ = new_n1372_ & ~new_n6522_;
  assign new_n6524_ = new_n1376_ & ~new_n6523_;
  assign new_n6525_ = new_n1380_ & ~new_n6524_;
  assign new_n6526_ = new_n1384_ & ~new_n6525_;
  assign new_n6527_ = new_n1388_ & ~new_n6526_;
  assign new_n6528_ = new_n1392_ & ~new_n6527_;
  assign new_n6529_ = new_n1396_ & ~new_n6528_;
  assign new_n6530_ = new_n1663_ & ~new_n6529_;
  assign new_n6531_ = new_n392_ & ~new_n6530_;
  assign new_n6532_ = new_n396_ & ~new_n6531_;
  assign new_n6533_ = new_n400_ & ~new_n6532_;
  assign new_n6534_ = new_n404_ & ~new_n6533_;
  assign new_n6535_ = new_n408_ & ~new_n6534_;
  assign new_n6536_ = new_n412_ & ~new_n6535_;
  assign new_n6537_ = new_n416_ & ~new_n6536_;
  assign new_n6538_ = new_n420_ & ~new_n6537_;
  assign new_n6539_ = new_n424_ & ~new_n6538_;
  assign new_n6540_ = new_n428_ & ~new_n6539_;
  assign new_n6541_ = new_n432_ & ~new_n6540_;
  assign new_n6542_ = new_n436_ & ~new_n6541_;
  assign new_n6543_ = new_n440_ & ~new_n6542_;
  assign new_n6544_ = new_n444_ & ~new_n6543_;
  assign new_n6545_ = new_n448_ & ~new_n6544_;
  assign new_n6546_ = new_n452_ & ~new_n6545_;
  assign new_n6547_ = new_n456_ & ~new_n6546_;
  assign new_n6548_ = new_n460_ & ~new_n6547_;
  assign new_n6549_ = new_n464_ & ~new_n6548_;
  assign new_n6550_ = new_n468_ & ~new_n6549_;
  assign new_n6551_ = new_n472_ & ~new_n6550_;
  assign new_n6552_ = new_n476_ & ~new_n6551_;
  assign new_n6553_ = new_n480_ & ~new_n6552_;
  assign new_n6554_ = new_n484_ & ~new_n6553_;
  assign new_n6555_ = new_n488_ & ~new_n6554_;
  assign new_n6556_ = new_n492_ & ~new_n6555_;
  assign new_n6557_ = new_n496_ & ~new_n6556_;
  assign new_n6558_ = new_n500_ & ~new_n6557_;
  assign new_n6559_ = new_n504_ & ~new_n6558_;
  assign new_n6560_ = new_n508_ & ~new_n6559_;
  assign new_n6561_ = new_n512_ & ~new_n6560_;
  assign new_n6562_ = new_n516_ & ~new_n6561_;
  assign new_n6563_ = new_n520_ & ~new_n6562_;
  assign new_n6564_ = new_n524_ & ~new_n6563_;
  assign new_n6565_ = new_n528_ & ~new_n6564_;
  assign new_n6566_ = new_n532_ & ~new_n6565_;
  assign new_n6567_ = new_n536_ & ~new_n6566_;
  assign new_n6568_ = new_n540_ & ~new_n6567_;
  assign new_n6569_ = new_n544_ & ~new_n6568_;
  assign new_n6570_ = \req[62]  & ~new_n546_;
  assign \grant[62]  = ~new_n6569_ & new_n6570_;
  assign new_n6572_ = new_n555_ & ~new_n890_;
  assign new_n6573_ = new_n560_ & ~new_n6572_;
  assign new_n6574_ = new_n564_ & ~new_n6573_;
  assign new_n6575_ = new_n568_ & ~new_n6574_;
  assign new_n6576_ = new_n572_ & ~new_n6575_;
  assign new_n6577_ = new_n576_ & ~new_n6576_;
  assign new_n6578_ = new_n580_ & ~new_n6577_;
  assign new_n6579_ = new_n584_ & ~new_n6578_;
  assign new_n6580_ = new_n588_ & ~new_n6579_;
  assign new_n6581_ = new_n592_ & ~new_n6580_;
  assign new_n6582_ = new_n596_ & ~new_n6581_;
  assign new_n6583_ = new_n600_ & ~new_n6582_;
  assign new_n6584_ = new_n604_ & ~new_n6583_;
  assign new_n6585_ = new_n608_ & ~new_n6584_;
  assign new_n6586_ = new_n612_ & ~new_n6585_;
  assign new_n6587_ = new_n616_ & ~new_n6586_;
  assign new_n6588_ = new_n620_ & ~new_n6587_;
  assign new_n6589_ = new_n624_ & ~new_n6588_;
  assign new_n6590_ = new_n628_ & ~new_n6589_;
  assign new_n6591_ = new_n632_ & ~new_n6590_;
  assign new_n6592_ = new_n636_ & ~new_n6591_;
  assign new_n6593_ = new_n640_ & ~new_n6592_;
  assign new_n6594_ = new_n644_ & ~new_n6593_;
  assign new_n6595_ = new_n648_ & ~new_n6594_;
  assign new_n6596_ = new_n652_ & ~new_n6595_;
  assign new_n6597_ = new_n656_ & ~new_n6596_;
  assign new_n6598_ = new_n660_ & ~new_n6597_;
  assign new_n6599_ = new_n664_ & ~new_n6598_;
  assign new_n6600_ = new_n668_ & ~new_n6599_;
  assign new_n6601_ = new_n672_ & ~new_n6600_;
  assign new_n6602_ = new_n676_ & ~new_n6601_;
  assign new_n6603_ = new_n680_ & ~new_n6602_;
  assign new_n6604_ = new_n684_ & ~new_n6603_;
  assign new_n6605_ = new_n688_ & ~new_n6604_;
  assign new_n6606_ = new_n692_ & ~new_n6605_;
  assign new_n6607_ = new_n696_ & ~new_n6606_;
  assign new_n6608_ = new_n700_ & ~new_n6607_;
  assign new_n6609_ = new_n704_ & ~new_n6608_;
  assign new_n6610_ = new_n708_ & ~new_n6609_;
  assign new_n6611_ = new_n712_ & ~new_n6610_;
  assign new_n6612_ = new_n716_ & ~new_n6611_;
  assign new_n6613_ = new_n720_ & ~new_n6612_;
  assign new_n6614_ = new_n1484_ & ~new_n6613_;
  assign new_n6615_ = new_n1486_ & ~new_n6614_;
  assign new_n6616_ = new_n1750_ & ~new_n6615_;
  assign new_n6617_ = new_n731_ & ~new_n6616_;
  assign new_n6618_ = new_n735_ & ~new_n6617_;
  assign new_n6619_ = new_n739_ & ~new_n6618_;
  assign new_n6620_ = new_n743_ & ~new_n6619_;
  assign new_n6621_ = new_n747_ & ~new_n6620_;
  assign new_n6622_ = new_n751_ & ~new_n6621_;
  assign new_n6623_ = new_n755_ & ~new_n6622_;
  assign new_n6624_ = new_n759_ & ~new_n6623_;
  assign new_n6625_ = new_n763_ & ~new_n6624_;
  assign new_n6626_ = new_n767_ & ~new_n6625_;
  assign new_n6627_ = new_n771_ & ~new_n6626_;
  assign new_n6628_ = new_n775_ & ~new_n6627_;
  assign new_n6629_ = new_n779_ & ~new_n6628_;
  assign new_n6630_ = new_n783_ & ~new_n6629_;
  assign new_n6631_ = new_n787_ & ~new_n6630_;
  assign new_n6632_ = new_n791_ & ~new_n6631_;
  assign new_n6633_ = new_n795_ & ~new_n6632_;
  assign new_n6634_ = new_n799_ & ~new_n6633_;
  assign new_n6635_ = new_n803_ & ~new_n6634_;
  assign new_n6636_ = new_n807_ & ~new_n6635_;
  assign new_n6637_ = new_n811_ & ~new_n6636_;
  assign new_n6638_ = new_n815_ & ~new_n6637_;
  assign new_n6639_ = new_n819_ & ~new_n6638_;
  assign new_n6640_ = new_n823_ & ~new_n6639_;
  assign new_n6641_ = new_n827_ & ~new_n6640_;
  assign new_n6642_ = new_n831_ & ~new_n6641_;
  assign new_n6643_ = new_n835_ & ~new_n6642_;
  assign new_n6644_ = new_n839_ & ~new_n6643_;
  assign new_n6645_ = new_n843_ & ~new_n6644_;
  assign new_n6646_ = new_n847_ & ~new_n6645_;
  assign new_n6647_ = new_n851_ & ~new_n6646_;
  assign new_n6648_ = new_n855_ & ~new_n6647_;
  assign new_n6649_ = new_n859_ & ~new_n6648_;
  assign new_n6650_ = new_n863_ & ~new_n6649_;
  assign new_n6651_ = new_n867_ & ~new_n6650_;
  assign new_n6652_ = new_n871_ & ~new_n6651_;
  assign new_n6653_ = new_n875_ & ~new_n6652_;
  assign new_n6654_ = new_n879_ & ~new_n6653_;
  assign new_n6655_ = new_n883_ & ~new_n6654_;
  assign new_n6656_ = \req[63]  & ~new_n885_;
  assign \grant[63]  = ~new_n6655_ & new_n6656_;
  assign new_n6658_ = new_n894_ & ~new_n1227_;
  assign new_n6659_ = new_n899_ & ~new_n6658_;
  assign new_n6660_ = new_n903_ & ~new_n6659_;
  assign new_n6661_ = new_n907_ & ~new_n6660_;
  assign new_n6662_ = new_n911_ & ~new_n6661_;
  assign new_n6663_ = new_n915_ & ~new_n6662_;
  assign new_n6664_ = new_n919_ & ~new_n6663_;
  assign new_n6665_ = new_n923_ & ~new_n6664_;
  assign new_n6666_ = new_n927_ & ~new_n6665_;
  assign new_n6667_ = new_n931_ & ~new_n6666_;
  assign new_n6668_ = new_n935_ & ~new_n6667_;
  assign new_n6669_ = new_n939_ & ~new_n6668_;
  assign new_n6670_ = new_n943_ & ~new_n6669_;
  assign new_n6671_ = new_n947_ & ~new_n6670_;
  assign new_n6672_ = new_n951_ & ~new_n6671_;
  assign new_n6673_ = new_n955_ & ~new_n6672_;
  assign new_n6674_ = new_n959_ & ~new_n6673_;
  assign new_n6675_ = new_n963_ & ~new_n6674_;
  assign new_n6676_ = new_n967_ & ~new_n6675_;
  assign new_n6677_ = new_n971_ & ~new_n6676_;
  assign new_n6678_ = new_n975_ & ~new_n6677_;
  assign new_n6679_ = new_n979_ & ~new_n6678_;
  assign new_n6680_ = new_n983_ & ~new_n6679_;
  assign new_n6681_ = new_n987_ & ~new_n6680_;
  assign new_n6682_ = new_n991_ & ~new_n6681_;
  assign new_n6683_ = new_n995_ & ~new_n6682_;
  assign new_n6684_ = new_n999_ & ~new_n6683_;
  assign new_n6685_ = new_n1003_ & ~new_n6684_;
  assign new_n6686_ = new_n1007_ & ~new_n6685_;
  assign new_n6687_ = new_n1011_ & ~new_n6686_;
  assign new_n6688_ = new_n1015_ & ~new_n6687_;
  assign new_n6689_ = new_n1019_ & ~new_n6688_;
  assign new_n6690_ = new_n1023_ & ~new_n6689_;
  assign new_n6691_ = new_n1027_ & ~new_n6690_;
  assign new_n6692_ = new_n1031_ & ~new_n6691_;
  assign new_n6693_ = new_n1035_ & ~new_n6692_;
  assign new_n6694_ = new_n1039_ & ~new_n6693_;
  assign new_n6695_ = new_n1043_ & ~new_n6694_;
  assign new_n6696_ = new_n1047_ & ~new_n6695_;
  assign new_n6697_ = new_n1051_ & ~new_n6696_;
  assign new_n6698_ = new_n1055_ & ~new_n6697_;
  assign new_n6699_ = new_n1059_ & ~new_n6698_;
  assign new_n6700_ = new_n1574_ & ~new_n6699_;
  assign new_n6701_ = new_n1576_ & ~new_n6700_;
  assign new_n6702_ = new_n1837_ & ~new_n6701_;
  assign new_n6703_ = new_n1068_ & ~new_n6702_;
  assign new_n6704_ = new_n1072_ & ~new_n6703_;
  assign new_n6705_ = new_n1076_ & ~new_n6704_;
  assign new_n6706_ = new_n1080_ & ~new_n6705_;
  assign new_n6707_ = new_n1084_ & ~new_n6706_;
  assign new_n6708_ = new_n1088_ & ~new_n6707_;
  assign new_n6709_ = new_n1092_ & ~new_n6708_;
  assign new_n6710_ = new_n1096_ & ~new_n6709_;
  assign new_n6711_ = new_n1100_ & ~new_n6710_;
  assign new_n6712_ = new_n1104_ & ~new_n6711_;
  assign new_n6713_ = new_n1108_ & ~new_n6712_;
  assign new_n6714_ = new_n1112_ & ~new_n6713_;
  assign new_n6715_ = new_n1116_ & ~new_n6714_;
  assign new_n6716_ = new_n1120_ & ~new_n6715_;
  assign new_n6717_ = new_n1124_ & ~new_n6716_;
  assign new_n6718_ = new_n1128_ & ~new_n6717_;
  assign new_n6719_ = new_n1132_ & ~new_n6718_;
  assign new_n6720_ = new_n1136_ & ~new_n6719_;
  assign new_n6721_ = new_n1140_ & ~new_n6720_;
  assign new_n6722_ = new_n1144_ & ~new_n6721_;
  assign new_n6723_ = new_n1148_ & ~new_n6722_;
  assign new_n6724_ = new_n1152_ & ~new_n6723_;
  assign new_n6725_ = new_n1156_ & ~new_n6724_;
  assign new_n6726_ = new_n1160_ & ~new_n6725_;
  assign new_n6727_ = new_n1164_ & ~new_n6726_;
  assign new_n6728_ = new_n1168_ & ~new_n6727_;
  assign new_n6729_ = new_n1172_ & ~new_n6728_;
  assign new_n6730_ = new_n1176_ & ~new_n6729_;
  assign new_n6731_ = new_n1180_ & ~new_n6730_;
  assign new_n6732_ = new_n1184_ & ~new_n6731_;
  assign new_n6733_ = new_n1188_ & ~new_n6732_;
  assign new_n6734_ = new_n1192_ & ~new_n6733_;
  assign new_n6735_ = new_n1196_ & ~new_n6734_;
  assign new_n6736_ = new_n1200_ & ~new_n6735_;
  assign new_n6737_ = new_n1204_ & ~new_n6736_;
  assign new_n6738_ = new_n1208_ & ~new_n6737_;
  assign new_n6739_ = new_n1212_ & ~new_n6738_;
  assign new_n6740_ = new_n1216_ & ~new_n6739_;
  assign new_n6741_ = new_n1220_ & ~new_n6740_;
  assign new_n6742_ = \req[64]  & ~new_n1222_;
  assign \grant[64]  = ~new_n6741_ & new_n6742_;
  assign new_n6744_ = ~new_n559_ & new_n1231_;
  assign new_n6745_ = new_n1236_ & ~new_n6744_;
  assign new_n6746_ = new_n1240_ & ~new_n6745_;
  assign new_n6747_ = new_n1244_ & ~new_n6746_;
  assign new_n6748_ = new_n1248_ & ~new_n6747_;
  assign new_n6749_ = new_n1252_ & ~new_n6748_;
  assign new_n6750_ = new_n1256_ & ~new_n6749_;
  assign new_n6751_ = new_n1260_ & ~new_n6750_;
  assign new_n6752_ = new_n1264_ & ~new_n6751_;
  assign new_n6753_ = new_n1268_ & ~new_n6752_;
  assign new_n6754_ = new_n1272_ & ~new_n6753_;
  assign new_n6755_ = new_n1276_ & ~new_n6754_;
  assign new_n6756_ = new_n1280_ & ~new_n6755_;
  assign new_n6757_ = new_n1284_ & ~new_n6756_;
  assign new_n6758_ = new_n1288_ & ~new_n6757_;
  assign new_n6759_ = new_n1292_ & ~new_n6758_;
  assign new_n6760_ = new_n1296_ & ~new_n6759_;
  assign new_n6761_ = new_n1300_ & ~new_n6760_;
  assign new_n6762_ = new_n1304_ & ~new_n6761_;
  assign new_n6763_ = new_n1308_ & ~new_n6762_;
  assign new_n6764_ = new_n1312_ & ~new_n6763_;
  assign new_n6765_ = new_n1316_ & ~new_n6764_;
  assign new_n6766_ = new_n1320_ & ~new_n6765_;
  assign new_n6767_ = new_n1324_ & ~new_n6766_;
  assign new_n6768_ = new_n1328_ & ~new_n6767_;
  assign new_n6769_ = new_n1332_ & ~new_n6768_;
  assign new_n6770_ = new_n1336_ & ~new_n6769_;
  assign new_n6771_ = new_n1340_ & ~new_n6770_;
  assign new_n6772_ = new_n1344_ & ~new_n6771_;
  assign new_n6773_ = new_n1348_ & ~new_n6772_;
  assign new_n6774_ = new_n1352_ & ~new_n6773_;
  assign new_n6775_ = new_n1356_ & ~new_n6774_;
  assign new_n6776_ = new_n1360_ & ~new_n6775_;
  assign new_n6777_ = new_n1364_ & ~new_n6776_;
  assign new_n6778_ = new_n1368_ & ~new_n6777_;
  assign new_n6779_ = new_n1372_ & ~new_n6778_;
  assign new_n6780_ = new_n1376_ & ~new_n6779_;
  assign new_n6781_ = new_n1380_ & ~new_n6780_;
  assign new_n6782_ = new_n1384_ & ~new_n6781_;
  assign new_n6783_ = new_n1388_ & ~new_n6782_;
  assign new_n6784_ = new_n1392_ & ~new_n6783_;
  assign new_n6785_ = new_n1396_ & ~new_n6784_;
  assign new_n6786_ = new_n1663_ & ~new_n6785_;
  assign new_n6787_ = new_n392_ & ~new_n6786_;
  assign new_n6788_ = new_n396_ & ~new_n6787_;
  assign new_n6789_ = new_n400_ & ~new_n6788_;
  assign new_n6790_ = new_n404_ & ~new_n6789_;
  assign new_n6791_ = new_n408_ & ~new_n6790_;
  assign new_n6792_ = new_n412_ & ~new_n6791_;
  assign new_n6793_ = new_n416_ & ~new_n6792_;
  assign new_n6794_ = new_n420_ & ~new_n6793_;
  assign new_n6795_ = new_n424_ & ~new_n6794_;
  assign new_n6796_ = new_n428_ & ~new_n6795_;
  assign new_n6797_ = new_n432_ & ~new_n6796_;
  assign new_n6798_ = new_n436_ & ~new_n6797_;
  assign new_n6799_ = new_n440_ & ~new_n6798_;
  assign new_n6800_ = new_n444_ & ~new_n6799_;
  assign new_n6801_ = new_n448_ & ~new_n6800_;
  assign new_n6802_ = new_n452_ & ~new_n6801_;
  assign new_n6803_ = new_n456_ & ~new_n6802_;
  assign new_n6804_ = new_n460_ & ~new_n6803_;
  assign new_n6805_ = new_n464_ & ~new_n6804_;
  assign new_n6806_ = new_n468_ & ~new_n6805_;
  assign new_n6807_ = new_n472_ & ~new_n6806_;
  assign new_n6808_ = new_n476_ & ~new_n6807_;
  assign new_n6809_ = new_n480_ & ~new_n6808_;
  assign new_n6810_ = new_n484_ & ~new_n6809_;
  assign new_n6811_ = new_n488_ & ~new_n6810_;
  assign new_n6812_ = new_n492_ & ~new_n6811_;
  assign new_n6813_ = new_n496_ & ~new_n6812_;
  assign new_n6814_ = new_n500_ & ~new_n6813_;
  assign new_n6815_ = new_n504_ & ~new_n6814_;
  assign new_n6816_ = new_n508_ & ~new_n6815_;
  assign new_n6817_ = new_n512_ & ~new_n6816_;
  assign new_n6818_ = new_n516_ & ~new_n6817_;
  assign new_n6819_ = new_n520_ & ~new_n6818_;
  assign new_n6820_ = new_n524_ & ~new_n6819_;
  assign new_n6821_ = new_n528_ & ~new_n6820_;
  assign new_n6822_ = new_n532_ & ~new_n6821_;
  assign new_n6823_ = new_n536_ & ~new_n6822_;
  assign new_n6824_ = new_n540_ & ~new_n6823_;
  assign new_n6825_ = new_n544_ & ~new_n6824_;
  assign new_n6826_ = new_n548_ & ~new_n6825_;
  assign new_n6827_ = new_n552_ & ~new_n6826_;
  assign new_n6828_ = \req[65]  & ~new_n554_;
  assign \grant[65]  = ~new_n6827_ & new_n6828_;
  assign new_n6830_ = new_n563_ & ~new_n898_;
  assign new_n6831_ = new_n568_ & ~new_n6830_;
  assign new_n6832_ = new_n572_ & ~new_n6831_;
  assign new_n6833_ = new_n576_ & ~new_n6832_;
  assign new_n6834_ = new_n580_ & ~new_n6833_;
  assign new_n6835_ = new_n584_ & ~new_n6834_;
  assign new_n6836_ = new_n588_ & ~new_n6835_;
  assign new_n6837_ = new_n592_ & ~new_n6836_;
  assign new_n6838_ = new_n596_ & ~new_n6837_;
  assign new_n6839_ = new_n600_ & ~new_n6838_;
  assign new_n6840_ = new_n604_ & ~new_n6839_;
  assign new_n6841_ = new_n608_ & ~new_n6840_;
  assign new_n6842_ = new_n612_ & ~new_n6841_;
  assign new_n6843_ = new_n616_ & ~new_n6842_;
  assign new_n6844_ = new_n620_ & ~new_n6843_;
  assign new_n6845_ = new_n624_ & ~new_n6844_;
  assign new_n6846_ = new_n628_ & ~new_n6845_;
  assign new_n6847_ = new_n632_ & ~new_n6846_;
  assign new_n6848_ = new_n636_ & ~new_n6847_;
  assign new_n6849_ = new_n640_ & ~new_n6848_;
  assign new_n6850_ = new_n644_ & ~new_n6849_;
  assign new_n6851_ = new_n648_ & ~new_n6850_;
  assign new_n6852_ = new_n652_ & ~new_n6851_;
  assign new_n6853_ = new_n656_ & ~new_n6852_;
  assign new_n6854_ = new_n660_ & ~new_n6853_;
  assign new_n6855_ = new_n664_ & ~new_n6854_;
  assign new_n6856_ = new_n668_ & ~new_n6855_;
  assign new_n6857_ = new_n672_ & ~new_n6856_;
  assign new_n6858_ = new_n676_ & ~new_n6857_;
  assign new_n6859_ = new_n680_ & ~new_n6858_;
  assign new_n6860_ = new_n684_ & ~new_n6859_;
  assign new_n6861_ = new_n688_ & ~new_n6860_;
  assign new_n6862_ = new_n692_ & ~new_n6861_;
  assign new_n6863_ = new_n696_ & ~new_n6862_;
  assign new_n6864_ = new_n700_ & ~new_n6863_;
  assign new_n6865_ = new_n704_ & ~new_n6864_;
  assign new_n6866_ = new_n708_ & ~new_n6865_;
  assign new_n6867_ = new_n712_ & ~new_n6866_;
  assign new_n6868_ = new_n716_ & ~new_n6867_;
  assign new_n6869_ = new_n720_ & ~new_n6868_;
  assign new_n6870_ = new_n1484_ & ~new_n6869_;
  assign new_n6871_ = new_n1486_ & ~new_n6870_;
  assign new_n6872_ = new_n1750_ & ~new_n6871_;
  assign new_n6873_ = new_n731_ & ~new_n6872_;
  assign new_n6874_ = new_n735_ & ~new_n6873_;
  assign new_n6875_ = new_n739_ & ~new_n6874_;
  assign new_n6876_ = new_n743_ & ~new_n6875_;
  assign new_n6877_ = new_n747_ & ~new_n6876_;
  assign new_n6878_ = new_n751_ & ~new_n6877_;
  assign new_n6879_ = new_n755_ & ~new_n6878_;
  assign new_n6880_ = new_n759_ & ~new_n6879_;
  assign new_n6881_ = new_n763_ & ~new_n6880_;
  assign new_n6882_ = new_n767_ & ~new_n6881_;
  assign new_n6883_ = new_n771_ & ~new_n6882_;
  assign new_n6884_ = new_n775_ & ~new_n6883_;
  assign new_n6885_ = new_n779_ & ~new_n6884_;
  assign new_n6886_ = new_n783_ & ~new_n6885_;
  assign new_n6887_ = new_n787_ & ~new_n6886_;
  assign new_n6888_ = new_n791_ & ~new_n6887_;
  assign new_n6889_ = new_n795_ & ~new_n6888_;
  assign new_n6890_ = new_n799_ & ~new_n6889_;
  assign new_n6891_ = new_n803_ & ~new_n6890_;
  assign new_n6892_ = new_n807_ & ~new_n6891_;
  assign new_n6893_ = new_n811_ & ~new_n6892_;
  assign new_n6894_ = new_n815_ & ~new_n6893_;
  assign new_n6895_ = new_n819_ & ~new_n6894_;
  assign new_n6896_ = new_n823_ & ~new_n6895_;
  assign new_n6897_ = new_n827_ & ~new_n6896_;
  assign new_n6898_ = new_n831_ & ~new_n6897_;
  assign new_n6899_ = new_n835_ & ~new_n6898_;
  assign new_n6900_ = new_n839_ & ~new_n6899_;
  assign new_n6901_ = new_n843_ & ~new_n6900_;
  assign new_n6902_ = new_n847_ & ~new_n6901_;
  assign new_n6903_ = new_n851_ & ~new_n6902_;
  assign new_n6904_ = new_n855_ & ~new_n6903_;
  assign new_n6905_ = new_n859_ & ~new_n6904_;
  assign new_n6906_ = new_n863_ & ~new_n6905_;
  assign new_n6907_ = new_n867_ & ~new_n6906_;
  assign new_n6908_ = new_n871_ & ~new_n6907_;
  assign new_n6909_ = new_n875_ & ~new_n6908_;
  assign new_n6910_ = new_n879_ & ~new_n6909_;
  assign new_n6911_ = new_n883_ & ~new_n6910_;
  assign new_n6912_ = new_n887_ & ~new_n6911_;
  assign new_n6913_ = new_n891_ & ~new_n6912_;
  assign new_n6914_ = \req[66]  & ~new_n893_;
  assign \grant[66]  = ~new_n6913_ & new_n6914_;
  assign new_n6916_ = new_n902_ & ~new_n1235_;
  assign new_n6917_ = new_n907_ & ~new_n6916_;
  assign new_n6918_ = new_n911_ & ~new_n6917_;
  assign new_n6919_ = new_n915_ & ~new_n6918_;
  assign new_n6920_ = new_n919_ & ~new_n6919_;
  assign new_n6921_ = new_n923_ & ~new_n6920_;
  assign new_n6922_ = new_n927_ & ~new_n6921_;
  assign new_n6923_ = new_n931_ & ~new_n6922_;
  assign new_n6924_ = new_n935_ & ~new_n6923_;
  assign new_n6925_ = new_n939_ & ~new_n6924_;
  assign new_n6926_ = new_n943_ & ~new_n6925_;
  assign new_n6927_ = new_n947_ & ~new_n6926_;
  assign new_n6928_ = new_n951_ & ~new_n6927_;
  assign new_n6929_ = new_n955_ & ~new_n6928_;
  assign new_n6930_ = new_n959_ & ~new_n6929_;
  assign new_n6931_ = new_n963_ & ~new_n6930_;
  assign new_n6932_ = new_n967_ & ~new_n6931_;
  assign new_n6933_ = new_n971_ & ~new_n6932_;
  assign new_n6934_ = new_n975_ & ~new_n6933_;
  assign new_n6935_ = new_n979_ & ~new_n6934_;
  assign new_n6936_ = new_n983_ & ~new_n6935_;
  assign new_n6937_ = new_n987_ & ~new_n6936_;
  assign new_n6938_ = new_n991_ & ~new_n6937_;
  assign new_n6939_ = new_n995_ & ~new_n6938_;
  assign new_n6940_ = new_n999_ & ~new_n6939_;
  assign new_n6941_ = new_n1003_ & ~new_n6940_;
  assign new_n6942_ = new_n1007_ & ~new_n6941_;
  assign new_n6943_ = new_n1011_ & ~new_n6942_;
  assign new_n6944_ = new_n1015_ & ~new_n6943_;
  assign new_n6945_ = new_n1019_ & ~new_n6944_;
  assign new_n6946_ = new_n1023_ & ~new_n6945_;
  assign new_n6947_ = new_n1027_ & ~new_n6946_;
  assign new_n6948_ = new_n1031_ & ~new_n6947_;
  assign new_n6949_ = new_n1035_ & ~new_n6948_;
  assign new_n6950_ = new_n1039_ & ~new_n6949_;
  assign new_n6951_ = new_n1043_ & ~new_n6950_;
  assign new_n6952_ = new_n1047_ & ~new_n6951_;
  assign new_n6953_ = new_n1051_ & ~new_n6952_;
  assign new_n6954_ = new_n1055_ & ~new_n6953_;
  assign new_n6955_ = new_n1059_ & ~new_n6954_;
  assign new_n6956_ = new_n1574_ & ~new_n6955_;
  assign new_n6957_ = new_n1576_ & ~new_n6956_;
  assign new_n6958_ = new_n1837_ & ~new_n6957_;
  assign new_n6959_ = new_n1068_ & ~new_n6958_;
  assign new_n6960_ = new_n1072_ & ~new_n6959_;
  assign new_n6961_ = new_n1076_ & ~new_n6960_;
  assign new_n6962_ = new_n1080_ & ~new_n6961_;
  assign new_n6963_ = new_n1084_ & ~new_n6962_;
  assign new_n6964_ = new_n1088_ & ~new_n6963_;
  assign new_n6965_ = new_n1092_ & ~new_n6964_;
  assign new_n6966_ = new_n1096_ & ~new_n6965_;
  assign new_n6967_ = new_n1100_ & ~new_n6966_;
  assign new_n6968_ = new_n1104_ & ~new_n6967_;
  assign new_n6969_ = new_n1108_ & ~new_n6968_;
  assign new_n6970_ = new_n1112_ & ~new_n6969_;
  assign new_n6971_ = new_n1116_ & ~new_n6970_;
  assign new_n6972_ = new_n1120_ & ~new_n6971_;
  assign new_n6973_ = new_n1124_ & ~new_n6972_;
  assign new_n6974_ = new_n1128_ & ~new_n6973_;
  assign new_n6975_ = new_n1132_ & ~new_n6974_;
  assign new_n6976_ = new_n1136_ & ~new_n6975_;
  assign new_n6977_ = new_n1140_ & ~new_n6976_;
  assign new_n6978_ = new_n1144_ & ~new_n6977_;
  assign new_n6979_ = new_n1148_ & ~new_n6978_;
  assign new_n6980_ = new_n1152_ & ~new_n6979_;
  assign new_n6981_ = new_n1156_ & ~new_n6980_;
  assign new_n6982_ = new_n1160_ & ~new_n6981_;
  assign new_n6983_ = new_n1164_ & ~new_n6982_;
  assign new_n6984_ = new_n1168_ & ~new_n6983_;
  assign new_n6985_ = new_n1172_ & ~new_n6984_;
  assign new_n6986_ = new_n1176_ & ~new_n6985_;
  assign new_n6987_ = new_n1180_ & ~new_n6986_;
  assign new_n6988_ = new_n1184_ & ~new_n6987_;
  assign new_n6989_ = new_n1188_ & ~new_n6988_;
  assign new_n6990_ = new_n1192_ & ~new_n6989_;
  assign new_n6991_ = new_n1196_ & ~new_n6990_;
  assign new_n6992_ = new_n1200_ & ~new_n6991_;
  assign new_n6993_ = new_n1204_ & ~new_n6992_;
  assign new_n6994_ = new_n1208_ & ~new_n6993_;
  assign new_n6995_ = new_n1212_ & ~new_n6994_;
  assign new_n6996_ = new_n1216_ & ~new_n6995_;
  assign new_n6997_ = new_n1220_ & ~new_n6996_;
  assign new_n6998_ = new_n1224_ & ~new_n6997_;
  assign new_n6999_ = new_n1228_ & ~new_n6998_;
  assign new_n7000_ = \req[67]  & ~new_n1230_;
  assign \grant[67]  = ~new_n6999_ & new_n7000_;
  assign new_n7002_ = ~new_n567_ & new_n1239_;
  assign new_n7003_ = new_n1244_ & ~new_n7002_;
  assign new_n7004_ = new_n1248_ & ~new_n7003_;
  assign new_n7005_ = new_n1252_ & ~new_n7004_;
  assign new_n7006_ = new_n1256_ & ~new_n7005_;
  assign new_n7007_ = new_n1260_ & ~new_n7006_;
  assign new_n7008_ = new_n1264_ & ~new_n7007_;
  assign new_n7009_ = new_n1268_ & ~new_n7008_;
  assign new_n7010_ = new_n1272_ & ~new_n7009_;
  assign new_n7011_ = new_n1276_ & ~new_n7010_;
  assign new_n7012_ = new_n1280_ & ~new_n7011_;
  assign new_n7013_ = new_n1284_ & ~new_n7012_;
  assign new_n7014_ = new_n1288_ & ~new_n7013_;
  assign new_n7015_ = new_n1292_ & ~new_n7014_;
  assign new_n7016_ = new_n1296_ & ~new_n7015_;
  assign new_n7017_ = new_n1300_ & ~new_n7016_;
  assign new_n7018_ = new_n1304_ & ~new_n7017_;
  assign new_n7019_ = new_n1308_ & ~new_n7018_;
  assign new_n7020_ = new_n1312_ & ~new_n7019_;
  assign new_n7021_ = new_n1316_ & ~new_n7020_;
  assign new_n7022_ = new_n1320_ & ~new_n7021_;
  assign new_n7023_ = new_n1324_ & ~new_n7022_;
  assign new_n7024_ = new_n1328_ & ~new_n7023_;
  assign new_n7025_ = new_n1332_ & ~new_n7024_;
  assign new_n7026_ = new_n1336_ & ~new_n7025_;
  assign new_n7027_ = new_n1340_ & ~new_n7026_;
  assign new_n7028_ = new_n1344_ & ~new_n7027_;
  assign new_n7029_ = new_n1348_ & ~new_n7028_;
  assign new_n7030_ = new_n1352_ & ~new_n7029_;
  assign new_n7031_ = new_n1356_ & ~new_n7030_;
  assign new_n7032_ = new_n1360_ & ~new_n7031_;
  assign new_n7033_ = new_n1364_ & ~new_n7032_;
  assign new_n7034_ = new_n1368_ & ~new_n7033_;
  assign new_n7035_ = new_n1372_ & ~new_n7034_;
  assign new_n7036_ = new_n1376_ & ~new_n7035_;
  assign new_n7037_ = new_n1380_ & ~new_n7036_;
  assign new_n7038_ = new_n1384_ & ~new_n7037_;
  assign new_n7039_ = new_n1388_ & ~new_n7038_;
  assign new_n7040_ = new_n1392_ & ~new_n7039_;
  assign new_n7041_ = new_n1396_ & ~new_n7040_;
  assign new_n7042_ = new_n1663_ & ~new_n7041_;
  assign new_n7043_ = new_n392_ & ~new_n7042_;
  assign new_n7044_ = new_n396_ & ~new_n7043_;
  assign new_n7045_ = new_n400_ & ~new_n7044_;
  assign new_n7046_ = new_n404_ & ~new_n7045_;
  assign new_n7047_ = new_n408_ & ~new_n7046_;
  assign new_n7048_ = new_n412_ & ~new_n7047_;
  assign new_n7049_ = new_n416_ & ~new_n7048_;
  assign new_n7050_ = new_n420_ & ~new_n7049_;
  assign new_n7051_ = new_n424_ & ~new_n7050_;
  assign new_n7052_ = new_n428_ & ~new_n7051_;
  assign new_n7053_ = new_n432_ & ~new_n7052_;
  assign new_n7054_ = new_n436_ & ~new_n7053_;
  assign new_n7055_ = new_n440_ & ~new_n7054_;
  assign new_n7056_ = new_n444_ & ~new_n7055_;
  assign new_n7057_ = new_n448_ & ~new_n7056_;
  assign new_n7058_ = new_n452_ & ~new_n7057_;
  assign new_n7059_ = new_n456_ & ~new_n7058_;
  assign new_n7060_ = new_n460_ & ~new_n7059_;
  assign new_n7061_ = new_n464_ & ~new_n7060_;
  assign new_n7062_ = new_n468_ & ~new_n7061_;
  assign new_n7063_ = new_n472_ & ~new_n7062_;
  assign new_n7064_ = new_n476_ & ~new_n7063_;
  assign new_n7065_ = new_n480_ & ~new_n7064_;
  assign new_n7066_ = new_n484_ & ~new_n7065_;
  assign new_n7067_ = new_n488_ & ~new_n7066_;
  assign new_n7068_ = new_n492_ & ~new_n7067_;
  assign new_n7069_ = new_n496_ & ~new_n7068_;
  assign new_n7070_ = new_n500_ & ~new_n7069_;
  assign new_n7071_ = new_n504_ & ~new_n7070_;
  assign new_n7072_ = new_n508_ & ~new_n7071_;
  assign new_n7073_ = new_n512_ & ~new_n7072_;
  assign new_n7074_ = new_n516_ & ~new_n7073_;
  assign new_n7075_ = new_n520_ & ~new_n7074_;
  assign new_n7076_ = new_n524_ & ~new_n7075_;
  assign new_n7077_ = new_n528_ & ~new_n7076_;
  assign new_n7078_ = new_n532_ & ~new_n7077_;
  assign new_n7079_ = new_n536_ & ~new_n7078_;
  assign new_n7080_ = new_n540_ & ~new_n7079_;
  assign new_n7081_ = new_n544_ & ~new_n7080_;
  assign new_n7082_ = new_n548_ & ~new_n7081_;
  assign new_n7083_ = new_n552_ & ~new_n7082_;
  assign new_n7084_ = new_n556_ & ~new_n7083_;
  assign new_n7085_ = new_n560_ & ~new_n7084_;
  assign new_n7086_ = \req[68]  & ~new_n562_;
  assign \grant[68]  = ~new_n7085_ & new_n7086_;
  assign new_n7088_ = new_n571_ & ~new_n906_;
  assign new_n7089_ = new_n576_ & ~new_n7088_;
  assign new_n7090_ = new_n580_ & ~new_n7089_;
  assign new_n7091_ = new_n584_ & ~new_n7090_;
  assign new_n7092_ = new_n588_ & ~new_n7091_;
  assign new_n7093_ = new_n592_ & ~new_n7092_;
  assign new_n7094_ = new_n596_ & ~new_n7093_;
  assign new_n7095_ = new_n600_ & ~new_n7094_;
  assign new_n7096_ = new_n604_ & ~new_n7095_;
  assign new_n7097_ = new_n608_ & ~new_n7096_;
  assign new_n7098_ = new_n612_ & ~new_n7097_;
  assign new_n7099_ = new_n616_ & ~new_n7098_;
  assign new_n7100_ = new_n620_ & ~new_n7099_;
  assign new_n7101_ = new_n624_ & ~new_n7100_;
  assign new_n7102_ = new_n628_ & ~new_n7101_;
  assign new_n7103_ = new_n632_ & ~new_n7102_;
  assign new_n7104_ = new_n636_ & ~new_n7103_;
  assign new_n7105_ = new_n640_ & ~new_n7104_;
  assign new_n7106_ = new_n644_ & ~new_n7105_;
  assign new_n7107_ = new_n648_ & ~new_n7106_;
  assign new_n7108_ = new_n652_ & ~new_n7107_;
  assign new_n7109_ = new_n656_ & ~new_n7108_;
  assign new_n7110_ = new_n660_ & ~new_n7109_;
  assign new_n7111_ = new_n664_ & ~new_n7110_;
  assign new_n7112_ = new_n668_ & ~new_n7111_;
  assign new_n7113_ = new_n672_ & ~new_n7112_;
  assign new_n7114_ = new_n676_ & ~new_n7113_;
  assign new_n7115_ = new_n680_ & ~new_n7114_;
  assign new_n7116_ = new_n684_ & ~new_n7115_;
  assign new_n7117_ = new_n688_ & ~new_n7116_;
  assign new_n7118_ = new_n692_ & ~new_n7117_;
  assign new_n7119_ = new_n696_ & ~new_n7118_;
  assign new_n7120_ = new_n700_ & ~new_n7119_;
  assign new_n7121_ = new_n704_ & ~new_n7120_;
  assign new_n7122_ = new_n708_ & ~new_n7121_;
  assign new_n7123_ = new_n712_ & ~new_n7122_;
  assign new_n7124_ = new_n716_ & ~new_n7123_;
  assign new_n7125_ = new_n720_ & ~new_n7124_;
  assign new_n7126_ = new_n1484_ & ~new_n7125_;
  assign new_n7127_ = new_n1486_ & ~new_n7126_;
  assign new_n7128_ = new_n1750_ & ~new_n7127_;
  assign new_n7129_ = new_n731_ & ~new_n7128_;
  assign new_n7130_ = new_n735_ & ~new_n7129_;
  assign new_n7131_ = new_n739_ & ~new_n7130_;
  assign new_n7132_ = new_n743_ & ~new_n7131_;
  assign new_n7133_ = new_n747_ & ~new_n7132_;
  assign new_n7134_ = new_n751_ & ~new_n7133_;
  assign new_n7135_ = new_n755_ & ~new_n7134_;
  assign new_n7136_ = new_n759_ & ~new_n7135_;
  assign new_n7137_ = new_n763_ & ~new_n7136_;
  assign new_n7138_ = new_n767_ & ~new_n7137_;
  assign new_n7139_ = new_n771_ & ~new_n7138_;
  assign new_n7140_ = new_n775_ & ~new_n7139_;
  assign new_n7141_ = new_n779_ & ~new_n7140_;
  assign new_n7142_ = new_n783_ & ~new_n7141_;
  assign new_n7143_ = new_n787_ & ~new_n7142_;
  assign new_n7144_ = new_n791_ & ~new_n7143_;
  assign new_n7145_ = new_n795_ & ~new_n7144_;
  assign new_n7146_ = new_n799_ & ~new_n7145_;
  assign new_n7147_ = new_n803_ & ~new_n7146_;
  assign new_n7148_ = new_n807_ & ~new_n7147_;
  assign new_n7149_ = new_n811_ & ~new_n7148_;
  assign new_n7150_ = new_n815_ & ~new_n7149_;
  assign new_n7151_ = new_n819_ & ~new_n7150_;
  assign new_n7152_ = new_n823_ & ~new_n7151_;
  assign new_n7153_ = new_n827_ & ~new_n7152_;
  assign new_n7154_ = new_n831_ & ~new_n7153_;
  assign new_n7155_ = new_n835_ & ~new_n7154_;
  assign new_n7156_ = new_n839_ & ~new_n7155_;
  assign new_n7157_ = new_n843_ & ~new_n7156_;
  assign new_n7158_ = new_n847_ & ~new_n7157_;
  assign new_n7159_ = new_n851_ & ~new_n7158_;
  assign new_n7160_ = new_n855_ & ~new_n7159_;
  assign new_n7161_ = new_n859_ & ~new_n7160_;
  assign new_n7162_ = new_n863_ & ~new_n7161_;
  assign new_n7163_ = new_n867_ & ~new_n7162_;
  assign new_n7164_ = new_n871_ & ~new_n7163_;
  assign new_n7165_ = new_n875_ & ~new_n7164_;
  assign new_n7166_ = new_n879_ & ~new_n7165_;
  assign new_n7167_ = new_n883_ & ~new_n7166_;
  assign new_n7168_ = new_n887_ & ~new_n7167_;
  assign new_n7169_ = new_n891_ & ~new_n7168_;
  assign new_n7170_ = new_n895_ & ~new_n7169_;
  assign new_n7171_ = new_n899_ & ~new_n7170_;
  assign new_n7172_ = \req[69]  & ~new_n901_;
  assign \grant[69]  = ~new_n7171_ & new_n7172_;
  assign new_n7174_ = new_n910_ & ~new_n1243_;
  assign new_n7175_ = new_n915_ & ~new_n7174_;
  assign new_n7176_ = new_n919_ & ~new_n7175_;
  assign new_n7177_ = new_n923_ & ~new_n7176_;
  assign new_n7178_ = new_n927_ & ~new_n7177_;
  assign new_n7179_ = new_n931_ & ~new_n7178_;
  assign new_n7180_ = new_n935_ & ~new_n7179_;
  assign new_n7181_ = new_n939_ & ~new_n7180_;
  assign new_n7182_ = new_n943_ & ~new_n7181_;
  assign new_n7183_ = new_n947_ & ~new_n7182_;
  assign new_n7184_ = new_n951_ & ~new_n7183_;
  assign new_n7185_ = new_n955_ & ~new_n7184_;
  assign new_n7186_ = new_n959_ & ~new_n7185_;
  assign new_n7187_ = new_n963_ & ~new_n7186_;
  assign new_n7188_ = new_n967_ & ~new_n7187_;
  assign new_n7189_ = new_n971_ & ~new_n7188_;
  assign new_n7190_ = new_n975_ & ~new_n7189_;
  assign new_n7191_ = new_n979_ & ~new_n7190_;
  assign new_n7192_ = new_n983_ & ~new_n7191_;
  assign new_n7193_ = new_n987_ & ~new_n7192_;
  assign new_n7194_ = new_n991_ & ~new_n7193_;
  assign new_n7195_ = new_n995_ & ~new_n7194_;
  assign new_n7196_ = new_n999_ & ~new_n7195_;
  assign new_n7197_ = new_n1003_ & ~new_n7196_;
  assign new_n7198_ = new_n1007_ & ~new_n7197_;
  assign new_n7199_ = new_n1011_ & ~new_n7198_;
  assign new_n7200_ = new_n1015_ & ~new_n7199_;
  assign new_n7201_ = new_n1019_ & ~new_n7200_;
  assign new_n7202_ = new_n1023_ & ~new_n7201_;
  assign new_n7203_ = new_n1027_ & ~new_n7202_;
  assign new_n7204_ = new_n1031_ & ~new_n7203_;
  assign new_n7205_ = new_n1035_ & ~new_n7204_;
  assign new_n7206_ = new_n1039_ & ~new_n7205_;
  assign new_n7207_ = new_n1043_ & ~new_n7206_;
  assign new_n7208_ = new_n1047_ & ~new_n7207_;
  assign new_n7209_ = new_n1051_ & ~new_n7208_;
  assign new_n7210_ = new_n1055_ & ~new_n7209_;
  assign new_n7211_ = new_n1059_ & ~new_n7210_;
  assign new_n7212_ = new_n1574_ & ~new_n7211_;
  assign new_n7213_ = new_n1576_ & ~new_n7212_;
  assign new_n7214_ = new_n1837_ & ~new_n7213_;
  assign new_n7215_ = new_n1068_ & ~new_n7214_;
  assign new_n7216_ = new_n1072_ & ~new_n7215_;
  assign new_n7217_ = new_n1076_ & ~new_n7216_;
  assign new_n7218_ = new_n1080_ & ~new_n7217_;
  assign new_n7219_ = new_n1084_ & ~new_n7218_;
  assign new_n7220_ = new_n1088_ & ~new_n7219_;
  assign new_n7221_ = new_n1092_ & ~new_n7220_;
  assign new_n7222_ = new_n1096_ & ~new_n7221_;
  assign new_n7223_ = new_n1100_ & ~new_n7222_;
  assign new_n7224_ = new_n1104_ & ~new_n7223_;
  assign new_n7225_ = new_n1108_ & ~new_n7224_;
  assign new_n7226_ = new_n1112_ & ~new_n7225_;
  assign new_n7227_ = new_n1116_ & ~new_n7226_;
  assign new_n7228_ = new_n1120_ & ~new_n7227_;
  assign new_n7229_ = new_n1124_ & ~new_n7228_;
  assign new_n7230_ = new_n1128_ & ~new_n7229_;
  assign new_n7231_ = new_n1132_ & ~new_n7230_;
  assign new_n7232_ = new_n1136_ & ~new_n7231_;
  assign new_n7233_ = new_n1140_ & ~new_n7232_;
  assign new_n7234_ = new_n1144_ & ~new_n7233_;
  assign new_n7235_ = new_n1148_ & ~new_n7234_;
  assign new_n7236_ = new_n1152_ & ~new_n7235_;
  assign new_n7237_ = new_n1156_ & ~new_n7236_;
  assign new_n7238_ = new_n1160_ & ~new_n7237_;
  assign new_n7239_ = new_n1164_ & ~new_n7238_;
  assign new_n7240_ = new_n1168_ & ~new_n7239_;
  assign new_n7241_ = new_n1172_ & ~new_n7240_;
  assign new_n7242_ = new_n1176_ & ~new_n7241_;
  assign new_n7243_ = new_n1180_ & ~new_n7242_;
  assign new_n7244_ = new_n1184_ & ~new_n7243_;
  assign new_n7245_ = new_n1188_ & ~new_n7244_;
  assign new_n7246_ = new_n1192_ & ~new_n7245_;
  assign new_n7247_ = new_n1196_ & ~new_n7246_;
  assign new_n7248_ = new_n1200_ & ~new_n7247_;
  assign new_n7249_ = new_n1204_ & ~new_n7248_;
  assign new_n7250_ = new_n1208_ & ~new_n7249_;
  assign new_n7251_ = new_n1212_ & ~new_n7250_;
  assign new_n7252_ = new_n1216_ & ~new_n7251_;
  assign new_n7253_ = new_n1220_ & ~new_n7252_;
  assign new_n7254_ = new_n1224_ & ~new_n7253_;
  assign new_n7255_ = new_n1228_ & ~new_n7254_;
  assign new_n7256_ = new_n1232_ & ~new_n7255_;
  assign new_n7257_ = new_n1236_ & ~new_n7256_;
  assign new_n7258_ = \req[70]  & ~new_n1238_;
  assign \grant[70]  = ~new_n7257_ & new_n7258_;
  assign new_n7260_ = ~new_n575_ & new_n1247_;
  assign new_n7261_ = new_n1252_ & ~new_n7260_;
  assign new_n7262_ = new_n1256_ & ~new_n7261_;
  assign new_n7263_ = new_n1260_ & ~new_n7262_;
  assign new_n7264_ = new_n1264_ & ~new_n7263_;
  assign new_n7265_ = new_n1268_ & ~new_n7264_;
  assign new_n7266_ = new_n1272_ & ~new_n7265_;
  assign new_n7267_ = new_n1276_ & ~new_n7266_;
  assign new_n7268_ = new_n1280_ & ~new_n7267_;
  assign new_n7269_ = new_n1284_ & ~new_n7268_;
  assign new_n7270_ = new_n1288_ & ~new_n7269_;
  assign new_n7271_ = new_n1292_ & ~new_n7270_;
  assign new_n7272_ = new_n1296_ & ~new_n7271_;
  assign new_n7273_ = new_n1300_ & ~new_n7272_;
  assign new_n7274_ = new_n1304_ & ~new_n7273_;
  assign new_n7275_ = new_n1308_ & ~new_n7274_;
  assign new_n7276_ = new_n1312_ & ~new_n7275_;
  assign new_n7277_ = new_n1316_ & ~new_n7276_;
  assign new_n7278_ = new_n1320_ & ~new_n7277_;
  assign new_n7279_ = new_n1324_ & ~new_n7278_;
  assign new_n7280_ = new_n1328_ & ~new_n7279_;
  assign new_n7281_ = new_n1332_ & ~new_n7280_;
  assign new_n7282_ = new_n1336_ & ~new_n7281_;
  assign new_n7283_ = new_n1340_ & ~new_n7282_;
  assign new_n7284_ = new_n1344_ & ~new_n7283_;
  assign new_n7285_ = new_n1348_ & ~new_n7284_;
  assign new_n7286_ = new_n1352_ & ~new_n7285_;
  assign new_n7287_ = new_n1356_ & ~new_n7286_;
  assign new_n7288_ = new_n1360_ & ~new_n7287_;
  assign new_n7289_ = new_n1364_ & ~new_n7288_;
  assign new_n7290_ = new_n1368_ & ~new_n7289_;
  assign new_n7291_ = new_n1372_ & ~new_n7290_;
  assign new_n7292_ = new_n1376_ & ~new_n7291_;
  assign new_n7293_ = new_n1380_ & ~new_n7292_;
  assign new_n7294_ = new_n1384_ & ~new_n7293_;
  assign new_n7295_ = new_n1388_ & ~new_n7294_;
  assign new_n7296_ = new_n1392_ & ~new_n7295_;
  assign new_n7297_ = new_n1396_ & ~new_n7296_;
  assign new_n7298_ = new_n1663_ & ~new_n7297_;
  assign new_n7299_ = new_n392_ & ~new_n7298_;
  assign new_n7300_ = new_n396_ & ~new_n7299_;
  assign new_n7301_ = new_n400_ & ~new_n7300_;
  assign new_n7302_ = new_n404_ & ~new_n7301_;
  assign new_n7303_ = new_n408_ & ~new_n7302_;
  assign new_n7304_ = new_n412_ & ~new_n7303_;
  assign new_n7305_ = new_n416_ & ~new_n7304_;
  assign new_n7306_ = new_n420_ & ~new_n7305_;
  assign new_n7307_ = new_n424_ & ~new_n7306_;
  assign new_n7308_ = new_n428_ & ~new_n7307_;
  assign new_n7309_ = new_n432_ & ~new_n7308_;
  assign new_n7310_ = new_n436_ & ~new_n7309_;
  assign new_n7311_ = new_n440_ & ~new_n7310_;
  assign new_n7312_ = new_n444_ & ~new_n7311_;
  assign new_n7313_ = new_n448_ & ~new_n7312_;
  assign new_n7314_ = new_n452_ & ~new_n7313_;
  assign new_n7315_ = new_n456_ & ~new_n7314_;
  assign new_n7316_ = new_n460_ & ~new_n7315_;
  assign new_n7317_ = new_n464_ & ~new_n7316_;
  assign new_n7318_ = new_n468_ & ~new_n7317_;
  assign new_n7319_ = new_n472_ & ~new_n7318_;
  assign new_n7320_ = new_n476_ & ~new_n7319_;
  assign new_n7321_ = new_n480_ & ~new_n7320_;
  assign new_n7322_ = new_n484_ & ~new_n7321_;
  assign new_n7323_ = new_n488_ & ~new_n7322_;
  assign new_n7324_ = new_n492_ & ~new_n7323_;
  assign new_n7325_ = new_n496_ & ~new_n7324_;
  assign new_n7326_ = new_n500_ & ~new_n7325_;
  assign new_n7327_ = new_n504_ & ~new_n7326_;
  assign new_n7328_ = new_n508_ & ~new_n7327_;
  assign new_n7329_ = new_n512_ & ~new_n7328_;
  assign new_n7330_ = new_n516_ & ~new_n7329_;
  assign new_n7331_ = new_n520_ & ~new_n7330_;
  assign new_n7332_ = new_n524_ & ~new_n7331_;
  assign new_n7333_ = new_n528_ & ~new_n7332_;
  assign new_n7334_ = new_n532_ & ~new_n7333_;
  assign new_n7335_ = new_n536_ & ~new_n7334_;
  assign new_n7336_ = new_n540_ & ~new_n7335_;
  assign new_n7337_ = new_n544_ & ~new_n7336_;
  assign new_n7338_ = new_n548_ & ~new_n7337_;
  assign new_n7339_ = new_n552_ & ~new_n7338_;
  assign new_n7340_ = new_n556_ & ~new_n7339_;
  assign new_n7341_ = new_n560_ & ~new_n7340_;
  assign new_n7342_ = new_n564_ & ~new_n7341_;
  assign new_n7343_ = new_n568_ & ~new_n7342_;
  assign new_n7344_ = \req[71]  & ~new_n570_;
  assign \grant[71]  = ~new_n7343_ & new_n7344_;
  assign new_n7346_ = new_n579_ & ~new_n914_;
  assign new_n7347_ = new_n584_ & ~new_n7346_;
  assign new_n7348_ = new_n588_ & ~new_n7347_;
  assign new_n7349_ = new_n592_ & ~new_n7348_;
  assign new_n7350_ = new_n596_ & ~new_n7349_;
  assign new_n7351_ = new_n600_ & ~new_n7350_;
  assign new_n7352_ = new_n604_ & ~new_n7351_;
  assign new_n7353_ = new_n608_ & ~new_n7352_;
  assign new_n7354_ = new_n612_ & ~new_n7353_;
  assign new_n7355_ = new_n616_ & ~new_n7354_;
  assign new_n7356_ = new_n620_ & ~new_n7355_;
  assign new_n7357_ = new_n624_ & ~new_n7356_;
  assign new_n7358_ = new_n628_ & ~new_n7357_;
  assign new_n7359_ = new_n632_ & ~new_n7358_;
  assign new_n7360_ = new_n636_ & ~new_n7359_;
  assign new_n7361_ = new_n640_ & ~new_n7360_;
  assign new_n7362_ = new_n644_ & ~new_n7361_;
  assign new_n7363_ = new_n648_ & ~new_n7362_;
  assign new_n7364_ = new_n652_ & ~new_n7363_;
  assign new_n7365_ = new_n656_ & ~new_n7364_;
  assign new_n7366_ = new_n660_ & ~new_n7365_;
  assign new_n7367_ = new_n664_ & ~new_n7366_;
  assign new_n7368_ = new_n668_ & ~new_n7367_;
  assign new_n7369_ = new_n672_ & ~new_n7368_;
  assign new_n7370_ = new_n676_ & ~new_n7369_;
  assign new_n7371_ = new_n680_ & ~new_n7370_;
  assign new_n7372_ = new_n684_ & ~new_n7371_;
  assign new_n7373_ = new_n688_ & ~new_n7372_;
  assign new_n7374_ = new_n692_ & ~new_n7373_;
  assign new_n7375_ = new_n696_ & ~new_n7374_;
  assign new_n7376_ = new_n700_ & ~new_n7375_;
  assign new_n7377_ = new_n704_ & ~new_n7376_;
  assign new_n7378_ = new_n708_ & ~new_n7377_;
  assign new_n7379_ = new_n712_ & ~new_n7378_;
  assign new_n7380_ = new_n716_ & ~new_n7379_;
  assign new_n7381_ = new_n720_ & ~new_n7380_;
  assign new_n7382_ = new_n1484_ & ~new_n7381_;
  assign new_n7383_ = new_n1486_ & ~new_n7382_;
  assign new_n7384_ = new_n1750_ & ~new_n7383_;
  assign new_n7385_ = new_n731_ & ~new_n7384_;
  assign new_n7386_ = new_n735_ & ~new_n7385_;
  assign new_n7387_ = new_n739_ & ~new_n7386_;
  assign new_n7388_ = new_n743_ & ~new_n7387_;
  assign new_n7389_ = new_n747_ & ~new_n7388_;
  assign new_n7390_ = new_n751_ & ~new_n7389_;
  assign new_n7391_ = new_n755_ & ~new_n7390_;
  assign new_n7392_ = new_n759_ & ~new_n7391_;
  assign new_n7393_ = new_n763_ & ~new_n7392_;
  assign new_n7394_ = new_n767_ & ~new_n7393_;
  assign new_n7395_ = new_n771_ & ~new_n7394_;
  assign new_n7396_ = new_n775_ & ~new_n7395_;
  assign new_n7397_ = new_n779_ & ~new_n7396_;
  assign new_n7398_ = new_n783_ & ~new_n7397_;
  assign new_n7399_ = new_n787_ & ~new_n7398_;
  assign new_n7400_ = new_n791_ & ~new_n7399_;
  assign new_n7401_ = new_n795_ & ~new_n7400_;
  assign new_n7402_ = new_n799_ & ~new_n7401_;
  assign new_n7403_ = new_n803_ & ~new_n7402_;
  assign new_n7404_ = new_n807_ & ~new_n7403_;
  assign new_n7405_ = new_n811_ & ~new_n7404_;
  assign new_n7406_ = new_n815_ & ~new_n7405_;
  assign new_n7407_ = new_n819_ & ~new_n7406_;
  assign new_n7408_ = new_n823_ & ~new_n7407_;
  assign new_n7409_ = new_n827_ & ~new_n7408_;
  assign new_n7410_ = new_n831_ & ~new_n7409_;
  assign new_n7411_ = new_n835_ & ~new_n7410_;
  assign new_n7412_ = new_n839_ & ~new_n7411_;
  assign new_n7413_ = new_n843_ & ~new_n7412_;
  assign new_n7414_ = new_n847_ & ~new_n7413_;
  assign new_n7415_ = new_n851_ & ~new_n7414_;
  assign new_n7416_ = new_n855_ & ~new_n7415_;
  assign new_n7417_ = new_n859_ & ~new_n7416_;
  assign new_n7418_ = new_n863_ & ~new_n7417_;
  assign new_n7419_ = new_n867_ & ~new_n7418_;
  assign new_n7420_ = new_n871_ & ~new_n7419_;
  assign new_n7421_ = new_n875_ & ~new_n7420_;
  assign new_n7422_ = new_n879_ & ~new_n7421_;
  assign new_n7423_ = new_n883_ & ~new_n7422_;
  assign new_n7424_ = new_n887_ & ~new_n7423_;
  assign new_n7425_ = new_n891_ & ~new_n7424_;
  assign new_n7426_ = new_n895_ & ~new_n7425_;
  assign new_n7427_ = new_n899_ & ~new_n7426_;
  assign new_n7428_ = new_n903_ & ~new_n7427_;
  assign new_n7429_ = new_n907_ & ~new_n7428_;
  assign new_n7430_ = \req[72]  & ~new_n909_;
  assign \grant[72]  = ~new_n7429_ & new_n7430_;
  assign new_n7432_ = new_n918_ & ~new_n1251_;
  assign new_n7433_ = new_n923_ & ~new_n7432_;
  assign new_n7434_ = new_n927_ & ~new_n7433_;
  assign new_n7435_ = new_n931_ & ~new_n7434_;
  assign new_n7436_ = new_n935_ & ~new_n7435_;
  assign new_n7437_ = new_n939_ & ~new_n7436_;
  assign new_n7438_ = new_n943_ & ~new_n7437_;
  assign new_n7439_ = new_n947_ & ~new_n7438_;
  assign new_n7440_ = new_n951_ & ~new_n7439_;
  assign new_n7441_ = new_n955_ & ~new_n7440_;
  assign new_n7442_ = new_n959_ & ~new_n7441_;
  assign new_n7443_ = new_n963_ & ~new_n7442_;
  assign new_n7444_ = new_n967_ & ~new_n7443_;
  assign new_n7445_ = new_n971_ & ~new_n7444_;
  assign new_n7446_ = new_n975_ & ~new_n7445_;
  assign new_n7447_ = new_n979_ & ~new_n7446_;
  assign new_n7448_ = new_n983_ & ~new_n7447_;
  assign new_n7449_ = new_n987_ & ~new_n7448_;
  assign new_n7450_ = new_n991_ & ~new_n7449_;
  assign new_n7451_ = new_n995_ & ~new_n7450_;
  assign new_n7452_ = new_n999_ & ~new_n7451_;
  assign new_n7453_ = new_n1003_ & ~new_n7452_;
  assign new_n7454_ = new_n1007_ & ~new_n7453_;
  assign new_n7455_ = new_n1011_ & ~new_n7454_;
  assign new_n7456_ = new_n1015_ & ~new_n7455_;
  assign new_n7457_ = new_n1019_ & ~new_n7456_;
  assign new_n7458_ = new_n1023_ & ~new_n7457_;
  assign new_n7459_ = new_n1027_ & ~new_n7458_;
  assign new_n7460_ = new_n1031_ & ~new_n7459_;
  assign new_n7461_ = new_n1035_ & ~new_n7460_;
  assign new_n7462_ = new_n1039_ & ~new_n7461_;
  assign new_n7463_ = new_n1043_ & ~new_n7462_;
  assign new_n7464_ = new_n1047_ & ~new_n7463_;
  assign new_n7465_ = new_n1051_ & ~new_n7464_;
  assign new_n7466_ = new_n1055_ & ~new_n7465_;
  assign new_n7467_ = new_n1059_ & ~new_n7466_;
  assign new_n7468_ = new_n1574_ & ~new_n7467_;
  assign new_n7469_ = new_n1576_ & ~new_n7468_;
  assign new_n7470_ = new_n1837_ & ~new_n7469_;
  assign new_n7471_ = new_n1068_ & ~new_n7470_;
  assign new_n7472_ = new_n1072_ & ~new_n7471_;
  assign new_n7473_ = new_n1076_ & ~new_n7472_;
  assign new_n7474_ = new_n1080_ & ~new_n7473_;
  assign new_n7475_ = new_n1084_ & ~new_n7474_;
  assign new_n7476_ = new_n1088_ & ~new_n7475_;
  assign new_n7477_ = new_n1092_ & ~new_n7476_;
  assign new_n7478_ = new_n1096_ & ~new_n7477_;
  assign new_n7479_ = new_n1100_ & ~new_n7478_;
  assign new_n7480_ = new_n1104_ & ~new_n7479_;
  assign new_n7481_ = new_n1108_ & ~new_n7480_;
  assign new_n7482_ = new_n1112_ & ~new_n7481_;
  assign new_n7483_ = new_n1116_ & ~new_n7482_;
  assign new_n7484_ = new_n1120_ & ~new_n7483_;
  assign new_n7485_ = new_n1124_ & ~new_n7484_;
  assign new_n7486_ = new_n1128_ & ~new_n7485_;
  assign new_n7487_ = new_n1132_ & ~new_n7486_;
  assign new_n7488_ = new_n1136_ & ~new_n7487_;
  assign new_n7489_ = new_n1140_ & ~new_n7488_;
  assign new_n7490_ = new_n1144_ & ~new_n7489_;
  assign new_n7491_ = new_n1148_ & ~new_n7490_;
  assign new_n7492_ = new_n1152_ & ~new_n7491_;
  assign new_n7493_ = new_n1156_ & ~new_n7492_;
  assign new_n7494_ = new_n1160_ & ~new_n7493_;
  assign new_n7495_ = new_n1164_ & ~new_n7494_;
  assign new_n7496_ = new_n1168_ & ~new_n7495_;
  assign new_n7497_ = new_n1172_ & ~new_n7496_;
  assign new_n7498_ = new_n1176_ & ~new_n7497_;
  assign new_n7499_ = new_n1180_ & ~new_n7498_;
  assign new_n7500_ = new_n1184_ & ~new_n7499_;
  assign new_n7501_ = new_n1188_ & ~new_n7500_;
  assign new_n7502_ = new_n1192_ & ~new_n7501_;
  assign new_n7503_ = new_n1196_ & ~new_n7502_;
  assign new_n7504_ = new_n1200_ & ~new_n7503_;
  assign new_n7505_ = new_n1204_ & ~new_n7504_;
  assign new_n7506_ = new_n1208_ & ~new_n7505_;
  assign new_n7507_ = new_n1212_ & ~new_n7506_;
  assign new_n7508_ = new_n1216_ & ~new_n7507_;
  assign new_n7509_ = new_n1220_ & ~new_n7508_;
  assign new_n7510_ = new_n1224_ & ~new_n7509_;
  assign new_n7511_ = new_n1228_ & ~new_n7510_;
  assign new_n7512_ = new_n1232_ & ~new_n7511_;
  assign new_n7513_ = new_n1236_ & ~new_n7512_;
  assign new_n7514_ = new_n1240_ & ~new_n7513_;
  assign new_n7515_ = new_n1244_ & ~new_n7514_;
  assign new_n7516_ = \req[73]  & ~new_n1246_;
  assign \grant[73]  = ~new_n7515_ & new_n7516_;
  assign new_n7518_ = ~new_n583_ & new_n1255_;
  assign new_n7519_ = new_n1260_ & ~new_n7518_;
  assign new_n7520_ = new_n1264_ & ~new_n7519_;
  assign new_n7521_ = new_n1268_ & ~new_n7520_;
  assign new_n7522_ = new_n1272_ & ~new_n7521_;
  assign new_n7523_ = new_n1276_ & ~new_n7522_;
  assign new_n7524_ = new_n1280_ & ~new_n7523_;
  assign new_n7525_ = new_n1284_ & ~new_n7524_;
  assign new_n7526_ = new_n1288_ & ~new_n7525_;
  assign new_n7527_ = new_n1292_ & ~new_n7526_;
  assign new_n7528_ = new_n1296_ & ~new_n7527_;
  assign new_n7529_ = new_n1300_ & ~new_n7528_;
  assign new_n7530_ = new_n1304_ & ~new_n7529_;
  assign new_n7531_ = new_n1308_ & ~new_n7530_;
  assign new_n7532_ = new_n1312_ & ~new_n7531_;
  assign new_n7533_ = new_n1316_ & ~new_n7532_;
  assign new_n7534_ = new_n1320_ & ~new_n7533_;
  assign new_n7535_ = new_n1324_ & ~new_n7534_;
  assign new_n7536_ = new_n1328_ & ~new_n7535_;
  assign new_n7537_ = new_n1332_ & ~new_n7536_;
  assign new_n7538_ = new_n1336_ & ~new_n7537_;
  assign new_n7539_ = new_n1340_ & ~new_n7538_;
  assign new_n7540_ = new_n1344_ & ~new_n7539_;
  assign new_n7541_ = new_n1348_ & ~new_n7540_;
  assign new_n7542_ = new_n1352_ & ~new_n7541_;
  assign new_n7543_ = new_n1356_ & ~new_n7542_;
  assign new_n7544_ = new_n1360_ & ~new_n7543_;
  assign new_n7545_ = new_n1364_ & ~new_n7544_;
  assign new_n7546_ = new_n1368_ & ~new_n7545_;
  assign new_n7547_ = new_n1372_ & ~new_n7546_;
  assign new_n7548_ = new_n1376_ & ~new_n7547_;
  assign new_n7549_ = new_n1380_ & ~new_n7548_;
  assign new_n7550_ = new_n1384_ & ~new_n7549_;
  assign new_n7551_ = new_n1388_ & ~new_n7550_;
  assign new_n7552_ = new_n1392_ & ~new_n7551_;
  assign new_n7553_ = new_n1396_ & ~new_n7552_;
  assign new_n7554_ = new_n1663_ & ~new_n7553_;
  assign new_n7555_ = new_n392_ & ~new_n7554_;
  assign new_n7556_ = new_n396_ & ~new_n7555_;
  assign new_n7557_ = new_n400_ & ~new_n7556_;
  assign new_n7558_ = new_n404_ & ~new_n7557_;
  assign new_n7559_ = new_n408_ & ~new_n7558_;
  assign new_n7560_ = new_n412_ & ~new_n7559_;
  assign new_n7561_ = new_n416_ & ~new_n7560_;
  assign new_n7562_ = new_n420_ & ~new_n7561_;
  assign new_n7563_ = new_n424_ & ~new_n7562_;
  assign new_n7564_ = new_n428_ & ~new_n7563_;
  assign new_n7565_ = new_n432_ & ~new_n7564_;
  assign new_n7566_ = new_n436_ & ~new_n7565_;
  assign new_n7567_ = new_n440_ & ~new_n7566_;
  assign new_n7568_ = new_n444_ & ~new_n7567_;
  assign new_n7569_ = new_n448_ & ~new_n7568_;
  assign new_n7570_ = new_n452_ & ~new_n7569_;
  assign new_n7571_ = new_n456_ & ~new_n7570_;
  assign new_n7572_ = new_n460_ & ~new_n7571_;
  assign new_n7573_ = new_n464_ & ~new_n7572_;
  assign new_n7574_ = new_n468_ & ~new_n7573_;
  assign new_n7575_ = new_n472_ & ~new_n7574_;
  assign new_n7576_ = new_n476_ & ~new_n7575_;
  assign new_n7577_ = new_n480_ & ~new_n7576_;
  assign new_n7578_ = new_n484_ & ~new_n7577_;
  assign new_n7579_ = new_n488_ & ~new_n7578_;
  assign new_n7580_ = new_n492_ & ~new_n7579_;
  assign new_n7581_ = new_n496_ & ~new_n7580_;
  assign new_n7582_ = new_n500_ & ~new_n7581_;
  assign new_n7583_ = new_n504_ & ~new_n7582_;
  assign new_n7584_ = new_n508_ & ~new_n7583_;
  assign new_n7585_ = new_n512_ & ~new_n7584_;
  assign new_n7586_ = new_n516_ & ~new_n7585_;
  assign new_n7587_ = new_n520_ & ~new_n7586_;
  assign new_n7588_ = new_n524_ & ~new_n7587_;
  assign new_n7589_ = new_n528_ & ~new_n7588_;
  assign new_n7590_ = new_n532_ & ~new_n7589_;
  assign new_n7591_ = new_n536_ & ~new_n7590_;
  assign new_n7592_ = new_n540_ & ~new_n7591_;
  assign new_n7593_ = new_n544_ & ~new_n7592_;
  assign new_n7594_ = new_n548_ & ~new_n7593_;
  assign new_n7595_ = new_n552_ & ~new_n7594_;
  assign new_n7596_ = new_n556_ & ~new_n7595_;
  assign new_n7597_ = new_n560_ & ~new_n7596_;
  assign new_n7598_ = new_n564_ & ~new_n7597_;
  assign new_n7599_ = new_n568_ & ~new_n7598_;
  assign new_n7600_ = new_n572_ & ~new_n7599_;
  assign new_n7601_ = new_n576_ & ~new_n7600_;
  assign new_n7602_ = \req[74]  & ~new_n578_;
  assign \grant[74]  = ~new_n7601_ & new_n7602_;
  assign new_n7604_ = new_n587_ & ~new_n922_;
  assign new_n7605_ = new_n592_ & ~new_n7604_;
  assign new_n7606_ = new_n596_ & ~new_n7605_;
  assign new_n7607_ = new_n600_ & ~new_n7606_;
  assign new_n7608_ = new_n604_ & ~new_n7607_;
  assign new_n7609_ = new_n608_ & ~new_n7608_;
  assign new_n7610_ = new_n612_ & ~new_n7609_;
  assign new_n7611_ = new_n616_ & ~new_n7610_;
  assign new_n7612_ = new_n620_ & ~new_n7611_;
  assign new_n7613_ = new_n624_ & ~new_n7612_;
  assign new_n7614_ = new_n628_ & ~new_n7613_;
  assign new_n7615_ = new_n632_ & ~new_n7614_;
  assign new_n7616_ = new_n636_ & ~new_n7615_;
  assign new_n7617_ = new_n640_ & ~new_n7616_;
  assign new_n7618_ = new_n644_ & ~new_n7617_;
  assign new_n7619_ = new_n648_ & ~new_n7618_;
  assign new_n7620_ = new_n652_ & ~new_n7619_;
  assign new_n7621_ = new_n656_ & ~new_n7620_;
  assign new_n7622_ = new_n660_ & ~new_n7621_;
  assign new_n7623_ = new_n664_ & ~new_n7622_;
  assign new_n7624_ = new_n668_ & ~new_n7623_;
  assign new_n7625_ = new_n672_ & ~new_n7624_;
  assign new_n7626_ = new_n676_ & ~new_n7625_;
  assign new_n7627_ = new_n680_ & ~new_n7626_;
  assign new_n7628_ = new_n684_ & ~new_n7627_;
  assign new_n7629_ = new_n688_ & ~new_n7628_;
  assign new_n7630_ = new_n692_ & ~new_n7629_;
  assign new_n7631_ = new_n696_ & ~new_n7630_;
  assign new_n7632_ = new_n700_ & ~new_n7631_;
  assign new_n7633_ = new_n704_ & ~new_n7632_;
  assign new_n7634_ = new_n708_ & ~new_n7633_;
  assign new_n7635_ = new_n712_ & ~new_n7634_;
  assign new_n7636_ = new_n716_ & ~new_n7635_;
  assign new_n7637_ = new_n720_ & ~new_n7636_;
  assign new_n7638_ = new_n1484_ & ~new_n7637_;
  assign new_n7639_ = new_n1486_ & ~new_n7638_;
  assign new_n7640_ = new_n1750_ & ~new_n7639_;
  assign new_n7641_ = new_n731_ & ~new_n7640_;
  assign new_n7642_ = new_n735_ & ~new_n7641_;
  assign new_n7643_ = new_n739_ & ~new_n7642_;
  assign new_n7644_ = new_n743_ & ~new_n7643_;
  assign new_n7645_ = new_n747_ & ~new_n7644_;
  assign new_n7646_ = new_n751_ & ~new_n7645_;
  assign new_n7647_ = new_n755_ & ~new_n7646_;
  assign new_n7648_ = new_n759_ & ~new_n7647_;
  assign new_n7649_ = new_n763_ & ~new_n7648_;
  assign new_n7650_ = new_n767_ & ~new_n7649_;
  assign new_n7651_ = new_n771_ & ~new_n7650_;
  assign new_n7652_ = new_n775_ & ~new_n7651_;
  assign new_n7653_ = new_n779_ & ~new_n7652_;
  assign new_n7654_ = new_n783_ & ~new_n7653_;
  assign new_n7655_ = new_n787_ & ~new_n7654_;
  assign new_n7656_ = new_n791_ & ~new_n7655_;
  assign new_n7657_ = new_n795_ & ~new_n7656_;
  assign new_n7658_ = new_n799_ & ~new_n7657_;
  assign new_n7659_ = new_n803_ & ~new_n7658_;
  assign new_n7660_ = new_n807_ & ~new_n7659_;
  assign new_n7661_ = new_n811_ & ~new_n7660_;
  assign new_n7662_ = new_n815_ & ~new_n7661_;
  assign new_n7663_ = new_n819_ & ~new_n7662_;
  assign new_n7664_ = new_n823_ & ~new_n7663_;
  assign new_n7665_ = new_n827_ & ~new_n7664_;
  assign new_n7666_ = new_n831_ & ~new_n7665_;
  assign new_n7667_ = new_n835_ & ~new_n7666_;
  assign new_n7668_ = new_n839_ & ~new_n7667_;
  assign new_n7669_ = new_n843_ & ~new_n7668_;
  assign new_n7670_ = new_n847_ & ~new_n7669_;
  assign new_n7671_ = new_n851_ & ~new_n7670_;
  assign new_n7672_ = new_n855_ & ~new_n7671_;
  assign new_n7673_ = new_n859_ & ~new_n7672_;
  assign new_n7674_ = new_n863_ & ~new_n7673_;
  assign new_n7675_ = new_n867_ & ~new_n7674_;
  assign new_n7676_ = new_n871_ & ~new_n7675_;
  assign new_n7677_ = new_n875_ & ~new_n7676_;
  assign new_n7678_ = new_n879_ & ~new_n7677_;
  assign new_n7679_ = new_n883_ & ~new_n7678_;
  assign new_n7680_ = new_n887_ & ~new_n7679_;
  assign new_n7681_ = new_n891_ & ~new_n7680_;
  assign new_n7682_ = new_n895_ & ~new_n7681_;
  assign new_n7683_ = new_n899_ & ~new_n7682_;
  assign new_n7684_ = new_n903_ & ~new_n7683_;
  assign new_n7685_ = new_n907_ & ~new_n7684_;
  assign new_n7686_ = new_n911_ & ~new_n7685_;
  assign new_n7687_ = new_n915_ & ~new_n7686_;
  assign new_n7688_ = \req[75]  & ~new_n917_;
  assign \grant[75]  = ~new_n7687_ & new_n7688_;
  assign new_n7690_ = new_n926_ & ~new_n1259_;
  assign new_n7691_ = new_n931_ & ~new_n7690_;
  assign new_n7692_ = new_n935_ & ~new_n7691_;
  assign new_n7693_ = new_n939_ & ~new_n7692_;
  assign new_n7694_ = new_n943_ & ~new_n7693_;
  assign new_n7695_ = new_n947_ & ~new_n7694_;
  assign new_n7696_ = new_n951_ & ~new_n7695_;
  assign new_n7697_ = new_n955_ & ~new_n7696_;
  assign new_n7698_ = new_n959_ & ~new_n7697_;
  assign new_n7699_ = new_n963_ & ~new_n7698_;
  assign new_n7700_ = new_n967_ & ~new_n7699_;
  assign new_n7701_ = new_n971_ & ~new_n7700_;
  assign new_n7702_ = new_n975_ & ~new_n7701_;
  assign new_n7703_ = new_n979_ & ~new_n7702_;
  assign new_n7704_ = new_n983_ & ~new_n7703_;
  assign new_n7705_ = new_n987_ & ~new_n7704_;
  assign new_n7706_ = new_n991_ & ~new_n7705_;
  assign new_n7707_ = new_n995_ & ~new_n7706_;
  assign new_n7708_ = new_n999_ & ~new_n7707_;
  assign new_n7709_ = new_n1003_ & ~new_n7708_;
  assign new_n7710_ = new_n1007_ & ~new_n7709_;
  assign new_n7711_ = new_n1011_ & ~new_n7710_;
  assign new_n7712_ = new_n1015_ & ~new_n7711_;
  assign new_n7713_ = new_n1019_ & ~new_n7712_;
  assign new_n7714_ = new_n1023_ & ~new_n7713_;
  assign new_n7715_ = new_n1027_ & ~new_n7714_;
  assign new_n7716_ = new_n1031_ & ~new_n7715_;
  assign new_n7717_ = new_n1035_ & ~new_n7716_;
  assign new_n7718_ = new_n1039_ & ~new_n7717_;
  assign new_n7719_ = new_n1043_ & ~new_n7718_;
  assign new_n7720_ = new_n1047_ & ~new_n7719_;
  assign new_n7721_ = new_n1051_ & ~new_n7720_;
  assign new_n7722_ = new_n1055_ & ~new_n7721_;
  assign new_n7723_ = new_n1059_ & ~new_n7722_;
  assign new_n7724_ = new_n1574_ & ~new_n7723_;
  assign new_n7725_ = new_n1576_ & ~new_n7724_;
  assign new_n7726_ = new_n1837_ & ~new_n7725_;
  assign new_n7727_ = new_n1068_ & ~new_n7726_;
  assign new_n7728_ = new_n1072_ & ~new_n7727_;
  assign new_n7729_ = new_n1076_ & ~new_n7728_;
  assign new_n7730_ = new_n1080_ & ~new_n7729_;
  assign new_n7731_ = new_n1084_ & ~new_n7730_;
  assign new_n7732_ = new_n1088_ & ~new_n7731_;
  assign new_n7733_ = new_n1092_ & ~new_n7732_;
  assign new_n7734_ = new_n1096_ & ~new_n7733_;
  assign new_n7735_ = new_n1100_ & ~new_n7734_;
  assign new_n7736_ = new_n1104_ & ~new_n7735_;
  assign new_n7737_ = new_n1108_ & ~new_n7736_;
  assign new_n7738_ = new_n1112_ & ~new_n7737_;
  assign new_n7739_ = new_n1116_ & ~new_n7738_;
  assign new_n7740_ = new_n1120_ & ~new_n7739_;
  assign new_n7741_ = new_n1124_ & ~new_n7740_;
  assign new_n7742_ = new_n1128_ & ~new_n7741_;
  assign new_n7743_ = new_n1132_ & ~new_n7742_;
  assign new_n7744_ = new_n1136_ & ~new_n7743_;
  assign new_n7745_ = new_n1140_ & ~new_n7744_;
  assign new_n7746_ = new_n1144_ & ~new_n7745_;
  assign new_n7747_ = new_n1148_ & ~new_n7746_;
  assign new_n7748_ = new_n1152_ & ~new_n7747_;
  assign new_n7749_ = new_n1156_ & ~new_n7748_;
  assign new_n7750_ = new_n1160_ & ~new_n7749_;
  assign new_n7751_ = new_n1164_ & ~new_n7750_;
  assign new_n7752_ = new_n1168_ & ~new_n7751_;
  assign new_n7753_ = new_n1172_ & ~new_n7752_;
  assign new_n7754_ = new_n1176_ & ~new_n7753_;
  assign new_n7755_ = new_n1180_ & ~new_n7754_;
  assign new_n7756_ = new_n1184_ & ~new_n7755_;
  assign new_n7757_ = new_n1188_ & ~new_n7756_;
  assign new_n7758_ = new_n1192_ & ~new_n7757_;
  assign new_n7759_ = new_n1196_ & ~new_n7758_;
  assign new_n7760_ = new_n1200_ & ~new_n7759_;
  assign new_n7761_ = new_n1204_ & ~new_n7760_;
  assign new_n7762_ = new_n1208_ & ~new_n7761_;
  assign new_n7763_ = new_n1212_ & ~new_n7762_;
  assign new_n7764_ = new_n1216_ & ~new_n7763_;
  assign new_n7765_ = new_n1220_ & ~new_n7764_;
  assign new_n7766_ = new_n1224_ & ~new_n7765_;
  assign new_n7767_ = new_n1228_ & ~new_n7766_;
  assign new_n7768_ = new_n1232_ & ~new_n7767_;
  assign new_n7769_ = new_n1236_ & ~new_n7768_;
  assign new_n7770_ = new_n1240_ & ~new_n7769_;
  assign new_n7771_ = new_n1244_ & ~new_n7770_;
  assign new_n7772_ = new_n1248_ & ~new_n7771_;
  assign new_n7773_ = new_n1252_ & ~new_n7772_;
  assign new_n7774_ = \req[76]  & ~new_n1254_;
  assign \grant[76]  = ~new_n7773_ & new_n7774_;
  assign new_n7776_ = ~new_n591_ & new_n1263_;
  assign new_n7777_ = new_n1268_ & ~new_n7776_;
  assign new_n7778_ = new_n1272_ & ~new_n7777_;
  assign new_n7779_ = new_n1276_ & ~new_n7778_;
  assign new_n7780_ = new_n1280_ & ~new_n7779_;
  assign new_n7781_ = new_n1284_ & ~new_n7780_;
  assign new_n7782_ = new_n1288_ & ~new_n7781_;
  assign new_n7783_ = new_n1292_ & ~new_n7782_;
  assign new_n7784_ = new_n1296_ & ~new_n7783_;
  assign new_n7785_ = new_n1300_ & ~new_n7784_;
  assign new_n7786_ = new_n1304_ & ~new_n7785_;
  assign new_n7787_ = new_n1308_ & ~new_n7786_;
  assign new_n7788_ = new_n1312_ & ~new_n7787_;
  assign new_n7789_ = new_n1316_ & ~new_n7788_;
  assign new_n7790_ = new_n1320_ & ~new_n7789_;
  assign new_n7791_ = new_n1324_ & ~new_n7790_;
  assign new_n7792_ = new_n1328_ & ~new_n7791_;
  assign new_n7793_ = new_n1332_ & ~new_n7792_;
  assign new_n7794_ = new_n1336_ & ~new_n7793_;
  assign new_n7795_ = new_n1340_ & ~new_n7794_;
  assign new_n7796_ = new_n1344_ & ~new_n7795_;
  assign new_n7797_ = new_n1348_ & ~new_n7796_;
  assign new_n7798_ = new_n1352_ & ~new_n7797_;
  assign new_n7799_ = new_n1356_ & ~new_n7798_;
  assign new_n7800_ = new_n1360_ & ~new_n7799_;
  assign new_n7801_ = new_n1364_ & ~new_n7800_;
  assign new_n7802_ = new_n1368_ & ~new_n7801_;
  assign new_n7803_ = new_n1372_ & ~new_n7802_;
  assign new_n7804_ = new_n1376_ & ~new_n7803_;
  assign new_n7805_ = new_n1380_ & ~new_n7804_;
  assign new_n7806_ = new_n1384_ & ~new_n7805_;
  assign new_n7807_ = new_n1388_ & ~new_n7806_;
  assign new_n7808_ = new_n1392_ & ~new_n7807_;
  assign new_n7809_ = new_n1396_ & ~new_n7808_;
  assign new_n7810_ = new_n1663_ & ~new_n7809_;
  assign new_n7811_ = new_n392_ & ~new_n7810_;
  assign new_n7812_ = new_n396_ & ~new_n7811_;
  assign new_n7813_ = new_n400_ & ~new_n7812_;
  assign new_n7814_ = new_n404_ & ~new_n7813_;
  assign new_n7815_ = new_n408_ & ~new_n7814_;
  assign new_n7816_ = new_n412_ & ~new_n7815_;
  assign new_n7817_ = new_n416_ & ~new_n7816_;
  assign new_n7818_ = new_n420_ & ~new_n7817_;
  assign new_n7819_ = new_n424_ & ~new_n7818_;
  assign new_n7820_ = new_n428_ & ~new_n7819_;
  assign new_n7821_ = new_n432_ & ~new_n7820_;
  assign new_n7822_ = new_n436_ & ~new_n7821_;
  assign new_n7823_ = new_n440_ & ~new_n7822_;
  assign new_n7824_ = new_n444_ & ~new_n7823_;
  assign new_n7825_ = new_n448_ & ~new_n7824_;
  assign new_n7826_ = new_n452_ & ~new_n7825_;
  assign new_n7827_ = new_n456_ & ~new_n7826_;
  assign new_n7828_ = new_n460_ & ~new_n7827_;
  assign new_n7829_ = new_n464_ & ~new_n7828_;
  assign new_n7830_ = new_n468_ & ~new_n7829_;
  assign new_n7831_ = new_n472_ & ~new_n7830_;
  assign new_n7832_ = new_n476_ & ~new_n7831_;
  assign new_n7833_ = new_n480_ & ~new_n7832_;
  assign new_n7834_ = new_n484_ & ~new_n7833_;
  assign new_n7835_ = new_n488_ & ~new_n7834_;
  assign new_n7836_ = new_n492_ & ~new_n7835_;
  assign new_n7837_ = new_n496_ & ~new_n7836_;
  assign new_n7838_ = new_n500_ & ~new_n7837_;
  assign new_n7839_ = new_n504_ & ~new_n7838_;
  assign new_n7840_ = new_n508_ & ~new_n7839_;
  assign new_n7841_ = new_n512_ & ~new_n7840_;
  assign new_n7842_ = new_n516_ & ~new_n7841_;
  assign new_n7843_ = new_n520_ & ~new_n7842_;
  assign new_n7844_ = new_n524_ & ~new_n7843_;
  assign new_n7845_ = new_n528_ & ~new_n7844_;
  assign new_n7846_ = new_n532_ & ~new_n7845_;
  assign new_n7847_ = new_n536_ & ~new_n7846_;
  assign new_n7848_ = new_n540_ & ~new_n7847_;
  assign new_n7849_ = new_n544_ & ~new_n7848_;
  assign new_n7850_ = new_n548_ & ~new_n7849_;
  assign new_n7851_ = new_n552_ & ~new_n7850_;
  assign new_n7852_ = new_n556_ & ~new_n7851_;
  assign new_n7853_ = new_n560_ & ~new_n7852_;
  assign new_n7854_ = new_n564_ & ~new_n7853_;
  assign new_n7855_ = new_n568_ & ~new_n7854_;
  assign new_n7856_ = new_n572_ & ~new_n7855_;
  assign new_n7857_ = new_n576_ & ~new_n7856_;
  assign new_n7858_ = new_n580_ & ~new_n7857_;
  assign new_n7859_ = new_n584_ & ~new_n7858_;
  assign new_n7860_ = \req[77]  & ~new_n586_;
  assign \grant[77]  = ~new_n7859_ & new_n7860_;
  assign new_n7862_ = new_n595_ & ~new_n930_;
  assign new_n7863_ = new_n600_ & ~new_n7862_;
  assign new_n7864_ = new_n604_ & ~new_n7863_;
  assign new_n7865_ = new_n608_ & ~new_n7864_;
  assign new_n7866_ = new_n612_ & ~new_n7865_;
  assign new_n7867_ = new_n616_ & ~new_n7866_;
  assign new_n7868_ = new_n620_ & ~new_n7867_;
  assign new_n7869_ = new_n624_ & ~new_n7868_;
  assign new_n7870_ = new_n628_ & ~new_n7869_;
  assign new_n7871_ = new_n632_ & ~new_n7870_;
  assign new_n7872_ = new_n636_ & ~new_n7871_;
  assign new_n7873_ = new_n640_ & ~new_n7872_;
  assign new_n7874_ = new_n644_ & ~new_n7873_;
  assign new_n7875_ = new_n648_ & ~new_n7874_;
  assign new_n7876_ = new_n652_ & ~new_n7875_;
  assign new_n7877_ = new_n656_ & ~new_n7876_;
  assign new_n7878_ = new_n660_ & ~new_n7877_;
  assign new_n7879_ = new_n664_ & ~new_n7878_;
  assign new_n7880_ = new_n668_ & ~new_n7879_;
  assign new_n7881_ = new_n672_ & ~new_n7880_;
  assign new_n7882_ = new_n676_ & ~new_n7881_;
  assign new_n7883_ = new_n680_ & ~new_n7882_;
  assign new_n7884_ = new_n684_ & ~new_n7883_;
  assign new_n7885_ = new_n688_ & ~new_n7884_;
  assign new_n7886_ = new_n692_ & ~new_n7885_;
  assign new_n7887_ = new_n696_ & ~new_n7886_;
  assign new_n7888_ = new_n700_ & ~new_n7887_;
  assign new_n7889_ = new_n704_ & ~new_n7888_;
  assign new_n7890_ = new_n708_ & ~new_n7889_;
  assign new_n7891_ = new_n712_ & ~new_n7890_;
  assign new_n7892_ = new_n716_ & ~new_n7891_;
  assign new_n7893_ = new_n720_ & ~new_n7892_;
  assign new_n7894_ = new_n1484_ & ~new_n7893_;
  assign new_n7895_ = new_n1486_ & ~new_n7894_;
  assign new_n7896_ = new_n1750_ & ~new_n7895_;
  assign new_n7897_ = new_n731_ & ~new_n7896_;
  assign new_n7898_ = new_n735_ & ~new_n7897_;
  assign new_n7899_ = new_n739_ & ~new_n7898_;
  assign new_n7900_ = new_n743_ & ~new_n7899_;
  assign new_n7901_ = new_n747_ & ~new_n7900_;
  assign new_n7902_ = new_n751_ & ~new_n7901_;
  assign new_n7903_ = new_n755_ & ~new_n7902_;
  assign new_n7904_ = new_n759_ & ~new_n7903_;
  assign new_n7905_ = new_n763_ & ~new_n7904_;
  assign new_n7906_ = new_n767_ & ~new_n7905_;
  assign new_n7907_ = new_n771_ & ~new_n7906_;
  assign new_n7908_ = new_n775_ & ~new_n7907_;
  assign new_n7909_ = new_n779_ & ~new_n7908_;
  assign new_n7910_ = new_n783_ & ~new_n7909_;
  assign new_n7911_ = new_n787_ & ~new_n7910_;
  assign new_n7912_ = new_n791_ & ~new_n7911_;
  assign new_n7913_ = new_n795_ & ~new_n7912_;
  assign new_n7914_ = new_n799_ & ~new_n7913_;
  assign new_n7915_ = new_n803_ & ~new_n7914_;
  assign new_n7916_ = new_n807_ & ~new_n7915_;
  assign new_n7917_ = new_n811_ & ~new_n7916_;
  assign new_n7918_ = new_n815_ & ~new_n7917_;
  assign new_n7919_ = new_n819_ & ~new_n7918_;
  assign new_n7920_ = new_n823_ & ~new_n7919_;
  assign new_n7921_ = new_n827_ & ~new_n7920_;
  assign new_n7922_ = new_n831_ & ~new_n7921_;
  assign new_n7923_ = new_n835_ & ~new_n7922_;
  assign new_n7924_ = new_n839_ & ~new_n7923_;
  assign new_n7925_ = new_n843_ & ~new_n7924_;
  assign new_n7926_ = new_n847_ & ~new_n7925_;
  assign new_n7927_ = new_n851_ & ~new_n7926_;
  assign new_n7928_ = new_n855_ & ~new_n7927_;
  assign new_n7929_ = new_n859_ & ~new_n7928_;
  assign new_n7930_ = new_n863_ & ~new_n7929_;
  assign new_n7931_ = new_n867_ & ~new_n7930_;
  assign new_n7932_ = new_n871_ & ~new_n7931_;
  assign new_n7933_ = new_n875_ & ~new_n7932_;
  assign new_n7934_ = new_n879_ & ~new_n7933_;
  assign new_n7935_ = new_n883_ & ~new_n7934_;
  assign new_n7936_ = new_n887_ & ~new_n7935_;
  assign new_n7937_ = new_n891_ & ~new_n7936_;
  assign new_n7938_ = new_n895_ & ~new_n7937_;
  assign new_n7939_ = new_n899_ & ~new_n7938_;
  assign new_n7940_ = new_n903_ & ~new_n7939_;
  assign new_n7941_ = new_n907_ & ~new_n7940_;
  assign new_n7942_ = new_n911_ & ~new_n7941_;
  assign new_n7943_ = new_n915_ & ~new_n7942_;
  assign new_n7944_ = new_n919_ & ~new_n7943_;
  assign new_n7945_ = new_n923_ & ~new_n7944_;
  assign new_n7946_ = \req[78]  & ~new_n925_;
  assign \grant[78]  = ~new_n7945_ & new_n7946_;
  assign new_n7948_ = new_n934_ & ~new_n1267_;
  assign new_n7949_ = new_n939_ & ~new_n7948_;
  assign new_n7950_ = new_n943_ & ~new_n7949_;
  assign new_n7951_ = new_n947_ & ~new_n7950_;
  assign new_n7952_ = new_n951_ & ~new_n7951_;
  assign new_n7953_ = new_n955_ & ~new_n7952_;
  assign new_n7954_ = new_n959_ & ~new_n7953_;
  assign new_n7955_ = new_n963_ & ~new_n7954_;
  assign new_n7956_ = new_n967_ & ~new_n7955_;
  assign new_n7957_ = new_n971_ & ~new_n7956_;
  assign new_n7958_ = new_n975_ & ~new_n7957_;
  assign new_n7959_ = new_n979_ & ~new_n7958_;
  assign new_n7960_ = new_n983_ & ~new_n7959_;
  assign new_n7961_ = new_n987_ & ~new_n7960_;
  assign new_n7962_ = new_n991_ & ~new_n7961_;
  assign new_n7963_ = new_n995_ & ~new_n7962_;
  assign new_n7964_ = new_n999_ & ~new_n7963_;
  assign new_n7965_ = new_n1003_ & ~new_n7964_;
  assign new_n7966_ = new_n1007_ & ~new_n7965_;
  assign new_n7967_ = new_n1011_ & ~new_n7966_;
  assign new_n7968_ = new_n1015_ & ~new_n7967_;
  assign new_n7969_ = new_n1019_ & ~new_n7968_;
  assign new_n7970_ = new_n1023_ & ~new_n7969_;
  assign new_n7971_ = new_n1027_ & ~new_n7970_;
  assign new_n7972_ = new_n1031_ & ~new_n7971_;
  assign new_n7973_ = new_n1035_ & ~new_n7972_;
  assign new_n7974_ = new_n1039_ & ~new_n7973_;
  assign new_n7975_ = new_n1043_ & ~new_n7974_;
  assign new_n7976_ = new_n1047_ & ~new_n7975_;
  assign new_n7977_ = new_n1051_ & ~new_n7976_;
  assign new_n7978_ = new_n1055_ & ~new_n7977_;
  assign new_n7979_ = new_n1059_ & ~new_n7978_;
  assign new_n7980_ = new_n1574_ & ~new_n7979_;
  assign new_n7981_ = new_n1576_ & ~new_n7980_;
  assign new_n7982_ = new_n1837_ & ~new_n7981_;
  assign new_n7983_ = new_n1068_ & ~new_n7982_;
  assign new_n7984_ = new_n1072_ & ~new_n7983_;
  assign new_n7985_ = new_n1076_ & ~new_n7984_;
  assign new_n7986_ = new_n1080_ & ~new_n7985_;
  assign new_n7987_ = new_n1084_ & ~new_n7986_;
  assign new_n7988_ = new_n1088_ & ~new_n7987_;
  assign new_n7989_ = new_n1092_ & ~new_n7988_;
  assign new_n7990_ = new_n1096_ & ~new_n7989_;
  assign new_n7991_ = new_n1100_ & ~new_n7990_;
  assign new_n7992_ = new_n1104_ & ~new_n7991_;
  assign new_n7993_ = new_n1108_ & ~new_n7992_;
  assign new_n7994_ = new_n1112_ & ~new_n7993_;
  assign new_n7995_ = new_n1116_ & ~new_n7994_;
  assign new_n7996_ = new_n1120_ & ~new_n7995_;
  assign new_n7997_ = new_n1124_ & ~new_n7996_;
  assign new_n7998_ = new_n1128_ & ~new_n7997_;
  assign new_n7999_ = new_n1132_ & ~new_n7998_;
  assign new_n8000_ = new_n1136_ & ~new_n7999_;
  assign new_n8001_ = new_n1140_ & ~new_n8000_;
  assign new_n8002_ = new_n1144_ & ~new_n8001_;
  assign new_n8003_ = new_n1148_ & ~new_n8002_;
  assign new_n8004_ = new_n1152_ & ~new_n8003_;
  assign new_n8005_ = new_n1156_ & ~new_n8004_;
  assign new_n8006_ = new_n1160_ & ~new_n8005_;
  assign new_n8007_ = new_n1164_ & ~new_n8006_;
  assign new_n8008_ = new_n1168_ & ~new_n8007_;
  assign new_n8009_ = new_n1172_ & ~new_n8008_;
  assign new_n8010_ = new_n1176_ & ~new_n8009_;
  assign new_n8011_ = new_n1180_ & ~new_n8010_;
  assign new_n8012_ = new_n1184_ & ~new_n8011_;
  assign new_n8013_ = new_n1188_ & ~new_n8012_;
  assign new_n8014_ = new_n1192_ & ~new_n8013_;
  assign new_n8015_ = new_n1196_ & ~new_n8014_;
  assign new_n8016_ = new_n1200_ & ~new_n8015_;
  assign new_n8017_ = new_n1204_ & ~new_n8016_;
  assign new_n8018_ = new_n1208_ & ~new_n8017_;
  assign new_n8019_ = new_n1212_ & ~new_n8018_;
  assign new_n8020_ = new_n1216_ & ~new_n8019_;
  assign new_n8021_ = new_n1220_ & ~new_n8020_;
  assign new_n8022_ = new_n1224_ & ~new_n8021_;
  assign new_n8023_ = new_n1228_ & ~new_n8022_;
  assign new_n8024_ = new_n1232_ & ~new_n8023_;
  assign new_n8025_ = new_n1236_ & ~new_n8024_;
  assign new_n8026_ = new_n1240_ & ~new_n8025_;
  assign new_n8027_ = new_n1244_ & ~new_n8026_;
  assign new_n8028_ = new_n1248_ & ~new_n8027_;
  assign new_n8029_ = new_n1252_ & ~new_n8028_;
  assign new_n8030_ = new_n1256_ & ~new_n8029_;
  assign new_n8031_ = new_n1260_ & ~new_n8030_;
  assign new_n8032_ = \req[79]  & ~new_n1262_;
  assign \grant[79]  = ~new_n8031_ & new_n8032_;
  assign new_n8034_ = ~new_n599_ & new_n1271_;
  assign new_n8035_ = new_n1276_ & ~new_n8034_;
  assign new_n8036_ = new_n1280_ & ~new_n8035_;
  assign new_n8037_ = new_n1284_ & ~new_n8036_;
  assign new_n8038_ = new_n1288_ & ~new_n8037_;
  assign new_n8039_ = new_n1292_ & ~new_n8038_;
  assign new_n8040_ = new_n1296_ & ~new_n8039_;
  assign new_n8041_ = new_n1300_ & ~new_n8040_;
  assign new_n8042_ = new_n1304_ & ~new_n8041_;
  assign new_n8043_ = new_n1308_ & ~new_n8042_;
  assign new_n8044_ = new_n1312_ & ~new_n8043_;
  assign new_n8045_ = new_n1316_ & ~new_n8044_;
  assign new_n8046_ = new_n1320_ & ~new_n8045_;
  assign new_n8047_ = new_n1324_ & ~new_n8046_;
  assign new_n8048_ = new_n1328_ & ~new_n8047_;
  assign new_n8049_ = new_n1332_ & ~new_n8048_;
  assign new_n8050_ = new_n1336_ & ~new_n8049_;
  assign new_n8051_ = new_n1340_ & ~new_n8050_;
  assign new_n8052_ = new_n1344_ & ~new_n8051_;
  assign new_n8053_ = new_n1348_ & ~new_n8052_;
  assign new_n8054_ = new_n1352_ & ~new_n8053_;
  assign new_n8055_ = new_n1356_ & ~new_n8054_;
  assign new_n8056_ = new_n1360_ & ~new_n8055_;
  assign new_n8057_ = new_n1364_ & ~new_n8056_;
  assign new_n8058_ = new_n1368_ & ~new_n8057_;
  assign new_n8059_ = new_n1372_ & ~new_n8058_;
  assign new_n8060_ = new_n1376_ & ~new_n8059_;
  assign new_n8061_ = new_n1380_ & ~new_n8060_;
  assign new_n8062_ = new_n1384_ & ~new_n8061_;
  assign new_n8063_ = new_n1388_ & ~new_n8062_;
  assign new_n8064_ = new_n1392_ & ~new_n8063_;
  assign new_n8065_ = new_n1396_ & ~new_n8064_;
  assign new_n8066_ = new_n1663_ & ~new_n8065_;
  assign new_n8067_ = new_n392_ & ~new_n8066_;
  assign new_n8068_ = new_n396_ & ~new_n8067_;
  assign new_n8069_ = new_n400_ & ~new_n8068_;
  assign new_n8070_ = new_n404_ & ~new_n8069_;
  assign new_n8071_ = new_n408_ & ~new_n8070_;
  assign new_n8072_ = new_n412_ & ~new_n8071_;
  assign new_n8073_ = new_n416_ & ~new_n8072_;
  assign new_n8074_ = new_n420_ & ~new_n8073_;
  assign new_n8075_ = new_n424_ & ~new_n8074_;
  assign new_n8076_ = new_n428_ & ~new_n8075_;
  assign new_n8077_ = new_n432_ & ~new_n8076_;
  assign new_n8078_ = new_n436_ & ~new_n8077_;
  assign new_n8079_ = new_n440_ & ~new_n8078_;
  assign new_n8080_ = new_n444_ & ~new_n8079_;
  assign new_n8081_ = new_n448_ & ~new_n8080_;
  assign new_n8082_ = new_n452_ & ~new_n8081_;
  assign new_n8083_ = new_n456_ & ~new_n8082_;
  assign new_n8084_ = new_n460_ & ~new_n8083_;
  assign new_n8085_ = new_n464_ & ~new_n8084_;
  assign new_n8086_ = new_n468_ & ~new_n8085_;
  assign new_n8087_ = new_n472_ & ~new_n8086_;
  assign new_n8088_ = new_n476_ & ~new_n8087_;
  assign new_n8089_ = new_n480_ & ~new_n8088_;
  assign new_n8090_ = new_n484_ & ~new_n8089_;
  assign new_n8091_ = new_n488_ & ~new_n8090_;
  assign new_n8092_ = new_n492_ & ~new_n8091_;
  assign new_n8093_ = new_n496_ & ~new_n8092_;
  assign new_n8094_ = new_n500_ & ~new_n8093_;
  assign new_n8095_ = new_n504_ & ~new_n8094_;
  assign new_n8096_ = new_n508_ & ~new_n8095_;
  assign new_n8097_ = new_n512_ & ~new_n8096_;
  assign new_n8098_ = new_n516_ & ~new_n8097_;
  assign new_n8099_ = new_n520_ & ~new_n8098_;
  assign new_n8100_ = new_n524_ & ~new_n8099_;
  assign new_n8101_ = new_n528_ & ~new_n8100_;
  assign new_n8102_ = new_n532_ & ~new_n8101_;
  assign new_n8103_ = new_n536_ & ~new_n8102_;
  assign new_n8104_ = new_n540_ & ~new_n8103_;
  assign new_n8105_ = new_n544_ & ~new_n8104_;
  assign new_n8106_ = new_n548_ & ~new_n8105_;
  assign new_n8107_ = new_n552_ & ~new_n8106_;
  assign new_n8108_ = new_n556_ & ~new_n8107_;
  assign new_n8109_ = new_n560_ & ~new_n8108_;
  assign new_n8110_ = new_n564_ & ~new_n8109_;
  assign new_n8111_ = new_n568_ & ~new_n8110_;
  assign new_n8112_ = new_n572_ & ~new_n8111_;
  assign new_n8113_ = new_n576_ & ~new_n8112_;
  assign new_n8114_ = new_n580_ & ~new_n8113_;
  assign new_n8115_ = new_n584_ & ~new_n8114_;
  assign new_n8116_ = new_n588_ & ~new_n8115_;
  assign new_n8117_ = new_n592_ & ~new_n8116_;
  assign new_n8118_ = \req[80]  & ~new_n594_;
  assign \grant[80]  = ~new_n8117_ & new_n8118_;
  assign new_n8120_ = new_n603_ & ~new_n938_;
  assign new_n8121_ = new_n608_ & ~new_n8120_;
  assign new_n8122_ = new_n612_ & ~new_n8121_;
  assign new_n8123_ = new_n616_ & ~new_n8122_;
  assign new_n8124_ = new_n620_ & ~new_n8123_;
  assign new_n8125_ = new_n624_ & ~new_n8124_;
  assign new_n8126_ = new_n628_ & ~new_n8125_;
  assign new_n8127_ = new_n632_ & ~new_n8126_;
  assign new_n8128_ = new_n636_ & ~new_n8127_;
  assign new_n8129_ = new_n640_ & ~new_n8128_;
  assign new_n8130_ = new_n644_ & ~new_n8129_;
  assign new_n8131_ = new_n648_ & ~new_n8130_;
  assign new_n8132_ = new_n652_ & ~new_n8131_;
  assign new_n8133_ = new_n656_ & ~new_n8132_;
  assign new_n8134_ = new_n660_ & ~new_n8133_;
  assign new_n8135_ = new_n664_ & ~new_n8134_;
  assign new_n8136_ = new_n668_ & ~new_n8135_;
  assign new_n8137_ = new_n672_ & ~new_n8136_;
  assign new_n8138_ = new_n676_ & ~new_n8137_;
  assign new_n8139_ = new_n680_ & ~new_n8138_;
  assign new_n8140_ = new_n684_ & ~new_n8139_;
  assign new_n8141_ = new_n688_ & ~new_n8140_;
  assign new_n8142_ = new_n692_ & ~new_n8141_;
  assign new_n8143_ = new_n696_ & ~new_n8142_;
  assign new_n8144_ = new_n700_ & ~new_n8143_;
  assign new_n8145_ = new_n704_ & ~new_n8144_;
  assign new_n8146_ = new_n708_ & ~new_n8145_;
  assign new_n8147_ = new_n712_ & ~new_n8146_;
  assign new_n8148_ = new_n716_ & ~new_n8147_;
  assign new_n8149_ = new_n720_ & ~new_n8148_;
  assign new_n8150_ = new_n1484_ & ~new_n8149_;
  assign new_n8151_ = new_n1486_ & ~new_n8150_;
  assign new_n8152_ = new_n1750_ & ~new_n8151_;
  assign new_n8153_ = new_n731_ & ~new_n8152_;
  assign new_n8154_ = new_n735_ & ~new_n8153_;
  assign new_n8155_ = new_n739_ & ~new_n8154_;
  assign new_n8156_ = new_n743_ & ~new_n8155_;
  assign new_n8157_ = new_n747_ & ~new_n8156_;
  assign new_n8158_ = new_n751_ & ~new_n8157_;
  assign new_n8159_ = new_n755_ & ~new_n8158_;
  assign new_n8160_ = new_n759_ & ~new_n8159_;
  assign new_n8161_ = new_n763_ & ~new_n8160_;
  assign new_n8162_ = new_n767_ & ~new_n8161_;
  assign new_n8163_ = new_n771_ & ~new_n8162_;
  assign new_n8164_ = new_n775_ & ~new_n8163_;
  assign new_n8165_ = new_n779_ & ~new_n8164_;
  assign new_n8166_ = new_n783_ & ~new_n8165_;
  assign new_n8167_ = new_n787_ & ~new_n8166_;
  assign new_n8168_ = new_n791_ & ~new_n8167_;
  assign new_n8169_ = new_n795_ & ~new_n8168_;
  assign new_n8170_ = new_n799_ & ~new_n8169_;
  assign new_n8171_ = new_n803_ & ~new_n8170_;
  assign new_n8172_ = new_n807_ & ~new_n8171_;
  assign new_n8173_ = new_n811_ & ~new_n8172_;
  assign new_n8174_ = new_n815_ & ~new_n8173_;
  assign new_n8175_ = new_n819_ & ~new_n8174_;
  assign new_n8176_ = new_n823_ & ~new_n8175_;
  assign new_n8177_ = new_n827_ & ~new_n8176_;
  assign new_n8178_ = new_n831_ & ~new_n8177_;
  assign new_n8179_ = new_n835_ & ~new_n8178_;
  assign new_n8180_ = new_n839_ & ~new_n8179_;
  assign new_n8181_ = new_n843_ & ~new_n8180_;
  assign new_n8182_ = new_n847_ & ~new_n8181_;
  assign new_n8183_ = new_n851_ & ~new_n8182_;
  assign new_n8184_ = new_n855_ & ~new_n8183_;
  assign new_n8185_ = new_n859_ & ~new_n8184_;
  assign new_n8186_ = new_n863_ & ~new_n8185_;
  assign new_n8187_ = new_n867_ & ~new_n8186_;
  assign new_n8188_ = new_n871_ & ~new_n8187_;
  assign new_n8189_ = new_n875_ & ~new_n8188_;
  assign new_n8190_ = new_n879_ & ~new_n8189_;
  assign new_n8191_ = new_n883_ & ~new_n8190_;
  assign new_n8192_ = new_n887_ & ~new_n8191_;
  assign new_n8193_ = new_n891_ & ~new_n8192_;
  assign new_n8194_ = new_n895_ & ~new_n8193_;
  assign new_n8195_ = new_n899_ & ~new_n8194_;
  assign new_n8196_ = new_n903_ & ~new_n8195_;
  assign new_n8197_ = new_n907_ & ~new_n8196_;
  assign new_n8198_ = new_n911_ & ~new_n8197_;
  assign new_n8199_ = new_n915_ & ~new_n8198_;
  assign new_n8200_ = new_n919_ & ~new_n8199_;
  assign new_n8201_ = new_n923_ & ~new_n8200_;
  assign new_n8202_ = new_n927_ & ~new_n8201_;
  assign new_n8203_ = new_n931_ & ~new_n8202_;
  assign new_n8204_ = \req[81]  & ~new_n933_;
  assign \grant[81]  = ~new_n8203_ & new_n8204_;
  assign new_n8206_ = new_n942_ & ~new_n1275_;
  assign new_n8207_ = new_n947_ & ~new_n8206_;
  assign new_n8208_ = new_n951_ & ~new_n8207_;
  assign new_n8209_ = new_n955_ & ~new_n8208_;
  assign new_n8210_ = new_n959_ & ~new_n8209_;
  assign new_n8211_ = new_n963_ & ~new_n8210_;
  assign new_n8212_ = new_n967_ & ~new_n8211_;
  assign new_n8213_ = new_n971_ & ~new_n8212_;
  assign new_n8214_ = new_n975_ & ~new_n8213_;
  assign new_n8215_ = new_n979_ & ~new_n8214_;
  assign new_n8216_ = new_n983_ & ~new_n8215_;
  assign new_n8217_ = new_n987_ & ~new_n8216_;
  assign new_n8218_ = new_n991_ & ~new_n8217_;
  assign new_n8219_ = new_n995_ & ~new_n8218_;
  assign new_n8220_ = new_n999_ & ~new_n8219_;
  assign new_n8221_ = new_n1003_ & ~new_n8220_;
  assign new_n8222_ = new_n1007_ & ~new_n8221_;
  assign new_n8223_ = new_n1011_ & ~new_n8222_;
  assign new_n8224_ = new_n1015_ & ~new_n8223_;
  assign new_n8225_ = new_n1019_ & ~new_n8224_;
  assign new_n8226_ = new_n1023_ & ~new_n8225_;
  assign new_n8227_ = new_n1027_ & ~new_n8226_;
  assign new_n8228_ = new_n1031_ & ~new_n8227_;
  assign new_n8229_ = new_n1035_ & ~new_n8228_;
  assign new_n8230_ = new_n1039_ & ~new_n8229_;
  assign new_n8231_ = new_n1043_ & ~new_n8230_;
  assign new_n8232_ = new_n1047_ & ~new_n8231_;
  assign new_n8233_ = new_n1051_ & ~new_n8232_;
  assign new_n8234_ = new_n1055_ & ~new_n8233_;
  assign new_n8235_ = new_n1059_ & ~new_n8234_;
  assign new_n8236_ = new_n1574_ & ~new_n8235_;
  assign new_n8237_ = new_n1576_ & ~new_n8236_;
  assign new_n8238_ = new_n1837_ & ~new_n8237_;
  assign new_n8239_ = new_n1068_ & ~new_n8238_;
  assign new_n8240_ = new_n1072_ & ~new_n8239_;
  assign new_n8241_ = new_n1076_ & ~new_n8240_;
  assign new_n8242_ = new_n1080_ & ~new_n8241_;
  assign new_n8243_ = new_n1084_ & ~new_n8242_;
  assign new_n8244_ = new_n1088_ & ~new_n8243_;
  assign new_n8245_ = new_n1092_ & ~new_n8244_;
  assign new_n8246_ = new_n1096_ & ~new_n8245_;
  assign new_n8247_ = new_n1100_ & ~new_n8246_;
  assign new_n8248_ = new_n1104_ & ~new_n8247_;
  assign new_n8249_ = new_n1108_ & ~new_n8248_;
  assign new_n8250_ = new_n1112_ & ~new_n8249_;
  assign new_n8251_ = new_n1116_ & ~new_n8250_;
  assign new_n8252_ = new_n1120_ & ~new_n8251_;
  assign new_n8253_ = new_n1124_ & ~new_n8252_;
  assign new_n8254_ = new_n1128_ & ~new_n8253_;
  assign new_n8255_ = new_n1132_ & ~new_n8254_;
  assign new_n8256_ = new_n1136_ & ~new_n8255_;
  assign new_n8257_ = new_n1140_ & ~new_n8256_;
  assign new_n8258_ = new_n1144_ & ~new_n8257_;
  assign new_n8259_ = new_n1148_ & ~new_n8258_;
  assign new_n8260_ = new_n1152_ & ~new_n8259_;
  assign new_n8261_ = new_n1156_ & ~new_n8260_;
  assign new_n8262_ = new_n1160_ & ~new_n8261_;
  assign new_n8263_ = new_n1164_ & ~new_n8262_;
  assign new_n8264_ = new_n1168_ & ~new_n8263_;
  assign new_n8265_ = new_n1172_ & ~new_n8264_;
  assign new_n8266_ = new_n1176_ & ~new_n8265_;
  assign new_n8267_ = new_n1180_ & ~new_n8266_;
  assign new_n8268_ = new_n1184_ & ~new_n8267_;
  assign new_n8269_ = new_n1188_ & ~new_n8268_;
  assign new_n8270_ = new_n1192_ & ~new_n8269_;
  assign new_n8271_ = new_n1196_ & ~new_n8270_;
  assign new_n8272_ = new_n1200_ & ~new_n8271_;
  assign new_n8273_ = new_n1204_ & ~new_n8272_;
  assign new_n8274_ = new_n1208_ & ~new_n8273_;
  assign new_n8275_ = new_n1212_ & ~new_n8274_;
  assign new_n8276_ = new_n1216_ & ~new_n8275_;
  assign new_n8277_ = new_n1220_ & ~new_n8276_;
  assign new_n8278_ = new_n1224_ & ~new_n8277_;
  assign new_n8279_ = new_n1228_ & ~new_n8278_;
  assign new_n8280_ = new_n1232_ & ~new_n8279_;
  assign new_n8281_ = new_n1236_ & ~new_n8280_;
  assign new_n8282_ = new_n1240_ & ~new_n8281_;
  assign new_n8283_ = new_n1244_ & ~new_n8282_;
  assign new_n8284_ = new_n1248_ & ~new_n8283_;
  assign new_n8285_ = new_n1252_ & ~new_n8284_;
  assign new_n8286_ = new_n1256_ & ~new_n8285_;
  assign new_n8287_ = new_n1260_ & ~new_n8286_;
  assign new_n8288_ = new_n1264_ & ~new_n8287_;
  assign new_n8289_ = new_n1268_ & ~new_n8288_;
  assign new_n8290_ = \req[82]  & ~new_n1270_;
  assign \grant[82]  = ~new_n8289_ & new_n8290_;
  assign new_n8292_ = ~new_n607_ & new_n1279_;
  assign new_n8293_ = new_n1284_ & ~new_n8292_;
  assign new_n8294_ = new_n1288_ & ~new_n8293_;
  assign new_n8295_ = new_n1292_ & ~new_n8294_;
  assign new_n8296_ = new_n1296_ & ~new_n8295_;
  assign new_n8297_ = new_n1300_ & ~new_n8296_;
  assign new_n8298_ = new_n1304_ & ~new_n8297_;
  assign new_n8299_ = new_n1308_ & ~new_n8298_;
  assign new_n8300_ = new_n1312_ & ~new_n8299_;
  assign new_n8301_ = new_n1316_ & ~new_n8300_;
  assign new_n8302_ = new_n1320_ & ~new_n8301_;
  assign new_n8303_ = new_n1324_ & ~new_n8302_;
  assign new_n8304_ = new_n1328_ & ~new_n8303_;
  assign new_n8305_ = new_n1332_ & ~new_n8304_;
  assign new_n8306_ = new_n1336_ & ~new_n8305_;
  assign new_n8307_ = new_n1340_ & ~new_n8306_;
  assign new_n8308_ = new_n1344_ & ~new_n8307_;
  assign new_n8309_ = new_n1348_ & ~new_n8308_;
  assign new_n8310_ = new_n1352_ & ~new_n8309_;
  assign new_n8311_ = new_n1356_ & ~new_n8310_;
  assign new_n8312_ = new_n1360_ & ~new_n8311_;
  assign new_n8313_ = new_n1364_ & ~new_n8312_;
  assign new_n8314_ = new_n1368_ & ~new_n8313_;
  assign new_n8315_ = new_n1372_ & ~new_n8314_;
  assign new_n8316_ = new_n1376_ & ~new_n8315_;
  assign new_n8317_ = new_n1380_ & ~new_n8316_;
  assign new_n8318_ = new_n1384_ & ~new_n8317_;
  assign new_n8319_ = new_n1388_ & ~new_n8318_;
  assign new_n8320_ = new_n1392_ & ~new_n8319_;
  assign new_n8321_ = new_n1396_ & ~new_n8320_;
  assign new_n8322_ = new_n1663_ & ~new_n8321_;
  assign new_n8323_ = new_n392_ & ~new_n8322_;
  assign new_n8324_ = new_n396_ & ~new_n8323_;
  assign new_n8325_ = new_n400_ & ~new_n8324_;
  assign new_n8326_ = new_n404_ & ~new_n8325_;
  assign new_n8327_ = new_n408_ & ~new_n8326_;
  assign new_n8328_ = new_n412_ & ~new_n8327_;
  assign new_n8329_ = new_n416_ & ~new_n8328_;
  assign new_n8330_ = new_n420_ & ~new_n8329_;
  assign new_n8331_ = new_n424_ & ~new_n8330_;
  assign new_n8332_ = new_n428_ & ~new_n8331_;
  assign new_n8333_ = new_n432_ & ~new_n8332_;
  assign new_n8334_ = new_n436_ & ~new_n8333_;
  assign new_n8335_ = new_n440_ & ~new_n8334_;
  assign new_n8336_ = new_n444_ & ~new_n8335_;
  assign new_n8337_ = new_n448_ & ~new_n8336_;
  assign new_n8338_ = new_n452_ & ~new_n8337_;
  assign new_n8339_ = new_n456_ & ~new_n8338_;
  assign new_n8340_ = new_n460_ & ~new_n8339_;
  assign new_n8341_ = new_n464_ & ~new_n8340_;
  assign new_n8342_ = new_n468_ & ~new_n8341_;
  assign new_n8343_ = new_n472_ & ~new_n8342_;
  assign new_n8344_ = new_n476_ & ~new_n8343_;
  assign new_n8345_ = new_n480_ & ~new_n8344_;
  assign new_n8346_ = new_n484_ & ~new_n8345_;
  assign new_n8347_ = new_n488_ & ~new_n8346_;
  assign new_n8348_ = new_n492_ & ~new_n8347_;
  assign new_n8349_ = new_n496_ & ~new_n8348_;
  assign new_n8350_ = new_n500_ & ~new_n8349_;
  assign new_n8351_ = new_n504_ & ~new_n8350_;
  assign new_n8352_ = new_n508_ & ~new_n8351_;
  assign new_n8353_ = new_n512_ & ~new_n8352_;
  assign new_n8354_ = new_n516_ & ~new_n8353_;
  assign new_n8355_ = new_n520_ & ~new_n8354_;
  assign new_n8356_ = new_n524_ & ~new_n8355_;
  assign new_n8357_ = new_n528_ & ~new_n8356_;
  assign new_n8358_ = new_n532_ & ~new_n8357_;
  assign new_n8359_ = new_n536_ & ~new_n8358_;
  assign new_n8360_ = new_n540_ & ~new_n8359_;
  assign new_n8361_ = new_n544_ & ~new_n8360_;
  assign new_n8362_ = new_n548_ & ~new_n8361_;
  assign new_n8363_ = new_n552_ & ~new_n8362_;
  assign new_n8364_ = new_n556_ & ~new_n8363_;
  assign new_n8365_ = new_n560_ & ~new_n8364_;
  assign new_n8366_ = new_n564_ & ~new_n8365_;
  assign new_n8367_ = new_n568_ & ~new_n8366_;
  assign new_n8368_ = new_n572_ & ~new_n8367_;
  assign new_n8369_ = new_n576_ & ~new_n8368_;
  assign new_n8370_ = new_n580_ & ~new_n8369_;
  assign new_n8371_ = new_n584_ & ~new_n8370_;
  assign new_n8372_ = new_n588_ & ~new_n8371_;
  assign new_n8373_ = new_n592_ & ~new_n8372_;
  assign new_n8374_ = new_n596_ & ~new_n8373_;
  assign new_n8375_ = new_n600_ & ~new_n8374_;
  assign new_n8376_ = \req[83]  & ~new_n602_;
  assign \grant[83]  = ~new_n8375_ & new_n8376_;
  assign new_n8378_ = new_n611_ & ~new_n946_;
  assign new_n8379_ = new_n616_ & ~new_n8378_;
  assign new_n8380_ = new_n620_ & ~new_n8379_;
  assign new_n8381_ = new_n624_ & ~new_n8380_;
  assign new_n8382_ = new_n628_ & ~new_n8381_;
  assign new_n8383_ = new_n632_ & ~new_n8382_;
  assign new_n8384_ = new_n636_ & ~new_n8383_;
  assign new_n8385_ = new_n640_ & ~new_n8384_;
  assign new_n8386_ = new_n644_ & ~new_n8385_;
  assign new_n8387_ = new_n648_ & ~new_n8386_;
  assign new_n8388_ = new_n652_ & ~new_n8387_;
  assign new_n8389_ = new_n656_ & ~new_n8388_;
  assign new_n8390_ = new_n660_ & ~new_n8389_;
  assign new_n8391_ = new_n664_ & ~new_n8390_;
  assign new_n8392_ = new_n668_ & ~new_n8391_;
  assign new_n8393_ = new_n672_ & ~new_n8392_;
  assign new_n8394_ = new_n676_ & ~new_n8393_;
  assign new_n8395_ = new_n680_ & ~new_n8394_;
  assign new_n8396_ = new_n684_ & ~new_n8395_;
  assign new_n8397_ = new_n688_ & ~new_n8396_;
  assign new_n8398_ = new_n692_ & ~new_n8397_;
  assign new_n8399_ = new_n696_ & ~new_n8398_;
  assign new_n8400_ = new_n700_ & ~new_n8399_;
  assign new_n8401_ = new_n704_ & ~new_n8400_;
  assign new_n8402_ = new_n708_ & ~new_n8401_;
  assign new_n8403_ = new_n712_ & ~new_n8402_;
  assign new_n8404_ = new_n716_ & ~new_n8403_;
  assign new_n8405_ = new_n720_ & ~new_n8404_;
  assign new_n8406_ = new_n1484_ & ~new_n8405_;
  assign new_n8407_ = new_n1486_ & ~new_n8406_;
  assign new_n8408_ = new_n1750_ & ~new_n8407_;
  assign new_n8409_ = new_n731_ & ~new_n8408_;
  assign new_n8410_ = new_n735_ & ~new_n8409_;
  assign new_n8411_ = new_n739_ & ~new_n8410_;
  assign new_n8412_ = new_n743_ & ~new_n8411_;
  assign new_n8413_ = new_n747_ & ~new_n8412_;
  assign new_n8414_ = new_n751_ & ~new_n8413_;
  assign new_n8415_ = new_n755_ & ~new_n8414_;
  assign new_n8416_ = new_n759_ & ~new_n8415_;
  assign new_n8417_ = new_n763_ & ~new_n8416_;
  assign new_n8418_ = new_n767_ & ~new_n8417_;
  assign new_n8419_ = new_n771_ & ~new_n8418_;
  assign new_n8420_ = new_n775_ & ~new_n8419_;
  assign new_n8421_ = new_n779_ & ~new_n8420_;
  assign new_n8422_ = new_n783_ & ~new_n8421_;
  assign new_n8423_ = new_n787_ & ~new_n8422_;
  assign new_n8424_ = new_n791_ & ~new_n8423_;
  assign new_n8425_ = new_n795_ & ~new_n8424_;
  assign new_n8426_ = new_n799_ & ~new_n8425_;
  assign new_n8427_ = new_n803_ & ~new_n8426_;
  assign new_n8428_ = new_n807_ & ~new_n8427_;
  assign new_n8429_ = new_n811_ & ~new_n8428_;
  assign new_n8430_ = new_n815_ & ~new_n8429_;
  assign new_n8431_ = new_n819_ & ~new_n8430_;
  assign new_n8432_ = new_n823_ & ~new_n8431_;
  assign new_n8433_ = new_n827_ & ~new_n8432_;
  assign new_n8434_ = new_n831_ & ~new_n8433_;
  assign new_n8435_ = new_n835_ & ~new_n8434_;
  assign new_n8436_ = new_n839_ & ~new_n8435_;
  assign new_n8437_ = new_n843_ & ~new_n8436_;
  assign new_n8438_ = new_n847_ & ~new_n8437_;
  assign new_n8439_ = new_n851_ & ~new_n8438_;
  assign new_n8440_ = new_n855_ & ~new_n8439_;
  assign new_n8441_ = new_n859_ & ~new_n8440_;
  assign new_n8442_ = new_n863_ & ~new_n8441_;
  assign new_n8443_ = new_n867_ & ~new_n8442_;
  assign new_n8444_ = new_n871_ & ~new_n8443_;
  assign new_n8445_ = new_n875_ & ~new_n8444_;
  assign new_n8446_ = new_n879_ & ~new_n8445_;
  assign new_n8447_ = new_n883_ & ~new_n8446_;
  assign new_n8448_ = new_n887_ & ~new_n8447_;
  assign new_n8449_ = new_n891_ & ~new_n8448_;
  assign new_n8450_ = new_n895_ & ~new_n8449_;
  assign new_n8451_ = new_n899_ & ~new_n8450_;
  assign new_n8452_ = new_n903_ & ~new_n8451_;
  assign new_n8453_ = new_n907_ & ~new_n8452_;
  assign new_n8454_ = new_n911_ & ~new_n8453_;
  assign new_n8455_ = new_n915_ & ~new_n8454_;
  assign new_n8456_ = new_n919_ & ~new_n8455_;
  assign new_n8457_ = new_n923_ & ~new_n8456_;
  assign new_n8458_ = new_n927_ & ~new_n8457_;
  assign new_n8459_ = new_n931_ & ~new_n8458_;
  assign new_n8460_ = new_n935_ & ~new_n8459_;
  assign new_n8461_ = new_n939_ & ~new_n8460_;
  assign new_n8462_ = \req[84]  & ~new_n941_;
  assign \grant[84]  = ~new_n8461_ & new_n8462_;
  assign new_n8464_ = new_n950_ & ~new_n1283_;
  assign new_n8465_ = new_n955_ & ~new_n8464_;
  assign new_n8466_ = new_n959_ & ~new_n8465_;
  assign new_n8467_ = new_n963_ & ~new_n8466_;
  assign new_n8468_ = new_n967_ & ~new_n8467_;
  assign new_n8469_ = new_n971_ & ~new_n8468_;
  assign new_n8470_ = new_n975_ & ~new_n8469_;
  assign new_n8471_ = new_n979_ & ~new_n8470_;
  assign new_n8472_ = new_n983_ & ~new_n8471_;
  assign new_n8473_ = new_n987_ & ~new_n8472_;
  assign new_n8474_ = new_n991_ & ~new_n8473_;
  assign new_n8475_ = new_n995_ & ~new_n8474_;
  assign new_n8476_ = new_n999_ & ~new_n8475_;
  assign new_n8477_ = new_n1003_ & ~new_n8476_;
  assign new_n8478_ = new_n1007_ & ~new_n8477_;
  assign new_n8479_ = new_n1011_ & ~new_n8478_;
  assign new_n8480_ = new_n1015_ & ~new_n8479_;
  assign new_n8481_ = new_n1019_ & ~new_n8480_;
  assign new_n8482_ = new_n1023_ & ~new_n8481_;
  assign new_n8483_ = new_n1027_ & ~new_n8482_;
  assign new_n8484_ = new_n1031_ & ~new_n8483_;
  assign new_n8485_ = new_n1035_ & ~new_n8484_;
  assign new_n8486_ = new_n1039_ & ~new_n8485_;
  assign new_n8487_ = new_n1043_ & ~new_n8486_;
  assign new_n8488_ = new_n1047_ & ~new_n8487_;
  assign new_n8489_ = new_n1051_ & ~new_n8488_;
  assign new_n8490_ = new_n1055_ & ~new_n8489_;
  assign new_n8491_ = new_n1059_ & ~new_n8490_;
  assign new_n8492_ = new_n1574_ & ~new_n8491_;
  assign new_n8493_ = new_n1576_ & ~new_n8492_;
  assign new_n8494_ = new_n1837_ & ~new_n8493_;
  assign new_n8495_ = new_n1068_ & ~new_n8494_;
  assign new_n8496_ = new_n1072_ & ~new_n8495_;
  assign new_n8497_ = new_n1076_ & ~new_n8496_;
  assign new_n8498_ = new_n1080_ & ~new_n8497_;
  assign new_n8499_ = new_n1084_ & ~new_n8498_;
  assign new_n8500_ = new_n1088_ & ~new_n8499_;
  assign new_n8501_ = new_n1092_ & ~new_n8500_;
  assign new_n8502_ = new_n1096_ & ~new_n8501_;
  assign new_n8503_ = new_n1100_ & ~new_n8502_;
  assign new_n8504_ = new_n1104_ & ~new_n8503_;
  assign new_n8505_ = new_n1108_ & ~new_n8504_;
  assign new_n8506_ = new_n1112_ & ~new_n8505_;
  assign new_n8507_ = new_n1116_ & ~new_n8506_;
  assign new_n8508_ = new_n1120_ & ~new_n8507_;
  assign new_n8509_ = new_n1124_ & ~new_n8508_;
  assign new_n8510_ = new_n1128_ & ~new_n8509_;
  assign new_n8511_ = new_n1132_ & ~new_n8510_;
  assign new_n8512_ = new_n1136_ & ~new_n8511_;
  assign new_n8513_ = new_n1140_ & ~new_n8512_;
  assign new_n8514_ = new_n1144_ & ~new_n8513_;
  assign new_n8515_ = new_n1148_ & ~new_n8514_;
  assign new_n8516_ = new_n1152_ & ~new_n8515_;
  assign new_n8517_ = new_n1156_ & ~new_n8516_;
  assign new_n8518_ = new_n1160_ & ~new_n8517_;
  assign new_n8519_ = new_n1164_ & ~new_n8518_;
  assign new_n8520_ = new_n1168_ & ~new_n8519_;
  assign new_n8521_ = new_n1172_ & ~new_n8520_;
  assign new_n8522_ = new_n1176_ & ~new_n8521_;
  assign new_n8523_ = new_n1180_ & ~new_n8522_;
  assign new_n8524_ = new_n1184_ & ~new_n8523_;
  assign new_n8525_ = new_n1188_ & ~new_n8524_;
  assign new_n8526_ = new_n1192_ & ~new_n8525_;
  assign new_n8527_ = new_n1196_ & ~new_n8526_;
  assign new_n8528_ = new_n1200_ & ~new_n8527_;
  assign new_n8529_ = new_n1204_ & ~new_n8528_;
  assign new_n8530_ = new_n1208_ & ~new_n8529_;
  assign new_n8531_ = new_n1212_ & ~new_n8530_;
  assign new_n8532_ = new_n1216_ & ~new_n8531_;
  assign new_n8533_ = new_n1220_ & ~new_n8532_;
  assign new_n8534_ = new_n1224_ & ~new_n8533_;
  assign new_n8535_ = new_n1228_ & ~new_n8534_;
  assign new_n8536_ = new_n1232_ & ~new_n8535_;
  assign new_n8537_ = new_n1236_ & ~new_n8536_;
  assign new_n8538_ = new_n1240_ & ~new_n8537_;
  assign new_n8539_ = new_n1244_ & ~new_n8538_;
  assign new_n8540_ = new_n1248_ & ~new_n8539_;
  assign new_n8541_ = new_n1252_ & ~new_n8540_;
  assign new_n8542_ = new_n1256_ & ~new_n8541_;
  assign new_n8543_ = new_n1260_ & ~new_n8542_;
  assign new_n8544_ = new_n1264_ & ~new_n8543_;
  assign new_n8545_ = new_n1268_ & ~new_n8544_;
  assign new_n8546_ = new_n1272_ & ~new_n8545_;
  assign new_n8547_ = new_n1276_ & ~new_n8546_;
  assign new_n8548_ = \req[85]  & ~new_n1278_;
  assign \grant[85]  = ~new_n8547_ & new_n8548_;
  assign new_n8550_ = ~new_n615_ & new_n1287_;
  assign new_n8551_ = new_n1292_ & ~new_n8550_;
  assign new_n8552_ = new_n1296_ & ~new_n8551_;
  assign new_n8553_ = new_n1300_ & ~new_n8552_;
  assign new_n8554_ = new_n1304_ & ~new_n8553_;
  assign new_n8555_ = new_n1308_ & ~new_n8554_;
  assign new_n8556_ = new_n1312_ & ~new_n8555_;
  assign new_n8557_ = new_n1316_ & ~new_n8556_;
  assign new_n8558_ = new_n1320_ & ~new_n8557_;
  assign new_n8559_ = new_n1324_ & ~new_n8558_;
  assign new_n8560_ = new_n1328_ & ~new_n8559_;
  assign new_n8561_ = new_n1332_ & ~new_n8560_;
  assign new_n8562_ = new_n1336_ & ~new_n8561_;
  assign new_n8563_ = new_n1340_ & ~new_n8562_;
  assign new_n8564_ = new_n1344_ & ~new_n8563_;
  assign new_n8565_ = new_n1348_ & ~new_n8564_;
  assign new_n8566_ = new_n1352_ & ~new_n8565_;
  assign new_n8567_ = new_n1356_ & ~new_n8566_;
  assign new_n8568_ = new_n1360_ & ~new_n8567_;
  assign new_n8569_ = new_n1364_ & ~new_n8568_;
  assign new_n8570_ = new_n1368_ & ~new_n8569_;
  assign new_n8571_ = new_n1372_ & ~new_n8570_;
  assign new_n8572_ = new_n1376_ & ~new_n8571_;
  assign new_n8573_ = new_n1380_ & ~new_n8572_;
  assign new_n8574_ = new_n1384_ & ~new_n8573_;
  assign new_n8575_ = new_n1388_ & ~new_n8574_;
  assign new_n8576_ = new_n1392_ & ~new_n8575_;
  assign new_n8577_ = new_n1396_ & ~new_n8576_;
  assign new_n8578_ = new_n1663_ & ~new_n8577_;
  assign new_n8579_ = new_n392_ & ~new_n8578_;
  assign new_n8580_ = new_n396_ & ~new_n8579_;
  assign new_n8581_ = new_n400_ & ~new_n8580_;
  assign new_n8582_ = new_n404_ & ~new_n8581_;
  assign new_n8583_ = new_n408_ & ~new_n8582_;
  assign new_n8584_ = new_n412_ & ~new_n8583_;
  assign new_n8585_ = new_n416_ & ~new_n8584_;
  assign new_n8586_ = new_n420_ & ~new_n8585_;
  assign new_n8587_ = new_n424_ & ~new_n8586_;
  assign new_n8588_ = new_n428_ & ~new_n8587_;
  assign new_n8589_ = new_n432_ & ~new_n8588_;
  assign new_n8590_ = new_n436_ & ~new_n8589_;
  assign new_n8591_ = new_n440_ & ~new_n8590_;
  assign new_n8592_ = new_n444_ & ~new_n8591_;
  assign new_n8593_ = new_n448_ & ~new_n8592_;
  assign new_n8594_ = new_n452_ & ~new_n8593_;
  assign new_n8595_ = new_n456_ & ~new_n8594_;
  assign new_n8596_ = new_n460_ & ~new_n8595_;
  assign new_n8597_ = new_n464_ & ~new_n8596_;
  assign new_n8598_ = new_n468_ & ~new_n8597_;
  assign new_n8599_ = new_n472_ & ~new_n8598_;
  assign new_n8600_ = new_n476_ & ~new_n8599_;
  assign new_n8601_ = new_n480_ & ~new_n8600_;
  assign new_n8602_ = new_n484_ & ~new_n8601_;
  assign new_n8603_ = new_n488_ & ~new_n8602_;
  assign new_n8604_ = new_n492_ & ~new_n8603_;
  assign new_n8605_ = new_n496_ & ~new_n8604_;
  assign new_n8606_ = new_n500_ & ~new_n8605_;
  assign new_n8607_ = new_n504_ & ~new_n8606_;
  assign new_n8608_ = new_n508_ & ~new_n8607_;
  assign new_n8609_ = new_n512_ & ~new_n8608_;
  assign new_n8610_ = new_n516_ & ~new_n8609_;
  assign new_n8611_ = new_n520_ & ~new_n8610_;
  assign new_n8612_ = new_n524_ & ~new_n8611_;
  assign new_n8613_ = new_n528_ & ~new_n8612_;
  assign new_n8614_ = new_n532_ & ~new_n8613_;
  assign new_n8615_ = new_n536_ & ~new_n8614_;
  assign new_n8616_ = new_n540_ & ~new_n8615_;
  assign new_n8617_ = new_n544_ & ~new_n8616_;
  assign new_n8618_ = new_n548_ & ~new_n8617_;
  assign new_n8619_ = new_n552_ & ~new_n8618_;
  assign new_n8620_ = new_n556_ & ~new_n8619_;
  assign new_n8621_ = new_n560_ & ~new_n8620_;
  assign new_n8622_ = new_n564_ & ~new_n8621_;
  assign new_n8623_ = new_n568_ & ~new_n8622_;
  assign new_n8624_ = new_n572_ & ~new_n8623_;
  assign new_n8625_ = new_n576_ & ~new_n8624_;
  assign new_n8626_ = new_n580_ & ~new_n8625_;
  assign new_n8627_ = new_n584_ & ~new_n8626_;
  assign new_n8628_ = new_n588_ & ~new_n8627_;
  assign new_n8629_ = new_n592_ & ~new_n8628_;
  assign new_n8630_ = new_n596_ & ~new_n8629_;
  assign new_n8631_ = new_n600_ & ~new_n8630_;
  assign new_n8632_ = new_n604_ & ~new_n8631_;
  assign new_n8633_ = new_n608_ & ~new_n8632_;
  assign new_n8634_ = \req[86]  & ~new_n610_;
  assign \grant[86]  = ~new_n8633_ & new_n8634_;
  assign new_n8636_ = new_n619_ & ~new_n954_;
  assign new_n8637_ = new_n624_ & ~new_n8636_;
  assign new_n8638_ = new_n628_ & ~new_n8637_;
  assign new_n8639_ = new_n632_ & ~new_n8638_;
  assign new_n8640_ = new_n636_ & ~new_n8639_;
  assign new_n8641_ = new_n640_ & ~new_n8640_;
  assign new_n8642_ = new_n644_ & ~new_n8641_;
  assign new_n8643_ = new_n648_ & ~new_n8642_;
  assign new_n8644_ = new_n652_ & ~new_n8643_;
  assign new_n8645_ = new_n656_ & ~new_n8644_;
  assign new_n8646_ = new_n660_ & ~new_n8645_;
  assign new_n8647_ = new_n664_ & ~new_n8646_;
  assign new_n8648_ = new_n668_ & ~new_n8647_;
  assign new_n8649_ = new_n672_ & ~new_n8648_;
  assign new_n8650_ = new_n676_ & ~new_n8649_;
  assign new_n8651_ = new_n680_ & ~new_n8650_;
  assign new_n8652_ = new_n684_ & ~new_n8651_;
  assign new_n8653_ = new_n688_ & ~new_n8652_;
  assign new_n8654_ = new_n692_ & ~new_n8653_;
  assign new_n8655_ = new_n696_ & ~new_n8654_;
  assign new_n8656_ = new_n700_ & ~new_n8655_;
  assign new_n8657_ = new_n704_ & ~new_n8656_;
  assign new_n8658_ = new_n708_ & ~new_n8657_;
  assign new_n8659_ = new_n712_ & ~new_n8658_;
  assign new_n8660_ = new_n716_ & ~new_n8659_;
  assign new_n8661_ = new_n720_ & ~new_n8660_;
  assign new_n8662_ = new_n1484_ & ~new_n8661_;
  assign new_n8663_ = new_n1486_ & ~new_n8662_;
  assign new_n8664_ = new_n1750_ & ~new_n8663_;
  assign new_n8665_ = new_n731_ & ~new_n8664_;
  assign new_n8666_ = new_n735_ & ~new_n8665_;
  assign new_n8667_ = new_n739_ & ~new_n8666_;
  assign new_n8668_ = new_n743_ & ~new_n8667_;
  assign new_n8669_ = new_n747_ & ~new_n8668_;
  assign new_n8670_ = new_n751_ & ~new_n8669_;
  assign new_n8671_ = new_n755_ & ~new_n8670_;
  assign new_n8672_ = new_n759_ & ~new_n8671_;
  assign new_n8673_ = new_n763_ & ~new_n8672_;
  assign new_n8674_ = new_n767_ & ~new_n8673_;
  assign new_n8675_ = new_n771_ & ~new_n8674_;
  assign new_n8676_ = new_n775_ & ~new_n8675_;
  assign new_n8677_ = new_n779_ & ~new_n8676_;
  assign new_n8678_ = new_n783_ & ~new_n8677_;
  assign new_n8679_ = new_n787_ & ~new_n8678_;
  assign new_n8680_ = new_n791_ & ~new_n8679_;
  assign new_n8681_ = new_n795_ & ~new_n8680_;
  assign new_n8682_ = new_n799_ & ~new_n8681_;
  assign new_n8683_ = new_n803_ & ~new_n8682_;
  assign new_n8684_ = new_n807_ & ~new_n8683_;
  assign new_n8685_ = new_n811_ & ~new_n8684_;
  assign new_n8686_ = new_n815_ & ~new_n8685_;
  assign new_n8687_ = new_n819_ & ~new_n8686_;
  assign new_n8688_ = new_n823_ & ~new_n8687_;
  assign new_n8689_ = new_n827_ & ~new_n8688_;
  assign new_n8690_ = new_n831_ & ~new_n8689_;
  assign new_n8691_ = new_n835_ & ~new_n8690_;
  assign new_n8692_ = new_n839_ & ~new_n8691_;
  assign new_n8693_ = new_n843_ & ~new_n8692_;
  assign new_n8694_ = new_n847_ & ~new_n8693_;
  assign new_n8695_ = new_n851_ & ~new_n8694_;
  assign new_n8696_ = new_n855_ & ~new_n8695_;
  assign new_n8697_ = new_n859_ & ~new_n8696_;
  assign new_n8698_ = new_n863_ & ~new_n8697_;
  assign new_n8699_ = new_n867_ & ~new_n8698_;
  assign new_n8700_ = new_n871_ & ~new_n8699_;
  assign new_n8701_ = new_n875_ & ~new_n8700_;
  assign new_n8702_ = new_n879_ & ~new_n8701_;
  assign new_n8703_ = new_n883_ & ~new_n8702_;
  assign new_n8704_ = new_n887_ & ~new_n8703_;
  assign new_n8705_ = new_n891_ & ~new_n8704_;
  assign new_n8706_ = new_n895_ & ~new_n8705_;
  assign new_n8707_ = new_n899_ & ~new_n8706_;
  assign new_n8708_ = new_n903_ & ~new_n8707_;
  assign new_n8709_ = new_n907_ & ~new_n8708_;
  assign new_n8710_ = new_n911_ & ~new_n8709_;
  assign new_n8711_ = new_n915_ & ~new_n8710_;
  assign new_n8712_ = new_n919_ & ~new_n8711_;
  assign new_n8713_ = new_n923_ & ~new_n8712_;
  assign new_n8714_ = new_n927_ & ~new_n8713_;
  assign new_n8715_ = new_n931_ & ~new_n8714_;
  assign new_n8716_ = new_n935_ & ~new_n8715_;
  assign new_n8717_ = new_n939_ & ~new_n8716_;
  assign new_n8718_ = new_n943_ & ~new_n8717_;
  assign new_n8719_ = new_n947_ & ~new_n8718_;
  assign new_n8720_ = \req[87]  & ~new_n949_;
  assign \grant[87]  = ~new_n8719_ & new_n8720_;
  assign new_n8722_ = new_n958_ & ~new_n1291_;
  assign new_n8723_ = new_n963_ & ~new_n8722_;
  assign new_n8724_ = new_n967_ & ~new_n8723_;
  assign new_n8725_ = new_n971_ & ~new_n8724_;
  assign new_n8726_ = new_n975_ & ~new_n8725_;
  assign new_n8727_ = new_n979_ & ~new_n8726_;
  assign new_n8728_ = new_n983_ & ~new_n8727_;
  assign new_n8729_ = new_n987_ & ~new_n8728_;
  assign new_n8730_ = new_n991_ & ~new_n8729_;
  assign new_n8731_ = new_n995_ & ~new_n8730_;
  assign new_n8732_ = new_n999_ & ~new_n8731_;
  assign new_n8733_ = new_n1003_ & ~new_n8732_;
  assign new_n8734_ = new_n1007_ & ~new_n8733_;
  assign new_n8735_ = new_n1011_ & ~new_n8734_;
  assign new_n8736_ = new_n1015_ & ~new_n8735_;
  assign new_n8737_ = new_n1019_ & ~new_n8736_;
  assign new_n8738_ = new_n1023_ & ~new_n8737_;
  assign new_n8739_ = new_n1027_ & ~new_n8738_;
  assign new_n8740_ = new_n1031_ & ~new_n8739_;
  assign new_n8741_ = new_n1035_ & ~new_n8740_;
  assign new_n8742_ = new_n1039_ & ~new_n8741_;
  assign new_n8743_ = new_n1043_ & ~new_n8742_;
  assign new_n8744_ = new_n1047_ & ~new_n8743_;
  assign new_n8745_ = new_n1051_ & ~new_n8744_;
  assign new_n8746_ = new_n1055_ & ~new_n8745_;
  assign new_n8747_ = new_n1059_ & ~new_n8746_;
  assign new_n8748_ = new_n1574_ & ~new_n8747_;
  assign new_n8749_ = new_n1576_ & ~new_n8748_;
  assign new_n8750_ = new_n1837_ & ~new_n8749_;
  assign new_n8751_ = new_n1068_ & ~new_n8750_;
  assign new_n8752_ = new_n1072_ & ~new_n8751_;
  assign new_n8753_ = new_n1076_ & ~new_n8752_;
  assign new_n8754_ = new_n1080_ & ~new_n8753_;
  assign new_n8755_ = new_n1084_ & ~new_n8754_;
  assign new_n8756_ = new_n1088_ & ~new_n8755_;
  assign new_n8757_ = new_n1092_ & ~new_n8756_;
  assign new_n8758_ = new_n1096_ & ~new_n8757_;
  assign new_n8759_ = new_n1100_ & ~new_n8758_;
  assign new_n8760_ = new_n1104_ & ~new_n8759_;
  assign new_n8761_ = new_n1108_ & ~new_n8760_;
  assign new_n8762_ = new_n1112_ & ~new_n8761_;
  assign new_n8763_ = new_n1116_ & ~new_n8762_;
  assign new_n8764_ = new_n1120_ & ~new_n8763_;
  assign new_n8765_ = new_n1124_ & ~new_n8764_;
  assign new_n8766_ = new_n1128_ & ~new_n8765_;
  assign new_n8767_ = new_n1132_ & ~new_n8766_;
  assign new_n8768_ = new_n1136_ & ~new_n8767_;
  assign new_n8769_ = new_n1140_ & ~new_n8768_;
  assign new_n8770_ = new_n1144_ & ~new_n8769_;
  assign new_n8771_ = new_n1148_ & ~new_n8770_;
  assign new_n8772_ = new_n1152_ & ~new_n8771_;
  assign new_n8773_ = new_n1156_ & ~new_n8772_;
  assign new_n8774_ = new_n1160_ & ~new_n8773_;
  assign new_n8775_ = new_n1164_ & ~new_n8774_;
  assign new_n8776_ = new_n1168_ & ~new_n8775_;
  assign new_n8777_ = new_n1172_ & ~new_n8776_;
  assign new_n8778_ = new_n1176_ & ~new_n8777_;
  assign new_n8779_ = new_n1180_ & ~new_n8778_;
  assign new_n8780_ = new_n1184_ & ~new_n8779_;
  assign new_n8781_ = new_n1188_ & ~new_n8780_;
  assign new_n8782_ = new_n1192_ & ~new_n8781_;
  assign new_n8783_ = new_n1196_ & ~new_n8782_;
  assign new_n8784_ = new_n1200_ & ~new_n8783_;
  assign new_n8785_ = new_n1204_ & ~new_n8784_;
  assign new_n8786_ = new_n1208_ & ~new_n8785_;
  assign new_n8787_ = new_n1212_ & ~new_n8786_;
  assign new_n8788_ = new_n1216_ & ~new_n8787_;
  assign new_n8789_ = new_n1220_ & ~new_n8788_;
  assign new_n8790_ = new_n1224_ & ~new_n8789_;
  assign new_n8791_ = new_n1228_ & ~new_n8790_;
  assign new_n8792_ = new_n1232_ & ~new_n8791_;
  assign new_n8793_ = new_n1236_ & ~new_n8792_;
  assign new_n8794_ = new_n1240_ & ~new_n8793_;
  assign new_n8795_ = new_n1244_ & ~new_n8794_;
  assign new_n8796_ = new_n1248_ & ~new_n8795_;
  assign new_n8797_ = new_n1252_ & ~new_n8796_;
  assign new_n8798_ = new_n1256_ & ~new_n8797_;
  assign new_n8799_ = new_n1260_ & ~new_n8798_;
  assign new_n8800_ = new_n1264_ & ~new_n8799_;
  assign new_n8801_ = new_n1268_ & ~new_n8800_;
  assign new_n8802_ = new_n1272_ & ~new_n8801_;
  assign new_n8803_ = new_n1276_ & ~new_n8802_;
  assign new_n8804_ = new_n1280_ & ~new_n8803_;
  assign new_n8805_ = new_n1284_ & ~new_n8804_;
  assign new_n8806_ = \req[88]  & ~new_n1286_;
  assign \grant[88]  = ~new_n8805_ & new_n8806_;
  assign new_n8808_ = ~new_n623_ & new_n1295_;
  assign new_n8809_ = new_n1300_ & ~new_n8808_;
  assign new_n8810_ = new_n1304_ & ~new_n8809_;
  assign new_n8811_ = new_n1308_ & ~new_n8810_;
  assign new_n8812_ = new_n1312_ & ~new_n8811_;
  assign new_n8813_ = new_n1316_ & ~new_n8812_;
  assign new_n8814_ = new_n1320_ & ~new_n8813_;
  assign new_n8815_ = new_n1324_ & ~new_n8814_;
  assign new_n8816_ = new_n1328_ & ~new_n8815_;
  assign new_n8817_ = new_n1332_ & ~new_n8816_;
  assign new_n8818_ = new_n1336_ & ~new_n8817_;
  assign new_n8819_ = new_n1340_ & ~new_n8818_;
  assign new_n8820_ = new_n1344_ & ~new_n8819_;
  assign new_n8821_ = new_n1348_ & ~new_n8820_;
  assign new_n8822_ = new_n1352_ & ~new_n8821_;
  assign new_n8823_ = new_n1356_ & ~new_n8822_;
  assign new_n8824_ = new_n1360_ & ~new_n8823_;
  assign new_n8825_ = new_n1364_ & ~new_n8824_;
  assign new_n8826_ = new_n1368_ & ~new_n8825_;
  assign new_n8827_ = new_n1372_ & ~new_n8826_;
  assign new_n8828_ = new_n1376_ & ~new_n8827_;
  assign new_n8829_ = new_n1380_ & ~new_n8828_;
  assign new_n8830_ = new_n1384_ & ~new_n8829_;
  assign new_n8831_ = new_n1388_ & ~new_n8830_;
  assign new_n8832_ = new_n1392_ & ~new_n8831_;
  assign new_n8833_ = new_n1396_ & ~new_n8832_;
  assign new_n8834_ = new_n1663_ & ~new_n8833_;
  assign new_n8835_ = new_n392_ & ~new_n8834_;
  assign new_n8836_ = new_n396_ & ~new_n8835_;
  assign new_n8837_ = new_n400_ & ~new_n8836_;
  assign new_n8838_ = new_n404_ & ~new_n8837_;
  assign new_n8839_ = new_n408_ & ~new_n8838_;
  assign new_n8840_ = new_n412_ & ~new_n8839_;
  assign new_n8841_ = new_n416_ & ~new_n8840_;
  assign new_n8842_ = new_n420_ & ~new_n8841_;
  assign new_n8843_ = new_n424_ & ~new_n8842_;
  assign new_n8844_ = new_n428_ & ~new_n8843_;
  assign new_n8845_ = new_n432_ & ~new_n8844_;
  assign new_n8846_ = new_n436_ & ~new_n8845_;
  assign new_n8847_ = new_n440_ & ~new_n8846_;
  assign new_n8848_ = new_n444_ & ~new_n8847_;
  assign new_n8849_ = new_n448_ & ~new_n8848_;
  assign new_n8850_ = new_n452_ & ~new_n8849_;
  assign new_n8851_ = new_n456_ & ~new_n8850_;
  assign new_n8852_ = new_n460_ & ~new_n8851_;
  assign new_n8853_ = new_n464_ & ~new_n8852_;
  assign new_n8854_ = new_n468_ & ~new_n8853_;
  assign new_n8855_ = new_n472_ & ~new_n8854_;
  assign new_n8856_ = new_n476_ & ~new_n8855_;
  assign new_n8857_ = new_n480_ & ~new_n8856_;
  assign new_n8858_ = new_n484_ & ~new_n8857_;
  assign new_n8859_ = new_n488_ & ~new_n8858_;
  assign new_n8860_ = new_n492_ & ~new_n8859_;
  assign new_n8861_ = new_n496_ & ~new_n8860_;
  assign new_n8862_ = new_n500_ & ~new_n8861_;
  assign new_n8863_ = new_n504_ & ~new_n8862_;
  assign new_n8864_ = new_n508_ & ~new_n8863_;
  assign new_n8865_ = new_n512_ & ~new_n8864_;
  assign new_n8866_ = new_n516_ & ~new_n8865_;
  assign new_n8867_ = new_n520_ & ~new_n8866_;
  assign new_n8868_ = new_n524_ & ~new_n8867_;
  assign new_n8869_ = new_n528_ & ~new_n8868_;
  assign new_n8870_ = new_n532_ & ~new_n8869_;
  assign new_n8871_ = new_n536_ & ~new_n8870_;
  assign new_n8872_ = new_n540_ & ~new_n8871_;
  assign new_n8873_ = new_n544_ & ~new_n8872_;
  assign new_n8874_ = new_n548_ & ~new_n8873_;
  assign new_n8875_ = new_n552_ & ~new_n8874_;
  assign new_n8876_ = new_n556_ & ~new_n8875_;
  assign new_n8877_ = new_n560_ & ~new_n8876_;
  assign new_n8878_ = new_n564_ & ~new_n8877_;
  assign new_n8879_ = new_n568_ & ~new_n8878_;
  assign new_n8880_ = new_n572_ & ~new_n8879_;
  assign new_n8881_ = new_n576_ & ~new_n8880_;
  assign new_n8882_ = new_n580_ & ~new_n8881_;
  assign new_n8883_ = new_n584_ & ~new_n8882_;
  assign new_n8884_ = new_n588_ & ~new_n8883_;
  assign new_n8885_ = new_n592_ & ~new_n8884_;
  assign new_n8886_ = new_n596_ & ~new_n8885_;
  assign new_n8887_ = new_n600_ & ~new_n8886_;
  assign new_n8888_ = new_n604_ & ~new_n8887_;
  assign new_n8889_ = new_n608_ & ~new_n8888_;
  assign new_n8890_ = new_n612_ & ~new_n8889_;
  assign new_n8891_ = new_n616_ & ~new_n8890_;
  assign new_n8892_ = \req[89]  & ~new_n618_;
  assign \grant[89]  = ~new_n8891_ & new_n8892_;
  assign new_n8894_ = new_n627_ & ~new_n962_;
  assign new_n8895_ = new_n632_ & ~new_n8894_;
  assign new_n8896_ = new_n636_ & ~new_n8895_;
  assign new_n8897_ = new_n640_ & ~new_n8896_;
  assign new_n8898_ = new_n644_ & ~new_n8897_;
  assign new_n8899_ = new_n648_ & ~new_n8898_;
  assign new_n8900_ = new_n652_ & ~new_n8899_;
  assign new_n8901_ = new_n656_ & ~new_n8900_;
  assign new_n8902_ = new_n660_ & ~new_n8901_;
  assign new_n8903_ = new_n664_ & ~new_n8902_;
  assign new_n8904_ = new_n668_ & ~new_n8903_;
  assign new_n8905_ = new_n672_ & ~new_n8904_;
  assign new_n8906_ = new_n676_ & ~new_n8905_;
  assign new_n8907_ = new_n680_ & ~new_n8906_;
  assign new_n8908_ = new_n684_ & ~new_n8907_;
  assign new_n8909_ = new_n688_ & ~new_n8908_;
  assign new_n8910_ = new_n692_ & ~new_n8909_;
  assign new_n8911_ = new_n696_ & ~new_n8910_;
  assign new_n8912_ = new_n700_ & ~new_n8911_;
  assign new_n8913_ = new_n704_ & ~new_n8912_;
  assign new_n8914_ = new_n708_ & ~new_n8913_;
  assign new_n8915_ = new_n712_ & ~new_n8914_;
  assign new_n8916_ = new_n716_ & ~new_n8915_;
  assign new_n8917_ = new_n720_ & ~new_n8916_;
  assign new_n8918_ = new_n1484_ & ~new_n8917_;
  assign new_n8919_ = new_n1486_ & ~new_n8918_;
  assign new_n8920_ = new_n1750_ & ~new_n8919_;
  assign new_n8921_ = new_n731_ & ~new_n8920_;
  assign new_n8922_ = new_n735_ & ~new_n8921_;
  assign new_n8923_ = new_n739_ & ~new_n8922_;
  assign new_n8924_ = new_n743_ & ~new_n8923_;
  assign new_n8925_ = new_n747_ & ~new_n8924_;
  assign new_n8926_ = new_n751_ & ~new_n8925_;
  assign new_n8927_ = new_n755_ & ~new_n8926_;
  assign new_n8928_ = new_n759_ & ~new_n8927_;
  assign new_n8929_ = new_n763_ & ~new_n8928_;
  assign new_n8930_ = new_n767_ & ~new_n8929_;
  assign new_n8931_ = new_n771_ & ~new_n8930_;
  assign new_n8932_ = new_n775_ & ~new_n8931_;
  assign new_n8933_ = new_n779_ & ~new_n8932_;
  assign new_n8934_ = new_n783_ & ~new_n8933_;
  assign new_n8935_ = new_n787_ & ~new_n8934_;
  assign new_n8936_ = new_n791_ & ~new_n8935_;
  assign new_n8937_ = new_n795_ & ~new_n8936_;
  assign new_n8938_ = new_n799_ & ~new_n8937_;
  assign new_n8939_ = new_n803_ & ~new_n8938_;
  assign new_n8940_ = new_n807_ & ~new_n8939_;
  assign new_n8941_ = new_n811_ & ~new_n8940_;
  assign new_n8942_ = new_n815_ & ~new_n8941_;
  assign new_n8943_ = new_n819_ & ~new_n8942_;
  assign new_n8944_ = new_n823_ & ~new_n8943_;
  assign new_n8945_ = new_n827_ & ~new_n8944_;
  assign new_n8946_ = new_n831_ & ~new_n8945_;
  assign new_n8947_ = new_n835_ & ~new_n8946_;
  assign new_n8948_ = new_n839_ & ~new_n8947_;
  assign new_n8949_ = new_n843_ & ~new_n8948_;
  assign new_n8950_ = new_n847_ & ~new_n8949_;
  assign new_n8951_ = new_n851_ & ~new_n8950_;
  assign new_n8952_ = new_n855_ & ~new_n8951_;
  assign new_n8953_ = new_n859_ & ~new_n8952_;
  assign new_n8954_ = new_n863_ & ~new_n8953_;
  assign new_n8955_ = new_n867_ & ~new_n8954_;
  assign new_n8956_ = new_n871_ & ~new_n8955_;
  assign new_n8957_ = new_n875_ & ~new_n8956_;
  assign new_n8958_ = new_n879_ & ~new_n8957_;
  assign new_n8959_ = new_n883_ & ~new_n8958_;
  assign new_n8960_ = new_n887_ & ~new_n8959_;
  assign new_n8961_ = new_n891_ & ~new_n8960_;
  assign new_n8962_ = new_n895_ & ~new_n8961_;
  assign new_n8963_ = new_n899_ & ~new_n8962_;
  assign new_n8964_ = new_n903_ & ~new_n8963_;
  assign new_n8965_ = new_n907_ & ~new_n8964_;
  assign new_n8966_ = new_n911_ & ~new_n8965_;
  assign new_n8967_ = new_n915_ & ~new_n8966_;
  assign new_n8968_ = new_n919_ & ~new_n8967_;
  assign new_n8969_ = new_n923_ & ~new_n8968_;
  assign new_n8970_ = new_n927_ & ~new_n8969_;
  assign new_n8971_ = new_n931_ & ~new_n8970_;
  assign new_n8972_ = new_n935_ & ~new_n8971_;
  assign new_n8973_ = new_n939_ & ~new_n8972_;
  assign new_n8974_ = new_n943_ & ~new_n8973_;
  assign new_n8975_ = new_n947_ & ~new_n8974_;
  assign new_n8976_ = new_n951_ & ~new_n8975_;
  assign new_n8977_ = new_n955_ & ~new_n8976_;
  assign new_n8978_ = \req[90]  & ~new_n957_;
  assign \grant[90]  = ~new_n8977_ & new_n8978_;
  assign new_n8980_ = new_n966_ & ~new_n1299_;
  assign new_n8981_ = new_n971_ & ~new_n8980_;
  assign new_n8982_ = new_n975_ & ~new_n8981_;
  assign new_n8983_ = new_n979_ & ~new_n8982_;
  assign new_n8984_ = new_n983_ & ~new_n8983_;
  assign new_n8985_ = new_n987_ & ~new_n8984_;
  assign new_n8986_ = new_n991_ & ~new_n8985_;
  assign new_n8987_ = new_n995_ & ~new_n8986_;
  assign new_n8988_ = new_n999_ & ~new_n8987_;
  assign new_n8989_ = new_n1003_ & ~new_n8988_;
  assign new_n8990_ = new_n1007_ & ~new_n8989_;
  assign new_n8991_ = new_n1011_ & ~new_n8990_;
  assign new_n8992_ = new_n1015_ & ~new_n8991_;
  assign new_n8993_ = new_n1019_ & ~new_n8992_;
  assign new_n8994_ = new_n1023_ & ~new_n8993_;
  assign new_n8995_ = new_n1027_ & ~new_n8994_;
  assign new_n8996_ = new_n1031_ & ~new_n8995_;
  assign new_n8997_ = new_n1035_ & ~new_n8996_;
  assign new_n8998_ = new_n1039_ & ~new_n8997_;
  assign new_n8999_ = new_n1043_ & ~new_n8998_;
  assign new_n9000_ = new_n1047_ & ~new_n8999_;
  assign new_n9001_ = new_n1051_ & ~new_n9000_;
  assign new_n9002_ = new_n1055_ & ~new_n9001_;
  assign new_n9003_ = new_n1059_ & ~new_n9002_;
  assign new_n9004_ = new_n1574_ & ~new_n9003_;
  assign new_n9005_ = new_n1576_ & ~new_n9004_;
  assign new_n9006_ = new_n1837_ & ~new_n9005_;
  assign new_n9007_ = new_n1068_ & ~new_n9006_;
  assign new_n9008_ = new_n1072_ & ~new_n9007_;
  assign new_n9009_ = new_n1076_ & ~new_n9008_;
  assign new_n9010_ = new_n1080_ & ~new_n9009_;
  assign new_n9011_ = new_n1084_ & ~new_n9010_;
  assign new_n9012_ = new_n1088_ & ~new_n9011_;
  assign new_n9013_ = new_n1092_ & ~new_n9012_;
  assign new_n9014_ = new_n1096_ & ~new_n9013_;
  assign new_n9015_ = new_n1100_ & ~new_n9014_;
  assign new_n9016_ = new_n1104_ & ~new_n9015_;
  assign new_n9017_ = new_n1108_ & ~new_n9016_;
  assign new_n9018_ = new_n1112_ & ~new_n9017_;
  assign new_n9019_ = new_n1116_ & ~new_n9018_;
  assign new_n9020_ = new_n1120_ & ~new_n9019_;
  assign new_n9021_ = new_n1124_ & ~new_n9020_;
  assign new_n9022_ = new_n1128_ & ~new_n9021_;
  assign new_n9023_ = new_n1132_ & ~new_n9022_;
  assign new_n9024_ = new_n1136_ & ~new_n9023_;
  assign new_n9025_ = new_n1140_ & ~new_n9024_;
  assign new_n9026_ = new_n1144_ & ~new_n9025_;
  assign new_n9027_ = new_n1148_ & ~new_n9026_;
  assign new_n9028_ = new_n1152_ & ~new_n9027_;
  assign new_n9029_ = new_n1156_ & ~new_n9028_;
  assign new_n9030_ = new_n1160_ & ~new_n9029_;
  assign new_n9031_ = new_n1164_ & ~new_n9030_;
  assign new_n9032_ = new_n1168_ & ~new_n9031_;
  assign new_n9033_ = new_n1172_ & ~new_n9032_;
  assign new_n9034_ = new_n1176_ & ~new_n9033_;
  assign new_n9035_ = new_n1180_ & ~new_n9034_;
  assign new_n9036_ = new_n1184_ & ~new_n9035_;
  assign new_n9037_ = new_n1188_ & ~new_n9036_;
  assign new_n9038_ = new_n1192_ & ~new_n9037_;
  assign new_n9039_ = new_n1196_ & ~new_n9038_;
  assign new_n9040_ = new_n1200_ & ~new_n9039_;
  assign new_n9041_ = new_n1204_ & ~new_n9040_;
  assign new_n9042_ = new_n1208_ & ~new_n9041_;
  assign new_n9043_ = new_n1212_ & ~new_n9042_;
  assign new_n9044_ = new_n1216_ & ~new_n9043_;
  assign new_n9045_ = new_n1220_ & ~new_n9044_;
  assign new_n9046_ = new_n1224_ & ~new_n9045_;
  assign new_n9047_ = new_n1228_ & ~new_n9046_;
  assign new_n9048_ = new_n1232_ & ~new_n9047_;
  assign new_n9049_ = new_n1236_ & ~new_n9048_;
  assign new_n9050_ = new_n1240_ & ~new_n9049_;
  assign new_n9051_ = new_n1244_ & ~new_n9050_;
  assign new_n9052_ = new_n1248_ & ~new_n9051_;
  assign new_n9053_ = new_n1252_ & ~new_n9052_;
  assign new_n9054_ = new_n1256_ & ~new_n9053_;
  assign new_n9055_ = new_n1260_ & ~new_n9054_;
  assign new_n9056_ = new_n1264_ & ~new_n9055_;
  assign new_n9057_ = new_n1268_ & ~new_n9056_;
  assign new_n9058_ = new_n1272_ & ~new_n9057_;
  assign new_n9059_ = new_n1276_ & ~new_n9058_;
  assign new_n9060_ = new_n1280_ & ~new_n9059_;
  assign new_n9061_ = new_n1284_ & ~new_n9060_;
  assign new_n9062_ = new_n1288_ & ~new_n9061_;
  assign new_n9063_ = new_n1292_ & ~new_n9062_;
  assign new_n9064_ = \req[91]  & ~new_n1294_;
  assign \grant[91]  = ~new_n9063_ & new_n9064_;
  assign new_n9066_ = ~new_n631_ & new_n1303_;
  assign new_n9067_ = new_n1308_ & ~new_n9066_;
  assign new_n9068_ = new_n1312_ & ~new_n9067_;
  assign new_n9069_ = new_n1316_ & ~new_n9068_;
  assign new_n9070_ = new_n1320_ & ~new_n9069_;
  assign new_n9071_ = new_n1324_ & ~new_n9070_;
  assign new_n9072_ = new_n1328_ & ~new_n9071_;
  assign new_n9073_ = new_n1332_ & ~new_n9072_;
  assign new_n9074_ = new_n1336_ & ~new_n9073_;
  assign new_n9075_ = new_n1340_ & ~new_n9074_;
  assign new_n9076_ = new_n1344_ & ~new_n9075_;
  assign new_n9077_ = new_n1348_ & ~new_n9076_;
  assign new_n9078_ = new_n1352_ & ~new_n9077_;
  assign new_n9079_ = new_n1356_ & ~new_n9078_;
  assign new_n9080_ = new_n1360_ & ~new_n9079_;
  assign new_n9081_ = new_n1364_ & ~new_n9080_;
  assign new_n9082_ = new_n1368_ & ~new_n9081_;
  assign new_n9083_ = new_n1372_ & ~new_n9082_;
  assign new_n9084_ = new_n1376_ & ~new_n9083_;
  assign new_n9085_ = new_n1380_ & ~new_n9084_;
  assign new_n9086_ = new_n1384_ & ~new_n9085_;
  assign new_n9087_ = new_n1388_ & ~new_n9086_;
  assign new_n9088_ = new_n1392_ & ~new_n9087_;
  assign new_n9089_ = new_n1396_ & ~new_n9088_;
  assign new_n9090_ = new_n1663_ & ~new_n9089_;
  assign new_n9091_ = new_n392_ & ~new_n9090_;
  assign new_n9092_ = new_n396_ & ~new_n9091_;
  assign new_n9093_ = new_n400_ & ~new_n9092_;
  assign new_n9094_ = new_n404_ & ~new_n9093_;
  assign new_n9095_ = new_n408_ & ~new_n9094_;
  assign new_n9096_ = new_n412_ & ~new_n9095_;
  assign new_n9097_ = new_n416_ & ~new_n9096_;
  assign new_n9098_ = new_n420_ & ~new_n9097_;
  assign new_n9099_ = new_n424_ & ~new_n9098_;
  assign new_n9100_ = new_n428_ & ~new_n9099_;
  assign new_n9101_ = new_n432_ & ~new_n9100_;
  assign new_n9102_ = new_n436_ & ~new_n9101_;
  assign new_n9103_ = new_n440_ & ~new_n9102_;
  assign new_n9104_ = new_n444_ & ~new_n9103_;
  assign new_n9105_ = new_n448_ & ~new_n9104_;
  assign new_n9106_ = new_n452_ & ~new_n9105_;
  assign new_n9107_ = new_n456_ & ~new_n9106_;
  assign new_n9108_ = new_n460_ & ~new_n9107_;
  assign new_n9109_ = new_n464_ & ~new_n9108_;
  assign new_n9110_ = new_n468_ & ~new_n9109_;
  assign new_n9111_ = new_n472_ & ~new_n9110_;
  assign new_n9112_ = new_n476_ & ~new_n9111_;
  assign new_n9113_ = new_n480_ & ~new_n9112_;
  assign new_n9114_ = new_n484_ & ~new_n9113_;
  assign new_n9115_ = new_n488_ & ~new_n9114_;
  assign new_n9116_ = new_n492_ & ~new_n9115_;
  assign new_n9117_ = new_n496_ & ~new_n9116_;
  assign new_n9118_ = new_n500_ & ~new_n9117_;
  assign new_n9119_ = new_n504_ & ~new_n9118_;
  assign new_n9120_ = new_n508_ & ~new_n9119_;
  assign new_n9121_ = new_n512_ & ~new_n9120_;
  assign new_n9122_ = new_n516_ & ~new_n9121_;
  assign new_n9123_ = new_n520_ & ~new_n9122_;
  assign new_n9124_ = new_n524_ & ~new_n9123_;
  assign new_n9125_ = new_n528_ & ~new_n9124_;
  assign new_n9126_ = new_n532_ & ~new_n9125_;
  assign new_n9127_ = new_n536_ & ~new_n9126_;
  assign new_n9128_ = new_n540_ & ~new_n9127_;
  assign new_n9129_ = new_n544_ & ~new_n9128_;
  assign new_n9130_ = new_n548_ & ~new_n9129_;
  assign new_n9131_ = new_n552_ & ~new_n9130_;
  assign new_n9132_ = new_n556_ & ~new_n9131_;
  assign new_n9133_ = new_n560_ & ~new_n9132_;
  assign new_n9134_ = new_n564_ & ~new_n9133_;
  assign new_n9135_ = new_n568_ & ~new_n9134_;
  assign new_n9136_ = new_n572_ & ~new_n9135_;
  assign new_n9137_ = new_n576_ & ~new_n9136_;
  assign new_n9138_ = new_n580_ & ~new_n9137_;
  assign new_n9139_ = new_n584_ & ~new_n9138_;
  assign new_n9140_ = new_n588_ & ~new_n9139_;
  assign new_n9141_ = new_n592_ & ~new_n9140_;
  assign new_n9142_ = new_n596_ & ~new_n9141_;
  assign new_n9143_ = new_n600_ & ~new_n9142_;
  assign new_n9144_ = new_n604_ & ~new_n9143_;
  assign new_n9145_ = new_n608_ & ~new_n9144_;
  assign new_n9146_ = new_n612_ & ~new_n9145_;
  assign new_n9147_ = new_n616_ & ~new_n9146_;
  assign new_n9148_ = new_n620_ & ~new_n9147_;
  assign new_n9149_ = new_n624_ & ~new_n9148_;
  assign new_n9150_ = \req[92]  & ~new_n626_;
  assign \grant[92]  = ~new_n9149_ & new_n9150_;
  assign new_n9152_ = new_n635_ & ~new_n970_;
  assign new_n9153_ = new_n640_ & ~new_n9152_;
  assign new_n9154_ = new_n644_ & ~new_n9153_;
  assign new_n9155_ = new_n648_ & ~new_n9154_;
  assign new_n9156_ = new_n652_ & ~new_n9155_;
  assign new_n9157_ = new_n656_ & ~new_n9156_;
  assign new_n9158_ = new_n660_ & ~new_n9157_;
  assign new_n9159_ = new_n664_ & ~new_n9158_;
  assign new_n9160_ = new_n668_ & ~new_n9159_;
  assign new_n9161_ = new_n672_ & ~new_n9160_;
  assign new_n9162_ = new_n676_ & ~new_n9161_;
  assign new_n9163_ = new_n680_ & ~new_n9162_;
  assign new_n9164_ = new_n684_ & ~new_n9163_;
  assign new_n9165_ = new_n688_ & ~new_n9164_;
  assign new_n9166_ = new_n692_ & ~new_n9165_;
  assign new_n9167_ = new_n696_ & ~new_n9166_;
  assign new_n9168_ = new_n700_ & ~new_n9167_;
  assign new_n9169_ = new_n704_ & ~new_n9168_;
  assign new_n9170_ = new_n708_ & ~new_n9169_;
  assign new_n9171_ = new_n712_ & ~new_n9170_;
  assign new_n9172_ = new_n716_ & ~new_n9171_;
  assign new_n9173_ = new_n720_ & ~new_n9172_;
  assign new_n9174_ = new_n1484_ & ~new_n9173_;
  assign new_n9175_ = new_n1486_ & ~new_n9174_;
  assign new_n9176_ = new_n1750_ & ~new_n9175_;
  assign new_n9177_ = new_n731_ & ~new_n9176_;
  assign new_n9178_ = new_n735_ & ~new_n9177_;
  assign new_n9179_ = new_n739_ & ~new_n9178_;
  assign new_n9180_ = new_n743_ & ~new_n9179_;
  assign new_n9181_ = new_n747_ & ~new_n9180_;
  assign new_n9182_ = new_n751_ & ~new_n9181_;
  assign new_n9183_ = new_n755_ & ~new_n9182_;
  assign new_n9184_ = new_n759_ & ~new_n9183_;
  assign new_n9185_ = new_n763_ & ~new_n9184_;
  assign new_n9186_ = new_n767_ & ~new_n9185_;
  assign new_n9187_ = new_n771_ & ~new_n9186_;
  assign new_n9188_ = new_n775_ & ~new_n9187_;
  assign new_n9189_ = new_n779_ & ~new_n9188_;
  assign new_n9190_ = new_n783_ & ~new_n9189_;
  assign new_n9191_ = new_n787_ & ~new_n9190_;
  assign new_n9192_ = new_n791_ & ~new_n9191_;
  assign new_n9193_ = new_n795_ & ~new_n9192_;
  assign new_n9194_ = new_n799_ & ~new_n9193_;
  assign new_n9195_ = new_n803_ & ~new_n9194_;
  assign new_n9196_ = new_n807_ & ~new_n9195_;
  assign new_n9197_ = new_n811_ & ~new_n9196_;
  assign new_n9198_ = new_n815_ & ~new_n9197_;
  assign new_n9199_ = new_n819_ & ~new_n9198_;
  assign new_n9200_ = new_n823_ & ~new_n9199_;
  assign new_n9201_ = new_n827_ & ~new_n9200_;
  assign new_n9202_ = new_n831_ & ~new_n9201_;
  assign new_n9203_ = new_n835_ & ~new_n9202_;
  assign new_n9204_ = new_n839_ & ~new_n9203_;
  assign new_n9205_ = new_n843_ & ~new_n9204_;
  assign new_n9206_ = new_n847_ & ~new_n9205_;
  assign new_n9207_ = new_n851_ & ~new_n9206_;
  assign new_n9208_ = new_n855_ & ~new_n9207_;
  assign new_n9209_ = new_n859_ & ~new_n9208_;
  assign new_n9210_ = new_n863_ & ~new_n9209_;
  assign new_n9211_ = new_n867_ & ~new_n9210_;
  assign new_n9212_ = new_n871_ & ~new_n9211_;
  assign new_n9213_ = new_n875_ & ~new_n9212_;
  assign new_n9214_ = new_n879_ & ~new_n9213_;
  assign new_n9215_ = new_n883_ & ~new_n9214_;
  assign new_n9216_ = new_n887_ & ~new_n9215_;
  assign new_n9217_ = new_n891_ & ~new_n9216_;
  assign new_n9218_ = new_n895_ & ~new_n9217_;
  assign new_n9219_ = new_n899_ & ~new_n9218_;
  assign new_n9220_ = new_n903_ & ~new_n9219_;
  assign new_n9221_ = new_n907_ & ~new_n9220_;
  assign new_n9222_ = new_n911_ & ~new_n9221_;
  assign new_n9223_ = new_n915_ & ~new_n9222_;
  assign new_n9224_ = new_n919_ & ~new_n9223_;
  assign new_n9225_ = new_n923_ & ~new_n9224_;
  assign new_n9226_ = new_n927_ & ~new_n9225_;
  assign new_n9227_ = new_n931_ & ~new_n9226_;
  assign new_n9228_ = new_n935_ & ~new_n9227_;
  assign new_n9229_ = new_n939_ & ~new_n9228_;
  assign new_n9230_ = new_n943_ & ~new_n9229_;
  assign new_n9231_ = new_n947_ & ~new_n9230_;
  assign new_n9232_ = new_n951_ & ~new_n9231_;
  assign new_n9233_ = new_n955_ & ~new_n9232_;
  assign new_n9234_ = new_n959_ & ~new_n9233_;
  assign new_n9235_ = new_n963_ & ~new_n9234_;
  assign new_n9236_ = \req[93]  & ~new_n965_;
  assign \grant[93]  = ~new_n9235_ & new_n9236_;
  assign new_n9238_ = new_n974_ & ~new_n1307_;
  assign new_n9239_ = new_n979_ & ~new_n9238_;
  assign new_n9240_ = new_n983_ & ~new_n9239_;
  assign new_n9241_ = new_n987_ & ~new_n9240_;
  assign new_n9242_ = new_n991_ & ~new_n9241_;
  assign new_n9243_ = new_n995_ & ~new_n9242_;
  assign new_n9244_ = new_n999_ & ~new_n9243_;
  assign new_n9245_ = new_n1003_ & ~new_n9244_;
  assign new_n9246_ = new_n1007_ & ~new_n9245_;
  assign new_n9247_ = new_n1011_ & ~new_n9246_;
  assign new_n9248_ = new_n1015_ & ~new_n9247_;
  assign new_n9249_ = new_n1019_ & ~new_n9248_;
  assign new_n9250_ = new_n1023_ & ~new_n9249_;
  assign new_n9251_ = new_n1027_ & ~new_n9250_;
  assign new_n9252_ = new_n1031_ & ~new_n9251_;
  assign new_n9253_ = new_n1035_ & ~new_n9252_;
  assign new_n9254_ = new_n1039_ & ~new_n9253_;
  assign new_n9255_ = new_n1043_ & ~new_n9254_;
  assign new_n9256_ = new_n1047_ & ~new_n9255_;
  assign new_n9257_ = new_n1051_ & ~new_n9256_;
  assign new_n9258_ = new_n1055_ & ~new_n9257_;
  assign new_n9259_ = new_n1059_ & ~new_n9258_;
  assign new_n9260_ = new_n1574_ & ~new_n9259_;
  assign new_n9261_ = new_n1576_ & ~new_n9260_;
  assign new_n9262_ = new_n1837_ & ~new_n9261_;
  assign new_n9263_ = new_n1068_ & ~new_n9262_;
  assign new_n9264_ = new_n1072_ & ~new_n9263_;
  assign new_n9265_ = new_n1076_ & ~new_n9264_;
  assign new_n9266_ = new_n1080_ & ~new_n9265_;
  assign new_n9267_ = new_n1084_ & ~new_n9266_;
  assign new_n9268_ = new_n1088_ & ~new_n9267_;
  assign new_n9269_ = new_n1092_ & ~new_n9268_;
  assign new_n9270_ = new_n1096_ & ~new_n9269_;
  assign new_n9271_ = new_n1100_ & ~new_n9270_;
  assign new_n9272_ = new_n1104_ & ~new_n9271_;
  assign new_n9273_ = new_n1108_ & ~new_n9272_;
  assign new_n9274_ = new_n1112_ & ~new_n9273_;
  assign new_n9275_ = new_n1116_ & ~new_n9274_;
  assign new_n9276_ = new_n1120_ & ~new_n9275_;
  assign new_n9277_ = new_n1124_ & ~new_n9276_;
  assign new_n9278_ = new_n1128_ & ~new_n9277_;
  assign new_n9279_ = new_n1132_ & ~new_n9278_;
  assign new_n9280_ = new_n1136_ & ~new_n9279_;
  assign new_n9281_ = new_n1140_ & ~new_n9280_;
  assign new_n9282_ = new_n1144_ & ~new_n9281_;
  assign new_n9283_ = new_n1148_ & ~new_n9282_;
  assign new_n9284_ = new_n1152_ & ~new_n9283_;
  assign new_n9285_ = new_n1156_ & ~new_n9284_;
  assign new_n9286_ = new_n1160_ & ~new_n9285_;
  assign new_n9287_ = new_n1164_ & ~new_n9286_;
  assign new_n9288_ = new_n1168_ & ~new_n9287_;
  assign new_n9289_ = new_n1172_ & ~new_n9288_;
  assign new_n9290_ = new_n1176_ & ~new_n9289_;
  assign new_n9291_ = new_n1180_ & ~new_n9290_;
  assign new_n9292_ = new_n1184_ & ~new_n9291_;
  assign new_n9293_ = new_n1188_ & ~new_n9292_;
  assign new_n9294_ = new_n1192_ & ~new_n9293_;
  assign new_n9295_ = new_n1196_ & ~new_n9294_;
  assign new_n9296_ = new_n1200_ & ~new_n9295_;
  assign new_n9297_ = new_n1204_ & ~new_n9296_;
  assign new_n9298_ = new_n1208_ & ~new_n9297_;
  assign new_n9299_ = new_n1212_ & ~new_n9298_;
  assign new_n9300_ = new_n1216_ & ~new_n9299_;
  assign new_n9301_ = new_n1220_ & ~new_n9300_;
  assign new_n9302_ = new_n1224_ & ~new_n9301_;
  assign new_n9303_ = new_n1228_ & ~new_n9302_;
  assign new_n9304_ = new_n1232_ & ~new_n9303_;
  assign new_n9305_ = new_n1236_ & ~new_n9304_;
  assign new_n9306_ = new_n1240_ & ~new_n9305_;
  assign new_n9307_ = new_n1244_ & ~new_n9306_;
  assign new_n9308_ = new_n1248_ & ~new_n9307_;
  assign new_n9309_ = new_n1252_ & ~new_n9308_;
  assign new_n9310_ = new_n1256_ & ~new_n9309_;
  assign new_n9311_ = new_n1260_ & ~new_n9310_;
  assign new_n9312_ = new_n1264_ & ~new_n9311_;
  assign new_n9313_ = new_n1268_ & ~new_n9312_;
  assign new_n9314_ = new_n1272_ & ~new_n9313_;
  assign new_n9315_ = new_n1276_ & ~new_n9314_;
  assign new_n9316_ = new_n1280_ & ~new_n9315_;
  assign new_n9317_ = new_n1284_ & ~new_n9316_;
  assign new_n9318_ = new_n1288_ & ~new_n9317_;
  assign new_n9319_ = new_n1292_ & ~new_n9318_;
  assign new_n9320_ = new_n1296_ & ~new_n9319_;
  assign new_n9321_ = new_n1300_ & ~new_n9320_;
  assign new_n9322_ = \req[94]  & ~new_n1302_;
  assign \grant[94]  = ~new_n9321_ & new_n9322_;
  assign new_n9324_ = ~new_n639_ & new_n1311_;
  assign new_n9325_ = new_n1316_ & ~new_n9324_;
  assign new_n9326_ = new_n1320_ & ~new_n9325_;
  assign new_n9327_ = new_n1324_ & ~new_n9326_;
  assign new_n9328_ = new_n1328_ & ~new_n9327_;
  assign new_n9329_ = new_n1332_ & ~new_n9328_;
  assign new_n9330_ = new_n1336_ & ~new_n9329_;
  assign new_n9331_ = new_n1340_ & ~new_n9330_;
  assign new_n9332_ = new_n1344_ & ~new_n9331_;
  assign new_n9333_ = new_n1348_ & ~new_n9332_;
  assign new_n9334_ = new_n1352_ & ~new_n9333_;
  assign new_n9335_ = new_n1356_ & ~new_n9334_;
  assign new_n9336_ = new_n1360_ & ~new_n9335_;
  assign new_n9337_ = new_n1364_ & ~new_n9336_;
  assign new_n9338_ = new_n1368_ & ~new_n9337_;
  assign new_n9339_ = new_n1372_ & ~new_n9338_;
  assign new_n9340_ = new_n1376_ & ~new_n9339_;
  assign new_n9341_ = new_n1380_ & ~new_n9340_;
  assign new_n9342_ = new_n1384_ & ~new_n9341_;
  assign new_n9343_ = new_n1388_ & ~new_n9342_;
  assign new_n9344_ = new_n1392_ & ~new_n9343_;
  assign new_n9345_ = new_n1396_ & ~new_n9344_;
  assign new_n9346_ = new_n1663_ & ~new_n9345_;
  assign new_n9347_ = new_n392_ & ~new_n9346_;
  assign new_n9348_ = new_n396_ & ~new_n9347_;
  assign new_n9349_ = new_n400_ & ~new_n9348_;
  assign new_n9350_ = new_n404_ & ~new_n9349_;
  assign new_n9351_ = new_n408_ & ~new_n9350_;
  assign new_n9352_ = new_n412_ & ~new_n9351_;
  assign new_n9353_ = new_n416_ & ~new_n9352_;
  assign new_n9354_ = new_n420_ & ~new_n9353_;
  assign new_n9355_ = new_n424_ & ~new_n9354_;
  assign new_n9356_ = new_n428_ & ~new_n9355_;
  assign new_n9357_ = new_n432_ & ~new_n9356_;
  assign new_n9358_ = new_n436_ & ~new_n9357_;
  assign new_n9359_ = new_n440_ & ~new_n9358_;
  assign new_n9360_ = new_n444_ & ~new_n9359_;
  assign new_n9361_ = new_n448_ & ~new_n9360_;
  assign new_n9362_ = new_n452_ & ~new_n9361_;
  assign new_n9363_ = new_n456_ & ~new_n9362_;
  assign new_n9364_ = new_n460_ & ~new_n9363_;
  assign new_n9365_ = new_n464_ & ~new_n9364_;
  assign new_n9366_ = new_n468_ & ~new_n9365_;
  assign new_n9367_ = new_n472_ & ~new_n9366_;
  assign new_n9368_ = new_n476_ & ~new_n9367_;
  assign new_n9369_ = new_n480_ & ~new_n9368_;
  assign new_n9370_ = new_n484_ & ~new_n9369_;
  assign new_n9371_ = new_n488_ & ~new_n9370_;
  assign new_n9372_ = new_n492_ & ~new_n9371_;
  assign new_n9373_ = new_n496_ & ~new_n9372_;
  assign new_n9374_ = new_n500_ & ~new_n9373_;
  assign new_n9375_ = new_n504_ & ~new_n9374_;
  assign new_n9376_ = new_n508_ & ~new_n9375_;
  assign new_n9377_ = new_n512_ & ~new_n9376_;
  assign new_n9378_ = new_n516_ & ~new_n9377_;
  assign new_n9379_ = new_n520_ & ~new_n9378_;
  assign new_n9380_ = new_n524_ & ~new_n9379_;
  assign new_n9381_ = new_n528_ & ~new_n9380_;
  assign new_n9382_ = new_n532_ & ~new_n9381_;
  assign new_n9383_ = new_n536_ & ~new_n9382_;
  assign new_n9384_ = new_n540_ & ~new_n9383_;
  assign new_n9385_ = new_n544_ & ~new_n9384_;
  assign new_n9386_ = new_n548_ & ~new_n9385_;
  assign new_n9387_ = new_n552_ & ~new_n9386_;
  assign new_n9388_ = new_n556_ & ~new_n9387_;
  assign new_n9389_ = new_n560_ & ~new_n9388_;
  assign new_n9390_ = new_n564_ & ~new_n9389_;
  assign new_n9391_ = new_n568_ & ~new_n9390_;
  assign new_n9392_ = new_n572_ & ~new_n9391_;
  assign new_n9393_ = new_n576_ & ~new_n9392_;
  assign new_n9394_ = new_n580_ & ~new_n9393_;
  assign new_n9395_ = new_n584_ & ~new_n9394_;
  assign new_n9396_ = new_n588_ & ~new_n9395_;
  assign new_n9397_ = new_n592_ & ~new_n9396_;
  assign new_n9398_ = new_n596_ & ~new_n9397_;
  assign new_n9399_ = new_n600_ & ~new_n9398_;
  assign new_n9400_ = new_n604_ & ~new_n9399_;
  assign new_n9401_ = new_n608_ & ~new_n9400_;
  assign new_n9402_ = new_n612_ & ~new_n9401_;
  assign new_n9403_ = new_n616_ & ~new_n9402_;
  assign new_n9404_ = new_n620_ & ~new_n9403_;
  assign new_n9405_ = new_n624_ & ~new_n9404_;
  assign new_n9406_ = new_n628_ & ~new_n9405_;
  assign new_n9407_ = new_n632_ & ~new_n9406_;
  assign new_n9408_ = \req[95]  & ~new_n634_;
  assign \grant[95]  = ~new_n9407_ & new_n9408_;
  assign new_n9410_ = new_n643_ & ~new_n978_;
  assign new_n9411_ = new_n648_ & ~new_n9410_;
  assign new_n9412_ = new_n652_ & ~new_n9411_;
  assign new_n9413_ = new_n656_ & ~new_n9412_;
  assign new_n9414_ = new_n660_ & ~new_n9413_;
  assign new_n9415_ = new_n664_ & ~new_n9414_;
  assign new_n9416_ = new_n668_ & ~new_n9415_;
  assign new_n9417_ = new_n672_ & ~new_n9416_;
  assign new_n9418_ = new_n676_ & ~new_n9417_;
  assign new_n9419_ = new_n680_ & ~new_n9418_;
  assign new_n9420_ = new_n684_ & ~new_n9419_;
  assign new_n9421_ = new_n688_ & ~new_n9420_;
  assign new_n9422_ = new_n692_ & ~new_n9421_;
  assign new_n9423_ = new_n696_ & ~new_n9422_;
  assign new_n9424_ = new_n700_ & ~new_n9423_;
  assign new_n9425_ = new_n704_ & ~new_n9424_;
  assign new_n9426_ = new_n708_ & ~new_n9425_;
  assign new_n9427_ = new_n712_ & ~new_n9426_;
  assign new_n9428_ = new_n716_ & ~new_n9427_;
  assign new_n9429_ = new_n720_ & ~new_n9428_;
  assign new_n9430_ = new_n1484_ & ~new_n9429_;
  assign new_n9431_ = new_n1486_ & ~new_n9430_;
  assign new_n9432_ = new_n1750_ & ~new_n9431_;
  assign new_n9433_ = new_n731_ & ~new_n9432_;
  assign new_n9434_ = new_n735_ & ~new_n9433_;
  assign new_n9435_ = new_n739_ & ~new_n9434_;
  assign new_n9436_ = new_n743_ & ~new_n9435_;
  assign new_n9437_ = new_n747_ & ~new_n9436_;
  assign new_n9438_ = new_n751_ & ~new_n9437_;
  assign new_n9439_ = new_n755_ & ~new_n9438_;
  assign new_n9440_ = new_n759_ & ~new_n9439_;
  assign new_n9441_ = new_n763_ & ~new_n9440_;
  assign new_n9442_ = new_n767_ & ~new_n9441_;
  assign new_n9443_ = new_n771_ & ~new_n9442_;
  assign new_n9444_ = new_n775_ & ~new_n9443_;
  assign new_n9445_ = new_n779_ & ~new_n9444_;
  assign new_n9446_ = new_n783_ & ~new_n9445_;
  assign new_n9447_ = new_n787_ & ~new_n9446_;
  assign new_n9448_ = new_n791_ & ~new_n9447_;
  assign new_n9449_ = new_n795_ & ~new_n9448_;
  assign new_n9450_ = new_n799_ & ~new_n9449_;
  assign new_n9451_ = new_n803_ & ~new_n9450_;
  assign new_n9452_ = new_n807_ & ~new_n9451_;
  assign new_n9453_ = new_n811_ & ~new_n9452_;
  assign new_n9454_ = new_n815_ & ~new_n9453_;
  assign new_n9455_ = new_n819_ & ~new_n9454_;
  assign new_n9456_ = new_n823_ & ~new_n9455_;
  assign new_n9457_ = new_n827_ & ~new_n9456_;
  assign new_n9458_ = new_n831_ & ~new_n9457_;
  assign new_n9459_ = new_n835_ & ~new_n9458_;
  assign new_n9460_ = new_n839_ & ~new_n9459_;
  assign new_n9461_ = new_n843_ & ~new_n9460_;
  assign new_n9462_ = new_n847_ & ~new_n9461_;
  assign new_n9463_ = new_n851_ & ~new_n9462_;
  assign new_n9464_ = new_n855_ & ~new_n9463_;
  assign new_n9465_ = new_n859_ & ~new_n9464_;
  assign new_n9466_ = new_n863_ & ~new_n9465_;
  assign new_n9467_ = new_n867_ & ~new_n9466_;
  assign new_n9468_ = new_n871_ & ~new_n9467_;
  assign new_n9469_ = new_n875_ & ~new_n9468_;
  assign new_n9470_ = new_n879_ & ~new_n9469_;
  assign new_n9471_ = new_n883_ & ~new_n9470_;
  assign new_n9472_ = new_n887_ & ~new_n9471_;
  assign new_n9473_ = new_n891_ & ~new_n9472_;
  assign new_n9474_ = new_n895_ & ~new_n9473_;
  assign new_n9475_ = new_n899_ & ~new_n9474_;
  assign new_n9476_ = new_n903_ & ~new_n9475_;
  assign new_n9477_ = new_n907_ & ~new_n9476_;
  assign new_n9478_ = new_n911_ & ~new_n9477_;
  assign new_n9479_ = new_n915_ & ~new_n9478_;
  assign new_n9480_ = new_n919_ & ~new_n9479_;
  assign new_n9481_ = new_n923_ & ~new_n9480_;
  assign new_n9482_ = new_n927_ & ~new_n9481_;
  assign new_n9483_ = new_n931_ & ~new_n9482_;
  assign new_n9484_ = new_n935_ & ~new_n9483_;
  assign new_n9485_ = new_n939_ & ~new_n9484_;
  assign new_n9486_ = new_n943_ & ~new_n9485_;
  assign new_n9487_ = new_n947_ & ~new_n9486_;
  assign new_n9488_ = new_n951_ & ~new_n9487_;
  assign new_n9489_ = new_n955_ & ~new_n9488_;
  assign new_n9490_ = new_n959_ & ~new_n9489_;
  assign new_n9491_ = new_n963_ & ~new_n9490_;
  assign new_n9492_ = new_n967_ & ~new_n9491_;
  assign new_n9493_ = new_n971_ & ~new_n9492_;
  assign new_n9494_ = \req[96]  & ~new_n973_;
  assign \grant[96]  = ~new_n9493_ & new_n9494_;
  assign new_n9496_ = new_n982_ & ~new_n1315_;
  assign new_n9497_ = new_n987_ & ~new_n9496_;
  assign new_n9498_ = new_n991_ & ~new_n9497_;
  assign new_n9499_ = new_n995_ & ~new_n9498_;
  assign new_n9500_ = new_n999_ & ~new_n9499_;
  assign new_n9501_ = new_n1003_ & ~new_n9500_;
  assign new_n9502_ = new_n1007_ & ~new_n9501_;
  assign new_n9503_ = new_n1011_ & ~new_n9502_;
  assign new_n9504_ = new_n1015_ & ~new_n9503_;
  assign new_n9505_ = new_n1019_ & ~new_n9504_;
  assign new_n9506_ = new_n1023_ & ~new_n9505_;
  assign new_n9507_ = new_n1027_ & ~new_n9506_;
  assign new_n9508_ = new_n1031_ & ~new_n9507_;
  assign new_n9509_ = new_n1035_ & ~new_n9508_;
  assign new_n9510_ = new_n1039_ & ~new_n9509_;
  assign new_n9511_ = new_n1043_ & ~new_n9510_;
  assign new_n9512_ = new_n1047_ & ~new_n9511_;
  assign new_n9513_ = new_n1051_ & ~new_n9512_;
  assign new_n9514_ = new_n1055_ & ~new_n9513_;
  assign new_n9515_ = new_n1059_ & ~new_n9514_;
  assign new_n9516_ = new_n1574_ & ~new_n9515_;
  assign new_n9517_ = new_n1576_ & ~new_n9516_;
  assign new_n9518_ = new_n1837_ & ~new_n9517_;
  assign new_n9519_ = new_n1068_ & ~new_n9518_;
  assign new_n9520_ = new_n1072_ & ~new_n9519_;
  assign new_n9521_ = new_n1076_ & ~new_n9520_;
  assign new_n9522_ = new_n1080_ & ~new_n9521_;
  assign new_n9523_ = new_n1084_ & ~new_n9522_;
  assign new_n9524_ = new_n1088_ & ~new_n9523_;
  assign new_n9525_ = new_n1092_ & ~new_n9524_;
  assign new_n9526_ = new_n1096_ & ~new_n9525_;
  assign new_n9527_ = new_n1100_ & ~new_n9526_;
  assign new_n9528_ = new_n1104_ & ~new_n9527_;
  assign new_n9529_ = new_n1108_ & ~new_n9528_;
  assign new_n9530_ = new_n1112_ & ~new_n9529_;
  assign new_n9531_ = new_n1116_ & ~new_n9530_;
  assign new_n9532_ = new_n1120_ & ~new_n9531_;
  assign new_n9533_ = new_n1124_ & ~new_n9532_;
  assign new_n9534_ = new_n1128_ & ~new_n9533_;
  assign new_n9535_ = new_n1132_ & ~new_n9534_;
  assign new_n9536_ = new_n1136_ & ~new_n9535_;
  assign new_n9537_ = new_n1140_ & ~new_n9536_;
  assign new_n9538_ = new_n1144_ & ~new_n9537_;
  assign new_n9539_ = new_n1148_ & ~new_n9538_;
  assign new_n9540_ = new_n1152_ & ~new_n9539_;
  assign new_n9541_ = new_n1156_ & ~new_n9540_;
  assign new_n9542_ = new_n1160_ & ~new_n9541_;
  assign new_n9543_ = new_n1164_ & ~new_n9542_;
  assign new_n9544_ = new_n1168_ & ~new_n9543_;
  assign new_n9545_ = new_n1172_ & ~new_n9544_;
  assign new_n9546_ = new_n1176_ & ~new_n9545_;
  assign new_n9547_ = new_n1180_ & ~new_n9546_;
  assign new_n9548_ = new_n1184_ & ~new_n9547_;
  assign new_n9549_ = new_n1188_ & ~new_n9548_;
  assign new_n9550_ = new_n1192_ & ~new_n9549_;
  assign new_n9551_ = new_n1196_ & ~new_n9550_;
  assign new_n9552_ = new_n1200_ & ~new_n9551_;
  assign new_n9553_ = new_n1204_ & ~new_n9552_;
  assign new_n9554_ = new_n1208_ & ~new_n9553_;
  assign new_n9555_ = new_n1212_ & ~new_n9554_;
  assign new_n9556_ = new_n1216_ & ~new_n9555_;
  assign new_n9557_ = new_n1220_ & ~new_n9556_;
  assign new_n9558_ = new_n1224_ & ~new_n9557_;
  assign new_n9559_ = new_n1228_ & ~new_n9558_;
  assign new_n9560_ = new_n1232_ & ~new_n9559_;
  assign new_n9561_ = new_n1236_ & ~new_n9560_;
  assign new_n9562_ = new_n1240_ & ~new_n9561_;
  assign new_n9563_ = new_n1244_ & ~new_n9562_;
  assign new_n9564_ = new_n1248_ & ~new_n9563_;
  assign new_n9565_ = new_n1252_ & ~new_n9564_;
  assign new_n9566_ = new_n1256_ & ~new_n9565_;
  assign new_n9567_ = new_n1260_ & ~new_n9566_;
  assign new_n9568_ = new_n1264_ & ~new_n9567_;
  assign new_n9569_ = new_n1268_ & ~new_n9568_;
  assign new_n9570_ = new_n1272_ & ~new_n9569_;
  assign new_n9571_ = new_n1276_ & ~new_n9570_;
  assign new_n9572_ = new_n1280_ & ~new_n9571_;
  assign new_n9573_ = new_n1284_ & ~new_n9572_;
  assign new_n9574_ = new_n1288_ & ~new_n9573_;
  assign new_n9575_ = new_n1292_ & ~new_n9574_;
  assign new_n9576_ = new_n1296_ & ~new_n9575_;
  assign new_n9577_ = new_n1300_ & ~new_n9576_;
  assign new_n9578_ = new_n1304_ & ~new_n9577_;
  assign new_n9579_ = new_n1308_ & ~new_n9578_;
  assign new_n9580_ = \req[97]  & ~new_n1310_;
  assign \grant[97]  = ~new_n9579_ & new_n9580_;
  assign new_n9582_ = ~new_n647_ & new_n1319_;
  assign new_n9583_ = new_n1324_ & ~new_n9582_;
  assign new_n9584_ = new_n1328_ & ~new_n9583_;
  assign new_n9585_ = new_n1332_ & ~new_n9584_;
  assign new_n9586_ = new_n1336_ & ~new_n9585_;
  assign new_n9587_ = new_n1340_ & ~new_n9586_;
  assign new_n9588_ = new_n1344_ & ~new_n9587_;
  assign new_n9589_ = new_n1348_ & ~new_n9588_;
  assign new_n9590_ = new_n1352_ & ~new_n9589_;
  assign new_n9591_ = new_n1356_ & ~new_n9590_;
  assign new_n9592_ = new_n1360_ & ~new_n9591_;
  assign new_n9593_ = new_n1364_ & ~new_n9592_;
  assign new_n9594_ = new_n1368_ & ~new_n9593_;
  assign new_n9595_ = new_n1372_ & ~new_n9594_;
  assign new_n9596_ = new_n1376_ & ~new_n9595_;
  assign new_n9597_ = new_n1380_ & ~new_n9596_;
  assign new_n9598_ = new_n1384_ & ~new_n9597_;
  assign new_n9599_ = new_n1388_ & ~new_n9598_;
  assign new_n9600_ = new_n1392_ & ~new_n9599_;
  assign new_n9601_ = new_n1396_ & ~new_n9600_;
  assign new_n9602_ = new_n1663_ & ~new_n9601_;
  assign new_n9603_ = new_n392_ & ~new_n9602_;
  assign new_n9604_ = new_n396_ & ~new_n9603_;
  assign new_n9605_ = new_n400_ & ~new_n9604_;
  assign new_n9606_ = new_n404_ & ~new_n9605_;
  assign new_n9607_ = new_n408_ & ~new_n9606_;
  assign new_n9608_ = new_n412_ & ~new_n9607_;
  assign new_n9609_ = new_n416_ & ~new_n9608_;
  assign new_n9610_ = new_n420_ & ~new_n9609_;
  assign new_n9611_ = new_n424_ & ~new_n9610_;
  assign new_n9612_ = new_n428_ & ~new_n9611_;
  assign new_n9613_ = new_n432_ & ~new_n9612_;
  assign new_n9614_ = new_n436_ & ~new_n9613_;
  assign new_n9615_ = new_n440_ & ~new_n9614_;
  assign new_n9616_ = new_n444_ & ~new_n9615_;
  assign new_n9617_ = new_n448_ & ~new_n9616_;
  assign new_n9618_ = new_n452_ & ~new_n9617_;
  assign new_n9619_ = new_n456_ & ~new_n9618_;
  assign new_n9620_ = new_n460_ & ~new_n9619_;
  assign new_n9621_ = new_n464_ & ~new_n9620_;
  assign new_n9622_ = new_n468_ & ~new_n9621_;
  assign new_n9623_ = new_n472_ & ~new_n9622_;
  assign new_n9624_ = new_n476_ & ~new_n9623_;
  assign new_n9625_ = new_n480_ & ~new_n9624_;
  assign new_n9626_ = new_n484_ & ~new_n9625_;
  assign new_n9627_ = new_n488_ & ~new_n9626_;
  assign new_n9628_ = new_n492_ & ~new_n9627_;
  assign new_n9629_ = new_n496_ & ~new_n9628_;
  assign new_n9630_ = new_n500_ & ~new_n9629_;
  assign new_n9631_ = new_n504_ & ~new_n9630_;
  assign new_n9632_ = new_n508_ & ~new_n9631_;
  assign new_n9633_ = new_n512_ & ~new_n9632_;
  assign new_n9634_ = new_n516_ & ~new_n9633_;
  assign new_n9635_ = new_n520_ & ~new_n9634_;
  assign new_n9636_ = new_n524_ & ~new_n9635_;
  assign new_n9637_ = new_n528_ & ~new_n9636_;
  assign new_n9638_ = new_n532_ & ~new_n9637_;
  assign new_n9639_ = new_n536_ & ~new_n9638_;
  assign new_n9640_ = new_n540_ & ~new_n9639_;
  assign new_n9641_ = new_n544_ & ~new_n9640_;
  assign new_n9642_ = new_n548_ & ~new_n9641_;
  assign new_n9643_ = new_n552_ & ~new_n9642_;
  assign new_n9644_ = new_n556_ & ~new_n9643_;
  assign new_n9645_ = new_n560_ & ~new_n9644_;
  assign new_n9646_ = new_n564_ & ~new_n9645_;
  assign new_n9647_ = new_n568_ & ~new_n9646_;
  assign new_n9648_ = new_n572_ & ~new_n9647_;
  assign new_n9649_ = new_n576_ & ~new_n9648_;
  assign new_n9650_ = new_n580_ & ~new_n9649_;
  assign new_n9651_ = new_n584_ & ~new_n9650_;
  assign new_n9652_ = new_n588_ & ~new_n9651_;
  assign new_n9653_ = new_n592_ & ~new_n9652_;
  assign new_n9654_ = new_n596_ & ~new_n9653_;
  assign new_n9655_ = new_n600_ & ~new_n9654_;
  assign new_n9656_ = new_n604_ & ~new_n9655_;
  assign new_n9657_ = new_n608_ & ~new_n9656_;
  assign new_n9658_ = new_n612_ & ~new_n9657_;
  assign new_n9659_ = new_n616_ & ~new_n9658_;
  assign new_n9660_ = new_n620_ & ~new_n9659_;
  assign new_n9661_ = new_n624_ & ~new_n9660_;
  assign new_n9662_ = new_n628_ & ~new_n9661_;
  assign new_n9663_ = new_n632_ & ~new_n9662_;
  assign new_n9664_ = new_n636_ & ~new_n9663_;
  assign new_n9665_ = new_n640_ & ~new_n9664_;
  assign new_n9666_ = \req[98]  & ~new_n642_;
  assign \grant[98]  = ~new_n9665_ & new_n9666_;
  assign new_n9668_ = new_n651_ & ~new_n986_;
  assign new_n9669_ = new_n656_ & ~new_n9668_;
  assign new_n9670_ = new_n660_ & ~new_n9669_;
  assign new_n9671_ = new_n664_ & ~new_n9670_;
  assign new_n9672_ = new_n668_ & ~new_n9671_;
  assign new_n9673_ = new_n672_ & ~new_n9672_;
  assign new_n9674_ = new_n676_ & ~new_n9673_;
  assign new_n9675_ = new_n680_ & ~new_n9674_;
  assign new_n9676_ = new_n684_ & ~new_n9675_;
  assign new_n9677_ = new_n688_ & ~new_n9676_;
  assign new_n9678_ = new_n692_ & ~new_n9677_;
  assign new_n9679_ = new_n696_ & ~new_n9678_;
  assign new_n9680_ = new_n700_ & ~new_n9679_;
  assign new_n9681_ = new_n704_ & ~new_n9680_;
  assign new_n9682_ = new_n708_ & ~new_n9681_;
  assign new_n9683_ = new_n712_ & ~new_n9682_;
  assign new_n9684_ = new_n716_ & ~new_n9683_;
  assign new_n9685_ = new_n720_ & ~new_n9684_;
  assign new_n9686_ = new_n1484_ & ~new_n9685_;
  assign new_n9687_ = new_n1486_ & ~new_n9686_;
  assign new_n9688_ = new_n1750_ & ~new_n9687_;
  assign new_n9689_ = new_n731_ & ~new_n9688_;
  assign new_n9690_ = new_n735_ & ~new_n9689_;
  assign new_n9691_ = new_n739_ & ~new_n9690_;
  assign new_n9692_ = new_n743_ & ~new_n9691_;
  assign new_n9693_ = new_n747_ & ~new_n9692_;
  assign new_n9694_ = new_n751_ & ~new_n9693_;
  assign new_n9695_ = new_n755_ & ~new_n9694_;
  assign new_n9696_ = new_n759_ & ~new_n9695_;
  assign new_n9697_ = new_n763_ & ~new_n9696_;
  assign new_n9698_ = new_n767_ & ~new_n9697_;
  assign new_n9699_ = new_n771_ & ~new_n9698_;
  assign new_n9700_ = new_n775_ & ~new_n9699_;
  assign new_n9701_ = new_n779_ & ~new_n9700_;
  assign new_n9702_ = new_n783_ & ~new_n9701_;
  assign new_n9703_ = new_n787_ & ~new_n9702_;
  assign new_n9704_ = new_n791_ & ~new_n9703_;
  assign new_n9705_ = new_n795_ & ~new_n9704_;
  assign new_n9706_ = new_n799_ & ~new_n9705_;
  assign new_n9707_ = new_n803_ & ~new_n9706_;
  assign new_n9708_ = new_n807_ & ~new_n9707_;
  assign new_n9709_ = new_n811_ & ~new_n9708_;
  assign new_n9710_ = new_n815_ & ~new_n9709_;
  assign new_n9711_ = new_n819_ & ~new_n9710_;
  assign new_n9712_ = new_n823_ & ~new_n9711_;
  assign new_n9713_ = new_n827_ & ~new_n9712_;
  assign new_n9714_ = new_n831_ & ~new_n9713_;
  assign new_n9715_ = new_n835_ & ~new_n9714_;
  assign new_n9716_ = new_n839_ & ~new_n9715_;
  assign new_n9717_ = new_n843_ & ~new_n9716_;
  assign new_n9718_ = new_n847_ & ~new_n9717_;
  assign new_n9719_ = new_n851_ & ~new_n9718_;
  assign new_n9720_ = new_n855_ & ~new_n9719_;
  assign new_n9721_ = new_n859_ & ~new_n9720_;
  assign new_n9722_ = new_n863_ & ~new_n9721_;
  assign new_n9723_ = new_n867_ & ~new_n9722_;
  assign new_n9724_ = new_n871_ & ~new_n9723_;
  assign new_n9725_ = new_n875_ & ~new_n9724_;
  assign new_n9726_ = new_n879_ & ~new_n9725_;
  assign new_n9727_ = new_n883_ & ~new_n9726_;
  assign new_n9728_ = new_n887_ & ~new_n9727_;
  assign new_n9729_ = new_n891_ & ~new_n9728_;
  assign new_n9730_ = new_n895_ & ~new_n9729_;
  assign new_n9731_ = new_n899_ & ~new_n9730_;
  assign new_n9732_ = new_n903_ & ~new_n9731_;
  assign new_n9733_ = new_n907_ & ~new_n9732_;
  assign new_n9734_ = new_n911_ & ~new_n9733_;
  assign new_n9735_ = new_n915_ & ~new_n9734_;
  assign new_n9736_ = new_n919_ & ~new_n9735_;
  assign new_n9737_ = new_n923_ & ~new_n9736_;
  assign new_n9738_ = new_n927_ & ~new_n9737_;
  assign new_n9739_ = new_n931_ & ~new_n9738_;
  assign new_n9740_ = new_n935_ & ~new_n9739_;
  assign new_n9741_ = new_n939_ & ~new_n9740_;
  assign new_n9742_ = new_n943_ & ~new_n9741_;
  assign new_n9743_ = new_n947_ & ~new_n9742_;
  assign new_n9744_ = new_n951_ & ~new_n9743_;
  assign new_n9745_ = new_n955_ & ~new_n9744_;
  assign new_n9746_ = new_n959_ & ~new_n9745_;
  assign new_n9747_ = new_n963_ & ~new_n9746_;
  assign new_n9748_ = new_n967_ & ~new_n9747_;
  assign new_n9749_ = new_n971_ & ~new_n9748_;
  assign new_n9750_ = new_n975_ & ~new_n9749_;
  assign new_n9751_ = new_n979_ & ~new_n9750_;
  assign new_n9752_ = \req[99]  & ~new_n981_;
  assign \grant[99]  = ~new_n9751_ & new_n9752_;
  assign new_n9754_ = new_n990_ & ~new_n1323_;
  assign new_n9755_ = new_n995_ & ~new_n9754_;
  assign new_n9756_ = new_n999_ & ~new_n9755_;
  assign new_n9757_ = new_n1003_ & ~new_n9756_;
  assign new_n9758_ = new_n1007_ & ~new_n9757_;
  assign new_n9759_ = new_n1011_ & ~new_n9758_;
  assign new_n9760_ = new_n1015_ & ~new_n9759_;
  assign new_n9761_ = new_n1019_ & ~new_n9760_;
  assign new_n9762_ = new_n1023_ & ~new_n9761_;
  assign new_n9763_ = new_n1027_ & ~new_n9762_;
  assign new_n9764_ = new_n1031_ & ~new_n9763_;
  assign new_n9765_ = new_n1035_ & ~new_n9764_;
  assign new_n9766_ = new_n1039_ & ~new_n9765_;
  assign new_n9767_ = new_n1043_ & ~new_n9766_;
  assign new_n9768_ = new_n1047_ & ~new_n9767_;
  assign new_n9769_ = new_n1051_ & ~new_n9768_;
  assign new_n9770_ = new_n1055_ & ~new_n9769_;
  assign new_n9771_ = new_n1059_ & ~new_n9770_;
  assign new_n9772_ = new_n1574_ & ~new_n9771_;
  assign new_n9773_ = new_n1576_ & ~new_n9772_;
  assign new_n9774_ = new_n1837_ & ~new_n9773_;
  assign new_n9775_ = new_n1068_ & ~new_n9774_;
  assign new_n9776_ = new_n1072_ & ~new_n9775_;
  assign new_n9777_ = new_n1076_ & ~new_n9776_;
  assign new_n9778_ = new_n1080_ & ~new_n9777_;
  assign new_n9779_ = new_n1084_ & ~new_n9778_;
  assign new_n9780_ = new_n1088_ & ~new_n9779_;
  assign new_n9781_ = new_n1092_ & ~new_n9780_;
  assign new_n9782_ = new_n1096_ & ~new_n9781_;
  assign new_n9783_ = new_n1100_ & ~new_n9782_;
  assign new_n9784_ = new_n1104_ & ~new_n9783_;
  assign new_n9785_ = new_n1108_ & ~new_n9784_;
  assign new_n9786_ = new_n1112_ & ~new_n9785_;
  assign new_n9787_ = new_n1116_ & ~new_n9786_;
  assign new_n9788_ = new_n1120_ & ~new_n9787_;
  assign new_n9789_ = new_n1124_ & ~new_n9788_;
  assign new_n9790_ = new_n1128_ & ~new_n9789_;
  assign new_n9791_ = new_n1132_ & ~new_n9790_;
  assign new_n9792_ = new_n1136_ & ~new_n9791_;
  assign new_n9793_ = new_n1140_ & ~new_n9792_;
  assign new_n9794_ = new_n1144_ & ~new_n9793_;
  assign new_n9795_ = new_n1148_ & ~new_n9794_;
  assign new_n9796_ = new_n1152_ & ~new_n9795_;
  assign new_n9797_ = new_n1156_ & ~new_n9796_;
  assign new_n9798_ = new_n1160_ & ~new_n9797_;
  assign new_n9799_ = new_n1164_ & ~new_n9798_;
  assign new_n9800_ = new_n1168_ & ~new_n9799_;
  assign new_n9801_ = new_n1172_ & ~new_n9800_;
  assign new_n9802_ = new_n1176_ & ~new_n9801_;
  assign new_n9803_ = new_n1180_ & ~new_n9802_;
  assign new_n9804_ = new_n1184_ & ~new_n9803_;
  assign new_n9805_ = new_n1188_ & ~new_n9804_;
  assign new_n9806_ = new_n1192_ & ~new_n9805_;
  assign new_n9807_ = new_n1196_ & ~new_n9806_;
  assign new_n9808_ = new_n1200_ & ~new_n9807_;
  assign new_n9809_ = new_n1204_ & ~new_n9808_;
  assign new_n9810_ = new_n1208_ & ~new_n9809_;
  assign new_n9811_ = new_n1212_ & ~new_n9810_;
  assign new_n9812_ = new_n1216_ & ~new_n9811_;
  assign new_n9813_ = new_n1220_ & ~new_n9812_;
  assign new_n9814_ = new_n1224_ & ~new_n9813_;
  assign new_n9815_ = new_n1228_ & ~new_n9814_;
  assign new_n9816_ = new_n1232_ & ~new_n9815_;
  assign new_n9817_ = new_n1236_ & ~new_n9816_;
  assign new_n9818_ = new_n1240_ & ~new_n9817_;
  assign new_n9819_ = new_n1244_ & ~new_n9818_;
  assign new_n9820_ = new_n1248_ & ~new_n9819_;
  assign new_n9821_ = new_n1252_ & ~new_n9820_;
  assign new_n9822_ = new_n1256_ & ~new_n9821_;
  assign new_n9823_ = new_n1260_ & ~new_n9822_;
  assign new_n9824_ = new_n1264_ & ~new_n9823_;
  assign new_n9825_ = new_n1268_ & ~new_n9824_;
  assign new_n9826_ = new_n1272_ & ~new_n9825_;
  assign new_n9827_ = new_n1276_ & ~new_n9826_;
  assign new_n9828_ = new_n1280_ & ~new_n9827_;
  assign new_n9829_ = new_n1284_ & ~new_n9828_;
  assign new_n9830_ = new_n1288_ & ~new_n9829_;
  assign new_n9831_ = new_n1292_ & ~new_n9830_;
  assign new_n9832_ = new_n1296_ & ~new_n9831_;
  assign new_n9833_ = new_n1300_ & ~new_n9832_;
  assign new_n9834_ = new_n1304_ & ~new_n9833_;
  assign new_n9835_ = new_n1308_ & ~new_n9834_;
  assign new_n9836_ = new_n1312_ & ~new_n9835_;
  assign new_n9837_ = new_n1316_ & ~new_n9836_;
  assign new_n9838_ = \req[100]  & ~new_n1318_;
  assign \grant[100]  = ~new_n9837_ & new_n9838_;
  assign new_n9840_ = ~new_n655_ & new_n1327_;
  assign new_n9841_ = new_n1332_ & ~new_n9840_;
  assign new_n9842_ = new_n1336_ & ~new_n9841_;
  assign new_n9843_ = new_n1340_ & ~new_n9842_;
  assign new_n9844_ = new_n1344_ & ~new_n9843_;
  assign new_n9845_ = new_n1348_ & ~new_n9844_;
  assign new_n9846_ = new_n1352_ & ~new_n9845_;
  assign new_n9847_ = new_n1356_ & ~new_n9846_;
  assign new_n9848_ = new_n1360_ & ~new_n9847_;
  assign new_n9849_ = new_n1364_ & ~new_n9848_;
  assign new_n9850_ = new_n1368_ & ~new_n9849_;
  assign new_n9851_ = new_n1372_ & ~new_n9850_;
  assign new_n9852_ = new_n1376_ & ~new_n9851_;
  assign new_n9853_ = new_n1380_ & ~new_n9852_;
  assign new_n9854_ = new_n1384_ & ~new_n9853_;
  assign new_n9855_ = new_n1388_ & ~new_n9854_;
  assign new_n9856_ = new_n1392_ & ~new_n9855_;
  assign new_n9857_ = new_n1396_ & ~new_n9856_;
  assign new_n9858_ = new_n1663_ & ~new_n9857_;
  assign new_n9859_ = new_n392_ & ~new_n9858_;
  assign new_n9860_ = new_n396_ & ~new_n9859_;
  assign new_n9861_ = new_n400_ & ~new_n9860_;
  assign new_n9862_ = new_n404_ & ~new_n9861_;
  assign new_n9863_ = new_n408_ & ~new_n9862_;
  assign new_n9864_ = new_n412_ & ~new_n9863_;
  assign new_n9865_ = new_n416_ & ~new_n9864_;
  assign new_n9866_ = new_n420_ & ~new_n9865_;
  assign new_n9867_ = new_n424_ & ~new_n9866_;
  assign new_n9868_ = new_n428_ & ~new_n9867_;
  assign new_n9869_ = new_n432_ & ~new_n9868_;
  assign new_n9870_ = new_n436_ & ~new_n9869_;
  assign new_n9871_ = new_n440_ & ~new_n9870_;
  assign new_n9872_ = new_n444_ & ~new_n9871_;
  assign new_n9873_ = new_n448_ & ~new_n9872_;
  assign new_n9874_ = new_n452_ & ~new_n9873_;
  assign new_n9875_ = new_n456_ & ~new_n9874_;
  assign new_n9876_ = new_n460_ & ~new_n9875_;
  assign new_n9877_ = new_n464_ & ~new_n9876_;
  assign new_n9878_ = new_n468_ & ~new_n9877_;
  assign new_n9879_ = new_n472_ & ~new_n9878_;
  assign new_n9880_ = new_n476_ & ~new_n9879_;
  assign new_n9881_ = new_n480_ & ~new_n9880_;
  assign new_n9882_ = new_n484_ & ~new_n9881_;
  assign new_n9883_ = new_n488_ & ~new_n9882_;
  assign new_n9884_ = new_n492_ & ~new_n9883_;
  assign new_n9885_ = new_n496_ & ~new_n9884_;
  assign new_n9886_ = new_n500_ & ~new_n9885_;
  assign new_n9887_ = new_n504_ & ~new_n9886_;
  assign new_n9888_ = new_n508_ & ~new_n9887_;
  assign new_n9889_ = new_n512_ & ~new_n9888_;
  assign new_n9890_ = new_n516_ & ~new_n9889_;
  assign new_n9891_ = new_n520_ & ~new_n9890_;
  assign new_n9892_ = new_n524_ & ~new_n9891_;
  assign new_n9893_ = new_n528_ & ~new_n9892_;
  assign new_n9894_ = new_n532_ & ~new_n9893_;
  assign new_n9895_ = new_n536_ & ~new_n9894_;
  assign new_n9896_ = new_n540_ & ~new_n9895_;
  assign new_n9897_ = new_n544_ & ~new_n9896_;
  assign new_n9898_ = new_n548_ & ~new_n9897_;
  assign new_n9899_ = new_n552_ & ~new_n9898_;
  assign new_n9900_ = new_n556_ & ~new_n9899_;
  assign new_n9901_ = new_n560_ & ~new_n9900_;
  assign new_n9902_ = new_n564_ & ~new_n9901_;
  assign new_n9903_ = new_n568_ & ~new_n9902_;
  assign new_n9904_ = new_n572_ & ~new_n9903_;
  assign new_n9905_ = new_n576_ & ~new_n9904_;
  assign new_n9906_ = new_n580_ & ~new_n9905_;
  assign new_n9907_ = new_n584_ & ~new_n9906_;
  assign new_n9908_ = new_n588_ & ~new_n9907_;
  assign new_n9909_ = new_n592_ & ~new_n9908_;
  assign new_n9910_ = new_n596_ & ~new_n9909_;
  assign new_n9911_ = new_n600_ & ~new_n9910_;
  assign new_n9912_ = new_n604_ & ~new_n9911_;
  assign new_n9913_ = new_n608_ & ~new_n9912_;
  assign new_n9914_ = new_n612_ & ~new_n9913_;
  assign new_n9915_ = new_n616_ & ~new_n9914_;
  assign new_n9916_ = new_n620_ & ~new_n9915_;
  assign new_n9917_ = new_n624_ & ~new_n9916_;
  assign new_n9918_ = new_n628_ & ~new_n9917_;
  assign new_n9919_ = new_n632_ & ~new_n9918_;
  assign new_n9920_ = new_n636_ & ~new_n9919_;
  assign new_n9921_ = new_n640_ & ~new_n9920_;
  assign new_n9922_ = new_n644_ & ~new_n9921_;
  assign new_n9923_ = new_n648_ & ~new_n9922_;
  assign new_n9924_ = \req[101]  & ~new_n650_;
  assign \grant[101]  = ~new_n9923_ & new_n9924_;
  assign new_n9926_ = new_n659_ & ~new_n994_;
  assign new_n9927_ = new_n664_ & ~new_n9926_;
  assign new_n9928_ = new_n668_ & ~new_n9927_;
  assign new_n9929_ = new_n672_ & ~new_n9928_;
  assign new_n9930_ = new_n676_ & ~new_n9929_;
  assign new_n9931_ = new_n680_ & ~new_n9930_;
  assign new_n9932_ = new_n684_ & ~new_n9931_;
  assign new_n9933_ = new_n688_ & ~new_n9932_;
  assign new_n9934_ = new_n692_ & ~new_n9933_;
  assign new_n9935_ = new_n696_ & ~new_n9934_;
  assign new_n9936_ = new_n700_ & ~new_n9935_;
  assign new_n9937_ = new_n704_ & ~new_n9936_;
  assign new_n9938_ = new_n708_ & ~new_n9937_;
  assign new_n9939_ = new_n712_ & ~new_n9938_;
  assign new_n9940_ = new_n716_ & ~new_n9939_;
  assign new_n9941_ = new_n720_ & ~new_n9940_;
  assign new_n9942_ = new_n1484_ & ~new_n9941_;
  assign new_n9943_ = new_n1486_ & ~new_n9942_;
  assign new_n9944_ = new_n1750_ & ~new_n9943_;
  assign new_n9945_ = new_n731_ & ~new_n9944_;
  assign new_n9946_ = new_n735_ & ~new_n9945_;
  assign new_n9947_ = new_n739_ & ~new_n9946_;
  assign new_n9948_ = new_n743_ & ~new_n9947_;
  assign new_n9949_ = new_n747_ & ~new_n9948_;
  assign new_n9950_ = new_n751_ & ~new_n9949_;
  assign new_n9951_ = new_n755_ & ~new_n9950_;
  assign new_n9952_ = new_n759_ & ~new_n9951_;
  assign new_n9953_ = new_n763_ & ~new_n9952_;
  assign new_n9954_ = new_n767_ & ~new_n9953_;
  assign new_n9955_ = new_n771_ & ~new_n9954_;
  assign new_n9956_ = new_n775_ & ~new_n9955_;
  assign new_n9957_ = new_n779_ & ~new_n9956_;
  assign new_n9958_ = new_n783_ & ~new_n9957_;
  assign new_n9959_ = new_n787_ & ~new_n9958_;
  assign new_n9960_ = new_n791_ & ~new_n9959_;
  assign new_n9961_ = new_n795_ & ~new_n9960_;
  assign new_n9962_ = new_n799_ & ~new_n9961_;
  assign new_n9963_ = new_n803_ & ~new_n9962_;
  assign new_n9964_ = new_n807_ & ~new_n9963_;
  assign new_n9965_ = new_n811_ & ~new_n9964_;
  assign new_n9966_ = new_n815_ & ~new_n9965_;
  assign new_n9967_ = new_n819_ & ~new_n9966_;
  assign new_n9968_ = new_n823_ & ~new_n9967_;
  assign new_n9969_ = new_n827_ & ~new_n9968_;
  assign new_n9970_ = new_n831_ & ~new_n9969_;
  assign new_n9971_ = new_n835_ & ~new_n9970_;
  assign new_n9972_ = new_n839_ & ~new_n9971_;
  assign new_n9973_ = new_n843_ & ~new_n9972_;
  assign new_n9974_ = new_n847_ & ~new_n9973_;
  assign new_n9975_ = new_n851_ & ~new_n9974_;
  assign new_n9976_ = new_n855_ & ~new_n9975_;
  assign new_n9977_ = new_n859_ & ~new_n9976_;
  assign new_n9978_ = new_n863_ & ~new_n9977_;
  assign new_n9979_ = new_n867_ & ~new_n9978_;
  assign new_n9980_ = new_n871_ & ~new_n9979_;
  assign new_n9981_ = new_n875_ & ~new_n9980_;
  assign new_n9982_ = new_n879_ & ~new_n9981_;
  assign new_n9983_ = new_n883_ & ~new_n9982_;
  assign new_n9984_ = new_n887_ & ~new_n9983_;
  assign new_n9985_ = new_n891_ & ~new_n9984_;
  assign new_n9986_ = new_n895_ & ~new_n9985_;
  assign new_n9987_ = new_n899_ & ~new_n9986_;
  assign new_n9988_ = new_n903_ & ~new_n9987_;
  assign new_n9989_ = new_n907_ & ~new_n9988_;
  assign new_n9990_ = new_n911_ & ~new_n9989_;
  assign new_n9991_ = new_n915_ & ~new_n9990_;
  assign new_n9992_ = new_n919_ & ~new_n9991_;
  assign new_n9993_ = new_n923_ & ~new_n9992_;
  assign new_n9994_ = new_n927_ & ~new_n9993_;
  assign new_n9995_ = new_n931_ & ~new_n9994_;
  assign new_n9996_ = new_n935_ & ~new_n9995_;
  assign new_n9997_ = new_n939_ & ~new_n9996_;
  assign new_n9998_ = new_n943_ & ~new_n9997_;
  assign new_n9999_ = new_n947_ & ~new_n9998_;
  assign new_n10000_ = new_n951_ & ~new_n9999_;
  assign new_n10001_ = new_n955_ & ~new_n10000_;
  assign new_n10002_ = new_n959_ & ~new_n10001_;
  assign new_n10003_ = new_n963_ & ~new_n10002_;
  assign new_n10004_ = new_n967_ & ~new_n10003_;
  assign new_n10005_ = new_n971_ & ~new_n10004_;
  assign new_n10006_ = new_n975_ & ~new_n10005_;
  assign new_n10007_ = new_n979_ & ~new_n10006_;
  assign new_n10008_ = new_n983_ & ~new_n10007_;
  assign new_n10009_ = new_n987_ & ~new_n10008_;
  assign new_n10010_ = \req[102]  & ~new_n989_;
  assign \grant[102]  = ~new_n10009_ & new_n10010_;
  assign new_n10012_ = new_n998_ & ~new_n1331_;
  assign new_n10013_ = new_n1003_ & ~new_n10012_;
  assign new_n10014_ = new_n1007_ & ~new_n10013_;
  assign new_n10015_ = new_n1011_ & ~new_n10014_;
  assign new_n10016_ = new_n1015_ & ~new_n10015_;
  assign new_n10017_ = new_n1019_ & ~new_n10016_;
  assign new_n10018_ = new_n1023_ & ~new_n10017_;
  assign new_n10019_ = new_n1027_ & ~new_n10018_;
  assign new_n10020_ = new_n1031_ & ~new_n10019_;
  assign new_n10021_ = new_n1035_ & ~new_n10020_;
  assign new_n10022_ = new_n1039_ & ~new_n10021_;
  assign new_n10023_ = new_n1043_ & ~new_n10022_;
  assign new_n10024_ = new_n1047_ & ~new_n10023_;
  assign new_n10025_ = new_n1051_ & ~new_n10024_;
  assign new_n10026_ = new_n1055_ & ~new_n10025_;
  assign new_n10027_ = new_n1059_ & ~new_n10026_;
  assign new_n10028_ = new_n1574_ & ~new_n10027_;
  assign new_n10029_ = new_n1576_ & ~new_n10028_;
  assign new_n10030_ = new_n1837_ & ~new_n10029_;
  assign new_n10031_ = new_n1068_ & ~new_n10030_;
  assign new_n10032_ = new_n1072_ & ~new_n10031_;
  assign new_n10033_ = new_n1076_ & ~new_n10032_;
  assign new_n10034_ = new_n1080_ & ~new_n10033_;
  assign new_n10035_ = new_n1084_ & ~new_n10034_;
  assign new_n10036_ = new_n1088_ & ~new_n10035_;
  assign new_n10037_ = new_n1092_ & ~new_n10036_;
  assign new_n10038_ = new_n1096_ & ~new_n10037_;
  assign new_n10039_ = new_n1100_ & ~new_n10038_;
  assign new_n10040_ = new_n1104_ & ~new_n10039_;
  assign new_n10041_ = new_n1108_ & ~new_n10040_;
  assign new_n10042_ = new_n1112_ & ~new_n10041_;
  assign new_n10043_ = new_n1116_ & ~new_n10042_;
  assign new_n10044_ = new_n1120_ & ~new_n10043_;
  assign new_n10045_ = new_n1124_ & ~new_n10044_;
  assign new_n10046_ = new_n1128_ & ~new_n10045_;
  assign new_n10047_ = new_n1132_ & ~new_n10046_;
  assign new_n10048_ = new_n1136_ & ~new_n10047_;
  assign new_n10049_ = new_n1140_ & ~new_n10048_;
  assign new_n10050_ = new_n1144_ & ~new_n10049_;
  assign new_n10051_ = new_n1148_ & ~new_n10050_;
  assign new_n10052_ = new_n1152_ & ~new_n10051_;
  assign new_n10053_ = new_n1156_ & ~new_n10052_;
  assign new_n10054_ = new_n1160_ & ~new_n10053_;
  assign new_n10055_ = new_n1164_ & ~new_n10054_;
  assign new_n10056_ = new_n1168_ & ~new_n10055_;
  assign new_n10057_ = new_n1172_ & ~new_n10056_;
  assign new_n10058_ = new_n1176_ & ~new_n10057_;
  assign new_n10059_ = new_n1180_ & ~new_n10058_;
  assign new_n10060_ = new_n1184_ & ~new_n10059_;
  assign new_n10061_ = new_n1188_ & ~new_n10060_;
  assign new_n10062_ = new_n1192_ & ~new_n10061_;
  assign new_n10063_ = new_n1196_ & ~new_n10062_;
  assign new_n10064_ = new_n1200_ & ~new_n10063_;
  assign new_n10065_ = new_n1204_ & ~new_n10064_;
  assign new_n10066_ = new_n1208_ & ~new_n10065_;
  assign new_n10067_ = new_n1212_ & ~new_n10066_;
  assign new_n10068_ = new_n1216_ & ~new_n10067_;
  assign new_n10069_ = new_n1220_ & ~new_n10068_;
  assign new_n10070_ = new_n1224_ & ~new_n10069_;
  assign new_n10071_ = new_n1228_ & ~new_n10070_;
  assign new_n10072_ = new_n1232_ & ~new_n10071_;
  assign new_n10073_ = new_n1236_ & ~new_n10072_;
  assign new_n10074_ = new_n1240_ & ~new_n10073_;
  assign new_n10075_ = new_n1244_ & ~new_n10074_;
  assign new_n10076_ = new_n1248_ & ~new_n10075_;
  assign new_n10077_ = new_n1252_ & ~new_n10076_;
  assign new_n10078_ = new_n1256_ & ~new_n10077_;
  assign new_n10079_ = new_n1260_ & ~new_n10078_;
  assign new_n10080_ = new_n1264_ & ~new_n10079_;
  assign new_n10081_ = new_n1268_ & ~new_n10080_;
  assign new_n10082_ = new_n1272_ & ~new_n10081_;
  assign new_n10083_ = new_n1276_ & ~new_n10082_;
  assign new_n10084_ = new_n1280_ & ~new_n10083_;
  assign new_n10085_ = new_n1284_ & ~new_n10084_;
  assign new_n10086_ = new_n1288_ & ~new_n10085_;
  assign new_n10087_ = new_n1292_ & ~new_n10086_;
  assign new_n10088_ = new_n1296_ & ~new_n10087_;
  assign new_n10089_ = new_n1300_ & ~new_n10088_;
  assign new_n10090_ = new_n1304_ & ~new_n10089_;
  assign new_n10091_ = new_n1308_ & ~new_n10090_;
  assign new_n10092_ = new_n1312_ & ~new_n10091_;
  assign new_n10093_ = new_n1316_ & ~new_n10092_;
  assign new_n10094_ = new_n1320_ & ~new_n10093_;
  assign new_n10095_ = new_n1324_ & ~new_n10094_;
  assign new_n10096_ = \req[103]  & ~new_n1326_;
  assign \grant[103]  = ~new_n10095_ & new_n10096_;
  assign new_n10098_ = ~new_n663_ & new_n1335_;
  assign new_n10099_ = new_n1340_ & ~new_n10098_;
  assign new_n10100_ = new_n1344_ & ~new_n10099_;
  assign new_n10101_ = new_n1348_ & ~new_n10100_;
  assign new_n10102_ = new_n1352_ & ~new_n10101_;
  assign new_n10103_ = new_n1356_ & ~new_n10102_;
  assign new_n10104_ = new_n1360_ & ~new_n10103_;
  assign new_n10105_ = new_n1364_ & ~new_n10104_;
  assign new_n10106_ = new_n1368_ & ~new_n10105_;
  assign new_n10107_ = new_n1372_ & ~new_n10106_;
  assign new_n10108_ = new_n1376_ & ~new_n10107_;
  assign new_n10109_ = new_n1380_ & ~new_n10108_;
  assign new_n10110_ = new_n1384_ & ~new_n10109_;
  assign new_n10111_ = new_n1388_ & ~new_n10110_;
  assign new_n10112_ = new_n1392_ & ~new_n10111_;
  assign new_n10113_ = new_n1396_ & ~new_n10112_;
  assign new_n10114_ = new_n1663_ & ~new_n10113_;
  assign new_n10115_ = new_n392_ & ~new_n10114_;
  assign new_n10116_ = new_n396_ & ~new_n10115_;
  assign new_n10117_ = new_n400_ & ~new_n10116_;
  assign new_n10118_ = new_n404_ & ~new_n10117_;
  assign new_n10119_ = new_n408_ & ~new_n10118_;
  assign new_n10120_ = new_n412_ & ~new_n10119_;
  assign new_n10121_ = new_n416_ & ~new_n10120_;
  assign new_n10122_ = new_n420_ & ~new_n10121_;
  assign new_n10123_ = new_n424_ & ~new_n10122_;
  assign new_n10124_ = new_n428_ & ~new_n10123_;
  assign new_n10125_ = new_n432_ & ~new_n10124_;
  assign new_n10126_ = new_n436_ & ~new_n10125_;
  assign new_n10127_ = new_n440_ & ~new_n10126_;
  assign new_n10128_ = new_n444_ & ~new_n10127_;
  assign new_n10129_ = new_n448_ & ~new_n10128_;
  assign new_n10130_ = new_n452_ & ~new_n10129_;
  assign new_n10131_ = new_n456_ & ~new_n10130_;
  assign new_n10132_ = new_n460_ & ~new_n10131_;
  assign new_n10133_ = new_n464_ & ~new_n10132_;
  assign new_n10134_ = new_n468_ & ~new_n10133_;
  assign new_n10135_ = new_n472_ & ~new_n10134_;
  assign new_n10136_ = new_n476_ & ~new_n10135_;
  assign new_n10137_ = new_n480_ & ~new_n10136_;
  assign new_n10138_ = new_n484_ & ~new_n10137_;
  assign new_n10139_ = new_n488_ & ~new_n10138_;
  assign new_n10140_ = new_n492_ & ~new_n10139_;
  assign new_n10141_ = new_n496_ & ~new_n10140_;
  assign new_n10142_ = new_n500_ & ~new_n10141_;
  assign new_n10143_ = new_n504_ & ~new_n10142_;
  assign new_n10144_ = new_n508_ & ~new_n10143_;
  assign new_n10145_ = new_n512_ & ~new_n10144_;
  assign new_n10146_ = new_n516_ & ~new_n10145_;
  assign new_n10147_ = new_n520_ & ~new_n10146_;
  assign new_n10148_ = new_n524_ & ~new_n10147_;
  assign new_n10149_ = new_n528_ & ~new_n10148_;
  assign new_n10150_ = new_n532_ & ~new_n10149_;
  assign new_n10151_ = new_n536_ & ~new_n10150_;
  assign new_n10152_ = new_n540_ & ~new_n10151_;
  assign new_n10153_ = new_n544_ & ~new_n10152_;
  assign new_n10154_ = new_n548_ & ~new_n10153_;
  assign new_n10155_ = new_n552_ & ~new_n10154_;
  assign new_n10156_ = new_n556_ & ~new_n10155_;
  assign new_n10157_ = new_n560_ & ~new_n10156_;
  assign new_n10158_ = new_n564_ & ~new_n10157_;
  assign new_n10159_ = new_n568_ & ~new_n10158_;
  assign new_n10160_ = new_n572_ & ~new_n10159_;
  assign new_n10161_ = new_n576_ & ~new_n10160_;
  assign new_n10162_ = new_n580_ & ~new_n10161_;
  assign new_n10163_ = new_n584_ & ~new_n10162_;
  assign new_n10164_ = new_n588_ & ~new_n10163_;
  assign new_n10165_ = new_n592_ & ~new_n10164_;
  assign new_n10166_ = new_n596_ & ~new_n10165_;
  assign new_n10167_ = new_n600_ & ~new_n10166_;
  assign new_n10168_ = new_n604_ & ~new_n10167_;
  assign new_n10169_ = new_n608_ & ~new_n10168_;
  assign new_n10170_ = new_n612_ & ~new_n10169_;
  assign new_n10171_ = new_n616_ & ~new_n10170_;
  assign new_n10172_ = new_n620_ & ~new_n10171_;
  assign new_n10173_ = new_n624_ & ~new_n10172_;
  assign new_n10174_ = new_n628_ & ~new_n10173_;
  assign new_n10175_ = new_n632_ & ~new_n10174_;
  assign new_n10176_ = new_n636_ & ~new_n10175_;
  assign new_n10177_ = new_n640_ & ~new_n10176_;
  assign new_n10178_ = new_n644_ & ~new_n10177_;
  assign new_n10179_ = new_n648_ & ~new_n10178_;
  assign new_n10180_ = new_n652_ & ~new_n10179_;
  assign new_n10181_ = new_n656_ & ~new_n10180_;
  assign new_n10182_ = \req[104]  & ~new_n658_;
  assign \grant[104]  = ~new_n10181_ & new_n10182_;
  assign new_n10184_ = new_n667_ & ~new_n1002_;
  assign new_n10185_ = new_n672_ & ~new_n10184_;
  assign new_n10186_ = new_n676_ & ~new_n10185_;
  assign new_n10187_ = new_n680_ & ~new_n10186_;
  assign new_n10188_ = new_n684_ & ~new_n10187_;
  assign new_n10189_ = new_n688_ & ~new_n10188_;
  assign new_n10190_ = new_n692_ & ~new_n10189_;
  assign new_n10191_ = new_n696_ & ~new_n10190_;
  assign new_n10192_ = new_n700_ & ~new_n10191_;
  assign new_n10193_ = new_n704_ & ~new_n10192_;
  assign new_n10194_ = new_n708_ & ~new_n10193_;
  assign new_n10195_ = new_n712_ & ~new_n10194_;
  assign new_n10196_ = new_n716_ & ~new_n10195_;
  assign new_n10197_ = new_n720_ & ~new_n10196_;
  assign new_n10198_ = new_n1484_ & ~new_n10197_;
  assign new_n10199_ = new_n1486_ & ~new_n10198_;
  assign new_n10200_ = new_n1750_ & ~new_n10199_;
  assign new_n10201_ = new_n731_ & ~new_n10200_;
  assign new_n10202_ = new_n735_ & ~new_n10201_;
  assign new_n10203_ = new_n739_ & ~new_n10202_;
  assign new_n10204_ = new_n743_ & ~new_n10203_;
  assign new_n10205_ = new_n747_ & ~new_n10204_;
  assign new_n10206_ = new_n751_ & ~new_n10205_;
  assign new_n10207_ = new_n755_ & ~new_n10206_;
  assign new_n10208_ = new_n759_ & ~new_n10207_;
  assign new_n10209_ = new_n763_ & ~new_n10208_;
  assign new_n10210_ = new_n767_ & ~new_n10209_;
  assign new_n10211_ = new_n771_ & ~new_n10210_;
  assign new_n10212_ = new_n775_ & ~new_n10211_;
  assign new_n10213_ = new_n779_ & ~new_n10212_;
  assign new_n10214_ = new_n783_ & ~new_n10213_;
  assign new_n10215_ = new_n787_ & ~new_n10214_;
  assign new_n10216_ = new_n791_ & ~new_n10215_;
  assign new_n10217_ = new_n795_ & ~new_n10216_;
  assign new_n10218_ = new_n799_ & ~new_n10217_;
  assign new_n10219_ = new_n803_ & ~new_n10218_;
  assign new_n10220_ = new_n807_ & ~new_n10219_;
  assign new_n10221_ = new_n811_ & ~new_n10220_;
  assign new_n10222_ = new_n815_ & ~new_n10221_;
  assign new_n10223_ = new_n819_ & ~new_n10222_;
  assign new_n10224_ = new_n823_ & ~new_n10223_;
  assign new_n10225_ = new_n827_ & ~new_n10224_;
  assign new_n10226_ = new_n831_ & ~new_n10225_;
  assign new_n10227_ = new_n835_ & ~new_n10226_;
  assign new_n10228_ = new_n839_ & ~new_n10227_;
  assign new_n10229_ = new_n843_ & ~new_n10228_;
  assign new_n10230_ = new_n847_ & ~new_n10229_;
  assign new_n10231_ = new_n851_ & ~new_n10230_;
  assign new_n10232_ = new_n855_ & ~new_n10231_;
  assign new_n10233_ = new_n859_ & ~new_n10232_;
  assign new_n10234_ = new_n863_ & ~new_n10233_;
  assign new_n10235_ = new_n867_ & ~new_n10234_;
  assign new_n10236_ = new_n871_ & ~new_n10235_;
  assign new_n10237_ = new_n875_ & ~new_n10236_;
  assign new_n10238_ = new_n879_ & ~new_n10237_;
  assign new_n10239_ = new_n883_ & ~new_n10238_;
  assign new_n10240_ = new_n887_ & ~new_n10239_;
  assign new_n10241_ = new_n891_ & ~new_n10240_;
  assign new_n10242_ = new_n895_ & ~new_n10241_;
  assign new_n10243_ = new_n899_ & ~new_n10242_;
  assign new_n10244_ = new_n903_ & ~new_n10243_;
  assign new_n10245_ = new_n907_ & ~new_n10244_;
  assign new_n10246_ = new_n911_ & ~new_n10245_;
  assign new_n10247_ = new_n915_ & ~new_n10246_;
  assign new_n10248_ = new_n919_ & ~new_n10247_;
  assign new_n10249_ = new_n923_ & ~new_n10248_;
  assign new_n10250_ = new_n927_ & ~new_n10249_;
  assign new_n10251_ = new_n931_ & ~new_n10250_;
  assign new_n10252_ = new_n935_ & ~new_n10251_;
  assign new_n10253_ = new_n939_ & ~new_n10252_;
  assign new_n10254_ = new_n943_ & ~new_n10253_;
  assign new_n10255_ = new_n947_ & ~new_n10254_;
  assign new_n10256_ = new_n951_ & ~new_n10255_;
  assign new_n10257_ = new_n955_ & ~new_n10256_;
  assign new_n10258_ = new_n959_ & ~new_n10257_;
  assign new_n10259_ = new_n963_ & ~new_n10258_;
  assign new_n10260_ = new_n967_ & ~new_n10259_;
  assign new_n10261_ = new_n971_ & ~new_n10260_;
  assign new_n10262_ = new_n975_ & ~new_n10261_;
  assign new_n10263_ = new_n979_ & ~new_n10262_;
  assign new_n10264_ = new_n983_ & ~new_n10263_;
  assign new_n10265_ = new_n987_ & ~new_n10264_;
  assign new_n10266_ = new_n991_ & ~new_n10265_;
  assign new_n10267_ = new_n995_ & ~new_n10266_;
  assign new_n10268_ = \req[105]  & ~new_n997_;
  assign \grant[105]  = ~new_n10267_ & new_n10268_;
  assign new_n10270_ = new_n1006_ & ~new_n1339_;
  assign new_n10271_ = new_n1011_ & ~new_n10270_;
  assign new_n10272_ = new_n1015_ & ~new_n10271_;
  assign new_n10273_ = new_n1019_ & ~new_n10272_;
  assign new_n10274_ = new_n1023_ & ~new_n10273_;
  assign new_n10275_ = new_n1027_ & ~new_n10274_;
  assign new_n10276_ = new_n1031_ & ~new_n10275_;
  assign new_n10277_ = new_n1035_ & ~new_n10276_;
  assign new_n10278_ = new_n1039_ & ~new_n10277_;
  assign new_n10279_ = new_n1043_ & ~new_n10278_;
  assign new_n10280_ = new_n1047_ & ~new_n10279_;
  assign new_n10281_ = new_n1051_ & ~new_n10280_;
  assign new_n10282_ = new_n1055_ & ~new_n10281_;
  assign new_n10283_ = new_n1059_ & ~new_n10282_;
  assign new_n10284_ = new_n1574_ & ~new_n10283_;
  assign new_n10285_ = new_n1576_ & ~new_n10284_;
  assign new_n10286_ = new_n1837_ & ~new_n10285_;
  assign new_n10287_ = new_n1068_ & ~new_n10286_;
  assign new_n10288_ = new_n1072_ & ~new_n10287_;
  assign new_n10289_ = new_n1076_ & ~new_n10288_;
  assign new_n10290_ = new_n1080_ & ~new_n10289_;
  assign new_n10291_ = new_n1084_ & ~new_n10290_;
  assign new_n10292_ = new_n1088_ & ~new_n10291_;
  assign new_n10293_ = new_n1092_ & ~new_n10292_;
  assign new_n10294_ = new_n1096_ & ~new_n10293_;
  assign new_n10295_ = new_n1100_ & ~new_n10294_;
  assign new_n10296_ = new_n1104_ & ~new_n10295_;
  assign new_n10297_ = new_n1108_ & ~new_n10296_;
  assign new_n10298_ = new_n1112_ & ~new_n10297_;
  assign new_n10299_ = new_n1116_ & ~new_n10298_;
  assign new_n10300_ = new_n1120_ & ~new_n10299_;
  assign new_n10301_ = new_n1124_ & ~new_n10300_;
  assign new_n10302_ = new_n1128_ & ~new_n10301_;
  assign new_n10303_ = new_n1132_ & ~new_n10302_;
  assign new_n10304_ = new_n1136_ & ~new_n10303_;
  assign new_n10305_ = new_n1140_ & ~new_n10304_;
  assign new_n10306_ = new_n1144_ & ~new_n10305_;
  assign new_n10307_ = new_n1148_ & ~new_n10306_;
  assign new_n10308_ = new_n1152_ & ~new_n10307_;
  assign new_n10309_ = new_n1156_ & ~new_n10308_;
  assign new_n10310_ = new_n1160_ & ~new_n10309_;
  assign new_n10311_ = new_n1164_ & ~new_n10310_;
  assign new_n10312_ = new_n1168_ & ~new_n10311_;
  assign new_n10313_ = new_n1172_ & ~new_n10312_;
  assign new_n10314_ = new_n1176_ & ~new_n10313_;
  assign new_n10315_ = new_n1180_ & ~new_n10314_;
  assign new_n10316_ = new_n1184_ & ~new_n10315_;
  assign new_n10317_ = new_n1188_ & ~new_n10316_;
  assign new_n10318_ = new_n1192_ & ~new_n10317_;
  assign new_n10319_ = new_n1196_ & ~new_n10318_;
  assign new_n10320_ = new_n1200_ & ~new_n10319_;
  assign new_n10321_ = new_n1204_ & ~new_n10320_;
  assign new_n10322_ = new_n1208_ & ~new_n10321_;
  assign new_n10323_ = new_n1212_ & ~new_n10322_;
  assign new_n10324_ = new_n1216_ & ~new_n10323_;
  assign new_n10325_ = new_n1220_ & ~new_n10324_;
  assign new_n10326_ = new_n1224_ & ~new_n10325_;
  assign new_n10327_ = new_n1228_ & ~new_n10326_;
  assign new_n10328_ = new_n1232_ & ~new_n10327_;
  assign new_n10329_ = new_n1236_ & ~new_n10328_;
  assign new_n10330_ = new_n1240_ & ~new_n10329_;
  assign new_n10331_ = new_n1244_ & ~new_n10330_;
  assign new_n10332_ = new_n1248_ & ~new_n10331_;
  assign new_n10333_ = new_n1252_ & ~new_n10332_;
  assign new_n10334_ = new_n1256_ & ~new_n10333_;
  assign new_n10335_ = new_n1260_ & ~new_n10334_;
  assign new_n10336_ = new_n1264_ & ~new_n10335_;
  assign new_n10337_ = new_n1268_ & ~new_n10336_;
  assign new_n10338_ = new_n1272_ & ~new_n10337_;
  assign new_n10339_ = new_n1276_ & ~new_n10338_;
  assign new_n10340_ = new_n1280_ & ~new_n10339_;
  assign new_n10341_ = new_n1284_ & ~new_n10340_;
  assign new_n10342_ = new_n1288_ & ~new_n10341_;
  assign new_n10343_ = new_n1292_ & ~new_n10342_;
  assign new_n10344_ = new_n1296_ & ~new_n10343_;
  assign new_n10345_ = new_n1300_ & ~new_n10344_;
  assign new_n10346_ = new_n1304_ & ~new_n10345_;
  assign new_n10347_ = new_n1308_ & ~new_n10346_;
  assign new_n10348_ = new_n1312_ & ~new_n10347_;
  assign new_n10349_ = new_n1316_ & ~new_n10348_;
  assign new_n10350_ = new_n1320_ & ~new_n10349_;
  assign new_n10351_ = new_n1324_ & ~new_n10350_;
  assign new_n10352_ = new_n1328_ & ~new_n10351_;
  assign new_n10353_ = new_n1332_ & ~new_n10352_;
  assign new_n10354_ = \req[106]  & ~new_n1334_;
  assign \grant[106]  = ~new_n10353_ & new_n10354_;
  assign new_n10356_ = ~new_n671_ & new_n1343_;
  assign new_n10357_ = new_n1348_ & ~new_n10356_;
  assign new_n10358_ = new_n1352_ & ~new_n10357_;
  assign new_n10359_ = new_n1356_ & ~new_n10358_;
  assign new_n10360_ = new_n1360_ & ~new_n10359_;
  assign new_n10361_ = new_n1364_ & ~new_n10360_;
  assign new_n10362_ = new_n1368_ & ~new_n10361_;
  assign new_n10363_ = new_n1372_ & ~new_n10362_;
  assign new_n10364_ = new_n1376_ & ~new_n10363_;
  assign new_n10365_ = new_n1380_ & ~new_n10364_;
  assign new_n10366_ = new_n1384_ & ~new_n10365_;
  assign new_n10367_ = new_n1388_ & ~new_n10366_;
  assign new_n10368_ = new_n1392_ & ~new_n10367_;
  assign new_n10369_ = new_n1396_ & ~new_n10368_;
  assign new_n10370_ = new_n1663_ & ~new_n10369_;
  assign new_n10371_ = new_n392_ & ~new_n10370_;
  assign new_n10372_ = new_n396_ & ~new_n10371_;
  assign new_n10373_ = new_n400_ & ~new_n10372_;
  assign new_n10374_ = new_n404_ & ~new_n10373_;
  assign new_n10375_ = new_n408_ & ~new_n10374_;
  assign new_n10376_ = new_n412_ & ~new_n10375_;
  assign new_n10377_ = new_n416_ & ~new_n10376_;
  assign new_n10378_ = new_n420_ & ~new_n10377_;
  assign new_n10379_ = new_n424_ & ~new_n10378_;
  assign new_n10380_ = new_n428_ & ~new_n10379_;
  assign new_n10381_ = new_n432_ & ~new_n10380_;
  assign new_n10382_ = new_n436_ & ~new_n10381_;
  assign new_n10383_ = new_n440_ & ~new_n10382_;
  assign new_n10384_ = new_n444_ & ~new_n10383_;
  assign new_n10385_ = new_n448_ & ~new_n10384_;
  assign new_n10386_ = new_n452_ & ~new_n10385_;
  assign new_n10387_ = new_n456_ & ~new_n10386_;
  assign new_n10388_ = new_n460_ & ~new_n10387_;
  assign new_n10389_ = new_n464_ & ~new_n10388_;
  assign new_n10390_ = new_n468_ & ~new_n10389_;
  assign new_n10391_ = new_n472_ & ~new_n10390_;
  assign new_n10392_ = new_n476_ & ~new_n10391_;
  assign new_n10393_ = new_n480_ & ~new_n10392_;
  assign new_n10394_ = new_n484_ & ~new_n10393_;
  assign new_n10395_ = new_n488_ & ~new_n10394_;
  assign new_n10396_ = new_n492_ & ~new_n10395_;
  assign new_n10397_ = new_n496_ & ~new_n10396_;
  assign new_n10398_ = new_n500_ & ~new_n10397_;
  assign new_n10399_ = new_n504_ & ~new_n10398_;
  assign new_n10400_ = new_n508_ & ~new_n10399_;
  assign new_n10401_ = new_n512_ & ~new_n10400_;
  assign new_n10402_ = new_n516_ & ~new_n10401_;
  assign new_n10403_ = new_n520_ & ~new_n10402_;
  assign new_n10404_ = new_n524_ & ~new_n10403_;
  assign new_n10405_ = new_n528_ & ~new_n10404_;
  assign new_n10406_ = new_n532_ & ~new_n10405_;
  assign new_n10407_ = new_n536_ & ~new_n10406_;
  assign new_n10408_ = new_n540_ & ~new_n10407_;
  assign new_n10409_ = new_n544_ & ~new_n10408_;
  assign new_n10410_ = new_n548_ & ~new_n10409_;
  assign new_n10411_ = new_n552_ & ~new_n10410_;
  assign new_n10412_ = new_n556_ & ~new_n10411_;
  assign new_n10413_ = new_n560_ & ~new_n10412_;
  assign new_n10414_ = new_n564_ & ~new_n10413_;
  assign new_n10415_ = new_n568_ & ~new_n10414_;
  assign new_n10416_ = new_n572_ & ~new_n10415_;
  assign new_n10417_ = new_n576_ & ~new_n10416_;
  assign new_n10418_ = new_n580_ & ~new_n10417_;
  assign new_n10419_ = new_n584_ & ~new_n10418_;
  assign new_n10420_ = new_n588_ & ~new_n10419_;
  assign new_n10421_ = new_n592_ & ~new_n10420_;
  assign new_n10422_ = new_n596_ & ~new_n10421_;
  assign new_n10423_ = new_n600_ & ~new_n10422_;
  assign new_n10424_ = new_n604_ & ~new_n10423_;
  assign new_n10425_ = new_n608_ & ~new_n10424_;
  assign new_n10426_ = new_n612_ & ~new_n10425_;
  assign new_n10427_ = new_n616_ & ~new_n10426_;
  assign new_n10428_ = new_n620_ & ~new_n10427_;
  assign new_n10429_ = new_n624_ & ~new_n10428_;
  assign new_n10430_ = new_n628_ & ~new_n10429_;
  assign new_n10431_ = new_n632_ & ~new_n10430_;
  assign new_n10432_ = new_n636_ & ~new_n10431_;
  assign new_n10433_ = new_n640_ & ~new_n10432_;
  assign new_n10434_ = new_n644_ & ~new_n10433_;
  assign new_n10435_ = new_n648_ & ~new_n10434_;
  assign new_n10436_ = new_n652_ & ~new_n10435_;
  assign new_n10437_ = new_n656_ & ~new_n10436_;
  assign new_n10438_ = new_n660_ & ~new_n10437_;
  assign new_n10439_ = new_n664_ & ~new_n10438_;
  assign new_n10440_ = \req[107]  & ~new_n666_;
  assign \grant[107]  = ~new_n10439_ & new_n10440_;
  assign new_n10442_ = new_n675_ & ~new_n1010_;
  assign new_n10443_ = new_n680_ & ~new_n10442_;
  assign new_n10444_ = new_n684_ & ~new_n10443_;
  assign new_n10445_ = new_n688_ & ~new_n10444_;
  assign new_n10446_ = new_n692_ & ~new_n10445_;
  assign new_n10447_ = new_n696_ & ~new_n10446_;
  assign new_n10448_ = new_n700_ & ~new_n10447_;
  assign new_n10449_ = new_n704_ & ~new_n10448_;
  assign new_n10450_ = new_n708_ & ~new_n10449_;
  assign new_n10451_ = new_n712_ & ~new_n10450_;
  assign new_n10452_ = new_n716_ & ~new_n10451_;
  assign new_n10453_ = new_n720_ & ~new_n10452_;
  assign new_n10454_ = new_n1484_ & ~new_n10453_;
  assign new_n10455_ = new_n1486_ & ~new_n10454_;
  assign new_n10456_ = new_n1750_ & ~new_n10455_;
  assign new_n10457_ = new_n731_ & ~new_n10456_;
  assign new_n10458_ = new_n735_ & ~new_n10457_;
  assign new_n10459_ = new_n739_ & ~new_n10458_;
  assign new_n10460_ = new_n743_ & ~new_n10459_;
  assign new_n10461_ = new_n747_ & ~new_n10460_;
  assign new_n10462_ = new_n751_ & ~new_n10461_;
  assign new_n10463_ = new_n755_ & ~new_n10462_;
  assign new_n10464_ = new_n759_ & ~new_n10463_;
  assign new_n10465_ = new_n763_ & ~new_n10464_;
  assign new_n10466_ = new_n767_ & ~new_n10465_;
  assign new_n10467_ = new_n771_ & ~new_n10466_;
  assign new_n10468_ = new_n775_ & ~new_n10467_;
  assign new_n10469_ = new_n779_ & ~new_n10468_;
  assign new_n10470_ = new_n783_ & ~new_n10469_;
  assign new_n10471_ = new_n787_ & ~new_n10470_;
  assign new_n10472_ = new_n791_ & ~new_n10471_;
  assign new_n10473_ = new_n795_ & ~new_n10472_;
  assign new_n10474_ = new_n799_ & ~new_n10473_;
  assign new_n10475_ = new_n803_ & ~new_n10474_;
  assign new_n10476_ = new_n807_ & ~new_n10475_;
  assign new_n10477_ = new_n811_ & ~new_n10476_;
  assign new_n10478_ = new_n815_ & ~new_n10477_;
  assign new_n10479_ = new_n819_ & ~new_n10478_;
  assign new_n10480_ = new_n823_ & ~new_n10479_;
  assign new_n10481_ = new_n827_ & ~new_n10480_;
  assign new_n10482_ = new_n831_ & ~new_n10481_;
  assign new_n10483_ = new_n835_ & ~new_n10482_;
  assign new_n10484_ = new_n839_ & ~new_n10483_;
  assign new_n10485_ = new_n843_ & ~new_n10484_;
  assign new_n10486_ = new_n847_ & ~new_n10485_;
  assign new_n10487_ = new_n851_ & ~new_n10486_;
  assign new_n10488_ = new_n855_ & ~new_n10487_;
  assign new_n10489_ = new_n859_ & ~new_n10488_;
  assign new_n10490_ = new_n863_ & ~new_n10489_;
  assign new_n10491_ = new_n867_ & ~new_n10490_;
  assign new_n10492_ = new_n871_ & ~new_n10491_;
  assign new_n10493_ = new_n875_ & ~new_n10492_;
  assign new_n10494_ = new_n879_ & ~new_n10493_;
  assign new_n10495_ = new_n883_ & ~new_n10494_;
  assign new_n10496_ = new_n887_ & ~new_n10495_;
  assign new_n10497_ = new_n891_ & ~new_n10496_;
  assign new_n10498_ = new_n895_ & ~new_n10497_;
  assign new_n10499_ = new_n899_ & ~new_n10498_;
  assign new_n10500_ = new_n903_ & ~new_n10499_;
  assign new_n10501_ = new_n907_ & ~new_n10500_;
  assign new_n10502_ = new_n911_ & ~new_n10501_;
  assign new_n10503_ = new_n915_ & ~new_n10502_;
  assign new_n10504_ = new_n919_ & ~new_n10503_;
  assign new_n10505_ = new_n923_ & ~new_n10504_;
  assign new_n10506_ = new_n927_ & ~new_n10505_;
  assign new_n10507_ = new_n931_ & ~new_n10506_;
  assign new_n10508_ = new_n935_ & ~new_n10507_;
  assign new_n10509_ = new_n939_ & ~new_n10508_;
  assign new_n10510_ = new_n943_ & ~new_n10509_;
  assign new_n10511_ = new_n947_ & ~new_n10510_;
  assign new_n10512_ = new_n951_ & ~new_n10511_;
  assign new_n10513_ = new_n955_ & ~new_n10512_;
  assign new_n10514_ = new_n959_ & ~new_n10513_;
  assign new_n10515_ = new_n963_ & ~new_n10514_;
  assign new_n10516_ = new_n967_ & ~new_n10515_;
  assign new_n10517_ = new_n971_ & ~new_n10516_;
  assign new_n10518_ = new_n975_ & ~new_n10517_;
  assign new_n10519_ = new_n979_ & ~new_n10518_;
  assign new_n10520_ = new_n983_ & ~new_n10519_;
  assign new_n10521_ = new_n987_ & ~new_n10520_;
  assign new_n10522_ = new_n991_ & ~new_n10521_;
  assign new_n10523_ = new_n995_ & ~new_n10522_;
  assign new_n10524_ = new_n999_ & ~new_n10523_;
  assign new_n10525_ = new_n1003_ & ~new_n10524_;
  assign new_n10526_ = \req[108]  & ~new_n1005_;
  assign \grant[108]  = ~new_n10525_ & new_n10526_;
  assign new_n10528_ = new_n1014_ & ~new_n1347_;
  assign new_n10529_ = new_n1019_ & ~new_n10528_;
  assign new_n10530_ = new_n1023_ & ~new_n10529_;
  assign new_n10531_ = new_n1027_ & ~new_n10530_;
  assign new_n10532_ = new_n1031_ & ~new_n10531_;
  assign new_n10533_ = new_n1035_ & ~new_n10532_;
  assign new_n10534_ = new_n1039_ & ~new_n10533_;
  assign new_n10535_ = new_n1043_ & ~new_n10534_;
  assign new_n10536_ = new_n1047_ & ~new_n10535_;
  assign new_n10537_ = new_n1051_ & ~new_n10536_;
  assign new_n10538_ = new_n1055_ & ~new_n10537_;
  assign new_n10539_ = new_n1059_ & ~new_n10538_;
  assign new_n10540_ = new_n1574_ & ~new_n10539_;
  assign new_n10541_ = new_n1576_ & ~new_n10540_;
  assign new_n10542_ = new_n1837_ & ~new_n10541_;
  assign new_n10543_ = new_n1068_ & ~new_n10542_;
  assign new_n10544_ = new_n1072_ & ~new_n10543_;
  assign new_n10545_ = new_n1076_ & ~new_n10544_;
  assign new_n10546_ = new_n1080_ & ~new_n10545_;
  assign new_n10547_ = new_n1084_ & ~new_n10546_;
  assign new_n10548_ = new_n1088_ & ~new_n10547_;
  assign new_n10549_ = new_n1092_ & ~new_n10548_;
  assign new_n10550_ = new_n1096_ & ~new_n10549_;
  assign new_n10551_ = new_n1100_ & ~new_n10550_;
  assign new_n10552_ = new_n1104_ & ~new_n10551_;
  assign new_n10553_ = new_n1108_ & ~new_n10552_;
  assign new_n10554_ = new_n1112_ & ~new_n10553_;
  assign new_n10555_ = new_n1116_ & ~new_n10554_;
  assign new_n10556_ = new_n1120_ & ~new_n10555_;
  assign new_n10557_ = new_n1124_ & ~new_n10556_;
  assign new_n10558_ = new_n1128_ & ~new_n10557_;
  assign new_n10559_ = new_n1132_ & ~new_n10558_;
  assign new_n10560_ = new_n1136_ & ~new_n10559_;
  assign new_n10561_ = new_n1140_ & ~new_n10560_;
  assign new_n10562_ = new_n1144_ & ~new_n10561_;
  assign new_n10563_ = new_n1148_ & ~new_n10562_;
  assign new_n10564_ = new_n1152_ & ~new_n10563_;
  assign new_n10565_ = new_n1156_ & ~new_n10564_;
  assign new_n10566_ = new_n1160_ & ~new_n10565_;
  assign new_n10567_ = new_n1164_ & ~new_n10566_;
  assign new_n10568_ = new_n1168_ & ~new_n10567_;
  assign new_n10569_ = new_n1172_ & ~new_n10568_;
  assign new_n10570_ = new_n1176_ & ~new_n10569_;
  assign new_n10571_ = new_n1180_ & ~new_n10570_;
  assign new_n10572_ = new_n1184_ & ~new_n10571_;
  assign new_n10573_ = new_n1188_ & ~new_n10572_;
  assign new_n10574_ = new_n1192_ & ~new_n10573_;
  assign new_n10575_ = new_n1196_ & ~new_n10574_;
  assign new_n10576_ = new_n1200_ & ~new_n10575_;
  assign new_n10577_ = new_n1204_ & ~new_n10576_;
  assign new_n10578_ = new_n1208_ & ~new_n10577_;
  assign new_n10579_ = new_n1212_ & ~new_n10578_;
  assign new_n10580_ = new_n1216_ & ~new_n10579_;
  assign new_n10581_ = new_n1220_ & ~new_n10580_;
  assign new_n10582_ = new_n1224_ & ~new_n10581_;
  assign new_n10583_ = new_n1228_ & ~new_n10582_;
  assign new_n10584_ = new_n1232_ & ~new_n10583_;
  assign new_n10585_ = new_n1236_ & ~new_n10584_;
  assign new_n10586_ = new_n1240_ & ~new_n10585_;
  assign new_n10587_ = new_n1244_ & ~new_n10586_;
  assign new_n10588_ = new_n1248_ & ~new_n10587_;
  assign new_n10589_ = new_n1252_ & ~new_n10588_;
  assign new_n10590_ = new_n1256_ & ~new_n10589_;
  assign new_n10591_ = new_n1260_ & ~new_n10590_;
  assign new_n10592_ = new_n1264_ & ~new_n10591_;
  assign new_n10593_ = new_n1268_ & ~new_n10592_;
  assign new_n10594_ = new_n1272_ & ~new_n10593_;
  assign new_n10595_ = new_n1276_ & ~new_n10594_;
  assign new_n10596_ = new_n1280_ & ~new_n10595_;
  assign new_n10597_ = new_n1284_ & ~new_n10596_;
  assign new_n10598_ = new_n1288_ & ~new_n10597_;
  assign new_n10599_ = new_n1292_ & ~new_n10598_;
  assign new_n10600_ = new_n1296_ & ~new_n10599_;
  assign new_n10601_ = new_n1300_ & ~new_n10600_;
  assign new_n10602_ = new_n1304_ & ~new_n10601_;
  assign new_n10603_ = new_n1308_ & ~new_n10602_;
  assign new_n10604_ = new_n1312_ & ~new_n10603_;
  assign new_n10605_ = new_n1316_ & ~new_n10604_;
  assign new_n10606_ = new_n1320_ & ~new_n10605_;
  assign new_n10607_ = new_n1324_ & ~new_n10606_;
  assign new_n10608_ = new_n1328_ & ~new_n10607_;
  assign new_n10609_ = new_n1332_ & ~new_n10608_;
  assign new_n10610_ = new_n1336_ & ~new_n10609_;
  assign new_n10611_ = new_n1340_ & ~new_n10610_;
  assign new_n10612_ = \req[109]  & ~new_n1342_;
  assign \grant[109]  = ~new_n10611_ & new_n10612_;
  assign new_n10614_ = ~new_n679_ & new_n1351_;
  assign new_n10615_ = new_n1356_ & ~new_n10614_;
  assign new_n10616_ = new_n1360_ & ~new_n10615_;
  assign new_n10617_ = new_n1364_ & ~new_n10616_;
  assign new_n10618_ = new_n1368_ & ~new_n10617_;
  assign new_n10619_ = new_n1372_ & ~new_n10618_;
  assign new_n10620_ = new_n1376_ & ~new_n10619_;
  assign new_n10621_ = new_n1380_ & ~new_n10620_;
  assign new_n10622_ = new_n1384_ & ~new_n10621_;
  assign new_n10623_ = new_n1388_ & ~new_n10622_;
  assign new_n10624_ = new_n1392_ & ~new_n10623_;
  assign new_n10625_ = new_n1396_ & ~new_n10624_;
  assign new_n10626_ = new_n1663_ & ~new_n10625_;
  assign new_n10627_ = new_n392_ & ~new_n10626_;
  assign new_n10628_ = new_n396_ & ~new_n10627_;
  assign new_n10629_ = new_n400_ & ~new_n10628_;
  assign new_n10630_ = new_n404_ & ~new_n10629_;
  assign new_n10631_ = new_n408_ & ~new_n10630_;
  assign new_n10632_ = new_n412_ & ~new_n10631_;
  assign new_n10633_ = new_n416_ & ~new_n10632_;
  assign new_n10634_ = new_n420_ & ~new_n10633_;
  assign new_n10635_ = new_n424_ & ~new_n10634_;
  assign new_n10636_ = new_n428_ & ~new_n10635_;
  assign new_n10637_ = new_n432_ & ~new_n10636_;
  assign new_n10638_ = new_n436_ & ~new_n10637_;
  assign new_n10639_ = new_n440_ & ~new_n10638_;
  assign new_n10640_ = new_n444_ & ~new_n10639_;
  assign new_n10641_ = new_n448_ & ~new_n10640_;
  assign new_n10642_ = new_n452_ & ~new_n10641_;
  assign new_n10643_ = new_n456_ & ~new_n10642_;
  assign new_n10644_ = new_n460_ & ~new_n10643_;
  assign new_n10645_ = new_n464_ & ~new_n10644_;
  assign new_n10646_ = new_n468_ & ~new_n10645_;
  assign new_n10647_ = new_n472_ & ~new_n10646_;
  assign new_n10648_ = new_n476_ & ~new_n10647_;
  assign new_n10649_ = new_n480_ & ~new_n10648_;
  assign new_n10650_ = new_n484_ & ~new_n10649_;
  assign new_n10651_ = new_n488_ & ~new_n10650_;
  assign new_n10652_ = new_n492_ & ~new_n10651_;
  assign new_n10653_ = new_n496_ & ~new_n10652_;
  assign new_n10654_ = new_n500_ & ~new_n10653_;
  assign new_n10655_ = new_n504_ & ~new_n10654_;
  assign new_n10656_ = new_n508_ & ~new_n10655_;
  assign new_n10657_ = new_n512_ & ~new_n10656_;
  assign new_n10658_ = new_n516_ & ~new_n10657_;
  assign new_n10659_ = new_n520_ & ~new_n10658_;
  assign new_n10660_ = new_n524_ & ~new_n10659_;
  assign new_n10661_ = new_n528_ & ~new_n10660_;
  assign new_n10662_ = new_n532_ & ~new_n10661_;
  assign new_n10663_ = new_n536_ & ~new_n10662_;
  assign new_n10664_ = new_n540_ & ~new_n10663_;
  assign new_n10665_ = new_n544_ & ~new_n10664_;
  assign new_n10666_ = new_n548_ & ~new_n10665_;
  assign new_n10667_ = new_n552_ & ~new_n10666_;
  assign new_n10668_ = new_n556_ & ~new_n10667_;
  assign new_n10669_ = new_n560_ & ~new_n10668_;
  assign new_n10670_ = new_n564_ & ~new_n10669_;
  assign new_n10671_ = new_n568_ & ~new_n10670_;
  assign new_n10672_ = new_n572_ & ~new_n10671_;
  assign new_n10673_ = new_n576_ & ~new_n10672_;
  assign new_n10674_ = new_n580_ & ~new_n10673_;
  assign new_n10675_ = new_n584_ & ~new_n10674_;
  assign new_n10676_ = new_n588_ & ~new_n10675_;
  assign new_n10677_ = new_n592_ & ~new_n10676_;
  assign new_n10678_ = new_n596_ & ~new_n10677_;
  assign new_n10679_ = new_n600_ & ~new_n10678_;
  assign new_n10680_ = new_n604_ & ~new_n10679_;
  assign new_n10681_ = new_n608_ & ~new_n10680_;
  assign new_n10682_ = new_n612_ & ~new_n10681_;
  assign new_n10683_ = new_n616_ & ~new_n10682_;
  assign new_n10684_ = new_n620_ & ~new_n10683_;
  assign new_n10685_ = new_n624_ & ~new_n10684_;
  assign new_n10686_ = new_n628_ & ~new_n10685_;
  assign new_n10687_ = new_n632_ & ~new_n10686_;
  assign new_n10688_ = new_n636_ & ~new_n10687_;
  assign new_n10689_ = new_n640_ & ~new_n10688_;
  assign new_n10690_ = new_n644_ & ~new_n10689_;
  assign new_n10691_ = new_n648_ & ~new_n10690_;
  assign new_n10692_ = new_n652_ & ~new_n10691_;
  assign new_n10693_ = new_n656_ & ~new_n10692_;
  assign new_n10694_ = new_n660_ & ~new_n10693_;
  assign new_n10695_ = new_n664_ & ~new_n10694_;
  assign new_n10696_ = new_n668_ & ~new_n10695_;
  assign new_n10697_ = new_n672_ & ~new_n10696_;
  assign new_n10698_ = \req[110]  & ~new_n674_;
  assign \grant[110]  = ~new_n10697_ & new_n10698_;
  assign new_n10700_ = new_n683_ & ~new_n1018_;
  assign new_n10701_ = new_n688_ & ~new_n10700_;
  assign new_n10702_ = new_n692_ & ~new_n10701_;
  assign new_n10703_ = new_n696_ & ~new_n10702_;
  assign new_n10704_ = new_n700_ & ~new_n10703_;
  assign new_n10705_ = new_n704_ & ~new_n10704_;
  assign new_n10706_ = new_n708_ & ~new_n10705_;
  assign new_n10707_ = new_n712_ & ~new_n10706_;
  assign new_n10708_ = new_n716_ & ~new_n10707_;
  assign new_n10709_ = new_n720_ & ~new_n10708_;
  assign new_n10710_ = new_n1484_ & ~new_n10709_;
  assign new_n10711_ = new_n1486_ & ~new_n10710_;
  assign new_n10712_ = new_n1750_ & ~new_n10711_;
  assign new_n10713_ = new_n731_ & ~new_n10712_;
  assign new_n10714_ = new_n735_ & ~new_n10713_;
  assign new_n10715_ = new_n739_ & ~new_n10714_;
  assign new_n10716_ = new_n743_ & ~new_n10715_;
  assign new_n10717_ = new_n747_ & ~new_n10716_;
  assign new_n10718_ = new_n751_ & ~new_n10717_;
  assign new_n10719_ = new_n755_ & ~new_n10718_;
  assign new_n10720_ = new_n759_ & ~new_n10719_;
  assign new_n10721_ = new_n763_ & ~new_n10720_;
  assign new_n10722_ = new_n767_ & ~new_n10721_;
  assign new_n10723_ = new_n771_ & ~new_n10722_;
  assign new_n10724_ = new_n775_ & ~new_n10723_;
  assign new_n10725_ = new_n779_ & ~new_n10724_;
  assign new_n10726_ = new_n783_ & ~new_n10725_;
  assign new_n10727_ = new_n787_ & ~new_n10726_;
  assign new_n10728_ = new_n791_ & ~new_n10727_;
  assign new_n10729_ = new_n795_ & ~new_n10728_;
  assign new_n10730_ = new_n799_ & ~new_n10729_;
  assign new_n10731_ = new_n803_ & ~new_n10730_;
  assign new_n10732_ = new_n807_ & ~new_n10731_;
  assign new_n10733_ = new_n811_ & ~new_n10732_;
  assign new_n10734_ = new_n815_ & ~new_n10733_;
  assign new_n10735_ = new_n819_ & ~new_n10734_;
  assign new_n10736_ = new_n823_ & ~new_n10735_;
  assign new_n10737_ = new_n827_ & ~new_n10736_;
  assign new_n10738_ = new_n831_ & ~new_n10737_;
  assign new_n10739_ = new_n835_ & ~new_n10738_;
  assign new_n10740_ = new_n839_ & ~new_n10739_;
  assign new_n10741_ = new_n843_ & ~new_n10740_;
  assign new_n10742_ = new_n847_ & ~new_n10741_;
  assign new_n10743_ = new_n851_ & ~new_n10742_;
  assign new_n10744_ = new_n855_ & ~new_n10743_;
  assign new_n10745_ = new_n859_ & ~new_n10744_;
  assign new_n10746_ = new_n863_ & ~new_n10745_;
  assign new_n10747_ = new_n867_ & ~new_n10746_;
  assign new_n10748_ = new_n871_ & ~new_n10747_;
  assign new_n10749_ = new_n875_ & ~new_n10748_;
  assign new_n10750_ = new_n879_ & ~new_n10749_;
  assign new_n10751_ = new_n883_ & ~new_n10750_;
  assign new_n10752_ = new_n887_ & ~new_n10751_;
  assign new_n10753_ = new_n891_ & ~new_n10752_;
  assign new_n10754_ = new_n895_ & ~new_n10753_;
  assign new_n10755_ = new_n899_ & ~new_n10754_;
  assign new_n10756_ = new_n903_ & ~new_n10755_;
  assign new_n10757_ = new_n907_ & ~new_n10756_;
  assign new_n10758_ = new_n911_ & ~new_n10757_;
  assign new_n10759_ = new_n915_ & ~new_n10758_;
  assign new_n10760_ = new_n919_ & ~new_n10759_;
  assign new_n10761_ = new_n923_ & ~new_n10760_;
  assign new_n10762_ = new_n927_ & ~new_n10761_;
  assign new_n10763_ = new_n931_ & ~new_n10762_;
  assign new_n10764_ = new_n935_ & ~new_n10763_;
  assign new_n10765_ = new_n939_ & ~new_n10764_;
  assign new_n10766_ = new_n943_ & ~new_n10765_;
  assign new_n10767_ = new_n947_ & ~new_n10766_;
  assign new_n10768_ = new_n951_ & ~new_n10767_;
  assign new_n10769_ = new_n955_ & ~new_n10768_;
  assign new_n10770_ = new_n959_ & ~new_n10769_;
  assign new_n10771_ = new_n963_ & ~new_n10770_;
  assign new_n10772_ = new_n967_ & ~new_n10771_;
  assign new_n10773_ = new_n971_ & ~new_n10772_;
  assign new_n10774_ = new_n975_ & ~new_n10773_;
  assign new_n10775_ = new_n979_ & ~new_n10774_;
  assign new_n10776_ = new_n983_ & ~new_n10775_;
  assign new_n10777_ = new_n987_ & ~new_n10776_;
  assign new_n10778_ = new_n991_ & ~new_n10777_;
  assign new_n10779_ = new_n995_ & ~new_n10778_;
  assign new_n10780_ = new_n999_ & ~new_n10779_;
  assign new_n10781_ = new_n1003_ & ~new_n10780_;
  assign new_n10782_ = new_n1007_ & ~new_n10781_;
  assign new_n10783_ = new_n1011_ & ~new_n10782_;
  assign new_n10784_ = \req[111]  & ~new_n1013_;
  assign \grant[111]  = ~new_n10783_ & new_n10784_;
  assign new_n10786_ = new_n1022_ & ~new_n1355_;
  assign new_n10787_ = new_n1027_ & ~new_n10786_;
  assign new_n10788_ = new_n1031_ & ~new_n10787_;
  assign new_n10789_ = new_n1035_ & ~new_n10788_;
  assign new_n10790_ = new_n1039_ & ~new_n10789_;
  assign new_n10791_ = new_n1043_ & ~new_n10790_;
  assign new_n10792_ = new_n1047_ & ~new_n10791_;
  assign new_n10793_ = new_n1051_ & ~new_n10792_;
  assign new_n10794_ = new_n1055_ & ~new_n10793_;
  assign new_n10795_ = new_n1059_ & ~new_n10794_;
  assign new_n10796_ = new_n1574_ & ~new_n10795_;
  assign new_n10797_ = new_n1576_ & ~new_n10796_;
  assign new_n10798_ = new_n1837_ & ~new_n10797_;
  assign new_n10799_ = new_n1068_ & ~new_n10798_;
  assign new_n10800_ = new_n1072_ & ~new_n10799_;
  assign new_n10801_ = new_n1076_ & ~new_n10800_;
  assign new_n10802_ = new_n1080_ & ~new_n10801_;
  assign new_n10803_ = new_n1084_ & ~new_n10802_;
  assign new_n10804_ = new_n1088_ & ~new_n10803_;
  assign new_n10805_ = new_n1092_ & ~new_n10804_;
  assign new_n10806_ = new_n1096_ & ~new_n10805_;
  assign new_n10807_ = new_n1100_ & ~new_n10806_;
  assign new_n10808_ = new_n1104_ & ~new_n10807_;
  assign new_n10809_ = new_n1108_ & ~new_n10808_;
  assign new_n10810_ = new_n1112_ & ~new_n10809_;
  assign new_n10811_ = new_n1116_ & ~new_n10810_;
  assign new_n10812_ = new_n1120_ & ~new_n10811_;
  assign new_n10813_ = new_n1124_ & ~new_n10812_;
  assign new_n10814_ = new_n1128_ & ~new_n10813_;
  assign new_n10815_ = new_n1132_ & ~new_n10814_;
  assign new_n10816_ = new_n1136_ & ~new_n10815_;
  assign new_n10817_ = new_n1140_ & ~new_n10816_;
  assign new_n10818_ = new_n1144_ & ~new_n10817_;
  assign new_n10819_ = new_n1148_ & ~new_n10818_;
  assign new_n10820_ = new_n1152_ & ~new_n10819_;
  assign new_n10821_ = new_n1156_ & ~new_n10820_;
  assign new_n10822_ = new_n1160_ & ~new_n10821_;
  assign new_n10823_ = new_n1164_ & ~new_n10822_;
  assign new_n10824_ = new_n1168_ & ~new_n10823_;
  assign new_n10825_ = new_n1172_ & ~new_n10824_;
  assign new_n10826_ = new_n1176_ & ~new_n10825_;
  assign new_n10827_ = new_n1180_ & ~new_n10826_;
  assign new_n10828_ = new_n1184_ & ~new_n10827_;
  assign new_n10829_ = new_n1188_ & ~new_n10828_;
  assign new_n10830_ = new_n1192_ & ~new_n10829_;
  assign new_n10831_ = new_n1196_ & ~new_n10830_;
  assign new_n10832_ = new_n1200_ & ~new_n10831_;
  assign new_n10833_ = new_n1204_ & ~new_n10832_;
  assign new_n10834_ = new_n1208_ & ~new_n10833_;
  assign new_n10835_ = new_n1212_ & ~new_n10834_;
  assign new_n10836_ = new_n1216_ & ~new_n10835_;
  assign new_n10837_ = new_n1220_ & ~new_n10836_;
  assign new_n10838_ = new_n1224_ & ~new_n10837_;
  assign new_n10839_ = new_n1228_ & ~new_n10838_;
  assign new_n10840_ = new_n1232_ & ~new_n10839_;
  assign new_n10841_ = new_n1236_ & ~new_n10840_;
  assign new_n10842_ = new_n1240_ & ~new_n10841_;
  assign new_n10843_ = new_n1244_ & ~new_n10842_;
  assign new_n10844_ = new_n1248_ & ~new_n10843_;
  assign new_n10845_ = new_n1252_ & ~new_n10844_;
  assign new_n10846_ = new_n1256_ & ~new_n10845_;
  assign new_n10847_ = new_n1260_ & ~new_n10846_;
  assign new_n10848_ = new_n1264_ & ~new_n10847_;
  assign new_n10849_ = new_n1268_ & ~new_n10848_;
  assign new_n10850_ = new_n1272_ & ~new_n10849_;
  assign new_n10851_ = new_n1276_ & ~new_n10850_;
  assign new_n10852_ = new_n1280_ & ~new_n10851_;
  assign new_n10853_ = new_n1284_ & ~new_n10852_;
  assign new_n10854_ = new_n1288_ & ~new_n10853_;
  assign new_n10855_ = new_n1292_ & ~new_n10854_;
  assign new_n10856_ = new_n1296_ & ~new_n10855_;
  assign new_n10857_ = new_n1300_ & ~new_n10856_;
  assign new_n10858_ = new_n1304_ & ~new_n10857_;
  assign new_n10859_ = new_n1308_ & ~new_n10858_;
  assign new_n10860_ = new_n1312_ & ~new_n10859_;
  assign new_n10861_ = new_n1316_ & ~new_n10860_;
  assign new_n10862_ = new_n1320_ & ~new_n10861_;
  assign new_n10863_ = new_n1324_ & ~new_n10862_;
  assign new_n10864_ = new_n1328_ & ~new_n10863_;
  assign new_n10865_ = new_n1332_ & ~new_n10864_;
  assign new_n10866_ = new_n1336_ & ~new_n10865_;
  assign new_n10867_ = new_n1340_ & ~new_n10866_;
  assign new_n10868_ = new_n1344_ & ~new_n10867_;
  assign new_n10869_ = new_n1348_ & ~new_n10868_;
  assign new_n10870_ = \req[112]  & ~new_n1350_;
  assign \grant[112]  = ~new_n10869_ & new_n10870_;
  assign new_n10872_ = ~new_n687_ & new_n1359_;
  assign new_n10873_ = new_n1364_ & ~new_n10872_;
  assign new_n10874_ = new_n1368_ & ~new_n10873_;
  assign new_n10875_ = new_n1372_ & ~new_n10874_;
  assign new_n10876_ = new_n1376_ & ~new_n10875_;
  assign new_n10877_ = new_n1380_ & ~new_n10876_;
  assign new_n10878_ = new_n1384_ & ~new_n10877_;
  assign new_n10879_ = new_n1388_ & ~new_n10878_;
  assign new_n10880_ = new_n1392_ & ~new_n10879_;
  assign new_n10881_ = new_n1396_ & ~new_n10880_;
  assign new_n10882_ = new_n1663_ & ~new_n10881_;
  assign new_n10883_ = new_n392_ & ~new_n10882_;
  assign new_n10884_ = new_n396_ & ~new_n10883_;
  assign new_n10885_ = new_n400_ & ~new_n10884_;
  assign new_n10886_ = new_n404_ & ~new_n10885_;
  assign new_n10887_ = new_n408_ & ~new_n10886_;
  assign new_n10888_ = new_n412_ & ~new_n10887_;
  assign new_n10889_ = new_n416_ & ~new_n10888_;
  assign new_n10890_ = new_n420_ & ~new_n10889_;
  assign new_n10891_ = new_n424_ & ~new_n10890_;
  assign new_n10892_ = new_n428_ & ~new_n10891_;
  assign new_n10893_ = new_n432_ & ~new_n10892_;
  assign new_n10894_ = new_n436_ & ~new_n10893_;
  assign new_n10895_ = new_n440_ & ~new_n10894_;
  assign new_n10896_ = new_n444_ & ~new_n10895_;
  assign new_n10897_ = new_n448_ & ~new_n10896_;
  assign new_n10898_ = new_n452_ & ~new_n10897_;
  assign new_n10899_ = new_n456_ & ~new_n10898_;
  assign new_n10900_ = new_n460_ & ~new_n10899_;
  assign new_n10901_ = new_n464_ & ~new_n10900_;
  assign new_n10902_ = new_n468_ & ~new_n10901_;
  assign new_n10903_ = new_n472_ & ~new_n10902_;
  assign new_n10904_ = new_n476_ & ~new_n10903_;
  assign new_n10905_ = new_n480_ & ~new_n10904_;
  assign new_n10906_ = new_n484_ & ~new_n10905_;
  assign new_n10907_ = new_n488_ & ~new_n10906_;
  assign new_n10908_ = new_n492_ & ~new_n10907_;
  assign new_n10909_ = new_n496_ & ~new_n10908_;
  assign new_n10910_ = new_n500_ & ~new_n10909_;
  assign new_n10911_ = new_n504_ & ~new_n10910_;
  assign new_n10912_ = new_n508_ & ~new_n10911_;
  assign new_n10913_ = new_n512_ & ~new_n10912_;
  assign new_n10914_ = new_n516_ & ~new_n10913_;
  assign new_n10915_ = new_n520_ & ~new_n10914_;
  assign new_n10916_ = new_n524_ & ~new_n10915_;
  assign new_n10917_ = new_n528_ & ~new_n10916_;
  assign new_n10918_ = new_n532_ & ~new_n10917_;
  assign new_n10919_ = new_n536_ & ~new_n10918_;
  assign new_n10920_ = new_n540_ & ~new_n10919_;
  assign new_n10921_ = new_n544_ & ~new_n10920_;
  assign new_n10922_ = new_n548_ & ~new_n10921_;
  assign new_n10923_ = new_n552_ & ~new_n10922_;
  assign new_n10924_ = new_n556_ & ~new_n10923_;
  assign new_n10925_ = new_n560_ & ~new_n10924_;
  assign new_n10926_ = new_n564_ & ~new_n10925_;
  assign new_n10927_ = new_n568_ & ~new_n10926_;
  assign new_n10928_ = new_n572_ & ~new_n10927_;
  assign new_n10929_ = new_n576_ & ~new_n10928_;
  assign new_n10930_ = new_n580_ & ~new_n10929_;
  assign new_n10931_ = new_n584_ & ~new_n10930_;
  assign new_n10932_ = new_n588_ & ~new_n10931_;
  assign new_n10933_ = new_n592_ & ~new_n10932_;
  assign new_n10934_ = new_n596_ & ~new_n10933_;
  assign new_n10935_ = new_n600_ & ~new_n10934_;
  assign new_n10936_ = new_n604_ & ~new_n10935_;
  assign new_n10937_ = new_n608_ & ~new_n10936_;
  assign new_n10938_ = new_n612_ & ~new_n10937_;
  assign new_n10939_ = new_n616_ & ~new_n10938_;
  assign new_n10940_ = new_n620_ & ~new_n10939_;
  assign new_n10941_ = new_n624_ & ~new_n10940_;
  assign new_n10942_ = new_n628_ & ~new_n10941_;
  assign new_n10943_ = new_n632_ & ~new_n10942_;
  assign new_n10944_ = new_n636_ & ~new_n10943_;
  assign new_n10945_ = new_n640_ & ~new_n10944_;
  assign new_n10946_ = new_n644_ & ~new_n10945_;
  assign new_n10947_ = new_n648_ & ~new_n10946_;
  assign new_n10948_ = new_n652_ & ~new_n10947_;
  assign new_n10949_ = new_n656_ & ~new_n10948_;
  assign new_n10950_ = new_n660_ & ~new_n10949_;
  assign new_n10951_ = new_n664_ & ~new_n10950_;
  assign new_n10952_ = new_n668_ & ~new_n10951_;
  assign new_n10953_ = new_n672_ & ~new_n10952_;
  assign new_n10954_ = new_n676_ & ~new_n10953_;
  assign new_n10955_ = new_n680_ & ~new_n10954_;
  assign new_n10956_ = \req[113]  & ~new_n682_;
  assign \grant[113]  = ~new_n10955_ & new_n10956_;
  assign new_n10958_ = new_n691_ & ~new_n1026_;
  assign new_n10959_ = new_n696_ & ~new_n10958_;
  assign new_n10960_ = new_n700_ & ~new_n10959_;
  assign new_n10961_ = new_n704_ & ~new_n10960_;
  assign new_n10962_ = new_n708_ & ~new_n10961_;
  assign new_n10963_ = new_n712_ & ~new_n10962_;
  assign new_n10964_ = new_n716_ & ~new_n10963_;
  assign new_n10965_ = new_n720_ & ~new_n10964_;
  assign new_n10966_ = new_n1484_ & ~new_n10965_;
  assign new_n10967_ = new_n1486_ & ~new_n10966_;
  assign new_n10968_ = new_n1750_ & ~new_n10967_;
  assign new_n10969_ = new_n731_ & ~new_n10968_;
  assign new_n10970_ = new_n735_ & ~new_n10969_;
  assign new_n10971_ = new_n739_ & ~new_n10970_;
  assign new_n10972_ = new_n743_ & ~new_n10971_;
  assign new_n10973_ = new_n747_ & ~new_n10972_;
  assign new_n10974_ = new_n751_ & ~new_n10973_;
  assign new_n10975_ = new_n755_ & ~new_n10974_;
  assign new_n10976_ = new_n759_ & ~new_n10975_;
  assign new_n10977_ = new_n763_ & ~new_n10976_;
  assign new_n10978_ = new_n767_ & ~new_n10977_;
  assign new_n10979_ = new_n771_ & ~new_n10978_;
  assign new_n10980_ = new_n775_ & ~new_n10979_;
  assign new_n10981_ = new_n779_ & ~new_n10980_;
  assign new_n10982_ = new_n783_ & ~new_n10981_;
  assign new_n10983_ = new_n787_ & ~new_n10982_;
  assign new_n10984_ = new_n791_ & ~new_n10983_;
  assign new_n10985_ = new_n795_ & ~new_n10984_;
  assign new_n10986_ = new_n799_ & ~new_n10985_;
  assign new_n10987_ = new_n803_ & ~new_n10986_;
  assign new_n10988_ = new_n807_ & ~new_n10987_;
  assign new_n10989_ = new_n811_ & ~new_n10988_;
  assign new_n10990_ = new_n815_ & ~new_n10989_;
  assign new_n10991_ = new_n819_ & ~new_n10990_;
  assign new_n10992_ = new_n823_ & ~new_n10991_;
  assign new_n10993_ = new_n827_ & ~new_n10992_;
  assign new_n10994_ = new_n831_ & ~new_n10993_;
  assign new_n10995_ = new_n835_ & ~new_n10994_;
  assign new_n10996_ = new_n839_ & ~new_n10995_;
  assign new_n10997_ = new_n843_ & ~new_n10996_;
  assign new_n10998_ = new_n847_ & ~new_n10997_;
  assign new_n10999_ = new_n851_ & ~new_n10998_;
  assign new_n11000_ = new_n855_ & ~new_n10999_;
  assign new_n11001_ = new_n859_ & ~new_n11000_;
  assign new_n11002_ = new_n863_ & ~new_n11001_;
  assign new_n11003_ = new_n867_ & ~new_n11002_;
  assign new_n11004_ = new_n871_ & ~new_n11003_;
  assign new_n11005_ = new_n875_ & ~new_n11004_;
  assign new_n11006_ = new_n879_ & ~new_n11005_;
  assign new_n11007_ = new_n883_ & ~new_n11006_;
  assign new_n11008_ = new_n887_ & ~new_n11007_;
  assign new_n11009_ = new_n891_ & ~new_n11008_;
  assign new_n11010_ = new_n895_ & ~new_n11009_;
  assign new_n11011_ = new_n899_ & ~new_n11010_;
  assign new_n11012_ = new_n903_ & ~new_n11011_;
  assign new_n11013_ = new_n907_ & ~new_n11012_;
  assign new_n11014_ = new_n911_ & ~new_n11013_;
  assign new_n11015_ = new_n915_ & ~new_n11014_;
  assign new_n11016_ = new_n919_ & ~new_n11015_;
  assign new_n11017_ = new_n923_ & ~new_n11016_;
  assign new_n11018_ = new_n927_ & ~new_n11017_;
  assign new_n11019_ = new_n931_ & ~new_n11018_;
  assign new_n11020_ = new_n935_ & ~new_n11019_;
  assign new_n11021_ = new_n939_ & ~new_n11020_;
  assign new_n11022_ = new_n943_ & ~new_n11021_;
  assign new_n11023_ = new_n947_ & ~new_n11022_;
  assign new_n11024_ = new_n951_ & ~new_n11023_;
  assign new_n11025_ = new_n955_ & ~new_n11024_;
  assign new_n11026_ = new_n959_ & ~new_n11025_;
  assign new_n11027_ = new_n963_ & ~new_n11026_;
  assign new_n11028_ = new_n967_ & ~new_n11027_;
  assign new_n11029_ = new_n971_ & ~new_n11028_;
  assign new_n11030_ = new_n975_ & ~new_n11029_;
  assign new_n11031_ = new_n979_ & ~new_n11030_;
  assign new_n11032_ = new_n983_ & ~new_n11031_;
  assign new_n11033_ = new_n987_ & ~new_n11032_;
  assign new_n11034_ = new_n991_ & ~new_n11033_;
  assign new_n11035_ = new_n995_ & ~new_n11034_;
  assign new_n11036_ = new_n999_ & ~new_n11035_;
  assign new_n11037_ = new_n1003_ & ~new_n11036_;
  assign new_n11038_ = new_n1007_ & ~new_n11037_;
  assign new_n11039_ = new_n1011_ & ~new_n11038_;
  assign new_n11040_ = new_n1015_ & ~new_n11039_;
  assign new_n11041_ = new_n1019_ & ~new_n11040_;
  assign new_n11042_ = \req[114]  & ~new_n1021_;
  assign \grant[114]  = ~new_n11041_ & new_n11042_;
  assign new_n11044_ = new_n1030_ & ~new_n1363_;
  assign new_n11045_ = new_n1035_ & ~new_n11044_;
  assign new_n11046_ = new_n1039_ & ~new_n11045_;
  assign new_n11047_ = new_n1043_ & ~new_n11046_;
  assign new_n11048_ = new_n1047_ & ~new_n11047_;
  assign new_n11049_ = new_n1051_ & ~new_n11048_;
  assign new_n11050_ = new_n1055_ & ~new_n11049_;
  assign new_n11051_ = new_n1059_ & ~new_n11050_;
  assign new_n11052_ = new_n1574_ & ~new_n11051_;
  assign new_n11053_ = new_n1576_ & ~new_n11052_;
  assign new_n11054_ = new_n1837_ & ~new_n11053_;
  assign new_n11055_ = new_n1068_ & ~new_n11054_;
  assign new_n11056_ = new_n1072_ & ~new_n11055_;
  assign new_n11057_ = new_n1076_ & ~new_n11056_;
  assign new_n11058_ = new_n1080_ & ~new_n11057_;
  assign new_n11059_ = new_n1084_ & ~new_n11058_;
  assign new_n11060_ = new_n1088_ & ~new_n11059_;
  assign new_n11061_ = new_n1092_ & ~new_n11060_;
  assign new_n11062_ = new_n1096_ & ~new_n11061_;
  assign new_n11063_ = new_n1100_ & ~new_n11062_;
  assign new_n11064_ = new_n1104_ & ~new_n11063_;
  assign new_n11065_ = new_n1108_ & ~new_n11064_;
  assign new_n11066_ = new_n1112_ & ~new_n11065_;
  assign new_n11067_ = new_n1116_ & ~new_n11066_;
  assign new_n11068_ = new_n1120_ & ~new_n11067_;
  assign new_n11069_ = new_n1124_ & ~new_n11068_;
  assign new_n11070_ = new_n1128_ & ~new_n11069_;
  assign new_n11071_ = new_n1132_ & ~new_n11070_;
  assign new_n11072_ = new_n1136_ & ~new_n11071_;
  assign new_n11073_ = new_n1140_ & ~new_n11072_;
  assign new_n11074_ = new_n1144_ & ~new_n11073_;
  assign new_n11075_ = new_n1148_ & ~new_n11074_;
  assign new_n11076_ = new_n1152_ & ~new_n11075_;
  assign new_n11077_ = new_n1156_ & ~new_n11076_;
  assign new_n11078_ = new_n1160_ & ~new_n11077_;
  assign new_n11079_ = new_n1164_ & ~new_n11078_;
  assign new_n11080_ = new_n1168_ & ~new_n11079_;
  assign new_n11081_ = new_n1172_ & ~new_n11080_;
  assign new_n11082_ = new_n1176_ & ~new_n11081_;
  assign new_n11083_ = new_n1180_ & ~new_n11082_;
  assign new_n11084_ = new_n1184_ & ~new_n11083_;
  assign new_n11085_ = new_n1188_ & ~new_n11084_;
  assign new_n11086_ = new_n1192_ & ~new_n11085_;
  assign new_n11087_ = new_n1196_ & ~new_n11086_;
  assign new_n11088_ = new_n1200_ & ~new_n11087_;
  assign new_n11089_ = new_n1204_ & ~new_n11088_;
  assign new_n11090_ = new_n1208_ & ~new_n11089_;
  assign new_n11091_ = new_n1212_ & ~new_n11090_;
  assign new_n11092_ = new_n1216_ & ~new_n11091_;
  assign new_n11093_ = new_n1220_ & ~new_n11092_;
  assign new_n11094_ = new_n1224_ & ~new_n11093_;
  assign new_n11095_ = new_n1228_ & ~new_n11094_;
  assign new_n11096_ = new_n1232_ & ~new_n11095_;
  assign new_n11097_ = new_n1236_ & ~new_n11096_;
  assign new_n11098_ = new_n1240_ & ~new_n11097_;
  assign new_n11099_ = new_n1244_ & ~new_n11098_;
  assign new_n11100_ = new_n1248_ & ~new_n11099_;
  assign new_n11101_ = new_n1252_ & ~new_n11100_;
  assign new_n11102_ = new_n1256_ & ~new_n11101_;
  assign new_n11103_ = new_n1260_ & ~new_n11102_;
  assign new_n11104_ = new_n1264_ & ~new_n11103_;
  assign new_n11105_ = new_n1268_ & ~new_n11104_;
  assign new_n11106_ = new_n1272_ & ~new_n11105_;
  assign new_n11107_ = new_n1276_ & ~new_n11106_;
  assign new_n11108_ = new_n1280_ & ~new_n11107_;
  assign new_n11109_ = new_n1284_ & ~new_n11108_;
  assign new_n11110_ = new_n1288_ & ~new_n11109_;
  assign new_n11111_ = new_n1292_ & ~new_n11110_;
  assign new_n11112_ = new_n1296_ & ~new_n11111_;
  assign new_n11113_ = new_n1300_ & ~new_n11112_;
  assign new_n11114_ = new_n1304_ & ~new_n11113_;
  assign new_n11115_ = new_n1308_ & ~new_n11114_;
  assign new_n11116_ = new_n1312_ & ~new_n11115_;
  assign new_n11117_ = new_n1316_ & ~new_n11116_;
  assign new_n11118_ = new_n1320_ & ~new_n11117_;
  assign new_n11119_ = new_n1324_ & ~new_n11118_;
  assign new_n11120_ = new_n1328_ & ~new_n11119_;
  assign new_n11121_ = new_n1332_ & ~new_n11120_;
  assign new_n11122_ = new_n1336_ & ~new_n11121_;
  assign new_n11123_ = new_n1340_ & ~new_n11122_;
  assign new_n11124_ = new_n1344_ & ~new_n11123_;
  assign new_n11125_ = new_n1348_ & ~new_n11124_;
  assign new_n11126_ = new_n1352_ & ~new_n11125_;
  assign new_n11127_ = new_n1356_ & ~new_n11126_;
  assign new_n11128_ = \req[115]  & ~new_n1358_;
  assign \grant[115]  = ~new_n11127_ & new_n11128_;
  assign new_n11130_ = ~new_n695_ & new_n1367_;
  assign new_n11131_ = new_n1372_ & ~new_n11130_;
  assign new_n11132_ = new_n1376_ & ~new_n11131_;
  assign new_n11133_ = new_n1380_ & ~new_n11132_;
  assign new_n11134_ = new_n1384_ & ~new_n11133_;
  assign new_n11135_ = new_n1388_ & ~new_n11134_;
  assign new_n11136_ = new_n1392_ & ~new_n11135_;
  assign new_n11137_ = new_n1396_ & ~new_n11136_;
  assign new_n11138_ = new_n1663_ & ~new_n11137_;
  assign new_n11139_ = new_n392_ & ~new_n11138_;
  assign new_n11140_ = new_n396_ & ~new_n11139_;
  assign new_n11141_ = new_n400_ & ~new_n11140_;
  assign new_n11142_ = new_n404_ & ~new_n11141_;
  assign new_n11143_ = new_n408_ & ~new_n11142_;
  assign new_n11144_ = new_n412_ & ~new_n11143_;
  assign new_n11145_ = new_n416_ & ~new_n11144_;
  assign new_n11146_ = new_n420_ & ~new_n11145_;
  assign new_n11147_ = new_n424_ & ~new_n11146_;
  assign new_n11148_ = new_n428_ & ~new_n11147_;
  assign new_n11149_ = new_n432_ & ~new_n11148_;
  assign new_n11150_ = new_n436_ & ~new_n11149_;
  assign new_n11151_ = new_n440_ & ~new_n11150_;
  assign new_n11152_ = new_n444_ & ~new_n11151_;
  assign new_n11153_ = new_n448_ & ~new_n11152_;
  assign new_n11154_ = new_n452_ & ~new_n11153_;
  assign new_n11155_ = new_n456_ & ~new_n11154_;
  assign new_n11156_ = new_n460_ & ~new_n11155_;
  assign new_n11157_ = new_n464_ & ~new_n11156_;
  assign new_n11158_ = new_n468_ & ~new_n11157_;
  assign new_n11159_ = new_n472_ & ~new_n11158_;
  assign new_n11160_ = new_n476_ & ~new_n11159_;
  assign new_n11161_ = new_n480_ & ~new_n11160_;
  assign new_n11162_ = new_n484_ & ~new_n11161_;
  assign new_n11163_ = new_n488_ & ~new_n11162_;
  assign new_n11164_ = new_n492_ & ~new_n11163_;
  assign new_n11165_ = new_n496_ & ~new_n11164_;
  assign new_n11166_ = new_n500_ & ~new_n11165_;
  assign new_n11167_ = new_n504_ & ~new_n11166_;
  assign new_n11168_ = new_n508_ & ~new_n11167_;
  assign new_n11169_ = new_n512_ & ~new_n11168_;
  assign new_n11170_ = new_n516_ & ~new_n11169_;
  assign new_n11171_ = new_n520_ & ~new_n11170_;
  assign new_n11172_ = new_n524_ & ~new_n11171_;
  assign new_n11173_ = new_n528_ & ~new_n11172_;
  assign new_n11174_ = new_n532_ & ~new_n11173_;
  assign new_n11175_ = new_n536_ & ~new_n11174_;
  assign new_n11176_ = new_n540_ & ~new_n11175_;
  assign new_n11177_ = new_n544_ & ~new_n11176_;
  assign new_n11178_ = new_n548_ & ~new_n11177_;
  assign new_n11179_ = new_n552_ & ~new_n11178_;
  assign new_n11180_ = new_n556_ & ~new_n11179_;
  assign new_n11181_ = new_n560_ & ~new_n11180_;
  assign new_n11182_ = new_n564_ & ~new_n11181_;
  assign new_n11183_ = new_n568_ & ~new_n11182_;
  assign new_n11184_ = new_n572_ & ~new_n11183_;
  assign new_n11185_ = new_n576_ & ~new_n11184_;
  assign new_n11186_ = new_n580_ & ~new_n11185_;
  assign new_n11187_ = new_n584_ & ~new_n11186_;
  assign new_n11188_ = new_n588_ & ~new_n11187_;
  assign new_n11189_ = new_n592_ & ~new_n11188_;
  assign new_n11190_ = new_n596_ & ~new_n11189_;
  assign new_n11191_ = new_n600_ & ~new_n11190_;
  assign new_n11192_ = new_n604_ & ~new_n11191_;
  assign new_n11193_ = new_n608_ & ~new_n11192_;
  assign new_n11194_ = new_n612_ & ~new_n11193_;
  assign new_n11195_ = new_n616_ & ~new_n11194_;
  assign new_n11196_ = new_n620_ & ~new_n11195_;
  assign new_n11197_ = new_n624_ & ~new_n11196_;
  assign new_n11198_ = new_n628_ & ~new_n11197_;
  assign new_n11199_ = new_n632_ & ~new_n11198_;
  assign new_n11200_ = new_n636_ & ~new_n11199_;
  assign new_n11201_ = new_n640_ & ~new_n11200_;
  assign new_n11202_ = new_n644_ & ~new_n11201_;
  assign new_n11203_ = new_n648_ & ~new_n11202_;
  assign new_n11204_ = new_n652_ & ~new_n11203_;
  assign new_n11205_ = new_n656_ & ~new_n11204_;
  assign new_n11206_ = new_n660_ & ~new_n11205_;
  assign new_n11207_ = new_n664_ & ~new_n11206_;
  assign new_n11208_ = new_n668_ & ~new_n11207_;
  assign new_n11209_ = new_n672_ & ~new_n11208_;
  assign new_n11210_ = new_n676_ & ~new_n11209_;
  assign new_n11211_ = new_n680_ & ~new_n11210_;
  assign new_n11212_ = new_n684_ & ~new_n11211_;
  assign new_n11213_ = new_n688_ & ~new_n11212_;
  assign new_n11214_ = \req[116]  & ~new_n690_;
  assign \grant[116]  = ~new_n11213_ & new_n11214_;
  assign new_n11216_ = new_n699_ & ~new_n1034_;
  assign new_n11217_ = new_n704_ & ~new_n11216_;
  assign new_n11218_ = new_n708_ & ~new_n11217_;
  assign new_n11219_ = new_n712_ & ~new_n11218_;
  assign new_n11220_ = new_n716_ & ~new_n11219_;
  assign new_n11221_ = new_n720_ & ~new_n11220_;
  assign new_n11222_ = new_n1484_ & ~new_n11221_;
  assign new_n11223_ = new_n1486_ & ~new_n11222_;
  assign new_n11224_ = new_n1750_ & ~new_n11223_;
  assign new_n11225_ = new_n731_ & ~new_n11224_;
  assign new_n11226_ = new_n735_ & ~new_n11225_;
  assign new_n11227_ = new_n739_ & ~new_n11226_;
  assign new_n11228_ = new_n743_ & ~new_n11227_;
  assign new_n11229_ = new_n747_ & ~new_n11228_;
  assign new_n11230_ = new_n751_ & ~new_n11229_;
  assign new_n11231_ = new_n755_ & ~new_n11230_;
  assign new_n11232_ = new_n759_ & ~new_n11231_;
  assign new_n11233_ = new_n763_ & ~new_n11232_;
  assign new_n11234_ = new_n767_ & ~new_n11233_;
  assign new_n11235_ = new_n771_ & ~new_n11234_;
  assign new_n11236_ = new_n775_ & ~new_n11235_;
  assign new_n11237_ = new_n779_ & ~new_n11236_;
  assign new_n11238_ = new_n783_ & ~new_n11237_;
  assign new_n11239_ = new_n787_ & ~new_n11238_;
  assign new_n11240_ = new_n791_ & ~new_n11239_;
  assign new_n11241_ = new_n795_ & ~new_n11240_;
  assign new_n11242_ = new_n799_ & ~new_n11241_;
  assign new_n11243_ = new_n803_ & ~new_n11242_;
  assign new_n11244_ = new_n807_ & ~new_n11243_;
  assign new_n11245_ = new_n811_ & ~new_n11244_;
  assign new_n11246_ = new_n815_ & ~new_n11245_;
  assign new_n11247_ = new_n819_ & ~new_n11246_;
  assign new_n11248_ = new_n823_ & ~new_n11247_;
  assign new_n11249_ = new_n827_ & ~new_n11248_;
  assign new_n11250_ = new_n831_ & ~new_n11249_;
  assign new_n11251_ = new_n835_ & ~new_n11250_;
  assign new_n11252_ = new_n839_ & ~new_n11251_;
  assign new_n11253_ = new_n843_ & ~new_n11252_;
  assign new_n11254_ = new_n847_ & ~new_n11253_;
  assign new_n11255_ = new_n851_ & ~new_n11254_;
  assign new_n11256_ = new_n855_ & ~new_n11255_;
  assign new_n11257_ = new_n859_ & ~new_n11256_;
  assign new_n11258_ = new_n863_ & ~new_n11257_;
  assign new_n11259_ = new_n867_ & ~new_n11258_;
  assign new_n11260_ = new_n871_ & ~new_n11259_;
  assign new_n11261_ = new_n875_ & ~new_n11260_;
  assign new_n11262_ = new_n879_ & ~new_n11261_;
  assign new_n11263_ = new_n883_ & ~new_n11262_;
  assign new_n11264_ = new_n887_ & ~new_n11263_;
  assign new_n11265_ = new_n891_ & ~new_n11264_;
  assign new_n11266_ = new_n895_ & ~new_n11265_;
  assign new_n11267_ = new_n899_ & ~new_n11266_;
  assign new_n11268_ = new_n903_ & ~new_n11267_;
  assign new_n11269_ = new_n907_ & ~new_n11268_;
  assign new_n11270_ = new_n911_ & ~new_n11269_;
  assign new_n11271_ = new_n915_ & ~new_n11270_;
  assign new_n11272_ = new_n919_ & ~new_n11271_;
  assign new_n11273_ = new_n923_ & ~new_n11272_;
  assign new_n11274_ = new_n927_ & ~new_n11273_;
  assign new_n11275_ = new_n931_ & ~new_n11274_;
  assign new_n11276_ = new_n935_ & ~new_n11275_;
  assign new_n11277_ = new_n939_ & ~new_n11276_;
  assign new_n11278_ = new_n943_ & ~new_n11277_;
  assign new_n11279_ = new_n947_ & ~new_n11278_;
  assign new_n11280_ = new_n951_ & ~new_n11279_;
  assign new_n11281_ = new_n955_ & ~new_n11280_;
  assign new_n11282_ = new_n959_ & ~new_n11281_;
  assign new_n11283_ = new_n963_ & ~new_n11282_;
  assign new_n11284_ = new_n967_ & ~new_n11283_;
  assign new_n11285_ = new_n971_ & ~new_n11284_;
  assign new_n11286_ = new_n975_ & ~new_n11285_;
  assign new_n11287_ = new_n979_ & ~new_n11286_;
  assign new_n11288_ = new_n983_ & ~new_n11287_;
  assign new_n11289_ = new_n987_ & ~new_n11288_;
  assign new_n11290_ = new_n991_ & ~new_n11289_;
  assign new_n11291_ = new_n995_ & ~new_n11290_;
  assign new_n11292_ = new_n999_ & ~new_n11291_;
  assign new_n11293_ = new_n1003_ & ~new_n11292_;
  assign new_n11294_ = new_n1007_ & ~new_n11293_;
  assign new_n11295_ = new_n1011_ & ~new_n11294_;
  assign new_n11296_ = new_n1015_ & ~new_n11295_;
  assign new_n11297_ = new_n1019_ & ~new_n11296_;
  assign new_n11298_ = new_n1023_ & ~new_n11297_;
  assign new_n11299_ = new_n1027_ & ~new_n11298_;
  assign new_n11300_ = \req[117]  & ~new_n1029_;
  assign \grant[117]  = ~new_n11299_ & new_n11300_;
  assign new_n11302_ = new_n1038_ & ~new_n1371_;
  assign new_n11303_ = new_n1043_ & ~new_n11302_;
  assign new_n11304_ = new_n1047_ & ~new_n11303_;
  assign new_n11305_ = new_n1051_ & ~new_n11304_;
  assign new_n11306_ = new_n1055_ & ~new_n11305_;
  assign new_n11307_ = new_n1059_ & ~new_n11306_;
  assign new_n11308_ = new_n1574_ & ~new_n11307_;
  assign new_n11309_ = new_n1576_ & ~new_n11308_;
  assign new_n11310_ = new_n1837_ & ~new_n11309_;
  assign new_n11311_ = new_n1068_ & ~new_n11310_;
  assign new_n11312_ = new_n1072_ & ~new_n11311_;
  assign new_n11313_ = new_n1076_ & ~new_n11312_;
  assign new_n11314_ = new_n1080_ & ~new_n11313_;
  assign new_n11315_ = new_n1084_ & ~new_n11314_;
  assign new_n11316_ = new_n1088_ & ~new_n11315_;
  assign new_n11317_ = new_n1092_ & ~new_n11316_;
  assign new_n11318_ = new_n1096_ & ~new_n11317_;
  assign new_n11319_ = new_n1100_ & ~new_n11318_;
  assign new_n11320_ = new_n1104_ & ~new_n11319_;
  assign new_n11321_ = new_n1108_ & ~new_n11320_;
  assign new_n11322_ = new_n1112_ & ~new_n11321_;
  assign new_n11323_ = new_n1116_ & ~new_n11322_;
  assign new_n11324_ = new_n1120_ & ~new_n11323_;
  assign new_n11325_ = new_n1124_ & ~new_n11324_;
  assign new_n11326_ = new_n1128_ & ~new_n11325_;
  assign new_n11327_ = new_n1132_ & ~new_n11326_;
  assign new_n11328_ = new_n1136_ & ~new_n11327_;
  assign new_n11329_ = new_n1140_ & ~new_n11328_;
  assign new_n11330_ = new_n1144_ & ~new_n11329_;
  assign new_n11331_ = new_n1148_ & ~new_n11330_;
  assign new_n11332_ = new_n1152_ & ~new_n11331_;
  assign new_n11333_ = new_n1156_ & ~new_n11332_;
  assign new_n11334_ = new_n1160_ & ~new_n11333_;
  assign new_n11335_ = new_n1164_ & ~new_n11334_;
  assign new_n11336_ = new_n1168_ & ~new_n11335_;
  assign new_n11337_ = new_n1172_ & ~new_n11336_;
  assign new_n11338_ = new_n1176_ & ~new_n11337_;
  assign new_n11339_ = new_n1180_ & ~new_n11338_;
  assign new_n11340_ = new_n1184_ & ~new_n11339_;
  assign new_n11341_ = new_n1188_ & ~new_n11340_;
  assign new_n11342_ = new_n1192_ & ~new_n11341_;
  assign new_n11343_ = new_n1196_ & ~new_n11342_;
  assign new_n11344_ = new_n1200_ & ~new_n11343_;
  assign new_n11345_ = new_n1204_ & ~new_n11344_;
  assign new_n11346_ = new_n1208_ & ~new_n11345_;
  assign new_n11347_ = new_n1212_ & ~new_n11346_;
  assign new_n11348_ = new_n1216_ & ~new_n11347_;
  assign new_n11349_ = new_n1220_ & ~new_n11348_;
  assign new_n11350_ = new_n1224_ & ~new_n11349_;
  assign new_n11351_ = new_n1228_ & ~new_n11350_;
  assign new_n11352_ = new_n1232_ & ~new_n11351_;
  assign new_n11353_ = new_n1236_ & ~new_n11352_;
  assign new_n11354_ = new_n1240_ & ~new_n11353_;
  assign new_n11355_ = new_n1244_ & ~new_n11354_;
  assign new_n11356_ = new_n1248_ & ~new_n11355_;
  assign new_n11357_ = new_n1252_ & ~new_n11356_;
  assign new_n11358_ = new_n1256_ & ~new_n11357_;
  assign new_n11359_ = new_n1260_ & ~new_n11358_;
  assign new_n11360_ = new_n1264_ & ~new_n11359_;
  assign new_n11361_ = new_n1268_ & ~new_n11360_;
  assign new_n11362_ = new_n1272_ & ~new_n11361_;
  assign new_n11363_ = new_n1276_ & ~new_n11362_;
  assign new_n11364_ = new_n1280_ & ~new_n11363_;
  assign new_n11365_ = new_n1284_ & ~new_n11364_;
  assign new_n11366_ = new_n1288_ & ~new_n11365_;
  assign new_n11367_ = new_n1292_ & ~new_n11366_;
  assign new_n11368_ = new_n1296_ & ~new_n11367_;
  assign new_n11369_ = new_n1300_ & ~new_n11368_;
  assign new_n11370_ = new_n1304_ & ~new_n11369_;
  assign new_n11371_ = new_n1308_ & ~new_n11370_;
  assign new_n11372_ = new_n1312_ & ~new_n11371_;
  assign new_n11373_ = new_n1316_ & ~new_n11372_;
  assign new_n11374_ = new_n1320_ & ~new_n11373_;
  assign new_n11375_ = new_n1324_ & ~new_n11374_;
  assign new_n11376_ = new_n1328_ & ~new_n11375_;
  assign new_n11377_ = new_n1332_ & ~new_n11376_;
  assign new_n11378_ = new_n1336_ & ~new_n11377_;
  assign new_n11379_ = new_n1340_ & ~new_n11378_;
  assign new_n11380_ = new_n1344_ & ~new_n11379_;
  assign new_n11381_ = new_n1348_ & ~new_n11380_;
  assign new_n11382_ = new_n1352_ & ~new_n11381_;
  assign new_n11383_ = new_n1356_ & ~new_n11382_;
  assign new_n11384_ = new_n1360_ & ~new_n11383_;
  assign new_n11385_ = new_n1364_ & ~new_n11384_;
  assign new_n11386_ = \req[118]  & ~new_n1366_;
  assign \grant[118]  = ~new_n11385_ & new_n11386_;
  assign new_n11388_ = ~new_n703_ & new_n1375_;
  assign new_n11389_ = new_n1380_ & ~new_n11388_;
  assign new_n11390_ = new_n1384_ & ~new_n11389_;
  assign new_n11391_ = new_n1388_ & ~new_n11390_;
  assign new_n11392_ = new_n1392_ & ~new_n11391_;
  assign new_n11393_ = new_n1396_ & ~new_n11392_;
  assign new_n11394_ = new_n1663_ & ~new_n11393_;
  assign new_n11395_ = new_n392_ & ~new_n11394_;
  assign new_n11396_ = new_n396_ & ~new_n11395_;
  assign new_n11397_ = new_n400_ & ~new_n11396_;
  assign new_n11398_ = new_n404_ & ~new_n11397_;
  assign new_n11399_ = new_n408_ & ~new_n11398_;
  assign new_n11400_ = new_n412_ & ~new_n11399_;
  assign new_n11401_ = new_n416_ & ~new_n11400_;
  assign new_n11402_ = new_n420_ & ~new_n11401_;
  assign new_n11403_ = new_n424_ & ~new_n11402_;
  assign new_n11404_ = new_n428_ & ~new_n11403_;
  assign new_n11405_ = new_n432_ & ~new_n11404_;
  assign new_n11406_ = new_n436_ & ~new_n11405_;
  assign new_n11407_ = new_n440_ & ~new_n11406_;
  assign new_n11408_ = new_n444_ & ~new_n11407_;
  assign new_n11409_ = new_n448_ & ~new_n11408_;
  assign new_n11410_ = new_n452_ & ~new_n11409_;
  assign new_n11411_ = new_n456_ & ~new_n11410_;
  assign new_n11412_ = new_n460_ & ~new_n11411_;
  assign new_n11413_ = new_n464_ & ~new_n11412_;
  assign new_n11414_ = new_n468_ & ~new_n11413_;
  assign new_n11415_ = new_n472_ & ~new_n11414_;
  assign new_n11416_ = new_n476_ & ~new_n11415_;
  assign new_n11417_ = new_n480_ & ~new_n11416_;
  assign new_n11418_ = new_n484_ & ~new_n11417_;
  assign new_n11419_ = new_n488_ & ~new_n11418_;
  assign new_n11420_ = new_n492_ & ~new_n11419_;
  assign new_n11421_ = new_n496_ & ~new_n11420_;
  assign new_n11422_ = new_n500_ & ~new_n11421_;
  assign new_n11423_ = new_n504_ & ~new_n11422_;
  assign new_n11424_ = new_n508_ & ~new_n11423_;
  assign new_n11425_ = new_n512_ & ~new_n11424_;
  assign new_n11426_ = new_n516_ & ~new_n11425_;
  assign new_n11427_ = new_n520_ & ~new_n11426_;
  assign new_n11428_ = new_n524_ & ~new_n11427_;
  assign new_n11429_ = new_n528_ & ~new_n11428_;
  assign new_n11430_ = new_n532_ & ~new_n11429_;
  assign new_n11431_ = new_n536_ & ~new_n11430_;
  assign new_n11432_ = new_n540_ & ~new_n11431_;
  assign new_n11433_ = new_n544_ & ~new_n11432_;
  assign new_n11434_ = new_n548_ & ~new_n11433_;
  assign new_n11435_ = new_n552_ & ~new_n11434_;
  assign new_n11436_ = new_n556_ & ~new_n11435_;
  assign new_n11437_ = new_n560_ & ~new_n11436_;
  assign new_n11438_ = new_n564_ & ~new_n11437_;
  assign new_n11439_ = new_n568_ & ~new_n11438_;
  assign new_n11440_ = new_n572_ & ~new_n11439_;
  assign new_n11441_ = new_n576_ & ~new_n11440_;
  assign new_n11442_ = new_n580_ & ~new_n11441_;
  assign new_n11443_ = new_n584_ & ~new_n11442_;
  assign new_n11444_ = new_n588_ & ~new_n11443_;
  assign new_n11445_ = new_n592_ & ~new_n11444_;
  assign new_n11446_ = new_n596_ & ~new_n11445_;
  assign new_n11447_ = new_n600_ & ~new_n11446_;
  assign new_n11448_ = new_n604_ & ~new_n11447_;
  assign new_n11449_ = new_n608_ & ~new_n11448_;
  assign new_n11450_ = new_n612_ & ~new_n11449_;
  assign new_n11451_ = new_n616_ & ~new_n11450_;
  assign new_n11452_ = new_n620_ & ~new_n11451_;
  assign new_n11453_ = new_n624_ & ~new_n11452_;
  assign new_n11454_ = new_n628_ & ~new_n11453_;
  assign new_n11455_ = new_n632_ & ~new_n11454_;
  assign new_n11456_ = new_n636_ & ~new_n11455_;
  assign new_n11457_ = new_n640_ & ~new_n11456_;
  assign new_n11458_ = new_n644_ & ~new_n11457_;
  assign new_n11459_ = new_n648_ & ~new_n11458_;
  assign new_n11460_ = new_n652_ & ~new_n11459_;
  assign new_n11461_ = new_n656_ & ~new_n11460_;
  assign new_n11462_ = new_n660_ & ~new_n11461_;
  assign new_n11463_ = new_n664_ & ~new_n11462_;
  assign new_n11464_ = new_n668_ & ~new_n11463_;
  assign new_n11465_ = new_n672_ & ~new_n11464_;
  assign new_n11466_ = new_n676_ & ~new_n11465_;
  assign new_n11467_ = new_n680_ & ~new_n11466_;
  assign new_n11468_ = new_n684_ & ~new_n11467_;
  assign new_n11469_ = new_n688_ & ~new_n11468_;
  assign new_n11470_ = new_n692_ & ~new_n11469_;
  assign new_n11471_ = new_n696_ & ~new_n11470_;
  assign new_n11472_ = \req[119]  & ~new_n698_;
  assign \grant[119]  = ~new_n11471_ & new_n11472_;
  assign new_n11474_ = new_n707_ & ~new_n1042_;
  assign new_n11475_ = new_n712_ & ~new_n11474_;
  assign new_n11476_ = new_n716_ & ~new_n11475_;
  assign new_n11477_ = new_n720_ & ~new_n11476_;
  assign new_n11478_ = new_n1484_ & ~new_n11477_;
  assign new_n11479_ = new_n1486_ & ~new_n11478_;
  assign new_n11480_ = new_n1750_ & ~new_n11479_;
  assign new_n11481_ = new_n731_ & ~new_n11480_;
  assign new_n11482_ = new_n735_ & ~new_n11481_;
  assign new_n11483_ = new_n739_ & ~new_n11482_;
  assign new_n11484_ = new_n743_ & ~new_n11483_;
  assign new_n11485_ = new_n747_ & ~new_n11484_;
  assign new_n11486_ = new_n751_ & ~new_n11485_;
  assign new_n11487_ = new_n755_ & ~new_n11486_;
  assign new_n11488_ = new_n759_ & ~new_n11487_;
  assign new_n11489_ = new_n763_ & ~new_n11488_;
  assign new_n11490_ = new_n767_ & ~new_n11489_;
  assign new_n11491_ = new_n771_ & ~new_n11490_;
  assign new_n11492_ = new_n775_ & ~new_n11491_;
  assign new_n11493_ = new_n779_ & ~new_n11492_;
  assign new_n11494_ = new_n783_ & ~new_n11493_;
  assign new_n11495_ = new_n787_ & ~new_n11494_;
  assign new_n11496_ = new_n791_ & ~new_n11495_;
  assign new_n11497_ = new_n795_ & ~new_n11496_;
  assign new_n11498_ = new_n799_ & ~new_n11497_;
  assign new_n11499_ = new_n803_ & ~new_n11498_;
  assign new_n11500_ = new_n807_ & ~new_n11499_;
  assign new_n11501_ = new_n811_ & ~new_n11500_;
  assign new_n11502_ = new_n815_ & ~new_n11501_;
  assign new_n11503_ = new_n819_ & ~new_n11502_;
  assign new_n11504_ = new_n823_ & ~new_n11503_;
  assign new_n11505_ = new_n827_ & ~new_n11504_;
  assign new_n11506_ = new_n831_ & ~new_n11505_;
  assign new_n11507_ = new_n835_ & ~new_n11506_;
  assign new_n11508_ = new_n839_ & ~new_n11507_;
  assign new_n11509_ = new_n843_ & ~new_n11508_;
  assign new_n11510_ = new_n847_ & ~new_n11509_;
  assign new_n11511_ = new_n851_ & ~new_n11510_;
  assign new_n11512_ = new_n855_ & ~new_n11511_;
  assign new_n11513_ = new_n859_ & ~new_n11512_;
  assign new_n11514_ = new_n863_ & ~new_n11513_;
  assign new_n11515_ = new_n867_ & ~new_n11514_;
  assign new_n11516_ = new_n871_ & ~new_n11515_;
  assign new_n11517_ = new_n875_ & ~new_n11516_;
  assign new_n11518_ = new_n879_ & ~new_n11517_;
  assign new_n11519_ = new_n883_ & ~new_n11518_;
  assign new_n11520_ = new_n887_ & ~new_n11519_;
  assign new_n11521_ = new_n891_ & ~new_n11520_;
  assign new_n11522_ = new_n895_ & ~new_n11521_;
  assign new_n11523_ = new_n899_ & ~new_n11522_;
  assign new_n11524_ = new_n903_ & ~new_n11523_;
  assign new_n11525_ = new_n907_ & ~new_n11524_;
  assign new_n11526_ = new_n911_ & ~new_n11525_;
  assign new_n11527_ = new_n915_ & ~new_n11526_;
  assign new_n11528_ = new_n919_ & ~new_n11527_;
  assign new_n11529_ = new_n923_ & ~new_n11528_;
  assign new_n11530_ = new_n927_ & ~new_n11529_;
  assign new_n11531_ = new_n931_ & ~new_n11530_;
  assign new_n11532_ = new_n935_ & ~new_n11531_;
  assign new_n11533_ = new_n939_ & ~new_n11532_;
  assign new_n11534_ = new_n943_ & ~new_n11533_;
  assign new_n11535_ = new_n947_ & ~new_n11534_;
  assign new_n11536_ = new_n951_ & ~new_n11535_;
  assign new_n11537_ = new_n955_ & ~new_n11536_;
  assign new_n11538_ = new_n959_ & ~new_n11537_;
  assign new_n11539_ = new_n963_ & ~new_n11538_;
  assign new_n11540_ = new_n967_ & ~new_n11539_;
  assign new_n11541_ = new_n971_ & ~new_n11540_;
  assign new_n11542_ = new_n975_ & ~new_n11541_;
  assign new_n11543_ = new_n979_ & ~new_n11542_;
  assign new_n11544_ = new_n983_ & ~new_n11543_;
  assign new_n11545_ = new_n987_ & ~new_n11544_;
  assign new_n11546_ = new_n991_ & ~new_n11545_;
  assign new_n11547_ = new_n995_ & ~new_n11546_;
  assign new_n11548_ = new_n999_ & ~new_n11547_;
  assign new_n11549_ = new_n1003_ & ~new_n11548_;
  assign new_n11550_ = new_n1007_ & ~new_n11549_;
  assign new_n11551_ = new_n1011_ & ~new_n11550_;
  assign new_n11552_ = new_n1015_ & ~new_n11551_;
  assign new_n11553_ = new_n1019_ & ~new_n11552_;
  assign new_n11554_ = new_n1023_ & ~new_n11553_;
  assign new_n11555_ = new_n1027_ & ~new_n11554_;
  assign new_n11556_ = new_n1031_ & ~new_n11555_;
  assign new_n11557_ = new_n1035_ & ~new_n11556_;
  assign new_n11558_ = \req[120]  & ~new_n1037_;
  assign \grant[120]  = ~new_n11557_ & new_n11558_;
  assign new_n11560_ = new_n1046_ & ~new_n1379_;
  assign new_n11561_ = new_n1051_ & ~new_n11560_;
  assign new_n11562_ = new_n1055_ & ~new_n11561_;
  assign new_n11563_ = new_n1059_ & ~new_n11562_;
  assign new_n11564_ = new_n1574_ & ~new_n11563_;
  assign new_n11565_ = new_n1576_ & ~new_n11564_;
  assign new_n11566_ = new_n1837_ & ~new_n11565_;
  assign new_n11567_ = new_n1068_ & ~new_n11566_;
  assign new_n11568_ = new_n1072_ & ~new_n11567_;
  assign new_n11569_ = new_n1076_ & ~new_n11568_;
  assign new_n11570_ = new_n1080_ & ~new_n11569_;
  assign new_n11571_ = new_n1084_ & ~new_n11570_;
  assign new_n11572_ = new_n1088_ & ~new_n11571_;
  assign new_n11573_ = new_n1092_ & ~new_n11572_;
  assign new_n11574_ = new_n1096_ & ~new_n11573_;
  assign new_n11575_ = new_n1100_ & ~new_n11574_;
  assign new_n11576_ = new_n1104_ & ~new_n11575_;
  assign new_n11577_ = new_n1108_ & ~new_n11576_;
  assign new_n11578_ = new_n1112_ & ~new_n11577_;
  assign new_n11579_ = new_n1116_ & ~new_n11578_;
  assign new_n11580_ = new_n1120_ & ~new_n11579_;
  assign new_n11581_ = new_n1124_ & ~new_n11580_;
  assign new_n11582_ = new_n1128_ & ~new_n11581_;
  assign new_n11583_ = new_n1132_ & ~new_n11582_;
  assign new_n11584_ = new_n1136_ & ~new_n11583_;
  assign new_n11585_ = new_n1140_ & ~new_n11584_;
  assign new_n11586_ = new_n1144_ & ~new_n11585_;
  assign new_n11587_ = new_n1148_ & ~new_n11586_;
  assign new_n11588_ = new_n1152_ & ~new_n11587_;
  assign new_n11589_ = new_n1156_ & ~new_n11588_;
  assign new_n11590_ = new_n1160_ & ~new_n11589_;
  assign new_n11591_ = new_n1164_ & ~new_n11590_;
  assign new_n11592_ = new_n1168_ & ~new_n11591_;
  assign new_n11593_ = new_n1172_ & ~new_n11592_;
  assign new_n11594_ = new_n1176_ & ~new_n11593_;
  assign new_n11595_ = new_n1180_ & ~new_n11594_;
  assign new_n11596_ = new_n1184_ & ~new_n11595_;
  assign new_n11597_ = new_n1188_ & ~new_n11596_;
  assign new_n11598_ = new_n1192_ & ~new_n11597_;
  assign new_n11599_ = new_n1196_ & ~new_n11598_;
  assign new_n11600_ = new_n1200_ & ~new_n11599_;
  assign new_n11601_ = new_n1204_ & ~new_n11600_;
  assign new_n11602_ = new_n1208_ & ~new_n11601_;
  assign new_n11603_ = new_n1212_ & ~new_n11602_;
  assign new_n11604_ = new_n1216_ & ~new_n11603_;
  assign new_n11605_ = new_n1220_ & ~new_n11604_;
  assign new_n11606_ = new_n1224_ & ~new_n11605_;
  assign new_n11607_ = new_n1228_ & ~new_n11606_;
  assign new_n11608_ = new_n1232_ & ~new_n11607_;
  assign new_n11609_ = new_n1236_ & ~new_n11608_;
  assign new_n11610_ = new_n1240_ & ~new_n11609_;
  assign new_n11611_ = new_n1244_ & ~new_n11610_;
  assign new_n11612_ = new_n1248_ & ~new_n11611_;
  assign new_n11613_ = new_n1252_ & ~new_n11612_;
  assign new_n11614_ = new_n1256_ & ~new_n11613_;
  assign new_n11615_ = new_n1260_ & ~new_n11614_;
  assign new_n11616_ = new_n1264_ & ~new_n11615_;
  assign new_n11617_ = new_n1268_ & ~new_n11616_;
  assign new_n11618_ = new_n1272_ & ~new_n11617_;
  assign new_n11619_ = new_n1276_ & ~new_n11618_;
  assign new_n11620_ = new_n1280_ & ~new_n11619_;
  assign new_n11621_ = new_n1284_ & ~new_n11620_;
  assign new_n11622_ = new_n1288_ & ~new_n11621_;
  assign new_n11623_ = new_n1292_ & ~new_n11622_;
  assign new_n11624_ = new_n1296_ & ~new_n11623_;
  assign new_n11625_ = new_n1300_ & ~new_n11624_;
  assign new_n11626_ = new_n1304_ & ~new_n11625_;
  assign new_n11627_ = new_n1308_ & ~new_n11626_;
  assign new_n11628_ = new_n1312_ & ~new_n11627_;
  assign new_n11629_ = new_n1316_ & ~new_n11628_;
  assign new_n11630_ = new_n1320_ & ~new_n11629_;
  assign new_n11631_ = new_n1324_ & ~new_n11630_;
  assign new_n11632_ = new_n1328_ & ~new_n11631_;
  assign new_n11633_ = new_n1332_ & ~new_n11632_;
  assign new_n11634_ = new_n1336_ & ~new_n11633_;
  assign new_n11635_ = new_n1340_ & ~new_n11634_;
  assign new_n11636_ = new_n1344_ & ~new_n11635_;
  assign new_n11637_ = new_n1348_ & ~new_n11636_;
  assign new_n11638_ = new_n1352_ & ~new_n11637_;
  assign new_n11639_ = new_n1356_ & ~new_n11638_;
  assign new_n11640_ = new_n1360_ & ~new_n11639_;
  assign new_n11641_ = new_n1364_ & ~new_n11640_;
  assign new_n11642_ = new_n1368_ & ~new_n11641_;
  assign new_n11643_ = new_n1372_ & ~new_n11642_;
  assign new_n11644_ = \req[121]  & ~new_n1374_;
  assign \grant[121]  = ~new_n11643_ & new_n11644_;
  assign new_n11646_ = ~new_n711_ & new_n1383_;
  assign new_n11647_ = new_n1388_ & ~new_n11646_;
  assign new_n11648_ = new_n1392_ & ~new_n11647_;
  assign new_n11649_ = new_n1396_ & ~new_n11648_;
  assign new_n11650_ = new_n1663_ & ~new_n11649_;
  assign new_n11651_ = new_n392_ & ~new_n11650_;
  assign new_n11652_ = new_n396_ & ~new_n11651_;
  assign new_n11653_ = new_n400_ & ~new_n11652_;
  assign new_n11654_ = new_n404_ & ~new_n11653_;
  assign new_n11655_ = new_n408_ & ~new_n11654_;
  assign new_n11656_ = new_n412_ & ~new_n11655_;
  assign new_n11657_ = new_n416_ & ~new_n11656_;
  assign new_n11658_ = new_n420_ & ~new_n11657_;
  assign new_n11659_ = new_n424_ & ~new_n11658_;
  assign new_n11660_ = new_n428_ & ~new_n11659_;
  assign new_n11661_ = new_n432_ & ~new_n11660_;
  assign new_n11662_ = new_n436_ & ~new_n11661_;
  assign new_n11663_ = new_n440_ & ~new_n11662_;
  assign new_n11664_ = new_n444_ & ~new_n11663_;
  assign new_n11665_ = new_n448_ & ~new_n11664_;
  assign new_n11666_ = new_n452_ & ~new_n11665_;
  assign new_n11667_ = new_n456_ & ~new_n11666_;
  assign new_n11668_ = new_n460_ & ~new_n11667_;
  assign new_n11669_ = new_n464_ & ~new_n11668_;
  assign new_n11670_ = new_n468_ & ~new_n11669_;
  assign new_n11671_ = new_n472_ & ~new_n11670_;
  assign new_n11672_ = new_n476_ & ~new_n11671_;
  assign new_n11673_ = new_n480_ & ~new_n11672_;
  assign new_n11674_ = new_n484_ & ~new_n11673_;
  assign new_n11675_ = new_n488_ & ~new_n11674_;
  assign new_n11676_ = new_n492_ & ~new_n11675_;
  assign new_n11677_ = new_n496_ & ~new_n11676_;
  assign new_n11678_ = new_n500_ & ~new_n11677_;
  assign new_n11679_ = new_n504_ & ~new_n11678_;
  assign new_n11680_ = new_n508_ & ~new_n11679_;
  assign new_n11681_ = new_n512_ & ~new_n11680_;
  assign new_n11682_ = new_n516_ & ~new_n11681_;
  assign new_n11683_ = new_n520_ & ~new_n11682_;
  assign new_n11684_ = new_n524_ & ~new_n11683_;
  assign new_n11685_ = new_n528_ & ~new_n11684_;
  assign new_n11686_ = new_n532_ & ~new_n11685_;
  assign new_n11687_ = new_n536_ & ~new_n11686_;
  assign new_n11688_ = new_n540_ & ~new_n11687_;
  assign new_n11689_ = new_n544_ & ~new_n11688_;
  assign new_n11690_ = new_n548_ & ~new_n11689_;
  assign new_n11691_ = new_n552_ & ~new_n11690_;
  assign new_n11692_ = new_n556_ & ~new_n11691_;
  assign new_n11693_ = new_n560_ & ~new_n11692_;
  assign new_n11694_ = new_n564_ & ~new_n11693_;
  assign new_n11695_ = new_n568_ & ~new_n11694_;
  assign new_n11696_ = new_n572_ & ~new_n11695_;
  assign new_n11697_ = new_n576_ & ~new_n11696_;
  assign new_n11698_ = new_n580_ & ~new_n11697_;
  assign new_n11699_ = new_n584_ & ~new_n11698_;
  assign new_n11700_ = new_n588_ & ~new_n11699_;
  assign new_n11701_ = new_n592_ & ~new_n11700_;
  assign new_n11702_ = new_n596_ & ~new_n11701_;
  assign new_n11703_ = new_n600_ & ~new_n11702_;
  assign new_n11704_ = new_n604_ & ~new_n11703_;
  assign new_n11705_ = new_n608_ & ~new_n11704_;
  assign new_n11706_ = new_n612_ & ~new_n11705_;
  assign new_n11707_ = new_n616_ & ~new_n11706_;
  assign new_n11708_ = new_n620_ & ~new_n11707_;
  assign new_n11709_ = new_n624_ & ~new_n11708_;
  assign new_n11710_ = new_n628_ & ~new_n11709_;
  assign new_n11711_ = new_n632_ & ~new_n11710_;
  assign new_n11712_ = new_n636_ & ~new_n11711_;
  assign new_n11713_ = new_n640_ & ~new_n11712_;
  assign new_n11714_ = new_n644_ & ~new_n11713_;
  assign new_n11715_ = new_n648_ & ~new_n11714_;
  assign new_n11716_ = new_n652_ & ~new_n11715_;
  assign new_n11717_ = new_n656_ & ~new_n11716_;
  assign new_n11718_ = new_n660_ & ~new_n11717_;
  assign new_n11719_ = new_n664_ & ~new_n11718_;
  assign new_n11720_ = new_n668_ & ~new_n11719_;
  assign new_n11721_ = new_n672_ & ~new_n11720_;
  assign new_n11722_ = new_n676_ & ~new_n11721_;
  assign new_n11723_ = new_n680_ & ~new_n11722_;
  assign new_n11724_ = new_n684_ & ~new_n11723_;
  assign new_n11725_ = new_n688_ & ~new_n11724_;
  assign new_n11726_ = new_n692_ & ~new_n11725_;
  assign new_n11727_ = new_n696_ & ~new_n11726_;
  assign new_n11728_ = new_n700_ & ~new_n11727_;
  assign new_n11729_ = new_n704_ & ~new_n11728_;
  assign new_n11730_ = \req[122]  & ~new_n706_;
  assign \grant[122]  = ~new_n11729_ & new_n11730_;
  assign new_n11732_ = new_n715_ & ~new_n1050_;
  assign new_n11733_ = new_n720_ & ~new_n11732_;
  assign new_n11734_ = new_n1484_ & ~new_n11733_;
  assign new_n11735_ = new_n1486_ & ~new_n11734_;
  assign new_n11736_ = new_n1750_ & ~new_n11735_;
  assign new_n11737_ = new_n731_ & ~new_n11736_;
  assign new_n11738_ = new_n735_ & ~new_n11737_;
  assign new_n11739_ = new_n739_ & ~new_n11738_;
  assign new_n11740_ = new_n743_ & ~new_n11739_;
  assign new_n11741_ = new_n747_ & ~new_n11740_;
  assign new_n11742_ = new_n751_ & ~new_n11741_;
  assign new_n11743_ = new_n755_ & ~new_n11742_;
  assign new_n11744_ = new_n759_ & ~new_n11743_;
  assign new_n11745_ = new_n763_ & ~new_n11744_;
  assign new_n11746_ = new_n767_ & ~new_n11745_;
  assign new_n11747_ = new_n771_ & ~new_n11746_;
  assign new_n11748_ = new_n775_ & ~new_n11747_;
  assign new_n11749_ = new_n779_ & ~new_n11748_;
  assign new_n11750_ = new_n783_ & ~new_n11749_;
  assign new_n11751_ = new_n787_ & ~new_n11750_;
  assign new_n11752_ = new_n791_ & ~new_n11751_;
  assign new_n11753_ = new_n795_ & ~new_n11752_;
  assign new_n11754_ = new_n799_ & ~new_n11753_;
  assign new_n11755_ = new_n803_ & ~new_n11754_;
  assign new_n11756_ = new_n807_ & ~new_n11755_;
  assign new_n11757_ = new_n811_ & ~new_n11756_;
  assign new_n11758_ = new_n815_ & ~new_n11757_;
  assign new_n11759_ = new_n819_ & ~new_n11758_;
  assign new_n11760_ = new_n823_ & ~new_n11759_;
  assign new_n11761_ = new_n827_ & ~new_n11760_;
  assign new_n11762_ = new_n831_ & ~new_n11761_;
  assign new_n11763_ = new_n835_ & ~new_n11762_;
  assign new_n11764_ = new_n839_ & ~new_n11763_;
  assign new_n11765_ = new_n843_ & ~new_n11764_;
  assign new_n11766_ = new_n847_ & ~new_n11765_;
  assign new_n11767_ = new_n851_ & ~new_n11766_;
  assign new_n11768_ = new_n855_ & ~new_n11767_;
  assign new_n11769_ = new_n859_ & ~new_n11768_;
  assign new_n11770_ = new_n863_ & ~new_n11769_;
  assign new_n11771_ = new_n867_ & ~new_n11770_;
  assign new_n11772_ = new_n871_ & ~new_n11771_;
  assign new_n11773_ = new_n875_ & ~new_n11772_;
  assign new_n11774_ = new_n879_ & ~new_n11773_;
  assign new_n11775_ = new_n883_ & ~new_n11774_;
  assign new_n11776_ = new_n887_ & ~new_n11775_;
  assign new_n11777_ = new_n891_ & ~new_n11776_;
  assign new_n11778_ = new_n895_ & ~new_n11777_;
  assign new_n11779_ = new_n899_ & ~new_n11778_;
  assign new_n11780_ = new_n903_ & ~new_n11779_;
  assign new_n11781_ = new_n907_ & ~new_n11780_;
  assign new_n11782_ = new_n911_ & ~new_n11781_;
  assign new_n11783_ = new_n915_ & ~new_n11782_;
  assign new_n11784_ = new_n919_ & ~new_n11783_;
  assign new_n11785_ = new_n923_ & ~new_n11784_;
  assign new_n11786_ = new_n927_ & ~new_n11785_;
  assign new_n11787_ = new_n931_ & ~new_n11786_;
  assign new_n11788_ = new_n935_ & ~new_n11787_;
  assign new_n11789_ = new_n939_ & ~new_n11788_;
  assign new_n11790_ = new_n943_ & ~new_n11789_;
  assign new_n11791_ = new_n947_ & ~new_n11790_;
  assign new_n11792_ = new_n951_ & ~new_n11791_;
  assign new_n11793_ = new_n955_ & ~new_n11792_;
  assign new_n11794_ = new_n959_ & ~new_n11793_;
  assign new_n11795_ = new_n963_ & ~new_n11794_;
  assign new_n11796_ = new_n967_ & ~new_n11795_;
  assign new_n11797_ = new_n971_ & ~new_n11796_;
  assign new_n11798_ = new_n975_ & ~new_n11797_;
  assign new_n11799_ = new_n979_ & ~new_n11798_;
  assign new_n11800_ = new_n983_ & ~new_n11799_;
  assign new_n11801_ = new_n987_ & ~new_n11800_;
  assign new_n11802_ = new_n991_ & ~new_n11801_;
  assign new_n11803_ = new_n995_ & ~new_n11802_;
  assign new_n11804_ = new_n999_ & ~new_n11803_;
  assign new_n11805_ = new_n1003_ & ~new_n11804_;
  assign new_n11806_ = new_n1007_ & ~new_n11805_;
  assign new_n11807_ = new_n1011_ & ~new_n11806_;
  assign new_n11808_ = new_n1015_ & ~new_n11807_;
  assign new_n11809_ = new_n1019_ & ~new_n11808_;
  assign new_n11810_ = new_n1023_ & ~new_n11809_;
  assign new_n11811_ = new_n1027_ & ~new_n11810_;
  assign new_n11812_ = new_n1031_ & ~new_n11811_;
  assign new_n11813_ = new_n1035_ & ~new_n11812_;
  assign new_n11814_ = new_n1039_ & ~new_n11813_;
  assign new_n11815_ = new_n1043_ & ~new_n11814_;
  assign new_n11816_ = \req[123]  & ~new_n1045_;
  assign \grant[123]  = ~new_n11815_ & new_n11816_;
  assign new_n11818_ = new_n1054_ & ~new_n1387_;
  assign new_n11819_ = new_n1059_ & ~new_n11818_;
  assign new_n11820_ = new_n1574_ & ~new_n11819_;
  assign new_n11821_ = new_n1576_ & ~new_n11820_;
  assign new_n11822_ = new_n1837_ & ~new_n11821_;
  assign new_n11823_ = new_n1068_ & ~new_n11822_;
  assign new_n11824_ = new_n1072_ & ~new_n11823_;
  assign new_n11825_ = new_n1076_ & ~new_n11824_;
  assign new_n11826_ = new_n1080_ & ~new_n11825_;
  assign new_n11827_ = new_n1084_ & ~new_n11826_;
  assign new_n11828_ = new_n1088_ & ~new_n11827_;
  assign new_n11829_ = new_n1092_ & ~new_n11828_;
  assign new_n11830_ = new_n1096_ & ~new_n11829_;
  assign new_n11831_ = new_n1100_ & ~new_n11830_;
  assign new_n11832_ = new_n1104_ & ~new_n11831_;
  assign new_n11833_ = new_n1108_ & ~new_n11832_;
  assign new_n11834_ = new_n1112_ & ~new_n11833_;
  assign new_n11835_ = new_n1116_ & ~new_n11834_;
  assign new_n11836_ = new_n1120_ & ~new_n11835_;
  assign new_n11837_ = new_n1124_ & ~new_n11836_;
  assign new_n11838_ = new_n1128_ & ~new_n11837_;
  assign new_n11839_ = new_n1132_ & ~new_n11838_;
  assign new_n11840_ = new_n1136_ & ~new_n11839_;
  assign new_n11841_ = new_n1140_ & ~new_n11840_;
  assign new_n11842_ = new_n1144_ & ~new_n11841_;
  assign new_n11843_ = new_n1148_ & ~new_n11842_;
  assign new_n11844_ = new_n1152_ & ~new_n11843_;
  assign new_n11845_ = new_n1156_ & ~new_n11844_;
  assign new_n11846_ = new_n1160_ & ~new_n11845_;
  assign new_n11847_ = new_n1164_ & ~new_n11846_;
  assign new_n11848_ = new_n1168_ & ~new_n11847_;
  assign new_n11849_ = new_n1172_ & ~new_n11848_;
  assign new_n11850_ = new_n1176_ & ~new_n11849_;
  assign new_n11851_ = new_n1180_ & ~new_n11850_;
  assign new_n11852_ = new_n1184_ & ~new_n11851_;
  assign new_n11853_ = new_n1188_ & ~new_n11852_;
  assign new_n11854_ = new_n1192_ & ~new_n11853_;
  assign new_n11855_ = new_n1196_ & ~new_n11854_;
  assign new_n11856_ = new_n1200_ & ~new_n11855_;
  assign new_n11857_ = new_n1204_ & ~new_n11856_;
  assign new_n11858_ = new_n1208_ & ~new_n11857_;
  assign new_n11859_ = new_n1212_ & ~new_n11858_;
  assign new_n11860_ = new_n1216_ & ~new_n11859_;
  assign new_n11861_ = new_n1220_ & ~new_n11860_;
  assign new_n11862_ = new_n1224_ & ~new_n11861_;
  assign new_n11863_ = new_n1228_ & ~new_n11862_;
  assign new_n11864_ = new_n1232_ & ~new_n11863_;
  assign new_n11865_ = new_n1236_ & ~new_n11864_;
  assign new_n11866_ = new_n1240_ & ~new_n11865_;
  assign new_n11867_ = new_n1244_ & ~new_n11866_;
  assign new_n11868_ = new_n1248_ & ~new_n11867_;
  assign new_n11869_ = new_n1252_ & ~new_n11868_;
  assign new_n11870_ = new_n1256_ & ~new_n11869_;
  assign new_n11871_ = new_n1260_ & ~new_n11870_;
  assign new_n11872_ = new_n1264_ & ~new_n11871_;
  assign new_n11873_ = new_n1268_ & ~new_n11872_;
  assign new_n11874_ = new_n1272_ & ~new_n11873_;
  assign new_n11875_ = new_n1276_ & ~new_n11874_;
  assign new_n11876_ = new_n1280_ & ~new_n11875_;
  assign new_n11877_ = new_n1284_ & ~new_n11876_;
  assign new_n11878_ = new_n1288_ & ~new_n11877_;
  assign new_n11879_ = new_n1292_ & ~new_n11878_;
  assign new_n11880_ = new_n1296_ & ~new_n11879_;
  assign new_n11881_ = new_n1300_ & ~new_n11880_;
  assign new_n11882_ = new_n1304_ & ~new_n11881_;
  assign new_n11883_ = new_n1308_ & ~new_n11882_;
  assign new_n11884_ = new_n1312_ & ~new_n11883_;
  assign new_n11885_ = new_n1316_ & ~new_n11884_;
  assign new_n11886_ = new_n1320_ & ~new_n11885_;
  assign new_n11887_ = new_n1324_ & ~new_n11886_;
  assign new_n11888_ = new_n1328_ & ~new_n11887_;
  assign new_n11889_ = new_n1332_ & ~new_n11888_;
  assign new_n11890_ = new_n1336_ & ~new_n11889_;
  assign new_n11891_ = new_n1340_ & ~new_n11890_;
  assign new_n11892_ = new_n1344_ & ~new_n11891_;
  assign new_n11893_ = new_n1348_ & ~new_n11892_;
  assign new_n11894_ = new_n1352_ & ~new_n11893_;
  assign new_n11895_ = new_n1356_ & ~new_n11894_;
  assign new_n11896_ = new_n1360_ & ~new_n11895_;
  assign new_n11897_ = new_n1364_ & ~new_n11896_;
  assign new_n11898_ = new_n1368_ & ~new_n11897_;
  assign new_n11899_ = new_n1372_ & ~new_n11898_;
  assign new_n11900_ = new_n1376_ & ~new_n11899_;
  assign new_n11901_ = new_n1380_ & ~new_n11900_;
  assign new_n11902_ = \req[124]  & ~new_n1382_;
  assign \grant[124]  = ~new_n11901_ & new_n11902_;
  assign new_n11904_ = ~new_n719_ & new_n1391_;
  assign new_n11905_ = new_n1396_ & ~new_n11904_;
  assign new_n11906_ = new_n1663_ & ~new_n11905_;
  assign new_n11907_ = new_n392_ & ~new_n11906_;
  assign new_n11908_ = new_n396_ & ~new_n11907_;
  assign new_n11909_ = new_n400_ & ~new_n11908_;
  assign new_n11910_ = new_n404_ & ~new_n11909_;
  assign new_n11911_ = new_n408_ & ~new_n11910_;
  assign new_n11912_ = new_n412_ & ~new_n11911_;
  assign new_n11913_ = new_n416_ & ~new_n11912_;
  assign new_n11914_ = new_n420_ & ~new_n11913_;
  assign new_n11915_ = new_n424_ & ~new_n11914_;
  assign new_n11916_ = new_n428_ & ~new_n11915_;
  assign new_n11917_ = new_n432_ & ~new_n11916_;
  assign new_n11918_ = new_n436_ & ~new_n11917_;
  assign new_n11919_ = new_n440_ & ~new_n11918_;
  assign new_n11920_ = new_n444_ & ~new_n11919_;
  assign new_n11921_ = new_n448_ & ~new_n11920_;
  assign new_n11922_ = new_n452_ & ~new_n11921_;
  assign new_n11923_ = new_n456_ & ~new_n11922_;
  assign new_n11924_ = new_n460_ & ~new_n11923_;
  assign new_n11925_ = new_n464_ & ~new_n11924_;
  assign new_n11926_ = new_n468_ & ~new_n11925_;
  assign new_n11927_ = new_n472_ & ~new_n11926_;
  assign new_n11928_ = new_n476_ & ~new_n11927_;
  assign new_n11929_ = new_n480_ & ~new_n11928_;
  assign new_n11930_ = new_n484_ & ~new_n11929_;
  assign new_n11931_ = new_n488_ & ~new_n11930_;
  assign new_n11932_ = new_n492_ & ~new_n11931_;
  assign new_n11933_ = new_n496_ & ~new_n11932_;
  assign new_n11934_ = new_n500_ & ~new_n11933_;
  assign new_n11935_ = new_n504_ & ~new_n11934_;
  assign new_n11936_ = new_n508_ & ~new_n11935_;
  assign new_n11937_ = new_n512_ & ~new_n11936_;
  assign new_n11938_ = new_n516_ & ~new_n11937_;
  assign new_n11939_ = new_n520_ & ~new_n11938_;
  assign new_n11940_ = new_n524_ & ~new_n11939_;
  assign new_n11941_ = new_n528_ & ~new_n11940_;
  assign new_n11942_ = new_n532_ & ~new_n11941_;
  assign new_n11943_ = new_n536_ & ~new_n11942_;
  assign new_n11944_ = new_n540_ & ~new_n11943_;
  assign new_n11945_ = new_n544_ & ~new_n11944_;
  assign new_n11946_ = new_n548_ & ~new_n11945_;
  assign new_n11947_ = new_n552_ & ~new_n11946_;
  assign new_n11948_ = new_n556_ & ~new_n11947_;
  assign new_n11949_ = new_n560_ & ~new_n11948_;
  assign new_n11950_ = new_n564_ & ~new_n11949_;
  assign new_n11951_ = new_n568_ & ~new_n11950_;
  assign new_n11952_ = new_n572_ & ~new_n11951_;
  assign new_n11953_ = new_n576_ & ~new_n11952_;
  assign new_n11954_ = new_n580_ & ~new_n11953_;
  assign new_n11955_ = new_n584_ & ~new_n11954_;
  assign new_n11956_ = new_n588_ & ~new_n11955_;
  assign new_n11957_ = new_n592_ & ~new_n11956_;
  assign new_n11958_ = new_n596_ & ~new_n11957_;
  assign new_n11959_ = new_n600_ & ~new_n11958_;
  assign new_n11960_ = new_n604_ & ~new_n11959_;
  assign new_n11961_ = new_n608_ & ~new_n11960_;
  assign new_n11962_ = new_n612_ & ~new_n11961_;
  assign new_n11963_ = new_n616_ & ~new_n11962_;
  assign new_n11964_ = new_n620_ & ~new_n11963_;
  assign new_n11965_ = new_n624_ & ~new_n11964_;
  assign new_n11966_ = new_n628_ & ~new_n11965_;
  assign new_n11967_ = new_n632_ & ~new_n11966_;
  assign new_n11968_ = new_n636_ & ~new_n11967_;
  assign new_n11969_ = new_n640_ & ~new_n11968_;
  assign new_n11970_ = new_n644_ & ~new_n11969_;
  assign new_n11971_ = new_n648_ & ~new_n11970_;
  assign new_n11972_ = new_n652_ & ~new_n11971_;
  assign new_n11973_ = new_n656_ & ~new_n11972_;
  assign new_n11974_ = new_n660_ & ~new_n11973_;
  assign new_n11975_ = new_n664_ & ~new_n11974_;
  assign new_n11976_ = new_n668_ & ~new_n11975_;
  assign new_n11977_ = new_n672_ & ~new_n11976_;
  assign new_n11978_ = new_n676_ & ~new_n11977_;
  assign new_n11979_ = new_n680_ & ~new_n11978_;
  assign new_n11980_ = new_n684_ & ~new_n11979_;
  assign new_n11981_ = new_n688_ & ~new_n11980_;
  assign new_n11982_ = new_n692_ & ~new_n11981_;
  assign new_n11983_ = new_n696_ & ~new_n11982_;
  assign new_n11984_ = new_n700_ & ~new_n11983_;
  assign new_n11985_ = new_n704_ & ~new_n11984_;
  assign new_n11986_ = new_n708_ & ~new_n11985_;
  assign new_n11987_ = new_n712_ & ~new_n11986_;
  assign new_n11988_ = \req[125]  & ~new_n714_;
  assign \grant[125]  = ~new_n11987_ & new_n11988_;
  assign new_n11990_ = ~new_n1058_ & new_n1483_;
  assign new_n11991_ = new_n1486_ & ~new_n11990_;
  assign new_n11992_ = new_n1750_ & ~new_n11991_;
  assign new_n11993_ = new_n731_ & ~new_n11992_;
  assign new_n11994_ = new_n735_ & ~new_n11993_;
  assign new_n11995_ = new_n739_ & ~new_n11994_;
  assign new_n11996_ = new_n743_ & ~new_n11995_;
  assign new_n11997_ = new_n747_ & ~new_n11996_;
  assign new_n11998_ = new_n751_ & ~new_n11997_;
  assign new_n11999_ = new_n755_ & ~new_n11998_;
  assign new_n12000_ = new_n759_ & ~new_n11999_;
  assign new_n12001_ = new_n763_ & ~new_n12000_;
  assign new_n12002_ = new_n767_ & ~new_n12001_;
  assign new_n12003_ = new_n771_ & ~new_n12002_;
  assign new_n12004_ = new_n775_ & ~new_n12003_;
  assign new_n12005_ = new_n779_ & ~new_n12004_;
  assign new_n12006_ = new_n783_ & ~new_n12005_;
  assign new_n12007_ = new_n787_ & ~new_n12006_;
  assign new_n12008_ = new_n791_ & ~new_n12007_;
  assign new_n12009_ = new_n795_ & ~new_n12008_;
  assign new_n12010_ = new_n799_ & ~new_n12009_;
  assign new_n12011_ = new_n803_ & ~new_n12010_;
  assign new_n12012_ = new_n807_ & ~new_n12011_;
  assign new_n12013_ = new_n811_ & ~new_n12012_;
  assign new_n12014_ = new_n815_ & ~new_n12013_;
  assign new_n12015_ = new_n819_ & ~new_n12014_;
  assign new_n12016_ = new_n823_ & ~new_n12015_;
  assign new_n12017_ = new_n827_ & ~new_n12016_;
  assign new_n12018_ = new_n831_ & ~new_n12017_;
  assign new_n12019_ = new_n835_ & ~new_n12018_;
  assign new_n12020_ = new_n839_ & ~new_n12019_;
  assign new_n12021_ = new_n843_ & ~new_n12020_;
  assign new_n12022_ = new_n847_ & ~new_n12021_;
  assign new_n12023_ = new_n851_ & ~new_n12022_;
  assign new_n12024_ = new_n855_ & ~new_n12023_;
  assign new_n12025_ = new_n859_ & ~new_n12024_;
  assign new_n12026_ = new_n863_ & ~new_n12025_;
  assign new_n12027_ = new_n867_ & ~new_n12026_;
  assign new_n12028_ = new_n871_ & ~new_n12027_;
  assign new_n12029_ = new_n875_ & ~new_n12028_;
  assign new_n12030_ = new_n879_ & ~new_n12029_;
  assign new_n12031_ = new_n883_ & ~new_n12030_;
  assign new_n12032_ = new_n887_ & ~new_n12031_;
  assign new_n12033_ = new_n891_ & ~new_n12032_;
  assign new_n12034_ = new_n895_ & ~new_n12033_;
  assign new_n12035_ = new_n899_ & ~new_n12034_;
  assign new_n12036_ = new_n903_ & ~new_n12035_;
  assign new_n12037_ = new_n907_ & ~new_n12036_;
  assign new_n12038_ = new_n911_ & ~new_n12037_;
  assign new_n12039_ = new_n915_ & ~new_n12038_;
  assign new_n12040_ = new_n919_ & ~new_n12039_;
  assign new_n12041_ = new_n923_ & ~new_n12040_;
  assign new_n12042_ = new_n927_ & ~new_n12041_;
  assign new_n12043_ = new_n931_ & ~new_n12042_;
  assign new_n12044_ = new_n935_ & ~new_n12043_;
  assign new_n12045_ = new_n939_ & ~new_n12044_;
  assign new_n12046_ = new_n943_ & ~new_n12045_;
  assign new_n12047_ = new_n947_ & ~new_n12046_;
  assign new_n12048_ = new_n951_ & ~new_n12047_;
  assign new_n12049_ = new_n955_ & ~new_n12048_;
  assign new_n12050_ = new_n959_ & ~new_n12049_;
  assign new_n12051_ = new_n963_ & ~new_n12050_;
  assign new_n12052_ = new_n967_ & ~new_n12051_;
  assign new_n12053_ = new_n971_ & ~new_n12052_;
  assign new_n12054_ = new_n975_ & ~new_n12053_;
  assign new_n12055_ = new_n979_ & ~new_n12054_;
  assign new_n12056_ = new_n983_ & ~new_n12055_;
  assign new_n12057_ = new_n987_ & ~new_n12056_;
  assign new_n12058_ = new_n991_ & ~new_n12057_;
  assign new_n12059_ = new_n995_ & ~new_n12058_;
  assign new_n12060_ = new_n999_ & ~new_n12059_;
  assign new_n12061_ = new_n1003_ & ~new_n12060_;
  assign new_n12062_ = new_n1007_ & ~new_n12061_;
  assign new_n12063_ = new_n1011_ & ~new_n12062_;
  assign new_n12064_ = new_n1015_ & ~new_n12063_;
  assign new_n12065_ = new_n1019_ & ~new_n12064_;
  assign new_n12066_ = new_n1023_ & ~new_n12065_;
  assign new_n12067_ = new_n1027_ & ~new_n12066_;
  assign new_n12068_ = new_n1031_ & ~new_n12067_;
  assign new_n12069_ = new_n1035_ & ~new_n12068_;
  assign new_n12070_ = new_n1039_ & ~new_n12069_;
  assign new_n12071_ = new_n1043_ & ~new_n12070_;
  assign new_n12072_ = new_n1047_ & ~new_n12071_;
  assign new_n12073_ = new_n1051_ & ~new_n12072_;
  assign new_n12074_ = \req[126]  & ~new_n1053_;
  assign \grant[126]  = ~new_n12073_ & new_n12074_;
  assign new_n12076_ = ~new_n1395_ & new_n1573_;
  assign new_n12077_ = new_n1576_ & ~new_n12076_;
  assign new_n12078_ = new_n1837_ & ~new_n12077_;
  assign new_n12079_ = new_n1068_ & ~new_n12078_;
  assign new_n12080_ = new_n1072_ & ~new_n12079_;
  assign new_n12081_ = new_n1076_ & ~new_n12080_;
  assign new_n12082_ = new_n1080_ & ~new_n12081_;
  assign new_n12083_ = new_n1084_ & ~new_n12082_;
  assign new_n12084_ = new_n1088_ & ~new_n12083_;
  assign new_n12085_ = new_n1092_ & ~new_n12084_;
  assign new_n12086_ = new_n1096_ & ~new_n12085_;
  assign new_n12087_ = new_n1100_ & ~new_n12086_;
  assign new_n12088_ = new_n1104_ & ~new_n12087_;
  assign new_n12089_ = new_n1108_ & ~new_n12088_;
  assign new_n12090_ = new_n1112_ & ~new_n12089_;
  assign new_n12091_ = new_n1116_ & ~new_n12090_;
  assign new_n12092_ = new_n1120_ & ~new_n12091_;
  assign new_n12093_ = new_n1124_ & ~new_n12092_;
  assign new_n12094_ = new_n1128_ & ~new_n12093_;
  assign new_n12095_ = new_n1132_ & ~new_n12094_;
  assign new_n12096_ = new_n1136_ & ~new_n12095_;
  assign new_n12097_ = new_n1140_ & ~new_n12096_;
  assign new_n12098_ = new_n1144_ & ~new_n12097_;
  assign new_n12099_ = new_n1148_ & ~new_n12098_;
  assign new_n12100_ = new_n1152_ & ~new_n12099_;
  assign new_n12101_ = new_n1156_ & ~new_n12100_;
  assign new_n12102_ = new_n1160_ & ~new_n12101_;
  assign new_n12103_ = new_n1164_ & ~new_n12102_;
  assign new_n12104_ = new_n1168_ & ~new_n12103_;
  assign new_n12105_ = new_n1172_ & ~new_n12104_;
  assign new_n12106_ = new_n1176_ & ~new_n12105_;
  assign new_n12107_ = new_n1180_ & ~new_n12106_;
  assign new_n12108_ = new_n1184_ & ~new_n12107_;
  assign new_n12109_ = new_n1188_ & ~new_n12108_;
  assign new_n12110_ = new_n1192_ & ~new_n12109_;
  assign new_n12111_ = new_n1196_ & ~new_n12110_;
  assign new_n12112_ = new_n1200_ & ~new_n12111_;
  assign new_n12113_ = new_n1204_ & ~new_n12112_;
  assign new_n12114_ = new_n1208_ & ~new_n12113_;
  assign new_n12115_ = new_n1212_ & ~new_n12114_;
  assign new_n12116_ = new_n1216_ & ~new_n12115_;
  assign new_n12117_ = new_n1220_ & ~new_n12116_;
  assign new_n12118_ = new_n1224_ & ~new_n12117_;
  assign new_n12119_ = new_n1228_ & ~new_n12118_;
  assign new_n12120_ = new_n1232_ & ~new_n12119_;
  assign new_n12121_ = new_n1236_ & ~new_n12120_;
  assign new_n12122_ = new_n1240_ & ~new_n12121_;
  assign new_n12123_ = new_n1244_ & ~new_n12122_;
  assign new_n12124_ = new_n1248_ & ~new_n12123_;
  assign new_n12125_ = new_n1252_ & ~new_n12124_;
  assign new_n12126_ = new_n1256_ & ~new_n12125_;
  assign new_n12127_ = new_n1260_ & ~new_n12126_;
  assign new_n12128_ = new_n1264_ & ~new_n12127_;
  assign new_n12129_ = new_n1268_ & ~new_n12128_;
  assign new_n12130_ = new_n1272_ & ~new_n12129_;
  assign new_n12131_ = new_n1276_ & ~new_n12130_;
  assign new_n12132_ = new_n1280_ & ~new_n12131_;
  assign new_n12133_ = new_n1284_ & ~new_n12132_;
  assign new_n12134_ = new_n1288_ & ~new_n12133_;
  assign new_n12135_ = new_n1292_ & ~new_n12134_;
  assign new_n12136_ = new_n1296_ & ~new_n12135_;
  assign new_n12137_ = new_n1300_ & ~new_n12136_;
  assign new_n12138_ = new_n1304_ & ~new_n12137_;
  assign new_n12139_ = new_n1308_ & ~new_n12138_;
  assign new_n12140_ = new_n1312_ & ~new_n12139_;
  assign new_n12141_ = new_n1316_ & ~new_n12140_;
  assign new_n12142_ = new_n1320_ & ~new_n12141_;
  assign new_n12143_ = new_n1324_ & ~new_n12142_;
  assign new_n12144_ = new_n1328_ & ~new_n12143_;
  assign new_n12145_ = new_n1332_ & ~new_n12144_;
  assign new_n12146_ = new_n1336_ & ~new_n12145_;
  assign new_n12147_ = new_n1340_ & ~new_n12146_;
  assign new_n12148_ = new_n1344_ & ~new_n12147_;
  assign new_n12149_ = new_n1348_ & ~new_n12148_;
  assign new_n12150_ = new_n1352_ & ~new_n12149_;
  assign new_n12151_ = new_n1356_ & ~new_n12150_;
  assign new_n12152_ = new_n1360_ & ~new_n12151_;
  assign new_n12153_ = new_n1364_ & ~new_n12152_;
  assign new_n12154_ = new_n1368_ & ~new_n12153_;
  assign new_n12155_ = new_n1372_ & ~new_n12154_;
  assign new_n12156_ = new_n1376_ & ~new_n12155_;
  assign new_n12157_ = new_n1380_ & ~new_n12156_;
  assign new_n12158_ = new_n1384_ & ~new_n12157_;
  assign new_n12159_ = new_n1388_ & ~new_n12158_;
  assign new_n12160_ = \req[127]  & ~new_n1390_;
  assign \grant[127]  = ~new_n12159_ & new_n12160_;
  assign new_n12162_ = new_n388_ & new_n403_;
  assign new_n12163_ = new_n419_ & new_n435_;
  assign new_n12164_ = new_n451_ & new_n467_;
  assign new_n12165_ = new_n483_ & new_n499_;
  assign new_n12166_ = new_n515_ & new_n531_;
  assign new_n12167_ = new_n547_ & new_n563_;
  assign new_n12168_ = new_n579_ & new_n595_;
  assign new_n12169_ = new_n611_ & new_n627_;
  assign new_n12170_ = new_n643_ & new_n659_;
  assign new_n12171_ = new_n675_ & new_n691_;
  assign new_n12172_ = new_n707_ & new_n734_;
  assign new_n12173_ = new_n750_ & new_n766_;
  assign new_n12174_ = new_n782_ & new_n798_;
  assign new_n12175_ = new_n814_ & new_n830_;
  assign new_n12176_ = new_n846_ & new_n862_;
  assign new_n12177_ = new_n878_ & new_n894_;
  assign new_n12178_ = new_n910_ & new_n926_;
  assign new_n12179_ = new_n942_ & new_n958_;
  assign new_n12180_ = new_n974_ & new_n990_;
  assign new_n12181_ = new_n1006_ & new_n1022_;
  assign new_n12182_ = new_n1038_ & new_n1054_;
  assign new_n12183_ = new_n1064_ & new_n1079_;
  assign new_n12184_ = new_n1095_ & new_n1111_;
  assign new_n12185_ = new_n1127_ & new_n1143_;
  assign new_n12186_ = new_n1159_ & new_n1175_;
  assign new_n12187_ = new_n1191_ & new_n1207_;
  assign new_n12188_ = new_n1223_ & new_n1239_;
  assign new_n12189_ = new_n1255_ & new_n1271_;
  assign new_n12190_ = new_n1287_ & new_n1303_;
  assign new_n12191_ = new_n1319_ & new_n1335_;
  assign new_n12192_ = new_n1351_ & new_n1367_;
  assign new_n12193_ = new_n1383_ & new_n1483_;
  assign new_n12194_ = new_n12192_ & new_n12193_;
  assign new_n12195_ = new_n12190_ & new_n12191_;
  assign new_n12196_ = new_n12188_ & new_n12189_;
  assign new_n12197_ = new_n12186_ & new_n12187_;
  assign new_n12198_ = new_n12184_ & new_n12185_;
  assign new_n12199_ = new_n12182_ & new_n12183_;
  assign new_n12200_ = new_n12180_ & new_n12181_;
  assign new_n12201_ = new_n12178_ & new_n12179_;
  assign new_n12202_ = new_n12176_ & new_n12177_;
  assign new_n12203_ = new_n12174_ & new_n12175_;
  assign new_n12204_ = new_n12172_ & new_n12173_;
  assign new_n12205_ = new_n12170_ & new_n12171_;
  assign new_n12206_ = new_n12168_ & new_n12169_;
  assign new_n12207_ = new_n12166_ & new_n12167_;
  assign new_n12208_ = new_n12164_ & new_n12165_;
  assign new_n12209_ = new_n12162_ & new_n12163_;
  assign new_n12210_ = new_n12208_ & new_n12209_;
  assign new_n12211_ = new_n12206_ & new_n12207_;
  assign new_n12212_ = new_n12204_ & new_n12205_;
  assign new_n12213_ = new_n12202_ & new_n12203_;
  assign new_n12214_ = new_n12200_ & new_n12201_;
  assign new_n12215_ = new_n12198_ & new_n12199_;
  assign new_n12216_ = new_n12196_ & new_n12197_;
  assign new_n12217_ = new_n12194_ & new_n12195_;
  assign new_n12218_ = new_n12216_ & new_n12217_;
  assign new_n12219_ = new_n12214_ & new_n12215_;
  assign new_n12220_ = new_n12212_ & new_n12213_;
  assign new_n12221_ = new_n12210_ & new_n12211_;
  assign new_n12222_ = new_n12220_ & new_n12221_;
  assign new_n12223_ = new_n12218_ & new_n12219_;
  assign anyGrant = ~new_n12222_ | ~new_n12223_;
endmodule


