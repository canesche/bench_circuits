module MinMax30 ( clock, 
    \1 , 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19,
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33,
    124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137,
    138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151,
    152, 153  );
  input  clock;
  input  \1 , 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18,
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33;
  output 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137,
    138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151,
    152, 153;
  reg 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50,
    51, 52, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68,
    69, 70, 71, 72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86,
    87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103,
    104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117,
    118, 119, 120, 121, 122, 123;
  wire new_n334_, new_n335_, new_n336_, new_n337_, new_n338_1_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_1_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_1_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_1_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_1_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_1_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_1_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_1_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_1_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_1_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_1_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_1_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_1_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_1_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_1_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_1_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_1_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_1_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_1_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_1_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_1_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_1_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_1_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_1_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_1_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_1_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_1_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_1_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_1_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_1_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_1_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_1_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_1_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_1_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_1_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_1_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_1_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_1_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_1_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_1_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_1_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_1_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_1_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_1_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_1_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_1_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_1_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_1_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1464_, new_n1466_, new_n1468_, new_n1470_,
    new_n1472_, new_n1474_, new_n1476_, new_n1478_, new_n1480_, new_n1482_,
    new_n1484_, new_n1486_, new_n1488_, new_n1490_, new_n1492_, new_n1494_,
    new_n1496_, new_n1498_, new_n1500_, new_n1502_, new_n1504_, new_n1506_,
    new_n1508_, new_n1510_, new_n1512_, new_n1514_, new_n1516_, new_n1518_,
    new_n1520_, new_n1522_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1584_, new_n1585_,
    new_n1586_, new_n1587_, new_n1588_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1656_, new_n1657_,
    new_n1658_, new_n1659_, new_n1660_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1704_, new_n1705_, new_n1707_, new_n1708_,
    new_n1710_, new_n1711_, new_n1713_, new_n1714_, new_n1716_, new_n1717_,
    new_n1719_, new_n1720_, new_n1722_, new_n1723_, new_n1725_, new_n1726_,
    new_n1728_, new_n1729_, new_n1731_, new_n1732_, new_n1734_, new_n1735_,
    new_n1737_, new_n1738_, new_n1740_, new_n1741_, new_n1743_, new_n1744_,
    new_n1746_, new_n1747_, new_n1749_, new_n1750_, new_n1752_, new_n1753_,
    new_n1755_, new_n1756_, new_n1758_, new_n1759_, new_n1761_, new_n1762_,
    new_n1764_, new_n1765_, new_n1767_, new_n1768_, new_n1770_, new_n1771_,
    new_n1773_, new_n1774_, new_n1776_, new_n1777_, new_n1779_, new_n1780_,
    new_n1782_, new_n1783_, new_n1785_, new_n1786_, new_n1788_, new_n1789_,
    new_n1791_, new_n1792_, n128, n133, n138, n143, n148, n153, n158, n163,
    n168, n173, n178, n183, n188, n193, n198, n203, n208, n213, n218, n223,
    n228, n233, n238, n243, n248, n253, n258, n263, n268, n273, n278, n283,
    n288, n293, n298, n303, n308, n313, n318, n323, n328, n333, n338, n343,
    n348, n353, n358, n363, n368, n373, n378, n383, n388, n393, n398, n403,
    n408, n413, n418, n423, n428, n433, n438, n443, n448, n453, n458, n463,
    n468, n473, n478, n483, n488, n493, n498, n503, n508, n513, n518, n523,
    n528, n533, n538, n543, n548, n553, n558, n563, n568, n573;
  assign new_n334_ = 33 & ~123;
  assign new_n335_ = ~33 & 123;
  assign new_n336_ = ~new_n334_ & ~new_n335_;
  assign new_n337_ = 32 & ~122;
  assign new_n338_1_ = ~32 & 122;
  assign new_n339_ = ~new_n337_ & ~new_n338_1_;
  assign new_n340_ = 31 & ~121;
  assign new_n341_ = ~31 & 121;
  assign new_n342_ = ~new_n340_ & ~new_n341_;
  assign new_n343_1_ = 30 & ~120;
  assign new_n344_ = ~30 & 120;
  assign new_n345_ = ~new_n343_1_ & ~new_n344_;
  assign new_n346_ = 29 & ~119;
  assign new_n347_ = ~29 & 119;
  assign new_n348_1_ = ~new_n346_ & ~new_n347_;
  assign new_n349_ = 28 & ~118;
  assign new_n350_ = ~28 & 118;
  assign new_n351_ = ~new_n349_ & ~new_n350_;
  assign new_n352_ = 27 & ~117;
  assign new_n353_1_ = ~27 & 117;
  assign new_n354_ = ~new_n352_ & ~new_n353_1_;
  assign new_n355_ = 26 & ~116;
  assign new_n356_ = ~26 & 116;
  assign new_n357_ = ~new_n355_ & ~new_n356_;
  assign new_n358_1_ = 25 & ~115;
  assign new_n359_ = ~25 & 115;
  assign new_n360_ = ~new_n358_1_ & ~new_n359_;
  assign new_n361_ = 24 & ~114;
  assign new_n362_ = ~24 & 114;
  assign new_n363_1_ = ~new_n361_ & ~new_n362_;
  assign new_n364_ = 23 & ~113;
  assign new_n365_ = ~23 & 113;
  assign new_n366_ = ~new_n364_ & ~new_n365_;
  assign new_n367_ = 22 & ~112;
  assign new_n368_1_ = ~22 & 112;
  assign new_n369_ = ~new_n367_ & ~new_n368_1_;
  assign new_n370_ = 21 & ~111;
  assign new_n371_ = ~21 & 111;
  assign new_n372_ = ~new_n370_ & ~new_n371_;
  assign new_n373_1_ = 20 & ~110;
  assign new_n374_ = ~20 & 110;
  assign new_n375_ = ~new_n373_1_ & ~new_n374_;
  assign new_n376_ = 19 & ~109;
  assign new_n377_ = ~19 & 109;
  assign new_n378_1_ = ~new_n376_ & ~new_n377_;
  assign new_n379_ = 18 & ~108;
  assign new_n380_ = ~18 & 108;
  assign new_n381_ = ~new_n379_ & ~new_n380_;
  assign new_n382_ = 17 & ~107;
  assign new_n383_1_ = ~17 & 107;
  assign new_n384_ = ~new_n382_ & ~new_n383_1_;
  assign new_n385_ = 16 & ~106;
  assign new_n386_ = ~16 & 106;
  assign new_n387_ = ~new_n385_ & ~new_n386_;
  assign new_n388_1_ = 15 & ~105;
  assign new_n389_ = ~15 & 105;
  assign new_n390_ = ~new_n388_1_ & ~new_n389_;
  assign new_n391_ = 14 & ~104;
  assign new_n392_ = ~14 & 104;
  assign new_n393_1_ = ~new_n391_ & ~new_n392_;
  assign new_n394_ = 13 & ~103;
  assign new_n395_ = ~13 & 103;
  assign new_n396_ = ~new_n394_ & ~new_n395_;
  assign new_n397_ = 12 & ~102;
  assign new_n398_1_ = ~12 & 102;
  assign new_n399_ = ~new_n397_ & ~new_n398_1_;
  assign new_n400_ = 11 & ~101;
  assign new_n401_ = ~11 & 101;
  assign new_n402_ = ~new_n400_ & ~new_n401_;
  assign new_n403_1_ = 10 & ~100;
  assign new_n404_ = ~10 & 100;
  assign new_n405_ = ~new_n403_1_ & ~new_n404_;
  assign new_n406_ = 9 & ~99;
  assign new_n407_ = ~9 & 99;
  assign new_n408_1_ = ~new_n406_ & ~new_n407_;
  assign new_n409_ = 8 & ~98;
  assign new_n410_ = ~8 & 98;
  assign new_n411_ = ~new_n409_ & ~new_n410_;
  assign new_n412_ = 7 & ~97;
  assign new_n413_1_ = ~7 & 97;
  assign new_n414_ = ~new_n412_ & ~new_n413_1_;
  assign new_n415_ = 6 & ~96;
  assign new_n416_ = ~6 & 96;
  assign new_n417_ = ~new_n415_ & ~new_n416_;
  assign new_n418_1_ = 5 & ~95;
  assign new_n419_ = ~5 & 95;
  assign new_n420_ = ~new_n418_1_ & ~new_n419_;
  assign new_n421_ = 4 & ~94;
  assign new_n422_ = ~4 & 94;
  assign new_n423_1_ = ~new_n421_ & ~new_n422_;
  assign new_n424_ = 4 & ~new_n423_1_;
  assign new_n425_ = new_n420_ & new_n424_;
  assign new_n426_ = 5 & ~new_n420_;
  assign new_n427_ = ~new_n425_ & ~new_n426_;
  assign new_n428_1_ = new_n417_ & ~new_n427_;
  assign new_n429_ = 6 & ~new_n417_;
  assign new_n430_ = ~new_n428_1_ & ~new_n429_;
  assign new_n431_ = new_n414_ & ~new_n430_;
  assign new_n432_ = 7 & ~new_n414_;
  assign new_n433_1_ = ~new_n431_ & ~new_n432_;
  assign new_n434_ = new_n411_ & ~new_n433_1_;
  assign new_n435_ = 8 & ~new_n411_;
  assign new_n436_ = ~new_n434_ & ~new_n435_;
  assign new_n437_ = new_n408_1_ & ~new_n436_;
  assign new_n438_1_ = 9 & ~new_n408_1_;
  assign new_n439_ = ~new_n437_ & ~new_n438_1_;
  assign new_n440_ = new_n405_ & ~new_n439_;
  assign new_n441_ = 10 & ~new_n405_;
  assign new_n442_ = ~new_n440_ & ~new_n441_;
  assign new_n443_1_ = new_n402_ & ~new_n442_;
  assign new_n444_ = 11 & ~new_n402_;
  assign new_n445_ = ~new_n443_1_ & ~new_n444_;
  assign new_n446_ = new_n399_ & ~new_n445_;
  assign new_n447_ = 12 & ~new_n399_;
  assign new_n448_1_ = ~new_n446_ & ~new_n447_;
  assign new_n449_ = new_n396_ & ~new_n448_1_;
  assign new_n450_ = 13 & ~new_n396_;
  assign new_n451_ = ~new_n449_ & ~new_n450_;
  assign new_n452_ = new_n393_1_ & ~new_n451_;
  assign new_n453_1_ = 14 & ~new_n393_1_;
  assign new_n454_ = ~new_n452_ & ~new_n453_1_;
  assign new_n455_ = new_n390_ & ~new_n454_;
  assign new_n456_ = 15 & ~new_n390_;
  assign new_n457_ = ~new_n455_ & ~new_n456_;
  assign new_n458_1_ = new_n387_ & ~new_n457_;
  assign new_n459_ = 16 & ~new_n387_;
  assign new_n460_ = ~new_n458_1_ & ~new_n459_;
  assign new_n461_ = new_n384_ & ~new_n460_;
  assign new_n462_ = 17 & ~new_n384_;
  assign new_n463_1_ = ~new_n461_ & ~new_n462_;
  assign new_n464_ = new_n381_ & ~new_n463_1_;
  assign new_n465_ = 18 & ~new_n381_;
  assign new_n466_ = ~new_n464_ & ~new_n465_;
  assign new_n467_ = new_n378_1_ & ~new_n466_;
  assign new_n468_1_ = 19 & ~new_n378_1_;
  assign new_n469_ = ~new_n467_ & ~new_n468_1_;
  assign new_n470_ = new_n375_ & ~new_n469_;
  assign new_n471_ = 20 & ~new_n375_;
  assign new_n472_ = ~new_n470_ & ~new_n471_;
  assign new_n473_1_ = new_n372_ & ~new_n472_;
  assign new_n474_ = 21 & ~new_n372_;
  assign new_n475_ = ~new_n473_1_ & ~new_n474_;
  assign new_n476_ = new_n369_ & ~new_n475_;
  assign new_n477_ = 22 & ~new_n369_;
  assign new_n478_1_ = ~new_n476_ & ~new_n477_;
  assign new_n479_ = new_n366_ & ~new_n478_1_;
  assign new_n480_ = 23 & ~new_n366_;
  assign new_n481_ = ~new_n479_ & ~new_n480_;
  assign new_n482_ = new_n363_1_ & ~new_n481_;
  assign new_n483_1_ = 24 & ~new_n363_1_;
  assign new_n484_ = ~new_n482_ & ~new_n483_1_;
  assign new_n485_ = new_n360_ & ~new_n484_;
  assign new_n486_ = 25 & ~new_n360_;
  assign new_n487_ = ~new_n485_ & ~new_n486_;
  assign new_n488_1_ = new_n357_ & ~new_n487_;
  assign new_n489_ = 26 & ~new_n357_;
  assign new_n490_ = ~new_n488_1_ & ~new_n489_;
  assign new_n491_ = new_n354_ & ~new_n490_;
  assign new_n492_ = 27 & ~new_n354_;
  assign new_n493_1_ = ~new_n491_ & ~new_n492_;
  assign new_n494_ = new_n351_ & ~new_n493_1_;
  assign new_n495_ = 28 & ~new_n351_;
  assign new_n496_ = ~new_n494_ & ~new_n495_;
  assign new_n497_ = new_n348_1_ & ~new_n496_;
  assign new_n498_1_ = 29 & ~new_n348_1_;
  assign new_n499_ = ~new_n497_ & ~new_n498_1_;
  assign new_n500_ = new_n345_ & ~new_n499_;
  assign new_n501_ = 30 & ~new_n345_;
  assign new_n502_ = ~new_n500_ & ~new_n501_;
  assign new_n503_1_ = new_n342_ & ~new_n502_;
  assign new_n504_ = 31 & ~new_n342_;
  assign new_n505_ = ~new_n503_1_ & ~new_n504_;
  assign new_n506_ = new_n339_ & ~new_n505_;
  assign new_n507_ = 32 & ~new_n339_;
  assign new_n508_1_ = ~new_n506_ & ~new_n507_;
  assign new_n509_ = new_n336_ & ~new_n508_1_;
  assign new_n510_ = 33 & ~new_n336_;
  assign new_n511_ = ~new_n509_ & ~new_n510_;
  assign new_n512_ = 2 & ~3;
  assign new_n513_1_ = ~\1  & new_n512_;
  assign new_n514_ = ~new_n511_ & new_n513_1_;
  assign new_n515_ = 94 & ~new_n514_;
  assign new_n516_ = 4 & new_n514_;
  assign new_n517_ = ~new_n515_ & ~new_n516_;
  assign new_n518_1_ = new_n513_1_ & ~new_n517_;
  assign new_n519_ = 33 & ~93;
  assign new_n520_ = ~33 & 93;
  assign new_n521_ = ~new_n519_ & ~new_n520_;
  assign new_n522_ = 32 & ~92;
  assign new_n523_1_ = ~32 & 92;
  assign new_n524_ = ~new_n522_ & ~new_n523_1_;
  assign new_n525_ = 31 & ~91;
  assign new_n526_ = ~31 & 91;
  assign new_n527_ = ~new_n525_ & ~new_n526_;
  assign new_n528_1_ = 30 & ~90;
  assign new_n529_ = ~30 & 90;
  assign new_n530_ = ~new_n528_1_ & ~new_n529_;
  assign new_n531_ = 29 & ~89;
  assign new_n532_ = ~29 & 89;
  assign new_n533_1_ = ~new_n531_ & ~new_n532_;
  assign new_n534_ = 28 & ~88;
  assign new_n535_ = ~28 & 88;
  assign new_n536_ = ~new_n534_ & ~new_n535_;
  assign new_n537_ = 27 & ~87;
  assign new_n538_1_ = ~27 & 87;
  assign new_n539_ = ~new_n537_ & ~new_n538_1_;
  assign new_n540_ = 26 & ~86;
  assign new_n541_ = ~26 & 86;
  assign new_n542_ = ~new_n540_ & ~new_n541_;
  assign new_n543_1_ = 25 & ~85;
  assign new_n544_ = ~25 & 85;
  assign new_n545_ = ~new_n543_1_ & ~new_n544_;
  assign new_n546_ = 24 & ~84;
  assign new_n547_ = ~24 & 84;
  assign new_n548_1_ = ~new_n546_ & ~new_n547_;
  assign new_n549_ = 23 & ~83;
  assign new_n550_ = ~23 & 83;
  assign new_n551_ = ~new_n549_ & ~new_n550_;
  assign new_n552_ = 22 & ~82;
  assign new_n553_1_ = ~22 & 82;
  assign new_n554_ = ~new_n552_ & ~new_n553_1_;
  assign new_n555_ = 21 & ~81;
  assign new_n556_ = ~21 & 81;
  assign new_n557_ = ~new_n555_ & ~new_n556_;
  assign new_n558_1_ = 20 & ~80;
  assign new_n559_ = ~20 & 80;
  assign new_n560_ = ~new_n558_1_ & ~new_n559_;
  assign new_n561_ = 19 & ~79;
  assign new_n562_ = ~19 & 79;
  assign new_n563_1_ = ~new_n561_ & ~new_n562_;
  assign new_n564_ = 18 & ~78;
  assign new_n565_ = ~18 & 78;
  assign new_n566_ = ~new_n564_ & ~new_n565_;
  assign new_n567_ = 17 & ~77;
  assign new_n568_1_ = ~17 & 77;
  assign new_n569_ = ~new_n567_ & ~new_n568_1_;
  assign new_n570_ = 16 & ~76;
  assign new_n571_ = ~16 & 76;
  assign new_n572_ = ~new_n570_ & ~new_n571_;
  assign new_n573_1_ = 15 & ~75;
  assign new_n574_ = ~15 & 75;
  assign new_n575_ = ~new_n573_1_ & ~new_n574_;
  assign new_n576_ = 14 & ~74;
  assign new_n577_ = ~14 & 74;
  assign new_n578_ = ~new_n576_ & ~new_n577_;
  assign new_n579_ = 13 & ~73;
  assign new_n580_ = ~13 & 73;
  assign new_n581_ = ~new_n579_ & ~new_n580_;
  assign new_n582_ = 12 & ~72;
  assign new_n583_ = ~12 & 72;
  assign new_n584_ = ~new_n582_ & ~new_n583_;
  assign new_n585_ = 11 & ~71;
  assign new_n586_ = ~11 & 71;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = 10 & ~70;
  assign new_n589_ = ~10 & 70;
  assign new_n590_ = ~new_n588_ & ~new_n589_;
  assign new_n591_ = 9 & ~69;
  assign new_n592_ = ~9 & 69;
  assign new_n593_ = ~new_n591_ & ~new_n592_;
  assign new_n594_ = 8 & ~68;
  assign new_n595_ = ~8 & 68;
  assign new_n596_ = ~new_n594_ & ~new_n595_;
  assign new_n597_ = 7 & ~67;
  assign new_n598_ = ~7 & 67;
  assign new_n599_ = ~new_n597_ & ~new_n598_;
  assign new_n600_ = 6 & ~66;
  assign new_n601_ = ~6 & 66;
  assign new_n602_ = ~new_n600_ & ~new_n601_;
  assign new_n603_ = 5 & ~65;
  assign new_n604_ = ~5 & 65;
  assign new_n605_ = ~new_n603_ & ~new_n604_;
  assign new_n606_ = 4 & ~64;
  assign new_n607_ = ~4 & 64;
  assign new_n608_ = ~new_n606_ & ~new_n607_;
  assign new_n609_ = 4 & ~new_n608_;
  assign new_n610_ = new_n605_ & new_n609_;
  assign new_n611_ = 5 & ~new_n605_;
  assign new_n612_ = ~new_n610_ & ~new_n611_;
  assign new_n613_ = new_n602_ & ~new_n612_;
  assign new_n614_ = 6 & ~new_n602_;
  assign new_n615_ = ~new_n613_ & ~new_n614_;
  assign new_n616_ = new_n599_ & ~new_n615_;
  assign new_n617_ = 7 & ~new_n599_;
  assign new_n618_ = ~new_n616_ & ~new_n617_;
  assign new_n619_ = new_n596_ & ~new_n618_;
  assign new_n620_ = 8 & ~new_n596_;
  assign new_n621_ = ~new_n619_ & ~new_n620_;
  assign new_n622_ = new_n593_ & ~new_n621_;
  assign new_n623_ = 9 & ~new_n593_;
  assign new_n624_ = ~new_n622_ & ~new_n623_;
  assign new_n625_ = new_n590_ & ~new_n624_;
  assign new_n626_ = 10 & ~new_n590_;
  assign new_n627_ = ~new_n625_ & ~new_n626_;
  assign new_n628_ = new_n587_ & ~new_n627_;
  assign new_n629_ = 11 & ~new_n587_;
  assign new_n630_ = ~new_n628_ & ~new_n629_;
  assign new_n631_ = new_n584_ & ~new_n630_;
  assign new_n632_ = 12 & ~new_n584_;
  assign new_n633_ = ~new_n631_ & ~new_n632_;
  assign new_n634_ = new_n581_ & ~new_n633_;
  assign new_n635_ = 13 & ~new_n581_;
  assign new_n636_ = ~new_n634_ & ~new_n635_;
  assign new_n637_ = new_n578_ & ~new_n636_;
  assign new_n638_ = 14 & ~new_n578_;
  assign new_n639_ = ~new_n637_ & ~new_n638_;
  assign new_n640_ = new_n575_ & ~new_n639_;
  assign new_n641_ = 15 & ~new_n575_;
  assign new_n642_ = ~new_n640_ & ~new_n641_;
  assign new_n643_ = new_n572_ & ~new_n642_;
  assign new_n644_ = 16 & ~new_n572_;
  assign new_n645_ = ~new_n643_ & ~new_n644_;
  assign new_n646_ = new_n569_ & ~new_n645_;
  assign new_n647_ = 17 & ~new_n569_;
  assign new_n648_ = ~new_n646_ & ~new_n647_;
  assign new_n649_ = new_n566_ & ~new_n648_;
  assign new_n650_ = 18 & ~new_n566_;
  assign new_n651_ = ~new_n649_ & ~new_n650_;
  assign new_n652_ = new_n563_1_ & ~new_n651_;
  assign new_n653_ = 19 & ~new_n563_1_;
  assign new_n654_ = ~new_n652_ & ~new_n653_;
  assign new_n655_ = new_n560_ & ~new_n654_;
  assign new_n656_ = 20 & ~new_n560_;
  assign new_n657_ = ~new_n655_ & ~new_n656_;
  assign new_n658_ = new_n557_ & ~new_n657_;
  assign new_n659_ = 21 & ~new_n557_;
  assign new_n660_ = ~new_n658_ & ~new_n659_;
  assign new_n661_ = new_n554_ & ~new_n660_;
  assign new_n662_ = 22 & ~new_n554_;
  assign new_n663_ = ~new_n661_ & ~new_n662_;
  assign new_n664_ = new_n551_ & ~new_n663_;
  assign new_n665_ = 23 & ~new_n551_;
  assign new_n666_ = ~new_n664_ & ~new_n665_;
  assign new_n667_ = new_n548_1_ & ~new_n666_;
  assign new_n668_ = 24 & ~new_n548_1_;
  assign new_n669_ = ~new_n667_ & ~new_n668_;
  assign new_n670_ = new_n545_ & ~new_n669_;
  assign new_n671_ = 25 & ~new_n545_;
  assign new_n672_ = ~new_n670_ & ~new_n671_;
  assign new_n673_ = new_n542_ & ~new_n672_;
  assign new_n674_ = 26 & ~new_n542_;
  assign new_n675_ = ~new_n673_ & ~new_n674_;
  assign new_n676_ = new_n539_ & ~new_n675_;
  assign new_n677_ = 27 & ~new_n539_;
  assign new_n678_ = ~new_n676_ & ~new_n677_;
  assign new_n679_ = new_n536_ & ~new_n678_;
  assign new_n680_ = 28 & ~new_n536_;
  assign new_n681_ = ~new_n679_ & ~new_n680_;
  assign new_n682_ = new_n533_1_ & ~new_n681_;
  assign new_n683_ = 29 & ~new_n533_1_;
  assign new_n684_ = ~new_n682_ & ~new_n683_;
  assign new_n685_ = new_n530_ & ~new_n684_;
  assign new_n686_ = 30 & ~new_n530_;
  assign new_n687_ = ~new_n685_ & ~new_n686_;
  assign new_n688_ = new_n527_ & ~new_n687_;
  assign new_n689_ = 31 & ~new_n527_;
  assign new_n690_ = ~new_n688_ & ~new_n689_;
  assign new_n691_ = new_n524_ & ~new_n690_;
  assign new_n692_ = 32 & ~new_n524_;
  assign new_n693_ = ~new_n691_ & ~new_n692_;
  assign new_n694_ = new_n521_ & ~new_n693_;
  assign new_n695_ = 33 & ~new_n521_;
  assign new_n696_ = ~new_n694_ & ~new_n695_;
  assign new_n697_ = new_n513_1_ & ~new_n696_;
  assign new_n698_ = 64 & new_n697_;
  assign new_n699_ = 4 & ~new_n697_;
  assign new_n700_ = ~new_n698_ & ~new_n699_;
  assign new_n701_ = new_n513_1_ & ~new_n700_;
  assign new_n702_ = new_n518_1_ & new_n701_;
  assign new_n703_ = 95 & ~new_n514_;
  assign new_n704_ = 5 & new_n514_;
  assign new_n705_ = ~new_n703_ & ~new_n704_;
  assign new_n706_ = new_n513_1_ & ~new_n705_;
  assign new_n707_ = 65 & new_n697_;
  assign new_n708_ = 5 & ~new_n697_;
  assign new_n709_ = ~new_n707_ & ~new_n708_;
  assign new_n710_ = new_n513_1_ & ~new_n709_;
  assign new_n711_ = ~new_n706_ & ~new_n710_;
  assign new_n712_ = new_n706_ & new_n710_;
  assign new_n713_ = ~new_n711_ & ~new_n712_;
  assign new_n714_ = new_n702_ & ~new_n713_;
  assign new_n715_ = ~new_n706_ & new_n710_;
  assign new_n716_ = new_n706_ & ~new_n710_;
  assign new_n717_ = ~new_n715_ & ~new_n716_;
  assign new_n718_ = ~new_n702_ & ~new_n717_;
  assign new_n719_ = ~new_n714_ & ~new_n718_;
  assign new_n720_ = ~3 & ~new_n719_;
  assign new_n721_ = 3 & 4;
  assign new_n722_ = ~new_n720_ & ~new_n721_;
  assign new_n723_ = 2 & ~new_n722_;
  assign new_n724_ = ~2 & 34;
  assign new_n725_ = ~new_n723_ & ~new_n724_;
  assign 124 = ~\1  & ~new_n725_;
  assign new_n727_ = new_n702_ & ~new_n711_;
  assign new_n728_ = ~new_n712_ & ~new_n727_;
  assign new_n729_ = 96 & ~new_n514_;
  assign new_n730_ = 6 & new_n514_;
  assign new_n731_ = ~new_n729_ & ~new_n730_;
  assign new_n732_ = new_n513_1_ & ~new_n731_;
  assign new_n733_ = 66 & new_n697_;
  assign new_n734_ = 6 & ~new_n697_;
  assign new_n735_ = ~new_n733_ & ~new_n734_;
  assign new_n736_ = new_n513_1_ & ~new_n735_;
  assign new_n737_ = ~new_n732_ & ~new_n736_;
  assign new_n738_ = new_n732_ & new_n736_;
  assign new_n739_ = ~new_n737_ & ~new_n738_;
  assign new_n740_ = ~new_n728_ & ~new_n739_;
  assign new_n741_ = ~new_n732_ & new_n736_;
  assign new_n742_ = new_n732_ & ~new_n736_;
  assign new_n743_ = ~new_n741_ & ~new_n742_;
  assign new_n744_ = new_n728_ & ~new_n743_;
  assign new_n745_ = ~new_n740_ & ~new_n744_;
  assign new_n746_ = ~3 & ~new_n745_;
  assign new_n747_ = 3 & 5;
  assign new_n748_ = ~new_n746_ & ~new_n747_;
  assign new_n749_ = 2 & ~new_n748_;
  assign new_n750_ = ~2 & 35;
  assign new_n751_ = ~new_n749_ & ~new_n750_;
  assign 125 = ~\1  & ~new_n751_;
  assign new_n753_ = ~new_n728_ & ~new_n737_;
  assign new_n754_ = ~new_n738_ & ~new_n753_;
  assign new_n755_ = 97 & ~new_n514_;
  assign new_n756_ = 7 & new_n514_;
  assign new_n757_ = ~new_n755_ & ~new_n756_;
  assign new_n758_ = new_n513_1_ & ~new_n757_;
  assign new_n759_ = 67 & new_n697_;
  assign new_n760_ = 7 & ~new_n697_;
  assign new_n761_ = ~new_n759_ & ~new_n760_;
  assign new_n762_ = new_n513_1_ & ~new_n761_;
  assign new_n763_ = ~new_n758_ & ~new_n762_;
  assign new_n764_ = new_n758_ & new_n762_;
  assign new_n765_ = ~new_n763_ & ~new_n764_;
  assign new_n766_ = ~new_n754_ & ~new_n765_;
  assign new_n767_ = ~new_n758_ & new_n762_;
  assign new_n768_ = new_n758_ & ~new_n762_;
  assign new_n769_ = ~new_n767_ & ~new_n768_;
  assign new_n770_ = new_n754_ & ~new_n769_;
  assign new_n771_ = ~new_n766_ & ~new_n770_;
  assign new_n772_ = ~3 & ~new_n771_;
  assign new_n773_ = 3 & 6;
  assign new_n774_ = ~new_n772_ & ~new_n773_;
  assign new_n775_ = 2 & ~new_n774_;
  assign new_n776_ = ~2 & 36;
  assign new_n777_ = ~new_n775_ & ~new_n776_;
  assign 126 = ~\1  & ~new_n777_;
  assign new_n779_ = ~new_n754_ & ~new_n763_;
  assign new_n780_ = ~new_n764_ & ~new_n779_;
  assign new_n781_ = 98 & ~new_n514_;
  assign new_n782_ = 8 & new_n514_;
  assign new_n783_ = ~new_n781_ & ~new_n782_;
  assign new_n784_ = new_n513_1_ & ~new_n783_;
  assign new_n785_ = 68 & new_n697_;
  assign new_n786_ = 8 & ~new_n697_;
  assign new_n787_ = ~new_n785_ & ~new_n786_;
  assign new_n788_ = new_n513_1_ & ~new_n787_;
  assign new_n789_ = ~new_n784_ & ~new_n788_;
  assign new_n790_ = new_n784_ & new_n788_;
  assign new_n791_ = ~new_n789_ & ~new_n790_;
  assign new_n792_ = ~new_n780_ & ~new_n791_;
  assign new_n793_ = ~new_n784_ & new_n788_;
  assign new_n794_ = new_n784_ & ~new_n788_;
  assign new_n795_ = ~new_n793_ & ~new_n794_;
  assign new_n796_ = new_n780_ & ~new_n795_;
  assign new_n797_ = ~new_n792_ & ~new_n796_;
  assign new_n798_ = ~3 & ~new_n797_;
  assign new_n799_ = 3 & 7;
  assign new_n800_ = ~new_n798_ & ~new_n799_;
  assign new_n801_ = 2 & ~new_n800_;
  assign new_n802_ = ~2 & 37;
  assign new_n803_ = ~new_n801_ & ~new_n802_;
  assign 127 = ~\1  & ~new_n803_;
  assign new_n805_ = ~new_n780_ & ~new_n789_;
  assign new_n806_ = ~new_n790_ & ~new_n805_;
  assign new_n807_ = 99 & ~new_n514_;
  assign new_n808_ = 9 & new_n514_;
  assign new_n809_ = ~new_n807_ & ~new_n808_;
  assign new_n810_ = new_n513_1_ & ~new_n809_;
  assign new_n811_ = 69 & new_n697_;
  assign new_n812_ = 9 & ~new_n697_;
  assign new_n813_ = ~new_n811_ & ~new_n812_;
  assign new_n814_ = new_n513_1_ & ~new_n813_;
  assign new_n815_ = ~new_n810_ & ~new_n814_;
  assign new_n816_ = new_n810_ & new_n814_;
  assign new_n817_ = ~new_n815_ & ~new_n816_;
  assign new_n818_ = ~new_n806_ & ~new_n817_;
  assign new_n819_ = ~new_n810_ & new_n814_;
  assign new_n820_ = new_n810_ & ~new_n814_;
  assign new_n821_ = ~new_n819_ & ~new_n820_;
  assign new_n822_ = new_n806_ & ~new_n821_;
  assign new_n823_ = ~new_n818_ & ~new_n822_;
  assign new_n824_ = ~3 & ~new_n823_;
  assign new_n825_ = 3 & 8;
  assign new_n826_ = ~new_n824_ & ~new_n825_;
  assign new_n827_ = 2 & ~new_n826_;
  assign new_n828_ = ~2 & 38;
  assign new_n829_ = ~new_n827_ & ~new_n828_;
  assign 128 = ~\1  & ~new_n829_;
  assign new_n831_ = ~new_n806_ & ~new_n815_;
  assign new_n832_ = ~new_n816_ & ~new_n831_;
  assign new_n833_ = 100 & ~new_n514_;
  assign new_n834_ = 10 & new_n514_;
  assign new_n835_ = ~new_n833_ & ~new_n834_;
  assign new_n836_ = new_n513_1_ & ~new_n835_;
  assign new_n837_ = 70 & new_n697_;
  assign new_n838_ = 10 & ~new_n697_;
  assign new_n839_ = ~new_n837_ & ~new_n838_;
  assign new_n840_ = new_n513_1_ & ~new_n839_;
  assign new_n841_ = ~new_n836_ & ~new_n840_;
  assign new_n842_ = new_n836_ & new_n840_;
  assign new_n843_ = ~new_n841_ & ~new_n842_;
  assign new_n844_ = ~new_n832_ & ~new_n843_;
  assign new_n845_ = ~new_n836_ & new_n840_;
  assign new_n846_ = new_n836_ & ~new_n840_;
  assign new_n847_ = ~new_n845_ & ~new_n846_;
  assign new_n848_ = new_n832_ & ~new_n847_;
  assign new_n849_ = ~new_n844_ & ~new_n848_;
  assign new_n850_ = ~3 & ~new_n849_;
  assign new_n851_ = 3 & 9;
  assign new_n852_ = ~new_n850_ & ~new_n851_;
  assign new_n853_ = 2 & ~new_n852_;
  assign new_n854_ = ~2 & 39;
  assign new_n855_ = ~new_n853_ & ~new_n854_;
  assign 129 = ~\1  & ~new_n855_;
  assign new_n857_ = ~new_n832_ & ~new_n841_;
  assign new_n858_ = ~new_n842_ & ~new_n857_;
  assign new_n859_ = 101 & ~new_n514_;
  assign new_n860_ = 11 & new_n514_;
  assign new_n861_ = ~new_n859_ & ~new_n860_;
  assign new_n862_ = new_n513_1_ & ~new_n861_;
  assign new_n863_ = 71 & new_n697_;
  assign new_n864_ = 11 & ~new_n697_;
  assign new_n865_ = ~new_n863_ & ~new_n864_;
  assign new_n866_ = new_n513_1_ & ~new_n865_;
  assign new_n867_ = ~new_n862_ & ~new_n866_;
  assign new_n868_ = new_n862_ & new_n866_;
  assign new_n869_ = ~new_n867_ & ~new_n868_;
  assign new_n870_ = ~new_n858_ & ~new_n869_;
  assign new_n871_ = ~new_n862_ & new_n866_;
  assign new_n872_ = new_n862_ & ~new_n866_;
  assign new_n873_ = ~new_n871_ & ~new_n872_;
  assign new_n874_ = new_n858_ & ~new_n873_;
  assign new_n875_ = ~new_n870_ & ~new_n874_;
  assign new_n876_ = ~3 & ~new_n875_;
  assign new_n877_ = 3 & 10;
  assign new_n878_ = ~new_n876_ & ~new_n877_;
  assign new_n879_ = 2 & ~new_n878_;
  assign new_n880_ = ~2 & 40;
  assign new_n881_ = ~new_n879_ & ~new_n880_;
  assign 130 = ~\1  & ~new_n881_;
  assign new_n883_ = ~new_n858_ & ~new_n867_;
  assign new_n884_ = ~new_n868_ & ~new_n883_;
  assign new_n885_ = 102 & ~new_n514_;
  assign new_n886_ = 12 & new_n514_;
  assign new_n887_ = ~new_n885_ & ~new_n886_;
  assign new_n888_ = new_n513_1_ & ~new_n887_;
  assign new_n889_ = 72 & new_n697_;
  assign new_n890_ = 12 & ~new_n697_;
  assign new_n891_ = ~new_n889_ & ~new_n890_;
  assign new_n892_ = new_n513_1_ & ~new_n891_;
  assign new_n893_ = ~new_n888_ & ~new_n892_;
  assign new_n894_ = new_n888_ & new_n892_;
  assign new_n895_ = ~new_n893_ & ~new_n894_;
  assign new_n896_ = ~new_n884_ & ~new_n895_;
  assign new_n897_ = ~new_n888_ & new_n892_;
  assign new_n898_ = new_n888_ & ~new_n892_;
  assign new_n899_ = ~new_n897_ & ~new_n898_;
  assign new_n900_ = new_n884_ & ~new_n899_;
  assign new_n901_ = ~new_n896_ & ~new_n900_;
  assign new_n902_ = ~3 & ~new_n901_;
  assign new_n903_ = 3 & 11;
  assign new_n904_ = ~new_n902_ & ~new_n903_;
  assign new_n905_ = 2 & ~new_n904_;
  assign new_n906_ = ~2 & 41;
  assign new_n907_ = ~new_n905_ & ~new_n906_;
  assign 131 = ~\1  & ~new_n907_;
  assign new_n909_ = ~new_n884_ & ~new_n893_;
  assign new_n910_ = ~new_n894_ & ~new_n909_;
  assign new_n911_ = 103 & ~new_n514_;
  assign new_n912_ = 13 & new_n514_;
  assign new_n913_ = ~new_n911_ & ~new_n912_;
  assign new_n914_ = new_n513_1_ & ~new_n913_;
  assign new_n915_ = 73 & new_n697_;
  assign new_n916_ = 13 & ~new_n697_;
  assign new_n917_ = ~new_n915_ & ~new_n916_;
  assign new_n918_ = new_n513_1_ & ~new_n917_;
  assign new_n919_ = ~new_n914_ & ~new_n918_;
  assign new_n920_ = new_n914_ & new_n918_;
  assign new_n921_ = ~new_n919_ & ~new_n920_;
  assign new_n922_ = ~new_n910_ & ~new_n921_;
  assign new_n923_ = ~new_n914_ & new_n918_;
  assign new_n924_ = new_n914_ & ~new_n918_;
  assign new_n925_ = ~new_n923_ & ~new_n924_;
  assign new_n926_ = new_n910_ & ~new_n925_;
  assign new_n927_ = ~new_n922_ & ~new_n926_;
  assign new_n928_ = ~3 & ~new_n927_;
  assign new_n929_ = 3 & 12;
  assign new_n930_ = ~new_n928_ & ~new_n929_;
  assign new_n931_ = 2 & ~new_n930_;
  assign new_n932_ = ~2 & 42;
  assign new_n933_ = ~new_n931_ & ~new_n932_;
  assign 132 = ~\1  & ~new_n933_;
  assign new_n935_ = ~new_n910_ & ~new_n919_;
  assign new_n936_ = ~new_n920_ & ~new_n935_;
  assign new_n937_ = 104 & ~new_n514_;
  assign new_n938_ = 14 & new_n514_;
  assign new_n939_ = ~new_n937_ & ~new_n938_;
  assign new_n940_ = new_n513_1_ & ~new_n939_;
  assign new_n941_ = 74 & new_n697_;
  assign new_n942_ = 14 & ~new_n697_;
  assign new_n943_ = ~new_n941_ & ~new_n942_;
  assign new_n944_ = new_n513_1_ & ~new_n943_;
  assign new_n945_ = ~new_n940_ & ~new_n944_;
  assign new_n946_ = new_n940_ & new_n944_;
  assign new_n947_ = ~new_n945_ & ~new_n946_;
  assign new_n948_ = ~new_n936_ & ~new_n947_;
  assign new_n949_ = ~new_n940_ & new_n944_;
  assign new_n950_ = new_n940_ & ~new_n944_;
  assign new_n951_ = ~new_n949_ & ~new_n950_;
  assign new_n952_ = new_n936_ & ~new_n951_;
  assign new_n953_ = ~new_n948_ & ~new_n952_;
  assign new_n954_ = ~3 & ~new_n953_;
  assign new_n955_ = 3 & 13;
  assign new_n956_ = ~new_n954_ & ~new_n955_;
  assign new_n957_ = 2 & ~new_n956_;
  assign new_n958_ = ~2 & 43;
  assign new_n959_ = ~new_n957_ & ~new_n958_;
  assign 133 = ~\1  & ~new_n959_;
  assign new_n961_ = ~new_n936_ & ~new_n945_;
  assign new_n962_ = ~new_n946_ & ~new_n961_;
  assign new_n963_ = 105 & ~new_n514_;
  assign new_n964_ = 15 & new_n514_;
  assign new_n965_ = ~new_n963_ & ~new_n964_;
  assign new_n966_ = new_n513_1_ & ~new_n965_;
  assign new_n967_ = 75 & new_n697_;
  assign new_n968_ = 15 & ~new_n697_;
  assign new_n969_ = ~new_n967_ & ~new_n968_;
  assign new_n970_ = new_n513_1_ & ~new_n969_;
  assign new_n971_ = ~new_n966_ & ~new_n970_;
  assign new_n972_ = new_n966_ & new_n970_;
  assign new_n973_ = ~new_n971_ & ~new_n972_;
  assign new_n974_ = ~new_n962_ & ~new_n973_;
  assign new_n975_ = ~new_n966_ & new_n970_;
  assign new_n976_ = new_n966_ & ~new_n970_;
  assign new_n977_ = ~new_n975_ & ~new_n976_;
  assign new_n978_ = new_n962_ & ~new_n977_;
  assign new_n979_ = ~new_n974_ & ~new_n978_;
  assign new_n980_ = ~3 & ~new_n979_;
  assign new_n981_ = 3 & 14;
  assign new_n982_ = ~new_n980_ & ~new_n981_;
  assign new_n983_ = 2 & ~new_n982_;
  assign new_n984_ = ~2 & 44;
  assign new_n985_ = ~new_n983_ & ~new_n984_;
  assign 134 = ~\1  & ~new_n985_;
  assign new_n987_ = ~new_n962_ & ~new_n971_;
  assign new_n988_ = ~new_n972_ & ~new_n987_;
  assign new_n989_ = 106 & ~new_n514_;
  assign new_n990_ = 16 & new_n514_;
  assign new_n991_ = ~new_n989_ & ~new_n990_;
  assign new_n992_ = new_n513_1_ & ~new_n991_;
  assign new_n993_ = 76 & new_n697_;
  assign new_n994_ = 16 & ~new_n697_;
  assign new_n995_ = ~new_n993_ & ~new_n994_;
  assign new_n996_ = new_n513_1_ & ~new_n995_;
  assign new_n997_ = ~new_n992_ & ~new_n996_;
  assign new_n998_ = new_n992_ & new_n996_;
  assign new_n999_ = ~new_n997_ & ~new_n998_;
  assign new_n1000_ = ~new_n988_ & ~new_n999_;
  assign new_n1001_ = ~new_n992_ & new_n996_;
  assign new_n1002_ = new_n992_ & ~new_n996_;
  assign new_n1003_ = ~new_n1001_ & ~new_n1002_;
  assign new_n1004_ = new_n988_ & ~new_n1003_;
  assign new_n1005_ = ~new_n1000_ & ~new_n1004_;
  assign new_n1006_ = ~3 & ~new_n1005_;
  assign new_n1007_ = 3 & 15;
  assign new_n1008_ = ~new_n1006_ & ~new_n1007_;
  assign new_n1009_ = 2 & ~new_n1008_;
  assign new_n1010_ = ~2 & 45;
  assign new_n1011_ = ~new_n1009_ & ~new_n1010_;
  assign 135 = ~\1  & ~new_n1011_;
  assign new_n1013_ = ~new_n988_ & ~new_n997_;
  assign new_n1014_ = ~new_n998_ & ~new_n1013_;
  assign new_n1015_ = 107 & ~new_n514_;
  assign new_n1016_ = 17 & new_n514_;
  assign new_n1017_ = ~new_n1015_ & ~new_n1016_;
  assign new_n1018_ = new_n513_1_ & ~new_n1017_;
  assign new_n1019_ = 77 & new_n697_;
  assign new_n1020_ = 17 & ~new_n697_;
  assign new_n1021_ = ~new_n1019_ & ~new_n1020_;
  assign new_n1022_ = new_n513_1_ & ~new_n1021_;
  assign new_n1023_ = ~new_n1018_ & ~new_n1022_;
  assign new_n1024_ = new_n1018_ & new_n1022_;
  assign new_n1025_ = ~new_n1023_ & ~new_n1024_;
  assign new_n1026_ = ~new_n1014_ & ~new_n1025_;
  assign new_n1027_ = ~new_n1018_ & new_n1022_;
  assign new_n1028_ = new_n1018_ & ~new_n1022_;
  assign new_n1029_ = ~new_n1027_ & ~new_n1028_;
  assign new_n1030_ = new_n1014_ & ~new_n1029_;
  assign new_n1031_ = ~new_n1026_ & ~new_n1030_;
  assign new_n1032_ = ~3 & ~new_n1031_;
  assign new_n1033_ = 3 & 16;
  assign new_n1034_ = ~new_n1032_ & ~new_n1033_;
  assign new_n1035_ = 2 & ~new_n1034_;
  assign new_n1036_ = ~2 & 46;
  assign new_n1037_ = ~new_n1035_ & ~new_n1036_;
  assign 136 = ~\1  & ~new_n1037_;
  assign new_n1039_ = ~new_n1014_ & ~new_n1023_;
  assign new_n1040_ = ~new_n1024_ & ~new_n1039_;
  assign new_n1041_ = 108 & ~new_n514_;
  assign new_n1042_ = 18 & new_n514_;
  assign new_n1043_ = ~new_n1041_ & ~new_n1042_;
  assign new_n1044_ = new_n513_1_ & ~new_n1043_;
  assign new_n1045_ = 78 & new_n697_;
  assign new_n1046_ = 18 & ~new_n697_;
  assign new_n1047_ = ~new_n1045_ & ~new_n1046_;
  assign new_n1048_ = new_n513_1_ & ~new_n1047_;
  assign new_n1049_ = ~new_n1044_ & ~new_n1048_;
  assign new_n1050_ = new_n1044_ & new_n1048_;
  assign new_n1051_ = ~new_n1049_ & ~new_n1050_;
  assign new_n1052_ = ~new_n1040_ & ~new_n1051_;
  assign new_n1053_ = ~new_n1044_ & new_n1048_;
  assign new_n1054_ = new_n1044_ & ~new_n1048_;
  assign new_n1055_ = ~new_n1053_ & ~new_n1054_;
  assign new_n1056_ = new_n1040_ & ~new_n1055_;
  assign new_n1057_ = ~new_n1052_ & ~new_n1056_;
  assign new_n1058_ = ~3 & ~new_n1057_;
  assign new_n1059_ = 3 & 17;
  assign new_n1060_ = ~new_n1058_ & ~new_n1059_;
  assign new_n1061_ = 2 & ~new_n1060_;
  assign new_n1062_ = ~2 & 47;
  assign new_n1063_ = ~new_n1061_ & ~new_n1062_;
  assign 137 = ~\1  & ~new_n1063_;
  assign new_n1065_ = ~new_n1040_ & ~new_n1049_;
  assign new_n1066_ = ~new_n1050_ & ~new_n1065_;
  assign new_n1067_ = 109 & ~new_n514_;
  assign new_n1068_ = 19 & new_n514_;
  assign new_n1069_ = ~new_n1067_ & ~new_n1068_;
  assign new_n1070_ = new_n513_1_ & ~new_n1069_;
  assign new_n1071_ = 79 & new_n697_;
  assign new_n1072_ = 19 & ~new_n697_;
  assign new_n1073_ = ~new_n1071_ & ~new_n1072_;
  assign new_n1074_ = new_n513_1_ & ~new_n1073_;
  assign new_n1075_ = ~new_n1070_ & ~new_n1074_;
  assign new_n1076_ = new_n1070_ & new_n1074_;
  assign new_n1077_ = ~new_n1075_ & ~new_n1076_;
  assign new_n1078_ = ~new_n1066_ & ~new_n1077_;
  assign new_n1079_ = ~new_n1070_ & new_n1074_;
  assign new_n1080_ = new_n1070_ & ~new_n1074_;
  assign new_n1081_ = ~new_n1079_ & ~new_n1080_;
  assign new_n1082_ = new_n1066_ & ~new_n1081_;
  assign new_n1083_ = ~new_n1078_ & ~new_n1082_;
  assign new_n1084_ = ~3 & ~new_n1083_;
  assign new_n1085_ = 3 & 18;
  assign new_n1086_ = ~new_n1084_ & ~new_n1085_;
  assign new_n1087_ = 2 & ~new_n1086_;
  assign new_n1088_ = ~2 & 48;
  assign new_n1089_ = ~new_n1087_ & ~new_n1088_;
  assign 138 = ~\1  & ~new_n1089_;
  assign new_n1091_ = ~new_n1066_ & ~new_n1075_;
  assign new_n1092_ = ~new_n1076_ & ~new_n1091_;
  assign new_n1093_ = 110 & ~new_n514_;
  assign new_n1094_ = 20 & new_n514_;
  assign new_n1095_ = ~new_n1093_ & ~new_n1094_;
  assign new_n1096_ = new_n513_1_ & ~new_n1095_;
  assign new_n1097_ = 80 & new_n697_;
  assign new_n1098_ = 20 & ~new_n697_;
  assign new_n1099_ = ~new_n1097_ & ~new_n1098_;
  assign new_n1100_ = new_n513_1_ & ~new_n1099_;
  assign new_n1101_ = ~new_n1096_ & ~new_n1100_;
  assign new_n1102_ = new_n1096_ & new_n1100_;
  assign new_n1103_ = ~new_n1101_ & ~new_n1102_;
  assign new_n1104_ = ~new_n1092_ & ~new_n1103_;
  assign new_n1105_ = ~new_n1096_ & new_n1100_;
  assign new_n1106_ = new_n1096_ & ~new_n1100_;
  assign new_n1107_ = ~new_n1105_ & ~new_n1106_;
  assign new_n1108_ = new_n1092_ & ~new_n1107_;
  assign new_n1109_ = ~new_n1104_ & ~new_n1108_;
  assign new_n1110_ = ~3 & ~new_n1109_;
  assign new_n1111_ = 3 & 19;
  assign new_n1112_ = ~new_n1110_ & ~new_n1111_;
  assign new_n1113_ = 2 & ~new_n1112_;
  assign new_n1114_ = ~2 & 49;
  assign new_n1115_ = ~new_n1113_ & ~new_n1114_;
  assign 139 = ~\1  & ~new_n1115_;
  assign new_n1117_ = ~new_n1092_ & ~new_n1101_;
  assign new_n1118_ = ~new_n1102_ & ~new_n1117_;
  assign new_n1119_ = 111 & ~new_n514_;
  assign new_n1120_ = 21 & new_n514_;
  assign new_n1121_ = ~new_n1119_ & ~new_n1120_;
  assign new_n1122_ = new_n513_1_ & ~new_n1121_;
  assign new_n1123_ = 81 & new_n697_;
  assign new_n1124_ = 21 & ~new_n697_;
  assign new_n1125_ = ~new_n1123_ & ~new_n1124_;
  assign new_n1126_ = new_n513_1_ & ~new_n1125_;
  assign new_n1127_ = ~new_n1122_ & ~new_n1126_;
  assign new_n1128_ = new_n1122_ & new_n1126_;
  assign new_n1129_ = ~new_n1127_ & ~new_n1128_;
  assign new_n1130_ = ~new_n1118_ & ~new_n1129_;
  assign new_n1131_ = ~new_n1122_ & new_n1126_;
  assign new_n1132_ = new_n1122_ & ~new_n1126_;
  assign new_n1133_ = ~new_n1131_ & ~new_n1132_;
  assign new_n1134_ = new_n1118_ & ~new_n1133_;
  assign new_n1135_ = ~new_n1130_ & ~new_n1134_;
  assign new_n1136_ = ~3 & ~new_n1135_;
  assign new_n1137_ = 3 & 20;
  assign new_n1138_ = ~new_n1136_ & ~new_n1137_;
  assign new_n1139_ = 2 & ~new_n1138_;
  assign new_n1140_ = ~2 & 50;
  assign new_n1141_ = ~new_n1139_ & ~new_n1140_;
  assign 140 = ~\1  & ~new_n1141_;
  assign new_n1143_ = ~new_n1118_ & ~new_n1127_;
  assign new_n1144_ = ~new_n1128_ & ~new_n1143_;
  assign new_n1145_ = 112 & ~new_n514_;
  assign new_n1146_ = 22 & new_n514_;
  assign new_n1147_ = ~new_n1145_ & ~new_n1146_;
  assign new_n1148_ = new_n513_1_ & ~new_n1147_;
  assign new_n1149_ = 82 & new_n697_;
  assign new_n1150_ = 22 & ~new_n697_;
  assign new_n1151_ = ~new_n1149_ & ~new_n1150_;
  assign new_n1152_ = new_n513_1_ & ~new_n1151_;
  assign new_n1153_ = ~new_n1148_ & ~new_n1152_;
  assign new_n1154_ = new_n1148_ & new_n1152_;
  assign new_n1155_ = ~new_n1153_ & ~new_n1154_;
  assign new_n1156_ = ~new_n1144_ & ~new_n1155_;
  assign new_n1157_ = ~new_n1148_ & new_n1152_;
  assign new_n1158_ = new_n1148_ & ~new_n1152_;
  assign new_n1159_ = ~new_n1157_ & ~new_n1158_;
  assign new_n1160_ = new_n1144_ & ~new_n1159_;
  assign new_n1161_ = ~new_n1156_ & ~new_n1160_;
  assign new_n1162_ = ~3 & ~new_n1161_;
  assign new_n1163_ = 3 & 21;
  assign new_n1164_ = ~new_n1162_ & ~new_n1163_;
  assign new_n1165_ = 2 & ~new_n1164_;
  assign new_n1166_ = ~2 & 51;
  assign new_n1167_ = ~new_n1165_ & ~new_n1166_;
  assign 141 = ~\1  & ~new_n1167_;
  assign new_n1169_ = ~new_n1144_ & ~new_n1153_;
  assign new_n1170_ = ~new_n1154_ & ~new_n1169_;
  assign new_n1171_ = 113 & ~new_n514_;
  assign new_n1172_ = 23 & new_n514_;
  assign new_n1173_ = ~new_n1171_ & ~new_n1172_;
  assign new_n1174_ = new_n513_1_ & ~new_n1173_;
  assign new_n1175_ = 83 & new_n697_;
  assign new_n1176_ = 23 & ~new_n697_;
  assign new_n1177_ = ~new_n1175_ & ~new_n1176_;
  assign new_n1178_ = new_n513_1_ & ~new_n1177_;
  assign new_n1179_ = ~new_n1174_ & ~new_n1178_;
  assign new_n1180_ = new_n1174_ & new_n1178_;
  assign new_n1181_ = ~new_n1179_ & ~new_n1180_;
  assign new_n1182_ = ~new_n1170_ & ~new_n1181_;
  assign new_n1183_ = ~new_n1174_ & new_n1178_;
  assign new_n1184_ = new_n1174_ & ~new_n1178_;
  assign new_n1185_ = ~new_n1183_ & ~new_n1184_;
  assign new_n1186_ = new_n1170_ & ~new_n1185_;
  assign new_n1187_ = ~new_n1182_ & ~new_n1186_;
  assign new_n1188_ = ~3 & ~new_n1187_;
  assign new_n1189_ = 3 & 22;
  assign new_n1190_ = ~new_n1188_ & ~new_n1189_;
  assign new_n1191_ = 2 & ~new_n1190_;
  assign new_n1192_ = ~2 & 52;
  assign new_n1193_ = ~new_n1191_ & ~new_n1192_;
  assign 142 = ~\1  & ~new_n1193_;
  assign new_n1195_ = ~new_n1170_ & ~new_n1179_;
  assign new_n1196_ = ~new_n1180_ & ~new_n1195_;
  assign new_n1197_ = 114 & ~new_n514_;
  assign new_n1198_ = 24 & new_n514_;
  assign new_n1199_ = ~new_n1197_ & ~new_n1198_;
  assign new_n1200_ = new_n513_1_ & ~new_n1199_;
  assign new_n1201_ = 84 & new_n697_;
  assign new_n1202_ = 24 & ~new_n697_;
  assign new_n1203_ = ~new_n1201_ & ~new_n1202_;
  assign new_n1204_ = new_n513_1_ & ~new_n1203_;
  assign new_n1205_ = ~new_n1200_ & ~new_n1204_;
  assign new_n1206_ = new_n1200_ & new_n1204_;
  assign new_n1207_ = ~new_n1205_ & ~new_n1206_;
  assign new_n1208_ = ~new_n1196_ & ~new_n1207_;
  assign new_n1209_ = ~new_n1200_ & new_n1204_;
  assign new_n1210_ = new_n1200_ & ~new_n1204_;
  assign new_n1211_ = ~new_n1209_ & ~new_n1210_;
  assign new_n1212_ = new_n1196_ & ~new_n1211_;
  assign new_n1213_ = ~new_n1208_ & ~new_n1212_;
  assign new_n1214_ = ~3 & ~new_n1213_;
  assign new_n1215_ = 3 & 23;
  assign new_n1216_ = ~new_n1214_ & ~new_n1215_;
  assign new_n1217_ = 2 & ~new_n1216_;
  assign new_n1218_ = ~2 & 53;
  assign new_n1219_ = ~new_n1217_ & ~new_n1218_;
  assign 143 = ~\1  & ~new_n1219_;
  assign new_n1221_ = ~new_n1196_ & ~new_n1205_;
  assign new_n1222_ = ~new_n1206_ & ~new_n1221_;
  assign new_n1223_ = 115 & ~new_n514_;
  assign new_n1224_ = 25 & new_n514_;
  assign new_n1225_ = ~new_n1223_ & ~new_n1224_;
  assign new_n1226_ = new_n513_1_ & ~new_n1225_;
  assign new_n1227_ = 85 & new_n697_;
  assign new_n1228_ = 25 & ~new_n697_;
  assign new_n1229_ = ~new_n1227_ & ~new_n1228_;
  assign new_n1230_ = new_n513_1_ & ~new_n1229_;
  assign new_n1231_ = ~new_n1226_ & ~new_n1230_;
  assign new_n1232_ = new_n1226_ & new_n1230_;
  assign new_n1233_ = ~new_n1231_ & ~new_n1232_;
  assign new_n1234_ = ~new_n1222_ & ~new_n1233_;
  assign new_n1235_ = ~new_n1226_ & new_n1230_;
  assign new_n1236_ = new_n1226_ & ~new_n1230_;
  assign new_n1237_ = ~new_n1235_ & ~new_n1236_;
  assign new_n1238_ = new_n1222_ & ~new_n1237_;
  assign new_n1239_ = ~new_n1234_ & ~new_n1238_;
  assign new_n1240_ = ~3 & ~new_n1239_;
  assign new_n1241_ = 3 & 24;
  assign new_n1242_ = ~new_n1240_ & ~new_n1241_;
  assign new_n1243_ = 2 & ~new_n1242_;
  assign new_n1244_ = ~2 & 54;
  assign new_n1245_ = ~new_n1243_ & ~new_n1244_;
  assign 144 = ~\1  & ~new_n1245_;
  assign new_n1247_ = ~new_n1222_ & ~new_n1231_;
  assign new_n1248_ = ~new_n1232_ & ~new_n1247_;
  assign new_n1249_ = 116 & ~new_n514_;
  assign new_n1250_ = 26 & new_n514_;
  assign new_n1251_ = ~new_n1249_ & ~new_n1250_;
  assign new_n1252_ = new_n513_1_ & ~new_n1251_;
  assign new_n1253_ = 86 & new_n697_;
  assign new_n1254_ = 26 & ~new_n697_;
  assign new_n1255_ = ~new_n1253_ & ~new_n1254_;
  assign new_n1256_ = new_n513_1_ & ~new_n1255_;
  assign new_n1257_ = ~new_n1252_ & ~new_n1256_;
  assign new_n1258_ = new_n1252_ & new_n1256_;
  assign new_n1259_ = ~new_n1257_ & ~new_n1258_;
  assign new_n1260_ = ~new_n1248_ & ~new_n1259_;
  assign new_n1261_ = ~new_n1252_ & new_n1256_;
  assign new_n1262_ = new_n1252_ & ~new_n1256_;
  assign new_n1263_ = ~new_n1261_ & ~new_n1262_;
  assign new_n1264_ = new_n1248_ & ~new_n1263_;
  assign new_n1265_ = ~new_n1260_ & ~new_n1264_;
  assign new_n1266_ = ~3 & ~new_n1265_;
  assign new_n1267_ = 3 & 25;
  assign new_n1268_ = ~new_n1266_ & ~new_n1267_;
  assign new_n1269_ = 2 & ~new_n1268_;
  assign new_n1270_ = ~2 & 55;
  assign new_n1271_ = ~new_n1269_ & ~new_n1270_;
  assign 145 = ~\1  & ~new_n1271_;
  assign new_n1273_ = ~new_n1248_ & ~new_n1257_;
  assign new_n1274_ = ~new_n1258_ & ~new_n1273_;
  assign new_n1275_ = 117 & ~new_n514_;
  assign new_n1276_ = 27 & new_n514_;
  assign new_n1277_ = ~new_n1275_ & ~new_n1276_;
  assign new_n1278_ = new_n513_1_ & ~new_n1277_;
  assign new_n1279_ = 87 & new_n697_;
  assign new_n1280_ = 27 & ~new_n697_;
  assign new_n1281_ = ~new_n1279_ & ~new_n1280_;
  assign new_n1282_ = new_n513_1_ & ~new_n1281_;
  assign new_n1283_ = ~new_n1278_ & ~new_n1282_;
  assign new_n1284_ = new_n1278_ & new_n1282_;
  assign new_n1285_ = ~new_n1283_ & ~new_n1284_;
  assign new_n1286_ = ~new_n1274_ & ~new_n1285_;
  assign new_n1287_ = ~new_n1278_ & new_n1282_;
  assign new_n1288_ = new_n1278_ & ~new_n1282_;
  assign new_n1289_ = ~new_n1287_ & ~new_n1288_;
  assign new_n1290_ = new_n1274_ & ~new_n1289_;
  assign new_n1291_ = ~new_n1286_ & ~new_n1290_;
  assign new_n1292_ = ~3 & ~new_n1291_;
  assign new_n1293_ = 3 & 26;
  assign new_n1294_ = ~new_n1292_ & ~new_n1293_;
  assign new_n1295_ = 2 & ~new_n1294_;
  assign new_n1296_ = ~2 & 56;
  assign new_n1297_ = ~new_n1295_ & ~new_n1296_;
  assign 146 = ~\1  & ~new_n1297_;
  assign new_n1299_ = ~new_n1274_ & ~new_n1283_;
  assign new_n1300_ = ~new_n1284_ & ~new_n1299_;
  assign new_n1301_ = 118 & ~new_n514_;
  assign new_n1302_ = 28 & new_n514_;
  assign new_n1303_ = ~new_n1301_ & ~new_n1302_;
  assign new_n1304_ = new_n513_1_ & ~new_n1303_;
  assign new_n1305_ = 88 & new_n697_;
  assign new_n1306_ = 28 & ~new_n697_;
  assign new_n1307_ = ~new_n1305_ & ~new_n1306_;
  assign new_n1308_ = new_n513_1_ & ~new_n1307_;
  assign new_n1309_ = ~new_n1304_ & ~new_n1308_;
  assign new_n1310_ = new_n1304_ & new_n1308_;
  assign new_n1311_ = ~new_n1309_ & ~new_n1310_;
  assign new_n1312_ = ~new_n1300_ & ~new_n1311_;
  assign new_n1313_ = ~new_n1304_ & new_n1308_;
  assign new_n1314_ = new_n1304_ & ~new_n1308_;
  assign new_n1315_ = ~new_n1313_ & ~new_n1314_;
  assign new_n1316_ = new_n1300_ & ~new_n1315_;
  assign new_n1317_ = ~new_n1312_ & ~new_n1316_;
  assign new_n1318_ = ~3 & ~new_n1317_;
  assign new_n1319_ = 3 & 27;
  assign new_n1320_ = ~new_n1318_ & ~new_n1319_;
  assign new_n1321_ = 2 & ~new_n1320_;
  assign new_n1322_ = ~2 & 57;
  assign new_n1323_ = ~new_n1321_ & ~new_n1322_;
  assign 147 = ~\1  & ~new_n1323_;
  assign new_n1325_ = ~new_n1300_ & ~new_n1309_;
  assign new_n1326_ = ~new_n1310_ & ~new_n1325_;
  assign new_n1327_ = 119 & ~new_n514_;
  assign new_n1328_ = 29 & new_n514_;
  assign new_n1329_ = ~new_n1327_ & ~new_n1328_;
  assign new_n1330_ = new_n513_1_ & ~new_n1329_;
  assign new_n1331_ = 89 & new_n697_;
  assign new_n1332_ = 29 & ~new_n697_;
  assign new_n1333_ = ~new_n1331_ & ~new_n1332_;
  assign new_n1334_ = new_n513_1_ & ~new_n1333_;
  assign new_n1335_ = ~new_n1330_ & ~new_n1334_;
  assign new_n1336_ = new_n1330_ & new_n1334_;
  assign new_n1337_ = ~new_n1335_ & ~new_n1336_;
  assign new_n1338_ = ~new_n1326_ & ~new_n1337_;
  assign new_n1339_ = ~new_n1330_ & new_n1334_;
  assign new_n1340_ = new_n1330_ & ~new_n1334_;
  assign new_n1341_ = ~new_n1339_ & ~new_n1340_;
  assign new_n1342_ = new_n1326_ & ~new_n1341_;
  assign new_n1343_ = ~new_n1338_ & ~new_n1342_;
  assign new_n1344_ = ~3 & ~new_n1343_;
  assign new_n1345_ = 3 & 28;
  assign new_n1346_ = ~new_n1344_ & ~new_n1345_;
  assign new_n1347_ = 2 & ~new_n1346_;
  assign new_n1348_ = ~2 & 58;
  assign new_n1349_ = ~new_n1347_ & ~new_n1348_;
  assign 148 = ~\1  & ~new_n1349_;
  assign new_n1351_ = ~new_n1326_ & ~new_n1335_;
  assign new_n1352_ = ~new_n1336_ & ~new_n1351_;
  assign new_n1353_ = 120 & ~new_n514_;
  assign new_n1354_ = 30 & new_n514_;
  assign new_n1355_ = ~new_n1353_ & ~new_n1354_;
  assign new_n1356_ = new_n513_1_ & ~new_n1355_;
  assign new_n1357_ = 90 & new_n697_;
  assign new_n1358_ = 30 & ~new_n697_;
  assign new_n1359_ = ~new_n1357_ & ~new_n1358_;
  assign new_n1360_ = new_n513_1_ & ~new_n1359_;
  assign new_n1361_ = ~new_n1356_ & ~new_n1360_;
  assign new_n1362_ = new_n1356_ & new_n1360_;
  assign new_n1363_ = ~new_n1361_ & ~new_n1362_;
  assign new_n1364_ = ~new_n1352_ & ~new_n1363_;
  assign new_n1365_ = ~new_n1356_ & new_n1360_;
  assign new_n1366_ = new_n1356_ & ~new_n1360_;
  assign new_n1367_ = ~new_n1365_ & ~new_n1366_;
  assign new_n1368_ = new_n1352_ & ~new_n1367_;
  assign new_n1369_ = ~new_n1364_ & ~new_n1368_;
  assign new_n1370_ = ~3 & ~new_n1369_;
  assign new_n1371_ = 3 & 29;
  assign new_n1372_ = ~new_n1370_ & ~new_n1371_;
  assign new_n1373_ = 2 & ~new_n1372_;
  assign new_n1374_ = ~2 & 59;
  assign new_n1375_ = ~new_n1373_ & ~new_n1374_;
  assign 149 = ~\1  & ~new_n1375_;
  assign new_n1377_ = ~new_n1352_ & ~new_n1361_;
  assign new_n1378_ = ~new_n1362_ & ~new_n1377_;
  assign new_n1379_ = 121 & ~new_n514_;
  assign new_n1380_ = 31 & new_n514_;
  assign new_n1381_ = ~new_n1379_ & ~new_n1380_;
  assign new_n1382_ = new_n513_1_ & ~new_n1381_;
  assign new_n1383_ = 91 & new_n697_;
  assign new_n1384_ = 31 & ~new_n697_;
  assign new_n1385_ = ~new_n1383_ & ~new_n1384_;
  assign new_n1386_ = new_n513_1_ & ~new_n1385_;
  assign new_n1387_ = ~new_n1382_ & ~new_n1386_;
  assign new_n1388_ = new_n1382_ & new_n1386_;
  assign new_n1389_ = ~new_n1387_ & ~new_n1388_;
  assign new_n1390_ = ~new_n1378_ & ~new_n1389_;
  assign new_n1391_ = ~new_n1382_ & new_n1386_;
  assign new_n1392_ = new_n1382_ & ~new_n1386_;
  assign new_n1393_ = ~new_n1391_ & ~new_n1392_;
  assign new_n1394_ = new_n1378_ & ~new_n1393_;
  assign new_n1395_ = ~new_n1390_ & ~new_n1394_;
  assign new_n1396_ = ~3 & ~new_n1395_;
  assign new_n1397_ = 3 & 30;
  assign new_n1398_ = ~new_n1396_ & ~new_n1397_;
  assign new_n1399_ = 2 & ~new_n1398_;
  assign new_n1400_ = ~2 & 60;
  assign new_n1401_ = ~new_n1399_ & ~new_n1400_;
  assign 150 = ~\1  & ~new_n1401_;
  assign new_n1403_ = ~new_n1378_ & ~new_n1387_;
  assign new_n1404_ = ~new_n1388_ & ~new_n1403_;
  assign new_n1405_ = 122 & ~new_n514_;
  assign new_n1406_ = 32 & new_n514_;
  assign new_n1407_ = ~new_n1405_ & ~new_n1406_;
  assign new_n1408_ = new_n513_1_ & ~new_n1407_;
  assign new_n1409_ = 92 & new_n697_;
  assign new_n1410_ = 32 & ~new_n697_;
  assign new_n1411_ = ~new_n1409_ & ~new_n1410_;
  assign new_n1412_ = new_n513_1_ & ~new_n1411_;
  assign new_n1413_ = ~new_n1408_ & ~new_n1412_;
  assign new_n1414_ = new_n1408_ & new_n1412_;
  assign new_n1415_ = ~new_n1413_ & ~new_n1414_;
  assign new_n1416_ = ~new_n1404_ & ~new_n1415_;
  assign new_n1417_ = ~new_n1408_ & new_n1412_;
  assign new_n1418_ = new_n1408_ & ~new_n1412_;
  assign new_n1419_ = ~new_n1417_ & ~new_n1418_;
  assign new_n1420_ = new_n1404_ & ~new_n1419_;
  assign new_n1421_ = ~new_n1416_ & ~new_n1420_;
  assign new_n1422_ = ~3 & ~new_n1421_;
  assign new_n1423_ = 3 & 31;
  assign new_n1424_ = ~new_n1422_ & ~new_n1423_;
  assign new_n1425_ = 2 & ~new_n1424_;
  assign new_n1426_ = ~2 & 61;
  assign new_n1427_ = ~new_n1425_ & ~new_n1426_;
  assign 151 = ~\1  & ~new_n1427_;
  assign new_n1429_ = ~new_n1404_ & ~new_n1413_;
  assign new_n1430_ = ~new_n1414_ & ~new_n1429_;
  assign new_n1431_ = 123 & ~new_n514_;
  assign new_n1432_ = 33 & new_n514_;
  assign new_n1433_ = ~new_n1431_ & ~new_n1432_;
  assign new_n1434_ = new_n513_1_ & ~new_n1433_;
  assign new_n1435_ = 93 & new_n697_;
  assign new_n1436_ = 33 & ~new_n697_;
  assign new_n1437_ = ~new_n1435_ & ~new_n1436_;
  assign new_n1438_ = new_n513_1_ & ~new_n1437_;
  assign new_n1439_ = ~new_n1434_ & ~new_n1438_;
  assign new_n1440_ = new_n1434_ & new_n1438_;
  assign new_n1441_ = ~new_n1439_ & ~new_n1440_;
  assign new_n1442_ = ~new_n1430_ & ~new_n1441_;
  assign new_n1443_ = ~new_n1434_ & new_n1438_;
  assign new_n1444_ = new_n1434_ & ~new_n1438_;
  assign new_n1445_ = ~new_n1443_ & ~new_n1444_;
  assign new_n1446_ = new_n1430_ & ~new_n1445_;
  assign new_n1447_ = ~new_n1442_ & ~new_n1446_;
  assign new_n1448_ = ~3 & ~new_n1447_;
  assign new_n1449_ = 3 & 32;
  assign new_n1450_ = ~new_n1448_ & ~new_n1449_;
  assign new_n1451_ = 2 & ~new_n1450_;
  assign new_n1452_ = ~2 & 62;
  assign new_n1453_ = ~new_n1451_ & ~new_n1452_;
  assign 152 = ~\1  & ~new_n1453_;
  assign new_n1455_ = ~new_n1430_ & ~new_n1439_;
  assign new_n1456_ = ~new_n1440_ & ~new_n1455_;
  assign new_n1457_ = ~3 & ~new_n1456_;
  assign new_n1458_ = 3 & 33;
  assign new_n1459_ = ~new_n1457_ & ~new_n1458_;
  assign new_n1460_ = 2 & ~new_n1459_;
  assign new_n1461_ = ~2 & 63;
  assign new_n1462_ = ~new_n1460_ & ~new_n1461_;
  assign 153 = ~\1  & ~new_n1462_;
  assign new_n1464_ = 2 & 4;
  assign n128 = ~\1  & new_n1464_;
  assign new_n1466_ = 2 & 5;
  assign n133 = ~\1  & new_n1466_;
  assign new_n1468_ = 2 & 6;
  assign n138 = ~\1  & new_n1468_;
  assign new_n1470_ = 2 & 7;
  assign n143 = ~\1  & new_n1470_;
  assign new_n1472_ = 2 & 8;
  assign n148 = ~\1  & new_n1472_;
  assign new_n1474_ = 2 & 9;
  assign n153 = ~\1  & new_n1474_;
  assign new_n1476_ = 2 & 10;
  assign n158 = ~\1  & new_n1476_;
  assign new_n1478_ = 2 & 11;
  assign n163 = ~\1  & new_n1478_;
  assign new_n1480_ = 2 & 12;
  assign n168 = ~\1  & new_n1480_;
  assign new_n1482_ = 2 & 13;
  assign n173 = ~\1  & new_n1482_;
  assign new_n1484_ = 2 & 14;
  assign n178 = ~\1  & new_n1484_;
  assign new_n1486_ = 2 & 15;
  assign n183 = ~\1  & new_n1486_;
  assign new_n1488_ = 2 & 16;
  assign n188 = ~\1  & new_n1488_;
  assign new_n1490_ = 2 & 17;
  assign n193 = ~\1  & new_n1490_;
  assign new_n1492_ = 2 & 18;
  assign n198 = ~\1  & new_n1492_;
  assign new_n1494_ = 2 & 19;
  assign n203 = ~\1  & new_n1494_;
  assign new_n1496_ = 2 & 20;
  assign n208 = ~\1  & new_n1496_;
  assign new_n1498_ = 2 & 21;
  assign n213 = ~\1  & new_n1498_;
  assign new_n1500_ = 2 & 22;
  assign n218 = ~\1  & new_n1500_;
  assign new_n1502_ = 2 & 23;
  assign n223 = ~\1  & new_n1502_;
  assign new_n1504_ = 2 & 24;
  assign n228 = ~\1  & new_n1504_;
  assign new_n1506_ = 2 & 25;
  assign n233 = ~\1  & new_n1506_;
  assign new_n1508_ = 2 & 26;
  assign n238 = ~\1  & new_n1508_;
  assign new_n1510_ = 2 & 27;
  assign n243 = ~\1  & new_n1510_;
  assign new_n1512_ = 2 & 28;
  assign n248 = ~\1  & new_n1512_;
  assign new_n1514_ = 2 & 29;
  assign n253 = ~\1  & new_n1514_;
  assign new_n1516_ = 2 & 30;
  assign n258 = ~\1  & new_n1516_;
  assign new_n1518_ = 2 & 31;
  assign n263 = ~\1  & new_n1518_;
  assign new_n1520_ = 2 & 32;
  assign n268 = ~\1  & new_n1520_;
  assign new_n1522_ = 2 & 33;
  assign n273 = ~\1  & new_n1522_;
  assign new_n1524_ = ~3 & new_n701_;
  assign new_n1525_ = ~3 & ~new_n1524_;
  assign new_n1526_ = 2 & ~new_n1525_;
  assign new_n1527_ = 2 & ~new_n1526_;
  assign new_n1528_ = ~\1  & ~new_n1527_;
  assign n278 = \1  | new_n1528_;
  assign new_n1530_ = ~3 & new_n710_;
  assign new_n1531_ = ~3 & ~new_n1530_;
  assign new_n1532_ = 2 & ~new_n1531_;
  assign new_n1533_ = 2 & ~new_n1532_;
  assign new_n1534_ = ~\1  & ~new_n1533_;
  assign n283 = \1  | new_n1534_;
  assign new_n1536_ = ~3 & new_n736_;
  assign new_n1537_ = ~3 & ~new_n1536_;
  assign new_n1538_ = 2 & ~new_n1537_;
  assign new_n1539_ = 2 & ~new_n1538_;
  assign new_n1540_ = ~\1  & ~new_n1539_;
  assign n288 = \1  | new_n1540_;
  assign new_n1542_ = ~3 & new_n762_;
  assign new_n1543_ = ~3 & ~new_n1542_;
  assign new_n1544_ = 2 & ~new_n1543_;
  assign new_n1545_ = 2 & ~new_n1544_;
  assign new_n1546_ = ~\1  & ~new_n1545_;
  assign n293 = \1  | new_n1546_;
  assign new_n1548_ = ~3 & new_n788_;
  assign new_n1549_ = ~3 & ~new_n1548_;
  assign new_n1550_ = 2 & ~new_n1549_;
  assign new_n1551_ = 2 & ~new_n1550_;
  assign new_n1552_ = ~\1  & ~new_n1551_;
  assign n298 = \1  | new_n1552_;
  assign new_n1554_ = ~3 & new_n814_;
  assign new_n1555_ = ~3 & ~new_n1554_;
  assign new_n1556_ = 2 & ~new_n1555_;
  assign new_n1557_ = 2 & ~new_n1556_;
  assign new_n1558_ = ~\1  & ~new_n1557_;
  assign n303 = \1  | new_n1558_;
  assign new_n1560_ = ~3 & new_n840_;
  assign new_n1561_ = ~3 & ~new_n1560_;
  assign new_n1562_ = 2 & ~new_n1561_;
  assign new_n1563_ = 2 & ~new_n1562_;
  assign new_n1564_ = ~\1  & ~new_n1563_;
  assign n308 = \1  | new_n1564_;
  assign new_n1566_ = ~3 & new_n866_;
  assign new_n1567_ = ~3 & ~new_n1566_;
  assign new_n1568_ = 2 & ~new_n1567_;
  assign new_n1569_ = 2 & ~new_n1568_;
  assign new_n1570_ = ~\1  & ~new_n1569_;
  assign n313 = \1  | new_n1570_;
  assign new_n1572_ = ~3 & new_n892_;
  assign new_n1573_ = ~3 & ~new_n1572_;
  assign new_n1574_ = 2 & ~new_n1573_;
  assign new_n1575_ = 2 & ~new_n1574_;
  assign new_n1576_ = ~\1  & ~new_n1575_;
  assign n318 = \1  | new_n1576_;
  assign new_n1578_ = ~3 & new_n918_;
  assign new_n1579_ = ~3 & ~new_n1578_;
  assign new_n1580_ = 2 & ~new_n1579_;
  assign new_n1581_ = 2 & ~new_n1580_;
  assign new_n1582_ = ~\1  & ~new_n1581_;
  assign n323 = \1  | new_n1582_;
  assign new_n1584_ = ~3 & new_n944_;
  assign new_n1585_ = ~3 & ~new_n1584_;
  assign new_n1586_ = 2 & ~new_n1585_;
  assign new_n1587_ = 2 & ~new_n1586_;
  assign new_n1588_ = ~\1  & ~new_n1587_;
  assign n328 = \1  | new_n1588_;
  assign new_n1590_ = ~3 & new_n970_;
  assign new_n1591_ = ~3 & ~new_n1590_;
  assign new_n1592_ = 2 & ~new_n1591_;
  assign new_n1593_ = 2 & ~new_n1592_;
  assign new_n1594_ = ~\1  & ~new_n1593_;
  assign n333 = \1  | new_n1594_;
  assign new_n1596_ = ~3 & new_n996_;
  assign new_n1597_ = ~3 & ~new_n1596_;
  assign new_n1598_ = 2 & ~new_n1597_;
  assign new_n1599_ = 2 & ~new_n1598_;
  assign new_n1600_ = ~\1  & ~new_n1599_;
  assign n338 = \1  | new_n1600_;
  assign new_n1602_ = ~3 & new_n1022_;
  assign new_n1603_ = ~3 & ~new_n1602_;
  assign new_n1604_ = 2 & ~new_n1603_;
  assign new_n1605_ = 2 & ~new_n1604_;
  assign new_n1606_ = ~\1  & ~new_n1605_;
  assign n343 = \1  | new_n1606_;
  assign new_n1608_ = ~3 & new_n1048_;
  assign new_n1609_ = ~3 & ~new_n1608_;
  assign new_n1610_ = 2 & ~new_n1609_;
  assign new_n1611_ = 2 & ~new_n1610_;
  assign new_n1612_ = ~\1  & ~new_n1611_;
  assign n348 = \1  | new_n1612_;
  assign new_n1614_ = ~3 & new_n1074_;
  assign new_n1615_ = ~3 & ~new_n1614_;
  assign new_n1616_ = 2 & ~new_n1615_;
  assign new_n1617_ = 2 & ~new_n1616_;
  assign new_n1618_ = ~\1  & ~new_n1617_;
  assign n353 = \1  | new_n1618_;
  assign new_n1620_ = ~3 & new_n1100_;
  assign new_n1621_ = ~3 & ~new_n1620_;
  assign new_n1622_ = 2 & ~new_n1621_;
  assign new_n1623_ = 2 & ~new_n1622_;
  assign new_n1624_ = ~\1  & ~new_n1623_;
  assign n358 = \1  | new_n1624_;
  assign new_n1626_ = ~3 & new_n1126_;
  assign new_n1627_ = ~3 & ~new_n1626_;
  assign new_n1628_ = 2 & ~new_n1627_;
  assign new_n1629_ = 2 & ~new_n1628_;
  assign new_n1630_ = ~\1  & ~new_n1629_;
  assign n363 = \1  | new_n1630_;
  assign new_n1632_ = ~3 & new_n1152_;
  assign new_n1633_ = ~3 & ~new_n1632_;
  assign new_n1634_ = 2 & ~new_n1633_;
  assign new_n1635_ = 2 & ~new_n1634_;
  assign new_n1636_ = ~\1  & ~new_n1635_;
  assign n368 = \1  | new_n1636_;
  assign new_n1638_ = ~3 & new_n1178_;
  assign new_n1639_ = ~3 & ~new_n1638_;
  assign new_n1640_ = 2 & ~new_n1639_;
  assign new_n1641_ = 2 & ~new_n1640_;
  assign new_n1642_ = ~\1  & ~new_n1641_;
  assign n373 = \1  | new_n1642_;
  assign new_n1644_ = ~3 & new_n1204_;
  assign new_n1645_ = ~3 & ~new_n1644_;
  assign new_n1646_ = 2 & ~new_n1645_;
  assign new_n1647_ = 2 & ~new_n1646_;
  assign new_n1648_ = ~\1  & ~new_n1647_;
  assign n378 = \1  | new_n1648_;
  assign new_n1650_ = ~3 & new_n1230_;
  assign new_n1651_ = ~3 & ~new_n1650_;
  assign new_n1652_ = 2 & ~new_n1651_;
  assign new_n1653_ = 2 & ~new_n1652_;
  assign new_n1654_ = ~\1  & ~new_n1653_;
  assign n383 = \1  | new_n1654_;
  assign new_n1656_ = ~3 & new_n1256_;
  assign new_n1657_ = ~3 & ~new_n1656_;
  assign new_n1658_ = 2 & ~new_n1657_;
  assign new_n1659_ = 2 & ~new_n1658_;
  assign new_n1660_ = ~\1  & ~new_n1659_;
  assign n388 = \1  | new_n1660_;
  assign new_n1662_ = ~3 & new_n1282_;
  assign new_n1663_ = ~3 & ~new_n1662_;
  assign new_n1664_ = 2 & ~new_n1663_;
  assign new_n1665_ = 2 & ~new_n1664_;
  assign new_n1666_ = ~\1  & ~new_n1665_;
  assign n393 = \1  | new_n1666_;
  assign new_n1668_ = ~3 & new_n1308_;
  assign new_n1669_ = ~3 & ~new_n1668_;
  assign new_n1670_ = 2 & ~new_n1669_;
  assign new_n1671_ = 2 & ~new_n1670_;
  assign new_n1672_ = ~\1  & ~new_n1671_;
  assign n398 = \1  | new_n1672_;
  assign new_n1674_ = ~3 & new_n1334_;
  assign new_n1675_ = ~3 & ~new_n1674_;
  assign new_n1676_ = 2 & ~new_n1675_;
  assign new_n1677_ = 2 & ~new_n1676_;
  assign new_n1678_ = ~\1  & ~new_n1677_;
  assign n403 = \1  | new_n1678_;
  assign new_n1680_ = ~3 & new_n1360_;
  assign new_n1681_ = ~3 & ~new_n1680_;
  assign new_n1682_ = 2 & ~new_n1681_;
  assign new_n1683_ = 2 & ~new_n1682_;
  assign new_n1684_ = ~\1  & ~new_n1683_;
  assign n408 = \1  | new_n1684_;
  assign new_n1686_ = ~3 & new_n1386_;
  assign new_n1687_ = ~3 & ~new_n1686_;
  assign new_n1688_ = 2 & ~new_n1687_;
  assign new_n1689_ = 2 & ~new_n1688_;
  assign new_n1690_ = ~\1  & ~new_n1689_;
  assign n413 = \1  | new_n1690_;
  assign new_n1692_ = ~3 & new_n1412_;
  assign new_n1693_ = ~3 & ~new_n1692_;
  assign new_n1694_ = 2 & ~new_n1693_;
  assign new_n1695_ = 2 & ~new_n1694_;
  assign new_n1696_ = ~\1  & ~new_n1695_;
  assign n418 = \1  | new_n1696_;
  assign new_n1698_ = ~3 & new_n1438_;
  assign new_n1699_ = ~3 & ~new_n1698_;
  assign new_n1700_ = 2 & ~new_n1699_;
  assign new_n1701_ = 2 & ~new_n1700_;
  assign new_n1702_ = ~\1  & ~new_n1701_;
  assign n423 = \1  | new_n1702_;
  assign new_n1704_ = ~3 & new_n518_1_;
  assign new_n1705_ = 2 & new_n1704_;
  assign n428 = ~\1  & new_n1705_;
  assign new_n1707_ = ~3 & new_n706_;
  assign new_n1708_ = 2 & new_n1707_;
  assign n433 = ~\1  & new_n1708_;
  assign new_n1710_ = ~3 & new_n732_;
  assign new_n1711_ = 2 & new_n1710_;
  assign n438 = ~\1  & new_n1711_;
  assign new_n1713_ = ~3 & new_n758_;
  assign new_n1714_ = 2 & new_n1713_;
  assign n443 = ~\1  & new_n1714_;
  assign new_n1716_ = ~3 & new_n784_;
  assign new_n1717_ = 2 & new_n1716_;
  assign n448 = ~\1  & new_n1717_;
  assign new_n1719_ = ~3 & new_n810_;
  assign new_n1720_ = 2 & new_n1719_;
  assign n453 = ~\1  & new_n1720_;
  assign new_n1722_ = ~3 & new_n836_;
  assign new_n1723_ = 2 & new_n1722_;
  assign n458 = ~\1  & new_n1723_;
  assign new_n1725_ = ~3 & new_n862_;
  assign new_n1726_ = 2 & new_n1725_;
  assign n463 = ~\1  & new_n1726_;
  assign new_n1728_ = ~3 & new_n888_;
  assign new_n1729_ = 2 & new_n1728_;
  assign n468 = ~\1  & new_n1729_;
  assign new_n1731_ = ~3 & new_n914_;
  assign new_n1732_ = 2 & new_n1731_;
  assign n473 = ~\1  & new_n1732_;
  assign new_n1734_ = ~3 & new_n940_;
  assign new_n1735_ = 2 & new_n1734_;
  assign n478 = ~\1  & new_n1735_;
  assign new_n1737_ = ~3 & new_n966_;
  assign new_n1738_ = 2 & new_n1737_;
  assign n483 = ~\1  & new_n1738_;
  assign new_n1740_ = ~3 & new_n992_;
  assign new_n1741_ = 2 & new_n1740_;
  assign n488 = ~\1  & new_n1741_;
  assign new_n1743_ = ~3 & new_n1018_;
  assign new_n1744_ = 2 & new_n1743_;
  assign n493 = ~\1  & new_n1744_;
  assign new_n1746_ = ~3 & new_n1044_;
  assign new_n1747_ = 2 & new_n1746_;
  assign n498 = ~\1  & new_n1747_;
  assign new_n1749_ = ~3 & new_n1070_;
  assign new_n1750_ = 2 & new_n1749_;
  assign n503 = ~\1  & new_n1750_;
  assign new_n1752_ = ~3 & new_n1096_;
  assign new_n1753_ = 2 & new_n1752_;
  assign n508 = ~\1  & new_n1753_;
  assign new_n1755_ = ~3 & new_n1122_;
  assign new_n1756_ = 2 & new_n1755_;
  assign n513 = ~\1  & new_n1756_;
  assign new_n1758_ = ~3 & new_n1148_;
  assign new_n1759_ = 2 & new_n1758_;
  assign n518 = ~\1  & new_n1759_;
  assign new_n1761_ = ~3 & new_n1174_;
  assign new_n1762_ = 2 & new_n1761_;
  assign n523 = ~\1  & new_n1762_;
  assign new_n1764_ = ~3 & new_n1200_;
  assign new_n1765_ = 2 & new_n1764_;
  assign n528 = ~\1  & new_n1765_;
  assign new_n1767_ = ~3 & new_n1226_;
  assign new_n1768_ = 2 & new_n1767_;
  assign n533 = ~\1  & new_n1768_;
  assign new_n1770_ = ~3 & new_n1252_;
  assign new_n1771_ = 2 & new_n1770_;
  assign n538 = ~\1  & new_n1771_;
  assign new_n1773_ = ~3 & new_n1278_;
  assign new_n1774_ = 2 & new_n1773_;
  assign n543 = ~\1  & new_n1774_;
  assign new_n1776_ = ~3 & new_n1304_;
  assign new_n1777_ = 2 & new_n1776_;
  assign n548 = ~\1  & new_n1777_;
  assign new_n1779_ = ~3 & new_n1330_;
  assign new_n1780_ = 2 & new_n1779_;
  assign n553 = ~\1  & new_n1780_;
  assign new_n1782_ = ~3 & new_n1356_;
  assign new_n1783_ = 2 & new_n1782_;
  assign n558 = ~\1  & new_n1783_;
  assign new_n1785_ = ~3 & new_n1382_;
  assign new_n1786_ = 2 & new_n1785_;
  assign n563 = ~\1  & new_n1786_;
  assign new_n1788_ = ~3 & new_n1408_;
  assign new_n1789_ = 2 & new_n1788_;
  assign n568 = ~\1  & new_n1789_;
  assign new_n1791_ = ~3 & new_n1434_;
  assign new_n1792_ = 2 & new_n1791_;
  assign n573 = ~\1  & new_n1792_;
  always @ (posedge clock) begin
    34 <= n128;
    35 <= n133;
    36 <= n138;
    37 <= n143;
    38 <= n148;
    39 <= n153;
    40 <= n158;
    41 <= n163;
    42 <= n168;
    43 <= n173;
    44 <= n178;
    45 <= n183;
    46 <= n188;
    47 <= n193;
    48 <= n198;
    49 <= n203;
    50 <= n208;
    51 <= n213;
    52 <= n218;
    53 <= n223;
    54 <= n228;
    55 <= n233;
    56 <= n238;
    57 <= n243;
    58 <= n248;
    59 <= n253;
    60 <= n258;
    61 <= n263;
    62 <= n268;
    63 <= n273;
    64 <= n278;
    65 <= n283;
    66 <= n288;
    67 <= n293;
    68 <= n298;
    69 <= n303;
    70 <= n308;
    71 <= n313;
    72 <= n318;
    73 <= n323;
    74 <= n328;
    75 <= n333;
    76 <= n338;
    77 <= n343;
    78 <= n348;
    79 <= n353;
    80 <= n358;
    81 <= n363;
    82 <= n368;
    83 <= n373;
    84 <= n378;
    85 <= n383;
    86 <= n388;
    87 <= n393;
    88 <= n398;
    89 <= n403;
    90 <= n408;
    91 <= n413;
    92 <= n418;
    93 <= n423;
    94 <= n428;
    95 <= n433;
    96 <= n438;
    97 <= n443;
    98 <= n448;
    99 <= n453;
    100 <= n458;
    101 <= n463;
    102 <= n468;
    103 <= n473;
    104 <= n478;
    105 <= n483;
    106 <= n488;
    107 <= n493;
    108 <= n498;
    109 <= n503;
    110 <= n508;
    111 <= n513;
    112 <= n518;
    113 <= n523;
    114 <= n528;
    115 <= n533;
    116 <= n538;
    117 <= n543;
    118 <= n548;
    119 <= n553;
    120 <= n558;
    121 <= n563;
    122 <= n568;
    123 <= n573;
  end
  initial begin
    64 <= 1'b1;
    65 <= 1'b1;
    66 <= 1'b1;
    67 <= 1'b1;
    68 <= 1'b1;
    69 <= 1'b1;
    70 <= 1'b1;
    71 <= 1'b1;
    72 <= 1'b1;
    73 <= 1'b1;
    74 <= 1'b1;
    75 <= 1'b1;
    76 <= 1'b1;
    77 <= 1'b1;
    78 <= 1'b1;
    79 <= 1'b1;
    80 <= 1'b1;
    81 <= 1'b1;
    82 <= 1'b1;
    83 <= 1'b1;
    84 <= 1'b1;
    85 <= 1'b1;
    86 <= 1'b1;
    87 <= 1'b1;
    88 <= 1'b1;
    89 <= 1'b1;
    90 <= 1'b1;
    91 <= 1'b1;
    92 <= 1'b1;
    93 <= 1'b1;
    94 <= 1'b0;
    95 <= 1'b0;
    96 <= 1'b0;
    97 <= 1'b0;
    98 <= 1'b0;
    99 <= 1'b0;
    100 <= 1'b0;
    101 <= 1'b0;
    102 <= 1'b0;
    103 <= 1'b0;
    104 <= 1'b0;
    105 <= 1'b0;
    106 <= 1'b0;
    107 <= 1'b0;
    108 <= 1'b0;
    109 <= 1'b0;
    110 <= 1'b0;
    111 <= 1'b0;
    112 <= 1'b0;
    113 <= 1'b0;
    114 <= 1'b0;
    115 <= 1'b0;
    116 <= 1'b0;
    117 <= 1'b0;
    118 <= 1'b0;
    119 <= 1'b0;
    120 <= 1'b0;
    121 <= 1'b0;
    122 <= 1'b0;
    123 <= 1'b0;
  end
endmodule

