module top ( 
    _1gat_0_, _11gat_3_, _17gat_5_, _95gat_29_, _112gat_34_, _4gat_1_,
    _30gat_9_, _27gat_8_, _8gat_2_, _40gat_12_, _47gat_14_, _69gat_21_,
    _73gat_22_, _89gat_27_, _53gat_16_, _115gat_35_, _37gat_11_,
    _63gat_19_, _99gat_30_, _79gat_24_, _14gat_4_, _102gat_31_, _24gat_7_,
    _82gat_25_, _66gat_20_, _43gat_13_, _92gat_28_, _76gat_23_, _86gat_26_,
    _50gat_15_, _108gat_33_, _21gat_6_, _60gat_18_, _56gat_17_,
    _105gat_32_, _34gat_10_,
    _421gat_188_, _329gat_133_, _223gat_84_, _370gat_163_, _431gat_194_,
    _432gat_195_, _430gat_193_  );
  input  _1gat_0_, _11gat_3_, _17gat_5_, _95gat_29_, _112gat_34_,
    _4gat_1_, _30gat_9_, _27gat_8_, _8gat_2_, _40gat_12_, _47gat_14_,
    _69gat_21_, _73gat_22_, _89gat_27_, _53gat_16_, _115gat_35_,
    _37gat_11_, _63gat_19_, _99gat_30_, _79gat_24_, _14gat_4_, _102gat_31_,
    _24gat_7_, _82gat_25_, _66gat_20_, _43gat_13_, _92gat_28_, _76gat_23_,
    _86gat_26_, _50gat_15_, _108gat_33_, _21gat_6_, _60gat_18_, _56gat_17_,
    _105gat_32_, _34gat_10_;
  output _421gat_188_, _329gat_133_, _223gat_84_, _370gat_163_, _431gat_194_,
    _432gat_195_, _430gat_193_;
  wire new_n44_, new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_,
    new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_,
    new_n58_, new_n59_, new_n60_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n253_, new_n254_;
  assign new_n44_ = ~_47gat_14_ & _43gat_13_;
  assign new_n45_ = ~_37gat_11_ & _43gat_13_;
  assign new_n46_ = ~_50gat_15_ & _56gat_17_;
  assign new_n47_ = ~_11gat_3_ & _17gat_5_;
  assign new_n48_ = _30gat_9_ & ~_24gat_7_;
  assign new_n49_ = ~_1gat_0_ & _4gat_1_;
  assign new_n50_ = _95gat_29_ & ~_89gat_27_;
  assign new_n51_ = ~_102gat_31_ & _108gat_33_;
  assign new_n52_ = _69gat_21_ & ~_63gat_19_;
  assign new_n53_ = _82gat_25_ & ~_76gat_23_;
  assign new_n54_ = ~new_n45_ & ~new_n46_;
  assign new_n55_ = ~new_n47_ & new_n54_;
  assign new_n56_ = ~new_n48_ & new_n55_;
  assign new_n57_ = ~new_n49_ & new_n56_;
  assign new_n58_ = ~new_n50_ & new_n57_;
  assign new_n59_ = ~new_n51_ & new_n58_;
  assign new_n60_ = ~new_n52_ & new_n59_;
  assign _223gat_84_ = new_n53_ | ~new_n60_;
  assign new_n62_ = new_n45_ & _223gat_84_;
  assign new_n63_ = ~new_n45_ & ~_223gat_84_;
  assign new_n64_ = ~new_n62_ & ~new_n63_;
  assign new_n65_ = new_n44_ & ~new_n64_;
  assign new_n66_ = ~_60gat_18_ & _56gat_17_;
  assign new_n67_ = new_n46_ & _223gat_84_;
  assign new_n68_ = ~new_n46_ & ~_223gat_84_;
  assign new_n69_ = ~new_n67_ & ~new_n68_;
  assign new_n70_ = new_n66_ & ~new_n69_;
  assign new_n71_ = _17gat_5_ & ~_21gat_6_;
  assign new_n72_ = new_n47_ & _223gat_84_;
  assign new_n73_ = ~new_n47_ & ~_223gat_84_;
  assign new_n74_ = ~new_n72_ & ~new_n73_;
  assign new_n75_ = new_n71_ & ~new_n74_;
  assign new_n76_ = _30gat_9_ & ~_34gat_10_;
  assign new_n77_ = new_n48_ & _223gat_84_;
  assign new_n78_ = ~new_n48_ & ~_223gat_84_;
  assign new_n79_ = ~new_n77_ & ~new_n78_;
  assign new_n80_ = new_n76_ & ~new_n79_;
  assign new_n81_ = _4gat_1_ & ~_8gat_2_;
  assign new_n82_ = new_n49_ & _223gat_84_;
  assign new_n83_ = ~new_n49_ & ~_223gat_84_;
  assign new_n84_ = ~new_n82_ & ~new_n83_;
  assign new_n85_ = new_n81_ & ~new_n84_;
  assign new_n86_ = _95gat_29_ & ~_99gat_30_;
  assign new_n87_ = new_n50_ & _223gat_84_;
  assign new_n88_ = ~new_n50_ & ~_223gat_84_;
  assign new_n89_ = ~new_n87_ & ~new_n88_;
  assign new_n90_ = new_n86_ & ~new_n89_;
  assign new_n91_ = ~_112gat_34_ & _108gat_33_;
  assign new_n92_ = new_n51_ & _223gat_84_;
  assign new_n93_ = ~new_n51_ & ~_223gat_84_;
  assign new_n94_ = ~new_n92_ & ~new_n93_;
  assign new_n95_ = new_n91_ & ~new_n94_;
  assign new_n96_ = _69gat_21_ & ~_73gat_22_;
  assign new_n97_ = new_n52_ & _223gat_84_;
  assign new_n98_ = ~new_n52_ & ~_223gat_84_;
  assign new_n99_ = ~new_n97_ & ~new_n98_;
  assign new_n100_ = new_n96_ & ~new_n99_;
  assign new_n101_ = _82gat_25_ & ~_86gat_26_;
  assign new_n102_ = new_n53_ & _223gat_84_;
  assign new_n103_ = ~new_n53_ & ~_223gat_84_;
  assign new_n104_ = ~new_n102_ & ~new_n103_;
  assign new_n105_ = new_n101_ & ~new_n104_;
  assign new_n106_ = ~new_n65_ & ~new_n70_;
  assign new_n107_ = ~new_n75_ & new_n106_;
  assign new_n108_ = ~new_n80_ & new_n107_;
  assign new_n109_ = ~new_n85_ & new_n108_;
  assign new_n110_ = ~new_n90_ & new_n109_;
  assign new_n111_ = ~new_n95_ & new_n110_;
  assign new_n112_ = ~new_n100_ & new_n111_;
  assign _329gat_133_ = new_n105_ | ~new_n112_;
  assign new_n114_ = _60gat_18_ & _329gat_133_;
  assign new_n115_ = ~_53gat_16_ & _43gat_13_;
  assign new_n116_ = ~new_n64_ & new_n115_;
  assign new_n117_ = new_n65_ & _329gat_133_;
  assign new_n118_ = ~new_n65_ & ~_329gat_133_;
  assign new_n119_ = ~new_n117_ & ~new_n118_;
  assign new_n120_ = new_n116_ & ~new_n119_;
  assign new_n121_ = ~_66gat_20_ & _56gat_17_;
  assign new_n122_ = ~new_n69_ & new_n121_;
  assign new_n123_ = new_n70_ & _329gat_133_;
  assign new_n124_ = ~new_n70_ & ~_329gat_133_;
  assign new_n125_ = ~new_n123_ & ~new_n124_;
  assign new_n126_ = new_n122_ & ~new_n125_;
  assign new_n127_ = _17gat_5_ & ~_27gat_8_;
  assign new_n128_ = ~new_n74_ & new_n127_;
  assign new_n129_ = new_n75_ & _329gat_133_;
  assign new_n130_ = ~new_n75_ & ~_329gat_133_;
  assign new_n131_ = ~new_n129_ & ~new_n130_;
  assign new_n132_ = new_n128_ & ~new_n131_;
  assign new_n133_ = _30gat_9_ & ~_40gat_12_;
  assign new_n134_ = ~new_n79_ & new_n133_;
  assign new_n135_ = new_n80_ & _329gat_133_;
  assign new_n136_ = ~new_n80_ & ~_329gat_133_;
  assign new_n137_ = ~new_n135_ & ~new_n136_;
  assign new_n138_ = new_n134_ & ~new_n137_;
  assign new_n139_ = _4gat_1_ & ~_14gat_4_;
  assign new_n140_ = ~new_n84_ & new_n139_;
  assign new_n141_ = new_n85_ & _329gat_133_;
  assign new_n142_ = ~new_n85_ & ~_329gat_133_;
  assign new_n143_ = ~new_n141_ & ~new_n142_;
  assign new_n144_ = new_n140_ & ~new_n143_;
  assign new_n145_ = _95gat_29_ & ~_105gat_32_;
  assign new_n146_ = ~new_n89_ & new_n145_;
  assign new_n147_ = new_n90_ & _329gat_133_;
  assign new_n148_ = ~new_n90_ & ~_329gat_133_;
  assign new_n149_ = ~new_n147_ & ~new_n148_;
  assign new_n150_ = new_n146_ & ~new_n149_;
  assign new_n151_ = ~_115gat_35_ & _108gat_33_;
  assign new_n152_ = ~new_n94_ & new_n151_;
  assign new_n153_ = new_n95_ & _329gat_133_;
  assign new_n154_ = ~new_n95_ & ~_329gat_133_;
  assign new_n155_ = ~new_n153_ & ~new_n154_;
  assign new_n156_ = new_n152_ & ~new_n155_;
  assign new_n157_ = _69gat_21_ & ~_79gat_24_;
  assign new_n158_ = ~new_n99_ & new_n157_;
  assign new_n159_ = new_n100_ & _329gat_133_;
  assign new_n160_ = ~new_n100_ & ~_329gat_133_;
  assign new_n161_ = ~new_n159_ & ~new_n160_;
  assign new_n162_ = new_n158_ & ~new_n161_;
  assign new_n163_ = _82gat_25_ & ~_92gat_28_;
  assign new_n164_ = ~new_n104_ & new_n163_;
  assign new_n165_ = new_n105_ & _329gat_133_;
  assign new_n166_ = ~new_n105_ & ~_329gat_133_;
  assign new_n167_ = ~new_n165_ & ~new_n166_;
  assign new_n168_ = new_n164_ & ~new_n167_;
  assign new_n169_ = ~new_n120_ & ~new_n126_;
  assign new_n170_ = ~new_n132_ & new_n169_;
  assign new_n171_ = ~new_n138_ & new_n170_;
  assign new_n172_ = ~new_n144_ & new_n171_;
  assign new_n173_ = ~new_n150_ & new_n172_;
  assign new_n174_ = ~new_n156_ & new_n173_;
  assign new_n175_ = ~new_n162_ & new_n174_;
  assign _370gat_163_ = new_n168_ | ~new_n175_;
  assign new_n177_ = _66gat_20_ & _370gat_163_;
  assign new_n178_ = _50gat_15_ & _223gat_84_;
  assign new_n179_ = _56gat_17_ & ~new_n114_;
  assign new_n180_ = ~new_n177_ & new_n179_;
  assign new_n181_ = ~new_n178_ & new_n180_;
  assign new_n182_ = _73gat_22_ & _329gat_133_;
  assign new_n183_ = _79gat_24_ & _370gat_163_;
  assign new_n184_ = _63gat_19_ & _223gat_84_;
  assign new_n185_ = _69gat_21_ & ~new_n182_;
  assign new_n186_ = ~new_n183_ & new_n185_;
  assign new_n187_ = ~new_n184_ & new_n186_;
  assign new_n188_ = _34gat_10_ & _329gat_133_;
  assign new_n189_ = _40gat_12_ & _370gat_163_;
  assign new_n190_ = _24gat_7_ & _223gat_84_;
  assign new_n191_ = _30gat_9_ & ~new_n188_;
  assign new_n192_ = ~new_n189_ & new_n191_;
  assign new_n193_ = ~new_n190_ & new_n192_;
  assign new_n194_ = _47gat_14_ & _329gat_133_;
  assign new_n195_ = _53gat_16_ & _370gat_163_;
  assign new_n196_ = _37gat_11_ & _223gat_84_;
  assign new_n197_ = _43gat_13_ & ~new_n194_;
  assign new_n198_ = ~new_n195_ & new_n197_;
  assign new_n199_ = ~new_n196_ & new_n198_;
  assign new_n200_ = _21gat_6_ & _329gat_133_;
  assign new_n201_ = _27gat_8_ & _370gat_163_;
  assign new_n202_ = _11gat_3_ & _223gat_84_;
  assign new_n203_ = _17gat_5_ & ~new_n200_;
  assign new_n204_ = ~new_n201_ & new_n203_;
  assign new_n205_ = ~new_n202_ & new_n204_;
  assign new_n206_ = _112gat_34_ & _329gat_133_;
  assign new_n207_ = _115gat_35_ & _370gat_163_;
  assign new_n208_ = _102gat_31_ & _223gat_84_;
  assign new_n209_ = _108gat_33_ & ~new_n206_;
  assign new_n210_ = ~new_n207_ & new_n209_;
  assign new_n211_ = ~new_n208_ & new_n210_;
  assign new_n212_ = _86gat_26_ & _329gat_133_;
  assign new_n213_ = _92gat_28_ & _370gat_163_;
  assign new_n214_ = _76gat_23_ & _223gat_84_;
  assign new_n215_ = _82gat_25_ & ~new_n212_;
  assign new_n216_ = ~new_n213_ & new_n215_;
  assign new_n217_ = ~new_n214_ & new_n216_;
  assign new_n218_ = _99gat_30_ & _329gat_133_;
  assign new_n219_ = _105gat_32_ & _370gat_163_;
  assign new_n220_ = _89gat_27_ & _223gat_84_;
  assign new_n221_ = _95gat_29_ & ~new_n218_;
  assign new_n222_ = ~new_n219_ & new_n221_;
  assign new_n223_ = ~new_n220_ & new_n222_;
  assign new_n224_ = ~new_n181_ & ~new_n187_;
  assign new_n225_ = ~new_n193_ & new_n224_;
  assign new_n226_ = ~new_n199_ & new_n225_;
  assign new_n227_ = ~new_n205_ & new_n226_;
  assign new_n228_ = ~new_n211_ & new_n227_;
  assign new_n229_ = ~new_n217_ & new_n228_;
  assign new_n230_ = ~new_n223_ & new_n229_;
  assign new_n231_ = _14gat_4_ & _370gat_163_;
  assign new_n232_ = _1gat_0_ & _223gat_84_;
  assign new_n233_ = _8gat_2_ & _329gat_133_;
  assign new_n234_ = ~new_n231_ & ~new_n232_;
  assign new_n235_ = ~new_n233_ & new_n234_;
  assign new_n236_ = _4gat_1_ & new_n235_;
  assign _421gat_188_ = ~new_n230_ & ~new_n236_;
  assign new_n238_ = ~new_n199_ & new_n217_;
  assign new_n239_ = ~new_n181_ & new_n238_;
  assign new_n240_ = ~new_n181_ & ~new_n199_;
  assign new_n241_ = new_n187_ & new_n240_;
  assign new_n242_ = ~new_n193_ & new_n241_;
  assign new_n243_ = ~new_n193_ & ~new_n239_;
  assign new_n244_ = ~new_n242_ & new_n243_;
  assign _431gat_194_ = new_n205_ | ~new_n244_;
  assign new_n246_ = ~new_n199_ & new_n223_;
  assign new_n247_ = ~new_n217_ & new_n246_;
  assign new_n248_ = ~new_n193_ & new_n247_;
  assign new_n249_ = ~new_n193_ & new_n199_;
  assign new_n250_ = ~new_n248_ & ~new_n249_;
  assign new_n251_ = ~new_n242_ & new_n250_;
  assign _432gat_195_ = new_n205_ | ~new_n251_;
  assign new_n253_ = ~new_n181_ & ~new_n193_;
  assign new_n254_ = ~new_n249_ & new_n253_;
  assign _430gat_193_ = new_n205_ | ~new_n254_;
endmodule

