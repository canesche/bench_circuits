module top ( 
    p_4_1_, p_26_9_, p_130_58_, p_53_19_, p_64_22_, p_67_23_, p_91_35_,
    p_94_36_, p_136_62_, p_173_76_, p_293_112_, p_545_150_, p_2174_161_,
    p_3717_169_, p_25_8_, p_106_40_, p_14_3_, p_52_18_, p_113_43_,
    p_117_47_, p_534_149_, p_24_7_, p_272_105_, p_302_114_, p_4091_175_,
    p_61_21_, p_100_38_, p_170_75_, p_210_89_, p_226_93_, p_373_133_,
    p_23_6_, p_167_74_, p_206_87_, p_400_137_, p_457_142_, p_1694_160_,
    p_4090_174_, p_11_2_, p_123_53_, p_315_117_, p_514_147_, p_1690_158_,
    p_4115_177_, p_109_41_, p_257_102_, p_323_119_, p_435_140_, p_559_154_,
    p_31_11_, p_34_12_, p_114_44_, p_118_48_, p_120_50_, p_176_77_,
    p_324_120_, p_552_152_, p_20_5_, p_40_14_, p_140_64_, p_549_151_,
    p_4092_176_, p_146_67_, p_242_97_, p_374_134_, p_4089_173_, p_203_86_,
    p_254_101_, p_308_116_, p_331_121_, p_37_13_, p_97_37_, p_127_55_,
    p_179_78_, p_468_143_, p_3552_168_, p_4088_172_, p_1_0_, p_182_79_,
    p_200_85_, p_233_94_, p_273_106_, p_490_145_, p_3550_167_, p_17_4_,
    p_137_63_, p_2824_163_, p_4087_171_, p_49_17_, p_70_24_, p_86_32_,
    p_87_33_, p_88_34_, p_217_90_, p_251_100_, p_351_127_, p_358_128_,
    p_369_131_, p_3173_164_, p_145_66_, p_241_96_, p_341_125_, p_348_126_,
    p_411_138_, p_46_16_, p_73_25_, p_83_31_, p_141_65_, p_152_69_,
    p_191_82_, p_234_95_, p_338_124_, p_121_51_, p_158_71_, p_248_99_,
    p_264_103_, p_361_129_, p_389_136_, p_446_141_, p_43_15_, p_76_26_,
    p_164_73_, p_556_153_, p_3548_166_, p_280_107_, p_82_30_, p_307_115_,
    p_335_123_, p_115_45_, p_128_56_, p_149_68_, p_245_98_, p_386_135_,
    p_3546_165_, p_131_59_, p_209_88_, p_218_91_, p_422_139_, p_1497_156_,
    p_1689_157_, p_27_10_, p_103_39_, p_112_42_, p_116_46_, p_122_52_,
    p_185_80_, p_265_104_, p_562_155_, p_1691_159_, p_79_27_, p_197_84_,
    p_299_113_, p_332_122_, p_503_146_, p_126_54_, p_135_61_, p_292_111_,
    p_194_83_, p_289_110_, p_366_130_, p_479_144_, p_2358_162_, p_80_28_,
    p_129_57_, p_188_81_, p_316_118_, p_54_20_, p_161_72_, p_523_148_,
    p_81_29_, p_119_49_, p_132_60_, p_155_70_, p_225_92_, p_281_108_,
    p_288_109_, p_372_132_, p_3724_170_,
    p_591_1894_, p_604_223_, p_664_2223_, p_690_2484_, p_699_2227_,
    p_618_1925_, p_588_1696_, p_615_1750_, p_688_2317_, p_704_1281_,
    p_818_2273_, p_869_2181_, p_973_202_, p_593_733_, p_600_259_,
    p_611_275_, p_648_2295_, p_822_1933_, p_757_2190_, p_722_2131_,
    p_802_2183_, p_1000_2168_, p_606_407_, p_682_2296_, p_792_2188_,
    p_838_2064_, p_603_225_, p_921_664_, p_629_1926_, p_892_408_,
    p_949_852_, p_612_263_, p_772_2299_, p_797_2191_, p_661_2178_,
    p_727_2298_, p_849_219_, p_939_853_, p_598_1623_, p_634_665_,
    p_636_1280_, p_742_2238_, p_767_2479_, p_836_2128_, p_693_2179_,
    p_702_2228_, p_807_2480_, p_594_224_, p_654_2315_, p_658_2483_,
    p_820_1283_, p_861_2070_, p_875_2125_, p_978_851_, p_685_2316_,
    p_815_627_, p_834_2123_, p_882_2456_, p_926_624_, p_621_1893_,
    p_676_2229_, p_667_2224_, p_696_2226_, p_787_2186_, p_877_2126_,
    p_1002_1920_, p_1004_1977_, p_670_2225_, p_712_2297_, p_298_299_,
    p_715_1278_, p_809_655_, p_843_2455_, p_867_2237_, p_602_222_,
    p_859_2132_, p_863_2276_, p_623_2152_, p_810_356_, p_642_2222_,
    p_777_2278_, p_830_2182_, p_626_1752_, p_632_1692_, p_645_2271_,
    p_679_2272_, p_707_1277_, p_737_2279_, p_782_2239_, p_850_217_,
    p_717_1282_, p_747_2187_, p_826_2275_, p_845_845_, p_871_2127_,
    p_585_2236_, p_865_2277_, p_673_1276_, p_887_528_, p_923_619_,
    p_144_354_, p_732_2300_, p_854_2268_, p_873_2124_, p_889_734_,
    p_599_269_, p_752_2189_, p_610_1519_, p_824_2274_, p_851_218_,
    p_813_2260_, p_832_2133_, p_848_330_, p_993_850_, p_575_2240_,
    p_601_220_, p_639_1275_, p_651_2314_, p_656_621_, p_762_2184_,
    p_828_2233_, p_847_465_, p_998_2163_  );
  input  p_4_1_, p_26_9_, p_130_58_, p_53_19_, p_64_22_, p_67_23_,
    p_91_35_, p_94_36_, p_136_62_, p_173_76_, p_293_112_, p_545_150_,
    p_2174_161_, p_3717_169_, p_25_8_, p_106_40_, p_14_3_, p_52_18_,
    p_113_43_, p_117_47_, p_534_149_, p_24_7_, p_272_105_, p_302_114_,
    p_4091_175_, p_61_21_, p_100_38_, p_170_75_, p_210_89_, p_226_93_,
    p_373_133_, p_23_6_, p_167_74_, p_206_87_, p_400_137_, p_457_142_,
    p_1694_160_, p_4090_174_, p_11_2_, p_123_53_, p_315_117_, p_514_147_,
    p_1690_158_, p_4115_177_, p_109_41_, p_257_102_, p_323_119_,
    p_435_140_, p_559_154_, p_31_11_, p_34_12_, p_114_44_, p_118_48_,
    p_120_50_, p_176_77_, p_324_120_, p_552_152_, p_20_5_, p_40_14_,
    p_140_64_, p_549_151_, p_4092_176_, p_146_67_, p_242_97_, p_374_134_,
    p_4089_173_, p_203_86_, p_254_101_, p_308_116_, p_331_121_, p_37_13_,
    p_97_37_, p_127_55_, p_179_78_, p_468_143_, p_3552_168_, p_4088_172_,
    p_1_0_, p_182_79_, p_200_85_, p_233_94_, p_273_106_, p_490_145_,
    p_3550_167_, p_17_4_, p_137_63_, p_2824_163_, p_4087_171_, p_49_17_,
    p_70_24_, p_86_32_, p_87_33_, p_88_34_, p_217_90_, p_251_100_,
    p_351_127_, p_358_128_, p_369_131_, p_3173_164_, p_145_66_, p_241_96_,
    p_341_125_, p_348_126_, p_411_138_, p_46_16_, p_73_25_, p_83_31_,
    p_141_65_, p_152_69_, p_191_82_, p_234_95_, p_338_124_, p_121_51_,
    p_158_71_, p_248_99_, p_264_103_, p_361_129_, p_389_136_, p_446_141_,
    p_43_15_, p_76_26_, p_164_73_, p_556_153_, p_3548_166_, p_280_107_,
    p_82_30_, p_307_115_, p_335_123_, p_115_45_, p_128_56_, p_149_68_,
    p_245_98_, p_386_135_, p_3546_165_, p_131_59_, p_209_88_, p_218_91_,
    p_422_139_, p_1497_156_, p_1689_157_, p_27_10_, p_103_39_, p_112_42_,
    p_116_46_, p_122_52_, p_185_80_, p_265_104_, p_562_155_, p_1691_159_,
    p_79_27_, p_197_84_, p_299_113_, p_332_122_, p_503_146_, p_126_54_,
    p_135_61_, p_292_111_, p_194_83_, p_289_110_, p_366_130_, p_479_144_,
    p_2358_162_, p_80_28_, p_129_57_, p_188_81_, p_316_118_, p_54_20_,
    p_161_72_, p_523_148_, p_81_29_, p_119_49_, p_132_60_, p_155_70_,
    p_225_92_, p_281_108_, p_288_109_, p_372_132_, p_3724_170_;
  output p_591_1894_, p_604_223_, p_664_2223_, p_690_2484_, p_699_2227_,
    p_618_1925_, p_588_1696_, p_615_1750_, p_688_2317_, p_704_1281_,
    p_818_2273_, p_869_2181_, p_973_202_, p_593_733_, p_600_259_,
    p_611_275_, p_648_2295_, p_822_1933_, p_757_2190_, p_722_2131_,
    p_802_2183_, p_1000_2168_, p_606_407_, p_682_2296_, p_792_2188_,
    p_838_2064_, p_603_225_, p_921_664_, p_629_1926_, p_892_408_,
    p_949_852_, p_612_263_, p_772_2299_, p_797_2191_, p_661_2178_,
    p_727_2298_, p_849_219_, p_939_853_, p_598_1623_, p_634_665_,
    p_636_1280_, p_742_2238_, p_767_2479_, p_836_2128_, p_693_2179_,
    p_702_2228_, p_807_2480_, p_594_224_, p_654_2315_, p_658_2483_,
    p_820_1283_, p_861_2070_, p_875_2125_, p_978_851_, p_685_2316_,
    p_815_627_, p_834_2123_, p_882_2456_, p_926_624_, p_621_1893_,
    p_676_2229_, p_667_2224_, p_696_2226_, p_787_2186_, p_877_2126_,
    p_1002_1920_, p_1004_1977_, p_670_2225_, p_712_2297_, p_298_299_,
    p_715_1278_, p_809_655_, p_843_2455_, p_867_2237_, p_602_222_,
    p_859_2132_, p_863_2276_, p_623_2152_, p_810_356_, p_642_2222_,
    p_777_2278_, p_830_2182_, p_626_1752_, p_632_1692_, p_645_2271_,
    p_679_2272_, p_707_1277_, p_737_2279_, p_782_2239_, p_850_217_,
    p_717_1282_, p_747_2187_, p_826_2275_, p_845_845_, p_871_2127_,
    p_585_2236_, p_865_2277_, p_673_1276_, p_887_528_, p_923_619_,
    p_144_354_, p_732_2300_, p_854_2268_, p_873_2124_, p_889_734_,
    p_599_269_, p_752_2189_, p_610_1519_, p_824_2274_, p_851_218_,
    p_813_2260_, p_832_2133_, p_848_330_, p_993_850_, p_575_2240_,
    p_601_220_, p_639_1275_, p_651_2314_, p_656_621_, p_762_2184_,
    p_828_2233_, p_847_465_, p_998_2163_;
  wire new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1159_, new_n1160_, new_n1161_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1180_, new_n1181_, new_n1182_, new_n1183_,
    new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_,
    new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_,
    new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1380_, new_n1381_, new_n1382_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1433_, new_n1434_,
    new_n1435_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1477_, new_n1478_, new_n1479_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1492_, new_n1493_, new_n1494_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1542_, new_n1543_, new_n1544_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_,
    new_n1696_, new_n1697_, new_n1698_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1761_, new_n1762_, new_n1764_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1769_, new_n1770_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1800_, new_n1801_, new_n1802_, new_n1803_,
    new_n1804_, new_n1805_, new_n1806_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1855_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_, new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_,
    new_n1869_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1879_, new_n1880_, new_n1881_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1898_,
    new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_,
    new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_;
  assign new_n302_ = p_264_103_ & p_335_123_;
  assign new_n303_ = p_257_102_ & ~p_335_123_;
  assign new_n304_ = ~new_n302_ & ~new_n303_;
  assign new_n305_ = p_389_136_ & new_n304_;
  assign new_n306_ = ~p_389_136_ & ~new_n304_;
  assign new_n307_ = ~new_n305_ & ~new_n306_;
  assign new_n308_ = p_241_96_ & p_335_123_;
  assign new_n309_ = p_234_95_ & ~p_335_123_;
  assign new_n310_ = ~new_n308_ & ~new_n309_;
  assign new_n311_ = p_435_140_ & new_n310_;
  assign new_n312_ = ~p_435_140_ & ~new_n310_;
  assign new_n313_ = ~new_n311_ & ~new_n312_;
  assign new_n314_ = p_280_107_ & p_335_123_;
  assign new_n315_ = p_273_106_ & ~p_335_123_;
  assign new_n316_ = ~new_n314_ & ~new_n315_;
  assign new_n317_ = p_411_138_ & ~new_n316_;
  assign new_n318_ = p_272_105_ & p_335_123_;
  assign new_n319_ = ~p_335_123_ & p_265_104_;
  assign new_n320_ = ~new_n318_ & ~new_n319_;
  assign new_n321_ = p_400_137_ & new_n320_;
  assign new_n322_ = ~p_400_137_ & ~new_n320_;
  assign new_n323_ = ~new_n321_ & ~new_n322_;
  assign new_n324_ = ~new_n307_ & ~new_n313_;
  assign new_n325_ = new_n317_ & new_n324_;
  assign new_n326_ = ~new_n323_ & new_n325_;
  assign new_n327_ = p_335_123_ & p_288_109_;
  assign new_n328_ = ~p_335_123_ & p_281_108_;
  assign new_n329_ = ~new_n327_ & ~new_n328_;
  assign new_n330_ = p_374_134_ & ~new_n329_;
  assign new_n331_ = p_411_138_ & new_n316_;
  assign new_n332_ = ~p_411_138_ & ~new_n316_;
  assign new_n333_ = ~new_n331_ & ~new_n332_;
  assign new_n334_ = ~new_n307_ & new_n330_;
  assign new_n335_ = ~new_n323_ & new_n334_;
  assign new_n336_ = ~new_n313_ & new_n335_;
  assign new_n337_ = ~new_n333_ & new_n336_;
  assign new_n338_ = p_389_136_ & ~new_n304_;
  assign new_n339_ = ~new_n313_ & new_n338_;
  assign new_n340_ = p_400_137_ & ~new_n320_;
  assign new_n341_ = ~new_n313_ & new_n340_;
  assign new_n342_ = ~new_n307_ & new_n341_;
  assign new_n343_ = p_435_140_ & ~new_n310_;
  assign new_n344_ = ~new_n326_ & ~new_n337_;
  assign new_n345_ = ~new_n339_ & new_n344_;
  assign new_n346_ = ~new_n342_ & new_n345_;
  assign new_n347_ = ~new_n343_ & new_n346_;
  assign new_n348_ = p_335_123_ & p_209_88_;
  assign new_n349_ = p_206_87_ & ~p_335_123_;
  assign new_n350_ = ~new_n348_ & ~new_n349_;
  assign new_n351_ = p_446_141_ & new_n350_;
  assign new_n352_ = ~p_446_141_ & ~new_n350_;
  assign new_n353_ = ~new_n351_ & ~new_n352_;
  assign new_n354_ = p_335_123_ & p_225_92_;
  assign new_n355_ = ~p_335_123_ & p_218_91_;
  assign new_n356_ = ~new_n354_ & ~new_n355_;
  assign new_n357_ = p_468_143_ & new_n356_;
  assign new_n358_ = ~p_468_143_ & ~new_n356_;
  assign new_n359_ = ~new_n357_ & ~new_n358_;
  assign new_n360_ = p_217_90_ & p_335_123_;
  assign new_n361_ = p_210_89_ & ~p_335_123_;
  assign new_n362_ = ~new_n360_ & ~new_n361_;
  assign new_n363_ = p_457_142_ & new_n362_;
  assign new_n364_ = ~p_457_142_ & ~new_n362_;
  assign new_n365_ = ~new_n363_ & ~new_n364_;
  assign new_n366_ = p_233_94_ & p_335_123_;
  assign new_n367_ = p_226_93_ & ~p_335_123_;
  assign new_n368_ = ~new_n366_ & ~new_n367_;
  assign new_n369_ = p_422_139_ & new_n368_;
  assign new_n370_ = ~p_422_139_ & ~new_n368_;
  assign new_n371_ = ~new_n369_ & ~new_n370_;
  assign new_n372_ = ~new_n353_ & ~new_n359_;
  assign new_n373_ = ~new_n365_ & new_n372_;
  assign new_n374_ = ~new_n371_ & new_n373_;
  assign new_n375_ = ~new_n347_ & new_n374_;
  assign new_n376_ = p_422_139_ & ~new_n368_;
  assign new_n377_ = ~new_n353_ & ~new_n365_;
  assign new_n378_ = new_n376_ & new_n377_;
  assign new_n379_ = ~new_n359_ & new_n378_;
  assign new_n380_ = p_457_142_ & ~new_n362_;
  assign new_n381_ = ~new_n353_ & new_n380_;
  assign new_n382_ = p_468_143_ & ~new_n356_;
  assign new_n383_ = ~new_n353_ & new_n382_;
  assign new_n384_ = ~new_n365_ & new_n383_;
  assign new_n385_ = p_446_141_ & ~new_n350_;
  assign new_n386_ = ~new_n379_ & ~new_n381_;
  assign new_n387_ = ~new_n384_ & new_n386_;
  assign new_n388_ = ~new_n385_ & new_n387_;
  assign p_591_1894_ = new_n375_ | ~new_n388_;
  assign new_n390_ = p_1690_158_ & p_1689_157_;
  assign new_n391_ = p_158_71_ & new_n390_;
  assign new_n392_ = ~p_374_134_ & ~new_n329_;
  assign new_n393_ = p_374_134_ & new_n329_;
  assign new_n394_ = ~new_n392_ & ~new_n393_;
  assign new_n395_ = p_4_1_ & ~new_n394_;
  assign new_n396_ = ~new_n330_ & ~new_n395_;
  assign new_n397_ = new_n333_ & ~new_n396_;
  assign new_n398_ = ~new_n333_ & new_n396_;
  assign new_n399_ = ~new_n397_ & ~new_n398_;
  assign new_n400_ = p_4091_175_ & ~p_4092_176_;
  assign new_n401_ = ~new_n399_ & new_n400_;
  assign new_n402_ = ~p_4091_175_ & p_4092_176_;
  assign new_n403_ = p_126_54_ & new_n402_;
  assign new_n404_ = ~p_273_106_ & ~p_3548_166_;
  assign new_n405_ = p_273_106_ & ~p_3546_165_;
  assign new_n406_ = ~p_411_138_ & ~new_n404_;
  assign new_n407_ = ~new_n405_ & new_n406_;
  assign new_n408_ = ~p_273_106_ & ~p_3550_167_;
  assign new_n409_ = p_411_138_ & new_n408_;
  assign new_n410_ = p_273_106_ & p_411_138_;
  assign new_n411_ = ~p_3552_168_ & new_n410_;
  assign new_n412_ = ~new_n409_ & ~new_n411_;
  assign new_n413_ = ~new_n407_ & new_n412_;
  assign new_n414_ = ~p_4091_175_ & ~p_4092_176_;
  assign new_n415_ = new_n413_ & new_n414_;
  assign new_n416_ = ~new_n401_ & ~new_n403_;
  assign p_877_2126_ = ~new_n415_ & new_n416_;
  assign new_n418_ = ~p_1690_158_ & p_1689_157_;
  assign new_n419_ = ~p_877_2126_ & new_n418_;
  assign new_n420_ = p_1690_158_ & ~p_1689_157_;
  assign new_n421_ = p_188_81_ & new_n420_;
  assign new_n422_ = p_358_128_ & p_332_122_;
  assign new_n423_ = p_351_127_ & ~p_332_122_;
  assign new_n424_ = ~new_n422_ & ~new_n423_;
  assign new_n425_ = ~p_534_149_ & ~new_n424_;
  assign new_n426_ = p_534_149_ & new_n424_;
  assign new_n427_ = ~new_n425_ & ~new_n426_;
  assign new_n428_ = p_332_122_ & p_366_130_;
  assign new_n429_ = p_361_129_ & ~p_332_122_;
  assign new_n430_ = ~new_n428_ & ~new_n429_;
  assign new_n431_ = p_54_20_ & new_n430_;
  assign new_n432_ = new_n430_ & ~new_n431_;
  assign new_n433_ = new_n427_ & ~new_n432_;
  assign new_n434_ = ~new_n427_ & new_n432_;
  assign new_n435_ = ~new_n433_ & ~new_n434_;
  assign new_n436_ = new_n400_ & ~new_n435_;
  assign new_n437_ = p_129_57_ & new_n402_;
  assign new_n438_ = ~p_351_127_ & ~p_3548_166_;
  assign new_n439_ = p_351_127_ & ~p_3546_165_;
  assign new_n440_ = ~p_534_149_ & ~new_n438_;
  assign new_n441_ = ~new_n439_ & new_n440_;
  assign new_n442_ = ~p_3550_167_ & ~p_351_127_;
  assign new_n443_ = p_534_149_ & new_n442_;
  assign new_n444_ = p_534_149_ & p_351_127_;
  assign new_n445_ = ~p_3552_168_ & new_n444_;
  assign new_n446_ = ~new_n443_ & ~new_n445_;
  assign new_n447_ = ~new_n441_ & new_n446_;
  assign new_n448_ = new_n414_ & new_n447_;
  assign new_n449_ = ~new_n436_ & ~new_n437_;
  assign p_838_2064_ = ~new_n448_ & new_n449_;
  assign new_n451_ = ~p_1690_158_ & ~p_1689_157_;
  assign new_n452_ = ~p_838_2064_ & new_n451_;
  assign new_n453_ = ~new_n391_ & ~new_n419_;
  assign new_n454_ = ~new_n421_ & new_n453_;
  assign new_n455_ = ~new_n452_ & new_n454_;
  assign p_664_2223_ = p_137_63_ & ~new_n455_;
  assign new_n457_ = p_1694_160_ & p_1691_159_;
  assign new_n458_ = p_179_78_ & new_n457_;
  assign new_n459_ = p_4092_176_ & p_97_37_;
  assign new_n460_ = ~new_n307_ & ~new_n323_;
  assign new_n461_ = new_n330_ & new_n460_;
  assign new_n462_ = ~new_n333_ & new_n461_;
  assign new_n463_ = ~new_n323_ & ~new_n333_;
  assign new_n464_ = ~new_n307_ & new_n463_;
  assign new_n465_ = ~new_n394_ & new_n464_;
  assign new_n466_ = ~new_n307_ & new_n340_;
  assign new_n467_ = ~new_n307_ & new_n317_;
  assign new_n468_ = ~new_n323_ & new_n467_;
  assign new_n469_ = ~new_n462_ & ~new_n465_;
  assign new_n470_ = ~new_n466_ & new_n469_;
  assign new_n471_ = ~new_n468_ & new_n470_;
  assign new_n472_ = ~new_n338_ & new_n471_;
  assign new_n473_ = ~new_n333_ & ~new_n394_;
  assign new_n474_ = new_n330_ & ~new_n333_;
  assign new_n475_ = ~new_n317_ & ~new_n474_;
  assign new_n476_ = ~new_n473_ & new_n475_;
  assign new_n477_ = ~new_n394_ & new_n463_;
  assign new_n478_ = new_n317_ & ~new_n323_;
  assign new_n479_ = ~new_n323_ & new_n330_;
  assign new_n480_ = ~new_n333_ & new_n479_;
  assign new_n481_ = ~new_n477_ & ~new_n478_;
  assign new_n482_ = ~new_n480_ & new_n481_;
  assign new_n483_ = ~new_n340_ & new_n482_;
  assign new_n484_ = ~p_374_134_ & new_n329_;
  assign new_n485_ = new_n483_ & new_n484_;
  assign new_n486_ = ~new_n483_ & ~new_n484_;
  assign new_n487_ = ~new_n485_ & ~new_n486_;
  assign new_n488_ = new_n476_ & ~new_n487_;
  assign new_n489_ = ~new_n476_ & new_n487_;
  assign new_n490_ = ~new_n488_ & ~new_n489_;
  assign new_n491_ = new_n472_ & ~new_n490_;
  assign new_n492_ = ~new_n472_ & new_n490_;
  assign new_n493_ = ~new_n491_ & ~new_n492_;
  assign new_n494_ = new_n394_ & ~new_n493_;
  assign new_n495_ = ~new_n394_ & new_n493_;
  assign new_n496_ = ~new_n494_ & ~new_n495_;
  assign new_n497_ = new_n333_ & ~new_n496_;
  assign new_n498_ = ~new_n333_ & new_n496_;
  assign new_n499_ = ~new_n497_ & ~new_n498_;
  assign new_n500_ = new_n313_ & ~new_n499_;
  assign new_n501_ = ~new_n313_ & new_n499_;
  assign new_n502_ = ~new_n500_ & ~new_n501_;
  assign new_n503_ = new_n323_ & ~new_n502_;
  assign new_n504_ = ~new_n323_ & new_n502_;
  assign new_n505_ = ~new_n503_ & ~new_n504_;
  assign new_n506_ = new_n307_ & ~new_n505_;
  assign new_n507_ = ~new_n307_ & new_n505_;
  assign new_n508_ = ~new_n506_ & ~new_n507_;
  assign new_n509_ = p_1497_156_ & ~new_n508_;
  assign new_n510_ = ~new_n462_ & ~new_n466_;
  assign new_n511_ = ~new_n468_ & new_n510_;
  assign new_n512_ = ~new_n338_ & new_n511_;
  assign new_n513_ = ~new_n478_ & ~new_n480_;
  assign new_n514_ = ~new_n340_ & new_n513_;
  assign new_n515_ = new_n330_ & ~new_n514_;
  assign new_n516_ = ~new_n330_ & new_n514_;
  assign new_n517_ = ~new_n515_ & ~new_n516_;
  assign new_n518_ = ~new_n475_ & ~new_n517_;
  assign new_n519_ = new_n475_ & new_n517_;
  assign new_n520_ = ~new_n518_ & ~new_n519_;
  assign new_n521_ = ~new_n512_ & ~new_n520_;
  assign new_n522_ = new_n512_ & new_n520_;
  assign new_n523_ = ~new_n521_ & ~new_n522_;
  assign new_n524_ = new_n394_ & ~new_n523_;
  assign new_n525_ = ~new_n394_ & new_n523_;
  assign new_n526_ = ~new_n524_ & ~new_n525_;
  assign new_n527_ = new_n333_ & ~new_n526_;
  assign new_n528_ = ~new_n333_ & new_n526_;
  assign new_n529_ = ~new_n527_ & ~new_n528_;
  assign new_n530_ = new_n313_ & ~new_n529_;
  assign new_n531_ = ~new_n313_ & new_n529_;
  assign new_n532_ = ~new_n530_ & ~new_n531_;
  assign new_n533_ = new_n323_ & ~new_n532_;
  assign new_n534_ = ~new_n323_ & new_n532_;
  assign new_n535_ = ~new_n533_ & ~new_n534_;
  assign new_n536_ = new_n307_ & ~new_n535_;
  assign new_n537_ = ~new_n307_ & new_n535_;
  assign new_n538_ = ~new_n536_ & ~new_n537_;
  assign new_n539_ = ~p_1497_156_ & new_n538_;
  assign new_n540_ = ~new_n509_ & ~new_n539_;
  assign new_n541_ = new_n324_ & ~new_n333_;
  assign new_n542_ = ~new_n323_ & new_n541_;
  assign new_n543_ = ~new_n394_ & new_n542_;
  assign new_n544_ = new_n347_ & ~new_n543_;
  assign new_n545_ = ~new_n359_ & ~new_n365_;
  assign new_n546_ = ~new_n371_ & new_n545_;
  assign new_n547_ = ~new_n365_ & new_n382_;
  assign new_n548_ = ~new_n365_ & new_n376_;
  assign new_n549_ = ~new_n359_ & new_n548_;
  assign new_n550_ = ~new_n546_ & ~new_n547_;
  assign new_n551_ = ~new_n549_ & new_n550_;
  assign new_n552_ = ~new_n380_ & new_n551_;
  assign new_n553_ = ~new_n359_ & ~new_n371_;
  assign new_n554_ = ~new_n359_ & new_n376_;
  assign new_n555_ = ~new_n382_ & ~new_n554_;
  assign new_n556_ = ~new_n553_ & new_n555_;
  assign new_n557_ = ~p_422_139_ & new_n368_;
  assign new_n558_ = new_n556_ & new_n557_;
  assign new_n559_ = ~new_n556_ & ~new_n557_;
  assign new_n560_ = ~new_n558_ & ~new_n559_;
  assign new_n561_ = new_n552_ & ~new_n560_;
  assign new_n562_ = ~new_n552_ & new_n560_;
  assign new_n563_ = ~new_n561_ & ~new_n562_;
  assign new_n564_ = new_n371_ & ~new_n563_;
  assign new_n565_ = ~new_n371_ & new_n563_;
  assign new_n566_ = ~new_n564_ & ~new_n565_;
  assign new_n567_ = new_n359_ & ~new_n566_;
  assign new_n568_ = ~new_n359_ & new_n566_;
  assign new_n569_ = ~new_n567_ & ~new_n568_;
  assign new_n570_ = new_n353_ & ~new_n569_;
  assign new_n571_ = ~new_n353_ & new_n569_;
  assign new_n572_ = ~new_n570_ & ~new_n571_;
  assign new_n573_ = new_n365_ & ~new_n572_;
  assign new_n574_ = ~new_n365_ & new_n572_;
  assign new_n575_ = ~new_n573_ & ~new_n574_;
  assign new_n576_ = p_1497_156_ & ~new_n544_;
  assign new_n577_ = ~new_n575_ & new_n576_;
  assign new_n578_ = ~p_1497_156_ & ~new_n347_;
  assign new_n579_ = ~new_n575_ & new_n578_;
  assign new_n580_ = ~new_n547_ & ~new_n549_;
  assign new_n581_ = ~new_n380_ & new_n580_;
  assign new_n582_ = new_n376_ & ~new_n555_;
  assign new_n583_ = ~new_n376_ & new_n555_;
  assign new_n584_ = ~new_n582_ & ~new_n583_;
  assign new_n585_ = ~new_n581_ & ~new_n584_;
  assign new_n586_ = new_n581_ & new_n584_;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = new_n371_ & ~new_n587_;
  assign new_n589_ = ~new_n371_ & new_n587_;
  assign new_n590_ = ~new_n588_ & ~new_n589_;
  assign new_n591_ = new_n359_ & ~new_n590_;
  assign new_n592_ = ~new_n359_ & new_n590_;
  assign new_n593_ = ~new_n591_ & ~new_n592_;
  assign new_n594_ = new_n353_ & ~new_n593_;
  assign new_n595_ = ~new_n353_ & new_n593_;
  assign new_n596_ = ~new_n594_ & ~new_n595_;
  assign new_n597_ = new_n365_ & ~new_n596_;
  assign new_n598_ = ~new_n365_ & new_n596_;
  assign new_n599_ = ~new_n597_ & ~new_n598_;
  assign new_n600_ = p_1497_156_ & new_n544_;
  assign new_n601_ = ~new_n599_ & new_n600_;
  assign new_n602_ = ~p_1497_156_ & new_n347_;
  assign new_n603_ = ~new_n599_ & new_n602_;
  assign new_n604_ = ~new_n577_ & ~new_n579_;
  assign new_n605_ = ~new_n601_ & new_n604_;
  assign new_n606_ = ~new_n603_ & new_n605_;
  assign new_n607_ = new_n540_ & ~new_n606_;
  assign new_n608_ = ~new_n540_ & new_n606_;
  assign new_n609_ = ~new_n607_ & ~new_n608_;
  assign new_n610_ = p_4091_175_ & new_n609_;
  assign new_n611_ = ~p_226_93_ & p_254_101_;
  assign new_n612_ = p_226_93_ & p_242_97_;
  assign new_n613_ = ~p_422_139_ & ~new_n611_;
  assign new_n614_ = ~new_n612_ & new_n613_;
  assign new_n615_ = ~p_226_93_ & p_251_100_;
  assign new_n616_ = p_422_139_ & new_n615_;
  assign new_n617_ = p_226_93_ & p_422_139_;
  assign new_n618_ = p_248_99_ & new_n617_;
  assign new_n619_ = ~new_n616_ & ~new_n618_;
  assign new_n620_ = ~new_n614_ & new_n619_;
  assign new_n621_ = p_254_101_ & ~p_218_91_;
  assign new_n622_ = p_242_97_ & p_218_91_;
  assign new_n623_ = ~p_468_143_ & ~new_n621_;
  assign new_n624_ = ~new_n622_ & new_n623_;
  assign new_n625_ = p_251_100_ & ~p_218_91_;
  assign new_n626_ = p_468_143_ & new_n625_;
  assign new_n627_ = p_468_143_ & p_218_91_;
  assign new_n628_ = p_248_99_ & new_n627_;
  assign new_n629_ = ~new_n626_ & ~new_n628_;
  assign new_n630_ = ~new_n624_ & new_n629_;
  assign new_n631_ = ~new_n620_ & new_n630_;
  assign new_n632_ = new_n620_ & ~new_n630_;
  assign new_n633_ = ~new_n631_ & ~new_n632_;
  assign new_n634_ = ~p_210_89_ & p_254_101_;
  assign new_n635_ = p_210_89_ & p_242_97_;
  assign new_n636_ = ~p_457_142_ & ~new_n634_;
  assign new_n637_ = ~new_n635_ & new_n636_;
  assign new_n638_ = ~p_210_89_ & p_251_100_;
  assign new_n639_ = p_457_142_ & new_n638_;
  assign new_n640_ = p_210_89_ & p_457_142_;
  assign new_n641_ = p_248_99_ & new_n640_;
  assign new_n642_ = ~new_n639_ & ~new_n641_;
  assign new_n643_ = ~new_n637_ & new_n642_;
  assign new_n644_ = ~p_206_87_ & p_254_101_;
  assign new_n645_ = p_206_87_ & p_242_97_;
  assign new_n646_ = ~p_446_141_ & ~new_n644_;
  assign new_n647_ = ~new_n645_ & new_n646_;
  assign new_n648_ = ~p_206_87_ & p_251_100_;
  assign new_n649_ = p_446_141_ & new_n648_;
  assign new_n650_ = p_206_87_ & p_446_141_;
  assign new_n651_ = p_248_99_ & new_n650_;
  assign new_n652_ = ~new_n649_ & ~new_n651_;
  assign new_n653_ = ~new_n647_ & new_n652_;
  assign new_n654_ = ~new_n643_ & new_n653_;
  assign new_n655_ = new_n643_ & ~new_n653_;
  assign new_n656_ = ~new_n654_ & ~new_n655_;
  assign new_n657_ = new_n633_ & ~new_n656_;
  assign new_n658_ = ~new_n633_ & new_n656_;
  assign new_n659_ = ~new_n657_ & ~new_n658_;
  assign new_n660_ = p_254_101_ & ~p_281_108_;
  assign new_n661_ = p_242_97_ & p_281_108_;
  assign new_n662_ = ~p_374_134_ & ~new_n660_;
  assign new_n663_ = ~new_n661_ & new_n662_;
  assign new_n664_ = p_251_100_ & ~p_281_108_;
  assign new_n665_ = p_374_134_ & new_n664_;
  assign new_n666_ = p_374_134_ & p_281_108_;
  assign new_n667_ = p_248_99_ & new_n666_;
  assign new_n668_ = ~new_n665_ & ~new_n667_;
  assign new_n669_ = ~new_n663_ & new_n668_;
  assign new_n670_ = ~p_257_102_ & p_254_101_;
  assign new_n671_ = p_257_102_ & p_242_97_;
  assign new_n672_ = ~p_389_136_ & ~new_n670_;
  assign new_n673_ = ~new_n671_ & new_n672_;
  assign new_n674_ = ~p_257_102_ & p_251_100_;
  assign new_n675_ = p_389_136_ & new_n674_;
  assign new_n676_ = p_257_102_ & p_389_136_;
  assign new_n677_ = p_248_99_ & new_n676_;
  assign new_n678_ = ~new_n675_ & ~new_n677_;
  assign new_n679_ = ~new_n673_ & new_n678_;
  assign new_n680_ = p_254_101_ & ~p_234_95_;
  assign new_n681_ = p_242_97_ & p_234_95_;
  assign new_n682_ = ~p_435_140_ & ~new_n680_;
  assign new_n683_ = ~new_n681_ & new_n682_;
  assign new_n684_ = p_251_100_ & ~p_234_95_;
  assign new_n685_ = p_435_140_ & new_n684_;
  assign new_n686_ = p_435_140_ & p_234_95_;
  assign new_n687_ = p_248_99_ & new_n686_;
  assign new_n688_ = ~new_n685_ & ~new_n687_;
  assign new_n689_ = ~new_n683_ & new_n688_;
  assign new_n690_ = ~new_n679_ & new_n689_;
  assign new_n691_ = new_n679_ & ~new_n689_;
  assign new_n692_ = ~new_n690_ & ~new_n691_;
  assign new_n693_ = p_254_101_ & ~p_273_106_;
  assign new_n694_ = p_242_97_ & p_273_106_;
  assign new_n695_ = ~p_411_138_ & ~new_n693_;
  assign new_n696_ = ~new_n694_ & new_n695_;
  assign new_n697_ = ~p_273_106_ & p_251_100_;
  assign new_n698_ = p_411_138_ & new_n697_;
  assign new_n699_ = p_248_99_ & new_n410_;
  assign new_n700_ = ~new_n698_ & ~new_n699_;
  assign new_n701_ = ~new_n696_ & new_n700_;
  assign new_n702_ = p_254_101_ & ~p_265_104_;
  assign new_n703_ = p_242_97_ & p_265_104_;
  assign new_n704_ = ~p_400_137_ & ~new_n702_;
  assign new_n705_ = ~new_n703_ & new_n704_;
  assign new_n706_ = p_251_100_ & ~p_265_104_;
  assign new_n707_ = p_400_137_ & new_n706_;
  assign new_n708_ = p_400_137_ & p_265_104_;
  assign new_n709_ = p_248_99_ & new_n708_;
  assign new_n710_ = ~new_n707_ & ~new_n709_;
  assign new_n711_ = ~new_n705_ & new_n710_;
  assign new_n712_ = ~new_n701_ & new_n711_;
  assign new_n713_ = new_n701_ & ~new_n711_;
  assign new_n714_ = ~new_n712_ & ~new_n713_;
  assign new_n715_ = ~new_n669_ & ~new_n692_;
  assign new_n716_ = ~new_n714_ & new_n715_;
  assign new_n717_ = new_n692_ & ~new_n714_;
  assign new_n718_ = new_n669_ & new_n717_;
  assign new_n719_ = ~new_n716_ & ~new_n718_;
  assign new_n720_ = new_n669_ & ~new_n692_;
  assign new_n721_ = new_n714_ & new_n720_;
  assign new_n722_ = new_n692_ & new_n714_;
  assign new_n723_ = ~new_n669_ & new_n722_;
  assign new_n724_ = ~new_n721_ & ~new_n723_;
  assign new_n725_ = new_n719_ & new_n724_;
  assign new_n726_ = new_n659_ & ~new_n725_;
  assign new_n727_ = ~new_n659_ & new_n725_;
  assign new_n728_ = ~new_n726_ & ~new_n727_;
  assign new_n729_ = ~p_4091_175_ & ~new_n728_;
  assign new_n730_ = ~new_n610_ & ~new_n729_;
  assign new_n731_ = ~p_4092_176_ & ~new_n730_;
  assign new_n732_ = ~new_n459_ & ~new_n731_;
  assign new_n733_ = ~p_1694_160_ & p_1691_159_;
  assign new_n734_ = ~new_n732_ & new_n733_;
  assign new_n735_ = p_1694_160_ & ~p_1691_159_;
  assign new_n736_ = p_176_77_ & new_n735_;
  assign new_n737_ = p_94_36_ & p_4092_176_;
  assign new_n738_ = p_338_124_ & p_332_122_;
  assign new_n739_ = p_332_122_ & ~new_n738_;
  assign new_n740_ = p_514_147_ & new_n739_;
  assign new_n741_ = ~p_514_147_ & ~new_n739_;
  assign new_n742_ = ~new_n740_ & ~new_n741_;
  assign new_n743_ = p_348_126_ & p_332_122_;
  assign new_n744_ = p_341_125_ & ~p_332_122_;
  assign new_n745_ = ~new_n743_ & ~new_n744_;
  assign new_n746_ = p_523_148_ & new_n745_;
  assign new_n747_ = ~p_523_148_ & ~new_n745_;
  assign new_n748_ = ~new_n746_ & ~new_n747_;
  assign new_n749_ = p_331_121_ & p_332_122_;
  assign new_n750_ = p_324_120_ & ~p_332_122_;
  assign new_n751_ = ~new_n749_ & ~new_n750_;
  assign new_n752_ = p_503_146_ & new_n751_;
  assign new_n753_ = ~p_503_146_ & ~new_n751_;
  assign new_n754_ = ~new_n752_ & ~new_n753_;
  assign new_n755_ = ~new_n742_ & ~new_n748_;
  assign new_n756_ = ~new_n430_ & new_n755_;
  assign new_n757_ = ~new_n427_ & new_n756_;
  assign new_n758_ = ~new_n427_ & ~new_n748_;
  assign new_n759_ = ~new_n742_ & new_n758_;
  assign new_n760_ = new_n430_ & new_n759_;
  assign new_n761_ = p_523_148_ & ~new_n745_;
  assign new_n762_ = ~new_n742_ & new_n761_;
  assign new_n763_ = p_534_149_ & ~new_n424_;
  assign new_n764_ = ~new_n742_ & new_n763_;
  assign new_n765_ = ~new_n748_ & new_n764_;
  assign new_n766_ = p_514_147_ & ~new_n739_;
  assign new_n767_ = ~new_n757_ & ~new_n760_;
  assign new_n768_ = ~new_n762_ & new_n767_;
  assign new_n769_ = ~new_n765_ & new_n768_;
  assign new_n770_ = ~new_n766_ & new_n769_;
  assign new_n771_ = ~new_n427_ & new_n430_;
  assign new_n772_ = ~new_n427_ & ~new_n430_;
  assign new_n773_ = ~new_n763_ & ~new_n772_;
  assign new_n774_ = ~new_n771_ & new_n773_;
  assign new_n775_ = new_n430_ & new_n758_;
  assign new_n776_ = ~new_n748_ & new_n763_;
  assign new_n777_ = ~new_n430_ & ~new_n748_;
  assign new_n778_ = ~new_n427_ & new_n777_;
  assign new_n779_ = ~new_n775_ & ~new_n776_;
  assign new_n780_ = ~new_n778_ & new_n779_;
  assign new_n781_ = ~new_n761_ & new_n780_;
  assign new_n782_ = new_n774_ & ~new_n781_;
  assign new_n783_ = ~new_n774_ & new_n781_;
  assign new_n784_ = ~new_n782_ & ~new_n783_;
  assign new_n785_ = new_n770_ & ~new_n784_;
  assign new_n786_ = ~new_n770_ & new_n784_;
  assign new_n787_ = ~new_n785_ & ~new_n786_;
  assign new_n788_ = ~new_n430_ & ~new_n787_;
  assign new_n789_ = new_n430_ & new_n787_;
  assign new_n790_ = ~new_n788_ & ~new_n789_;
  assign new_n791_ = new_n427_ & ~new_n790_;
  assign new_n792_ = ~new_n427_ & new_n790_;
  assign new_n793_ = ~new_n791_ & ~new_n792_;
  assign new_n794_ = new_n754_ & ~new_n793_;
  assign new_n795_ = ~new_n754_ & new_n793_;
  assign new_n796_ = ~new_n794_ & ~new_n795_;
  assign new_n797_ = new_n748_ & ~new_n796_;
  assign new_n798_ = ~new_n748_ & new_n796_;
  assign new_n799_ = ~new_n797_ & ~new_n798_;
  assign new_n800_ = new_n742_ & ~new_n799_;
  assign new_n801_ = ~new_n742_ & new_n799_;
  assign new_n802_ = ~new_n800_ & ~new_n801_;
  assign new_n803_ = p_2174_161_ & ~new_n802_;
  assign new_n804_ = ~new_n757_ & ~new_n762_;
  assign new_n805_ = ~new_n765_ & new_n804_;
  assign new_n806_ = ~new_n766_ & new_n805_;
  assign new_n807_ = ~new_n776_ & ~new_n778_;
  assign new_n808_ = ~new_n761_ & new_n807_;
  assign new_n809_ = ~new_n430_ & ~new_n808_;
  assign new_n810_ = new_n430_ & new_n808_;
  assign new_n811_ = ~new_n809_ & ~new_n810_;
  assign new_n812_ = ~new_n773_ & ~new_n811_;
  assign new_n813_ = new_n773_ & new_n811_;
  assign new_n814_ = ~new_n812_ & ~new_n813_;
  assign new_n815_ = ~new_n806_ & ~new_n814_;
  assign new_n816_ = new_n806_ & new_n814_;
  assign new_n817_ = ~new_n815_ & ~new_n816_;
  assign new_n818_ = ~new_n430_ & ~new_n817_;
  assign new_n819_ = new_n430_ & new_n817_;
  assign new_n820_ = ~new_n818_ & ~new_n819_;
  assign new_n821_ = new_n427_ & ~new_n820_;
  assign new_n822_ = ~new_n427_ & new_n820_;
  assign new_n823_ = ~new_n821_ & ~new_n822_;
  assign new_n824_ = new_n754_ & ~new_n823_;
  assign new_n825_ = ~new_n754_ & new_n823_;
  assign new_n826_ = ~new_n824_ & ~new_n825_;
  assign new_n827_ = new_n748_ & ~new_n826_;
  assign new_n828_ = ~new_n748_ & new_n826_;
  assign new_n829_ = ~new_n827_ & ~new_n828_;
  assign new_n830_ = new_n742_ & ~new_n829_;
  assign new_n831_ = ~new_n742_ & new_n829_;
  assign new_n832_ = ~new_n830_ & ~new_n831_;
  assign new_n833_ = ~p_2174_161_ & new_n832_;
  assign new_n834_ = ~new_n803_ & ~new_n833_;
  assign new_n835_ = ~new_n742_ & ~new_n754_;
  assign new_n836_ = ~new_n427_ & new_n835_;
  assign new_n837_ = ~new_n748_ & new_n836_;
  assign new_n838_ = new_n430_ & new_n837_;
  assign new_n839_ = new_n763_ & new_n835_;
  assign new_n840_ = ~new_n748_ & new_n839_;
  assign new_n841_ = ~new_n430_ & ~new_n742_;
  assign new_n842_ = ~new_n748_ & new_n841_;
  assign new_n843_ = ~new_n754_ & new_n842_;
  assign new_n844_ = ~new_n427_ & new_n843_;
  assign new_n845_ = ~new_n754_ & new_n766_;
  assign new_n846_ = ~new_n754_ & new_n761_;
  assign new_n847_ = ~new_n742_ & new_n846_;
  assign new_n848_ = p_503_146_ & ~new_n751_;
  assign new_n849_ = ~new_n840_ & ~new_n844_;
  assign new_n850_ = ~new_n845_ & new_n849_;
  assign new_n851_ = ~new_n847_ & new_n850_;
  assign new_n852_ = ~new_n848_ & new_n851_;
  assign new_n853_ = ~new_n838_ & new_n852_;
  assign new_n854_ = p_307_115_ & p_332_122_;
  assign new_n855_ = p_302_114_ & ~p_332_122_;
  assign new_n856_ = ~new_n854_ & ~new_n855_;
  assign new_n857_ = p_299_113_ & p_332_122_;
  assign new_n858_ = p_293_112_ & ~p_332_122_;
  assign new_n859_ = ~new_n857_ & ~new_n858_;
  assign new_n860_ = p_315_117_ & p_332_122_;
  assign new_n861_ = p_308_116_ & ~p_332_122_;
  assign new_n862_ = ~new_n860_ & ~new_n861_;
  assign new_n863_ = p_479_144_ & new_n862_;
  assign new_n864_ = ~p_479_144_ & ~new_n862_;
  assign new_n865_ = ~new_n863_ & ~new_n864_;
  assign new_n866_ = p_323_119_ & p_332_122_;
  assign new_n867_ = ~p_332_122_ & p_316_118_;
  assign new_n868_ = ~new_n866_ & ~new_n867_;
  assign new_n869_ = p_490_145_ & new_n868_;
  assign new_n870_ = ~p_490_145_ & ~new_n868_;
  assign new_n871_ = ~new_n869_ & ~new_n870_;
  assign new_n872_ = new_n856_ & ~new_n865_;
  assign new_n873_ = ~new_n871_ & new_n872_;
  assign new_n874_ = p_479_144_ & ~new_n862_;
  assign new_n875_ = new_n856_ & new_n874_;
  assign new_n876_ = p_490_145_ & ~new_n868_;
  assign new_n877_ = new_n856_ & new_n876_;
  assign new_n878_ = ~new_n865_ & new_n877_;
  assign new_n879_ = ~new_n873_ & ~new_n875_;
  assign new_n880_ = ~new_n878_ & new_n879_;
  assign new_n881_ = new_n856_ & new_n880_;
  assign new_n882_ = ~new_n865_ & ~new_n871_;
  assign new_n883_ = ~new_n865_ & new_n876_;
  assign new_n884_ = ~new_n874_ & ~new_n883_;
  assign new_n885_ = ~new_n882_ & new_n884_;
  assign new_n886_ = ~p_490_145_ & new_n868_;
  assign new_n887_ = new_n885_ & new_n886_;
  assign new_n888_ = ~new_n885_ & ~new_n886_;
  assign new_n889_ = ~new_n887_ & ~new_n888_;
  assign new_n890_ = new_n881_ & ~new_n889_;
  assign new_n891_ = ~new_n881_ & new_n889_;
  assign new_n892_ = ~new_n890_ & ~new_n891_;
  assign new_n893_ = new_n871_ & ~new_n892_;
  assign new_n894_ = ~new_n871_ & new_n892_;
  assign new_n895_ = ~new_n893_ & ~new_n894_;
  assign new_n896_ = new_n865_ & ~new_n895_;
  assign new_n897_ = ~new_n865_ & new_n895_;
  assign new_n898_ = ~new_n896_ & ~new_n897_;
  assign new_n899_ = ~new_n859_ & ~new_n898_;
  assign new_n900_ = new_n859_ & new_n898_;
  assign new_n901_ = ~new_n899_ & ~new_n900_;
  assign new_n902_ = ~new_n856_ & ~new_n901_;
  assign new_n903_ = new_n856_ & new_n901_;
  assign new_n904_ = ~new_n902_ & ~new_n903_;
  assign new_n905_ = p_2174_161_ & ~new_n853_;
  assign new_n906_ = ~new_n904_ & new_n905_;
  assign new_n907_ = ~p_2174_161_ & ~new_n852_;
  assign new_n908_ = ~new_n904_ & new_n907_;
  assign new_n909_ = ~new_n875_ & ~new_n878_;
  assign new_n910_ = new_n856_ & new_n909_;
  assign new_n911_ = new_n876_ & ~new_n884_;
  assign new_n912_ = ~new_n876_ & new_n884_;
  assign new_n913_ = ~new_n911_ & ~new_n912_;
  assign new_n914_ = ~new_n910_ & ~new_n913_;
  assign new_n915_ = new_n910_ & new_n913_;
  assign new_n916_ = ~new_n914_ & ~new_n915_;
  assign new_n917_ = new_n871_ & ~new_n916_;
  assign new_n918_ = ~new_n871_ & new_n916_;
  assign new_n919_ = ~new_n917_ & ~new_n918_;
  assign new_n920_ = new_n865_ & ~new_n919_;
  assign new_n921_ = ~new_n865_ & new_n919_;
  assign new_n922_ = ~new_n920_ & ~new_n921_;
  assign new_n923_ = ~new_n859_ & ~new_n922_;
  assign new_n924_ = new_n859_ & new_n922_;
  assign new_n925_ = ~new_n923_ & ~new_n924_;
  assign new_n926_ = ~new_n856_ & ~new_n925_;
  assign new_n927_ = new_n856_ & new_n925_;
  assign new_n928_ = ~new_n926_ & ~new_n927_;
  assign new_n929_ = p_2174_161_ & new_n853_;
  assign new_n930_ = ~new_n928_ & new_n929_;
  assign new_n931_ = ~p_2174_161_ & new_n852_;
  assign new_n932_ = ~new_n928_ & new_n931_;
  assign new_n933_ = ~new_n906_ & ~new_n908_;
  assign new_n934_ = ~new_n930_ & new_n933_;
  assign new_n935_ = ~new_n932_ & new_n934_;
  assign new_n936_ = new_n834_ & ~new_n935_;
  assign new_n937_ = ~new_n834_ & new_n935_;
  assign new_n938_ = ~new_n936_ & ~new_n937_;
  assign new_n939_ = p_4091_175_ & new_n938_;
  assign new_n940_ = p_254_101_ & ~p_316_118_;
  assign new_n941_ = p_242_97_ & p_316_118_;
  assign new_n942_ = ~p_490_145_ & ~new_n940_;
  assign new_n943_ = ~new_n941_ & new_n942_;
  assign new_n944_ = p_251_100_ & ~p_316_118_;
  assign new_n945_ = p_490_145_ & new_n944_;
  assign new_n946_ = p_490_145_ & p_316_118_;
  assign new_n947_ = p_248_99_ & new_n946_;
  assign new_n948_ = ~new_n945_ & ~new_n947_;
  assign new_n949_ = ~new_n943_ & new_n948_;
  assign new_n950_ = p_254_101_ & ~p_308_116_;
  assign new_n951_ = p_242_97_ & p_308_116_;
  assign new_n952_ = ~p_479_144_ & ~new_n950_;
  assign new_n953_ = ~new_n951_ & new_n952_;
  assign new_n954_ = ~p_308_116_ & p_251_100_;
  assign new_n955_ = p_479_144_ & new_n954_;
  assign new_n956_ = p_308_116_ & p_479_144_;
  assign new_n957_ = p_248_99_ & new_n956_;
  assign new_n958_ = ~new_n955_ & ~new_n957_;
  assign new_n959_ = ~new_n953_ & new_n958_;
  assign new_n960_ = ~new_n949_ & new_n959_;
  assign new_n961_ = new_n949_ & ~new_n959_;
  assign new_n962_ = ~new_n960_ & ~new_n961_;
  assign new_n963_ = ~p_302_114_ & p_251_100_;
  assign new_n964_ = p_302_114_ & p_248_99_;
  assign new_n965_ = ~new_n963_ & ~new_n964_;
  assign new_n966_ = ~p_293_112_ & p_254_101_;
  assign new_n967_ = p_293_112_ & p_242_97_;
  assign new_n968_ = ~new_n966_ & ~new_n967_;
  assign new_n969_ = ~new_n965_ & ~new_n968_;
  assign new_n970_ = new_n965_ & new_n968_;
  assign new_n971_ = ~new_n969_ & ~new_n970_;
  assign new_n972_ = new_n962_ & ~new_n971_;
  assign new_n973_ = ~new_n962_ & new_n971_;
  assign new_n974_ = ~new_n972_ & ~new_n973_;
  assign new_n975_ = p_251_100_ & ~p_361_129_;
  assign new_n976_ = p_248_99_ & p_361_129_;
  assign new_n977_ = ~new_n975_ & ~new_n976_;
  assign new_n978_ = ~p_514_147_ & ~p_242_97_;
  assign new_n979_ = p_514_147_ & p_248_99_;
  assign new_n980_ = ~new_n978_ & ~new_n979_;
  assign new_n981_ = ~p_324_120_ & p_254_101_;
  assign new_n982_ = p_324_120_ & p_242_97_;
  assign new_n983_ = ~p_503_146_ & ~new_n981_;
  assign new_n984_ = ~new_n982_ & new_n983_;
  assign new_n985_ = ~p_324_120_ & p_251_100_;
  assign new_n986_ = p_503_146_ & new_n985_;
  assign new_n987_ = p_324_120_ & p_503_146_;
  assign new_n988_ = p_248_99_ & new_n987_;
  assign new_n989_ = ~new_n986_ & ~new_n988_;
  assign new_n990_ = ~new_n984_ & new_n989_;
  assign new_n991_ = ~new_n980_ & new_n990_;
  assign new_n992_ = new_n980_ & ~new_n990_;
  assign new_n993_ = ~new_n991_ & ~new_n992_;
  assign new_n994_ = p_254_101_ & ~p_351_127_;
  assign new_n995_ = p_242_97_ & p_351_127_;
  assign new_n996_ = ~p_534_149_ & ~new_n994_;
  assign new_n997_ = ~new_n995_ & new_n996_;
  assign new_n998_ = p_251_100_ & ~p_351_127_;
  assign new_n999_ = p_534_149_ & new_n998_;
  assign new_n1000_ = p_248_99_ & new_n444_;
  assign new_n1001_ = ~new_n999_ & ~new_n1000_;
  assign new_n1002_ = ~new_n997_ & new_n1001_;
  assign new_n1003_ = p_254_101_ & ~p_341_125_;
  assign new_n1004_ = p_242_97_ & p_341_125_;
  assign new_n1005_ = ~p_523_148_ & ~new_n1003_;
  assign new_n1006_ = ~new_n1004_ & new_n1005_;
  assign new_n1007_ = p_251_100_ & ~p_341_125_;
  assign new_n1008_ = p_523_148_ & new_n1007_;
  assign new_n1009_ = p_341_125_ & p_523_148_;
  assign new_n1010_ = p_248_99_ & new_n1009_;
  assign new_n1011_ = ~new_n1008_ & ~new_n1010_;
  assign new_n1012_ = ~new_n1006_ & new_n1011_;
  assign new_n1013_ = ~new_n1002_ & new_n1012_;
  assign new_n1014_ = new_n1002_ & ~new_n1012_;
  assign new_n1015_ = ~new_n1013_ & ~new_n1014_;
  assign new_n1016_ = ~new_n977_ & ~new_n993_;
  assign new_n1017_ = ~new_n1015_ & new_n1016_;
  assign new_n1018_ = new_n993_ & ~new_n1015_;
  assign new_n1019_ = new_n977_ & new_n1018_;
  assign new_n1020_ = ~new_n1017_ & ~new_n1019_;
  assign new_n1021_ = new_n977_ & ~new_n993_;
  assign new_n1022_ = new_n1015_ & new_n1021_;
  assign new_n1023_ = new_n993_ & new_n1015_;
  assign new_n1024_ = ~new_n977_ & new_n1023_;
  assign new_n1025_ = ~new_n1022_ & ~new_n1024_;
  assign new_n1026_ = new_n1020_ & new_n1025_;
  assign new_n1027_ = new_n974_ & ~new_n1026_;
  assign new_n1028_ = ~new_n974_ & new_n1026_;
  assign new_n1029_ = ~new_n1027_ & ~new_n1028_;
  assign new_n1030_ = ~p_4091_175_ & ~new_n1029_;
  assign new_n1031_ = ~new_n939_ & ~new_n1030_;
  assign new_n1032_ = ~p_4092_176_ & ~new_n1031_;
  assign new_n1033_ = ~new_n737_ & ~new_n1032_;
  assign new_n1034_ = ~p_1694_160_ & ~p_1691_159_;
  assign new_n1035_ = ~new_n1033_ & new_n1034_;
  assign new_n1036_ = ~new_n458_ & ~new_n734_;
  assign new_n1037_ = ~new_n736_ & new_n1036_;
  assign new_n1038_ = ~new_n1035_ & new_n1037_;
  assign p_690_2484_ = ~p_137_63_ | new_n1038_;
  assign new_n1040_ = p_152_69_ & new_n457_;
  assign new_n1041_ = p_4_1_ & new_n473_;
  assign new_n1042_ = ~new_n474_ & ~new_n1041_;
  assign new_n1043_ = ~new_n317_ & new_n1042_;
  assign new_n1044_ = new_n323_ & ~new_n1043_;
  assign new_n1045_ = ~new_n323_ & new_n1043_;
  assign new_n1046_ = ~new_n1044_ & ~new_n1045_;
  assign new_n1047_ = new_n400_ & ~new_n1046_;
  assign new_n1048_ = p_127_55_ & new_n402_;
  assign new_n1049_ = ~p_3548_166_ & ~p_265_104_;
  assign new_n1050_ = ~p_3546_165_ & p_265_104_;
  assign new_n1051_ = ~p_400_137_ & ~new_n1049_;
  assign new_n1052_ = ~new_n1050_ & new_n1051_;
  assign new_n1053_ = ~p_3550_167_ & ~p_265_104_;
  assign new_n1054_ = p_400_137_ & new_n1053_;
  assign new_n1055_ = ~p_3552_168_ & new_n708_;
  assign new_n1056_ = ~new_n1054_ & ~new_n1055_;
  assign new_n1057_ = ~new_n1052_ & new_n1056_;
  assign new_n1058_ = new_n414_ & new_n1057_;
  assign new_n1059_ = ~new_n1047_ & ~new_n1048_;
  assign p_875_2125_ = ~new_n1058_ & new_n1059_;
  assign new_n1061_ = new_n733_ & ~p_875_2125_;
  assign new_n1062_ = p_155_70_ & new_n735_;
  assign new_n1063_ = p_54_20_ & new_n771_;
  assign new_n1064_ = ~new_n772_ & ~new_n1063_;
  assign new_n1065_ = ~new_n763_ & new_n1064_;
  assign new_n1066_ = new_n748_ & ~new_n1065_;
  assign new_n1067_ = ~new_n748_ & new_n1065_;
  assign new_n1068_ = ~new_n1066_ & ~new_n1067_;
  assign new_n1069_ = new_n400_ & ~new_n1068_;
  assign new_n1070_ = p_119_49_ & new_n402_;
  assign new_n1071_ = ~p_341_125_ & ~p_3548_166_;
  assign new_n1072_ = p_341_125_ & ~p_3546_165_;
  assign new_n1073_ = ~p_523_148_ & ~new_n1071_;
  assign new_n1074_ = ~new_n1072_ & new_n1073_;
  assign new_n1075_ = ~p_3550_167_ & ~p_341_125_;
  assign new_n1076_ = p_523_148_ & new_n1075_;
  assign new_n1077_ = ~p_3552_168_ & new_n1009_;
  assign new_n1078_ = ~new_n1076_ & ~new_n1077_;
  assign new_n1079_ = ~new_n1074_ & new_n1078_;
  assign new_n1080_ = new_n414_ & new_n1079_;
  assign new_n1081_ = ~new_n1069_ & ~new_n1070_;
  assign p_836_2128_ = ~new_n1080_ & new_n1081_;
  assign new_n1083_ = new_n1034_ & ~p_836_2128_;
  assign new_n1084_ = ~new_n1040_ & ~new_n1061_;
  assign new_n1085_ = ~new_n1062_ & new_n1084_;
  assign new_n1086_ = ~new_n1083_ & new_n1085_;
  assign p_699_2227_ = p_137_63_ & ~new_n1086_;
  assign new_n1088_ = new_n859_ & ~new_n871_;
  assign new_n1089_ = ~new_n865_ & new_n1088_;
  assign new_n1090_ = new_n856_ & new_n1089_;
  assign new_n1091_ = ~new_n852_ & new_n1090_;
  assign new_n1092_ = new_n856_ & new_n859_;
  assign new_n1093_ = new_n876_ & new_n1092_;
  assign new_n1094_ = ~new_n865_ & new_n1093_;
  assign new_n1095_ = ~new_n856_ & new_n859_;
  assign new_n1096_ = new_n859_ & new_n874_;
  assign new_n1097_ = new_n856_ & new_n1096_;
  assign new_n1098_ = ~new_n1094_ & ~new_n1095_;
  assign new_n1099_ = ~new_n1097_ & new_n1098_;
  assign new_n1100_ = new_n859_ & new_n1099_;
  assign p_618_1925_ = new_n1091_ | ~new_n1100_;
  assign p_588_1696_ = new_n374_ & new_n543_;
  assign new_n1103_ = ~new_n427_ & ~new_n754_;
  assign new_n1104_ = new_n430_ & new_n1103_;
  assign new_n1105_ = ~new_n748_ & new_n1104_;
  assign new_n1106_ = ~new_n742_ & new_n1105_;
  assign p_615_1750_ = new_n1090_ & new_n1106_;
  assign new_n1108_ = p_161_72_ & new_n457_;
  assign new_n1109_ = new_n353_ & ~new_n552_;
  assign new_n1110_ = ~new_n353_ & new_n552_;
  assign new_n1111_ = ~new_n1109_ & ~new_n1110_;
  assign new_n1112_ = ~new_n313_ & ~new_n333_;
  assign new_n1113_ = ~new_n394_ & new_n1112_;
  assign new_n1114_ = ~new_n323_ & new_n1113_;
  assign new_n1115_ = ~new_n307_ & new_n1114_;
  assign new_n1116_ = p_4_1_ & new_n1115_;
  assign new_n1117_ = new_n347_ & ~new_n1116_;
  assign new_n1118_ = ~new_n1111_ & ~new_n1117_;
  assign new_n1119_ = new_n376_ & new_n545_;
  assign new_n1120_ = ~new_n547_ & ~new_n1119_;
  assign new_n1121_ = ~new_n380_ & new_n1120_;
  assign new_n1122_ = new_n353_ & new_n1121_;
  assign new_n1123_ = ~new_n353_ & ~new_n1121_;
  assign new_n1124_ = ~new_n1122_ & ~new_n1123_;
  assign new_n1125_ = new_n1117_ & new_n1124_;
  assign new_n1126_ = ~new_n1118_ & ~new_n1125_;
  assign new_n1127_ = new_n400_ & ~new_n1126_;
  assign new_n1128_ = p_115_45_ & new_n402_;
  assign new_n1129_ = new_n414_ & new_n653_;
  assign new_n1130_ = ~new_n1127_ & ~new_n1128_;
  assign p_863_2276_ = ~new_n1129_ & new_n1130_;
  assign new_n1132_ = new_n733_ & ~p_863_2276_;
  assign new_n1133_ = p_191_82_ & new_n735_;
  assign new_n1134_ = ~new_n859_ & ~new_n881_;
  assign new_n1135_ = new_n859_ & new_n881_;
  assign new_n1136_ = ~new_n1134_ & ~new_n1135_;
  assign new_n1137_ = p_54_20_ & new_n1106_;
  assign new_n1138_ = new_n852_ & ~new_n1137_;
  assign new_n1139_ = ~new_n1136_ & ~new_n1138_;
  assign new_n1140_ = new_n872_ & new_n876_;
  assign new_n1141_ = ~new_n875_ & ~new_n1140_;
  assign new_n1142_ = new_n856_ & new_n1141_;
  assign new_n1143_ = ~new_n859_ & new_n1142_;
  assign new_n1144_ = new_n859_ & ~new_n1142_;
  assign new_n1145_ = ~new_n1143_ & ~new_n1144_;
  assign new_n1146_ = new_n1138_ & new_n1145_;
  assign p_623_2152_ = ~new_n1139_ & ~new_n1146_;
  assign new_n1148_ = new_n400_ & ~p_623_2152_;
  assign new_n1149_ = p_123_53_ & new_n402_;
  assign new_n1150_ = new_n414_ & ~new_n968_;
  assign new_n1151_ = ~new_n1148_ & ~new_n1149_;
  assign p_824_2274_ = ~new_n1150_ & new_n1151_;
  assign new_n1153_ = new_n1034_ & ~p_824_2274_;
  assign new_n1154_ = ~new_n1108_ & ~new_n1132_;
  assign new_n1155_ = ~new_n1133_ & new_n1154_;
  assign new_n1156_ = ~new_n1153_ & new_n1155_;
  assign p_688_2317_ = p_137_63_ & ~new_n1156_;
  assign p_809_655_ = ~p_31_11_ | ~p_27_10_;
  assign new_n1159_ = p_88_34_ & ~p_2358_162_;
  assign new_n1160_ = p_34_12_ & p_2358_162_;
  assign new_n1161_ = ~new_n1159_ & ~new_n1160_;
  assign p_704_1281_ = p_809_655_ | new_n1161_;
  assign new_n1163_ = p_3717_169_ & p_3724_170_;
  assign new_n1164_ = ~p_623_2152_ & new_n1163_;
  assign new_n1165_ = p_132_60_ & new_n859_;
  assign new_n1166_ = p_132_60_ & ~new_n1165_;
  assign new_n1167_ = new_n859_ & ~new_n1165_;
  assign new_n1168_ = ~new_n1166_ & ~new_n1167_;
  assign new_n1169_ = ~p_3717_169_ & p_3724_170_;
  assign new_n1170_ = ~new_n1168_ & new_n1169_;
  assign new_n1171_ = p_3717_169_ & ~p_3724_170_;
  assign new_n1172_ = p_123_53_ & new_n1171_;
  assign new_n1173_ = ~p_3717_169_ & ~p_3724_170_;
  assign new_n1174_ = ~new_n968_ & new_n1173_;
  assign new_n1175_ = ~new_n1164_ & ~new_n1170_;
  assign new_n1176_ = ~new_n1172_ & new_n1175_;
  assign new_n1177_ = ~new_n1174_ & new_n1176_;
  assign new_n1178_ = p_4115_177_ & p_135_61_;
  assign p_818_2273_ = ~new_n1177_ & ~new_n1178_;
  assign new_n1180_ = new_n371_ & ~new_n1117_;
  assign new_n1181_ = ~new_n371_ & new_n1117_;
  assign new_n1182_ = ~new_n1180_ & ~new_n1181_;
  assign new_n1183_ = new_n400_ & ~new_n1182_;
  assign new_n1184_ = p_113_43_ & new_n402_;
  assign new_n1185_ = ~p_226_93_ & ~p_3548_166_;
  assign new_n1186_ = p_226_93_ & ~p_3546_165_;
  assign new_n1187_ = ~p_422_139_ & ~new_n1185_;
  assign new_n1188_ = ~new_n1186_ & new_n1187_;
  assign new_n1189_ = ~p_226_93_ & ~p_3550_167_;
  assign new_n1190_ = p_422_139_ & new_n1189_;
  assign new_n1191_ = ~p_3552_168_ & new_n617_;
  assign new_n1192_ = ~new_n1190_ & ~new_n1191_;
  assign new_n1193_ = ~new_n1188_ & new_n1192_;
  assign new_n1194_ = new_n414_ & new_n1193_;
  assign new_n1195_ = ~new_n1183_ & ~new_n1184_;
  assign p_869_2181_ = ~new_n1194_ & new_n1195_;
  assign new_n1197_ = p_167_74_ & new_n390_;
  assign new_n1198_ = new_n359_ & new_n557_;
  assign new_n1199_ = ~new_n359_ & ~new_n557_;
  assign new_n1200_ = ~new_n1198_ & ~new_n1199_;
  assign new_n1201_ = ~new_n1117_ & new_n1200_;
  assign new_n1202_ = new_n359_ & new_n376_;
  assign new_n1203_ = ~new_n359_ & ~new_n376_;
  assign new_n1204_ = ~new_n1202_ & ~new_n1203_;
  assign new_n1205_ = new_n1117_ & ~new_n1204_;
  assign new_n1206_ = ~new_n1201_ & ~new_n1205_;
  assign new_n1207_ = new_n400_ & ~new_n1206_;
  assign new_n1208_ = p_53_19_ & new_n402_;
  assign new_n1209_ = ~p_3548_166_ & ~p_218_91_;
  assign new_n1210_ = ~p_3546_165_ & p_218_91_;
  assign new_n1211_ = ~p_468_143_ & ~new_n1209_;
  assign new_n1212_ = ~new_n1210_ & new_n1211_;
  assign new_n1213_ = ~p_3550_167_ & ~p_218_91_;
  assign new_n1214_ = p_468_143_ & new_n1213_;
  assign new_n1215_ = ~p_3552_168_ & new_n627_;
  assign new_n1216_ = ~new_n1214_ & ~new_n1215_;
  assign new_n1217_ = ~new_n1212_ & new_n1216_;
  assign new_n1218_ = new_n414_ & new_n1217_;
  assign new_n1219_ = ~new_n1207_ & ~new_n1208_;
  assign p_867_2237_ = ~new_n1218_ & new_n1219_;
  assign new_n1221_ = new_n418_ & ~p_867_2237_;
  assign new_n1222_ = p_197_84_ & new_n420_;
  assign new_n1223_ = new_n865_ & new_n886_;
  assign new_n1224_ = ~new_n865_ & ~new_n886_;
  assign new_n1225_ = ~new_n1223_ & ~new_n1224_;
  assign new_n1226_ = ~new_n1138_ & new_n1225_;
  assign new_n1227_ = new_n865_ & new_n876_;
  assign new_n1228_ = ~new_n865_ & ~new_n876_;
  assign new_n1229_ = ~new_n1227_ & ~new_n1228_;
  assign new_n1230_ = new_n1138_ & ~new_n1229_;
  assign new_n1231_ = ~new_n1226_ & ~new_n1230_;
  assign new_n1232_ = new_n400_ & ~new_n1231_;
  assign new_n1233_ = p_116_46_ & new_n402_;
  assign new_n1234_ = new_n414_ & new_n959_;
  assign new_n1235_ = ~new_n1232_ & ~new_n1233_;
  assign p_828_2233_ = ~new_n1234_ & new_n1235_;
  assign new_n1237_ = new_n451_ & ~p_828_2233_;
  assign new_n1238_ = ~new_n1197_ & ~new_n1221_;
  assign new_n1239_ = ~new_n1222_ & new_n1238_;
  assign new_n1240_ = ~new_n1237_ & new_n1239_;
  assign p_648_2295_ = p_137_63_ & ~new_n1240_;
  assign new_n1242_ = p_54_20_ & ~new_n430_;
  assign new_n1243_ = ~p_54_20_ & new_n430_;
  assign new_n1244_ = ~new_n1242_ & ~new_n1243_;
  assign new_n1245_ = new_n400_ & ~new_n1244_;
  assign new_n1246_ = p_131_59_ & new_n402_;
  assign new_n1247_ = new_n414_ & new_n977_;
  assign new_n1248_ = ~new_n1245_ & ~new_n1246_;
  assign p_822_1933_ = ~new_n1247_ & new_n1248_;
  assign new_n1250_ = p_4088_172_ & p_4087_171_;
  assign new_n1251_ = p_17_4_ & new_n1250_;
  assign new_n1252_ = p_4088_172_ & ~p_4087_171_;
  assign new_n1253_ = ~p_875_2125_ & new_n1252_;
  assign new_n1254_ = ~p_4088_172_ & p_4087_171_;
  assign new_n1255_ = p_73_25_ & new_n1254_;
  assign new_n1256_ = ~p_4088_172_ & ~p_4087_171_;
  assign new_n1257_ = ~p_836_2128_ & new_n1256_;
  assign new_n1258_ = ~new_n1251_ & ~new_n1253_;
  assign new_n1259_ = ~new_n1255_ & new_n1258_;
  assign p_757_2190_ = new_n1257_ | ~new_n1259_;
  assign new_n1261_ = p_61_21_ & new_n1250_;
  assign new_n1262_ = p_4_1_ & new_n394_;
  assign new_n1263_ = ~p_4_1_ & ~new_n394_;
  assign new_n1264_ = ~new_n1262_ & ~new_n1263_;
  assign new_n1265_ = new_n400_ & ~new_n1264_;
  assign new_n1266_ = p_117_47_ & new_n402_;
  assign new_n1267_ = ~p_3548_166_ & ~p_281_108_;
  assign new_n1268_ = ~p_3546_165_ & p_281_108_;
  assign new_n1269_ = ~p_374_134_ & ~new_n1267_;
  assign new_n1270_ = ~new_n1268_ & new_n1269_;
  assign new_n1271_ = ~p_3550_167_ & ~p_281_108_;
  assign new_n1272_ = p_374_134_ & new_n1271_;
  assign new_n1273_ = ~p_3552_168_ & new_n666_;
  assign new_n1274_ = ~new_n1272_ & ~new_n1273_;
  assign new_n1275_ = ~new_n1270_ & new_n1274_;
  assign new_n1276_ = new_n414_ & new_n1275_;
  assign new_n1277_ = ~new_n1265_ & ~new_n1266_;
  assign p_861_2070_ = ~new_n1276_ & new_n1277_;
  assign new_n1279_ = new_n1252_ & ~p_861_2070_;
  assign new_n1280_ = p_11_2_ & new_n1254_;
  assign new_n1281_ = ~p_822_1933_ & new_n1256_;
  assign new_n1282_ = ~new_n1261_ & ~new_n1279_;
  assign new_n1283_ = ~new_n1280_ & new_n1282_;
  assign p_722_2131_ = new_n1281_ | ~new_n1283_;
  assign new_n1285_ = p_4090_174_ & p_4089_173_;
  assign new_n1286_ = p_70_24_ & new_n1285_;
  assign new_n1287_ = ~p_4090_174_ & p_4089_173_;
  assign new_n1288_ = ~p_877_2126_ & new_n1287_;
  assign new_n1289_ = p_4090_174_ & ~p_4089_173_;
  assign new_n1290_ = p_67_23_ & new_n1289_;
  assign new_n1291_ = ~p_4090_174_ & ~p_4089_173_;
  assign new_n1292_ = ~p_838_2064_ & new_n1291_;
  assign new_n1293_ = ~new_n1286_ & ~new_n1288_;
  assign new_n1294_ = ~new_n1290_ & new_n1293_;
  assign p_802_2183_ = new_n1292_ | ~new_n1294_;
  assign new_n1296_ = ~new_n316_ & new_n329_;
  assign new_n1297_ = new_n316_ & ~new_n329_;
  assign new_n1298_ = ~new_n1296_ & ~new_n1297_;
  assign new_n1299_ = ~new_n304_ & new_n320_;
  assign new_n1300_ = new_n304_ & ~new_n320_;
  assign new_n1301_ = ~new_n1299_ & ~new_n1300_;
  assign new_n1302_ = new_n1298_ & ~new_n1301_;
  assign new_n1303_ = ~new_n1298_ & new_n1301_;
  assign new_n1304_ = ~new_n1302_ & ~new_n1303_;
  assign new_n1305_ = new_n310_ & ~new_n368_;
  assign new_n1306_ = ~new_n310_ & new_n368_;
  assign new_n1307_ = ~new_n1305_ & ~new_n1306_;
  assign new_n1308_ = p_335_123_ & p_292_111_;
  assign new_n1309_ = ~p_335_123_ & p_289_110_;
  assign new_n1310_ = ~new_n1308_ & ~new_n1309_;
  assign new_n1311_ = new_n350_ & ~new_n1310_;
  assign new_n1312_ = ~new_n350_ & new_n1310_;
  assign new_n1313_ = ~new_n1311_ & ~new_n1312_;
  assign new_n1314_ = new_n356_ & ~new_n362_;
  assign new_n1315_ = ~new_n356_ & new_n362_;
  assign new_n1316_ = ~new_n1314_ & ~new_n1315_;
  assign new_n1317_ = ~new_n1307_ & ~new_n1313_;
  assign new_n1318_ = ~new_n1316_ & new_n1317_;
  assign new_n1319_ = new_n1313_ & ~new_n1316_;
  assign new_n1320_ = new_n1307_ & new_n1319_;
  assign new_n1321_ = ~new_n1318_ & ~new_n1320_;
  assign new_n1322_ = new_n1307_ & ~new_n1313_;
  assign new_n1323_ = new_n1316_ & new_n1322_;
  assign new_n1324_ = new_n1313_ & new_n1316_;
  assign new_n1325_ = ~new_n1307_ & new_n1324_;
  assign new_n1326_ = ~new_n1323_ & ~new_n1325_;
  assign new_n1327_ = new_n1321_ & new_n1326_;
  assign new_n1328_ = new_n1304_ & ~new_n1327_;
  assign new_n1329_ = ~new_n1304_ & new_n1327_;
  assign p_1000_2168_ = new_n1328_ | new_n1329_;
  assign new_n1331_ = p_167_74_ & new_n457_;
  assign new_n1332_ = new_n733_ & ~p_867_2237_;
  assign new_n1333_ = p_197_84_ & new_n735_;
  assign new_n1334_ = new_n1034_ & ~p_828_2233_;
  assign new_n1335_ = ~new_n1331_ & ~new_n1332_;
  assign new_n1336_ = ~new_n1333_ & new_n1335_;
  assign new_n1337_ = ~new_n1334_ & new_n1336_;
  assign p_682_2296_ = p_137_63_ & ~new_n1337_;
  assign new_n1339_ = p_20_5_ & new_n1285_;
  assign new_n1340_ = ~new_n323_ & new_n473_;
  assign new_n1341_ = p_4_1_ & new_n1340_;
  assign new_n1342_ = ~new_n478_ & ~new_n1341_;
  assign new_n1343_ = ~new_n480_ & new_n1342_;
  assign new_n1344_ = ~new_n340_ & new_n1343_;
  assign new_n1345_ = new_n307_ & ~new_n1344_;
  assign new_n1346_ = ~new_n307_ & new_n1344_;
  assign new_n1347_ = ~new_n1345_ & ~new_n1346_;
  assign new_n1348_ = new_n400_ & ~new_n1347_;
  assign new_n1349_ = p_128_56_ & new_n402_;
  assign new_n1350_ = ~p_257_102_ & ~p_3548_166_;
  assign new_n1351_ = p_257_102_ & ~p_3546_165_;
  assign new_n1352_ = ~p_389_136_ & ~new_n1350_;
  assign new_n1353_ = ~new_n1351_ & new_n1352_;
  assign new_n1354_ = ~p_257_102_ & ~p_3550_167_;
  assign new_n1355_ = p_389_136_ & new_n1354_;
  assign new_n1356_ = ~p_3552_168_ & new_n676_;
  assign new_n1357_ = ~new_n1355_ & ~new_n1356_;
  assign new_n1358_ = ~new_n1353_ & new_n1357_;
  assign new_n1359_ = new_n414_ & new_n1358_;
  assign new_n1360_ = ~new_n1348_ & ~new_n1349_;
  assign p_873_2124_ = ~new_n1359_ & new_n1360_;
  assign new_n1362_ = new_n1287_ & ~p_873_2124_;
  assign new_n1363_ = p_76_26_ & new_n1289_;
  assign new_n1364_ = ~new_n748_ & new_n771_;
  assign new_n1365_ = p_54_20_ & new_n1364_;
  assign new_n1366_ = ~new_n776_ & ~new_n1365_;
  assign new_n1367_ = ~new_n778_ & new_n1366_;
  assign new_n1368_ = ~new_n761_ & new_n1367_;
  assign new_n1369_ = new_n742_ & ~new_n1368_;
  assign new_n1370_ = ~new_n742_ & new_n1368_;
  assign new_n1371_ = ~new_n1369_ & ~new_n1370_;
  assign new_n1372_ = new_n400_ & ~new_n1371_;
  assign new_n1373_ = p_130_58_ & new_n402_;
  assign new_n1374_ = ~p_514_147_ & p_3546_165_;
  assign new_n1375_ = p_514_147_ & ~p_3552_168_;
  assign new_n1376_ = ~new_n1374_ & ~new_n1375_;
  assign new_n1377_ = new_n414_ & new_n1376_;
  assign new_n1378_ = ~new_n1372_ & ~new_n1373_;
  assign p_834_2123_ = ~new_n1377_ & new_n1378_;
  assign new_n1380_ = new_n1291_ & ~p_834_2123_;
  assign new_n1381_ = ~new_n1339_ & ~new_n1362_;
  assign new_n1382_ = ~new_n1363_ & new_n1381_;
  assign p_792_2188_ = new_n1380_ | ~new_n1382_;
  assign new_n1384_ = new_n859_ & ~new_n865_;
  assign new_n1385_ = new_n856_ & new_n1384_;
  assign new_n1386_ = ~new_n871_ & new_n1385_;
  assign new_n1387_ = ~new_n852_ & new_n1386_;
  assign p_629_1926_ = ~new_n1100_ | new_n1387_;
  assign new_n1389_ = p_49_17_ & new_n1285_;
  assign new_n1390_ = ~new_n553_ & ~new_n554_;
  assign new_n1391_ = ~new_n382_ & new_n1390_;
  assign new_n1392_ = new_n365_ & ~new_n1391_;
  assign new_n1393_ = ~new_n365_ & new_n1391_;
  assign new_n1394_ = ~new_n1392_ & ~new_n1393_;
  assign new_n1395_ = ~new_n1117_ & ~new_n1394_;
  assign new_n1396_ = new_n365_ & new_n555_;
  assign new_n1397_ = ~new_n365_ & ~new_n555_;
  assign new_n1398_ = ~new_n1396_ & ~new_n1397_;
  assign new_n1399_ = new_n1117_ & new_n1398_;
  assign new_n1400_ = ~new_n1395_ & ~new_n1399_;
  assign new_n1401_ = new_n400_ & ~new_n1400_;
  assign new_n1402_ = p_114_44_ & new_n402_;
  assign new_n1403_ = ~p_210_89_ & ~p_3548_166_;
  assign new_n1404_ = p_210_89_ & ~p_3546_165_;
  assign new_n1405_ = ~p_457_142_ & ~new_n1403_;
  assign new_n1406_ = ~new_n1404_ & new_n1405_;
  assign new_n1407_ = ~p_210_89_ & ~p_3550_167_;
  assign new_n1408_ = p_457_142_ & new_n1407_;
  assign new_n1409_ = ~p_3552_168_ & new_n640_;
  assign new_n1410_ = ~new_n1408_ & ~new_n1409_;
  assign new_n1411_ = ~new_n1406_ & new_n1410_;
  assign new_n1412_ = new_n414_ & new_n1411_;
  assign new_n1413_ = ~new_n1401_ & ~new_n1402_;
  assign p_865_2277_ = ~new_n1412_ & new_n1413_;
  assign new_n1415_ = new_n1287_ & ~p_865_2277_;
  assign new_n1416_ = p_46_16_ & new_n1289_;
  assign new_n1417_ = ~new_n882_ & ~new_n883_;
  assign new_n1418_ = ~new_n874_ & new_n1417_;
  assign new_n1419_ = ~new_n856_ & ~new_n1418_;
  assign new_n1420_ = new_n856_ & new_n1418_;
  assign new_n1421_ = ~new_n1419_ & ~new_n1420_;
  assign new_n1422_ = ~new_n1138_ & ~new_n1421_;
  assign new_n1423_ = ~new_n856_ & new_n884_;
  assign new_n1424_ = new_n856_ & ~new_n884_;
  assign new_n1425_ = ~new_n1423_ & ~new_n1424_;
  assign new_n1426_ = new_n1138_ & new_n1425_;
  assign new_n1427_ = ~new_n1422_ & ~new_n1426_;
  assign new_n1428_ = new_n400_ & ~new_n1427_;
  assign new_n1429_ = p_121_51_ & new_n402_;
  assign new_n1430_ = new_n414_ & new_n965_;
  assign new_n1431_ = ~new_n1428_ & ~new_n1429_;
  assign p_826_2275_ = ~new_n1430_ & new_n1431_;
  assign new_n1433_ = new_n1291_ & ~p_826_2275_;
  assign new_n1434_ = ~new_n1389_ & ~new_n1415_;
  assign new_n1435_ = ~new_n1416_ & new_n1434_;
  assign p_772_2299_ = new_n1433_ | ~new_n1435_;
  assign new_n1437_ = p_17_4_ & new_n1285_;
  assign new_n1438_ = ~p_875_2125_ & new_n1287_;
  assign new_n1439_ = p_73_25_ & new_n1289_;
  assign new_n1440_ = ~p_836_2128_ & new_n1291_;
  assign new_n1441_ = ~new_n1437_ & ~new_n1438_;
  assign new_n1442_ = ~new_n1439_ & new_n1441_;
  assign p_797_2191_ = new_n1440_ | ~new_n1442_;
  assign new_n1444_ = p_185_80_ & new_n390_;
  assign new_n1445_ = new_n418_ & ~p_861_2070_;
  assign new_n1446_ = p_182_79_ & new_n420_;
  assign new_n1447_ = new_n451_ & ~p_822_1933_;
  assign new_n1448_ = ~new_n1444_ & ~new_n1445_;
  assign new_n1449_ = ~new_n1446_ & new_n1448_;
  assign new_n1450_ = ~new_n1447_ & new_n1449_;
  assign p_661_2178_ = p_137_63_ & ~new_n1450_;
  assign new_n1452_ = p_106_40_ & new_n1250_;
  assign new_n1453_ = ~p_863_2276_ & new_n1252_;
  assign new_n1454_ = p_109_41_ & new_n1254_;
  assign new_n1455_ = ~p_824_2274_ & new_n1256_;
  assign new_n1456_ = ~new_n1452_ & ~new_n1453_;
  assign new_n1457_ = ~new_n1454_ & new_n1456_;
  assign p_727_2298_ = new_n1455_ | ~new_n1457_;
  assign new_n1459_ = ~p_324_120_ & ~p_3548_166_;
  assign new_n1460_ = p_324_120_ & ~p_3546_165_;
  assign new_n1461_ = ~p_503_146_ & ~new_n1459_;
  assign new_n1462_ = ~new_n1460_ & new_n1461_;
  assign new_n1463_ = ~p_324_120_ & ~p_3550_167_;
  assign new_n1464_ = p_503_146_ & new_n1463_;
  assign new_n1465_ = ~p_3552_168_ & new_n987_;
  assign new_n1466_ = ~new_n1464_ & ~new_n1465_;
  assign new_n1467_ = ~new_n1462_ & new_n1466_;
  assign new_n1468_ = ~new_n1079_ & ~new_n1467_;
  assign new_n1469_ = ~new_n1376_ & new_n1468_;
  assign new_n1470_ = ~new_n447_ & new_n1469_;
  assign new_n1471_ = ~new_n959_ & new_n968_;
  assign new_n1472_ = ~new_n965_ & new_n1471_;
  assign new_n1473_ = ~new_n949_ & new_n1472_;
  assign new_n1474_ = ~new_n977_ & new_n1470_;
  assign p_598_1623_ = new_n1473_ & new_n1474_;
  assign p_634_665_ = p_373_133_ & p_1_0_;
  assign new_n1477_ = p_86_32_ & ~p_2358_162_;
  assign new_n1478_ = p_87_33_ & p_2358_162_;
  assign new_n1479_ = ~new_n1477_ & ~new_n1478_;
  assign p_636_1280_ = p_809_655_ | new_n1479_;
  assign new_n1481_ = p_40_14_ & new_n1250_;
  assign new_n1482_ = ~p_869_2181_ & new_n1252_;
  assign new_n1483_ = p_91_35_ & new_n1254_;
  assign new_n1484_ = new_n871_ & ~new_n1138_;
  assign new_n1485_ = ~new_n871_ & new_n1138_;
  assign new_n1486_ = ~new_n1484_ & ~new_n1485_;
  assign new_n1487_ = new_n400_ & ~new_n1486_;
  assign new_n1488_ = p_112_42_ & new_n402_;
  assign new_n1489_ = new_n414_ & new_n949_;
  assign new_n1490_ = ~new_n1487_ & ~new_n1488_;
  assign p_830_2182_ = ~new_n1489_ & new_n1490_;
  assign new_n1492_ = new_n1256_ & ~p_830_2182_;
  assign new_n1493_ = ~new_n1481_ & ~new_n1482_;
  assign new_n1494_ = ~new_n1483_ & new_n1493_;
  assign p_742_2238_ = new_n1492_ | ~new_n1494_;
  assign new_n1496_ = p_64_22_ & new_n1250_;
  assign new_n1497_ = ~new_n732_ & new_n1252_;
  assign new_n1498_ = p_14_3_ & new_n1254_;
  assign new_n1499_ = ~new_n1033_ & new_n1256_;
  assign new_n1500_ = ~new_n1496_ & ~new_n1497_;
  assign new_n1501_ = ~new_n1498_ & new_n1500_;
  assign p_767_2479_ = new_n1499_ | ~new_n1501_;
  assign new_n1503_ = p_185_80_ & new_n457_;
  assign new_n1504_ = new_n733_ & ~p_861_2070_;
  assign new_n1505_ = p_182_79_ & new_n735_;
  assign new_n1506_ = new_n1034_ & ~p_822_1933_;
  assign new_n1507_ = ~new_n1503_ & ~new_n1504_;
  assign new_n1508_ = ~new_n1505_ & new_n1507_;
  assign new_n1509_ = ~new_n1506_ & new_n1508_;
  assign p_693_2179_ = p_137_63_ & ~new_n1509_;
  assign new_n1511_ = p_146_67_ & new_n457_;
  assign new_n1512_ = new_n733_ & ~p_873_2124_;
  assign new_n1513_ = p_149_68_ & new_n735_;
  assign new_n1514_ = new_n1034_ & ~p_834_2123_;
  assign new_n1515_ = ~new_n1511_ & ~new_n1512_;
  assign new_n1516_ = ~new_n1513_ & new_n1515_;
  assign new_n1517_ = ~new_n1514_ & new_n1516_;
  assign p_702_2228_ = p_137_63_ & ~new_n1517_;
  assign new_n1519_ = p_64_22_ & new_n1285_;
  assign new_n1520_ = ~new_n732_ & new_n1287_;
  assign new_n1521_ = p_14_3_ & new_n1289_;
  assign new_n1522_ = ~new_n1033_ & new_n1291_;
  assign new_n1523_ = ~new_n1519_ & ~new_n1520_;
  assign new_n1524_ = ~new_n1521_ & new_n1523_;
  assign p_807_2480_ = new_n1522_ | ~new_n1524_;
  assign new_n1526_ = p_161_72_ & new_n390_;
  assign new_n1527_ = new_n418_ & ~p_863_2276_;
  assign new_n1528_ = p_191_82_ & new_n420_;
  assign new_n1529_ = new_n451_ & ~p_824_2274_;
  assign new_n1530_ = ~new_n1526_ & ~new_n1527_;
  assign new_n1531_ = ~new_n1528_ & new_n1530_;
  assign new_n1532_ = ~new_n1529_ & new_n1531_;
  assign p_654_2315_ = p_137_63_ & ~new_n1532_;
  assign new_n1534_ = p_179_78_ & new_n390_;
  assign new_n1535_ = new_n418_ & ~new_n732_;
  assign new_n1536_ = p_176_77_ & new_n420_;
  assign new_n1537_ = new_n451_ & ~new_n1033_;
  assign new_n1538_ = ~new_n1534_ & ~new_n1535_;
  assign new_n1539_ = ~new_n1536_ & new_n1538_;
  assign new_n1540_ = ~new_n1537_ & new_n1539_;
  assign p_658_2483_ = ~p_137_63_ | new_n1540_;
  assign new_n1542_ = p_83_31_ & ~p_2358_162_;
  assign new_n1543_ = p_83_31_ & p_2358_162_;
  assign new_n1544_ = ~new_n1542_ & ~new_n1543_;
  assign p_820_1283_ = p_809_655_ | new_n1544_;
  assign new_n1546_ = p_164_73_ & new_n457_;
  assign new_n1547_ = new_n733_ & ~p_865_2277_;
  assign new_n1548_ = p_194_83_ & new_n735_;
  assign new_n1549_ = new_n1034_ & ~p_826_2275_;
  assign new_n1550_ = ~new_n1546_ & ~new_n1547_;
  assign new_n1551_ = ~new_n1548_ & new_n1550_;
  assign new_n1552_ = ~new_n1549_ & new_n1551_;
  assign p_685_2316_ = p_137_63_ & ~new_n1552_;
  assign p_815_627_ = p_136_62_ & ~p_3173_164_;
  assign new_n1555_ = p_4091_175_ & p_4092_176_;
  assign new_n1556_ = new_n400_ & ~new_n609_;
  assign new_n1557_ = p_118_48_ & new_n402_;
  assign new_n1558_ = new_n414_ & new_n728_;
  assign new_n1559_ = ~new_n1555_ & ~new_n1556_;
  assign new_n1560_ = ~new_n1557_ & new_n1559_;
  assign p_882_2456_ = new_n1558_ | ~new_n1560_;
  assign new_n1562_ = ~new_n353_ & ~new_n371_;
  assign new_n1563_ = ~new_n359_ & new_n1562_;
  assign new_n1564_ = ~new_n365_ & new_n1563_;
  assign new_n1565_ = ~new_n347_ & new_n1564_;
  assign p_621_1893_ = ~new_n388_ | new_n1565_;
  assign new_n1567_ = p_170_75_ & new_n457_;
  assign new_n1568_ = ~new_n307_ & ~new_n333_;
  assign new_n1569_ = ~new_n394_ & new_n1568_;
  assign new_n1570_ = ~new_n323_ & new_n1569_;
  assign new_n1571_ = p_4_1_ & new_n1570_;
  assign new_n1572_ = ~new_n462_ & ~new_n1571_;
  assign new_n1573_ = ~new_n466_ & new_n1572_;
  assign new_n1574_ = ~new_n468_ & new_n1573_;
  assign new_n1575_ = ~new_n338_ & new_n1574_;
  assign new_n1576_ = new_n313_ & ~new_n1575_;
  assign new_n1577_ = ~new_n313_ & new_n1575_;
  assign new_n1578_ = ~new_n1576_ & ~new_n1577_;
  assign new_n1579_ = new_n400_ & ~new_n1578_;
  assign new_n1580_ = p_122_52_ & new_n402_;
  assign new_n1581_ = ~p_234_95_ & ~p_3548_166_;
  assign new_n1582_ = p_234_95_ & ~p_3546_165_;
  assign new_n1583_ = ~p_435_140_ & ~new_n1581_;
  assign new_n1584_ = ~new_n1582_ & new_n1583_;
  assign new_n1585_ = ~p_3550_167_ & ~p_234_95_;
  assign new_n1586_ = p_435_140_ & new_n1585_;
  assign new_n1587_ = ~p_3552_168_ & new_n686_;
  assign new_n1588_ = ~new_n1586_ & ~new_n1587_;
  assign new_n1589_ = ~new_n1584_ & new_n1588_;
  assign new_n1590_ = new_n414_ & new_n1589_;
  assign new_n1591_ = ~new_n1579_ & ~new_n1580_;
  assign p_871_2127_ = ~new_n1590_ & new_n1591_;
  assign new_n1593_ = new_n733_ & ~p_871_2127_;
  assign new_n1594_ = p_200_85_ & new_n735_;
  assign new_n1595_ = ~new_n427_ & ~new_n742_;
  assign new_n1596_ = new_n430_ & new_n1595_;
  assign new_n1597_ = ~new_n748_ & new_n1596_;
  assign new_n1598_ = p_54_20_ & new_n1597_;
  assign new_n1599_ = ~new_n757_ & ~new_n1598_;
  assign new_n1600_ = ~new_n762_ & new_n1599_;
  assign new_n1601_ = ~new_n765_ & new_n1600_;
  assign new_n1602_ = ~new_n766_ & new_n1601_;
  assign new_n1603_ = new_n754_ & ~new_n1602_;
  assign new_n1604_ = ~new_n754_ & new_n1602_;
  assign new_n1605_ = ~new_n1603_ & ~new_n1604_;
  assign new_n1606_ = new_n400_ & ~new_n1605_;
  assign new_n1607_ = p_52_18_ & new_n402_;
  assign new_n1608_ = new_n414_ & new_n1467_;
  assign new_n1609_ = ~new_n1606_ & ~new_n1607_;
  assign p_832_2133_ = ~new_n1608_ & new_n1609_;
  assign new_n1611_ = new_n1034_ & ~p_832_2133_;
  assign new_n1612_ = ~new_n1567_ & ~new_n1593_;
  assign new_n1613_ = ~new_n1594_ & new_n1612_;
  assign new_n1614_ = ~new_n1611_ & new_n1613_;
  assign p_676_2229_ = p_137_63_ & ~new_n1614_;
  assign new_n1616_ = p_152_69_ & new_n390_;
  assign new_n1617_ = new_n418_ & ~p_875_2125_;
  assign new_n1618_ = p_155_70_ & new_n420_;
  assign new_n1619_ = new_n451_ & ~p_836_2128_;
  assign new_n1620_ = ~new_n1616_ & ~new_n1617_;
  assign new_n1621_ = ~new_n1618_ & new_n1620_;
  assign new_n1622_ = ~new_n1619_ & new_n1621_;
  assign p_667_2224_ = p_137_63_ & ~new_n1622_;
  assign new_n1624_ = p_158_71_ & new_n457_;
  assign new_n1625_ = ~p_877_2126_ & new_n733_;
  assign new_n1626_ = p_188_81_ & new_n735_;
  assign new_n1627_ = ~p_838_2064_ & new_n1034_;
  assign new_n1628_ = ~new_n1624_ & ~new_n1625_;
  assign new_n1629_ = ~new_n1626_ & new_n1628_;
  assign new_n1630_ = ~new_n1627_ & new_n1629_;
  assign p_696_2226_ = p_137_63_ & ~new_n1630_;
  assign new_n1632_ = p_37_13_ & new_n1285_;
  assign new_n1633_ = new_n1287_ & ~p_871_2127_;
  assign new_n1634_ = p_43_15_ & new_n1289_;
  assign new_n1635_ = new_n1291_ & ~p_832_2133_;
  assign new_n1636_ = ~new_n1632_ & ~new_n1633_;
  assign new_n1637_ = ~new_n1634_ & new_n1636_;
  assign p_787_2186_ = new_n1635_ | ~new_n1637_;
  assign new_n1639_ = p_308_116_ & ~p_316_118_;
  assign new_n1640_ = ~p_308_116_ & p_316_118_;
  assign new_n1641_ = ~new_n1639_ & ~new_n1640_;
  assign new_n1642_ = p_293_112_ & ~p_302_114_;
  assign new_n1643_ = ~p_293_112_ & p_302_114_;
  assign new_n1644_ = ~new_n1642_ & ~new_n1643_;
  assign new_n1645_ = new_n1641_ & ~new_n1644_;
  assign new_n1646_ = ~new_n1641_ & new_n1644_;
  assign new_n1647_ = ~new_n1645_ & ~new_n1646_;
  assign new_n1648_ = ~p_369_131_ & p_361_129_;
  assign new_n1649_ = p_369_131_ & ~p_361_129_;
  assign new_n1650_ = ~new_n1648_ & ~new_n1649_;
  assign new_n1651_ = ~p_351_127_ & p_341_125_;
  assign new_n1652_ = p_351_127_ & ~p_341_125_;
  assign new_n1653_ = ~new_n1651_ & ~new_n1652_;
  assign new_n1654_ = ~p_324_120_ & ~new_n1650_;
  assign new_n1655_ = ~new_n1653_ & new_n1654_;
  assign new_n1656_ = p_324_120_ & ~new_n1653_;
  assign new_n1657_ = new_n1650_ & new_n1656_;
  assign new_n1658_ = ~new_n1655_ & ~new_n1657_;
  assign new_n1659_ = ~p_324_120_ & new_n1650_;
  assign new_n1660_ = new_n1653_ & new_n1659_;
  assign new_n1661_ = p_324_120_ & new_n1653_;
  assign new_n1662_ = ~new_n1650_ & new_n1661_;
  assign new_n1663_ = ~new_n1660_ & ~new_n1662_;
  assign new_n1664_ = new_n1658_ & new_n1663_;
  assign new_n1665_ = new_n1647_ & ~new_n1664_;
  assign new_n1666_ = ~new_n1647_ & new_n1664_;
  assign p_1002_1920_ = new_n1665_ | new_n1666_;
  assign new_n1668_ = ~p_226_93_ & p_218_91_;
  assign new_n1669_ = p_226_93_ & ~p_218_91_;
  assign new_n1670_ = ~new_n1668_ & ~new_n1669_;
  assign new_n1671_ = ~p_210_89_ & p_206_87_;
  assign new_n1672_ = p_210_89_ & ~p_206_87_;
  assign new_n1673_ = ~new_n1671_ & ~new_n1672_;
  assign new_n1674_ = new_n1670_ & ~new_n1673_;
  assign new_n1675_ = ~new_n1670_ & new_n1673_;
  assign new_n1676_ = ~new_n1674_ & ~new_n1675_;
  assign new_n1677_ = ~p_289_110_ & p_281_108_;
  assign new_n1678_ = p_289_110_ & ~p_281_108_;
  assign new_n1679_ = ~new_n1677_ & ~new_n1678_;
  assign new_n1680_ = ~p_257_102_ & p_234_95_;
  assign new_n1681_ = p_257_102_ & ~p_234_95_;
  assign new_n1682_ = ~new_n1680_ & ~new_n1681_;
  assign new_n1683_ = ~p_273_106_ & p_265_104_;
  assign new_n1684_ = p_273_106_ & ~p_265_104_;
  assign new_n1685_ = ~new_n1683_ & ~new_n1684_;
  assign new_n1686_ = ~new_n1679_ & ~new_n1682_;
  assign new_n1687_ = ~new_n1685_ & new_n1686_;
  assign new_n1688_ = new_n1682_ & ~new_n1685_;
  assign new_n1689_ = new_n1679_ & new_n1688_;
  assign new_n1690_ = ~new_n1687_ & ~new_n1689_;
  assign new_n1691_ = new_n1679_ & ~new_n1682_;
  assign new_n1692_ = new_n1685_ & new_n1691_;
  assign new_n1693_ = new_n1682_ & new_n1685_;
  assign new_n1694_ = ~new_n1679_ & new_n1693_;
  assign new_n1695_ = ~new_n1692_ & ~new_n1694_;
  assign new_n1696_ = new_n1690_ & new_n1695_;
  assign new_n1697_ = new_n1676_ & ~new_n1696_;
  assign new_n1698_ = ~new_n1676_ & new_n1696_;
  assign p_1004_1977_ = new_n1697_ | new_n1698_;
  assign new_n1700_ = p_146_67_ & new_n390_;
  assign new_n1701_ = new_n418_ & ~p_873_2124_;
  assign new_n1702_ = p_149_68_ & new_n420_;
  assign new_n1703_ = new_n451_ & ~p_834_2123_;
  assign new_n1704_ = ~new_n1700_ & ~new_n1701_;
  assign new_n1705_ = ~new_n1702_ & new_n1704_;
  assign new_n1706_ = ~new_n1703_ & new_n1705_;
  assign p_670_2225_ = p_137_63_ & ~new_n1706_;
  assign new_n1708_ = p_106_40_ & new_n1285_;
  assign new_n1709_ = ~p_863_2276_ & new_n1287_;
  assign new_n1710_ = p_109_41_ & new_n1289_;
  assign new_n1711_ = ~p_824_2274_ & new_n1291_;
  assign new_n1712_ = ~new_n1708_ & ~new_n1709_;
  assign new_n1713_ = ~new_n1710_ & new_n1712_;
  assign p_712_2297_ = new_n1711_ | ~new_n1713_;
  assign new_n1715_ = p_2358_162_ & p_809_655_;
  assign new_n1716_ = p_2358_162_ & ~p_809_655_;
  assign new_n1717_ = p_80_28_ & new_n1716_;
  assign new_n1718_ = ~p_2358_162_ & p_809_655_;
  assign new_n1719_ = ~p_2358_162_ & ~p_809_655_;
  assign new_n1720_ = p_82_30_ & new_n1719_;
  assign new_n1721_ = ~new_n1715_ & ~new_n1717_;
  assign new_n1722_ = ~new_n1718_ & new_n1721_;
  assign new_n1723_ = ~new_n1720_ & new_n1722_;
  assign p_715_1278_ = p_141_65_ & ~new_n1723_;
  assign new_n1725_ = new_n400_ & ~new_n938_;
  assign new_n1726_ = p_120_50_ & new_n402_;
  assign new_n1727_ = new_n414_ & new_n1029_;
  assign new_n1728_ = ~new_n1555_ & ~new_n1725_;
  assign new_n1729_ = ~new_n1726_ & new_n1728_;
  assign p_843_2455_ = new_n1727_ | ~new_n1729_;
  assign new_n1731_ = p_61_21_ & new_n1285_;
  assign new_n1732_ = ~p_861_2070_ & new_n1287_;
  assign new_n1733_ = p_11_2_ & new_n1289_;
  assign new_n1734_ = ~p_822_1933_ & new_n1291_;
  assign new_n1735_ = ~new_n1731_ & ~new_n1732_;
  assign new_n1736_ = ~new_n1733_ & new_n1735_;
  assign p_859_2132_ = new_n1734_ | ~new_n1736_;
  assign p_810_356_ = p_145_66_ & p_141_65_;
  assign new_n1739_ = p_170_75_ & new_n390_;
  assign new_n1740_ = new_n418_ & ~p_871_2127_;
  assign new_n1741_ = p_200_85_ & new_n420_;
  assign new_n1742_ = new_n451_ & ~p_832_2133_;
  assign new_n1743_ = ~new_n1739_ & ~new_n1740_;
  assign new_n1744_ = ~new_n1741_ & new_n1743_;
  assign new_n1745_ = ~new_n1742_ & new_n1744_;
  assign p_642_2222_ = p_137_63_ & ~new_n1745_;
  assign new_n1747_ = p_103_39_ & new_n1285_;
  assign new_n1748_ = ~p_867_2237_ & new_n1287_;
  assign new_n1749_ = p_100_38_ & new_n1289_;
  assign new_n1750_ = ~p_828_2233_ & new_n1291_;
  assign new_n1751_ = ~new_n1747_ & ~new_n1748_;
  assign new_n1752_ = ~new_n1749_ & new_n1751_;
  assign p_777_2278_ = new_n1750_ | ~new_n1752_;
  assign p_626_1752_ = new_n838_ & new_n1386_;
  assign p_632_1692_ = new_n1115_ & new_n1564_;
  assign new_n1756_ = p_173_76_ & new_n390_;
  assign new_n1757_ = new_n418_ & ~p_869_2181_;
  assign new_n1758_ = p_203_86_ & new_n420_;
  assign new_n1759_ = new_n451_ & ~p_830_2182_;
  assign new_n1760_ = ~new_n1756_ & ~new_n1757_;
  assign new_n1761_ = ~new_n1758_ & new_n1760_;
  assign new_n1762_ = ~new_n1759_ & new_n1761_;
  assign p_645_2271_ = p_137_63_ & ~new_n1762_;
  assign new_n1764_ = p_173_76_ & new_n457_;
  assign new_n1765_ = new_n733_ & ~p_869_2181_;
  assign new_n1766_ = p_203_86_ & new_n735_;
  assign new_n1767_ = new_n1034_ & ~p_830_2182_;
  assign new_n1768_ = ~new_n1764_ & ~new_n1765_;
  assign new_n1769_ = ~new_n1766_ & new_n1768_;
  assign new_n1770_ = ~new_n1767_ & new_n1769_;
  assign p_679_2272_ = p_137_63_ & ~new_n1770_;
  assign new_n1772_ = p_23_6_ & new_n1716_;
  assign new_n1773_ = p_79_27_ & new_n1719_;
  assign new_n1774_ = ~new_n1715_ & ~new_n1772_;
  assign new_n1775_ = ~new_n1718_ & new_n1774_;
  assign new_n1776_ = ~new_n1773_ & new_n1775_;
  assign p_707_1277_ = p_141_65_ & ~new_n1776_;
  assign new_n1778_ = p_103_39_ & new_n1250_;
  assign new_n1779_ = ~p_867_2237_ & new_n1252_;
  assign new_n1780_ = p_100_38_ & new_n1254_;
  assign new_n1781_ = ~p_828_2233_ & new_n1256_;
  assign new_n1782_ = ~new_n1778_ & ~new_n1779_;
  assign new_n1783_ = ~new_n1780_ & new_n1782_;
  assign p_737_2279_ = new_n1781_ | ~new_n1783_;
  assign new_n1785_ = p_40_14_ & new_n1285_;
  assign new_n1786_ = ~p_869_2181_ & new_n1287_;
  assign new_n1787_ = p_91_35_ & new_n1289_;
  assign new_n1788_ = new_n1291_ & ~p_830_2182_;
  assign new_n1789_ = ~new_n1785_ & ~new_n1786_;
  assign new_n1790_ = ~new_n1787_ & new_n1789_;
  assign p_782_2239_ = new_n1788_ | ~new_n1790_;
  assign new_n1792_ = p_37_13_ & new_n1250_;
  assign new_n1793_ = new_n1252_ & ~p_871_2127_;
  assign new_n1794_ = p_43_15_ & new_n1254_;
  assign new_n1795_ = new_n1256_ & ~p_832_2133_;
  assign new_n1796_ = ~new_n1792_ & ~new_n1793_;
  assign new_n1797_ = ~new_n1794_ & new_n1796_;
  assign p_747_2187_ = new_n1795_ | ~new_n1797_;
  assign p_845_845_ = p_2824_163_ | ~p_27_10_;
  assign new_n1800_ = new_n1371_ & new_n1605_;
  assign new_n1801_ = new_n435_ & new_n1800_;
  assign new_n1802_ = new_n1068_ & new_n1801_;
  assign new_n1803_ = new_n1244_ & new_n1802_;
  assign new_n1804_ = new_n1427_ & new_n1803_;
  assign new_n1805_ = p_623_2152_ & new_n1804_;
  assign new_n1806_ = new_n1486_ & new_n1805_;
  assign p_585_2236_ = new_n1231_ & new_n1806_;
  assign new_n1808_ = p_81_29_ & new_n1716_;
  assign new_n1809_ = p_26_9_ & new_n1719_;
  assign new_n1810_ = ~new_n1715_ & ~new_n1808_;
  assign new_n1811_ = ~new_n1718_ & new_n1810_;
  assign new_n1812_ = ~new_n1809_ & new_n1811_;
  assign p_673_1276_ = p_141_65_ & ~new_n1812_;
  assign new_n1814_ = p_49_17_ & new_n1250_;
  assign new_n1815_ = new_n1252_ & ~p_865_2277_;
  assign new_n1816_ = p_46_16_ & new_n1254_;
  assign new_n1817_ = new_n1256_ & ~p_826_2275_;
  assign new_n1818_ = ~new_n1814_ & ~new_n1815_;
  assign new_n1819_ = ~new_n1816_ & new_n1818_;
  assign p_732_2300_ = new_n1817_ | ~new_n1819_;
  assign new_n1821_ = ~new_n862_ & new_n868_;
  assign new_n1822_ = new_n862_ & ~new_n868_;
  assign new_n1823_ = ~new_n1821_ & ~new_n1822_;
  assign new_n1824_ = new_n856_ & ~new_n859_;
  assign new_n1825_ = ~new_n1095_ & ~new_n1824_;
  assign new_n1826_ = new_n1823_ & ~new_n1825_;
  assign new_n1827_ = ~new_n1823_ & new_n1825_;
  assign new_n1828_ = ~new_n1826_ & ~new_n1827_;
  assign new_n1829_ = ~new_n424_ & new_n745_;
  assign new_n1830_ = new_n424_ & ~new_n745_;
  assign new_n1831_ = ~new_n1829_ & ~new_n1830_;
  assign new_n1832_ = new_n739_ & ~new_n751_;
  assign new_n1833_ = ~new_n739_ & new_n751_;
  assign new_n1834_ = ~new_n1832_ & ~new_n1833_;
  assign new_n1835_ = p_332_122_ & p_372_132_;
  assign new_n1836_ = p_369_131_ & ~p_332_122_;
  assign new_n1837_ = ~new_n1835_ & ~new_n1836_;
  assign new_n1838_ = new_n430_ & ~new_n1837_;
  assign new_n1839_ = ~new_n430_ & new_n1837_;
  assign new_n1840_ = ~new_n1838_ & ~new_n1839_;
  assign new_n1841_ = ~new_n1831_ & ~new_n1834_;
  assign new_n1842_ = ~new_n1840_ & new_n1841_;
  assign new_n1843_ = new_n1834_ & ~new_n1840_;
  assign new_n1844_ = new_n1831_ & new_n1843_;
  assign new_n1845_ = ~new_n1842_ & ~new_n1844_;
  assign new_n1846_ = new_n1831_ & ~new_n1834_;
  assign new_n1847_ = new_n1840_ & new_n1846_;
  assign new_n1848_ = new_n1834_ & new_n1840_;
  assign new_n1849_ = ~new_n1831_ & new_n1848_;
  assign new_n1850_ = ~new_n1847_ & ~new_n1849_;
  assign new_n1851_ = new_n1845_ & new_n1850_;
  assign new_n1852_ = new_n1828_ & ~new_n1851_;
  assign new_n1853_ = ~new_n1828_ & new_n1851_;
  assign p_998_2163_ = new_n1852_ | new_n1853_;
  assign new_n1855_ = ~p_1002_1920_ & ~p_1004_1977_;
  assign new_n1856_ = ~p_998_2163_ & new_n1855_;
  assign new_n1857_ = ~p_1000_2168_ & new_n1856_;
  assign new_n1858_ = p_562_155_ & new_n1857_;
  assign new_n1859_ = p_559_154_ & p_552_152_;
  assign new_n1860_ = p_556_153_ & new_n1859_;
  assign new_n1861_ = p_386_135_ & new_n1860_;
  assign new_n1862_ = p_245_98_ & new_n1858_;
  assign p_854_2268_ = new_n1861_ & new_n1862_;
  assign new_n1864_ = p_20_5_ & new_n1250_;
  assign new_n1865_ = new_n1252_ & ~p_873_2124_;
  assign new_n1866_ = p_76_26_ & new_n1254_;
  assign new_n1867_ = new_n1256_ & ~p_834_2123_;
  assign new_n1868_ = ~new_n1864_ & ~new_n1865_;
  assign new_n1869_ = ~new_n1866_ & new_n1868_;
  assign p_752_2189_ = new_n1867_ | ~new_n1869_;
  assign new_n1871_ = ~new_n413_ & ~new_n1358_;
  assign new_n1872_ = ~new_n1057_ & new_n1871_;
  assign new_n1873_ = ~new_n1275_ & new_n1872_;
  assign new_n1874_ = ~new_n1193_ & ~new_n1411_;
  assign new_n1875_ = ~new_n1217_ & new_n1874_;
  assign new_n1876_ = ~new_n1589_ & new_n1875_;
  assign new_n1877_ = ~new_n653_ & new_n1873_;
  assign p_610_1519_ = new_n1876_ & new_n1877_;
  assign new_n1879_ = ~p_623_2152_ & ~new_n1168_;
  assign new_n1880_ = ~p_623_2152_ & ~new_n1879_;
  assign new_n1881_ = ~new_n1168_ & ~new_n1879_;
  assign p_813_2260_ = new_n1880_ | new_n1881_;
  assign new_n1883_ = new_n1347_ & new_n1578_;
  assign new_n1884_ = new_n399_ & new_n1883_;
  assign new_n1885_ = new_n1046_ & new_n1884_;
  assign new_n1886_ = new_n1264_ & new_n1885_;
  assign new_n1887_ = new_n1400_ & new_n1886_;
  assign new_n1888_ = new_n1126_ & new_n1887_;
  assign new_n1889_ = new_n1182_ & new_n1888_;
  assign p_575_2240_ = new_n1206_ & new_n1889_;
  assign p_601_220_ = p_552_152_ & p_562_155_;
  assign new_n1892_ = p_25_8_ & new_n1716_;
  assign new_n1893_ = p_24_7_ & new_n1719_;
  assign new_n1894_ = ~new_n1715_ & ~new_n1892_;
  assign new_n1895_ = ~new_n1718_ & new_n1894_;
  assign new_n1896_ = ~new_n1893_ & new_n1895_;
  assign p_639_1275_ = p_141_65_ & ~new_n1896_;
  assign new_n1898_ = p_164_73_ & new_n390_;
  assign new_n1899_ = new_n418_ & ~p_865_2277_;
  assign new_n1900_ = p_194_83_ & new_n420_;
  assign new_n1901_ = new_n451_ & ~p_826_2275_;
  assign new_n1902_ = ~new_n1898_ & ~new_n1899_;
  assign new_n1903_ = ~new_n1900_ & new_n1902_;
  assign new_n1904_ = ~new_n1901_ & new_n1903_;
  assign p_651_2314_ = p_137_63_ & ~new_n1904_;
  assign p_656_621_ = ~p_140_64_ | p_809_655_;
  assign new_n1907_ = p_70_24_ & new_n1250_;
  assign new_n1908_ = ~p_877_2126_ & new_n1252_;
  assign new_n1909_ = p_67_23_ & new_n1254_;
  assign new_n1910_ = ~p_838_2064_ & new_n1256_;
  assign new_n1911_ = ~new_n1907_ & ~new_n1908_;
  assign new_n1912_ = ~new_n1909_ & new_n1911_;
  assign p_762_2184_ = new_n1910_ | ~new_n1912_;
  assign p_847_465_ = ~p_556_153_ | ~p_386_135_;
  assign p_604_223_ = ~p_545_150_;
  assign p_593_733_ = ~p_299_113_;
  assign p_600_259_ = ~p_366_130_;
  assign p_611_275_ = ~p_338_124_;
  assign p_606_407_ = ~p_549_151_;
  assign p_612_263_ = ~p_358_128_;
  assign p_849_219_ = ~p_552_152_;
  assign p_850_217_ = ~p_562_155_;
  assign p_599_269_ = ~p_348_126_;
  assign p_851_218_ = ~p_559_154_;
  assign p_848_330_ = ~p_245_98_;
  assign p_973_202_ = p_3173_164_;
  assign p_603_225_ = p_604_223_;
  assign p_921_664_ = p_1_0_;
  assign p_892_408_ = p_549_151_;
  assign p_949_852_ = p_1_0_;
  assign p_939_853_ = p_1_0_;
  assign p_594_224_ = p_604_223_;
  assign p_978_851_ = p_1_0_;
  assign p_926_624_ = p_137_63_;
  assign p_298_299_ = p_293_112_;
  assign p_602_222_ = p_606_407_;
  assign p_717_1282_ = p_704_1281_;
  assign p_887_528_ = p_299_113_;
  assign p_923_619_ = p_141_65_;
  assign p_144_354_ = p_141_65_;
  assign p_889_734_ = p_299_113_;
  assign p_993_850_ = p_1_0_;
endmodule

