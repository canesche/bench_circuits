// Benchmark "testing" written by ABC on Thu Oct  8 22:16:32 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A41  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A41;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[351]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[360]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[370]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[380]_ , \new_[381]_ , \new_[385]_ , \new_[386]_ ,
    \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[392]_ , \new_[396]_ ,
    \new_[397]_ , \new_[398]_ , \new_[402]_ , \new_[403]_ , \new_[407]_ ,
    \new_[408]_ , \new_[409]_ , \new_[410]_ , \new_[413]_ , \new_[417]_ ,
    \new_[418]_ , \new_[419]_ , \new_[423]_ , \new_[424]_ , \new_[428]_ ,
    \new_[429]_ , \new_[430]_ , \new_[431]_ , \new_[432]_ , \new_[433]_ ,
    \new_[436]_ , \new_[440]_ , \new_[441]_ , \new_[442]_ , \new_[446]_ ,
    \new_[447]_ , \new_[451]_ , \new_[452]_ , \new_[453]_ , \new_[454]_ ,
    \new_[457]_ , \new_[461]_ , \new_[462]_ , \new_[463]_ , \new_[467]_ ,
    \new_[468]_ , \new_[472]_ , \new_[473]_ , \new_[474]_ , \new_[475]_ ,
    \new_[476]_ , \new_[479]_ , \new_[483]_ , \new_[484]_ , \new_[485]_ ,
    \new_[489]_ , \new_[490]_ , \new_[494]_ , \new_[495]_ , \new_[496]_ ,
    \new_[497]_ , \new_[500]_ , \new_[504]_ , \new_[505]_ , \new_[506]_ ,
    \new_[510]_ , \new_[511]_ , \new_[515]_ , \new_[516]_ , \new_[517]_ ,
    \new_[518]_ , \new_[519]_ , \new_[520]_ , \new_[521]_ , \new_[524]_ ,
    \new_[528]_ , \new_[529]_ , \new_[530]_ , \new_[533]_ , \new_[537]_ ,
    \new_[538]_ , \new_[539]_ , \new_[540]_ , \new_[543]_ , \new_[547]_ ,
    \new_[548]_ , \new_[549]_ , \new_[553]_ , \new_[554]_ , \new_[558]_ ,
    \new_[559]_ , \new_[560]_ , \new_[561]_ , \new_[562]_ , \new_[565]_ ,
    \new_[569]_ , \new_[570]_ , \new_[571]_ , \new_[575]_ , \new_[576]_ ,
    \new_[580]_ , \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[586]_ ,
    \new_[590]_ , \new_[591]_ , \new_[592]_ , \new_[596]_ , \new_[597]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[609]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[619]_ , \new_[620]_ , \new_[624]_ , \new_[625]_ , \new_[626]_ ,
    \new_[627]_ , \new_[630]_ , \new_[634]_ , \new_[635]_ , \new_[636]_ ,
    \new_[640]_ , \new_[641]_ , \new_[645]_ , \new_[646]_ , \new_[647]_ ,
    \new_[648]_ , \new_[649]_ , \new_[652]_ , \new_[656]_ , \new_[657]_ ,
    \new_[658]_ , \new_[662]_ , \new_[663]_ , \new_[667]_ , \new_[668]_ ,
    \new_[669]_ , \new_[670]_ , \new_[673]_ , \new_[677]_ , \new_[678]_ ,
    \new_[679]_ , \new_[683]_ , \new_[684]_ , \new_[688]_ , \new_[689]_ ,
    \new_[690]_ , \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[694]_ ,
    \new_[695]_ , \new_[698]_ , \new_[702]_ , \new_[703]_ , \new_[704]_ ,
    \new_[707]_ , \new_[711]_ , \new_[712]_ , \new_[713]_ , \new_[714]_ ,
    \new_[717]_ , \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[727]_ ,
    \new_[728]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[736]_ , \new_[739]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ ,
    \new_[749]_ , \new_[750]_ , \new_[754]_ , \new_[755]_ , \new_[756]_ ,
    \new_[757]_ , \new_[760]_ , \new_[764]_ , \new_[765]_ , \new_[766]_ ,
    \new_[770]_ , \new_[771]_ , \new_[775]_ , \new_[776]_ , \new_[777]_ ,
    \new_[778]_ , \new_[779]_ , \new_[780]_ , \new_[783]_ , \new_[787]_ ,
    \new_[788]_ , \new_[789]_ , \new_[793]_ , \new_[794]_ , \new_[798]_ ,
    \new_[799]_ , \new_[800]_ , \new_[801]_ , \new_[804]_ , \new_[808]_ ,
    \new_[809]_ , \new_[810]_ , \new_[814]_ , \new_[815]_ , \new_[819]_ ,
    \new_[820]_ , \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[826]_ ,
    \new_[830]_ , \new_[831]_ , \new_[832]_ , \new_[836]_ , \new_[837]_ ,
    \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[847]_ ,
    \new_[851]_ , \new_[852]_ , \new_[853]_ , \new_[857]_ , \new_[858]_ ,
    \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[865]_ , \new_[866]_ ,
    \new_[867]_ , \new_[868]_ , \new_[871]_ , \new_[875]_ , \new_[876]_ ,
    \new_[877]_ , \new_[880]_ , \new_[884]_ , \new_[885]_ , \new_[886]_ ,
    \new_[887]_ , \new_[890]_ , \new_[894]_ , \new_[895]_ , \new_[896]_ ,
    \new_[900]_ , \new_[901]_ , \new_[905]_ , \new_[906]_ , \new_[907]_ ,
    \new_[908]_ , \new_[909]_ , \new_[912]_ , \new_[916]_ , \new_[917]_ ,
    \new_[918]_ , \new_[922]_ , \new_[923]_ , \new_[927]_ , \new_[928]_ ,
    \new_[929]_ , \new_[930]_ , \new_[933]_ , \new_[937]_ , \new_[938]_ ,
    \new_[939]_ , \new_[943]_ , \new_[944]_ , \new_[948]_ , \new_[949]_ ,
    \new_[950]_ , \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[956]_ ,
    \new_[960]_ , \new_[961]_ , \new_[962]_ , \new_[966]_ , \new_[967]_ ,
    \new_[971]_ , \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[977]_ ,
    \new_[981]_ , \new_[982]_ , \new_[983]_ , \new_[987]_ , \new_[988]_ ,
    \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ , \new_[996]_ ,
    \new_[999]_ , \new_[1003]_ , \new_[1004]_ , \new_[1005]_ ,
    \new_[1009]_ , \new_[1010]_ , \new_[1014]_ , \new_[1015]_ ,
    \new_[1016]_ , \new_[1017]_ , \new_[1020]_ , \new_[1024]_ ,
    \new_[1025]_ , \new_[1026]_ , \new_[1030]_ , \new_[1031]_ ,
    \new_[1035]_ , \new_[1036]_ , \new_[1037]_ , \new_[1038]_ ,
    \new_[1039]_ , \new_[1040]_ , \new_[1041]_ , \new_[1042]_ ,
    \new_[1049]_ , \new_[1052]_ , \new_[1055]_ , \new_[1058]_ ,
    \new_[1061]_ , \new_[1064]_ , \new_[1067]_ , \new_[1070]_ ,
    \new_[1073]_ , \new_[1076]_ , \new_[1079]_ , \new_[1082]_ ,
    \new_[1085]_ , \new_[1088]_ , \new_[1091]_ , \new_[1094]_ ,
    \new_[1097]_ , \new_[1100]_ , \new_[1103]_ , \new_[1106]_ ,
    \new_[1110]_ , \new_[1111]_ , \new_[1115]_ , \new_[1116]_ ,
    \new_[1120]_ , \new_[1121]_ , \new_[1125]_ , \new_[1126]_ ,
    \new_[1130]_ , \new_[1131]_ , \new_[1135]_ , \new_[1136]_ ,
    \new_[1140]_ , \new_[1141]_ , \new_[1145]_ , \new_[1146]_ ,
    \new_[1150]_ , \new_[1151]_ , \new_[1155]_ , \new_[1156]_ ,
    \new_[1160]_ , \new_[1161]_ , \new_[1165]_ , \new_[1166]_ ,
    \new_[1170]_ , \new_[1171]_ , \new_[1175]_ , \new_[1176]_ ,
    \new_[1180]_ , \new_[1181]_ , \new_[1185]_ , \new_[1186]_ ,
    \new_[1190]_ , \new_[1191]_ , \new_[1195]_ , \new_[1196]_ ,
    \new_[1200]_ , \new_[1201]_ , \new_[1205]_ , \new_[1206]_ ,
    \new_[1210]_ , \new_[1211]_ , \new_[1215]_ , \new_[1216]_ ,
    \new_[1220]_ , \new_[1221]_ , \new_[1225]_ , \new_[1226]_ ,
    \new_[1230]_ , \new_[1231]_ , \new_[1235]_ , \new_[1236]_ ,
    \new_[1240]_ , \new_[1241]_ , \new_[1245]_ , \new_[1246]_ ,
    \new_[1250]_ , \new_[1251]_ , \new_[1255]_ , \new_[1256]_ ,
    \new_[1260]_ , \new_[1261]_ , \new_[1265]_ , \new_[1266]_ ,
    \new_[1270]_ , \new_[1271]_ , \new_[1275]_ , \new_[1276]_ ,
    \new_[1280]_ , \new_[1281]_ , \new_[1285]_ , \new_[1286]_ ,
    \new_[1290]_ , \new_[1291]_ , \new_[1295]_ , \new_[1296]_ ,
    \new_[1300]_ , \new_[1301]_ , \new_[1305]_ , \new_[1306]_ ,
    \new_[1310]_ , \new_[1311]_ , \new_[1315]_ , \new_[1316]_ ,
    \new_[1320]_ , \new_[1321]_ , \new_[1325]_ , \new_[1326]_ ,
    \new_[1330]_ , \new_[1331]_ , \new_[1335]_ , \new_[1336]_ ,
    \new_[1340]_ , \new_[1341]_ , \new_[1345]_ , \new_[1346]_ ,
    \new_[1350]_ , \new_[1351]_ , \new_[1355]_ , \new_[1356]_ ,
    \new_[1360]_ , \new_[1361]_ , \new_[1365]_ , \new_[1366]_ ,
    \new_[1370]_ , \new_[1371]_ , \new_[1375]_ , \new_[1376]_ ,
    \new_[1380]_ , \new_[1381]_ , \new_[1385]_ , \new_[1386]_ ,
    \new_[1390]_ , \new_[1391]_ , \new_[1395]_ , \new_[1396]_ ,
    \new_[1400]_ , \new_[1401]_ , \new_[1405]_ , \new_[1406]_ ,
    \new_[1410]_ , \new_[1411]_ , \new_[1415]_ , \new_[1416]_ ,
    \new_[1420]_ , \new_[1421]_ , \new_[1425]_ , \new_[1426]_ ,
    \new_[1430]_ , \new_[1431]_ , \new_[1435]_ , \new_[1436]_ ,
    \new_[1440]_ , \new_[1441]_ , \new_[1445]_ , \new_[1446]_ ,
    \new_[1450]_ , \new_[1451]_ , \new_[1455]_ , \new_[1456]_ ,
    \new_[1460]_ , \new_[1461]_ , \new_[1465]_ , \new_[1466]_ ,
    \new_[1470]_ , \new_[1471]_ , \new_[1474]_ , \new_[1477]_ ,
    \new_[1478]_ , \new_[1482]_ , \new_[1483]_ , \new_[1486]_ ,
    \new_[1489]_ , \new_[1490]_ , \new_[1494]_ , \new_[1495]_ ,
    \new_[1498]_ , \new_[1501]_ , \new_[1502]_ , \new_[1506]_ ,
    \new_[1507]_ , \new_[1510]_ , \new_[1513]_ , \new_[1514]_ ,
    \new_[1518]_ , \new_[1519]_ , \new_[1522]_ , \new_[1525]_ ,
    \new_[1526]_ , \new_[1530]_ , \new_[1531]_ , \new_[1534]_ ,
    \new_[1537]_ , \new_[1538]_ , \new_[1542]_ , \new_[1543]_ ,
    \new_[1546]_ , \new_[1549]_ , \new_[1550]_ , \new_[1554]_ ,
    \new_[1555]_ , \new_[1558]_ , \new_[1561]_ , \new_[1562]_ ,
    \new_[1565]_ , \new_[1568]_ , \new_[1569]_ , \new_[1572]_ ,
    \new_[1575]_ , \new_[1576]_ , \new_[1579]_ , \new_[1582]_ ,
    \new_[1583]_ , \new_[1586]_ , \new_[1589]_ , \new_[1590]_ ,
    \new_[1593]_ , \new_[1596]_ , \new_[1597]_ , \new_[1600]_ ,
    \new_[1603]_ , \new_[1604]_ , \new_[1607]_ , \new_[1610]_ ,
    \new_[1611]_ , \new_[1614]_ , \new_[1617]_ , \new_[1618]_ ,
    \new_[1621]_ , \new_[1624]_ , \new_[1625]_ , \new_[1628]_ ,
    \new_[1631]_ , \new_[1632]_ , \new_[1635]_ , \new_[1638]_ ,
    \new_[1639]_ , \new_[1642]_ , \new_[1645]_ , \new_[1646]_ ,
    \new_[1649]_ , \new_[1652]_ , \new_[1653]_ , \new_[1656]_ ,
    \new_[1659]_ , \new_[1660]_ , \new_[1663]_ , \new_[1666]_ ,
    \new_[1667]_ , \new_[1670]_ , \new_[1673]_ , \new_[1674]_ ,
    \new_[1677]_ , \new_[1680]_ , \new_[1681]_ , \new_[1684]_ ,
    \new_[1687]_ , \new_[1688]_ , \new_[1691]_ , \new_[1694]_ ,
    \new_[1695]_ , \new_[1698]_ , \new_[1701]_ , \new_[1702]_ ,
    \new_[1705]_ , \new_[1708]_ , \new_[1709]_ , \new_[1712]_ ,
    \new_[1715]_ , \new_[1716]_ , \new_[1719]_ , \new_[1722]_ ,
    \new_[1723]_ , \new_[1726]_ , \new_[1729]_ , \new_[1730]_ ,
    \new_[1733]_ , \new_[1736]_ , \new_[1737]_ , \new_[1740]_ ,
    \new_[1743]_ , \new_[1744]_ , \new_[1747]_ , \new_[1750]_ ,
    \new_[1751]_ , \new_[1754]_ , \new_[1757]_ , \new_[1758]_ ,
    \new_[1761]_ , \new_[1764]_ , \new_[1765]_ , \new_[1768]_ ,
    \new_[1771]_ , \new_[1772]_ , \new_[1775]_ , \new_[1778]_ ,
    \new_[1779]_ , \new_[1782]_ , \new_[1785]_ , \new_[1786]_ ,
    \new_[1789]_ , \new_[1792]_ , \new_[1793]_ , \new_[1796]_ ,
    \new_[1799]_ , \new_[1800]_ , \new_[1803]_ , \new_[1806]_ ,
    \new_[1807]_ , \new_[1810]_ , \new_[1813]_ , \new_[1814]_ ,
    \new_[1817]_ , \new_[1820]_ , \new_[1821]_ , \new_[1824]_ ,
    \new_[1827]_ , \new_[1828]_ , \new_[1831]_ , \new_[1834]_ ,
    \new_[1835]_ , \new_[1838]_ , \new_[1841]_ , \new_[1842]_ ,
    \new_[1845]_ , \new_[1848]_ , \new_[1849]_ , \new_[1852]_ ,
    \new_[1855]_ , \new_[1856]_ , \new_[1859]_ , \new_[1862]_ ,
    \new_[1863]_ , \new_[1866]_ , \new_[1869]_ , \new_[1870]_ ,
    \new_[1873]_ , \new_[1876]_ , \new_[1877]_ , \new_[1880]_ ,
    \new_[1883]_ , \new_[1884]_ , \new_[1887]_ , \new_[1890]_ ,
    \new_[1891]_ , \new_[1894]_ , \new_[1897]_ , \new_[1898]_ ,
    \new_[1901]_ , \new_[1904]_ , \new_[1905]_ , \new_[1908]_ ,
    \new_[1911]_ , \new_[1912]_ , \new_[1915]_ , \new_[1918]_ ,
    \new_[1919]_ , \new_[1922]_ , \new_[1925]_ , \new_[1926]_ ,
    \new_[1929]_ , \new_[1932]_ , \new_[1933]_ , \new_[1936]_ ,
    \new_[1939]_ , \new_[1940]_ , \new_[1943]_ , \new_[1946]_ ,
    \new_[1947]_ , \new_[1950]_ , \new_[1953]_ , \new_[1954]_ ,
    \new_[1957]_ , \new_[1960]_ , \new_[1961]_ , \new_[1964]_ ,
    \new_[1967]_ , \new_[1968]_ , \new_[1971]_ , \new_[1974]_ ,
    \new_[1975]_ , \new_[1978]_ , \new_[1981]_ , \new_[1982]_ ,
    \new_[1985]_ , \new_[1988]_ , \new_[1989]_ , \new_[1992]_ ,
    \new_[1995]_ , \new_[1996]_ , \new_[1999]_ , \new_[2002]_ ,
    \new_[2003]_ , \new_[2006]_ , \new_[2009]_ , \new_[2010]_ ,
    \new_[2013]_ , \new_[2016]_ , \new_[2017]_ , \new_[2020]_ ,
    \new_[2023]_ , \new_[2024]_ , \new_[2027]_ , \new_[2030]_ ,
    \new_[2031]_ , \new_[2034]_ , \new_[2037]_ , \new_[2038]_ ,
    \new_[2041]_ , \new_[2044]_ , \new_[2045]_ , \new_[2048]_ ,
    \new_[2051]_ , \new_[2052]_ , \new_[2055]_ , \new_[2058]_ ,
    \new_[2059]_ , \new_[2062]_ , \new_[2065]_ , \new_[2066]_ ,
    \new_[2069]_ , \new_[2072]_ , \new_[2073]_ , \new_[2076]_ ,
    \new_[2079]_ , \new_[2080]_ , \new_[2083]_ , \new_[2086]_ ,
    \new_[2087]_ , \new_[2090]_ , \new_[2093]_ , \new_[2094]_ ,
    \new_[2097]_ , \new_[2100]_ , \new_[2101]_ , \new_[2104]_ ,
    \new_[2107]_ , \new_[2108]_ , \new_[2111]_ , \new_[2114]_ ,
    \new_[2115]_ , \new_[2118]_ , \new_[2121]_ , \new_[2122]_ ,
    \new_[2125]_ , \new_[2128]_ , \new_[2129]_ , \new_[2132]_ ,
    \new_[2135]_ , \new_[2136]_ , \new_[2139]_ , \new_[2142]_ ,
    \new_[2143]_ , \new_[2146]_ , \new_[2149]_ , \new_[2150]_ ,
    \new_[2153]_ , \new_[2156]_ , \new_[2157]_ , \new_[2160]_ ,
    \new_[2163]_ , \new_[2164]_ , \new_[2167]_ , \new_[2170]_ ,
    \new_[2171]_ , \new_[2174]_ , \new_[2177]_ , \new_[2178]_ ,
    \new_[2181]_ , \new_[2184]_ , \new_[2185]_ , \new_[2188]_ ,
    \new_[2191]_ , \new_[2192]_ , \new_[2195]_ , \new_[2198]_ ,
    \new_[2199]_ , \new_[2202]_ , \new_[2205]_ , \new_[2206]_ ,
    \new_[2209]_ , \new_[2212]_ , \new_[2213]_ , \new_[2216]_ ,
    \new_[2219]_ , \new_[2220]_ , \new_[2223]_ , \new_[2226]_ ,
    \new_[2227]_ , \new_[2230]_ , \new_[2233]_ , \new_[2234]_ ,
    \new_[2237]_ , \new_[2240]_ , \new_[2241]_ , \new_[2244]_ ,
    \new_[2247]_ , \new_[2248]_ , \new_[2251]_ , \new_[2254]_ ,
    \new_[2255]_ , \new_[2258]_ , \new_[2261]_ , \new_[2262]_ ,
    \new_[2265]_ , \new_[2268]_ , \new_[2269]_ , \new_[2272]_ ,
    \new_[2275]_ , \new_[2276]_ , \new_[2279]_ , \new_[2282]_ ,
    \new_[2283]_ , \new_[2286]_ , \new_[2289]_ , \new_[2290]_ ,
    \new_[2293]_ , \new_[2296]_ , \new_[2297]_ , \new_[2300]_ ,
    \new_[2303]_ , \new_[2304]_ , \new_[2307]_ , \new_[2310]_ ,
    \new_[2311]_ , \new_[2314]_ , \new_[2317]_ , \new_[2318]_ ,
    \new_[2321]_ , \new_[2324]_ , \new_[2325]_ , \new_[2328]_ ,
    \new_[2331]_ , \new_[2332]_ , \new_[2335]_ , \new_[2338]_ ,
    \new_[2339]_ , \new_[2342]_ , \new_[2345]_ , \new_[2346]_ ,
    \new_[2349]_ , \new_[2352]_ , \new_[2353]_ , \new_[2356]_ ,
    \new_[2359]_ , \new_[2360]_ , \new_[2363]_ , \new_[2366]_ ,
    \new_[2367]_ , \new_[2370]_ , \new_[2373]_ , \new_[2374]_ ,
    \new_[2377]_ , \new_[2380]_ , \new_[2381]_ , \new_[2384]_ ,
    \new_[2387]_ , \new_[2388]_ , \new_[2391]_ , \new_[2394]_ ,
    \new_[2395]_ , \new_[2398]_ , \new_[2401]_ , \new_[2402]_ ,
    \new_[2405]_ , \new_[2408]_ , \new_[2409]_ , \new_[2412]_ ,
    \new_[2415]_ , \new_[2416]_ , \new_[2419]_ , \new_[2422]_ ,
    \new_[2423]_ , \new_[2426]_ , \new_[2429]_ , \new_[2430]_ ,
    \new_[2433]_ , \new_[2436]_ , \new_[2437]_ , \new_[2440]_ ,
    \new_[2443]_ , \new_[2444]_ , \new_[2447]_ , \new_[2450]_ ,
    \new_[2451]_ , \new_[2454]_ , \new_[2457]_ , \new_[2458]_ ,
    \new_[2461]_ , \new_[2464]_ , \new_[2465]_ , \new_[2468]_ ,
    \new_[2471]_ , \new_[2472]_ , \new_[2475]_ , \new_[2478]_ ,
    \new_[2479]_ , \new_[2482]_ , \new_[2485]_ , \new_[2486]_ ,
    \new_[2489]_ , \new_[2492]_ , \new_[2493]_ , \new_[2496]_ ,
    \new_[2499]_ , \new_[2500]_ , \new_[2503]_ , \new_[2506]_ ,
    \new_[2507]_ , \new_[2510]_ , \new_[2513]_ , \new_[2514]_ ,
    \new_[2517]_ , \new_[2520]_ , \new_[2521]_ , \new_[2524]_ ,
    \new_[2527]_ , \new_[2528]_ , \new_[2531]_ , \new_[2534]_ ,
    \new_[2535]_ , \new_[2538]_ , \new_[2541]_ , \new_[2542]_ ,
    \new_[2545]_ , \new_[2548]_ , \new_[2549]_ , \new_[2552]_ ,
    \new_[2555]_ , \new_[2556]_ , \new_[2559]_ , \new_[2562]_ ,
    \new_[2563]_ , \new_[2566]_ , \new_[2569]_ , \new_[2570]_ ,
    \new_[2573]_ , \new_[2576]_ , \new_[2577]_ , \new_[2580]_ ,
    \new_[2583]_ , \new_[2584]_ , \new_[2587]_ , \new_[2590]_ ,
    \new_[2591]_ , \new_[2594]_ , \new_[2597]_ , \new_[2598]_ ,
    \new_[2601]_ , \new_[2604]_ , \new_[2605]_ , \new_[2608]_ ,
    \new_[2611]_ , \new_[2612]_ , \new_[2615]_ , \new_[2618]_ ,
    \new_[2619]_ , \new_[2622]_ , \new_[2625]_ , \new_[2626]_ ,
    \new_[2629]_ , \new_[2632]_ , \new_[2633]_ , \new_[2636]_ ,
    \new_[2639]_ , \new_[2640]_ , \new_[2643]_ , \new_[2646]_ ,
    \new_[2647]_ , \new_[2650]_ , \new_[2653]_ , \new_[2654]_ ,
    \new_[2657]_ , \new_[2660]_ , \new_[2661]_ , \new_[2664]_ ,
    \new_[2667]_ , \new_[2668]_ , \new_[2671]_ , \new_[2674]_ ,
    \new_[2675]_ , \new_[2678]_ , \new_[2681]_ , \new_[2682]_ ,
    \new_[2685]_ , \new_[2688]_ , \new_[2689]_ , \new_[2692]_ ,
    \new_[2695]_ , \new_[2696]_ , \new_[2699]_ , \new_[2702]_ ,
    \new_[2703]_ , \new_[2706]_ , \new_[2709]_ , \new_[2710]_ ,
    \new_[2713]_ , \new_[2716]_ , \new_[2717]_ , \new_[2720]_ ,
    \new_[2723]_ , \new_[2724]_ , \new_[2727]_ , \new_[2730]_ ,
    \new_[2731]_ , \new_[2734]_ , \new_[2737]_ , \new_[2738]_ ,
    \new_[2741]_ , \new_[2744]_ , \new_[2745]_ , \new_[2748]_ ,
    \new_[2752]_ , \new_[2753]_ , \new_[2754]_ , \new_[2757]_ ,
    \new_[2760]_ , \new_[2761]_ , \new_[2764]_ , \new_[2768]_ ,
    \new_[2769]_ , \new_[2770]_ , \new_[2773]_ , \new_[2776]_ ,
    \new_[2777]_ , \new_[2780]_ , \new_[2784]_ , \new_[2785]_ ,
    \new_[2786]_ , \new_[2789]_ , \new_[2792]_ , \new_[2793]_ ,
    \new_[2796]_ , \new_[2800]_ , \new_[2801]_ , \new_[2802]_ ,
    \new_[2805]_ , \new_[2808]_ , \new_[2809]_ , \new_[2812]_ ,
    \new_[2816]_ , \new_[2817]_ , \new_[2818]_ , \new_[2821]_ ,
    \new_[2824]_ , \new_[2825]_ , \new_[2828]_ , \new_[2832]_ ,
    \new_[2833]_ , \new_[2834]_ , \new_[2837]_ , \new_[2840]_ ,
    \new_[2841]_ , \new_[2844]_ , \new_[2848]_ , \new_[2849]_ ,
    \new_[2850]_ , \new_[2853]_ , \new_[2856]_ , \new_[2857]_ ,
    \new_[2860]_ , \new_[2864]_ , \new_[2865]_ , \new_[2866]_ ,
    \new_[2869]_ , \new_[2872]_ , \new_[2873]_ , \new_[2876]_ ,
    \new_[2880]_ , \new_[2881]_ , \new_[2882]_ , \new_[2885]_ ,
    \new_[2888]_ , \new_[2889]_ , \new_[2892]_ , \new_[2896]_ ,
    \new_[2897]_ , \new_[2898]_ , \new_[2901]_ , \new_[2904]_ ,
    \new_[2905]_ , \new_[2908]_ , \new_[2912]_ , \new_[2913]_ ,
    \new_[2914]_ , \new_[2917]_ , \new_[2920]_ , \new_[2921]_ ,
    \new_[2924]_ , \new_[2928]_ , \new_[2929]_ , \new_[2930]_ ,
    \new_[2933]_ , \new_[2936]_ , \new_[2937]_ , \new_[2940]_ ,
    \new_[2944]_ , \new_[2945]_ , \new_[2946]_ , \new_[2949]_ ,
    \new_[2952]_ , \new_[2953]_ , \new_[2956]_ , \new_[2960]_ ,
    \new_[2961]_ , \new_[2962]_ , \new_[2965]_ , \new_[2968]_ ,
    \new_[2969]_ , \new_[2972]_ , \new_[2976]_ , \new_[2977]_ ,
    \new_[2978]_ , \new_[2981]_ , \new_[2984]_ , \new_[2985]_ ,
    \new_[2988]_ , \new_[2992]_ , \new_[2993]_ , \new_[2994]_ ,
    \new_[2997]_ , \new_[3000]_ , \new_[3001]_ , \new_[3004]_ ,
    \new_[3008]_ , \new_[3009]_ , \new_[3010]_ , \new_[3013]_ ,
    \new_[3016]_ , \new_[3017]_ , \new_[3020]_ , \new_[3024]_ ,
    \new_[3025]_ , \new_[3026]_ , \new_[3029]_ , \new_[3032]_ ,
    \new_[3033]_ , \new_[3036]_ , \new_[3040]_ , \new_[3041]_ ,
    \new_[3042]_ , \new_[3045]_ , \new_[3048]_ , \new_[3049]_ ,
    \new_[3052]_ , \new_[3056]_ , \new_[3057]_ , \new_[3058]_ ,
    \new_[3061]_ , \new_[3064]_ , \new_[3065]_ , \new_[3068]_ ,
    \new_[3072]_ , \new_[3073]_ , \new_[3074]_ , \new_[3077]_ ,
    \new_[3080]_ , \new_[3081]_ , \new_[3084]_ , \new_[3088]_ ,
    \new_[3089]_ , \new_[3090]_ , \new_[3093]_ , \new_[3096]_ ,
    \new_[3097]_ , \new_[3100]_ , \new_[3104]_ , \new_[3105]_ ,
    \new_[3106]_ , \new_[3109]_ , \new_[3112]_ , \new_[3113]_ ,
    \new_[3116]_ , \new_[3120]_ , \new_[3121]_ , \new_[3122]_ ,
    \new_[3125]_ , \new_[3128]_ , \new_[3129]_ , \new_[3132]_ ,
    \new_[3136]_ , \new_[3137]_ , \new_[3138]_ , \new_[3141]_ ,
    \new_[3144]_ , \new_[3145]_ , \new_[3148]_ , \new_[3152]_ ,
    \new_[3153]_ , \new_[3154]_ , \new_[3157]_ , \new_[3160]_ ,
    \new_[3161]_ , \new_[3164]_ , \new_[3168]_ , \new_[3169]_ ,
    \new_[3170]_ , \new_[3173]_ , \new_[3176]_ , \new_[3177]_ ,
    \new_[3180]_ , \new_[3184]_ , \new_[3185]_ , \new_[3186]_ ,
    \new_[3189]_ , \new_[3192]_ , \new_[3193]_ , \new_[3196]_ ,
    \new_[3200]_ , \new_[3201]_ , \new_[3202]_ , \new_[3205]_ ,
    \new_[3208]_ , \new_[3209]_ , \new_[3212]_ , \new_[3216]_ ,
    \new_[3217]_ , \new_[3218]_ , \new_[3221]_ , \new_[3224]_ ,
    \new_[3225]_ , \new_[3228]_ , \new_[3232]_ , \new_[3233]_ ,
    \new_[3234]_ , \new_[3237]_ , \new_[3240]_ , \new_[3241]_ ,
    \new_[3244]_ , \new_[3248]_ , \new_[3249]_ , \new_[3250]_ ,
    \new_[3253]_ , \new_[3257]_ , \new_[3258]_ , \new_[3259]_ ,
    \new_[3262]_ , \new_[3266]_ , \new_[3267]_ , \new_[3268]_ ,
    \new_[3271]_ , \new_[3275]_ , \new_[3276]_ , \new_[3277]_ ,
    \new_[3280]_ , \new_[3284]_ , \new_[3285]_ , \new_[3286]_ ,
    \new_[3289]_ , \new_[3293]_ , \new_[3294]_ , \new_[3295]_ ,
    \new_[3298]_ , \new_[3302]_ , \new_[3303]_ , \new_[3304]_ ,
    \new_[3307]_ , \new_[3311]_ , \new_[3312]_ , \new_[3313]_ ,
    \new_[3316]_ , \new_[3320]_ , \new_[3321]_ , \new_[3322]_ ,
    \new_[3325]_ , \new_[3329]_ , \new_[3330]_ , \new_[3331]_ ,
    \new_[3334]_ , \new_[3338]_ , \new_[3339]_ , \new_[3340]_ ,
    \new_[3343]_ , \new_[3347]_ , \new_[3348]_ , \new_[3349]_ ,
    \new_[3352]_ , \new_[3356]_ , \new_[3357]_ , \new_[3358]_ ,
    \new_[3361]_ , \new_[3365]_ , \new_[3366]_ , \new_[3367]_ ,
    \new_[3370]_ , \new_[3374]_ , \new_[3375]_ , \new_[3376]_ ,
    \new_[3379]_ , \new_[3383]_ , \new_[3384]_ , \new_[3385]_ ,
    \new_[3388]_ , \new_[3392]_ , \new_[3393]_ , \new_[3394]_ ,
    \new_[3397]_ , \new_[3401]_ , \new_[3402]_ , \new_[3403]_ ,
    \new_[3406]_ , \new_[3410]_ , \new_[3411]_ , \new_[3412]_ ,
    \new_[3415]_ , \new_[3419]_ , \new_[3420]_ , \new_[3421]_ ,
    \new_[3424]_ , \new_[3428]_ , \new_[3429]_ , \new_[3430]_ ,
    \new_[3433]_ , \new_[3437]_ , \new_[3438]_ , \new_[3439]_ ,
    \new_[3442]_ , \new_[3446]_ , \new_[3447]_ , \new_[3448]_ ,
    \new_[3451]_ , \new_[3455]_ , \new_[3456]_ , \new_[3457]_ ,
    \new_[3460]_ , \new_[3464]_ , \new_[3465]_ , \new_[3466]_ ,
    \new_[3469]_ , \new_[3473]_ , \new_[3474]_ , \new_[3475]_ ,
    \new_[3478]_ , \new_[3482]_ , \new_[3483]_ , \new_[3484]_ ,
    \new_[3487]_ , \new_[3491]_ , \new_[3492]_ , \new_[3493]_ ,
    \new_[3496]_ , \new_[3500]_ , \new_[3501]_ , \new_[3502]_ ,
    \new_[3505]_ , \new_[3509]_ , \new_[3510]_ , \new_[3511]_ ,
    \new_[3514]_ , \new_[3518]_ , \new_[3519]_ , \new_[3520]_ ,
    \new_[3523]_ , \new_[3527]_ , \new_[3528]_ , \new_[3529]_ ,
    \new_[3532]_ , \new_[3536]_ , \new_[3537]_ , \new_[3538]_ ,
    \new_[3541]_ , \new_[3545]_ , \new_[3546]_ , \new_[3547]_ ,
    \new_[3550]_ , \new_[3554]_ , \new_[3555]_ , \new_[3556]_ ,
    \new_[3559]_ , \new_[3563]_ , \new_[3564]_ , \new_[3565]_ ,
    \new_[3568]_ , \new_[3572]_ , \new_[3573]_ , \new_[3574]_ ,
    \new_[3577]_ , \new_[3581]_ , \new_[3582]_ , \new_[3583]_ ,
    \new_[3586]_ , \new_[3590]_ , \new_[3591]_ , \new_[3592]_ ,
    \new_[3595]_ , \new_[3599]_ , \new_[3600]_ , \new_[3601]_ ,
    \new_[3604]_ , \new_[3608]_ , \new_[3609]_ , \new_[3610]_ ,
    \new_[3613]_ , \new_[3617]_ , \new_[3618]_ , \new_[3619]_ ,
    \new_[3622]_ , \new_[3626]_ , \new_[3627]_ , \new_[3628]_ ,
    \new_[3631]_ , \new_[3635]_ , \new_[3636]_ , \new_[3637]_ ,
    \new_[3640]_ , \new_[3644]_ , \new_[3645]_ , \new_[3646]_ ,
    \new_[3649]_ , \new_[3653]_ , \new_[3654]_ , \new_[3655]_ ,
    \new_[3658]_ , \new_[3662]_ , \new_[3663]_ , \new_[3664]_ ,
    \new_[3667]_ , \new_[3671]_ , \new_[3672]_ , \new_[3673]_ ,
    \new_[3676]_ , \new_[3680]_ , \new_[3681]_ , \new_[3682]_ ,
    \new_[3685]_ , \new_[3689]_ , \new_[3690]_ , \new_[3691]_ ,
    \new_[3694]_ , \new_[3698]_ , \new_[3699]_ , \new_[3700]_ ,
    \new_[3703]_ , \new_[3707]_ , \new_[3708]_ , \new_[3709]_ ,
    \new_[3712]_ , \new_[3716]_ , \new_[3717]_ , \new_[3718]_ ,
    \new_[3721]_ , \new_[3725]_ , \new_[3726]_ , \new_[3727]_ ,
    \new_[3730]_ , \new_[3734]_ , \new_[3735]_ , \new_[3736]_ ,
    \new_[3739]_ , \new_[3743]_ , \new_[3744]_ , \new_[3745]_ ,
    \new_[3748]_ , \new_[3752]_ , \new_[3753]_ , \new_[3754]_ ,
    \new_[3757]_ , \new_[3761]_ , \new_[3762]_ , \new_[3763]_ ,
    \new_[3766]_ , \new_[3770]_ , \new_[3771]_ , \new_[3772]_ ,
    \new_[3775]_ , \new_[3779]_ , \new_[3780]_ , \new_[3781]_ ,
    \new_[3784]_ , \new_[3788]_ , \new_[3789]_ , \new_[3790]_ ,
    \new_[3793]_ , \new_[3797]_ , \new_[3798]_ , \new_[3799]_ ,
    \new_[3802]_ , \new_[3806]_ , \new_[3807]_ , \new_[3808]_ ,
    \new_[3811]_ , \new_[3815]_ , \new_[3816]_ , \new_[3817]_ ,
    \new_[3820]_ , \new_[3824]_ , \new_[3825]_ , \new_[3826]_ ,
    \new_[3829]_ , \new_[3833]_ , \new_[3834]_ , \new_[3835]_ ,
    \new_[3838]_ , \new_[3842]_ , \new_[3843]_ , \new_[3844]_ ,
    \new_[3847]_ , \new_[3851]_ , \new_[3852]_ , \new_[3853]_ ,
    \new_[3856]_ , \new_[3860]_ , \new_[3861]_ , \new_[3862]_ ,
    \new_[3865]_ , \new_[3869]_ , \new_[3870]_ , \new_[3871]_ ,
    \new_[3874]_ , \new_[3878]_ , \new_[3879]_ , \new_[3880]_ ,
    \new_[3883]_ , \new_[3887]_ , \new_[3888]_ , \new_[3889]_ ,
    \new_[3892]_ , \new_[3896]_ , \new_[3897]_ , \new_[3898]_ ,
    \new_[3901]_ , \new_[3905]_ , \new_[3906]_ , \new_[3907]_ ,
    \new_[3910]_ , \new_[3914]_ , \new_[3915]_ , \new_[3916]_ ,
    \new_[3919]_ , \new_[3923]_ , \new_[3924]_ , \new_[3925]_ ,
    \new_[3928]_ , \new_[3932]_ , \new_[3933]_ , \new_[3934]_ ,
    \new_[3937]_ , \new_[3941]_ , \new_[3942]_ , \new_[3943]_ ,
    \new_[3946]_ , \new_[3950]_ , \new_[3951]_ , \new_[3952]_ ,
    \new_[3955]_ , \new_[3959]_ , \new_[3960]_ , \new_[3961]_ ,
    \new_[3964]_ , \new_[3968]_ , \new_[3969]_ , \new_[3970]_ ,
    \new_[3973]_ , \new_[3977]_ , \new_[3978]_ , \new_[3979]_ ,
    \new_[3982]_ , \new_[3986]_ , \new_[3987]_ , \new_[3988]_ ,
    \new_[3991]_ , \new_[3995]_ , \new_[3996]_ , \new_[3997]_ ,
    \new_[4000]_ , \new_[4004]_ , \new_[4005]_ , \new_[4006]_ ,
    \new_[4009]_ , \new_[4013]_ , \new_[4014]_ , \new_[4015]_ ,
    \new_[4018]_ , \new_[4022]_ , \new_[4023]_ , \new_[4024]_ ,
    \new_[4027]_ , \new_[4031]_ , \new_[4032]_ , \new_[4033]_ ,
    \new_[4036]_ , \new_[4040]_ , \new_[4041]_ , \new_[4042]_ ,
    \new_[4045]_ , \new_[4049]_ , \new_[4050]_ , \new_[4051]_ ,
    \new_[4054]_ , \new_[4058]_ , \new_[4059]_ , \new_[4060]_ ,
    \new_[4063]_ , \new_[4067]_ , \new_[4068]_ , \new_[4069]_ ,
    \new_[4072]_ , \new_[4076]_ , \new_[4077]_ , \new_[4078]_ ,
    \new_[4081]_ , \new_[4085]_ , \new_[4086]_ , \new_[4087]_ ,
    \new_[4090]_ , \new_[4094]_ , \new_[4095]_ , \new_[4096]_ ,
    \new_[4099]_ , \new_[4103]_ , \new_[4104]_ , \new_[4105]_ ,
    \new_[4108]_ , \new_[4112]_ , \new_[4113]_ , \new_[4114]_ ,
    \new_[4117]_ , \new_[4121]_ , \new_[4122]_ , \new_[4123]_ ,
    \new_[4126]_ , \new_[4130]_ , \new_[4131]_ , \new_[4132]_ ,
    \new_[4135]_ , \new_[4139]_ , \new_[4140]_ , \new_[4141]_ ,
    \new_[4144]_ , \new_[4148]_ , \new_[4149]_ , \new_[4150]_ ,
    \new_[4153]_ , \new_[4157]_ , \new_[4158]_ , \new_[4159]_ ,
    \new_[4162]_ , \new_[4166]_ , \new_[4167]_ , \new_[4168]_ ,
    \new_[4171]_ , \new_[4175]_ , \new_[4176]_ , \new_[4177]_ ,
    \new_[4180]_ , \new_[4184]_ , \new_[4185]_ , \new_[4186]_ ,
    \new_[4189]_ , \new_[4193]_ , \new_[4194]_ , \new_[4195]_ ,
    \new_[4198]_ , \new_[4202]_ , \new_[4203]_ , \new_[4204]_ ,
    \new_[4207]_ , \new_[4211]_ , \new_[4212]_ , \new_[4213]_ ,
    \new_[4216]_ , \new_[4220]_ , \new_[4221]_ , \new_[4222]_ ,
    \new_[4225]_ , \new_[4229]_ , \new_[4230]_ , \new_[4231]_ ,
    \new_[4234]_ , \new_[4238]_ , \new_[4239]_ , \new_[4240]_ ,
    \new_[4243]_ , \new_[4247]_ , \new_[4248]_ , \new_[4249]_ ,
    \new_[4252]_ , \new_[4256]_ , \new_[4257]_ , \new_[4258]_ ,
    \new_[4261]_ , \new_[4265]_ , \new_[4266]_ , \new_[4267]_ ,
    \new_[4270]_ , \new_[4274]_ , \new_[4275]_ , \new_[4276]_ ,
    \new_[4279]_ , \new_[4283]_ , \new_[4284]_ , \new_[4285]_ ,
    \new_[4288]_ , \new_[4292]_ , \new_[4293]_ , \new_[4294]_ ,
    \new_[4297]_ , \new_[4301]_ , \new_[4302]_ , \new_[4303]_ ,
    \new_[4306]_ , \new_[4310]_ , \new_[4311]_ , \new_[4312]_ ,
    \new_[4315]_ , \new_[4319]_ , \new_[4320]_ , \new_[4321]_ ,
    \new_[4324]_ , \new_[4328]_ , \new_[4329]_ , \new_[4330]_ ,
    \new_[4333]_ , \new_[4337]_ , \new_[4338]_ , \new_[4339]_ ,
    \new_[4342]_ , \new_[4346]_ , \new_[4347]_ , \new_[4348]_ ,
    \new_[4351]_ , \new_[4355]_ , \new_[4356]_ , \new_[4357]_ ,
    \new_[4360]_ , \new_[4364]_ , \new_[4365]_ , \new_[4366]_ ,
    \new_[4369]_ , \new_[4373]_ , \new_[4374]_ , \new_[4375]_ ,
    \new_[4378]_ , \new_[4382]_ , \new_[4383]_ , \new_[4384]_ ,
    \new_[4387]_ , \new_[4391]_ , \new_[4392]_ , \new_[4393]_ ,
    \new_[4396]_ , \new_[4400]_ , \new_[4401]_ , \new_[4402]_ ,
    \new_[4405]_ , \new_[4409]_ , \new_[4410]_ , \new_[4411]_ ,
    \new_[4414]_ , \new_[4418]_ , \new_[4419]_ , \new_[4420]_ ,
    \new_[4423]_ , \new_[4427]_ , \new_[4428]_ , \new_[4429]_ ,
    \new_[4432]_ , \new_[4436]_ , \new_[4437]_ , \new_[4438]_ ,
    \new_[4441]_ , \new_[4445]_ , \new_[4446]_ , \new_[4447]_ ,
    \new_[4450]_ , \new_[4454]_ , \new_[4455]_ , \new_[4456]_ ,
    \new_[4459]_ , \new_[4463]_ , \new_[4464]_ , \new_[4465]_ ,
    \new_[4468]_ , \new_[4472]_ , \new_[4473]_ , \new_[4474]_ ,
    \new_[4477]_ , \new_[4481]_ , \new_[4482]_ , \new_[4483]_ ,
    \new_[4486]_ , \new_[4490]_ , \new_[4491]_ , \new_[4492]_ ,
    \new_[4495]_ , \new_[4499]_ , \new_[4500]_ , \new_[4501]_ ,
    \new_[4504]_ , \new_[4508]_ , \new_[4509]_ , \new_[4510]_ ,
    \new_[4513]_ , \new_[4517]_ , \new_[4518]_ , \new_[4519]_ ,
    \new_[4522]_ , \new_[4526]_ , \new_[4527]_ , \new_[4528]_ ,
    \new_[4531]_ , \new_[4535]_ , \new_[4536]_ , \new_[4537]_ ,
    \new_[4540]_ , \new_[4544]_ , \new_[4545]_ , \new_[4546]_ ,
    \new_[4549]_ , \new_[4553]_ , \new_[4554]_ , \new_[4555]_ ,
    \new_[4558]_ , \new_[4562]_ , \new_[4563]_ , \new_[4564]_ ,
    \new_[4567]_ , \new_[4571]_ , \new_[4572]_ , \new_[4573]_ ,
    \new_[4576]_ , \new_[4580]_ , \new_[4581]_ , \new_[4582]_ ,
    \new_[4585]_ , \new_[4589]_ , \new_[4590]_ , \new_[4591]_ ,
    \new_[4594]_ , \new_[4598]_ , \new_[4599]_ , \new_[4600]_ ,
    \new_[4603]_ , \new_[4607]_ , \new_[4608]_ , \new_[4609]_ ,
    \new_[4612]_ , \new_[4616]_ , \new_[4617]_ , \new_[4618]_ ,
    \new_[4621]_ , \new_[4625]_ , \new_[4626]_ , \new_[4627]_ ,
    \new_[4630]_ , \new_[4634]_ , \new_[4635]_ , \new_[4636]_ ,
    \new_[4639]_ , \new_[4643]_ , \new_[4644]_ , \new_[4645]_ ,
    \new_[4648]_ , \new_[4652]_ , \new_[4653]_ , \new_[4654]_ ,
    \new_[4657]_ , \new_[4661]_ , \new_[4662]_ , \new_[4663]_ ,
    \new_[4666]_ , \new_[4670]_ , \new_[4671]_ , \new_[4672]_ ,
    \new_[4675]_ , \new_[4679]_ , \new_[4680]_ , \new_[4681]_ ,
    \new_[4684]_ , \new_[4688]_ , \new_[4689]_ , \new_[4690]_ ,
    \new_[4693]_ , \new_[4697]_ , \new_[4698]_ , \new_[4699]_ ,
    \new_[4702]_ , \new_[4706]_ , \new_[4707]_ , \new_[4708]_ ,
    \new_[4711]_ , \new_[4715]_ , \new_[4716]_ , \new_[4717]_ ,
    \new_[4720]_ , \new_[4724]_ , \new_[4725]_ , \new_[4726]_ ,
    \new_[4729]_ , \new_[4733]_ , \new_[4734]_ , \new_[4735]_ ,
    \new_[4738]_ , \new_[4742]_ , \new_[4743]_ , \new_[4744]_ ,
    \new_[4747]_ , \new_[4751]_ , \new_[4752]_ , \new_[4753]_ ,
    \new_[4756]_ , \new_[4760]_ , \new_[4761]_ , \new_[4762]_ ,
    \new_[4765]_ , \new_[4769]_ , \new_[4770]_ , \new_[4771]_ ,
    \new_[4774]_ , \new_[4778]_ , \new_[4779]_ , \new_[4780]_ ,
    \new_[4783]_ , \new_[4787]_ , \new_[4788]_ , \new_[4789]_ ,
    \new_[4792]_ , \new_[4796]_ , \new_[4797]_ , \new_[4798]_ ,
    \new_[4801]_ , \new_[4805]_ , \new_[4806]_ , \new_[4807]_ ,
    \new_[4810]_ , \new_[4814]_ , \new_[4815]_ , \new_[4816]_ ,
    \new_[4819]_ , \new_[4823]_ , \new_[4824]_ , \new_[4825]_ ,
    \new_[4828]_ , \new_[4832]_ , \new_[4833]_ , \new_[4834]_ ,
    \new_[4837]_ , \new_[4841]_ , \new_[4842]_ , \new_[4843]_ ,
    \new_[4846]_ , \new_[4850]_ , \new_[4851]_ , \new_[4852]_ ,
    \new_[4855]_ , \new_[4859]_ , \new_[4860]_ , \new_[4861]_ ,
    \new_[4864]_ , \new_[4868]_ , \new_[4869]_ , \new_[4870]_ ,
    \new_[4873]_ , \new_[4877]_ , \new_[4878]_ , \new_[4879]_ ,
    \new_[4882]_ , \new_[4886]_ , \new_[4887]_ , \new_[4888]_ ,
    \new_[4891]_ , \new_[4895]_ , \new_[4896]_ , \new_[4897]_ ,
    \new_[4900]_ , \new_[4904]_ , \new_[4905]_ , \new_[4906]_ ,
    \new_[4909]_ , \new_[4913]_ , \new_[4914]_ , \new_[4915]_ ,
    \new_[4918]_ , \new_[4922]_ , \new_[4923]_ , \new_[4924]_ ,
    \new_[4927]_ , \new_[4931]_ , \new_[4932]_ , \new_[4933]_ ,
    \new_[4936]_ , \new_[4940]_ , \new_[4941]_ , \new_[4942]_ ,
    \new_[4945]_ , \new_[4949]_ , \new_[4950]_ , \new_[4951]_ ,
    \new_[4954]_ , \new_[4958]_ , \new_[4959]_ , \new_[4960]_ ,
    \new_[4963]_ , \new_[4967]_ , \new_[4968]_ , \new_[4969]_ ,
    \new_[4972]_ , \new_[4976]_ , \new_[4977]_ , \new_[4978]_ ,
    \new_[4981]_ , \new_[4985]_ , \new_[4986]_ , \new_[4987]_ ,
    \new_[4991]_ , \new_[4992]_ , \new_[4996]_ , \new_[4997]_ ,
    \new_[4998]_ , \new_[5001]_ , \new_[5005]_ , \new_[5006]_ ,
    \new_[5007]_ , \new_[5011]_ , \new_[5012]_ , \new_[5016]_ ,
    \new_[5017]_ , \new_[5018]_ , \new_[5021]_ , \new_[5025]_ ,
    \new_[5026]_ , \new_[5027]_ , \new_[5031]_ , \new_[5032]_ ,
    \new_[5036]_ , \new_[5037]_ , \new_[5038]_ , \new_[5041]_ ,
    \new_[5045]_ , \new_[5046]_ , \new_[5047]_ , \new_[5051]_ ,
    \new_[5052]_ , \new_[5056]_ , \new_[5057]_ , \new_[5058]_ ,
    \new_[5061]_ , \new_[5065]_ , \new_[5066]_ , \new_[5067]_ ,
    \new_[5071]_ , \new_[5072]_ , \new_[5076]_ , \new_[5077]_ ,
    \new_[5078]_ , \new_[5081]_ , \new_[5085]_ , \new_[5086]_ ,
    \new_[5087]_ , \new_[5091]_ , \new_[5092]_ , \new_[5096]_ ,
    \new_[5097]_ , \new_[5098]_ , \new_[5101]_ , \new_[5105]_ ,
    \new_[5106]_ , \new_[5107]_ , \new_[5111]_ , \new_[5112]_ ,
    \new_[5116]_ , \new_[5117]_ , \new_[5118]_ , \new_[5121]_ ,
    \new_[5125]_ , \new_[5126]_ , \new_[5127]_ , \new_[5131]_ ,
    \new_[5132]_ , \new_[5136]_ , \new_[5137]_ , \new_[5138]_ ,
    \new_[5141]_ , \new_[5145]_ , \new_[5146]_ , \new_[5147]_ ,
    \new_[5151]_ , \new_[5152]_ , \new_[5156]_ , \new_[5157]_ ,
    \new_[5158]_ , \new_[5161]_ , \new_[5165]_ , \new_[5166]_ ,
    \new_[5167]_ , \new_[5171]_ , \new_[5172]_ , \new_[5176]_ ,
    \new_[5177]_ , \new_[5178]_ , \new_[5181]_ , \new_[5185]_ ,
    \new_[5186]_ , \new_[5187]_ , \new_[5191]_ , \new_[5192]_ ,
    \new_[5196]_ , \new_[5197]_ , \new_[5198]_ , \new_[5201]_ ,
    \new_[5205]_ , \new_[5206]_ , \new_[5207]_ , \new_[5211]_ ,
    \new_[5212]_ , \new_[5216]_ , \new_[5217]_ , \new_[5218]_ ,
    \new_[5221]_ , \new_[5225]_ , \new_[5226]_ , \new_[5227]_ ,
    \new_[5231]_ , \new_[5232]_ , \new_[5236]_ , \new_[5237]_ ,
    \new_[5238]_ , \new_[5241]_ , \new_[5245]_ , \new_[5246]_ ,
    \new_[5247]_ , \new_[5251]_ , \new_[5252]_ , \new_[5256]_ ,
    \new_[5257]_ , \new_[5258]_ , \new_[5261]_ , \new_[5265]_ ,
    \new_[5266]_ , \new_[5267]_ , \new_[5271]_ , \new_[5272]_ ,
    \new_[5276]_ , \new_[5277]_ , \new_[5278]_ , \new_[5281]_ ,
    \new_[5285]_ , \new_[5286]_ , \new_[5287]_ , \new_[5291]_ ,
    \new_[5292]_ , \new_[5296]_ , \new_[5297]_ , \new_[5298]_ ,
    \new_[5301]_ , \new_[5305]_ , \new_[5306]_ , \new_[5307]_ ,
    \new_[5311]_ , \new_[5312]_ , \new_[5316]_ , \new_[5317]_ ,
    \new_[5318]_ , \new_[5321]_ , \new_[5325]_ , \new_[5326]_ ,
    \new_[5327]_ , \new_[5331]_ , \new_[5332]_ , \new_[5336]_ ,
    \new_[5337]_ , \new_[5338]_ , \new_[5341]_ , \new_[5345]_ ,
    \new_[5346]_ , \new_[5347]_ , \new_[5351]_ , \new_[5352]_ ,
    \new_[5356]_ , \new_[5357]_ , \new_[5358]_ , \new_[5361]_ ,
    \new_[5365]_ , \new_[5366]_ , \new_[5367]_ , \new_[5371]_ ,
    \new_[5372]_ , \new_[5376]_ , \new_[5377]_ , \new_[5378]_ ,
    \new_[5381]_ , \new_[5385]_ , \new_[5386]_ , \new_[5387]_ ,
    \new_[5391]_ , \new_[5392]_ , \new_[5396]_ , \new_[5397]_ ,
    \new_[5398]_ , \new_[5401]_ , \new_[5405]_ , \new_[5406]_ ,
    \new_[5407]_ , \new_[5411]_ , \new_[5412]_ , \new_[5416]_ ,
    \new_[5417]_ , \new_[5418]_ , \new_[5421]_ , \new_[5425]_ ,
    \new_[5426]_ , \new_[5427]_ , \new_[5431]_ , \new_[5432]_ ,
    \new_[5436]_ , \new_[5437]_ , \new_[5438]_ , \new_[5441]_ ,
    \new_[5445]_ , \new_[5446]_ , \new_[5447]_ , \new_[5451]_ ,
    \new_[5452]_ , \new_[5456]_ , \new_[5457]_ , \new_[5458]_ ,
    \new_[5461]_ , \new_[5465]_ , \new_[5466]_ , \new_[5467]_ ,
    \new_[5471]_ , \new_[5472]_ , \new_[5476]_ , \new_[5477]_ ,
    \new_[5478]_ , \new_[5481]_ , \new_[5485]_ , \new_[5486]_ ,
    \new_[5487]_ , \new_[5491]_ , \new_[5492]_ , \new_[5496]_ ,
    \new_[5497]_ , \new_[5498]_ , \new_[5501]_ , \new_[5505]_ ,
    \new_[5506]_ , \new_[5507]_ , \new_[5511]_ , \new_[5512]_ ,
    \new_[5516]_ , \new_[5517]_ , \new_[5518]_ , \new_[5521]_ ,
    \new_[5525]_ , \new_[5526]_ , \new_[5527]_ , \new_[5531]_ ,
    \new_[5532]_ , \new_[5536]_ , \new_[5537]_ , \new_[5538]_ ,
    \new_[5541]_ , \new_[5545]_ , \new_[5546]_ , \new_[5547]_ ,
    \new_[5551]_ , \new_[5552]_ , \new_[5556]_ , \new_[5557]_ ,
    \new_[5558]_ , \new_[5561]_ , \new_[5565]_ , \new_[5566]_ ,
    \new_[5567]_ , \new_[5571]_ , \new_[5572]_ , \new_[5576]_ ,
    \new_[5577]_ , \new_[5578]_ , \new_[5581]_ , \new_[5585]_ ,
    \new_[5586]_ , \new_[5587]_ , \new_[5591]_ , \new_[5592]_ ,
    \new_[5596]_ , \new_[5597]_ , \new_[5598]_ , \new_[5601]_ ,
    \new_[5605]_ , \new_[5606]_ , \new_[5607]_ , \new_[5611]_ ,
    \new_[5612]_ , \new_[5616]_ , \new_[5617]_ , \new_[5618]_ ,
    \new_[5622]_ , \new_[5623]_ , \new_[5627]_ , \new_[5628]_ ,
    \new_[5629]_ , \new_[5633]_ , \new_[5634]_ , \new_[5638]_ ,
    \new_[5639]_ , \new_[5640]_ , \new_[5644]_ , \new_[5645]_ ,
    \new_[5649]_ , \new_[5650]_ , \new_[5651]_ , \new_[5655]_ ,
    \new_[5656]_ , \new_[5660]_ , \new_[5661]_ , \new_[5662]_ ,
    \new_[5666]_ , \new_[5667]_ , \new_[5671]_ , \new_[5672]_ ,
    \new_[5673]_ , \new_[5677]_ , \new_[5678]_ , \new_[5682]_ ,
    \new_[5683]_ , \new_[5684]_ , \new_[5688]_ , \new_[5689]_ ,
    \new_[5693]_ , \new_[5694]_ , \new_[5695]_ , \new_[5699]_ ,
    \new_[5700]_ , \new_[5704]_ , \new_[5705]_ , \new_[5706]_ ,
    \new_[5710]_ , \new_[5711]_ , \new_[5715]_ , \new_[5716]_ ,
    \new_[5717]_ , \new_[5721]_ , \new_[5722]_ , \new_[5726]_ ,
    \new_[5727]_ , \new_[5728]_ , \new_[5732]_ , \new_[5733]_ ,
    \new_[5737]_ , \new_[5738]_ , \new_[5739]_ , \new_[5743]_ ,
    \new_[5744]_ , \new_[5748]_ , \new_[5749]_ , \new_[5750]_ ,
    \new_[5754]_ , \new_[5755]_ , \new_[5759]_ , \new_[5760]_ ,
    \new_[5761]_ , \new_[5765]_ , \new_[5766]_ , \new_[5770]_ ,
    \new_[5771]_ , \new_[5772]_ , \new_[5776]_ , \new_[5777]_ ,
    \new_[5781]_ , \new_[5782]_ , \new_[5783]_ , \new_[5787]_ ,
    \new_[5788]_ , \new_[5792]_ , \new_[5793]_ , \new_[5794]_ ,
    \new_[5798]_ , \new_[5799]_ , \new_[5803]_ , \new_[5804]_ ,
    \new_[5805]_ , \new_[5809]_ , \new_[5810]_ , \new_[5814]_ ,
    \new_[5815]_ , \new_[5816]_ , \new_[5820]_ , \new_[5821]_ ,
    \new_[5825]_ , \new_[5826]_ , \new_[5827]_ , \new_[5831]_ ,
    \new_[5832]_ , \new_[5836]_ , \new_[5837]_ , \new_[5838]_ ,
    \new_[5842]_ , \new_[5843]_ , \new_[5847]_ , \new_[5848]_ ,
    \new_[5849]_ , \new_[5853]_ , \new_[5854]_ , \new_[5858]_ ,
    \new_[5859]_ , \new_[5860]_ , \new_[5864]_ , \new_[5865]_ ,
    \new_[5869]_ , \new_[5870]_ , \new_[5871]_ , \new_[5875]_ ,
    \new_[5876]_ , \new_[5880]_ , \new_[5881]_ , \new_[5882]_ ,
    \new_[5886]_ , \new_[5887]_ , \new_[5891]_ , \new_[5892]_ ,
    \new_[5893]_ , \new_[5897]_ , \new_[5898]_ , \new_[5902]_ ,
    \new_[5903]_ , \new_[5904]_ , \new_[5908]_ , \new_[5909]_ ,
    \new_[5913]_ , \new_[5914]_ , \new_[5915]_ , \new_[5919]_ ,
    \new_[5920]_ , \new_[5924]_ , \new_[5925]_ , \new_[5926]_ ,
    \new_[5930]_ , \new_[5931]_ , \new_[5935]_ , \new_[5936]_ ,
    \new_[5937]_ , \new_[5941]_ , \new_[5942]_ , \new_[5946]_ ,
    \new_[5947]_ , \new_[5948]_ , \new_[5952]_ , \new_[5953]_ ,
    \new_[5957]_ , \new_[5958]_ , \new_[5959]_ , \new_[5963]_ ,
    \new_[5964]_ , \new_[5968]_ , \new_[5969]_ , \new_[5970]_ ,
    \new_[5974]_ , \new_[5975]_ , \new_[5979]_ , \new_[5980]_ ,
    \new_[5981]_ , \new_[5985]_ , \new_[5986]_ , \new_[5990]_ ,
    \new_[5991]_ , \new_[5992]_ , \new_[5996]_ , \new_[5997]_ ,
    \new_[6001]_ , \new_[6002]_ , \new_[6003]_ , \new_[6007]_ ,
    \new_[6008]_ , \new_[6012]_ , \new_[6013]_ , \new_[6014]_ ,
    \new_[6018]_ , \new_[6019]_ , \new_[6023]_ , \new_[6024]_ ,
    \new_[6025]_ , \new_[6029]_ , \new_[6030]_ , \new_[6034]_ ,
    \new_[6035]_ , \new_[6036]_ , \new_[6040]_ , \new_[6041]_ ,
    \new_[6045]_ , \new_[6046]_ , \new_[6047]_ , \new_[6051]_ ,
    \new_[6052]_ , \new_[6056]_ , \new_[6057]_ , \new_[6058]_ ,
    \new_[6062]_ , \new_[6063]_ , \new_[6067]_ , \new_[6068]_ ,
    \new_[6069]_ , \new_[6073]_ , \new_[6074]_ , \new_[6078]_ ,
    \new_[6079]_ , \new_[6080]_ , \new_[6084]_ , \new_[6085]_ ,
    \new_[6089]_ , \new_[6090]_ , \new_[6091]_ , \new_[6095]_ ,
    \new_[6096]_ , \new_[6100]_ , \new_[6101]_ , \new_[6102]_ ,
    \new_[6106]_ , \new_[6107]_ , \new_[6111]_ , \new_[6112]_ ,
    \new_[6113]_ , \new_[6117]_ , \new_[6118]_ , \new_[6122]_ ,
    \new_[6123]_ , \new_[6124]_ , \new_[6128]_ , \new_[6129]_ ,
    \new_[6133]_ , \new_[6134]_ , \new_[6135]_ , \new_[6139]_ ,
    \new_[6140]_ , \new_[6144]_ , \new_[6145]_ , \new_[6146]_ ,
    \new_[6150]_ , \new_[6151]_ , \new_[6155]_ , \new_[6156]_ ,
    \new_[6157]_ , \new_[6161]_ , \new_[6162]_ , \new_[6166]_ ,
    \new_[6167]_ , \new_[6168]_ , \new_[6172]_ , \new_[6173]_ ,
    \new_[6177]_ , \new_[6178]_ , \new_[6179]_ , \new_[6183]_ ,
    \new_[6184]_ , \new_[6188]_ , \new_[6189]_ , \new_[6190]_ ,
    \new_[6194]_ , \new_[6195]_ , \new_[6199]_ , \new_[6200]_ ,
    \new_[6201]_ , \new_[6205]_ , \new_[6206]_ , \new_[6210]_ ,
    \new_[6211]_ , \new_[6212]_ , \new_[6216]_ , \new_[6217]_ ,
    \new_[6221]_ , \new_[6222]_ , \new_[6223]_ , \new_[6227]_ ,
    \new_[6228]_ , \new_[6232]_ , \new_[6233]_ , \new_[6234]_ ,
    \new_[6238]_ , \new_[6239]_ , \new_[6243]_ , \new_[6244]_ ,
    \new_[6245]_ , \new_[6249]_ , \new_[6250]_ , \new_[6254]_ ,
    \new_[6255]_ , \new_[6256]_ , \new_[6260]_ , \new_[6261]_ ,
    \new_[6265]_ , \new_[6266]_ , \new_[6267]_ , \new_[6271]_ ,
    \new_[6272]_ , \new_[6276]_ , \new_[6277]_ , \new_[6278]_ ,
    \new_[6282]_ , \new_[6283]_ , \new_[6287]_ , \new_[6288]_ ,
    \new_[6289]_ , \new_[6293]_ , \new_[6294]_ , \new_[6298]_ ,
    \new_[6299]_ , \new_[6300]_ , \new_[6304]_ , \new_[6305]_ ,
    \new_[6309]_ , \new_[6310]_ , \new_[6311]_ , \new_[6315]_ ,
    \new_[6316]_ , \new_[6320]_ , \new_[6321]_ , \new_[6322]_ ,
    \new_[6326]_ , \new_[6327]_ , \new_[6331]_ , \new_[6332]_ ,
    \new_[6333]_ , \new_[6337]_ , \new_[6338]_ , \new_[6342]_ ,
    \new_[6343]_ , \new_[6344]_ , \new_[6348]_ , \new_[6349]_ ,
    \new_[6353]_ , \new_[6354]_ , \new_[6355]_ , \new_[6359]_ ,
    \new_[6360]_ , \new_[6364]_ , \new_[6365]_ , \new_[6366]_ ,
    \new_[6370]_ , \new_[6371]_ , \new_[6375]_ , \new_[6376]_ ,
    \new_[6377]_ , \new_[6381]_ , \new_[6382]_ , \new_[6386]_ ,
    \new_[6387]_ , \new_[6388]_ , \new_[6392]_ , \new_[6393]_ ,
    \new_[6397]_ , \new_[6398]_ , \new_[6399]_ , \new_[6403]_ ,
    \new_[6404]_ , \new_[6408]_ , \new_[6409]_ , \new_[6410]_ ,
    \new_[6414]_ , \new_[6415]_ , \new_[6419]_ , \new_[6420]_ ,
    \new_[6421]_ , \new_[6425]_ , \new_[6426]_ , \new_[6430]_ ,
    \new_[6431]_ , \new_[6432]_ , \new_[6436]_ , \new_[6437]_ ,
    \new_[6441]_ , \new_[6442]_ , \new_[6443]_ , \new_[6447]_ ,
    \new_[6448]_ , \new_[6452]_ , \new_[6453]_ , \new_[6454]_ ,
    \new_[6458]_ , \new_[6459]_ , \new_[6463]_ , \new_[6464]_ ,
    \new_[6465]_ , \new_[6469]_ , \new_[6470]_ , \new_[6474]_ ,
    \new_[6475]_ , \new_[6476]_ , \new_[6480]_ , \new_[6481]_ ,
    \new_[6485]_ , \new_[6486]_ , \new_[6487]_ , \new_[6491]_ ,
    \new_[6492]_ , \new_[6496]_ , \new_[6497]_ , \new_[6498]_ ,
    \new_[6502]_ , \new_[6503]_ , \new_[6507]_ , \new_[6508]_ ,
    \new_[6509]_ , \new_[6513]_ , \new_[6514]_ , \new_[6518]_ ,
    \new_[6519]_ , \new_[6520]_ , \new_[6524]_ , \new_[6525]_ ,
    \new_[6529]_ , \new_[6530]_ , \new_[6531]_ , \new_[6535]_ ,
    \new_[6536]_ , \new_[6540]_ , \new_[6541]_ , \new_[6542]_ ,
    \new_[6546]_ , \new_[6547]_ , \new_[6551]_ , \new_[6552]_ ,
    \new_[6553]_ , \new_[6557]_ , \new_[6558]_ , \new_[6562]_ ,
    \new_[6563]_ , \new_[6564]_ , \new_[6568]_ , \new_[6569]_ ,
    \new_[6573]_ , \new_[6574]_ , \new_[6575]_ , \new_[6579]_ ,
    \new_[6580]_ , \new_[6584]_ , \new_[6585]_ , \new_[6586]_ ,
    \new_[6590]_ , \new_[6591]_ , \new_[6595]_ , \new_[6596]_ ,
    \new_[6597]_ , \new_[6601]_ , \new_[6602]_ , \new_[6606]_ ,
    \new_[6607]_ , \new_[6608]_ , \new_[6612]_ , \new_[6613]_ ,
    \new_[6617]_ , \new_[6618]_ , \new_[6619]_ , \new_[6623]_ ,
    \new_[6624]_ , \new_[6628]_ , \new_[6629]_ , \new_[6630]_ ,
    \new_[6634]_ , \new_[6635]_ , \new_[6639]_ , \new_[6640]_ ,
    \new_[6641]_ , \new_[6645]_ , \new_[6646]_ , \new_[6650]_ ,
    \new_[6651]_ , \new_[6652]_ , \new_[6656]_ , \new_[6657]_ ,
    \new_[6661]_ , \new_[6662]_ , \new_[6663]_ , \new_[6667]_ ,
    \new_[6668]_ , \new_[6672]_ , \new_[6673]_ , \new_[6674]_ ;
  assign A41 = \new_[1042]_  | \new_[695]_ ;
  assign \new_[1]_  = \new_[6674]_  & \new_[6663]_ ;
  assign \new_[2]_  = \new_[6652]_  & \new_[6641]_ ;
  assign \new_[3]_  = \new_[6630]_  & \new_[6619]_ ;
  assign \new_[4]_  = \new_[6608]_  & \new_[6597]_ ;
  assign \new_[5]_  = \new_[6586]_  & \new_[6575]_ ;
  assign \new_[6]_  = \new_[6564]_  & \new_[6553]_ ;
  assign \new_[7]_  = \new_[6542]_  & \new_[6531]_ ;
  assign \new_[8]_  = \new_[6520]_  & \new_[6509]_ ;
  assign \new_[9]_  = \new_[6498]_  & \new_[6487]_ ;
  assign \new_[10]_  = \new_[6476]_  & \new_[6465]_ ;
  assign \new_[11]_  = \new_[6454]_  & \new_[6443]_ ;
  assign \new_[12]_  = \new_[6432]_  & \new_[6421]_ ;
  assign \new_[13]_  = \new_[6410]_  & \new_[6399]_ ;
  assign \new_[14]_  = \new_[6388]_  & \new_[6377]_ ;
  assign \new_[15]_  = \new_[6366]_  & \new_[6355]_ ;
  assign \new_[16]_  = \new_[6344]_  & \new_[6333]_ ;
  assign \new_[17]_  = \new_[6322]_  & \new_[6311]_ ;
  assign \new_[18]_  = \new_[6300]_  & \new_[6289]_ ;
  assign \new_[19]_  = \new_[6278]_  & \new_[6267]_ ;
  assign \new_[20]_  = \new_[6256]_  & \new_[6245]_ ;
  assign \new_[21]_  = \new_[6234]_  & \new_[6223]_ ;
  assign \new_[22]_  = \new_[6212]_  & \new_[6201]_ ;
  assign \new_[23]_  = \new_[6190]_  & \new_[6179]_ ;
  assign \new_[24]_  = \new_[6168]_  & \new_[6157]_ ;
  assign \new_[25]_  = \new_[6146]_  & \new_[6135]_ ;
  assign \new_[26]_  = \new_[6124]_  & \new_[6113]_ ;
  assign \new_[27]_  = \new_[6102]_  & \new_[6091]_ ;
  assign \new_[28]_  = \new_[6080]_  & \new_[6069]_ ;
  assign \new_[29]_  = \new_[6058]_  & \new_[6047]_ ;
  assign \new_[30]_  = \new_[6036]_  & \new_[6025]_ ;
  assign \new_[31]_  = \new_[6014]_  & \new_[6003]_ ;
  assign \new_[32]_  = \new_[5992]_  & \new_[5981]_ ;
  assign \new_[33]_  = \new_[5970]_  & \new_[5959]_ ;
  assign \new_[34]_  = \new_[5948]_  & \new_[5937]_ ;
  assign \new_[35]_  = \new_[5926]_  & \new_[5915]_ ;
  assign \new_[36]_  = \new_[5904]_  & \new_[5893]_ ;
  assign \new_[37]_  = \new_[5882]_  & \new_[5871]_ ;
  assign \new_[38]_  = \new_[5860]_  & \new_[5849]_ ;
  assign \new_[39]_  = \new_[5838]_  & \new_[5827]_ ;
  assign \new_[40]_  = \new_[5816]_  & \new_[5805]_ ;
  assign \new_[41]_  = \new_[5794]_  & \new_[5783]_ ;
  assign \new_[42]_  = \new_[5772]_  & \new_[5761]_ ;
  assign \new_[43]_  = \new_[5750]_  & \new_[5739]_ ;
  assign \new_[44]_  = \new_[5728]_  & \new_[5717]_ ;
  assign \new_[45]_  = \new_[5706]_  & \new_[5695]_ ;
  assign \new_[46]_  = \new_[5684]_  & \new_[5673]_ ;
  assign \new_[47]_  = \new_[5662]_  & \new_[5651]_ ;
  assign \new_[48]_  = \new_[5640]_  & \new_[5629]_ ;
  assign \new_[49]_  = \new_[5618]_  & \new_[5607]_ ;
  assign \new_[50]_  = \new_[5598]_  & \new_[5587]_ ;
  assign \new_[51]_  = \new_[5578]_  & \new_[5567]_ ;
  assign \new_[52]_  = \new_[5558]_  & \new_[5547]_ ;
  assign \new_[53]_  = \new_[5538]_  & \new_[5527]_ ;
  assign \new_[54]_  = \new_[5518]_  & \new_[5507]_ ;
  assign \new_[55]_  = \new_[5498]_  & \new_[5487]_ ;
  assign \new_[56]_  = \new_[5478]_  & \new_[5467]_ ;
  assign \new_[57]_  = \new_[5458]_  & \new_[5447]_ ;
  assign \new_[58]_  = \new_[5438]_  & \new_[5427]_ ;
  assign \new_[59]_  = \new_[5418]_  & \new_[5407]_ ;
  assign \new_[60]_  = \new_[5398]_  & \new_[5387]_ ;
  assign \new_[61]_  = \new_[5378]_  & \new_[5367]_ ;
  assign \new_[62]_  = \new_[5358]_  & \new_[5347]_ ;
  assign \new_[63]_  = \new_[5338]_  & \new_[5327]_ ;
  assign \new_[64]_  = \new_[5318]_  & \new_[5307]_ ;
  assign \new_[65]_  = \new_[5298]_  & \new_[5287]_ ;
  assign \new_[66]_  = \new_[5278]_  & \new_[5267]_ ;
  assign \new_[67]_  = \new_[5258]_  & \new_[5247]_ ;
  assign \new_[68]_  = \new_[5238]_  & \new_[5227]_ ;
  assign \new_[69]_  = \new_[5218]_  & \new_[5207]_ ;
  assign \new_[70]_  = \new_[5198]_  & \new_[5187]_ ;
  assign \new_[71]_  = \new_[5178]_  & \new_[5167]_ ;
  assign \new_[72]_  = \new_[5158]_  & \new_[5147]_ ;
  assign \new_[73]_  = \new_[5138]_  & \new_[5127]_ ;
  assign \new_[74]_  = \new_[5118]_  & \new_[5107]_ ;
  assign \new_[75]_  = \new_[5098]_  & \new_[5087]_ ;
  assign \new_[76]_  = \new_[5078]_  & \new_[5067]_ ;
  assign \new_[77]_  = \new_[5058]_  & \new_[5047]_ ;
  assign \new_[78]_  = \new_[5038]_  & \new_[5027]_ ;
  assign \new_[79]_  = \new_[5018]_  & \new_[5007]_ ;
  assign \new_[80]_  = \new_[4998]_  & \new_[4987]_ ;
  assign \new_[81]_  = \new_[4978]_  & \new_[4969]_ ;
  assign \new_[82]_  = \new_[4960]_  & \new_[4951]_ ;
  assign \new_[83]_  = \new_[4942]_  & \new_[4933]_ ;
  assign \new_[84]_  = \new_[4924]_  & \new_[4915]_ ;
  assign \new_[85]_  = \new_[4906]_  & \new_[4897]_ ;
  assign \new_[86]_  = \new_[4888]_  & \new_[4879]_ ;
  assign \new_[87]_  = \new_[4870]_  & \new_[4861]_ ;
  assign \new_[88]_  = \new_[4852]_  & \new_[4843]_ ;
  assign \new_[89]_  = \new_[4834]_  & \new_[4825]_ ;
  assign \new_[90]_  = \new_[4816]_  & \new_[4807]_ ;
  assign \new_[91]_  = \new_[4798]_  & \new_[4789]_ ;
  assign \new_[92]_  = \new_[4780]_  & \new_[4771]_ ;
  assign \new_[93]_  = \new_[4762]_  & \new_[4753]_ ;
  assign \new_[94]_  = \new_[4744]_  & \new_[4735]_ ;
  assign \new_[95]_  = \new_[4726]_  & \new_[4717]_ ;
  assign \new_[96]_  = \new_[4708]_  & \new_[4699]_ ;
  assign \new_[97]_  = \new_[4690]_  & \new_[4681]_ ;
  assign \new_[98]_  = \new_[4672]_  & \new_[4663]_ ;
  assign \new_[99]_  = \new_[4654]_  & \new_[4645]_ ;
  assign \new_[100]_  = \new_[4636]_  & \new_[4627]_ ;
  assign \new_[101]_  = \new_[4618]_  & \new_[4609]_ ;
  assign \new_[102]_  = \new_[4600]_  & \new_[4591]_ ;
  assign \new_[103]_  = \new_[4582]_  & \new_[4573]_ ;
  assign \new_[104]_  = \new_[4564]_  & \new_[4555]_ ;
  assign \new_[105]_  = \new_[4546]_  & \new_[4537]_ ;
  assign \new_[106]_  = \new_[4528]_  & \new_[4519]_ ;
  assign \new_[107]_  = \new_[4510]_  & \new_[4501]_ ;
  assign \new_[108]_  = \new_[4492]_  & \new_[4483]_ ;
  assign \new_[109]_  = \new_[4474]_  & \new_[4465]_ ;
  assign \new_[110]_  = \new_[4456]_  & \new_[4447]_ ;
  assign \new_[111]_  = \new_[4438]_  & \new_[4429]_ ;
  assign \new_[112]_  = \new_[4420]_  & \new_[4411]_ ;
  assign \new_[113]_  = \new_[4402]_  & \new_[4393]_ ;
  assign \new_[114]_  = \new_[4384]_  & \new_[4375]_ ;
  assign \new_[115]_  = \new_[4366]_  & \new_[4357]_ ;
  assign \new_[116]_  = \new_[4348]_  & \new_[4339]_ ;
  assign \new_[117]_  = \new_[4330]_  & \new_[4321]_ ;
  assign \new_[118]_  = \new_[4312]_  & \new_[4303]_ ;
  assign \new_[119]_  = \new_[4294]_  & \new_[4285]_ ;
  assign \new_[120]_  = \new_[4276]_  & \new_[4267]_ ;
  assign \new_[121]_  = \new_[4258]_  & \new_[4249]_ ;
  assign \new_[122]_  = \new_[4240]_  & \new_[4231]_ ;
  assign \new_[123]_  = \new_[4222]_  & \new_[4213]_ ;
  assign \new_[124]_  = \new_[4204]_  & \new_[4195]_ ;
  assign \new_[125]_  = \new_[4186]_  & \new_[4177]_ ;
  assign \new_[126]_  = \new_[4168]_  & \new_[4159]_ ;
  assign \new_[127]_  = \new_[4150]_  & \new_[4141]_ ;
  assign \new_[128]_  = \new_[4132]_  & \new_[4123]_ ;
  assign \new_[129]_  = \new_[4114]_  & \new_[4105]_ ;
  assign \new_[130]_  = \new_[4096]_  & \new_[4087]_ ;
  assign \new_[131]_  = \new_[4078]_  & \new_[4069]_ ;
  assign \new_[132]_  = \new_[4060]_  & \new_[4051]_ ;
  assign \new_[133]_  = \new_[4042]_  & \new_[4033]_ ;
  assign \new_[134]_  = \new_[4024]_  & \new_[4015]_ ;
  assign \new_[135]_  = \new_[4006]_  & \new_[3997]_ ;
  assign \new_[136]_  = \new_[3988]_  & \new_[3979]_ ;
  assign \new_[137]_  = \new_[3970]_  & \new_[3961]_ ;
  assign \new_[138]_  = \new_[3952]_  & \new_[3943]_ ;
  assign \new_[139]_  = \new_[3934]_  & \new_[3925]_ ;
  assign \new_[140]_  = \new_[3916]_  & \new_[3907]_ ;
  assign \new_[141]_  = \new_[3898]_  & \new_[3889]_ ;
  assign \new_[142]_  = \new_[3880]_  & \new_[3871]_ ;
  assign \new_[143]_  = \new_[3862]_  & \new_[3853]_ ;
  assign \new_[144]_  = \new_[3844]_  & \new_[3835]_ ;
  assign \new_[145]_  = \new_[3826]_  & \new_[3817]_ ;
  assign \new_[146]_  = \new_[3808]_  & \new_[3799]_ ;
  assign \new_[147]_  = \new_[3790]_  & \new_[3781]_ ;
  assign \new_[148]_  = \new_[3772]_  & \new_[3763]_ ;
  assign \new_[149]_  = \new_[3754]_  & \new_[3745]_ ;
  assign \new_[150]_  = \new_[3736]_  & \new_[3727]_ ;
  assign \new_[151]_  = \new_[3718]_  & \new_[3709]_ ;
  assign \new_[152]_  = \new_[3700]_  & \new_[3691]_ ;
  assign \new_[153]_  = \new_[3682]_  & \new_[3673]_ ;
  assign \new_[154]_  = \new_[3664]_  & \new_[3655]_ ;
  assign \new_[155]_  = \new_[3646]_  & \new_[3637]_ ;
  assign \new_[156]_  = \new_[3628]_  & \new_[3619]_ ;
  assign \new_[157]_  = \new_[3610]_  & \new_[3601]_ ;
  assign \new_[158]_  = \new_[3592]_  & \new_[3583]_ ;
  assign \new_[159]_  = \new_[3574]_  & \new_[3565]_ ;
  assign \new_[160]_  = \new_[3556]_  & \new_[3547]_ ;
  assign \new_[161]_  = \new_[3538]_  & \new_[3529]_ ;
  assign \new_[162]_  = \new_[3520]_  & \new_[3511]_ ;
  assign \new_[163]_  = \new_[3502]_  & \new_[3493]_ ;
  assign \new_[164]_  = \new_[3484]_  & \new_[3475]_ ;
  assign \new_[165]_  = \new_[3466]_  & \new_[3457]_ ;
  assign \new_[166]_  = \new_[3448]_  & \new_[3439]_ ;
  assign \new_[167]_  = \new_[3430]_  & \new_[3421]_ ;
  assign \new_[168]_  = \new_[3412]_  & \new_[3403]_ ;
  assign \new_[169]_  = \new_[3394]_  & \new_[3385]_ ;
  assign \new_[170]_  = \new_[3376]_  & \new_[3367]_ ;
  assign \new_[171]_  = \new_[3358]_  & \new_[3349]_ ;
  assign \new_[172]_  = \new_[3340]_  & \new_[3331]_ ;
  assign \new_[173]_  = \new_[3322]_  & \new_[3313]_ ;
  assign \new_[174]_  = \new_[3304]_  & \new_[3295]_ ;
  assign \new_[175]_  = \new_[3286]_  & \new_[3277]_ ;
  assign \new_[176]_  = \new_[3268]_  & \new_[3259]_ ;
  assign \new_[177]_  = \new_[3250]_  & \new_[3241]_ ;
  assign \new_[178]_  = \new_[3234]_  & \new_[3225]_ ;
  assign \new_[179]_  = \new_[3218]_  & \new_[3209]_ ;
  assign \new_[180]_  = \new_[3202]_  & \new_[3193]_ ;
  assign \new_[181]_  = \new_[3186]_  & \new_[3177]_ ;
  assign \new_[182]_  = \new_[3170]_  & \new_[3161]_ ;
  assign \new_[183]_  = \new_[3154]_  & \new_[3145]_ ;
  assign \new_[184]_  = \new_[3138]_  & \new_[3129]_ ;
  assign \new_[185]_  = \new_[3122]_  & \new_[3113]_ ;
  assign \new_[186]_  = \new_[3106]_  & \new_[3097]_ ;
  assign \new_[187]_  = \new_[3090]_  & \new_[3081]_ ;
  assign \new_[188]_  = \new_[3074]_  & \new_[3065]_ ;
  assign \new_[189]_  = \new_[3058]_  & \new_[3049]_ ;
  assign \new_[190]_  = \new_[3042]_  & \new_[3033]_ ;
  assign \new_[191]_  = \new_[3026]_  & \new_[3017]_ ;
  assign \new_[192]_  = \new_[3010]_  & \new_[3001]_ ;
  assign \new_[193]_  = \new_[2994]_  & \new_[2985]_ ;
  assign \new_[194]_  = \new_[2978]_  & \new_[2969]_ ;
  assign \new_[195]_  = \new_[2962]_  & \new_[2953]_ ;
  assign \new_[196]_  = \new_[2946]_  & \new_[2937]_ ;
  assign \new_[197]_  = \new_[2930]_  & \new_[2921]_ ;
  assign \new_[198]_  = \new_[2914]_  & \new_[2905]_ ;
  assign \new_[199]_  = \new_[2898]_  & \new_[2889]_ ;
  assign \new_[200]_  = \new_[2882]_  & \new_[2873]_ ;
  assign \new_[201]_  = \new_[2866]_  & \new_[2857]_ ;
  assign \new_[202]_  = \new_[2850]_  & \new_[2841]_ ;
  assign \new_[203]_  = \new_[2834]_  & \new_[2825]_ ;
  assign \new_[204]_  = \new_[2818]_  & \new_[2809]_ ;
  assign \new_[205]_  = \new_[2802]_  & \new_[2793]_ ;
  assign \new_[206]_  = \new_[2786]_  & \new_[2777]_ ;
  assign \new_[207]_  = \new_[2770]_  & \new_[2761]_ ;
  assign \new_[208]_  = \new_[2754]_  & \new_[2745]_ ;
  assign \new_[209]_  = \new_[2738]_  & \new_[2731]_ ;
  assign \new_[210]_  = \new_[2724]_  & \new_[2717]_ ;
  assign \new_[211]_  = \new_[2710]_  & \new_[2703]_ ;
  assign \new_[212]_  = \new_[2696]_  & \new_[2689]_ ;
  assign \new_[213]_  = \new_[2682]_  & \new_[2675]_ ;
  assign \new_[214]_  = \new_[2668]_  & \new_[2661]_ ;
  assign \new_[215]_  = \new_[2654]_  & \new_[2647]_ ;
  assign \new_[216]_  = \new_[2640]_  & \new_[2633]_ ;
  assign \new_[217]_  = \new_[2626]_  & \new_[2619]_ ;
  assign \new_[218]_  = \new_[2612]_  & \new_[2605]_ ;
  assign \new_[219]_  = \new_[2598]_  & \new_[2591]_ ;
  assign \new_[220]_  = \new_[2584]_  & \new_[2577]_ ;
  assign \new_[221]_  = \new_[2570]_  & \new_[2563]_ ;
  assign \new_[222]_  = \new_[2556]_  & \new_[2549]_ ;
  assign \new_[223]_  = \new_[2542]_  & \new_[2535]_ ;
  assign \new_[224]_  = \new_[2528]_  & \new_[2521]_ ;
  assign \new_[225]_  = \new_[2514]_  & \new_[2507]_ ;
  assign \new_[226]_  = \new_[2500]_  & \new_[2493]_ ;
  assign \new_[227]_  = \new_[2486]_  & \new_[2479]_ ;
  assign \new_[228]_  = \new_[2472]_  & \new_[2465]_ ;
  assign \new_[229]_  = \new_[2458]_  & \new_[2451]_ ;
  assign \new_[230]_  = \new_[2444]_  & \new_[2437]_ ;
  assign \new_[231]_  = \new_[2430]_  & \new_[2423]_ ;
  assign \new_[232]_  = \new_[2416]_  & \new_[2409]_ ;
  assign \new_[233]_  = \new_[2402]_  & \new_[2395]_ ;
  assign \new_[234]_  = \new_[2388]_  & \new_[2381]_ ;
  assign \new_[235]_  = \new_[2374]_  & \new_[2367]_ ;
  assign \new_[236]_  = \new_[2360]_  & \new_[2353]_ ;
  assign \new_[237]_  = \new_[2346]_  & \new_[2339]_ ;
  assign \new_[238]_  = \new_[2332]_  & \new_[2325]_ ;
  assign \new_[239]_  = \new_[2318]_  & \new_[2311]_ ;
  assign \new_[240]_  = \new_[2304]_  & \new_[2297]_ ;
  assign \new_[241]_  = \new_[2290]_  & \new_[2283]_ ;
  assign \new_[242]_  = \new_[2276]_  & \new_[2269]_ ;
  assign \new_[243]_  = \new_[2262]_  & \new_[2255]_ ;
  assign \new_[244]_  = \new_[2248]_  & \new_[2241]_ ;
  assign \new_[245]_  = \new_[2234]_  & \new_[2227]_ ;
  assign \new_[246]_  = \new_[2220]_  & \new_[2213]_ ;
  assign \new_[247]_  = \new_[2206]_  & \new_[2199]_ ;
  assign \new_[248]_  = \new_[2192]_  & \new_[2185]_ ;
  assign \new_[249]_  = \new_[2178]_  & \new_[2171]_ ;
  assign \new_[250]_  = \new_[2164]_  & \new_[2157]_ ;
  assign \new_[251]_  = \new_[2150]_  & \new_[2143]_ ;
  assign \new_[252]_  = \new_[2136]_  & \new_[2129]_ ;
  assign \new_[253]_  = \new_[2122]_  & \new_[2115]_ ;
  assign \new_[254]_  = \new_[2108]_  & \new_[2101]_ ;
  assign \new_[255]_  = \new_[2094]_  & \new_[2087]_ ;
  assign \new_[256]_  = \new_[2080]_  & \new_[2073]_ ;
  assign \new_[257]_  = \new_[2066]_  & \new_[2059]_ ;
  assign \new_[258]_  = \new_[2052]_  & \new_[2045]_ ;
  assign \new_[259]_  = \new_[2038]_  & \new_[2031]_ ;
  assign \new_[260]_  = \new_[2024]_  & \new_[2017]_ ;
  assign \new_[261]_  = \new_[2010]_  & \new_[2003]_ ;
  assign \new_[262]_  = \new_[1996]_  & \new_[1989]_ ;
  assign \new_[263]_  = \new_[1982]_  & \new_[1975]_ ;
  assign \new_[264]_  = \new_[1968]_  & \new_[1961]_ ;
  assign \new_[265]_  = \new_[1954]_  & \new_[1947]_ ;
  assign \new_[266]_  = \new_[1940]_  & \new_[1933]_ ;
  assign \new_[267]_  = \new_[1926]_  & \new_[1919]_ ;
  assign \new_[268]_  = \new_[1912]_  & \new_[1905]_ ;
  assign \new_[269]_  = \new_[1898]_  & \new_[1891]_ ;
  assign \new_[270]_  = \new_[1884]_  & \new_[1877]_ ;
  assign \new_[271]_  = \new_[1870]_  & \new_[1863]_ ;
  assign \new_[272]_  = \new_[1856]_  & \new_[1849]_ ;
  assign \new_[273]_  = \new_[1842]_  & \new_[1835]_ ;
  assign \new_[274]_  = \new_[1828]_  & \new_[1821]_ ;
  assign \new_[275]_  = \new_[1814]_  & \new_[1807]_ ;
  assign \new_[276]_  = \new_[1800]_  & \new_[1793]_ ;
  assign \new_[277]_  = \new_[1786]_  & \new_[1779]_ ;
  assign \new_[278]_  = \new_[1772]_  & \new_[1765]_ ;
  assign \new_[279]_  = \new_[1758]_  & \new_[1751]_ ;
  assign \new_[280]_  = \new_[1744]_  & \new_[1737]_ ;
  assign \new_[281]_  = \new_[1730]_  & \new_[1723]_ ;
  assign \new_[282]_  = \new_[1716]_  & \new_[1709]_ ;
  assign \new_[283]_  = \new_[1702]_  & \new_[1695]_ ;
  assign \new_[284]_  = \new_[1688]_  & \new_[1681]_ ;
  assign \new_[285]_  = \new_[1674]_  & \new_[1667]_ ;
  assign \new_[286]_  = \new_[1660]_  & \new_[1653]_ ;
  assign \new_[287]_  = \new_[1646]_  & \new_[1639]_ ;
  assign \new_[288]_  = \new_[1632]_  & \new_[1625]_ ;
  assign \new_[289]_  = \new_[1618]_  & \new_[1611]_ ;
  assign \new_[290]_  = \new_[1604]_  & \new_[1597]_ ;
  assign \new_[291]_  = \new_[1590]_  & \new_[1583]_ ;
  assign \new_[292]_  = \new_[1576]_  & \new_[1569]_ ;
  assign \new_[293]_  = \new_[1562]_  & \new_[1555]_ ;
  assign \new_[294]_  = \new_[1550]_  & \new_[1543]_ ;
  assign \new_[295]_  = \new_[1538]_  & \new_[1531]_ ;
  assign \new_[296]_  = \new_[1526]_  & \new_[1519]_ ;
  assign \new_[297]_  = \new_[1514]_  & \new_[1507]_ ;
  assign \new_[298]_  = \new_[1502]_  & \new_[1495]_ ;
  assign \new_[299]_  = \new_[1490]_  & \new_[1483]_ ;
  assign \new_[300]_  = \new_[1478]_  & \new_[1471]_ ;
  assign \new_[301]_  = \new_[1466]_  & \new_[1461]_ ;
  assign \new_[302]_  = \new_[1456]_  & \new_[1451]_ ;
  assign \new_[303]_  = \new_[1446]_  & \new_[1441]_ ;
  assign \new_[304]_  = \new_[1436]_  & \new_[1431]_ ;
  assign \new_[305]_  = \new_[1426]_  & \new_[1421]_ ;
  assign \new_[306]_  = \new_[1416]_  & \new_[1411]_ ;
  assign \new_[307]_  = \new_[1406]_  & \new_[1401]_ ;
  assign \new_[308]_  = \new_[1396]_  & \new_[1391]_ ;
  assign \new_[309]_  = \new_[1386]_  & \new_[1381]_ ;
  assign \new_[310]_  = \new_[1376]_  & \new_[1371]_ ;
  assign \new_[311]_  = \new_[1366]_  & \new_[1361]_ ;
  assign \new_[312]_  = \new_[1356]_  & \new_[1351]_ ;
  assign \new_[313]_  = \new_[1346]_  & \new_[1341]_ ;
  assign \new_[314]_  = \new_[1336]_  & \new_[1331]_ ;
  assign \new_[315]_  = \new_[1326]_  & \new_[1321]_ ;
  assign \new_[316]_  = \new_[1316]_  & \new_[1311]_ ;
  assign \new_[317]_  = \new_[1306]_  & \new_[1301]_ ;
  assign \new_[318]_  = \new_[1296]_  & \new_[1291]_ ;
  assign \new_[319]_  = \new_[1286]_  & \new_[1281]_ ;
  assign \new_[320]_  = \new_[1276]_  & \new_[1271]_ ;
  assign \new_[321]_  = \new_[1266]_  & \new_[1261]_ ;
  assign \new_[322]_  = \new_[1256]_  & \new_[1251]_ ;
  assign \new_[323]_  = \new_[1246]_  & \new_[1241]_ ;
  assign \new_[324]_  = \new_[1236]_  & \new_[1231]_ ;
  assign \new_[325]_  = \new_[1226]_  & \new_[1221]_ ;
  assign \new_[326]_  = \new_[1216]_  & \new_[1211]_ ;
  assign \new_[327]_  = \new_[1206]_  & \new_[1201]_ ;
  assign \new_[328]_  = \new_[1196]_  & \new_[1191]_ ;
  assign \new_[329]_  = \new_[1186]_  & \new_[1181]_ ;
  assign \new_[330]_  = \new_[1176]_  & \new_[1171]_ ;
  assign \new_[331]_  = \new_[1166]_  & \new_[1161]_ ;
  assign \new_[332]_  = \new_[1156]_  & \new_[1151]_ ;
  assign \new_[333]_  = \new_[1146]_  & \new_[1141]_ ;
  assign \new_[334]_  = \new_[1136]_  & \new_[1131]_ ;
  assign \new_[335]_  = \new_[1126]_  & \new_[1121]_ ;
  assign \new_[336]_  = \new_[1116]_  & \new_[1111]_ ;
  assign \new_[337]_  = \new_[1106]_  & \new_[1103]_ ;
  assign \new_[338]_  = \new_[1100]_  & \new_[1097]_ ;
  assign \new_[339]_  = \new_[1094]_  & \new_[1091]_ ;
  assign \new_[340]_  = \new_[1088]_  & \new_[1085]_ ;
  assign \new_[341]_  = \new_[1082]_  & \new_[1079]_ ;
  assign \new_[342]_  = \new_[1076]_  & \new_[1073]_ ;
  assign \new_[343]_  = \new_[1070]_  & \new_[1067]_ ;
  assign \new_[344]_  = \new_[1064]_  & \new_[1061]_ ;
  assign \new_[345]_  = \new_[1058]_  & \new_[1055]_ ;
  assign \new_[346]_  = \new_[1052]_  & \new_[1049]_ ;
  assign \new_[347]_  = A267 & A266;
  assign \new_[348]_  = A267 & A265;
  assign \new_[351]_  = \new_[347]_  | \new_[348]_ ;
  assign \new_[355]_  = \new_[344]_  | \new_[345]_ ;
  assign \new_[356]_  = \new_[346]_  | \new_[355]_ ;
  assign \new_[357]_  = \new_[356]_  | \new_[351]_ ;
  assign \new_[360]_  = \new_[342]_  | \new_[343]_ ;
  assign \new_[364]_  = \new_[339]_  | \new_[340]_ ;
  assign \new_[365]_  = \new_[341]_  | \new_[364]_ ;
  assign \new_[366]_  = \new_[365]_  | \new_[360]_ ;
  assign \new_[367]_  = \new_[366]_  | \new_[357]_ ;
  assign \new_[370]_  = \new_[337]_  | \new_[338]_ ;
  assign \new_[374]_  = \new_[334]_  | \new_[335]_ ;
  assign \new_[375]_  = \new_[336]_  | \new_[374]_ ;
  assign \new_[376]_  = \new_[375]_  | \new_[370]_ ;
  assign \new_[380]_  = \new_[331]_  | \new_[332]_ ;
  assign \new_[381]_  = \new_[333]_  | \new_[380]_ ;
  assign \new_[385]_  = \new_[328]_  | \new_[329]_ ;
  assign \new_[386]_  = \new_[330]_  | \new_[385]_ ;
  assign \new_[387]_  = \new_[386]_  | \new_[381]_ ;
  assign \new_[388]_  = \new_[387]_  | \new_[376]_ ;
  assign \new_[389]_  = \new_[388]_  | \new_[367]_ ;
  assign \new_[392]_  = \new_[326]_  | \new_[327]_ ;
  assign \new_[396]_  = \new_[323]_  | \new_[324]_ ;
  assign \new_[397]_  = \new_[325]_  | \new_[396]_ ;
  assign \new_[398]_  = \new_[397]_  | \new_[392]_ ;
  assign \new_[402]_  = \new_[320]_  | \new_[321]_ ;
  assign \new_[403]_  = \new_[322]_  | \new_[402]_ ;
  assign \new_[407]_  = \new_[317]_  | \new_[318]_ ;
  assign \new_[408]_  = \new_[319]_  | \new_[407]_ ;
  assign \new_[409]_  = \new_[408]_  | \new_[403]_ ;
  assign \new_[410]_  = \new_[409]_  | \new_[398]_ ;
  assign \new_[413]_  = \new_[315]_  | \new_[316]_ ;
  assign \new_[417]_  = \new_[312]_  | \new_[313]_ ;
  assign \new_[418]_  = \new_[314]_  | \new_[417]_ ;
  assign \new_[419]_  = \new_[418]_  | \new_[413]_ ;
  assign \new_[423]_  = \new_[309]_  | \new_[310]_ ;
  assign \new_[424]_  = \new_[311]_  | \new_[423]_ ;
  assign \new_[428]_  = \new_[306]_  | \new_[307]_ ;
  assign \new_[429]_  = \new_[308]_  | \new_[428]_ ;
  assign \new_[430]_  = \new_[429]_  | \new_[424]_ ;
  assign \new_[431]_  = \new_[430]_  | \new_[419]_ ;
  assign \new_[432]_  = \new_[431]_  | \new_[410]_ ;
  assign \new_[433]_  = \new_[432]_  | \new_[389]_ ;
  assign \new_[436]_  = \new_[304]_  | \new_[305]_ ;
  assign \new_[440]_  = \new_[301]_  | \new_[302]_ ;
  assign \new_[441]_  = \new_[303]_  | \new_[440]_ ;
  assign \new_[442]_  = \new_[441]_  | \new_[436]_ ;
  assign \new_[446]_  = \new_[298]_  | \new_[299]_ ;
  assign \new_[447]_  = \new_[300]_  | \new_[446]_ ;
  assign \new_[451]_  = \new_[295]_  | \new_[296]_ ;
  assign \new_[452]_  = \new_[297]_  | \new_[451]_ ;
  assign \new_[453]_  = \new_[452]_  | \new_[447]_ ;
  assign \new_[454]_  = \new_[453]_  | \new_[442]_ ;
  assign \new_[457]_  = \new_[293]_  | \new_[294]_ ;
  assign \new_[461]_  = \new_[290]_  | \new_[291]_ ;
  assign \new_[462]_  = \new_[292]_  | \new_[461]_ ;
  assign \new_[463]_  = \new_[462]_  | \new_[457]_ ;
  assign \new_[467]_  = \new_[287]_  | \new_[288]_ ;
  assign \new_[468]_  = \new_[289]_  | \new_[467]_ ;
  assign \new_[472]_  = \new_[284]_  | \new_[285]_ ;
  assign \new_[473]_  = \new_[286]_  | \new_[472]_ ;
  assign \new_[474]_  = \new_[473]_  | \new_[468]_ ;
  assign \new_[475]_  = \new_[474]_  | \new_[463]_ ;
  assign \new_[476]_  = \new_[475]_  | \new_[454]_ ;
  assign \new_[479]_  = \new_[282]_  | \new_[283]_ ;
  assign \new_[483]_  = \new_[279]_  | \new_[280]_ ;
  assign \new_[484]_  = \new_[281]_  | \new_[483]_ ;
  assign \new_[485]_  = \new_[484]_  | \new_[479]_ ;
  assign \new_[489]_  = \new_[276]_  | \new_[277]_ ;
  assign \new_[490]_  = \new_[278]_  | \new_[489]_ ;
  assign \new_[494]_  = \new_[273]_  | \new_[274]_ ;
  assign \new_[495]_  = \new_[275]_  | \new_[494]_ ;
  assign \new_[496]_  = \new_[495]_  | \new_[490]_ ;
  assign \new_[497]_  = \new_[496]_  | \new_[485]_ ;
  assign \new_[500]_  = \new_[271]_  | \new_[272]_ ;
  assign \new_[504]_  = \new_[268]_  | \new_[269]_ ;
  assign \new_[505]_  = \new_[270]_  | \new_[504]_ ;
  assign \new_[506]_  = \new_[505]_  | \new_[500]_ ;
  assign \new_[510]_  = \new_[265]_  | \new_[266]_ ;
  assign \new_[511]_  = \new_[267]_  | \new_[510]_ ;
  assign \new_[515]_  = \new_[262]_  | \new_[263]_ ;
  assign \new_[516]_  = \new_[264]_  | \new_[515]_ ;
  assign \new_[517]_  = \new_[516]_  | \new_[511]_ ;
  assign \new_[518]_  = \new_[517]_  | \new_[506]_ ;
  assign \new_[519]_  = \new_[518]_  | \new_[497]_ ;
  assign \new_[520]_  = \new_[519]_  | \new_[476]_ ;
  assign \new_[521]_  = \new_[520]_  | \new_[433]_ ;
  assign \new_[524]_  = \new_[260]_  | \new_[261]_ ;
  assign \new_[528]_  = \new_[257]_  | \new_[258]_ ;
  assign \new_[529]_  = \new_[259]_  | \new_[528]_ ;
  assign \new_[530]_  = \new_[529]_  | \new_[524]_ ;
  assign \new_[533]_  = \new_[255]_  | \new_[256]_ ;
  assign \new_[537]_  = \new_[252]_  | \new_[253]_ ;
  assign \new_[538]_  = \new_[254]_  | \new_[537]_ ;
  assign \new_[539]_  = \new_[538]_  | \new_[533]_ ;
  assign \new_[540]_  = \new_[539]_  | \new_[530]_ ;
  assign \new_[543]_  = \new_[250]_  | \new_[251]_ ;
  assign \new_[547]_  = \new_[247]_  | \new_[248]_ ;
  assign \new_[548]_  = \new_[249]_  | \new_[547]_ ;
  assign \new_[549]_  = \new_[548]_  | \new_[543]_ ;
  assign \new_[553]_  = \new_[244]_  | \new_[245]_ ;
  assign \new_[554]_  = \new_[246]_  | \new_[553]_ ;
  assign \new_[558]_  = \new_[241]_  | \new_[242]_ ;
  assign \new_[559]_  = \new_[243]_  | \new_[558]_ ;
  assign \new_[560]_  = \new_[559]_  | \new_[554]_ ;
  assign \new_[561]_  = \new_[560]_  | \new_[549]_ ;
  assign \new_[562]_  = \new_[561]_  | \new_[540]_ ;
  assign \new_[565]_  = \new_[239]_  | \new_[240]_ ;
  assign \new_[569]_  = \new_[236]_  | \new_[237]_ ;
  assign \new_[570]_  = \new_[238]_  | \new_[569]_ ;
  assign \new_[571]_  = \new_[570]_  | \new_[565]_ ;
  assign \new_[575]_  = \new_[233]_  | \new_[234]_ ;
  assign \new_[576]_  = \new_[235]_  | \new_[575]_ ;
  assign \new_[580]_  = \new_[230]_  | \new_[231]_ ;
  assign \new_[581]_  = \new_[232]_  | \new_[580]_ ;
  assign \new_[582]_  = \new_[581]_  | \new_[576]_ ;
  assign \new_[583]_  = \new_[582]_  | \new_[571]_ ;
  assign \new_[586]_  = \new_[228]_  | \new_[229]_ ;
  assign \new_[590]_  = \new_[225]_  | \new_[226]_ ;
  assign \new_[591]_  = \new_[227]_  | \new_[590]_ ;
  assign \new_[592]_  = \new_[591]_  | \new_[586]_ ;
  assign \new_[596]_  = \new_[222]_  | \new_[223]_ ;
  assign \new_[597]_  = \new_[224]_  | \new_[596]_ ;
  assign \new_[601]_  = \new_[219]_  | \new_[220]_ ;
  assign \new_[602]_  = \new_[221]_  | \new_[601]_ ;
  assign \new_[603]_  = \new_[602]_  | \new_[597]_ ;
  assign \new_[604]_  = \new_[603]_  | \new_[592]_ ;
  assign \new_[605]_  = \new_[604]_  | \new_[583]_ ;
  assign \new_[606]_  = \new_[605]_  | \new_[562]_ ;
  assign \new_[609]_  = \new_[217]_  | \new_[218]_ ;
  assign \new_[613]_  = \new_[214]_  | \new_[215]_ ;
  assign \new_[614]_  = \new_[216]_  | \new_[613]_ ;
  assign \new_[615]_  = \new_[614]_  | \new_[609]_ ;
  assign \new_[619]_  = \new_[211]_  | \new_[212]_ ;
  assign \new_[620]_  = \new_[213]_  | \new_[619]_ ;
  assign \new_[624]_  = \new_[208]_  | \new_[209]_ ;
  assign \new_[625]_  = \new_[210]_  | \new_[624]_ ;
  assign \new_[626]_  = \new_[625]_  | \new_[620]_ ;
  assign \new_[627]_  = \new_[626]_  | \new_[615]_ ;
  assign \new_[630]_  = \new_[206]_  | \new_[207]_ ;
  assign \new_[634]_  = \new_[203]_  | \new_[204]_ ;
  assign \new_[635]_  = \new_[205]_  | \new_[634]_ ;
  assign \new_[636]_  = \new_[635]_  | \new_[630]_ ;
  assign \new_[640]_  = \new_[200]_  | \new_[201]_ ;
  assign \new_[641]_  = \new_[202]_  | \new_[640]_ ;
  assign \new_[645]_  = \new_[197]_  | \new_[198]_ ;
  assign \new_[646]_  = \new_[199]_  | \new_[645]_ ;
  assign \new_[647]_  = \new_[646]_  | \new_[641]_ ;
  assign \new_[648]_  = \new_[647]_  | \new_[636]_ ;
  assign \new_[649]_  = \new_[648]_  | \new_[627]_ ;
  assign \new_[652]_  = \new_[195]_  | \new_[196]_ ;
  assign \new_[656]_  = \new_[192]_  | \new_[193]_ ;
  assign \new_[657]_  = \new_[194]_  | \new_[656]_ ;
  assign \new_[658]_  = \new_[657]_  | \new_[652]_ ;
  assign \new_[662]_  = \new_[189]_  | \new_[190]_ ;
  assign \new_[663]_  = \new_[191]_  | \new_[662]_ ;
  assign \new_[667]_  = \new_[186]_  | \new_[187]_ ;
  assign \new_[668]_  = \new_[188]_  | \new_[667]_ ;
  assign \new_[669]_  = \new_[668]_  | \new_[663]_ ;
  assign \new_[670]_  = \new_[669]_  | \new_[658]_ ;
  assign \new_[673]_  = \new_[184]_  | \new_[185]_ ;
  assign \new_[677]_  = \new_[181]_  | \new_[182]_ ;
  assign \new_[678]_  = \new_[183]_  | \new_[677]_ ;
  assign \new_[679]_  = \new_[678]_  | \new_[673]_ ;
  assign \new_[683]_  = \new_[178]_  | \new_[179]_ ;
  assign \new_[684]_  = \new_[180]_  | \new_[683]_ ;
  assign \new_[688]_  = \new_[175]_  | \new_[176]_ ;
  assign \new_[689]_  = \new_[177]_  | \new_[688]_ ;
  assign \new_[690]_  = \new_[689]_  | \new_[684]_ ;
  assign \new_[691]_  = \new_[690]_  | \new_[679]_ ;
  assign \new_[692]_  = \new_[691]_  | \new_[670]_ ;
  assign \new_[693]_  = \new_[692]_  | \new_[649]_ ;
  assign \new_[694]_  = \new_[693]_  | \new_[606]_ ;
  assign \new_[695]_  = \new_[694]_  | \new_[521]_ ;
  assign \new_[698]_  = \new_[173]_  | \new_[174]_ ;
  assign \new_[702]_  = \new_[170]_  | \new_[171]_ ;
  assign \new_[703]_  = \new_[172]_  | \new_[702]_ ;
  assign \new_[704]_  = \new_[703]_  | \new_[698]_ ;
  assign \new_[707]_  = \new_[168]_  | \new_[169]_ ;
  assign \new_[711]_  = \new_[165]_  | \new_[166]_ ;
  assign \new_[712]_  = \new_[167]_  | \new_[711]_ ;
  assign \new_[713]_  = \new_[712]_  | \new_[707]_ ;
  assign \new_[714]_  = \new_[713]_  | \new_[704]_ ;
  assign \new_[717]_  = \new_[163]_  | \new_[164]_ ;
  assign \new_[721]_  = \new_[160]_  | \new_[161]_ ;
  assign \new_[722]_  = \new_[162]_  | \new_[721]_ ;
  assign \new_[723]_  = \new_[722]_  | \new_[717]_ ;
  assign \new_[727]_  = \new_[157]_  | \new_[158]_ ;
  assign \new_[728]_  = \new_[159]_  | \new_[727]_ ;
  assign \new_[732]_  = \new_[154]_  | \new_[155]_ ;
  assign \new_[733]_  = \new_[156]_  | \new_[732]_ ;
  assign \new_[734]_  = \new_[733]_  | \new_[728]_ ;
  assign \new_[735]_  = \new_[734]_  | \new_[723]_ ;
  assign \new_[736]_  = \new_[735]_  | \new_[714]_ ;
  assign \new_[739]_  = \new_[152]_  | \new_[153]_ ;
  assign \new_[743]_  = \new_[149]_  | \new_[150]_ ;
  assign \new_[744]_  = \new_[151]_  | \new_[743]_ ;
  assign \new_[745]_  = \new_[744]_  | \new_[739]_ ;
  assign \new_[749]_  = \new_[146]_  | \new_[147]_ ;
  assign \new_[750]_  = \new_[148]_  | \new_[749]_ ;
  assign \new_[754]_  = \new_[143]_  | \new_[144]_ ;
  assign \new_[755]_  = \new_[145]_  | \new_[754]_ ;
  assign \new_[756]_  = \new_[755]_  | \new_[750]_ ;
  assign \new_[757]_  = \new_[756]_  | \new_[745]_ ;
  assign \new_[760]_  = \new_[141]_  | \new_[142]_ ;
  assign \new_[764]_  = \new_[138]_  | \new_[139]_ ;
  assign \new_[765]_  = \new_[140]_  | \new_[764]_ ;
  assign \new_[766]_  = \new_[765]_  | \new_[760]_ ;
  assign \new_[770]_  = \new_[135]_  | \new_[136]_ ;
  assign \new_[771]_  = \new_[137]_  | \new_[770]_ ;
  assign \new_[775]_  = \new_[132]_  | \new_[133]_ ;
  assign \new_[776]_  = \new_[134]_  | \new_[775]_ ;
  assign \new_[777]_  = \new_[776]_  | \new_[771]_ ;
  assign \new_[778]_  = \new_[777]_  | \new_[766]_ ;
  assign \new_[779]_  = \new_[778]_  | \new_[757]_ ;
  assign \new_[780]_  = \new_[779]_  | \new_[736]_ ;
  assign \new_[783]_  = \new_[130]_  | \new_[131]_ ;
  assign \new_[787]_  = \new_[127]_  | \new_[128]_ ;
  assign \new_[788]_  = \new_[129]_  | \new_[787]_ ;
  assign \new_[789]_  = \new_[788]_  | \new_[783]_ ;
  assign \new_[793]_  = \new_[124]_  | \new_[125]_ ;
  assign \new_[794]_  = \new_[126]_  | \new_[793]_ ;
  assign \new_[798]_  = \new_[121]_  | \new_[122]_ ;
  assign \new_[799]_  = \new_[123]_  | \new_[798]_ ;
  assign \new_[800]_  = \new_[799]_  | \new_[794]_ ;
  assign \new_[801]_  = \new_[800]_  | \new_[789]_ ;
  assign \new_[804]_  = \new_[119]_  | \new_[120]_ ;
  assign \new_[808]_  = \new_[116]_  | \new_[117]_ ;
  assign \new_[809]_  = \new_[118]_  | \new_[808]_ ;
  assign \new_[810]_  = \new_[809]_  | \new_[804]_ ;
  assign \new_[814]_  = \new_[113]_  | \new_[114]_ ;
  assign \new_[815]_  = \new_[115]_  | \new_[814]_ ;
  assign \new_[819]_  = \new_[110]_  | \new_[111]_ ;
  assign \new_[820]_  = \new_[112]_  | \new_[819]_ ;
  assign \new_[821]_  = \new_[820]_  | \new_[815]_ ;
  assign \new_[822]_  = \new_[821]_  | \new_[810]_ ;
  assign \new_[823]_  = \new_[822]_  | \new_[801]_ ;
  assign \new_[826]_  = \new_[108]_  | \new_[109]_ ;
  assign \new_[830]_  = \new_[105]_  | \new_[106]_ ;
  assign \new_[831]_  = \new_[107]_  | \new_[830]_ ;
  assign \new_[832]_  = \new_[831]_  | \new_[826]_ ;
  assign \new_[836]_  = \new_[102]_  | \new_[103]_ ;
  assign \new_[837]_  = \new_[104]_  | \new_[836]_ ;
  assign \new_[841]_  = \new_[99]_  | \new_[100]_ ;
  assign \new_[842]_  = \new_[101]_  | \new_[841]_ ;
  assign \new_[843]_  = \new_[842]_  | \new_[837]_ ;
  assign \new_[844]_  = \new_[843]_  | \new_[832]_ ;
  assign \new_[847]_  = \new_[97]_  | \new_[98]_ ;
  assign \new_[851]_  = \new_[94]_  | \new_[95]_ ;
  assign \new_[852]_  = \new_[96]_  | \new_[851]_ ;
  assign \new_[853]_  = \new_[852]_  | \new_[847]_ ;
  assign \new_[857]_  = \new_[91]_  | \new_[92]_ ;
  assign \new_[858]_  = \new_[93]_  | \new_[857]_ ;
  assign \new_[862]_  = \new_[88]_  | \new_[89]_ ;
  assign \new_[863]_  = \new_[90]_  | \new_[862]_ ;
  assign \new_[864]_  = \new_[863]_  | \new_[858]_ ;
  assign \new_[865]_  = \new_[864]_  | \new_[853]_ ;
  assign \new_[866]_  = \new_[865]_  | \new_[844]_ ;
  assign \new_[867]_  = \new_[866]_  | \new_[823]_ ;
  assign \new_[868]_  = \new_[867]_  | \new_[780]_ ;
  assign \new_[871]_  = \new_[86]_  | \new_[87]_ ;
  assign \new_[875]_  = \new_[83]_  | \new_[84]_ ;
  assign \new_[876]_  = \new_[85]_  | \new_[875]_ ;
  assign \new_[877]_  = \new_[876]_  | \new_[871]_ ;
  assign \new_[880]_  = \new_[81]_  | \new_[82]_ ;
  assign \new_[884]_  = \new_[78]_  | \new_[79]_ ;
  assign \new_[885]_  = \new_[80]_  | \new_[884]_ ;
  assign \new_[886]_  = \new_[885]_  | \new_[880]_ ;
  assign \new_[887]_  = \new_[886]_  | \new_[877]_ ;
  assign \new_[890]_  = \new_[76]_  | \new_[77]_ ;
  assign \new_[894]_  = \new_[73]_  | \new_[74]_ ;
  assign \new_[895]_  = \new_[75]_  | \new_[894]_ ;
  assign \new_[896]_  = \new_[895]_  | \new_[890]_ ;
  assign \new_[900]_  = \new_[70]_  | \new_[71]_ ;
  assign \new_[901]_  = \new_[72]_  | \new_[900]_ ;
  assign \new_[905]_  = \new_[67]_  | \new_[68]_ ;
  assign \new_[906]_  = \new_[69]_  | \new_[905]_ ;
  assign \new_[907]_  = \new_[906]_  | \new_[901]_ ;
  assign \new_[908]_  = \new_[907]_  | \new_[896]_ ;
  assign \new_[909]_  = \new_[908]_  | \new_[887]_ ;
  assign \new_[912]_  = \new_[65]_  | \new_[66]_ ;
  assign \new_[916]_  = \new_[62]_  | \new_[63]_ ;
  assign \new_[917]_  = \new_[64]_  | \new_[916]_ ;
  assign \new_[918]_  = \new_[917]_  | \new_[912]_ ;
  assign \new_[922]_  = \new_[59]_  | \new_[60]_ ;
  assign \new_[923]_  = \new_[61]_  | \new_[922]_ ;
  assign \new_[927]_  = \new_[56]_  | \new_[57]_ ;
  assign \new_[928]_  = \new_[58]_  | \new_[927]_ ;
  assign \new_[929]_  = \new_[928]_  | \new_[923]_ ;
  assign \new_[930]_  = \new_[929]_  | \new_[918]_ ;
  assign \new_[933]_  = \new_[54]_  | \new_[55]_ ;
  assign \new_[937]_  = \new_[51]_  | \new_[52]_ ;
  assign \new_[938]_  = \new_[53]_  | \new_[937]_ ;
  assign \new_[939]_  = \new_[938]_  | \new_[933]_ ;
  assign \new_[943]_  = \new_[48]_  | \new_[49]_ ;
  assign \new_[944]_  = \new_[50]_  | \new_[943]_ ;
  assign \new_[948]_  = \new_[45]_  | \new_[46]_ ;
  assign \new_[949]_  = \new_[47]_  | \new_[948]_ ;
  assign \new_[950]_  = \new_[949]_  | \new_[944]_ ;
  assign \new_[951]_  = \new_[950]_  | \new_[939]_ ;
  assign \new_[952]_  = \new_[951]_  | \new_[930]_ ;
  assign \new_[953]_  = \new_[952]_  | \new_[909]_ ;
  assign \new_[956]_  = \new_[43]_  | \new_[44]_ ;
  assign \new_[960]_  = \new_[40]_  | \new_[41]_ ;
  assign \new_[961]_  = \new_[42]_  | \new_[960]_ ;
  assign \new_[962]_  = \new_[961]_  | \new_[956]_ ;
  assign \new_[966]_  = \new_[37]_  | \new_[38]_ ;
  assign \new_[967]_  = \new_[39]_  | \new_[966]_ ;
  assign \new_[971]_  = \new_[34]_  | \new_[35]_ ;
  assign \new_[972]_  = \new_[36]_  | \new_[971]_ ;
  assign \new_[973]_  = \new_[972]_  | \new_[967]_ ;
  assign \new_[974]_  = \new_[973]_  | \new_[962]_ ;
  assign \new_[977]_  = \new_[32]_  | \new_[33]_ ;
  assign \new_[981]_  = \new_[29]_  | \new_[30]_ ;
  assign \new_[982]_  = \new_[31]_  | \new_[981]_ ;
  assign \new_[983]_  = \new_[982]_  | \new_[977]_ ;
  assign \new_[987]_  = \new_[26]_  | \new_[27]_ ;
  assign \new_[988]_  = \new_[28]_  | \new_[987]_ ;
  assign \new_[992]_  = \new_[23]_  | \new_[24]_ ;
  assign \new_[993]_  = \new_[25]_  | \new_[992]_ ;
  assign \new_[994]_  = \new_[993]_  | \new_[988]_ ;
  assign \new_[995]_  = \new_[994]_  | \new_[983]_ ;
  assign \new_[996]_  = \new_[995]_  | \new_[974]_ ;
  assign \new_[999]_  = \new_[21]_  | \new_[22]_ ;
  assign \new_[1003]_  = \new_[18]_  | \new_[19]_ ;
  assign \new_[1004]_  = \new_[20]_  | \new_[1003]_ ;
  assign \new_[1005]_  = \new_[1004]_  | \new_[999]_ ;
  assign \new_[1009]_  = \new_[15]_  | \new_[16]_ ;
  assign \new_[1010]_  = \new_[17]_  | \new_[1009]_ ;
  assign \new_[1014]_  = \new_[12]_  | \new_[13]_ ;
  assign \new_[1015]_  = \new_[14]_  | \new_[1014]_ ;
  assign \new_[1016]_  = \new_[1015]_  | \new_[1010]_ ;
  assign \new_[1017]_  = \new_[1016]_  | \new_[1005]_ ;
  assign \new_[1020]_  = \new_[10]_  | \new_[11]_ ;
  assign \new_[1024]_  = \new_[7]_  | \new_[8]_ ;
  assign \new_[1025]_  = \new_[9]_  | \new_[1024]_ ;
  assign \new_[1026]_  = \new_[1025]_  | \new_[1020]_ ;
  assign \new_[1030]_  = \new_[4]_  | \new_[5]_ ;
  assign \new_[1031]_  = \new_[6]_  | \new_[1030]_ ;
  assign \new_[1035]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[1036]_  = \new_[3]_  | \new_[1035]_ ;
  assign \new_[1037]_  = \new_[1036]_  | \new_[1031]_ ;
  assign \new_[1038]_  = \new_[1037]_  | \new_[1026]_ ;
  assign \new_[1039]_  = \new_[1038]_  | \new_[1017]_ ;
  assign \new_[1040]_  = \new_[1039]_  | \new_[996]_ ;
  assign \new_[1041]_  = \new_[1040]_  | \new_[953]_ ;
  assign \new_[1042]_  = \new_[1041]_  | \new_[868]_ ;
  assign \new_[1049]_  = A266 & A265;
  assign \new_[1052]_  = ~A269 & A268;
  assign \new_[1055]_  = A266 & ~A265;
  assign \new_[1058]_  = A269 & ~A268;
  assign \new_[1061]_  = ~A266 & A265;
  assign \new_[1064]_  = A269 & ~A268;
  assign \new_[1067]_  = ~A266 & ~A265;
  assign \new_[1070]_  = ~A269 & A268;
  assign \new_[1073]_  = A201 & A199;
  assign \new_[1076]_  = A234 & A232;
  assign \new_[1079]_  = A201 & A199;
  assign \new_[1082]_  = A234 & A233;
  assign \new_[1085]_  = A201 & A200;
  assign \new_[1088]_  = A234 & A232;
  assign \new_[1091]_  = A201 & A200;
  assign \new_[1094]_  = A234 & A233;
  assign \new_[1097]_  = ~A166 & A167;
  assign \new_[1100]_  = A234 & A232;
  assign \new_[1103]_  = ~A166 & A167;
  assign \new_[1106]_  = A234 & A233;
  assign \new_[1110]_  = A232 & A201;
  assign \new_[1111]_  = A199 & \new_[1110]_ ;
  assign \new_[1115]_  = ~A236 & A235;
  assign \new_[1116]_  = A233 & \new_[1115]_ ;
  assign \new_[1120]_  = ~A232 & A201;
  assign \new_[1121]_  = A199 & \new_[1120]_ ;
  assign \new_[1125]_  = A236 & ~A235;
  assign \new_[1126]_  = A233 & \new_[1125]_ ;
  assign \new_[1130]_  = A232 & A201;
  assign \new_[1131]_  = A199 & \new_[1130]_ ;
  assign \new_[1135]_  = A236 & ~A235;
  assign \new_[1136]_  = ~A233 & \new_[1135]_ ;
  assign \new_[1140]_  = ~A232 & A201;
  assign \new_[1141]_  = A199 & \new_[1140]_ ;
  assign \new_[1145]_  = ~A236 & A235;
  assign \new_[1146]_  = ~A233 & \new_[1145]_ ;
  assign \new_[1150]_  = A232 & A201;
  assign \new_[1151]_  = A200 & \new_[1150]_ ;
  assign \new_[1155]_  = ~A236 & A235;
  assign \new_[1156]_  = A233 & \new_[1155]_ ;
  assign \new_[1160]_  = ~A232 & A201;
  assign \new_[1161]_  = A200 & \new_[1160]_ ;
  assign \new_[1165]_  = A236 & ~A235;
  assign \new_[1166]_  = A233 & \new_[1165]_ ;
  assign \new_[1170]_  = A232 & A201;
  assign \new_[1171]_  = A200 & \new_[1170]_ ;
  assign \new_[1175]_  = A236 & ~A235;
  assign \new_[1176]_  = ~A233 & \new_[1175]_ ;
  assign \new_[1180]_  = ~A232 & A201;
  assign \new_[1181]_  = A200 & \new_[1180]_ ;
  assign \new_[1185]_  = ~A236 & A235;
  assign \new_[1186]_  = ~A233 & \new_[1185]_ ;
  assign \new_[1190]_  = A202 & A200;
  assign \new_[1191]_  = A199 & \new_[1190]_ ;
  assign \new_[1195]_  = A234 & A232;
  assign \new_[1196]_  = ~A203 & \new_[1195]_ ;
  assign \new_[1200]_  = A202 & A200;
  assign \new_[1201]_  = A199 & \new_[1200]_ ;
  assign \new_[1205]_  = A234 & A233;
  assign \new_[1206]_  = ~A203 & \new_[1205]_ ;
  assign \new_[1210]_  = ~A202 & A200;
  assign \new_[1211]_  = ~A199 & \new_[1210]_ ;
  assign \new_[1215]_  = A234 & A232;
  assign \new_[1216]_  = A203 & \new_[1215]_ ;
  assign \new_[1220]_  = ~A202 & A200;
  assign \new_[1221]_  = ~A199 & \new_[1220]_ ;
  assign \new_[1225]_  = A234 & A233;
  assign \new_[1226]_  = A203 & \new_[1225]_ ;
  assign \new_[1230]_  = ~A202 & ~A200;
  assign \new_[1231]_  = A199 & \new_[1230]_ ;
  assign \new_[1235]_  = A234 & A232;
  assign \new_[1236]_  = A203 & \new_[1235]_ ;
  assign \new_[1240]_  = ~A202 & ~A200;
  assign \new_[1241]_  = A199 & \new_[1240]_ ;
  assign \new_[1245]_  = A234 & A233;
  assign \new_[1246]_  = A203 & \new_[1245]_ ;
  assign \new_[1250]_  = A202 & ~A200;
  assign \new_[1251]_  = ~A199 & \new_[1250]_ ;
  assign \new_[1255]_  = A234 & A232;
  assign \new_[1256]_  = ~A203 & \new_[1255]_ ;
  assign \new_[1260]_  = A202 & ~A200;
  assign \new_[1261]_  = ~A199 & \new_[1260]_ ;
  assign \new_[1265]_  = A234 & A233;
  assign \new_[1266]_  = ~A203 & \new_[1265]_ ;
  assign \new_[1270]_  = A199 & A166;
  assign \new_[1271]_  = A167 & \new_[1270]_ ;
  assign \new_[1275]_  = A300 & A299;
  assign \new_[1276]_  = A201 & \new_[1275]_ ;
  assign \new_[1280]_  = A199 & A166;
  assign \new_[1281]_  = A167 & \new_[1280]_ ;
  assign \new_[1285]_  = A300 & A298;
  assign \new_[1286]_  = A201 & \new_[1285]_ ;
  assign \new_[1290]_  = A200 & A166;
  assign \new_[1291]_  = A167 & \new_[1290]_ ;
  assign \new_[1295]_  = A300 & A299;
  assign \new_[1296]_  = A201 & \new_[1295]_ ;
  assign \new_[1300]_  = A200 & A166;
  assign \new_[1301]_  = A167 & \new_[1300]_ ;
  assign \new_[1305]_  = A300 & A298;
  assign \new_[1306]_  = A201 & \new_[1305]_ ;
  assign \new_[1310]_  = A232 & ~A166;
  assign \new_[1311]_  = A167 & \new_[1310]_ ;
  assign \new_[1315]_  = ~A236 & A235;
  assign \new_[1316]_  = A233 & \new_[1315]_ ;
  assign \new_[1320]_  = ~A232 & ~A166;
  assign \new_[1321]_  = A167 & \new_[1320]_ ;
  assign \new_[1325]_  = A236 & ~A235;
  assign \new_[1326]_  = A233 & \new_[1325]_ ;
  assign \new_[1330]_  = A232 & ~A166;
  assign \new_[1331]_  = A167 & \new_[1330]_ ;
  assign \new_[1335]_  = A236 & ~A235;
  assign \new_[1336]_  = ~A233 & \new_[1335]_ ;
  assign \new_[1340]_  = ~A232 & ~A166;
  assign \new_[1341]_  = A167 & \new_[1340]_ ;
  assign \new_[1345]_  = ~A236 & A235;
  assign \new_[1346]_  = ~A233 & \new_[1345]_ ;
  assign \new_[1350]_  = A199 & ~A166;
  assign \new_[1351]_  = ~A167 & \new_[1350]_ ;
  assign \new_[1355]_  = A300 & A299;
  assign \new_[1356]_  = A201 & \new_[1355]_ ;
  assign \new_[1360]_  = A199 & ~A166;
  assign \new_[1361]_  = ~A167 & \new_[1360]_ ;
  assign \new_[1365]_  = A300 & A298;
  assign \new_[1366]_  = A201 & \new_[1365]_ ;
  assign \new_[1370]_  = A200 & ~A166;
  assign \new_[1371]_  = ~A167 & \new_[1370]_ ;
  assign \new_[1375]_  = A300 & A299;
  assign \new_[1376]_  = A201 & \new_[1375]_ ;
  assign \new_[1380]_  = A200 & ~A166;
  assign \new_[1381]_  = ~A167 & \new_[1380]_ ;
  assign \new_[1385]_  = A300 & A298;
  assign \new_[1386]_  = A201 & \new_[1385]_ ;
  assign \new_[1390]_  = A199 & ~A167;
  assign \new_[1391]_  = ~A168 & \new_[1390]_ ;
  assign \new_[1395]_  = A300 & A299;
  assign \new_[1396]_  = A201 & \new_[1395]_ ;
  assign \new_[1400]_  = A199 & ~A167;
  assign \new_[1401]_  = ~A168 & \new_[1400]_ ;
  assign \new_[1405]_  = A300 & A298;
  assign \new_[1406]_  = A201 & \new_[1405]_ ;
  assign \new_[1410]_  = A200 & ~A167;
  assign \new_[1411]_  = ~A168 & \new_[1410]_ ;
  assign \new_[1415]_  = A300 & A299;
  assign \new_[1416]_  = A201 & \new_[1415]_ ;
  assign \new_[1420]_  = A200 & ~A167;
  assign \new_[1421]_  = ~A168 & \new_[1420]_ ;
  assign \new_[1425]_  = A300 & A298;
  assign \new_[1426]_  = A201 & \new_[1425]_ ;
  assign \new_[1430]_  = ~A167 & A168;
  assign \new_[1431]_  = A170 & \new_[1430]_ ;
  assign \new_[1435]_  = A234 & A232;
  assign \new_[1436]_  = A166 & \new_[1435]_ ;
  assign \new_[1440]_  = ~A167 & A168;
  assign \new_[1441]_  = A170 & \new_[1440]_ ;
  assign \new_[1445]_  = A234 & A233;
  assign \new_[1446]_  = A166 & \new_[1445]_ ;
  assign \new_[1450]_  = ~A167 & A168;
  assign \new_[1451]_  = A169 & \new_[1450]_ ;
  assign \new_[1455]_  = A234 & A232;
  assign \new_[1456]_  = A166 & \new_[1455]_ ;
  assign \new_[1460]_  = ~A167 & A168;
  assign \new_[1461]_  = A169 & \new_[1460]_ ;
  assign \new_[1465]_  = A234 & A233;
  assign \new_[1466]_  = A166 & \new_[1465]_ ;
  assign \new_[1470]_  = ~A199 & ~A166;
  assign \new_[1471]_  = A167 & \new_[1470]_ ;
  assign \new_[1474]_  = ~A202 & ~A200;
  assign \new_[1477]_  = A300 & A299;
  assign \new_[1478]_  = \new_[1477]_  & \new_[1474]_ ;
  assign \new_[1482]_  = ~A199 & ~A166;
  assign \new_[1483]_  = A167 & \new_[1482]_ ;
  assign \new_[1486]_  = ~A202 & ~A200;
  assign \new_[1489]_  = A300 & A298;
  assign \new_[1490]_  = \new_[1489]_  & \new_[1486]_ ;
  assign \new_[1494]_  = ~A199 & ~A166;
  assign \new_[1495]_  = A167 & \new_[1494]_ ;
  assign \new_[1498]_  = A203 & ~A200;
  assign \new_[1501]_  = A300 & A299;
  assign \new_[1502]_  = \new_[1501]_  & \new_[1498]_ ;
  assign \new_[1506]_  = ~A199 & ~A166;
  assign \new_[1507]_  = A167 & \new_[1506]_ ;
  assign \new_[1510]_  = A203 & ~A200;
  assign \new_[1513]_  = A300 & A298;
  assign \new_[1514]_  = \new_[1513]_  & \new_[1510]_ ;
  assign \new_[1518]_  = ~A167 & ~A169;
  assign \new_[1519]_  = ~A170 & \new_[1518]_ ;
  assign \new_[1522]_  = A201 & A199;
  assign \new_[1525]_  = A300 & A299;
  assign \new_[1526]_  = \new_[1525]_  & \new_[1522]_ ;
  assign \new_[1530]_  = ~A167 & ~A169;
  assign \new_[1531]_  = ~A170 & \new_[1530]_ ;
  assign \new_[1534]_  = A201 & A199;
  assign \new_[1537]_  = A300 & A298;
  assign \new_[1538]_  = \new_[1537]_  & \new_[1534]_ ;
  assign \new_[1542]_  = ~A167 & ~A169;
  assign \new_[1543]_  = ~A170 & \new_[1542]_ ;
  assign \new_[1546]_  = A201 & A200;
  assign \new_[1549]_  = A300 & A299;
  assign \new_[1550]_  = \new_[1549]_  & \new_[1546]_ ;
  assign \new_[1554]_  = ~A167 & ~A169;
  assign \new_[1555]_  = ~A170 & \new_[1554]_ ;
  assign \new_[1558]_  = A201 & A200;
  assign \new_[1561]_  = A300 & A298;
  assign \new_[1562]_  = \new_[1561]_  & \new_[1558]_ ;
  assign \new_[1565]_  = A200 & A199;
  assign \new_[1568]_  = ~A203 & A202;
  assign \new_[1569]_  = \new_[1568]_  & \new_[1565]_ ;
  assign \new_[1572]_  = A233 & A232;
  assign \new_[1575]_  = ~A236 & A235;
  assign \new_[1576]_  = \new_[1575]_  & \new_[1572]_ ;
  assign \new_[1579]_  = A200 & A199;
  assign \new_[1582]_  = ~A203 & A202;
  assign \new_[1583]_  = \new_[1582]_  & \new_[1579]_ ;
  assign \new_[1586]_  = A233 & ~A232;
  assign \new_[1589]_  = A236 & ~A235;
  assign \new_[1590]_  = \new_[1589]_  & \new_[1586]_ ;
  assign \new_[1593]_  = A200 & A199;
  assign \new_[1596]_  = ~A203 & A202;
  assign \new_[1597]_  = \new_[1596]_  & \new_[1593]_ ;
  assign \new_[1600]_  = ~A233 & A232;
  assign \new_[1603]_  = A236 & ~A235;
  assign \new_[1604]_  = \new_[1603]_  & \new_[1600]_ ;
  assign \new_[1607]_  = A200 & A199;
  assign \new_[1610]_  = ~A203 & A202;
  assign \new_[1611]_  = \new_[1610]_  & \new_[1607]_ ;
  assign \new_[1614]_  = ~A233 & ~A232;
  assign \new_[1617]_  = ~A236 & A235;
  assign \new_[1618]_  = \new_[1617]_  & \new_[1614]_ ;
  assign \new_[1621]_  = A200 & ~A199;
  assign \new_[1624]_  = A203 & ~A202;
  assign \new_[1625]_  = \new_[1624]_  & \new_[1621]_ ;
  assign \new_[1628]_  = A233 & A232;
  assign \new_[1631]_  = ~A236 & A235;
  assign \new_[1632]_  = \new_[1631]_  & \new_[1628]_ ;
  assign \new_[1635]_  = A200 & ~A199;
  assign \new_[1638]_  = A203 & ~A202;
  assign \new_[1639]_  = \new_[1638]_  & \new_[1635]_ ;
  assign \new_[1642]_  = A233 & ~A232;
  assign \new_[1645]_  = A236 & ~A235;
  assign \new_[1646]_  = \new_[1645]_  & \new_[1642]_ ;
  assign \new_[1649]_  = A200 & ~A199;
  assign \new_[1652]_  = A203 & ~A202;
  assign \new_[1653]_  = \new_[1652]_  & \new_[1649]_ ;
  assign \new_[1656]_  = ~A233 & A232;
  assign \new_[1659]_  = A236 & ~A235;
  assign \new_[1660]_  = \new_[1659]_  & \new_[1656]_ ;
  assign \new_[1663]_  = A200 & ~A199;
  assign \new_[1666]_  = A203 & ~A202;
  assign \new_[1667]_  = \new_[1666]_  & \new_[1663]_ ;
  assign \new_[1670]_  = ~A233 & ~A232;
  assign \new_[1673]_  = ~A236 & A235;
  assign \new_[1674]_  = \new_[1673]_  & \new_[1670]_ ;
  assign \new_[1677]_  = ~A200 & A199;
  assign \new_[1680]_  = A203 & ~A202;
  assign \new_[1681]_  = \new_[1680]_  & \new_[1677]_ ;
  assign \new_[1684]_  = A233 & A232;
  assign \new_[1687]_  = ~A236 & A235;
  assign \new_[1688]_  = \new_[1687]_  & \new_[1684]_ ;
  assign \new_[1691]_  = ~A200 & A199;
  assign \new_[1694]_  = A203 & ~A202;
  assign \new_[1695]_  = \new_[1694]_  & \new_[1691]_ ;
  assign \new_[1698]_  = A233 & ~A232;
  assign \new_[1701]_  = A236 & ~A235;
  assign \new_[1702]_  = \new_[1701]_  & \new_[1698]_ ;
  assign \new_[1705]_  = ~A200 & A199;
  assign \new_[1708]_  = A203 & ~A202;
  assign \new_[1709]_  = \new_[1708]_  & \new_[1705]_ ;
  assign \new_[1712]_  = ~A233 & A232;
  assign \new_[1715]_  = A236 & ~A235;
  assign \new_[1716]_  = \new_[1715]_  & \new_[1712]_ ;
  assign \new_[1719]_  = ~A200 & A199;
  assign \new_[1722]_  = A203 & ~A202;
  assign \new_[1723]_  = \new_[1722]_  & \new_[1719]_ ;
  assign \new_[1726]_  = ~A233 & ~A232;
  assign \new_[1729]_  = ~A236 & A235;
  assign \new_[1730]_  = \new_[1729]_  & \new_[1726]_ ;
  assign \new_[1733]_  = ~A200 & ~A199;
  assign \new_[1736]_  = ~A203 & A202;
  assign \new_[1737]_  = \new_[1736]_  & \new_[1733]_ ;
  assign \new_[1740]_  = A233 & A232;
  assign \new_[1743]_  = ~A236 & A235;
  assign \new_[1744]_  = \new_[1743]_  & \new_[1740]_ ;
  assign \new_[1747]_  = ~A200 & ~A199;
  assign \new_[1750]_  = ~A203 & A202;
  assign \new_[1751]_  = \new_[1750]_  & \new_[1747]_ ;
  assign \new_[1754]_  = A233 & ~A232;
  assign \new_[1757]_  = A236 & ~A235;
  assign \new_[1758]_  = \new_[1757]_  & \new_[1754]_ ;
  assign \new_[1761]_  = ~A200 & ~A199;
  assign \new_[1764]_  = ~A203 & A202;
  assign \new_[1765]_  = \new_[1764]_  & \new_[1761]_ ;
  assign \new_[1768]_  = ~A233 & A232;
  assign \new_[1771]_  = A236 & ~A235;
  assign \new_[1772]_  = \new_[1771]_  & \new_[1768]_ ;
  assign \new_[1775]_  = ~A200 & ~A199;
  assign \new_[1778]_  = ~A203 & A202;
  assign \new_[1779]_  = \new_[1778]_  & \new_[1775]_ ;
  assign \new_[1782]_  = ~A233 & ~A232;
  assign \new_[1785]_  = ~A236 & A235;
  assign \new_[1786]_  = \new_[1785]_  & \new_[1782]_ ;
  assign \new_[1789]_  = A166 & A167;
  assign \new_[1792]_  = A201 & A199;
  assign \new_[1793]_  = \new_[1792]_  & \new_[1789]_ ;
  assign \new_[1796]_  = A299 & A298;
  assign \new_[1799]_  = ~A302 & A301;
  assign \new_[1800]_  = \new_[1799]_  & \new_[1796]_ ;
  assign \new_[1803]_  = A166 & A167;
  assign \new_[1806]_  = A201 & A199;
  assign \new_[1807]_  = \new_[1806]_  & \new_[1803]_ ;
  assign \new_[1810]_  = ~A299 & A298;
  assign \new_[1813]_  = A302 & ~A301;
  assign \new_[1814]_  = \new_[1813]_  & \new_[1810]_ ;
  assign \new_[1817]_  = A166 & A167;
  assign \new_[1820]_  = A201 & A199;
  assign \new_[1821]_  = \new_[1820]_  & \new_[1817]_ ;
  assign \new_[1824]_  = A299 & ~A298;
  assign \new_[1827]_  = A302 & ~A301;
  assign \new_[1828]_  = \new_[1827]_  & \new_[1824]_ ;
  assign \new_[1831]_  = A166 & A167;
  assign \new_[1834]_  = A201 & A199;
  assign \new_[1835]_  = \new_[1834]_  & \new_[1831]_ ;
  assign \new_[1838]_  = ~A299 & ~A298;
  assign \new_[1841]_  = ~A302 & A301;
  assign \new_[1842]_  = \new_[1841]_  & \new_[1838]_ ;
  assign \new_[1845]_  = A166 & A167;
  assign \new_[1848]_  = A201 & A200;
  assign \new_[1849]_  = \new_[1848]_  & \new_[1845]_ ;
  assign \new_[1852]_  = A299 & A298;
  assign \new_[1855]_  = ~A302 & A301;
  assign \new_[1856]_  = \new_[1855]_  & \new_[1852]_ ;
  assign \new_[1859]_  = A166 & A167;
  assign \new_[1862]_  = A201 & A200;
  assign \new_[1863]_  = \new_[1862]_  & \new_[1859]_ ;
  assign \new_[1866]_  = ~A299 & A298;
  assign \new_[1869]_  = A302 & ~A301;
  assign \new_[1870]_  = \new_[1869]_  & \new_[1866]_ ;
  assign \new_[1873]_  = A166 & A167;
  assign \new_[1876]_  = A201 & A200;
  assign \new_[1877]_  = \new_[1876]_  & \new_[1873]_ ;
  assign \new_[1880]_  = A299 & ~A298;
  assign \new_[1883]_  = A302 & ~A301;
  assign \new_[1884]_  = \new_[1883]_  & \new_[1880]_ ;
  assign \new_[1887]_  = A166 & A167;
  assign \new_[1890]_  = A201 & A200;
  assign \new_[1891]_  = \new_[1890]_  & \new_[1887]_ ;
  assign \new_[1894]_  = ~A299 & ~A298;
  assign \new_[1897]_  = ~A302 & A301;
  assign \new_[1898]_  = \new_[1897]_  & \new_[1894]_ ;
  assign \new_[1901]_  = A166 & A167;
  assign \new_[1904]_  = A200 & A199;
  assign \new_[1905]_  = \new_[1904]_  & \new_[1901]_ ;
  assign \new_[1908]_  = ~A203 & A202;
  assign \new_[1911]_  = A300 & A299;
  assign \new_[1912]_  = \new_[1911]_  & \new_[1908]_ ;
  assign \new_[1915]_  = A166 & A167;
  assign \new_[1918]_  = A200 & A199;
  assign \new_[1919]_  = \new_[1918]_  & \new_[1915]_ ;
  assign \new_[1922]_  = ~A203 & A202;
  assign \new_[1925]_  = A300 & A298;
  assign \new_[1926]_  = \new_[1925]_  & \new_[1922]_ ;
  assign \new_[1929]_  = A166 & A167;
  assign \new_[1932]_  = A200 & ~A199;
  assign \new_[1933]_  = \new_[1932]_  & \new_[1929]_ ;
  assign \new_[1936]_  = A203 & ~A202;
  assign \new_[1939]_  = A300 & A299;
  assign \new_[1940]_  = \new_[1939]_  & \new_[1936]_ ;
  assign \new_[1943]_  = A166 & A167;
  assign \new_[1946]_  = A200 & ~A199;
  assign \new_[1947]_  = \new_[1946]_  & \new_[1943]_ ;
  assign \new_[1950]_  = A203 & ~A202;
  assign \new_[1953]_  = A300 & A298;
  assign \new_[1954]_  = \new_[1953]_  & \new_[1950]_ ;
  assign \new_[1957]_  = A166 & A167;
  assign \new_[1960]_  = ~A200 & A199;
  assign \new_[1961]_  = \new_[1960]_  & \new_[1957]_ ;
  assign \new_[1964]_  = A203 & ~A202;
  assign \new_[1967]_  = A300 & A299;
  assign \new_[1968]_  = \new_[1967]_  & \new_[1964]_ ;
  assign \new_[1971]_  = A166 & A167;
  assign \new_[1974]_  = ~A200 & A199;
  assign \new_[1975]_  = \new_[1974]_  & \new_[1971]_ ;
  assign \new_[1978]_  = A203 & ~A202;
  assign \new_[1981]_  = A300 & A298;
  assign \new_[1982]_  = \new_[1981]_  & \new_[1978]_ ;
  assign \new_[1985]_  = A166 & A167;
  assign \new_[1988]_  = ~A200 & ~A199;
  assign \new_[1989]_  = \new_[1988]_  & \new_[1985]_ ;
  assign \new_[1992]_  = ~A203 & A202;
  assign \new_[1995]_  = A300 & A299;
  assign \new_[1996]_  = \new_[1995]_  & \new_[1992]_ ;
  assign \new_[1999]_  = A166 & A167;
  assign \new_[2002]_  = ~A200 & ~A199;
  assign \new_[2003]_  = \new_[2002]_  & \new_[1999]_ ;
  assign \new_[2006]_  = ~A203 & A202;
  assign \new_[2009]_  = A300 & A298;
  assign \new_[2010]_  = \new_[2009]_  & \new_[2006]_ ;
  assign \new_[2013]_  = ~A166 & A167;
  assign \new_[2016]_  = A200 & A199;
  assign \new_[2017]_  = \new_[2016]_  & \new_[2013]_ ;
  assign \new_[2020]_  = ~A202 & ~A201;
  assign \new_[2023]_  = A300 & A299;
  assign \new_[2024]_  = \new_[2023]_  & \new_[2020]_ ;
  assign \new_[2027]_  = ~A166 & A167;
  assign \new_[2030]_  = A200 & A199;
  assign \new_[2031]_  = \new_[2030]_  & \new_[2027]_ ;
  assign \new_[2034]_  = ~A202 & ~A201;
  assign \new_[2037]_  = A300 & A298;
  assign \new_[2038]_  = \new_[2037]_  & \new_[2034]_ ;
  assign \new_[2041]_  = ~A166 & A167;
  assign \new_[2044]_  = A200 & A199;
  assign \new_[2045]_  = \new_[2044]_  & \new_[2041]_ ;
  assign \new_[2048]_  = A203 & ~A201;
  assign \new_[2051]_  = A300 & A299;
  assign \new_[2052]_  = \new_[2051]_  & \new_[2048]_ ;
  assign \new_[2055]_  = ~A166 & A167;
  assign \new_[2058]_  = A200 & A199;
  assign \new_[2059]_  = \new_[2058]_  & \new_[2055]_ ;
  assign \new_[2062]_  = A203 & ~A201;
  assign \new_[2065]_  = A300 & A298;
  assign \new_[2066]_  = \new_[2065]_  & \new_[2062]_ ;
  assign \new_[2069]_  = ~A166 & A167;
  assign \new_[2072]_  = A200 & ~A199;
  assign \new_[2073]_  = \new_[2072]_  & \new_[2069]_ ;
  assign \new_[2076]_  = A202 & ~A201;
  assign \new_[2079]_  = A300 & A299;
  assign \new_[2080]_  = \new_[2079]_  & \new_[2076]_ ;
  assign \new_[2083]_  = ~A166 & A167;
  assign \new_[2086]_  = A200 & ~A199;
  assign \new_[2087]_  = \new_[2086]_  & \new_[2083]_ ;
  assign \new_[2090]_  = A202 & ~A201;
  assign \new_[2093]_  = A300 & A298;
  assign \new_[2094]_  = \new_[2093]_  & \new_[2090]_ ;
  assign \new_[2097]_  = ~A166 & A167;
  assign \new_[2100]_  = A200 & ~A199;
  assign \new_[2101]_  = \new_[2100]_  & \new_[2097]_ ;
  assign \new_[2104]_  = ~A203 & ~A201;
  assign \new_[2107]_  = A300 & A299;
  assign \new_[2108]_  = \new_[2107]_  & \new_[2104]_ ;
  assign \new_[2111]_  = ~A166 & A167;
  assign \new_[2114]_  = A200 & ~A199;
  assign \new_[2115]_  = \new_[2114]_  & \new_[2111]_ ;
  assign \new_[2118]_  = ~A203 & ~A201;
  assign \new_[2121]_  = A300 & A298;
  assign \new_[2122]_  = \new_[2121]_  & \new_[2118]_ ;
  assign \new_[2125]_  = ~A166 & A167;
  assign \new_[2128]_  = ~A200 & A199;
  assign \new_[2129]_  = \new_[2128]_  & \new_[2125]_ ;
  assign \new_[2132]_  = A202 & ~A201;
  assign \new_[2135]_  = A300 & A299;
  assign \new_[2136]_  = \new_[2135]_  & \new_[2132]_ ;
  assign \new_[2139]_  = ~A166 & A167;
  assign \new_[2142]_  = ~A200 & A199;
  assign \new_[2143]_  = \new_[2142]_  & \new_[2139]_ ;
  assign \new_[2146]_  = A202 & ~A201;
  assign \new_[2149]_  = A300 & A298;
  assign \new_[2150]_  = \new_[2149]_  & \new_[2146]_ ;
  assign \new_[2153]_  = ~A166 & A167;
  assign \new_[2156]_  = ~A200 & A199;
  assign \new_[2157]_  = \new_[2156]_  & \new_[2153]_ ;
  assign \new_[2160]_  = ~A203 & ~A201;
  assign \new_[2163]_  = A300 & A299;
  assign \new_[2164]_  = \new_[2163]_  & \new_[2160]_ ;
  assign \new_[2167]_  = ~A166 & A167;
  assign \new_[2170]_  = ~A200 & A199;
  assign \new_[2171]_  = \new_[2170]_  & \new_[2167]_ ;
  assign \new_[2174]_  = ~A203 & ~A201;
  assign \new_[2177]_  = A300 & A298;
  assign \new_[2178]_  = \new_[2177]_  & \new_[2174]_ ;
  assign \new_[2181]_  = ~A166 & ~A167;
  assign \new_[2184]_  = A201 & A199;
  assign \new_[2185]_  = \new_[2184]_  & \new_[2181]_ ;
  assign \new_[2188]_  = A299 & A298;
  assign \new_[2191]_  = ~A302 & A301;
  assign \new_[2192]_  = \new_[2191]_  & \new_[2188]_ ;
  assign \new_[2195]_  = ~A166 & ~A167;
  assign \new_[2198]_  = A201 & A199;
  assign \new_[2199]_  = \new_[2198]_  & \new_[2195]_ ;
  assign \new_[2202]_  = ~A299 & A298;
  assign \new_[2205]_  = A302 & ~A301;
  assign \new_[2206]_  = \new_[2205]_  & \new_[2202]_ ;
  assign \new_[2209]_  = ~A166 & ~A167;
  assign \new_[2212]_  = A201 & A199;
  assign \new_[2213]_  = \new_[2212]_  & \new_[2209]_ ;
  assign \new_[2216]_  = A299 & ~A298;
  assign \new_[2219]_  = A302 & ~A301;
  assign \new_[2220]_  = \new_[2219]_  & \new_[2216]_ ;
  assign \new_[2223]_  = ~A166 & ~A167;
  assign \new_[2226]_  = A201 & A199;
  assign \new_[2227]_  = \new_[2226]_  & \new_[2223]_ ;
  assign \new_[2230]_  = ~A299 & ~A298;
  assign \new_[2233]_  = ~A302 & A301;
  assign \new_[2234]_  = \new_[2233]_  & \new_[2230]_ ;
  assign \new_[2237]_  = ~A166 & ~A167;
  assign \new_[2240]_  = A201 & A200;
  assign \new_[2241]_  = \new_[2240]_  & \new_[2237]_ ;
  assign \new_[2244]_  = A299 & A298;
  assign \new_[2247]_  = ~A302 & A301;
  assign \new_[2248]_  = \new_[2247]_  & \new_[2244]_ ;
  assign \new_[2251]_  = ~A166 & ~A167;
  assign \new_[2254]_  = A201 & A200;
  assign \new_[2255]_  = \new_[2254]_  & \new_[2251]_ ;
  assign \new_[2258]_  = ~A299 & A298;
  assign \new_[2261]_  = A302 & ~A301;
  assign \new_[2262]_  = \new_[2261]_  & \new_[2258]_ ;
  assign \new_[2265]_  = ~A166 & ~A167;
  assign \new_[2268]_  = A201 & A200;
  assign \new_[2269]_  = \new_[2268]_  & \new_[2265]_ ;
  assign \new_[2272]_  = A299 & ~A298;
  assign \new_[2275]_  = A302 & ~A301;
  assign \new_[2276]_  = \new_[2275]_  & \new_[2272]_ ;
  assign \new_[2279]_  = ~A166 & ~A167;
  assign \new_[2282]_  = A201 & A200;
  assign \new_[2283]_  = \new_[2282]_  & \new_[2279]_ ;
  assign \new_[2286]_  = ~A299 & ~A298;
  assign \new_[2289]_  = ~A302 & A301;
  assign \new_[2290]_  = \new_[2289]_  & \new_[2286]_ ;
  assign \new_[2293]_  = ~A166 & ~A167;
  assign \new_[2296]_  = A200 & A199;
  assign \new_[2297]_  = \new_[2296]_  & \new_[2293]_ ;
  assign \new_[2300]_  = ~A203 & A202;
  assign \new_[2303]_  = A300 & A299;
  assign \new_[2304]_  = \new_[2303]_  & \new_[2300]_ ;
  assign \new_[2307]_  = ~A166 & ~A167;
  assign \new_[2310]_  = A200 & A199;
  assign \new_[2311]_  = \new_[2310]_  & \new_[2307]_ ;
  assign \new_[2314]_  = ~A203 & A202;
  assign \new_[2317]_  = A300 & A298;
  assign \new_[2318]_  = \new_[2317]_  & \new_[2314]_ ;
  assign \new_[2321]_  = ~A166 & ~A167;
  assign \new_[2324]_  = A200 & ~A199;
  assign \new_[2325]_  = \new_[2324]_  & \new_[2321]_ ;
  assign \new_[2328]_  = A203 & ~A202;
  assign \new_[2331]_  = A300 & A299;
  assign \new_[2332]_  = \new_[2331]_  & \new_[2328]_ ;
  assign \new_[2335]_  = ~A166 & ~A167;
  assign \new_[2338]_  = A200 & ~A199;
  assign \new_[2339]_  = \new_[2338]_  & \new_[2335]_ ;
  assign \new_[2342]_  = A203 & ~A202;
  assign \new_[2345]_  = A300 & A298;
  assign \new_[2346]_  = \new_[2345]_  & \new_[2342]_ ;
  assign \new_[2349]_  = ~A166 & ~A167;
  assign \new_[2352]_  = ~A200 & A199;
  assign \new_[2353]_  = \new_[2352]_  & \new_[2349]_ ;
  assign \new_[2356]_  = A203 & ~A202;
  assign \new_[2359]_  = A300 & A299;
  assign \new_[2360]_  = \new_[2359]_  & \new_[2356]_ ;
  assign \new_[2363]_  = ~A166 & ~A167;
  assign \new_[2366]_  = ~A200 & A199;
  assign \new_[2367]_  = \new_[2366]_  & \new_[2363]_ ;
  assign \new_[2370]_  = A203 & ~A202;
  assign \new_[2373]_  = A300 & A298;
  assign \new_[2374]_  = \new_[2373]_  & \new_[2370]_ ;
  assign \new_[2377]_  = ~A166 & ~A167;
  assign \new_[2380]_  = ~A200 & ~A199;
  assign \new_[2381]_  = \new_[2380]_  & \new_[2377]_ ;
  assign \new_[2384]_  = ~A203 & A202;
  assign \new_[2387]_  = A300 & A299;
  assign \new_[2388]_  = \new_[2387]_  & \new_[2384]_ ;
  assign \new_[2391]_  = ~A166 & ~A167;
  assign \new_[2394]_  = ~A200 & ~A199;
  assign \new_[2395]_  = \new_[2394]_  & \new_[2391]_ ;
  assign \new_[2398]_  = ~A203 & A202;
  assign \new_[2401]_  = A300 & A298;
  assign \new_[2402]_  = \new_[2401]_  & \new_[2398]_ ;
  assign \new_[2405]_  = ~A167 & ~A168;
  assign \new_[2408]_  = A201 & A199;
  assign \new_[2409]_  = \new_[2408]_  & \new_[2405]_ ;
  assign \new_[2412]_  = A299 & A298;
  assign \new_[2415]_  = ~A302 & A301;
  assign \new_[2416]_  = \new_[2415]_  & \new_[2412]_ ;
  assign \new_[2419]_  = ~A167 & ~A168;
  assign \new_[2422]_  = A201 & A199;
  assign \new_[2423]_  = \new_[2422]_  & \new_[2419]_ ;
  assign \new_[2426]_  = ~A299 & A298;
  assign \new_[2429]_  = A302 & ~A301;
  assign \new_[2430]_  = \new_[2429]_  & \new_[2426]_ ;
  assign \new_[2433]_  = ~A167 & ~A168;
  assign \new_[2436]_  = A201 & A199;
  assign \new_[2437]_  = \new_[2436]_  & \new_[2433]_ ;
  assign \new_[2440]_  = A299 & ~A298;
  assign \new_[2443]_  = A302 & ~A301;
  assign \new_[2444]_  = \new_[2443]_  & \new_[2440]_ ;
  assign \new_[2447]_  = ~A167 & ~A168;
  assign \new_[2450]_  = A201 & A199;
  assign \new_[2451]_  = \new_[2450]_  & \new_[2447]_ ;
  assign \new_[2454]_  = ~A299 & ~A298;
  assign \new_[2457]_  = ~A302 & A301;
  assign \new_[2458]_  = \new_[2457]_  & \new_[2454]_ ;
  assign \new_[2461]_  = ~A167 & ~A168;
  assign \new_[2464]_  = A201 & A200;
  assign \new_[2465]_  = \new_[2464]_  & \new_[2461]_ ;
  assign \new_[2468]_  = A299 & A298;
  assign \new_[2471]_  = ~A302 & A301;
  assign \new_[2472]_  = \new_[2471]_  & \new_[2468]_ ;
  assign \new_[2475]_  = ~A167 & ~A168;
  assign \new_[2478]_  = A201 & A200;
  assign \new_[2479]_  = \new_[2478]_  & \new_[2475]_ ;
  assign \new_[2482]_  = ~A299 & A298;
  assign \new_[2485]_  = A302 & ~A301;
  assign \new_[2486]_  = \new_[2485]_  & \new_[2482]_ ;
  assign \new_[2489]_  = ~A167 & ~A168;
  assign \new_[2492]_  = A201 & A200;
  assign \new_[2493]_  = \new_[2492]_  & \new_[2489]_ ;
  assign \new_[2496]_  = A299 & ~A298;
  assign \new_[2499]_  = A302 & ~A301;
  assign \new_[2500]_  = \new_[2499]_  & \new_[2496]_ ;
  assign \new_[2503]_  = ~A167 & ~A168;
  assign \new_[2506]_  = A201 & A200;
  assign \new_[2507]_  = \new_[2506]_  & \new_[2503]_ ;
  assign \new_[2510]_  = ~A299 & ~A298;
  assign \new_[2513]_  = ~A302 & A301;
  assign \new_[2514]_  = \new_[2513]_  & \new_[2510]_ ;
  assign \new_[2517]_  = ~A167 & ~A168;
  assign \new_[2520]_  = A200 & A199;
  assign \new_[2521]_  = \new_[2520]_  & \new_[2517]_ ;
  assign \new_[2524]_  = ~A203 & A202;
  assign \new_[2527]_  = A300 & A299;
  assign \new_[2528]_  = \new_[2527]_  & \new_[2524]_ ;
  assign \new_[2531]_  = ~A167 & ~A168;
  assign \new_[2534]_  = A200 & A199;
  assign \new_[2535]_  = \new_[2534]_  & \new_[2531]_ ;
  assign \new_[2538]_  = ~A203 & A202;
  assign \new_[2541]_  = A300 & A298;
  assign \new_[2542]_  = \new_[2541]_  & \new_[2538]_ ;
  assign \new_[2545]_  = ~A167 & ~A168;
  assign \new_[2548]_  = A200 & ~A199;
  assign \new_[2549]_  = \new_[2548]_  & \new_[2545]_ ;
  assign \new_[2552]_  = A203 & ~A202;
  assign \new_[2555]_  = A300 & A299;
  assign \new_[2556]_  = \new_[2555]_  & \new_[2552]_ ;
  assign \new_[2559]_  = ~A167 & ~A168;
  assign \new_[2562]_  = A200 & ~A199;
  assign \new_[2563]_  = \new_[2562]_  & \new_[2559]_ ;
  assign \new_[2566]_  = A203 & ~A202;
  assign \new_[2569]_  = A300 & A298;
  assign \new_[2570]_  = \new_[2569]_  & \new_[2566]_ ;
  assign \new_[2573]_  = ~A167 & ~A168;
  assign \new_[2576]_  = ~A200 & A199;
  assign \new_[2577]_  = \new_[2576]_  & \new_[2573]_ ;
  assign \new_[2580]_  = A203 & ~A202;
  assign \new_[2583]_  = A300 & A299;
  assign \new_[2584]_  = \new_[2583]_  & \new_[2580]_ ;
  assign \new_[2587]_  = ~A167 & ~A168;
  assign \new_[2590]_  = ~A200 & A199;
  assign \new_[2591]_  = \new_[2590]_  & \new_[2587]_ ;
  assign \new_[2594]_  = A203 & ~A202;
  assign \new_[2597]_  = A300 & A298;
  assign \new_[2598]_  = \new_[2597]_  & \new_[2594]_ ;
  assign \new_[2601]_  = ~A167 & ~A168;
  assign \new_[2604]_  = ~A200 & ~A199;
  assign \new_[2605]_  = \new_[2604]_  & \new_[2601]_ ;
  assign \new_[2608]_  = ~A203 & A202;
  assign \new_[2611]_  = A300 & A299;
  assign \new_[2612]_  = \new_[2611]_  & \new_[2608]_ ;
  assign \new_[2615]_  = ~A167 & ~A168;
  assign \new_[2618]_  = ~A200 & ~A199;
  assign \new_[2619]_  = \new_[2618]_  & \new_[2615]_ ;
  assign \new_[2622]_  = ~A203 & A202;
  assign \new_[2625]_  = A300 & A298;
  assign \new_[2626]_  = \new_[2625]_  & \new_[2622]_ ;
  assign \new_[2629]_  = A168 & A170;
  assign \new_[2632]_  = A166 & ~A167;
  assign \new_[2633]_  = \new_[2632]_  & \new_[2629]_ ;
  assign \new_[2636]_  = A233 & A232;
  assign \new_[2639]_  = ~A236 & A235;
  assign \new_[2640]_  = \new_[2639]_  & \new_[2636]_ ;
  assign \new_[2643]_  = A168 & A170;
  assign \new_[2646]_  = A166 & ~A167;
  assign \new_[2647]_  = \new_[2646]_  & \new_[2643]_ ;
  assign \new_[2650]_  = A233 & ~A232;
  assign \new_[2653]_  = A236 & ~A235;
  assign \new_[2654]_  = \new_[2653]_  & \new_[2650]_ ;
  assign \new_[2657]_  = A168 & A170;
  assign \new_[2660]_  = A166 & ~A167;
  assign \new_[2661]_  = \new_[2660]_  & \new_[2657]_ ;
  assign \new_[2664]_  = ~A233 & A232;
  assign \new_[2667]_  = A236 & ~A235;
  assign \new_[2668]_  = \new_[2667]_  & \new_[2664]_ ;
  assign \new_[2671]_  = A168 & A170;
  assign \new_[2674]_  = A166 & ~A167;
  assign \new_[2675]_  = \new_[2674]_  & \new_[2671]_ ;
  assign \new_[2678]_  = ~A233 & ~A232;
  assign \new_[2681]_  = ~A236 & A235;
  assign \new_[2682]_  = \new_[2681]_  & \new_[2678]_ ;
  assign \new_[2685]_  = A168 & A169;
  assign \new_[2688]_  = A166 & ~A167;
  assign \new_[2689]_  = \new_[2688]_  & \new_[2685]_ ;
  assign \new_[2692]_  = A233 & A232;
  assign \new_[2695]_  = ~A236 & A235;
  assign \new_[2696]_  = \new_[2695]_  & \new_[2692]_ ;
  assign \new_[2699]_  = A168 & A169;
  assign \new_[2702]_  = A166 & ~A167;
  assign \new_[2703]_  = \new_[2702]_  & \new_[2699]_ ;
  assign \new_[2706]_  = A233 & ~A232;
  assign \new_[2709]_  = A236 & ~A235;
  assign \new_[2710]_  = \new_[2709]_  & \new_[2706]_ ;
  assign \new_[2713]_  = A168 & A169;
  assign \new_[2716]_  = A166 & ~A167;
  assign \new_[2717]_  = \new_[2716]_  & \new_[2713]_ ;
  assign \new_[2720]_  = ~A233 & A232;
  assign \new_[2723]_  = A236 & ~A235;
  assign \new_[2724]_  = \new_[2723]_  & \new_[2720]_ ;
  assign \new_[2727]_  = A168 & A169;
  assign \new_[2730]_  = A166 & ~A167;
  assign \new_[2731]_  = \new_[2730]_  & \new_[2727]_ ;
  assign \new_[2734]_  = ~A233 & ~A232;
  assign \new_[2737]_  = ~A236 & A235;
  assign \new_[2738]_  = \new_[2737]_  & \new_[2734]_ ;
  assign \new_[2741]_  = ~A166 & A167;
  assign \new_[2744]_  = ~A200 & ~A199;
  assign \new_[2745]_  = \new_[2744]_  & \new_[2741]_ ;
  assign \new_[2748]_  = A298 & ~A202;
  assign \new_[2752]_  = ~A302 & A301;
  assign \new_[2753]_  = A299 & \new_[2752]_ ;
  assign \new_[2754]_  = \new_[2753]_  & \new_[2748]_ ;
  assign \new_[2757]_  = ~A166 & A167;
  assign \new_[2760]_  = ~A200 & ~A199;
  assign \new_[2761]_  = \new_[2760]_  & \new_[2757]_ ;
  assign \new_[2764]_  = A298 & ~A202;
  assign \new_[2768]_  = A302 & ~A301;
  assign \new_[2769]_  = ~A299 & \new_[2768]_ ;
  assign \new_[2770]_  = \new_[2769]_  & \new_[2764]_ ;
  assign \new_[2773]_  = ~A166 & A167;
  assign \new_[2776]_  = ~A200 & ~A199;
  assign \new_[2777]_  = \new_[2776]_  & \new_[2773]_ ;
  assign \new_[2780]_  = ~A298 & ~A202;
  assign \new_[2784]_  = A302 & ~A301;
  assign \new_[2785]_  = A299 & \new_[2784]_ ;
  assign \new_[2786]_  = \new_[2785]_  & \new_[2780]_ ;
  assign \new_[2789]_  = ~A166 & A167;
  assign \new_[2792]_  = ~A200 & ~A199;
  assign \new_[2793]_  = \new_[2792]_  & \new_[2789]_ ;
  assign \new_[2796]_  = ~A298 & ~A202;
  assign \new_[2800]_  = ~A302 & A301;
  assign \new_[2801]_  = ~A299 & \new_[2800]_ ;
  assign \new_[2802]_  = \new_[2801]_  & \new_[2796]_ ;
  assign \new_[2805]_  = ~A166 & A167;
  assign \new_[2808]_  = ~A200 & ~A199;
  assign \new_[2809]_  = \new_[2808]_  & \new_[2805]_ ;
  assign \new_[2812]_  = A298 & A203;
  assign \new_[2816]_  = ~A302 & A301;
  assign \new_[2817]_  = A299 & \new_[2816]_ ;
  assign \new_[2818]_  = \new_[2817]_  & \new_[2812]_ ;
  assign \new_[2821]_  = ~A166 & A167;
  assign \new_[2824]_  = ~A200 & ~A199;
  assign \new_[2825]_  = \new_[2824]_  & \new_[2821]_ ;
  assign \new_[2828]_  = A298 & A203;
  assign \new_[2832]_  = A302 & ~A301;
  assign \new_[2833]_  = ~A299 & \new_[2832]_ ;
  assign \new_[2834]_  = \new_[2833]_  & \new_[2828]_ ;
  assign \new_[2837]_  = ~A166 & A167;
  assign \new_[2840]_  = ~A200 & ~A199;
  assign \new_[2841]_  = \new_[2840]_  & \new_[2837]_ ;
  assign \new_[2844]_  = ~A298 & A203;
  assign \new_[2848]_  = A302 & ~A301;
  assign \new_[2849]_  = A299 & \new_[2848]_ ;
  assign \new_[2850]_  = \new_[2849]_  & \new_[2844]_ ;
  assign \new_[2853]_  = ~A166 & A167;
  assign \new_[2856]_  = ~A200 & ~A199;
  assign \new_[2857]_  = \new_[2856]_  & \new_[2853]_ ;
  assign \new_[2860]_  = ~A298 & A203;
  assign \new_[2864]_  = ~A302 & A301;
  assign \new_[2865]_  = ~A299 & \new_[2864]_ ;
  assign \new_[2866]_  = \new_[2865]_  & \new_[2860]_ ;
  assign \new_[2869]_  = A168 & A170;
  assign \new_[2872]_  = A166 & ~A167;
  assign \new_[2873]_  = \new_[2872]_  & \new_[2869]_ ;
  assign \new_[2876]_  = ~A200 & ~A199;
  assign \new_[2880]_  = A300 & A299;
  assign \new_[2881]_  = ~A202 & \new_[2880]_ ;
  assign \new_[2882]_  = \new_[2881]_  & \new_[2876]_ ;
  assign \new_[2885]_  = A168 & A170;
  assign \new_[2888]_  = A166 & ~A167;
  assign \new_[2889]_  = \new_[2888]_  & \new_[2885]_ ;
  assign \new_[2892]_  = ~A200 & ~A199;
  assign \new_[2896]_  = A300 & A298;
  assign \new_[2897]_  = ~A202 & \new_[2896]_ ;
  assign \new_[2898]_  = \new_[2897]_  & \new_[2892]_ ;
  assign \new_[2901]_  = A168 & A170;
  assign \new_[2904]_  = A166 & ~A167;
  assign \new_[2905]_  = \new_[2904]_  & \new_[2901]_ ;
  assign \new_[2908]_  = ~A200 & ~A199;
  assign \new_[2912]_  = A300 & A299;
  assign \new_[2913]_  = A203 & \new_[2912]_ ;
  assign \new_[2914]_  = \new_[2913]_  & \new_[2908]_ ;
  assign \new_[2917]_  = A168 & A170;
  assign \new_[2920]_  = A166 & ~A167;
  assign \new_[2921]_  = \new_[2920]_  & \new_[2917]_ ;
  assign \new_[2924]_  = ~A200 & ~A199;
  assign \new_[2928]_  = A300 & A298;
  assign \new_[2929]_  = A203 & \new_[2928]_ ;
  assign \new_[2930]_  = \new_[2929]_  & \new_[2924]_ ;
  assign \new_[2933]_  = A168 & A169;
  assign \new_[2936]_  = A166 & ~A167;
  assign \new_[2937]_  = \new_[2936]_  & \new_[2933]_ ;
  assign \new_[2940]_  = ~A200 & ~A199;
  assign \new_[2944]_  = A300 & A299;
  assign \new_[2945]_  = ~A202 & \new_[2944]_ ;
  assign \new_[2946]_  = \new_[2945]_  & \new_[2940]_ ;
  assign \new_[2949]_  = A168 & A169;
  assign \new_[2952]_  = A166 & ~A167;
  assign \new_[2953]_  = \new_[2952]_  & \new_[2949]_ ;
  assign \new_[2956]_  = ~A200 & ~A199;
  assign \new_[2960]_  = A300 & A298;
  assign \new_[2961]_  = ~A202 & \new_[2960]_ ;
  assign \new_[2962]_  = \new_[2961]_  & \new_[2956]_ ;
  assign \new_[2965]_  = A168 & A169;
  assign \new_[2968]_  = A166 & ~A167;
  assign \new_[2969]_  = \new_[2968]_  & \new_[2965]_ ;
  assign \new_[2972]_  = ~A200 & ~A199;
  assign \new_[2976]_  = A300 & A299;
  assign \new_[2977]_  = A203 & \new_[2976]_ ;
  assign \new_[2978]_  = \new_[2977]_  & \new_[2972]_ ;
  assign \new_[2981]_  = A168 & A169;
  assign \new_[2984]_  = A166 & ~A167;
  assign \new_[2985]_  = \new_[2984]_  & \new_[2981]_ ;
  assign \new_[2988]_  = ~A200 & ~A199;
  assign \new_[2992]_  = A300 & A298;
  assign \new_[2993]_  = A203 & \new_[2992]_ ;
  assign \new_[2994]_  = \new_[2993]_  & \new_[2988]_ ;
  assign \new_[2997]_  = ~A169 & ~A170;
  assign \new_[3000]_  = A199 & ~A167;
  assign \new_[3001]_  = \new_[3000]_  & \new_[2997]_ ;
  assign \new_[3004]_  = A298 & A201;
  assign \new_[3008]_  = ~A302 & A301;
  assign \new_[3009]_  = A299 & \new_[3008]_ ;
  assign \new_[3010]_  = \new_[3009]_  & \new_[3004]_ ;
  assign \new_[3013]_  = ~A169 & ~A170;
  assign \new_[3016]_  = A199 & ~A167;
  assign \new_[3017]_  = \new_[3016]_  & \new_[3013]_ ;
  assign \new_[3020]_  = A298 & A201;
  assign \new_[3024]_  = A302 & ~A301;
  assign \new_[3025]_  = ~A299 & \new_[3024]_ ;
  assign \new_[3026]_  = \new_[3025]_  & \new_[3020]_ ;
  assign \new_[3029]_  = ~A169 & ~A170;
  assign \new_[3032]_  = A199 & ~A167;
  assign \new_[3033]_  = \new_[3032]_  & \new_[3029]_ ;
  assign \new_[3036]_  = ~A298 & A201;
  assign \new_[3040]_  = A302 & ~A301;
  assign \new_[3041]_  = A299 & \new_[3040]_ ;
  assign \new_[3042]_  = \new_[3041]_  & \new_[3036]_ ;
  assign \new_[3045]_  = ~A169 & ~A170;
  assign \new_[3048]_  = A199 & ~A167;
  assign \new_[3049]_  = \new_[3048]_  & \new_[3045]_ ;
  assign \new_[3052]_  = ~A298 & A201;
  assign \new_[3056]_  = ~A302 & A301;
  assign \new_[3057]_  = ~A299 & \new_[3056]_ ;
  assign \new_[3058]_  = \new_[3057]_  & \new_[3052]_ ;
  assign \new_[3061]_  = ~A169 & ~A170;
  assign \new_[3064]_  = A200 & ~A167;
  assign \new_[3065]_  = \new_[3064]_  & \new_[3061]_ ;
  assign \new_[3068]_  = A298 & A201;
  assign \new_[3072]_  = ~A302 & A301;
  assign \new_[3073]_  = A299 & \new_[3072]_ ;
  assign \new_[3074]_  = \new_[3073]_  & \new_[3068]_ ;
  assign \new_[3077]_  = ~A169 & ~A170;
  assign \new_[3080]_  = A200 & ~A167;
  assign \new_[3081]_  = \new_[3080]_  & \new_[3077]_ ;
  assign \new_[3084]_  = A298 & A201;
  assign \new_[3088]_  = A302 & ~A301;
  assign \new_[3089]_  = ~A299 & \new_[3088]_ ;
  assign \new_[3090]_  = \new_[3089]_  & \new_[3084]_ ;
  assign \new_[3093]_  = ~A169 & ~A170;
  assign \new_[3096]_  = A200 & ~A167;
  assign \new_[3097]_  = \new_[3096]_  & \new_[3093]_ ;
  assign \new_[3100]_  = ~A298 & A201;
  assign \new_[3104]_  = A302 & ~A301;
  assign \new_[3105]_  = A299 & \new_[3104]_ ;
  assign \new_[3106]_  = \new_[3105]_  & \new_[3100]_ ;
  assign \new_[3109]_  = ~A169 & ~A170;
  assign \new_[3112]_  = A200 & ~A167;
  assign \new_[3113]_  = \new_[3112]_  & \new_[3109]_ ;
  assign \new_[3116]_  = ~A298 & A201;
  assign \new_[3120]_  = ~A302 & A301;
  assign \new_[3121]_  = ~A299 & \new_[3120]_ ;
  assign \new_[3122]_  = \new_[3121]_  & \new_[3116]_ ;
  assign \new_[3125]_  = ~A169 & ~A170;
  assign \new_[3128]_  = A199 & ~A167;
  assign \new_[3129]_  = \new_[3128]_  & \new_[3125]_ ;
  assign \new_[3132]_  = A202 & A200;
  assign \new_[3136]_  = A300 & A299;
  assign \new_[3137]_  = ~A203 & \new_[3136]_ ;
  assign \new_[3138]_  = \new_[3137]_  & \new_[3132]_ ;
  assign \new_[3141]_  = ~A169 & ~A170;
  assign \new_[3144]_  = A199 & ~A167;
  assign \new_[3145]_  = \new_[3144]_  & \new_[3141]_ ;
  assign \new_[3148]_  = A202 & A200;
  assign \new_[3152]_  = A300 & A298;
  assign \new_[3153]_  = ~A203 & \new_[3152]_ ;
  assign \new_[3154]_  = \new_[3153]_  & \new_[3148]_ ;
  assign \new_[3157]_  = ~A169 & ~A170;
  assign \new_[3160]_  = ~A199 & ~A167;
  assign \new_[3161]_  = \new_[3160]_  & \new_[3157]_ ;
  assign \new_[3164]_  = ~A202 & A200;
  assign \new_[3168]_  = A300 & A299;
  assign \new_[3169]_  = A203 & \new_[3168]_ ;
  assign \new_[3170]_  = \new_[3169]_  & \new_[3164]_ ;
  assign \new_[3173]_  = ~A169 & ~A170;
  assign \new_[3176]_  = ~A199 & ~A167;
  assign \new_[3177]_  = \new_[3176]_  & \new_[3173]_ ;
  assign \new_[3180]_  = ~A202 & A200;
  assign \new_[3184]_  = A300 & A298;
  assign \new_[3185]_  = A203 & \new_[3184]_ ;
  assign \new_[3186]_  = \new_[3185]_  & \new_[3180]_ ;
  assign \new_[3189]_  = ~A169 & ~A170;
  assign \new_[3192]_  = A199 & ~A167;
  assign \new_[3193]_  = \new_[3192]_  & \new_[3189]_ ;
  assign \new_[3196]_  = ~A202 & ~A200;
  assign \new_[3200]_  = A300 & A299;
  assign \new_[3201]_  = A203 & \new_[3200]_ ;
  assign \new_[3202]_  = \new_[3201]_  & \new_[3196]_ ;
  assign \new_[3205]_  = ~A169 & ~A170;
  assign \new_[3208]_  = A199 & ~A167;
  assign \new_[3209]_  = \new_[3208]_  & \new_[3205]_ ;
  assign \new_[3212]_  = ~A202 & ~A200;
  assign \new_[3216]_  = A300 & A298;
  assign \new_[3217]_  = A203 & \new_[3216]_ ;
  assign \new_[3218]_  = \new_[3217]_  & \new_[3212]_ ;
  assign \new_[3221]_  = ~A169 & ~A170;
  assign \new_[3224]_  = ~A199 & ~A167;
  assign \new_[3225]_  = \new_[3224]_  & \new_[3221]_ ;
  assign \new_[3228]_  = A202 & ~A200;
  assign \new_[3232]_  = A300 & A299;
  assign \new_[3233]_  = ~A203 & \new_[3232]_ ;
  assign \new_[3234]_  = \new_[3233]_  & \new_[3228]_ ;
  assign \new_[3237]_  = ~A169 & ~A170;
  assign \new_[3240]_  = ~A199 & ~A167;
  assign \new_[3241]_  = \new_[3240]_  & \new_[3237]_ ;
  assign \new_[3244]_  = A202 & ~A200;
  assign \new_[3248]_  = A300 & A298;
  assign \new_[3249]_  = ~A203 & \new_[3248]_ ;
  assign \new_[3250]_  = \new_[3249]_  & \new_[3244]_ ;
  assign \new_[3253]_  = A166 & A167;
  assign \new_[3257]_  = A202 & A200;
  assign \new_[3258]_  = A199 & \new_[3257]_ ;
  assign \new_[3259]_  = \new_[3258]_  & \new_[3253]_ ;
  assign \new_[3262]_  = A298 & ~A203;
  assign \new_[3266]_  = ~A302 & A301;
  assign \new_[3267]_  = A299 & \new_[3266]_ ;
  assign \new_[3268]_  = \new_[3267]_  & \new_[3262]_ ;
  assign \new_[3271]_  = A166 & A167;
  assign \new_[3275]_  = A202 & A200;
  assign \new_[3276]_  = A199 & \new_[3275]_ ;
  assign \new_[3277]_  = \new_[3276]_  & \new_[3271]_ ;
  assign \new_[3280]_  = A298 & ~A203;
  assign \new_[3284]_  = A302 & ~A301;
  assign \new_[3285]_  = ~A299 & \new_[3284]_ ;
  assign \new_[3286]_  = \new_[3285]_  & \new_[3280]_ ;
  assign \new_[3289]_  = A166 & A167;
  assign \new_[3293]_  = A202 & A200;
  assign \new_[3294]_  = A199 & \new_[3293]_ ;
  assign \new_[3295]_  = \new_[3294]_  & \new_[3289]_ ;
  assign \new_[3298]_  = ~A298 & ~A203;
  assign \new_[3302]_  = A302 & ~A301;
  assign \new_[3303]_  = A299 & \new_[3302]_ ;
  assign \new_[3304]_  = \new_[3303]_  & \new_[3298]_ ;
  assign \new_[3307]_  = A166 & A167;
  assign \new_[3311]_  = A202 & A200;
  assign \new_[3312]_  = A199 & \new_[3311]_ ;
  assign \new_[3313]_  = \new_[3312]_  & \new_[3307]_ ;
  assign \new_[3316]_  = ~A298 & ~A203;
  assign \new_[3320]_  = ~A302 & A301;
  assign \new_[3321]_  = ~A299 & \new_[3320]_ ;
  assign \new_[3322]_  = \new_[3321]_  & \new_[3316]_ ;
  assign \new_[3325]_  = A166 & A167;
  assign \new_[3329]_  = ~A202 & A200;
  assign \new_[3330]_  = ~A199 & \new_[3329]_ ;
  assign \new_[3331]_  = \new_[3330]_  & \new_[3325]_ ;
  assign \new_[3334]_  = A298 & A203;
  assign \new_[3338]_  = ~A302 & A301;
  assign \new_[3339]_  = A299 & \new_[3338]_ ;
  assign \new_[3340]_  = \new_[3339]_  & \new_[3334]_ ;
  assign \new_[3343]_  = A166 & A167;
  assign \new_[3347]_  = ~A202 & A200;
  assign \new_[3348]_  = ~A199 & \new_[3347]_ ;
  assign \new_[3349]_  = \new_[3348]_  & \new_[3343]_ ;
  assign \new_[3352]_  = A298 & A203;
  assign \new_[3356]_  = A302 & ~A301;
  assign \new_[3357]_  = ~A299 & \new_[3356]_ ;
  assign \new_[3358]_  = \new_[3357]_  & \new_[3352]_ ;
  assign \new_[3361]_  = A166 & A167;
  assign \new_[3365]_  = ~A202 & A200;
  assign \new_[3366]_  = ~A199 & \new_[3365]_ ;
  assign \new_[3367]_  = \new_[3366]_  & \new_[3361]_ ;
  assign \new_[3370]_  = ~A298 & A203;
  assign \new_[3374]_  = A302 & ~A301;
  assign \new_[3375]_  = A299 & \new_[3374]_ ;
  assign \new_[3376]_  = \new_[3375]_  & \new_[3370]_ ;
  assign \new_[3379]_  = A166 & A167;
  assign \new_[3383]_  = ~A202 & A200;
  assign \new_[3384]_  = ~A199 & \new_[3383]_ ;
  assign \new_[3385]_  = \new_[3384]_  & \new_[3379]_ ;
  assign \new_[3388]_  = ~A298 & A203;
  assign \new_[3392]_  = ~A302 & A301;
  assign \new_[3393]_  = ~A299 & \new_[3392]_ ;
  assign \new_[3394]_  = \new_[3393]_  & \new_[3388]_ ;
  assign \new_[3397]_  = A166 & A167;
  assign \new_[3401]_  = ~A202 & ~A200;
  assign \new_[3402]_  = A199 & \new_[3401]_ ;
  assign \new_[3403]_  = \new_[3402]_  & \new_[3397]_ ;
  assign \new_[3406]_  = A298 & A203;
  assign \new_[3410]_  = ~A302 & A301;
  assign \new_[3411]_  = A299 & \new_[3410]_ ;
  assign \new_[3412]_  = \new_[3411]_  & \new_[3406]_ ;
  assign \new_[3415]_  = A166 & A167;
  assign \new_[3419]_  = ~A202 & ~A200;
  assign \new_[3420]_  = A199 & \new_[3419]_ ;
  assign \new_[3421]_  = \new_[3420]_  & \new_[3415]_ ;
  assign \new_[3424]_  = A298 & A203;
  assign \new_[3428]_  = A302 & ~A301;
  assign \new_[3429]_  = ~A299 & \new_[3428]_ ;
  assign \new_[3430]_  = \new_[3429]_  & \new_[3424]_ ;
  assign \new_[3433]_  = A166 & A167;
  assign \new_[3437]_  = ~A202 & ~A200;
  assign \new_[3438]_  = A199 & \new_[3437]_ ;
  assign \new_[3439]_  = \new_[3438]_  & \new_[3433]_ ;
  assign \new_[3442]_  = ~A298 & A203;
  assign \new_[3446]_  = A302 & ~A301;
  assign \new_[3447]_  = A299 & \new_[3446]_ ;
  assign \new_[3448]_  = \new_[3447]_  & \new_[3442]_ ;
  assign \new_[3451]_  = A166 & A167;
  assign \new_[3455]_  = ~A202 & ~A200;
  assign \new_[3456]_  = A199 & \new_[3455]_ ;
  assign \new_[3457]_  = \new_[3456]_  & \new_[3451]_ ;
  assign \new_[3460]_  = ~A298 & A203;
  assign \new_[3464]_  = ~A302 & A301;
  assign \new_[3465]_  = ~A299 & \new_[3464]_ ;
  assign \new_[3466]_  = \new_[3465]_  & \new_[3460]_ ;
  assign \new_[3469]_  = A166 & A167;
  assign \new_[3473]_  = A202 & ~A200;
  assign \new_[3474]_  = ~A199 & \new_[3473]_ ;
  assign \new_[3475]_  = \new_[3474]_  & \new_[3469]_ ;
  assign \new_[3478]_  = A298 & ~A203;
  assign \new_[3482]_  = ~A302 & A301;
  assign \new_[3483]_  = A299 & \new_[3482]_ ;
  assign \new_[3484]_  = \new_[3483]_  & \new_[3478]_ ;
  assign \new_[3487]_  = A166 & A167;
  assign \new_[3491]_  = A202 & ~A200;
  assign \new_[3492]_  = ~A199 & \new_[3491]_ ;
  assign \new_[3493]_  = \new_[3492]_  & \new_[3487]_ ;
  assign \new_[3496]_  = A298 & ~A203;
  assign \new_[3500]_  = A302 & ~A301;
  assign \new_[3501]_  = ~A299 & \new_[3500]_ ;
  assign \new_[3502]_  = \new_[3501]_  & \new_[3496]_ ;
  assign \new_[3505]_  = A166 & A167;
  assign \new_[3509]_  = A202 & ~A200;
  assign \new_[3510]_  = ~A199 & \new_[3509]_ ;
  assign \new_[3511]_  = \new_[3510]_  & \new_[3505]_ ;
  assign \new_[3514]_  = ~A298 & ~A203;
  assign \new_[3518]_  = A302 & ~A301;
  assign \new_[3519]_  = A299 & \new_[3518]_ ;
  assign \new_[3520]_  = \new_[3519]_  & \new_[3514]_ ;
  assign \new_[3523]_  = A166 & A167;
  assign \new_[3527]_  = A202 & ~A200;
  assign \new_[3528]_  = ~A199 & \new_[3527]_ ;
  assign \new_[3529]_  = \new_[3528]_  & \new_[3523]_ ;
  assign \new_[3532]_  = ~A298 & ~A203;
  assign \new_[3536]_  = ~A302 & A301;
  assign \new_[3537]_  = ~A299 & \new_[3536]_ ;
  assign \new_[3538]_  = \new_[3537]_  & \new_[3532]_ ;
  assign \new_[3541]_  = ~A166 & A167;
  assign \new_[3545]_  = ~A201 & A200;
  assign \new_[3546]_  = A199 & \new_[3545]_ ;
  assign \new_[3547]_  = \new_[3546]_  & \new_[3541]_ ;
  assign \new_[3550]_  = A298 & ~A202;
  assign \new_[3554]_  = ~A302 & A301;
  assign \new_[3555]_  = A299 & \new_[3554]_ ;
  assign \new_[3556]_  = \new_[3555]_  & \new_[3550]_ ;
  assign \new_[3559]_  = ~A166 & A167;
  assign \new_[3563]_  = ~A201 & A200;
  assign \new_[3564]_  = A199 & \new_[3563]_ ;
  assign \new_[3565]_  = \new_[3564]_  & \new_[3559]_ ;
  assign \new_[3568]_  = A298 & ~A202;
  assign \new_[3572]_  = A302 & ~A301;
  assign \new_[3573]_  = ~A299 & \new_[3572]_ ;
  assign \new_[3574]_  = \new_[3573]_  & \new_[3568]_ ;
  assign \new_[3577]_  = ~A166 & A167;
  assign \new_[3581]_  = ~A201 & A200;
  assign \new_[3582]_  = A199 & \new_[3581]_ ;
  assign \new_[3583]_  = \new_[3582]_  & \new_[3577]_ ;
  assign \new_[3586]_  = ~A298 & ~A202;
  assign \new_[3590]_  = A302 & ~A301;
  assign \new_[3591]_  = A299 & \new_[3590]_ ;
  assign \new_[3592]_  = \new_[3591]_  & \new_[3586]_ ;
  assign \new_[3595]_  = ~A166 & A167;
  assign \new_[3599]_  = ~A201 & A200;
  assign \new_[3600]_  = A199 & \new_[3599]_ ;
  assign \new_[3601]_  = \new_[3600]_  & \new_[3595]_ ;
  assign \new_[3604]_  = ~A298 & ~A202;
  assign \new_[3608]_  = ~A302 & A301;
  assign \new_[3609]_  = ~A299 & \new_[3608]_ ;
  assign \new_[3610]_  = \new_[3609]_  & \new_[3604]_ ;
  assign \new_[3613]_  = ~A166 & A167;
  assign \new_[3617]_  = ~A201 & A200;
  assign \new_[3618]_  = A199 & \new_[3617]_ ;
  assign \new_[3619]_  = \new_[3618]_  & \new_[3613]_ ;
  assign \new_[3622]_  = A298 & A203;
  assign \new_[3626]_  = ~A302 & A301;
  assign \new_[3627]_  = A299 & \new_[3626]_ ;
  assign \new_[3628]_  = \new_[3627]_  & \new_[3622]_ ;
  assign \new_[3631]_  = ~A166 & A167;
  assign \new_[3635]_  = ~A201 & A200;
  assign \new_[3636]_  = A199 & \new_[3635]_ ;
  assign \new_[3637]_  = \new_[3636]_  & \new_[3631]_ ;
  assign \new_[3640]_  = A298 & A203;
  assign \new_[3644]_  = A302 & ~A301;
  assign \new_[3645]_  = ~A299 & \new_[3644]_ ;
  assign \new_[3646]_  = \new_[3645]_  & \new_[3640]_ ;
  assign \new_[3649]_  = ~A166 & A167;
  assign \new_[3653]_  = ~A201 & A200;
  assign \new_[3654]_  = A199 & \new_[3653]_ ;
  assign \new_[3655]_  = \new_[3654]_  & \new_[3649]_ ;
  assign \new_[3658]_  = ~A298 & A203;
  assign \new_[3662]_  = A302 & ~A301;
  assign \new_[3663]_  = A299 & \new_[3662]_ ;
  assign \new_[3664]_  = \new_[3663]_  & \new_[3658]_ ;
  assign \new_[3667]_  = ~A166 & A167;
  assign \new_[3671]_  = ~A201 & A200;
  assign \new_[3672]_  = A199 & \new_[3671]_ ;
  assign \new_[3673]_  = \new_[3672]_  & \new_[3667]_ ;
  assign \new_[3676]_  = ~A298 & A203;
  assign \new_[3680]_  = ~A302 & A301;
  assign \new_[3681]_  = ~A299 & \new_[3680]_ ;
  assign \new_[3682]_  = \new_[3681]_  & \new_[3676]_ ;
  assign \new_[3685]_  = ~A166 & A167;
  assign \new_[3689]_  = ~A201 & A200;
  assign \new_[3690]_  = ~A199 & \new_[3689]_ ;
  assign \new_[3691]_  = \new_[3690]_  & \new_[3685]_ ;
  assign \new_[3694]_  = A298 & A202;
  assign \new_[3698]_  = ~A302 & A301;
  assign \new_[3699]_  = A299 & \new_[3698]_ ;
  assign \new_[3700]_  = \new_[3699]_  & \new_[3694]_ ;
  assign \new_[3703]_  = ~A166 & A167;
  assign \new_[3707]_  = ~A201 & A200;
  assign \new_[3708]_  = ~A199 & \new_[3707]_ ;
  assign \new_[3709]_  = \new_[3708]_  & \new_[3703]_ ;
  assign \new_[3712]_  = A298 & A202;
  assign \new_[3716]_  = A302 & ~A301;
  assign \new_[3717]_  = ~A299 & \new_[3716]_ ;
  assign \new_[3718]_  = \new_[3717]_  & \new_[3712]_ ;
  assign \new_[3721]_  = ~A166 & A167;
  assign \new_[3725]_  = ~A201 & A200;
  assign \new_[3726]_  = ~A199 & \new_[3725]_ ;
  assign \new_[3727]_  = \new_[3726]_  & \new_[3721]_ ;
  assign \new_[3730]_  = ~A298 & A202;
  assign \new_[3734]_  = A302 & ~A301;
  assign \new_[3735]_  = A299 & \new_[3734]_ ;
  assign \new_[3736]_  = \new_[3735]_  & \new_[3730]_ ;
  assign \new_[3739]_  = ~A166 & A167;
  assign \new_[3743]_  = ~A201 & A200;
  assign \new_[3744]_  = ~A199 & \new_[3743]_ ;
  assign \new_[3745]_  = \new_[3744]_  & \new_[3739]_ ;
  assign \new_[3748]_  = ~A298 & A202;
  assign \new_[3752]_  = ~A302 & A301;
  assign \new_[3753]_  = ~A299 & \new_[3752]_ ;
  assign \new_[3754]_  = \new_[3753]_  & \new_[3748]_ ;
  assign \new_[3757]_  = ~A166 & A167;
  assign \new_[3761]_  = ~A201 & A200;
  assign \new_[3762]_  = ~A199 & \new_[3761]_ ;
  assign \new_[3763]_  = \new_[3762]_  & \new_[3757]_ ;
  assign \new_[3766]_  = A298 & ~A203;
  assign \new_[3770]_  = ~A302 & A301;
  assign \new_[3771]_  = A299 & \new_[3770]_ ;
  assign \new_[3772]_  = \new_[3771]_  & \new_[3766]_ ;
  assign \new_[3775]_  = ~A166 & A167;
  assign \new_[3779]_  = ~A201 & A200;
  assign \new_[3780]_  = ~A199 & \new_[3779]_ ;
  assign \new_[3781]_  = \new_[3780]_  & \new_[3775]_ ;
  assign \new_[3784]_  = A298 & ~A203;
  assign \new_[3788]_  = A302 & ~A301;
  assign \new_[3789]_  = ~A299 & \new_[3788]_ ;
  assign \new_[3790]_  = \new_[3789]_  & \new_[3784]_ ;
  assign \new_[3793]_  = ~A166 & A167;
  assign \new_[3797]_  = ~A201 & A200;
  assign \new_[3798]_  = ~A199 & \new_[3797]_ ;
  assign \new_[3799]_  = \new_[3798]_  & \new_[3793]_ ;
  assign \new_[3802]_  = ~A298 & ~A203;
  assign \new_[3806]_  = A302 & ~A301;
  assign \new_[3807]_  = A299 & \new_[3806]_ ;
  assign \new_[3808]_  = \new_[3807]_  & \new_[3802]_ ;
  assign \new_[3811]_  = ~A166 & A167;
  assign \new_[3815]_  = ~A201 & A200;
  assign \new_[3816]_  = ~A199 & \new_[3815]_ ;
  assign \new_[3817]_  = \new_[3816]_  & \new_[3811]_ ;
  assign \new_[3820]_  = ~A298 & ~A203;
  assign \new_[3824]_  = ~A302 & A301;
  assign \new_[3825]_  = ~A299 & \new_[3824]_ ;
  assign \new_[3826]_  = \new_[3825]_  & \new_[3820]_ ;
  assign \new_[3829]_  = ~A166 & A167;
  assign \new_[3833]_  = ~A201 & ~A200;
  assign \new_[3834]_  = A199 & \new_[3833]_ ;
  assign \new_[3835]_  = \new_[3834]_  & \new_[3829]_ ;
  assign \new_[3838]_  = A298 & A202;
  assign \new_[3842]_  = ~A302 & A301;
  assign \new_[3843]_  = A299 & \new_[3842]_ ;
  assign \new_[3844]_  = \new_[3843]_  & \new_[3838]_ ;
  assign \new_[3847]_  = ~A166 & A167;
  assign \new_[3851]_  = ~A201 & ~A200;
  assign \new_[3852]_  = A199 & \new_[3851]_ ;
  assign \new_[3853]_  = \new_[3852]_  & \new_[3847]_ ;
  assign \new_[3856]_  = A298 & A202;
  assign \new_[3860]_  = A302 & ~A301;
  assign \new_[3861]_  = ~A299 & \new_[3860]_ ;
  assign \new_[3862]_  = \new_[3861]_  & \new_[3856]_ ;
  assign \new_[3865]_  = ~A166 & A167;
  assign \new_[3869]_  = ~A201 & ~A200;
  assign \new_[3870]_  = A199 & \new_[3869]_ ;
  assign \new_[3871]_  = \new_[3870]_  & \new_[3865]_ ;
  assign \new_[3874]_  = ~A298 & A202;
  assign \new_[3878]_  = A302 & ~A301;
  assign \new_[3879]_  = A299 & \new_[3878]_ ;
  assign \new_[3880]_  = \new_[3879]_  & \new_[3874]_ ;
  assign \new_[3883]_  = ~A166 & A167;
  assign \new_[3887]_  = ~A201 & ~A200;
  assign \new_[3888]_  = A199 & \new_[3887]_ ;
  assign \new_[3889]_  = \new_[3888]_  & \new_[3883]_ ;
  assign \new_[3892]_  = ~A298 & A202;
  assign \new_[3896]_  = ~A302 & A301;
  assign \new_[3897]_  = ~A299 & \new_[3896]_ ;
  assign \new_[3898]_  = \new_[3897]_  & \new_[3892]_ ;
  assign \new_[3901]_  = ~A166 & A167;
  assign \new_[3905]_  = ~A201 & ~A200;
  assign \new_[3906]_  = A199 & \new_[3905]_ ;
  assign \new_[3907]_  = \new_[3906]_  & \new_[3901]_ ;
  assign \new_[3910]_  = A298 & ~A203;
  assign \new_[3914]_  = ~A302 & A301;
  assign \new_[3915]_  = A299 & \new_[3914]_ ;
  assign \new_[3916]_  = \new_[3915]_  & \new_[3910]_ ;
  assign \new_[3919]_  = ~A166 & A167;
  assign \new_[3923]_  = ~A201 & ~A200;
  assign \new_[3924]_  = A199 & \new_[3923]_ ;
  assign \new_[3925]_  = \new_[3924]_  & \new_[3919]_ ;
  assign \new_[3928]_  = A298 & ~A203;
  assign \new_[3932]_  = A302 & ~A301;
  assign \new_[3933]_  = ~A299 & \new_[3932]_ ;
  assign \new_[3934]_  = \new_[3933]_  & \new_[3928]_ ;
  assign \new_[3937]_  = ~A166 & A167;
  assign \new_[3941]_  = ~A201 & ~A200;
  assign \new_[3942]_  = A199 & \new_[3941]_ ;
  assign \new_[3943]_  = \new_[3942]_  & \new_[3937]_ ;
  assign \new_[3946]_  = ~A298 & ~A203;
  assign \new_[3950]_  = A302 & ~A301;
  assign \new_[3951]_  = A299 & \new_[3950]_ ;
  assign \new_[3952]_  = \new_[3951]_  & \new_[3946]_ ;
  assign \new_[3955]_  = ~A166 & A167;
  assign \new_[3959]_  = ~A201 & ~A200;
  assign \new_[3960]_  = A199 & \new_[3959]_ ;
  assign \new_[3961]_  = \new_[3960]_  & \new_[3955]_ ;
  assign \new_[3964]_  = ~A298 & ~A203;
  assign \new_[3968]_  = ~A302 & A301;
  assign \new_[3969]_  = ~A299 & \new_[3968]_ ;
  assign \new_[3970]_  = \new_[3969]_  & \new_[3964]_ ;
  assign \new_[3973]_  = ~A166 & ~A167;
  assign \new_[3977]_  = A202 & A200;
  assign \new_[3978]_  = A199 & \new_[3977]_ ;
  assign \new_[3979]_  = \new_[3978]_  & \new_[3973]_ ;
  assign \new_[3982]_  = A298 & ~A203;
  assign \new_[3986]_  = ~A302 & A301;
  assign \new_[3987]_  = A299 & \new_[3986]_ ;
  assign \new_[3988]_  = \new_[3987]_  & \new_[3982]_ ;
  assign \new_[3991]_  = ~A166 & ~A167;
  assign \new_[3995]_  = A202 & A200;
  assign \new_[3996]_  = A199 & \new_[3995]_ ;
  assign \new_[3997]_  = \new_[3996]_  & \new_[3991]_ ;
  assign \new_[4000]_  = A298 & ~A203;
  assign \new_[4004]_  = A302 & ~A301;
  assign \new_[4005]_  = ~A299 & \new_[4004]_ ;
  assign \new_[4006]_  = \new_[4005]_  & \new_[4000]_ ;
  assign \new_[4009]_  = ~A166 & ~A167;
  assign \new_[4013]_  = A202 & A200;
  assign \new_[4014]_  = A199 & \new_[4013]_ ;
  assign \new_[4015]_  = \new_[4014]_  & \new_[4009]_ ;
  assign \new_[4018]_  = ~A298 & ~A203;
  assign \new_[4022]_  = A302 & ~A301;
  assign \new_[4023]_  = A299 & \new_[4022]_ ;
  assign \new_[4024]_  = \new_[4023]_  & \new_[4018]_ ;
  assign \new_[4027]_  = ~A166 & ~A167;
  assign \new_[4031]_  = A202 & A200;
  assign \new_[4032]_  = A199 & \new_[4031]_ ;
  assign \new_[4033]_  = \new_[4032]_  & \new_[4027]_ ;
  assign \new_[4036]_  = ~A298 & ~A203;
  assign \new_[4040]_  = ~A302 & A301;
  assign \new_[4041]_  = ~A299 & \new_[4040]_ ;
  assign \new_[4042]_  = \new_[4041]_  & \new_[4036]_ ;
  assign \new_[4045]_  = ~A166 & ~A167;
  assign \new_[4049]_  = ~A202 & A200;
  assign \new_[4050]_  = ~A199 & \new_[4049]_ ;
  assign \new_[4051]_  = \new_[4050]_  & \new_[4045]_ ;
  assign \new_[4054]_  = A298 & A203;
  assign \new_[4058]_  = ~A302 & A301;
  assign \new_[4059]_  = A299 & \new_[4058]_ ;
  assign \new_[4060]_  = \new_[4059]_  & \new_[4054]_ ;
  assign \new_[4063]_  = ~A166 & ~A167;
  assign \new_[4067]_  = ~A202 & A200;
  assign \new_[4068]_  = ~A199 & \new_[4067]_ ;
  assign \new_[4069]_  = \new_[4068]_  & \new_[4063]_ ;
  assign \new_[4072]_  = A298 & A203;
  assign \new_[4076]_  = A302 & ~A301;
  assign \new_[4077]_  = ~A299 & \new_[4076]_ ;
  assign \new_[4078]_  = \new_[4077]_  & \new_[4072]_ ;
  assign \new_[4081]_  = ~A166 & ~A167;
  assign \new_[4085]_  = ~A202 & A200;
  assign \new_[4086]_  = ~A199 & \new_[4085]_ ;
  assign \new_[4087]_  = \new_[4086]_  & \new_[4081]_ ;
  assign \new_[4090]_  = ~A298 & A203;
  assign \new_[4094]_  = A302 & ~A301;
  assign \new_[4095]_  = A299 & \new_[4094]_ ;
  assign \new_[4096]_  = \new_[4095]_  & \new_[4090]_ ;
  assign \new_[4099]_  = ~A166 & ~A167;
  assign \new_[4103]_  = ~A202 & A200;
  assign \new_[4104]_  = ~A199 & \new_[4103]_ ;
  assign \new_[4105]_  = \new_[4104]_  & \new_[4099]_ ;
  assign \new_[4108]_  = ~A298 & A203;
  assign \new_[4112]_  = ~A302 & A301;
  assign \new_[4113]_  = ~A299 & \new_[4112]_ ;
  assign \new_[4114]_  = \new_[4113]_  & \new_[4108]_ ;
  assign \new_[4117]_  = ~A166 & ~A167;
  assign \new_[4121]_  = ~A202 & ~A200;
  assign \new_[4122]_  = A199 & \new_[4121]_ ;
  assign \new_[4123]_  = \new_[4122]_  & \new_[4117]_ ;
  assign \new_[4126]_  = A298 & A203;
  assign \new_[4130]_  = ~A302 & A301;
  assign \new_[4131]_  = A299 & \new_[4130]_ ;
  assign \new_[4132]_  = \new_[4131]_  & \new_[4126]_ ;
  assign \new_[4135]_  = ~A166 & ~A167;
  assign \new_[4139]_  = ~A202 & ~A200;
  assign \new_[4140]_  = A199 & \new_[4139]_ ;
  assign \new_[4141]_  = \new_[4140]_  & \new_[4135]_ ;
  assign \new_[4144]_  = A298 & A203;
  assign \new_[4148]_  = A302 & ~A301;
  assign \new_[4149]_  = ~A299 & \new_[4148]_ ;
  assign \new_[4150]_  = \new_[4149]_  & \new_[4144]_ ;
  assign \new_[4153]_  = ~A166 & ~A167;
  assign \new_[4157]_  = ~A202 & ~A200;
  assign \new_[4158]_  = A199 & \new_[4157]_ ;
  assign \new_[4159]_  = \new_[4158]_  & \new_[4153]_ ;
  assign \new_[4162]_  = ~A298 & A203;
  assign \new_[4166]_  = A302 & ~A301;
  assign \new_[4167]_  = A299 & \new_[4166]_ ;
  assign \new_[4168]_  = \new_[4167]_  & \new_[4162]_ ;
  assign \new_[4171]_  = ~A166 & ~A167;
  assign \new_[4175]_  = ~A202 & ~A200;
  assign \new_[4176]_  = A199 & \new_[4175]_ ;
  assign \new_[4177]_  = \new_[4176]_  & \new_[4171]_ ;
  assign \new_[4180]_  = ~A298 & A203;
  assign \new_[4184]_  = ~A302 & A301;
  assign \new_[4185]_  = ~A299 & \new_[4184]_ ;
  assign \new_[4186]_  = \new_[4185]_  & \new_[4180]_ ;
  assign \new_[4189]_  = ~A166 & ~A167;
  assign \new_[4193]_  = A202 & ~A200;
  assign \new_[4194]_  = ~A199 & \new_[4193]_ ;
  assign \new_[4195]_  = \new_[4194]_  & \new_[4189]_ ;
  assign \new_[4198]_  = A298 & ~A203;
  assign \new_[4202]_  = ~A302 & A301;
  assign \new_[4203]_  = A299 & \new_[4202]_ ;
  assign \new_[4204]_  = \new_[4203]_  & \new_[4198]_ ;
  assign \new_[4207]_  = ~A166 & ~A167;
  assign \new_[4211]_  = A202 & ~A200;
  assign \new_[4212]_  = ~A199 & \new_[4211]_ ;
  assign \new_[4213]_  = \new_[4212]_  & \new_[4207]_ ;
  assign \new_[4216]_  = A298 & ~A203;
  assign \new_[4220]_  = A302 & ~A301;
  assign \new_[4221]_  = ~A299 & \new_[4220]_ ;
  assign \new_[4222]_  = \new_[4221]_  & \new_[4216]_ ;
  assign \new_[4225]_  = ~A166 & ~A167;
  assign \new_[4229]_  = A202 & ~A200;
  assign \new_[4230]_  = ~A199 & \new_[4229]_ ;
  assign \new_[4231]_  = \new_[4230]_  & \new_[4225]_ ;
  assign \new_[4234]_  = ~A298 & ~A203;
  assign \new_[4238]_  = A302 & ~A301;
  assign \new_[4239]_  = A299 & \new_[4238]_ ;
  assign \new_[4240]_  = \new_[4239]_  & \new_[4234]_ ;
  assign \new_[4243]_  = ~A166 & ~A167;
  assign \new_[4247]_  = A202 & ~A200;
  assign \new_[4248]_  = ~A199 & \new_[4247]_ ;
  assign \new_[4249]_  = \new_[4248]_  & \new_[4243]_ ;
  assign \new_[4252]_  = ~A298 & ~A203;
  assign \new_[4256]_  = ~A302 & A301;
  assign \new_[4257]_  = ~A299 & \new_[4256]_ ;
  assign \new_[4258]_  = \new_[4257]_  & \new_[4252]_ ;
  assign \new_[4261]_  = ~A167 & ~A168;
  assign \new_[4265]_  = A202 & A200;
  assign \new_[4266]_  = A199 & \new_[4265]_ ;
  assign \new_[4267]_  = \new_[4266]_  & \new_[4261]_ ;
  assign \new_[4270]_  = A298 & ~A203;
  assign \new_[4274]_  = ~A302 & A301;
  assign \new_[4275]_  = A299 & \new_[4274]_ ;
  assign \new_[4276]_  = \new_[4275]_  & \new_[4270]_ ;
  assign \new_[4279]_  = ~A167 & ~A168;
  assign \new_[4283]_  = A202 & A200;
  assign \new_[4284]_  = A199 & \new_[4283]_ ;
  assign \new_[4285]_  = \new_[4284]_  & \new_[4279]_ ;
  assign \new_[4288]_  = A298 & ~A203;
  assign \new_[4292]_  = A302 & ~A301;
  assign \new_[4293]_  = ~A299 & \new_[4292]_ ;
  assign \new_[4294]_  = \new_[4293]_  & \new_[4288]_ ;
  assign \new_[4297]_  = ~A167 & ~A168;
  assign \new_[4301]_  = A202 & A200;
  assign \new_[4302]_  = A199 & \new_[4301]_ ;
  assign \new_[4303]_  = \new_[4302]_  & \new_[4297]_ ;
  assign \new_[4306]_  = ~A298 & ~A203;
  assign \new_[4310]_  = A302 & ~A301;
  assign \new_[4311]_  = A299 & \new_[4310]_ ;
  assign \new_[4312]_  = \new_[4311]_  & \new_[4306]_ ;
  assign \new_[4315]_  = ~A167 & ~A168;
  assign \new_[4319]_  = A202 & A200;
  assign \new_[4320]_  = A199 & \new_[4319]_ ;
  assign \new_[4321]_  = \new_[4320]_  & \new_[4315]_ ;
  assign \new_[4324]_  = ~A298 & ~A203;
  assign \new_[4328]_  = ~A302 & A301;
  assign \new_[4329]_  = ~A299 & \new_[4328]_ ;
  assign \new_[4330]_  = \new_[4329]_  & \new_[4324]_ ;
  assign \new_[4333]_  = ~A167 & ~A168;
  assign \new_[4337]_  = ~A202 & A200;
  assign \new_[4338]_  = ~A199 & \new_[4337]_ ;
  assign \new_[4339]_  = \new_[4338]_  & \new_[4333]_ ;
  assign \new_[4342]_  = A298 & A203;
  assign \new_[4346]_  = ~A302 & A301;
  assign \new_[4347]_  = A299 & \new_[4346]_ ;
  assign \new_[4348]_  = \new_[4347]_  & \new_[4342]_ ;
  assign \new_[4351]_  = ~A167 & ~A168;
  assign \new_[4355]_  = ~A202 & A200;
  assign \new_[4356]_  = ~A199 & \new_[4355]_ ;
  assign \new_[4357]_  = \new_[4356]_  & \new_[4351]_ ;
  assign \new_[4360]_  = A298 & A203;
  assign \new_[4364]_  = A302 & ~A301;
  assign \new_[4365]_  = ~A299 & \new_[4364]_ ;
  assign \new_[4366]_  = \new_[4365]_  & \new_[4360]_ ;
  assign \new_[4369]_  = ~A167 & ~A168;
  assign \new_[4373]_  = ~A202 & A200;
  assign \new_[4374]_  = ~A199 & \new_[4373]_ ;
  assign \new_[4375]_  = \new_[4374]_  & \new_[4369]_ ;
  assign \new_[4378]_  = ~A298 & A203;
  assign \new_[4382]_  = A302 & ~A301;
  assign \new_[4383]_  = A299 & \new_[4382]_ ;
  assign \new_[4384]_  = \new_[4383]_  & \new_[4378]_ ;
  assign \new_[4387]_  = ~A167 & ~A168;
  assign \new_[4391]_  = ~A202 & A200;
  assign \new_[4392]_  = ~A199 & \new_[4391]_ ;
  assign \new_[4393]_  = \new_[4392]_  & \new_[4387]_ ;
  assign \new_[4396]_  = ~A298 & A203;
  assign \new_[4400]_  = ~A302 & A301;
  assign \new_[4401]_  = ~A299 & \new_[4400]_ ;
  assign \new_[4402]_  = \new_[4401]_  & \new_[4396]_ ;
  assign \new_[4405]_  = ~A167 & ~A168;
  assign \new_[4409]_  = ~A202 & ~A200;
  assign \new_[4410]_  = A199 & \new_[4409]_ ;
  assign \new_[4411]_  = \new_[4410]_  & \new_[4405]_ ;
  assign \new_[4414]_  = A298 & A203;
  assign \new_[4418]_  = ~A302 & A301;
  assign \new_[4419]_  = A299 & \new_[4418]_ ;
  assign \new_[4420]_  = \new_[4419]_  & \new_[4414]_ ;
  assign \new_[4423]_  = ~A167 & ~A168;
  assign \new_[4427]_  = ~A202 & ~A200;
  assign \new_[4428]_  = A199 & \new_[4427]_ ;
  assign \new_[4429]_  = \new_[4428]_  & \new_[4423]_ ;
  assign \new_[4432]_  = A298 & A203;
  assign \new_[4436]_  = A302 & ~A301;
  assign \new_[4437]_  = ~A299 & \new_[4436]_ ;
  assign \new_[4438]_  = \new_[4437]_  & \new_[4432]_ ;
  assign \new_[4441]_  = ~A167 & ~A168;
  assign \new_[4445]_  = ~A202 & ~A200;
  assign \new_[4446]_  = A199 & \new_[4445]_ ;
  assign \new_[4447]_  = \new_[4446]_  & \new_[4441]_ ;
  assign \new_[4450]_  = ~A298 & A203;
  assign \new_[4454]_  = A302 & ~A301;
  assign \new_[4455]_  = A299 & \new_[4454]_ ;
  assign \new_[4456]_  = \new_[4455]_  & \new_[4450]_ ;
  assign \new_[4459]_  = ~A167 & ~A168;
  assign \new_[4463]_  = ~A202 & ~A200;
  assign \new_[4464]_  = A199 & \new_[4463]_ ;
  assign \new_[4465]_  = \new_[4464]_  & \new_[4459]_ ;
  assign \new_[4468]_  = ~A298 & A203;
  assign \new_[4472]_  = ~A302 & A301;
  assign \new_[4473]_  = ~A299 & \new_[4472]_ ;
  assign \new_[4474]_  = \new_[4473]_  & \new_[4468]_ ;
  assign \new_[4477]_  = ~A167 & ~A168;
  assign \new_[4481]_  = A202 & ~A200;
  assign \new_[4482]_  = ~A199 & \new_[4481]_ ;
  assign \new_[4483]_  = \new_[4482]_  & \new_[4477]_ ;
  assign \new_[4486]_  = A298 & ~A203;
  assign \new_[4490]_  = ~A302 & A301;
  assign \new_[4491]_  = A299 & \new_[4490]_ ;
  assign \new_[4492]_  = \new_[4491]_  & \new_[4486]_ ;
  assign \new_[4495]_  = ~A167 & ~A168;
  assign \new_[4499]_  = A202 & ~A200;
  assign \new_[4500]_  = ~A199 & \new_[4499]_ ;
  assign \new_[4501]_  = \new_[4500]_  & \new_[4495]_ ;
  assign \new_[4504]_  = A298 & ~A203;
  assign \new_[4508]_  = A302 & ~A301;
  assign \new_[4509]_  = ~A299 & \new_[4508]_ ;
  assign \new_[4510]_  = \new_[4509]_  & \new_[4504]_ ;
  assign \new_[4513]_  = ~A167 & ~A168;
  assign \new_[4517]_  = A202 & ~A200;
  assign \new_[4518]_  = ~A199 & \new_[4517]_ ;
  assign \new_[4519]_  = \new_[4518]_  & \new_[4513]_ ;
  assign \new_[4522]_  = ~A298 & ~A203;
  assign \new_[4526]_  = A302 & ~A301;
  assign \new_[4527]_  = A299 & \new_[4526]_ ;
  assign \new_[4528]_  = \new_[4527]_  & \new_[4522]_ ;
  assign \new_[4531]_  = ~A167 & ~A168;
  assign \new_[4535]_  = A202 & ~A200;
  assign \new_[4536]_  = ~A199 & \new_[4535]_ ;
  assign \new_[4537]_  = \new_[4536]_  & \new_[4531]_ ;
  assign \new_[4540]_  = ~A298 & ~A203;
  assign \new_[4544]_  = ~A302 & A301;
  assign \new_[4545]_  = ~A299 & \new_[4544]_ ;
  assign \new_[4546]_  = \new_[4545]_  & \new_[4540]_ ;
  assign \new_[4549]_  = A168 & A170;
  assign \new_[4553]_  = A199 & A166;
  assign \new_[4554]_  = ~A167 & \new_[4553]_ ;
  assign \new_[4555]_  = \new_[4554]_  & \new_[4549]_ ;
  assign \new_[4558]_  = ~A201 & A200;
  assign \new_[4562]_  = A300 & A299;
  assign \new_[4563]_  = ~A202 & \new_[4562]_ ;
  assign \new_[4564]_  = \new_[4563]_  & \new_[4558]_ ;
  assign \new_[4567]_  = A168 & A170;
  assign \new_[4571]_  = A199 & A166;
  assign \new_[4572]_  = ~A167 & \new_[4571]_ ;
  assign \new_[4573]_  = \new_[4572]_  & \new_[4567]_ ;
  assign \new_[4576]_  = ~A201 & A200;
  assign \new_[4580]_  = A300 & A298;
  assign \new_[4581]_  = ~A202 & \new_[4580]_ ;
  assign \new_[4582]_  = \new_[4581]_  & \new_[4576]_ ;
  assign \new_[4585]_  = A168 & A170;
  assign \new_[4589]_  = A199 & A166;
  assign \new_[4590]_  = ~A167 & \new_[4589]_ ;
  assign \new_[4591]_  = \new_[4590]_  & \new_[4585]_ ;
  assign \new_[4594]_  = ~A201 & A200;
  assign \new_[4598]_  = A300 & A299;
  assign \new_[4599]_  = A203 & \new_[4598]_ ;
  assign \new_[4600]_  = \new_[4599]_  & \new_[4594]_ ;
  assign \new_[4603]_  = A168 & A170;
  assign \new_[4607]_  = A199 & A166;
  assign \new_[4608]_  = ~A167 & \new_[4607]_ ;
  assign \new_[4609]_  = \new_[4608]_  & \new_[4603]_ ;
  assign \new_[4612]_  = ~A201 & A200;
  assign \new_[4616]_  = A300 & A298;
  assign \new_[4617]_  = A203 & \new_[4616]_ ;
  assign \new_[4618]_  = \new_[4617]_  & \new_[4612]_ ;
  assign \new_[4621]_  = A168 & A170;
  assign \new_[4625]_  = ~A199 & A166;
  assign \new_[4626]_  = ~A167 & \new_[4625]_ ;
  assign \new_[4627]_  = \new_[4626]_  & \new_[4621]_ ;
  assign \new_[4630]_  = ~A201 & A200;
  assign \new_[4634]_  = A300 & A299;
  assign \new_[4635]_  = A202 & \new_[4634]_ ;
  assign \new_[4636]_  = \new_[4635]_  & \new_[4630]_ ;
  assign \new_[4639]_  = A168 & A170;
  assign \new_[4643]_  = ~A199 & A166;
  assign \new_[4644]_  = ~A167 & \new_[4643]_ ;
  assign \new_[4645]_  = \new_[4644]_  & \new_[4639]_ ;
  assign \new_[4648]_  = ~A201 & A200;
  assign \new_[4652]_  = A300 & A298;
  assign \new_[4653]_  = A202 & \new_[4652]_ ;
  assign \new_[4654]_  = \new_[4653]_  & \new_[4648]_ ;
  assign \new_[4657]_  = A168 & A170;
  assign \new_[4661]_  = ~A199 & A166;
  assign \new_[4662]_  = ~A167 & \new_[4661]_ ;
  assign \new_[4663]_  = \new_[4662]_  & \new_[4657]_ ;
  assign \new_[4666]_  = ~A201 & A200;
  assign \new_[4670]_  = A300 & A299;
  assign \new_[4671]_  = ~A203 & \new_[4670]_ ;
  assign \new_[4672]_  = \new_[4671]_  & \new_[4666]_ ;
  assign \new_[4675]_  = A168 & A170;
  assign \new_[4679]_  = ~A199 & A166;
  assign \new_[4680]_  = ~A167 & \new_[4679]_ ;
  assign \new_[4681]_  = \new_[4680]_  & \new_[4675]_ ;
  assign \new_[4684]_  = ~A201 & A200;
  assign \new_[4688]_  = A300 & A298;
  assign \new_[4689]_  = ~A203 & \new_[4688]_ ;
  assign \new_[4690]_  = \new_[4689]_  & \new_[4684]_ ;
  assign \new_[4693]_  = A168 & A170;
  assign \new_[4697]_  = A199 & A166;
  assign \new_[4698]_  = ~A167 & \new_[4697]_ ;
  assign \new_[4699]_  = \new_[4698]_  & \new_[4693]_ ;
  assign \new_[4702]_  = ~A201 & ~A200;
  assign \new_[4706]_  = A300 & A299;
  assign \new_[4707]_  = A202 & \new_[4706]_ ;
  assign \new_[4708]_  = \new_[4707]_  & \new_[4702]_ ;
  assign \new_[4711]_  = A168 & A170;
  assign \new_[4715]_  = A199 & A166;
  assign \new_[4716]_  = ~A167 & \new_[4715]_ ;
  assign \new_[4717]_  = \new_[4716]_  & \new_[4711]_ ;
  assign \new_[4720]_  = ~A201 & ~A200;
  assign \new_[4724]_  = A300 & A298;
  assign \new_[4725]_  = A202 & \new_[4724]_ ;
  assign \new_[4726]_  = \new_[4725]_  & \new_[4720]_ ;
  assign \new_[4729]_  = A168 & A170;
  assign \new_[4733]_  = A199 & A166;
  assign \new_[4734]_  = ~A167 & \new_[4733]_ ;
  assign \new_[4735]_  = \new_[4734]_  & \new_[4729]_ ;
  assign \new_[4738]_  = ~A201 & ~A200;
  assign \new_[4742]_  = A300 & A299;
  assign \new_[4743]_  = ~A203 & \new_[4742]_ ;
  assign \new_[4744]_  = \new_[4743]_  & \new_[4738]_ ;
  assign \new_[4747]_  = A168 & A170;
  assign \new_[4751]_  = A199 & A166;
  assign \new_[4752]_  = ~A167 & \new_[4751]_ ;
  assign \new_[4753]_  = \new_[4752]_  & \new_[4747]_ ;
  assign \new_[4756]_  = ~A201 & ~A200;
  assign \new_[4760]_  = A300 & A298;
  assign \new_[4761]_  = ~A203 & \new_[4760]_ ;
  assign \new_[4762]_  = \new_[4761]_  & \new_[4756]_ ;
  assign \new_[4765]_  = A168 & A169;
  assign \new_[4769]_  = A199 & A166;
  assign \new_[4770]_  = ~A167 & \new_[4769]_ ;
  assign \new_[4771]_  = \new_[4770]_  & \new_[4765]_ ;
  assign \new_[4774]_  = ~A201 & A200;
  assign \new_[4778]_  = A300 & A299;
  assign \new_[4779]_  = ~A202 & \new_[4778]_ ;
  assign \new_[4780]_  = \new_[4779]_  & \new_[4774]_ ;
  assign \new_[4783]_  = A168 & A169;
  assign \new_[4787]_  = A199 & A166;
  assign \new_[4788]_  = ~A167 & \new_[4787]_ ;
  assign \new_[4789]_  = \new_[4788]_  & \new_[4783]_ ;
  assign \new_[4792]_  = ~A201 & A200;
  assign \new_[4796]_  = A300 & A298;
  assign \new_[4797]_  = ~A202 & \new_[4796]_ ;
  assign \new_[4798]_  = \new_[4797]_  & \new_[4792]_ ;
  assign \new_[4801]_  = A168 & A169;
  assign \new_[4805]_  = A199 & A166;
  assign \new_[4806]_  = ~A167 & \new_[4805]_ ;
  assign \new_[4807]_  = \new_[4806]_  & \new_[4801]_ ;
  assign \new_[4810]_  = ~A201 & A200;
  assign \new_[4814]_  = A300 & A299;
  assign \new_[4815]_  = A203 & \new_[4814]_ ;
  assign \new_[4816]_  = \new_[4815]_  & \new_[4810]_ ;
  assign \new_[4819]_  = A168 & A169;
  assign \new_[4823]_  = A199 & A166;
  assign \new_[4824]_  = ~A167 & \new_[4823]_ ;
  assign \new_[4825]_  = \new_[4824]_  & \new_[4819]_ ;
  assign \new_[4828]_  = ~A201 & A200;
  assign \new_[4832]_  = A300 & A298;
  assign \new_[4833]_  = A203 & \new_[4832]_ ;
  assign \new_[4834]_  = \new_[4833]_  & \new_[4828]_ ;
  assign \new_[4837]_  = A168 & A169;
  assign \new_[4841]_  = ~A199 & A166;
  assign \new_[4842]_  = ~A167 & \new_[4841]_ ;
  assign \new_[4843]_  = \new_[4842]_  & \new_[4837]_ ;
  assign \new_[4846]_  = ~A201 & A200;
  assign \new_[4850]_  = A300 & A299;
  assign \new_[4851]_  = A202 & \new_[4850]_ ;
  assign \new_[4852]_  = \new_[4851]_  & \new_[4846]_ ;
  assign \new_[4855]_  = A168 & A169;
  assign \new_[4859]_  = ~A199 & A166;
  assign \new_[4860]_  = ~A167 & \new_[4859]_ ;
  assign \new_[4861]_  = \new_[4860]_  & \new_[4855]_ ;
  assign \new_[4864]_  = ~A201 & A200;
  assign \new_[4868]_  = A300 & A298;
  assign \new_[4869]_  = A202 & \new_[4868]_ ;
  assign \new_[4870]_  = \new_[4869]_  & \new_[4864]_ ;
  assign \new_[4873]_  = A168 & A169;
  assign \new_[4877]_  = ~A199 & A166;
  assign \new_[4878]_  = ~A167 & \new_[4877]_ ;
  assign \new_[4879]_  = \new_[4878]_  & \new_[4873]_ ;
  assign \new_[4882]_  = ~A201 & A200;
  assign \new_[4886]_  = A300 & A299;
  assign \new_[4887]_  = ~A203 & \new_[4886]_ ;
  assign \new_[4888]_  = \new_[4887]_  & \new_[4882]_ ;
  assign \new_[4891]_  = A168 & A169;
  assign \new_[4895]_  = ~A199 & A166;
  assign \new_[4896]_  = ~A167 & \new_[4895]_ ;
  assign \new_[4897]_  = \new_[4896]_  & \new_[4891]_ ;
  assign \new_[4900]_  = ~A201 & A200;
  assign \new_[4904]_  = A300 & A298;
  assign \new_[4905]_  = ~A203 & \new_[4904]_ ;
  assign \new_[4906]_  = \new_[4905]_  & \new_[4900]_ ;
  assign \new_[4909]_  = A168 & A169;
  assign \new_[4913]_  = A199 & A166;
  assign \new_[4914]_  = ~A167 & \new_[4913]_ ;
  assign \new_[4915]_  = \new_[4914]_  & \new_[4909]_ ;
  assign \new_[4918]_  = ~A201 & ~A200;
  assign \new_[4922]_  = A300 & A299;
  assign \new_[4923]_  = A202 & \new_[4922]_ ;
  assign \new_[4924]_  = \new_[4923]_  & \new_[4918]_ ;
  assign \new_[4927]_  = A168 & A169;
  assign \new_[4931]_  = A199 & A166;
  assign \new_[4932]_  = ~A167 & \new_[4931]_ ;
  assign \new_[4933]_  = \new_[4932]_  & \new_[4927]_ ;
  assign \new_[4936]_  = ~A201 & ~A200;
  assign \new_[4940]_  = A300 & A298;
  assign \new_[4941]_  = A202 & \new_[4940]_ ;
  assign \new_[4942]_  = \new_[4941]_  & \new_[4936]_ ;
  assign \new_[4945]_  = A168 & A169;
  assign \new_[4949]_  = A199 & A166;
  assign \new_[4950]_  = ~A167 & \new_[4949]_ ;
  assign \new_[4951]_  = \new_[4950]_  & \new_[4945]_ ;
  assign \new_[4954]_  = ~A201 & ~A200;
  assign \new_[4958]_  = A300 & A299;
  assign \new_[4959]_  = ~A203 & \new_[4958]_ ;
  assign \new_[4960]_  = \new_[4959]_  & \new_[4954]_ ;
  assign \new_[4963]_  = A168 & A169;
  assign \new_[4967]_  = A199 & A166;
  assign \new_[4968]_  = ~A167 & \new_[4967]_ ;
  assign \new_[4969]_  = \new_[4968]_  & \new_[4963]_ ;
  assign \new_[4972]_  = ~A201 & ~A200;
  assign \new_[4976]_  = A300 & A298;
  assign \new_[4977]_  = ~A203 & \new_[4976]_ ;
  assign \new_[4978]_  = \new_[4977]_  & \new_[4972]_ ;
  assign \new_[4981]_  = A168 & A170;
  assign \new_[4985]_  = ~A199 & A166;
  assign \new_[4986]_  = ~A167 & \new_[4985]_ ;
  assign \new_[4987]_  = \new_[4986]_  & \new_[4981]_ ;
  assign \new_[4991]_  = A298 & ~A202;
  assign \new_[4992]_  = ~A200 & \new_[4991]_ ;
  assign \new_[4996]_  = ~A302 & A301;
  assign \new_[4997]_  = A299 & \new_[4996]_ ;
  assign \new_[4998]_  = \new_[4997]_  & \new_[4992]_ ;
  assign \new_[5001]_  = A168 & A170;
  assign \new_[5005]_  = ~A199 & A166;
  assign \new_[5006]_  = ~A167 & \new_[5005]_ ;
  assign \new_[5007]_  = \new_[5006]_  & \new_[5001]_ ;
  assign \new_[5011]_  = A298 & ~A202;
  assign \new_[5012]_  = ~A200 & \new_[5011]_ ;
  assign \new_[5016]_  = A302 & ~A301;
  assign \new_[5017]_  = ~A299 & \new_[5016]_ ;
  assign \new_[5018]_  = \new_[5017]_  & \new_[5012]_ ;
  assign \new_[5021]_  = A168 & A170;
  assign \new_[5025]_  = ~A199 & A166;
  assign \new_[5026]_  = ~A167 & \new_[5025]_ ;
  assign \new_[5027]_  = \new_[5026]_  & \new_[5021]_ ;
  assign \new_[5031]_  = ~A298 & ~A202;
  assign \new_[5032]_  = ~A200 & \new_[5031]_ ;
  assign \new_[5036]_  = A302 & ~A301;
  assign \new_[5037]_  = A299 & \new_[5036]_ ;
  assign \new_[5038]_  = \new_[5037]_  & \new_[5032]_ ;
  assign \new_[5041]_  = A168 & A170;
  assign \new_[5045]_  = ~A199 & A166;
  assign \new_[5046]_  = ~A167 & \new_[5045]_ ;
  assign \new_[5047]_  = \new_[5046]_  & \new_[5041]_ ;
  assign \new_[5051]_  = ~A298 & ~A202;
  assign \new_[5052]_  = ~A200 & \new_[5051]_ ;
  assign \new_[5056]_  = ~A302 & A301;
  assign \new_[5057]_  = ~A299 & \new_[5056]_ ;
  assign \new_[5058]_  = \new_[5057]_  & \new_[5052]_ ;
  assign \new_[5061]_  = A168 & A170;
  assign \new_[5065]_  = ~A199 & A166;
  assign \new_[5066]_  = ~A167 & \new_[5065]_ ;
  assign \new_[5067]_  = \new_[5066]_  & \new_[5061]_ ;
  assign \new_[5071]_  = A298 & A203;
  assign \new_[5072]_  = ~A200 & \new_[5071]_ ;
  assign \new_[5076]_  = ~A302 & A301;
  assign \new_[5077]_  = A299 & \new_[5076]_ ;
  assign \new_[5078]_  = \new_[5077]_  & \new_[5072]_ ;
  assign \new_[5081]_  = A168 & A170;
  assign \new_[5085]_  = ~A199 & A166;
  assign \new_[5086]_  = ~A167 & \new_[5085]_ ;
  assign \new_[5087]_  = \new_[5086]_  & \new_[5081]_ ;
  assign \new_[5091]_  = A298 & A203;
  assign \new_[5092]_  = ~A200 & \new_[5091]_ ;
  assign \new_[5096]_  = A302 & ~A301;
  assign \new_[5097]_  = ~A299 & \new_[5096]_ ;
  assign \new_[5098]_  = \new_[5097]_  & \new_[5092]_ ;
  assign \new_[5101]_  = A168 & A170;
  assign \new_[5105]_  = ~A199 & A166;
  assign \new_[5106]_  = ~A167 & \new_[5105]_ ;
  assign \new_[5107]_  = \new_[5106]_  & \new_[5101]_ ;
  assign \new_[5111]_  = ~A298 & A203;
  assign \new_[5112]_  = ~A200 & \new_[5111]_ ;
  assign \new_[5116]_  = A302 & ~A301;
  assign \new_[5117]_  = A299 & \new_[5116]_ ;
  assign \new_[5118]_  = \new_[5117]_  & \new_[5112]_ ;
  assign \new_[5121]_  = A168 & A170;
  assign \new_[5125]_  = ~A199 & A166;
  assign \new_[5126]_  = ~A167 & \new_[5125]_ ;
  assign \new_[5127]_  = \new_[5126]_  & \new_[5121]_ ;
  assign \new_[5131]_  = ~A298 & A203;
  assign \new_[5132]_  = ~A200 & \new_[5131]_ ;
  assign \new_[5136]_  = ~A302 & A301;
  assign \new_[5137]_  = ~A299 & \new_[5136]_ ;
  assign \new_[5138]_  = \new_[5137]_  & \new_[5132]_ ;
  assign \new_[5141]_  = A168 & A169;
  assign \new_[5145]_  = ~A199 & A166;
  assign \new_[5146]_  = ~A167 & \new_[5145]_ ;
  assign \new_[5147]_  = \new_[5146]_  & \new_[5141]_ ;
  assign \new_[5151]_  = A298 & ~A202;
  assign \new_[5152]_  = ~A200 & \new_[5151]_ ;
  assign \new_[5156]_  = ~A302 & A301;
  assign \new_[5157]_  = A299 & \new_[5156]_ ;
  assign \new_[5158]_  = \new_[5157]_  & \new_[5152]_ ;
  assign \new_[5161]_  = A168 & A169;
  assign \new_[5165]_  = ~A199 & A166;
  assign \new_[5166]_  = ~A167 & \new_[5165]_ ;
  assign \new_[5167]_  = \new_[5166]_  & \new_[5161]_ ;
  assign \new_[5171]_  = A298 & ~A202;
  assign \new_[5172]_  = ~A200 & \new_[5171]_ ;
  assign \new_[5176]_  = A302 & ~A301;
  assign \new_[5177]_  = ~A299 & \new_[5176]_ ;
  assign \new_[5178]_  = \new_[5177]_  & \new_[5172]_ ;
  assign \new_[5181]_  = A168 & A169;
  assign \new_[5185]_  = ~A199 & A166;
  assign \new_[5186]_  = ~A167 & \new_[5185]_ ;
  assign \new_[5187]_  = \new_[5186]_  & \new_[5181]_ ;
  assign \new_[5191]_  = ~A298 & ~A202;
  assign \new_[5192]_  = ~A200 & \new_[5191]_ ;
  assign \new_[5196]_  = A302 & ~A301;
  assign \new_[5197]_  = A299 & \new_[5196]_ ;
  assign \new_[5198]_  = \new_[5197]_  & \new_[5192]_ ;
  assign \new_[5201]_  = A168 & A169;
  assign \new_[5205]_  = ~A199 & A166;
  assign \new_[5206]_  = ~A167 & \new_[5205]_ ;
  assign \new_[5207]_  = \new_[5206]_  & \new_[5201]_ ;
  assign \new_[5211]_  = ~A298 & ~A202;
  assign \new_[5212]_  = ~A200 & \new_[5211]_ ;
  assign \new_[5216]_  = ~A302 & A301;
  assign \new_[5217]_  = ~A299 & \new_[5216]_ ;
  assign \new_[5218]_  = \new_[5217]_  & \new_[5212]_ ;
  assign \new_[5221]_  = A168 & A169;
  assign \new_[5225]_  = ~A199 & A166;
  assign \new_[5226]_  = ~A167 & \new_[5225]_ ;
  assign \new_[5227]_  = \new_[5226]_  & \new_[5221]_ ;
  assign \new_[5231]_  = A298 & A203;
  assign \new_[5232]_  = ~A200 & \new_[5231]_ ;
  assign \new_[5236]_  = ~A302 & A301;
  assign \new_[5237]_  = A299 & \new_[5236]_ ;
  assign \new_[5238]_  = \new_[5237]_  & \new_[5232]_ ;
  assign \new_[5241]_  = A168 & A169;
  assign \new_[5245]_  = ~A199 & A166;
  assign \new_[5246]_  = ~A167 & \new_[5245]_ ;
  assign \new_[5247]_  = \new_[5246]_  & \new_[5241]_ ;
  assign \new_[5251]_  = A298 & A203;
  assign \new_[5252]_  = ~A200 & \new_[5251]_ ;
  assign \new_[5256]_  = A302 & ~A301;
  assign \new_[5257]_  = ~A299 & \new_[5256]_ ;
  assign \new_[5258]_  = \new_[5257]_  & \new_[5252]_ ;
  assign \new_[5261]_  = A168 & A169;
  assign \new_[5265]_  = ~A199 & A166;
  assign \new_[5266]_  = ~A167 & \new_[5265]_ ;
  assign \new_[5267]_  = \new_[5266]_  & \new_[5261]_ ;
  assign \new_[5271]_  = ~A298 & A203;
  assign \new_[5272]_  = ~A200 & \new_[5271]_ ;
  assign \new_[5276]_  = A302 & ~A301;
  assign \new_[5277]_  = A299 & \new_[5276]_ ;
  assign \new_[5278]_  = \new_[5277]_  & \new_[5272]_ ;
  assign \new_[5281]_  = A168 & A169;
  assign \new_[5285]_  = ~A199 & A166;
  assign \new_[5286]_  = ~A167 & \new_[5285]_ ;
  assign \new_[5287]_  = \new_[5286]_  & \new_[5281]_ ;
  assign \new_[5291]_  = ~A298 & A203;
  assign \new_[5292]_  = ~A200 & \new_[5291]_ ;
  assign \new_[5296]_  = ~A302 & A301;
  assign \new_[5297]_  = ~A299 & \new_[5296]_ ;
  assign \new_[5298]_  = \new_[5297]_  & \new_[5292]_ ;
  assign \new_[5301]_  = ~A169 & ~A170;
  assign \new_[5305]_  = A200 & A199;
  assign \new_[5306]_  = ~A167 & \new_[5305]_ ;
  assign \new_[5307]_  = \new_[5306]_  & \new_[5301]_ ;
  assign \new_[5311]_  = A298 & ~A203;
  assign \new_[5312]_  = A202 & \new_[5311]_ ;
  assign \new_[5316]_  = ~A302 & A301;
  assign \new_[5317]_  = A299 & \new_[5316]_ ;
  assign \new_[5318]_  = \new_[5317]_  & \new_[5312]_ ;
  assign \new_[5321]_  = ~A169 & ~A170;
  assign \new_[5325]_  = A200 & A199;
  assign \new_[5326]_  = ~A167 & \new_[5325]_ ;
  assign \new_[5327]_  = \new_[5326]_  & \new_[5321]_ ;
  assign \new_[5331]_  = A298 & ~A203;
  assign \new_[5332]_  = A202 & \new_[5331]_ ;
  assign \new_[5336]_  = A302 & ~A301;
  assign \new_[5337]_  = ~A299 & \new_[5336]_ ;
  assign \new_[5338]_  = \new_[5337]_  & \new_[5332]_ ;
  assign \new_[5341]_  = ~A169 & ~A170;
  assign \new_[5345]_  = A200 & A199;
  assign \new_[5346]_  = ~A167 & \new_[5345]_ ;
  assign \new_[5347]_  = \new_[5346]_  & \new_[5341]_ ;
  assign \new_[5351]_  = ~A298 & ~A203;
  assign \new_[5352]_  = A202 & \new_[5351]_ ;
  assign \new_[5356]_  = A302 & ~A301;
  assign \new_[5357]_  = A299 & \new_[5356]_ ;
  assign \new_[5358]_  = \new_[5357]_  & \new_[5352]_ ;
  assign \new_[5361]_  = ~A169 & ~A170;
  assign \new_[5365]_  = A200 & A199;
  assign \new_[5366]_  = ~A167 & \new_[5365]_ ;
  assign \new_[5367]_  = \new_[5366]_  & \new_[5361]_ ;
  assign \new_[5371]_  = ~A298 & ~A203;
  assign \new_[5372]_  = A202 & \new_[5371]_ ;
  assign \new_[5376]_  = ~A302 & A301;
  assign \new_[5377]_  = ~A299 & \new_[5376]_ ;
  assign \new_[5378]_  = \new_[5377]_  & \new_[5372]_ ;
  assign \new_[5381]_  = ~A169 & ~A170;
  assign \new_[5385]_  = A200 & ~A199;
  assign \new_[5386]_  = ~A167 & \new_[5385]_ ;
  assign \new_[5387]_  = \new_[5386]_  & \new_[5381]_ ;
  assign \new_[5391]_  = A298 & A203;
  assign \new_[5392]_  = ~A202 & \new_[5391]_ ;
  assign \new_[5396]_  = ~A302 & A301;
  assign \new_[5397]_  = A299 & \new_[5396]_ ;
  assign \new_[5398]_  = \new_[5397]_  & \new_[5392]_ ;
  assign \new_[5401]_  = ~A169 & ~A170;
  assign \new_[5405]_  = A200 & ~A199;
  assign \new_[5406]_  = ~A167 & \new_[5405]_ ;
  assign \new_[5407]_  = \new_[5406]_  & \new_[5401]_ ;
  assign \new_[5411]_  = A298 & A203;
  assign \new_[5412]_  = ~A202 & \new_[5411]_ ;
  assign \new_[5416]_  = A302 & ~A301;
  assign \new_[5417]_  = ~A299 & \new_[5416]_ ;
  assign \new_[5418]_  = \new_[5417]_  & \new_[5412]_ ;
  assign \new_[5421]_  = ~A169 & ~A170;
  assign \new_[5425]_  = A200 & ~A199;
  assign \new_[5426]_  = ~A167 & \new_[5425]_ ;
  assign \new_[5427]_  = \new_[5426]_  & \new_[5421]_ ;
  assign \new_[5431]_  = ~A298 & A203;
  assign \new_[5432]_  = ~A202 & \new_[5431]_ ;
  assign \new_[5436]_  = A302 & ~A301;
  assign \new_[5437]_  = A299 & \new_[5436]_ ;
  assign \new_[5438]_  = \new_[5437]_  & \new_[5432]_ ;
  assign \new_[5441]_  = ~A169 & ~A170;
  assign \new_[5445]_  = A200 & ~A199;
  assign \new_[5446]_  = ~A167 & \new_[5445]_ ;
  assign \new_[5447]_  = \new_[5446]_  & \new_[5441]_ ;
  assign \new_[5451]_  = ~A298 & A203;
  assign \new_[5452]_  = ~A202 & \new_[5451]_ ;
  assign \new_[5456]_  = ~A302 & A301;
  assign \new_[5457]_  = ~A299 & \new_[5456]_ ;
  assign \new_[5458]_  = \new_[5457]_  & \new_[5452]_ ;
  assign \new_[5461]_  = ~A169 & ~A170;
  assign \new_[5465]_  = ~A200 & A199;
  assign \new_[5466]_  = ~A167 & \new_[5465]_ ;
  assign \new_[5467]_  = \new_[5466]_  & \new_[5461]_ ;
  assign \new_[5471]_  = A298 & A203;
  assign \new_[5472]_  = ~A202 & \new_[5471]_ ;
  assign \new_[5476]_  = ~A302 & A301;
  assign \new_[5477]_  = A299 & \new_[5476]_ ;
  assign \new_[5478]_  = \new_[5477]_  & \new_[5472]_ ;
  assign \new_[5481]_  = ~A169 & ~A170;
  assign \new_[5485]_  = ~A200 & A199;
  assign \new_[5486]_  = ~A167 & \new_[5485]_ ;
  assign \new_[5487]_  = \new_[5486]_  & \new_[5481]_ ;
  assign \new_[5491]_  = A298 & A203;
  assign \new_[5492]_  = ~A202 & \new_[5491]_ ;
  assign \new_[5496]_  = A302 & ~A301;
  assign \new_[5497]_  = ~A299 & \new_[5496]_ ;
  assign \new_[5498]_  = \new_[5497]_  & \new_[5492]_ ;
  assign \new_[5501]_  = ~A169 & ~A170;
  assign \new_[5505]_  = ~A200 & A199;
  assign \new_[5506]_  = ~A167 & \new_[5505]_ ;
  assign \new_[5507]_  = \new_[5506]_  & \new_[5501]_ ;
  assign \new_[5511]_  = ~A298 & A203;
  assign \new_[5512]_  = ~A202 & \new_[5511]_ ;
  assign \new_[5516]_  = A302 & ~A301;
  assign \new_[5517]_  = A299 & \new_[5516]_ ;
  assign \new_[5518]_  = \new_[5517]_  & \new_[5512]_ ;
  assign \new_[5521]_  = ~A169 & ~A170;
  assign \new_[5525]_  = ~A200 & A199;
  assign \new_[5526]_  = ~A167 & \new_[5525]_ ;
  assign \new_[5527]_  = \new_[5526]_  & \new_[5521]_ ;
  assign \new_[5531]_  = ~A298 & A203;
  assign \new_[5532]_  = ~A202 & \new_[5531]_ ;
  assign \new_[5536]_  = ~A302 & A301;
  assign \new_[5537]_  = ~A299 & \new_[5536]_ ;
  assign \new_[5538]_  = \new_[5537]_  & \new_[5532]_ ;
  assign \new_[5541]_  = ~A169 & ~A170;
  assign \new_[5545]_  = ~A200 & ~A199;
  assign \new_[5546]_  = ~A167 & \new_[5545]_ ;
  assign \new_[5547]_  = \new_[5546]_  & \new_[5541]_ ;
  assign \new_[5551]_  = A298 & ~A203;
  assign \new_[5552]_  = A202 & \new_[5551]_ ;
  assign \new_[5556]_  = ~A302 & A301;
  assign \new_[5557]_  = A299 & \new_[5556]_ ;
  assign \new_[5558]_  = \new_[5557]_  & \new_[5552]_ ;
  assign \new_[5561]_  = ~A169 & ~A170;
  assign \new_[5565]_  = ~A200 & ~A199;
  assign \new_[5566]_  = ~A167 & \new_[5565]_ ;
  assign \new_[5567]_  = \new_[5566]_  & \new_[5561]_ ;
  assign \new_[5571]_  = A298 & ~A203;
  assign \new_[5572]_  = A202 & \new_[5571]_ ;
  assign \new_[5576]_  = A302 & ~A301;
  assign \new_[5577]_  = ~A299 & \new_[5576]_ ;
  assign \new_[5578]_  = \new_[5577]_  & \new_[5572]_ ;
  assign \new_[5581]_  = ~A169 & ~A170;
  assign \new_[5585]_  = ~A200 & ~A199;
  assign \new_[5586]_  = ~A167 & \new_[5585]_ ;
  assign \new_[5587]_  = \new_[5586]_  & \new_[5581]_ ;
  assign \new_[5591]_  = ~A298 & ~A203;
  assign \new_[5592]_  = A202 & \new_[5591]_ ;
  assign \new_[5596]_  = A302 & ~A301;
  assign \new_[5597]_  = A299 & \new_[5596]_ ;
  assign \new_[5598]_  = \new_[5597]_  & \new_[5592]_ ;
  assign \new_[5601]_  = ~A169 & ~A170;
  assign \new_[5605]_  = ~A200 & ~A199;
  assign \new_[5606]_  = ~A167 & \new_[5605]_ ;
  assign \new_[5607]_  = \new_[5606]_  & \new_[5601]_ ;
  assign \new_[5611]_  = ~A298 & ~A203;
  assign \new_[5612]_  = A202 & \new_[5611]_ ;
  assign \new_[5616]_  = ~A302 & A301;
  assign \new_[5617]_  = ~A299 & \new_[5616]_ ;
  assign \new_[5618]_  = \new_[5617]_  & \new_[5612]_ ;
  assign \new_[5622]_  = ~A167 & A168;
  assign \new_[5623]_  = A170 & \new_[5622]_ ;
  assign \new_[5627]_  = A200 & A199;
  assign \new_[5628]_  = A166 & \new_[5627]_ ;
  assign \new_[5629]_  = \new_[5628]_  & \new_[5623]_ ;
  assign \new_[5633]_  = A298 & ~A202;
  assign \new_[5634]_  = ~A201 & \new_[5633]_ ;
  assign \new_[5638]_  = ~A302 & A301;
  assign \new_[5639]_  = A299 & \new_[5638]_ ;
  assign \new_[5640]_  = \new_[5639]_  & \new_[5634]_ ;
  assign \new_[5644]_  = ~A167 & A168;
  assign \new_[5645]_  = A170 & \new_[5644]_ ;
  assign \new_[5649]_  = A200 & A199;
  assign \new_[5650]_  = A166 & \new_[5649]_ ;
  assign \new_[5651]_  = \new_[5650]_  & \new_[5645]_ ;
  assign \new_[5655]_  = A298 & ~A202;
  assign \new_[5656]_  = ~A201 & \new_[5655]_ ;
  assign \new_[5660]_  = A302 & ~A301;
  assign \new_[5661]_  = ~A299 & \new_[5660]_ ;
  assign \new_[5662]_  = \new_[5661]_  & \new_[5656]_ ;
  assign \new_[5666]_  = ~A167 & A168;
  assign \new_[5667]_  = A170 & \new_[5666]_ ;
  assign \new_[5671]_  = A200 & A199;
  assign \new_[5672]_  = A166 & \new_[5671]_ ;
  assign \new_[5673]_  = \new_[5672]_  & \new_[5667]_ ;
  assign \new_[5677]_  = ~A298 & ~A202;
  assign \new_[5678]_  = ~A201 & \new_[5677]_ ;
  assign \new_[5682]_  = A302 & ~A301;
  assign \new_[5683]_  = A299 & \new_[5682]_ ;
  assign \new_[5684]_  = \new_[5683]_  & \new_[5678]_ ;
  assign \new_[5688]_  = ~A167 & A168;
  assign \new_[5689]_  = A170 & \new_[5688]_ ;
  assign \new_[5693]_  = A200 & A199;
  assign \new_[5694]_  = A166 & \new_[5693]_ ;
  assign \new_[5695]_  = \new_[5694]_  & \new_[5689]_ ;
  assign \new_[5699]_  = ~A298 & ~A202;
  assign \new_[5700]_  = ~A201 & \new_[5699]_ ;
  assign \new_[5704]_  = ~A302 & A301;
  assign \new_[5705]_  = ~A299 & \new_[5704]_ ;
  assign \new_[5706]_  = \new_[5705]_  & \new_[5700]_ ;
  assign \new_[5710]_  = ~A167 & A168;
  assign \new_[5711]_  = A170 & \new_[5710]_ ;
  assign \new_[5715]_  = A200 & A199;
  assign \new_[5716]_  = A166 & \new_[5715]_ ;
  assign \new_[5717]_  = \new_[5716]_  & \new_[5711]_ ;
  assign \new_[5721]_  = A298 & A203;
  assign \new_[5722]_  = ~A201 & \new_[5721]_ ;
  assign \new_[5726]_  = ~A302 & A301;
  assign \new_[5727]_  = A299 & \new_[5726]_ ;
  assign \new_[5728]_  = \new_[5727]_  & \new_[5722]_ ;
  assign \new_[5732]_  = ~A167 & A168;
  assign \new_[5733]_  = A170 & \new_[5732]_ ;
  assign \new_[5737]_  = A200 & A199;
  assign \new_[5738]_  = A166 & \new_[5737]_ ;
  assign \new_[5739]_  = \new_[5738]_  & \new_[5733]_ ;
  assign \new_[5743]_  = A298 & A203;
  assign \new_[5744]_  = ~A201 & \new_[5743]_ ;
  assign \new_[5748]_  = A302 & ~A301;
  assign \new_[5749]_  = ~A299 & \new_[5748]_ ;
  assign \new_[5750]_  = \new_[5749]_  & \new_[5744]_ ;
  assign \new_[5754]_  = ~A167 & A168;
  assign \new_[5755]_  = A170 & \new_[5754]_ ;
  assign \new_[5759]_  = A200 & A199;
  assign \new_[5760]_  = A166 & \new_[5759]_ ;
  assign \new_[5761]_  = \new_[5760]_  & \new_[5755]_ ;
  assign \new_[5765]_  = ~A298 & A203;
  assign \new_[5766]_  = ~A201 & \new_[5765]_ ;
  assign \new_[5770]_  = A302 & ~A301;
  assign \new_[5771]_  = A299 & \new_[5770]_ ;
  assign \new_[5772]_  = \new_[5771]_  & \new_[5766]_ ;
  assign \new_[5776]_  = ~A167 & A168;
  assign \new_[5777]_  = A170 & \new_[5776]_ ;
  assign \new_[5781]_  = A200 & A199;
  assign \new_[5782]_  = A166 & \new_[5781]_ ;
  assign \new_[5783]_  = \new_[5782]_  & \new_[5777]_ ;
  assign \new_[5787]_  = ~A298 & A203;
  assign \new_[5788]_  = ~A201 & \new_[5787]_ ;
  assign \new_[5792]_  = ~A302 & A301;
  assign \new_[5793]_  = ~A299 & \new_[5792]_ ;
  assign \new_[5794]_  = \new_[5793]_  & \new_[5788]_ ;
  assign \new_[5798]_  = ~A167 & A168;
  assign \new_[5799]_  = A170 & \new_[5798]_ ;
  assign \new_[5803]_  = A200 & ~A199;
  assign \new_[5804]_  = A166 & \new_[5803]_ ;
  assign \new_[5805]_  = \new_[5804]_  & \new_[5799]_ ;
  assign \new_[5809]_  = A298 & A202;
  assign \new_[5810]_  = ~A201 & \new_[5809]_ ;
  assign \new_[5814]_  = ~A302 & A301;
  assign \new_[5815]_  = A299 & \new_[5814]_ ;
  assign \new_[5816]_  = \new_[5815]_  & \new_[5810]_ ;
  assign \new_[5820]_  = ~A167 & A168;
  assign \new_[5821]_  = A170 & \new_[5820]_ ;
  assign \new_[5825]_  = A200 & ~A199;
  assign \new_[5826]_  = A166 & \new_[5825]_ ;
  assign \new_[5827]_  = \new_[5826]_  & \new_[5821]_ ;
  assign \new_[5831]_  = A298 & A202;
  assign \new_[5832]_  = ~A201 & \new_[5831]_ ;
  assign \new_[5836]_  = A302 & ~A301;
  assign \new_[5837]_  = ~A299 & \new_[5836]_ ;
  assign \new_[5838]_  = \new_[5837]_  & \new_[5832]_ ;
  assign \new_[5842]_  = ~A167 & A168;
  assign \new_[5843]_  = A170 & \new_[5842]_ ;
  assign \new_[5847]_  = A200 & ~A199;
  assign \new_[5848]_  = A166 & \new_[5847]_ ;
  assign \new_[5849]_  = \new_[5848]_  & \new_[5843]_ ;
  assign \new_[5853]_  = ~A298 & A202;
  assign \new_[5854]_  = ~A201 & \new_[5853]_ ;
  assign \new_[5858]_  = A302 & ~A301;
  assign \new_[5859]_  = A299 & \new_[5858]_ ;
  assign \new_[5860]_  = \new_[5859]_  & \new_[5854]_ ;
  assign \new_[5864]_  = ~A167 & A168;
  assign \new_[5865]_  = A170 & \new_[5864]_ ;
  assign \new_[5869]_  = A200 & ~A199;
  assign \new_[5870]_  = A166 & \new_[5869]_ ;
  assign \new_[5871]_  = \new_[5870]_  & \new_[5865]_ ;
  assign \new_[5875]_  = ~A298 & A202;
  assign \new_[5876]_  = ~A201 & \new_[5875]_ ;
  assign \new_[5880]_  = ~A302 & A301;
  assign \new_[5881]_  = ~A299 & \new_[5880]_ ;
  assign \new_[5882]_  = \new_[5881]_  & \new_[5876]_ ;
  assign \new_[5886]_  = ~A167 & A168;
  assign \new_[5887]_  = A170 & \new_[5886]_ ;
  assign \new_[5891]_  = A200 & ~A199;
  assign \new_[5892]_  = A166 & \new_[5891]_ ;
  assign \new_[5893]_  = \new_[5892]_  & \new_[5887]_ ;
  assign \new_[5897]_  = A298 & ~A203;
  assign \new_[5898]_  = ~A201 & \new_[5897]_ ;
  assign \new_[5902]_  = ~A302 & A301;
  assign \new_[5903]_  = A299 & \new_[5902]_ ;
  assign \new_[5904]_  = \new_[5903]_  & \new_[5898]_ ;
  assign \new_[5908]_  = ~A167 & A168;
  assign \new_[5909]_  = A170 & \new_[5908]_ ;
  assign \new_[5913]_  = A200 & ~A199;
  assign \new_[5914]_  = A166 & \new_[5913]_ ;
  assign \new_[5915]_  = \new_[5914]_  & \new_[5909]_ ;
  assign \new_[5919]_  = A298 & ~A203;
  assign \new_[5920]_  = ~A201 & \new_[5919]_ ;
  assign \new_[5924]_  = A302 & ~A301;
  assign \new_[5925]_  = ~A299 & \new_[5924]_ ;
  assign \new_[5926]_  = \new_[5925]_  & \new_[5920]_ ;
  assign \new_[5930]_  = ~A167 & A168;
  assign \new_[5931]_  = A170 & \new_[5930]_ ;
  assign \new_[5935]_  = A200 & ~A199;
  assign \new_[5936]_  = A166 & \new_[5935]_ ;
  assign \new_[5937]_  = \new_[5936]_  & \new_[5931]_ ;
  assign \new_[5941]_  = ~A298 & ~A203;
  assign \new_[5942]_  = ~A201 & \new_[5941]_ ;
  assign \new_[5946]_  = A302 & ~A301;
  assign \new_[5947]_  = A299 & \new_[5946]_ ;
  assign \new_[5948]_  = \new_[5947]_  & \new_[5942]_ ;
  assign \new_[5952]_  = ~A167 & A168;
  assign \new_[5953]_  = A170 & \new_[5952]_ ;
  assign \new_[5957]_  = A200 & ~A199;
  assign \new_[5958]_  = A166 & \new_[5957]_ ;
  assign \new_[5959]_  = \new_[5958]_  & \new_[5953]_ ;
  assign \new_[5963]_  = ~A298 & ~A203;
  assign \new_[5964]_  = ~A201 & \new_[5963]_ ;
  assign \new_[5968]_  = ~A302 & A301;
  assign \new_[5969]_  = ~A299 & \new_[5968]_ ;
  assign \new_[5970]_  = \new_[5969]_  & \new_[5964]_ ;
  assign \new_[5974]_  = ~A167 & A168;
  assign \new_[5975]_  = A170 & \new_[5974]_ ;
  assign \new_[5979]_  = ~A200 & A199;
  assign \new_[5980]_  = A166 & \new_[5979]_ ;
  assign \new_[5981]_  = \new_[5980]_  & \new_[5975]_ ;
  assign \new_[5985]_  = A298 & A202;
  assign \new_[5986]_  = ~A201 & \new_[5985]_ ;
  assign \new_[5990]_  = ~A302 & A301;
  assign \new_[5991]_  = A299 & \new_[5990]_ ;
  assign \new_[5992]_  = \new_[5991]_  & \new_[5986]_ ;
  assign \new_[5996]_  = ~A167 & A168;
  assign \new_[5997]_  = A170 & \new_[5996]_ ;
  assign \new_[6001]_  = ~A200 & A199;
  assign \new_[6002]_  = A166 & \new_[6001]_ ;
  assign \new_[6003]_  = \new_[6002]_  & \new_[5997]_ ;
  assign \new_[6007]_  = A298 & A202;
  assign \new_[6008]_  = ~A201 & \new_[6007]_ ;
  assign \new_[6012]_  = A302 & ~A301;
  assign \new_[6013]_  = ~A299 & \new_[6012]_ ;
  assign \new_[6014]_  = \new_[6013]_  & \new_[6008]_ ;
  assign \new_[6018]_  = ~A167 & A168;
  assign \new_[6019]_  = A170 & \new_[6018]_ ;
  assign \new_[6023]_  = ~A200 & A199;
  assign \new_[6024]_  = A166 & \new_[6023]_ ;
  assign \new_[6025]_  = \new_[6024]_  & \new_[6019]_ ;
  assign \new_[6029]_  = ~A298 & A202;
  assign \new_[6030]_  = ~A201 & \new_[6029]_ ;
  assign \new_[6034]_  = A302 & ~A301;
  assign \new_[6035]_  = A299 & \new_[6034]_ ;
  assign \new_[6036]_  = \new_[6035]_  & \new_[6030]_ ;
  assign \new_[6040]_  = ~A167 & A168;
  assign \new_[6041]_  = A170 & \new_[6040]_ ;
  assign \new_[6045]_  = ~A200 & A199;
  assign \new_[6046]_  = A166 & \new_[6045]_ ;
  assign \new_[6047]_  = \new_[6046]_  & \new_[6041]_ ;
  assign \new_[6051]_  = ~A298 & A202;
  assign \new_[6052]_  = ~A201 & \new_[6051]_ ;
  assign \new_[6056]_  = ~A302 & A301;
  assign \new_[6057]_  = ~A299 & \new_[6056]_ ;
  assign \new_[6058]_  = \new_[6057]_  & \new_[6052]_ ;
  assign \new_[6062]_  = ~A167 & A168;
  assign \new_[6063]_  = A170 & \new_[6062]_ ;
  assign \new_[6067]_  = ~A200 & A199;
  assign \new_[6068]_  = A166 & \new_[6067]_ ;
  assign \new_[6069]_  = \new_[6068]_  & \new_[6063]_ ;
  assign \new_[6073]_  = A298 & ~A203;
  assign \new_[6074]_  = ~A201 & \new_[6073]_ ;
  assign \new_[6078]_  = ~A302 & A301;
  assign \new_[6079]_  = A299 & \new_[6078]_ ;
  assign \new_[6080]_  = \new_[6079]_  & \new_[6074]_ ;
  assign \new_[6084]_  = ~A167 & A168;
  assign \new_[6085]_  = A170 & \new_[6084]_ ;
  assign \new_[6089]_  = ~A200 & A199;
  assign \new_[6090]_  = A166 & \new_[6089]_ ;
  assign \new_[6091]_  = \new_[6090]_  & \new_[6085]_ ;
  assign \new_[6095]_  = A298 & ~A203;
  assign \new_[6096]_  = ~A201 & \new_[6095]_ ;
  assign \new_[6100]_  = A302 & ~A301;
  assign \new_[6101]_  = ~A299 & \new_[6100]_ ;
  assign \new_[6102]_  = \new_[6101]_  & \new_[6096]_ ;
  assign \new_[6106]_  = ~A167 & A168;
  assign \new_[6107]_  = A170 & \new_[6106]_ ;
  assign \new_[6111]_  = ~A200 & A199;
  assign \new_[6112]_  = A166 & \new_[6111]_ ;
  assign \new_[6113]_  = \new_[6112]_  & \new_[6107]_ ;
  assign \new_[6117]_  = ~A298 & ~A203;
  assign \new_[6118]_  = ~A201 & \new_[6117]_ ;
  assign \new_[6122]_  = A302 & ~A301;
  assign \new_[6123]_  = A299 & \new_[6122]_ ;
  assign \new_[6124]_  = \new_[6123]_  & \new_[6118]_ ;
  assign \new_[6128]_  = ~A167 & A168;
  assign \new_[6129]_  = A170 & \new_[6128]_ ;
  assign \new_[6133]_  = ~A200 & A199;
  assign \new_[6134]_  = A166 & \new_[6133]_ ;
  assign \new_[6135]_  = \new_[6134]_  & \new_[6129]_ ;
  assign \new_[6139]_  = ~A298 & ~A203;
  assign \new_[6140]_  = ~A201 & \new_[6139]_ ;
  assign \new_[6144]_  = ~A302 & A301;
  assign \new_[6145]_  = ~A299 & \new_[6144]_ ;
  assign \new_[6146]_  = \new_[6145]_  & \new_[6140]_ ;
  assign \new_[6150]_  = ~A167 & A168;
  assign \new_[6151]_  = A169 & \new_[6150]_ ;
  assign \new_[6155]_  = A200 & A199;
  assign \new_[6156]_  = A166 & \new_[6155]_ ;
  assign \new_[6157]_  = \new_[6156]_  & \new_[6151]_ ;
  assign \new_[6161]_  = A298 & ~A202;
  assign \new_[6162]_  = ~A201 & \new_[6161]_ ;
  assign \new_[6166]_  = ~A302 & A301;
  assign \new_[6167]_  = A299 & \new_[6166]_ ;
  assign \new_[6168]_  = \new_[6167]_  & \new_[6162]_ ;
  assign \new_[6172]_  = ~A167 & A168;
  assign \new_[6173]_  = A169 & \new_[6172]_ ;
  assign \new_[6177]_  = A200 & A199;
  assign \new_[6178]_  = A166 & \new_[6177]_ ;
  assign \new_[6179]_  = \new_[6178]_  & \new_[6173]_ ;
  assign \new_[6183]_  = A298 & ~A202;
  assign \new_[6184]_  = ~A201 & \new_[6183]_ ;
  assign \new_[6188]_  = A302 & ~A301;
  assign \new_[6189]_  = ~A299 & \new_[6188]_ ;
  assign \new_[6190]_  = \new_[6189]_  & \new_[6184]_ ;
  assign \new_[6194]_  = ~A167 & A168;
  assign \new_[6195]_  = A169 & \new_[6194]_ ;
  assign \new_[6199]_  = A200 & A199;
  assign \new_[6200]_  = A166 & \new_[6199]_ ;
  assign \new_[6201]_  = \new_[6200]_  & \new_[6195]_ ;
  assign \new_[6205]_  = ~A298 & ~A202;
  assign \new_[6206]_  = ~A201 & \new_[6205]_ ;
  assign \new_[6210]_  = A302 & ~A301;
  assign \new_[6211]_  = A299 & \new_[6210]_ ;
  assign \new_[6212]_  = \new_[6211]_  & \new_[6206]_ ;
  assign \new_[6216]_  = ~A167 & A168;
  assign \new_[6217]_  = A169 & \new_[6216]_ ;
  assign \new_[6221]_  = A200 & A199;
  assign \new_[6222]_  = A166 & \new_[6221]_ ;
  assign \new_[6223]_  = \new_[6222]_  & \new_[6217]_ ;
  assign \new_[6227]_  = ~A298 & ~A202;
  assign \new_[6228]_  = ~A201 & \new_[6227]_ ;
  assign \new_[6232]_  = ~A302 & A301;
  assign \new_[6233]_  = ~A299 & \new_[6232]_ ;
  assign \new_[6234]_  = \new_[6233]_  & \new_[6228]_ ;
  assign \new_[6238]_  = ~A167 & A168;
  assign \new_[6239]_  = A169 & \new_[6238]_ ;
  assign \new_[6243]_  = A200 & A199;
  assign \new_[6244]_  = A166 & \new_[6243]_ ;
  assign \new_[6245]_  = \new_[6244]_  & \new_[6239]_ ;
  assign \new_[6249]_  = A298 & A203;
  assign \new_[6250]_  = ~A201 & \new_[6249]_ ;
  assign \new_[6254]_  = ~A302 & A301;
  assign \new_[6255]_  = A299 & \new_[6254]_ ;
  assign \new_[6256]_  = \new_[6255]_  & \new_[6250]_ ;
  assign \new_[6260]_  = ~A167 & A168;
  assign \new_[6261]_  = A169 & \new_[6260]_ ;
  assign \new_[6265]_  = A200 & A199;
  assign \new_[6266]_  = A166 & \new_[6265]_ ;
  assign \new_[6267]_  = \new_[6266]_  & \new_[6261]_ ;
  assign \new_[6271]_  = A298 & A203;
  assign \new_[6272]_  = ~A201 & \new_[6271]_ ;
  assign \new_[6276]_  = A302 & ~A301;
  assign \new_[6277]_  = ~A299 & \new_[6276]_ ;
  assign \new_[6278]_  = \new_[6277]_  & \new_[6272]_ ;
  assign \new_[6282]_  = ~A167 & A168;
  assign \new_[6283]_  = A169 & \new_[6282]_ ;
  assign \new_[6287]_  = A200 & A199;
  assign \new_[6288]_  = A166 & \new_[6287]_ ;
  assign \new_[6289]_  = \new_[6288]_  & \new_[6283]_ ;
  assign \new_[6293]_  = ~A298 & A203;
  assign \new_[6294]_  = ~A201 & \new_[6293]_ ;
  assign \new_[6298]_  = A302 & ~A301;
  assign \new_[6299]_  = A299 & \new_[6298]_ ;
  assign \new_[6300]_  = \new_[6299]_  & \new_[6294]_ ;
  assign \new_[6304]_  = ~A167 & A168;
  assign \new_[6305]_  = A169 & \new_[6304]_ ;
  assign \new_[6309]_  = A200 & A199;
  assign \new_[6310]_  = A166 & \new_[6309]_ ;
  assign \new_[6311]_  = \new_[6310]_  & \new_[6305]_ ;
  assign \new_[6315]_  = ~A298 & A203;
  assign \new_[6316]_  = ~A201 & \new_[6315]_ ;
  assign \new_[6320]_  = ~A302 & A301;
  assign \new_[6321]_  = ~A299 & \new_[6320]_ ;
  assign \new_[6322]_  = \new_[6321]_  & \new_[6316]_ ;
  assign \new_[6326]_  = ~A167 & A168;
  assign \new_[6327]_  = A169 & \new_[6326]_ ;
  assign \new_[6331]_  = A200 & ~A199;
  assign \new_[6332]_  = A166 & \new_[6331]_ ;
  assign \new_[6333]_  = \new_[6332]_  & \new_[6327]_ ;
  assign \new_[6337]_  = A298 & A202;
  assign \new_[6338]_  = ~A201 & \new_[6337]_ ;
  assign \new_[6342]_  = ~A302 & A301;
  assign \new_[6343]_  = A299 & \new_[6342]_ ;
  assign \new_[6344]_  = \new_[6343]_  & \new_[6338]_ ;
  assign \new_[6348]_  = ~A167 & A168;
  assign \new_[6349]_  = A169 & \new_[6348]_ ;
  assign \new_[6353]_  = A200 & ~A199;
  assign \new_[6354]_  = A166 & \new_[6353]_ ;
  assign \new_[6355]_  = \new_[6354]_  & \new_[6349]_ ;
  assign \new_[6359]_  = A298 & A202;
  assign \new_[6360]_  = ~A201 & \new_[6359]_ ;
  assign \new_[6364]_  = A302 & ~A301;
  assign \new_[6365]_  = ~A299 & \new_[6364]_ ;
  assign \new_[6366]_  = \new_[6365]_  & \new_[6360]_ ;
  assign \new_[6370]_  = ~A167 & A168;
  assign \new_[6371]_  = A169 & \new_[6370]_ ;
  assign \new_[6375]_  = A200 & ~A199;
  assign \new_[6376]_  = A166 & \new_[6375]_ ;
  assign \new_[6377]_  = \new_[6376]_  & \new_[6371]_ ;
  assign \new_[6381]_  = ~A298 & A202;
  assign \new_[6382]_  = ~A201 & \new_[6381]_ ;
  assign \new_[6386]_  = A302 & ~A301;
  assign \new_[6387]_  = A299 & \new_[6386]_ ;
  assign \new_[6388]_  = \new_[6387]_  & \new_[6382]_ ;
  assign \new_[6392]_  = ~A167 & A168;
  assign \new_[6393]_  = A169 & \new_[6392]_ ;
  assign \new_[6397]_  = A200 & ~A199;
  assign \new_[6398]_  = A166 & \new_[6397]_ ;
  assign \new_[6399]_  = \new_[6398]_  & \new_[6393]_ ;
  assign \new_[6403]_  = ~A298 & A202;
  assign \new_[6404]_  = ~A201 & \new_[6403]_ ;
  assign \new_[6408]_  = ~A302 & A301;
  assign \new_[6409]_  = ~A299 & \new_[6408]_ ;
  assign \new_[6410]_  = \new_[6409]_  & \new_[6404]_ ;
  assign \new_[6414]_  = ~A167 & A168;
  assign \new_[6415]_  = A169 & \new_[6414]_ ;
  assign \new_[6419]_  = A200 & ~A199;
  assign \new_[6420]_  = A166 & \new_[6419]_ ;
  assign \new_[6421]_  = \new_[6420]_  & \new_[6415]_ ;
  assign \new_[6425]_  = A298 & ~A203;
  assign \new_[6426]_  = ~A201 & \new_[6425]_ ;
  assign \new_[6430]_  = ~A302 & A301;
  assign \new_[6431]_  = A299 & \new_[6430]_ ;
  assign \new_[6432]_  = \new_[6431]_  & \new_[6426]_ ;
  assign \new_[6436]_  = ~A167 & A168;
  assign \new_[6437]_  = A169 & \new_[6436]_ ;
  assign \new_[6441]_  = A200 & ~A199;
  assign \new_[6442]_  = A166 & \new_[6441]_ ;
  assign \new_[6443]_  = \new_[6442]_  & \new_[6437]_ ;
  assign \new_[6447]_  = A298 & ~A203;
  assign \new_[6448]_  = ~A201 & \new_[6447]_ ;
  assign \new_[6452]_  = A302 & ~A301;
  assign \new_[6453]_  = ~A299 & \new_[6452]_ ;
  assign \new_[6454]_  = \new_[6453]_  & \new_[6448]_ ;
  assign \new_[6458]_  = ~A167 & A168;
  assign \new_[6459]_  = A169 & \new_[6458]_ ;
  assign \new_[6463]_  = A200 & ~A199;
  assign \new_[6464]_  = A166 & \new_[6463]_ ;
  assign \new_[6465]_  = \new_[6464]_  & \new_[6459]_ ;
  assign \new_[6469]_  = ~A298 & ~A203;
  assign \new_[6470]_  = ~A201 & \new_[6469]_ ;
  assign \new_[6474]_  = A302 & ~A301;
  assign \new_[6475]_  = A299 & \new_[6474]_ ;
  assign \new_[6476]_  = \new_[6475]_  & \new_[6470]_ ;
  assign \new_[6480]_  = ~A167 & A168;
  assign \new_[6481]_  = A169 & \new_[6480]_ ;
  assign \new_[6485]_  = A200 & ~A199;
  assign \new_[6486]_  = A166 & \new_[6485]_ ;
  assign \new_[6487]_  = \new_[6486]_  & \new_[6481]_ ;
  assign \new_[6491]_  = ~A298 & ~A203;
  assign \new_[6492]_  = ~A201 & \new_[6491]_ ;
  assign \new_[6496]_  = ~A302 & A301;
  assign \new_[6497]_  = ~A299 & \new_[6496]_ ;
  assign \new_[6498]_  = \new_[6497]_  & \new_[6492]_ ;
  assign \new_[6502]_  = ~A167 & A168;
  assign \new_[6503]_  = A169 & \new_[6502]_ ;
  assign \new_[6507]_  = ~A200 & A199;
  assign \new_[6508]_  = A166 & \new_[6507]_ ;
  assign \new_[6509]_  = \new_[6508]_  & \new_[6503]_ ;
  assign \new_[6513]_  = A298 & A202;
  assign \new_[6514]_  = ~A201 & \new_[6513]_ ;
  assign \new_[6518]_  = ~A302 & A301;
  assign \new_[6519]_  = A299 & \new_[6518]_ ;
  assign \new_[6520]_  = \new_[6519]_  & \new_[6514]_ ;
  assign \new_[6524]_  = ~A167 & A168;
  assign \new_[6525]_  = A169 & \new_[6524]_ ;
  assign \new_[6529]_  = ~A200 & A199;
  assign \new_[6530]_  = A166 & \new_[6529]_ ;
  assign \new_[6531]_  = \new_[6530]_  & \new_[6525]_ ;
  assign \new_[6535]_  = A298 & A202;
  assign \new_[6536]_  = ~A201 & \new_[6535]_ ;
  assign \new_[6540]_  = A302 & ~A301;
  assign \new_[6541]_  = ~A299 & \new_[6540]_ ;
  assign \new_[6542]_  = \new_[6541]_  & \new_[6536]_ ;
  assign \new_[6546]_  = ~A167 & A168;
  assign \new_[6547]_  = A169 & \new_[6546]_ ;
  assign \new_[6551]_  = ~A200 & A199;
  assign \new_[6552]_  = A166 & \new_[6551]_ ;
  assign \new_[6553]_  = \new_[6552]_  & \new_[6547]_ ;
  assign \new_[6557]_  = ~A298 & A202;
  assign \new_[6558]_  = ~A201 & \new_[6557]_ ;
  assign \new_[6562]_  = A302 & ~A301;
  assign \new_[6563]_  = A299 & \new_[6562]_ ;
  assign \new_[6564]_  = \new_[6563]_  & \new_[6558]_ ;
  assign \new_[6568]_  = ~A167 & A168;
  assign \new_[6569]_  = A169 & \new_[6568]_ ;
  assign \new_[6573]_  = ~A200 & A199;
  assign \new_[6574]_  = A166 & \new_[6573]_ ;
  assign \new_[6575]_  = \new_[6574]_  & \new_[6569]_ ;
  assign \new_[6579]_  = ~A298 & A202;
  assign \new_[6580]_  = ~A201 & \new_[6579]_ ;
  assign \new_[6584]_  = ~A302 & A301;
  assign \new_[6585]_  = ~A299 & \new_[6584]_ ;
  assign \new_[6586]_  = \new_[6585]_  & \new_[6580]_ ;
  assign \new_[6590]_  = ~A167 & A168;
  assign \new_[6591]_  = A169 & \new_[6590]_ ;
  assign \new_[6595]_  = ~A200 & A199;
  assign \new_[6596]_  = A166 & \new_[6595]_ ;
  assign \new_[6597]_  = \new_[6596]_  & \new_[6591]_ ;
  assign \new_[6601]_  = A298 & ~A203;
  assign \new_[6602]_  = ~A201 & \new_[6601]_ ;
  assign \new_[6606]_  = ~A302 & A301;
  assign \new_[6607]_  = A299 & \new_[6606]_ ;
  assign \new_[6608]_  = \new_[6607]_  & \new_[6602]_ ;
  assign \new_[6612]_  = ~A167 & A168;
  assign \new_[6613]_  = A169 & \new_[6612]_ ;
  assign \new_[6617]_  = ~A200 & A199;
  assign \new_[6618]_  = A166 & \new_[6617]_ ;
  assign \new_[6619]_  = \new_[6618]_  & \new_[6613]_ ;
  assign \new_[6623]_  = A298 & ~A203;
  assign \new_[6624]_  = ~A201 & \new_[6623]_ ;
  assign \new_[6628]_  = A302 & ~A301;
  assign \new_[6629]_  = ~A299 & \new_[6628]_ ;
  assign \new_[6630]_  = \new_[6629]_  & \new_[6624]_ ;
  assign \new_[6634]_  = ~A167 & A168;
  assign \new_[6635]_  = A169 & \new_[6634]_ ;
  assign \new_[6639]_  = ~A200 & A199;
  assign \new_[6640]_  = A166 & \new_[6639]_ ;
  assign \new_[6641]_  = \new_[6640]_  & \new_[6635]_ ;
  assign \new_[6645]_  = ~A298 & ~A203;
  assign \new_[6646]_  = ~A201 & \new_[6645]_ ;
  assign \new_[6650]_  = A302 & ~A301;
  assign \new_[6651]_  = A299 & \new_[6650]_ ;
  assign \new_[6652]_  = \new_[6651]_  & \new_[6646]_ ;
  assign \new_[6656]_  = ~A167 & A168;
  assign \new_[6657]_  = A169 & \new_[6656]_ ;
  assign \new_[6661]_  = ~A200 & A199;
  assign \new_[6662]_  = A166 & \new_[6661]_ ;
  assign \new_[6663]_  = \new_[6662]_  & \new_[6657]_ ;
  assign \new_[6667]_  = ~A298 & ~A203;
  assign \new_[6668]_  = ~A201 & \new_[6667]_ ;
  assign \new_[6672]_  = ~A302 & A301;
  assign \new_[6673]_  = ~A299 & \new_[6672]_ ;
  assign \new_[6674]_  = \new_[6673]_  & \new_[6668]_ ;
endmodule


