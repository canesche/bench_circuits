module top ( 
    pa1, pb2, pp, pa0, pc2, pq, pb0, pc1, pr, pa2, pb1, pc0, ps, pd0, pe1,
    pf2, pt, pd1, pe0, pg2, pu, pd2, pf0, pg1, pv, pe2, pf1, pg0, pw, ph0,
    pi1, px, ph1, pi0, py, ph2, pj0, pk1, pz, pj1, pk0, pl0, pm1, pl1, pm0,
    pn0, po1, pn1, po0, pp0, pq1, pa, pp1, pq0, pb, pr0, ps1, pr1, ps0, pd,
    pt0, pu1, pe, pt1, pu0, pf, pv0, pw1, pg, pv1, pw0, ph, px0, py1, pi,
    px1, py0, pj, pz0, pk, pz1, pl, pm, pn, po,
    pc3, pd4, pb3, pe4, pa3, pf4, pg4, pg3, pa4, pf3, pb4, pe3, pc4, pd3,
    pj2, pk3, pl4, pj3, pk2, pm4, pi3, pn4, ph3, pi2, po4, ph4, pn2, po3,
    pi4, pn3, po2, pj4, pl2, pm3, pk4, pl3, pm2, pr2, ps3, pt4, pr3, ps2,
    pu4, pp2, pq3, pv4, pp3, pq2, pp4, pv2, pw3, pq4, pv3, pw2, pr4, pt2,
    pu3, ps4, pt3, pu2, pz2, pz3, px2, py3, px3, py2  );
  input  pa1, pb2, pp, pa0, pc2, pq, pb0, pc1, pr, pa2, pb1, pc0, ps,
    pd0, pe1, pf2, pt, pd1, pe0, pg2, pu, pd2, pf0, pg1, pv, pe2, pf1, pg0,
    pw, ph0, pi1, px, ph1, pi0, py, ph2, pj0, pk1, pz, pj1, pk0, pl0, pm1,
    pl1, pm0, pn0, po1, pn1, po0, pp0, pq1, pa, pp1, pq0, pb, pr0, ps1,
    pr1, ps0, pd, pt0, pu1, pe, pt1, pu0, pf, pv0, pw1, pg, pv1, pw0, ph,
    px0, py1, pi, px1, py0, pj, pz0, pk, pz1, pl, pm, pn, po;
  output pc3, pd4, pb3, pe4, pa3, pf4, pg4, pg3, pa4, pf3, pb4, pe3, pc4, pd3,
    pj2, pk3, pl4, pj3, pk2, pm4, pi3, pn4, ph3, pi2, po4, ph4, pn2, po3,
    pi4, pn3, po2, pj4, pl2, pm3, pk4, pl3, pm2, pr2, ps3, pt4, pr3, ps2,
    pu4, pp2, pq3, pv4, pp3, pq2, pp4, pv2, pw3, pq4, pv3, pw2, pr4, pt2,
    pu3, ps4, pt3, pu2, pz2, pz3, px2, py3, px3, py2;
  wire new_n152_, new_n153_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n195_, new_n196_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n206_, new_n207_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n214_, new_n215_, new_n216_, new_n217_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n251_,
    new_n252_, new_n253_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n279_, new_n280_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n288_, new_n289_,
    new_n290_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n318_, new_n319_, new_n322_, new_n323_, new_n325_, new_n326_,
    new_n327_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n348_, new_n349_, new_n350_, new_n351_, new_n353_,
    new_n354_, new_n357_, new_n358_, new_n359_, new_n360_, new_n363_,
    new_n364_, new_n366_, new_n367_, new_n368_, new_n369_, new_n372_,
    new_n373_, new_n376_, new_n377_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n387_, new_n388_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n395_, new_n396_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n405_, new_n406_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n422_,
    new_n423_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n443_, new_n444_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n456_, new_n457_, new_n460_,
    new_n463_, new_n464_, new_n466_, new_n467_, new_n470_, new_n471_,
    new_n475_, new_n476_;
  assign new_n152_ = pp0 & pu0;
  assign new_n153_ = pn0 & ~pp0;
  assign pc3 = new_n152_ | new_n153_;
  assign new_n155_ = pe2 & ~ph2;
  assign new_n156_ = ~pe2 & ph2;
  assign new_n157_ = ~new_n155_ & ~new_n156_;
  assign new_n158_ = ~pb2 & pa2;
  assign new_n159_ = py1 & new_n157_;
  assign new_n160_ = ~pb & new_n159_;
  assign new_n161_ = pc2 & new_n160_;
  assign new_n162_ = new_n158_ & new_n161_;
  assign new_n163_ = ~pf2 & ~pe2;
  assign new_n164_ = ~ph2 & new_n163_;
  assign new_n165_ = ~pg2 & new_n164_;
  assign new_n166_ = ~new_n157_ & new_n165_;
  assign new_n167_ = ~pb & new_n166_;
  assign new_n168_ = pc2 & new_n167_;
  assign new_n169_ = new_n158_ & new_n168_;
  assign new_n170_ = pp1 & new_n169_;
  assign new_n171_ = pd2 & new_n170_;
  assign new_n172_ = pq0 & new_n171_;
  assign new_n173_ = pb2 & ~pc2;
  assign new_n174_ = ~pb & new_n173_;
  assign pl2 = pb1 & new_n174_;
  assign new_n176_ = ~pa2 & pf;
  assign new_n177_ = pl2 & new_n176_;
  assign new_n178_ = pq & new_n177_;
  assign new_n179_ = pq1 & new_n157_;
  assign new_n180_ = ~pb & new_n179_;
  assign new_n181_ = pc2 & new_n180_;
  assign new_n182_ = new_n158_ & new_n181_;
  assign new_n183_ = ~pb & new_n176_;
  assign new_n184_ = new_n173_ & new_n183_;
  assign new_n185_ = ~pb1 & new_n184_;
  assign new_n186_ = pi & new_n185_;
  assign new_n187_ = ~pp1 & new_n169_;
  assign new_n188_ = pd2 & new_n187_;
  assign new_n189_ = ~pq0 & new_n188_;
  assign new_n190_ = ~new_n182_ & ~new_n186_;
  assign new_n191_ = ~new_n189_ & new_n190_;
  assign new_n192_ = ~new_n162_ & ~new_n172_;
  assign new_n193_ = ~new_n178_ & new_n192_;
  assign pd4 = ~new_n191_ | ~new_n193_;
  assign new_n195_ = pp0 & pv0;
  assign new_n196_ = pm0 & ~pp0;
  assign pb3 = new_n195_ | new_n196_;
  assign new_n198_ = pj & new_n185_;
  assign new_n199_ = ~pb & new_n158_;
  assign new_n200_ = pc2 & new_n199_;
  assign new_n201_ = new_n157_ & new_n200_;
  assign new_n202_ = pr1 & new_n201_;
  assign new_n203_ = pr & new_n177_;
  assign new_n204_ = ~new_n198_ & ~new_n202_;
  assign pe4 = new_n203_ | ~new_n204_;
  assign new_n206_ = pp0 & pw0;
  assign new_n207_ = pl0 & ~pp0;
  assign pa3 = new_n206_ | new_n207_;
  assign new_n209_ = pk & new_n185_;
  assign new_n210_ = ps1 & new_n201_;
  assign new_n211_ = ps & new_n177_;
  assign new_n212_ = ~new_n209_ & ~new_n210_;
  assign pf4 = new_n211_ | ~new_n212_;
  assign new_n214_ = pl & new_n185_;
  assign new_n215_ = pt1 & new_n201_;
  assign new_n216_ = pt & new_n177_;
  assign new_n217_ = ~new_n214_ & ~new_n215_;
  assign pg4 = new_n216_ | ~new_n217_;
  assign new_n219_ = pb2 & pa2;
  assign new_n220_ = ~ps0 & new_n219_;
  assign new_n221_ = pg & new_n220_;
  assign new_n222_ = ~pf & new_n221_;
  assign new_n223_ = ~pb & new_n222_;
  assign new_n224_ = ~pc2 & ~ps0;
  assign new_n225_ = pg & new_n224_;
  assign new_n226_ = ~pf & new_n225_;
  assign new_n227_ = ~pb & new_n226_;
  assign pg3 = new_n223_ | new_n227_;
  assign new_n229_ = pf2 & pe2;
  assign new_n230_ = ~new_n163_ & ~new_n229_;
  assign new_n231_ = ~pg2 & new_n230_;
  assign new_n232_ = pg2 & ~new_n230_;
  assign new_n233_ = ~new_n231_ & ~new_n232_;
  assign new_n234_ = ph2 & new_n233_;
  assign new_n235_ = ~ph2 & ~new_n233_;
  assign new_n236_ = ~new_n234_ & ~new_n235_;
  assign new_n237_ = pc2 & ~pb;
  assign new_n238_ = ~pf & new_n219_;
  assign new_n239_ = new_n237_ & new_n238_;
  assign new_n240_ = pr0 & ~new_n236_;
  assign new_n241_ = new_n239_ & new_n240_;
  assign new_n242_ = ~pr0 & new_n230_;
  assign new_n243_ = ~ph2 & new_n242_;
  assign new_n244_ = new_n239_ & new_n243_;
  assign new_n245_ = ~pr0 & ~new_n230_;
  assign new_n246_ = ph2 & new_n245_;
  assign new_n247_ = new_n239_ & new_n246_;
  assign new_n248_ = ~new_n244_ & ~new_n247_;
  assign new_n249_ = ~new_n241_ & new_n248_;
  assign pa4 = pl1 & ~new_n249_;
  assign new_n251_ = ~pc2 & ~pf;
  assign new_n252_ = pg & new_n251_;
  assign new_n253_ = ~pb & ~new_n252_;
  assign pf3 = ~pa | ~new_n253_;
  assign pb4 = pm1 & ~new_n249_;
  assign new_n256_ = pb2 & ~pa2;
  assign new_n257_ = py1 & new_n256_;
  assign new_n258_ = new_n237_ & new_n257_;
  assign new_n259_ = pp1 & new_n158_;
  assign new_n260_ = new_n237_ & new_n259_;
  assign pk2 = new_n258_ | new_n260_;
  assign new_n262_ = new_n157_ & pk2;
  assign new_n263_ = ~pq0 & new_n262_;
  assign new_n264_ = pd2 & ~px1;
  assign new_n265_ = new_n229_ & new_n264_;
  assign new_n266_ = ~pg2 & ps0;
  assign new_n267_ = ph2 & new_n266_;
  assign new_n268_ = new_n265_ & new_n267_;
  assign new_n269_ = pa2 & ~new_n268_;
  assign new_n270_ = ~pr0 & new_n269_;
  assign new_n271_ = pb2 & pf;
  assign new_n272_ = ~pb & new_n270_;
  assign new_n273_ = new_n271_ & new_n272_;
  assign new_n274_ = ~pc2 & ~pb;
  assign new_n275_ = new_n271_ & new_n274_;
  assign new_n276_ = ~new_n273_ & ~new_n275_;
  assign pe3 = new_n263_ | ~new_n276_;
  assign pc4 = pn1 & ~new_n249_;
  assign new_n279_ = pp0 & pt0;
  assign new_n280_ = po0 & ~pp0;
  assign pd3 = new_n279_ | new_n280_;
  assign new_n282_ = ~pb & new_n219_;
  assign new_n283_ = ~pb2 & ~pa2;
  assign new_n284_ = ~pb & new_n283_;
  assign new_n285_ = ~new_n282_ & ~new_n284_;
  assign pj2 = new_n274_ | ~new_n285_;
  assign pk3 = pv0 & ~new_n248_;
  assign new_n288_ = new_n163_ & new_n239_;
  assign new_n289_ = pg2 & new_n288_;
  assign new_n290_ = ph2 & new_n289_;
  assign pl4 = ~pd2 & new_n290_;
  assign pj3 = pu0 & ~new_n248_;
  assign new_n293_ = pz1 & ~new_n219_;
  assign new_n294_ = new_n157_ & new_n293_;
  assign new_n295_ = pc2 & new_n294_;
  assign new_n296_ = ~pd2 & ~new_n219_;
  assign new_n297_ = ~new_n157_ & new_n296_;
  assign new_n298_ = pc2 & new_n297_;
  assign new_n299_ = ~pq0 & ~py1;
  assign new_n300_ = pc2 & new_n299_;
  assign new_n301_ = ~new_n157_ & new_n300_;
  assign new_n302_ = ~pa2 & new_n301_;
  assign new_n303_ = ~new_n165_ & ~new_n219_;
  assign new_n304_ = ~new_n157_ & new_n303_;
  assign new_n305_ = pc2 & new_n304_;
  assign new_n306_ = pq0 & py1;
  assign new_n307_ = pc2 & new_n306_;
  assign new_n308_ = ~new_n157_ & new_n307_;
  assign new_n309_ = ~pa2 & new_n308_;
  assign new_n310_ = ~new_n305_ & ~new_n309_;
  assign new_n311_ = ~pb & ~new_n302_;
  assign new_n312_ = new_n310_ & new_n311_;
  assign new_n313_ = ~new_n295_ & ~new_n298_;
  assign new_n314_ = pa & ~new_n283_;
  assign new_n315_ = new_n313_ & new_n314_;
  assign pm4 = ~new_n312_ | ~new_n315_;
  assign pi3 = pt0 & ~new_n248_;
  assign new_n318_ = ~pb & pe;
  assign new_n319_ = ~pd & new_n318_;
  assign pn4 = pa & new_n319_;
  assign ph3 = pg & ~new_n248_;
  assign new_n322_ = pb1 & pp0;
  assign new_n323_ = ~pb & ~new_n219_;
  assign pm2 = new_n237_ | new_n323_;
  assign new_n325_ = pp0 & pm2;
  assign new_n326_ = ~pp0 & ph;
  assign new_n327_ = ~new_n322_ & ~new_n325_;
  assign pi2 = new_n326_ | ~new_n327_;
  assign new_n329_ = ~pr0 & new_n158_;
  assign new_n330_ = ~pc2 & new_n329_;
  assign new_n331_ = pp0 & new_n330_;
  assign new_n332_ = ~pb & new_n331_;
  assign new_n333_ = ~pr0 & new_n268_;
  assign new_n334_ = new_n237_ & new_n333_;
  assign new_n335_ = pa2 & new_n334_;
  assign new_n336_ = new_n271_ & new_n335_;
  assign new_n337_ = ~pc2 & new_n256_;
  assign new_n338_ = ~pb & new_n337_;
  assign new_n339_ = ~pp0 & pr0;
  assign new_n340_ = new_n237_ & new_n339_;
  assign new_n341_ = pa2 & new_n340_;
  assign new_n342_ = new_n271_ & new_n341_;
  assign new_n343_ = ~pb & new_n251_;
  assign new_n344_ = ~new_n342_ & ~new_n343_;
  assign new_n345_ = ~new_n332_ & ~new_n336_;
  assign new_n346_ = ~new_n338_ & new_n345_;
  assign po4 = ~new_n344_ | ~new_n346_;
  assign new_n348_ = pm & new_n185_;
  assign new_n349_ = pu1 & new_n201_;
  assign new_n350_ = pu & new_n177_;
  assign new_n351_ = ~new_n348_ & ~new_n349_;
  assign ph4 = new_n350_ | ~new_n351_;
  assign new_n353_ = po1 & pp0;
  assign new_n354_ = py & ~pp0;
  assign pn2 = new_n353_ | new_n354_;
  assign po3 = pz0 & ~new_n248_;
  assign new_n357_ = pn & new_n185_;
  assign new_n358_ = pv1 & new_n201_;
  assign new_n359_ = pv & new_n177_;
  assign new_n360_ = ~new_n357_ & ~new_n358_;
  assign pi4 = new_n359_ | ~new_n360_;
  assign pn3 = py0 & ~new_n248_;
  assign new_n363_ = pn1 & pp0;
  assign new_n364_ = pz & ~pp0;
  assign po2 = new_n363_ | new_n364_;
  assign new_n366_ = po & new_n185_;
  assign new_n367_ = pw1 & new_n201_;
  assign new_n368_ = pw & new_n177_;
  assign new_n369_ = ~new_n366_ & ~new_n367_;
  assign pj4 = new_n368_ | ~new_n369_;
  assign pm3 = px0 & ~new_n248_;
  assign new_n372_ = pp & new_n185_;
  assign new_n373_ = px & new_n177_;
  assign pk4 = new_n372_ | new_n373_;
  assign pl3 = pw0 & ~new_n248_;
  assign new_n376_ = pk1 & pp0;
  assign new_n377_ = pc0 & ~pp0;
  assign pr2 = new_n376_ | new_n377_;
  assign ps3 = pd1 & ~new_n249_;
  assign new_n380_ = new_n157_ & new_n158_;
  assign new_n381_ = new_n157_ & new_n256_;
  assign new_n382_ = ~new_n380_ & ~new_n381_;
  assign new_n383_ = ~new_n238_ & new_n382_;
  assign new_n384_ = new_n237_ & ~new_n383_;
  assign pt4 = pf2 & new_n384_;
  assign pr3 = pc1 & ~new_n249_;
  assign new_n387_ = pj1 & pp0;
  assign new_n388_ = pd0 & ~pp0;
  assign ps2 = new_n387_ | new_n388_;
  assign new_n390_ = ~pa2 & new_n173_;
  assign new_n391_ = pf & new_n390_;
  assign new_n392_ = ~pb & new_n391_;
  assign new_n393_ = pg2 & new_n384_;
  assign pu4 = new_n392_ | new_n393_;
  assign new_n395_ = pm1 & pp0;
  assign new_n396_ = pa0 & ~pp0;
  assign pp2 = new_n395_ | new_n396_;
  assign pq3 = pb1 & ~new_n249_;
  assign pv4 = ph2 & new_n384_;
  assign new_n400_ = pr0 & new_n239_;
  assign new_n401_ = ~new_n236_ & new_n400_;
  assign new_n402_ = pg & new_n401_;
  assign new_n403_ = pa1 & ~new_n248_;
  assign pp3 = new_n402_ | new_n403_;
  assign new_n405_ = pl1 & pp0;
  assign new_n406_ = pb0 & ~pp0;
  assign pq2 = new_n405_ | new_n406_;
  assign new_n408_ = pa2 & new_n271_;
  assign new_n409_ = pp0 & new_n408_;
  assign new_n410_ = ~pb & new_n409_;
  assign new_n411_ = pa2 & new_n173_;
  assign new_n412_ = ~pb & new_n411_;
  assign new_n413_ = ~pc2 & pa2;
  assign new_n414_ = pp0 & new_n413_;
  assign new_n415_ = ~pb & new_n414_;
  assign new_n416_ = new_n270_ & new_n271_;
  assign new_n417_ = ~new_n251_ & ~new_n416_;
  assign new_n418_ = ~pb & ~new_n417_;
  assign new_n419_ = ~new_n410_ & ~new_n412_;
  assign new_n420_ = ~new_n415_ & ~new_n418_;
  assign pp4 = ~new_n419_ | ~new_n420_;
  assign new_n422_ = pg1 & pp0;
  assign new_n423_ = pg0 & ~pp0;
  assign pv2 = new_n422_ | new_n423_;
  assign pw3 = ph1 & ~new_n249_;
  assign new_n426_ = ~new_n157_ & new_n256_;
  assign new_n427_ = ~pd2 & new_n426_;
  assign new_n428_ = ~pb & new_n427_;
  assign new_n429_ = pc2 & new_n158_;
  assign new_n430_ = ~new_n157_ & new_n429_;
  assign new_n431_ = ~new_n165_ & new_n430_;
  assign new_n432_ = ~pb & new_n431_;
  assign new_n433_ = ~new_n165_ & new_n426_;
  assign new_n434_ = ~pb & new_n433_;
  assign new_n435_ = ~pd2 & new_n430_;
  assign new_n436_ = ~pb & new_n435_;
  assign new_n437_ = ~new_n418_ & ~new_n434_;
  assign new_n438_ = ~new_n436_ & new_n437_;
  assign new_n439_ = ~new_n428_ & ~new_n432_;
  assign new_n440_ = ~new_n174_ & new_n439_;
  assign pq4 = ~new_n438_ | ~new_n440_;
  assign pv3 = pg1 & ~new_n249_;
  assign new_n443_ = pa1 & pp0;
  assign new_n444_ = ph0 & ~pp0;
  assign pw2 = new_n443_ | new_n444_;
  assign new_n446_ = pd2 & new_n158_;
  assign new_n447_ = new_n165_ & new_n446_;
  assign new_n448_ = new_n237_ & new_n447_;
  assign new_n449_ = pd2 & new_n256_;
  assign new_n450_ = new_n165_ & new_n449_;
  assign new_n451_ = new_n237_ & new_n450_;
  assign new_n452_ = pd2 & ~new_n383_;
  assign new_n453_ = new_n237_ & new_n452_;
  assign new_n454_ = ~new_n448_ & ~new_n451_;
  assign pr4 = new_n453_ | ~new_n454_;
  assign new_n456_ = pi1 & pp0;
  assign new_n457_ = pe0 & ~pp0;
  assign pt2 = new_n456_ | new_n457_;
  assign pu3 = pf1 & ~new_n249_;
  assign new_n460_ = pe2 & new_n384_;
  assign ps4 = ~new_n276_ | new_n460_;
  assign pt3 = pe1 & ~new_n249_;
  assign new_n463_ = ph1 & pp0;
  assign new_n464_ = pf0 & ~pp0;
  assign pu2 = new_n463_ | new_n464_;
  assign new_n466_ = pp0 & px0;
  assign new_n467_ = pk0 & ~pp0;
  assign pz2 = new_n466_ | new_n467_;
  assign pz3 = pk1 & ~new_n249_;
  assign new_n470_ = pp0 & pz0;
  assign new_n471_ = pi0 & ~pp0;
  assign px2 = new_n470_ | new_n471_;
  assign py3 = pj1 & ~new_n249_;
  assign px3 = pi1 & ~new_n249_;
  assign new_n475_ = pp0 & py0;
  assign new_n476_ = pj0 & ~pp0;
  assign py2 = new_n475_ | new_n476_;
endmodule

