module top ( 
    pp, pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw, ph0,
    px, pi0, py, pj0, pz, pk0, pl0, pm0, pn0, po0, pp0, pa, pq0, pr0, pc,
    ps0, pd, pt0, pe, pu0, pf, pv0, pg, ph, pi, pj, pk, pl, pm, pn, po,
    pa1, pb2, pc2, pc1, pa2, pb1, pe1, pf2, pd1, pd2, pg1, pe2, pf1, pi1,
    ph1, pk1, pj1, pm1, pl1, po1, pn1, pq1, pp1, ps1, pr1, pu1, pt1, pw1,
    pv1, pw0, px0, py1, px1, py0, pz0, pz1  );
  input  pp, pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0,
    pw, ph0, px, pi0, py, pj0, pz, pk0, pl0, pm0, pn0, po0, pp0, pa, pq0,
    pr0, pc, ps0, pd, pt0, pe, pu0, pf, pv0, pg, ph, pi, pj, pk, pl, pm,
    pn, po;
  output pa1, pb2, pc2, pc1, pa2, pb1, pe1, pf2, pd1, pd2, pg1, pe2, pf1, pi1,
    ph1, pk1, pj1, pm1, pl1, po1, pn1, pq1, pp1, ps1, pr1, pu1, pt1, pw1,
    pv1, pw0, px0, py1, px1, py0, pz0, pz1;
  wire new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_,
    new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_,
    new_n99_, new_n100_, new_n101_, new_n102_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n142_, new_n143_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n148_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_;
  assign new_n84_ = pd & ~pl;
  assign new_n85_ = pi & new_n84_;
  assign new_n86_ = pq & pd;
  assign new_n87_ = ~pl & new_n86_;
  assign new_n88_ = pq & ~pl;
  assign new_n89_ = ~pi & new_n88_;
  assign new_n90_ = ~new_n85_ & ~new_n87_;
  assign pa1 = new_n89_ | ~new_n90_;
  assign new_n92_ = ps0 & ~pl;
  assign new_n93_ = ~pp & new_n92_;
  assign new_n94_ = pk & new_n93_;
  assign new_n95_ = pp & pr0;
  assign new_n96_ = ~pl & new_n95_;
  assign new_n97_ = pr0 & ps0;
  assign new_n98_ = ~pl & new_n97_;
  assign new_n99_ = pr0 & ~pl;
  assign new_n100_ = ~pk & new_n99_;
  assign new_n101_ = ~new_n94_ & ~new_n96_;
  assign new_n102_ = ~new_n98_ & ~new_n100_;
  assign pb2 = ~new_n101_ | ~new_n102_;
  assign new_n104_ = pt0 & ~pl;
  assign new_n105_ = ~pp & new_n104_;
  assign new_n106_ = pk & new_n105_;
  assign new_n107_ = pp & ps0;
  assign new_n108_ = ~pl & new_n107_;
  assign new_n109_ = ps0 & pt0;
  assign new_n110_ = ~pl & new_n109_;
  assign new_n111_ = ~pk & new_n92_;
  assign new_n112_ = ~new_n106_ & ~new_n108_;
  assign new_n113_ = ~new_n110_ & ~new_n111_;
  assign pc2 = ~new_n112_ | ~new_n113_;
  assign new_n115_ = ps & ~pl;
  assign new_n116_ = ~pj & new_n115_;
  assign new_n117_ = ps & pt;
  assign new_n118_ = ~pl & new_n117_;
  assign new_n119_ = pt & ~pl;
  assign new_n120_ = pj & new_n119_;
  assign new_n121_ = ~new_n116_ & ~new_n118_;
  assign pc1 = new_n120_ | ~new_n121_;
  assign new_n123_ = ~pp & new_n99_;
  assign new_n124_ = pk & new_n123_;
  assign new_n125_ = pp & pq0;
  assign new_n126_ = ~pl & new_n125_;
  assign new_n127_ = pq0 & pr0;
  assign new_n128_ = ~pl & new_n127_;
  assign new_n129_ = pq0 & ~pl;
  assign new_n130_ = ~pk & new_n129_;
  assign new_n131_ = ~new_n124_ & ~new_n126_;
  assign new_n132_ = ~new_n128_ & ~new_n130_;
  assign pa2 = ~new_n131_ | ~new_n132_;
  assign new_n134_ = pe & ~pl;
  assign new_n135_ = pi & new_n134_;
  assign new_n136_ = pr & pe;
  assign new_n137_ = ~pl & new_n136_;
  assign new_n138_ = pr & ~pl;
  assign new_n139_ = ~pi & new_n138_;
  assign new_n140_ = ~new_n135_ & ~new_n137_;
  assign pb1 = new_n139_ | ~new_n140_;
  assign new_n142_ = pu & ~pl;
  assign new_n143_ = ~pj & new_n142_;
  assign new_n144_ = pu & pv;
  assign new_n145_ = ~pl & new_n144_;
  assign new_n146_ = pv & ~pl;
  assign new_n147_ = pj & new_n146_;
  assign new_n148_ = ~new_n143_ & ~new_n145_;
  assign pe1 = new_n147_ | ~new_n148_;
  assign new_n150_ = ~pp & pk;
  assign new_n151_ = ~pl & new_n150_;
  assign new_n152_ = pa & new_n151_;
  assign new_n153_ = pv0 & ~pl;
  assign new_n154_ = ~pk & new_n153_;
  assign new_n155_ = pp & pv0;
  assign new_n156_ = ~pl & new_n155_;
  assign new_n157_ = pa & new_n153_;
  assign new_n158_ = ~new_n152_ & ~new_n154_;
  assign new_n159_ = ~new_n156_ & ~new_n157_;
  assign pf2 = ~new_n158_ | ~new_n159_;
  assign new_n161_ = ~pj & new_n119_;
  assign new_n162_ = pt & pu;
  assign new_n163_ = ~pl & new_n162_;
  assign new_n164_ = pj & new_n142_;
  assign new_n165_ = ~new_n161_ & ~new_n163_;
  assign pd1 = new_n164_ | ~new_n165_;
  assign new_n167_ = pu0 & ~pl;
  assign new_n168_ = ~pp & new_n167_;
  assign new_n169_ = pk & new_n168_;
  assign new_n170_ = pp & pt0;
  assign new_n171_ = ~pl & new_n170_;
  assign new_n172_ = pt0 & pu0;
  assign new_n173_ = ~pl & new_n172_;
  assign new_n174_ = ~pk & new_n104_;
  assign new_n175_ = ~new_n169_ & ~new_n171_;
  assign new_n176_ = ~new_n173_ & ~new_n174_;
  assign pd2 = ~new_n175_ | ~new_n176_;
  assign new_n178_ = pw & ~pl;
  assign new_n179_ = ~pj & new_n178_;
  assign new_n180_ = pw & px;
  assign new_n181_ = ~pl & new_n180_;
  assign new_n182_ = px & ~pl;
  assign new_n183_ = pj & new_n182_;
  assign new_n184_ = ~new_n179_ & ~new_n181_;
  assign pg1 = new_n183_ | ~new_n184_;
  assign new_n186_ = ~pp & new_n153_;
  assign new_n187_ = pk & new_n186_;
  assign new_n188_ = pp & pu0;
  assign new_n189_ = ~pl & new_n188_;
  assign new_n190_ = pu0 & pv0;
  assign new_n191_ = ~pl & new_n190_;
  assign new_n192_ = ~pk & new_n167_;
  assign new_n193_ = ~new_n187_ & ~new_n189_;
  assign new_n194_ = ~new_n191_ & ~new_n192_;
  assign pe2 = ~new_n193_ | ~new_n194_;
  assign new_n196_ = ~pj & new_n146_;
  assign new_n197_ = pv & pw;
  assign new_n198_ = ~pl & new_n197_;
  assign new_n199_ = pj & new_n178_;
  assign new_n200_ = ~new_n196_ & ~new_n198_;
  assign pf1 = new_n199_ | ~new_n200_;
  assign new_n202_ = py & ~pl;
  assign new_n203_ = ~pj & new_n202_;
  assign new_n204_ = py & pz;
  assign new_n205_ = ~pl & new_n204_;
  assign new_n206_ = pz & ~pl;
  assign new_n207_ = pj & new_n206_;
  assign new_n208_ = ~new_n203_ & ~new_n205_;
  assign pi1 = new_n207_ | ~new_n208_;
  assign new_n210_ = ~pj & new_n182_;
  assign new_n211_ = px & py;
  assign new_n212_ = ~pl & new_n211_;
  assign new_n213_ = pj & new_n202_;
  assign new_n214_ = ~new_n210_ & ~new_n212_;
  assign ph1 = new_n213_ | ~new_n214_;
  assign new_n216_ = pa0 & ~pl;
  assign new_n217_ = ~pj & new_n216_;
  assign new_n218_ = pa0 & pb0;
  assign new_n219_ = ~pl & new_n218_;
  assign new_n220_ = pb0 & ~pl;
  assign new_n221_ = pj & new_n220_;
  assign new_n222_ = ~new_n217_ & ~new_n219_;
  assign pk1 = new_n221_ | ~new_n222_;
  assign new_n224_ = ~pj & new_n206_;
  assign new_n225_ = pa0 & pz;
  assign new_n226_ = ~pl & new_n225_;
  assign new_n227_ = pj & new_n216_;
  assign new_n228_ = ~new_n224_ & ~new_n226_;
  assign pj1 = new_n227_ | ~new_n228_;
  assign new_n230_ = pc0 & ~pl;
  assign new_n231_ = ~pj & new_n230_;
  assign new_n232_ = pc0 & pd0;
  assign new_n233_ = ~pl & new_n232_;
  assign new_n234_ = pd0 & ~pl;
  assign new_n235_ = pj & new_n234_;
  assign new_n236_ = ~new_n231_ & ~new_n233_;
  assign pm1 = new_n235_ | ~new_n236_;
  assign new_n238_ = ~pj & new_n220_;
  assign new_n239_ = pb0 & pc0;
  assign new_n240_ = ~pl & new_n239_;
  assign new_n241_ = pj & new_n230_;
  assign new_n242_ = ~new_n238_ & ~new_n240_;
  assign pl1 = new_n241_ | ~new_n242_;
  assign new_n244_ = pe0 & ~pl;
  assign new_n245_ = ~pj & new_n244_;
  assign new_n246_ = pe0 & pf0;
  assign new_n247_ = ~pl & new_n246_;
  assign new_n248_ = pf0 & ~pl;
  assign new_n249_ = pj & new_n248_;
  assign new_n250_ = ~new_n245_ & ~new_n247_;
  assign po1 = new_n249_ | ~new_n250_;
  assign new_n252_ = ~pj & new_n234_;
  assign new_n253_ = pd0 & pe0;
  assign new_n254_ = ~pl & new_n253_;
  assign new_n255_ = pj & new_n244_;
  assign new_n256_ = ~new_n252_ & ~new_n254_;
  assign pn1 = new_n255_ | ~new_n256_;
  assign new_n258_ = pg0 & ~pl;
  assign new_n259_ = ~pk & new_n258_;
  assign new_n260_ = pg0 & ph0;
  assign new_n261_ = ~pl & new_n260_;
  assign new_n262_ = ph0 & ~pl;
  assign new_n263_ = pk & new_n262_;
  assign new_n264_ = ~new_n259_ & ~new_n261_;
  assign pq1 = new_n263_ | ~new_n264_;
  assign new_n266_ = pa & ~pl;
  assign new_n267_ = pj & new_n266_;
  assign new_n268_ = pf0 & pa;
  assign new_n269_ = ~pl & new_n268_;
  assign new_n270_ = ~pj & new_n248_;
  assign new_n271_ = ~new_n267_ & ~new_n269_;
  assign pp1 = new_n270_ | ~new_n271_;
  assign new_n273_ = pi0 & ~pl;
  assign new_n274_ = ~pk & new_n273_;
  assign new_n275_ = pi0 & pj0;
  assign new_n276_ = ~pl & new_n275_;
  assign new_n277_ = pj0 & ~pl;
  assign new_n278_ = pk & new_n277_;
  assign new_n279_ = ~new_n274_ & ~new_n276_;
  assign ps1 = new_n278_ | ~new_n279_;
  assign new_n281_ = ~pk & new_n262_;
  assign new_n282_ = ph0 & pi0;
  assign new_n283_ = ~pl & new_n282_;
  assign new_n284_ = pk & new_n273_;
  assign new_n285_ = ~new_n281_ & ~new_n283_;
  assign pr1 = new_n284_ | ~new_n285_;
  assign new_n287_ = pk0 & ~pl;
  assign new_n288_ = ~pk & new_n287_;
  assign new_n289_ = pk0 & pl0;
  assign new_n290_ = ~pl & new_n289_;
  assign new_n291_ = pl0 & ~pl;
  assign new_n292_ = pk & new_n291_;
  assign new_n293_ = ~new_n288_ & ~new_n290_;
  assign pu1 = new_n292_ | ~new_n293_;
  assign new_n295_ = ~pk & new_n277_;
  assign new_n296_ = pj0 & pk0;
  assign new_n297_ = ~pl & new_n296_;
  assign new_n298_ = pk & new_n287_;
  assign new_n299_ = ~new_n295_ & ~new_n297_;
  assign pt1 = new_n298_ | ~new_n299_;
  assign new_n301_ = pm0 & ~pl;
  assign new_n302_ = ~pk & new_n301_;
  assign new_n303_ = pm0 & pn0;
  assign new_n304_ = ~pl & new_n303_;
  assign new_n305_ = pn0 & ~pl;
  assign new_n306_ = pk & new_n305_;
  assign new_n307_ = ~new_n302_ & ~new_n304_;
  assign pw1 = new_n306_ | ~new_n307_;
  assign new_n309_ = ~pk & new_n291_;
  assign new_n310_ = pl0 & pm0;
  assign new_n311_ = ~pl & new_n310_;
  assign new_n312_ = pk & new_n301_;
  assign new_n313_ = ~new_n309_ & ~new_n311_;
  assign pv1 = new_n312_ | ~new_n313_;
  assign new_n315_ = pf & ~pl;
  assign new_n316_ = pi & new_n315_;
  assign new_n317_ = pf & pm;
  assign new_n318_ = ~pl & new_n317_;
  assign new_n319_ = ~pl & pm;
  assign new_n320_ = ~pi & new_n319_;
  assign new_n321_ = ~new_n316_ & ~new_n318_;
  assign pw0 = new_n320_ | ~new_n321_;
  assign new_n323_ = pg & ~pl;
  assign new_n324_ = pi & new_n323_;
  assign new_n325_ = pg & pn;
  assign new_n326_ = ~pl & new_n325_;
  assign new_n327_ = ~pl & pn;
  assign new_n328_ = ~pi & new_n327_;
  assign new_n329_ = ~new_n324_ & ~new_n326_;
  assign px0 = new_n328_ | ~new_n329_;
  assign new_n331_ = pp0 & ~pl;
  assign new_n332_ = ~pp & new_n331_;
  assign new_n333_ = pk & new_n332_;
  assign new_n334_ = pp & po0;
  assign new_n335_ = ~pl & new_n334_;
  assign new_n336_ = po0 & pp0;
  assign new_n337_ = ~pl & new_n336_;
  assign new_n338_ = po0 & ~pl;
  assign new_n339_ = ~pk & new_n338_;
  assign new_n340_ = ~new_n333_ & ~new_n335_;
  assign new_n341_ = ~new_n337_ & ~new_n339_;
  assign py1 = ~new_n340_ | ~new_n341_;
  assign new_n343_ = po0 & pk;
  assign new_n344_ = ~pl & new_n343_;
  assign new_n345_ = pa & new_n344_;
  assign new_n346_ = ~pp & new_n338_;
  assign new_n347_ = pk & new_n346_;
  assign new_n348_ = pp & pk;
  assign new_n349_ = ~pl & new_n348_;
  assign new_n350_ = pa & new_n349_;
  assign new_n351_ = pp & new_n305_;
  assign new_n352_ = pa & new_n351_;
  assign new_n353_ = ~pk & new_n305_;
  assign new_n354_ = pn0 & new_n338_;
  assign new_n355_ = pa & new_n354_;
  assign new_n356_ = ~pp & po0;
  assign new_n357_ = pn0 & new_n356_;
  assign new_n358_ = ~pl & new_n357_;
  assign new_n359_ = ~new_n345_ & ~new_n347_;
  assign new_n360_ = ~new_n350_ & ~new_n352_;
  assign new_n361_ = new_n359_ & new_n360_;
  assign new_n362_ = ~new_n353_ & ~new_n355_;
  assign new_n363_ = ~new_n358_ & new_n362_;
  assign px1 = ~new_n361_ | ~new_n363_;
  assign new_n365_ = ph & ~pl;
  assign new_n366_ = pi & new_n365_;
  assign new_n367_ = ph & po;
  assign new_n368_ = ~pl & new_n367_;
  assign new_n369_ = ~pl & po;
  assign new_n370_ = ~pi & new_n369_;
  assign new_n371_ = ~new_n366_ & ~new_n368_;
  assign py0 = new_n370_ | ~new_n371_;
  assign new_n373_ = pc & ~pl;
  assign new_n374_ = pi & new_n373_;
  assign new_n375_ = pp & pc;
  assign new_n376_ = ~pl & new_n375_;
  assign new_n377_ = pp & ~pl;
  assign new_n378_ = ~pi & new_n377_;
  assign new_n379_ = ~new_n374_ & ~new_n376_;
  assign pz0 = new_n378_ | ~new_n379_;
  assign new_n381_ = ~pp & new_n129_;
  assign new_n382_ = pk & new_n381_;
  assign new_n383_ = pp & pp0;
  assign new_n384_ = ~pl & new_n383_;
  assign new_n385_ = pp0 & pq0;
  assign new_n386_ = ~pl & new_n385_;
  assign new_n387_ = ~pk & new_n331_;
  assign new_n388_ = ~new_n382_ & ~new_n384_;
  assign new_n389_ = ~new_n386_ & ~new_n387_;
  assign pz1 = ~new_n388_ | ~new_n389_;
endmodule

