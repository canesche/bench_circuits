// Benchmark "testing" written by ABC on Thu Oct  8 22:16:32 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A42  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A42;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ , \new_[350]_ ,
    \new_[351]_ , \new_[352]_ , \new_[353]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[405]_ ,
    \new_[406]_ , \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ ,
    \new_[411]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[436]_ , \new_[437]_ , \new_[438]_ , \new_[439]_ , \new_[440]_ ,
    \new_[441]_ , \new_[442]_ , \new_[443]_ , \new_[444]_ , \new_[445]_ ,
    \new_[446]_ , \new_[447]_ , \new_[448]_ , \new_[449]_ , \new_[450]_ ,
    \new_[451]_ , \new_[452]_ , \new_[453]_ , \new_[454]_ , \new_[455]_ ,
    \new_[456]_ , \new_[457]_ , \new_[458]_ , \new_[459]_ , \new_[460]_ ,
    \new_[461]_ , \new_[462]_ , \new_[463]_ , \new_[464]_ , \new_[465]_ ,
    \new_[466]_ , \new_[467]_ , \new_[468]_ , \new_[469]_ , \new_[470]_ ,
    \new_[471]_ , \new_[472]_ , \new_[473]_ , \new_[474]_ , \new_[475]_ ,
    \new_[476]_ , \new_[477]_ , \new_[478]_ , \new_[479]_ , \new_[480]_ ,
    \new_[481]_ , \new_[482]_ , \new_[483]_ , \new_[484]_ , \new_[485]_ ,
    \new_[486]_ , \new_[487]_ , \new_[488]_ , \new_[489]_ , \new_[490]_ ,
    \new_[491]_ , \new_[492]_ , \new_[493]_ , \new_[494]_ , \new_[495]_ ,
    \new_[496]_ , \new_[497]_ , \new_[498]_ , \new_[499]_ , \new_[500]_ ,
    \new_[501]_ , \new_[502]_ , \new_[503]_ , \new_[504]_ , \new_[505]_ ,
    \new_[506]_ , \new_[507]_ , \new_[508]_ , \new_[509]_ , \new_[510]_ ,
    \new_[511]_ , \new_[512]_ , \new_[513]_ , \new_[514]_ , \new_[515]_ ,
    \new_[516]_ , \new_[517]_ , \new_[518]_ , \new_[519]_ , \new_[520]_ ,
    \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[525]_ ,
    \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ , \new_[530]_ ,
    \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ , \new_[535]_ ,
    \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ , \new_[540]_ ,
    \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ , \new_[545]_ ,
    \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ , \new_[550]_ ,
    \new_[551]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[566]_ , \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ ,
    \new_[571]_ , \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ ,
    \new_[576]_ , \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ ,
    \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[584]_ , \new_[585]_ ,
    \new_[586]_ , \new_[587]_ , \new_[588]_ , \new_[589]_ , \new_[590]_ ,
    \new_[591]_ , \new_[592]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[598]_ , \new_[599]_ , \new_[600]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ ,
    \new_[611]_ , \new_[612]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[616]_ , \new_[617]_ , \new_[618]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[626]_ , \new_[627]_ , \new_[628]_ , \new_[629]_ , \new_[630]_ ,
    \new_[631]_ , \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ ,
    \new_[636]_ , \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ ,
    \new_[641]_ , \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ ,
    \new_[646]_ , \new_[647]_ , \new_[648]_ , \new_[649]_ , \new_[650]_ ,
    \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[655]_ ,
    \new_[656]_ , \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ ,
    \new_[661]_ , \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ ,
    \new_[666]_ , \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ ,
    \new_[671]_ , \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ ,
    \new_[676]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ ,
    \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ ,
    \new_[686]_ , \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ ,
    \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ ,
    \new_[696]_ , \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ ,
    \new_[701]_ , \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ ,
    \new_[706]_ , \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ ,
    \new_[711]_ , \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ ,
    \new_[716]_ , \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ ,
    \new_[726]_ , \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ ,
    \new_[731]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[736]_ , \new_[737]_ , \new_[738]_ , \new_[739]_ , \new_[740]_ ,
    \new_[741]_ , \new_[742]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ ,
    \new_[746]_ , \new_[747]_ , \new_[748]_ , \new_[749]_ , \new_[750]_ ,
    \new_[751]_ , \new_[752]_ , \new_[753]_ , \new_[754]_ , \new_[755]_ ,
    \new_[756]_ , \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ ,
    \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ ,
    \new_[766]_ , \new_[767]_ , \new_[768]_ , \new_[769]_ , \new_[770]_ ,
    \new_[771]_ , \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ ,
    \new_[776]_ , \new_[777]_ , \new_[778]_ , \new_[779]_ , \new_[780]_ ,
    \new_[781]_ , \new_[782]_ , \new_[783]_ , \new_[784]_ , \new_[785]_ ,
    \new_[786]_ , \new_[787]_ , \new_[788]_ , \new_[789]_ , \new_[790]_ ,
    \new_[791]_ , \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ ,
    \new_[796]_ , \new_[797]_ , \new_[798]_ , \new_[799]_ , \new_[800]_ ,
    \new_[801]_ , \new_[802]_ , \new_[803]_ , \new_[804]_ , \new_[805]_ ,
    \new_[806]_ , \new_[807]_ , \new_[808]_ , \new_[809]_ , \new_[810]_ ,
    \new_[811]_ , \new_[812]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ ,
    \new_[816]_ , \new_[817]_ , \new_[818]_ , \new_[819]_ , \new_[820]_ ,
    \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[824]_ , \new_[825]_ ,
    \new_[826]_ , \new_[827]_ , \new_[828]_ , \new_[829]_ , \new_[830]_ ,
    \new_[831]_ , \new_[832]_ , \new_[833]_ , \new_[834]_ , \new_[835]_ ,
    \new_[836]_ , \new_[837]_ , \new_[838]_ , \new_[839]_ , \new_[840]_ ,
    \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[845]_ ,
    \new_[846]_ , \new_[847]_ , \new_[848]_ , \new_[849]_ , \new_[850]_ ,
    \new_[851]_ , \new_[852]_ , \new_[853]_ , \new_[854]_ , \new_[855]_ ,
    \new_[856]_ , \new_[857]_ , \new_[858]_ , \new_[859]_ , \new_[860]_ ,
    \new_[861]_ , \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[865]_ ,
    \new_[866]_ , \new_[867]_ , \new_[868]_ , \new_[869]_ , \new_[870]_ ,
    \new_[871]_ , \new_[872]_ , \new_[873]_ , \new_[874]_ , \new_[875]_ ,
    \new_[876]_ , \new_[877]_ , \new_[878]_ , \new_[879]_ , \new_[880]_ ,
    \new_[881]_ , \new_[882]_ , \new_[883]_ , \new_[884]_ , \new_[885]_ ,
    \new_[886]_ , \new_[887]_ , \new_[888]_ , \new_[889]_ , \new_[890]_ ,
    \new_[891]_ , \new_[892]_ , \new_[893]_ , \new_[894]_ , \new_[895]_ ,
    \new_[896]_ , \new_[897]_ , \new_[898]_ , \new_[899]_ , \new_[900]_ ,
    \new_[901]_ , \new_[902]_ , \new_[903]_ , \new_[904]_ , \new_[905]_ ,
    \new_[906]_ , \new_[907]_ , \new_[908]_ , \new_[909]_ , \new_[910]_ ,
    \new_[911]_ , \new_[912]_ , \new_[913]_ , \new_[914]_ , \new_[915]_ ,
    \new_[916]_ , \new_[917]_ , \new_[918]_ , \new_[919]_ , \new_[920]_ ,
    \new_[921]_ , \new_[922]_ , \new_[923]_ , \new_[924]_ , \new_[925]_ ,
    \new_[926]_ , \new_[927]_ , \new_[928]_ , \new_[929]_ , \new_[930]_ ,
    \new_[931]_ , \new_[932]_ , \new_[933]_ , \new_[934]_ , \new_[935]_ ,
    \new_[936]_ , \new_[937]_ , \new_[938]_ , \new_[939]_ , \new_[940]_ ,
    \new_[941]_ , \new_[942]_ , \new_[943]_ , \new_[944]_ , \new_[945]_ ,
    \new_[946]_ , \new_[947]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ ,
    \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[955]_ ,
    \new_[956]_ , \new_[957]_ , \new_[958]_ , \new_[959]_ , \new_[960]_ ,
    \new_[961]_ , \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ ,
    \new_[966]_ , \new_[967]_ , \new_[968]_ , \new_[969]_ , \new_[970]_ ,
    \new_[971]_ , \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[975]_ ,
    \new_[976]_ , \new_[977]_ , \new_[978]_ , \new_[979]_ , \new_[980]_ ,
    \new_[981]_ , \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ ,
    \new_[986]_ , \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ ,
    \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ ,
    \new_[996]_ , \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ ,
    \new_[1001]_ , \new_[1002]_ , \new_[1003]_ , \new_[1004]_ ,
    \new_[1005]_ , \new_[1006]_ , \new_[1007]_ , \new_[1008]_ ,
    \new_[1009]_ , \new_[1010]_ , \new_[1011]_ , \new_[1012]_ ,
    \new_[1013]_ , \new_[1014]_ , \new_[1015]_ , \new_[1016]_ ,
    \new_[1017]_ , \new_[1018]_ , \new_[1019]_ , \new_[1020]_ ,
    \new_[1021]_ , \new_[1022]_ , \new_[1023]_ , \new_[1024]_ ,
    \new_[1025]_ , \new_[1026]_ , \new_[1027]_ , \new_[1028]_ ,
    \new_[1029]_ , \new_[1030]_ , \new_[1031]_ , \new_[1032]_ ,
    \new_[1033]_ , \new_[1034]_ , \new_[1035]_ , \new_[1036]_ ,
    \new_[1037]_ , \new_[1038]_ , \new_[1039]_ , \new_[1040]_ ,
    \new_[1041]_ , \new_[1042]_ , \new_[1043]_ , \new_[1044]_ ,
    \new_[1045]_ , \new_[1046]_ , \new_[1047]_ , \new_[1048]_ ,
    \new_[1049]_ , \new_[1050]_ , \new_[1051]_ , \new_[1052]_ ,
    \new_[1053]_ , \new_[1054]_ , \new_[1055]_ , \new_[1056]_ ,
    \new_[1057]_ , \new_[1058]_ , \new_[1059]_ , \new_[1060]_ ,
    \new_[1061]_ , \new_[1062]_ , \new_[1063]_ , \new_[1064]_ ,
    \new_[1065]_ , \new_[1066]_ , \new_[1067]_ , \new_[1068]_ ,
    \new_[1069]_ , \new_[1070]_ , \new_[1071]_ , \new_[1072]_ ,
    \new_[1073]_ , \new_[1074]_ , \new_[1075]_ , \new_[1076]_ ,
    \new_[1077]_ , \new_[1078]_ , \new_[1079]_ , \new_[1080]_ ,
    \new_[1081]_ , \new_[1082]_ , \new_[1083]_ , \new_[1084]_ ,
    \new_[1085]_ , \new_[1086]_ , \new_[1087]_ , \new_[1088]_ ,
    \new_[1089]_ , \new_[1090]_ , \new_[1091]_ , \new_[1092]_ ,
    \new_[1093]_ , \new_[1094]_ , \new_[1095]_ , \new_[1096]_ ,
    \new_[1097]_ , \new_[1098]_ , \new_[1099]_ , \new_[1100]_ ,
    \new_[1101]_ , \new_[1102]_ , \new_[1103]_ , \new_[1104]_ ,
    \new_[1105]_ , \new_[1106]_ , \new_[1107]_ , \new_[1108]_ ,
    \new_[1109]_ , \new_[1110]_ , \new_[1111]_ , \new_[1112]_ ,
    \new_[1113]_ , \new_[1114]_ , \new_[1115]_ , \new_[1116]_ ,
    \new_[1117]_ , \new_[1118]_ , \new_[1119]_ , \new_[1120]_ ,
    \new_[1121]_ , \new_[1122]_ , \new_[1123]_ , \new_[1124]_ ,
    \new_[1125]_ , \new_[1126]_ , \new_[1127]_ , \new_[1128]_ ,
    \new_[1129]_ , \new_[1130]_ , \new_[1131]_ , \new_[1132]_ ,
    \new_[1133]_ , \new_[1134]_ , \new_[1135]_ , \new_[1136]_ ,
    \new_[1137]_ , \new_[1138]_ , \new_[1139]_ , \new_[1140]_ ,
    \new_[1141]_ , \new_[1142]_ , \new_[1143]_ , \new_[1144]_ ,
    \new_[1145]_ , \new_[1146]_ , \new_[1147]_ , \new_[1148]_ ,
    \new_[1149]_ , \new_[1150]_ , \new_[1151]_ , \new_[1152]_ ,
    \new_[1153]_ , \new_[1154]_ , \new_[1155]_ , \new_[1156]_ ,
    \new_[1157]_ , \new_[1158]_ , \new_[1159]_ , \new_[1160]_ ,
    \new_[1161]_ , \new_[1162]_ , \new_[1163]_ , \new_[1164]_ ,
    \new_[1165]_ , \new_[1166]_ , \new_[1167]_ , \new_[1168]_ ,
    \new_[1169]_ , \new_[1170]_ , \new_[1171]_ , \new_[1172]_ ,
    \new_[1173]_ , \new_[1174]_ , \new_[1175]_ , \new_[1176]_ ,
    \new_[1177]_ , \new_[1178]_ , \new_[1179]_ , \new_[1180]_ ,
    \new_[1181]_ , \new_[1182]_ , \new_[1183]_ , \new_[1184]_ ,
    \new_[1185]_ , \new_[1186]_ , \new_[1187]_ , \new_[1188]_ ,
    \new_[1189]_ , \new_[1190]_ , \new_[1191]_ , \new_[1192]_ ,
    \new_[1193]_ , \new_[1194]_ , \new_[1195]_ , \new_[1196]_ ,
    \new_[1197]_ , \new_[1198]_ , \new_[1199]_ , \new_[1200]_ ,
    \new_[1201]_ , \new_[1202]_ , \new_[1203]_ , \new_[1204]_ ,
    \new_[1205]_ , \new_[1206]_ , \new_[1207]_ , \new_[1208]_ ,
    \new_[1209]_ , \new_[1210]_ , \new_[1211]_ , \new_[1212]_ ,
    \new_[1213]_ , \new_[1214]_ , \new_[1215]_ , \new_[1216]_ ,
    \new_[1217]_ , \new_[1218]_ , \new_[1219]_ , \new_[1220]_ ,
    \new_[1221]_ , \new_[1222]_ , \new_[1223]_ , \new_[1224]_ ,
    \new_[1225]_ , \new_[1226]_ , \new_[1227]_ , \new_[1228]_ ,
    \new_[1229]_ , \new_[1230]_ , \new_[1231]_ , \new_[1232]_ ,
    \new_[1233]_ , \new_[1234]_ , \new_[1235]_ , \new_[1236]_ ,
    \new_[1237]_ , \new_[1238]_ , \new_[1239]_ , \new_[1240]_ ,
    \new_[1241]_ , \new_[1242]_ , \new_[1243]_ , \new_[1244]_ ,
    \new_[1245]_ , \new_[1246]_ , \new_[1247]_ , \new_[1248]_ ,
    \new_[1249]_ , \new_[1250]_ , \new_[1251]_ , \new_[1252]_ ,
    \new_[1253]_ , \new_[1254]_ , \new_[1255]_ , \new_[1256]_ ,
    \new_[1257]_ , \new_[1258]_ , \new_[1259]_ , \new_[1260]_ ,
    \new_[1261]_ , \new_[1262]_ , \new_[1263]_ , \new_[1264]_ ,
    \new_[1265]_ , \new_[1266]_ , \new_[1267]_ , \new_[1268]_ ,
    \new_[1269]_ , \new_[1270]_ , \new_[1271]_ , \new_[1272]_ ,
    \new_[1273]_ , \new_[1274]_ , \new_[1275]_ , \new_[1276]_ ,
    \new_[1277]_ , \new_[1278]_ , \new_[1279]_ , \new_[1280]_ ,
    \new_[1281]_ , \new_[1282]_ , \new_[1283]_ , \new_[1284]_ ,
    \new_[1285]_ , \new_[1286]_ , \new_[1287]_ , \new_[1288]_ ,
    \new_[1289]_ , \new_[1290]_ , \new_[1291]_ , \new_[1292]_ ,
    \new_[1293]_ , \new_[1294]_ , \new_[1295]_ , \new_[1296]_ ,
    \new_[1297]_ , \new_[1298]_ , \new_[1299]_ , \new_[1300]_ ,
    \new_[1301]_ , \new_[1302]_ , \new_[1303]_ , \new_[1304]_ ,
    \new_[1305]_ , \new_[1306]_ , \new_[1307]_ , \new_[1308]_ ,
    \new_[1309]_ , \new_[1310]_ , \new_[1311]_ , \new_[1312]_ ,
    \new_[1313]_ , \new_[1314]_ , \new_[1315]_ , \new_[1316]_ ,
    \new_[1317]_ , \new_[1318]_ , \new_[1319]_ , \new_[1320]_ ,
    \new_[1321]_ , \new_[1322]_ , \new_[1323]_ , \new_[1324]_ ,
    \new_[1325]_ , \new_[1326]_ , \new_[1327]_ , \new_[1328]_ ,
    \new_[1329]_ , \new_[1330]_ , \new_[1331]_ , \new_[1332]_ ,
    \new_[1333]_ , \new_[1334]_ , \new_[1335]_ , \new_[1336]_ ,
    \new_[1337]_ , \new_[1338]_ , \new_[1339]_ , \new_[1340]_ ,
    \new_[1341]_ , \new_[1342]_ , \new_[1343]_ , \new_[1344]_ ,
    \new_[1345]_ , \new_[1346]_ , \new_[1347]_ , \new_[1348]_ ,
    \new_[1349]_ , \new_[1350]_ , \new_[1351]_ , \new_[1352]_ ,
    \new_[1353]_ , \new_[1354]_ , \new_[1355]_ , \new_[1356]_ ,
    \new_[1357]_ , \new_[1358]_ , \new_[1359]_ , \new_[1360]_ ,
    \new_[1361]_ , \new_[1362]_ , \new_[1363]_ , \new_[1364]_ ,
    \new_[1365]_ , \new_[1366]_ , \new_[1367]_ , \new_[1368]_ ,
    \new_[1369]_ , \new_[1370]_ , \new_[1371]_ , \new_[1372]_ ,
    \new_[1373]_ , \new_[1374]_ , \new_[1375]_ , \new_[1376]_ ,
    \new_[1377]_ , \new_[1378]_ , \new_[1379]_ , \new_[1380]_ ,
    \new_[1381]_ , \new_[1382]_ , \new_[1383]_ , \new_[1384]_ ,
    \new_[1385]_ , \new_[1386]_ , \new_[1387]_ , \new_[1388]_ ,
    \new_[1389]_ , \new_[1390]_ , \new_[1391]_ , \new_[1392]_ ,
    \new_[1393]_ , \new_[1394]_ , \new_[1395]_ , \new_[1396]_ ,
    \new_[1397]_ , \new_[1398]_ , \new_[1399]_ , \new_[1400]_ ,
    \new_[1401]_ , \new_[1402]_ , \new_[1403]_ , \new_[1404]_ ,
    \new_[1405]_ , \new_[1406]_ , \new_[1407]_ , \new_[1408]_ ,
    \new_[1409]_ , \new_[1410]_ , \new_[1411]_ , \new_[1412]_ ,
    \new_[1413]_ , \new_[1414]_ , \new_[1415]_ , \new_[1416]_ ,
    \new_[1417]_ , \new_[1418]_ , \new_[1419]_ , \new_[1420]_ ,
    \new_[1421]_ , \new_[1422]_ , \new_[1423]_ , \new_[1424]_ ,
    \new_[1425]_ , \new_[1426]_ , \new_[1427]_ , \new_[1428]_ ,
    \new_[1429]_ , \new_[1430]_ , \new_[1431]_ , \new_[1432]_ ,
    \new_[1433]_ , \new_[1434]_ , \new_[1435]_ , \new_[1436]_ ,
    \new_[1437]_ , \new_[1438]_ , \new_[1439]_ , \new_[1440]_ ,
    \new_[1441]_ , \new_[1442]_ , \new_[1443]_ , \new_[1444]_ ,
    \new_[1445]_ , \new_[1446]_ , \new_[1447]_ , \new_[1448]_ ,
    \new_[1449]_ , \new_[1450]_ , \new_[1451]_ , \new_[1452]_ ,
    \new_[1453]_ , \new_[1454]_ , \new_[1455]_ , \new_[1456]_ ,
    \new_[1457]_ , \new_[1458]_ , \new_[1459]_ , \new_[1460]_ ,
    \new_[1461]_ , \new_[1462]_ , \new_[1463]_ , \new_[1464]_ ,
    \new_[1465]_ , \new_[1466]_ , \new_[1467]_ , \new_[1468]_ ,
    \new_[1469]_ , \new_[1470]_ , \new_[1471]_ , \new_[1472]_ ,
    \new_[1473]_ , \new_[1474]_ , \new_[1475]_ , \new_[1476]_ ,
    \new_[1477]_ , \new_[1478]_ , \new_[1479]_ , \new_[1480]_ ,
    \new_[1481]_ , \new_[1482]_ , \new_[1483]_ , \new_[1484]_ ,
    \new_[1485]_ , \new_[1486]_ , \new_[1487]_ , \new_[1488]_ ,
    \new_[1489]_ , \new_[1490]_ , \new_[1491]_ , \new_[1492]_ ,
    \new_[1493]_ , \new_[1494]_ , \new_[1495]_ , \new_[1496]_ ,
    \new_[1497]_ , \new_[1498]_ , \new_[1499]_ , \new_[1500]_ ,
    \new_[1501]_ , \new_[1502]_ , \new_[1503]_ , \new_[1504]_ ,
    \new_[1505]_ , \new_[1506]_ , \new_[1507]_ , \new_[1508]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1512]_ ,
    \new_[1513]_ , \new_[1514]_ , \new_[1515]_ , \new_[1516]_ ,
    \new_[1517]_ , \new_[1518]_ , \new_[1519]_ , \new_[1520]_ ,
    \new_[1521]_ , \new_[1522]_ , \new_[1523]_ , \new_[1524]_ ,
    \new_[1525]_ , \new_[1526]_ , \new_[1527]_ , \new_[1528]_ ,
    \new_[1529]_ , \new_[1530]_ , \new_[1531]_ , \new_[1532]_ ,
    \new_[1533]_ , \new_[1534]_ , \new_[1535]_ , \new_[1536]_ ,
    \new_[1537]_ , \new_[1538]_ , \new_[1539]_ , \new_[1540]_ ,
    \new_[1541]_ , \new_[1542]_ , \new_[1543]_ , \new_[1544]_ ,
    \new_[1545]_ , \new_[1546]_ , \new_[1547]_ , \new_[1548]_ ,
    \new_[1549]_ , \new_[1550]_ , \new_[1551]_ , \new_[1552]_ ,
    \new_[1553]_ , \new_[1554]_ , \new_[1555]_ , \new_[1556]_ ,
    \new_[1557]_ , \new_[1558]_ , \new_[1559]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1562]_ , \new_[1563]_ , \new_[1564]_ ,
    \new_[1565]_ , \new_[1566]_ , \new_[1567]_ , \new_[1568]_ ,
    \new_[1569]_ , \new_[1570]_ , \new_[1571]_ , \new_[1572]_ ,
    \new_[1573]_ , \new_[1574]_ , \new_[1575]_ , \new_[1576]_ ,
    \new_[1577]_ , \new_[1578]_ , \new_[1579]_ , \new_[1580]_ ,
    \new_[1581]_ , \new_[1582]_ , \new_[1583]_ , \new_[1584]_ ,
    \new_[1585]_ , \new_[1586]_ , \new_[1587]_ , \new_[1588]_ ,
    \new_[1589]_ , \new_[1590]_ , \new_[1591]_ , \new_[1592]_ ,
    \new_[1593]_ , \new_[1594]_ , \new_[1595]_ , \new_[1596]_ ,
    \new_[1597]_ , \new_[1598]_ , \new_[1599]_ , \new_[1600]_ ,
    \new_[1601]_ , \new_[1602]_ , \new_[1603]_ , \new_[1604]_ ,
    \new_[1605]_ , \new_[1606]_ , \new_[1607]_ , \new_[1608]_ ,
    \new_[1609]_ , \new_[1610]_ , \new_[1611]_ , \new_[1612]_ ,
    \new_[1613]_ , \new_[1614]_ , \new_[1615]_ , \new_[1616]_ ,
    \new_[1617]_ , \new_[1618]_ , \new_[1619]_ , \new_[1620]_ ,
    \new_[1621]_ , \new_[1622]_ , \new_[1623]_ , \new_[1624]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1627]_ , \new_[1628]_ ,
    \new_[1629]_ , \new_[1630]_ , \new_[1631]_ , \new_[1632]_ ,
    \new_[1633]_ , \new_[1634]_ , \new_[1635]_ , \new_[1636]_ ,
    \new_[1637]_ , \new_[1638]_ , \new_[1639]_ , \new_[1640]_ ,
    \new_[1641]_ , \new_[1642]_ , \new_[1643]_ , \new_[1644]_ ,
    \new_[1645]_ , \new_[1646]_ , \new_[1647]_ , \new_[1648]_ ,
    \new_[1649]_ , \new_[1650]_ , \new_[1651]_ , \new_[1652]_ ,
    \new_[1653]_ , \new_[1654]_ , \new_[1655]_ , \new_[1656]_ ,
    \new_[1657]_ , \new_[1658]_ , \new_[1659]_ , \new_[1660]_ ,
    \new_[1661]_ , \new_[1662]_ , \new_[1663]_ , \new_[1664]_ ,
    \new_[1665]_ , \new_[1666]_ , \new_[1667]_ , \new_[1668]_ ,
    \new_[1669]_ , \new_[1670]_ , \new_[1671]_ , \new_[1672]_ ,
    \new_[1673]_ , \new_[1674]_ , \new_[1675]_ , \new_[1676]_ ,
    \new_[1677]_ , \new_[1678]_ , \new_[1679]_ , \new_[1680]_ ,
    \new_[1681]_ , \new_[1682]_ , \new_[1683]_ , \new_[1684]_ ,
    \new_[1685]_ , \new_[1686]_ , \new_[1687]_ , \new_[1688]_ ,
    \new_[1689]_ , \new_[1690]_ , \new_[1691]_ , \new_[1692]_ ,
    \new_[1693]_ , \new_[1694]_ , \new_[1695]_ , \new_[1696]_ ,
    \new_[1697]_ , \new_[1698]_ , \new_[1699]_ , \new_[1700]_ ,
    \new_[1701]_ , \new_[1702]_ , \new_[1703]_ , \new_[1704]_ ,
    \new_[1705]_ , \new_[1706]_ , \new_[1707]_ , \new_[1708]_ ,
    \new_[1709]_ , \new_[1710]_ , \new_[1711]_ , \new_[1712]_ ,
    \new_[1713]_ , \new_[1714]_ , \new_[1715]_ , \new_[1716]_ ,
    \new_[1717]_ , \new_[1718]_ , \new_[1719]_ , \new_[1720]_ ,
    \new_[1721]_ , \new_[1722]_ , \new_[1723]_ , \new_[1724]_ ,
    \new_[1725]_ , \new_[1726]_ , \new_[1727]_ , \new_[1728]_ ,
    \new_[1729]_ , \new_[1730]_ , \new_[1731]_ , \new_[1732]_ ,
    \new_[1733]_ , \new_[1734]_ , \new_[1735]_ , \new_[1736]_ ,
    \new_[1737]_ , \new_[1738]_ , \new_[1739]_ , \new_[1740]_ ,
    \new_[1741]_ , \new_[1742]_ , \new_[1743]_ , \new_[1744]_ ,
    \new_[1745]_ , \new_[1746]_ , \new_[1747]_ , \new_[1748]_ ,
    \new_[1749]_ , \new_[1750]_ , \new_[1751]_ , \new_[1752]_ ,
    \new_[1756]_ , \new_[1757]_ , \new_[1761]_ , \new_[1762]_ ,
    \new_[1763]_ , \new_[1767]_ , \new_[1768]_ , \new_[1771]_ ,
    \new_[1774]_ , \new_[1775]_ , \new_[1776]_ , \new_[1777]_ ,
    \new_[1781]_ , \new_[1782]_ , \new_[1785]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1794]_ , \new_[1795]_ ,
    \new_[1798]_ , \new_[1801]_ , \new_[1802]_ , \new_[1803]_ ,
    \new_[1804]_ , \new_[1805]_ , \new_[1809]_ , \new_[1810]_ ,
    \new_[1814]_ , \new_[1815]_ , \new_[1816]_ , \new_[1820]_ ,
    \new_[1821]_ , \new_[1824]_ , \new_[1827]_ , \new_[1828]_ ,
    \new_[1829]_ , \new_[1830]_ , \new_[1834]_ , \new_[1835]_ ,
    \new_[1838]_ , \new_[1841]_ , \new_[1842]_ , \new_[1843]_ ,
    \new_[1847]_ , \new_[1848]_ , \new_[1851]_ , \new_[1854]_ ,
    \new_[1855]_ , \new_[1856]_ , \new_[1857]_ , \new_[1858]_ ,
    \new_[1859]_ , \new_[1863]_ , \new_[1864]_ , \new_[1868]_ ,
    \new_[1869]_ , \new_[1870]_ , \new_[1874]_ , \new_[1875]_ ,
    \new_[1878]_ , \new_[1881]_ , \new_[1882]_ , \new_[1883]_ ,
    \new_[1884]_ , \new_[1888]_ , \new_[1889]_ , \new_[1892]_ ,
    \new_[1895]_ , \new_[1896]_ , \new_[1897]_ , \new_[1901]_ ,
    \new_[1902]_ , \new_[1905]_ , \new_[1908]_ , \new_[1909]_ ,
    \new_[1910]_ , \new_[1911]_ , \new_[1912]_ , \new_[1916]_ ,
    \new_[1917]_ , \new_[1920]_ , \new_[1923]_ , \new_[1924]_ ,
    \new_[1925]_ , \new_[1929]_ , \new_[1930]_ , \new_[1933]_ ,
    \new_[1936]_ , \new_[1937]_ , \new_[1938]_ , \new_[1939]_ ,
    \new_[1943]_ , \new_[1944]_ , \new_[1947]_ , \new_[1950]_ ,
    \new_[1951]_ , \new_[1952]_ , \new_[1956]_ , \new_[1957]_ ,
    \new_[1960]_ , \new_[1963]_ , \new_[1964]_ , \new_[1965]_ ,
    \new_[1966]_ , \new_[1967]_ , \new_[1968]_ , \new_[1969]_ ,
    \new_[1973]_ , \new_[1974]_ , \new_[1978]_ , \new_[1979]_ ,
    \new_[1980]_ , \new_[1984]_ , \new_[1985]_ , \new_[1988]_ ,
    \new_[1991]_ , \new_[1992]_ , \new_[1993]_ , \new_[1994]_ ,
    \new_[1998]_ , \new_[1999]_ , \new_[2002]_ , \new_[2005]_ ,
    \new_[2006]_ , \new_[2007]_ , \new_[2011]_ , \new_[2012]_ ,
    \new_[2015]_ , \new_[2018]_ , \new_[2019]_ , \new_[2020]_ ,
    \new_[2021]_ , \new_[2022]_ , \new_[2026]_ , \new_[2027]_ ,
    \new_[2030]_ , \new_[2033]_ , \new_[2034]_ , \new_[2035]_ ,
    \new_[2039]_ , \new_[2040]_ , \new_[2043]_ , \new_[2046]_ ,
    \new_[2047]_ , \new_[2048]_ , \new_[2049]_ , \new_[2053]_ ,
    \new_[2054]_ , \new_[2057]_ , \new_[2060]_ , \new_[2061]_ ,
    \new_[2062]_ , \new_[2066]_ , \new_[2067]_ , \new_[2070]_ ,
    \new_[2073]_ , \new_[2074]_ , \new_[2075]_ , \new_[2076]_ ,
    \new_[2077]_ , \new_[2078]_ , \new_[2082]_ , \new_[2083]_ ,
    \new_[2087]_ , \new_[2088]_ , \new_[2089]_ , \new_[2093]_ ,
    \new_[2094]_ , \new_[2097]_ , \new_[2100]_ , \new_[2101]_ ,
    \new_[2102]_ , \new_[2103]_ , \new_[2107]_ , \new_[2108]_ ,
    \new_[2111]_ , \new_[2114]_ , \new_[2115]_ , \new_[2116]_ ,
    \new_[2120]_ , \new_[2121]_ , \new_[2124]_ , \new_[2127]_ ,
    \new_[2128]_ , \new_[2129]_ , \new_[2130]_ , \new_[2131]_ ,
    \new_[2135]_ , \new_[2136]_ , \new_[2139]_ , \new_[2142]_ ,
    \new_[2143]_ , \new_[2144]_ , \new_[2148]_ , \new_[2149]_ ,
    \new_[2152]_ , \new_[2155]_ , \new_[2156]_ , \new_[2157]_ ,
    \new_[2158]_ , \new_[2162]_ , \new_[2163]_ , \new_[2166]_ ,
    \new_[2169]_ , \new_[2170]_ , \new_[2171]_ , \new_[2175]_ ,
    \new_[2176]_ , \new_[2179]_ , \new_[2182]_ , \new_[2183]_ ,
    \new_[2184]_ , \new_[2185]_ , \new_[2186]_ , \new_[2187]_ ,
    \new_[2188]_ , \new_[2189]_ , \new_[2193]_ , \new_[2194]_ ,
    \new_[2198]_ , \new_[2199]_ , \new_[2200]_ , \new_[2204]_ ,
    \new_[2205]_ , \new_[2208]_ , \new_[2211]_ , \new_[2212]_ ,
    \new_[2213]_ , \new_[2214]_ , \new_[2218]_ , \new_[2219]_ ,
    \new_[2222]_ , \new_[2225]_ , \new_[2226]_ , \new_[2227]_ ,
    \new_[2231]_ , \new_[2232]_ , \new_[2235]_ , \new_[2238]_ ,
    \new_[2239]_ , \new_[2240]_ , \new_[2241]_ , \new_[2242]_ ,
    \new_[2246]_ , \new_[2247]_ , \new_[2251]_ , \new_[2252]_ ,
    \new_[2253]_ , \new_[2257]_ , \new_[2258]_ , \new_[2261]_ ,
    \new_[2264]_ , \new_[2265]_ , \new_[2266]_ , \new_[2267]_ ,
    \new_[2271]_ , \new_[2272]_ , \new_[2275]_ , \new_[2278]_ ,
    \new_[2279]_ , \new_[2280]_ , \new_[2284]_ , \new_[2285]_ ,
    \new_[2288]_ , \new_[2291]_ , \new_[2292]_ , \new_[2293]_ ,
    \new_[2294]_ , \new_[2295]_ , \new_[2296]_ , \new_[2300]_ ,
    \new_[2301]_ , \new_[2305]_ , \new_[2306]_ , \new_[2307]_ ,
    \new_[2311]_ , \new_[2312]_ , \new_[2315]_ , \new_[2318]_ ,
    \new_[2319]_ , \new_[2320]_ , \new_[2321]_ , \new_[2325]_ ,
    \new_[2326]_ , \new_[2329]_ , \new_[2332]_ , \new_[2333]_ ,
    \new_[2334]_ , \new_[2338]_ , \new_[2339]_ , \new_[2342]_ ,
    \new_[2345]_ , \new_[2346]_ , \new_[2347]_ , \new_[2348]_ ,
    \new_[2349]_ , \new_[2353]_ , \new_[2354]_ , \new_[2357]_ ,
    \new_[2360]_ , \new_[2361]_ , \new_[2362]_ , \new_[2366]_ ,
    \new_[2367]_ , \new_[2370]_ , \new_[2373]_ , \new_[2374]_ ,
    \new_[2375]_ , \new_[2376]_ , \new_[2380]_ , \new_[2381]_ ,
    \new_[2384]_ , \new_[2387]_ , \new_[2388]_ , \new_[2389]_ ,
    \new_[2393]_ , \new_[2394]_ , \new_[2397]_ , \new_[2400]_ ,
    \new_[2401]_ , \new_[2402]_ , \new_[2403]_ , \new_[2404]_ ,
    \new_[2405]_ , \new_[2406]_ , \new_[2410]_ , \new_[2411]_ ,
    \new_[2415]_ , \new_[2416]_ , \new_[2417]_ , \new_[2421]_ ,
    \new_[2422]_ , \new_[2425]_ , \new_[2428]_ , \new_[2429]_ ,
    \new_[2430]_ , \new_[2431]_ , \new_[2435]_ , \new_[2436]_ ,
    \new_[2439]_ , \new_[2442]_ , \new_[2443]_ , \new_[2444]_ ,
    \new_[2448]_ , \new_[2449]_ , \new_[2452]_ , \new_[2455]_ ,
    \new_[2456]_ , \new_[2457]_ , \new_[2458]_ , \new_[2459]_ ,
    \new_[2463]_ , \new_[2464]_ , \new_[2467]_ , \new_[2470]_ ,
    \new_[2471]_ , \new_[2472]_ , \new_[2476]_ , \new_[2477]_ ,
    \new_[2480]_ , \new_[2483]_ , \new_[2484]_ , \new_[2485]_ ,
    \new_[2486]_ , \new_[2490]_ , \new_[2491]_ , \new_[2494]_ ,
    \new_[2497]_ , \new_[2498]_ , \new_[2499]_ , \new_[2503]_ ,
    \new_[2504]_ , \new_[2507]_ , \new_[2510]_ , \new_[2511]_ ,
    \new_[2512]_ , \new_[2513]_ , \new_[2514]_ , \new_[2515]_ ,
    \new_[2519]_ , \new_[2520]_ , \new_[2524]_ , \new_[2525]_ ,
    \new_[2526]_ , \new_[2530]_ , \new_[2531]_ , \new_[2534]_ ,
    \new_[2537]_ , \new_[2538]_ , \new_[2539]_ , \new_[2540]_ ,
    \new_[2544]_ , \new_[2545]_ , \new_[2548]_ , \new_[2551]_ ,
    \new_[2552]_ , \new_[2553]_ , \new_[2557]_ , \new_[2558]_ ,
    \new_[2561]_ , \new_[2564]_ , \new_[2565]_ , \new_[2566]_ ,
    \new_[2567]_ , \new_[2568]_ , \new_[2572]_ , \new_[2573]_ ,
    \new_[2576]_ , \new_[2579]_ , \new_[2580]_ , \new_[2581]_ ,
    \new_[2585]_ , \new_[2586]_ , \new_[2589]_ , \new_[2592]_ ,
    \new_[2593]_ , \new_[2594]_ , \new_[2595]_ , \new_[2599]_ ,
    \new_[2600]_ , \new_[2603]_ , \new_[2606]_ , \new_[2607]_ ,
    \new_[2608]_ , \new_[2612]_ , \new_[2613]_ , \new_[2616]_ ,
    \new_[2619]_ , \new_[2620]_ , \new_[2621]_ , \new_[2622]_ ,
    \new_[2623]_ , \new_[2624]_ , \new_[2625]_ , \new_[2626]_ ,
    \new_[2627]_ , \new_[2631]_ , \new_[2632]_ , \new_[2636]_ ,
    \new_[2637]_ , \new_[2638]_ , \new_[2642]_ , \new_[2643]_ ,
    \new_[2646]_ , \new_[2649]_ , \new_[2650]_ , \new_[2651]_ ,
    \new_[2652]_ , \new_[2656]_ , \new_[2657]_ , \new_[2660]_ ,
    \new_[2663]_ , \new_[2664]_ , \new_[2665]_ , \new_[2669]_ ,
    \new_[2670]_ , \new_[2673]_ , \new_[2676]_ , \new_[2677]_ ,
    \new_[2678]_ , \new_[2679]_ , \new_[2680]_ , \new_[2684]_ ,
    \new_[2685]_ , \new_[2689]_ , \new_[2690]_ , \new_[2691]_ ,
    \new_[2695]_ , \new_[2696]_ , \new_[2699]_ , \new_[2702]_ ,
    \new_[2703]_ , \new_[2704]_ , \new_[2705]_ , \new_[2709]_ ,
    \new_[2710]_ , \new_[2713]_ , \new_[2716]_ , \new_[2717]_ ,
    \new_[2718]_ , \new_[2722]_ , \new_[2723]_ , \new_[2726]_ ,
    \new_[2729]_ , \new_[2730]_ , \new_[2731]_ , \new_[2732]_ ,
    \new_[2733]_ , \new_[2734]_ , \new_[2738]_ , \new_[2739]_ ,
    \new_[2743]_ , \new_[2744]_ , \new_[2745]_ , \new_[2749]_ ,
    \new_[2750]_ , \new_[2753]_ , \new_[2756]_ , \new_[2757]_ ,
    \new_[2758]_ , \new_[2759]_ , \new_[2763]_ , \new_[2764]_ ,
    \new_[2767]_ , \new_[2770]_ , \new_[2771]_ , \new_[2772]_ ,
    \new_[2776]_ , \new_[2777]_ , \new_[2780]_ , \new_[2783]_ ,
    \new_[2784]_ , \new_[2785]_ , \new_[2786]_ , \new_[2787]_ ,
    \new_[2791]_ , \new_[2792]_ , \new_[2795]_ , \new_[2798]_ ,
    \new_[2799]_ , \new_[2800]_ , \new_[2804]_ , \new_[2805]_ ,
    \new_[2808]_ , \new_[2811]_ , \new_[2812]_ , \new_[2813]_ ,
    \new_[2814]_ , \new_[2818]_ , \new_[2819]_ , \new_[2822]_ ,
    \new_[2825]_ , \new_[2826]_ , \new_[2827]_ , \new_[2831]_ ,
    \new_[2832]_ , \new_[2835]_ , \new_[2838]_ , \new_[2839]_ ,
    \new_[2840]_ , \new_[2841]_ , \new_[2842]_ , \new_[2843]_ ,
    \new_[2844]_ , \new_[2848]_ , \new_[2849]_ , \new_[2853]_ ,
    \new_[2854]_ , \new_[2855]_ , \new_[2859]_ , \new_[2860]_ ,
    \new_[2863]_ , \new_[2866]_ , \new_[2867]_ , \new_[2868]_ ,
    \new_[2869]_ , \new_[2873]_ , \new_[2874]_ , \new_[2877]_ ,
    \new_[2880]_ , \new_[2881]_ , \new_[2882]_ , \new_[2886]_ ,
    \new_[2887]_ , \new_[2890]_ , \new_[2893]_ , \new_[2894]_ ,
    \new_[2895]_ , \new_[2896]_ , \new_[2897]_ , \new_[2901]_ ,
    \new_[2902]_ , \new_[2905]_ , \new_[2908]_ , \new_[2909]_ ,
    \new_[2910]_ , \new_[2914]_ , \new_[2915]_ , \new_[2918]_ ,
    \new_[2921]_ , \new_[2922]_ , \new_[2923]_ , \new_[2924]_ ,
    \new_[2928]_ , \new_[2929]_ , \new_[2932]_ , \new_[2935]_ ,
    \new_[2936]_ , \new_[2937]_ , \new_[2941]_ , \new_[2942]_ ,
    \new_[2945]_ , \new_[2948]_ , \new_[2949]_ , \new_[2950]_ ,
    \new_[2951]_ , \new_[2952]_ , \new_[2953]_ , \new_[2957]_ ,
    \new_[2958]_ , \new_[2962]_ , \new_[2963]_ , \new_[2964]_ ,
    \new_[2968]_ , \new_[2969]_ , \new_[2972]_ , \new_[2975]_ ,
    \new_[2976]_ , \new_[2977]_ , \new_[2978]_ , \new_[2982]_ ,
    \new_[2983]_ , \new_[2986]_ , \new_[2989]_ , \new_[2990]_ ,
    \new_[2991]_ , \new_[2995]_ , \new_[2996]_ , \new_[2999]_ ,
    \new_[3002]_ , \new_[3003]_ , \new_[3004]_ , \new_[3005]_ ,
    \new_[3006]_ , \new_[3010]_ , \new_[3011]_ , \new_[3014]_ ,
    \new_[3017]_ , \new_[3018]_ , \new_[3019]_ , \new_[3023]_ ,
    \new_[3024]_ , \new_[3027]_ , \new_[3030]_ , \new_[3031]_ ,
    \new_[3032]_ , \new_[3033]_ , \new_[3037]_ , \new_[3038]_ ,
    \new_[3041]_ , \new_[3044]_ , \new_[3045]_ , \new_[3046]_ ,
    \new_[3050]_ , \new_[3051]_ , \new_[3054]_ , \new_[3057]_ ,
    \new_[3058]_ , \new_[3059]_ , \new_[3060]_ , \new_[3061]_ ,
    \new_[3062]_ , \new_[3063]_ , \new_[3064]_ , \new_[3068]_ ,
    \new_[3069]_ , \new_[3073]_ , \new_[3074]_ , \new_[3075]_ ,
    \new_[3079]_ , \new_[3080]_ , \new_[3083]_ , \new_[3086]_ ,
    \new_[3087]_ , \new_[3088]_ , \new_[3089]_ , \new_[3093]_ ,
    \new_[3094]_ , \new_[3097]_ , \new_[3100]_ , \new_[3101]_ ,
    \new_[3102]_ , \new_[3106]_ , \new_[3107]_ , \new_[3110]_ ,
    \new_[3113]_ , \new_[3114]_ , \new_[3115]_ , \new_[3116]_ ,
    \new_[3117]_ , \new_[3121]_ , \new_[3122]_ , \new_[3126]_ ,
    \new_[3127]_ , \new_[3128]_ , \new_[3132]_ , \new_[3133]_ ,
    \new_[3136]_ , \new_[3139]_ , \new_[3140]_ , \new_[3141]_ ,
    \new_[3142]_ , \new_[3146]_ , \new_[3147]_ , \new_[3150]_ ,
    \new_[3153]_ , \new_[3154]_ , \new_[3155]_ , \new_[3159]_ ,
    \new_[3160]_ , \new_[3163]_ , \new_[3166]_ , \new_[3167]_ ,
    \new_[3168]_ , \new_[3169]_ , \new_[3170]_ , \new_[3171]_ ,
    \new_[3175]_ , \new_[3176]_ , \new_[3180]_ , \new_[3181]_ ,
    \new_[3182]_ , \new_[3186]_ , \new_[3187]_ , \new_[3190]_ ,
    \new_[3193]_ , \new_[3194]_ , \new_[3195]_ , \new_[3196]_ ,
    \new_[3200]_ , \new_[3201]_ , \new_[3204]_ , \new_[3207]_ ,
    \new_[3208]_ , \new_[3209]_ , \new_[3213]_ , \new_[3214]_ ,
    \new_[3217]_ , \new_[3220]_ , \new_[3221]_ , \new_[3222]_ ,
    \new_[3223]_ , \new_[3224]_ , \new_[3228]_ , \new_[3229]_ ,
    \new_[3232]_ , \new_[3235]_ , \new_[3236]_ , \new_[3237]_ ,
    \new_[3241]_ , \new_[3242]_ , \new_[3245]_ , \new_[3248]_ ,
    \new_[3249]_ , \new_[3250]_ , \new_[3251]_ , \new_[3255]_ ,
    \new_[3256]_ , \new_[3259]_ , \new_[3262]_ , \new_[3263]_ ,
    \new_[3264]_ , \new_[3268]_ , \new_[3269]_ , \new_[3272]_ ,
    \new_[3275]_ , \new_[3276]_ , \new_[3277]_ , \new_[3278]_ ,
    \new_[3279]_ , \new_[3280]_ , \new_[3281]_ , \new_[3285]_ ,
    \new_[3286]_ , \new_[3290]_ , \new_[3291]_ , \new_[3292]_ ,
    \new_[3296]_ , \new_[3297]_ , \new_[3300]_ , \new_[3303]_ ,
    \new_[3304]_ , \new_[3305]_ , \new_[3306]_ , \new_[3310]_ ,
    \new_[3311]_ , \new_[3314]_ , \new_[3317]_ , \new_[3318]_ ,
    \new_[3319]_ , \new_[3323]_ , \new_[3324]_ , \new_[3327]_ ,
    \new_[3330]_ , \new_[3331]_ , \new_[3332]_ , \new_[3333]_ ,
    \new_[3334]_ , \new_[3338]_ , \new_[3339]_ , \new_[3342]_ ,
    \new_[3345]_ , \new_[3346]_ , \new_[3347]_ , \new_[3351]_ ,
    \new_[3352]_ , \new_[3355]_ , \new_[3358]_ , \new_[3359]_ ,
    \new_[3360]_ , \new_[3361]_ , \new_[3365]_ , \new_[3366]_ ,
    \new_[3369]_ , \new_[3372]_ , \new_[3373]_ , \new_[3374]_ ,
    \new_[3378]_ , \new_[3379]_ , \new_[3382]_ , \new_[3385]_ ,
    \new_[3386]_ , \new_[3387]_ , \new_[3388]_ , \new_[3389]_ ,
    \new_[3390]_ , \new_[3394]_ , \new_[3395]_ , \new_[3399]_ ,
    \new_[3400]_ , \new_[3401]_ , \new_[3405]_ , \new_[3406]_ ,
    \new_[3409]_ , \new_[3412]_ , \new_[3413]_ , \new_[3414]_ ,
    \new_[3415]_ , \new_[3419]_ , \new_[3420]_ , \new_[3423]_ ,
    \new_[3426]_ , \new_[3427]_ , \new_[3428]_ , \new_[3432]_ ,
    \new_[3433]_ , \new_[3436]_ , \new_[3439]_ , \new_[3440]_ ,
    \new_[3441]_ , \new_[3442]_ , \new_[3443]_ , \new_[3447]_ ,
    \new_[3448]_ , \new_[3451]_ , \new_[3454]_ , \new_[3455]_ ,
    \new_[3456]_ , \new_[3460]_ , \new_[3461]_ , \new_[3464]_ ,
    \new_[3467]_ , \new_[3468]_ , \new_[3469]_ , \new_[3470]_ ,
    \new_[3474]_ , \new_[3475]_ , \new_[3478]_ , \new_[3481]_ ,
    \new_[3482]_ , \new_[3483]_ , \new_[3487]_ , \new_[3488]_ ,
    \new_[3491]_ , \new_[3494]_ , \new_[3495]_ , \new_[3496]_ ,
    \new_[3497]_ , \new_[3498]_ , \new_[3499]_ , \new_[3500]_ ,
    \new_[3501]_ , \new_[3502]_ , \new_[3503]_ , \new_[3507]_ ,
    \new_[3508]_ , \new_[3512]_ , \new_[3513]_ , \new_[3514]_ ,
    \new_[3518]_ , \new_[3519]_ , \new_[3522]_ , \new_[3525]_ ,
    \new_[3526]_ , \new_[3527]_ , \new_[3528]_ , \new_[3532]_ ,
    \new_[3533]_ , \new_[3536]_ , \new_[3539]_ , \new_[3540]_ ,
    \new_[3541]_ , \new_[3545]_ , \new_[3546]_ , \new_[3549]_ ,
    \new_[3552]_ , \new_[3553]_ , \new_[3554]_ , \new_[3555]_ ,
    \new_[3556]_ , \new_[3560]_ , \new_[3561]_ , \new_[3565]_ ,
    \new_[3566]_ , \new_[3567]_ , \new_[3571]_ , \new_[3572]_ ,
    \new_[3575]_ , \new_[3578]_ , \new_[3579]_ , \new_[3580]_ ,
    \new_[3581]_ , \new_[3585]_ , \new_[3586]_ , \new_[3589]_ ,
    \new_[3592]_ , \new_[3593]_ , \new_[3594]_ , \new_[3598]_ ,
    \new_[3599]_ , \new_[3602]_ , \new_[3605]_ , \new_[3606]_ ,
    \new_[3607]_ , \new_[3608]_ , \new_[3609]_ , \new_[3610]_ ,
    \new_[3614]_ , \new_[3615]_ , \new_[3619]_ , \new_[3620]_ ,
    \new_[3621]_ , \new_[3625]_ , \new_[3626]_ , \new_[3629]_ ,
    \new_[3632]_ , \new_[3633]_ , \new_[3634]_ , \new_[3635]_ ,
    \new_[3639]_ , \new_[3640]_ , \new_[3643]_ , \new_[3646]_ ,
    \new_[3647]_ , \new_[3648]_ , \new_[3652]_ , \new_[3653]_ ,
    \new_[3656]_ , \new_[3659]_ , \new_[3660]_ , \new_[3661]_ ,
    \new_[3662]_ , \new_[3663]_ , \new_[3667]_ , \new_[3668]_ ,
    \new_[3671]_ , \new_[3674]_ , \new_[3675]_ , \new_[3676]_ ,
    \new_[3680]_ , \new_[3681]_ , \new_[3684]_ , \new_[3687]_ ,
    \new_[3688]_ , \new_[3689]_ , \new_[3690]_ , \new_[3694]_ ,
    \new_[3695]_ , \new_[3698]_ , \new_[3701]_ , \new_[3702]_ ,
    \new_[3703]_ , \new_[3707]_ , \new_[3708]_ , \new_[3711]_ ,
    \new_[3714]_ , \new_[3715]_ , \new_[3716]_ , \new_[3717]_ ,
    \new_[3718]_ , \new_[3719]_ , \new_[3720]_ , \new_[3724]_ ,
    \new_[3725]_ , \new_[3729]_ , \new_[3730]_ , \new_[3731]_ ,
    \new_[3735]_ , \new_[3736]_ , \new_[3739]_ , \new_[3742]_ ,
    \new_[3743]_ , \new_[3744]_ , \new_[3745]_ , \new_[3749]_ ,
    \new_[3750]_ , \new_[3753]_ , \new_[3756]_ , \new_[3757]_ ,
    \new_[3758]_ , \new_[3762]_ , \new_[3763]_ , \new_[3766]_ ,
    \new_[3769]_ , \new_[3770]_ , \new_[3771]_ , \new_[3772]_ ,
    \new_[3773]_ , \new_[3777]_ , \new_[3778]_ , \new_[3781]_ ,
    \new_[3784]_ , \new_[3785]_ , \new_[3786]_ , \new_[3790]_ ,
    \new_[3791]_ , \new_[3794]_ , \new_[3797]_ , \new_[3798]_ ,
    \new_[3799]_ , \new_[3800]_ , \new_[3804]_ , \new_[3805]_ ,
    \new_[3808]_ , \new_[3811]_ , \new_[3812]_ , \new_[3813]_ ,
    \new_[3817]_ , \new_[3818]_ , \new_[3821]_ , \new_[3824]_ ,
    \new_[3825]_ , \new_[3826]_ , \new_[3827]_ , \new_[3828]_ ,
    \new_[3829]_ , \new_[3833]_ , \new_[3834]_ , \new_[3838]_ ,
    \new_[3839]_ , \new_[3840]_ , \new_[3844]_ , \new_[3845]_ ,
    \new_[3848]_ , \new_[3851]_ , \new_[3852]_ , \new_[3853]_ ,
    \new_[3854]_ , \new_[3858]_ , \new_[3859]_ , \new_[3862]_ ,
    \new_[3865]_ , \new_[3866]_ , \new_[3867]_ , \new_[3871]_ ,
    \new_[3872]_ , \new_[3875]_ , \new_[3878]_ , \new_[3879]_ ,
    \new_[3880]_ , \new_[3881]_ , \new_[3882]_ , \new_[3886]_ ,
    \new_[3887]_ , \new_[3890]_ , \new_[3893]_ , \new_[3894]_ ,
    \new_[3895]_ , \new_[3899]_ , \new_[3900]_ , \new_[3903]_ ,
    \new_[3906]_ , \new_[3907]_ , \new_[3908]_ , \new_[3909]_ ,
    \new_[3913]_ , \new_[3914]_ , \new_[3917]_ , \new_[3920]_ ,
    \new_[3921]_ , \new_[3922]_ , \new_[3926]_ , \new_[3927]_ ,
    \new_[3930]_ , \new_[3933]_ , \new_[3934]_ , \new_[3935]_ ,
    \new_[3936]_ , \new_[3937]_ , \new_[3938]_ , \new_[3939]_ ,
    \new_[3940]_ , \new_[3944]_ , \new_[3945]_ , \new_[3949]_ ,
    \new_[3950]_ , \new_[3951]_ , \new_[3955]_ , \new_[3956]_ ,
    \new_[3959]_ , \new_[3962]_ , \new_[3963]_ , \new_[3964]_ ,
    \new_[3965]_ , \new_[3969]_ , \new_[3970]_ , \new_[3973]_ ,
    \new_[3976]_ , \new_[3977]_ , \new_[3978]_ , \new_[3982]_ ,
    \new_[3983]_ , \new_[3986]_ , \new_[3989]_ , \new_[3990]_ ,
    \new_[3991]_ , \new_[3992]_ , \new_[3993]_ , \new_[3997]_ ,
    \new_[3998]_ , \new_[4002]_ , \new_[4003]_ , \new_[4004]_ ,
    \new_[4008]_ , \new_[4009]_ , \new_[4012]_ , \new_[4015]_ ,
    \new_[4016]_ , \new_[4017]_ , \new_[4018]_ , \new_[4022]_ ,
    \new_[4023]_ , \new_[4026]_ , \new_[4029]_ , \new_[4030]_ ,
    \new_[4031]_ , \new_[4035]_ , \new_[4036]_ , \new_[4039]_ ,
    \new_[4042]_ , \new_[4043]_ , \new_[4044]_ , \new_[4045]_ ,
    \new_[4046]_ , \new_[4047]_ , \new_[4051]_ , \new_[4052]_ ,
    \new_[4056]_ , \new_[4057]_ , \new_[4058]_ , \new_[4062]_ ,
    \new_[4063]_ , \new_[4066]_ , \new_[4069]_ , \new_[4070]_ ,
    \new_[4071]_ , \new_[4072]_ , \new_[4076]_ , \new_[4077]_ ,
    \new_[4080]_ , \new_[4083]_ , \new_[4084]_ , \new_[4085]_ ,
    \new_[4089]_ , \new_[4090]_ , \new_[4093]_ , \new_[4096]_ ,
    \new_[4097]_ , \new_[4098]_ , \new_[4099]_ , \new_[4100]_ ,
    \new_[4104]_ , \new_[4105]_ , \new_[4108]_ , \new_[4111]_ ,
    \new_[4112]_ , \new_[4113]_ , \new_[4117]_ , \new_[4118]_ ,
    \new_[4121]_ , \new_[4124]_ , \new_[4125]_ , \new_[4126]_ ,
    \new_[4127]_ , \new_[4131]_ , \new_[4132]_ , \new_[4135]_ ,
    \new_[4138]_ , \new_[4139]_ , \new_[4140]_ , \new_[4144]_ ,
    \new_[4145]_ , \new_[4148]_ , \new_[4151]_ , \new_[4152]_ ,
    \new_[4153]_ , \new_[4154]_ , \new_[4155]_ , \new_[4156]_ ,
    \new_[4157]_ , \new_[4161]_ , \new_[4162]_ , \new_[4166]_ ,
    \new_[4167]_ , \new_[4168]_ , \new_[4172]_ , \new_[4173]_ ,
    \new_[4176]_ , \new_[4179]_ , \new_[4180]_ , \new_[4181]_ ,
    \new_[4182]_ , \new_[4186]_ , \new_[4187]_ , \new_[4190]_ ,
    \new_[4193]_ , \new_[4194]_ , \new_[4195]_ , \new_[4199]_ ,
    \new_[4200]_ , \new_[4203]_ , \new_[4206]_ , \new_[4207]_ ,
    \new_[4208]_ , \new_[4209]_ , \new_[4210]_ , \new_[4214]_ ,
    \new_[4215]_ , \new_[4218]_ , \new_[4221]_ , \new_[4222]_ ,
    \new_[4223]_ , \new_[4227]_ , \new_[4228]_ , \new_[4231]_ ,
    \new_[4234]_ , \new_[4235]_ , \new_[4236]_ , \new_[4237]_ ,
    \new_[4241]_ , \new_[4242]_ , \new_[4245]_ , \new_[4248]_ ,
    \new_[4249]_ , \new_[4250]_ , \new_[4254]_ , \new_[4255]_ ,
    \new_[4258]_ , \new_[4261]_ , \new_[4262]_ , \new_[4263]_ ,
    \new_[4264]_ , \new_[4265]_ , \new_[4266]_ , \new_[4270]_ ,
    \new_[4271]_ , \new_[4275]_ , \new_[4276]_ , \new_[4277]_ ,
    \new_[4281]_ , \new_[4282]_ , \new_[4285]_ , \new_[4288]_ ,
    \new_[4289]_ , \new_[4290]_ , \new_[4291]_ , \new_[4295]_ ,
    \new_[4296]_ , \new_[4299]_ , \new_[4302]_ , \new_[4303]_ ,
    \new_[4304]_ , \new_[4308]_ , \new_[4309]_ , \new_[4312]_ ,
    \new_[4315]_ , \new_[4316]_ , \new_[4317]_ , \new_[4318]_ ,
    \new_[4319]_ , \new_[4323]_ , \new_[4324]_ , \new_[4327]_ ,
    \new_[4330]_ , \new_[4331]_ , \new_[4332]_ , \new_[4336]_ ,
    \new_[4337]_ , \new_[4340]_ , \new_[4343]_ , \new_[4344]_ ,
    \new_[4345]_ , \new_[4346]_ , \new_[4350]_ , \new_[4351]_ ,
    \new_[4354]_ , \new_[4357]_ , \new_[4358]_ , \new_[4359]_ ,
    \new_[4363]_ , \new_[4364]_ , \new_[4367]_ , \new_[4370]_ ,
    \new_[4371]_ , \new_[4372]_ , \new_[4373]_ , \new_[4374]_ ,
    \new_[4375]_ , \new_[4376]_ , \new_[4377]_ , \new_[4378]_ ,
    \new_[4382]_ , \new_[4383]_ , \new_[4387]_ , \new_[4388]_ ,
    \new_[4389]_ , \new_[4393]_ , \new_[4394]_ , \new_[4397]_ ,
    \new_[4400]_ , \new_[4401]_ , \new_[4402]_ , \new_[4403]_ ,
    \new_[4407]_ , \new_[4408]_ , \new_[4411]_ , \new_[4414]_ ,
    \new_[4415]_ , \new_[4416]_ , \new_[4420]_ , \new_[4421]_ ,
    \new_[4424]_ , \new_[4427]_ , \new_[4428]_ , \new_[4429]_ ,
    \new_[4430]_ , \new_[4431]_ , \new_[4435]_ , \new_[4436]_ ,
    \new_[4440]_ , \new_[4441]_ , \new_[4442]_ , \new_[4446]_ ,
    \new_[4447]_ , \new_[4450]_ , \new_[4453]_ , \new_[4454]_ ,
    \new_[4455]_ , \new_[4456]_ , \new_[4460]_ , \new_[4461]_ ,
    \new_[4464]_ , \new_[4467]_ , \new_[4468]_ , \new_[4469]_ ,
    \new_[4473]_ , \new_[4474]_ , \new_[4477]_ , \new_[4480]_ ,
    \new_[4481]_ , \new_[4482]_ , \new_[4483]_ , \new_[4484]_ ,
    \new_[4485]_ , \new_[4489]_ , \new_[4490]_ , \new_[4494]_ ,
    \new_[4495]_ , \new_[4496]_ , \new_[4500]_ , \new_[4501]_ ,
    \new_[4504]_ , \new_[4507]_ , \new_[4508]_ , \new_[4509]_ ,
    \new_[4510]_ , \new_[4514]_ , \new_[4515]_ , \new_[4518]_ ,
    \new_[4521]_ , \new_[4522]_ , \new_[4523]_ , \new_[4527]_ ,
    \new_[4528]_ , \new_[4531]_ , \new_[4534]_ , \new_[4535]_ ,
    \new_[4536]_ , \new_[4537]_ , \new_[4538]_ , \new_[4542]_ ,
    \new_[4543]_ , \new_[4546]_ , \new_[4549]_ , \new_[4550]_ ,
    \new_[4551]_ , \new_[4555]_ , \new_[4556]_ , \new_[4559]_ ,
    \new_[4562]_ , \new_[4563]_ , \new_[4564]_ , \new_[4565]_ ,
    \new_[4569]_ , \new_[4570]_ , \new_[4573]_ , \new_[4576]_ ,
    \new_[4577]_ , \new_[4578]_ , \new_[4582]_ , \new_[4583]_ ,
    \new_[4586]_ , \new_[4589]_ , \new_[4590]_ , \new_[4591]_ ,
    \new_[4592]_ , \new_[4593]_ , \new_[4594]_ , \new_[4595]_ ,
    \new_[4599]_ , \new_[4600]_ , \new_[4604]_ , \new_[4605]_ ,
    \new_[4606]_ , \new_[4610]_ , \new_[4611]_ , \new_[4614]_ ,
    \new_[4617]_ , \new_[4618]_ , \new_[4619]_ , \new_[4620]_ ,
    \new_[4624]_ , \new_[4625]_ , \new_[4628]_ , \new_[4631]_ ,
    \new_[4632]_ , \new_[4633]_ , \new_[4637]_ , \new_[4638]_ ,
    \new_[4641]_ , \new_[4644]_ , \new_[4645]_ , \new_[4646]_ ,
    \new_[4647]_ , \new_[4648]_ , \new_[4652]_ , \new_[4653]_ ,
    \new_[4656]_ , \new_[4659]_ , \new_[4660]_ , \new_[4661]_ ,
    \new_[4665]_ , \new_[4666]_ , \new_[4669]_ , \new_[4672]_ ,
    \new_[4673]_ , \new_[4674]_ , \new_[4675]_ , \new_[4679]_ ,
    \new_[4680]_ , \new_[4683]_ , \new_[4686]_ , \new_[4687]_ ,
    \new_[4688]_ , \new_[4692]_ , \new_[4693]_ , \new_[4696]_ ,
    \new_[4699]_ , \new_[4700]_ , \new_[4701]_ , \new_[4702]_ ,
    \new_[4703]_ , \new_[4704]_ , \new_[4708]_ , \new_[4709]_ ,
    \new_[4713]_ , \new_[4714]_ , \new_[4715]_ , \new_[4719]_ ,
    \new_[4720]_ , \new_[4723]_ , \new_[4726]_ , \new_[4727]_ ,
    \new_[4728]_ , \new_[4729]_ , \new_[4733]_ , \new_[4734]_ ,
    \new_[4737]_ , \new_[4740]_ , \new_[4741]_ , \new_[4742]_ ,
    \new_[4746]_ , \new_[4747]_ , \new_[4750]_ , \new_[4753]_ ,
    \new_[4754]_ , \new_[4755]_ , \new_[4756]_ , \new_[4757]_ ,
    \new_[4761]_ , \new_[4762]_ , \new_[4765]_ , \new_[4768]_ ,
    \new_[4769]_ , \new_[4770]_ , \new_[4774]_ , \new_[4775]_ ,
    \new_[4778]_ , \new_[4781]_ , \new_[4782]_ , \new_[4783]_ ,
    \new_[4784]_ , \new_[4788]_ , \new_[4789]_ , \new_[4792]_ ,
    \new_[4795]_ , \new_[4796]_ , \new_[4797]_ , \new_[4801]_ ,
    \new_[4802]_ , \new_[4805]_ , \new_[4808]_ , \new_[4809]_ ,
    \new_[4810]_ , \new_[4811]_ , \new_[4812]_ , \new_[4813]_ ,
    \new_[4814]_ , \new_[4815]_ , \new_[4819]_ , \new_[4820]_ ,
    \new_[4824]_ , \new_[4825]_ , \new_[4826]_ , \new_[4830]_ ,
    \new_[4831]_ , \new_[4834]_ , \new_[4837]_ , \new_[4838]_ ,
    \new_[4839]_ , \new_[4840]_ , \new_[4844]_ , \new_[4845]_ ,
    \new_[4848]_ , \new_[4851]_ , \new_[4852]_ , \new_[4853]_ ,
    \new_[4857]_ , \new_[4858]_ , \new_[4861]_ , \new_[4864]_ ,
    \new_[4865]_ , \new_[4866]_ , \new_[4867]_ , \new_[4868]_ ,
    \new_[4872]_ , \new_[4873]_ , \new_[4877]_ , \new_[4878]_ ,
    \new_[4879]_ , \new_[4883]_ , \new_[4884]_ , \new_[4887]_ ,
    \new_[4890]_ , \new_[4891]_ , \new_[4892]_ , \new_[4893]_ ,
    \new_[4897]_ , \new_[4898]_ , \new_[4901]_ , \new_[4904]_ ,
    \new_[4905]_ , \new_[4906]_ , \new_[4910]_ , \new_[4911]_ ,
    \new_[4914]_ , \new_[4917]_ , \new_[4918]_ , \new_[4919]_ ,
    \new_[4920]_ , \new_[4921]_ , \new_[4922]_ , \new_[4926]_ ,
    \new_[4927]_ , \new_[4931]_ , \new_[4932]_ , \new_[4933]_ ,
    \new_[4937]_ , \new_[4938]_ , \new_[4941]_ , \new_[4944]_ ,
    \new_[4945]_ , \new_[4946]_ , \new_[4947]_ , \new_[4951]_ ,
    \new_[4952]_ , \new_[4955]_ , \new_[4958]_ , \new_[4959]_ ,
    \new_[4960]_ , \new_[4964]_ , \new_[4965]_ , \new_[4968]_ ,
    \new_[4971]_ , \new_[4972]_ , \new_[4973]_ , \new_[4974]_ ,
    \new_[4975]_ , \new_[4979]_ , \new_[4980]_ , \new_[4983]_ ,
    \new_[4986]_ , \new_[4987]_ , \new_[4988]_ , \new_[4992]_ ,
    \new_[4993]_ , \new_[4996]_ , \new_[4999]_ , \new_[5000]_ ,
    \new_[5001]_ , \new_[5002]_ , \new_[5006]_ , \new_[5007]_ ,
    \new_[5010]_ , \new_[5013]_ , \new_[5014]_ , \new_[5015]_ ,
    \new_[5019]_ , \new_[5020]_ , \new_[5023]_ , \new_[5026]_ ,
    \new_[5027]_ , \new_[5028]_ , \new_[5029]_ , \new_[5030]_ ,
    \new_[5031]_ , \new_[5032]_ , \new_[5036]_ , \new_[5037]_ ,
    \new_[5041]_ , \new_[5042]_ , \new_[5043]_ , \new_[5047]_ ,
    \new_[5048]_ , \new_[5051]_ , \new_[5054]_ , \new_[5055]_ ,
    \new_[5056]_ , \new_[5057]_ , \new_[5061]_ , \new_[5062]_ ,
    \new_[5065]_ , \new_[5068]_ , \new_[5069]_ , \new_[5070]_ ,
    \new_[5074]_ , \new_[5075]_ , \new_[5078]_ , \new_[5081]_ ,
    \new_[5082]_ , \new_[5083]_ , \new_[5084]_ , \new_[5085]_ ,
    \new_[5089]_ , \new_[5090]_ , \new_[5093]_ , \new_[5096]_ ,
    \new_[5097]_ , \new_[5098]_ , \new_[5102]_ , \new_[5103]_ ,
    \new_[5106]_ , \new_[5109]_ , \new_[5110]_ , \new_[5111]_ ,
    \new_[5112]_ , \new_[5116]_ , \new_[5117]_ , \new_[5120]_ ,
    \new_[5123]_ , \new_[5124]_ , \new_[5125]_ , \new_[5129]_ ,
    \new_[5130]_ , \new_[5133]_ , \new_[5136]_ , \new_[5137]_ ,
    \new_[5138]_ , \new_[5139]_ , \new_[5140]_ , \new_[5141]_ ,
    \new_[5145]_ , \new_[5146]_ , \new_[5150]_ , \new_[5151]_ ,
    \new_[5152]_ , \new_[5156]_ , \new_[5157]_ , \new_[5160]_ ,
    \new_[5163]_ , \new_[5164]_ , \new_[5165]_ , \new_[5166]_ ,
    \new_[5170]_ , \new_[5171]_ , \new_[5174]_ , \new_[5177]_ ,
    \new_[5178]_ , \new_[5179]_ , \new_[5183]_ , \new_[5184]_ ,
    \new_[5187]_ , \new_[5190]_ , \new_[5191]_ , \new_[5192]_ ,
    \new_[5193]_ , \new_[5194]_ , \new_[5198]_ , \new_[5199]_ ,
    \new_[5202]_ , \new_[5205]_ , \new_[5206]_ , \new_[5207]_ ,
    \new_[5211]_ , \new_[5212]_ , \new_[5215]_ , \new_[5218]_ ,
    \new_[5219]_ , \new_[5220]_ , \new_[5221]_ , \new_[5225]_ ,
    \new_[5226]_ , \new_[5229]_ , \new_[5232]_ , \new_[5233]_ ,
    \new_[5234]_ , \new_[5238]_ , \new_[5239]_ , \new_[5242]_ ,
    \new_[5245]_ , \new_[5246]_ , \new_[5247]_ , \new_[5248]_ ,
    \new_[5249]_ , \new_[5250]_ , \new_[5251]_ , \new_[5252]_ ,
    \new_[5253]_ , \new_[5254]_ , \new_[5257]_ , \new_[5260]_ ,
    \new_[5263]_ , \new_[5266]_ , \new_[5269]_ , \new_[5272]_ ,
    \new_[5275]_ , \new_[5278]_ , \new_[5281]_ , \new_[5284]_ ,
    \new_[5287]_ , \new_[5290]_ , \new_[5293]_ , \new_[5297]_ ,
    \new_[5298]_ , \new_[5301]_ , \new_[5305]_ , \new_[5306]_ ,
    \new_[5310]_ , \new_[5311]_ , \new_[5315]_ , \new_[5316]_ ,
    \new_[5320]_ , \new_[5321]_ , \new_[5325]_ , \new_[5326]_ ,
    \new_[5330]_ , \new_[5331]_ , \new_[5335]_ , \new_[5336]_ ,
    \new_[5340]_ , \new_[5341]_ , \new_[5345]_ , \new_[5346]_ ,
    \new_[5350]_ , \new_[5351]_ , \new_[5355]_ , \new_[5356]_ ,
    \new_[5360]_ , \new_[5361]_ , \new_[5365]_ , \new_[5366]_ ,
    \new_[5370]_ , \new_[5371]_ , \new_[5375]_ , \new_[5376]_ ,
    \new_[5380]_ , \new_[5381]_ , \new_[5385]_ , \new_[5386]_ ,
    \new_[5390]_ , \new_[5391]_ , \new_[5395]_ , \new_[5396]_ ,
    \new_[5400]_ , \new_[5401]_ , \new_[5405]_ , \new_[5406]_ ,
    \new_[5410]_ , \new_[5411]_ , \new_[5415]_ , \new_[5416]_ ,
    \new_[5420]_ , \new_[5421]_ , \new_[5425]_ , \new_[5426]_ ,
    \new_[5430]_ , \new_[5431]_ , \new_[5434]_ , \new_[5437]_ ,
    \new_[5438]_ , \new_[5442]_ , \new_[5443]_ , \new_[5446]_ ,
    \new_[5449]_ , \new_[5450]_ , \new_[5454]_ , \new_[5455]_ ,
    \new_[5458]_ , \new_[5461]_ , \new_[5462]_ , \new_[5466]_ ,
    \new_[5467]_ , \new_[5470]_ , \new_[5473]_ , \new_[5474]_ ,
    \new_[5477]_ , \new_[5480]_ , \new_[5481]_ , \new_[5484]_ ,
    \new_[5488]_ , \new_[5489]_ , \new_[5490]_ , \new_[5493]_ ,
    \new_[5496]_ , \new_[5497]_ , \new_[5500]_ , \new_[5504]_ ,
    \new_[5505]_ , \new_[5506]_ , \new_[5509]_ , \new_[5512]_ ,
    \new_[5513]_ , \new_[5516]_ , \new_[5520]_ , \new_[5521]_ ,
    \new_[5522]_ , \new_[5525]_ , \new_[5528]_ , \new_[5529]_ ,
    \new_[5532]_ , \new_[5536]_ , \new_[5537]_ , \new_[5538]_ ,
    \new_[5541]_ , \new_[5544]_ , \new_[5545]_ , \new_[5548]_ ,
    \new_[5552]_ , \new_[5553]_ , \new_[5554]_ , \new_[5557]_ ,
    \new_[5560]_ , \new_[5561]_ , \new_[5564]_ , \new_[5568]_ ,
    \new_[5569]_ , \new_[5570]_ , \new_[5573]_ , \new_[5576]_ ,
    \new_[5577]_ , \new_[5580]_ , \new_[5584]_ , \new_[5585]_ ,
    \new_[5586]_ , \new_[5589]_ , \new_[5592]_ , \new_[5593]_ ,
    \new_[5596]_ , \new_[5600]_ , \new_[5601]_ , \new_[5602]_ ,
    \new_[5605]_ , \new_[5608]_ , \new_[5609]_ , \new_[5612]_ ,
    \new_[5616]_ , \new_[5617]_ , \new_[5618]_ , \new_[5621]_ ,
    \new_[5624]_ , \new_[5625]_ , \new_[5628]_ , \new_[5632]_ ,
    \new_[5633]_ , \new_[5634]_ , \new_[5637]_ , \new_[5640]_ ,
    \new_[5641]_ , \new_[5644]_ , \new_[5648]_ , \new_[5649]_ ,
    \new_[5650]_ , \new_[5653]_ , \new_[5656]_ , \new_[5657]_ ,
    \new_[5660]_ , \new_[5664]_ , \new_[5665]_ , \new_[5666]_ ,
    \new_[5669]_ , \new_[5672]_ , \new_[5673]_ , \new_[5676]_ ,
    \new_[5680]_ , \new_[5681]_ , \new_[5682]_ , \new_[5685]_ ,
    \new_[5688]_ , \new_[5689]_ , \new_[5692]_ , \new_[5696]_ ,
    \new_[5697]_ , \new_[5698]_ , \new_[5701]_ , \new_[5704]_ ,
    \new_[5705]_ , \new_[5708]_ , \new_[5712]_ , \new_[5713]_ ,
    \new_[5714]_ , \new_[5717]_ , \new_[5720]_ , \new_[5721]_ ,
    \new_[5724]_ , \new_[5728]_ , \new_[5729]_ , \new_[5730]_ ,
    \new_[5733]_ , \new_[5737]_ , \new_[5738]_ , \new_[5739]_ ,
    \new_[5742]_ , \new_[5746]_ , \new_[5747]_ , \new_[5748]_ ,
    \new_[5751]_ , \new_[5755]_ , \new_[5756]_ , \new_[5757]_ ,
    \new_[5760]_ , \new_[5764]_ , \new_[5765]_ , \new_[5766]_ ,
    \new_[5769]_ , \new_[5773]_ , \new_[5774]_ , \new_[5775]_ ,
    \new_[5778]_ , \new_[5782]_ , \new_[5783]_ , \new_[5784]_ ,
    \new_[5787]_ , \new_[5791]_ , \new_[5792]_ , \new_[5793]_ ,
    \new_[5796]_ , \new_[5800]_ , \new_[5801]_ , \new_[5802]_ ,
    \new_[5805]_ , \new_[5809]_ , \new_[5810]_ , \new_[5811]_ ,
    \new_[5814]_ , \new_[5818]_ , \new_[5819]_ , \new_[5820]_ ,
    \new_[5823]_ , \new_[5827]_ , \new_[5828]_ , \new_[5829]_ ,
    \new_[5832]_ , \new_[5836]_ , \new_[5837]_ , \new_[5838]_ ,
    \new_[5841]_ , \new_[5845]_ , \new_[5846]_ , \new_[5847]_ ,
    \new_[5850]_ , \new_[5854]_ , \new_[5855]_ , \new_[5856]_ ,
    \new_[5859]_ , \new_[5863]_ , \new_[5864]_ , \new_[5865]_ ,
    \new_[5868]_ , \new_[5872]_ , \new_[5873]_ , \new_[5874]_ ,
    \new_[5877]_ , \new_[5881]_ , \new_[5882]_ , \new_[5883]_ ,
    \new_[5886]_ , \new_[5890]_ , \new_[5891]_ , \new_[5892]_ ,
    \new_[5895]_ , \new_[5899]_ , \new_[5900]_ , \new_[5901]_ ,
    \new_[5904]_ , \new_[5908]_ , \new_[5909]_ , \new_[5910]_ ,
    \new_[5913]_ , \new_[5917]_ , \new_[5918]_ , \new_[5919]_ ,
    \new_[5922]_ , \new_[5926]_ , \new_[5927]_ , \new_[5928]_ ,
    \new_[5931]_ , \new_[5935]_ , \new_[5936]_ , \new_[5937]_ ,
    \new_[5940]_ , \new_[5944]_ , \new_[5945]_ , \new_[5946]_ ,
    \new_[5949]_ , \new_[5953]_ , \new_[5954]_ , \new_[5955]_ ,
    \new_[5958]_ , \new_[5962]_ , \new_[5963]_ , \new_[5964]_ ,
    \new_[5967]_ , \new_[5971]_ , \new_[5972]_ , \new_[5973]_ ,
    \new_[5976]_ , \new_[5980]_ , \new_[5981]_ , \new_[5982]_ ,
    \new_[5985]_ , \new_[5989]_ , \new_[5990]_ , \new_[5991]_ ,
    \new_[5994]_ , \new_[5998]_ , \new_[5999]_ , \new_[6000]_ ,
    \new_[6003]_ , \new_[6007]_ , \new_[6008]_ , \new_[6009]_ ,
    \new_[6012]_ , \new_[6016]_ , \new_[6017]_ , \new_[6018]_ ,
    \new_[6021]_ , \new_[6025]_ , \new_[6026]_ , \new_[6027]_ ,
    \new_[6030]_ , \new_[6034]_ , \new_[6035]_ , \new_[6036]_ ,
    \new_[6039]_ , \new_[6043]_ , \new_[6044]_ , \new_[6045]_ ,
    \new_[6048]_ , \new_[6052]_ , \new_[6053]_ , \new_[6054]_ ,
    \new_[6057]_ , \new_[6061]_ , \new_[6062]_ , \new_[6063]_ ,
    \new_[6066]_ , \new_[6070]_ , \new_[6071]_ , \new_[6072]_ ,
    \new_[6075]_ , \new_[6079]_ , \new_[6080]_ , \new_[6081]_ ,
    \new_[6084]_ , \new_[6088]_ , \new_[6089]_ , \new_[6090]_ ,
    \new_[6093]_ , \new_[6097]_ , \new_[6098]_ , \new_[6099]_ ,
    \new_[6102]_ , \new_[6106]_ , \new_[6107]_ , \new_[6108]_ ,
    \new_[6111]_ , \new_[6115]_ , \new_[6116]_ , \new_[6117]_ ,
    \new_[6120]_ , \new_[6124]_ , \new_[6125]_ , \new_[6126]_ ,
    \new_[6129]_ , \new_[6133]_ , \new_[6134]_ , \new_[6135]_ ,
    \new_[6138]_ , \new_[6142]_ , \new_[6143]_ , \new_[6144]_ ,
    \new_[6147]_ , \new_[6151]_ , \new_[6152]_ , \new_[6153]_ ,
    \new_[6156]_ , \new_[6160]_ , \new_[6161]_ , \new_[6162]_ ,
    \new_[6165]_ , \new_[6169]_ , \new_[6170]_ , \new_[6171]_ ,
    \new_[6174]_ , \new_[6178]_ , \new_[6179]_ , \new_[6180]_ ,
    \new_[6183]_ , \new_[6187]_ , \new_[6188]_ , \new_[6189]_ ,
    \new_[6192]_ , \new_[6196]_ , \new_[6197]_ , \new_[6198]_ ,
    \new_[6201]_ , \new_[6205]_ , \new_[6206]_ , \new_[6207]_ ,
    \new_[6210]_ , \new_[6214]_ , \new_[6215]_ , \new_[6216]_ ,
    \new_[6219]_ , \new_[6223]_ , \new_[6224]_ , \new_[6225]_ ,
    \new_[6228]_ , \new_[6232]_ , \new_[6233]_ , \new_[6234]_ ,
    \new_[6237]_ , \new_[6241]_ , \new_[6242]_ , \new_[6243]_ ,
    \new_[6246]_ , \new_[6250]_ , \new_[6251]_ , \new_[6252]_ ,
    \new_[6255]_ , \new_[6259]_ , \new_[6260]_ , \new_[6261]_ ,
    \new_[6264]_ , \new_[6268]_ , \new_[6269]_ , \new_[6270]_ ,
    \new_[6273]_ , \new_[6277]_ , \new_[6278]_ , \new_[6279]_ ,
    \new_[6282]_ , \new_[6286]_ , \new_[6287]_ , \new_[6288]_ ,
    \new_[6291]_ , \new_[6295]_ , \new_[6296]_ , \new_[6297]_ ,
    \new_[6300]_ , \new_[6304]_ , \new_[6305]_ , \new_[6306]_ ,
    \new_[6309]_ , \new_[6313]_ , \new_[6314]_ , \new_[6315]_ ,
    \new_[6318]_ , \new_[6322]_ , \new_[6323]_ , \new_[6324]_ ,
    \new_[6327]_ , \new_[6331]_ , \new_[6332]_ , \new_[6333]_ ,
    \new_[6336]_ , \new_[6340]_ , \new_[6341]_ , \new_[6342]_ ,
    \new_[6345]_ , \new_[6349]_ , \new_[6350]_ , \new_[6351]_ ,
    \new_[6354]_ , \new_[6358]_ , \new_[6359]_ , \new_[6360]_ ,
    \new_[6363]_ , \new_[6367]_ , \new_[6368]_ , \new_[6369]_ ,
    \new_[6372]_ , \new_[6376]_ , \new_[6377]_ , \new_[6378]_ ,
    \new_[6381]_ , \new_[6385]_ , \new_[6386]_ , \new_[6387]_ ,
    \new_[6390]_ , \new_[6394]_ , \new_[6395]_ , \new_[6396]_ ,
    \new_[6399]_ , \new_[6403]_ , \new_[6404]_ , \new_[6405]_ ,
    \new_[6408]_ , \new_[6412]_ , \new_[6413]_ , \new_[6414]_ ,
    \new_[6417]_ , \new_[6421]_ , \new_[6422]_ , \new_[6423]_ ,
    \new_[6426]_ , \new_[6430]_ , \new_[6431]_ , \new_[6432]_ ,
    \new_[6435]_ , \new_[6439]_ , \new_[6440]_ , \new_[6441]_ ,
    \new_[6444]_ , \new_[6448]_ , \new_[6449]_ , \new_[6450]_ ,
    \new_[6453]_ , \new_[6457]_ , \new_[6458]_ , \new_[6459]_ ,
    \new_[6462]_ , \new_[6466]_ , \new_[6467]_ , \new_[6468]_ ,
    \new_[6471]_ , \new_[6475]_ , \new_[6476]_ , \new_[6477]_ ,
    \new_[6480]_ , \new_[6484]_ , \new_[6485]_ , \new_[6486]_ ,
    \new_[6489]_ , \new_[6493]_ , \new_[6494]_ , \new_[6495]_ ,
    \new_[6498]_ , \new_[6502]_ , \new_[6503]_ , \new_[6504]_ ,
    \new_[6507]_ , \new_[6511]_ , \new_[6512]_ , \new_[6513]_ ,
    \new_[6516]_ , \new_[6520]_ , \new_[6521]_ , \new_[6522]_ ,
    \new_[6525]_ , \new_[6529]_ , \new_[6530]_ , \new_[6531]_ ,
    \new_[6534]_ , \new_[6538]_ , \new_[6539]_ , \new_[6540]_ ,
    \new_[6543]_ , \new_[6547]_ , \new_[6548]_ , \new_[6549]_ ,
    \new_[6552]_ , \new_[6556]_ , \new_[6557]_ , \new_[6558]_ ,
    \new_[6561]_ , \new_[6565]_ , \new_[6566]_ , \new_[6567]_ ,
    \new_[6570]_ , \new_[6574]_ , \new_[6575]_ , \new_[6576]_ ,
    \new_[6579]_ , \new_[6583]_ , \new_[6584]_ , \new_[6585]_ ,
    \new_[6588]_ , \new_[6592]_ , \new_[6593]_ , \new_[6594]_ ,
    \new_[6597]_ , \new_[6601]_ , \new_[6602]_ , \new_[6603]_ ,
    \new_[6607]_ , \new_[6608]_ , \new_[6612]_ , \new_[6613]_ ,
    \new_[6614]_ , \new_[6617]_ , \new_[6621]_ , \new_[6622]_ ,
    \new_[6623]_ , \new_[6627]_ , \new_[6628]_ , \new_[6632]_ ,
    \new_[6633]_ , \new_[6634]_ , \new_[6637]_ , \new_[6641]_ ,
    \new_[6642]_ , \new_[6643]_ , \new_[6647]_ , \new_[6648]_ ,
    \new_[6652]_ , \new_[6653]_ , \new_[6654]_ , \new_[6657]_ ,
    \new_[6661]_ , \new_[6662]_ , \new_[6663]_ , \new_[6667]_ ,
    \new_[6668]_ , \new_[6672]_ , \new_[6673]_ , \new_[6674]_ ,
    \new_[6677]_ , \new_[6681]_ , \new_[6682]_ , \new_[6683]_ ,
    \new_[6687]_ , \new_[6688]_ , \new_[6692]_ , \new_[6693]_ ,
    \new_[6694]_ , \new_[6697]_ , \new_[6701]_ , \new_[6702]_ ,
    \new_[6703]_ , \new_[6707]_ , \new_[6708]_ , \new_[6712]_ ,
    \new_[6713]_ , \new_[6714]_ , \new_[6717]_ , \new_[6721]_ ,
    \new_[6722]_ , \new_[6723]_ , \new_[6727]_ , \new_[6728]_ ,
    \new_[6732]_ , \new_[6733]_ , \new_[6734]_ , \new_[6737]_ ,
    \new_[6741]_ , \new_[6742]_ , \new_[6743]_ , \new_[6747]_ ,
    \new_[6748]_ , \new_[6752]_ , \new_[6753]_ , \new_[6754]_ ,
    \new_[6757]_ , \new_[6761]_ , \new_[6762]_ , \new_[6763]_ ,
    \new_[6767]_ , \new_[6768]_ , \new_[6772]_ , \new_[6773]_ ,
    \new_[6774]_ , \new_[6777]_ , \new_[6781]_ , \new_[6782]_ ,
    \new_[6783]_ , \new_[6787]_ , \new_[6788]_ , \new_[6792]_ ,
    \new_[6793]_ , \new_[6794]_ , \new_[6797]_ , \new_[6801]_ ,
    \new_[6802]_ , \new_[6803]_ , \new_[6807]_ , \new_[6808]_ ,
    \new_[6812]_ , \new_[6813]_ , \new_[6814]_ , \new_[6817]_ ,
    \new_[6821]_ , \new_[6822]_ , \new_[6823]_ , \new_[6827]_ ,
    \new_[6828]_ , \new_[6832]_ , \new_[6833]_ , \new_[6834]_ ,
    \new_[6837]_ , \new_[6841]_ , \new_[6842]_ , \new_[6843]_ ,
    \new_[6847]_ , \new_[6848]_ , \new_[6852]_ , \new_[6853]_ ,
    \new_[6854]_ , \new_[6857]_ , \new_[6861]_ , \new_[6862]_ ,
    \new_[6863]_ , \new_[6867]_ , \new_[6868]_ , \new_[6872]_ ,
    \new_[6873]_ , \new_[6874]_ , \new_[6877]_ , \new_[6881]_ ,
    \new_[6882]_ , \new_[6883]_ , \new_[6887]_ , \new_[6888]_ ,
    \new_[6892]_ , \new_[6893]_ , \new_[6894]_ , \new_[6897]_ ,
    \new_[6901]_ , \new_[6902]_ , \new_[6903]_ , \new_[6907]_ ,
    \new_[6908]_ , \new_[6912]_ , \new_[6913]_ , \new_[6914]_ ,
    \new_[6917]_ , \new_[6921]_ , \new_[6922]_ , \new_[6923]_ ,
    \new_[6927]_ , \new_[6928]_ , \new_[6932]_ , \new_[6933]_ ,
    \new_[6934]_ , \new_[6937]_ , \new_[6941]_ , \new_[6942]_ ,
    \new_[6943]_ , \new_[6947]_ , \new_[6948]_ , \new_[6952]_ ,
    \new_[6953]_ , \new_[6954]_ , \new_[6957]_ , \new_[6961]_ ,
    \new_[6962]_ , \new_[6963]_ , \new_[6967]_ , \new_[6968]_ ,
    \new_[6972]_ , \new_[6973]_ , \new_[6974]_ , \new_[6977]_ ,
    \new_[6981]_ , \new_[6982]_ , \new_[6983]_ , \new_[6987]_ ,
    \new_[6988]_ , \new_[6992]_ , \new_[6993]_ , \new_[6994]_ ,
    \new_[6997]_ , \new_[7001]_ , \new_[7002]_ , \new_[7003]_ ,
    \new_[7007]_ , \new_[7008]_ , \new_[7012]_ , \new_[7013]_ ,
    \new_[7014]_ , \new_[7017]_ , \new_[7021]_ , \new_[7022]_ ,
    \new_[7023]_ , \new_[7027]_ , \new_[7028]_ , \new_[7032]_ ,
    \new_[7033]_ , \new_[7034]_ , \new_[7037]_ , \new_[7041]_ ,
    \new_[7042]_ , \new_[7043]_ , \new_[7047]_ , \new_[7048]_ ,
    \new_[7052]_ , \new_[7053]_ , \new_[7054]_ , \new_[7057]_ ,
    \new_[7061]_ , \new_[7062]_ , \new_[7063]_ , \new_[7067]_ ,
    \new_[7068]_ , \new_[7072]_ , \new_[7073]_ , \new_[7074]_ ,
    \new_[7077]_ , \new_[7081]_ , \new_[7082]_ , \new_[7083]_ ,
    \new_[7087]_ , \new_[7088]_ , \new_[7092]_ , \new_[7093]_ ,
    \new_[7094]_ , \new_[7097]_ , \new_[7101]_ , \new_[7102]_ ,
    \new_[7103]_ , \new_[7107]_ , \new_[7108]_ , \new_[7112]_ ,
    \new_[7113]_ , \new_[7114]_ , \new_[7117]_ , \new_[7121]_ ,
    \new_[7122]_ , \new_[7123]_ , \new_[7127]_ , \new_[7128]_ ,
    \new_[7132]_ , \new_[7133]_ , \new_[7134]_ , \new_[7137]_ ,
    \new_[7141]_ , \new_[7142]_ , \new_[7143]_ , \new_[7147]_ ,
    \new_[7148]_ , \new_[7152]_ , \new_[7153]_ , \new_[7154]_ ,
    \new_[7157]_ , \new_[7161]_ , \new_[7162]_ , \new_[7163]_ ,
    \new_[7167]_ , \new_[7168]_ , \new_[7172]_ , \new_[7173]_ ,
    \new_[7174]_ , \new_[7177]_ , \new_[7181]_ , \new_[7182]_ ,
    \new_[7183]_ , \new_[7187]_ , \new_[7188]_ , \new_[7192]_ ,
    \new_[7193]_ , \new_[7194]_ , \new_[7197]_ , \new_[7201]_ ,
    \new_[7202]_ , \new_[7203]_ , \new_[7207]_ , \new_[7208]_ ,
    \new_[7212]_ , \new_[7213]_ , \new_[7214]_ , \new_[7217]_ ,
    \new_[7221]_ , \new_[7222]_ , \new_[7223]_ , \new_[7227]_ ,
    \new_[7228]_ , \new_[7232]_ , \new_[7233]_ , \new_[7234]_ ,
    \new_[7237]_ , \new_[7241]_ , \new_[7242]_ , \new_[7243]_ ,
    \new_[7247]_ , \new_[7248]_ , \new_[7252]_ , \new_[7253]_ ,
    \new_[7254]_ , \new_[7257]_ , \new_[7261]_ , \new_[7262]_ ,
    \new_[7263]_ , \new_[7267]_ , \new_[7268]_ , \new_[7272]_ ,
    \new_[7273]_ , \new_[7274]_ , \new_[7277]_ , \new_[7281]_ ,
    \new_[7282]_ , \new_[7283]_ , \new_[7287]_ , \new_[7288]_ ,
    \new_[7292]_ , \new_[7293]_ , \new_[7294]_ , \new_[7297]_ ,
    \new_[7301]_ , \new_[7302]_ , \new_[7303]_ , \new_[7307]_ ,
    \new_[7308]_ , \new_[7312]_ , \new_[7313]_ , \new_[7314]_ ,
    \new_[7317]_ , \new_[7321]_ , \new_[7322]_ , \new_[7323]_ ,
    \new_[7327]_ , \new_[7328]_ , \new_[7332]_ , \new_[7333]_ ,
    \new_[7334]_ , \new_[7337]_ , \new_[7341]_ , \new_[7342]_ ,
    \new_[7343]_ , \new_[7347]_ , \new_[7348]_ , \new_[7352]_ ,
    \new_[7353]_ , \new_[7354]_ , \new_[7357]_ , \new_[7361]_ ,
    \new_[7362]_ , \new_[7363]_ , \new_[7367]_ , \new_[7368]_ ,
    \new_[7372]_ , \new_[7373]_ , \new_[7374]_ , \new_[7377]_ ,
    \new_[7381]_ , \new_[7382]_ , \new_[7383]_ , \new_[7387]_ ,
    \new_[7388]_ , \new_[7392]_ , \new_[7393]_ , \new_[7394]_ ,
    \new_[7397]_ , \new_[7401]_ , \new_[7402]_ , \new_[7403]_ ,
    \new_[7407]_ , \new_[7408]_ , \new_[7412]_ , \new_[7413]_ ,
    \new_[7414]_ , \new_[7417]_ , \new_[7421]_ , \new_[7422]_ ,
    \new_[7423]_ , \new_[7427]_ , \new_[7428]_ , \new_[7432]_ ,
    \new_[7433]_ , \new_[7434]_ , \new_[7437]_ , \new_[7441]_ ,
    \new_[7442]_ , \new_[7443]_ , \new_[7447]_ , \new_[7448]_ ,
    \new_[7452]_ , \new_[7453]_ , \new_[7454]_ , \new_[7457]_ ,
    \new_[7461]_ , \new_[7462]_ , \new_[7463]_ , \new_[7467]_ ,
    \new_[7468]_ , \new_[7472]_ , \new_[7473]_ , \new_[7474]_ ,
    \new_[7477]_ , \new_[7481]_ , \new_[7482]_ , \new_[7483]_ ,
    \new_[7487]_ , \new_[7488]_ , \new_[7492]_ , \new_[7493]_ ,
    \new_[7494]_ , \new_[7497]_ , \new_[7501]_ , \new_[7502]_ ,
    \new_[7503]_ , \new_[7507]_ , \new_[7508]_ , \new_[7512]_ ,
    \new_[7513]_ , \new_[7514]_ , \new_[7517]_ , \new_[7521]_ ,
    \new_[7522]_ , \new_[7523]_ , \new_[7527]_ , \new_[7528]_ ,
    \new_[7532]_ , \new_[7533]_ , \new_[7534]_ , \new_[7537]_ ,
    \new_[7541]_ , \new_[7542]_ , \new_[7543]_ , \new_[7547]_ ,
    \new_[7548]_ , \new_[7552]_ , \new_[7553]_ , \new_[7554]_ ,
    \new_[7557]_ , \new_[7561]_ , \new_[7562]_ , \new_[7563]_ ,
    \new_[7567]_ , \new_[7568]_ , \new_[7572]_ , \new_[7573]_ ,
    \new_[7574]_ , \new_[7577]_ , \new_[7581]_ , \new_[7582]_ ,
    \new_[7583]_ , \new_[7587]_ , \new_[7588]_ , \new_[7592]_ ,
    \new_[7593]_ , \new_[7594]_ , \new_[7597]_ , \new_[7601]_ ,
    \new_[7602]_ , \new_[7603]_ , \new_[7607]_ , \new_[7608]_ ,
    \new_[7612]_ , \new_[7613]_ , \new_[7614]_ , \new_[7617]_ ,
    \new_[7621]_ , \new_[7622]_ , \new_[7623]_ , \new_[7627]_ ,
    \new_[7628]_ , \new_[7632]_ , \new_[7633]_ , \new_[7634]_ ,
    \new_[7637]_ , \new_[7641]_ , \new_[7642]_ , \new_[7643]_ ,
    \new_[7647]_ , \new_[7648]_ , \new_[7652]_ , \new_[7653]_ ,
    \new_[7654]_ , \new_[7657]_ , \new_[7661]_ , \new_[7662]_ ,
    \new_[7663]_ , \new_[7667]_ , \new_[7668]_ , \new_[7672]_ ,
    \new_[7673]_ , \new_[7674]_ , \new_[7677]_ , \new_[7681]_ ,
    \new_[7682]_ , \new_[7683]_ , \new_[7687]_ , \new_[7688]_ ,
    \new_[7692]_ , \new_[7693]_ , \new_[7694]_ , \new_[7697]_ ,
    \new_[7701]_ , \new_[7702]_ , \new_[7703]_ , \new_[7707]_ ,
    \new_[7708]_ , \new_[7712]_ , \new_[7713]_ , \new_[7714]_ ,
    \new_[7717]_ , \new_[7721]_ , \new_[7722]_ , \new_[7723]_ ,
    \new_[7727]_ , \new_[7728]_ , \new_[7732]_ , \new_[7733]_ ,
    \new_[7734]_ , \new_[7737]_ , \new_[7741]_ , \new_[7742]_ ,
    \new_[7743]_ , \new_[7747]_ , \new_[7748]_ , \new_[7752]_ ,
    \new_[7753]_ , \new_[7754]_ , \new_[7757]_ , \new_[7761]_ ,
    \new_[7762]_ , \new_[7763]_ , \new_[7767]_ , \new_[7768]_ ,
    \new_[7772]_ , \new_[7773]_ , \new_[7774]_ , \new_[7777]_ ,
    \new_[7781]_ , \new_[7782]_ , \new_[7783]_ , \new_[7787]_ ,
    \new_[7788]_ , \new_[7792]_ , \new_[7793]_ , \new_[7794]_ ,
    \new_[7797]_ , \new_[7801]_ , \new_[7802]_ , \new_[7803]_ ,
    \new_[7807]_ , \new_[7808]_ , \new_[7812]_ , \new_[7813]_ ,
    \new_[7814]_ , \new_[7817]_ , \new_[7821]_ , \new_[7822]_ ,
    \new_[7823]_ , \new_[7827]_ , \new_[7828]_ , \new_[7832]_ ,
    \new_[7833]_ , \new_[7834]_ , \new_[7837]_ , \new_[7841]_ ,
    \new_[7842]_ , \new_[7843]_ , \new_[7847]_ , \new_[7848]_ ,
    \new_[7852]_ , \new_[7853]_ , \new_[7854]_ , \new_[7857]_ ,
    \new_[7861]_ , \new_[7862]_ , \new_[7863]_ , \new_[7867]_ ,
    \new_[7868]_ , \new_[7872]_ , \new_[7873]_ , \new_[7874]_ ,
    \new_[7877]_ , \new_[7881]_ , \new_[7882]_ , \new_[7883]_ ,
    \new_[7887]_ , \new_[7888]_ , \new_[7892]_ , \new_[7893]_ ,
    \new_[7894]_ , \new_[7897]_ , \new_[7901]_ , \new_[7902]_ ,
    \new_[7903]_ , \new_[7907]_ , \new_[7908]_ , \new_[7912]_ ,
    \new_[7913]_ , \new_[7914]_ , \new_[7917]_ , \new_[7921]_ ,
    \new_[7922]_ , \new_[7923]_ , \new_[7927]_ , \new_[7928]_ ,
    \new_[7932]_ , \new_[7933]_ , \new_[7934]_ , \new_[7937]_ ,
    \new_[7941]_ , \new_[7942]_ , \new_[7943]_ , \new_[7947]_ ,
    \new_[7948]_ , \new_[7952]_ , \new_[7953]_ , \new_[7954]_ ,
    \new_[7957]_ , \new_[7961]_ , \new_[7962]_ , \new_[7963]_ ,
    \new_[7967]_ , \new_[7968]_ , \new_[7972]_ , \new_[7973]_ ,
    \new_[7974]_ , \new_[7977]_ , \new_[7981]_ , \new_[7982]_ ,
    \new_[7983]_ , \new_[7987]_ , \new_[7988]_ , \new_[7992]_ ,
    \new_[7993]_ , \new_[7994]_ , \new_[7997]_ , \new_[8001]_ ,
    \new_[8002]_ , \new_[8003]_ , \new_[8007]_ , \new_[8008]_ ,
    \new_[8012]_ , \new_[8013]_ , \new_[8014]_ , \new_[8017]_ ,
    \new_[8021]_ , \new_[8022]_ , \new_[8023]_ , \new_[8027]_ ,
    \new_[8028]_ , \new_[8032]_ , \new_[8033]_ , \new_[8034]_ ,
    \new_[8037]_ , \new_[8041]_ , \new_[8042]_ , \new_[8043]_ ,
    \new_[8047]_ , \new_[8048]_ , \new_[8052]_ , \new_[8053]_ ,
    \new_[8054]_ , \new_[8057]_ , \new_[8061]_ , \new_[8062]_ ,
    \new_[8063]_ , \new_[8067]_ , \new_[8068]_ , \new_[8072]_ ,
    \new_[8073]_ , \new_[8074]_ , \new_[8077]_ , \new_[8081]_ ,
    \new_[8082]_ , \new_[8083]_ , \new_[8087]_ , \new_[8088]_ ,
    \new_[8092]_ , \new_[8093]_ , \new_[8094]_ , \new_[8097]_ ,
    \new_[8101]_ , \new_[8102]_ , \new_[8103]_ , \new_[8107]_ ,
    \new_[8108]_ , \new_[8112]_ , \new_[8113]_ , \new_[8114]_ ,
    \new_[8117]_ , \new_[8121]_ , \new_[8122]_ , \new_[8123]_ ,
    \new_[8127]_ , \new_[8128]_ , \new_[8132]_ , \new_[8133]_ ,
    \new_[8134]_ , \new_[8137]_ , \new_[8141]_ , \new_[8142]_ ,
    \new_[8143]_ , \new_[8147]_ , \new_[8148]_ , \new_[8152]_ ,
    \new_[8153]_ , \new_[8154]_ , \new_[8157]_ , \new_[8161]_ ,
    \new_[8162]_ , \new_[8163]_ , \new_[8167]_ , \new_[8168]_ ,
    \new_[8172]_ , \new_[8173]_ , \new_[8174]_ , \new_[8177]_ ,
    \new_[8181]_ , \new_[8182]_ , \new_[8183]_ , \new_[8187]_ ,
    \new_[8188]_ , \new_[8192]_ , \new_[8193]_ , \new_[8194]_ ,
    \new_[8197]_ , \new_[8201]_ , \new_[8202]_ , \new_[8203]_ ,
    \new_[8207]_ , \new_[8208]_ , \new_[8212]_ , \new_[8213]_ ,
    \new_[8214]_ , \new_[8217]_ , \new_[8221]_ , \new_[8222]_ ,
    \new_[8223]_ , \new_[8227]_ , \new_[8228]_ , \new_[8232]_ ,
    \new_[8233]_ , \new_[8234]_ , \new_[8237]_ , \new_[8241]_ ,
    \new_[8242]_ , \new_[8243]_ , \new_[8247]_ , \new_[8248]_ ,
    \new_[8252]_ , \new_[8253]_ , \new_[8254]_ , \new_[8257]_ ,
    \new_[8261]_ , \new_[8262]_ , \new_[8263]_ , \new_[8267]_ ,
    \new_[8268]_ , \new_[8272]_ , \new_[8273]_ , \new_[8274]_ ,
    \new_[8277]_ , \new_[8281]_ , \new_[8282]_ , \new_[8283]_ ,
    \new_[8287]_ , \new_[8288]_ , \new_[8292]_ , \new_[8293]_ ,
    \new_[8294]_ , \new_[8297]_ , \new_[8301]_ , \new_[8302]_ ,
    \new_[8303]_ , \new_[8307]_ , \new_[8308]_ , \new_[8312]_ ,
    \new_[8313]_ , \new_[8314]_ , \new_[8317]_ , \new_[8321]_ ,
    \new_[8322]_ , \new_[8323]_ , \new_[8327]_ , \new_[8328]_ ,
    \new_[8332]_ , \new_[8333]_ , \new_[8334]_ , \new_[8337]_ ,
    \new_[8341]_ , \new_[8342]_ , \new_[8343]_ , \new_[8347]_ ,
    \new_[8348]_ , \new_[8352]_ , \new_[8353]_ , \new_[8354]_ ,
    \new_[8357]_ , \new_[8361]_ , \new_[8362]_ , \new_[8363]_ ,
    \new_[8367]_ , \new_[8368]_ , \new_[8372]_ , \new_[8373]_ ,
    \new_[8374]_ , \new_[8377]_ , \new_[8381]_ , \new_[8382]_ ,
    \new_[8383]_ , \new_[8387]_ , \new_[8388]_ , \new_[8392]_ ,
    \new_[8393]_ , \new_[8394]_ , \new_[8397]_ , \new_[8401]_ ,
    \new_[8402]_ , \new_[8403]_ , \new_[8407]_ , \new_[8408]_ ,
    \new_[8412]_ , \new_[8413]_ , \new_[8414]_ , \new_[8417]_ ,
    \new_[8421]_ , \new_[8422]_ , \new_[8423]_ , \new_[8427]_ ,
    \new_[8428]_ , \new_[8432]_ , \new_[8433]_ , \new_[8434]_ ,
    \new_[8437]_ , \new_[8441]_ , \new_[8442]_ , \new_[8443]_ ,
    \new_[8447]_ , \new_[8448]_ , \new_[8452]_ , \new_[8453]_ ,
    \new_[8454]_ , \new_[8457]_ , \new_[8461]_ , \new_[8462]_ ,
    \new_[8463]_ , \new_[8467]_ , \new_[8468]_ , \new_[8472]_ ,
    \new_[8473]_ , \new_[8474]_ , \new_[8477]_ , \new_[8481]_ ,
    \new_[8482]_ , \new_[8483]_ , \new_[8487]_ , \new_[8488]_ ,
    \new_[8492]_ , \new_[8493]_ , \new_[8494]_ , \new_[8497]_ ,
    \new_[8501]_ , \new_[8502]_ , \new_[8503]_ , \new_[8507]_ ,
    \new_[8508]_ , \new_[8512]_ , \new_[8513]_ , \new_[8514]_ ,
    \new_[8518]_ , \new_[8519]_ , \new_[8523]_ , \new_[8524]_ ,
    \new_[8525]_ , \new_[8529]_ , \new_[8530]_ , \new_[8534]_ ,
    \new_[8535]_ , \new_[8536]_ , \new_[8540]_ , \new_[8541]_ ,
    \new_[8545]_ , \new_[8546]_ , \new_[8547]_ , \new_[8551]_ ,
    \new_[8552]_ , \new_[8556]_ , \new_[8557]_ , \new_[8558]_ ,
    \new_[8562]_ , \new_[8563]_ , \new_[8567]_ , \new_[8568]_ ,
    \new_[8569]_ , \new_[8573]_ , \new_[8574]_ , \new_[8578]_ ,
    \new_[8579]_ , \new_[8580]_ , \new_[8584]_ , \new_[8585]_ ,
    \new_[8589]_ , \new_[8590]_ , \new_[8591]_ , \new_[8595]_ ,
    \new_[8596]_ , \new_[8600]_ , \new_[8601]_ , \new_[8602]_ ,
    \new_[8606]_ , \new_[8607]_ , \new_[8611]_ , \new_[8612]_ ,
    \new_[8613]_ , \new_[8617]_ , \new_[8618]_ , \new_[8622]_ ,
    \new_[8623]_ , \new_[8624]_ , \new_[8628]_ , \new_[8629]_ ,
    \new_[8633]_ , \new_[8634]_ , \new_[8635]_ , \new_[8639]_ ,
    \new_[8640]_ , \new_[8644]_ , \new_[8645]_ , \new_[8646]_ ,
    \new_[8650]_ , \new_[8651]_ , \new_[8655]_ , \new_[8656]_ ,
    \new_[8657]_ , \new_[8661]_ , \new_[8662]_ , \new_[8666]_ ,
    \new_[8667]_ , \new_[8668]_ , \new_[8672]_ , \new_[8673]_ ,
    \new_[8677]_ , \new_[8678]_ , \new_[8679]_ , \new_[8683]_ ,
    \new_[8684]_ , \new_[8688]_ , \new_[8689]_ , \new_[8690]_ ,
    \new_[8694]_ , \new_[8695]_ , \new_[8699]_ , \new_[8700]_ ,
    \new_[8701]_ , \new_[8705]_ , \new_[8706]_ , \new_[8710]_ ,
    \new_[8711]_ , \new_[8712]_ , \new_[8716]_ , \new_[8717]_ ,
    \new_[8721]_ , \new_[8722]_ , \new_[8723]_ , \new_[8727]_ ,
    \new_[8728]_ , \new_[8732]_ , \new_[8733]_ , \new_[8734]_ ,
    \new_[8738]_ , \new_[8739]_ , \new_[8743]_ , \new_[8744]_ ,
    \new_[8745]_ , \new_[8749]_ , \new_[8750]_ , \new_[8754]_ ,
    \new_[8755]_ , \new_[8756]_ , \new_[8760]_ , \new_[8761]_ ,
    \new_[8765]_ , \new_[8766]_ , \new_[8767]_ , \new_[8771]_ ,
    \new_[8772]_ , \new_[8776]_ , \new_[8777]_ , \new_[8778]_ ,
    \new_[8782]_ , \new_[8783]_ , \new_[8787]_ , \new_[8788]_ ,
    \new_[8789]_ , \new_[8793]_ , \new_[8794]_ , \new_[8798]_ ,
    \new_[8799]_ , \new_[8800]_ , \new_[8804]_ , \new_[8805]_ ,
    \new_[8809]_ , \new_[8810]_ , \new_[8811]_ , \new_[8815]_ ,
    \new_[8816]_ , \new_[8820]_ , \new_[8821]_ , \new_[8822]_ ,
    \new_[8826]_ , \new_[8827]_ , \new_[8831]_ , \new_[8832]_ ,
    \new_[8833]_ , \new_[8837]_ , \new_[8838]_ , \new_[8842]_ ,
    \new_[8843]_ , \new_[8844]_ , \new_[8848]_ , \new_[8849]_ ,
    \new_[8853]_ , \new_[8854]_ , \new_[8855]_ , \new_[8859]_ ,
    \new_[8860]_ , \new_[8864]_ , \new_[8865]_ , \new_[8866]_ ,
    \new_[8870]_ , \new_[8871]_ , \new_[8875]_ , \new_[8876]_ ,
    \new_[8877]_ , \new_[8881]_ , \new_[8882]_ , \new_[8886]_ ,
    \new_[8887]_ , \new_[8888]_ , \new_[8892]_ , \new_[8893]_ ,
    \new_[8897]_ , \new_[8898]_ , \new_[8899]_ , \new_[8903]_ ,
    \new_[8904]_ , \new_[8908]_ , \new_[8909]_ , \new_[8910]_ ,
    \new_[8914]_ , \new_[8915]_ , \new_[8919]_ , \new_[8920]_ ,
    \new_[8921]_ , \new_[8925]_ , \new_[8926]_ , \new_[8930]_ ,
    \new_[8931]_ , \new_[8932]_ , \new_[8936]_ , \new_[8937]_ ,
    \new_[8941]_ , \new_[8942]_ , \new_[8943]_ , \new_[8947]_ ,
    \new_[8948]_ , \new_[8952]_ , \new_[8953]_ , \new_[8954]_ ,
    \new_[8958]_ , \new_[8959]_ , \new_[8963]_ , \new_[8964]_ ,
    \new_[8965]_ , \new_[8969]_ , \new_[8970]_ , \new_[8974]_ ,
    \new_[8975]_ , \new_[8976]_ , \new_[8980]_ , \new_[8981]_ ,
    \new_[8985]_ , \new_[8986]_ , \new_[8987]_ , \new_[8991]_ ,
    \new_[8992]_ , \new_[8996]_ , \new_[8997]_ , \new_[8998]_ ,
    \new_[9002]_ , \new_[9003]_ , \new_[9007]_ , \new_[9008]_ ,
    \new_[9009]_ , \new_[9013]_ , \new_[9014]_ , \new_[9018]_ ,
    \new_[9019]_ , \new_[9020]_ , \new_[9024]_ , \new_[9025]_ ,
    \new_[9029]_ , \new_[9030]_ , \new_[9031]_ , \new_[9035]_ ,
    \new_[9036]_ , \new_[9040]_ , \new_[9041]_ , \new_[9042]_ ,
    \new_[9046]_ , \new_[9047]_ , \new_[9051]_ , \new_[9052]_ ,
    \new_[9053]_ , \new_[9057]_ , \new_[9058]_ , \new_[9062]_ ,
    \new_[9063]_ , \new_[9064]_ , \new_[9068]_ , \new_[9069]_ ,
    \new_[9073]_ , \new_[9074]_ , \new_[9075]_ , \new_[9079]_ ,
    \new_[9080]_ , \new_[9084]_ , \new_[9085]_ , \new_[9086]_ ,
    \new_[9090]_ , \new_[9091]_ , \new_[9095]_ , \new_[9096]_ ,
    \new_[9097]_ , \new_[9101]_ , \new_[9102]_ , \new_[9106]_ ,
    \new_[9107]_ , \new_[9108]_ , \new_[9112]_ , \new_[9113]_ ,
    \new_[9117]_ , \new_[9118]_ , \new_[9119]_ , \new_[9123]_ ,
    \new_[9124]_ , \new_[9128]_ , \new_[9129]_ , \new_[9130]_ ,
    \new_[9134]_ , \new_[9135]_ , \new_[9139]_ , \new_[9140]_ ,
    \new_[9141]_ , \new_[9145]_ , \new_[9146]_ , \new_[9150]_ ,
    \new_[9151]_ , \new_[9152]_ , \new_[9156]_ , \new_[9157]_ ,
    \new_[9161]_ , \new_[9162]_ , \new_[9163]_ , \new_[9167]_ ,
    \new_[9168]_ , \new_[9172]_ , \new_[9173]_ , \new_[9174]_ ,
    \new_[9178]_ , \new_[9179]_ , \new_[9183]_ , \new_[9184]_ ,
    \new_[9185]_ , \new_[9189]_ , \new_[9190]_ , \new_[9194]_ ,
    \new_[9195]_ , \new_[9196]_ , \new_[9200]_ , \new_[9201]_ ,
    \new_[9205]_ , \new_[9206]_ , \new_[9207]_ , \new_[9211]_ ,
    \new_[9212]_ , \new_[9216]_ , \new_[9217]_ , \new_[9218]_ ,
    \new_[9222]_ , \new_[9223]_ , \new_[9227]_ , \new_[9228]_ ,
    \new_[9229]_ , \new_[9233]_ , \new_[9234]_ , \new_[9238]_ ,
    \new_[9239]_ , \new_[9240]_ , \new_[9244]_ , \new_[9245]_ ,
    \new_[9249]_ , \new_[9250]_ , \new_[9251]_ , \new_[9255]_ ,
    \new_[9256]_ , \new_[9260]_ , \new_[9261]_ , \new_[9262]_ ,
    \new_[9266]_ , \new_[9267]_ , \new_[9271]_ , \new_[9272]_ ,
    \new_[9273]_ , \new_[9277]_ , \new_[9278]_ , \new_[9282]_ ,
    \new_[9283]_ , \new_[9284]_ , \new_[9288]_ , \new_[9289]_ ,
    \new_[9293]_ , \new_[9294]_ , \new_[9295]_ , \new_[9299]_ ,
    \new_[9300]_ , \new_[9304]_ , \new_[9305]_ , \new_[9306]_ ,
    \new_[9310]_ , \new_[9311]_ , \new_[9315]_ , \new_[9316]_ ,
    \new_[9317]_ , \new_[9321]_ , \new_[9322]_ , \new_[9326]_ ,
    \new_[9327]_ , \new_[9328]_ , \new_[9332]_ , \new_[9333]_ ,
    \new_[9337]_ , \new_[9338]_ , \new_[9339]_ , \new_[9343]_ ,
    \new_[9344]_ , \new_[9348]_ , \new_[9349]_ , \new_[9350]_ ,
    \new_[9354]_ , \new_[9355]_ , \new_[9359]_ , \new_[9360]_ ,
    \new_[9361]_ , \new_[9365]_ , \new_[9366]_ , \new_[9370]_ ,
    \new_[9371]_ , \new_[9372]_ , \new_[9376]_ , \new_[9377]_ ,
    \new_[9381]_ , \new_[9382]_ , \new_[9383]_ , \new_[9387]_ ,
    \new_[9388]_ , \new_[9392]_ , \new_[9393]_ , \new_[9394]_ ,
    \new_[9398]_ , \new_[9399]_ , \new_[9403]_ , \new_[9404]_ ,
    \new_[9405]_ , \new_[9409]_ , \new_[9410]_ , \new_[9414]_ ,
    \new_[9415]_ , \new_[9416]_ , \new_[9420]_ , \new_[9421]_ ,
    \new_[9425]_ , \new_[9426]_ , \new_[9427]_ , \new_[9431]_ ,
    \new_[9432]_ , \new_[9436]_ , \new_[9437]_ , \new_[9438]_ ,
    \new_[9442]_ , \new_[9443]_ , \new_[9447]_ , \new_[9448]_ ,
    \new_[9449]_ , \new_[9453]_ , \new_[9454]_ , \new_[9458]_ ,
    \new_[9459]_ , \new_[9460]_ , \new_[9464]_ , \new_[9465]_ ,
    \new_[9469]_ , \new_[9470]_ , \new_[9471]_ , \new_[9475]_ ,
    \new_[9476]_ , \new_[9480]_ , \new_[9481]_ , \new_[9482]_ ,
    \new_[9486]_ , \new_[9487]_ , \new_[9491]_ , \new_[9492]_ ,
    \new_[9493]_ , \new_[9497]_ , \new_[9498]_ , \new_[9502]_ ,
    \new_[9503]_ , \new_[9504]_ , \new_[9508]_ , \new_[9509]_ ,
    \new_[9513]_ , \new_[9514]_ , \new_[9515]_ , \new_[9519]_ ,
    \new_[9520]_ , \new_[9524]_ , \new_[9525]_ , \new_[9526]_ ,
    \new_[9530]_ , \new_[9531]_ , \new_[9535]_ , \new_[9536]_ ,
    \new_[9537]_ , \new_[9541]_ , \new_[9542]_ , \new_[9546]_ ,
    \new_[9547]_ , \new_[9548]_ , \new_[9552]_ , \new_[9553]_ ,
    \new_[9557]_ , \new_[9558]_ , \new_[9559]_ , \new_[9563]_ ,
    \new_[9564]_ , \new_[9568]_ , \new_[9569]_ , \new_[9570]_ ,
    \new_[9574]_ , \new_[9575]_ , \new_[9579]_ , \new_[9580]_ ,
    \new_[9581]_ , \new_[9585]_ , \new_[9586]_ , \new_[9590]_ ,
    \new_[9591]_ , \new_[9592]_ , \new_[9596]_ , \new_[9597]_ ,
    \new_[9601]_ , \new_[9602]_ , \new_[9603]_ , \new_[9607]_ ,
    \new_[9608]_ , \new_[9612]_ , \new_[9613]_ , \new_[9614]_ ,
    \new_[9618]_ , \new_[9619]_ , \new_[9623]_ , \new_[9624]_ ,
    \new_[9625]_ , \new_[9629]_ , \new_[9630]_ , \new_[9634]_ ,
    \new_[9635]_ , \new_[9636]_ , \new_[9640]_ , \new_[9641]_ ,
    \new_[9645]_ , \new_[9646]_ , \new_[9647]_ , \new_[9651]_ ,
    \new_[9652]_ , \new_[9656]_ , \new_[9657]_ , \new_[9658]_ ,
    \new_[9662]_ , \new_[9663]_ , \new_[9667]_ , \new_[9668]_ ,
    \new_[9669]_ , \new_[9673]_ , \new_[9674]_ , \new_[9678]_ ,
    \new_[9679]_ , \new_[9680]_ , \new_[9684]_ , \new_[9685]_ ,
    \new_[9689]_ , \new_[9690]_ , \new_[9691]_ , \new_[9695]_ ,
    \new_[9696]_ , \new_[9700]_ , \new_[9701]_ , \new_[9702]_ ,
    \new_[9706]_ , \new_[9707]_ , \new_[9711]_ , \new_[9712]_ ,
    \new_[9713]_ , \new_[9717]_ , \new_[9718]_ , \new_[9722]_ ,
    \new_[9723]_ , \new_[9724]_ , \new_[9728]_ , \new_[9729]_ ,
    \new_[9733]_ , \new_[9734]_ , \new_[9735]_ , \new_[9739]_ ,
    \new_[9740]_ , \new_[9744]_ , \new_[9745]_ , \new_[9746]_ ,
    \new_[9750]_ , \new_[9751]_ , \new_[9755]_ , \new_[9756]_ ,
    \new_[9757]_ , \new_[9761]_ , \new_[9762]_ , \new_[9766]_ ,
    \new_[9767]_ , \new_[9768]_ , \new_[9772]_ , \new_[9773]_ ,
    \new_[9777]_ , \new_[9778]_ , \new_[9779]_ , \new_[9783]_ ,
    \new_[9784]_ , \new_[9788]_ , \new_[9789]_ , \new_[9790]_ ,
    \new_[9794]_ , \new_[9795]_ , \new_[9799]_ , \new_[9800]_ ,
    \new_[9801]_ , \new_[9805]_ , \new_[9806]_ , \new_[9810]_ ,
    \new_[9811]_ , \new_[9812]_ , \new_[9816]_ , \new_[9817]_ ,
    \new_[9821]_ , \new_[9822]_ , \new_[9823]_ , \new_[9827]_ ,
    \new_[9828]_ , \new_[9832]_ , \new_[9833]_ , \new_[9834]_ ,
    \new_[9838]_ , \new_[9839]_ , \new_[9843]_ , \new_[9844]_ ,
    \new_[9845]_ , \new_[9849]_ , \new_[9850]_ , \new_[9854]_ ,
    \new_[9855]_ , \new_[9856]_ , \new_[9860]_ , \new_[9861]_ ,
    \new_[9865]_ , \new_[9866]_ , \new_[9867]_ , \new_[9871]_ ,
    \new_[9872]_ , \new_[9876]_ , \new_[9877]_ , \new_[9878]_ ,
    \new_[9882]_ , \new_[9883]_ , \new_[9887]_ , \new_[9888]_ ,
    \new_[9889]_ , \new_[9893]_ , \new_[9894]_ , \new_[9898]_ ,
    \new_[9899]_ , \new_[9900]_ , \new_[9904]_ , \new_[9905]_ ,
    \new_[9909]_ , \new_[9910]_ , \new_[9911]_ , \new_[9915]_ ,
    \new_[9916]_ , \new_[9920]_ , \new_[9921]_ , \new_[9922]_ ,
    \new_[9926]_ , \new_[9927]_ , \new_[9931]_ , \new_[9932]_ ,
    \new_[9933]_ , \new_[9937]_ , \new_[9938]_ , \new_[9942]_ ,
    \new_[9943]_ , \new_[9944]_ , \new_[9948]_ , \new_[9949]_ ,
    \new_[9953]_ , \new_[9954]_ , \new_[9955]_ , \new_[9959]_ ,
    \new_[9960]_ , \new_[9964]_ , \new_[9965]_ , \new_[9966]_ ,
    \new_[9970]_ , \new_[9971]_ , \new_[9975]_ , \new_[9976]_ ,
    \new_[9977]_ , \new_[9981]_ , \new_[9982]_ , \new_[9986]_ ,
    \new_[9987]_ , \new_[9988]_ , \new_[9992]_ , \new_[9993]_ ,
    \new_[9997]_ , \new_[9998]_ , \new_[9999]_ , \new_[10003]_ ,
    \new_[10004]_ , \new_[10008]_ , \new_[10009]_ , \new_[10010]_ ,
    \new_[10014]_ , \new_[10015]_ , \new_[10019]_ , \new_[10020]_ ,
    \new_[10021]_ , \new_[10025]_ , \new_[10026]_ , \new_[10030]_ ,
    \new_[10031]_ , \new_[10032]_ , \new_[10036]_ , \new_[10037]_ ,
    \new_[10041]_ , \new_[10042]_ , \new_[10043]_ , \new_[10047]_ ,
    \new_[10048]_ , \new_[10052]_ , \new_[10053]_ , \new_[10054]_ ,
    \new_[10058]_ , \new_[10059]_ , \new_[10063]_ , \new_[10064]_ ,
    \new_[10065]_ , \new_[10069]_ , \new_[10070]_ , \new_[10074]_ ,
    \new_[10075]_ , \new_[10076]_ , \new_[10080]_ , \new_[10081]_ ,
    \new_[10085]_ , \new_[10086]_ , \new_[10087]_ , \new_[10091]_ ,
    \new_[10092]_ , \new_[10096]_ , \new_[10097]_ , \new_[10098]_ ,
    \new_[10102]_ , \new_[10103]_ , \new_[10107]_ , \new_[10108]_ ,
    \new_[10109]_ , \new_[10113]_ , \new_[10114]_ , \new_[10118]_ ,
    \new_[10119]_ , \new_[10120]_ , \new_[10124]_ , \new_[10125]_ ,
    \new_[10129]_ , \new_[10130]_ , \new_[10131]_ , \new_[10135]_ ,
    \new_[10136]_ , \new_[10140]_ , \new_[10141]_ , \new_[10142]_ ,
    \new_[10146]_ , \new_[10147]_ , \new_[10151]_ , \new_[10152]_ ,
    \new_[10153]_ , \new_[10157]_ , \new_[10158]_ , \new_[10162]_ ,
    \new_[10163]_ , \new_[10164]_ , \new_[10168]_ , \new_[10169]_ ,
    \new_[10173]_ , \new_[10174]_ , \new_[10175]_ , \new_[10179]_ ,
    \new_[10180]_ , \new_[10184]_ , \new_[10185]_ , \new_[10186]_ ,
    \new_[10190]_ , \new_[10191]_ , \new_[10195]_ , \new_[10196]_ ,
    \new_[10197]_ , \new_[10201]_ , \new_[10202]_ , \new_[10206]_ ,
    \new_[10207]_ , \new_[10208]_ , \new_[10212]_ , \new_[10213]_ ,
    \new_[10217]_ , \new_[10218]_ , \new_[10219]_ , \new_[10223]_ ,
    \new_[10224]_ , \new_[10228]_ , \new_[10229]_ , \new_[10230]_ ,
    \new_[10234]_ , \new_[10235]_ , \new_[10239]_ , \new_[10240]_ ,
    \new_[10241]_ , \new_[10245]_ , \new_[10246]_ , \new_[10250]_ ,
    \new_[10251]_ , \new_[10252]_ , \new_[10256]_ , \new_[10257]_ ,
    \new_[10261]_ , \new_[10262]_ , \new_[10263]_ , \new_[10267]_ ,
    \new_[10268]_ , \new_[10272]_ , \new_[10273]_ , \new_[10274]_ ,
    \new_[10278]_ , \new_[10279]_ , \new_[10283]_ , \new_[10284]_ ,
    \new_[10285]_ , \new_[10289]_ , \new_[10290]_ , \new_[10294]_ ,
    \new_[10295]_ , \new_[10296]_ , \new_[10300]_ , \new_[10301]_ ,
    \new_[10305]_ , \new_[10306]_ , \new_[10307]_ , \new_[10311]_ ,
    \new_[10312]_ , \new_[10316]_ , \new_[10317]_ , \new_[10318]_ ,
    \new_[10322]_ , \new_[10323]_ , \new_[10327]_ , \new_[10328]_ ,
    \new_[10329]_ , \new_[10333]_ , \new_[10334]_ , \new_[10338]_ ,
    \new_[10339]_ , \new_[10340]_ , \new_[10344]_ , \new_[10345]_ ,
    \new_[10349]_ , \new_[10350]_ , \new_[10351]_ , \new_[10355]_ ,
    \new_[10356]_ , \new_[10360]_ , \new_[10361]_ , \new_[10362]_ ,
    \new_[10366]_ , \new_[10367]_ , \new_[10371]_ , \new_[10372]_ ,
    \new_[10373]_ , \new_[10377]_ , \new_[10378]_ , \new_[10382]_ ,
    \new_[10383]_ , \new_[10384]_ , \new_[10388]_ , \new_[10389]_ ,
    \new_[10393]_ , \new_[10394]_ , \new_[10395]_ , \new_[10399]_ ,
    \new_[10400]_ , \new_[10404]_ , \new_[10405]_ , \new_[10406]_ ,
    \new_[10410]_ , \new_[10411]_ , \new_[10415]_ , \new_[10416]_ ,
    \new_[10417]_ , \new_[10421]_ , \new_[10422]_ , \new_[10426]_ ,
    \new_[10427]_ , \new_[10428]_ , \new_[10432]_ , \new_[10433]_ ,
    \new_[10437]_ , \new_[10438]_ , \new_[10439]_ , \new_[10443]_ ,
    \new_[10444]_ , \new_[10448]_ , \new_[10449]_ , \new_[10450]_ ,
    \new_[10454]_ , \new_[10455]_ , \new_[10459]_ , \new_[10460]_ ,
    \new_[10461]_ , \new_[10465]_ , \new_[10466]_ , \new_[10470]_ ,
    \new_[10471]_ , \new_[10472]_ , \new_[10476]_ , \new_[10477]_ ,
    \new_[10481]_ , \new_[10482]_ , \new_[10483]_ , \new_[10487]_ ,
    \new_[10488]_ , \new_[10492]_ , \new_[10493]_ , \new_[10494]_ ,
    \new_[10498]_ , \new_[10499]_ , \new_[10503]_ , \new_[10504]_ ,
    \new_[10505]_ , \new_[10509]_ , \new_[10510]_ , \new_[10514]_ ,
    \new_[10515]_ , \new_[10516]_ , \new_[10520]_ , \new_[10521]_ ,
    \new_[10525]_ , \new_[10526]_ , \new_[10527]_ , \new_[10531]_ ,
    \new_[10532]_ , \new_[10536]_ , \new_[10537]_ , \new_[10538]_ ,
    \new_[10542]_ , \new_[10543]_ , \new_[10547]_ , \new_[10548]_ ,
    \new_[10549]_ , \new_[10553]_ , \new_[10554]_ , \new_[10558]_ ,
    \new_[10559]_ , \new_[10560]_ , \new_[10564]_ , \new_[10565]_ ,
    \new_[10569]_ , \new_[10570]_ , \new_[10571]_ , \new_[10575]_ ,
    \new_[10576]_ , \new_[10580]_ , \new_[10581]_ , \new_[10582]_ ,
    \new_[10586]_ , \new_[10587]_ , \new_[10591]_ , \new_[10592]_ ,
    \new_[10593]_ , \new_[10597]_ , \new_[10598]_ , \new_[10602]_ ,
    \new_[10603]_ , \new_[10604]_ , \new_[10608]_ , \new_[10609]_ ,
    \new_[10613]_ , \new_[10614]_ , \new_[10615]_ , \new_[10619]_ ,
    \new_[10620]_ , \new_[10624]_ , \new_[10625]_ , \new_[10626]_ ,
    \new_[10630]_ , \new_[10631]_ , \new_[10635]_ , \new_[10636]_ ,
    \new_[10637]_ , \new_[10641]_ , \new_[10642]_ , \new_[10646]_ ,
    \new_[10647]_ , \new_[10648]_ , \new_[10652]_ , \new_[10653]_ ,
    \new_[10657]_ , \new_[10658]_ , \new_[10659]_ , \new_[10663]_ ,
    \new_[10664]_ , \new_[10668]_ , \new_[10669]_ , \new_[10670]_ ,
    \new_[10674]_ , \new_[10675]_ , \new_[10679]_ , \new_[10680]_ ,
    \new_[10681]_ , \new_[10685]_ , \new_[10686]_ , \new_[10690]_ ,
    \new_[10691]_ , \new_[10692]_ , \new_[10696]_ , \new_[10697]_ ,
    \new_[10701]_ , \new_[10702]_ , \new_[10703]_ , \new_[10707]_ ,
    \new_[10708]_ , \new_[10712]_ , \new_[10713]_ , \new_[10714]_ ,
    \new_[10718]_ , \new_[10719]_ , \new_[10723]_ , \new_[10724]_ ,
    \new_[10725]_ , \new_[10729]_ , \new_[10730]_ , \new_[10734]_ ,
    \new_[10735]_ , \new_[10736]_ , \new_[10740]_ , \new_[10741]_ ,
    \new_[10745]_ , \new_[10746]_ , \new_[10747]_ , \new_[10751]_ ,
    \new_[10752]_ , \new_[10756]_ , \new_[10757]_ , \new_[10758]_ ,
    \new_[10762]_ , \new_[10763]_ , \new_[10767]_ , \new_[10768]_ ,
    \new_[10769]_ , \new_[10773]_ , \new_[10774]_ , \new_[10778]_ ,
    \new_[10779]_ , \new_[10780]_ , \new_[10784]_ , \new_[10785]_ ,
    \new_[10789]_ , \new_[10790]_ , \new_[10791]_ , \new_[10795]_ ,
    \new_[10796]_ , \new_[10800]_ , \new_[10801]_ , \new_[10802]_ ,
    \new_[10806]_ , \new_[10807]_ , \new_[10811]_ , \new_[10812]_ ,
    \new_[10813]_ , \new_[10817]_ , \new_[10818]_ , \new_[10822]_ ,
    \new_[10823]_ , \new_[10824]_ , \new_[10828]_ , \new_[10829]_ ,
    \new_[10833]_ , \new_[10834]_ , \new_[10835]_ , \new_[10839]_ ,
    \new_[10840]_ , \new_[10844]_ , \new_[10845]_ , \new_[10846]_ ,
    \new_[10850]_ , \new_[10851]_ , \new_[10855]_ , \new_[10856]_ ,
    \new_[10857]_ , \new_[10861]_ , \new_[10862]_ , \new_[10866]_ ,
    \new_[10867]_ , \new_[10868]_ , \new_[10872]_ , \new_[10873]_ ,
    \new_[10877]_ , \new_[10878]_ , \new_[10879]_ , \new_[10883]_ ,
    \new_[10884]_ , \new_[10888]_ , \new_[10889]_ , \new_[10890]_ ,
    \new_[10894]_ , \new_[10895]_ , \new_[10899]_ , \new_[10900]_ ,
    \new_[10901]_ , \new_[10905]_ , \new_[10906]_ , \new_[10910]_ ,
    \new_[10911]_ , \new_[10912]_ , \new_[10916]_ , \new_[10917]_ ,
    \new_[10921]_ , \new_[10922]_ , \new_[10923]_ , \new_[10927]_ ,
    \new_[10928]_ , \new_[10932]_ , \new_[10933]_ , \new_[10934]_ ,
    \new_[10938]_ , \new_[10939]_ , \new_[10943]_ , \new_[10944]_ ,
    \new_[10945]_ , \new_[10949]_ , \new_[10950]_ , \new_[10954]_ ,
    \new_[10955]_ , \new_[10956]_ , \new_[10960]_ , \new_[10961]_ ,
    \new_[10965]_ , \new_[10966]_ , \new_[10967]_ , \new_[10971]_ ,
    \new_[10972]_ , \new_[10976]_ , \new_[10977]_ , \new_[10978]_ ,
    \new_[10982]_ , \new_[10983]_ , \new_[10987]_ , \new_[10988]_ ,
    \new_[10989]_ , \new_[10993]_ , \new_[10994]_ , \new_[10998]_ ,
    \new_[10999]_ , \new_[11000]_ , \new_[11004]_ , \new_[11005]_ ,
    \new_[11009]_ , \new_[11010]_ , \new_[11011]_ , \new_[11015]_ ,
    \new_[11016]_ , \new_[11020]_ , \new_[11021]_ , \new_[11022]_ ,
    \new_[11026]_ , \new_[11027]_ , \new_[11031]_ , \new_[11032]_ ,
    \new_[11033]_ , \new_[11037]_ , \new_[11038]_ , \new_[11042]_ ,
    \new_[11043]_ , \new_[11044]_ , \new_[11048]_ , \new_[11049]_ ,
    \new_[11053]_ , \new_[11054]_ , \new_[11055]_ , \new_[11059]_ ,
    \new_[11060]_ , \new_[11064]_ , \new_[11065]_ , \new_[11066]_ ,
    \new_[11070]_ , \new_[11071]_ , \new_[11075]_ , \new_[11076]_ ,
    \new_[11077]_ , \new_[11081]_ , \new_[11082]_ , \new_[11086]_ ,
    \new_[11087]_ , \new_[11088]_ , \new_[11092]_ , \new_[11093]_ ,
    \new_[11097]_ , \new_[11098]_ , \new_[11099]_ , \new_[11103]_ ,
    \new_[11104]_ , \new_[11108]_ , \new_[11109]_ , \new_[11110]_ ,
    \new_[11114]_ , \new_[11115]_ , \new_[11119]_ , \new_[11120]_ ,
    \new_[11121]_ , \new_[11125]_ , \new_[11126]_ , \new_[11130]_ ,
    \new_[11131]_ , \new_[11132]_ , \new_[11136]_ , \new_[11137]_ ,
    \new_[11141]_ , \new_[11142]_ , \new_[11143]_ , \new_[11147]_ ,
    \new_[11148]_ , \new_[11152]_ , \new_[11153]_ , \new_[11154]_ ,
    \new_[11158]_ , \new_[11159]_ , \new_[11163]_ , \new_[11164]_ ,
    \new_[11165]_ , \new_[11169]_ , \new_[11170]_ , \new_[11174]_ ,
    \new_[11175]_ , \new_[11176]_ , \new_[11180]_ , \new_[11181]_ ,
    \new_[11185]_ , \new_[11186]_ , \new_[11187]_ , \new_[11191]_ ,
    \new_[11192]_ , \new_[11196]_ , \new_[11197]_ , \new_[11198]_ ,
    \new_[11202]_ , \new_[11203]_ , \new_[11207]_ , \new_[11208]_ ,
    \new_[11209]_ , \new_[11213]_ , \new_[11214]_ , \new_[11218]_ ,
    \new_[11219]_ , \new_[11220]_ , \new_[11224]_ , \new_[11225]_ ,
    \new_[11229]_ , \new_[11230]_ , \new_[11231]_ , \new_[11235]_ ,
    \new_[11236]_ , \new_[11240]_ , \new_[11241]_ , \new_[11242]_ ,
    \new_[11246]_ , \new_[11247]_ , \new_[11251]_ , \new_[11252]_ ,
    \new_[11253]_ , \new_[11257]_ , \new_[11258]_ , \new_[11262]_ ,
    \new_[11263]_ , \new_[11264]_ , \new_[11268]_ , \new_[11269]_ ,
    \new_[11273]_ , \new_[11274]_ , \new_[11275]_ , \new_[11279]_ ,
    \new_[11280]_ , \new_[11284]_ , \new_[11285]_ , \new_[11286]_ ,
    \new_[11290]_ , \new_[11291]_ , \new_[11295]_ , \new_[11296]_ ,
    \new_[11297]_ , \new_[11301]_ , \new_[11302]_ , \new_[11306]_ ,
    \new_[11307]_ , \new_[11308]_ , \new_[11312]_ , \new_[11313]_ ,
    \new_[11317]_ , \new_[11318]_ , \new_[11319]_ , \new_[11323]_ ,
    \new_[11324]_ , \new_[11328]_ , \new_[11329]_ , \new_[11330]_ ,
    \new_[11334]_ , \new_[11335]_ , \new_[11339]_ , \new_[11340]_ ,
    \new_[11341]_ , \new_[11345]_ , \new_[11346]_ , \new_[11350]_ ,
    \new_[11351]_ , \new_[11352]_ , \new_[11356]_ , \new_[11357]_ ,
    \new_[11361]_ , \new_[11362]_ , \new_[11363]_ , \new_[11367]_ ,
    \new_[11368]_ , \new_[11372]_ , \new_[11373]_ , \new_[11374]_ ,
    \new_[11378]_ , \new_[11379]_ , \new_[11383]_ , \new_[11384]_ ,
    \new_[11385]_ , \new_[11389]_ , \new_[11390]_ , \new_[11394]_ ,
    \new_[11395]_ , \new_[11396]_ , \new_[11400]_ , \new_[11401]_ ,
    \new_[11405]_ , \new_[11406]_ , \new_[11407]_ , \new_[11411]_ ,
    \new_[11412]_ , \new_[11416]_ , \new_[11417]_ , \new_[11418]_ ,
    \new_[11422]_ , \new_[11423]_ , \new_[11427]_ , \new_[11428]_ ,
    \new_[11429]_ , \new_[11433]_ , \new_[11434]_ , \new_[11438]_ ,
    \new_[11439]_ , \new_[11440]_ , \new_[11444]_ , \new_[11445]_ ,
    \new_[11449]_ , \new_[11450]_ , \new_[11451]_ , \new_[11455]_ ,
    \new_[11456]_ , \new_[11460]_ , \new_[11461]_ , \new_[11462]_ ,
    \new_[11466]_ , \new_[11467]_ , \new_[11471]_ , \new_[11472]_ ,
    \new_[11473]_ , \new_[11477]_ , \new_[11478]_ , \new_[11482]_ ,
    \new_[11483]_ , \new_[11484]_ , \new_[11488]_ , \new_[11489]_ ,
    \new_[11493]_ , \new_[11494]_ , \new_[11495]_ , \new_[11499]_ ,
    \new_[11500]_ , \new_[11504]_ , \new_[11505]_ , \new_[11506]_ ,
    \new_[11510]_ , \new_[11511]_ , \new_[11515]_ , \new_[11516]_ ,
    \new_[11517]_ , \new_[11521]_ , \new_[11522]_ , \new_[11526]_ ,
    \new_[11527]_ , \new_[11528]_ , \new_[11532]_ , \new_[11533]_ ,
    \new_[11537]_ , \new_[11538]_ , \new_[11539]_ , \new_[11543]_ ,
    \new_[11544]_ , \new_[11548]_ , \new_[11549]_ , \new_[11550]_ ,
    \new_[11554]_ , \new_[11555]_ , \new_[11559]_ , \new_[11560]_ ,
    \new_[11561]_ , \new_[11565]_ , \new_[11566]_ , \new_[11570]_ ,
    \new_[11571]_ , \new_[11572]_ , \new_[11576]_ , \new_[11577]_ ,
    \new_[11581]_ , \new_[11582]_ , \new_[11583]_ , \new_[11587]_ ,
    \new_[11588]_ , \new_[11592]_ , \new_[11593]_ , \new_[11594]_ ,
    \new_[11598]_ , \new_[11599]_ , \new_[11603]_ , \new_[11604]_ ,
    \new_[11605]_ , \new_[11609]_ , \new_[11610]_ , \new_[11614]_ ,
    \new_[11615]_ , \new_[11616]_ , \new_[11620]_ , \new_[11621]_ ,
    \new_[11625]_ , \new_[11626]_ , \new_[11627]_ , \new_[11631]_ ,
    \new_[11632]_ , \new_[11636]_ , \new_[11637]_ , \new_[11638]_ ,
    \new_[11642]_ , \new_[11643]_ , \new_[11647]_ , \new_[11648]_ ,
    \new_[11649]_ , \new_[11653]_ , \new_[11654]_ , \new_[11658]_ ,
    \new_[11659]_ , \new_[11660]_ , \new_[11664]_ , \new_[11665]_ ,
    \new_[11669]_ , \new_[11670]_ , \new_[11671]_ , \new_[11675]_ ,
    \new_[11676]_ , \new_[11680]_ , \new_[11681]_ , \new_[11682]_ ,
    \new_[11686]_ , \new_[11687]_ , \new_[11691]_ , \new_[11692]_ ,
    \new_[11693]_ , \new_[11697]_ , \new_[11698]_ , \new_[11702]_ ,
    \new_[11703]_ , \new_[11704]_ , \new_[11708]_ , \new_[11709]_ ,
    \new_[11713]_ , \new_[11714]_ , \new_[11715]_ , \new_[11719]_ ,
    \new_[11720]_ , \new_[11724]_ , \new_[11725]_ , \new_[11726]_ ,
    \new_[11730]_ , \new_[11731]_ , \new_[11735]_ , \new_[11736]_ ,
    \new_[11737]_ , \new_[11741]_ , \new_[11742]_ , \new_[11746]_ ,
    \new_[11747]_ , \new_[11748]_ , \new_[11752]_ , \new_[11753]_ ,
    \new_[11757]_ , \new_[11758]_ , \new_[11759]_ , \new_[11763]_ ,
    \new_[11764]_ , \new_[11768]_ , \new_[11769]_ , \new_[11770]_ ,
    \new_[11774]_ , \new_[11775]_ , \new_[11779]_ , \new_[11780]_ ,
    \new_[11781]_ , \new_[11785]_ , \new_[11786]_ , \new_[11790]_ ,
    \new_[11791]_ , \new_[11792]_ , \new_[11796]_ , \new_[11797]_ ,
    \new_[11801]_ , \new_[11802]_ , \new_[11803]_ , \new_[11807]_ ,
    \new_[11808]_ , \new_[11812]_ , \new_[11813]_ , \new_[11814]_ ,
    \new_[11818]_ , \new_[11819]_ , \new_[11823]_ , \new_[11824]_ ,
    \new_[11825]_ , \new_[11829]_ , \new_[11830]_ , \new_[11834]_ ,
    \new_[11835]_ , \new_[11836]_ , \new_[11840]_ , \new_[11841]_ ,
    \new_[11845]_ , \new_[11846]_ , \new_[11847]_ , \new_[11851]_ ,
    \new_[11852]_ , \new_[11856]_ , \new_[11857]_ , \new_[11858]_ ,
    \new_[11862]_ , \new_[11863]_ , \new_[11867]_ , \new_[11868]_ ,
    \new_[11869]_ , \new_[11873]_ , \new_[11874]_ , \new_[11878]_ ,
    \new_[11879]_ , \new_[11880]_ , \new_[11884]_ , \new_[11885]_ ,
    \new_[11889]_ , \new_[11890]_ , \new_[11891]_ , \new_[11895]_ ,
    \new_[11896]_ , \new_[11900]_ , \new_[11901]_ , \new_[11902]_ ,
    \new_[11906]_ , \new_[11907]_ , \new_[11911]_ , \new_[11912]_ ,
    \new_[11913]_ , \new_[11917]_ , \new_[11918]_ , \new_[11922]_ ,
    \new_[11923]_ , \new_[11924]_ , \new_[11928]_ , \new_[11929]_ ,
    \new_[11933]_ , \new_[11934]_ , \new_[11935]_ , \new_[11939]_ ,
    \new_[11940]_ , \new_[11944]_ , \new_[11945]_ , \new_[11946]_ ,
    \new_[11950]_ , \new_[11951]_ , \new_[11955]_ , \new_[11956]_ ,
    \new_[11957]_ , \new_[11961]_ , \new_[11962]_ , \new_[11966]_ ,
    \new_[11967]_ , \new_[11968]_ , \new_[11972]_ , \new_[11973]_ ,
    \new_[11977]_ , \new_[11978]_ , \new_[11979]_ , \new_[11983]_ ,
    \new_[11984]_ , \new_[11988]_ , \new_[11989]_ , \new_[11990]_ ,
    \new_[11994]_ , \new_[11995]_ , \new_[11999]_ , \new_[12000]_ ,
    \new_[12001]_ , \new_[12005]_ , \new_[12006]_ , \new_[12010]_ ,
    \new_[12011]_ , \new_[12012]_ , \new_[12016]_ , \new_[12017]_ ,
    \new_[12021]_ , \new_[12022]_ , \new_[12023]_ , \new_[12027]_ ,
    \new_[12028]_ , \new_[12032]_ , \new_[12033]_ , \new_[12034]_ ,
    \new_[12038]_ , \new_[12039]_ , \new_[12043]_ , \new_[12044]_ ,
    \new_[12045]_ , \new_[12049]_ , \new_[12050]_ , \new_[12054]_ ,
    \new_[12055]_ , \new_[12056]_ , \new_[12060]_ , \new_[12061]_ ,
    \new_[12065]_ , \new_[12066]_ , \new_[12067]_ , \new_[12071]_ ,
    \new_[12072]_ , \new_[12076]_ , \new_[12077]_ , \new_[12078]_ ,
    \new_[12082]_ , \new_[12083]_ , \new_[12087]_ , \new_[12088]_ ,
    \new_[12089]_ , \new_[12093]_ , \new_[12094]_ , \new_[12098]_ ,
    \new_[12099]_ , \new_[12100]_ , \new_[12104]_ , \new_[12105]_ ,
    \new_[12109]_ , \new_[12110]_ , \new_[12111]_ , \new_[12115]_ ,
    \new_[12116]_ , \new_[12120]_ , \new_[12121]_ , \new_[12122]_ ,
    \new_[12126]_ , \new_[12127]_ , \new_[12131]_ , \new_[12132]_ ,
    \new_[12133]_ , \new_[12137]_ , \new_[12138]_ , \new_[12142]_ ,
    \new_[12143]_ , \new_[12144]_ , \new_[12148]_ , \new_[12149]_ ,
    \new_[12153]_ , \new_[12154]_ , \new_[12155]_ , \new_[12159]_ ,
    \new_[12160]_ , \new_[12164]_ , \new_[12165]_ , \new_[12166]_ ,
    \new_[12170]_ , \new_[12171]_ , \new_[12175]_ , \new_[12176]_ ,
    \new_[12177]_ , \new_[12181]_ , \new_[12182]_ , \new_[12186]_ ,
    \new_[12187]_ , \new_[12188]_ , \new_[12192]_ , \new_[12193]_ ,
    \new_[12197]_ , \new_[12198]_ , \new_[12199]_ , \new_[12203]_ ,
    \new_[12204]_ , \new_[12208]_ , \new_[12209]_ , \new_[12210]_ ,
    \new_[12214]_ , \new_[12215]_ , \new_[12219]_ , \new_[12220]_ ,
    \new_[12221]_ , \new_[12225]_ , \new_[12226]_ , \new_[12230]_ ,
    \new_[12231]_ , \new_[12232]_ , \new_[12236]_ , \new_[12237]_ ,
    \new_[12241]_ , \new_[12242]_ , \new_[12243]_ , \new_[12247]_ ,
    \new_[12248]_ , \new_[12252]_ , \new_[12253]_ , \new_[12254]_ ,
    \new_[12258]_ , \new_[12259]_ , \new_[12263]_ , \new_[12264]_ ,
    \new_[12265]_ , \new_[12269]_ , \new_[12270]_ , \new_[12274]_ ,
    \new_[12275]_ , \new_[12276]_ , \new_[12280]_ , \new_[12281]_ ,
    \new_[12285]_ , \new_[12286]_ , \new_[12287]_ , \new_[12291]_ ,
    \new_[12292]_ , \new_[12296]_ , \new_[12297]_ , \new_[12298]_ ,
    \new_[12302]_ , \new_[12303]_ , \new_[12307]_ , \new_[12308]_ ,
    \new_[12309]_ , \new_[12313]_ , \new_[12314]_ , \new_[12318]_ ,
    \new_[12319]_ , \new_[12320]_ , \new_[12324]_ , \new_[12325]_ ,
    \new_[12329]_ , \new_[12330]_ , \new_[12331]_ , \new_[12335]_ ,
    \new_[12336]_ , \new_[12340]_ , \new_[12341]_ , \new_[12342]_ ,
    \new_[12346]_ , \new_[12347]_ , \new_[12351]_ , \new_[12352]_ ,
    \new_[12353]_ , \new_[12357]_ , \new_[12358]_ , \new_[12362]_ ,
    \new_[12363]_ , \new_[12364]_ , \new_[12368]_ , \new_[12369]_ ,
    \new_[12373]_ , \new_[12374]_ , \new_[12375]_ , \new_[12379]_ ,
    \new_[12380]_ , \new_[12384]_ , \new_[12385]_ , \new_[12386]_ ,
    \new_[12390]_ , \new_[12391]_ , \new_[12395]_ , \new_[12396]_ ,
    \new_[12397]_ , \new_[12401]_ , \new_[12402]_ , \new_[12406]_ ,
    \new_[12407]_ , \new_[12408]_ , \new_[12412]_ , \new_[12413]_ ,
    \new_[12417]_ , \new_[12418]_ , \new_[12419]_ , \new_[12423]_ ,
    \new_[12424]_ , \new_[12428]_ , \new_[12429]_ , \new_[12430]_ ,
    \new_[12434]_ , \new_[12435]_ , \new_[12439]_ , \new_[12440]_ ,
    \new_[12441]_ , \new_[12445]_ , \new_[12446]_ , \new_[12450]_ ,
    \new_[12451]_ , \new_[12452]_ , \new_[12456]_ , \new_[12457]_ ,
    \new_[12461]_ , \new_[12462]_ , \new_[12463]_ , \new_[12467]_ ,
    \new_[12468]_ , \new_[12472]_ , \new_[12473]_ , \new_[12474]_ ,
    \new_[12478]_ , \new_[12479]_ , \new_[12483]_ , \new_[12484]_ ,
    \new_[12485]_ , \new_[12489]_ , \new_[12490]_ , \new_[12494]_ ,
    \new_[12495]_ , \new_[12496]_ , \new_[12500]_ , \new_[12501]_ ,
    \new_[12505]_ , \new_[12506]_ , \new_[12507]_ , \new_[12511]_ ,
    \new_[12512]_ , \new_[12516]_ , \new_[12517]_ , \new_[12518]_ ,
    \new_[12522]_ , \new_[12523]_ , \new_[12527]_ , \new_[12528]_ ,
    \new_[12529]_ , \new_[12533]_ , \new_[12534]_ , \new_[12538]_ ,
    \new_[12539]_ , \new_[12540]_ , \new_[12544]_ , \new_[12545]_ ,
    \new_[12549]_ , \new_[12550]_ , \new_[12551]_ , \new_[12555]_ ,
    \new_[12556]_ , \new_[12560]_ , \new_[12561]_ , \new_[12562]_ ,
    \new_[12566]_ , \new_[12567]_ , \new_[12571]_ , \new_[12572]_ ,
    \new_[12573]_ , \new_[12577]_ , \new_[12578]_ , \new_[12582]_ ,
    \new_[12583]_ , \new_[12584]_ , \new_[12588]_ , \new_[12589]_ ,
    \new_[12593]_ , \new_[12594]_ , \new_[12595]_ , \new_[12599]_ ,
    \new_[12600]_ , \new_[12604]_ , \new_[12605]_ , \new_[12606]_ ,
    \new_[12610]_ , \new_[12611]_ , \new_[12615]_ , \new_[12616]_ ,
    \new_[12617]_ , \new_[12621]_ , \new_[12622]_ , \new_[12626]_ ,
    \new_[12627]_ , \new_[12628]_ , \new_[12632]_ , \new_[12633]_ ,
    \new_[12637]_ , \new_[12638]_ , \new_[12639]_ , \new_[12643]_ ,
    \new_[12644]_ , \new_[12648]_ , \new_[12649]_ , \new_[12650]_ ,
    \new_[12654]_ , \new_[12655]_ , \new_[12659]_ , \new_[12660]_ ,
    \new_[12661]_ , \new_[12665]_ , \new_[12666]_ , \new_[12670]_ ,
    \new_[12671]_ , \new_[12672]_ , \new_[12676]_ , \new_[12677]_ ,
    \new_[12681]_ , \new_[12682]_ , \new_[12683]_ , \new_[12687]_ ,
    \new_[12688]_ , \new_[12692]_ , \new_[12693]_ , \new_[12694]_ ,
    \new_[12698]_ , \new_[12699]_ , \new_[12703]_ , \new_[12704]_ ,
    \new_[12705]_ , \new_[12709]_ , \new_[12710]_ , \new_[12714]_ ,
    \new_[12715]_ , \new_[12716]_ , \new_[12720]_ , \new_[12721]_ ,
    \new_[12725]_ , \new_[12726]_ , \new_[12727]_ , \new_[12731]_ ,
    \new_[12732]_ , \new_[12736]_ , \new_[12737]_ , \new_[12738]_ ,
    \new_[12742]_ , \new_[12743]_ , \new_[12747]_ , \new_[12748]_ ,
    \new_[12749]_ , \new_[12753]_ , \new_[12754]_ , \new_[12758]_ ,
    \new_[12759]_ , \new_[12760]_ , \new_[12764]_ , \new_[12765]_ ,
    \new_[12769]_ , \new_[12770]_ , \new_[12771]_ , \new_[12775]_ ,
    \new_[12776]_ , \new_[12780]_ , \new_[12781]_ , \new_[12782]_ ,
    \new_[12786]_ , \new_[12787]_ , \new_[12791]_ , \new_[12792]_ ,
    \new_[12793]_ , \new_[12797]_ , \new_[12798]_ , \new_[12802]_ ,
    \new_[12803]_ , \new_[12804]_ , \new_[12808]_ , \new_[12809]_ ,
    \new_[12813]_ , \new_[12814]_ , \new_[12815]_ , \new_[12819]_ ,
    \new_[12820]_ , \new_[12824]_ , \new_[12825]_ , \new_[12826]_ ,
    \new_[12830]_ , \new_[12831]_ , \new_[12835]_ , \new_[12836]_ ,
    \new_[12837]_ , \new_[12841]_ , \new_[12842]_ , \new_[12846]_ ,
    \new_[12847]_ , \new_[12848]_ , \new_[12852]_ , \new_[12853]_ ,
    \new_[12857]_ , \new_[12858]_ , \new_[12859]_ , \new_[12863]_ ,
    \new_[12864]_ , \new_[12868]_ , \new_[12869]_ , \new_[12870]_ ,
    \new_[12874]_ , \new_[12875]_ , \new_[12879]_ , \new_[12880]_ ,
    \new_[12881]_ , \new_[12885]_ , \new_[12886]_ , \new_[12890]_ ,
    \new_[12891]_ , \new_[12892]_ , \new_[12896]_ , \new_[12897]_ ,
    \new_[12901]_ , \new_[12902]_ , \new_[12903]_ , \new_[12907]_ ,
    \new_[12908]_ , \new_[12912]_ , \new_[12913]_ , \new_[12914]_ ,
    \new_[12918]_ , \new_[12919]_ , \new_[12923]_ , \new_[12924]_ ,
    \new_[12925]_ , \new_[12929]_ , \new_[12930]_ , \new_[12934]_ ,
    \new_[12935]_ , \new_[12936]_ , \new_[12940]_ , \new_[12941]_ ,
    \new_[12945]_ , \new_[12946]_ , \new_[12947]_ , \new_[12951]_ ,
    \new_[12952]_ , \new_[12956]_ , \new_[12957]_ , \new_[12958]_ ,
    \new_[12962]_ , \new_[12963]_ , \new_[12967]_ , \new_[12968]_ ,
    \new_[12969]_ , \new_[12973]_ , \new_[12974]_ , \new_[12978]_ ,
    \new_[12979]_ , \new_[12980]_ , \new_[12984]_ , \new_[12985]_ ,
    \new_[12989]_ , \new_[12990]_ , \new_[12991]_ , \new_[12995]_ ,
    \new_[12996]_ , \new_[13000]_ , \new_[13001]_ , \new_[13002]_ ,
    \new_[13006]_ , \new_[13007]_ , \new_[13011]_ , \new_[13012]_ ,
    \new_[13013]_ , \new_[13017]_ , \new_[13018]_ , \new_[13022]_ ,
    \new_[13023]_ , \new_[13024]_ , \new_[13028]_ , \new_[13029]_ ,
    \new_[13033]_ , \new_[13034]_ , \new_[13035]_ , \new_[13039]_ ,
    \new_[13040]_ , \new_[13044]_ , \new_[13045]_ , \new_[13046]_ ,
    \new_[13050]_ , \new_[13051]_ , \new_[13055]_ , \new_[13056]_ ,
    \new_[13057]_ , \new_[13061]_ , \new_[13062]_ , \new_[13066]_ ,
    \new_[13067]_ , \new_[13068]_ , \new_[13072]_ , \new_[13073]_ ,
    \new_[13077]_ , \new_[13078]_ , \new_[13079]_ , \new_[13083]_ ,
    \new_[13084]_ , \new_[13088]_ , \new_[13089]_ , \new_[13090]_ ,
    \new_[13094]_ , \new_[13095]_ , \new_[13099]_ , \new_[13100]_ ,
    \new_[13101]_ , \new_[13105]_ , \new_[13106]_ , \new_[13110]_ ,
    \new_[13111]_ , \new_[13112]_ , \new_[13116]_ , \new_[13117]_ ,
    \new_[13121]_ , \new_[13122]_ , \new_[13123]_ , \new_[13127]_ ,
    \new_[13128]_ , \new_[13132]_ , \new_[13133]_ , \new_[13134]_ ,
    \new_[13138]_ , \new_[13139]_ , \new_[13143]_ , \new_[13144]_ ,
    \new_[13145]_ , \new_[13149]_ , \new_[13150]_ , \new_[13154]_ ,
    \new_[13155]_ , \new_[13156]_ , \new_[13160]_ , \new_[13161]_ ,
    \new_[13165]_ , \new_[13166]_ , \new_[13167]_ , \new_[13171]_ ,
    \new_[13172]_ , \new_[13176]_ , \new_[13177]_ , \new_[13178]_ ,
    \new_[13182]_ , \new_[13183]_ , \new_[13187]_ , \new_[13188]_ ,
    \new_[13189]_ , \new_[13193]_ , \new_[13194]_ , \new_[13198]_ ,
    \new_[13199]_ , \new_[13200]_ , \new_[13204]_ , \new_[13205]_ ,
    \new_[13209]_ , \new_[13210]_ , \new_[13211]_ , \new_[13215]_ ,
    \new_[13216]_ , \new_[13220]_ , \new_[13221]_ , \new_[13222]_ ,
    \new_[13226]_ , \new_[13227]_ , \new_[13231]_ , \new_[13232]_ ,
    \new_[13233]_ , \new_[13237]_ , \new_[13238]_ , \new_[13242]_ ,
    \new_[13243]_ , \new_[13244]_ , \new_[13248]_ , \new_[13249]_ ,
    \new_[13253]_ , \new_[13254]_ , \new_[13255]_ , \new_[13259]_ ,
    \new_[13260]_ , \new_[13264]_ , \new_[13265]_ , \new_[13266]_ ,
    \new_[13270]_ , \new_[13271]_ , \new_[13275]_ , \new_[13276]_ ,
    \new_[13277]_ , \new_[13281]_ , \new_[13282]_ , \new_[13286]_ ,
    \new_[13287]_ , \new_[13288]_ , \new_[13292]_ , \new_[13293]_ ,
    \new_[13297]_ , \new_[13298]_ , \new_[13299]_ , \new_[13303]_ ,
    \new_[13304]_ , \new_[13308]_ , \new_[13309]_ , \new_[13310]_ ,
    \new_[13314]_ , \new_[13315]_ , \new_[13319]_ , \new_[13320]_ ,
    \new_[13321]_ , \new_[13325]_ , \new_[13326]_ , \new_[13330]_ ,
    \new_[13331]_ , \new_[13332]_ , \new_[13336]_ , \new_[13337]_ ,
    \new_[13341]_ , \new_[13342]_ , \new_[13343]_ , \new_[13347]_ ,
    \new_[13348]_ , \new_[13352]_ , \new_[13353]_ , \new_[13354]_ ,
    \new_[13358]_ , \new_[13359]_ , \new_[13363]_ , \new_[13364]_ ,
    \new_[13365]_ , \new_[13369]_ , \new_[13370]_ , \new_[13374]_ ,
    \new_[13375]_ , \new_[13376]_ , \new_[13380]_ , \new_[13381]_ ,
    \new_[13385]_ , \new_[13386]_ , \new_[13387]_ , \new_[13391]_ ,
    \new_[13392]_ , \new_[13396]_ , \new_[13397]_ , \new_[13398]_ ,
    \new_[13402]_ , \new_[13403]_ , \new_[13407]_ , \new_[13408]_ ,
    \new_[13409]_ , \new_[13413]_ , \new_[13414]_ , \new_[13418]_ ,
    \new_[13419]_ , \new_[13420]_ , \new_[13424]_ , \new_[13425]_ ,
    \new_[13429]_ , \new_[13430]_ , \new_[13431]_ , \new_[13435]_ ,
    \new_[13436]_ , \new_[13440]_ , \new_[13441]_ , \new_[13442]_ ,
    \new_[13446]_ , \new_[13447]_ , \new_[13451]_ , \new_[13452]_ ,
    \new_[13453]_ , \new_[13457]_ , \new_[13458]_ , \new_[13462]_ ,
    \new_[13463]_ , \new_[13464]_ , \new_[13468]_ , \new_[13469]_ ,
    \new_[13473]_ , \new_[13474]_ , \new_[13475]_ , \new_[13479]_ ,
    \new_[13480]_ , \new_[13484]_ , \new_[13485]_ , \new_[13486]_ ,
    \new_[13490]_ , \new_[13491]_ , \new_[13495]_ , \new_[13496]_ ,
    \new_[13497]_ , \new_[13501]_ , \new_[13502]_ , \new_[13506]_ ,
    \new_[13507]_ , \new_[13508]_ , \new_[13512]_ , \new_[13513]_ ,
    \new_[13517]_ , \new_[13518]_ , \new_[13519]_ , \new_[13523]_ ,
    \new_[13524]_ , \new_[13528]_ , \new_[13529]_ , \new_[13530]_ ,
    \new_[13534]_ , \new_[13535]_ , \new_[13539]_ , \new_[13540]_ ,
    \new_[13541]_ , \new_[13545]_ , \new_[13546]_ , \new_[13550]_ ,
    \new_[13551]_ , \new_[13552]_ , \new_[13556]_ , \new_[13557]_ ,
    \new_[13561]_ , \new_[13562]_ , \new_[13563]_ , \new_[13567]_ ,
    \new_[13568]_ , \new_[13572]_ , \new_[13573]_ , \new_[13574]_ ,
    \new_[13578]_ , \new_[13579]_ , \new_[13583]_ , \new_[13584]_ ,
    \new_[13585]_ , \new_[13589]_ , \new_[13590]_ , \new_[13594]_ ,
    \new_[13595]_ , \new_[13596]_ , \new_[13600]_ , \new_[13601]_ ,
    \new_[13605]_ , \new_[13606]_ , \new_[13607]_ , \new_[13611]_ ,
    \new_[13612]_ , \new_[13616]_ , \new_[13617]_ , \new_[13618]_ ,
    \new_[13622]_ , \new_[13623]_ , \new_[13627]_ , \new_[13628]_ ,
    \new_[13629]_ , \new_[13633]_ , \new_[13634]_ , \new_[13638]_ ,
    \new_[13639]_ , \new_[13640]_ , \new_[13644]_ , \new_[13645]_ ,
    \new_[13649]_ , \new_[13650]_ , \new_[13651]_ , \new_[13655]_ ,
    \new_[13656]_ , \new_[13660]_ , \new_[13661]_ , \new_[13662]_ ,
    \new_[13666]_ , \new_[13667]_ , \new_[13671]_ , \new_[13672]_ ,
    \new_[13673]_ , \new_[13677]_ , \new_[13678]_ , \new_[13682]_ ,
    \new_[13683]_ , \new_[13684]_ , \new_[13688]_ , \new_[13689]_ ,
    \new_[13693]_ , \new_[13694]_ , \new_[13695]_ , \new_[13699]_ ,
    \new_[13700]_ , \new_[13704]_ , \new_[13705]_ , \new_[13706]_ ,
    \new_[13710]_ , \new_[13711]_ , \new_[13715]_ , \new_[13716]_ ,
    \new_[13717]_ , \new_[13721]_ , \new_[13722]_ , \new_[13726]_ ,
    \new_[13727]_ , \new_[13728]_ , \new_[13732]_ , \new_[13733]_ ,
    \new_[13737]_ , \new_[13738]_ , \new_[13739]_ , \new_[13743]_ ,
    \new_[13744]_ , \new_[13748]_ , \new_[13749]_ , \new_[13750]_ ,
    \new_[13754]_ , \new_[13755]_ , \new_[13759]_ , \new_[13760]_ ,
    \new_[13761]_ , \new_[13765]_ , \new_[13766]_ , \new_[13770]_ ,
    \new_[13771]_ , \new_[13772]_ , \new_[13776]_ , \new_[13777]_ ,
    \new_[13781]_ , \new_[13782]_ , \new_[13783]_ , \new_[13787]_ ,
    \new_[13788]_ , \new_[13792]_ , \new_[13793]_ , \new_[13794]_ ,
    \new_[13798]_ , \new_[13799]_ , \new_[13803]_ , \new_[13804]_ ,
    \new_[13805]_ , \new_[13809]_ , \new_[13810]_ , \new_[13814]_ ,
    \new_[13815]_ , \new_[13816]_ , \new_[13820]_ , \new_[13821]_ ,
    \new_[13825]_ , \new_[13826]_ , \new_[13827]_ , \new_[13831]_ ,
    \new_[13832]_ , \new_[13836]_ , \new_[13837]_ , \new_[13838]_ ,
    \new_[13842]_ , \new_[13843]_ , \new_[13847]_ , \new_[13848]_ ,
    \new_[13849]_ , \new_[13853]_ , \new_[13854]_ , \new_[13858]_ ,
    \new_[13859]_ , \new_[13860]_ , \new_[13864]_ , \new_[13865]_ ,
    \new_[13869]_ , \new_[13870]_ , \new_[13871]_ , \new_[13875]_ ,
    \new_[13876]_ , \new_[13880]_ , \new_[13881]_ , \new_[13882]_ ,
    \new_[13886]_ , \new_[13887]_ , \new_[13891]_ , \new_[13892]_ ,
    \new_[13893]_ , \new_[13897]_ , \new_[13898]_ , \new_[13902]_ ,
    \new_[13903]_ , \new_[13904]_ , \new_[13908]_ , \new_[13909]_ ,
    \new_[13913]_ , \new_[13914]_ , \new_[13915]_ , \new_[13919]_ ,
    \new_[13920]_ , \new_[13924]_ , \new_[13925]_ , \new_[13926]_ ,
    \new_[13930]_ , \new_[13931]_ , \new_[13935]_ , \new_[13936]_ ,
    \new_[13937]_ , \new_[13941]_ , \new_[13942]_ , \new_[13946]_ ,
    \new_[13947]_ , \new_[13948]_ , \new_[13952]_ , \new_[13953]_ ,
    \new_[13957]_ , \new_[13958]_ , \new_[13959]_ , \new_[13963]_ ,
    \new_[13964]_ , \new_[13968]_ , \new_[13969]_ , \new_[13970]_ ,
    \new_[13974]_ , \new_[13975]_ , \new_[13979]_ , \new_[13980]_ ,
    \new_[13981]_ , \new_[13985]_ , \new_[13986]_ , \new_[13990]_ ,
    \new_[13991]_ , \new_[13992]_ , \new_[13996]_ , \new_[13997]_ ,
    \new_[14001]_ , \new_[14002]_ , \new_[14003]_ , \new_[14007]_ ,
    \new_[14008]_ , \new_[14012]_ , \new_[14013]_ , \new_[14014]_ ,
    \new_[14018]_ , \new_[14019]_ , \new_[14023]_ , \new_[14024]_ ,
    \new_[14025]_ , \new_[14029]_ , \new_[14030]_ , \new_[14034]_ ,
    \new_[14035]_ , \new_[14036]_ , \new_[14040]_ , \new_[14041]_ ,
    \new_[14045]_ , \new_[14046]_ , \new_[14047]_ , \new_[14051]_ ,
    \new_[14052]_ , \new_[14056]_ , \new_[14057]_ , \new_[14058]_ ,
    \new_[14062]_ , \new_[14063]_ , \new_[14067]_ , \new_[14068]_ ,
    \new_[14069]_ , \new_[14073]_ , \new_[14074]_ , \new_[14078]_ ,
    \new_[14079]_ , \new_[14080]_ , \new_[14084]_ , \new_[14085]_ ,
    \new_[14089]_ , \new_[14090]_ , \new_[14091]_ , \new_[14095]_ ,
    \new_[14096]_ , \new_[14100]_ , \new_[14101]_ , \new_[14102]_ ,
    \new_[14106]_ , \new_[14107]_ , \new_[14111]_ , \new_[14112]_ ,
    \new_[14113]_ , \new_[14117]_ , \new_[14118]_ , \new_[14122]_ ,
    \new_[14123]_ , \new_[14124]_ , \new_[14128]_ , \new_[14129]_ ,
    \new_[14133]_ , \new_[14134]_ , \new_[14135]_ , \new_[14139]_ ,
    \new_[14140]_ , \new_[14144]_ , \new_[14145]_ , \new_[14146]_ ,
    \new_[14150]_ , \new_[14151]_ , \new_[14155]_ , \new_[14156]_ ,
    \new_[14157]_ , \new_[14161]_ , \new_[14162]_ , \new_[14166]_ ,
    \new_[14167]_ , \new_[14168]_ , \new_[14172]_ , \new_[14173]_ ,
    \new_[14177]_ , \new_[14178]_ , \new_[14179]_ , \new_[14183]_ ,
    \new_[14184]_ , \new_[14188]_ , \new_[14189]_ , \new_[14190]_ ,
    \new_[14194]_ , \new_[14195]_ , \new_[14199]_ , \new_[14200]_ ,
    \new_[14201]_ , \new_[14205]_ , \new_[14206]_ , \new_[14210]_ ,
    \new_[14211]_ , \new_[14212]_ , \new_[14216]_ , \new_[14217]_ ,
    \new_[14221]_ , \new_[14222]_ , \new_[14223]_ , \new_[14227]_ ,
    \new_[14228]_ , \new_[14232]_ , \new_[14233]_ , \new_[14234]_ ,
    \new_[14238]_ , \new_[14239]_ , \new_[14243]_ , \new_[14244]_ ,
    \new_[14245]_ , \new_[14249]_ , \new_[14250]_ , \new_[14254]_ ,
    \new_[14255]_ , \new_[14256]_ , \new_[14260]_ , \new_[14261]_ ,
    \new_[14265]_ , \new_[14266]_ , \new_[14267]_ , \new_[14271]_ ,
    \new_[14272]_ , \new_[14276]_ , \new_[14277]_ , \new_[14278]_ ,
    \new_[14282]_ , \new_[14283]_ , \new_[14287]_ , \new_[14288]_ ,
    \new_[14289]_ , \new_[14293]_ , \new_[14294]_ , \new_[14298]_ ,
    \new_[14299]_ , \new_[14300]_ , \new_[14304]_ , \new_[14305]_ ,
    \new_[14309]_ , \new_[14310]_ , \new_[14311]_ , \new_[14315]_ ,
    \new_[14316]_ , \new_[14320]_ , \new_[14321]_ , \new_[14322]_ ,
    \new_[14326]_ , \new_[14327]_ , \new_[14331]_ , \new_[14332]_ ,
    \new_[14333]_ , \new_[14337]_ , \new_[14338]_ , \new_[14342]_ ,
    \new_[14343]_ , \new_[14344]_ , \new_[14348]_ , \new_[14349]_ ,
    \new_[14353]_ , \new_[14354]_ , \new_[14355]_ , \new_[14359]_ ,
    \new_[14360]_ , \new_[14364]_ , \new_[14365]_ , \new_[14366]_ ,
    \new_[14370]_ , \new_[14371]_ , \new_[14375]_ , \new_[14376]_ ,
    \new_[14377]_ , \new_[14381]_ , \new_[14382]_ , \new_[14386]_ ,
    \new_[14387]_ , \new_[14388]_ , \new_[14392]_ , \new_[14393]_ ,
    \new_[14397]_ , \new_[14398]_ , \new_[14399]_ , \new_[14403]_ ,
    \new_[14404]_ , \new_[14408]_ , \new_[14409]_ , \new_[14410]_ ,
    \new_[14414]_ , \new_[14415]_ , \new_[14419]_ , \new_[14420]_ ,
    \new_[14421]_ , \new_[14425]_ , \new_[14426]_ , \new_[14430]_ ,
    \new_[14431]_ , \new_[14432]_ , \new_[14436]_ , \new_[14437]_ ,
    \new_[14441]_ , \new_[14442]_ , \new_[14443]_ , \new_[14447]_ ,
    \new_[14448]_ , \new_[14452]_ , \new_[14453]_ , \new_[14454]_ ,
    \new_[14458]_ , \new_[14459]_ , \new_[14463]_ , \new_[14464]_ ,
    \new_[14465]_ , \new_[14469]_ , \new_[14470]_ , \new_[14474]_ ,
    \new_[14475]_ , \new_[14476]_ , \new_[14480]_ , \new_[14481]_ ,
    \new_[14485]_ , \new_[14486]_ , \new_[14487]_ , \new_[14491]_ ,
    \new_[14492]_ , \new_[14496]_ , \new_[14497]_ , \new_[14498]_ ,
    \new_[14502]_ , \new_[14503]_ , \new_[14507]_ , \new_[14508]_ ,
    \new_[14509]_ , \new_[14513]_ , \new_[14514]_ , \new_[14518]_ ,
    \new_[14519]_ , \new_[14520]_ , \new_[14524]_ , \new_[14525]_ ,
    \new_[14529]_ , \new_[14530]_ , \new_[14531]_ , \new_[14535]_ ,
    \new_[14536]_ , \new_[14540]_ , \new_[14541]_ , \new_[14542]_ ,
    \new_[14546]_ , \new_[14547]_ , \new_[14551]_ , \new_[14552]_ ,
    \new_[14553]_ , \new_[14557]_ , \new_[14558]_ , \new_[14562]_ ,
    \new_[14563]_ , \new_[14564]_ , \new_[14568]_ , \new_[14569]_ ,
    \new_[14573]_ , \new_[14574]_ , \new_[14575]_ , \new_[14579]_ ,
    \new_[14580]_ , \new_[14584]_ , \new_[14585]_ , \new_[14586]_ ,
    \new_[14590]_ , \new_[14591]_ , \new_[14595]_ , \new_[14596]_ ,
    \new_[14597]_ , \new_[14601]_ , \new_[14602]_ , \new_[14606]_ ,
    \new_[14607]_ , \new_[14608]_ , \new_[14612]_ , \new_[14613]_ ,
    \new_[14617]_ , \new_[14618]_ , \new_[14619]_ , \new_[14623]_ ,
    \new_[14624]_ , \new_[14628]_ , \new_[14629]_ , \new_[14630]_ ,
    \new_[14634]_ , \new_[14635]_ , \new_[14639]_ , \new_[14640]_ ,
    \new_[14641]_ , \new_[14645]_ , \new_[14646]_ , \new_[14650]_ ,
    \new_[14651]_ , \new_[14652]_ , \new_[14656]_ , \new_[14657]_ ,
    \new_[14661]_ , \new_[14662]_ , \new_[14663]_ , \new_[14667]_ ,
    \new_[14668]_ , \new_[14672]_ , \new_[14673]_ , \new_[14674]_ ,
    \new_[14678]_ , \new_[14679]_ , \new_[14683]_ , \new_[14684]_ ,
    \new_[14685]_ , \new_[14689]_ , \new_[14690]_ , \new_[14694]_ ,
    \new_[14695]_ , \new_[14696]_ , \new_[14700]_ , \new_[14701]_ ,
    \new_[14705]_ , \new_[14706]_ , \new_[14707]_ , \new_[14711]_ ,
    \new_[14712]_ , \new_[14716]_ , \new_[14717]_ , \new_[14718]_ ,
    \new_[14722]_ , \new_[14723]_ , \new_[14727]_ , \new_[14728]_ ,
    \new_[14729]_ , \new_[14733]_ , \new_[14734]_ , \new_[14738]_ ,
    \new_[14739]_ , \new_[14740]_ , \new_[14744]_ , \new_[14745]_ ,
    \new_[14749]_ , \new_[14750]_ , \new_[14751]_ , \new_[14755]_ ,
    \new_[14756]_ , \new_[14760]_ , \new_[14761]_ , \new_[14762]_ ,
    \new_[14766]_ , \new_[14767]_ , \new_[14771]_ , \new_[14772]_ ,
    \new_[14773]_ , \new_[14777]_ , \new_[14778]_ , \new_[14782]_ ,
    \new_[14783]_ , \new_[14784]_ , \new_[14788]_ , \new_[14789]_ ,
    \new_[14793]_ , \new_[14794]_ , \new_[14795]_ , \new_[14799]_ ,
    \new_[14800]_ , \new_[14804]_ , \new_[14805]_ , \new_[14806]_ ,
    \new_[14810]_ , \new_[14811]_ , \new_[14815]_ , \new_[14816]_ ,
    \new_[14817]_ , \new_[14821]_ , \new_[14822]_ , \new_[14826]_ ,
    \new_[14827]_ , \new_[14828]_ , \new_[14832]_ , \new_[14833]_ ,
    \new_[14837]_ , \new_[14838]_ , \new_[14839]_ , \new_[14843]_ ,
    \new_[14844]_ , \new_[14848]_ , \new_[14849]_ , \new_[14850]_ ,
    \new_[14854]_ , \new_[14855]_ , \new_[14859]_ , \new_[14860]_ ,
    \new_[14861]_ , \new_[14865]_ , \new_[14866]_ , \new_[14869]_ ,
    \new_[14872]_ , \new_[14873]_ , \new_[14874]_ , \new_[14878]_ ,
    \new_[14879]_ , \new_[14883]_ , \new_[14884]_ , \new_[14885]_ ,
    \new_[14889]_ , \new_[14890]_ , \new_[14893]_ , \new_[14896]_ ,
    \new_[14897]_ , \new_[14898]_ , \new_[14902]_ , \new_[14903]_ ,
    \new_[14907]_ , \new_[14908]_ , \new_[14909]_ , \new_[14913]_ ,
    \new_[14914]_ , \new_[14917]_ , \new_[14920]_ , \new_[14921]_ ,
    \new_[14922]_ , \new_[14926]_ , \new_[14927]_ , \new_[14931]_ ,
    \new_[14932]_ , \new_[14933]_ , \new_[14937]_ , \new_[14938]_ ,
    \new_[14941]_ , \new_[14944]_ , \new_[14945]_ , \new_[14946]_ ,
    \new_[14950]_ , \new_[14951]_ , \new_[14955]_ , \new_[14956]_ ,
    \new_[14957]_ , \new_[14961]_ , \new_[14962]_ , \new_[14965]_ ,
    \new_[14968]_ , \new_[14969]_ , \new_[14970]_ , \new_[14974]_ ,
    \new_[14975]_ , \new_[14979]_ , \new_[14980]_ , \new_[14981]_ ,
    \new_[14985]_ , \new_[14986]_ , \new_[14989]_ , \new_[14992]_ ,
    \new_[14993]_ , \new_[14994]_ , \new_[14998]_ , \new_[14999]_ ,
    \new_[15003]_ , \new_[15004]_ , \new_[15005]_ , \new_[15009]_ ,
    \new_[15010]_ , \new_[15013]_ , \new_[15016]_ , \new_[15017]_ ,
    \new_[15018]_ , \new_[15022]_ , \new_[15023]_ , \new_[15027]_ ,
    \new_[15028]_ , \new_[15029]_ , \new_[15033]_ , \new_[15034]_ ,
    \new_[15037]_ , \new_[15040]_ , \new_[15041]_ , \new_[15042]_ ,
    \new_[15046]_ , \new_[15047]_ , \new_[15051]_ , \new_[15052]_ ,
    \new_[15053]_ , \new_[15057]_ , \new_[15058]_ , \new_[15061]_ ,
    \new_[15064]_ , \new_[15065]_ , \new_[15066]_ , \new_[15070]_ ,
    \new_[15071]_ , \new_[15075]_ , \new_[15076]_ , \new_[15077]_ ,
    \new_[15081]_ , \new_[15082]_ , \new_[15085]_ , \new_[15088]_ ,
    \new_[15089]_ , \new_[15090]_ , \new_[15094]_ , \new_[15095]_ ,
    \new_[15099]_ , \new_[15100]_ , \new_[15101]_ , \new_[15105]_ ,
    \new_[15106]_ , \new_[15109]_ , \new_[15112]_ , \new_[15113]_ ,
    \new_[15114]_ , \new_[15118]_ , \new_[15119]_ , \new_[15123]_ ,
    \new_[15124]_ , \new_[15125]_ , \new_[15129]_ , \new_[15130]_ ,
    \new_[15133]_ , \new_[15136]_ , \new_[15137]_ , \new_[15138]_ ,
    \new_[15142]_ , \new_[15143]_ , \new_[15147]_ , \new_[15148]_ ,
    \new_[15149]_ , \new_[15153]_ , \new_[15154]_ , \new_[15157]_ ,
    \new_[15160]_ , \new_[15161]_ , \new_[15162]_ , \new_[15166]_ ,
    \new_[15167]_ , \new_[15171]_ , \new_[15172]_ , \new_[15173]_ ,
    \new_[15177]_ , \new_[15178]_ , \new_[15181]_ , \new_[15184]_ ,
    \new_[15185]_ , \new_[15186]_ , \new_[15190]_ , \new_[15191]_ ,
    \new_[15195]_ , \new_[15196]_ , \new_[15197]_ , \new_[15201]_ ,
    \new_[15202]_ , \new_[15205]_ , \new_[15208]_ , \new_[15209]_ ,
    \new_[15210]_ , \new_[15214]_ , \new_[15215]_ , \new_[15219]_ ,
    \new_[15220]_ , \new_[15221]_ , \new_[15225]_ , \new_[15226]_ ,
    \new_[15229]_ , \new_[15232]_ , \new_[15233]_ , \new_[15234]_ ,
    \new_[15238]_ , \new_[15239]_ , \new_[15243]_ , \new_[15244]_ ,
    \new_[15245]_ , \new_[15249]_ , \new_[15250]_ , \new_[15253]_ ,
    \new_[15256]_ , \new_[15257]_ , \new_[15258]_ , \new_[15262]_ ,
    \new_[15263]_ , \new_[15267]_ , \new_[15268]_ , \new_[15269]_ ,
    \new_[15273]_ , \new_[15274]_ , \new_[15277]_ , \new_[15280]_ ,
    \new_[15281]_ , \new_[15282]_ , \new_[15286]_ , \new_[15287]_ ,
    \new_[15291]_ , \new_[15292]_ , \new_[15293]_ , \new_[15297]_ ,
    \new_[15298]_ , \new_[15301]_ , \new_[15304]_ , \new_[15305]_ ,
    \new_[15306]_ , \new_[15310]_ , \new_[15311]_ , \new_[15315]_ ,
    \new_[15316]_ , \new_[15317]_ , \new_[15321]_ , \new_[15322]_ ,
    \new_[15325]_ , \new_[15328]_ , \new_[15329]_ , \new_[15330]_ ,
    \new_[15334]_ , \new_[15335]_ , \new_[15339]_ , \new_[15340]_ ,
    \new_[15341]_ , \new_[15345]_ , \new_[15346]_ , \new_[15349]_ ,
    \new_[15352]_ , \new_[15353]_ , \new_[15354]_ , \new_[15358]_ ,
    \new_[15359]_ , \new_[15363]_ , \new_[15364]_ , \new_[15365]_ ,
    \new_[15369]_ , \new_[15370]_ , \new_[15373]_ , \new_[15376]_ ,
    \new_[15377]_ , \new_[15378]_ , \new_[15382]_ , \new_[15383]_ ,
    \new_[15387]_ , \new_[15388]_ , \new_[15389]_ , \new_[15393]_ ,
    \new_[15394]_ , \new_[15397]_ , \new_[15400]_ , \new_[15401]_ ,
    \new_[15402]_ , \new_[15406]_ , \new_[15407]_ , \new_[15411]_ ,
    \new_[15412]_ , \new_[15413]_ , \new_[15417]_ , \new_[15418]_ ,
    \new_[15421]_ , \new_[15424]_ , \new_[15425]_ , \new_[15426]_ ,
    \new_[15430]_ , \new_[15431]_ , \new_[15435]_ , \new_[15436]_ ,
    \new_[15437]_ , \new_[15441]_ , \new_[15442]_ , \new_[15445]_ ,
    \new_[15448]_ , \new_[15449]_ , \new_[15450]_ , \new_[15454]_ ,
    \new_[15455]_ , \new_[15459]_ , \new_[15460]_ , \new_[15461]_ ,
    \new_[15465]_ , \new_[15466]_ , \new_[15469]_ , \new_[15472]_ ,
    \new_[15473]_ , \new_[15474]_ , \new_[15478]_ , \new_[15479]_ ,
    \new_[15483]_ , \new_[15484]_ , \new_[15485]_ , \new_[15489]_ ,
    \new_[15490]_ , \new_[15493]_ , \new_[15496]_ , \new_[15497]_ ,
    \new_[15498]_ , \new_[15502]_ , \new_[15503]_ , \new_[15507]_ ,
    \new_[15508]_ , \new_[15509]_ , \new_[15513]_ , \new_[15514]_ ,
    \new_[15517]_ , \new_[15520]_ , \new_[15521]_ , \new_[15522]_ ,
    \new_[15526]_ , \new_[15527]_ , \new_[15531]_ , \new_[15532]_ ,
    \new_[15533]_ , \new_[15537]_ , \new_[15538]_ , \new_[15541]_ ,
    \new_[15544]_ , \new_[15545]_ , \new_[15546]_ , \new_[15550]_ ,
    \new_[15551]_ , \new_[15555]_ , \new_[15556]_ , \new_[15557]_ ,
    \new_[15561]_ , \new_[15562]_ , \new_[15565]_ , \new_[15568]_ ,
    \new_[15569]_ , \new_[15570]_ , \new_[15574]_ , \new_[15575]_ ,
    \new_[15579]_ , \new_[15580]_ , \new_[15581]_ , \new_[15585]_ ,
    \new_[15586]_ , \new_[15589]_ , \new_[15592]_ , \new_[15593]_ ,
    \new_[15594]_ , \new_[15598]_ , \new_[15599]_ , \new_[15603]_ ,
    \new_[15604]_ , \new_[15605]_ , \new_[15609]_ , \new_[15610]_ ,
    \new_[15613]_ , \new_[15616]_ , \new_[15617]_ , \new_[15618]_ ,
    \new_[15622]_ , \new_[15623]_ , \new_[15627]_ , \new_[15628]_ ,
    \new_[15629]_ , \new_[15633]_ , \new_[15634]_ , \new_[15637]_ ,
    \new_[15640]_ , \new_[15641]_ , \new_[15642]_ , \new_[15646]_ ,
    \new_[15647]_ , \new_[15651]_ , \new_[15652]_ , \new_[15653]_ ,
    \new_[15657]_ , \new_[15658]_ , \new_[15661]_ , \new_[15664]_ ,
    \new_[15665]_ , \new_[15666]_ , \new_[15670]_ , \new_[15671]_ ,
    \new_[15675]_ , \new_[15676]_ , \new_[15677]_ , \new_[15681]_ ,
    \new_[15682]_ , \new_[15685]_ , \new_[15688]_ , \new_[15689]_ ,
    \new_[15690]_ , \new_[15694]_ , \new_[15695]_ , \new_[15699]_ ,
    \new_[15700]_ , \new_[15701]_ , \new_[15705]_ , \new_[15706]_ ,
    \new_[15709]_ , \new_[15712]_ , \new_[15713]_ , \new_[15714]_ ,
    \new_[15718]_ , \new_[15719]_ , \new_[15723]_ , \new_[15724]_ ,
    \new_[15725]_ , \new_[15729]_ , \new_[15730]_ , \new_[15733]_ ,
    \new_[15736]_ , \new_[15737]_ , \new_[15738]_ , \new_[15742]_ ,
    \new_[15743]_ , \new_[15747]_ , \new_[15748]_ , \new_[15749]_ ,
    \new_[15753]_ , \new_[15754]_ , \new_[15757]_ , \new_[15760]_ ,
    \new_[15761]_ , \new_[15762]_ , \new_[15766]_ , \new_[15767]_ ,
    \new_[15771]_ , \new_[15772]_ , \new_[15773]_ , \new_[15777]_ ,
    \new_[15778]_ , \new_[15781]_ , \new_[15784]_ , \new_[15785]_ ,
    \new_[15786]_ , \new_[15790]_ , \new_[15791]_ , \new_[15795]_ ,
    \new_[15796]_ , \new_[15797]_ , \new_[15801]_ , \new_[15802]_ ,
    \new_[15805]_ , \new_[15808]_ , \new_[15809]_ , \new_[15810]_ ,
    \new_[15814]_ , \new_[15815]_ , \new_[15819]_ , \new_[15820]_ ,
    \new_[15821]_ , \new_[15825]_ , \new_[15826]_ , \new_[15829]_ ,
    \new_[15832]_ , \new_[15833]_ , \new_[15834]_ , \new_[15838]_ ,
    \new_[15839]_ , \new_[15843]_ , \new_[15844]_ , \new_[15845]_ ,
    \new_[15849]_ , \new_[15850]_ , \new_[15853]_ , \new_[15856]_ ,
    \new_[15857]_ , \new_[15858]_ , \new_[15862]_ , \new_[15863]_ ,
    \new_[15867]_ , \new_[15868]_ , \new_[15869]_ , \new_[15873]_ ,
    \new_[15874]_ , \new_[15877]_ , \new_[15880]_ , \new_[15881]_ ,
    \new_[15882]_ , \new_[15886]_ , \new_[15887]_ , \new_[15891]_ ,
    \new_[15892]_ , \new_[15893]_ , \new_[15897]_ , \new_[15898]_ ,
    \new_[15901]_ , \new_[15904]_ , \new_[15905]_ , \new_[15906]_ ,
    \new_[15910]_ , \new_[15911]_ , \new_[15915]_ , \new_[15916]_ ,
    \new_[15917]_ , \new_[15921]_ , \new_[15922]_ , \new_[15925]_ ,
    \new_[15928]_ , \new_[15929]_ , \new_[15930]_ , \new_[15934]_ ,
    \new_[15935]_ , \new_[15939]_ , \new_[15940]_ , \new_[15941]_ ,
    \new_[15945]_ , \new_[15946]_ , \new_[15949]_ , \new_[15952]_ ,
    \new_[15953]_ , \new_[15954]_ , \new_[15958]_ , \new_[15959]_ ,
    \new_[15963]_ , \new_[15964]_ , \new_[15965]_ , \new_[15969]_ ,
    \new_[15970]_ , \new_[15973]_ , \new_[15976]_ , \new_[15977]_ ,
    \new_[15978]_ , \new_[15982]_ , \new_[15983]_ , \new_[15987]_ ,
    \new_[15988]_ , \new_[15989]_ , \new_[15993]_ , \new_[15994]_ ,
    \new_[15997]_ , \new_[16000]_ , \new_[16001]_ , \new_[16002]_ ,
    \new_[16006]_ , \new_[16007]_ , \new_[16011]_ , \new_[16012]_ ,
    \new_[16013]_ , \new_[16017]_ , \new_[16018]_ , \new_[16021]_ ,
    \new_[16024]_ , \new_[16025]_ , \new_[16026]_ , \new_[16030]_ ,
    \new_[16031]_ , \new_[16035]_ , \new_[16036]_ , \new_[16037]_ ,
    \new_[16041]_ , \new_[16042]_ , \new_[16045]_ , \new_[16048]_ ,
    \new_[16049]_ , \new_[16050]_ , \new_[16054]_ , \new_[16055]_ ,
    \new_[16059]_ , \new_[16060]_ , \new_[16061]_ , \new_[16065]_ ,
    \new_[16066]_ , \new_[16069]_ , \new_[16072]_ , \new_[16073]_ ,
    \new_[16074]_ , \new_[16078]_ , \new_[16079]_ , \new_[16083]_ ,
    \new_[16084]_ , \new_[16085]_ , \new_[16089]_ , \new_[16090]_ ,
    \new_[16093]_ , \new_[16096]_ , \new_[16097]_ , \new_[16098]_ ,
    \new_[16102]_ , \new_[16103]_ , \new_[16107]_ , \new_[16108]_ ,
    \new_[16109]_ , \new_[16113]_ , \new_[16114]_ , \new_[16117]_ ,
    \new_[16120]_ , \new_[16121]_ , \new_[16122]_ , \new_[16126]_ ,
    \new_[16127]_ , \new_[16131]_ , \new_[16132]_ , \new_[16133]_ ,
    \new_[16137]_ , \new_[16138]_ , \new_[16141]_ , \new_[16144]_ ,
    \new_[16145]_ , \new_[16146]_ , \new_[16150]_ , \new_[16151]_ ,
    \new_[16155]_ , \new_[16156]_ , \new_[16157]_ , \new_[16161]_ ,
    \new_[16162]_ , \new_[16165]_ , \new_[16168]_ , \new_[16169]_ ,
    \new_[16170]_ , \new_[16174]_ , \new_[16175]_ , \new_[16179]_ ,
    \new_[16180]_ , \new_[16181]_ , \new_[16185]_ , \new_[16186]_ ,
    \new_[16189]_ , \new_[16192]_ , \new_[16193]_ , \new_[16194]_ ,
    \new_[16198]_ , \new_[16199]_ , \new_[16203]_ , \new_[16204]_ ,
    \new_[16205]_ , \new_[16209]_ , \new_[16210]_ , \new_[16213]_ ,
    \new_[16216]_ , \new_[16217]_ , \new_[16218]_ , \new_[16222]_ ,
    \new_[16223]_ , \new_[16227]_ , \new_[16228]_ , \new_[16229]_ ,
    \new_[16233]_ , \new_[16234]_ , \new_[16237]_ , \new_[16240]_ ,
    \new_[16241]_ , \new_[16242]_ , \new_[16246]_ , \new_[16247]_ ,
    \new_[16251]_ , \new_[16252]_ , \new_[16253]_ , \new_[16257]_ ,
    \new_[16258]_ , \new_[16261]_ , \new_[16264]_ , \new_[16265]_ ,
    \new_[16266]_ , \new_[16270]_ , \new_[16271]_ , \new_[16275]_ ,
    \new_[16276]_ , \new_[16277]_ , \new_[16281]_ , \new_[16282]_ ,
    \new_[16285]_ , \new_[16288]_ , \new_[16289]_ , \new_[16290]_ ,
    \new_[16294]_ , \new_[16295]_ , \new_[16299]_ , \new_[16300]_ ,
    \new_[16301]_ , \new_[16305]_ , \new_[16306]_ , \new_[16309]_ ,
    \new_[16312]_ , \new_[16313]_ , \new_[16314]_ , \new_[16318]_ ,
    \new_[16319]_ , \new_[16323]_ , \new_[16324]_ , \new_[16325]_ ,
    \new_[16329]_ , \new_[16330]_ , \new_[16333]_ , \new_[16336]_ ,
    \new_[16337]_ , \new_[16338]_ , \new_[16342]_ , \new_[16343]_ ,
    \new_[16347]_ , \new_[16348]_ , \new_[16349]_ , \new_[16353]_ ,
    \new_[16354]_ , \new_[16357]_ , \new_[16360]_ , \new_[16361]_ ,
    \new_[16362]_ , \new_[16366]_ , \new_[16367]_ , \new_[16371]_ ,
    \new_[16372]_ , \new_[16373]_ , \new_[16377]_ , \new_[16378]_ ,
    \new_[16381]_ , \new_[16384]_ , \new_[16385]_ , \new_[16386]_ ,
    \new_[16390]_ , \new_[16391]_ , \new_[16395]_ , \new_[16396]_ ,
    \new_[16397]_ , \new_[16401]_ , \new_[16402]_ , \new_[16405]_ ,
    \new_[16408]_ , \new_[16409]_ , \new_[16410]_ , \new_[16414]_ ,
    \new_[16415]_ , \new_[16419]_ , \new_[16420]_ , \new_[16421]_ ,
    \new_[16425]_ , \new_[16426]_ , \new_[16429]_ , \new_[16432]_ ,
    \new_[16433]_ , \new_[16434]_ , \new_[16438]_ , \new_[16439]_ ,
    \new_[16443]_ , \new_[16444]_ , \new_[16445]_ , \new_[16449]_ ,
    \new_[16450]_ , \new_[16453]_ , \new_[16456]_ , \new_[16457]_ ,
    \new_[16458]_ , \new_[16462]_ , \new_[16463]_ , \new_[16467]_ ,
    \new_[16468]_ , \new_[16469]_ , \new_[16473]_ , \new_[16474]_ ,
    \new_[16477]_ , \new_[16480]_ , \new_[16481]_ , \new_[16482]_ ,
    \new_[16486]_ , \new_[16487]_ , \new_[16491]_ , \new_[16492]_ ,
    \new_[16493]_ , \new_[16497]_ , \new_[16498]_ , \new_[16501]_ ,
    \new_[16504]_ , \new_[16505]_ , \new_[16506]_ , \new_[16510]_ ,
    \new_[16511]_ , \new_[16515]_ , \new_[16516]_ , \new_[16517]_ ,
    \new_[16521]_ , \new_[16522]_ , \new_[16525]_ , \new_[16528]_ ,
    \new_[16529]_ , \new_[16530]_ , \new_[16534]_ , \new_[16535]_ ,
    \new_[16539]_ , \new_[16540]_ , \new_[16541]_ , \new_[16545]_ ,
    \new_[16546]_ , \new_[16549]_ , \new_[16552]_ , \new_[16553]_ ,
    \new_[16554]_ , \new_[16558]_ , \new_[16559]_ , \new_[16563]_ ,
    \new_[16564]_ , \new_[16565]_ , \new_[16569]_ , \new_[16570]_ ,
    \new_[16573]_ , \new_[16576]_ , \new_[16577]_ , \new_[16578]_ ,
    \new_[16582]_ , \new_[16583]_ , \new_[16587]_ , \new_[16588]_ ,
    \new_[16589]_ , \new_[16593]_ , \new_[16594]_ , \new_[16597]_ ,
    \new_[16600]_ , \new_[16601]_ , \new_[16602]_ , \new_[16606]_ ,
    \new_[16607]_ , \new_[16611]_ , \new_[16612]_ , \new_[16613]_ ,
    \new_[16617]_ , \new_[16618]_ , \new_[16621]_ , \new_[16624]_ ,
    \new_[16625]_ , \new_[16626]_ , \new_[16630]_ , \new_[16631]_ ,
    \new_[16635]_ , \new_[16636]_ , \new_[16637]_ , \new_[16641]_ ,
    \new_[16642]_ , \new_[16645]_ , \new_[16648]_ , \new_[16649]_ ,
    \new_[16650]_ , \new_[16654]_ , \new_[16655]_ , \new_[16659]_ ,
    \new_[16660]_ , \new_[16661]_ , \new_[16665]_ , \new_[16666]_ ,
    \new_[16669]_ , \new_[16672]_ , \new_[16673]_ , \new_[16674]_ ,
    \new_[16678]_ , \new_[16679]_ , \new_[16683]_ , \new_[16684]_ ,
    \new_[16685]_ , \new_[16689]_ , \new_[16690]_ , \new_[16693]_ ,
    \new_[16696]_ , \new_[16697]_ , \new_[16698]_ , \new_[16702]_ ,
    \new_[16703]_ , \new_[16707]_ , \new_[16708]_ , \new_[16709]_ ,
    \new_[16713]_ , \new_[16714]_ , \new_[16717]_ , \new_[16720]_ ,
    \new_[16721]_ , \new_[16722]_ , \new_[16726]_ , \new_[16727]_ ,
    \new_[16731]_ , \new_[16732]_ , \new_[16733]_ , \new_[16737]_ ,
    \new_[16738]_ , \new_[16741]_ , \new_[16744]_ , \new_[16745]_ ,
    \new_[16746]_ , \new_[16750]_ , \new_[16751]_ , \new_[16755]_ ,
    \new_[16756]_ , \new_[16757]_ , \new_[16761]_ , \new_[16762]_ ,
    \new_[16765]_ , \new_[16768]_ , \new_[16769]_ , \new_[16770]_ ,
    \new_[16774]_ , \new_[16775]_ , \new_[16779]_ , \new_[16780]_ ,
    \new_[16781]_ , \new_[16785]_ , \new_[16786]_ , \new_[16789]_ ,
    \new_[16792]_ , \new_[16793]_ , \new_[16794]_ , \new_[16798]_ ,
    \new_[16799]_ , \new_[16803]_ , \new_[16804]_ , \new_[16805]_ ,
    \new_[16809]_ , \new_[16810]_ , \new_[16813]_ , \new_[16816]_ ,
    \new_[16817]_ , \new_[16818]_ , \new_[16822]_ , \new_[16823]_ ,
    \new_[16827]_ , \new_[16828]_ , \new_[16829]_ , \new_[16833]_ ,
    \new_[16834]_ , \new_[16837]_ , \new_[16840]_ , \new_[16841]_ ,
    \new_[16842]_ , \new_[16846]_ , \new_[16847]_ , \new_[16851]_ ,
    \new_[16852]_ , \new_[16853]_ , \new_[16857]_ , \new_[16858]_ ,
    \new_[16861]_ , \new_[16864]_ , \new_[16865]_ , \new_[16866]_ ,
    \new_[16870]_ , \new_[16871]_ , \new_[16875]_ , \new_[16876]_ ,
    \new_[16877]_ , \new_[16881]_ , \new_[16882]_ , \new_[16885]_ ,
    \new_[16888]_ , \new_[16889]_ , \new_[16890]_ , \new_[16894]_ ,
    \new_[16895]_ , \new_[16899]_ , \new_[16900]_ , \new_[16901]_ ,
    \new_[16905]_ , \new_[16906]_ , \new_[16909]_ , \new_[16912]_ ,
    \new_[16913]_ , \new_[16914]_ , \new_[16918]_ , \new_[16919]_ ,
    \new_[16923]_ , \new_[16924]_ , \new_[16925]_ , \new_[16929]_ ,
    \new_[16930]_ , \new_[16933]_ , \new_[16936]_ , \new_[16937]_ ,
    \new_[16938]_ , \new_[16942]_ , \new_[16943]_ , \new_[16947]_ ,
    \new_[16948]_ , \new_[16949]_ , \new_[16953]_ , \new_[16954]_ ,
    \new_[16957]_ , \new_[16960]_ , \new_[16961]_ , \new_[16962]_ ,
    \new_[16966]_ , \new_[16967]_ , \new_[16971]_ , \new_[16972]_ ,
    \new_[16973]_ , \new_[16977]_ , \new_[16978]_ , \new_[16981]_ ,
    \new_[16984]_ , \new_[16985]_ , \new_[16986]_ , \new_[16990]_ ,
    \new_[16991]_ , \new_[16995]_ , \new_[16996]_ , \new_[16997]_ ,
    \new_[17001]_ , \new_[17002]_ , \new_[17005]_ , \new_[17008]_ ,
    \new_[17009]_ , \new_[17010]_ , \new_[17014]_ , \new_[17015]_ ,
    \new_[17019]_ , \new_[17020]_ , \new_[17021]_ , \new_[17025]_ ,
    \new_[17026]_ , \new_[17029]_ , \new_[17032]_ , \new_[17033]_ ,
    \new_[17034]_ , \new_[17038]_ , \new_[17039]_ , \new_[17043]_ ,
    \new_[17044]_ , \new_[17045]_ , \new_[17049]_ , \new_[17050]_ ,
    \new_[17053]_ , \new_[17056]_ , \new_[17057]_ , \new_[17058]_ ,
    \new_[17062]_ , \new_[17063]_ , \new_[17067]_ , \new_[17068]_ ,
    \new_[17069]_ , \new_[17073]_ , \new_[17074]_ , \new_[17077]_ ,
    \new_[17080]_ , \new_[17081]_ , \new_[17082]_ , \new_[17086]_ ,
    \new_[17087]_ , \new_[17091]_ , \new_[17092]_ , \new_[17093]_ ,
    \new_[17097]_ , \new_[17098]_ , \new_[17101]_ , \new_[17104]_ ,
    \new_[17105]_ , \new_[17106]_ , \new_[17110]_ , \new_[17111]_ ,
    \new_[17115]_ , \new_[17116]_ , \new_[17117]_ , \new_[17121]_ ,
    \new_[17122]_ , \new_[17125]_ , \new_[17128]_ , \new_[17129]_ ,
    \new_[17130]_ , \new_[17134]_ , \new_[17135]_ , \new_[17139]_ ,
    \new_[17140]_ , \new_[17141]_ , \new_[17145]_ , \new_[17146]_ ,
    \new_[17149]_ , \new_[17152]_ , \new_[17153]_ , \new_[17154]_ ,
    \new_[17158]_ , \new_[17159]_ , \new_[17163]_ , \new_[17164]_ ,
    \new_[17165]_ , \new_[17169]_ , \new_[17170]_ , \new_[17173]_ ,
    \new_[17176]_ , \new_[17177]_ , \new_[17178]_ , \new_[17182]_ ,
    \new_[17183]_ , \new_[17187]_ , \new_[17188]_ , \new_[17189]_ ,
    \new_[17193]_ , \new_[17194]_ , \new_[17197]_ , \new_[17200]_ ,
    \new_[17201]_ , \new_[17202]_ , \new_[17206]_ , \new_[17207]_ ,
    \new_[17211]_ , \new_[17212]_ , \new_[17213]_ , \new_[17217]_ ,
    \new_[17218]_ , \new_[17221]_ , \new_[17224]_ , \new_[17225]_ ,
    \new_[17226]_ , \new_[17230]_ , \new_[17231]_ , \new_[17235]_ ,
    \new_[17236]_ , \new_[17237]_ , \new_[17241]_ , \new_[17242]_ ,
    \new_[17245]_ , \new_[17248]_ , \new_[17249]_ , \new_[17250]_ ,
    \new_[17254]_ , \new_[17255]_ , \new_[17259]_ , \new_[17260]_ ,
    \new_[17261]_ , \new_[17265]_ , \new_[17266]_ , \new_[17269]_ ,
    \new_[17272]_ , \new_[17273]_ , \new_[17274]_ , \new_[17278]_ ,
    \new_[17279]_ , \new_[17283]_ , \new_[17284]_ , \new_[17285]_ ,
    \new_[17289]_ , \new_[17290]_ , \new_[17293]_ , \new_[17296]_ ,
    \new_[17297]_ , \new_[17298]_ , \new_[17302]_ , \new_[17303]_ ,
    \new_[17307]_ , \new_[17308]_ , \new_[17309]_ , \new_[17313]_ ,
    \new_[17314]_ , \new_[17317]_ , \new_[17320]_ , \new_[17321]_ ,
    \new_[17322]_ , \new_[17326]_ , \new_[17327]_ , \new_[17331]_ ,
    \new_[17332]_ , \new_[17333]_ , \new_[17337]_ , \new_[17338]_ ,
    \new_[17341]_ , \new_[17344]_ , \new_[17345]_ , \new_[17346]_ ,
    \new_[17350]_ , \new_[17351]_ , \new_[17355]_ , \new_[17356]_ ,
    \new_[17357]_ , \new_[17361]_ , \new_[17362]_ , \new_[17365]_ ,
    \new_[17368]_ , \new_[17369]_ , \new_[17370]_ , \new_[17374]_ ,
    \new_[17375]_ , \new_[17379]_ , \new_[17380]_ , \new_[17381]_ ,
    \new_[17385]_ , \new_[17386]_ , \new_[17389]_ , \new_[17392]_ ,
    \new_[17393]_ , \new_[17394]_ , \new_[17398]_ , \new_[17399]_ ,
    \new_[17403]_ , \new_[17404]_ , \new_[17405]_ , \new_[17409]_ ,
    \new_[17410]_ , \new_[17413]_ , \new_[17416]_ , \new_[17417]_ ,
    \new_[17418]_ , \new_[17422]_ , \new_[17423]_ , \new_[17427]_ ,
    \new_[17428]_ , \new_[17429]_ , \new_[17433]_ , \new_[17434]_ ,
    \new_[17437]_ , \new_[17440]_ , \new_[17441]_ , \new_[17442]_ ,
    \new_[17446]_ , \new_[17447]_ , \new_[17451]_ , \new_[17452]_ ,
    \new_[17453]_ , \new_[17457]_ , \new_[17458]_ , \new_[17461]_ ,
    \new_[17464]_ , \new_[17465]_ , \new_[17466]_ , \new_[17470]_ ,
    \new_[17471]_ , \new_[17475]_ , \new_[17476]_ , \new_[17477]_ ,
    \new_[17481]_ , \new_[17482]_ , \new_[17485]_ , \new_[17488]_ ,
    \new_[17489]_ , \new_[17490]_ , \new_[17494]_ , \new_[17495]_ ,
    \new_[17499]_ , \new_[17500]_ , \new_[17501]_ , \new_[17505]_ ,
    \new_[17506]_ , \new_[17509]_ , \new_[17512]_ , \new_[17513]_ ,
    \new_[17514]_ , \new_[17518]_ , \new_[17519]_ , \new_[17523]_ ,
    \new_[17524]_ , \new_[17525]_ , \new_[17529]_ , \new_[17530]_ ,
    \new_[17533]_ , \new_[17536]_ , \new_[17537]_ , \new_[17538]_ ,
    \new_[17542]_ , \new_[17543]_ , \new_[17547]_ , \new_[17548]_ ,
    \new_[17549]_ , \new_[17553]_ , \new_[17554]_ , \new_[17557]_ ,
    \new_[17560]_ , \new_[17561]_ , \new_[17562]_ , \new_[17566]_ ,
    \new_[17567]_ , \new_[17571]_ , \new_[17572]_ , \new_[17573]_ ,
    \new_[17577]_ , \new_[17578]_ , \new_[17581]_ , \new_[17584]_ ,
    \new_[17585]_ , \new_[17586]_ , \new_[17590]_ , \new_[17591]_ ,
    \new_[17595]_ , \new_[17596]_ , \new_[17597]_ , \new_[17601]_ ,
    \new_[17602]_ , \new_[17605]_ , \new_[17608]_ , \new_[17609]_ ,
    \new_[17610]_ , \new_[17614]_ , \new_[17615]_ , \new_[17619]_ ,
    \new_[17620]_ , \new_[17621]_ , \new_[17625]_ , \new_[17626]_ ,
    \new_[17629]_ , \new_[17632]_ , \new_[17633]_ , \new_[17634]_ ,
    \new_[17638]_ , \new_[17639]_ , \new_[17643]_ , \new_[17644]_ ,
    \new_[17645]_ , \new_[17649]_ , \new_[17650]_ , \new_[17653]_ ,
    \new_[17656]_ , \new_[17657]_ , \new_[17658]_ , \new_[17662]_ ,
    \new_[17663]_ , \new_[17667]_ , \new_[17668]_ , \new_[17669]_ ,
    \new_[17673]_ , \new_[17674]_ , \new_[17677]_ , \new_[17680]_ ,
    \new_[17681]_ , \new_[17682]_ , \new_[17686]_ , \new_[17687]_ ,
    \new_[17691]_ , \new_[17692]_ , \new_[17693]_ , \new_[17697]_ ,
    \new_[17698]_ , \new_[17701]_ , \new_[17704]_ , \new_[17705]_ ,
    \new_[17706]_ , \new_[17710]_ , \new_[17711]_ , \new_[17715]_ ,
    \new_[17716]_ , \new_[17717]_ , \new_[17721]_ , \new_[17722]_ ,
    \new_[17725]_ , \new_[17728]_ , \new_[17729]_ , \new_[17730]_ ,
    \new_[17734]_ , \new_[17735]_ , \new_[17739]_ , \new_[17740]_ ,
    \new_[17741]_ , \new_[17745]_ , \new_[17746]_ , \new_[17749]_ ,
    \new_[17752]_ , \new_[17753]_ , \new_[17754]_ , \new_[17758]_ ,
    \new_[17759]_ , \new_[17763]_ , \new_[17764]_ , \new_[17765]_ ,
    \new_[17769]_ , \new_[17770]_ , \new_[17773]_ , \new_[17776]_ ,
    \new_[17777]_ , \new_[17778]_ , \new_[17782]_ , \new_[17783]_ ,
    \new_[17787]_ , \new_[17788]_ , \new_[17789]_ , \new_[17793]_ ,
    \new_[17794]_ , \new_[17797]_ , \new_[17800]_ , \new_[17801]_ ,
    \new_[17802]_ , \new_[17806]_ , \new_[17807]_ , \new_[17811]_ ,
    \new_[17812]_ , \new_[17813]_ , \new_[17817]_ , \new_[17818]_ ,
    \new_[17821]_ , \new_[17824]_ , \new_[17825]_ , \new_[17826]_ ,
    \new_[17830]_ , \new_[17831]_ , \new_[17835]_ , \new_[17836]_ ,
    \new_[17837]_ , \new_[17841]_ , \new_[17842]_ , \new_[17845]_ ,
    \new_[17848]_ , \new_[17849]_ , \new_[17850]_ , \new_[17854]_ ,
    \new_[17855]_ , \new_[17859]_ , \new_[17860]_ , \new_[17861]_ ,
    \new_[17865]_ , \new_[17866]_ , \new_[17869]_ , \new_[17872]_ ,
    \new_[17873]_ , \new_[17874]_ , \new_[17878]_ , \new_[17879]_ ,
    \new_[17883]_ , \new_[17884]_ , \new_[17885]_ , \new_[17889]_ ,
    \new_[17890]_ , \new_[17893]_ , \new_[17896]_ , \new_[17897]_ ,
    \new_[17898]_ , \new_[17902]_ , \new_[17903]_ , \new_[17907]_ ,
    \new_[17908]_ , \new_[17909]_ , \new_[17913]_ , \new_[17914]_ ,
    \new_[17917]_ , \new_[17920]_ , \new_[17921]_ , \new_[17922]_ ,
    \new_[17926]_ , \new_[17927]_ , \new_[17931]_ , \new_[17932]_ ,
    \new_[17933]_ , \new_[17937]_ , \new_[17938]_ , \new_[17941]_ ,
    \new_[17944]_ , \new_[17945]_ , \new_[17946]_ , \new_[17950]_ ,
    \new_[17951]_ , \new_[17955]_ , \new_[17956]_ , \new_[17957]_ ,
    \new_[17961]_ , \new_[17962]_ , \new_[17965]_ , \new_[17968]_ ,
    \new_[17969]_ , \new_[17970]_ , \new_[17974]_ , \new_[17975]_ ,
    \new_[17979]_ , \new_[17980]_ , \new_[17981]_ , \new_[17985]_ ,
    \new_[17986]_ , \new_[17989]_ , \new_[17992]_ , \new_[17993]_ ,
    \new_[17994]_ , \new_[17998]_ , \new_[17999]_ , \new_[18003]_ ,
    \new_[18004]_ , \new_[18005]_ , \new_[18009]_ , \new_[18010]_ ,
    \new_[18013]_ , \new_[18016]_ , \new_[18017]_ , \new_[18018]_ ,
    \new_[18022]_ , \new_[18023]_ , \new_[18027]_ , \new_[18028]_ ,
    \new_[18029]_ , \new_[18033]_ , \new_[18034]_ , \new_[18037]_ ,
    \new_[18040]_ , \new_[18041]_ , \new_[18042]_ , \new_[18046]_ ,
    \new_[18047]_ , \new_[18051]_ , \new_[18052]_ , \new_[18053]_ ,
    \new_[18057]_ , \new_[18058]_ , \new_[18061]_ , \new_[18064]_ ,
    \new_[18065]_ , \new_[18066]_ , \new_[18070]_ , \new_[18071]_ ,
    \new_[18075]_ , \new_[18076]_ , \new_[18077]_ , \new_[18081]_ ,
    \new_[18082]_ , \new_[18085]_ , \new_[18088]_ , \new_[18089]_ ,
    \new_[18090]_ , \new_[18094]_ , \new_[18095]_ , \new_[18099]_ ,
    \new_[18100]_ , \new_[18101]_ , \new_[18105]_ , \new_[18106]_ ,
    \new_[18109]_ , \new_[18112]_ , \new_[18113]_ , \new_[18114]_ ,
    \new_[18118]_ , \new_[18119]_ , \new_[18123]_ , \new_[18124]_ ,
    \new_[18125]_ , \new_[18129]_ , \new_[18130]_ , \new_[18133]_ ,
    \new_[18136]_ , \new_[18137]_ , \new_[18138]_ , \new_[18142]_ ,
    \new_[18143]_ , \new_[18147]_ , \new_[18148]_ , \new_[18149]_ ,
    \new_[18153]_ , \new_[18154]_ , \new_[18157]_ , \new_[18160]_ ,
    \new_[18161]_ , \new_[18162]_ , \new_[18166]_ , \new_[18167]_ ,
    \new_[18171]_ , \new_[18172]_ , \new_[18173]_ , \new_[18177]_ ,
    \new_[18178]_ , \new_[18181]_ , \new_[18184]_ , \new_[18185]_ ,
    \new_[18186]_ , \new_[18190]_ , \new_[18191]_ , \new_[18195]_ ,
    \new_[18196]_ , \new_[18197]_ , \new_[18201]_ , \new_[18202]_ ,
    \new_[18205]_ , \new_[18208]_ , \new_[18209]_ , \new_[18210]_ ,
    \new_[18214]_ , \new_[18215]_ , \new_[18219]_ , \new_[18220]_ ,
    \new_[18221]_ , \new_[18225]_ , \new_[18226]_ , \new_[18229]_ ,
    \new_[18232]_ , \new_[18233]_ , \new_[18234]_ , \new_[18238]_ ,
    \new_[18239]_ , \new_[18243]_ , \new_[18244]_ , \new_[18245]_ ,
    \new_[18249]_ , \new_[18250]_ , \new_[18253]_ , \new_[18256]_ ,
    \new_[18257]_ , \new_[18258]_ , \new_[18262]_ , \new_[18263]_ ,
    \new_[18267]_ , \new_[18268]_ , \new_[18269]_ , \new_[18273]_ ,
    \new_[18274]_ , \new_[18277]_ , \new_[18280]_ , \new_[18281]_ ,
    \new_[18282]_ , \new_[18286]_ , \new_[18287]_ , \new_[18291]_ ,
    \new_[18292]_ , \new_[18293]_ , \new_[18297]_ , \new_[18298]_ ,
    \new_[18301]_ , \new_[18304]_ , \new_[18305]_ , \new_[18306]_ ,
    \new_[18310]_ , \new_[18311]_ , \new_[18315]_ , \new_[18316]_ ,
    \new_[18317]_ , \new_[18321]_ , \new_[18322]_ , \new_[18325]_ ,
    \new_[18328]_ , \new_[18329]_ , \new_[18330]_ , \new_[18334]_ ,
    \new_[18335]_ , \new_[18339]_ , \new_[18340]_ , \new_[18341]_ ,
    \new_[18345]_ , \new_[18346]_ , \new_[18349]_ , \new_[18352]_ ,
    \new_[18353]_ , \new_[18354]_ , \new_[18358]_ , \new_[18359]_ ,
    \new_[18363]_ , \new_[18364]_ , \new_[18365]_ , \new_[18369]_ ,
    \new_[18370]_ , \new_[18373]_ , \new_[18376]_ , \new_[18377]_ ,
    \new_[18378]_ , \new_[18382]_ , \new_[18383]_ , \new_[18387]_ ,
    \new_[18388]_ , \new_[18389]_ , \new_[18393]_ , \new_[18394]_ ,
    \new_[18397]_ , \new_[18400]_ , \new_[18401]_ , \new_[18402]_ ,
    \new_[18406]_ , \new_[18407]_ , \new_[18411]_ , \new_[18412]_ ,
    \new_[18413]_ , \new_[18417]_ , \new_[18418]_ , \new_[18421]_ ,
    \new_[18424]_ , \new_[18425]_ , \new_[18426]_ , \new_[18430]_ ,
    \new_[18431]_ , \new_[18435]_ , \new_[18436]_ , \new_[18437]_ ,
    \new_[18441]_ , \new_[18442]_ , \new_[18445]_ , \new_[18448]_ ,
    \new_[18449]_ , \new_[18450]_ , \new_[18454]_ , \new_[18455]_ ,
    \new_[18459]_ , \new_[18460]_ , \new_[18461]_ , \new_[18465]_ ,
    \new_[18466]_ , \new_[18469]_ , \new_[18472]_ , \new_[18473]_ ,
    \new_[18474]_ , \new_[18478]_ , \new_[18479]_ , \new_[18483]_ ,
    \new_[18484]_ , \new_[18485]_ , \new_[18489]_ , \new_[18490]_ ,
    \new_[18493]_ , \new_[18496]_ , \new_[18497]_ , \new_[18498]_ ,
    \new_[18502]_ , \new_[18503]_ , \new_[18507]_ , \new_[18508]_ ,
    \new_[18509]_ , \new_[18513]_ , \new_[18514]_ , \new_[18517]_ ,
    \new_[18520]_ , \new_[18521]_ , \new_[18522]_ , \new_[18526]_ ,
    \new_[18527]_ , \new_[18531]_ , \new_[18532]_ , \new_[18533]_ ,
    \new_[18537]_ , \new_[18538]_ , \new_[18541]_ , \new_[18544]_ ,
    \new_[18545]_ , \new_[18546]_ , \new_[18550]_ , \new_[18551]_ ,
    \new_[18555]_ , \new_[18556]_ , \new_[18557]_ , \new_[18561]_ ,
    \new_[18562]_ , \new_[18565]_ , \new_[18568]_ , \new_[18569]_ ,
    \new_[18570]_ , \new_[18574]_ , \new_[18575]_ , \new_[18579]_ ,
    \new_[18580]_ , \new_[18581]_ , \new_[18585]_ , \new_[18586]_ ,
    \new_[18589]_ , \new_[18592]_ , \new_[18593]_ , \new_[18594]_ ,
    \new_[18598]_ , \new_[18599]_ , \new_[18603]_ , \new_[18604]_ ,
    \new_[18605]_ , \new_[18609]_ , \new_[18610]_ , \new_[18613]_ ,
    \new_[18616]_ , \new_[18617]_ , \new_[18618]_ , \new_[18622]_ ,
    \new_[18623]_ , \new_[18627]_ , \new_[18628]_ , \new_[18629]_ ,
    \new_[18633]_ , \new_[18634]_ , \new_[18637]_ , \new_[18640]_ ,
    \new_[18641]_ , \new_[18642]_ , \new_[18646]_ , \new_[18647]_ ,
    \new_[18651]_ , \new_[18652]_ , \new_[18653]_ , \new_[18657]_ ,
    \new_[18658]_ , \new_[18661]_ , \new_[18664]_ , \new_[18665]_ ,
    \new_[18666]_ , \new_[18670]_ , \new_[18671]_ , \new_[18675]_ ,
    \new_[18676]_ , \new_[18677]_ , \new_[18681]_ , \new_[18682]_ ,
    \new_[18685]_ , \new_[18688]_ , \new_[18689]_ , \new_[18690]_ ,
    \new_[18694]_ , \new_[18695]_ , \new_[18699]_ , \new_[18700]_ ,
    \new_[18701]_ , \new_[18705]_ , \new_[18706]_ , \new_[18709]_ ,
    \new_[18712]_ , \new_[18713]_ , \new_[18714]_ , \new_[18718]_ ,
    \new_[18719]_ , \new_[18723]_ , \new_[18724]_ , \new_[18725]_ ,
    \new_[18729]_ , \new_[18730]_ , \new_[18733]_ , \new_[18736]_ ,
    \new_[18737]_ , \new_[18738]_ , \new_[18742]_ , \new_[18743]_ ,
    \new_[18747]_ , \new_[18748]_ , \new_[18749]_ , \new_[18753]_ ,
    \new_[18754]_ , \new_[18757]_ , \new_[18760]_ , \new_[18761]_ ,
    \new_[18762]_ , \new_[18766]_ , \new_[18767]_ , \new_[18771]_ ,
    \new_[18772]_ , \new_[18773]_ , \new_[18777]_ , \new_[18778]_ ,
    \new_[18781]_ , \new_[18784]_ , \new_[18785]_ , \new_[18786]_ ,
    \new_[18790]_ , \new_[18791]_ , \new_[18795]_ , \new_[18796]_ ,
    \new_[18797]_ , \new_[18801]_ , \new_[18802]_ , \new_[18805]_ ,
    \new_[18808]_ , \new_[18809]_ , \new_[18810]_ , \new_[18814]_ ,
    \new_[18815]_ , \new_[18819]_ , \new_[18820]_ , \new_[18821]_ ,
    \new_[18825]_ , \new_[18826]_ , \new_[18829]_ , \new_[18832]_ ,
    \new_[18833]_ , \new_[18834]_ , \new_[18838]_ , \new_[18839]_ ,
    \new_[18843]_ , \new_[18844]_ , \new_[18845]_ , \new_[18849]_ ,
    \new_[18850]_ , \new_[18853]_ , \new_[18856]_ , \new_[18857]_ ,
    \new_[18858]_ , \new_[18862]_ , \new_[18863]_ , \new_[18867]_ ,
    \new_[18868]_ , \new_[18869]_ , \new_[18873]_ , \new_[18874]_ ,
    \new_[18877]_ , \new_[18880]_ , \new_[18881]_ , \new_[18882]_ ,
    \new_[18886]_ , \new_[18887]_ , \new_[18891]_ , \new_[18892]_ ,
    \new_[18893]_ , \new_[18897]_ , \new_[18898]_ , \new_[18901]_ ,
    \new_[18904]_ , \new_[18905]_ , \new_[18906]_ , \new_[18910]_ ,
    \new_[18911]_ , \new_[18915]_ , \new_[18916]_ , \new_[18917]_ ,
    \new_[18921]_ , \new_[18922]_ , \new_[18925]_ , \new_[18928]_ ,
    \new_[18929]_ , \new_[18930]_ , \new_[18934]_ , \new_[18935]_ ,
    \new_[18939]_ , \new_[18940]_ , \new_[18941]_ , \new_[18945]_ ,
    \new_[18946]_ , \new_[18949]_ , \new_[18952]_ , \new_[18953]_ ,
    \new_[18954]_ , \new_[18958]_ , \new_[18959]_ , \new_[18963]_ ,
    \new_[18964]_ , \new_[18965]_ , \new_[18969]_ , \new_[18970]_ ,
    \new_[18973]_ , \new_[18976]_ , \new_[18977]_ , \new_[18978]_ ,
    \new_[18982]_ , \new_[18983]_ , \new_[18987]_ , \new_[18988]_ ,
    \new_[18989]_ , \new_[18993]_ , \new_[18994]_ , \new_[18997]_ ,
    \new_[19000]_ , \new_[19001]_ , \new_[19002]_ , \new_[19006]_ ,
    \new_[19007]_ , \new_[19011]_ , \new_[19012]_ , \new_[19013]_ ,
    \new_[19017]_ , \new_[19018]_ , \new_[19021]_ , \new_[19024]_ ,
    \new_[19025]_ , \new_[19026]_ , \new_[19030]_ , \new_[19031]_ ,
    \new_[19035]_ , \new_[19036]_ , \new_[19037]_ , \new_[19041]_ ,
    \new_[19042]_ , \new_[19045]_ , \new_[19048]_ , \new_[19049]_ ,
    \new_[19050]_ , \new_[19054]_ , \new_[19055]_ , \new_[19059]_ ,
    \new_[19060]_ , \new_[19061]_ , \new_[19065]_ , \new_[19066]_ ,
    \new_[19069]_ , \new_[19072]_ , \new_[19073]_ , \new_[19074]_ ,
    \new_[19078]_ , \new_[19079]_ , \new_[19083]_ , \new_[19084]_ ,
    \new_[19085]_ , \new_[19089]_ , \new_[19090]_ , \new_[19093]_ ,
    \new_[19096]_ , \new_[19097]_ , \new_[19098]_ , \new_[19102]_ ,
    \new_[19103]_ , \new_[19107]_ , \new_[19108]_ , \new_[19109]_ ,
    \new_[19113]_ , \new_[19114]_ , \new_[19117]_ , \new_[19120]_ ,
    \new_[19121]_ , \new_[19122]_ , \new_[19126]_ , \new_[19127]_ ,
    \new_[19131]_ , \new_[19132]_ , \new_[19133]_ , \new_[19137]_ ,
    \new_[19138]_ , \new_[19141]_ , \new_[19144]_ , \new_[19145]_ ,
    \new_[19146]_ , \new_[19150]_ , \new_[19151]_ , \new_[19155]_ ,
    \new_[19156]_ , \new_[19157]_ , \new_[19161]_ , \new_[19162]_ ,
    \new_[19165]_ , \new_[19168]_ , \new_[19169]_ , \new_[19170]_ ,
    \new_[19174]_ , \new_[19175]_ , \new_[19179]_ , \new_[19180]_ ,
    \new_[19181]_ , \new_[19185]_ , \new_[19186]_ , \new_[19189]_ ,
    \new_[19192]_ , \new_[19193]_ , \new_[19194]_ , \new_[19198]_ ,
    \new_[19199]_ , \new_[19203]_ , \new_[19204]_ , \new_[19205]_ ,
    \new_[19209]_ , \new_[19210]_ , \new_[19213]_ , \new_[19216]_ ,
    \new_[19217]_ , \new_[19218]_ , \new_[19222]_ , \new_[19223]_ ,
    \new_[19227]_ , \new_[19228]_ , \new_[19229]_ , \new_[19233]_ ,
    \new_[19234]_ , \new_[19237]_ , \new_[19240]_ , \new_[19241]_ ,
    \new_[19242]_ , \new_[19246]_ , \new_[19247]_ , \new_[19251]_ ,
    \new_[19252]_ , \new_[19253]_ , \new_[19257]_ , \new_[19258]_ ,
    \new_[19261]_ , \new_[19264]_ , \new_[19265]_ , \new_[19266]_ ,
    \new_[19270]_ , \new_[19271]_ , \new_[19275]_ , \new_[19276]_ ,
    \new_[19277]_ , \new_[19281]_ , \new_[19282]_ , \new_[19285]_ ,
    \new_[19288]_ , \new_[19289]_ , \new_[19290]_ , \new_[19294]_ ,
    \new_[19295]_ , \new_[19299]_ , \new_[19300]_ , \new_[19301]_ ,
    \new_[19305]_ , \new_[19306]_ , \new_[19309]_ , \new_[19312]_ ,
    \new_[19313]_ , \new_[19314]_ , \new_[19318]_ , \new_[19319]_ ,
    \new_[19323]_ , \new_[19324]_ , \new_[19325]_ , \new_[19329]_ ,
    \new_[19330]_ , \new_[19333]_ , \new_[19336]_ , \new_[19337]_ ,
    \new_[19338]_ , \new_[19342]_ , \new_[19343]_ , \new_[19347]_ ,
    \new_[19348]_ , \new_[19349]_ , \new_[19353]_ , \new_[19354]_ ,
    \new_[19357]_ , \new_[19360]_ , \new_[19361]_ , \new_[19362]_ ,
    \new_[19366]_ , \new_[19367]_ , \new_[19371]_ , \new_[19372]_ ,
    \new_[19373]_ , \new_[19377]_ , \new_[19378]_ , \new_[19381]_ ,
    \new_[19384]_ , \new_[19385]_ , \new_[19386]_ , \new_[19390]_ ,
    \new_[19391]_ , \new_[19395]_ , \new_[19396]_ , \new_[19397]_ ,
    \new_[19401]_ , \new_[19402]_ , \new_[19405]_ , \new_[19408]_ ,
    \new_[19409]_ , \new_[19410]_ , \new_[19414]_ , \new_[19415]_ ,
    \new_[19419]_ , \new_[19420]_ , \new_[19421]_ , \new_[19425]_ ,
    \new_[19426]_ , \new_[19429]_ , \new_[19432]_ , \new_[19433]_ ,
    \new_[19434]_ , \new_[19438]_ , \new_[19439]_ , \new_[19443]_ ,
    \new_[19444]_ , \new_[19445]_ , \new_[19449]_ , \new_[19450]_ ,
    \new_[19453]_ , \new_[19456]_ , \new_[19457]_ , \new_[19458]_ ,
    \new_[19462]_ , \new_[19463]_ , \new_[19466]_ , \new_[19469]_ ,
    \new_[19470]_ , \new_[19471]_ , \new_[19475]_ , \new_[19476]_ ,
    \new_[19479]_ , \new_[19482]_ , \new_[19483]_ , \new_[19484]_ ,
    \new_[19488]_ , \new_[19489]_ , \new_[19492]_ , \new_[19495]_ ,
    \new_[19496]_ , \new_[19497]_ , \new_[19501]_ , \new_[19502]_ ,
    \new_[19505]_ , \new_[19508]_ , \new_[19509]_ , \new_[19510]_ ,
    \new_[19514]_ , \new_[19515]_ , \new_[19518]_ , \new_[19521]_ ,
    \new_[19522]_ , \new_[19523]_ , \new_[19527]_ , \new_[19528]_ ,
    \new_[19531]_ , \new_[19534]_ , \new_[19535]_ , \new_[19536]_ ,
    \new_[19540]_ , \new_[19541]_ , \new_[19544]_ , \new_[19547]_ ,
    \new_[19548]_ , \new_[19549]_ , \new_[19553]_ , \new_[19554]_ ,
    \new_[19557]_ , \new_[19560]_ , \new_[19561]_ , \new_[19562]_ ,
    \new_[19566]_ , \new_[19567]_ , \new_[19570]_ , \new_[19573]_ ,
    \new_[19574]_ , \new_[19575]_ , \new_[19579]_ , \new_[19580]_ ,
    \new_[19583]_ , \new_[19586]_ , \new_[19587]_ , \new_[19588]_ ,
    \new_[19592]_ , \new_[19593]_ , \new_[19596]_ , \new_[19599]_ ,
    \new_[19600]_ , \new_[19601]_ , \new_[19605]_ , \new_[19606]_ ,
    \new_[19609]_ , \new_[19612]_ , \new_[19613]_ , \new_[19614]_ ,
    \new_[19618]_ , \new_[19619]_ , \new_[19622]_ , \new_[19625]_ ,
    \new_[19626]_ , \new_[19627]_ , \new_[19631]_ , \new_[19632]_ ,
    \new_[19635]_ , \new_[19638]_ , \new_[19639]_ , \new_[19640]_ ,
    \new_[19644]_ , \new_[19645]_ , \new_[19648]_ , \new_[19651]_ ,
    \new_[19652]_ , \new_[19653]_ , \new_[19657]_ , \new_[19658]_ ,
    \new_[19661]_ , \new_[19664]_ , \new_[19665]_ , \new_[19666]_ ,
    \new_[19670]_ , \new_[19671]_ , \new_[19674]_ , \new_[19677]_ ,
    \new_[19678]_ , \new_[19679]_ , \new_[19683]_ , \new_[19684]_ ,
    \new_[19687]_ , \new_[19690]_ , \new_[19691]_ , \new_[19692]_ ,
    \new_[19696]_ , \new_[19697]_ , \new_[19700]_ , \new_[19703]_ ,
    \new_[19704]_ , \new_[19705]_ , \new_[19709]_ , \new_[19710]_ ,
    \new_[19713]_ , \new_[19716]_ , \new_[19717]_ , \new_[19718]_ ,
    \new_[19722]_ , \new_[19723]_ , \new_[19726]_ , \new_[19729]_ ,
    \new_[19730]_ , \new_[19731]_ , \new_[19735]_ , \new_[19736]_ ,
    \new_[19739]_ , \new_[19742]_ , \new_[19743]_ , \new_[19744]_ ,
    \new_[19748]_ , \new_[19749]_ , \new_[19752]_ , \new_[19755]_ ,
    \new_[19756]_ , \new_[19757]_ , \new_[19761]_ , \new_[19762]_ ,
    \new_[19765]_ , \new_[19768]_ , \new_[19769]_ , \new_[19770]_ ,
    \new_[19774]_ , \new_[19775]_ , \new_[19778]_ , \new_[19781]_ ,
    \new_[19782]_ , \new_[19783]_ , \new_[19787]_ , \new_[19788]_ ,
    \new_[19791]_ , \new_[19794]_ , \new_[19795]_ , \new_[19796]_ ,
    \new_[19800]_ , \new_[19801]_ , \new_[19804]_ , \new_[19807]_ ,
    \new_[19808]_ , \new_[19809]_ , \new_[19813]_ , \new_[19814]_ ,
    \new_[19817]_ , \new_[19820]_ , \new_[19821]_ , \new_[19822]_ ,
    \new_[19826]_ , \new_[19827]_ , \new_[19830]_ , \new_[19833]_ ,
    \new_[19834]_ , \new_[19835]_ , \new_[19839]_ , \new_[19840]_ ,
    \new_[19843]_ , \new_[19846]_ , \new_[19847]_ , \new_[19848]_ ,
    \new_[19852]_ , \new_[19853]_ , \new_[19856]_ , \new_[19859]_ ,
    \new_[19860]_ , \new_[19861]_ , \new_[19865]_ , \new_[19866]_ ,
    \new_[19869]_ , \new_[19872]_ , \new_[19873]_ , \new_[19874]_ ,
    \new_[19878]_ , \new_[19879]_ , \new_[19882]_ , \new_[19885]_ ,
    \new_[19886]_ , \new_[19887]_ , \new_[19891]_ , \new_[19892]_ ,
    \new_[19895]_ , \new_[19898]_ , \new_[19899]_ , \new_[19900]_ ,
    \new_[19904]_ , \new_[19905]_ , \new_[19908]_ , \new_[19911]_ ,
    \new_[19912]_ , \new_[19913]_ , \new_[19917]_ , \new_[19918]_ ,
    \new_[19921]_ , \new_[19924]_ , \new_[19925]_ , \new_[19926]_ ,
    \new_[19930]_ , \new_[19931]_ , \new_[19934]_ , \new_[19937]_ ,
    \new_[19938]_ , \new_[19939]_ , \new_[19943]_ , \new_[19944]_ ,
    \new_[19947]_ , \new_[19950]_ , \new_[19951]_ , \new_[19952]_ ,
    \new_[19956]_ , \new_[19957]_ , \new_[19960]_ , \new_[19963]_ ,
    \new_[19964]_ , \new_[19965]_ , \new_[19969]_ , \new_[19970]_ ,
    \new_[19973]_ , \new_[19976]_ , \new_[19977]_ , \new_[19978]_ ,
    \new_[19982]_ , \new_[19983]_ , \new_[19986]_ , \new_[19989]_ ,
    \new_[19990]_ , \new_[19991]_ , \new_[19995]_ , \new_[19996]_ ,
    \new_[19999]_ , \new_[20002]_ , \new_[20003]_ , \new_[20004]_ ,
    \new_[20008]_ , \new_[20009]_ , \new_[20012]_ , \new_[20015]_ ,
    \new_[20016]_ , \new_[20017]_ , \new_[20021]_ , \new_[20022]_ ,
    \new_[20025]_ , \new_[20028]_ , \new_[20029]_ , \new_[20030]_ ,
    \new_[20034]_ , \new_[20035]_ , \new_[20038]_ , \new_[20041]_ ,
    \new_[20042]_ , \new_[20043]_ , \new_[20047]_ , \new_[20048]_ ,
    \new_[20051]_ , \new_[20054]_ , \new_[20055]_ , \new_[20056]_ ,
    \new_[20060]_ , \new_[20061]_ , \new_[20064]_ , \new_[20067]_ ,
    \new_[20068]_ , \new_[20069]_ , \new_[20073]_ , \new_[20074]_ ,
    \new_[20077]_ , \new_[20080]_ , \new_[20081]_ , \new_[20082]_ ,
    \new_[20086]_ , \new_[20087]_ , \new_[20090]_ , \new_[20093]_ ,
    \new_[20094]_ , \new_[20095]_ , \new_[20099]_ , \new_[20100]_ ,
    \new_[20103]_ , \new_[20106]_ , \new_[20107]_ , \new_[20108]_ ,
    \new_[20112]_ , \new_[20113]_ , \new_[20116]_ , \new_[20119]_ ,
    \new_[20120]_ , \new_[20121]_ , \new_[20125]_ , \new_[20126]_ ,
    \new_[20129]_ , \new_[20132]_ , \new_[20133]_ , \new_[20134]_ ,
    \new_[20138]_ , \new_[20139]_ , \new_[20142]_ , \new_[20145]_ ,
    \new_[20146]_ , \new_[20147]_ , \new_[20151]_ , \new_[20152]_ ,
    \new_[20155]_ , \new_[20158]_ , \new_[20159]_ , \new_[20160]_ ,
    \new_[20164]_ , \new_[20165]_ , \new_[20168]_ , \new_[20171]_ ,
    \new_[20172]_ , \new_[20173]_ , \new_[20177]_ , \new_[20178]_ ,
    \new_[20181]_ , \new_[20184]_ , \new_[20185]_ , \new_[20186]_ ,
    \new_[20190]_ , \new_[20191]_ , \new_[20194]_ , \new_[20197]_ ,
    \new_[20198]_ , \new_[20199]_ , \new_[20203]_ , \new_[20204]_ ,
    \new_[20207]_ , \new_[20210]_ , \new_[20211]_ , \new_[20212]_ ,
    \new_[20216]_ , \new_[20217]_ , \new_[20220]_ , \new_[20223]_ ,
    \new_[20224]_ , \new_[20225]_ , \new_[20229]_ , \new_[20230]_ ,
    \new_[20233]_ , \new_[20236]_ , \new_[20237]_ , \new_[20238]_ ,
    \new_[20242]_ , \new_[20243]_ , \new_[20246]_ , \new_[20249]_ ,
    \new_[20250]_ , \new_[20251]_ , \new_[20255]_ , \new_[20256]_ ,
    \new_[20259]_ , \new_[20262]_ , \new_[20263]_ , \new_[20264]_ ,
    \new_[20268]_ , \new_[20269]_ , \new_[20272]_ , \new_[20275]_ ,
    \new_[20276]_ , \new_[20277]_ , \new_[20281]_ , \new_[20282]_ ,
    \new_[20285]_ , \new_[20288]_ , \new_[20289]_ , \new_[20290]_ ,
    \new_[20294]_ , \new_[20295]_ , \new_[20298]_ , \new_[20301]_ ,
    \new_[20302]_ , \new_[20303]_ , \new_[20307]_ , \new_[20308]_ ,
    \new_[20311]_ , \new_[20314]_ , \new_[20315]_ , \new_[20316]_ ,
    \new_[20320]_ , \new_[20321]_ , \new_[20324]_ , \new_[20327]_ ,
    \new_[20328]_ , \new_[20329]_ , \new_[20333]_ , \new_[20334]_ ,
    \new_[20337]_ , \new_[20340]_ , \new_[20341]_ , \new_[20342]_ ,
    \new_[20346]_ , \new_[20347]_ , \new_[20350]_ , \new_[20353]_ ,
    \new_[20354]_ , \new_[20355]_ , \new_[20359]_ , \new_[20360]_ ,
    \new_[20363]_ , \new_[20366]_ , \new_[20367]_ , \new_[20368]_ ,
    \new_[20372]_ , \new_[20373]_ , \new_[20376]_ , \new_[20379]_ ,
    \new_[20380]_ , \new_[20381]_ , \new_[20385]_ , \new_[20386]_ ,
    \new_[20389]_ , \new_[20392]_ , \new_[20393]_ , \new_[20394]_ ,
    \new_[20398]_ , \new_[20399]_ , \new_[20402]_ , \new_[20405]_ ,
    \new_[20406]_ , \new_[20407]_ , \new_[20411]_ , \new_[20412]_ ,
    \new_[20415]_ , \new_[20418]_ , \new_[20419]_ , \new_[20420]_ ,
    \new_[20424]_ , \new_[20425]_ , \new_[20428]_ , \new_[20431]_ ,
    \new_[20432]_ , \new_[20433]_ , \new_[20437]_ , \new_[20438]_ ,
    \new_[20441]_ , \new_[20444]_ , \new_[20445]_ , \new_[20446]_ ,
    \new_[20450]_ , \new_[20451]_ , \new_[20454]_ , \new_[20457]_ ,
    \new_[20458]_ , \new_[20459]_ , \new_[20463]_ , \new_[20464]_ ,
    \new_[20467]_ , \new_[20470]_ , \new_[20471]_ , \new_[20472]_ ,
    \new_[20476]_ , \new_[20477]_ , \new_[20480]_ , \new_[20483]_ ,
    \new_[20484]_ , \new_[20485]_ , \new_[20489]_ , \new_[20490]_ ,
    \new_[20493]_ , \new_[20496]_ , \new_[20497]_ , \new_[20498]_ ,
    \new_[20502]_ , \new_[20503]_ , \new_[20506]_ , \new_[20509]_ ,
    \new_[20510]_ , \new_[20511]_ , \new_[20515]_ , \new_[20516]_ ,
    \new_[20519]_ , \new_[20522]_ , \new_[20523]_ , \new_[20524]_ ,
    \new_[20528]_ , \new_[20529]_ , \new_[20532]_ , \new_[20535]_ ,
    \new_[20536]_ , \new_[20537]_ , \new_[20541]_ , \new_[20542]_ ,
    \new_[20545]_ , \new_[20548]_ , \new_[20549]_ , \new_[20550]_ ,
    \new_[20554]_ , \new_[20555]_ , \new_[20558]_ , \new_[20561]_ ,
    \new_[20562]_ , \new_[20563]_ , \new_[20567]_ , \new_[20568]_ ,
    \new_[20571]_ , \new_[20574]_ , \new_[20575]_ , \new_[20576]_ ,
    \new_[20580]_ , \new_[20581]_ , \new_[20584]_ , \new_[20587]_ ,
    \new_[20588]_ , \new_[20589]_ , \new_[20593]_ , \new_[20594]_ ,
    \new_[20597]_ , \new_[20600]_ , \new_[20601]_ , \new_[20602]_ ,
    \new_[20606]_ , \new_[20607]_ , \new_[20610]_ , \new_[20613]_ ,
    \new_[20614]_ , \new_[20615]_ , \new_[20619]_ , \new_[20620]_ ,
    \new_[20623]_ , \new_[20626]_ , \new_[20627]_ , \new_[20628]_ ,
    \new_[20632]_ , \new_[20633]_ , \new_[20636]_ , \new_[20639]_ ,
    \new_[20640]_ , \new_[20641]_ , \new_[20645]_ , \new_[20646]_ ,
    \new_[20649]_ , \new_[20652]_ , \new_[20653]_ , \new_[20654]_ ,
    \new_[20658]_ , \new_[20659]_ , \new_[20662]_ , \new_[20665]_ ,
    \new_[20666]_ , \new_[20667]_ , \new_[20671]_ , \new_[20672]_ ,
    \new_[20675]_ , \new_[20678]_ , \new_[20679]_ , \new_[20680]_ ,
    \new_[20684]_ , \new_[20685]_ , \new_[20688]_ , \new_[20691]_ ,
    \new_[20692]_ , \new_[20693]_ , \new_[20697]_ , \new_[20698]_ ,
    \new_[20701]_ , \new_[20704]_ , \new_[20705]_ , \new_[20706]_ ,
    \new_[20710]_ , \new_[20711]_ , \new_[20714]_ , \new_[20717]_ ,
    \new_[20718]_ , \new_[20719]_ , \new_[20723]_ , \new_[20724]_ ,
    \new_[20727]_ , \new_[20730]_ , \new_[20731]_ , \new_[20732]_ ,
    \new_[20736]_ , \new_[20737]_ , \new_[20740]_ , \new_[20743]_ ,
    \new_[20744]_ , \new_[20745]_ , \new_[20749]_ , \new_[20750]_ ,
    \new_[20753]_ , \new_[20756]_ , \new_[20757]_ , \new_[20758]_ ,
    \new_[20762]_ , \new_[20763]_ , \new_[20766]_ , \new_[20769]_ ,
    \new_[20770]_ , \new_[20771]_ , \new_[20775]_ , \new_[20776]_ ,
    \new_[20779]_ , \new_[20782]_ , \new_[20783]_ , \new_[20784]_ ,
    \new_[20788]_ , \new_[20789]_ , \new_[20792]_ , \new_[20795]_ ,
    \new_[20796]_ , \new_[20797]_ , \new_[20801]_ , \new_[20802]_ ,
    \new_[20805]_ , \new_[20808]_ , \new_[20809]_ , \new_[20810]_ ,
    \new_[20814]_ , \new_[20815]_ , \new_[20818]_ , \new_[20821]_ ,
    \new_[20822]_ , \new_[20823]_ , \new_[20827]_ , \new_[20828]_ ,
    \new_[20831]_ , \new_[20834]_ , \new_[20835]_ , \new_[20836]_ ,
    \new_[20840]_ , \new_[20841]_ , \new_[20844]_ , \new_[20847]_ ,
    \new_[20848]_ , \new_[20849]_ , \new_[20853]_ , \new_[20854]_ ,
    \new_[20857]_ , \new_[20860]_ , \new_[20861]_ , \new_[20862]_ ,
    \new_[20866]_ , \new_[20867]_ , \new_[20870]_ , \new_[20873]_ ,
    \new_[20874]_ , \new_[20875]_ , \new_[20879]_ , \new_[20880]_ ,
    \new_[20883]_ , \new_[20886]_ , \new_[20887]_ , \new_[20888]_ ,
    \new_[20892]_ , \new_[20893]_ , \new_[20896]_ , \new_[20899]_ ,
    \new_[20900]_ , \new_[20901]_ , \new_[20905]_ , \new_[20906]_ ,
    \new_[20909]_ , \new_[20912]_ , \new_[20913]_ , \new_[20914]_ ,
    \new_[20918]_ , \new_[20919]_ , \new_[20922]_ , \new_[20925]_ ,
    \new_[20926]_ , \new_[20927]_ , \new_[20931]_ , \new_[20932]_ ,
    \new_[20935]_ , \new_[20938]_ , \new_[20939]_ , \new_[20940]_ ,
    \new_[20944]_ , \new_[20945]_ , \new_[20948]_ , \new_[20951]_ ,
    \new_[20952]_ , \new_[20953]_ , \new_[20957]_ , \new_[20958]_ ,
    \new_[20961]_ , \new_[20964]_ , \new_[20965]_ , \new_[20966]_ ,
    \new_[20970]_ , \new_[20971]_ , \new_[20974]_ , \new_[20977]_ ,
    \new_[20978]_ , \new_[20979]_ , \new_[20983]_ , \new_[20984]_ ,
    \new_[20987]_ , \new_[20990]_ , \new_[20991]_ , \new_[20992]_ ,
    \new_[20996]_ , \new_[20997]_ , \new_[21000]_ , \new_[21003]_ ,
    \new_[21004]_ , \new_[21005]_ , \new_[21009]_ , \new_[21010]_ ,
    \new_[21013]_ , \new_[21016]_ , \new_[21017]_ , \new_[21018]_ ,
    \new_[21022]_ , \new_[21023]_ , \new_[21026]_ , \new_[21029]_ ,
    \new_[21030]_ , \new_[21031]_ , \new_[21035]_ , \new_[21036]_ ,
    \new_[21039]_ , \new_[21042]_ , \new_[21043]_ , \new_[21044]_ ,
    \new_[21048]_ , \new_[21049]_ , \new_[21052]_ , \new_[21055]_ ,
    \new_[21056]_ , \new_[21057]_ , \new_[21061]_ , \new_[21062]_ ,
    \new_[21065]_ , \new_[21068]_ , \new_[21069]_ , \new_[21070]_ ,
    \new_[21074]_ , \new_[21075]_ , \new_[21078]_ , \new_[21081]_ ,
    \new_[21082]_ , \new_[21083]_ , \new_[21087]_ , \new_[21088]_ ,
    \new_[21091]_ , \new_[21094]_ , \new_[21095]_ , \new_[21096]_ ,
    \new_[21100]_ , \new_[21101]_ , \new_[21104]_ , \new_[21107]_ ,
    \new_[21108]_ , \new_[21109]_ , \new_[21113]_ , \new_[21114]_ ,
    \new_[21117]_ , \new_[21120]_ , \new_[21121]_ , \new_[21122]_ ,
    \new_[21126]_ , \new_[21127]_ , \new_[21130]_ , \new_[21133]_ ,
    \new_[21134]_ , \new_[21135]_ , \new_[21139]_ , \new_[21140]_ ,
    \new_[21143]_ , \new_[21146]_ , \new_[21147]_ , \new_[21148]_ ,
    \new_[21152]_ , \new_[21153]_ , \new_[21156]_ , \new_[21159]_ ,
    \new_[21160]_ , \new_[21161]_ , \new_[21165]_ , \new_[21166]_ ,
    \new_[21169]_ , \new_[21172]_ , \new_[21173]_ , \new_[21174]_ ,
    \new_[21178]_ , \new_[21179]_ , \new_[21182]_ , \new_[21185]_ ,
    \new_[21186]_ , \new_[21187]_ , \new_[21191]_ , \new_[21192]_ ,
    \new_[21195]_ , \new_[21198]_ , \new_[21199]_ , \new_[21200]_ ,
    \new_[21204]_ , \new_[21205]_ , \new_[21208]_ , \new_[21211]_ ,
    \new_[21212]_ , \new_[21213]_ , \new_[21217]_ , \new_[21218]_ ,
    \new_[21221]_ , \new_[21224]_ , \new_[21225]_ , \new_[21226]_ ,
    \new_[21230]_ , \new_[21231]_ , \new_[21234]_ , \new_[21237]_ ,
    \new_[21238]_ , \new_[21239]_ , \new_[21243]_ , \new_[21244]_ ,
    \new_[21247]_ , \new_[21250]_ , \new_[21251]_ , \new_[21252]_ ,
    \new_[21256]_ , \new_[21257]_ , \new_[21260]_ , \new_[21263]_ ,
    \new_[21264]_ , \new_[21265]_ , \new_[21269]_ , \new_[21270]_ ,
    \new_[21273]_ , \new_[21276]_ , \new_[21277]_ , \new_[21278]_ ,
    \new_[21282]_ , \new_[21283]_ , \new_[21286]_ , \new_[21289]_ ,
    \new_[21290]_ , \new_[21291]_ , \new_[21295]_ , \new_[21296]_ ,
    \new_[21299]_ , \new_[21302]_ , \new_[21303]_ , \new_[21304]_ ,
    \new_[21308]_ , \new_[21309]_ , \new_[21312]_ , \new_[21315]_ ,
    \new_[21316]_ , \new_[21317]_ , \new_[21321]_ , \new_[21322]_ ,
    \new_[21325]_ , \new_[21328]_ , \new_[21329]_ , \new_[21330]_ ,
    \new_[21334]_ , \new_[21335]_ , \new_[21338]_ , \new_[21341]_ ,
    \new_[21342]_ , \new_[21343]_ , \new_[21347]_ , \new_[21348]_ ,
    \new_[21351]_ , \new_[21354]_ , \new_[21355]_ , \new_[21356]_ ,
    \new_[21360]_ , \new_[21361]_ , \new_[21364]_ , \new_[21367]_ ,
    \new_[21368]_ , \new_[21369]_ , \new_[21373]_ , \new_[21374]_ ,
    \new_[21377]_ , \new_[21380]_ , \new_[21381]_ , \new_[21382]_ ,
    \new_[21386]_ , \new_[21387]_ , \new_[21390]_ , \new_[21393]_ ,
    \new_[21394]_ , \new_[21395]_ , \new_[21399]_ , \new_[21400]_ ,
    \new_[21403]_ , \new_[21406]_ , \new_[21407]_ , \new_[21408]_ ,
    \new_[21412]_ , \new_[21413]_ , \new_[21416]_ , \new_[21419]_ ,
    \new_[21420]_ , \new_[21421]_ , \new_[21425]_ , \new_[21426]_ ,
    \new_[21429]_ , \new_[21432]_ , \new_[21433]_ , \new_[21434]_ ,
    \new_[21438]_ , \new_[21439]_ , \new_[21442]_ , \new_[21445]_ ,
    \new_[21446]_ , \new_[21447]_ , \new_[21451]_ , \new_[21452]_ ,
    \new_[21455]_ , \new_[21458]_ , \new_[21459]_ , \new_[21460]_ ,
    \new_[21464]_ , \new_[21465]_ , \new_[21468]_ , \new_[21471]_ ,
    \new_[21472]_ , \new_[21473]_ , \new_[21477]_ , \new_[21478]_ ,
    \new_[21481]_ , \new_[21484]_ , \new_[21485]_ , \new_[21486]_ ,
    \new_[21490]_ , \new_[21491]_ , \new_[21494]_ , \new_[21497]_ ,
    \new_[21498]_ , \new_[21499]_ , \new_[21503]_ , \new_[21504]_ ,
    \new_[21507]_ , \new_[21510]_ , \new_[21511]_ , \new_[21512]_ ,
    \new_[21516]_ , \new_[21517]_ , \new_[21520]_ , \new_[21523]_ ,
    \new_[21524]_ , \new_[21525]_ , \new_[21529]_ , \new_[21530]_ ,
    \new_[21533]_ , \new_[21536]_ , \new_[21537]_ , \new_[21538]_ ,
    \new_[21542]_ , \new_[21543]_ , \new_[21546]_ , \new_[21549]_ ,
    \new_[21550]_ , \new_[21551]_ , \new_[21555]_ , \new_[21556]_ ,
    \new_[21559]_ , \new_[21562]_ , \new_[21563]_ , \new_[21564]_ ,
    \new_[21568]_ , \new_[21569]_ , \new_[21572]_ , \new_[21575]_ ,
    \new_[21576]_ , \new_[21577]_ , \new_[21581]_ , \new_[21582]_ ,
    \new_[21585]_ , \new_[21588]_ , \new_[21589]_ , \new_[21590]_ ,
    \new_[21594]_ , \new_[21595]_ , \new_[21598]_ , \new_[21601]_ ,
    \new_[21602]_ , \new_[21603]_ , \new_[21607]_ , \new_[21608]_ ,
    \new_[21611]_ , \new_[21614]_ , \new_[21615]_ , \new_[21616]_ ,
    \new_[21620]_ , \new_[21621]_ , \new_[21624]_ , \new_[21627]_ ,
    \new_[21628]_ , \new_[21629]_ , \new_[21633]_ , \new_[21634]_ ,
    \new_[21637]_ , \new_[21640]_ , \new_[21641]_ , \new_[21642]_ ,
    \new_[21646]_ , \new_[21647]_ , \new_[21650]_ , \new_[21653]_ ,
    \new_[21654]_ , \new_[21655]_ , \new_[21659]_ , \new_[21660]_ ,
    \new_[21663]_ , \new_[21666]_ , \new_[21667]_ , \new_[21668]_ ,
    \new_[21672]_ , \new_[21673]_ , \new_[21676]_ , \new_[21679]_ ,
    \new_[21680]_ , \new_[21681]_ , \new_[21685]_ , \new_[21686]_ ,
    \new_[21689]_ , \new_[21692]_ , \new_[21693]_ , \new_[21694]_ ,
    \new_[21698]_ , \new_[21699]_ , \new_[21702]_ , \new_[21705]_ ,
    \new_[21706]_ , \new_[21707]_ , \new_[21711]_ , \new_[21712]_ ,
    \new_[21715]_ , \new_[21718]_ , \new_[21719]_ , \new_[21720]_ ,
    \new_[21724]_ , \new_[21725]_ , \new_[21728]_ , \new_[21731]_ ,
    \new_[21732]_ , \new_[21733]_ , \new_[21737]_ , \new_[21738]_ ,
    \new_[21741]_ , \new_[21744]_ , \new_[21745]_ , \new_[21746]_ ,
    \new_[21750]_ , \new_[21751]_ , \new_[21754]_ , \new_[21757]_ ,
    \new_[21758]_ , \new_[21759]_ , \new_[21763]_ , \new_[21764]_ ,
    \new_[21767]_ , \new_[21770]_ , \new_[21771]_ , \new_[21772]_ ,
    \new_[21776]_ , \new_[21777]_ , \new_[21780]_ , \new_[21783]_ ,
    \new_[21784]_ , \new_[21785]_ , \new_[21789]_ , \new_[21790]_ ,
    \new_[21793]_ , \new_[21796]_ , \new_[21797]_ , \new_[21798]_ ,
    \new_[21802]_ , \new_[21803]_ , \new_[21806]_ , \new_[21809]_ ,
    \new_[21810]_ , \new_[21811]_ , \new_[21815]_ , \new_[21816]_ ,
    \new_[21819]_ , \new_[21822]_ , \new_[21823]_ , \new_[21824]_ ,
    \new_[21828]_ , \new_[21829]_ , \new_[21832]_ , \new_[21835]_ ,
    \new_[21836]_ , \new_[21837]_ , \new_[21841]_ , \new_[21842]_ ,
    \new_[21845]_ , \new_[21848]_ , \new_[21849]_ , \new_[21850]_ ,
    \new_[21854]_ , \new_[21855]_ , \new_[21858]_ , \new_[21861]_ ,
    \new_[21862]_ , \new_[21863]_ , \new_[21867]_ , \new_[21868]_ ,
    \new_[21871]_ , \new_[21874]_ , \new_[21875]_ , \new_[21876]_ ,
    \new_[21880]_ , \new_[21881]_ , \new_[21884]_ , \new_[21887]_ ,
    \new_[21888]_ , \new_[21889]_ , \new_[21893]_ , \new_[21894]_ ,
    \new_[21897]_ , \new_[21900]_ , \new_[21901]_ , \new_[21902]_ ,
    \new_[21906]_ , \new_[21907]_ , \new_[21910]_ , \new_[21913]_ ,
    \new_[21914]_ , \new_[21915]_ , \new_[21919]_ , \new_[21920]_ ,
    \new_[21923]_ , \new_[21926]_ , \new_[21927]_ , \new_[21928]_ ,
    \new_[21932]_ , \new_[21933]_ , \new_[21936]_ , \new_[21939]_ ,
    \new_[21940]_ , \new_[21941]_ , \new_[21945]_ , \new_[21946]_ ,
    \new_[21949]_ , \new_[21952]_ , \new_[21953]_ , \new_[21954]_ ,
    \new_[21958]_ , \new_[21959]_ , \new_[21962]_ , \new_[21965]_ ,
    \new_[21966]_ , \new_[21967]_ , \new_[21971]_ , \new_[21972]_ ,
    \new_[21975]_ , \new_[21978]_ , \new_[21979]_ , \new_[21980]_ ,
    \new_[21984]_ , \new_[21985]_ , \new_[21988]_ , \new_[21991]_ ,
    \new_[21992]_ , \new_[21993]_ , \new_[21997]_ , \new_[21998]_ ,
    \new_[22001]_ , \new_[22004]_ , \new_[22005]_ , \new_[22006]_ ,
    \new_[22010]_ , \new_[22011]_ , \new_[22014]_ , \new_[22017]_ ,
    \new_[22018]_ , \new_[22019]_ , \new_[22023]_ , \new_[22024]_ ,
    \new_[22027]_ , \new_[22030]_ , \new_[22031]_ , \new_[22032]_ ,
    \new_[22036]_ , \new_[22037]_ , \new_[22040]_ , \new_[22043]_ ,
    \new_[22044]_ , \new_[22045]_ , \new_[22049]_ , \new_[22050]_ ,
    \new_[22053]_ , \new_[22056]_ , \new_[22057]_ , \new_[22058]_ ,
    \new_[22062]_ , \new_[22063]_ , \new_[22066]_ , \new_[22069]_ ,
    \new_[22070]_ , \new_[22071]_ , \new_[22075]_ , \new_[22076]_ ,
    \new_[22079]_ , \new_[22082]_ , \new_[22083]_ , \new_[22084]_ ,
    \new_[22088]_ , \new_[22089]_ , \new_[22092]_ , \new_[22095]_ ,
    \new_[22096]_ , \new_[22097]_ , \new_[22101]_ , \new_[22102]_ ,
    \new_[22105]_ , \new_[22108]_ , \new_[22109]_ , \new_[22110]_ ,
    \new_[22114]_ , \new_[22115]_ , \new_[22118]_ , \new_[22121]_ ,
    \new_[22122]_ , \new_[22123]_ , \new_[22127]_ , \new_[22128]_ ,
    \new_[22131]_ , \new_[22134]_ , \new_[22135]_ , \new_[22136]_ ,
    \new_[22140]_ , \new_[22141]_ , \new_[22144]_ , \new_[22147]_ ,
    \new_[22148]_ , \new_[22149]_ , \new_[22153]_ , \new_[22154]_ ,
    \new_[22157]_ , \new_[22160]_ , \new_[22161]_ , \new_[22162]_ ,
    \new_[22166]_ , \new_[22167]_ , \new_[22170]_ , \new_[22173]_ ,
    \new_[22174]_ , \new_[22175]_ , \new_[22179]_ , \new_[22180]_ ,
    \new_[22183]_ , \new_[22186]_ , \new_[22187]_ , \new_[22188]_ ,
    \new_[22192]_ , \new_[22193]_ , \new_[22196]_ , \new_[22199]_ ,
    \new_[22200]_ , \new_[22201]_ , \new_[22205]_ , \new_[22206]_ ,
    \new_[22209]_ , \new_[22212]_ , \new_[22213]_ , \new_[22214]_ ,
    \new_[22218]_ , \new_[22219]_ , \new_[22222]_ , \new_[22225]_ ,
    \new_[22226]_ , \new_[22227]_ , \new_[22231]_ , \new_[22232]_ ,
    \new_[22235]_ , \new_[22238]_ , \new_[22239]_ , \new_[22240]_ ,
    \new_[22244]_ , \new_[22245]_ , \new_[22248]_ , \new_[22251]_ ,
    \new_[22252]_ , \new_[22253]_ , \new_[22257]_ , \new_[22258]_ ,
    \new_[22261]_ , \new_[22264]_ , \new_[22265]_ , \new_[22266]_ ,
    \new_[22270]_ , \new_[22271]_ , \new_[22274]_ , \new_[22277]_ ,
    \new_[22278]_ , \new_[22279]_ , \new_[22283]_ , \new_[22284]_ ,
    \new_[22287]_ , \new_[22290]_ , \new_[22291]_ , \new_[22292]_ ,
    \new_[22296]_ , \new_[22297]_ , \new_[22300]_ , \new_[22303]_ ,
    \new_[22304]_ , \new_[22305]_ , \new_[22309]_ , \new_[22310]_ ,
    \new_[22313]_ , \new_[22316]_ , \new_[22317]_ , \new_[22318]_ ,
    \new_[22322]_ , \new_[22323]_ , \new_[22326]_ , \new_[22329]_ ,
    \new_[22330]_ , \new_[22331]_ , \new_[22335]_ , \new_[22336]_ ,
    \new_[22339]_ , \new_[22342]_ , \new_[22343]_ , \new_[22344]_ ,
    \new_[22348]_ , \new_[22349]_ , \new_[22352]_ , \new_[22355]_ ,
    \new_[22356]_ , \new_[22357]_ , \new_[22361]_ , \new_[22362]_ ,
    \new_[22365]_ , \new_[22368]_ , \new_[22369]_ , \new_[22370]_ ,
    \new_[22374]_ , \new_[22375]_ , \new_[22378]_ , \new_[22381]_ ,
    \new_[22382]_ , \new_[22383]_ , \new_[22387]_ , \new_[22388]_ ,
    \new_[22391]_ , \new_[22394]_ , \new_[22395]_ , \new_[22396]_ ,
    \new_[22400]_ , \new_[22401]_ , \new_[22404]_ , \new_[22407]_ ,
    \new_[22408]_ , \new_[22409]_ , \new_[22413]_ , \new_[22414]_ ,
    \new_[22417]_ , \new_[22420]_ , \new_[22421]_ , \new_[22422]_ ,
    \new_[22426]_ , \new_[22427]_ , \new_[22430]_ , \new_[22433]_ ,
    \new_[22434]_ , \new_[22435]_ , \new_[22439]_ , \new_[22440]_ ,
    \new_[22443]_ , \new_[22446]_ , \new_[22447]_ , \new_[22448]_ ,
    \new_[22452]_ , \new_[22453]_ , \new_[22456]_ , \new_[22459]_ ,
    \new_[22460]_ , \new_[22461]_ , \new_[22465]_ , \new_[22466]_ ,
    \new_[22469]_ , \new_[22472]_ , \new_[22473]_ , \new_[22474]_ ,
    \new_[22478]_ , \new_[22479]_ , \new_[22482]_ , \new_[22485]_ ,
    \new_[22486]_ , \new_[22487]_ , \new_[22491]_ , \new_[22492]_ ,
    \new_[22495]_ , \new_[22498]_ , \new_[22499]_ , \new_[22500]_ ,
    \new_[22504]_ , \new_[22505]_ , \new_[22508]_ , \new_[22511]_ ,
    \new_[22512]_ , \new_[22513]_ , \new_[22517]_ , \new_[22518]_ ,
    \new_[22521]_ , \new_[22524]_ , \new_[22525]_ , \new_[22526]_ ,
    \new_[22530]_ , \new_[22531]_ , \new_[22534]_ , \new_[22537]_ ,
    \new_[22538]_ , \new_[22539]_ , \new_[22543]_ , \new_[22544]_ ,
    \new_[22547]_ , \new_[22550]_ , \new_[22551]_ , \new_[22552]_ ,
    \new_[22556]_ , \new_[22557]_ , \new_[22560]_ , \new_[22563]_ ,
    \new_[22564]_ , \new_[22565]_ , \new_[22569]_ , \new_[22570]_ ,
    \new_[22573]_ , \new_[22576]_ , \new_[22577]_ , \new_[22578]_ ,
    \new_[22582]_ , \new_[22583]_ , \new_[22586]_ , \new_[22589]_ ,
    \new_[22590]_ , \new_[22591]_ , \new_[22595]_ , \new_[22596]_ ,
    \new_[22599]_ , \new_[22602]_ , \new_[22603]_ , \new_[22604]_ ,
    \new_[22608]_ , \new_[22609]_ , \new_[22612]_ , \new_[22615]_ ,
    \new_[22616]_ , \new_[22617]_ , \new_[22621]_ , \new_[22622]_ ,
    \new_[22625]_ , \new_[22628]_ , \new_[22629]_ , \new_[22630]_ ,
    \new_[22634]_ , \new_[22635]_ , \new_[22638]_ , \new_[22641]_ ,
    \new_[22642]_ , \new_[22643]_ , \new_[22647]_ , \new_[22648]_ ,
    \new_[22651]_ , \new_[22654]_ , \new_[22655]_ , \new_[22656]_ ,
    \new_[22660]_ , \new_[22661]_ , \new_[22664]_ , \new_[22667]_ ,
    \new_[22668]_ , \new_[22669]_ , \new_[22673]_ , \new_[22674]_ ,
    \new_[22677]_ , \new_[22680]_ , \new_[22681]_ , \new_[22682]_ ,
    \new_[22686]_ , \new_[22687]_ , \new_[22690]_ , \new_[22693]_ ,
    \new_[22694]_ , \new_[22695]_ , \new_[22699]_ , \new_[22700]_ ,
    \new_[22703]_ , \new_[22706]_ , \new_[22707]_ , \new_[22708]_ ,
    \new_[22712]_ , \new_[22713]_ , \new_[22716]_ , \new_[22719]_ ,
    \new_[22720]_ , \new_[22721]_ , \new_[22725]_ , \new_[22726]_ ,
    \new_[22729]_ , \new_[22732]_ , \new_[22733]_ , \new_[22734]_ ,
    \new_[22738]_ , \new_[22739]_ , \new_[22742]_ , \new_[22745]_ ,
    \new_[22746]_ , \new_[22747]_ , \new_[22751]_ , \new_[22752]_ ,
    \new_[22755]_ , \new_[22758]_ , \new_[22759]_ , \new_[22760]_ ,
    \new_[22764]_ , \new_[22765]_ , \new_[22768]_ , \new_[22771]_ ,
    \new_[22772]_ , \new_[22773]_ , \new_[22777]_ , \new_[22778]_ ,
    \new_[22781]_ , \new_[22784]_ , \new_[22785]_ , \new_[22786]_ ,
    \new_[22790]_ , \new_[22791]_ , \new_[22794]_ , \new_[22797]_ ,
    \new_[22798]_ , \new_[22799]_ , \new_[22803]_ , \new_[22804]_ ,
    \new_[22807]_ , \new_[22810]_ , \new_[22811]_ , \new_[22812]_ ,
    \new_[22816]_ , \new_[22817]_ , \new_[22820]_ , \new_[22823]_ ,
    \new_[22824]_ , \new_[22825]_ , \new_[22829]_ , \new_[22830]_ ,
    \new_[22833]_ , \new_[22836]_ , \new_[22837]_ , \new_[22838]_ ,
    \new_[22842]_ , \new_[22843]_ , \new_[22846]_ , \new_[22849]_ ,
    \new_[22850]_ , \new_[22851]_ , \new_[22855]_ , \new_[22856]_ ,
    \new_[22859]_ , \new_[22862]_ , \new_[22863]_ , \new_[22864]_ ,
    \new_[22868]_ , \new_[22869]_ , \new_[22872]_ , \new_[22875]_ ,
    \new_[22876]_ , \new_[22877]_ , \new_[22881]_ , \new_[22882]_ ,
    \new_[22885]_ , \new_[22888]_ , \new_[22889]_ , \new_[22890]_ ,
    \new_[22894]_ , \new_[22895]_ , \new_[22898]_ , \new_[22901]_ ,
    \new_[22902]_ , \new_[22903]_ , \new_[22907]_ , \new_[22908]_ ,
    \new_[22911]_ , \new_[22914]_ , \new_[22915]_ , \new_[22916]_ ,
    \new_[22920]_ , \new_[22921]_ , \new_[22924]_ , \new_[22927]_ ,
    \new_[22928]_ , \new_[22929]_ , \new_[22933]_ , \new_[22934]_ ,
    \new_[22937]_ , \new_[22940]_ , \new_[22941]_ , \new_[22942]_ ,
    \new_[22946]_ , \new_[22947]_ , \new_[22950]_ , \new_[22953]_ ,
    \new_[22954]_ , \new_[22955]_ , \new_[22959]_ , \new_[22960]_ ,
    \new_[22963]_ , \new_[22966]_ , \new_[22967]_ , \new_[22968]_ ,
    \new_[22972]_ , \new_[22973]_ , \new_[22976]_ , \new_[22979]_ ,
    \new_[22980]_ , \new_[22981]_ , \new_[22985]_ , \new_[22986]_ ,
    \new_[22989]_ , \new_[22992]_ , \new_[22993]_ , \new_[22994]_ ,
    \new_[22998]_ , \new_[22999]_ , \new_[23002]_ , \new_[23005]_ ,
    \new_[23006]_ , \new_[23007]_ , \new_[23011]_ , \new_[23012]_ ,
    \new_[23015]_ , \new_[23018]_ , \new_[23019]_ , \new_[23020]_ ,
    \new_[23024]_ , \new_[23025]_ , \new_[23028]_ , \new_[23031]_ ,
    \new_[23032]_ , \new_[23033]_ , \new_[23037]_ , \new_[23038]_ ,
    \new_[23041]_ , \new_[23044]_ , \new_[23045]_ , \new_[23046]_ ,
    \new_[23050]_ , \new_[23051]_ , \new_[23054]_ , \new_[23057]_ ,
    \new_[23058]_ , \new_[23059]_ , \new_[23063]_ , \new_[23064]_ ,
    \new_[23067]_ , \new_[23070]_ , \new_[23071]_ , \new_[23072]_ ,
    \new_[23076]_ , \new_[23077]_ , \new_[23080]_ , \new_[23083]_ ,
    \new_[23084]_ , \new_[23085]_ , \new_[23089]_ , \new_[23090]_ ,
    \new_[23093]_ , \new_[23096]_ , \new_[23097]_ , \new_[23098]_ ,
    \new_[23102]_ , \new_[23103]_ , \new_[23106]_ , \new_[23109]_ ,
    \new_[23110]_ , \new_[23111]_ , \new_[23115]_ , \new_[23116]_ ,
    \new_[23119]_ , \new_[23122]_ , \new_[23123]_ , \new_[23124]_ ,
    \new_[23128]_ , \new_[23129]_ , \new_[23132]_ , \new_[23135]_ ,
    \new_[23136]_ , \new_[23137]_ , \new_[23141]_ , \new_[23142]_ ,
    \new_[23145]_ , \new_[23148]_ , \new_[23149]_ , \new_[23150]_ ,
    \new_[23154]_ , \new_[23155]_ , \new_[23158]_ , \new_[23161]_ ,
    \new_[23162]_ , \new_[23163]_ , \new_[23167]_ , \new_[23168]_ ,
    \new_[23171]_ , \new_[23174]_ , \new_[23175]_ , \new_[23176]_ ,
    \new_[23180]_ , \new_[23181]_ , \new_[23184]_ , \new_[23187]_ ,
    \new_[23188]_ , \new_[23189]_ , \new_[23193]_ , \new_[23194]_ ,
    \new_[23197]_ , \new_[23200]_ , \new_[23201]_ , \new_[23202]_ ,
    \new_[23206]_ , \new_[23207]_ , \new_[23210]_ , \new_[23213]_ ,
    \new_[23214]_ , \new_[23215]_ , \new_[23219]_ , \new_[23220]_ ,
    \new_[23223]_ , \new_[23226]_ , \new_[23227]_ , \new_[23228]_ ,
    \new_[23232]_ , \new_[23233]_ , \new_[23236]_ , \new_[23239]_ ,
    \new_[23240]_ , \new_[23241]_ , \new_[23245]_ , \new_[23246]_ ,
    \new_[23249]_ , \new_[23252]_ , \new_[23253]_ , \new_[23254]_ ,
    \new_[23258]_ , \new_[23259]_ , \new_[23262]_ , \new_[23265]_ ,
    \new_[23266]_ , \new_[23267]_ , \new_[23271]_ , \new_[23272]_ ,
    \new_[23275]_ , \new_[23278]_ , \new_[23279]_ , \new_[23280]_ ,
    \new_[23284]_ , \new_[23285]_ , \new_[23288]_ , \new_[23291]_ ,
    \new_[23292]_ , \new_[23293]_ , \new_[23297]_ , \new_[23298]_ ,
    \new_[23301]_ , \new_[23304]_ , \new_[23305]_ , \new_[23306]_ ,
    \new_[23310]_ , \new_[23311]_ , \new_[23314]_ , \new_[23317]_ ,
    \new_[23318]_ , \new_[23319]_ , \new_[23323]_ , \new_[23324]_ ,
    \new_[23327]_ , \new_[23330]_ , \new_[23331]_ , \new_[23332]_ ,
    \new_[23336]_ , \new_[23337]_ , \new_[23340]_ , \new_[23343]_ ,
    \new_[23344]_ , \new_[23345]_ , \new_[23349]_ , \new_[23350]_ ,
    \new_[23353]_ , \new_[23356]_ , \new_[23357]_ , \new_[23358]_ ,
    \new_[23362]_ , \new_[23363]_ , \new_[23366]_ , \new_[23369]_ ,
    \new_[23370]_ , \new_[23371]_ , \new_[23375]_ , \new_[23376]_ ,
    \new_[23379]_ , \new_[23382]_ , \new_[23383]_ , \new_[23384]_ ,
    \new_[23388]_ , \new_[23389]_ , \new_[23392]_ , \new_[23395]_ ,
    \new_[23396]_ , \new_[23397]_ , \new_[23401]_ , \new_[23402]_ ,
    \new_[23405]_ , \new_[23408]_ , \new_[23409]_ , \new_[23410]_ ,
    \new_[23414]_ , \new_[23415]_ , \new_[23418]_ , \new_[23421]_ ,
    \new_[23422]_ , \new_[23423]_ , \new_[23427]_ , \new_[23428]_ ,
    \new_[23431]_ , \new_[23434]_ , \new_[23435]_ , \new_[23436]_ ,
    \new_[23440]_ , \new_[23441]_ , \new_[23444]_ , \new_[23447]_ ,
    \new_[23448]_ , \new_[23449]_ , \new_[23453]_ , \new_[23454]_ ,
    \new_[23457]_ , \new_[23460]_ , \new_[23461]_ , \new_[23462]_ ,
    \new_[23466]_ , \new_[23467]_ , \new_[23470]_ , \new_[23473]_ ,
    \new_[23474]_ , \new_[23475]_ , \new_[23479]_ , \new_[23480]_ ,
    \new_[23483]_ , \new_[23486]_ , \new_[23487]_ , \new_[23488]_ ,
    \new_[23492]_ , \new_[23493]_ , \new_[23496]_ , \new_[23499]_ ,
    \new_[23500]_ , \new_[23501]_ , \new_[23505]_ , \new_[23506]_ ,
    \new_[23509]_ , \new_[23512]_ , \new_[23513]_ , \new_[23514]_ ,
    \new_[23518]_ , \new_[23519]_ , \new_[23522]_ , \new_[23525]_ ,
    \new_[23526]_ , \new_[23527]_ , \new_[23531]_ , \new_[23532]_ ,
    \new_[23535]_ , \new_[23538]_ , \new_[23539]_ , \new_[23540]_ ,
    \new_[23544]_ , \new_[23545]_ , \new_[23548]_ , \new_[23551]_ ,
    \new_[23552]_ , \new_[23553]_ , \new_[23557]_ , \new_[23558]_ ,
    \new_[23561]_ , \new_[23564]_ , \new_[23565]_ , \new_[23566]_ ,
    \new_[23570]_ , \new_[23571]_ , \new_[23574]_ , \new_[23577]_ ,
    \new_[23578]_ , \new_[23579]_ , \new_[23583]_ , \new_[23584]_ ,
    \new_[23587]_ , \new_[23590]_ , \new_[23591]_ , \new_[23592]_ ,
    \new_[23596]_ , \new_[23597]_ , \new_[23600]_ , \new_[23603]_ ,
    \new_[23604]_ , \new_[23605]_ , \new_[23609]_ , \new_[23610]_ ,
    \new_[23613]_ , \new_[23616]_ , \new_[23617]_ , \new_[23618]_ ,
    \new_[23622]_ , \new_[23623]_ , \new_[23626]_ , \new_[23629]_ ,
    \new_[23630]_ , \new_[23631]_ , \new_[23635]_ , \new_[23636]_ ,
    \new_[23639]_ , \new_[23642]_ , \new_[23643]_ , \new_[23644]_ ,
    \new_[23648]_ , \new_[23649]_ , \new_[23652]_ , \new_[23655]_ ,
    \new_[23656]_ , \new_[23657]_ , \new_[23661]_ , \new_[23662]_ ,
    \new_[23665]_ , \new_[23668]_ , \new_[23669]_ , \new_[23670]_ ,
    \new_[23674]_ , \new_[23675]_ , \new_[23678]_ , \new_[23681]_ ,
    \new_[23682]_ , \new_[23683]_ , \new_[23687]_ , \new_[23688]_ ,
    \new_[23691]_ , \new_[23694]_ , \new_[23695]_ , \new_[23696]_ ,
    \new_[23700]_ , \new_[23701]_ , \new_[23704]_ , \new_[23707]_ ,
    \new_[23708]_ , \new_[23709]_ , \new_[23713]_ , \new_[23714]_ ,
    \new_[23717]_ , \new_[23720]_ , \new_[23721]_ , \new_[23722]_ ,
    \new_[23726]_ , \new_[23727]_ , \new_[23730]_ , \new_[23733]_ ,
    \new_[23734]_ , \new_[23735]_ , \new_[23739]_ , \new_[23740]_ ,
    \new_[23743]_ , \new_[23746]_ , \new_[23747]_ , \new_[23748]_ ,
    \new_[23752]_ , \new_[23753]_ , \new_[23756]_ , \new_[23759]_ ,
    \new_[23760]_ , \new_[23761]_ , \new_[23765]_ , \new_[23766]_ ,
    \new_[23769]_ , \new_[23772]_ , \new_[23773]_ , \new_[23774]_ ,
    \new_[23778]_ , \new_[23779]_ , \new_[23782]_ , \new_[23785]_ ,
    \new_[23786]_ , \new_[23787]_ , \new_[23791]_ , \new_[23792]_ ,
    \new_[23795]_ , \new_[23798]_ , \new_[23799]_ , \new_[23800]_ ,
    \new_[23804]_ , \new_[23805]_ , \new_[23808]_ , \new_[23811]_ ,
    \new_[23812]_ , \new_[23813]_ , \new_[23817]_ , \new_[23818]_ ,
    \new_[23821]_ , \new_[23824]_ , \new_[23825]_ , \new_[23826]_ ,
    \new_[23830]_ , \new_[23831]_ , \new_[23834]_ , \new_[23837]_ ,
    \new_[23838]_ , \new_[23839]_ , \new_[23843]_ , \new_[23844]_ ,
    \new_[23847]_ , \new_[23850]_ , \new_[23851]_ , \new_[23852]_ ,
    \new_[23856]_ , \new_[23857]_ , \new_[23860]_ , \new_[23863]_ ,
    \new_[23864]_ , \new_[23865]_ , \new_[23869]_ , \new_[23870]_ ,
    \new_[23873]_ , \new_[23876]_ , \new_[23877]_ , \new_[23878]_ ,
    \new_[23882]_ , \new_[23883]_ , \new_[23886]_ , \new_[23889]_ ,
    \new_[23890]_ , \new_[23891]_ , \new_[23895]_ , \new_[23896]_ ,
    \new_[23899]_ , \new_[23902]_ , \new_[23903]_ , \new_[23904]_ ,
    \new_[23908]_ , \new_[23909]_ , \new_[23912]_ , \new_[23915]_ ,
    \new_[23916]_ , \new_[23917]_ , \new_[23921]_ , \new_[23922]_ ,
    \new_[23925]_ , \new_[23928]_ , \new_[23929]_ , \new_[23930]_ ,
    \new_[23934]_ , \new_[23935]_ , \new_[23938]_ , \new_[23941]_ ,
    \new_[23942]_ , \new_[23943]_ , \new_[23947]_ , \new_[23948]_ ,
    \new_[23951]_ , \new_[23954]_ , \new_[23955]_ , \new_[23956]_ ,
    \new_[23960]_ , \new_[23961]_ , \new_[23964]_ , \new_[23967]_ ,
    \new_[23968]_ , \new_[23969]_ , \new_[23973]_ , \new_[23974]_ ,
    \new_[23977]_ , \new_[23980]_ , \new_[23981]_ , \new_[23982]_ ,
    \new_[23986]_ , \new_[23987]_ , \new_[23990]_ , \new_[23993]_ ,
    \new_[23994]_ , \new_[23995]_ , \new_[23999]_ , \new_[24000]_ ,
    \new_[24003]_ , \new_[24006]_ , \new_[24007]_ , \new_[24008]_ ,
    \new_[24012]_ , \new_[24013]_ , \new_[24016]_ , \new_[24019]_ ,
    \new_[24020]_ , \new_[24021]_ , \new_[24025]_ , \new_[24026]_ ,
    \new_[24029]_ , \new_[24032]_ , \new_[24033]_ , \new_[24034]_ ,
    \new_[24038]_ , \new_[24039]_ , \new_[24042]_ , \new_[24045]_ ,
    \new_[24046]_ , \new_[24047]_ , \new_[24051]_ , \new_[24052]_ ,
    \new_[24055]_ , \new_[24058]_ , \new_[24059]_ , \new_[24060]_ ,
    \new_[24064]_ , \new_[24065]_ , \new_[24068]_ , \new_[24071]_ ,
    \new_[24072]_ , \new_[24073]_ , \new_[24077]_ , \new_[24078]_ ,
    \new_[24081]_ , \new_[24084]_ , \new_[24085]_ , \new_[24086]_ ,
    \new_[24090]_ , \new_[24091]_ , \new_[24094]_ , \new_[24097]_ ,
    \new_[24098]_ , \new_[24099]_ , \new_[24103]_ , \new_[24104]_ ,
    \new_[24107]_ , \new_[24110]_ , \new_[24111]_ , \new_[24112]_ ,
    \new_[24116]_ , \new_[24117]_ , \new_[24120]_ , \new_[24123]_ ,
    \new_[24124]_ , \new_[24125]_ , \new_[24129]_ , \new_[24130]_ ,
    \new_[24133]_ , \new_[24136]_ , \new_[24137]_ , \new_[24138]_ ,
    \new_[24142]_ , \new_[24143]_ , \new_[24146]_ , \new_[24149]_ ,
    \new_[24150]_ , \new_[24151]_ , \new_[24155]_ , \new_[24156]_ ,
    \new_[24159]_ , \new_[24162]_ , \new_[24163]_ , \new_[24164]_ ,
    \new_[24168]_ , \new_[24169]_ , \new_[24172]_ , \new_[24175]_ ,
    \new_[24176]_ , \new_[24177]_ , \new_[24181]_ , \new_[24182]_ ,
    \new_[24185]_ , \new_[24188]_ , \new_[24189]_ , \new_[24190]_ ,
    \new_[24194]_ , \new_[24195]_ , \new_[24198]_ , \new_[24201]_ ,
    \new_[24202]_ , \new_[24203]_ , \new_[24207]_ , \new_[24208]_ ,
    \new_[24211]_ , \new_[24214]_ , \new_[24215]_ , \new_[24216]_ ,
    \new_[24220]_ , \new_[24221]_ , \new_[24224]_ , \new_[24227]_ ,
    \new_[24228]_ , \new_[24229]_ , \new_[24233]_ , \new_[24234]_ ,
    \new_[24237]_ , \new_[24240]_ , \new_[24241]_ , \new_[24242]_ ,
    \new_[24246]_ , \new_[24247]_ , \new_[24250]_ , \new_[24253]_ ,
    \new_[24254]_ , \new_[24255]_ , \new_[24259]_ , \new_[24260]_ ,
    \new_[24263]_ , \new_[24266]_ , \new_[24267]_ , \new_[24268]_ ,
    \new_[24272]_ , \new_[24273]_ , \new_[24276]_ , \new_[24279]_ ,
    \new_[24280]_ , \new_[24281]_ , \new_[24285]_ , \new_[24286]_ ,
    \new_[24289]_ , \new_[24292]_ , \new_[24293]_ , \new_[24294]_ ,
    \new_[24298]_ , \new_[24299]_ , \new_[24302]_ , \new_[24305]_ ,
    \new_[24306]_ , \new_[24307]_ , \new_[24311]_ , \new_[24312]_ ,
    \new_[24315]_ , \new_[24318]_ , \new_[24319]_ , \new_[24320]_ ,
    \new_[24324]_ , \new_[24325]_ , \new_[24328]_ , \new_[24331]_ ,
    \new_[24332]_ , \new_[24333]_ , \new_[24337]_ , \new_[24338]_ ,
    \new_[24341]_ , \new_[24344]_ , \new_[24345]_ , \new_[24346]_ ,
    \new_[24350]_ , \new_[24351]_ , \new_[24354]_ , \new_[24357]_ ,
    \new_[24358]_ , \new_[24359]_ , \new_[24363]_ , \new_[24364]_ ,
    \new_[24367]_ , \new_[24370]_ , \new_[24371]_ , \new_[24372]_ ,
    \new_[24376]_ , \new_[24377]_ , \new_[24380]_ , \new_[24383]_ ,
    \new_[24384]_ , \new_[24385]_ , \new_[24389]_ , \new_[24390]_ ,
    \new_[24393]_ , \new_[24396]_ , \new_[24397]_ , \new_[24398]_ ,
    \new_[24402]_ , \new_[24403]_ , \new_[24406]_ , \new_[24409]_ ,
    \new_[24410]_ , \new_[24411]_ , \new_[24415]_ , \new_[24416]_ ,
    \new_[24419]_ , \new_[24422]_ , \new_[24423]_ , \new_[24424]_ ,
    \new_[24428]_ , \new_[24429]_ , \new_[24432]_ , \new_[24435]_ ,
    \new_[24436]_ , \new_[24437]_ , \new_[24441]_ , \new_[24442]_ ,
    \new_[24445]_ , \new_[24448]_ , \new_[24449]_ , \new_[24450]_ ,
    \new_[24454]_ , \new_[24455]_ , \new_[24458]_ , \new_[24461]_ ,
    \new_[24462]_ , \new_[24463]_ , \new_[24467]_ , \new_[24468]_ ,
    \new_[24471]_ , \new_[24474]_ , \new_[24475]_ , \new_[24476]_ ,
    \new_[24480]_ , \new_[24481]_ , \new_[24484]_ , \new_[24487]_ ,
    \new_[24488]_ , \new_[24489]_ , \new_[24493]_ , \new_[24494]_ ,
    \new_[24497]_ , \new_[24500]_ , \new_[24501]_ , \new_[24502]_ ,
    \new_[24506]_ , \new_[24507]_ , \new_[24510]_ , \new_[24513]_ ,
    \new_[24514]_ , \new_[24515]_ , \new_[24519]_ , \new_[24520]_ ,
    \new_[24523]_ , \new_[24526]_ , \new_[24527]_ , \new_[24528]_ ,
    \new_[24532]_ , \new_[24533]_ , \new_[24536]_ , \new_[24539]_ ,
    \new_[24540]_ , \new_[24541]_ , \new_[24545]_ , \new_[24546]_ ,
    \new_[24549]_ , \new_[24552]_ , \new_[24553]_ , \new_[24554]_ ,
    \new_[24558]_ , \new_[24559]_ , \new_[24562]_ , \new_[24565]_ ,
    \new_[24566]_ , \new_[24567]_ , \new_[24571]_ , \new_[24572]_ ,
    \new_[24575]_ , \new_[24578]_ , \new_[24579]_ , \new_[24580]_ ,
    \new_[24584]_ , \new_[24585]_ , \new_[24588]_ , \new_[24591]_ ,
    \new_[24592]_ , \new_[24593]_ , \new_[24597]_ , \new_[24598]_ ,
    \new_[24601]_ , \new_[24604]_ , \new_[24605]_ , \new_[24606]_ ,
    \new_[24610]_ , \new_[24611]_ , \new_[24614]_ , \new_[24617]_ ,
    \new_[24618]_ , \new_[24619]_ , \new_[24623]_ , \new_[24624]_ ,
    \new_[24627]_ , \new_[24630]_ , \new_[24631]_ , \new_[24632]_ ,
    \new_[24636]_ , \new_[24637]_ , \new_[24640]_ , \new_[24643]_ ,
    \new_[24644]_ , \new_[24645]_ , \new_[24649]_ , \new_[24650]_ ,
    \new_[24653]_ , \new_[24656]_ , \new_[24657]_ , \new_[24658]_ ,
    \new_[24662]_ , \new_[24663]_ , \new_[24666]_ , \new_[24669]_ ,
    \new_[24670]_ , \new_[24671]_ , \new_[24675]_ , \new_[24676]_ ,
    \new_[24679]_ , \new_[24682]_ , \new_[24683]_ , \new_[24684]_ ,
    \new_[24688]_ , \new_[24689]_ , \new_[24692]_ , \new_[24695]_ ,
    \new_[24696]_ , \new_[24697]_ , \new_[24701]_ , \new_[24702]_ ,
    \new_[24705]_ , \new_[24708]_ , \new_[24709]_ , \new_[24710]_ ,
    \new_[24714]_ , \new_[24715]_ , \new_[24718]_ , \new_[24721]_ ,
    \new_[24722]_ , \new_[24723]_ , \new_[24727]_ , \new_[24728]_ ,
    \new_[24731]_ , \new_[24734]_ , \new_[24735]_ , \new_[24736]_ ,
    \new_[24740]_ , \new_[24741]_ , \new_[24744]_ , \new_[24747]_ ,
    \new_[24748]_ , \new_[24749]_ , \new_[24753]_ , \new_[24754]_ ,
    \new_[24757]_ , \new_[24760]_ , \new_[24761]_ , \new_[24762]_ ,
    \new_[24766]_ , \new_[24767]_ , \new_[24770]_ , \new_[24773]_ ,
    \new_[24774]_ , \new_[24775]_ , \new_[24779]_ , \new_[24780]_ ,
    \new_[24783]_ , \new_[24786]_ , \new_[24787]_ , \new_[24788]_ ,
    \new_[24792]_ , \new_[24793]_ , \new_[24796]_ , \new_[24799]_ ,
    \new_[24800]_ , \new_[24801]_ , \new_[24805]_ , \new_[24806]_ ,
    \new_[24809]_ , \new_[24812]_ , \new_[24813]_ , \new_[24814]_ ,
    \new_[24818]_ , \new_[24819]_ , \new_[24822]_ , \new_[24825]_ ,
    \new_[24826]_ , \new_[24827]_ , \new_[24831]_ , \new_[24832]_ ,
    \new_[24835]_ , \new_[24838]_ , \new_[24839]_ , \new_[24840]_ ,
    \new_[24844]_ , \new_[24845]_ , \new_[24848]_ , \new_[24851]_ ,
    \new_[24852]_ , \new_[24853]_ , \new_[24857]_ , \new_[24858]_ ,
    \new_[24861]_ , \new_[24864]_ , \new_[24865]_ , \new_[24866]_ ,
    \new_[24870]_ , \new_[24871]_ , \new_[24874]_ , \new_[24877]_ ,
    \new_[24878]_ , \new_[24879]_ , \new_[24883]_ , \new_[24884]_ ,
    \new_[24887]_ , \new_[24890]_ , \new_[24891]_ , \new_[24892]_ ,
    \new_[24896]_ , \new_[24897]_ , \new_[24900]_ , \new_[24903]_ ,
    \new_[24904]_ , \new_[24905]_ , \new_[24909]_ , \new_[24910]_ ,
    \new_[24913]_ , \new_[24916]_ , \new_[24917]_ , \new_[24918]_ ,
    \new_[24922]_ , \new_[24923]_ , \new_[24926]_ , \new_[24929]_ ,
    \new_[24930]_ , \new_[24931]_ , \new_[24935]_ , \new_[24936]_ ,
    \new_[24939]_ , \new_[24942]_ , \new_[24943]_ , \new_[24944]_ ,
    \new_[24948]_ , \new_[24949]_ , \new_[24952]_ , \new_[24955]_ ,
    \new_[24956]_ , \new_[24957]_ , \new_[24961]_ , \new_[24962]_ ,
    \new_[24965]_ , \new_[24968]_ , \new_[24969]_ , \new_[24970]_ ,
    \new_[24974]_ , \new_[24975]_ , \new_[24978]_ , \new_[24981]_ ,
    \new_[24982]_ , \new_[24983]_ , \new_[24987]_ , \new_[24988]_ ,
    \new_[24991]_ , \new_[24994]_ , \new_[24995]_ , \new_[24996]_ ,
    \new_[25000]_ , \new_[25001]_ , \new_[25004]_ , \new_[25007]_ ,
    \new_[25008]_ , \new_[25009]_ , \new_[25013]_ , \new_[25014]_ ,
    \new_[25017]_ , \new_[25020]_ , \new_[25021]_ , \new_[25022]_ ,
    \new_[25026]_ , \new_[25027]_ , \new_[25030]_ , \new_[25033]_ ,
    \new_[25034]_ , \new_[25035]_ , \new_[25039]_ , \new_[25040]_ ,
    \new_[25043]_ , \new_[25046]_ , \new_[25047]_ , \new_[25048]_ ,
    \new_[25052]_ , \new_[25053]_ , \new_[25056]_ , \new_[25059]_ ,
    \new_[25060]_ , \new_[25061]_ , \new_[25065]_ , \new_[25066]_ ,
    \new_[25069]_ , \new_[25072]_ , \new_[25073]_ , \new_[25074]_ ,
    \new_[25078]_ , \new_[25079]_ , \new_[25082]_ , \new_[25085]_ ,
    \new_[25086]_ , \new_[25087]_ , \new_[25091]_ , \new_[25092]_ ,
    \new_[25095]_ , \new_[25098]_ , \new_[25099]_ , \new_[25100]_ ,
    \new_[25104]_ , \new_[25105]_ , \new_[25108]_ , \new_[25111]_ ,
    \new_[25112]_ , \new_[25113]_ , \new_[25117]_ , \new_[25118]_ ,
    \new_[25121]_ , \new_[25124]_ , \new_[25125]_ , \new_[25126]_ ,
    \new_[25130]_ , \new_[25131]_ , \new_[25134]_ , \new_[25137]_ ,
    \new_[25138]_ , \new_[25139]_ , \new_[25143]_ , \new_[25144]_ ,
    \new_[25147]_ , \new_[25150]_ , \new_[25151]_ , \new_[25152]_ ,
    \new_[25156]_ , \new_[25157]_ , \new_[25160]_ , \new_[25163]_ ,
    \new_[25164]_ , \new_[25165]_ , \new_[25169]_ , \new_[25170]_ ,
    \new_[25173]_ , \new_[25176]_ , \new_[25177]_ , \new_[25178]_ ,
    \new_[25182]_ , \new_[25183]_ , \new_[25186]_ , \new_[25189]_ ,
    \new_[25190]_ , \new_[25191]_ , \new_[25195]_ , \new_[25196]_ ,
    \new_[25199]_ , \new_[25202]_ , \new_[25203]_ , \new_[25204]_ ,
    \new_[25208]_ , \new_[25209]_ , \new_[25212]_ , \new_[25215]_ ,
    \new_[25216]_ , \new_[25217]_ , \new_[25221]_ , \new_[25222]_ ,
    \new_[25225]_ , \new_[25228]_ , \new_[25229]_ , \new_[25230]_ ,
    \new_[25234]_ , \new_[25235]_ , \new_[25238]_ , \new_[25241]_ ,
    \new_[25242]_ , \new_[25243]_ , \new_[25247]_ , \new_[25248]_ ,
    \new_[25251]_ , \new_[25254]_ , \new_[25255]_ , \new_[25256]_ ,
    \new_[25260]_ , \new_[25261]_ , \new_[25264]_ , \new_[25267]_ ,
    \new_[25268]_ , \new_[25269]_ , \new_[25273]_ , \new_[25274]_ ,
    \new_[25277]_ , \new_[25280]_ , \new_[25281]_ , \new_[25282]_ ,
    \new_[25286]_ , \new_[25287]_ , \new_[25290]_ , \new_[25293]_ ,
    \new_[25294]_ , \new_[25295]_ , \new_[25299]_ , \new_[25300]_ ,
    \new_[25303]_ , \new_[25306]_ , \new_[25307]_ , \new_[25308]_ ,
    \new_[25312]_ , \new_[25313]_ , \new_[25316]_ , \new_[25319]_ ,
    \new_[25320]_ , \new_[25321]_ , \new_[25325]_ , \new_[25326]_ ,
    \new_[25329]_ , \new_[25332]_ , \new_[25333]_ , \new_[25334]_ ,
    \new_[25338]_ , \new_[25339]_ , \new_[25342]_ , \new_[25345]_ ,
    \new_[25346]_ , \new_[25347]_ , \new_[25351]_ , \new_[25352]_ ,
    \new_[25355]_ , \new_[25358]_ , \new_[25359]_ , \new_[25360]_ ,
    \new_[25364]_ , \new_[25365]_ , \new_[25368]_ , \new_[25371]_ ,
    \new_[25372]_ , \new_[25373]_ , \new_[25377]_ , \new_[25378]_ ,
    \new_[25381]_ , \new_[25384]_ , \new_[25385]_ , \new_[25386]_ ,
    \new_[25390]_ , \new_[25391]_ , \new_[25394]_ , \new_[25397]_ ,
    \new_[25398]_ , \new_[25399]_ , \new_[25403]_ , \new_[25404]_ ,
    \new_[25407]_ , \new_[25410]_ , \new_[25411]_ , \new_[25412]_ ,
    \new_[25416]_ , \new_[25417]_ , \new_[25420]_ , \new_[25423]_ ,
    \new_[25424]_ , \new_[25425]_ , \new_[25429]_ , \new_[25430]_ ,
    \new_[25433]_ , \new_[25436]_ , \new_[25437]_ , \new_[25438]_ ,
    \new_[25442]_ , \new_[25443]_ , \new_[25446]_ , \new_[25449]_ ,
    \new_[25450]_ , \new_[25451]_ , \new_[25455]_ , \new_[25456]_ ,
    \new_[25459]_ , \new_[25462]_ , \new_[25463]_ , \new_[25464]_ ,
    \new_[25468]_ , \new_[25469]_ , \new_[25472]_ , \new_[25475]_ ,
    \new_[25476]_ , \new_[25477]_ , \new_[25481]_ , \new_[25482]_ ,
    \new_[25485]_ , \new_[25488]_ , \new_[25489]_ , \new_[25490]_ ,
    \new_[25494]_ , \new_[25495]_ , \new_[25498]_ , \new_[25501]_ ,
    \new_[25502]_ , \new_[25503]_ , \new_[25507]_ , \new_[25508]_ ,
    \new_[25511]_ , \new_[25514]_ , \new_[25515]_ , \new_[25516]_ ,
    \new_[25520]_ , \new_[25521]_ , \new_[25524]_ , \new_[25527]_ ,
    \new_[25528]_ , \new_[25529]_ , \new_[25533]_ , \new_[25534]_ ,
    \new_[25537]_ , \new_[25540]_ , \new_[25541]_ , \new_[25542]_ ,
    \new_[25546]_ , \new_[25547]_ , \new_[25550]_ , \new_[25553]_ ,
    \new_[25554]_ , \new_[25555]_ , \new_[25559]_ , \new_[25560]_ ,
    \new_[25563]_ , \new_[25566]_ , \new_[25567]_ , \new_[25568]_ ,
    \new_[25572]_ , \new_[25573]_ , \new_[25576]_ , \new_[25579]_ ,
    \new_[25580]_ , \new_[25581]_ , \new_[25585]_ , \new_[25586]_ ,
    \new_[25589]_ , \new_[25592]_ , \new_[25593]_ , \new_[25594]_ ,
    \new_[25598]_ , \new_[25599]_ , \new_[25602]_ , \new_[25605]_ ,
    \new_[25606]_ , \new_[25607]_ , \new_[25611]_ , \new_[25612]_ ,
    \new_[25615]_ , \new_[25618]_ , \new_[25619]_ , \new_[25620]_ ,
    \new_[25624]_ , \new_[25625]_ , \new_[25628]_ , \new_[25631]_ ,
    \new_[25632]_ , \new_[25633]_ , \new_[25637]_ , \new_[25638]_ ,
    \new_[25641]_ , \new_[25644]_ , \new_[25645]_ , \new_[25646]_ ,
    \new_[25650]_ , \new_[25651]_ , \new_[25654]_ , \new_[25657]_ ,
    \new_[25658]_ , \new_[25659]_ , \new_[25663]_ , \new_[25664]_ ,
    \new_[25667]_ , \new_[25670]_ , \new_[25671]_ , \new_[25672]_ ,
    \new_[25676]_ , \new_[25677]_ , \new_[25680]_ , \new_[25683]_ ,
    \new_[25684]_ , \new_[25685]_ , \new_[25689]_ , \new_[25690]_ ,
    \new_[25693]_ , \new_[25696]_ , \new_[25697]_ , \new_[25698]_ ,
    \new_[25702]_ , \new_[25703]_ , \new_[25706]_ , \new_[25709]_ ,
    \new_[25710]_ , \new_[25711]_ , \new_[25715]_ , \new_[25716]_ ,
    \new_[25719]_ , \new_[25722]_ , \new_[25723]_ , \new_[25724]_ ,
    \new_[25728]_ , \new_[25729]_ , \new_[25732]_ , \new_[25735]_ ,
    \new_[25736]_ , \new_[25737]_ , \new_[25741]_ , \new_[25742]_ ,
    \new_[25745]_ , \new_[25748]_ , \new_[25749]_ , \new_[25750]_ ,
    \new_[25754]_ , \new_[25755]_ , \new_[25758]_ , \new_[25761]_ ,
    \new_[25762]_ , \new_[25763]_ , \new_[25767]_ , \new_[25768]_ ,
    \new_[25771]_ , \new_[25774]_ , \new_[25775]_ , \new_[25776]_ ,
    \new_[25780]_ , \new_[25781]_ , \new_[25784]_ , \new_[25787]_ ,
    \new_[25788]_ , \new_[25789]_ , \new_[25793]_ , \new_[25794]_ ,
    \new_[25797]_ , \new_[25800]_ , \new_[25801]_ , \new_[25802]_ ,
    \new_[25806]_ , \new_[25807]_ , \new_[25810]_ , \new_[25813]_ ,
    \new_[25814]_ , \new_[25815]_ , \new_[25819]_ , \new_[25820]_ ,
    \new_[25823]_ , \new_[25826]_ , \new_[25827]_ , \new_[25828]_ ,
    \new_[25832]_ , \new_[25833]_ , \new_[25836]_ , \new_[25839]_ ,
    \new_[25840]_ , \new_[25841]_ , \new_[25845]_ , \new_[25846]_ ,
    \new_[25849]_ , \new_[25852]_ , \new_[25853]_ , \new_[25854]_ ,
    \new_[25858]_ , \new_[25859]_ , \new_[25862]_ , \new_[25865]_ ,
    \new_[25866]_ , \new_[25867]_ , \new_[25871]_ , \new_[25872]_ ,
    \new_[25875]_ , \new_[25878]_ , \new_[25879]_ , \new_[25880]_ ,
    \new_[25884]_ , \new_[25885]_ , \new_[25888]_ , \new_[25891]_ ,
    \new_[25892]_ , \new_[25893]_ , \new_[25897]_ , \new_[25898]_ ,
    \new_[25901]_ , \new_[25904]_ , \new_[25905]_ , \new_[25906]_ ,
    \new_[25910]_ , \new_[25911]_ , \new_[25914]_ , \new_[25917]_ ,
    \new_[25918]_ , \new_[25919]_ , \new_[25923]_ , \new_[25924]_ ,
    \new_[25927]_ , \new_[25930]_ , \new_[25931]_ , \new_[25932]_ ,
    \new_[25936]_ , \new_[25937]_ , \new_[25940]_ , \new_[25943]_ ,
    \new_[25944]_ , \new_[25945]_ , \new_[25949]_ , \new_[25950]_ ,
    \new_[25953]_ , \new_[25956]_ , \new_[25957]_ , \new_[25958]_ ,
    \new_[25962]_ , \new_[25963]_ , \new_[25966]_ , \new_[25969]_ ,
    \new_[25970]_ , \new_[25971]_ , \new_[25975]_ , \new_[25976]_ ,
    \new_[25979]_ , \new_[25982]_ , \new_[25983]_ , \new_[25984]_ ,
    \new_[25988]_ , \new_[25989]_ , \new_[25992]_ , \new_[25995]_ ,
    \new_[25996]_ , \new_[25997]_ , \new_[26001]_ , \new_[26002]_ ,
    \new_[26005]_ , \new_[26008]_ , \new_[26009]_ , \new_[26010]_ ,
    \new_[26014]_ , \new_[26015]_ , \new_[26018]_ , \new_[26021]_ ,
    \new_[26022]_ , \new_[26023]_ , \new_[26027]_ , \new_[26028]_ ,
    \new_[26031]_ , \new_[26034]_ , \new_[26035]_ , \new_[26036]_ ,
    \new_[26040]_ , \new_[26041]_ , \new_[26044]_ , \new_[26047]_ ,
    \new_[26048]_ , \new_[26049]_ , \new_[26053]_ , \new_[26054]_ ,
    \new_[26057]_ , \new_[26060]_ , \new_[26061]_ , \new_[26062]_ ,
    \new_[26066]_ , \new_[26067]_ , \new_[26070]_ , \new_[26073]_ ,
    \new_[26074]_ , \new_[26075]_ , \new_[26079]_ , \new_[26080]_ ,
    \new_[26083]_ , \new_[26086]_ , \new_[26087]_ , \new_[26088]_ ,
    \new_[26092]_ , \new_[26093]_ , \new_[26096]_ , \new_[26099]_ ,
    \new_[26100]_ , \new_[26101]_ , \new_[26105]_ , \new_[26106]_ ,
    \new_[26109]_ , \new_[26112]_ , \new_[26113]_ , \new_[26114]_ ,
    \new_[26118]_ , \new_[26119]_ , \new_[26122]_ , \new_[26125]_ ,
    \new_[26126]_ , \new_[26127]_ , \new_[26131]_ , \new_[26132]_ ,
    \new_[26135]_ , \new_[26138]_ , \new_[26139]_ , \new_[26140]_ ,
    \new_[26144]_ , \new_[26145]_ , \new_[26148]_ , \new_[26151]_ ,
    \new_[26152]_ , \new_[26153]_ , \new_[26157]_ , \new_[26158]_ ,
    \new_[26161]_ , \new_[26164]_ , \new_[26165]_ , \new_[26166]_ ,
    \new_[26170]_ , \new_[26171]_ , \new_[26174]_ , \new_[26177]_ ,
    \new_[26178]_ , \new_[26179]_ , \new_[26183]_ , \new_[26184]_ ,
    \new_[26187]_ , \new_[26190]_ , \new_[26191]_ , \new_[26192]_ ,
    \new_[26196]_ , \new_[26197]_ , \new_[26200]_ , \new_[26203]_ ,
    \new_[26204]_ , \new_[26205]_ , \new_[26209]_ , \new_[26210]_ ,
    \new_[26213]_ , \new_[26216]_ , \new_[26217]_ , \new_[26218]_ ,
    \new_[26222]_ , \new_[26223]_ , \new_[26226]_ , \new_[26229]_ ,
    \new_[26230]_ , \new_[26231]_ , \new_[26235]_ , \new_[26236]_ ,
    \new_[26239]_ , \new_[26242]_ , \new_[26243]_ , \new_[26244]_ ,
    \new_[26248]_ , \new_[26249]_ , \new_[26252]_ , \new_[26255]_ ,
    \new_[26256]_ , \new_[26257]_ , \new_[26261]_ , \new_[26262]_ ,
    \new_[26265]_ , \new_[26268]_ , \new_[26269]_ , \new_[26270]_ ,
    \new_[26274]_ , \new_[26275]_ , \new_[26278]_ , \new_[26281]_ ,
    \new_[26282]_ , \new_[26283]_ , \new_[26287]_ , \new_[26288]_ ,
    \new_[26291]_ , \new_[26294]_ , \new_[26295]_ , \new_[26296]_ ,
    \new_[26300]_ , \new_[26301]_ , \new_[26304]_ , \new_[26307]_ ,
    \new_[26308]_ , \new_[26309]_ , \new_[26313]_ , \new_[26314]_ ,
    \new_[26317]_ , \new_[26320]_ , \new_[26321]_ , \new_[26322]_ ,
    \new_[26326]_ , \new_[26327]_ , \new_[26330]_ , \new_[26333]_ ,
    \new_[26334]_ , \new_[26335]_ , \new_[26339]_ , \new_[26340]_ ,
    \new_[26343]_ , \new_[26346]_ , \new_[26347]_ , \new_[26348]_ ,
    \new_[26352]_ , \new_[26353]_ , \new_[26356]_ , \new_[26359]_ ,
    \new_[26360]_ , \new_[26361]_ , \new_[26365]_ , \new_[26366]_ ,
    \new_[26369]_ , \new_[26372]_ , \new_[26373]_ , \new_[26374]_ ,
    \new_[26378]_ , \new_[26379]_ , \new_[26382]_ , \new_[26385]_ ,
    \new_[26386]_ , \new_[26387]_ , \new_[26391]_ , \new_[26392]_ ,
    \new_[26395]_ , \new_[26398]_ , \new_[26399]_ , \new_[26400]_ ,
    \new_[26404]_ , \new_[26405]_ , \new_[26408]_ , \new_[26411]_ ,
    \new_[26412]_ , \new_[26413]_ , \new_[26417]_ , \new_[26418]_ ,
    \new_[26421]_ , \new_[26424]_ , \new_[26425]_ , \new_[26426]_ ,
    \new_[26430]_ , \new_[26431]_ , \new_[26434]_ , \new_[26437]_ ,
    \new_[26438]_ , \new_[26439]_ , \new_[26443]_ , \new_[26444]_ ,
    \new_[26447]_ , \new_[26450]_ , \new_[26451]_ , \new_[26452]_ ,
    \new_[26456]_ , \new_[26457]_ , \new_[26460]_ , \new_[26463]_ ,
    \new_[26464]_ , \new_[26465]_ , \new_[26469]_ , \new_[26470]_ ,
    \new_[26473]_ , \new_[26476]_ , \new_[26477]_ , \new_[26478]_ ,
    \new_[26482]_ , \new_[26483]_ , \new_[26486]_ , \new_[26489]_ ,
    \new_[26490]_ , \new_[26491]_ , \new_[26495]_ , \new_[26496]_ ,
    \new_[26499]_ , \new_[26502]_ , \new_[26503]_ , \new_[26504]_ ,
    \new_[26508]_ , \new_[26509]_ , \new_[26512]_ , \new_[26515]_ ,
    \new_[26516]_ , \new_[26517]_ , \new_[26521]_ , \new_[26522]_ ,
    \new_[26525]_ , \new_[26528]_ , \new_[26529]_ , \new_[26530]_ ,
    \new_[26534]_ , \new_[26535]_ , \new_[26538]_ , \new_[26541]_ ,
    \new_[26542]_ , \new_[26543]_ , \new_[26547]_ , \new_[26548]_ ,
    \new_[26551]_ , \new_[26554]_ , \new_[26555]_ , \new_[26556]_ ,
    \new_[26560]_ , \new_[26561]_ , \new_[26564]_ , \new_[26567]_ ,
    \new_[26568]_ , \new_[26569]_ , \new_[26573]_ , \new_[26574]_ ,
    \new_[26577]_ , \new_[26580]_ , \new_[26581]_ , \new_[26582]_ ,
    \new_[26586]_ , \new_[26587]_ , \new_[26590]_ , \new_[26593]_ ,
    \new_[26594]_ , \new_[26595]_ , \new_[26599]_ , \new_[26600]_ ,
    \new_[26603]_ , \new_[26606]_ , \new_[26607]_ , \new_[26608]_ ,
    \new_[26612]_ , \new_[26613]_ , \new_[26616]_ , \new_[26619]_ ,
    \new_[26620]_ , \new_[26621]_ , \new_[26625]_ , \new_[26626]_ ,
    \new_[26629]_ , \new_[26632]_ , \new_[26633]_ , \new_[26634]_ ,
    \new_[26638]_ , \new_[26639]_ , \new_[26642]_ , \new_[26645]_ ,
    \new_[26646]_ , \new_[26647]_ , \new_[26651]_ , \new_[26652]_ ,
    \new_[26655]_ , \new_[26658]_ , \new_[26659]_ , \new_[26660]_ ,
    \new_[26664]_ , \new_[26665]_ , \new_[26668]_ , \new_[26671]_ ,
    \new_[26672]_ , \new_[26673]_ , \new_[26677]_ , \new_[26678]_ ,
    \new_[26681]_ , \new_[26684]_ , \new_[26685]_ , \new_[26686]_ ,
    \new_[26690]_ , \new_[26691]_ , \new_[26694]_ , \new_[26697]_ ,
    \new_[26698]_ , \new_[26699]_ , \new_[26703]_ , \new_[26704]_ ,
    \new_[26707]_ , \new_[26710]_ , \new_[26711]_ , \new_[26712]_ ,
    \new_[26716]_ , \new_[26717]_ , \new_[26720]_ , \new_[26723]_ ,
    \new_[26724]_ , \new_[26725]_ , \new_[26729]_ , \new_[26730]_ ,
    \new_[26733]_ , \new_[26736]_ , \new_[26737]_ , \new_[26738]_ ,
    \new_[26742]_ , \new_[26743]_ , \new_[26746]_ , \new_[26749]_ ,
    \new_[26750]_ , \new_[26751]_ , \new_[26755]_ , \new_[26756]_ ,
    \new_[26759]_ , \new_[26762]_ , \new_[26763]_ , \new_[26764]_ ,
    \new_[26768]_ , \new_[26769]_ , \new_[26772]_ , \new_[26775]_ ,
    \new_[26776]_ , \new_[26777]_ , \new_[26781]_ , \new_[26782]_ ,
    \new_[26785]_ , \new_[26788]_ , \new_[26789]_ , \new_[26790]_ ,
    \new_[26794]_ , \new_[26795]_ , \new_[26798]_ , \new_[26801]_ ,
    \new_[26802]_ , \new_[26803]_ , \new_[26807]_ , \new_[26808]_ ,
    \new_[26811]_ , \new_[26814]_ , \new_[26815]_ , \new_[26816]_ ,
    \new_[26820]_ , \new_[26821]_ , \new_[26824]_ , \new_[26827]_ ,
    \new_[26828]_ , \new_[26829]_ , \new_[26833]_ , \new_[26834]_ ,
    \new_[26837]_ , \new_[26840]_ , \new_[26841]_ , \new_[26842]_ ,
    \new_[26846]_ , \new_[26847]_ , \new_[26850]_ , \new_[26853]_ ,
    \new_[26854]_ , \new_[26855]_ , \new_[26859]_ , \new_[26860]_ ,
    \new_[26863]_ , \new_[26866]_ , \new_[26867]_ , \new_[26868]_ ,
    \new_[26872]_ , \new_[26873]_ , \new_[26876]_ , \new_[26879]_ ,
    \new_[26880]_ , \new_[26881]_ , \new_[26885]_ , \new_[26886]_ ,
    \new_[26889]_ , \new_[26892]_ , \new_[26893]_ , \new_[26894]_ ,
    \new_[26898]_ , \new_[26899]_ , \new_[26902]_ , \new_[26905]_ ,
    \new_[26906]_ , \new_[26907]_ , \new_[26911]_ , \new_[26912]_ ,
    \new_[26915]_ , \new_[26918]_ , \new_[26919]_ , \new_[26920]_ ,
    \new_[26924]_ , \new_[26925]_ , \new_[26928]_ , \new_[26931]_ ,
    \new_[26932]_ , \new_[26933]_ , \new_[26937]_ , \new_[26938]_ ,
    \new_[26941]_ , \new_[26944]_ , \new_[26945]_ , \new_[26946]_ ,
    \new_[26950]_ , \new_[26951]_ , \new_[26954]_ , \new_[26957]_ ,
    \new_[26958]_ , \new_[26959]_ , \new_[26963]_ , \new_[26964]_ ,
    \new_[26967]_ , \new_[26970]_ , \new_[26971]_ , \new_[26972]_ ,
    \new_[26976]_ , \new_[26977]_ , \new_[26980]_ , \new_[26983]_ ,
    \new_[26984]_ , \new_[26985]_ , \new_[26989]_ , \new_[26990]_ ,
    \new_[26993]_ , \new_[26996]_ , \new_[26997]_ , \new_[26998]_ ,
    \new_[27002]_ , \new_[27003]_ , \new_[27006]_ , \new_[27009]_ ,
    \new_[27010]_ , \new_[27011]_ , \new_[27015]_ , \new_[27016]_ ,
    \new_[27019]_ , \new_[27022]_ , \new_[27023]_ , \new_[27024]_ ,
    \new_[27028]_ , \new_[27029]_ , \new_[27032]_ , \new_[27035]_ ,
    \new_[27036]_ , \new_[27037]_ , \new_[27041]_ , \new_[27042]_ ,
    \new_[27045]_ , \new_[27048]_ , \new_[27049]_ , \new_[27050]_ ,
    \new_[27054]_ , \new_[27055]_ , \new_[27058]_ , \new_[27061]_ ,
    \new_[27062]_ , \new_[27063]_ , \new_[27067]_ , \new_[27068]_ ,
    \new_[27071]_ , \new_[27074]_ , \new_[27075]_ , \new_[27076]_ ,
    \new_[27080]_ , \new_[27081]_ , \new_[27084]_ , \new_[27087]_ ,
    \new_[27088]_ , \new_[27089]_ , \new_[27093]_ , \new_[27094]_ ,
    \new_[27097]_ , \new_[27100]_ , \new_[27101]_ , \new_[27102]_ ,
    \new_[27106]_ , \new_[27107]_ , \new_[27110]_ , \new_[27113]_ ,
    \new_[27114]_ , \new_[27115]_ , \new_[27119]_ , \new_[27120]_ ,
    \new_[27123]_ , \new_[27126]_ , \new_[27127]_ , \new_[27128]_ ,
    \new_[27132]_ , \new_[27133]_ , \new_[27136]_ , \new_[27139]_ ,
    \new_[27140]_ , \new_[27141]_ , \new_[27145]_ , \new_[27146]_ ,
    \new_[27149]_ , \new_[27152]_ , \new_[27153]_ , \new_[27154]_ ,
    \new_[27158]_ , \new_[27159]_ , \new_[27162]_ , \new_[27165]_ ,
    \new_[27166]_ , \new_[27167]_ , \new_[27171]_ , \new_[27172]_ ,
    \new_[27175]_ , \new_[27178]_ , \new_[27179]_ , \new_[27180]_ ,
    \new_[27184]_ , \new_[27185]_ , \new_[27188]_ , \new_[27191]_ ,
    \new_[27192]_ , \new_[27193]_ , \new_[27197]_ , \new_[27198]_ ,
    \new_[27201]_ , \new_[27204]_ , \new_[27205]_ , \new_[27206]_ ,
    \new_[27210]_ , \new_[27211]_ , \new_[27214]_ , \new_[27217]_ ,
    \new_[27218]_ , \new_[27219]_ , \new_[27223]_ , \new_[27224]_ ,
    \new_[27227]_ , \new_[27230]_ , \new_[27231]_ , \new_[27232]_ ,
    \new_[27236]_ , \new_[27237]_ , \new_[27240]_ , \new_[27243]_ ,
    \new_[27244]_ , \new_[27245]_ , \new_[27249]_ , \new_[27250]_ ,
    \new_[27253]_ , \new_[27256]_ , \new_[27257]_ , \new_[27258]_ ,
    \new_[27262]_ , \new_[27263]_ , \new_[27266]_ , \new_[27269]_ ,
    \new_[27270]_ , \new_[27271]_ , \new_[27275]_ , \new_[27276]_ ,
    \new_[27279]_ , \new_[27282]_ , \new_[27283]_ , \new_[27284]_ ,
    \new_[27288]_ , \new_[27289]_ , \new_[27292]_ , \new_[27295]_ ,
    \new_[27296]_ , \new_[27297]_ , \new_[27301]_ , \new_[27302]_ ,
    \new_[27305]_ , \new_[27308]_ , \new_[27309]_ , \new_[27310]_ ,
    \new_[27314]_ , \new_[27315]_ , \new_[27318]_ , \new_[27321]_ ,
    \new_[27322]_ , \new_[27323]_ , \new_[27327]_ , \new_[27328]_ ,
    \new_[27331]_ , \new_[27334]_ , \new_[27335]_ , \new_[27336]_ ,
    \new_[27340]_ , \new_[27341]_ , \new_[27344]_ , \new_[27347]_ ,
    \new_[27348]_ , \new_[27349]_ , \new_[27353]_ , \new_[27354]_ ,
    \new_[27357]_ , \new_[27360]_ , \new_[27361]_ , \new_[27362]_ ,
    \new_[27366]_ , \new_[27367]_ , \new_[27370]_ , \new_[27373]_ ,
    \new_[27374]_ , \new_[27375]_ , \new_[27379]_ , \new_[27380]_ ,
    \new_[27383]_ , \new_[27386]_ , \new_[27387]_ , \new_[27388]_ ,
    \new_[27392]_ , \new_[27393]_ , \new_[27396]_ , \new_[27399]_ ,
    \new_[27400]_ , \new_[27401]_ , \new_[27405]_ , \new_[27406]_ ,
    \new_[27409]_ , \new_[27412]_ , \new_[27413]_ , \new_[27414]_ ,
    \new_[27418]_ , \new_[27419]_ , \new_[27422]_ , \new_[27425]_ ,
    \new_[27426]_ , \new_[27427]_ , \new_[27431]_ , \new_[27432]_ ,
    \new_[27435]_ , \new_[27438]_ , \new_[27439]_ , \new_[27440]_ ,
    \new_[27444]_ , \new_[27445]_ , \new_[27448]_ , \new_[27451]_ ,
    \new_[27452]_ , \new_[27453]_ , \new_[27457]_ , \new_[27458]_ ,
    \new_[27461]_ , \new_[27464]_ , \new_[27465]_ , \new_[27466]_ ,
    \new_[27470]_ , \new_[27471]_ , \new_[27474]_ , \new_[27477]_ ,
    \new_[27478]_ , \new_[27479]_ , \new_[27483]_ , \new_[27484]_ ,
    \new_[27487]_ , \new_[27490]_ , \new_[27491]_ , \new_[27492]_ ,
    \new_[27496]_ , \new_[27497]_ , \new_[27500]_ , \new_[27503]_ ,
    \new_[27504]_ , \new_[27505]_ , \new_[27509]_ , \new_[27510]_ ,
    \new_[27513]_ , \new_[27516]_ , \new_[27517]_ , \new_[27518]_ ,
    \new_[27522]_ , \new_[27523]_ , \new_[27526]_ , \new_[27529]_ ,
    \new_[27530]_ , \new_[27531]_ , \new_[27535]_ , \new_[27536]_ ,
    \new_[27539]_ , \new_[27542]_ , \new_[27543]_ , \new_[27544]_ ,
    \new_[27548]_ , \new_[27549]_ , \new_[27552]_ , \new_[27555]_ ,
    \new_[27556]_ , \new_[27557]_ , \new_[27561]_ , \new_[27562]_ ,
    \new_[27565]_ , \new_[27568]_ , \new_[27569]_ , \new_[27570]_ ,
    \new_[27574]_ , \new_[27575]_ , \new_[27578]_ , \new_[27581]_ ,
    \new_[27582]_ , \new_[27583]_ , \new_[27587]_ , \new_[27588]_ ,
    \new_[27591]_ , \new_[27594]_ , \new_[27595]_ , \new_[27596]_ ,
    \new_[27600]_ , \new_[27601]_ , \new_[27604]_ , \new_[27607]_ ,
    \new_[27608]_ , \new_[27609]_ , \new_[27613]_ , \new_[27614]_ ,
    \new_[27617]_ , \new_[27620]_ , \new_[27621]_ , \new_[27622]_ ,
    \new_[27626]_ , \new_[27627]_ , \new_[27630]_ , \new_[27633]_ ,
    \new_[27634]_ , \new_[27635]_ , \new_[27639]_ , \new_[27640]_ ,
    \new_[27643]_ , \new_[27646]_ , \new_[27647]_ , \new_[27648]_ ,
    \new_[27652]_ , \new_[27653]_ , \new_[27656]_ , \new_[27659]_ ,
    \new_[27660]_ , \new_[27661]_ , \new_[27665]_ , \new_[27666]_ ,
    \new_[27669]_ , \new_[27672]_ , \new_[27673]_ , \new_[27674]_ ,
    \new_[27678]_ , \new_[27679]_ , \new_[27682]_ , \new_[27685]_ ,
    \new_[27686]_ , \new_[27687]_ , \new_[27691]_ , \new_[27692]_ ,
    \new_[27695]_ , \new_[27698]_ , \new_[27699]_ , \new_[27700]_ ,
    \new_[27704]_ , \new_[27705]_ , \new_[27708]_ , \new_[27711]_ ,
    \new_[27712]_ , \new_[27713]_ , \new_[27717]_ , \new_[27718]_ ,
    \new_[27721]_ , \new_[27724]_ , \new_[27725]_ , \new_[27726]_ ,
    \new_[27730]_ , \new_[27731]_ , \new_[27734]_ , \new_[27737]_ ,
    \new_[27738]_ , \new_[27739]_ , \new_[27743]_ , \new_[27744]_ ,
    \new_[27747]_ , \new_[27750]_ , \new_[27751]_ , \new_[27752]_ ,
    \new_[27756]_ , \new_[27757]_ , \new_[27760]_ , \new_[27763]_ ,
    \new_[27764]_ , \new_[27765]_ , \new_[27769]_ , \new_[27770]_ ,
    \new_[27773]_ , \new_[27776]_ , \new_[27777]_ , \new_[27778]_ ,
    \new_[27782]_ , \new_[27783]_ , \new_[27786]_ , \new_[27789]_ ,
    \new_[27790]_ , \new_[27791]_ , \new_[27795]_ , \new_[27796]_ ,
    \new_[27799]_ , \new_[27802]_ , \new_[27803]_ , \new_[27804]_ ,
    \new_[27808]_ , \new_[27809]_ , \new_[27812]_ , \new_[27815]_ ,
    \new_[27816]_ , \new_[27817]_ , \new_[27821]_ , \new_[27822]_ ,
    \new_[27825]_ , \new_[27828]_ , \new_[27829]_ , \new_[27830]_ ,
    \new_[27834]_ , \new_[27835]_ , \new_[27838]_ , \new_[27841]_ ,
    \new_[27842]_ , \new_[27843]_ , \new_[27847]_ , \new_[27848]_ ,
    \new_[27851]_ , \new_[27854]_ , \new_[27855]_ , \new_[27856]_ ,
    \new_[27860]_ , \new_[27861]_ , \new_[27864]_ , \new_[27867]_ ,
    \new_[27868]_ , \new_[27869]_ , \new_[27873]_ , \new_[27874]_ ,
    \new_[27877]_ , \new_[27880]_ , \new_[27881]_ , \new_[27882]_ ,
    \new_[27886]_ , \new_[27887]_ , \new_[27890]_ , \new_[27893]_ ,
    \new_[27894]_ , \new_[27895]_ , \new_[27899]_ , \new_[27900]_ ,
    \new_[27903]_ , \new_[27906]_ , \new_[27907]_ , \new_[27908]_ ,
    \new_[27912]_ , \new_[27913]_ , \new_[27916]_ , \new_[27919]_ ,
    \new_[27920]_ , \new_[27921]_ , \new_[27925]_ , \new_[27926]_ ,
    \new_[27929]_ , \new_[27932]_ , \new_[27933]_ , \new_[27934]_ ,
    \new_[27938]_ , \new_[27939]_ , \new_[27942]_ , \new_[27945]_ ,
    \new_[27946]_ , \new_[27947]_ , \new_[27951]_ , \new_[27952]_ ,
    \new_[27955]_ , \new_[27958]_ , \new_[27959]_ , \new_[27960]_ ,
    \new_[27964]_ , \new_[27965]_ , \new_[27968]_ , \new_[27971]_ ,
    \new_[27972]_ , \new_[27973]_ , \new_[27977]_ , \new_[27978]_ ,
    \new_[27981]_ , \new_[27984]_ , \new_[27985]_ , \new_[27986]_ ,
    \new_[27990]_ , \new_[27991]_ , \new_[27994]_ , \new_[27997]_ ,
    \new_[27998]_ , \new_[27999]_ , \new_[28003]_ , \new_[28004]_ ,
    \new_[28007]_ , \new_[28010]_ , \new_[28011]_ , \new_[28012]_ ,
    \new_[28016]_ , \new_[28017]_ , \new_[28020]_ , \new_[28023]_ ,
    \new_[28024]_ , \new_[28025]_ , \new_[28029]_ , \new_[28030]_ ,
    \new_[28033]_ , \new_[28036]_ , \new_[28037]_ , \new_[28038]_ ,
    \new_[28042]_ , \new_[28043]_ , \new_[28046]_ , \new_[28049]_ ,
    \new_[28050]_ , \new_[28051]_ , \new_[28055]_ , \new_[28056]_ ,
    \new_[28059]_ , \new_[28062]_ , \new_[28063]_ , \new_[28064]_ ,
    \new_[28068]_ , \new_[28069]_ , \new_[28072]_ , \new_[28075]_ ,
    \new_[28076]_ , \new_[28077]_ , \new_[28081]_ , \new_[28082]_ ,
    \new_[28085]_ , \new_[28088]_ , \new_[28089]_ , \new_[28090]_ ,
    \new_[28094]_ , \new_[28095]_ , \new_[28098]_ , \new_[28101]_ ,
    \new_[28102]_ , \new_[28103]_ , \new_[28107]_ , \new_[28108]_ ,
    \new_[28111]_ , \new_[28114]_ , \new_[28115]_ , \new_[28116]_ ,
    \new_[28120]_ , \new_[28121]_ , \new_[28124]_ , \new_[28127]_ ,
    \new_[28128]_ , \new_[28129]_ , \new_[28133]_ , \new_[28134]_ ,
    \new_[28137]_ , \new_[28140]_ , \new_[28141]_ , \new_[28142]_ ,
    \new_[28146]_ , \new_[28147]_ , \new_[28150]_ , \new_[28153]_ ,
    \new_[28154]_ , \new_[28155]_ , \new_[28159]_ , \new_[28160]_ ,
    \new_[28163]_ , \new_[28166]_ , \new_[28167]_ , \new_[28168]_ ,
    \new_[28172]_ , \new_[28173]_ , \new_[28176]_ , \new_[28179]_ ,
    \new_[28180]_ , \new_[28181]_ , \new_[28185]_ , \new_[28186]_ ,
    \new_[28189]_ , \new_[28192]_ , \new_[28193]_ , \new_[28194]_ ,
    \new_[28198]_ , \new_[28199]_ , \new_[28202]_ , \new_[28205]_ ,
    \new_[28206]_ , \new_[28207]_ , \new_[28211]_ , \new_[28212]_ ,
    \new_[28215]_ , \new_[28218]_ , \new_[28219]_ , \new_[28220]_ ,
    \new_[28224]_ , \new_[28225]_ , \new_[28228]_ , \new_[28231]_ ,
    \new_[28232]_ , \new_[28233]_ , \new_[28237]_ , \new_[28238]_ ,
    \new_[28241]_ , \new_[28244]_ , \new_[28245]_ , \new_[28246]_ ,
    \new_[28250]_ , \new_[28251]_ , \new_[28254]_ , \new_[28257]_ ,
    \new_[28258]_ , \new_[28259]_ , \new_[28263]_ , \new_[28264]_ ,
    \new_[28267]_ , \new_[28270]_ , \new_[28271]_ , \new_[28272]_ ,
    \new_[28276]_ , \new_[28277]_ , \new_[28280]_ , \new_[28283]_ ,
    \new_[28284]_ , \new_[28285]_ , \new_[28289]_ , \new_[28290]_ ,
    \new_[28293]_ , \new_[28296]_ , \new_[28297]_ , \new_[28298]_ ,
    \new_[28302]_ , \new_[28303]_ , \new_[28306]_ , \new_[28309]_ ,
    \new_[28310]_ , \new_[28311]_ , \new_[28315]_ , \new_[28316]_ ,
    \new_[28319]_ , \new_[28322]_ , \new_[28323]_ , \new_[28324]_ ,
    \new_[28328]_ , \new_[28329]_ , \new_[28332]_ , \new_[28335]_ ,
    \new_[28336]_ , \new_[28337]_ , \new_[28341]_ , \new_[28342]_ ,
    \new_[28345]_ , \new_[28348]_ , \new_[28349]_ , \new_[28350]_ ,
    \new_[28354]_ , \new_[28355]_ , \new_[28358]_ , \new_[28361]_ ,
    \new_[28362]_ , \new_[28363]_ , \new_[28367]_ , \new_[28368]_ ,
    \new_[28371]_ , \new_[28374]_ , \new_[28375]_ , \new_[28376]_ ,
    \new_[28380]_ , \new_[28381]_ , \new_[28384]_ , \new_[28387]_ ,
    \new_[28388]_ , \new_[28389]_ , \new_[28393]_ , \new_[28394]_ ,
    \new_[28397]_ , \new_[28400]_ , \new_[28401]_ , \new_[28402]_ ,
    \new_[28406]_ , \new_[28407]_ , \new_[28410]_ , \new_[28413]_ ,
    \new_[28414]_ , \new_[28415]_ , \new_[28419]_ , \new_[28420]_ ,
    \new_[28423]_ , \new_[28426]_ , \new_[28427]_ , \new_[28428]_ ,
    \new_[28432]_ , \new_[28433]_ , \new_[28436]_ , \new_[28439]_ ,
    \new_[28440]_ , \new_[28441]_ , \new_[28445]_ , \new_[28446]_ ,
    \new_[28449]_ , \new_[28452]_ , \new_[28453]_ , \new_[28454]_ ,
    \new_[28458]_ , \new_[28459]_ , \new_[28462]_ , \new_[28465]_ ,
    \new_[28466]_ , \new_[28467]_ , \new_[28471]_ , \new_[28472]_ ,
    \new_[28475]_ , \new_[28478]_ , \new_[28479]_ , \new_[28480]_ ,
    \new_[28484]_ , \new_[28485]_ , \new_[28488]_ , \new_[28491]_ ,
    \new_[28492]_ , \new_[28493]_ , \new_[28497]_ , \new_[28498]_ ,
    \new_[28501]_ , \new_[28504]_ , \new_[28505]_ , \new_[28506]_ ,
    \new_[28510]_ , \new_[28511]_ , \new_[28514]_ , \new_[28517]_ ,
    \new_[28518]_ , \new_[28519]_ , \new_[28523]_ , \new_[28524]_ ,
    \new_[28527]_ , \new_[28530]_ , \new_[28531]_ , \new_[28532]_ ,
    \new_[28536]_ , \new_[28537]_ , \new_[28540]_ , \new_[28543]_ ,
    \new_[28544]_ , \new_[28545]_ , \new_[28549]_ , \new_[28550]_ ,
    \new_[28553]_ , \new_[28556]_ , \new_[28557]_ , \new_[28558]_ ,
    \new_[28562]_ , \new_[28563]_ , \new_[28566]_ , \new_[28569]_ ,
    \new_[28570]_ , \new_[28571]_ , \new_[28575]_ , \new_[28576]_ ,
    \new_[28579]_ , \new_[28582]_ , \new_[28583]_ , \new_[28584]_ ,
    \new_[28588]_ , \new_[28589]_ , \new_[28592]_ , \new_[28595]_ ,
    \new_[28596]_ , \new_[28597]_ , \new_[28601]_ , \new_[28602]_ ,
    \new_[28605]_ , \new_[28608]_ , \new_[28609]_ , \new_[28610]_ ,
    \new_[28614]_ , \new_[28615]_ , \new_[28618]_ , \new_[28621]_ ,
    \new_[28622]_ , \new_[28623]_ , \new_[28627]_ , \new_[28628]_ ,
    \new_[28631]_ , \new_[28634]_ , \new_[28635]_ , \new_[28636]_ ,
    \new_[28640]_ , \new_[28641]_ , \new_[28644]_ , \new_[28647]_ ,
    \new_[28648]_ , \new_[28649]_ , \new_[28653]_ , \new_[28654]_ ,
    \new_[28657]_ , \new_[28660]_ , \new_[28661]_ , \new_[28662]_ ,
    \new_[28666]_ , \new_[28667]_ , \new_[28670]_ , \new_[28673]_ ,
    \new_[28674]_ , \new_[28675]_ , \new_[28679]_ , \new_[28680]_ ,
    \new_[28683]_ , \new_[28686]_ , \new_[28687]_ , \new_[28688]_ ,
    \new_[28692]_ , \new_[28693]_ , \new_[28696]_ , \new_[28699]_ ,
    \new_[28700]_ , \new_[28701]_ , \new_[28705]_ , \new_[28706]_ ,
    \new_[28709]_ , \new_[28712]_ , \new_[28713]_ , \new_[28714]_ ,
    \new_[28718]_ , \new_[28719]_ , \new_[28722]_ , \new_[28725]_ ,
    \new_[28726]_ , \new_[28727]_ , \new_[28731]_ , \new_[28732]_ ,
    \new_[28735]_ , \new_[28738]_ , \new_[28739]_ , \new_[28740]_ ,
    \new_[28744]_ , \new_[28745]_ , \new_[28748]_ , \new_[28751]_ ,
    \new_[28752]_ , \new_[28753]_ , \new_[28757]_ , \new_[28758]_ ,
    \new_[28761]_ , \new_[28764]_ , \new_[28765]_ , \new_[28766]_ ,
    \new_[28770]_ , \new_[28771]_ , \new_[28774]_ , \new_[28777]_ ,
    \new_[28778]_ , \new_[28779]_ , \new_[28783]_ , \new_[28784]_ ,
    \new_[28787]_ , \new_[28790]_ , \new_[28791]_ , \new_[28792]_ ,
    \new_[28796]_ , \new_[28797]_ , \new_[28800]_ , \new_[28803]_ ,
    \new_[28804]_ , \new_[28805]_ , \new_[28809]_ , \new_[28810]_ ,
    \new_[28813]_ , \new_[28816]_ , \new_[28817]_ , \new_[28818]_ ,
    \new_[28822]_ , \new_[28823]_ , \new_[28826]_ , \new_[28829]_ ,
    \new_[28830]_ , \new_[28831]_ , \new_[28835]_ , \new_[28836]_ ,
    \new_[28839]_ , \new_[28842]_ , \new_[28843]_ , \new_[28844]_ ,
    \new_[28848]_ , \new_[28849]_ , \new_[28852]_ , \new_[28855]_ ,
    \new_[28856]_ , \new_[28857]_ , \new_[28861]_ , \new_[28862]_ ,
    \new_[28865]_ , \new_[28868]_ , \new_[28869]_ , \new_[28870]_ ,
    \new_[28874]_ , \new_[28875]_ , \new_[28878]_ , \new_[28881]_ ,
    \new_[28882]_ , \new_[28883]_ , \new_[28887]_ , \new_[28888]_ ,
    \new_[28891]_ , \new_[28894]_ , \new_[28895]_ , \new_[28896]_ ,
    \new_[28900]_ , \new_[28901]_ , \new_[28904]_ , \new_[28907]_ ,
    \new_[28908]_ , \new_[28909]_ , \new_[28913]_ , \new_[28914]_ ,
    \new_[28917]_ , \new_[28920]_ , \new_[28921]_ , \new_[28922]_ ,
    \new_[28926]_ , \new_[28927]_ , \new_[28930]_ , \new_[28933]_ ,
    \new_[28934]_ , \new_[28935]_ , \new_[28939]_ , \new_[28940]_ ,
    \new_[28943]_ , \new_[28946]_ , \new_[28947]_ , \new_[28948]_ ,
    \new_[28952]_ , \new_[28953]_ , \new_[28956]_ , \new_[28959]_ ,
    \new_[28960]_ , \new_[28961]_ , \new_[28965]_ , \new_[28966]_ ,
    \new_[28969]_ , \new_[28972]_ , \new_[28973]_ , \new_[28974]_ ,
    \new_[28978]_ , \new_[28979]_ , \new_[28982]_ , \new_[28985]_ ,
    \new_[28986]_ , \new_[28987]_ , \new_[28991]_ , \new_[28992]_ ,
    \new_[28995]_ , \new_[28998]_ , \new_[28999]_ , \new_[29000]_ ,
    \new_[29004]_ , \new_[29005]_ , \new_[29008]_ , \new_[29011]_ ,
    \new_[29012]_ , \new_[29013]_ , \new_[29017]_ , \new_[29018]_ ,
    \new_[29021]_ , \new_[29024]_ , \new_[29025]_ , \new_[29026]_ ,
    \new_[29030]_ , \new_[29031]_ , \new_[29034]_ , \new_[29037]_ ,
    \new_[29038]_ , \new_[29039]_ , \new_[29043]_ , \new_[29044]_ ,
    \new_[29047]_ , \new_[29050]_ , \new_[29051]_ , \new_[29052]_ ,
    \new_[29056]_ , \new_[29057]_ , \new_[29060]_ , \new_[29063]_ ,
    \new_[29064]_ , \new_[29065]_ , \new_[29069]_ , \new_[29070]_ ,
    \new_[29073]_ , \new_[29076]_ , \new_[29077]_ , \new_[29078]_ ,
    \new_[29082]_ , \new_[29083]_ , \new_[29086]_ , \new_[29089]_ ,
    \new_[29090]_ , \new_[29091]_ , \new_[29095]_ , \new_[29096]_ ,
    \new_[29099]_ , \new_[29102]_ , \new_[29103]_ , \new_[29104]_ ,
    \new_[29108]_ , \new_[29109]_ , \new_[29112]_ , \new_[29115]_ ,
    \new_[29116]_ , \new_[29117]_ , \new_[29121]_ , \new_[29122]_ ,
    \new_[29125]_ , \new_[29128]_ , \new_[29129]_ , \new_[29130]_ ,
    \new_[29134]_ , \new_[29135]_ , \new_[29138]_ , \new_[29141]_ ,
    \new_[29142]_ , \new_[29143]_ , \new_[29147]_ , \new_[29148]_ ,
    \new_[29151]_ , \new_[29154]_ , \new_[29155]_ , \new_[29156]_ ,
    \new_[29160]_ , \new_[29161]_ , \new_[29164]_ , \new_[29167]_ ,
    \new_[29168]_ , \new_[29169]_ , \new_[29173]_ , \new_[29174]_ ,
    \new_[29177]_ , \new_[29180]_ , \new_[29181]_ , \new_[29182]_ ,
    \new_[29186]_ , \new_[29187]_ , \new_[29190]_ , \new_[29193]_ ,
    \new_[29194]_ , \new_[29195]_ , \new_[29199]_ , \new_[29200]_ ,
    \new_[29203]_ , \new_[29206]_ , \new_[29207]_ , \new_[29208]_ ,
    \new_[29212]_ , \new_[29213]_ , \new_[29216]_ , \new_[29219]_ ,
    \new_[29220]_ , \new_[29221]_ , \new_[29225]_ , \new_[29226]_ ,
    \new_[29229]_ , \new_[29232]_ , \new_[29233]_ , \new_[29234]_ ,
    \new_[29238]_ , \new_[29239]_ , \new_[29242]_ , \new_[29245]_ ,
    \new_[29246]_ , \new_[29247]_ , \new_[29251]_ , \new_[29252]_ ,
    \new_[29255]_ , \new_[29258]_ , \new_[29259]_ , \new_[29260]_ ,
    \new_[29264]_ , \new_[29265]_ , \new_[29268]_ , \new_[29271]_ ,
    \new_[29272]_ , \new_[29273]_ , \new_[29277]_ , \new_[29278]_ ,
    \new_[29281]_ , \new_[29284]_ , \new_[29285]_ , \new_[29286]_ ,
    \new_[29290]_ , \new_[29291]_ , \new_[29294]_ , \new_[29297]_ ,
    \new_[29298]_ , \new_[29299]_ , \new_[29303]_ , \new_[29304]_ ,
    \new_[29307]_ , \new_[29310]_ , \new_[29311]_ , \new_[29312]_ ,
    \new_[29316]_ , \new_[29317]_ , \new_[29320]_ , \new_[29323]_ ,
    \new_[29324]_ , \new_[29325]_ , \new_[29329]_ , \new_[29330]_ ,
    \new_[29333]_ , \new_[29336]_ , \new_[29337]_ , \new_[29338]_ ,
    \new_[29342]_ , \new_[29343]_ , \new_[29346]_ , \new_[29349]_ ,
    \new_[29350]_ , \new_[29351]_ , \new_[29355]_ , \new_[29356]_ ,
    \new_[29359]_ , \new_[29362]_ , \new_[29363]_ , \new_[29364]_ ,
    \new_[29368]_ , \new_[29369]_ , \new_[29372]_ , \new_[29375]_ ,
    \new_[29376]_ , \new_[29377]_ , \new_[29381]_ , \new_[29382]_ ,
    \new_[29385]_ , \new_[29388]_ , \new_[29389]_ , \new_[29390]_ ,
    \new_[29394]_ , \new_[29395]_ , \new_[29398]_ , \new_[29401]_ ,
    \new_[29402]_ , \new_[29403]_ , \new_[29407]_ , \new_[29408]_ ,
    \new_[29411]_ , \new_[29414]_ , \new_[29415]_ , \new_[29416]_ ,
    \new_[29420]_ , \new_[29421]_ , \new_[29424]_ , \new_[29427]_ ,
    \new_[29428]_ , \new_[29429]_ , \new_[29433]_ , \new_[29434]_ ,
    \new_[29437]_ , \new_[29440]_ , \new_[29441]_ , \new_[29442]_ ,
    \new_[29446]_ , \new_[29447]_ , \new_[29450]_ , \new_[29453]_ ,
    \new_[29454]_ , \new_[29455]_ , \new_[29459]_ , \new_[29460]_ ,
    \new_[29463]_ , \new_[29466]_ , \new_[29467]_ , \new_[29468]_ ,
    \new_[29472]_ , \new_[29473]_ , \new_[29476]_ , \new_[29479]_ ,
    \new_[29480]_ , \new_[29481]_ , \new_[29485]_ , \new_[29486]_ ,
    \new_[29489]_ , \new_[29492]_ , \new_[29493]_ , \new_[29494]_ ,
    \new_[29498]_ , \new_[29499]_ , \new_[29502]_ , \new_[29505]_ ,
    \new_[29506]_ , \new_[29507]_ , \new_[29511]_ , \new_[29512]_ ,
    \new_[29515]_ , \new_[29518]_ , \new_[29519]_ , \new_[29520]_ ,
    \new_[29524]_ , \new_[29525]_ , \new_[29528]_ , \new_[29531]_ ,
    \new_[29532]_ , \new_[29533]_ , \new_[29537]_ , \new_[29538]_ ,
    \new_[29541]_ , \new_[29544]_ , \new_[29545]_ , \new_[29546]_ ,
    \new_[29550]_ , \new_[29551]_ , \new_[29554]_ , \new_[29557]_ ,
    \new_[29558]_ , \new_[29559]_ , \new_[29563]_ , \new_[29564]_ ,
    \new_[29567]_ , \new_[29570]_ , \new_[29571]_ , \new_[29572]_ ,
    \new_[29576]_ , \new_[29577]_ , \new_[29580]_ , \new_[29583]_ ,
    \new_[29584]_ , \new_[29585]_ , \new_[29589]_ , \new_[29590]_ ,
    \new_[29593]_ , \new_[29596]_ , \new_[29597]_ , \new_[29598]_ ,
    \new_[29602]_ , \new_[29603]_ , \new_[29606]_ , \new_[29609]_ ,
    \new_[29610]_ , \new_[29611]_ , \new_[29615]_ , \new_[29616]_ ,
    \new_[29619]_ , \new_[29622]_ , \new_[29623]_ , \new_[29624]_ ,
    \new_[29628]_ , \new_[29629]_ , \new_[29632]_ , \new_[29635]_ ,
    \new_[29636]_ , \new_[29637]_ , \new_[29641]_ , \new_[29642]_ ,
    \new_[29645]_ , \new_[29648]_ , \new_[29649]_ , \new_[29650]_ ,
    \new_[29654]_ , \new_[29655]_ , \new_[29658]_ , \new_[29661]_ ,
    \new_[29662]_ , \new_[29663]_ , \new_[29667]_ , \new_[29668]_ ,
    \new_[29671]_ , \new_[29674]_ , \new_[29675]_ , \new_[29676]_ ,
    \new_[29680]_ , \new_[29681]_ , \new_[29684]_ , \new_[29687]_ ,
    \new_[29688]_ , \new_[29689]_ , \new_[29693]_ , \new_[29694]_ ,
    \new_[29697]_ , \new_[29700]_ , \new_[29701]_ , \new_[29702]_ ,
    \new_[29706]_ , \new_[29707]_ , \new_[29710]_ , \new_[29713]_ ,
    \new_[29714]_ , \new_[29715]_ , \new_[29719]_ , \new_[29720]_ ,
    \new_[29723]_ , \new_[29726]_ , \new_[29727]_ , \new_[29728]_ ,
    \new_[29732]_ , \new_[29733]_ , \new_[29736]_ , \new_[29739]_ ,
    \new_[29740]_ , \new_[29741]_ , \new_[29745]_ , \new_[29746]_ ,
    \new_[29749]_ , \new_[29752]_ , \new_[29753]_ , \new_[29754]_ ,
    \new_[29758]_ , \new_[29759]_ , \new_[29762]_ , \new_[29765]_ ,
    \new_[29766]_ , \new_[29767]_ , \new_[29771]_ , \new_[29772]_ ,
    \new_[29775]_ , \new_[29778]_ , \new_[29779]_ , \new_[29780]_ ,
    \new_[29784]_ , \new_[29785]_ , \new_[29788]_ , \new_[29791]_ ,
    \new_[29792]_ , \new_[29793]_ , \new_[29797]_ , \new_[29798]_ ,
    \new_[29801]_ , \new_[29804]_ , \new_[29805]_ , \new_[29806]_ ,
    \new_[29810]_ , \new_[29811]_ , \new_[29814]_ , \new_[29817]_ ,
    \new_[29818]_ , \new_[29819]_ , \new_[29823]_ , \new_[29824]_ ,
    \new_[29827]_ , \new_[29830]_ , \new_[29831]_ , \new_[29832]_ ,
    \new_[29836]_ , \new_[29837]_ , \new_[29840]_ , \new_[29843]_ ,
    \new_[29844]_ , \new_[29845]_ , \new_[29849]_ , \new_[29850]_ ,
    \new_[29853]_ , \new_[29856]_ , \new_[29857]_ , \new_[29858]_ ,
    \new_[29862]_ , \new_[29863]_ , \new_[29866]_ , \new_[29869]_ ,
    \new_[29870]_ , \new_[29871]_ , \new_[29875]_ , \new_[29876]_ ,
    \new_[29879]_ , \new_[29882]_ , \new_[29883]_ , \new_[29884]_ ,
    \new_[29888]_ , \new_[29889]_ , \new_[29892]_ , \new_[29895]_ ,
    \new_[29896]_ , \new_[29897]_ , \new_[29901]_ , \new_[29902]_ ,
    \new_[29905]_ , \new_[29908]_ , \new_[29909]_ , \new_[29910]_ ,
    \new_[29914]_ , \new_[29915]_ , \new_[29918]_ , \new_[29921]_ ,
    \new_[29922]_ , \new_[29923]_ , \new_[29927]_ , \new_[29928]_ ,
    \new_[29931]_ , \new_[29934]_ , \new_[29935]_ , \new_[29936]_ ,
    \new_[29940]_ , \new_[29941]_ , \new_[29944]_ , \new_[29947]_ ,
    \new_[29948]_ , \new_[29949]_ , \new_[29953]_ , \new_[29954]_ ,
    \new_[29957]_ , \new_[29960]_ , \new_[29961]_ , \new_[29962]_ ,
    \new_[29966]_ , \new_[29967]_ , \new_[29970]_ , \new_[29973]_ ,
    \new_[29974]_ , \new_[29975]_ , \new_[29979]_ , \new_[29980]_ ,
    \new_[29983]_ , \new_[29986]_ , \new_[29987]_ , \new_[29988]_ ,
    \new_[29992]_ , \new_[29993]_ , \new_[29996]_ , \new_[29999]_ ,
    \new_[30000]_ , \new_[30001]_ , \new_[30005]_ , \new_[30006]_ ,
    \new_[30009]_ , \new_[30012]_ , \new_[30013]_ , \new_[30014]_ ,
    \new_[30018]_ , \new_[30019]_ , \new_[30022]_ , \new_[30025]_ ,
    \new_[30026]_ , \new_[30027]_ , \new_[30031]_ , \new_[30032]_ ,
    \new_[30035]_ , \new_[30038]_ , \new_[30039]_ , \new_[30040]_ ,
    \new_[30044]_ , \new_[30045]_ , \new_[30048]_ , \new_[30051]_ ,
    \new_[30052]_ , \new_[30053]_ , \new_[30057]_ , \new_[30058]_ ,
    \new_[30061]_ , \new_[30064]_ , \new_[30065]_ , \new_[30066]_ ,
    \new_[30070]_ , \new_[30071]_ , \new_[30074]_ , \new_[30077]_ ,
    \new_[30078]_ , \new_[30079]_ , \new_[30083]_ , \new_[30084]_ ,
    \new_[30087]_ , \new_[30090]_ , \new_[30091]_ , \new_[30092]_ ,
    \new_[30096]_ , \new_[30097]_ , \new_[30100]_ , \new_[30103]_ ,
    \new_[30104]_ , \new_[30105]_ , \new_[30109]_ , \new_[30110]_ ,
    \new_[30113]_ , \new_[30116]_ , \new_[30117]_ , \new_[30118]_ ,
    \new_[30122]_ , \new_[30123]_ , \new_[30126]_ , \new_[30129]_ ,
    \new_[30130]_ , \new_[30131]_ , \new_[30135]_ , \new_[30136]_ ,
    \new_[30139]_ , \new_[30142]_ , \new_[30143]_ , \new_[30144]_ ,
    \new_[30148]_ , \new_[30149]_ , \new_[30152]_ , \new_[30155]_ ,
    \new_[30156]_ , \new_[30157]_ , \new_[30161]_ , \new_[30162]_ ,
    \new_[30165]_ , \new_[30168]_ , \new_[30169]_ , \new_[30170]_ ,
    \new_[30174]_ , \new_[30175]_ , \new_[30178]_ , \new_[30181]_ ,
    \new_[30182]_ , \new_[30183]_ , \new_[30187]_ , \new_[30188]_ ,
    \new_[30191]_ , \new_[30194]_ , \new_[30195]_ , \new_[30196]_ ,
    \new_[30200]_ , \new_[30201]_ , \new_[30204]_ , \new_[30207]_ ,
    \new_[30208]_ , \new_[30209]_ , \new_[30213]_ , \new_[30214]_ ,
    \new_[30217]_ , \new_[30220]_ , \new_[30221]_ , \new_[30222]_ ,
    \new_[30226]_ , \new_[30227]_ , \new_[30230]_ , \new_[30233]_ ,
    \new_[30234]_ , \new_[30235]_ , \new_[30239]_ , \new_[30240]_ ,
    \new_[30243]_ , \new_[30246]_ , \new_[30247]_ , \new_[30248]_ ,
    \new_[30252]_ , \new_[30253]_ , \new_[30256]_ , \new_[30259]_ ,
    \new_[30260]_ , \new_[30261]_ , \new_[30265]_ , \new_[30266]_ ,
    \new_[30269]_ , \new_[30272]_ , \new_[30273]_ , \new_[30274]_ ,
    \new_[30278]_ , \new_[30279]_ , \new_[30282]_ , \new_[30285]_ ,
    \new_[30286]_ , \new_[30287]_ , \new_[30291]_ , \new_[30292]_ ,
    \new_[30295]_ , \new_[30298]_ , \new_[30299]_ , \new_[30300]_ ,
    \new_[30304]_ , \new_[30305]_ , \new_[30308]_ , \new_[30311]_ ,
    \new_[30312]_ , \new_[30313]_ , \new_[30317]_ , \new_[30318]_ ,
    \new_[30321]_ , \new_[30324]_ , \new_[30325]_ , \new_[30326]_ ,
    \new_[30330]_ , \new_[30331]_ , \new_[30334]_ , \new_[30337]_ ,
    \new_[30338]_ , \new_[30339]_ , \new_[30343]_ , \new_[30344]_ ,
    \new_[30347]_ , \new_[30350]_ , \new_[30351]_ , \new_[30352]_ ,
    \new_[30356]_ , \new_[30357]_ , \new_[30360]_ , \new_[30363]_ ,
    \new_[30364]_ , \new_[30365]_ , \new_[30369]_ , \new_[30370]_ ,
    \new_[30373]_ , \new_[30376]_ , \new_[30377]_ , \new_[30378]_ ,
    \new_[30382]_ , \new_[30383]_ , \new_[30386]_ , \new_[30389]_ ,
    \new_[30390]_ , \new_[30391]_ , \new_[30395]_ , \new_[30396]_ ,
    \new_[30399]_ , \new_[30402]_ , \new_[30403]_ , \new_[30404]_ ,
    \new_[30408]_ , \new_[30409]_ , \new_[30412]_ , \new_[30415]_ ,
    \new_[30416]_ , \new_[30417]_ , \new_[30421]_ , \new_[30422]_ ,
    \new_[30425]_ , \new_[30428]_ , \new_[30429]_ , \new_[30430]_ ,
    \new_[30434]_ , \new_[30435]_ , \new_[30438]_ , \new_[30441]_ ,
    \new_[30442]_ , \new_[30443]_ , \new_[30447]_ , \new_[30448]_ ,
    \new_[30451]_ , \new_[30454]_ , \new_[30455]_ , \new_[30456]_ ,
    \new_[30460]_ , \new_[30461]_ , \new_[30464]_ , \new_[30467]_ ,
    \new_[30468]_ , \new_[30469]_ , \new_[30473]_ , \new_[30474]_ ,
    \new_[30477]_ , \new_[30480]_ , \new_[30481]_ , \new_[30482]_ ,
    \new_[30486]_ , \new_[30487]_ , \new_[30490]_ , \new_[30493]_ ,
    \new_[30494]_ , \new_[30495]_ , \new_[30499]_ , \new_[30500]_ ,
    \new_[30503]_ , \new_[30506]_ , \new_[30507]_ , \new_[30508]_ ,
    \new_[30512]_ , \new_[30513]_ , \new_[30516]_ , \new_[30519]_ ,
    \new_[30520]_ , \new_[30521]_ , \new_[30525]_ , \new_[30526]_ ,
    \new_[30529]_ , \new_[30532]_ , \new_[30533]_ , \new_[30534]_ ,
    \new_[30538]_ , \new_[30539]_ , \new_[30542]_ , \new_[30545]_ ,
    \new_[30546]_ , \new_[30547]_ , \new_[30551]_ , \new_[30552]_ ,
    \new_[30555]_ , \new_[30558]_ , \new_[30559]_ , \new_[30560]_ ,
    \new_[30564]_ , \new_[30565]_ , \new_[30568]_ , \new_[30571]_ ,
    \new_[30572]_ , \new_[30573]_ , \new_[30577]_ , \new_[30578]_ ,
    \new_[30581]_ , \new_[30584]_ , \new_[30585]_ , \new_[30586]_ ,
    \new_[30590]_ , \new_[30591]_ , \new_[30594]_ , \new_[30597]_ ,
    \new_[30598]_ , \new_[30599]_ , \new_[30603]_ , \new_[30604]_ ,
    \new_[30607]_ , \new_[30610]_ , \new_[30611]_ , \new_[30612]_ ,
    \new_[30616]_ , \new_[30617]_ , \new_[30620]_ , \new_[30623]_ ,
    \new_[30624]_ , \new_[30625]_ , \new_[30629]_ , \new_[30630]_ ,
    \new_[30633]_ , \new_[30636]_ , \new_[30637]_ , \new_[30638]_ ,
    \new_[30642]_ , \new_[30643]_ , \new_[30646]_ , \new_[30649]_ ,
    \new_[30650]_ , \new_[30651]_ , \new_[30655]_ , \new_[30656]_ ,
    \new_[30659]_ , \new_[30662]_ , \new_[30663]_ , \new_[30664]_ ,
    \new_[30668]_ , \new_[30669]_ , \new_[30672]_ , \new_[30675]_ ,
    \new_[30676]_ , \new_[30677]_ , \new_[30681]_ , \new_[30682]_ ,
    \new_[30685]_ , \new_[30688]_ , \new_[30689]_ , \new_[30690]_ ,
    \new_[30694]_ , \new_[30695]_ , \new_[30698]_ , \new_[30701]_ ,
    \new_[30702]_ , \new_[30703]_ , \new_[30707]_ , \new_[30708]_ ,
    \new_[30711]_ , \new_[30714]_ , \new_[30715]_ , \new_[30716]_ ,
    \new_[30720]_ , \new_[30721]_ , \new_[30724]_ , \new_[30727]_ ,
    \new_[30728]_ , \new_[30729]_ , \new_[30733]_ , \new_[30734]_ ,
    \new_[30737]_ , \new_[30740]_ , \new_[30741]_ , \new_[30742]_ ,
    \new_[30746]_ , \new_[30747]_ , \new_[30750]_ , \new_[30753]_ ,
    \new_[30754]_ , \new_[30755]_ , \new_[30759]_ , \new_[30760]_ ,
    \new_[30763]_ , \new_[30766]_ , \new_[30767]_ , \new_[30768]_ ,
    \new_[30772]_ , \new_[30773]_ , \new_[30776]_ , \new_[30779]_ ,
    \new_[30780]_ , \new_[30781]_ , \new_[30785]_ , \new_[30786]_ ,
    \new_[30789]_ , \new_[30792]_ , \new_[30793]_ , \new_[30794]_ ,
    \new_[30798]_ , \new_[30799]_ , \new_[30802]_ , \new_[30805]_ ,
    \new_[30806]_ , \new_[30807]_ , \new_[30811]_ , \new_[30812]_ ,
    \new_[30815]_ , \new_[30818]_ , \new_[30819]_ , \new_[30820]_ ,
    \new_[30824]_ , \new_[30825]_ , \new_[30828]_ , \new_[30831]_ ,
    \new_[30832]_ , \new_[30833]_ , \new_[30837]_ , \new_[30838]_ ,
    \new_[30841]_ , \new_[30844]_ , \new_[30845]_ , \new_[30846]_ ,
    \new_[30850]_ , \new_[30851]_ , \new_[30854]_ , \new_[30857]_ ,
    \new_[30858]_ , \new_[30859]_ , \new_[30863]_ , \new_[30864]_ ,
    \new_[30867]_ , \new_[30870]_ , \new_[30871]_ , \new_[30872]_ ,
    \new_[30876]_ , \new_[30877]_ , \new_[30880]_ , \new_[30883]_ ,
    \new_[30884]_ , \new_[30885]_ , \new_[30889]_ , \new_[30890]_ ,
    \new_[30893]_ , \new_[30896]_ , \new_[30897]_ , \new_[30898]_ ,
    \new_[30902]_ , \new_[30903]_ , \new_[30906]_ , \new_[30909]_ ,
    \new_[30910]_ , \new_[30911]_ , \new_[30915]_ , \new_[30916]_ ,
    \new_[30919]_ , \new_[30922]_ , \new_[30923]_ , \new_[30924]_ ,
    \new_[30928]_ , \new_[30929]_ , \new_[30932]_ , \new_[30935]_ ,
    \new_[30936]_ , \new_[30937]_ , \new_[30941]_ , \new_[30942]_ ,
    \new_[30945]_ , \new_[30948]_ , \new_[30949]_ , \new_[30950]_ ,
    \new_[30954]_ , \new_[30955]_ , \new_[30958]_ , \new_[30961]_ ,
    \new_[30962]_ , \new_[30963]_ , \new_[30967]_ , \new_[30968]_ ,
    \new_[30971]_ , \new_[30974]_ , \new_[30975]_ , \new_[30976]_ ,
    \new_[30980]_ , \new_[30981]_ , \new_[30984]_ , \new_[30987]_ ,
    \new_[30988]_ , \new_[30989]_ , \new_[30993]_ , \new_[30994]_ ,
    \new_[30997]_ , \new_[31000]_ , \new_[31001]_ , \new_[31002]_ ,
    \new_[31006]_ , \new_[31007]_ , \new_[31010]_ , \new_[31013]_ ,
    \new_[31014]_ , \new_[31015]_ , \new_[31019]_ , \new_[31020]_ ,
    \new_[31023]_ , \new_[31026]_ , \new_[31027]_ , \new_[31028]_ ,
    \new_[31032]_ , \new_[31033]_ , \new_[31036]_ , \new_[31039]_ ,
    \new_[31040]_ , \new_[31041]_ , \new_[31045]_ , \new_[31046]_ ,
    \new_[31049]_ , \new_[31052]_ , \new_[31053]_ , \new_[31054]_ ,
    \new_[31058]_ , \new_[31059]_ , \new_[31062]_ , \new_[31065]_ ,
    \new_[31066]_ , \new_[31067]_ , \new_[31071]_ , \new_[31072]_ ,
    \new_[31075]_ , \new_[31078]_ , \new_[31079]_ , \new_[31080]_ ,
    \new_[31084]_ , \new_[31085]_ , \new_[31088]_ , \new_[31091]_ ,
    \new_[31092]_ , \new_[31093]_ , \new_[31097]_ , \new_[31098]_ ,
    \new_[31101]_ , \new_[31104]_ , \new_[31105]_ , \new_[31106]_ ,
    \new_[31110]_ , \new_[31111]_ , \new_[31114]_ , \new_[31117]_ ,
    \new_[31118]_ , \new_[31119]_ , \new_[31123]_ , \new_[31124]_ ,
    \new_[31127]_ , \new_[31130]_ , \new_[31131]_ , \new_[31132]_ ,
    \new_[31136]_ , \new_[31137]_ , \new_[31140]_ , \new_[31143]_ ,
    \new_[31144]_ , \new_[31145]_ , \new_[31149]_ , \new_[31150]_ ,
    \new_[31153]_ , \new_[31156]_ , \new_[31157]_ , \new_[31158]_ ,
    \new_[31162]_ , \new_[31163]_ , \new_[31166]_ , \new_[31169]_ ,
    \new_[31170]_ , \new_[31171]_ , \new_[31175]_ , \new_[31176]_ ,
    \new_[31179]_ , \new_[31182]_ , \new_[31183]_ , \new_[31184]_ ,
    \new_[31188]_ , \new_[31189]_ , \new_[31192]_ , \new_[31195]_ ,
    \new_[31196]_ , \new_[31197]_ , \new_[31201]_ , \new_[31202]_ ,
    \new_[31205]_ , \new_[31208]_ , \new_[31209]_ , \new_[31210]_ ,
    \new_[31214]_ , \new_[31215]_ , \new_[31218]_ , \new_[31221]_ ,
    \new_[31222]_ , \new_[31223]_ , \new_[31227]_ , \new_[31228]_ ,
    \new_[31231]_ , \new_[31234]_ , \new_[31235]_ , \new_[31236]_ ,
    \new_[31240]_ , \new_[31241]_ , \new_[31244]_ , \new_[31247]_ ,
    \new_[31248]_ , \new_[31249]_ , \new_[31253]_ , \new_[31254]_ ,
    \new_[31257]_ , \new_[31260]_ , \new_[31261]_ , \new_[31262]_ ,
    \new_[31266]_ , \new_[31267]_ , \new_[31270]_ , \new_[31273]_ ,
    \new_[31274]_ , \new_[31275]_ , \new_[31279]_ , \new_[31280]_ ,
    \new_[31283]_ , \new_[31286]_ , \new_[31287]_ , \new_[31288]_ ,
    \new_[31292]_ , \new_[31293]_ , \new_[31296]_ , \new_[31299]_ ,
    \new_[31300]_ , \new_[31301]_ , \new_[31305]_ , \new_[31306]_ ,
    \new_[31309]_ , \new_[31312]_ , \new_[31313]_ , \new_[31314]_ ,
    \new_[31318]_ , \new_[31319]_ , \new_[31322]_ , \new_[31325]_ ,
    \new_[31326]_ , \new_[31327]_ , \new_[31331]_ , \new_[31332]_ ,
    \new_[31335]_ , \new_[31338]_ , \new_[31339]_ , \new_[31340]_ ,
    \new_[31344]_ , \new_[31345]_ , \new_[31348]_ , \new_[31351]_ ,
    \new_[31352]_ , \new_[31353]_ , \new_[31357]_ , \new_[31358]_ ,
    \new_[31361]_ , \new_[31364]_ , \new_[31365]_ , \new_[31366]_ ,
    \new_[31370]_ , \new_[31371]_ , \new_[31374]_ , \new_[31377]_ ,
    \new_[31378]_ , \new_[31379]_ , \new_[31383]_ , \new_[31384]_ ,
    \new_[31387]_ , \new_[31390]_ , \new_[31391]_ , \new_[31392]_ ,
    \new_[31396]_ , \new_[31397]_ , \new_[31400]_ , \new_[31403]_ ,
    \new_[31404]_ , \new_[31405]_ , \new_[31409]_ , \new_[31410]_ ,
    \new_[31413]_ , \new_[31416]_ , \new_[31417]_ , \new_[31418]_ ,
    \new_[31422]_ , \new_[31423]_ , \new_[31426]_ , \new_[31429]_ ,
    \new_[31430]_ , \new_[31431]_ , \new_[31435]_ , \new_[31436]_ ,
    \new_[31439]_ , \new_[31442]_ , \new_[31443]_ , \new_[31444]_ ,
    \new_[31448]_ , \new_[31449]_ , \new_[31452]_ , \new_[31455]_ ,
    \new_[31456]_ , \new_[31457]_ , \new_[31461]_ , \new_[31462]_ ,
    \new_[31465]_ , \new_[31468]_ , \new_[31469]_ , \new_[31470]_ ,
    \new_[31474]_ , \new_[31475]_ , \new_[31478]_ , \new_[31481]_ ,
    \new_[31482]_ , \new_[31483]_ , \new_[31487]_ , \new_[31488]_ ,
    \new_[31491]_ , \new_[31494]_ , \new_[31495]_ , \new_[31496]_ ,
    \new_[31500]_ , \new_[31501]_ , \new_[31504]_ , \new_[31507]_ ,
    \new_[31508]_ , \new_[31509]_ , \new_[31513]_ , \new_[31514]_ ,
    \new_[31517]_ , \new_[31520]_ , \new_[31521]_ , \new_[31522]_ ,
    \new_[31526]_ , \new_[31527]_ , \new_[31530]_ , \new_[31533]_ ,
    \new_[31534]_ , \new_[31535]_ , \new_[31539]_ , \new_[31540]_ ,
    \new_[31543]_ , \new_[31546]_ , \new_[31547]_ , \new_[31548]_ ,
    \new_[31552]_ , \new_[31553]_ , \new_[31556]_ , \new_[31559]_ ,
    \new_[31560]_ , \new_[31561]_ , \new_[31565]_ , \new_[31566]_ ,
    \new_[31569]_ , \new_[31572]_ , \new_[31573]_ , \new_[31574]_ ,
    \new_[31578]_ , \new_[31579]_ , \new_[31582]_ , \new_[31585]_ ,
    \new_[31586]_ , \new_[31587]_ , \new_[31591]_ , \new_[31592]_ ,
    \new_[31595]_ , \new_[31598]_ , \new_[31599]_ , \new_[31600]_ ,
    \new_[31604]_ , \new_[31605]_ , \new_[31608]_ , \new_[31611]_ ,
    \new_[31612]_ , \new_[31613]_ , \new_[31617]_ , \new_[31618]_ ,
    \new_[31621]_ , \new_[31624]_ , \new_[31625]_ , \new_[31626]_ ,
    \new_[31630]_ , \new_[31631]_ , \new_[31634]_ , \new_[31637]_ ,
    \new_[31638]_ , \new_[31639]_ , \new_[31643]_ , \new_[31644]_ ,
    \new_[31647]_ , \new_[31650]_ , \new_[31651]_ , \new_[31652]_ ,
    \new_[31656]_ , \new_[31657]_ , \new_[31660]_ , \new_[31663]_ ,
    \new_[31664]_ , \new_[31665]_ , \new_[31669]_ , \new_[31670]_ ,
    \new_[31673]_ , \new_[31676]_ , \new_[31677]_ , \new_[31678]_ ,
    \new_[31682]_ , \new_[31683]_ , \new_[31686]_ , \new_[31689]_ ,
    \new_[31690]_ , \new_[31691]_ , \new_[31695]_ , \new_[31696]_ ,
    \new_[31699]_ , \new_[31702]_ , \new_[31703]_ , \new_[31704]_ ,
    \new_[31708]_ , \new_[31709]_ , \new_[31712]_ , \new_[31715]_ ,
    \new_[31716]_ , \new_[31717]_ , \new_[31721]_ , \new_[31722]_ ,
    \new_[31725]_ , \new_[31728]_ , \new_[31729]_ , \new_[31730]_ ,
    \new_[31734]_ , \new_[31735]_ , \new_[31738]_ , \new_[31741]_ ,
    \new_[31742]_ , \new_[31743]_ , \new_[31747]_ , \new_[31748]_ ,
    \new_[31751]_ , \new_[31754]_ , \new_[31755]_ , \new_[31756]_ ,
    \new_[31760]_ , \new_[31761]_ , \new_[31764]_ , \new_[31767]_ ,
    \new_[31768]_ , \new_[31769]_ , \new_[31773]_ , \new_[31774]_ ,
    \new_[31777]_ , \new_[31780]_ , \new_[31781]_ , \new_[31782]_ ,
    \new_[31786]_ , \new_[31787]_ , \new_[31790]_ , \new_[31793]_ ,
    \new_[31794]_ , \new_[31795]_ , \new_[31799]_ , \new_[31800]_ ,
    \new_[31803]_ , \new_[31806]_ , \new_[31807]_ , \new_[31808]_ ,
    \new_[31812]_ , \new_[31813]_ , \new_[31816]_ , \new_[31819]_ ,
    \new_[31820]_ , \new_[31821]_ , \new_[31825]_ , \new_[31826]_ ,
    \new_[31829]_ , \new_[31832]_ , \new_[31833]_ , \new_[31834]_ ,
    \new_[31838]_ , \new_[31839]_ , \new_[31842]_ , \new_[31845]_ ,
    \new_[31846]_ , \new_[31847]_ , \new_[31851]_ , \new_[31852]_ ,
    \new_[31855]_ , \new_[31858]_ , \new_[31859]_ , \new_[31860]_ ,
    \new_[31864]_ , \new_[31865]_ , \new_[31868]_ , \new_[31871]_ ,
    \new_[31872]_ , \new_[31873]_ , \new_[31877]_ , \new_[31878]_ ,
    \new_[31881]_ , \new_[31884]_ , \new_[31885]_ , \new_[31886]_ ,
    \new_[31890]_ , \new_[31891]_ , \new_[31894]_ , \new_[31897]_ ,
    \new_[31898]_ , \new_[31899]_ , \new_[31903]_ , \new_[31904]_ ,
    \new_[31907]_ , \new_[31910]_ , \new_[31911]_ , \new_[31912]_ ,
    \new_[31916]_ , \new_[31917]_ , \new_[31920]_ , \new_[31923]_ ,
    \new_[31924]_ , \new_[31925]_ , \new_[31929]_ , \new_[31930]_ ,
    \new_[31933]_ , \new_[31936]_ , \new_[31937]_ , \new_[31938]_ ,
    \new_[31942]_ , \new_[31943]_ , \new_[31946]_ , \new_[31949]_ ,
    \new_[31950]_ , \new_[31951]_ , \new_[31955]_ , \new_[31956]_ ,
    \new_[31959]_ , \new_[31962]_ , \new_[31963]_ , \new_[31964]_ ,
    \new_[31968]_ , \new_[31969]_ , \new_[31972]_ , \new_[31975]_ ,
    \new_[31976]_ , \new_[31977]_ , \new_[31981]_ , \new_[31982]_ ,
    \new_[31985]_ , \new_[31988]_ , \new_[31989]_ , \new_[31990]_ ,
    \new_[31994]_ , \new_[31995]_ , \new_[31998]_ , \new_[32001]_ ,
    \new_[32002]_ , \new_[32003]_ , \new_[32007]_ , \new_[32008]_ ,
    \new_[32011]_ , \new_[32014]_ , \new_[32015]_ , \new_[32016]_ ,
    \new_[32020]_ , \new_[32021]_ , \new_[32024]_ , \new_[32027]_ ,
    \new_[32028]_ , \new_[32029]_ , \new_[32033]_ , \new_[32034]_ ,
    \new_[32037]_ , \new_[32040]_ , \new_[32041]_ , \new_[32042]_ ,
    \new_[32046]_ , \new_[32047]_ , \new_[32050]_ , \new_[32053]_ ,
    \new_[32054]_ , \new_[32055]_ , \new_[32059]_ , \new_[32060]_ ,
    \new_[32063]_ , \new_[32066]_ , \new_[32067]_ , \new_[32068]_ ,
    \new_[32072]_ , \new_[32073]_ , \new_[32076]_ , \new_[32079]_ ,
    \new_[32080]_ , \new_[32081]_ , \new_[32085]_ , \new_[32086]_ ,
    \new_[32089]_ , \new_[32092]_ , \new_[32093]_ , \new_[32094]_ ,
    \new_[32098]_ , \new_[32099]_ , \new_[32102]_ , \new_[32105]_ ,
    \new_[32106]_ , \new_[32107]_ , \new_[32111]_ , \new_[32112]_ ,
    \new_[32115]_ , \new_[32118]_ , \new_[32119]_ , \new_[32120]_ ,
    \new_[32124]_ , \new_[32125]_ , \new_[32128]_ , \new_[32131]_ ,
    \new_[32132]_ , \new_[32133]_ , \new_[32137]_ , \new_[32138]_ ,
    \new_[32141]_ , \new_[32144]_ , \new_[32145]_ , \new_[32146]_ ,
    \new_[32150]_ , \new_[32151]_ , \new_[32154]_ , \new_[32157]_ ,
    \new_[32158]_ , \new_[32159]_ , \new_[32163]_ , \new_[32164]_ ,
    \new_[32167]_ , \new_[32170]_ , \new_[32171]_ , \new_[32172]_ ,
    \new_[32176]_ , \new_[32177]_ , \new_[32180]_ , \new_[32183]_ ,
    \new_[32184]_ , \new_[32185]_ , \new_[32189]_ , \new_[32190]_ ,
    \new_[32193]_ , \new_[32196]_ , \new_[32197]_ , \new_[32198]_ ,
    \new_[32202]_ , \new_[32203]_ , \new_[32206]_ , \new_[32209]_ ,
    \new_[32210]_ , \new_[32211]_ , \new_[32215]_ , \new_[32216]_ ,
    \new_[32219]_ , \new_[32222]_ , \new_[32223]_ , \new_[32224]_ ,
    \new_[32228]_ , \new_[32229]_ , \new_[32232]_ , \new_[32235]_ ,
    \new_[32236]_ , \new_[32237]_ , \new_[32241]_ , \new_[32242]_ ,
    \new_[32245]_ , \new_[32248]_ , \new_[32249]_ , \new_[32250]_ ,
    \new_[32254]_ , \new_[32255]_ , \new_[32258]_ , \new_[32261]_ ,
    \new_[32262]_ , \new_[32263]_ , \new_[32267]_ , \new_[32268]_ ,
    \new_[32271]_ , \new_[32274]_ , \new_[32275]_ , \new_[32276]_ ,
    \new_[32280]_ , \new_[32281]_ , \new_[32284]_ , \new_[32287]_ ,
    \new_[32288]_ , \new_[32289]_ , \new_[32293]_ , \new_[32294]_ ,
    \new_[32297]_ , \new_[32300]_ , \new_[32301]_ , \new_[32302]_ ,
    \new_[32306]_ , \new_[32307]_ , \new_[32310]_ , \new_[32313]_ ,
    \new_[32314]_ , \new_[32315]_ , \new_[32319]_ , \new_[32320]_ ,
    \new_[32323]_ , \new_[32326]_ , \new_[32327]_ , \new_[32328]_ ,
    \new_[32332]_ , \new_[32333]_ , \new_[32336]_ , \new_[32339]_ ,
    \new_[32340]_ , \new_[32341]_ , \new_[32345]_ , \new_[32346]_ ,
    \new_[32349]_ , \new_[32352]_ , \new_[32353]_ , \new_[32354]_ ,
    \new_[32358]_ , \new_[32359]_ , \new_[32362]_ , \new_[32365]_ ,
    \new_[32366]_ , \new_[32367]_ , \new_[32371]_ , \new_[32372]_ ,
    \new_[32375]_ , \new_[32378]_ , \new_[32379]_ , \new_[32380]_ ,
    \new_[32384]_ , \new_[32385]_ , \new_[32388]_ , \new_[32391]_ ,
    \new_[32392]_ , \new_[32393]_ , \new_[32397]_ , \new_[32398]_ ,
    \new_[32401]_ , \new_[32404]_ , \new_[32405]_ , \new_[32406]_ ,
    \new_[32410]_ , \new_[32411]_ , \new_[32414]_ , \new_[32417]_ ,
    \new_[32418]_ , \new_[32419]_ , \new_[32423]_ , \new_[32424]_ ,
    \new_[32427]_ , \new_[32430]_ , \new_[32431]_ , \new_[32432]_ ,
    \new_[32436]_ , \new_[32437]_ , \new_[32440]_ , \new_[32443]_ ,
    \new_[32444]_ , \new_[32445]_ , \new_[32449]_ , \new_[32450]_ ,
    \new_[32453]_ , \new_[32456]_ , \new_[32457]_ , \new_[32458]_ ,
    \new_[32462]_ , \new_[32463]_ , \new_[32466]_ , \new_[32469]_ ,
    \new_[32470]_ , \new_[32471]_ , \new_[32475]_ , \new_[32476]_ ,
    \new_[32479]_ , \new_[32482]_ , \new_[32483]_ , \new_[32484]_ ,
    \new_[32488]_ , \new_[32489]_ , \new_[32492]_ , \new_[32495]_ ,
    \new_[32496]_ , \new_[32497]_ , \new_[32501]_ , \new_[32502]_ ,
    \new_[32505]_ , \new_[32508]_ , \new_[32509]_ , \new_[32510]_ ,
    \new_[32514]_ , \new_[32515]_ , \new_[32518]_ , \new_[32521]_ ,
    \new_[32522]_ , \new_[32523]_ , \new_[32527]_ , \new_[32528]_ ,
    \new_[32531]_ , \new_[32534]_ , \new_[32535]_ , \new_[32536]_ ,
    \new_[32540]_ , \new_[32541]_ , \new_[32544]_ , \new_[32547]_ ,
    \new_[32548]_ , \new_[32549]_ , \new_[32553]_ , \new_[32554]_ ,
    \new_[32557]_ , \new_[32560]_ , \new_[32561]_ , \new_[32562]_ ,
    \new_[32566]_ , \new_[32567]_ , \new_[32570]_ , \new_[32573]_ ,
    \new_[32574]_ , \new_[32575]_ , \new_[32579]_ , \new_[32580]_ ,
    \new_[32583]_ , \new_[32586]_ , \new_[32587]_ , \new_[32588]_ ,
    \new_[32592]_ , \new_[32593]_ , \new_[32596]_ , \new_[32599]_ ,
    \new_[32600]_ , \new_[32601]_ , \new_[32605]_ , \new_[32606]_ ,
    \new_[32609]_ , \new_[32612]_ , \new_[32613]_ , \new_[32614]_ ,
    \new_[32618]_ , \new_[32619]_ , \new_[32622]_ , \new_[32625]_ ,
    \new_[32626]_ , \new_[32627]_ , \new_[32631]_ , \new_[32632]_ ,
    \new_[32635]_ , \new_[32638]_ , \new_[32639]_ , \new_[32640]_ ,
    \new_[32644]_ , \new_[32645]_ , \new_[32648]_ , \new_[32651]_ ,
    \new_[32652]_ , \new_[32653]_ , \new_[32657]_ , \new_[32658]_ ,
    \new_[32661]_ , \new_[32664]_ , \new_[32665]_ , \new_[32666]_ ,
    \new_[32670]_ , \new_[32671]_ , \new_[32674]_ , \new_[32677]_ ,
    \new_[32678]_ , \new_[32679]_ , \new_[32683]_ , \new_[32684]_ ,
    \new_[32687]_ , \new_[32690]_ , \new_[32691]_ , \new_[32692]_ ,
    \new_[32696]_ , \new_[32697]_ , \new_[32700]_ , \new_[32703]_ ,
    \new_[32704]_ , \new_[32705]_ , \new_[32709]_ , \new_[32710]_ ,
    \new_[32713]_ , \new_[32716]_ , \new_[32717]_ , \new_[32718]_ ,
    \new_[32722]_ , \new_[32723]_ , \new_[32726]_ , \new_[32729]_ ,
    \new_[32730]_ , \new_[32731]_ , \new_[32735]_ , \new_[32736]_ ,
    \new_[32739]_ , \new_[32742]_ , \new_[32743]_ , \new_[32744]_ ,
    \new_[32748]_ , \new_[32749]_ , \new_[32752]_ , \new_[32755]_ ,
    \new_[32756]_ , \new_[32757]_ , \new_[32761]_ , \new_[32762]_ ,
    \new_[32765]_ , \new_[32768]_ , \new_[32769]_ , \new_[32770]_ ,
    \new_[32774]_ , \new_[32775]_ , \new_[32778]_ , \new_[32781]_ ,
    \new_[32782]_ , \new_[32783]_ , \new_[32787]_ , \new_[32788]_ ,
    \new_[32791]_ , \new_[32794]_ , \new_[32795]_ , \new_[32796]_ ,
    \new_[32800]_ , \new_[32801]_ , \new_[32804]_ , \new_[32807]_ ,
    \new_[32808]_ , \new_[32809]_ , \new_[32813]_ , \new_[32814]_ ,
    \new_[32817]_ , \new_[32820]_ , \new_[32821]_ , \new_[32822]_ ,
    \new_[32826]_ , \new_[32827]_ , \new_[32830]_ , \new_[32833]_ ,
    \new_[32834]_ , \new_[32835]_ , \new_[32839]_ , \new_[32840]_ ,
    \new_[32843]_ , \new_[32846]_ , \new_[32847]_ , \new_[32848]_ ,
    \new_[32852]_ , \new_[32853]_ , \new_[32856]_ , \new_[32859]_ ,
    \new_[32860]_ , \new_[32861]_ , \new_[32865]_ , \new_[32866]_ ,
    \new_[32869]_ , \new_[32872]_ , \new_[32873]_ , \new_[32874]_ ,
    \new_[32878]_ , \new_[32879]_ , \new_[32882]_ , \new_[32885]_ ,
    \new_[32886]_ , \new_[32887]_ , \new_[32891]_ , \new_[32892]_ ,
    \new_[32895]_ , \new_[32898]_ , \new_[32899]_ , \new_[32900]_ ,
    \new_[32904]_ , \new_[32905]_ , \new_[32908]_ , \new_[32911]_ ,
    \new_[32912]_ , \new_[32913]_ , \new_[32917]_ , \new_[32918]_ ,
    \new_[32921]_ , \new_[32924]_ , \new_[32925]_ , \new_[32926]_ ,
    \new_[32930]_ , \new_[32931]_ , \new_[32934]_ , \new_[32937]_ ,
    \new_[32938]_ , \new_[32939]_ , \new_[32943]_ , \new_[32944]_ ,
    \new_[32947]_ , \new_[32950]_ , \new_[32951]_ , \new_[32952]_ ,
    \new_[32956]_ , \new_[32957]_ , \new_[32960]_ , \new_[32963]_ ,
    \new_[32964]_ , \new_[32965]_ , \new_[32969]_ , \new_[32970]_ ,
    \new_[32973]_ , \new_[32976]_ , \new_[32977]_ , \new_[32978]_ ,
    \new_[32982]_ , \new_[32983]_ , \new_[32986]_ , \new_[32989]_ ,
    \new_[32990]_ , \new_[32991]_ , \new_[32995]_ , \new_[32996]_ ,
    \new_[32999]_ , \new_[33002]_ , \new_[33003]_ , \new_[33004]_ ,
    \new_[33008]_ , \new_[33009]_ , \new_[33012]_ , \new_[33015]_ ,
    \new_[33016]_ , \new_[33017]_ , \new_[33021]_ , \new_[33022]_ ,
    \new_[33025]_ , \new_[33028]_ , \new_[33029]_ , \new_[33030]_ ,
    \new_[33034]_ , \new_[33035]_ , \new_[33038]_ , \new_[33041]_ ,
    \new_[33042]_ , \new_[33043]_ , \new_[33047]_ , \new_[33048]_ ,
    \new_[33051]_ , \new_[33054]_ , \new_[33055]_ , \new_[33056]_ ,
    \new_[33060]_ , \new_[33061]_ , \new_[33064]_ , \new_[33067]_ ,
    \new_[33068]_ , \new_[33069]_ , \new_[33073]_ , \new_[33074]_ ,
    \new_[33077]_ , \new_[33080]_ , \new_[33081]_ , \new_[33082]_ ,
    \new_[33086]_ , \new_[33087]_ , \new_[33090]_ , \new_[33093]_ ,
    \new_[33094]_ , \new_[33095]_ , \new_[33099]_ , \new_[33100]_ ,
    \new_[33103]_ , \new_[33106]_ , \new_[33107]_ , \new_[33108]_ ,
    \new_[33112]_ , \new_[33113]_ , \new_[33116]_ , \new_[33119]_ ,
    \new_[33120]_ , \new_[33121]_ , \new_[33125]_ , \new_[33126]_ ,
    \new_[33129]_ , \new_[33132]_ , \new_[33133]_ , \new_[33134]_ ,
    \new_[33138]_ , \new_[33139]_ , \new_[33142]_ , \new_[33145]_ ,
    \new_[33146]_ , \new_[33147]_ , \new_[33151]_ , \new_[33152]_ ,
    \new_[33155]_ , \new_[33158]_ , \new_[33159]_ , \new_[33160]_ ,
    \new_[33164]_ , \new_[33165]_ , \new_[33168]_ , \new_[33171]_ ,
    \new_[33172]_ , \new_[33173]_ , \new_[33177]_ , \new_[33178]_ ,
    \new_[33181]_ , \new_[33184]_ , \new_[33185]_ , \new_[33186]_ ,
    \new_[33190]_ , \new_[33191]_ , \new_[33194]_ , \new_[33197]_ ,
    \new_[33198]_ , \new_[33199]_ , \new_[33203]_ , \new_[33204]_ ,
    \new_[33207]_ , \new_[33210]_ , \new_[33211]_ , \new_[33212]_ ,
    \new_[33216]_ , \new_[33217]_ , \new_[33220]_ , \new_[33223]_ ,
    \new_[33224]_ , \new_[33225]_ , \new_[33229]_ , \new_[33230]_ ,
    \new_[33233]_ , \new_[33236]_ , \new_[33237]_ , \new_[33238]_ ,
    \new_[33242]_ , \new_[33243]_ , \new_[33246]_ , \new_[33249]_ ,
    \new_[33250]_ , \new_[33251]_ , \new_[33255]_ , \new_[33256]_ ,
    \new_[33259]_ , \new_[33262]_ , \new_[33263]_ , \new_[33264]_ ,
    \new_[33268]_ , \new_[33269]_ , \new_[33272]_ , \new_[33275]_ ,
    \new_[33276]_ , \new_[33277]_ , \new_[33281]_ , \new_[33282]_ ,
    \new_[33285]_ , \new_[33288]_ , \new_[33289]_ , \new_[33290]_ ,
    \new_[33294]_ , \new_[33295]_ , \new_[33298]_ , \new_[33301]_ ,
    \new_[33302]_ , \new_[33303]_ , \new_[33307]_ , \new_[33308]_ ,
    \new_[33311]_ , \new_[33314]_ , \new_[33315]_ , \new_[33316]_ ,
    \new_[33320]_ , \new_[33321]_ , \new_[33324]_ , \new_[33327]_ ,
    \new_[33328]_ , \new_[33329]_ , \new_[33333]_ , \new_[33334]_ ,
    \new_[33337]_ , \new_[33340]_ , \new_[33341]_ , \new_[33342]_ ,
    \new_[33346]_ , \new_[33347]_ , \new_[33350]_ , \new_[33353]_ ,
    \new_[33354]_ , \new_[33355]_ , \new_[33359]_ , \new_[33360]_ ,
    \new_[33363]_ , \new_[33366]_ , \new_[33367]_ , \new_[33368]_ ,
    \new_[33372]_ , \new_[33373]_ , \new_[33376]_ , \new_[33379]_ ,
    \new_[33380]_ , \new_[33381]_ , \new_[33385]_ , \new_[33386]_ ,
    \new_[33389]_ , \new_[33392]_ , \new_[33393]_ , \new_[33394]_ ,
    \new_[33398]_ , \new_[33399]_ , \new_[33402]_ , \new_[33405]_ ,
    \new_[33406]_ , \new_[33407]_ , \new_[33411]_ , \new_[33412]_ ,
    \new_[33415]_ , \new_[33418]_ , \new_[33419]_ , \new_[33420]_ ,
    \new_[33424]_ , \new_[33425]_ , \new_[33428]_ , \new_[33431]_ ,
    \new_[33432]_ , \new_[33433]_ , \new_[33437]_ , \new_[33438]_ ,
    \new_[33441]_ , \new_[33444]_ , \new_[33445]_ , \new_[33446]_ ,
    \new_[33450]_ , \new_[33451]_ , \new_[33454]_ , \new_[33457]_ ,
    \new_[33458]_ , \new_[33459]_ , \new_[33463]_ , \new_[33464]_ ,
    \new_[33467]_ , \new_[33470]_ , \new_[33471]_ , \new_[33472]_ ,
    \new_[33476]_ , \new_[33477]_ , \new_[33480]_ , \new_[33483]_ ,
    \new_[33484]_ , \new_[33485]_ , \new_[33489]_ , \new_[33490]_ ,
    \new_[33493]_ , \new_[33496]_ , \new_[33497]_ , \new_[33498]_ ,
    \new_[33502]_ , \new_[33503]_ , \new_[33506]_ , \new_[33509]_ ,
    \new_[33510]_ , \new_[33511]_ , \new_[33515]_ , \new_[33516]_ ,
    \new_[33519]_ , \new_[33522]_ , \new_[33523]_ , \new_[33524]_ ,
    \new_[33528]_ , \new_[33529]_ , \new_[33532]_ , \new_[33535]_ ,
    \new_[33536]_ , \new_[33537]_ , \new_[33541]_ , \new_[33542]_ ,
    \new_[33545]_ , \new_[33548]_ , \new_[33549]_ , \new_[33550]_ ,
    \new_[33554]_ , \new_[33555]_ , \new_[33558]_ , \new_[33561]_ ,
    \new_[33562]_ , \new_[33563]_ , \new_[33567]_ , \new_[33568]_ ,
    \new_[33571]_ , \new_[33574]_ , \new_[33575]_ , \new_[33576]_ ,
    \new_[33580]_ , \new_[33581]_ , \new_[33584]_ , \new_[33587]_ ,
    \new_[33588]_ , \new_[33589]_ , \new_[33593]_ , \new_[33594]_ ,
    \new_[33597]_ , \new_[33600]_ , \new_[33601]_ , \new_[33602]_ ,
    \new_[33606]_ , \new_[33607]_ , \new_[33610]_ , \new_[33613]_ ,
    \new_[33614]_ , \new_[33615]_ , \new_[33619]_ , \new_[33620]_ ,
    \new_[33623]_ , \new_[33626]_ , \new_[33627]_ , \new_[33628]_ ,
    \new_[33632]_ , \new_[33633]_ , \new_[33636]_ , \new_[33639]_ ,
    \new_[33640]_ , \new_[33641]_ , \new_[33645]_ , \new_[33646]_ ,
    \new_[33649]_ , \new_[33652]_ , \new_[33653]_ , \new_[33654]_ ,
    \new_[33658]_ , \new_[33659]_ , \new_[33662]_ , \new_[33665]_ ,
    \new_[33666]_ , \new_[33667]_ , \new_[33671]_ , \new_[33672]_ ,
    \new_[33675]_ , \new_[33678]_ , \new_[33679]_ , \new_[33680]_ ,
    \new_[33684]_ , \new_[33685]_ , \new_[33688]_ , \new_[33691]_ ,
    \new_[33692]_ , \new_[33693]_ , \new_[33697]_ , \new_[33698]_ ,
    \new_[33701]_ , \new_[33704]_ , \new_[33705]_ , \new_[33706]_ ,
    \new_[33710]_ , \new_[33711]_ , \new_[33714]_ , \new_[33717]_ ,
    \new_[33718]_ , \new_[33719]_ , \new_[33723]_ , \new_[33724]_ ,
    \new_[33727]_ , \new_[33730]_ , \new_[33731]_ , \new_[33732]_ ,
    \new_[33736]_ , \new_[33737]_ , \new_[33740]_ , \new_[33743]_ ,
    \new_[33744]_ , \new_[33745]_ , \new_[33749]_ , \new_[33750]_ ,
    \new_[33753]_ , \new_[33756]_ , \new_[33757]_ , \new_[33758]_ ,
    \new_[33762]_ , \new_[33763]_ , \new_[33766]_ , \new_[33769]_ ,
    \new_[33770]_ , \new_[33771]_ , \new_[33775]_ , \new_[33776]_ ,
    \new_[33779]_ , \new_[33782]_ , \new_[33783]_ , \new_[33784]_ ,
    \new_[33788]_ , \new_[33789]_ , \new_[33792]_ , \new_[33795]_ ,
    \new_[33796]_ , \new_[33797]_ , \new_[33801]_ , \new_[33802]_ ,
    \new_[33805]_ , \new_[33808]_ , \new_[33809]_ , \new_[33810]_ ,
    \new_[33814]_ , \new_[33815]_ , \new_[33818]_ , \new_[33821]_ ,
    \new_[33822]_ , \new_[33823]_ , \new_[33827]_ , \new_[33828]_ ,
    \new_[33831]_ , \new_[33834]_ , \new_[33835]_ , \new_[33836]_ ,
    \new_[33840]_ , \new_[33841]_ , \new_[33844]_ , \new_[33847]_ ,
    \new_[33848]_ , \new_[33849]_ , \new_[33853]_ , \new_[33854]_ ,
    \new_[33857]_ , \new_[33860]_ , \new_[33861]_ , \new_[33862]_ ,
    \new_[33866]_ , \new_[33867]_ , \new_[33870]_ , \new_[33873]_ ,
    \new_[33874]_ , \new_[33875]_ , \new_[33879]_ , \new_[33880]_ ,
    \new_[33883]_ , \new_[33886]_ , \new_[33887]_ , \new_[33888]_ ,
    \new_[33892]_ , \new_[33893]_ , \new_[33896]_ , \new_[33899]_ ,
    \new_[33900]_ , \new_[33901]_ , \new_[33905]_ , \new_[33906]_ ,
    \new_[33909]_ , \new_[33912]_ , \new_[33913]_ , \new_[33914]_ ,
    \new_[33918]_ , \new_[33919]_ , \new_[33922]_ , \new_[33925]_ ,
    \new_[33926]_ , \new_[33927]_ , \new_[33931]_ , \new_[33932]_ ,
    \new_[33935]_ , \new_[33938]_ , \new_[33939]_ , \new_[33940]_ ,
    \new_[33944]_ , \new_[33945]_ , \new_[33948]_ , \new_[33951]_ ,
    \new_[33952]_ , \new_[33953]_ , \new_[33957]_ , \new_[33958]_ ,
    \new_[33961]_ , \new_[33964]_ , \new_[33965]_ , \new_[33966]_ ,
    \new_[33970]_ , \new_[33971]_ , \new_[33974]_ , \new_[33977]_ ,
    \new_[33978]_ , \new_[33979]_ , \new_[33983]_ , \new_[33984]_ ,
    \new_[33987]_ , \new_[33990]_ , \new_[33991]_ , \new_[33992]_ ,
    \new_[33996]_ , \new_[33997]_ , \new_[34000]_ , \new_[34003]_ ,
    \new_[34004]_ , \new_[34005]_ , \new_[34009]_ , \new_[34010]_ ,
    \new_[34013]_ , \new_[34016]_ , \new_[34017]_ , \new_[34018]_ ,
    \new_[34022]_ , \new_[34023]_ , \new_[34026]_ , \new_[34029]_ ,
    \new_[34030]_ , \new_[34031]_ , \new_[34035]_ , \new_[34036]_ ,
    \new_[34039]_ , \new_[34042]_ , \new_[34043]_ , \new_[34044]_ ,
    \new_[34048]_ , \new_[34049]_ , \new_[34052]_ , \new_[34055]_ ,
    \new_[34056]_ , \new_[34057]_ , \new_[34061]_ , \new_[34062]_ ,
    \new_[34065]_ , \new_[34068]_ , \new_[34069]_ , \new_[34070]_ ,
    \new_[34074]_ , \new_[34075]_ , \new_[34078]_ , \new_[34081]_ ,
    \new_[34082]_ , \new_[34083]_ , \new_[34087]_ , \new_[34088]_ ,
    \new_[34091]_ , \new_[34094]_ , \new_[34095]_ , \new_[34096]_ ,
    \new_[34100]_ , \new_[34101]_ , \new_[34104]_ , \new_[34107]_ ,
    \new_[34108]_ , \new_[34109]_ , \new_[34113]_ , \new_[34114]_ ,
    \new_[34117]_ , \new_[34120]_ , \new_[34121]_ , \new_[34122]_ ,
    \new_[34126]_ , \new_[34127]_ , \new_[34130]_ , \new_[34133]_ ,
    \new_[34134]_ , \new_[34135]_ , \new_[34139]_ , \new_[34140]_ ,
    \new_[34143]_ , \new_[34146]_ , \new_[34147]_ , \new_[34148]_ ,
    \new_[34152]_ , \new_[34153]_ , \new_[34156]_ , \new_[34159]_ ,
    \new_[34160]_ , \new_[34161]_ , \new_[34165]_ , \new_[34166]_ ,
    \new_[34169]_ , \new_[34172]_ , \new_[34173]_ , \new_[34174]_ ,
    \new_[34178]_ , \new_[34179]_ , \new_[34182]_ , \new_[34185]_ ,
    \new_[34186]_ , \new_[34187]_ , \new_[34191]_ , \new_[34192]_ ,
    \new_[34195]_ , \new_[34198]_ , \new_[34199]_ , \new_[34200]_ ,
    \new_[34204]_ , \new_[34205]_ , \new_[34208]_ , \new_[34211]_ ,
    \new_[34212]_ , \new_[34213]_ , \new_[34217]_ , \new_[34218]_ ,
    \new_[34221]_ , \new_[34224]_ , \new_[34225]_ , \new_[34226]_ ,
    \new_[34230]_ , \new_[34231]_ , \new_[34234]_ , \new_[34237]_ ,
    \new_[34238]_ , \new_[34239]_ , \new_[34243]_ , \new_[34244]_ ,
    \new_[34247]_ , \new_[34250]_ , \new_[34251]_ , \new_[34252]_ ,
    \new_[34256]_ , \new_[34257]_ , \new_[34260]_ , \new_[34263]_ ,
    \new_[34264]_ , \new_[34265]_ , \new_[34269]_ , \new_[34270]_ ,
    \new_[34273]_ , \new_[34276]_ , \new_[34277]_ , \new_[34278]_ ,
    \new_[34282]_ , \new_[34283]_ , \new_[34286]_ , \new_[34289]_ ,
    \new_[34290]_ , \new_[34291]_ , \new_[34295]_ , \new_[34296]_ ,
    \new_[34299]_ , \new_[34302]_ , \new_[34303]_ , \new_[34304]_ ,
    \new_[34308]_ , \new_[34309]_ , \new_[34312]_ , \new_[34315]_ ,
    \new_[34316]_ , \new_[34317]_ , \new_[34321]_ , \new_[34322]_ ,
    \new_[34325]_ , \new_[34328]_ , \new_[34329]_ , \new_[34330]_ ,
    \new_[34334]_ , \new_[34335]_ , \new_[34338]_ , \new_[34341]_ ,
    \new_[34342]_ , \new_[34343]_ , \new_[34347]_ , \new_[34348]_ ,
    \new_[34351]_ , \new_[34354]_ , \new_[34355]_ , \new_[34356]_ ,
    \new_[34360]_ , \new_[34361]_ , \new_[34364]_ , \new_[34367]_ ,
    \new_[34368]_ , \new_[34369]_ , \new_[34373]_ , \new_[34374]_ ,
    \new_[34377]_ , \new_[34380]_ , \new_[34381]_ , \new_[34382]_ ,
    \new_[34386]_ , \new_[34387]_ , \new_[34390]_ , \new_[34393]_ ,
    \new_[34394]_ , \new_[34395]_ , \new_[34399]_ , \new_[34400]_ ,
    \new_[34403]_ , \new_[34406]_ , \new_[34407]_ , \new_[34408]_ ,
    \new_[34412]_ , \new_[34413]_ , \new_[34416]_ , \new_[34419]_ ,
    \new_[34420]_ , \new_[34421]_ , \new_[34425]_ , \new_[34426]_ ,
    \new_[34429]_ , \new_[34432]_ , \new_[34433]_ , \new_[34434]_ ,
    \new_[34438]_ , \new_[34439]_ , \new_[34442]_ , \new_[34445]_ ,
    \new_[34446]_ , \new_[34447]_ , \new_[34450]_ , \new_[34453]_ ,
    \new_[34454]_ , \new_[34457]_ , \new_[34460]_ , \new_[34461]_ ,
    \new_[34462]_ , \new_[34466]_ , \new_[34467]_ , \new_[34470]_ ,
    \new_[34473]_ , \new_[34474]_ , \new_[34475]_ , \new_[34478]_ ,
    \new_[34481]_ , \new_[34482]_ , \new_[34485]_ , \new_[34488]_ ,
    \new_[34489]_ , \new_[34490]_ , \new_[34494]_ , \new_[34495]_ ,
    \new_[34498]_ , \new_[34501]_ , \new_[34502]_ , \new_[34503]_ ,
    \new_[34506]_ , \new_[34509]_ , \new_[34510]_ , \new_[34513]_ ,
    \new_[34516]_ , \new_[34517]_ , \new_[34518]_ , \new_[34522]_ ,
    \new_[34523]_ , \new_[34526]_ , \new_[34529]_ , \new_[34530]_ ,
    \new_[34531]_ , \new_[34534]_ , \new_[34537]_ , \new_[34538]_ ,
    \new_[34541]_ , \new_[34544]_ , \new_[34545]_ , \new_[34546]_ ,
    \new_[34550]_ , \new_[34551]_ , \new_[34554]_ , \new_[34557]_ ,
    \new_[34558]_ , \new_[34559]_ , \new_[34562]_ , \new_[34565]_ ,
    \new_[34566]_ , \new_[34569]_ , \new_[34572]_ , \new_[34573]_ ,
    \new_[34574]_ , \new_[34578]_ , \new_[34579]_ , \new_[34582]_ ,
    \new_[34585]_ , \new_[34586]_ , \new_[34587]_ , \new_[34590]_ ,
    \new_[34593]_ , \new_[34594]_ , \new_[34597]_ , \new_[34600]_ ,
    \new_[34601]_ , \new_[34602]_ , \new_[34606]_ , \new_[34607]_ ,
    \new_[34610]_ , \new_[34613]_ , \new_[34614]_ , \new_[34615]_ ,
    \new_[34618]_ , \new_[34621]_ , \new_[34622]_ , \new_[34625]_ ,
    \new_[34628]_ , \new_[34629]_ , \new_[34630]_ , \new_[34634]_ ,
    \new_[34635]_ , \new_[34638]_ , \new_[34641]_ , \new_[34642]_ ,
    \new_[34643]_ , \new_[34646]_ , \new_[34649]_ , \new_[34650]_ ,
    \new_[34653]_ , \new_[34656]_ , \new_[34657]_ , \new_[34658]_ ,
    \new_[34662]_ , \new_[34663]_ , \new_[34666]_ , \new_[34669]_ ,
    \new_[34670]_ , \new_[34671]_ , \new_[34674]_ , \new_[34677]_ ,
    \new_[34678]_ , \new_[34681]_ , \new_[34684]_ , \new_[34685]_ ,
    \new_[34686]_ , \new_[34690]_ , \new_[34691]_ , \new_[34694]_ ,
    \new_[34697]_ , \new_[34698]_ , \new_[34699]_ , \new_[34702]_ ,
    \new_[34705]_ , \new_[34706]_ , \new_[34709]_ , \new_[34712]_ ,
    \new_[34713]_ , \new_[34714]_ , \new_[34718]_ , \new_[34719]_ ,
    \new_[34722]_ , \new_[34725]_ , \new_[34726]_ , \new_[34727]_ ,
    \new_[34730]_ , \new_[34733]_ , \new_[34734]_ , \new_[34737]_ ,
    \new_[34740]_ , \new_[34741]_ , \new_[34742]_ , \new_[34746]_ ,
    \new_[34747]_ , \new_[34750]_ , \new_[34753]_ , \new_[34754]_ ,
    \new_[34755]_ , \new_[34758]_ , \new_[34761]_ , \new_[34762]_ ,
    \new_[34765]_ , \new_[34768]_ , \new_[34769]_ , \new_[34770]_ ,
    \new_[34774]_ , \new_[34775]_ , \new_[34778]_ , \new_[34781]_ ,
    \new_[34782]_ , \new_[34783]_ , \new_[34786]_ , \new_[34789]_ ,
    \new_[34790]_ , \new_[34793]_ , \new_[34796]_ , \new_[34797]_ ,
    \new_[34798]_ , \new_[34802]_ , \new_[34803]_ , \new_[34806]_ ,
    \new_[34809]_ , \new_[34810]_ , \new_[34811]_ , \new_[34814]_ ,
    \new_[34817]_ , \new_[34818]_ , \new_[34821]_ , \new_[34824]_ ,
    \new_[34825]_ , \new_[34826]_ , \new_[34830]_ , \new_[34831]_ ,
    \new_[34834]_ , \new_[34837]_ , \new_[34838]_ , \new_[34839]_ ,
    \new_[34842]_ , \new_[34845]_ , \new_[34846]_ , \new_[34849]_ ,
    \new_[34852]_ , \new_[34853]_ , \new_[34854]_ , \new_[34858]_ ,
    \new_[34859]_ , \new_[34862]_ , \new_[34865]_ , \new_[34866]_ ,
    \new_[34867]_ , \new_[34870]_ , \new_[34873]_ , \new_[34874]_ ,
    \new_[34877]_ , \new_[34880]_ , \new_[34881]_ , \new_[34882]_ ,
    \new_[34886]_ , \new_[34887]_ , \new_[34890]_ , \new_[34893]_ ,
    \new_[34894]_ , \new_[34895]_ , \new_[34898]_ , \new_[34901]_ ,
    \new_[34902]_ , \new_[34905]_ , \new_[34908]_ , \new_[34909]_ ,
    \new_[34910]_ , \new_[34914]_ , \new_[34915]_ , \new_[34918]_ ,
    \new_[34921]_ , \new_[34922]_ , \new_[34923]_ , \new_[34926]_ ,
    \new_[34929]_ , \new_[34930]_ , \new_[34933]_ , \new_[34936]_ ,
    \new_[34937]_ , \new_[34938]_ , \new_[34942]_ , \new_[34943]_ ,
    \new_[34946]_ , \new_[34949]_ , \new_[34950]_ , \new_[34951]_ ,
    \new_[34954]_ , \new_[34957]_ , \new_[34958]_ , \new_[34961]_ ,
    \new_[34964]_ , \new_[34965]_ , \new_[34966]_ , \new_[34970]_ ,
    \new_[34971]_ , \new_[34974]_ , \new_[34977]_ , \new_[34978]_ ,
    \new_[34979]_ , \new_[34982]_ , \new_[34985]_ , \new_[34986]_ ,
    \new_[34989]_ , \new_[34992]_ , \new_[34993]_ , \new_[34994]_ ,
    \new_[34998]_ , \new_[34999]_ , \new_[35002]_ , \new_[35005]_ ,
    \new_[35006]_ , \new_[35007]_ , \new_[35010]_ , \new_[35013]_ ,
    \new_[35014]_ , \new_[35017]_ , \new_[35020]_ , \new_[35021]_ ,
    \new_[35022]_ , \new_[35026]_ , \new_[35027]_ , \new_[35030]_ ,
    \new_[35033]_ , \new_[35034]_ , \new_[35035]_ , \new_[35038]_ ,
    \new_[35041]_ , \new_[35042]_ , \new_[35045]_ , \new_[35048]_ ,
    \new_[35049]_ , \new_[35050]_ , \new_[35054]_ , \new_[35055]_ ,
    \new_[35058]_ , \new_[35061]_ , \new_[35062]_ , \new_[35063]_ ,
    \new_[35066]_ , \new_[35069]_ , \new_[35070]_ , \new_[35073]_ ,
    \new_[35076]_ , \new_[35077]_ , \new_[35078]_ , \new_[35082]_ ,
    \new_[35083]_ , \new_[35086]_ , \new_[35089]_ , \new_[35090]_ ,
    \new_[35091]_ , \new_[35094]_ , \new_[35097]_ , \new_[35098]_ ,
    \new_[35101]_ , \new_[35104]_ , \new_[35105]_ , \new_[35106]_ ,
    \new_[35110]_ , \new_[35111]_ , \new_[35114]_ , \new_[35117]_ ,
    \new_[35118]_ , \new_[35119]_ , \new_[35122]_ , \new_[35125]_ ,
    \new_[35126]_ , \new_[35129]_ , \new_[35132]_ , \new_[35133]_ ,
    \new_[35134]_ , \new_[35138]_ , \new_[35139]_ , \new_[35142]_ ,
    \new_[35145]_ , \new_[35146]_ , \new_[35147]_ , \new_[35150]_ ,
    \new_[35153]_ , \new_[35154]_ , \new_[35157]_ , \new_[35160]_ ,
    \new_[35161]_ , \new_[35162]_ , \new_[35166]_ , \new_[35167]_ ,
    \new_[35170]_ , \new_[35173]_ , \new_[35174]_ , \new_[35175]_ ,
    \new_[35178]_ , \new_[35181]_ , \new_[35182]_ , \new_[35185]_ ,
    \new_[35188]_ , \new_[35189]_ , \new_[35190]_ , \new_[35194]_ ,
    \new_[35195]_ , \new_[35198]_ , \new_[35201]_ , \new_[35202]_ ,
    \new_[35203]_ , \new_[35206]_ , \new_[35209]_ , \new_[35210]_ ,
    \new_[35213]_ , \new_[35216]_ , \new_[35217]_ , \new_[35218]_ ,
    \new_[35222]_ , \new_[35223]_ , \new_[35226]_ , \new_[35229]_ ,
    \new_[35230]_ , \new_[35231]_ , \new_[35234]_ , \new_[35237]_ ,
    \new_[35238]_ , \new_[35241]_ , \new_[35244]_ , \new_[35245]_ ,
    \new_[35246]_ , \new_[35250]_ , \new_[35251]_ , \new_[35254]_ ,
    \new_[35257]_ , \new_[35258]_ , \new_[35259]_ , \new_[35262]_ ,
    \new_[35265]_ , \new_[35266]_ , \new_[35269]_ , \new_[35272]_ ,
    \new_[35273]_ , \new_[35274]_ , \new_[35278]_ , \new_[35279]_ ,
    \new_[35282]_ , \new_[35285]_ , \new_[35286]_ , \new_[35287]_ ,
    \new_[35290]_ , \new_[35293]_ , \new_[35294]_ , \new_[35297]_ ,
    \new_[35300]_ , \new_[35301]_ , \new_[35302]_ , \new_[35306]_ ,
    \new_[35307]_ , \new_[35310]_ , \new_[35313]_ , \new_[35314]_ ,
    \new_[35315]_ , \new_[35318]_ , \new_[35321]_ , \new_[35322]_ ,
    \new_[35325]_ , \new_[35328]_ , \new_[35329]_ , \new_[35330]_ ,
    \new_[35334]_ , \new_[35335]_ , \new_[35338]_ , \new_[35341]_ ,
    \new_[35342]_ , \new_[35343]_ , \new_[35346]_ , \new_[35349]_ ,
    \new_[35350]_ , \new_[35353]_ , \new_[35356]_ , \new_[35357]_ ,
    \new_[35358]_ , \new_[35362]_ , \new_[35363]_ , \new_[35366]_ ,
    \new_[35369]_ , \new_[35370]_ , \new_[35371]_ , \new_[35374]_ ,
    \new_[35377]_ , \new_[35378]_ , \new_[35381]_ , \new_[35384]_ ,
    \new_[35385]_ , \new_[35386]_ , \new_[35390]_ , \new_[35391]_ ,
    \new_[35394]_ , \new_[35397]_ , \new_[35398]_ , \new_[35399]_ ,
    \new_[35402]_ , \new_[35405]_ , \new_[35406]_ , \new_[35409]_ ,
    \new_[35412]_ , \new_[35413]_ , \new_[35414]_ , \new_[35418]_ ,
    \new_[35419]_ , \new_[35422]_ , \new_[35425]_ , \new_[35426]_ ,
    \new_[35427]_ , \new_[35430]_ , \new_[35433]_ , \new_[35434]_ ,
    \new_[35437]_ , \new_[35440]_ , \new_[35441]_ , \new_[35442]_ ,
    \new_[35446]_ , \new_[35447]_ , \new_[35450]_ , \new_[35453]_ ,
    \new_[35454]_ , \new_[35455]_ , \new_[35458]_ , \new_[35461]_ ,
    \new_[35462]_ , \new_[35465]_ , \new_[35468]_ , \new_[35469]_ ,
    \new_[35470]_ , \new_[35474]_ , \new_[35475]_ , \new_[35478]_ ,
    \new_[35481]_ , \new_[35482]_ , \new_[35483]_ , \new_[35486]_ ,
    \new_[35489]_ , \new_[35490]_ , \new_[35493]_ , \new_[35496]_ ,
    \new_[35497]_ , \new_[35498]_ , \new_[35502]_ , \new_[35503]_ ,
    \new_[35506]_ , \new_[35509]_ , \new_[35510]_ , \new_[35511]_ ,
    \new_[35514]_ , \new_[35517]_ , \new_[35518]_ , \new_[35521]_ ,
    \new_[35524]_ , \new_[35525]_ , \new_[35526]_ , \new_[35530]_ ,
    \new_[35531]_ , \new_[35534]_ , \new_[35537]_ , \new_[35538]_ ,
    \new_[35539]_ , \new_[35542]_ , \new_[35545]_ , \new_[35546]_ ,
    \new_[35549]_ , \new_[35552]_ , \new_[35553]_ , \new_[35554]_ ,
    \new_[35558]_ , \new_[35559]_ , \new_[35562]_ , \new_[35565]_ ,
    \new_[35566]_ , \new_[35567]_ , \new_[35570]_ , \new_[35573]_ ,
    \new_[35574]_ , \new_[35577]_ , \new_[35580]_ , \new_[35581]_ ,
    \new_[35582]_ , \new_[35586]_ , \new_[35587]_ , \new_[35590]_ ,
    \new_[35593]_ , \new_[35594]_ , \new_[35595]_ , \new_[35598]_ ,
    \new_[35601]_ , \new_[35602]_ , \new_[35605]_ , \new_[35608]_ ,
    \new_[35609]_ , \new_[35610]_ , \new_[35614]_ , \new_[35615]_ ,
    \new_[35618]_ , \new_[35621]_ , \new_[35622]_ , \new_[35623]_ ,
    \new_[35626]_ , \new_[35629]_ , \new_[35630]_ , \new_[35633]_ ,
    \new_[35636]_ , \new_[35637]_ , \new_[35638]_ , \new_[35642]_ ,
    \new_[35643]_ , \new_[35646]_ , \new_[35649]_ , \new_[35650]_ ,
    \new_[35651]_ , \new_[35654]_ , \new_[35657]_ , \new_[35658]_ ,
    \new_[35661]_ , \new_[35664]_ , \new_[35665]_ , \new_[35666]_ ,
    \new_[35670]_ , \new_[35671]_ , \new_[35674]_ , \new_[35677]_ ,
    \new_[35678]_ , \new_[35679]_ , \new_[35682]_ , \new_[35685]_ ,
    \new_[35686]_ , \new_[35689]_ , \new_[35692]_ , \new_[35693]_ ,
    \new_[35694]_ , \new_[35698]_ , \new_[35699]_ , \new_[35702]_ ,
    \new_[35705]_ , \new_[35706]_ , \new_[35707]_ , \new_[35710]_ ,
    \new_[35713]_ , \new_[35714]_ , \new_[35717]_ , \new_[35720]_ ,
    \new_[35721]_ , \new_[35722]_ , \new_[35726]_ , \new_[35727]_ ,
    \new_[35730]_ , \new_[35733]_ , \new_[35734]_ , \new_[35735]_ ,
    \new_[35738]_ , \new_[35741]_ , \new_[35742]_ , \new_[35745]_ ,
    \new_[35748]_ , \new_[35749]_ , \new_[35750]_ , \new_[35754]_ ,
    \new_[35755]_ , \new_[35758]_ , \new_[35761]_ , \new_[35762]_ ,
    \new_[35763]_ , \new_[35766]_ , \new_[35769]_ , \new_[35770]_ ,
    \new_[35773]_ , \new_[35776]_ , \new_[35777]_ , \new_[35778]_ ,
    \new_[35782]_ , \new_[35783]_ , \new_[35786]_ , \new_[35789]_ ,
    \new_[35790]_ , \new_[35791]_ , \new_[35794]_ , \new_[35797]_ ,
    \new_[35798]_ , \new_[35801]_ , \new_[35804]_ , \new_[35805]_ ,
    \new_[35806]_ , \new_[35810]_ , \new_[35811]_ , \new_[35814]_ ,
    \new_[35817]_ , \new_[35818]_ , \new_[35819]_ , \new_[35822]_ ,
    \new_[35825]_ , \new_[35826]_ , \new_[35829]_ , \new_[35832]_ ,
    \new_[35833]_ , \new_[35834]_ , \new_[35838]_ , \new_[35839]_ ,
    \new_[35842]_ , \new_[35845]_ , \new_[35846]_ , \new_[35847]_ ,
    \new_[35850]_ , \new_[35853]_ , \new_[35854]_ , \new_[35857]_ ,
    \new_[35860]_ , \new_[35861]_ , \new_[35862]_ , \new_[35866]_ ,
    \new_[35867]_ , \new_[35870]_ , \new_[35873]_ , \new_[35874]_ ,
    \new_[35875]_ , \new_[35878]_ , \new_[35881]_ , \new_[35882]_ ,
    \new_[35885]_ , \new_[35888]_ , \new_[35889]_ , \new_[35890]_ ,
    \new_[35894]_ , \new_[35895]_ , \new_[35898]_ , \new_[35901]_ ,
    \new_[35902]_ , \new_[35903]_ , \new_[35906]_ , \new_[35909]_ ,
    \new_[35910]_ , \new_[35913]_ , \new_[35916]_ , \new_[35917]_ ,
    \new_[35918]_ , \new_[35922]_ , \new_[35923]_ , \new_[35926]_ ,
    \new_[35929]_ , \new_[35930]_ , \new_[35931]_ , \new_[35934]_ ,
    \new_[35937]_ , \new_[35938]_ , \new_[35941]_ , \new_[35944]_ ,
    \new_[35945]_ , \new_[35946]_ , \new_[35950]_ , \new_[35951]_ ,
    \new_[35954]_ , \new_[35957]_ , \new_[35958]_ , \new_[35959]_ ,
    \new_[35962]_ , \new_[35965]_ , \new_[35966]_ , \new_[35969]_ ,
    \new_[35972]_ , \new_[35973]_ , \new_[35974]_ , \new_[35978]_ ,
    \new_[35979]_ , \new_[35982]_ , \new_[35985]_ , \new_[35986]_ ,
    \new_[35987]_ , \new_[35990]_ , \new_[35993]_ , \new_[35994]_ ,
    \new_[35997]_ , \new_[36000]_ , \new_[36001]_ , \new_[36002]_ ,
    \new_[36006]_ , \new_[36007]_ , \new_[36010]_ , \new_[36013]_ ,
    \new_[36014]_ , \new_[36015]_ , \new_[36018]_ , \new_[36021]_ ,
    \new_[36022]_ , \new_[36025]_ , \new_[36028]_ , \new_[36029]_ ,
    \new_[36030]_ , \new_[36034]_ , \new_[36035]_ , \new_[36038]_ ,
    \new_[36041]_ , \new_[36042]_ , \new_[36043]_ , \new_[36046]_ ,
    \new_[36049]_ , \new_[36050]_ , \new_[36053]_ , \new_[36056]_ ,
    \new_[36057]_ , \new_[36058]_ , \new_[36062]_ , \new_[36063]_ ,
    \new_[36066]_ , \new_[36069]_ , \new_[36070]_ , \new_[36071]_ ,
    \new_[36074]_ , \new_[36077]_ , \new_[36078]_ , \new_[36081]_ ,
    \new_[36084]_ , \new_[36085]_ , \new_[36086]_ , \new_[36090]_ ,
    \new_[36091]_ , \new_[36094]_ , \new_[36097]_ , \new_[36098]_ ,
    \new_[36099]_ , \new_[36102]_ , \new_[36105]_ , \new_[36106]_ ,
    \new_[36109]_ , \new_[36112]_ , \new_[36113]_ , \new_[36114]_ ,
    \new_[36118]_ , \new_[36119]_ , \new_[36122]_ , \new_[36125]_ ,
    \new_[36126]_ , \new_[36127]_ , \new_[36130]_ , \new_[36133]_ ,
    \new_[36134]_ , \new_[36137]_ , \new_[36140]_ , \new_[36141]_ ,
    \new_[36142]_ , \new_[36146]_ , \new_[36147]_ , \new_[36150]_ ,
    \new_[36153]_ , \new_[36154]_ , \new_[36155]_ , \new_[36158]_ ,
    \new_[36161]_ , \new_[36162]_ , \new_[36165]_ , \new_[36168]_ ,
    \new_[36169]_ , \new_[36170]_ , \new_[36174]_ , \new_[36175]_ ,
    \new_[36178]_ , \new_[36181]_ , \new_[36182]_ , \new_[36183]_ ,
    \new_[36186]_ , \new_[36189]_ , \new_[36190]_ , \new_[36193]_ ,
    \new_[36196]_ , \new_[36197]_ , \new_[36198]_ , \new_[36202]_ ,
    \new_[36203]_ , \new_[36206]_ , \new_[36209]_ , \new_[36210]_ ,
    \new_[36211]_ , \new_[36214]_ , \new_[36217]_ , \new_[36218]_ ,
    \new_[36221]_ , \new_[36224]_ , \new_[36225]_ , \new_[36226]_ ,
    \new_[36230]_ , \new_[36231]_ , \new_[36234]_ , \new_[36237]_ ,
    \new_[36238]_ , \new_[36239]_ , \new_[36242]_ , \new_[36245]_ ,
    \new_[36246]_ , \new_[36249]_ , \new_[36252]_ , \new_[36253]_ ,
    \new_[36254]_ , \new_[36258]_ , \new_[36259]_ , \new_[36262]_ ,
    \new_[36265]_ , \new_[36266]_ , \new_[36267]_ , \new_[36270]_ ,
    \new_[36273]_ , \new_[36274]_ , \new_[36277]_ , \new_[36280]_ ,
    \new_[36281]_ , \new_[36282]_ , \new_[36286]_ , \new_[36287]_ ,
    \new_[36290]_ , \new_[36293]_ , \new_[36294]_ , \new_[36295]_ ,
    \new_[36298]_ , \new_[36301]_ , \new_[36302]_ , \new_[36305]_ ,
    \new_[36308]_ , \new_[36309]_ , \new_[36310]_ , \new_[36314]_ ,
    \new_[36315]_ , \new_[36318]_ , \new_[36321]_ , \new_[36322]_ ,
    \new_[36323]_ , \new_[36326]_ , \new_[36329]_ , \new_[36330]_ ,
    \new_[36333]_ , \new_[36336]_ , \new_[36337]_ , \new_[36338]_ ,
    \new_[36342]_ , \new_[36343]_ , \new_[36346]_ , \new_[36349]_ ,
    \new_[36350]_ , \new_[36351]_ , \new_[36354]_ , \new_[36357]_ ,
    \new_[36358]_ , \new_[36361]_ , \new_[36364]_ , \new_[36365]_ ,
    \new_[36366]_ , \new_[36370]_ , \new_[36371]_ , \new_[36374]_ ,
    \new_[36377]_ , \new_[36378]_ , \new_[36379]_ , \new_[36382]_ ,
    \new_[36385]_ , \new_[36386]_ , \new_[36389]_ , \new_[36392]_ ,
    \new_[36393]_ , \new_[36394]_ , \new_[36398]_ , \new_[36399]_ ,
    \new_[36402]_ , \new_[36405]_ , \new_[36406]_ , \new_[36407]_ ,
    \new_[36410]_ , \new_[36413]_ , \new_[36414]_ , \new_[36417]_ ,
    \new_[36420]_ , \new_[36421]_ , \new_[36422]_ , \new_[36426]_ ,
    \new_[36427]_ , \new_[36430]_ , \new_[36433]_ , \new_[36434]_ ,
    \new_[36435]_ , \new_[36438]_ , \new_[36441]_ , \new_[36442]_ ,
    \new_[36445]_ , \new_[36448]_ , \new_[36449]_ , \new_[36450]_ ,
    \new_[36454]_ , \new_[36455]_ , \new_[36458]_ , \new_[36461]_ ,
    \new_[36462]_ , \new_[36463]_ , \new_[36466]_ , \new_[36469]_ ,
    \new_[36470]_ , \new_[36473]_ , \new_[36476]_ , \new_[36477]_ ,
    \new_[36478]_ , \new_[36482]_ , \new_[36483]_ , \new_[36486]_ ,
    \new_[36489]_ , \new_[36490]_ , \new_[36491]_ , \new_[36494]_ ,
    \new_[36497]_ , \new_[36498]_ , \new_[36501]_ , \new_[36504]_ ,
    \new_[36505]_ , \new_[36506]_ , \new_[36510]_ , \new_[36511]_ ,
    \new_[36514]_ , \new_[36517]_ , \new_[36518]_ , \new_[36519]_ ,
    \new_[36522]_ , \new_[36525]_ , \new_[36526]_ , \new_[36529]_ ,
    \new_[36532]_ , \new_[36533]_ , \new_[36534]_ , \new_[36538]_ ,
    \new_[36539]_ , \new_[36542]_ , \new_[36545]_ , \new_[36546]_ ,
    \new_[36547]_ , \new_[36550]_ , \new_[36553]_ , \new_[36554]_ ,
    \new_[36557]_ , \new_[36560]_ , \new_[36561]_ , \new_[36562]_ ,
    \new_[36566]_ , \new_[36567]_ , \new_[36570]_ , \new_[36573]_ ,
    \new_[36574]_ , \new_[36575]_ , \new_[36578]_ , \new_[36581]_ ,
    \new_[36582]_ , \new_[36585]_ , \new_[36588]_ , \new_[36589]_ ,
    \new_[36590]_ , \new_[36594]_ , \new_[36595]_ , \new_[36598]_ ,
    \new_[36601]_ , \new_[36602]_ , \new_[36603]_ , \new_[36606]_ ,
    \new_[36609]_ , \new_[36610]_ , \new_[36613]_ , \new_[36616]_ ,
    \new_[36617]_ , \new_[36618]_ , \new_[36622]_ , \new_[36623]_ ,
    \new_[36626]_ , \new_[36629]_ , \new_[36630]_ , \new_[36631]_ ,
    \new_[36634]_ , \new_[36637]_ , \new_[36638]_ , \new_[36641]_ ,
    \new_[36644]_ , \new_[36645]_ , \new_[36646]_ , \new_[36650]_ ,
    \new_[36651]_ , \new_[36654]_ , \new_[36657]_ , \new_[36658]_ ,
    \new_[36659]_ , \new_[36662]_ , \new_[36665]_ , \new_[36666]_ ,
    \new_[36669]_ , \new_[36672]_ , \new_[36673]_ , \new_[36674]_ ,
    \new_[36678]_ , \new_[36679]_ , \new_[36682]_ , \new_[36685]_ ,
    \new_[36686]_ , \new_[36687]_ , \new_[36690]_ , \new_[36693]_ ,
    \new_[36694]_ , \new_[36697]_ , \new_[36700]_ , \new_[36701]_ ,
    \new_[36702]_ , \new_[36706]_ , \new_[36707]_ , \new_[36710]_ ,
    \new_[36713]_ , \new_[36714]_ , \new_[36715]_ , \new_[36718]_ ,
    \new_[36721]_ , \new_[36722]_ , \new_[36725]_ , \new_[36728]_ ,
    \new_[36729]_ , \new_[36730]_ , \new_[36734]_ , \new_[36735]_ ,
    \new_[36738]_ , \new_[36741]_ , \new_[36742]_ , \new_[36743]_ ,
    \new_[36746]_ , \new_[36749]_ , \new_[36750]_ , \new_[36753]_ ,
    \new_[36756]_ , \new_[36757]_ , \new_[36758]_ , \new_[36762]_ ,
    \new_[36763]_ , \new_[36766]_ , \new_[36769]_ , \new_[36770]_ ,
    \new_[36771]_ , \new_[36774]_ , \new_[36777]_ , \new_[36778]_ ,
    \new_[36781]_ , \new_[36784]_ , \new_[36785]_ , \new_[36786]_ ,
    \new_[36790]_ , \new_[36791]_ , \new_[36794]_ , \new_[36797]_ ,
    \new_[36798]_ , \new_[36799]_ , \new_[36802]_ , \new_[36805]_ ,
    \new_[36806]_ , \new_[36809]_ , \new_[36812]_ , \new_[36813]_ ,
    \new_[36814]_ , \new_[36818]_ , \new_[36819]_ , \new_[36822]_ ,
    \new_[36825]_ , \new_[36826]_ , \new_[36827]_ , \new_[36830]_ ,
    \new_[36833]_ , \new_[36834]_ , \new_[36837]_ , \new_[36840]_ ,
    \new_[36841]_ , \new_[36842]_ , \new_[36846]_ , \new_[36847]_ ,
    \new_[36850]_ , \new_[36853]_ , \new_[36854]_ , \new_[36855]_ ,
    \new_[36858]_ , \new_[36861]_ , \new_[36862]_ , \new_[36865]_ ,
    \new_[36868]_ , \new_[36869]_ , \new_[36870]_ , \new_[36874]_ ,
    \new_[36875]_ , \new_[36878]_ , \new_[36881]_ , \new_[36882]_ ,
    \new_[36883]_ , \new_[36886]_ , \new_[36889]_ , \new_[36890]_ ,
    \new_[36893]_ , \new_[36896]_ , \new_[36897]_ , \new_[36898]_ ,
    \new_[36902]_ , \new_[36903]_ , \new_[36906]_ , \new_[36909]_ ,
    \new_[36910]_ , \new_[36911]_ , \new_[36914]_ , \new_[36917]_ ,
    \new_[36918]_ , \new_[36921]_ , \new_[36924]_ , \new_[36925]_ ,
    \new_[36926]_ , \new_[36930]_ , \new_[36931]_ , \new_[36934]_ ,
    \new_[36937]_ , \new_[36938]_ , \new_[36939]_ , \new_[36942]_ ,
    \new_[36945]_ , \new_[36946]_ , \new_[36949]_ , \new_[36952]_ ,
    \new_[36953]_ , \new_[36954]_ , \new_[36958]_ , \new_[36959]_ ,
    \new_[36962]_ , \new_[36965]_ , \new_[36966]_ , \new_[36967]_ ,
    \new_[36970]_ , \new_[36973]_ , \new_[36974]_ , \new_[36977]_ ,
    \new_[36980]_ , \new_[36981]_ , \new_[36982]_ , \new_[36986]_ ,
    \new_[36987]_ , \new_[36990]_ , \new_[36993]_ , \new_[36994]_ ,
    \new_[36995]_ , \new_[36998]_ , \new_[37001]_ , \new_[37002]_ ,
    \new_[37005]_ , \new_[37008]_ , \new_[37009]_ , \new_[37010]_ ,
    \new_[37014]_ , \new_[37015]_ , \new_[37018]_ , \new_[37021]_ ,
    \new_[37022]_ , \new_[37023]_ , \new_[37026]_ , \new_[37029]_ ,
    \new_[37030]_ , \new_[37033]_ , \new_[37036]_ , \new_[37037]_ ,
    \new_[37038]_ , \new_[37042]_ , \new_[37043]_ , \new_[37046]_ ,
    \new_[37049]_ , \new_[37050]_ , \new_[37051]_ , \new_[37054]_ ,
    \new_[37057]_ , \new_[37058]_ , \new_[37061]_ , \new_[37064]_ ,
    \new_[37065]_ , \new_[37066]_ , \new_[37070]_ , \new_[37071]_ ,
    \new_[37074]_ , \new_[37077]_ , \new_[37078]_ , \new_[37079]_ ,
    \new_[37082]_ , \new_[37085]_ , \new_[37086]_ , \new_[37089]_ ,
    \new_[37092]_ , \new_[37093]_ , \new_[37094]_ , \new_[37098]_ ,
    \new_[37099]_ , \new_[37102]_ , \new_[37105]_ , \new_[37106]_ ,
    \new_[37107]_ , \new_[37110]_ , \new_[37113]_ , \new_[37114]_ ,
    \new_[37117]_ , \new_[37120]_ , \new_[37121]_ , \new_[37122]_ ,
    \new_[37126]_ , \new_[37127]_ , \new_[37130]_ , \new_[37133]_ ,
    \new_[37134]_ , \new_[37135]_ , \new_[37138]_ , \new_[37141]_ ,
    \new_[37142]_ , \new_[37145]_ , \new_[37148]_ , \new_[37149]_ ,
    \new_[37150]_ , \new_[37154]_ , \new_[37155]_ , \new_[37158]_ ,
    \new_[37161]_ , \new_[37162]_ , \new_[37163]_ , \new_[37166]_ ,
    \new_[37169]_ , \new_[37170]_ , \new_[37173]_ , \new_[37176]_ ,
    \new_[37177]_ , \new_[37178]_ , \new_[37182]_ , \new_[37183]_ ,
    \new_[37186]_ , \new_[37189]_ , \new_[37190]_ , \new_[37191]_ ,
    \new_[37194]_ , \new_[37197]_ , \new_[37198]_ , \new_[37201]_ ,
    \new_[37204]_ , \new_[37205]_ , \new_[37206]_ , \new_[37210]_ ,
    \new_[37211]_ , \new_[37214]_ , \new_[37217]_ , \new_[37218]_ ,
    \new_[37219]_ , \new_[37222]_ , \new_[37225]_ , \new_[37226]_ ,
    \new_[37229]_ , \new_[37232]_ , \new_[37233]_ , \new_[37234]_ ,
    \new_[37238]_ , \new_[37239]_ , \new_[37242]_ , \new_[37245]_ ,
    \new_[37246]_ , \new_[37247]_ , \new_[37250]_ , \new_[37253]_ ,
    \new_[37254]_ , \new_[37257]_ , \new_[37260]_ , \new_[37261]_ ,
    \new_[37262]_ , \new_[37266]_ , \new_[37267]_ , \new_[37270]_ ,
    \new_[37273]_ , \new_[37274]_ , \new_[37275]_ , \new_[37278]_ ,
    \new_[37281]_ , \new_[37282]_ , \new_[37285]_ , \new_[37288]_ ,
    \new_[37289]_ , \new_[37290]_ , \new_[37294]_ , \new_[37295]_ ,
    \new_[37298]_ , \new_[37301]_ , \new_[37302]_ , \new_[37303]_ ,
    \new_[37306]_ , \new_[37309]_ , \new_[37310]_ , \new_[37313]_ ,
    \new_[37316]_ , \new_[37317]_ , \new_[37318]_ , \new_[37322]_ ,
    \new_[37323]_ , \new_[37326]_ , \new_[37329]_ , \new_[37330]_ ,
    \new_[37331]_ , \new_[37334]_ , \new_[37337]_ , \new_[37338]_ ,
    \new_[37341]_ , \new_[37344]_ , \new_[37345]_ , \new_[37346]_ ,
    \new_[37350]_ , \new_[37351]_ , \new_[37354]_ , \new_[37357]_ ,
    \new_[37358]_ , \new_[37359]_ , \new_[37362]_ , \new_[37365]_ ,
    \new_[37366]_ , \new_[37369]_ , \new_[37372]_ , \new_[37373]_ ,
    \new_[37374]_ , \new_[37378]_ , \new_[37379]_ , \new_[37382]_ ,
    \new_[37385]_ , \new_[37386]_ , \new_[37387]_ , \new_[37390]_ ,
    \new_[37393]_ , \new_[37394]_ , \new_[37397]_ , \new_[37400]_ ,
    \new_[37401]_ , \new_[37402]_ , \new_[37406]_ , \new_[37407]_ ,
    \new_[37410]_ , \new_[37413]_ , \new_[37414]_ , \new_[37415]_ ,
    \new_[37418]_ , \new_[37421]_ , \new_[37422]_ , \new_[37425]_ ,
    \new_[37428]_ , \new_[37429]_ , \new_[37430]_ , \new_[37434]_ ,
    \new_[37435]_ , \new_[37438]_ , \new_[37441]_ , \new_[37442]_ ,
    \new_[37443]_ , \new_[37446]_ , \new_[37449]_ , \new_[37450]_ ,
    \new_[37453]_ , \new_[37456]_ , \new_[37457]_ , \new_[37458]_ ,
    \new_[37462]_ , \new_[37463]_ , \new_[37466]_ , \new_[37469]_ ,
    \new_[37470]_ , \new_[37471]_ , \new_[37474]_ , \new_[37477]_ ,
    \new_[37478]_ , \new_[37481]_ , \new_[37484]_ , \new_[37485]_ ,
    \new_[37486]_ , \new_[37490]_ , \new_[37491]_ , \new_[37494]_ ,
    \new_[37497]_ , \new_[37498]_ , \new_[37499]_ , \new_[37502]_ ,
    \new_[37505]_ , \new_[37506]_ , \new_[37509]_ , \new_[37512]_ ,
    \new_[37513]_ , \new_[37514]_ , \new_[37518]_ , \new_[37519]_ ,
    \new_[37522]_ , \new_[37525]_ , \new_[37526]_ , \new_[37527]_ ,
    \new_[37530]_ , \new_[37533]_ , \new_[37534]_ , \new_[37537]_ ,
    \new_[37540]_ , \new_[37541]_ , \new_[37542]_ , \new_[37546]_ ,
    \new_[37547]_ , \new_[37550]_ , \new_[37553]_ , \new_[37554]_ ,
    \new_[37555]_ , \new_[37558]_ , \new_[37561]_ , \new_[37562]_ ,
    \new_[37565]_ , \new_[37568]_ , \new_[37569]_ , \new_[37570]_ ,
    \new_[37574]_ , \new_[37575]_ , \new_[37578]_ , \new_[37581]_ ,
    \new_[37582]_ , \new_[37583]_ , \new_[37586]_ , \new_[37589]_ ,
    \new_[37590]_ , \new_[37593]_ , \new_[37596]_ , \new_[37597]_ ,
    \new_[37598]_ , \new_[37602]_ , \new_[37603]_ , \new_[37606]_ ,
    \new_[37609]_ , \new_[37610]_ , \new_[37611]_ , \new_[37614]_ ,
    \new_[37617]_ , \new_[37618]_ , \new_[37621]_ , \new_[37624]_ ,
    \new_[37625]_ , \new_[37626]_ , \new_[37630]_ , \new_[37631]_ ,
    \new_[37634]_ , \new_[37637]_ , \new_[37638]_ , \new_[37639]_ ,
    \new_[37642]_ , \new_[37645]_ , \new_[37646]_ , \new_[37649]_ ,
    \new_[37652]_ , \new_[37653]_ , \new_[37654]_ , \new_[37658]_ ,
    \new_[37659]_ , \new_[37662]_ , \new_[37665]_ , \new_[37666]_ ,
    \new_[37667]_ , \new_[37670]_ , \new_[37673]_ , \new_[37674]_ ,
    \new_[37677]_ , \new_[37680]_ , \new_[37681]_ , \new_[37682]_ ,
    \new_[37686]_ , \new_[37687]_ , \new_[37690]_ , \new_[37693]_ ,
    \new_[37694]_ , \new_[37695]_ , \new_[37698]_ , \new_[37701]_ ,
    \new_[37702]_ , \new_[37705]_ , \new_[37708]_ , \new_[37709]_ ,
    \new_[37710]_ , \new_[37714]_ , \new_[37715]_ , \new_[37718]_ ,
    \new_[37721]_ , \new_[37722]_ , \new_[37723]_ , \new_[37726]_ ,
    \new_[37729]_ , \new_[37730]_ , \new_[37733]_ , \new_[37736]_ ,
    \new_[37737]_ , \new_[37738]_ , \new_[37742]_ , \new_[37743]_ ,
    \new_[37746]_ , \new_[37749]_ , \new_[37750]_ , \new_[37751]_ ,
    \new_[37754]_ , \new_[37757]_ , \new_[37758]_ , \new_[37761]_ ,
    \new_[37764]_ , \new_[37765]_ , \new_[37766]_ , \new_[37770]_ ,
    \new_[37771]_ , \new_[37774]_ , \new_[37777]_ , \new_[37778]_ ,
    \new_[37779]_ , \new_[37782]_ , \new_[37785]_ , \new_[37786]_ ,
    \new_[37789]_ , \new_[37792]_ , \new_[37793]_ , \new_[37794]_ ,
    \new_[37798]_ , \new_[37799]_ , \new_[37802]_ , \new_[37805]_ ,
    \new_[37806]_ , \new_[37807]_ , \new_[37810]_ , \new_[37813]_ ,
    \new_[37814]_ , \new_[37817]_ , \new_[37820]_ , \new_[37821]_ ,
    \new_[37822]_ , \new_[37826]_ , \new_[37827]_ , \new_[37830]_ ,
    \new_[37833]_ , \new_[37834]_ , \new_[37835]_ , \new_[37838]_ ,
    \new_[37841]_ , \new_[37842]_ , \new_[37845]_ , \new_[37848]_ ,
    \new_[37849]_ , \new_[37850]_ , \new_[37854]_ , \new_[37855]_ ,
    \new_[37858]_ , \new_[37861]_ , \new_[37862]_ , \new_[37863]_ ,
    \new_[37866]_ , \new_[37869]_ , \new_[37870]_ , \new_[37873]_ ,
    \new_[37876]_ , \new_[37877]_ , \new_[37878]_ , \new_[37882]_ ,
    \new_[37883]_ , \new_[37886]_ , \new_[37889]_ , \new_[37890]_ ,
    \new_[37891]_ , \new_[37894]_ , \new_[37897]_ , \new_[37898]_ ,
    \new_[37901]_ , \new_[37904]_ , \new_[37905]_ , \new_[37906]_ ,
    \new_[37910]_ , \new_[37911]_ , \new_[37914]_ , \new_[37917]_ ,
    \new_[37918]_ , \new_[37919]_ , \new_[37922]_ , \new_[37925]_ ,
    \new_[37926]_ , \new_[37929]_ , \new_[37932]_ , \new_[37933]_ ,
    \new_[37934]_ , \new_[37938]_ , \new_[37939]_ , \new_[37942]_ ,
    \new_[37945]_ , \new_[37946]_ , \new_[37947]_ , \new_[37950]_ ,
    \new_[37953]_ , \new_[37954]_ , \new_[37957]_ , \new_[37960]_ ,
    \new_[37961]_ , \new_[37962]_ , \new_[37966]_ , \new_[37967]_ ,
    \new_[37970]_ , \new_[37973]_ , \new_[37974]_ , \new_[37975]_ ,
    \new_[37978]_ , \new_[37981]_ , \new_[37982]_ , \new_[37985]_ ,
    \new_[37988]_ , \new_[37989]_ , \new_[37990]_ , \new_[37994]_ ,
    \new_[37995]_ , \new_[37998]_ , \new_[38001]_ , \new_[38002]_ ,
    \new_[38003]_ , \new_[38006]_ , \new_[38009]_ , \new_[38010]_ ,
    \new_[38013]_ , \new_[38016]_ , \new_[38017]_ , \new_[38018]_ ,
    \new_[38021]_ , \new_[38024]_ , \new_[38025]_ , \new_[38028]_ ,
    \new_[38031]_ , \new_[38032]_ , \new_[38033]_ , \new_[38036]_ ,
    \new_[38039]_ , \new_[38040]_ , \new_[38043]_ , \new_[38046]_ ,
    \new_[38047]_ , \new_[38048]_ , \new_[38051]_ , \new_[38054]_ ,
    \new_[38055]_ , \new_[38058]_ , \new_[38061]_ , \new_[38062]_ ,
    \new_[38063]_ , \new_[38066]_ , \new_[38069]_ , \new_[38070]_ ,
    \new_[38073]_ , \new_[38076]_ , \new_[38077]_ , \new_[38078]_ ,
    \new_[38081]_ , \new_[38084]_ , \new_[38085]_ , \new_[38088]_ ,
    \new_[38091]_ , \new_[38092]_ , \new_[38093]_ , \new_[38096]_ ,
    \new_[38099]_ , \new_[38100]_ , \new_[38103]_ , \new_[38106]_ ,
    \new_[38107]_ , \new_[38108]_ , \new_[38111]_ , \new_[38114]_ ,
    \new_[38115]_ , \new_[38118]_ , \new_[38121]_ , \new_[38122]_ ,
    \new_[38123]_ , \new_[38126]_ , \new_[38129]_ , \new_[38130]_ ,
    \new_[38133]_ , \new_[38136]_ , \new_[38137]_ , \new_[38138]_ ,
    \new_[38141]_ , \new_[38144]_ , \new_[38145]_ , \new_[38148]_ ,
    \new_[38151]_ , \new_[38152]_ , \new_[38153]_ , \new_[38156]_ ,
    \new_[38159]_ , \new_[38160]_ , \new_[38163]_ , \new_[38166]_ ,
    \new_[38167]_ , \new_[38168]_ , \new_[38171]_ , \new_[38174]_ ,
    \new_[38175]_ , \new_[38178]_ , \new_[38181]_ , \new_[38182]_ ,
    \new_[38183]_ , \new_[38186]_ , \new_[38189]_ , \new_[38190]_ ,
    \new_[38193]_ , \new_[38196]_ , \new_[38197]_ , \new_[38198]_ ,
    \new_[38201]_ , \new_[38204]_ , \new_[38205]_ , \new_[38208]_ ,
    \new_[38211]_ , \new_[38212]_ , \new_[38213]_ , \new_[38216]_ ,
    \new_[38219]_ , \new_[38220]_ , \new_[38223]_ , \new_[38226]_ ,
    \new_[38227]_ , \new_[38228]_ , \new_[38231]_ , \new_[38234]_ ,
    \new_[38235]_ , \new_[38238]_ , \new_[38241]_ , \new_[38242]_ ,
    \new_[38243]_ , \new_[38246]_ , \new_[38249]_ , \new_[38250]_ ,
    \new_[38253]_ , \new_[38256]_ , \new_[38257]_ , \new_[38258]_ ,
    \new_[38261]_ , \new_[38264]_ , \new_[38265]_ , \new_[38268]_ ,
    \new_[38271]_ , \new_[38272]_ , \new_[38273]_ , \new_[38276]_ ,
    \new_[38279]_ , \new_[38280]_ , \new_[38283]_ , \new_[38286]_ ,
    \new_[38287]_ , \new_[38288]_ , \new_[38291]_ , \new_[38294]_ ,
    \new_[38295]_ , \new_[38298]_ , \new_[38301]_ , \new_[38302]_ ,
    \new_[38303]_ , \new_[38306]_ , \new_[38309]_ , \new_[38310]_ ,
    \new_[38313]_ , \new_[38316]_ , \new_[38317]_ , \new_[38318]_ ,
    \new_[38321]_ , \new_[38324]_ , \new_[38325]_ , \new_[38328]_ ,
    \new_[38331]_ , \new_[38332]_ , \new_[38333]_ , \new_[38336]_ ,
    \new_[38339]_ , \new_[38340]_ , \new_[38343]_ , \new_[38346]_ ,
    \new_[38347]_ , \new_[38348]_ , \new_[38351]_ , \new_[38354]_ ,
    \new_[38355]_ , \new_[38358]_ , \new_[38361]_ , \new_[38362]_ ,
    \new_[38363]_ , \new_[38366]_ , \new_[38369]_ , \new_[38370]_ ,
    \new_[38373]_ , \new_[38376]_ , \new_[38377]_ , \new_[38378]_ ,
    \new_[38381]_ , \new_[38384]_ , \new_[38385]_ , \new_[38388]_ ,
    \new_[38391]_ , \new_[38392]_ , \new_[38393]_ , \new_[38396]_ ,
    \new_[38399]_ , \new_[38400]_ , \new_[38403]_ , \new_[38406]_ ,
    \new_[38407]_ , \new_[38408]_ , \new_[38411]_ , \new_[38414]_ ,
    \new_[38415]_ , \new_[38418]_ , \new_[38421]_ , \new_[38422]_ ,
    \new_[38423]_ , \new_[38426]_ , \new_[38429]_ , \new_[38430]_ ,
    \new_[38433]_ , \new_[38436]_ , \new_[38437]_ , \new_[38438]_ ,
    \new_[38441]_ , \new_[38444]_ , \new_[38445]_ , \new_[38448]_ ,
    \new_[38451]_ , \new_[38452]_ , \new_[38453]_ , \new_[38456]_ ,
    \new_[38459]_ , \new_[38460]_ , \new_[38463]_ , \new_[38466]_ ,
    \new_[38467]_ , \new_[38468]_ , \new_[38471]_ , \new_[38474]_ ,
    \new_[38475]_ , \new_[38478]_ , \new_[38481]_ , \new_[38482]_ ,
    \new_[38483]_ , \new_[38486]_ , \new_[38489]_ , \new_[38490]_ ,
    \new_[38493]_ , \new_[38496]_ , \new_[38497]_ , \new_[38498]_ ,
    \new_[38501]_ , \new_[38504]_ , \new_[38505]_ , \new_[38508]_ ,
    \new_[38511]_ , \new_[38512]_ , \new_[38513]_ , \new_[38516]_ ,
    \new_[38519]_ , \new_[38520]_ , \new_[38523]_ , \new_[38526]_ ,
    \new_[38527]_ , \new_[38528]_ , \new_[38531]_ , \new_[38534]_ ,
    \new_[38535]_ , \new_[38538]_ , \new_[38541]_ , \new_[38542]_ ,
    \new_[38543]_ , \new_[38546]_ , \new_[38549]_ , \new_[38550]_ ,
    \new_[38553]_ , \new_[38556]_ , \new_[38557]_ , \new_[38558]_ ,
    \new_[38561]_ , \new_[38564]_ , \new_[38565]_ , \new_[38568]_ ,
    \new_[38571]_ , \new_[38572]_ , \new_[38573]_ , \new_[38576]_ ,
    \new_[38579]_ , \new_[38580]_ , \new_[38583]_ , \new_[38586]_ ,
    \new_[38587]_ , \new_[38588]_ , \new_[38591]_ , \new_[38594]_ ,
    \new_[38595]_ , \new_[38598]_ , \new_[38601]_ , \new_[38602]_ ,
    \new_[38603]_ , \new_[38606]_ , \new_[38609]_ , \new_[38610]_ ,
    \new_[38613]_ , \new_[38616]_ , \new_[38617]_ , \new_[38618]_ ,
    \new_[38621]_ , \new_[38624]_ , \new_[38625]_ , \new_[38628]_ ,
    \new_[38631]_ , \new_[38632]_ , \new_[38633]_ , \new_[38636]_ ,
    \new_[38639]_ , \new_[38640]_ , \new_[38643]_ , \new_[38646]_ ,
    \new_[38647]_ , \new_[38648]_ , \new_[38651]_ , \new_[38654]_ ,
    \new_[38655]_ , \new_[38658]_ , \new_[38661]_ , \new_[38662]_ ,
    \new_[38663]_ , \new_[38666]_ , \new_[38669]_ , \new_[38670]_ ,
    \new_[38673]_ , \new_[38676]_ , \new_[38677]_ , \new_[38678]_ ,
    \new_[38681]_ , \new_[38684]_ , \new_[38685]_ , \new_[38688]_ ,
    \new_[38691]_ , \new_[38692]_ , \new_[38693]_ , \new_[38696]_ ,
    \new_[38699]_ , \new_[38700]_ , \new_[38703]_ , \new_[38706]_ ,
    \new_[38707]_ , \new_[38708]_ , \new_[38711]_ , \new_[38714]_ ,
    \new_[38715]_ , \new_[38718]_ , \new_[38721]_ , \new_[38722]_ ,
    \new_[38723]_ , \new_[38726]_ , \new_[38729]_ , \new_[38730]_ ,
    \new_[38733]_ , \new_[38736]_ , \new_[38737]_ , \new_[38738]_ ,
    \new_[38741]_ , \new_[38744]_ , \new_[38745]_ , \new_[38748]_ ,
    \new_[38751]_ , \new_[38752]_ , \new_[38753]_ , \new_[38756]_ ,
    \new_[38759]_ , \new_[38760]_ , \new_[38763]_ , \new_[38766]_ ,
    \new_[38767]_ , \new_[38768]_ , \new_[38771]_ , \new_[38774]_ ,
    \new_[38775]_ , \new_[38778]_ , \new_[38781]_ , \new_[38782]_ ,
    \new_[38783]_ , \new_[38786]_ , \new_[38789]_ , \new_[38790]_ ,
    \new_[38793]_ , \new_[38796]_ , \new_[38797]_ , \new_[38798]_ ,
    \new_[38801]_ , \new_[38804]_ , \new_[38805]_ , \new_[38808]_ ,
    \new_[38811]_ , \new_[38812]_ , \new_[38813]_ , \new_[38816]_ ,
    \new_[38819]_ , \new_[38820]_ , \new_[38823]_ , \new_[38826]_ ,
    \new_[38827]_ , \new_[38828]_ , \new_[38831]_ , \new_[38834]_ ,
    \new_[38835]_ , \new_[38838]_ , \new_[38841]_ , \new_[38842]_ ,
    \new_[38843]_ , \new_[38846]_ , \new_[38849]_ , \new_[38850]_ ,
    \new_[38853]_ , \new_[38856]_ , \new_[38857]_ , \new_[38858]_ ,
    \new_[38861]_ , \new_[38864]_ , \new_[38865]_ , \new_[38868]_ ,
    \new_[38871]_ , \new_[38872]_ , \new_[38873]_ , \new_[38876]_ ,
    \new_[38879]_ , \new_[38880]_ , \new_[38883]_ , \new_[38886]_ ,
    \new_[38887]_ , \new_[38888]_ , \new_[38891]_ , \new_[38894]_ ,
    \new_[38895]_ , \new_[38898]_ , \new_[38901]_ , \new_[38902]_ ,
    \new_[38903]_ , \new_[38906]_ , \new_[38909]_ , \new_[38910]_ ,
    \new_[38913]_ , \new_[38916]_ , \new_[38917]_ , \new_[38918]_ ,
    \new_[38921]_ , \new_[38924]_ , \new_[38925]_ , \new_[38928]_ ,
    \new_[38931]_ , \new_[38932]_ , \new_[38933]_ , \new_[38936]_ ,
    \new_[38939]_ , \new_[38940]_ , \new_[38943]_ , \new_[38946]_ ,
    \new_[38947]_ , \new_[38948]_ , \new_[38951]_ , \new_[38954]_ ,
    \new_[38955]_ , \new_[38958]_ , \new_[38961]_ , \new_[38962]_ ,
    \new_[38963]_ , \new_[38966]_ , \new_[38969]_ , \new_[38970]_ ,
    \new_[38973]_ , \new_[38976]_ , \new_[38977]_ , \new_[38978]_ ,
    \new_[38981]_ , \new_[38984]_ , \new_[38985]_ , \new_[38988]_ ,
    \new_[38991]_ , \new_[38992]_ , \new_[38993]_ , \new_[38996]_ ,
    \new_[38999]_ , \new_[39000]_ , \new_[39003]_ , \new_[39006]_ ,
    \new_[39007]_ , \new_[39008]_ , \new_[39011]_ , \new_[39014]_ ,
    \new_[39015]_ , \new_[39018]_ , \new_[39021]_ , \new_[39022]_ ,
    \new_[39023]_ , \new_[39026]_ , \new_[39029]_ , \new_[39030]_ ,
    \new_[39033]_ , \new_[39036]_ , \new_[39037]_ , \new_[39038]_ ,
    \new_[39041]_ , \new_[39044]_ , \new_[39045]_ , \new_[39048]_ ,
    \new_[39051]_ , \new_[39052]_ , \new_[39053]_ , \new_[39056]_ ,
    \new_[39059]_ , \new_[39060]_ , \new_[39063]_ , \new_[39066]_ ,
    \new_[39067]_ , \new_[39068]_ , \new_[39071]_ , \new_[39074]_ ,
    \new_[39075]_ , \new_[39078]_ , \new_[39081]_ , \new_[39082]_ ,
    \new_[39083]_ , \new_[39086]_ , \new_[39089]_ , \new_[39090]_ ,
    \new_[39093]_ , \new_[39096]_ , \new_[39097]_ , \new_[39098]_ ,
    \new_[39101]_ , \new_[39104]_ , \new_[39105]_ , \new_[39108]_ ,
    \new_[39111]_ , \new_[39112]_ , \new_[39113]_ , \new_[39116]_ ,
    \new_[39119]_ , \new_[39120]_ , \new_[39123]_ , \new_[39126]_ ,
    \new_[39127]_ , \new_[39128]_ , \new_[39131]_ , \new_[39134]_ ,
    \new_[39135]_ , \new_[39138]_ , \new_[39141]_ , \new_[39142]_ ,
    \new_[39143]_ , \new_[39146]_ , \new_[39149]_ , \new_[39150]_ ,
    \new_[39153]_ , \new_[39156]_ , \new_[39157]_ , \new_[39158]_ ,
    \new_[39161]_ , \new_[39164]_ , \new_[39165]_ , \new_[39168]_ ,
    \new_[39171]_ , \new_[39172]_ , \new_[39173]_ , \new_[39176]_ ,
    \new_[39179]_ , \new_[39180]_ , \new_[39183]_ , \new_[39186]_ ,
    \new_[39187]_ , \new_[39188]_ , \new_[39191]_ , \new_[39194]_ ,
    \new_[39195]_ , \new_[39198]_ , \new_[39201]_ , \new_[39202]_ ,
    \new_[39203]_ , \new_[39206]_ , \new_[39209]_ , \new_[39210]_ ,
    \new_[39213]_ , \new_[39216]_ , \new_[39217]_ , \new_[39218]_ ,
    \new_[39221]_ , \new_[39224]_ , \new_[39225]_ , \new_[39228]_ ,
    \new_[39231]_ , \new_[39232]_ , \new_[39233]_ , \new_[39236]_ ,
    \new_[39239]_ , \new_[39240]_ , \new_[39243]_ , \new_[39246]_ ,
    \new_[39247]_ , \new_[39248]_ , \new_[39251]_ , \new_[39254]_ ,
    \new_[39255]_ , \new_[39258]_ , \new_[39261]_ , \new_[39262]_ ,
    \new_[39263]_ , \new_[39266]_ , \new_[39269]_ , \new_[39270]_ ,
    \new_[39273]_ , \new_[39276]_ , \new_[39277]_ , \new_[39278]_ ,
    \new_[39281]_ , \new_[39284]_ , \new_[39285]_ , \new_[39288]_ ,
    \new_[39291]_ , \new_[39292]_ , \new_[39293]_ , \new_[39296]_ ,
    \new_[39299]_ , \new_[39300]_ , \new_[39303]_ , \new_[39306]_ ,
    \new_[39307]_ , \new_[39308]_ , \new_[39311]_ , \new_[39314]_ ,
    \new_[39315]_ , \new_[39318]_ , \new_[39321]_ , \new_[39322]_ ,
    \new_[39323]_ , \new_[39326]_ , \new_[39329]_ , \new_[39330]_ ,
    \new_[39333]_ , \new_[39336]_ , \new_[39337]_ , \new_[39338]_ ,
    \new_[39341]_ , \new_[39344]_ , \new_[39345]_ , \new_[39348]_ ,
    \new_[39351]_ , \new_[39352]_ , \new_[39353]_ , \new_[39356]_ ,
    \new_[39359]_ , \new_[39360]_ , \new_[39363]_ , \new_[39366]_ ,
    \new_[39367]_ , \new_[39368]_ , \new_[39371]_ , \new_[39374]_ ,
    \new_[39375]_ , \new_[39378]_ , \new_[39381]_ , \new_[39382]_ ,
    \new_[39383]_ , \new_[39386]_ , \new_[39389]_ , \new_[39390]_ ,
    \new_[39393]_ , \new_[39396]_ , \new_[39397]_ , \new_[39398]_ ,
    \new_[39401]_ , \new_[39404]_ , \new_[39405]_ , \new_[39408]_ ,
    \new_[39411]_ , \new_[39412]_ , \new_[39413]_ , \new_[39416]_ ,
    \new_[39419]_ , \new_[39420]_ , \new_[39423]_ , \new_[39426]_ ,
    \new_[39427]_ , \new_[39428]_ , \new_[39431]_ , \new_[39434]_ ,
    \new_[39435]_ , \new_[39438]_ , \new_[39441]_ , \new_[39442]_ ,
    \new_[39443]_ , \new_[39446]_ , \new_[39449]_ , \new_[39450]_ ,
    \new_[39453]_ , \new_[39456]_ , \new_[39457]_ , \new_[39458]_ ,
    \new_[39461]_ , \new_[39464]_ , \new_[39465]_ , \new_[39468]_ ,
    \new_[39471]_ , \new_[39472]_ , \new_[39473]_ , \new_[39476]_ ,
    \new_[39479]_ , \new_[39480]_ , \new_[39483]_ , \new_[39486]_ ,
    \new_[39487]_ , \new_[39488]_ , \new_[39491]_ , \new_[39494]_ ,
    \new_[39495]_ , \new_[39498]_ , \new_[39501]_ , \new_[39502]_ ,
    \new_[39503]_ , \new_[39506]_ , \new_[39509]_ , \new_[39510]_ ,
    \new_[39513]_ , \new_[39516]_ , \new_[39517]_ , \new_[39518]_ ,
    \new_[39521]_ , \new_[39524]_ , \new_[39525]_ , \new_[39528]_ ,
    \new_[39531]_ , \new_[39532]_ , \new_[39533]_ , \new_[39536]_ ,
    \new_[39539]_ , \new_[39540]_ , \new_[39543]_ , \new_[39546]_ ,
    \new_[39547]_ , \new_[39548]_ , \new_[39551]_ , \new_[39554]_ ,
    \new_[39555]_ , \new_[39558]_ , \new_[39561]_ , \new_[39562]_ ,
    \new_[39563]_ , \new_[39566]_ , \new_[39569]_ , \new_[39570]_ ,
    \new_[39573]_ , \new_[39576]_ , \new_[39577]_ , \new_[39578]_ ,
    \new_[39581]_ , \new_[39584]_ , \new_[39585]_ , \new_[39588]_ ,
    \new_[39591]_ , \new_[39592]_ , \new_[39593]_ , \new_[39596]_ ,
    \new_[39599]_ , \new_[39600]_ , \new_[39603]_ , \new_[39606]_ ,
    \new_[39607]_ , \new_[39608]_ , \new_[39611]_ , \new_[39614]_ ,
    \new_[39615]_ , \new_[39618]_ , \new_[39621]_ , \new_[39622]_ ,
    \new_[39623]_ , \new_[39626]_ , \new_[39629]_ , \new_[39630]_ ,
    \new_[39633]_ , \new_[39636]_ , \new_[39637]_ , \new_[39638]_ ,
    \new_[39641]_ , \new_[39644]_ , \new_[39645]_ , \new_[39648]_ ,
    \new_[39651]_ , \new_[39652]_ , \new_[39653]_ , \new_[39656]_ ,
    \new_[39659]_ , \new_[39660]_ , \new_[39663]_ , \new_[39666]_ ,
    \new_[39667]_ , \new_[39668]_ , \new_[39671]_ , \new_[39674]_ ,
    \new_[39675]_ , \new_[39678]_ , \new_[39681]_ , \new_[39682]_ ,
    \new_[39683]_ , \new_[39686]_ , \new_[39689]_ , \new_[39690]_ ,
    \new_[39693]_ , \new_[39696]_ , \new_[39697]_ , \new_[39698]_ ,
    \new_[39701]_ , \new_[39704]_ , \new_[39705]_ , \new_[39708]_ ,
    \new_[39711]_ , \new_[39712]_ , \new_[39713]_ , \new_[39716]_ ,
    \new_[39719]_ , \new_[39720]_ , \new_[39723]_ , \new_[39726]_ ,
    \new_[39727]_ , \new_[39728]_ , \new_[39731]_ , \new_[39734]_ ,
    \new_[39735]_ , \new_[39738]_ , \new_[39741]_ , \new_[39742]_ ,
    \new_[39743]_ , \new_[39746]_ , \new_[39749]_ , \new_[39750]_ ,
    \new_[39753]_ , \new_[39756]_ , \new_[39757]_ , \new_[39758]_ ,
    \new_[39761]_ , \new_[39764]_ , \new_[39765]_ , \new_[39768]_ ,
    \new_[39771]_ , \new_[39772]_ , \new_[39773]_ , \new_[39776]_ ,
    \new_[39779]_ , \new_[39780]_ , \new_[39783]_ , \new_[39786]_ ,
    \new_[39787]_ , \new_[39788]_ , \new_[39791]_ , \new_[39794]_ ,
    \new_[39795]_ , \new_[39798]_ , \new_[39801]_ , \new_[39802]_ ,
    \new_[39803]_ , \new_[39806]_ , \new_[39809]_ , \new_[39810]_ ,
    \new_[39813]_ , \new_[39816]_ , \new_[39817]_ , \new_[39818]_ ,
    \new_[39821]_ , \new_[39824]_ , \new_[39825]_ , \new_[39828]_ ,
    \new_[39831]_ , \new_[39832]_ , \new_[39833]_ , \new_[39836]_ ,
    \new_[39839]_ , \new_[39840]_ , \new_[39843]_ , \new_[39846]_ ,
    \new_[39847]_ , \new_[39848]_ , \new_[39851]_ , \new_[39854]_ ,
    \new_[39855]_ , \new_[39858]_ , \new_[39861]_ , \new_[39862]_ ,
    \new_[39863]_ , \new_[39866]_ , \new_[39869]_ , \new_[39870]_ ,
    \new_[39873]_ , \new_[39876]_ , \new_[39877]_ , \new_[39878]_ ,
    \new_[39881]_ , \new_[39884]_ , \new_[39885]_ , \new_[39888]_ ,
    \new_[39891]_ , \new_[39892]_ , \new_[39893]_ , \new_[39896]_ ,
    \new_[39899]_ , \new_[39900]_ , \new_[39903]_ , \new_[39906]_ ,
    \new_[39907]_ , \new_[39908]_ , \new_[39911]_ , \new_[39914]_ ,
    \new_[39915]_ , \new_[39918]_ , \new_[39921]_ , \new_[39922]_ ,
    \new_[39923]_ , \new_[39926]_ , \new_[39929]_ , \new_[39930]_ ,
    \new_[39933]_ , \new_[39936]_ , \new_[39937]_ , \new_[39938]_ ,
    \new_[39941]_ , \new_[39944]_ , \new_[39945]_ , \new_[39948]_ ,
    \new_[39951]_ , \new_[39952]_ , \new_[39953]_ , \new_[39956]_ ,
    \new_[39959]_ , \new_[39960]_ , \new_[39963]_ , \new_[39966]_ ,
    \new_[39967]_ , \new_[39968]_ , \new_[39971]_ , \new_[39974]_ ,
    \new_[39975]_ , \new_[39978]_ , \new_[39981]_ , \new_[39982]_ ,
    \new_[39983]_ , \new_[39986]_ , \new_[39989]_ , \new_[39990]_ ,
    \new_[39993]_ , \new_[39996]_ , \new_[39997]_ , \new_[39998]_ ,
    \new_[40001]_ , \new_[40004]_ , \new_[40005]_ , \new_[40008]_ ,
    \new_[40011]_ , \new_[40012]_ , \new_[40013]_ , \new_[40016]_ ,
    \new_[40019]_ , \new_[40020]_ , \new_[40023]_ , \new_[40026]_ ,
    \new_[40027]_ , \new_[40028]_ , \new_[40031]_ , \new_[40034]_ ,
    \new_[40035]_ , \new_[40038]_ , \new_[40041]_ , \new_[40042]_ ,
    \new_[40043]_ , \new_[40046]_ , \new_[40049]_ , \new_[40050]_ ,
    \new_[40053]_ , \new_[40056]_ , \new_[40057]_ , \new_[40058]_ ,
    \new_[40061]_ , \new_[40064]_ , \new_[40065]_ , \new_[40068]_ ,
    \new_[40071]_ , \new_[40072]_ , \new_[40073]_ , \new_[40076]_ ,
    \new_[40079]_ , \new_[40080]_ , \new_[40083]_ , \new_[40086]_ ,
    \new_[40087]_ , \new_[40088]_ , \new_[40091]_ , \new_[40094]_ ,
    \new_[40095]_ , \new_[40098]_ , \new_[40101]_ , \new_[40102]_ ,
    \new_[40103]_ , \new_[40106]_ , \new_[40109]_ , \new_[40110]_ ,
    \new_[40113]_ , \new_[40116]_ , \new_[40117]_ , \new_[40118]_ ,
    \new_[40121]_ , \new_[40124]_ , \new_[40125]_ , \new_[40128]_ ,
    \new_[40131]_ , \new_[40132]_ , \new_[40133]_ , \new_[40136]_ ,
    \new_[40139]_ , \new_[40140]_ , \new_[40143]_ , \new_[40146]_ ,
    \new_[40147]_ , \new_[40148]_ , \new_[40151]_ , \new_[40154]_ ,
    \new_[40155]_ , \new_[40158]_ , \new_[40161]_ , \new_[40162]_ ,
    \new_[40163]_ , \new_[40166]_ , \new_[40169]_ , \new_[40170]_ ,
    \new_[40173]_ , \new_[40176]_ , \new_[40177]_ , \new_[40178]_ ,
    \new_[40181]_ , \new_[40184]_ , \new_[40185]_ , \new_[40188]_ ,
    \new_[40191]_ , \new_[40192]_ , \new_[40193]_ , \new_[40196]_ ,
    \new_[40199]_ , \new_[40200]_ , \new_[40203]_ , \new_[40206]_ ,
    \new_[40207]_ , \new_[40208]_ , \new_[40211]_ , \new_[40214]_ ,
    \new_[40215]_ , \new_[40218]_ , \new_[40221]_ , \new_[40222]_ ,
    \new_[40223]_ , \new_[40226]_ , \new_[40229]_ , \new_[40230]_ ,
    \new_[40233]_ , \new_[40236]_ , \new_[40237]_ , \new_[40238]_ ,
    \new_[40241]_ , \new_[40244]_ , \new_[40245]_ , \new_[40248]_ ,
    \new_[40251]_ , \new_[40252]_ , \new_[40253]_ , \new_[40256]_ ,
    \new_[40259]_ , \new_[40260]_ , \new_[40263]_ , \new_[40266]_ ,
    \new_[40267]_ , \new_[40268]_ , \new_[40271]_ , \new_[40274]_ ,
    \new_[40275]_ , \new_[40278]_ , \new_[40281]_ , \new_[40282]_ ,
    \new_[40283]_ , \new_[40286]_ , \new_[40289]_ , \new_[40290]_ ,
    \new_[40293]_ , \new_[40296]_ , \new_[40297]_ , \new_[40298]_ ,
    \new_[40301]_ , \new_[40304]_ , \new_[40305]_ , \new_[40308]_ ,
    \new_[40311]_ , \new_[40312]_ , \new_[40313]_ , \new_[40316]_ ,
    \new_[40319]_ , \new_[40320]_ , \new_[40323]_ , \new_[40326]_ ,
    \new_[40327]_ , \new_[40328]_ , \new_[40331]_ , \new_[40334]_ ,
    \new_[40335]_ , \new_[40338]_ , \new_[40341]_ , \new_[40342]_ ,
    \new_[40343]_ , \new_[40346]_ , \new_[40349]_ , \new_[40350]_ ,
    \new_[40353]_ , \new_[40356]_ , \new_[40357]_ , \new_[40358]_ ,
    \new_[40361]_ , \new_[40364]_ , \new_[40365]_ , \new_[40368]_ ,
    \new_[40371]_ , \new_[40372]_ , \new_[40373]_ , \new_[40376]_ ,
    \new_[40379]_ , \new_[40380]_ , \new_[40383]_ , \new_[40386]_ ,
    \new_[40387]_ , \new_[40388]_ , \new_[40391]_ , \new_[40394]_ ,
    \new_[40395]_ , \new_[40398]_ , \new_[40401]_ , \new_[40402]_ ,
    \new_[40403]_ , \new_[40406]_ , \new_[40409]_ , \new_[40410]_ ,
    \new_[40413]_ , \new_[40416]_ , \new_[40417]_ , \new_[40418]_ ,
    \new_[40421]_ , \new_[40424]_ , \new_[40425]_ , \new_[40428]_ ,
    \new_[40431]_ , \new_[40432]_ , \new_[40433]_ , \new_[40436]_ ,
    \new_[40439]_ , \new_[40440]_ , \new_[40443]_ , \new_[40446]_ ,
    \new_[40447]_ , \new_[40448]_ , \new_[40451]_ , \new_[40454]_ ,
    \new_[40455]_ , \new_[40458]_ , \new_[40461]_ , \new_[40462]_ ,
    \new_[40463]_ , \new_[40466]_ , \new_[40469]_ , \new_[40470]_ ,
    \new_[40473]_ , \new_[40476]_ , \new_[40477]_ , \new_[40478]_ ,
    \new_[40481]_ , \new_[40484]_ , \new_[40485]_ , \new_[40488]_ ,
    \new_[40491]_ , \new_[40492]_ , \new_[40493]_ , \new_[40496]_ ,
    \new_[40499]_ , \new_[40500]_ , \new_[40503]_ , \new_[40506]_ ,
    \new_[40507]_ , \new_[40508]_ , \new_[40511]_ , \new_[40514]_ ,
    \new_[40515]_ , \new_[40518]_ , \new_[40521]_ , \new_[40522]_ ,
    \new_[40523]_ , \new_[40526]_ , \new_[40529]_ , \new_[40530]_ ,
    \new_[40533]_ , \new_[40536]_ , \new_[40537]_ , \new_[40538]_ ,
    \new_[40541]_ , \new_[40544]_ , \new_[40545]_ , \new_[40548]_ ,
    \new_[40551]_ , \new_[40552]_ , \new_[40553]_ , \new_[40556]_ ,
    \new_[40559]_ , \new_[40560]_ , \new_[40563]_ , \new_[40566]_ ,
    \new_[40567]_ , \new_[40568]_ , \new_[40571]_ , \new_[40574]_ ,
    \new_[40575]_ , \new_[40578]_ , \new_[40581]_ , \new_[40582]_ ,
    \new_[40583]_ , \new_[40586]_ , \new_[40589]_ , \new_[40590]_ ,
    \new_[40593]_ , \new_[40596]_ , \new_[40597]_ , \new_[40598]_ ,
    \new_[40601]_ , \new_[40604]_ , \new_[40605]_ , \new_[40608]_ ,
    \new_[40611]_ , \new_[40612]_ , \new_[40613]_ , \new_[40616]_ ,
    \new_[40619]_ , \new_[40620]_ , \new_[40623]_ , \new_[40626]_ ,
    \new_[40627]_ , \new_[40628]_ , \new_[40631]_ , \new_[40634]_ ,
    \new_[40635]_ , \new_[40638]_ , \new_[40641]_ , \new_[40642]_ ,
    \new_[40643]_ , \new_[40646]_ , \new_[40649]_ , \new_[40650]_ ,
    \new_[40653]_ , \new_[40656]_ , \new_[40657]_ , \new_[40658]_ ,
    \new_[40661]_ , \new_[40664]_ , \new_[40665]_ , \new_[40668]_ ,
    \new_[40671]_ , \new_[40672]_ , \new_[40673]_ , \new_[40676]_ ,
    \new_[40679]_ , \new_[40680]_ , \new_[40683]_ , \new_[40686]_ ,
    \new_[40687]_ , \new_[40688]_ , \new_[40691]_ , \new_[40694]_ ,
    \new_[40695]_ , \new_[40698]_ , \new_[40701]_ , \new_[40702]_ ,
    \new_[40703]_ , \new_[40706]_ , \new_[40709]_ , \new_[40710]_ ,
    \new_[40713]_ , \new_[40716]_ , \new_[40717]_ , \new_[40718]_ ,
    \new_[40721]_ , \new_[40724]_ , \new_[40725]_ , \new_[40728]_ ,
    \new_[40731]_ , \new_[40732]_ , \new_[40733]_ , \new_[40736]_ ,
    \new_[40739]_ , \new_[40740]_ , \new_[40743]_ , \new_[40746]_ ,
    \new_[40747]_ , \new_[40748]_ , \new_[40751]_ , \new_[40754]_ ,
    \new_[40755]_ , \new_[40758]_ , \new_[40761]_ , \new_[40762]_ ,
    \new_[40763]_ , \new_[40766]_ , \new_[40769]_ , \new_[40770]_ ,
    \new_[40773]_ , \new_[40776]_ , \new_[40777]_ , \new_[40778]_ ,
    \new_[40781]_ , \new_[40784]_ , \new_[40785]_ , \new_[40788]_ ,
    \new_[40791]_ , \new_[40792]_ , \new_[40793]_ , \new_[40796]_ ,
    \new_[40799]_ , \new_[40800]_ , \new_[40803]_ , \new_[40806]_ ,
    \new_[40807]_ , \new_[40808]_ , \new_[40811]_ , \new_[40814]_ ,
    \new_[40815]_ , \new_[40818]_ , \new_[40821]_ , \new_[40822]_ ,
    \new_[40823]_ , \new_[40826]_ , \new_[40829]_ , \new_[40830]_ ,
    \new_[40833]_ , \new_[40836]_ , \new_[40837]_ , \new_[40838]_ ,
    \new_[40841]_ , \new_[40844]_ , \new_[40845]_ , \new_[40848]_ ,
    \new_[40851]_ , \new_[40852]_ , \new_[40853]_ , \new_[40856]_ ,
    \new_[40859]_ , \new_[40860]_ , \new_[40863]_ , \new_[40866]_ ,
    \new_[40867]_ , \new_[40868]_ , \new_[40871]_ , \new_[40874]_ ,
    \new_[40875]_ , \new_[40878]_ , \new_[40881]_ , \new_[40882]_ ,
    \new_[40883]_ , \new_[40886]_ , \new_[40889]_ , \new_[40890]_ ,
    \new_[40893]_ , \new_[40896]_ , \new_[40897]_ , \new_[40898]_ ,
    \new_[40901]_ , \new_[40904]_ , \new_[40905]_ , \new_[40908]_ ,
    \new_[40911]_ , \new_[40912]_ , \new_[40913]_ , \new_[40916]_ ,
    \new_[40919]_ , \new_[40920]_ , \new_[40923]_ , \new_[40926]_ ,
    \new_[40927]_ , \new_[40928]_ , \new_[40931]_ , \new_[40934]_ ,
    \new_[40935]_ , \new_[40938]_ , \new_[40941]_ , \new_[40942]_ ,
    \new_[40943]_ , \new_[40946]_ , \new_[40949]_ , \new_[40950]_ ,
    \new_[40953]_ , \new_[40956]_ , \new_[40957]_ , \new_[40958]_ ,
    \new_[40961]_ , \new_[40964]_ , \new_[40965]_ , \new_[40968]_ ,
    \new_[40971]_ , \new_[40972]_ , \new_[40973]_ , \new_[40976]_ ,
    \new_[40979]_ , \new_[40980]_ , \new_[40983]_ , \new_[40986]_ ,
    \new_[40987]_ , \new_[40988]_ , \new_[40991]_ , \new_[40994]_ ,
    \new_[40995]_ , \new_[40998]_ , \new_[41001]_ , \new_[41002]_ ,
    \new_[41003]_ , \new_[41006]_ , \new_[41009]_ , \new_[41010]_ ,
    \new_[41013]_ , \new_[41016]_ , \new_[41017]_ , \new_[41018]_ ,
    \new_[41021]_ , \new_[41024]_ , \new_[41025]_ , \new_[41028]_ ,
    \new_[41031]_ , \new_[41032]_ , \new_[41033]_ , \new_[41036]_ ,
    \new_[41039]_ , \new_[41040]_ , \new_[41043]_ , \new_[41046]_ ,
    \new_[41047]_ , \new_[41048]_ , \new_[41051]_ , \new_[41054]_ ,
    \new_[41055]_ , \new_[41058]_ , \new_[41061]_ , \new_[41062]_ ,
    \new_[41063]_ , \new_[41066]_ , \new_[41069]_ , \new_[41070]_ ,
    \new_[41073]_ , \new_[41076]_ , \new_[41077]_ , \new_[41078]_ ,
    \new_[41081]_ , \new_[41084]_ , \new_[41085]_ , \new_[41088]_ ,
    \new_[41091]_ , \new_[41092]_ , \new_[41093]_ , \new_[41096]_ ,
    \new_[41099]_ , \new_[41100]_ , \new_[41103]_ , \new_[41106]_ ,
    \new_[41107]_ , \new_[41108]_ , \new_[41111]_ , \new_[41114]_ ,
    \new_[41115]_ , \new_[41118]_ , \new_[41121]_ , \new_[41122]_ ,
    \new_[41123]_ , \new_[41126]_ , \new_[41129]_ , \new_[41130]_ ,
    \new_[41133]_ , \new_[41136]_ , \new_[41137]_ , \new_[41138]_ ,
    \new_[41141]_ , \new_[41144]_ , \new_[41145]_ , \new_[41148]_ ,
    \new_[41151]_ , \new_[41152]_ , \new_[41153]_ , \new_[41156]_ ,
    \new_[41159]_ , \new_[41160]_ , \new_[41163]_ , \new_[41166]_ ,
    \new_[41167]_ , \new_[41168]_ , \new_[41171]_ , \new_[41174]_ ,
    \new_[41175]_ , \new_[41178]_ , \new_[41181]_ , \new_[41182]_ ,
    \new_[41183]_ , \new_[41186]_ , \new_[41189]_ , \new_[41190]_ ,
    \new_[41193]_ , \new_[41196]_ , \new_[41197]_ , \new_[41198]_ ,
    \new_[41201]_ , \new_[41204]_ , \new_[41205]_ , \new_[41208]_ ,
    \new_[41211]_ , \new_[41212]_ , \new_[41213]_ , \new_[41216]_ ,
    \new_[41219]_ , \new_[41220]_ , \new_[41223]_ , \new_[41226]_ ,
    \new_[41227]_ , \new_[41228]_ , \new_[41231]_ , \new_[41234]_ ,
    \new_[41235]_ , \new_[41238]_ , \new_[41241]_ , \new_[41242]_ ,
    \new_[41243]_ , \new_[41246]_ , \new_[41249]_ , \new_[41250]_ ,
    \new_[41253]_ , \new_[41256]_ , \new_[41257]_ , \new_[41258]_ ,
    \new_[41261]_ , \new_[41264]_ , \new_[41265]_ , \new_[41268]_ ,
    \new_[41271]_ , \new_[41272]_ , \new_[41273]_ , \new_[41276]_ ,
    \new_[41279]_ , \new_[41280]_ , \new_[41283]_ , \new_[41286]_ ,
    \new_[41287]_ , \new_[41288]_ , \new_[41291]_ , \new_[41294]_ ,
    \new_[41295]_ , \new_[41298]_ , \new_[41301]_ , \new_[41302]_ ,
    \new_[41303]_ , \new_[41306]_ , \new_[41309]_ , \new_[41310]_ ,
    \new_[41313]_ , \new_[41316]_ , \new_[41317]_ , \new_[41318]_ ,
    \new_[41321]_ , \new_[41324]_ , \new_[41325]_ , \new_[41328]_ ,
    \new_[41331]_ , \new_[41332]_ , \new_[41333]_ , \new_[41336]_ ,
    \new_[41339]_ , \new_[41340]_ , \new_[41343]_ , \new_[41346]_ ,
    \new_[41347]_ , \new_[41348]_ , \new_[41351]_ , \new_[41354]_ ,
    \new_[41355]_ , \new_[41358]_ , \new_[41361]_ , \new_[41362]_ ,
    \new_[41363]_ , \new_[41366]_ , \new_[41369]_ , \new_[41370]_ ,
    \new_[41373]_ , \new_[41376]_ , \new_[41377]_ , \new_[41378]_ ,
    \new_[41381]_ , \new_[41384]_ , \new_[41385]_ , \new_[41388]_ ,
    \new_[41391]_ , \new_[41392]_ , \new_[41393]_ , \new_[41396]_ ,
    \new_[41399]_ , \new_[41400]_ , \new_[41403]_ , \new_[41406]_ ,
    \new_[41407]_ , \new_[41408]_ , \new_[41411]_ , \new_[41414]_ ,
    \new_[41415]_ , \new_[41418]_ , \new_[41421]_ , \new_[41422]_ ,
    \new_[41423]_ , \new_[41426]_ , \new_[41429]_ , \new_[41430]_ ,
    \new_[41433]_ , \new_[41436]_ , \new_[41437]_ , \new_[41438]_ ,
    \new_[41441]_ , \new_[41444]_ , \new_[41445]_ , \new_[41448]_ ,
    \new_[41451]_ , \new_[41452]_ , \new_[41453]_ , \new_[41456]_ ,
    \new_[41459]_ , \new_[41460]_ , \new_[41463]_ , \new_[41466]_ ,
    \new_[41467]_ , \new_[41468]_ , \new_[41471]_ , \new_[41474]_ ,
    \new_[41475]_ , \new_[41478]_ , \new_[41481]_ , \new_[41482]_ ,
    \new_[41483]_ , \new_[41486]_ , \new_[41489]_ , \new_[41490]_ ,
    \new_[41493]_ , \new_[41496]_ , \new_[41497]_ , \new_[41498]_ ,
    \new_[41501]_ , \new_[41504]_ , \new_[41505]_ , \new_[41508]_ ,
    \new_[41511]_ , \new_[41512]_ , \new_[41513]_ , \new_[41516]_ ,
    \new_[41519]_ , \new_[41520]_ , \new_[41523]_ , \new_[41526]_ ,
    \new_[41527]_ , \new_[41528]_ , \new_[41531]_ , \new_[41534]_ ,
    \new_[41535]_ , \new_[41538]_ , \new_[41541]_ , \new_[41542]_ ,
    \new_[41543]_ , \new_[41546]_ , \new_[41549]_ , \new_[41550]_ ,
    \new_[41553]_ , \new_[41556]_ , \new_[41557]_ , \new_[41558]_ ,
    \new_[41561]_ , \new_[41564]_ , \new_[41565]_ , \new_[41568]_ ,
    \new_[41571]_ , \new_[41572]_ , \new_[41573]_ , \new_[41576]_ ,
    \new_[41579]_ , \new_[41580]_ , \new_[41583]_ , \new_[41586]_ ,
    \new_[41587]_ , \new_[41588]_ , \new_[41591]_ , \new_[41594]_ ,
    \new_[41595]_ , \new_[41598]_ , \new_[41601]_ , \new_[41602]_ ,
    \new_[41603]_ , \new_[41606]_ , \new_[41609]_ , \new_[41610]_ ,
    \new_[41613]_ , \new_[41616]_ , \new_[41617]_ , \new_[41618]_ ,
    \new_[41621]_ , \new_[41624]_ , \new_[41625]_ , \new_[41628]_ ,
    \new_[41631]_ , \new_[41632]_ , \new_[41633]_ , \new_[41636]_ ,
    \new_[41639]_ , \new_[41640]_ , \new_[41643]_ , \new_[41646]_ ,
    \new_[41647]_ , \new_[41648]_ , \new_[41651]_ , \new_[41654]_ ,
    \new_[41655]_ , \new_[41658]_ , \new_[41661]_ , \new_[41662]_ ,
    \new_[41663]_ , \new_[41666]_ , \new_[41669]_ , \new_[41670]_ ,
    \new_[41673]_ , \new_[41676]_ , \new_[41677]_ , \new_[41678]_ ,
    \new_[41681]_ , \new_[41684]_ , \new_[41685]_ , \new_[41688]_ ,
    \new_[41691]_ , \new_[41692]_ , \new_[41693]_ , \new_[41696]_ ,
    \new_[41699]_ , \new_[41700]_ , \new_[41703]_ , \new_[41706]_ ,
    \new_[41707]_ , \new_[41708]_ , \new_[41711]_ , \new_[41714]_ ,
    \new_[41715]_ , \new_[41718]_ , \new_[41721]_ , \new_[41722]_ ,
    \new_[41723]_ , \new_[41726]_ , \new_[41729]_ , \new_[41730]_ ,
    \new_[41733]_ , \new_[41736]_ , \new_[41737]_ , \new_[41738]_ ,
    \new_[41741]_ , \new_[41744]_ , \new_[41745]_ , \new_[41748]_ ,
    \new_[41751]_ , \new_[41752]_ , \new_[41753]_ , \new_[41756]_ ,
    \new_[41759]_ , \new_[41760]_ , \new_[41763]_ , \new_[41766]_ ,
    \new_[41767]_ , \new_[41768]_ , \new_[41771]_ , \new_[41774]_ ,
    \new_[41775]_ , \new_[41778]_ , \new_[41781]_ , \new_[41782]_ ,
    \new_[41783]_ , \new_[41786]_ , \new_[41789]_ , \new_[41790]_ ,
    \new_[41793]_ , \new_[41796]_ , \new_[41797]_ , \new_[41798]_ ,
    \new_[41801]_ , \new_[41804]_ , \new_[41805]_ , \new_[41808]_ ,
    \new_[41811]_ , \new_[41812]_ , \new_[41813]_ , \new_[41816]_ ,
    \new_[41819]_ , \new_[41820]_ , \new_[41823]_ , \new_[41826]_ ,
    \new_[41827]_ , \new_[41828]_ , \new_[41831]_ , \new_[41834]_ ,
    \new_[41835]_ , \new_[41838]_ , \new_[41841]_ , \new_[41842]_ ,
    \new_[41843]_ , \new_[41846]_ , \new_[41849]_ , \new_[41850]_ ,
    \new_[41853]_ , \new_[41856]_ , \new_[41857]_ , \new_[41858]_ ,
    \new_[41861]_ , \new_[41864]_ , \new_[41865]_ , \new_[41868]_ ,
    \new_[41871]_ , \new_[41872]_ , \new_[41873]_ , \new_[41876]_ ,
    \new_[41879]_ , \new_[41880]_ , \new_[41883]_ , \new_[41886]_ ,
    \new_[41887]_ , \new_[41888]_ , \new_[41891]_ , \new_[41894]_ ,
    \new_[41895]_ , \new_[41898]_ , \new_[41901]_ , \new_[41902]_ ,
    \new_[41903]_ , \new_[41906]_ , \new_[41909]_ , \new_[41910]_ ,
    \new_[41913]_ , \new_[41916]_ , \new_[41917]_ , \new_[41918]_ ,
    \new_[41921]_ , \new_[41924]_ , \new_[41925]_ , \new_[41928]_ ,
    \new_[41931]_ , \new_[41932]_ , \new_[41933]_ , \new_[41936]_ ,
    \new_[41939]_ , \new_[41940]_ , \new_[41943]_ , \new_[41946]_ ,
    \new_[41947]_ , \new_[41948]_ , \new_[41951]_ , \new_[41954]_ ,
    \new_[41955]_ , \new_[41958]_ , \new_[41961]_ , \new_[41962]_ ,
    \new_[41963]_ , \new_[41966]_ , \new_[41969]_ , \new_[41970]_ ,
    \new_[41973]_ , \new_[41976]_ , \new_[41977]_ , \new_[41978]_ ,
    \new_[41981]_ , \new_[41984]_ , \new_[41985]_ , \new_[41988]_ ,
    \new_[41991]_ , \new_[41992]_ , \new_[41993]_ , \new_[41996]_ ,
    \new_[41999]_ , \new_[42000]_ , \new_[42003]_ , \new_[42006]_ ,
    \new_[42007]_ , \new_[42008]_ , \new_[42011]_ , \new_[42014]_ ,
    \new_[42015]_ , \new_[42018]_ , \new_[42021]_ , \new_[42022]_ ,
    \new_[42023]_ , \new_[42026]_ , \new_[42029]_ , \new_[42030]_ ,
    \new_[42033]_ , \new_[42036]_ , \new_[42037]_ , \new_[42038]_ ,
    \new_[42041]_ , \new_[42044]_ , \new_[42045]_ , \new_[42048]_ ,
    \new_[42051]_ , \new_[42052]_ , \new_[42053]_ , \new_[42056]_ ,
    \new_[42059]_ , \new_[42060]_ , \new_[42063]_ , \new_[42066]_ ,
    \new_[42067]_ , \new_[42068]_ , \new_[42071]_ , \new_[42074]_ ,
    \new_[42075]_ , \new_[42078]_ , \new_[42081]_ , \new_[42082]_ ,
    \new_[42083]_ , \new_[42086]_ , \new_[42089]_ , \new_[42090]_ ,
    \new_[42093]_ , \new_[42096]_ , \new_[42097]_ , \new_[42098]_ ,
    \new_[42101]_ , \new_[42104]_ , \new_[42105]_ , \new_[42108]_ ,
    \new_[42111]_ , \new_[42112]_ , \new_[42113]_ , \new_[42116]_ ,
    \new_[42119]_ , \new_[42120]_ , \new_[42123]_ , \new_[42126]_ ,
    \new_[42127]_ , \new_[42128]_ , \new_[42131]_ , \new_[42134]_ ,
    \new_[42135]_ , \new_[42138]_ , \new_[42141]_ , \new_[42142]_ ,
    \new_[42143]_ , \new_[42146]_ , \new_[42149]_ , \new_[42150]_ ,
    \new_[42153]_ , \new_[42156]_ , \new_[42157]_ , \new_[42158]_ ,
    \new_[42161]_ , \new_[42164]_ , \new_[42165]_ , \new_[42168]_ ,
    \new_[42171]_ , \new_[42172]_ , \new_[42173]_ , \new_[42176]_ ,
    \new_[42179]_ , \new_[42180]_ , \new_[42183]_ , \new_[42186]_ ,
    \new_[42187]_ , \new_[42188]_ , \new_[42191]_ , \new_[42194]_ ,
    \new_[42195]_ , \new_[42198]_ , \new_[42201]_ , \new_[42202]_ ,
    \new_[42203]_ , \new_[42206]_ , \new_[42209]_ , \new_[42210]_ ,
    \new_[42213]_ , \new_[42216]_ , \new_[42217]_ , \new_[42218]_ ,
    \new_[42221]_ , \new_[42224]_ , \new_[42225]_ , \new_[42228]_ ,
    \new_[42231]_ , \new_[42232]_ , \new_[42233]_ , \new_[42236]_ ,
    \new_[42239]_ , \new_[42240]_ , \new_[42243]_ , \new_[42246]_ ,
    \new_[42247]_ , \new_[42248]_ , \new_[42251]_ , \new_[42254]_ ,
    \new_[42255]_ , \new_[42258]_ , \new_[42261]_ , \new_[42262]_ ,
    \new_[42263]_ , \new_[42266]_ , \new_[42269]_ , \new_[42270]_ ,
    \new_[42273]_ , \new_[42276]_ , \new_[42277]_ , \new_[42278]_ ,
    \new_[42281]_ , \new_[42284]_ , \new_[42285]_ , \new_[42288]_ ,
    \new_[42291]_ , \new_[42292]_ , \new_[42293]_ , \new_[42296]_ ,
    \new_[42299]_ , \new_[42300]_ , \new_[42303]_ , \new_[42306]_ ,
    \new_[42307]_ , \new_[42308]_ , \new_[42311]_ , \new_[42314]_ ,
    \new_[42315]_ , \new_[42318]_ , \new_[42321]_ , \new_[42322]_ ,
    \new_[42323]_ , \new_[42326]_ , \new_[42329]_ , \new_[42330]_ ,
    \new_[42333]_ , \new_[42336]_ , \new_[42337]_ , \new_[42338]_ ,
    \new_[42341]_ , \new_[42344]_ , \new_[42345]_ , \new_[42348]_ ,
    \new_[42351]_ , \new_[42352]_ , \new_[42353]_ , \new_[42356]_ ,
    \new_[42359]_ , \new_[42360]_ , \new_[42363]_ , \new_[42366]_ ,
    \new_[42367]_ , \new_[42368]_ , \new_[42371]_ , \new_[42374]_ ,
    \new_[42375]_ , \new_[42378]_ , \new_[42381]_ , \new_[42382]_ ,
    \new_[42383]_ , \new_[42386]_ , \new_[42389]_ , \new_[42390]_ ,
    \new_[42393]_ , \new_[42396]_ , \new_[42397]_ , \new_[42398]_ ,
    \new_[42401]_ , \new_[42404]_ , \new_[42405]_ , \new_[42408]_ ,
    \new_[42411]_ , \new_[42412]_ , \new_[42413]_ , \new_[42416]_ ,
    \new_[42419]_ , \new_[42420]_ , \new_[42423]_ , \new_[42426]_ ,
    \new_[42427]_ , \new_[42428]_ , \new_[42431]_ , \new_[42434]_ ,
    \new_[42435]_ , \new_[42438]_ , \new_[42441]_ , \new_[42442]_ ,
    \new_[42443]_ , \new_[42446]_ , \new_[42449]_ , \new_[42450]_ ,
    \new_[42453]_ , \new_[42456]_ , \new_[42457]_ , \new_[42458]_ ,
    \new_[42461]_ , \new_[42464]_ , \new_[42465]_ , \new_[42468]_ ,
    \new_[42471]_ , \new_[42472]_ , \new_[42473]_ , \new_[42476]_ ,
    \new_[42479]_ , \new_[42480]_ , \new_[42483]_ , \new_[42486]_ ,
    \new_[42487]_ , \new_[42488]_ , \new_[42491]_ , \new_[42494]_ ,
    \new_[42495]_ , \new_[42498]_ , \new_[42501]_ , \new_[42502]_ ,
    \new_[42503]_ , \new_[42506]_ , \new_[42509]_ , \new_[42510]_ ,
    \new_[42513]_ , \new_[42516]_ , \new_[42517]_ , \new_[42518]_ ,
    \new_[42521]_ , \new_[42524]_ , \new_[42525]_ , \new_[42528]_ ,
    \new_[42531]_ , \new_[42532]_ , \new_[42533]_ , \new_[42536]_ ,
    \new_[42539]_ , \new_[42540]_ , \new_[42543]_ , \new_[42546]_ ,
    \new_[42547]_ , \new_[42548]_ , \new_[42551]_ , \new_[42554]_ ,
    \new_[42555]_ , \new_[42558]_ , \new_[42561]_ , \new_[42562]_ ,
    \new_[42563]_ , \new_[42566]_ , \new_[42569]_ , \new_[42570]_ ,
    \new_[42573]_ , \new_[42576]_ , \new_[42577]_ , \new_[42578]_ ,
    \new_[42581]_ , \new_[42584]_ , \new_[42585]_ , \new_[42588]_ ,
    \new_[42591]_ , \new_[42592]_ , \new_[42593]_ , \new_[42596]_ ,
    \new_[42599]_ , \new_[42600]_ , \new_[42603]_ , \new_[42606]_ ,
    \new_[42607]_ , \new_[42608]_ , \new_[42611]_ , \new_[42614]_ ,
    \new_[42615]_ , \new_[42618]_ , \new_[42621]_ , \new_[42622]_ ,
    \new_[42623]_ , \new_[42626]_ , \new_[42629]_ , \new_[42630]_ ,
    \new_[42633]_ , \new_[42636]_ , \new_[42637]_ , \new_[42638]_ ,
    \new_[42641]_ , \new_[42644]_ , \new_[42645]_ , \new_[42648]_ ,
    \new_[42651]_ , \new_[42652]_ , \new_[42653]_ , \new_[42656]_ ,
    \new_[42659]_ , \new_[42660]_ , \new_[42663]_ , \new_[42666]_ ,
    \new_[42667]_ , \new_[42668]_ , \new_[42671]_ , \new_[42674]_ ,
    \new_[42675]_ , \new_[42678]_ , \new_[42681]_ , \new_[42682]_ ,
    \new_[42683]_ , \new_[42686]_ , \new_[42689]_ , \new_[42690]_ ,
    \new_[42693]_ , \new_[42696]_ , \new_[42697]_ , \new_[42698]_ ,
    \new_[42701]_ , \new_[42704]_ , \new_[42705]_ , \new_[42708]_ ,
    \new_[42711]_ , \new_[42712]_ , \new_[42713]_ , \new_[42716]_ ,
    \new_[42719]_ , \new_[42720]_ , \new_[42723]_ , \new_[42726]_ ,
    \new_[42727]_ , \new_[42728]_ , \new_[42731]_ , \new_[42734]_ ,
    \new_[42735]_ , \new_[42738]_ , \new_[42741]_ , \new_[42742]_ ,
    \new_[42743]_ , \new_[42746]_ , \new_[42749]_ , \new_[42750]_ ,
    \new_[42753]_ , \new_[42756]_ , \new_[42757]_ , \new_[42758]_ ,
    \new_[42761]_ , \new_[42764]_ , \new_[42765]_ , \new_[42768]_ ,
    \new_[42771]_ , \new_[42772]_ , \new_[42773]_ , \new_[42776]_ ,
    \new_[42779]_ , \new_[42780]_ , \new_[42783]_ , \new_[42786]_ ,
    \new_[42787]_ , \new_[42788]_ , \new_[42791]_ , \new_[42794]_ ,
    \new_[42795]_ , \new_[42798]_ , \new_[42801]_ , \new_[42802]_ ,
    \new_[42803]_ , \new_[42806]_ , \new_[42809]_ , \new_[42810]_ ,
    \new_[42813]_ , \new_[42816]_ , \new_[42817]_ , \new_[42818]_ ,
    \new_[42821]_ , \new_[42824]_ , \new_[42825]_ , \new_[42828]_ ,
    \new_[42831]_ , \new_[42832]_ , \new_[42833]_ , \new_[42836]_ ,
    \new_[42839]_ , \new_[42840]_ , \new_[42843]_ , \new_[42846]_ ,
    \new_[42847]_ , \new_[42848]_ , \new_[42851]_ , \new_[42854]_ ,
    \new_[42855]_ , \new_[42858]_ , \new_[42861]_ , \new_[42862]_ ,
    \new_[42863]_ , \new_[42866]_ , \new_[42869]_ , \new_[42870]_ ,
    \new_[42873]_ , \new_[42876]_ , \new_[42877]_ , \new_[42878]_ ,
    \new_[42881]_ , \new_[42884]_ , \new_[42885]_ , \new_[42888]_ ,
    \new_[42891]_ , \new_[42892]_ , \new_[42893]_ , \new_[42896]_ ,
    \new_[42899]_ , \new_[42900]_ , \new_[42903]_ , \new_[42906]_ ,
    \new_[42907]_ , \new_[42908]_ , \new_[42911]_ , \new_[42914]_ ,
    \new_[42915]_ , \new_[42918]_ , \new_[42921]_ , \new_[42922]_ ,
    \new_[42923]_ , \new_[42926]_ , \new_[42929]_ , \new_[42930]_ ,
    \new_[42933]_ , \new_[42936]_ , \new_[42937]_ , \new_[42938]_ ,
    \new_[42941]_ , \new_[42944]_ , \new_[42945]_ , \new_[42948]_ ,
    \new_[42951]_ , \new_[42952]_ , \new_[42953]_ , \new_[42956]_ ,
    \new_[42959]_ , \new_[42960]_ , \new_[42963]_ , \new_[42966]_ ,
    \new_[42967]_ , \new_[42968]_ , \new_[42971]_ , \new_[42974]_ ,
    \new_[42975]_ , \new_[42978]_ , \new_[42981]_ , \new_[42982]_ ,
    \new_[42983]_ , \new_[42986]_ , \new_[42989]_ , \new_[42990]_ ,
    \new_[42993]_ , \new_[42996]_ , \new_[42997]_ , \new_[42998]_ ,
    \new_[43001]_ , \new_[43004]_ , \new_[43005]_ , \new_[43008]_ ,
    \new_[43011]_ , \new_[43012]_ , \new_[43013]_ , \new_[43016]_ ,
    \new_[43019]_ , \new_[43020]_ , \new_[43023]_ , \new_[43026]_ ,
    \new_[43027]_ , \new_[43028]_ , \new_[43031]_ , \new_[43034]_ ,
    \new_[43035]_ , \new_[43038]_ , \new_[43041]_ , \new_[43042]_ ,
    \new_[43043]_ , \new_[43046]_ , \new_[43049]_ , \new_[43050]_ ,
    \new_[43053]_ , \new_[43056]_ , \new_[43057]_ , \new_[43058]_ ,
    \new_[43061]_ , \new_[43064]_ , \new_[43065]_ , \new_[43068]_ ,
    \new_[43071]_ , \new_[43072]_ , \new_[43073]_ , \new_[43076]_ ,
    \new_[43079]_ , \new_[43080]_ , \new_[43083]_ , \new_[43086]_ ,
    \new_[43087]_ , \new_[43088]_ , \new_[43091]_ , \new_[43094]_ ,
    \new_[43095]_ , \new_[43098]_ , \new_[43101]_ , \new_[43102]_ ,
    \new_[43103]_ , \new_[43106]_ , \new_[43109]_ , \new_[43110]_ ,
    \new_[43113]_ , \new_[43116]_ , \new_[43117]_ , \new_[43118]_ ,
    \new_[43121]_ , \new_[43124]_ , \new_[43125]_ , \new_[43128]_ ,
    \new_[43131]_ , \new_[43132]_ , \new_[43133]_ , \new_[43136]_ ,
    \new_[43139]_ , \new_[43140]_ , \new_[43143]_ , \new_[43146]_ ,
    \new_[43147]_ , \new_[43148]_ , \new_[43151]_ , \new_[43154]_ ,
    \new_[43155]_ , \new_[43158]_ , \new_[43161]_ , \new_[43162]_ ,
    \new_[43163]_ , \new_[43166]_ , \new_[43169]_ , \new_[43170]_ ,
    \new_[43173]_ , \new_[43176]_ , \new_[43177]_ , \new_[43178]_ ,
    \new_[43181]_ , \new_[43184]_ , \new_[43185]_ , \new_[43188]_ ,
    \new_[43191]_ , \new_[43192]_ , \new_[43193]_ , \new_[43196]_ ,
    \new_[43199]_ , \new_[43200]_ , \new_[43203]_ , \new_[43206]_ ,
    \new_[43207]_ , \new_[43208]_ , \new_[43211]_ , \new_[43214]_ ,
    \new_[43215]_ , \new_[43218]_ , \new_[43221]_ , \new_[43222]_ ,
    \new_[43223]_ , \new_[43226]_ , \new_[43229]_ , \new_[43230]_ ,
    \new_[43233]_ , \new_[43236]_ , \new_[43237]_ , \new_[43238]_ ,
    \new_[43241]_ , \new_[43244]_ , \new_[43245]_ , \new_[43248]_ ,
    \new_[43251]_ , \new_[43252]_ , \new_[43253]_ , \new_[43256]_ ,
    \new_[43259]_ , \new_[43260]_ , \new_[43263]_ , \new_[43266]_ ,
    \new_[43267]_ , \new_[43268]_ , \new_[43271]_ , \new_[43274]_ ,
    \new_[43275]_ , \new_[43278]_ , \new_[43281]_ , \new_[43282]_ ,
    \new_[43283]_ , \new_[43286]_ , \new_[43289]_ , \new_[43290]_ ,
    \new_[43293]_ , \new_[43296]_ , \new_[43297]_ , \new_[43298]_ ,
    \new_[43301]_ , \new_[43304]_ , \new_[43305]_ , \new_[43308]_ ,
    \new_[43311]_ , \new_[43312]_ , \new_[43313]_ , \new_[43316]_ ,
    \new_[43319]_ , \new_[43320]_ , \new_[43323]_ , \new_[43326]_ ,
    \new_[43327]_ , \new_[43328]_ , \new_[43331]_ , \new_[43334]_ ,
    \new_[43335]_ , \new_[43338]_ , \new_[43341]_ , \new_[43342]_ ,
    \new_[43343]_ , \new_[43346]_ , \new_[43349]_ , \new_[43350]_ ,
    \new_[43353]_ , \new_[43356]_ , \new_[43357]_ , \new_[43358]_ ,
    \new_[43361]_ , \new_[43364]_ , \new_[43365]_ , \new_[43368]_ ,
    \new_[43371]_ , \new_[43372]_ , \new_[43373]_ , \new_[43376]_ ,
    \new_[43379]_ , \new_[43380]_ , \new_[43383]_ , \new_[43386]_ ,
    \new_[43387]_ , \new_[43388]_ , \new_[43391]_ , \new_[43394]_ ,
    \new_[43395]_ , \new_[43398]_ , \new_[43401]_ , \new_[43402]_ ,
    \new_[43403]_ , \new_[43406]_ , \new_[43409]_ , \new_[43410]_ ,
    \new_[43413]_ , \new_[43416]_ , \new_[43417]_ , \new_[43418]_ ,
    \new_[43421]_ , \new_[43424]_ , \new_[43425]_ , \new_[43428]_ ,
    \new_[43431]_ , \new_[43432]_ , \new_[43433]_ , \new_[43436]_ ,
    \new_[43439]_ , \new_[43440]_ , \new_[43443]_ , \new_[43446]_ ,
    \new_[43447]_ , \new_[43448]_ , \new_[43451]_ , \new_[43454]_ ,
    \new_[43455]_ , \new_[43458]_ , \new_[43461]_ , \new_[43462]_ ,
    \new_[43463]_ , \new_[43466]_ , \new_[43469]_ , \new_[43470]_ ,
    \new_[43473]_ , \new_[43476]_ , \new_[43477]_ , \new_[43478]_ ,
    \new_[43481]_ , \new_[43484]_ , \new_[43485]_ , \new_[43488]_ ,
    \new_[43491]_ , \new_[43492]_ , \new_[43493]_ , \new_[43496]_ ,
    \new_[43499]_ , \new_[43500]_ , \new_[43503]_ , \new_[43506]_ ,
    \new_[43507]_ , \new_[43508]_ , \new_[43511]_ , \new_[43514]_ ,
    \new_[43515]_ , \new_[43518]_ , \new_[43521]_ , \new_[43522]_ ,
    \new_[43523]_ , \new_[43526]_ , \new_[43529]_ , \new_[43530]_ ,
    \new_[43533]_ , \new_[43536]_ , \new_[43537]_ , \new_[43538]_ ,
    \new_[43541]_ , \new_[43544]_ , \new_[43545]_ , \new_[43548]_ ,
    \new_[43551]_ , \new_[43552]_ , \new_[43553]_ , \new_[43556]_ ,
    \new_[43559]_ , \new_[43560]_ , \new_[43563]_ , \new_[43566]_ ,
    \new_[43567]_ , \new_[43568]_ , \new_[43571]_ , \new_[43574]_ ,
    \new_[43575]_ , \new_[43578]_ , \new_[43581]_ , \new_[43582]_ ,
    \new_[43583]_ , \new_[43586]_ , \new_[43589]_ , \new_[43590]_ ,
    \new_[43593]_ , \new_[43596]_ , \new_[43597]_ , \new_[43598]_ ,
    \new_[43601]_ , \new_[43604]_ , \new_[43605]_ , \new_[43608]_ ,
    \new_[43611]_ , \new_[43612]_ , \new_[43613]_ , \new_[43616]_ ,
    \new_[43619]_ , \new_[43620]_ , \new_[43623]_ , \new_[43626]_ ,
    \new_[43627]_ , \new_[43628]_ , \new_[43631]_ , \new_[43634]_ ,
    \new_[43635]_ , \new_[43638]_ , \new_[43641]_ , \new_[43642]_ ,
    \new_[43643]_ , \new_[43646]_ , \new_[43649]_ , \new_[43650]_ ,
    \new_[43653]_ , \new_[43656]_ , \new_[43657]_ , \new_[43658]_ ,
    \new_[43661]_ , \new_[43664]_ , \new_[43665]_ , \new_[43668]_ ,
    \new_[43671]_ , \new_[43672]_ , \new_[43673]_ , \new_[43676]_ ,
    \new_[43679]_ , \new_[43680]_ , \new_[43683]_ , \new_[43686]_ ,
    \new_[43687]_ , \new_[43688]_ , \new_[43691]_ , \new_[43694]_ ,
    \new_[43695]_ , \new_[43698]_ , \new_[43701]_ , \new_[43702]_ ,
    \new_[43703]_ , \new_[43706]_ , \new_[43709]_ , \new_[43710]_ ,
    \new_[43713]_ , \new_[43716]_ , \new_[43717]_ , \new_[43718]_ ,
    \new_[43721]_ , \new_[43724]_ , \new_[43725]_ , \new_[43728]_ ,
    \new_[43731]_ , \new_[43732]_ , \new_[43733]_ , \new_[43736]_ ,
    \new_[43739]_ , \new_[43740]_ , \new_[43743]_ , \new_[43746]_ ,
    \new_[43747]_ , \new_[43748]_ , \new_[43751]_ , \new_[43754]_ ,
    \new_[43755]_ , \new_[43758]_ , \new_[43761]_ , \new_[43762]_ ,
    \new_[43763]_ , \new_[43766]_ , \new_[43769]_ , \new_[43770]_ ,
    \new_[43773]_ , \new_[43776]_ , \new_[43777]_ , \new_[43778]_ ,
    \new_[43781]_ , \new_[43784]_ , \new_[43785]_ , \new_[43788]_ ,
    \new_[43791]_ , \new_[43792]_ , \new_[43793]_ , \new_[43796]_ ,
    \new_[43799]_ , \new_[43800]_ , \new_[43803]_ , \new_[43806]_ ,
    \new_[43807]_ , \new_[43808]_ , \new_[43811]_ , \new_[43814]_ ,
    \new_[43815]_ , \new_[43818]_ , \new_[43821]_ , \new_[43822]_ ,
    \new_[43823]_ , \new_[43826]_ , \new_[43829]_ , \new_[43830]_ ,
    \new_[43833]_ , \new_[43836]_ , \new_[43837]_ , \new_[43838]_ ,
    \new_[43841]_ , \new_[43844]_ , \new_[43845]_ , \new_[43848]_ ,
    \new_[43851]_ , \new_[43852]_ , \new_[43853]_ , \new_[43856]_ ,
    \new_[43859]_ , \new_[43860]_ , \new_[43863]_ , \new_[43866]_ ,
    \new_[43867]_ , \new_[43868]_ , \new_[43871]_ , \new_[43874]_ ,
    \new_[43875]_ , \new_[43878]_ , \new_[43881]_ , \new_[43882]_ ,
    \new_[43883]_ , \new_[43886]_ , \new_[43889]_ , \new_[43890]_ ,
    \new_[43893]_ , \new_[43896]_ , \new_[43897]_ , \new_[43898]_ ,
    \new_[43901]_ , \new_[43904]_ , \new_[43905]_ , \new_[43908]_ ,
    \new_[43911]_ , \new_[43912]_ , \new_[43913]_ , \new_[43916]_ ,
    \new_[43919]_ , \new_[43920]_ , \new_[43923]_ , \new_[43926]_ ,
    \new_[43927]_ , \new_[43928]_ , \new_[43931]_ , \new_[43934]_ ,
    \new_[43935]_ , \new_[43938]_ , \new_[43941]_ , \new_[43942]_ ,
    \new_[43943]_ , \new_[43946]_ , \new_[43949]_ , \new_[43950]_ ,
    \new_[43953]_ , \new_[43956]_ , \new_[43957]_ , \new_[43958]_ ,
    \new_[43961]_ , \new_[43964]_ , \new_[43965]_ , \new_[43968]_ ,
    \new_[43971]_ , \new_[43972]_ , \new_[43973]_ , \new_[43976]_ ,
    \new_[43979]_ , \new_[43980]_ , \new_[43983]_ , \new_[43986]_ ,
    \new_[43987]_ , \new_[43988]_ , \new_[43991]_ , \new_[43994]_ ,
    \new_[43995]_ , \new_[43998]_ , \new_[44001]_ , \new_[44002]_ ,
    \new_[44003]_ , \new_[44006]_ , \new_[44009]_ , \new_[44010]_ ,
    \new_[44013]_ , \new_[44016]_ , \new_[44017]_ , \new_[44018]_ ,
    \new_[44021]_ , \new_[44024]_ , \new_[44025]_ , \new_[44028]_ ,
    \new_[44031]_ , \new_[44032]_ , \new_[44033]_ , \new_[44036]_ ,
    \new_[44039]_ , \new_[44040]_ , \new_[44043]_ , \new_[44046]_ ,
    \new_[44047]_ , \new_[44048]_ , \new_[44051]_ , \new_[44054]_ ,
    \new_[44055]_ , \new_[44058]_ , \new_[44061]_ , \new_[44062]_ ,
    \new_[44063]_ , \new_[44066]_ , \new_[44069]_ , \new_[44070]_ ,
    \new_[44073]_ , \new_[44076]_ , \new_[44077]_ , \new_[44078]_ ,
    \new_[44081]_ , \new_[44084]_ , \new_[44085]_ , \new_[44088]_ ,
    \new_[44091]_ , \new_[44092]_ , \new_[44093]_ , \new_[44096]_ ,
    \new_[44099]_ , \new_[44100]_ , \new_[44103]_ , \new_[44106]_ ,
    \new_[44107]_ , \new_[44108]_ , \new_[44111]_ , \new_[44114]_ ,
    \new_[44115]_ , \new_[44118]_ , \new_[44121]_ , \new_[44122]_ ,
    \new_[44123]_ , \new_[44126]_ , \new_[44129]_ , \new_[44130]_ ,
    \new_[44133]_ , \new_[44136]_ , \new_[44137]_ , \new_[44138]_ ,
    \new_[44141]_ , \new_[44144]_ , \new_[44145]_ , \new_[44148]_ ,
    \new_[44151]_ , \new_[44152]_ , \new_[44153]_ , \new_[44156]_ ,
    \new_[44159]_ , \new_[44160]_ , \new_[44163]_ , \new_[44166]_ ,
    \new_[44167]_ , \new_[44168]_ , \new_[44171]_ , \new_[44174]_ ,
    \new_[44175]_ , \new_[44178]_ , \new_[44181]_ , \new_[44182]_ ,
    \new_[44183]_ , \new_[44186]_ , \new_[44189]_ , \new_[44190]_ ,
    \new_[44193]_ , \new_[44196]_ , \new_[44197]_ , \new_[44198]_ ,
    \new_[44201]_ , \new_[44204]_ , \new_[44205]_ , \new_[44208]_ ,
    \new_[44211]_ , \new_[44212]_ , \new_[44213]_ , \new_[44216]_ ,
    \new_[44219]_ , \new_[44220]_ , \new_[44223]_ , \new_[44226]_ ,
    \new_[44227]_ , \new_[44228]_ , \new_[44231]_ , \new_[44234]_ ,
    \new_[44235]_ , \new_[44238]_ , \new_[44241]_ , \new_[44242]_ ,
    \new_[44243]_ , \new_[44246]_ , \new_[44249]_ , \new_[44250]_ ,
    \new_[44253]_ , \new_[44256]_ , \new_[44257]_ , \new_[44258]_ ,
    \new_[44261]_ , \new_[44264]_ , \new_[44265]_ , \new_[44268]_ ,
    \new_[44271]_ , \new_[44272]_ , \new_[44273]_ , \new_[44276]_ ,
    \new_[44279]_ , \new_[44280]_ , \new_[44283]_ , \new_[44286]_ ,
    \new_[44287]_ , \new_[44288]_ , \new_[44291]_ , \new_[44294]_ ,
    \new_[44295]_ , \new_[44298]_ , \new_[44301]_ , \new_[44302]_ ,
    \new_[44303]_ , \new_[44306]_ , \new_[44309]_ , \new_[44310]_ ,
    \new_[44313]_ , \new_[44316]_ , \new_[44317]_ , \new_[44318]_ ,
    \new_[44321]_ , \new_[44324]_ , \new_[44325]_ , \new_[44328]_ ,
    \new_[44331]_ , \new_[44332]_ , \new_[44333]_ , \new_[44336]_ ,
    \new_[44339]_ , \new_[44340]_ , \new_[44343]_ , \new_[44346]_ ,
    \new_[44347]_ , \new_[44348]_ , \new_[44351]_ , \new_[44354]_ ,
    \new_[44355]_ , \new_[44358]_ , \new_[44361]_ , \new_[44362]_ ,
    \new_[44363]_ , \new_[44366]_ , \new_[44369]_ , \new_[44370]_ ,
    \new_[44373]_ , \new_[44376]_ , \new_[44377]_ , \new_[44378]_ ,
    \new_[44381]_ , \new_[44384]_ , \new_[44385]_ , \new_[44388]_ ,
    \new_[44391]_ , \new_[44392]_ , \new_[44393]_ , \new_[44396]_ ,
    \new_[44399]_ , \new_[44400]_ , \new_[44403]_ , \new_[44406]_ ,
    \new_[44407]_ , \new_[44408]_ , \new_[44411]_ , \new_[44414]_ ,
    \new_[44415]_ , \new_[44418]_ , \new_[44421]_ , \new_[44422]_ ,
    \new_[44423]_ , \new_[44426]_ , \new_[44429]_ , \new_[44430]_ ,
    \new_[44433]_ , \new_[44436]_ , \new_[44437]_ , \new_[44438]_ ,
    \new_[44441]_ , \new_[44444]_ , \new_[44445]_ , \new_[44448]_ ,
    \new_[44451]_ , \new_[44452]_ , \new_[44453]_ , \new_[44456]_ ,
    \new_[44459]_ , \new_[44460]_ , \new_[44463]_ , \new_[44466]_ ,
    \new_[44467]_ , \new_[44468]_ , \new_[44471]_ , \new_[44474]_ ,
    \new_[44475]_ , \new_[44478]_ , \new_[44481]_ , \new_[44482]_ ,
    \new_[44483]_ , \new_[44486]_ , \new_[44489]_ , \new_[44490]_ ,
    \new_[44493]_ , \new_[44496]_ , \new_[44497]_ , \new_[44498]_ ,
    \new_[44501]_ , \new_[44504]_ , \new_[44505]_ , \new_[44508]_ ,
    \new_[44511]_ , \new_[44512]_ , \new_[44513]_ , \new_[44516]_ ,
    \new_[44519]_ , \new_[44520]_ , \new_[44523]_ , \new_[44526]_ ,
    \new_[44527]_ , \new_[44528]_ , \new_[44531]_ , \new_[44534]_ ,
    \new_[44535]_ , \new_[44538]_ , \new_[44541]_ , \new_[44542]_ ,
    \new_[44543]_ , \new_[44546]_ , \new_[44549]_ , \new_[44550]_ ,
    \new_[44553]_ , \new_[44556]_ , \new_[44557]_ , \new_[44558]_ ,
    \new_[44561]_ , \new_[44564]_ , \new_[44565]_ , \new_[44568]_ ,
    \new_[44571]_ , \new_[44572]_ , \new_[44573]_ , \new_[44576]_ ,
    \new_[44579]_ , \new_[44580]_ , \new_[44583]_ , \new_[44586]_ ,
    \new_[44587]_ , \new_[44588]_ , \new_[44591]_ , \new_[44594]_ ,
    \new_[44595]_ , \new_[44598]_ , \new_[44601]_ , \new_[44602]_ ,
    \new_[44603]_ , \new_[44606]_ , \new_[44609]_ , \new_[44610]_ ,
    \new_[44613]_ , \new_[44616]_ , \new_[44617]_ , \new_[44618]_ ,
    \new_[44621]_ , \new_[44624]_ , \new_[44625]_ , \new_[44628]_ ,
    \new_[44631]_ , \new_[44632]_ , \new_[44633]_ , \new_[44636]_ ,
    \new_[44639]_ , \new_[44640]_ , \new_[44643]_ , \new_[44646]_ ,
    \new_[44647]_ , \new_[44648]_ , \new_[44651]_ , \new_[44654]_ ,
    \new_[44655]_ , \new_[44658]_ , \new_[44661]_ , \new_[44662]_ ,
    \new_[44663]_ , \new_[44666]_ , \new_[44669]_ , \new_[44670]_ ,
    \new_[44673]_ , \new_[44676]_ , \new_[44677]_ , \new_[44678]_ ,
    \new_[44681]_ , \new_[44684]_ , \new_[44685]_ , \new_[44688]_ ,
    \new_[44691]_ , \new_[44692]_ , \new_[44693]_ , \new_[44696]_ ,
    \new_[44699]_ , \new_[44700]_ , \new_[44703]_ , \new_[44706]_ ,
    \new_[44707]_ , \new_[44708]_ , \new_[44711]_ , \new_[44714]_ ,
    \new_[44715]_ , \new_[44718]_ , \new_[44721]_ , \new_[44722]_ ,
    \new_[44723]_ , \new_[44726]_ , \new_[44729]_ , \new_[44730]_ ,
    \new_[44733]_ , \new_[44736]_ , \new_[44737]_ , \new_[44738]_ ,
    \new_[44741]_ , \new_[44744]_ , \new_[44745]_ , \new_[44748]_ ,
    \new_[44751]_ , \new_[44752]_ , \new_[44753]_ , \new_[44756]_ ,
    \new_[44759]_ , \new_[44760]_ , \new_[44763]_ , \new_[44766]_ ,
    \new_[44767]_ , \new_[44768]_ , \new_[44771]_ , \new_[44774]_ ,
    \new_[44775]_ , \new_[44778]_ , \new_[44781]_ , \new_[44782]_ ,
    \new_[44783]_ , \new_[44786]_ , \new_[44789]_ , \new_[44790]_ ,
    \new_[44793]_ , \new_[44796]_ , \new_[44797]_ , \new_[44798]_ ,
    \new_[44801]_ , \new_[44804]_ , \new_[44805]_ , \new_[44808]_ ,
    \new_[44811]_ , \new_[44812]_ , \new_[44813]_ , \new_[44816]_ ,
    \new_[44819]_ , \new_[44820]_ , \new_[44823]_ , \new_[44826]_ ,
    \new_[44827]_ , \new_[44828]_ , \new_[44831]_ , \new_[44834]_ ,
    \new_[44835]_ , \new_[44838]_ , \new_[44841]_ , \new_[44842]_ ,
    \new_[44843]_ , \new_[44846]_ , \new_[44849]_ , \new_[44850]_ ,
    \new_[44853]_ , \new_[44856]_ , \new_[44857]_ , \new_[44858]_ ,
    \new_[44861]_ , \new_[44864]_ , \new_[44865]_ , \new_[44868]_ ,
    \new_[44871]_ , \new_[44872]_ , \new_[44873]_ , \new_[44876]_ ,
    \new_[44879]_ , \new_[44880]_ , \new_[44883]_ , \new_[44886]_ ,
    \new_[44887]_ , \new_[44888]_ , \new_[44891]_ , \new_[44894]_ ,
    \new_[44895]_ , \new_[44898]_ , \new_[44901]_ , \new_[44902]_ ,
    \new_[44903]_ , \new_[44906]_ , \new_[44909]_ , \new_[44910]_ ,
    \new_[44913]_ , \new_[44916]_ , \new_[44917]_ , \new_[44918]_ ,
    \new_[44921]_ , \new_[44924]_ , \new_[44925]_ , \new_[44928]_ ,
    \new_[44931]_ , \new_[44932]_ , \new_[44933]_ , \new_[44936]_ ,
    \new_[44939]_ , \new_[44940]_ , \new_[44943]_ , \new_[44946]_ ,
    \new_[44947]_ , \new_[44948]_ , \new_[44951]_ , \new_[44954]_ ,
    \new_[44955]_ , \new_[44958]_ , \new_[44961]_ , \new_[44962]_ ,
    \new_[44963]_ , \new_[44966]_ , \new_[44969]_ , \new_[44970]_ ,
    \new_[44973]_ , \new_[44976]_ , \new_[44977]_ , \new_[44978]_ ,
    \new_[44981]_ , \new_[44984]_ , \new_[44985]_ , \new_[44988]_ ,
    \new_[44991]_ , \new_[44992]_ , \new_[44993]_ , \new_[44996]_ ,
    \new_[44999]_ , \new_[45000]_ , \new_[45003]_ , \new_[45006]_ ,
    \new_[45007]_ , \new_[45008]_ , \new_[45011]_ , \new_[45014]_ ,
    \new_[45015]_ , \new_[45018]_ , \new_[45021]_ , \new_[45022]_ ,
    \new_[45023]_ , \new_[45026]_ , \new_[45029]_ , \new_[45030]_ ,
    \new_[45033]_ , \new_[45036]_ , \new_[45037]_ , \new_[45038]_ ,
    \new_[45041]_ , \new_[45044]_ , \new_[45045]_ , \new_[45048]_ ,
    \new_[45051]_ , \new_[45052]_ , \new_[45053]_ , \new_[45056]_ ,
    \new_[45059]_ , \new_[45060]_ , \new_[45063]_ , \new_[45066]_ ,
    \new_[45067]_ , \new_[45068]_ , \new_[45071]_ , \new_[45074]_ ,
    \new_[45075]_ , \new_[45078]_ , \new_[45081]_ , \new_[45082]_ ,
    \new_[45083]_ , \new_[45086]_ , \new_[45089]_ , \new_[45090]_ ,
    \new_[45093]_ , \new_[45096]_ , \new_[45097]_ , \new_[45098]_ ,
    \new_[45101]_ , \new_[45104]_ , \new_[45105]_ , \new_[45108]_ ,
    \new_[45111]_ , \new_[45112]_ , \new_[45113]_ , \new_[45116]_ ,
    \new_[45119]_ , \new_[45120]_ , \new_[45123]_ , \new_[45126]_ ,
    \new_[45127]_ , \new_[45128]_ , \new_[45131]_ , \new_[45134]_ ,
    \new_[45135]_ , \new_[45138]_ , \new_[45141]_ , \new_[45142]_ ,
    \new_[45143]_ , \new_[45146]_ , \new_[45149]_ , \new_[45150]_ ,
    \new_[45153]_ , \new_[45156]_ , \new_[45157]_ , \new_[45158]_ ,
    \new_[45161]_ , \new_[45164]_ , \new_[45165]_ , \new_[45168]_ ,
    \new_[45171]_ , \new_[45172]_ , \new_[45173]_ , \new_[45176]_ ,
    \new_[45179]_ , \new_[45180]_ , \new_[45183]_ , \new_[45186]_ ,
    \new_[45187]_ , \new_[45188]_ , \new_[45191]_ , \new_[45194]_ ,
    \new_[45195]_ , \new_[45198]_ , \new_[45201]_ , \new_[45202]_ ,
    \new_[45203]_ , \new_[45206]_ , \new_[45209]_ , \new_[45210]_ ,
    \new_[45213]_ , \new_[45216]_ , \new_[45217]_ , \new_[45218]_ ,
    \new_[45221]_ , \new_[45224]_ , \new_[45225]_ , \new_[45228]_ ,
    \new_[45231]_ , \new_[45232]_ , \new_[45233]_ , \new_[45236]_ ,
    \new_[45239]_ , \new_[45240]_ , \new_[45243]_ , \new_[45246]_ ,
    \new_[45247]_ , \new_[45248]_ , \new_[45251]_ , \new_[45254]_ ,
    \new_[45255]_ , \new_[45258]_ , \new_[45261]_ , \new_[45262]_ ,
    \new_[45263]_ , \new_[45266]_ , \new_[45269]_ , \new_[45270]_ ,
    \new_[45273]_ , \new_[45276]_ , \new_[45277]_ , \new_[45278]_ ,
    \new_[45281]_ , \new_[45284]_ , \new_[45285]_ , \new_[45288]_ ,
    \new_[45291]_ , \new_[45292]_ , \new_[45293]_ , \new_[45296]_ ,
    \new_[45299]_ , \new_[45300]_ , \new_[45303]_ , \new_[45306]_ ,
    \new_[45307]_ , \new_[45308]_ , \new_[45311]_ , \new_[45314]_ ,
    \new_[45315]_ , \new_[45318]_ , \new_[45321]_ , \new_[45322]_ ,
    \new_[45323]_ , \new_[45326]_ , \new_[45329]_ , \new_[45330]_ ,
    \new_[45333]_ , \new_[45336]_ , \new_[45337]_ , \new_[45338]_ ,
    \new_[45341]_ , \new_[45344]_ , \new_[45345]_ , \new_[45348]_ ,
    \new_[45351]_ , \new_[45352]_ , \new_[45353]_ , \new_[45356]_ ,
    \new_[45359]_ , \new_[45360]_ , \new_[45363]_ , \new_[45366]_ ,
    \new_[45367]_ , \new_[45368]_ , \new_[45371]_ , \new_[45374]_ ,
    \new_[45375]_ , \new_[45378]_ , \new_[45381]_ , \new_[45382]_ ,
    \new_[45383]_ , \new_[45386]_ , \new_[45389]_ , \new_[45390]_ ,
    \new_[45393]_ , \new_[45396]_ , \new_[45397]_ , \new_[45398]_ ,
    \new_[45401]_ , \new_[45404]_ , \new_[45405]_ , \new_[45408]_ ,
    \new_[45411]_ , \new_[45412]_ , \new_[45413]_ , \new_[45416]_ ,
    \new_[45419]_ , \new_[45420]_ , \new_[45423]_ , \new_[45426]_ ,
    \new_[45427]_ , \new_[45428]_ , \new_[45431]_ , \new_[45434]_ ,
    \new_[45435]_ , \new_[45438]_ , \new_[45441]_ , \new_[45442]_ ,
    \new_[45443]_ , \new_[45446]_ , \new_[45449]_ , \new_[45450]_ ,
    \new_[45453]_ , \new_[45456]_ , \new_[45457]_ , \new_[45458]_ ,
    \new_[45461]_ , \new_[45464]_ , \new_[45465]_ , \new_[45468]_ ,
    \new_[45471]_ , \new_[45472]_ , \new_[45473]_ , \new_[45476]_ ,
    \new_[45479]_ , \new_[45480]_ , \new_[45483]_ , \new_[45486]_ ,
    \new_[45487]_ , \new_[45488]_ , \new_[45491]_ , \new_[45494]_ ,
    \new_[45495]_ , \new_[45498]_ , \new_[45501]_ , \new_[45502]_ ,
    \new_[45503]_ , \new_[45506]_ , \new_[45509]_ , \new_[45510]_ ,
    \new_[45513]_ , \new_[45516]_ , \new_[45517]_ , \new_[45518]_ ,
    \new_[45521]_ , \new_[45524]_ , \new_[45525]_ , \new_[45528]_ ,
    \new_[45531]_ , \new_[45532]_ , \new_[45533]_ , \new_[45536]_ ,
    \new_[45539]_ , \new_[45540]_ , \new_[45543]_ , \new_[45546]_ ,
    \new_[45547]_ , \new_[45548]_ , \new_[45551]_ , \new_[45554]_ ,
    \new_[45555]_ , \new_[45558]_ , \new_[45561]_ , \new_[45562]_ ,
    \new_[45563]_ , \new_[45566]_ , \new_[45569]_ , \new_[45570]_ ,
    \new_[45573]_ , \new_[45576]_ , \new_[45577]_ , \new_[45578]_ ,
    \new_[45581]_ , \new_[45584]_ , \new_[45585]_ , \new_[45588]_ ,
    \new_[45591]_ , \new_[45592]_ , \new_[45593]_ , \new_[45596]_ ,
    \new_[45599]_ , \new_[45600]_ , \new_[45603]_ , \new_[45606]_ ,
    \new_[45607]_ , \new_[45608]_ , \new_[45611]_ , \new_[45614]_ ,
    \new_[45615]_ , \new_[45618]_ , \new_[45621]_ , \new_[45622]_ ,
    \new_[45623]_ , \new_[45626]_ , \new_[45629]_ , \new_[45630]_ ,
    \new_[45633]_ , \new_[45636]_ , \new_[45637]_ , \new_[45638]_ ,
    \new_[45641]_ , \new_[45644]_ , \new_[45645]_ , \new_[45648]_ ,
    \new_[45651]_ , \new_[45652]_ , \new_[45653]_ , \new_[45656]_ ,
    \new_[45659]_ , \new_[45660]_ , \new_[45663]_ , \new_[45666]_ ,
    \new_[45667]_ , \new_[45668]_ , \new_[45671]_ , \new_[45674]_ ,
    \new_[45675]_ , \new_[45678]_ , \new_[45681]_ , \new_[45682]_ ,
    \new_[45683]_ , \new_[45686]_ , \new_[45689]_ , \new_[45690]_ ,
    \new_[45693]_ , \new_[45696]_ , \new_[45697]_ , \new_[45698]_ ,
    \new_[45701]_ , \new_[45704]_ , \new_[45705]_ , \new_[45708]_ ,
    \new_[45711]_ , \new_[45712]_ , \new_[45713]_ , \new_[45716]_ ,
    \new_[45719]_ , \new_[45720]_ , \new_[45723]_ , \new_[45726]_ ,
    \new_[45727]_ , \new_[45728]_ , \new_[45731]_ , \new_[45734]_ ,
    \new_[45735]_ , \new_[45738]_ , \new_[45741]_ , \new_[45742]_ ,
    \new_[45743]_ , \new_[45746]_ , \new_[45749]_ , \new_[45750]_ ,
    \new_[45753]_ , \new_[45756]_ , \new_[45757]_ , \new_[45758]_ ,
    \new_[45761]_ , \new_[45764]_ , \new_[45765]_ , \new_[45768]_ ,
    \new_[45771]_ , \new_[45772]_ , \new_[45773]_ , \new_[45776]_ ,
    \new_[45779]_ , \new_[45780]_ , \new_[45783]_ , \new_[45786]_ ,
    \new_[45787]_ , \new_[45788]_ , \new_[45791]_ , \new_[45794]_ ,
    \new_[45795]_ , \new_[45798]_ , \new_[45801]_ , \new_[45802]_ ,
    \new_[45803]_ , \new_[45806]_ , \new_[45809]_ , \new_[45810]_ ,
    \new_[45813]_ , \new_[45816]_ , \new_[45817]_ , \new_[45818]_ ,
    \new_[45821]_ , \new_[45824]_ , \new_[45825]_ , \new_[45828]_ ,
    \new_[45831]_ , \new_[45832]_ , \new_[45833]_ , \new_[45836]_ ,
    \new_[45839]_ , \new_[45840]_ , \new_[45843]_ , \new_[45846]_ ,
    \new_[45847]_ , \new_[45848]_ , \new_[45851]_ , \new_[45854]_ ,
    \new_[45855]_ , \new_[45858]_ , \new_[45861]_ , \new_[45862]_ ,
    \new_[45863]_ , \new_[45866]_ , \new_[45869]_ , \new_[45870]_ ,
    \new_[45873]_ , \new_[45876]_ , \new_[45877]_ , \new_[45878]_ ,
    \new_[45881]_ , \new_[45884]_ , \new_[45885]_ , \new_[45888]_ ,
    \new_[45891]_ , \new_[45892]_ , \new_[45893]_ , \new_[45896]_ ,
    \new_[45899]_ , \new_[45900]_ , \new_[45903]_ , \new_[45906]_ ,
    \new_[45907]_ , \new_[45908]_ , \new_[45911]_ , \new_[45914]_ ,
    \new_[45915]_ , \new_[45918]_ , \new_[45921]_ , \new_[45922]_ ,
    \new_[45923]_ , \new_[45926]_ , \new_[45929]_ , \new_[45930]_ ,
    \new_[45933]_ , \new_[45936]_ , \new_[45937]_ , \new_[45938]_ ,
    \new_[45941]_ , \new_[45944]_ , \new_[45945]_ , \new_[45948]_ ,
    \new_[45951]_ , \new_[45952]_ , \new_[45953]_ , \new_[45956]_ ,
    \new_[45959]_ , \new_[45960]_ , \new_[45963]_ , \new_[45966]_ ,
    \new_[45967]_ , \new_[45968]_ , \new_[45971]_ , \new_[45974]_ ,
    \new_[45975]_ , \new_[45978]_ , \new_[45981]_ , \new_[45982]_ ,
    \new_[45983]_ , \new_[45986]_ , \new_[45989]_ , \new_[45990]_ ,
    \new_[45993]_ , \new_[45996]_ , \new_[45997]_ , \new_[45998]_ ,
    \new_[46001]_ , \new_[46004]_ , \new_[46005]_ , \new_[46008]_ ,
    \new_[46011]_ , \new_[46012]_ , \new_[46013]_ , \new_[46016]_ ,
    \new_[46019]_ , \new_[46020]_ , \new_[46023]_ , \new_[46026]_ ,
    \new_[46027]_ , \new_[46028]_ , \new_[46031]_ , \new_[46034]_ ,
    \new_[46035]_ , \new_[46038]_ , \new_[46041]_ , \new_[46042]_ ,
    \new_[46043]_ , \new_[46046]_ , \new_[46049]_ , \new_[46050]_ ,
    \new_[46053]_ , \new_[46056]_ , \new_[46057]_ , \new_[46058]_ ,
    \new_[46061]_ , \new_[46064]_ , \new_[46065]_ , \new_[46068]_ ,
    \new_[46071]_ , \new_[46072]_ , \new_[46073]_ , \new_[46076]_ ,
    \new_[46079]_ , \new_[46080]_ , \new_[46083]_ , \new_[46086]_ ,
    \new_[46087]_ , \new_[46088]_ , \new_[46091]_ , \new_[46094]_ ,
    \new_[46095]_ , \new_[46098]_ , \new_[46101]_ , \new_[46102]_ ,
    \new_[46103]_ , \new_[46106]_ , \new_[46109]_ , \new_[46110]_ ,
    \new_[46113]_ , \new_[46116]_ , \new_[46117]_ , \new_[46118]_ ,
    \new_[46121]_ , \new_[46124]_ , \new_[46125]_ , \new_[46128]_ ,
    \new_[46131]_ , \new_[46132]_ , \new_[46133]_ , \new_[46136]_ ,
    \new_[46139]_ , \new_[46140]_ , \new_[46143]_ , \new_[46146]_ ,
    \new_[46147]_ , \new_[46148]_ , \new_[46151]_ , \new_[46154]_ ,
    \new_[46155]_ , \new_[46158]_ , \new_[46161]_ , \new_[46162]_ ,
    \new_[46163]_ , \new_[46166]_ , \new_[46169]_ , \new_[46170]_ ,
    \new_[46173]_ , \new_[46176]_ , \new_[46177]_ , \new_[46178]_ ,
    \new_[46181]_ , \new_[46184]_ , \new_[46185]_ , \new_[46188]_ ,
    \new_[46191]_ , \new_[46192]_ , \new_[46193]_ , \new_[46196]_ ,
    \new_[46199]_ , \new_[46200]_ , \new_[46203]_ , \new_[46206]_ ,
    \new_[46207]_ , \new_[46208]_ , \new_[46211]_ , \new_[46214]_ ,
    \new_[46215]_ , \new_[46218]_ , \new_[46221]_ , \new_[46222]_ ,
    \new_[46223]_ , \new_[46226]_ , \new_[46229]_ , \new_[46230]_ ,
    \new_[46233]_ , \new_[46236]_ , \new_[46237]_ , \new_[46238]_ ,
    \new_[46241]_ , \new_[46244]_ , \new_[46245]_ , \new_[46248]_ ,
    \new_[46251]_ , \new_[46252]_ , \new_[46253]_ , \new_[46256]_ ,
    \new_[46259]_ , \new_[46260]_ , \new_[46263]_ , \new_[46266]_ ,
    \new_[46267]_ , \new_[46268]_ , \new_[46271]_ , \new_[46274]_ ,
    \new_[46275]_ , \new_[46278]_ , \new_[46281]_ , \new_[46282]_ ,
    \new_[46283]_ , \new_[46286]_ , \new_[46289]_ , \new_[46290]_ ,
    \new_[46293]_ , \new_[46296]_ , \new_[46297]_ , \new_[46298]_ ,
    \new_[46301]_ , \new_[46304]_ , \new_[46305]_ , \new_[46308]_ ,
    \new_[46311]_ , \new_[46312]_ , \new_[46313]_ , \new_[46316]_ ,
    \new_[46319]_ , \new_[46320]_ , \new_[46323]_ , \new_[46326]_ ,
    \new_[46327]_ , \new_[46328]_ , \new_[46331]_ , \new_[46334]_ ,
    \new_[46335]_ , \new_[46338]_ , \new_[46341]_ , \new_[46342]_ ,
    \new_[46343]_ , \new_[46346]_ , \new_[46349]_ , \new_[46350]_ ,
    \new_[46353]_ , \new_[46356]_ , \new_[46357]_ , \new_[46358]_ ,
    \new_[46361]_ , \new_[46364]_ , \new_[46365]_ , \new_[46368]_ ,
    \new_[46371]_ , \new_[46372]_ , \new_[46373]_ , \new_[46376]_ ,
    \new_[46379]_ , \new_[46380]_ , \new_[46383]_ , \new_[46386]_ ,
    \new_[46387]_ , \new_[46388]_ , \new_[46391]_ , \new_[46394]_ ,
    \new_[46395]_ , \new_[46398]_ , \new_[46401]_ , \new_[46402]_ ,
    \new_[46403]_ , \new_[46406]_ , \new_[46409]_ , \new_[46410]_ ,
    \new_[46413]_ , \new_[46416]_ , \new_[46417]_ , \new_[46418]_ ,
    \new_[46421]_ , \new_[46424]_ , \new_[46425]_ , \new_[46428]_ ,
    \new_[46431]_ , \new_[46432]_ , \new_[46433]_ , \new_[46436]_ ,
    \new_[46439]_ , \new_[46440]_ , \new_[46443]_ , \new_[46446]_ ,
    \new_[46447]_ , \new_[46448]_ , \new_[46451]_ , \new_[46454]_ ,
    \new_[46455]_ , \new_[46458]_ , \new_[46461]_ , \new_[46462]_ ,
    \new_[46463]_ , \new_[46466]_ , \new_[46469]_ , \new_[46470]_ ,
    \new_[46473]_ , \new_[46476]_ , \new_[46477]_ , \new_[46478]_ ,
    \new_[46481]_ , \new_[46484]_ , \new_[46485]_ , \new_[46488]_ ,
    \new_[46491]_ , \new_[46492]_ , \new_[46493]_ , \new_[46496]_ ,
    \new_[46499]_ , \new_[46500]_ , \new_[46503]_ , \new_[46506]_ ,
    \new_[46507]_ , \new_[46508]_ , \new_[46511]_ , \new_[46514]_ ,
    \new_[46515]_ , \new_[46518]_ , \new_[46521]_ , \new_[46522]_ ,
    \new_[46523]_ , \new_[46526]_ , \new_[46529]_ , \new_[46530]_ ,
    \new_[46533]_ , \new_[46536]_ , \new_[46537]_ , \new_[46538]_ ,
    \new_[46541]_ , \new_[46544]_ , \new_[46545]_ , \new_[46548]_ ,
    \new_[46551]_ , \new_[46552]_ , \new_[46553]_ , \new_[46556]_ ,
    \new_[46559]_ , \new_[46560]_ , \new_[46563]_ , \new_[46566]_ ,
    \new_[46567]_ , \new_[46568]_ , \new_[46571]_ , \new_[46574]_ ,
    \new_[46575]_ , \new_[46578]_ , \new_[46581]_ , \new_[46582]_ ,
    \new_[46583]_ , \new_[46586]_ , \new_[46589]_ , \new_[46590]_ ,
    \new_[46593]_ , \new_[46596]_ , \new_[46597]_ , \new_[46598]_ ,
    \new_[46601]_ , \new_[46604]_ , \new_[46605]_ , \new_[46608]_ ,
    \new_[46611]_ , \new_[46612]_ , \new_[46613]_ , \new_[46616]_ ,
    \new_[46619]_ , \new_[46620]_ , \new_[46623]_ , \new_[46626]_ ,
    \new_[46627]_ , \new_[46628]_ , \new_[46631]_ , \new_[46634]_ ,
    \new_[46635]_ , \new_[46638]_ , \new_[46641]_ , \new_[46642]_ ,
    \new_[46643]_ , \new_[46646]_ , \new_[46649]_ , \new_[46650]_ ,
    \new_[46653]_ , \new_[46656]_ , \new_[46657]_ , \new_[46658]_ ,
    \new_[46661]_ , \new_[46664]_ , \new_[46665]_ , \new_[46668]_ ,
    \new_[46671]_ , \new_[46672]_ , \new_[46673]_ , \new_[46676]_ ,
    \new_[46679]_ , \new_[46680]_ , \new_[46683]_ , \new_[46686]_ ,
    \new_[46687]_ , \new_[46688]_ , \new_[46691]_ , \new_[46694]_ ,
    \new_[46695]_ , \new_[46698]_ , \new_[46701]_ , \new_[46702]_ ,
    \new_[46703]_ , \new_[46706]_ , \new_[46709]_ , \new_[46710]_ ,
    \new_[46713]_ , \new_[46716]_ , \new_[46717]_ , \new_[46718]_ ,
    \new_[46721]_ , \new_[46724]_ , \new_[46725]_ , \new_[46728]_ ,
    \new_[46731]_ , \new_[46732]_ , \new_[46733]_ , \new_[46736]_ ,
    \new_[46739]_ , \new_[46740]_ , \new_[46743]_ , \new_[46746]_ ,
    \new_[46747]_ , \new_[46748]_ , \new_[46751]_ , \new_[46754]_ ,
    \new_[46755]_ , \new_[46758]_ , \new_[46761]_ , \new_[46762]_ ,
    \new_[46763]_ , \new_[46766]_ , \new_[46769]_ , \new_[46770]_ ,
    \new_[46773]_ , \new_[46776]_ , \new_[46777]_ , \new_[46778]_ ,
    \new_[46781]_ , \new_[46784]_ , \new_[46785]_ , \new_[46788]_ ,
    \new_[46791]_ , \new_[46792]_ , \new_[46793]_ , \new_[46796]_ ,
    \new_[46799]_ , \new_[46800]_ , \new_[46803]_ , \new_[46806]_ ,
    \new_[46807]_ , \new_[46808]_ , \new_[46811]_ , \new_[46814]_ ,
    \new_[46815]_ , \new_[46818]_ , \new_[46821]_ , \new_[46822]_ ,
    \new_[46823]_ , \new_[46826]_ , \new_[46829]_ , \new_[46830]_ ,
    \new_[46833]_ , \new_[46836]_ , \new_[46837]_ , \new_[46838]_ ,
    \new_[46841]_ , \new_[46844]_ , \new_[46845]_ , \new_[46848]_ ,
    \new_[46851]_ , \new_[46852]_ , \new_[46853]_ , \new_[46856]_ ,
    \new_[46859]_ , \new_[46860]_ , \new_[46863]_ , \new_[46866]_ ,
    \new_[46867]_ , \new_[46868]_ , \new_[46871]_ , \new_[46874]_ ,
    \new_[46875]_ , \new_[46878]_ , \new_[46881]_ , \new_[46882]_ ,
    \new_[46883]_ , \new_[46886]_ , \new_[46889]_ , \new_[46890]_ ,
    \new_[46893]_ , \new_[46896]_ , \new_[46897]_ , \new_[46898]_ ,
    \new_[46901]_ , \new_[46904]_ , \new_[46905]_ , \new_[46908]_ ,
    \new_[46911]_ , \new_[46912]_ , \new_[46913]_ , \new_[46916]_ ,
    \new_[46919]_ , \new_[46920]_ , \new_[46923]_ , \new_[46926]_ ,
    \new_[46927]_ , \new_[46928]_ , \new_[46931]_ , \new_[46934]_ ,
    \new_[46935]_ , \new_[46938]_ , \new_[46941]_ , \new_[46942]_ ,
    \new_[46943]_ , \new_[46946]_ , \new_[46949]_ , \new_[46950]_ ,
    \new_[46953]_ , \new_[46956]_ , \new_[46957]_ , \new_[46958]_ ,
    \new_[46961]_ , \new_[46964]_ , \new_[46965]_ , \new_[46968]_ ,
    \new_[46971]_ , \new_[46972]_ , \new_[46973]_ , \new_[46976]_ ,
    \new_[46979]_ , \new_[46980]_ , \new_[46983]_ , \new_[46986]_ ,
    \new_[46987]_ , \new_[46988]_ , \new_[46991]_ , \new_[46994]_ ,
    \new_[46995]_ , \new_[46998]_ , \new_[47001]_ , \new_[47002]_ ,
    \new_[47003]_ , \new_[47006]_ , \new_[47009]_ , \new_[47010]_ ,
    \new_[47013]_ , \new_[47016]_ , \new_[47017]_ , \new_[47018]_ ,
    \new_[47021]_ , \new_[47024]_ , \new_[47025]_ , \new_[47028]_ ,
    \new_[47031]_ , \new_[47032]_ , \new_[47033]_ , \new_[47036]_ ,
    \new_[47039]_ , \new_[47040]_ , \new_[47043]_ , \new_[47046]_ ,
    \new_[47047]_ , \new_[47048]_ , \new_[47051]_ , \new_[47054]_ ,
    \new_[47055]_ , \new_[47058]_ , \new_[47061]_ , \new_[47062]_ ,
    \new_[47063]_ , \new_[47066]_ , \new_[47069]_ , \new_[47070]_ ,
    \new_[47073]_ , \new_[47076]_ , \new_[47077]_ , \new_[47078]_ ,
    \new_[47081]_ , \new_[47084]_ , \new_[47085]_ , \new_[47088]_ ,
    \new_[47091]_ , \new_[47092]_ , \new_[47093]_ , \new_[47096]_ ,
    \new_[47099]_ , \new_[47100]_ , \new_[47103]_ , \new_[47106]_ ,
    \new_[47107]_ , \new_[47108]_ , \new_[47111]_ , \new_[47114]_ ,
    \new_[47115]_ , \new_[47118]_ , \new_[47121]_ , \new_[47122]_ ,
    \new_[47123]_ , \new_[47126]_ , \new_[47129]_ , \new_[47130]_ ,
    \new_[47133]_ , \new_[47136]_ , \new_[47137]_ , \new_[47138]_ ,
    \new_[47141]_ , \new_[47144]_ , \new_[47145]_ , \new_[47148]_ ,
    \new_[47151]_ , \new_[47152]_ , \new_[47153]_ , \new_[47156]_ ,
    \new_[47159]_ , \new_[47160]_ , \new_[47163]_ , \new_[47166]_ ,
    \new_[47167]_ , \new_[47168]_ , \new_[47171]_ , \new_[47174]_ ,
    \new_[47175]_ , \new_[47178]_ , \new_[47181]_ , \new_[47182]_ ,
    \new_[47183]_ , \new_[47186]_ , \new_[47189]_ , \new_[47190]_ ,
    \new_[47193]_ , \new_[47196]_ , \new_[47197]_ , \new_[47198]_ ,
    \new_[47201]_ , \new_[47204]_ , \new_[47205]_ , \new_[47208]_ ,
    \new_[47211]_ , \new_[47212]_ , \new_[47213]_ , \new_[47216]_ ,
    \new_[47219]_ , \new_[47220]_ , \new_[47223]_ , \new_[47226]_ ,
    \new_[47227]_ , \new_[47228]_ , \new_[47231]_ , \new_[47234]_ ,
    \new_[47235]_ , \new_[47238]_ , \new_[47241]_ , \new_[47242]_ ,
    \new_[47243]_ , \new_[47246]_ , \new_[47249]_ , \new_[47250]_ ,
    \new_[47253]_ , \new_[47256]_ , \new_[47257]_ , \new_[47258]_ ,
    \new_[47261]_ , \new_[47264]_ , \new_[47265]_ , \new_[47268]_ ,
    \new_[47271]_ , \new_[47272]_ , \new_[47273]_ , \new_[47276]_ ,
    \new_[47279]_ , \new_[47280]_ , \new_[47283]_ , \new_[47286]_ ,
    \new_[47287]_ , \new_[47288]_ , \new_[47291]_ , \new_[47294]_ ,
    \new_[47295]_ , \new_[47298]_ , \new_[47301]_ , \new_[47302]_ ,
    \new_[47303]_ , \new_[47306]_ , \new_[47309]_ , \new_[47310]_ ,
    \new_[47313]_ , \new_[47316]_ , \new_[47317]_ , \new_[47318]_ ,
    \new_[47321]_ , \new_[47324]_ , \new_[47325]_ , \new_[47328]_ ,
    \new_[47331]_ , \new_[47332]_ , \new_[47333]_ , \new_[47336]_ ,
    \new_[47339]_ , \new_[47340]_ , \new_[47343]_ , \new_[47346]_ ,
    \new_[47347]_ , \new_[47348]_ , \new_[47351]_ , \new_[47354]_ ,
    \new_[47355]_ , \new_[47358]_ , \new_[47361]_ , \new_[47362]_ ,
    \new_[47363]_ , \new_[47366]_ , \new_[47369]_ , \new_[47370]_ ,
    \new_[47373]_ , \new_[47376]_ , \new_[47377]_ , \new_[47378]_ ,
    \new_[47381]_ , \new_[47384]_ , \new_[47385]_ , \new_[47388]_ ,
    \new_[47391]_ , \new_[47392]_ , \new_[47393]_ , \new_[47396]_ ,
    \new_[47399]_ , \new_[47400]_ , \new_[47403]_ , \new_[47406]_ ,
    \new_[47407]_ , \new_[47408]_ , \new_[47411]_ , \new_[47414]_ ,
    \new_[47415]_ , \new_[47418]_ , \new_[47421]_ , \new_[47422]_ ,
    \new_[47423]_ , \new_[47426]_ , \new_[47429]_ , \new_[47430]_ ,
    \new_[47433]_ , \new_[47436]_ , \new_[47437]_ , \new_[47438]_ ,
    \new_[47441]_ , \new_[47444]_ , \new_[47445]_ , \new_[47448]_ ,
    \new_[47451]_ , \new_[47452]_ , \new_[47453]_ , \new_[47456]_ ,
    \new_[47459]_ , \new_[47460]_ , \new_[47463]_ , \new_[47466]_ ,
    \new_[47467]_ , \new_[47468]_ , \new_[47471]_ , \new_[47474]_ ,
    \new_[47475]_ , \new_[47478]_ , \new_[47481]_ , \new_[47482]_ ,
    \new_[47483]_ , \new_[47486]_ , \new_[47489]_ , \new_[47490]_ ,
    \new_[47493]_ , \new_[47496]_ , \new_[47497]_ , \new_[47498]_ ,
    \new_[47501]_ , \new_[47504]_ , \new_[47505]_ , \new_[47508]_ ,
    \new_[47511]_ , \new_[47512]_ , \new_[47513]_ , \new_[47516]_ ,
    \new_[47519]_ , \new_[47520]_ , \new_[47523]_ , \new_[47526]_ ,
    \new_[47527]_ , \new_[47528]_ , \new_[47531]_ , \new_[47534]_ ,
    \new_[47535]_ , \new_[47538]_ , \new_[47541]_ , \new_[47542]_ ,
    \new_[47543]_ , \new_[47546]_ , \new_[47549]_ , \new_[47550]_ ,
    \new_[47553]_ , \new_[47556]_ , \new_[47557]_ , \new_[47558]_ ,
    \new_[47561]_ , \new_[47564]_ , \new_[47565]_ , \new_[47568]_ ,
    \new_[47571]_ , \new_[47572]_ , \new_[47573]_ , \new_[47576]_ ,
    \new_[47579]_ , \new_[47580]_ , \new_[47583]_ , \new_[47586]_ ,
    \new_[47587]_ , \new_[47588]_ , \new_[47591]_ , \new_[47594]_ ,
    \new_[47595]_ , \new_[47598]_ , \new_[47601]_ , \new_[47602]_ ,
    \new_[47603]_ , \new_[47606]_ , \new_[47609]_ , \new_[47610]_ ,
    \new_[47613]_ , \new_[47616]_ , \new_[47617]_ , \new_[47618]_ ,
    \new_[47621]_ , \new_[47624]_ , \new_[47625]_ , \new_[47628]_ ,
    \new_[47631]_ , \new_[47632]_ , \new_[47633]_ , \new_[47636]_ ,
    \new_[47639]_ , \new_[47640]_ , \new_[47643]_ , \new_[47646]_ ,
    \new_[47647]_ , \new_[47648]_ , \new_[47651]_ , \new_[47654]_ ,
    \new_[47655]_ , \new_[47658]_ , \new_[47661]_ , \new_[47662]_ ,
    \new_[47663]_ , \new_[47666]_ , \new_[47669]_ , \new_[47670]_ ,
    \new_[47673]_ , \new_[47676]_ , \new_[47677]_ , \new_[47678]_ ,
    \new_[47681]_ , \new_[47684]_ , \new_[47685]_ , \new_[47688]_ ,
    \new_[47691]_ , \new_[47692]_ , \new_[47693]_ , \new_[47696]_ ,
    \new_[47699]_ , \new_[47700]_ , \new_[47703]_ , \new_[47706]_ ,
    \new_[47707]_ , \new_[47708]_ , \new_[47711]_ , \new_[47714]_ ,
    \new_[47715]_ , \new_[47718]_ , \new_[47721]_ , \new_[47722]_ ,
    \new_[47723]_ , \new_[47726]_ , \new_[47729]_ , \new_[47730]_ ,
    \new_[47733]_ , \new_[47736]_ , \new_[47737]_ , \new_[47738]_ ,
    \new_[47741]_ , \new_[47744]_ , \new_[47745]_ , \new_[47748]_ ,
    \new_[47751]_ , \new_[47752]_ , \new_[47753]_ , \new_[47756]_ ,
    \new_[47759]_ , \new_[47760]_ , \new_[47763]_ , \new_[47766]_ ,
    \new_[47767]_ , \new_[47768]_ , \new_[47771]_ , \new_[47774]_ ,
    \new_[47775]_ , \new_[47778]_ , \new_[47781]_ , \new_[47782]_ ,
    \new_[47783]_ , \new_[47786]_ , \new_[47789]_ , \new_[47790]_ ,
    \new_[47793]_ , \new_[47796]_ , \new_[47797]_ , \new_[47798]_ ,
    \new_[47801]_ , \new_[47804]_ , \new_[47805]_ , \new_[47808]_ ,
    \new_[47811]_ , \new_[47812]_ , \new_[47813]_ , \new_[47816]_ ,
    \new_[47819]_ , \new_[47820]_ , \new_[47823]_ , \new_[47826]_ ,
    \new_[47827]_ , \new_[47828]_ , \new_[47831]_ , \new_[47834]_ ,
    \new_[47835]_ , \new_[47838]_ , \new_[47841]_ , \new_[47842]_ ,
    \new_[47843]_ , \new_[47846]_ , \new_[47849]_ , \new_[47850]_ ,
    \new_[47853]_ , \new_[47856]_ , \new_[47857]_ , \new_[47858]_ ,
    \new_[47861]_ , \new_[47864]_ , \new_[47865]_ , \new_[47868]_ ,
    \new_[47871]_ , \new_[47872]_ , \new_[47873]_ , \new_[47876]_ ,
    \new_[47879]_ , \new_[47880]_ , \new_[47883]_ , \new_[47886]_ ,
    \new_[47887]_ , \new_[47888]_ , \new_[47891]_ , \new_[47894]_ ,
    \new_[47895]_ , \new_[47898]_ , \new_[47901]_ , \new_[47902]_ ,
    \new_[47903]_ , \new_[47906]_ , \new_[47909]_ , \new_[47910]_ ,
    \new_[47913]_ , \new_[47916]_ , \new_[47917]_ , \new_[47918]_ ,
    \new_[47921]_ , \new_[47924]_ , \new_[47925]_ , \new_[47928]_ ,
    \new_[47931]_ , \new_[47932]_ , \new_[47933]_ , \new_[47936]_ ,
    \new_[47939]_ , \new_[47940]_ , \new_[47943]_ , \new_[47946]_ ,
    \new_[47947]_ , \new_[47948]_ , \new_[47951]_ , \new_[47954]_ ,
    \new_[47955]_ , \new_[47958]_ , \new_[47961]_ , \new_[47962]_ ,
    \new_[47963]_ , \new_[47966]_ , \new_[47969]_ , \new_[47970]_ ,
    \new_[47973]_ , \new_[47976]_ , \new_[47977]_ , \new_[47978]_ ,
    \new_[47981]_ , \new_[47984]_ , \new_[47985]_ , \new_[47988]_ ,
    \new_[47991]_ , \new_[47992]_ , \new_[47993]_ , \new_[47996]_ ,
    \new_[47999]_ , \new_[48000]_ , \new_[48003]_ , \new_[48006]_ ,
    \new_[48007]_ , \new_[48008]_ , \new_[48011]_ , \new_[48014]_ ,
    \new_[48015]_ , \new_[48018]_ , \new_[48021]_ , \new_[48022]_ ,
    \new_[48023]_ , \new_[48026]_ , \new_[48029]_ , \new_[48030]_ ,
    \new_[48033]_ , \new_[48036]_ , \new_[48037]_ , \new_[48038]_ ,
    \new_[48041]_ , \new_[48044]_ , \new_[48045]_ , \new_[48048]_ ,
    \new_[48051]_ , \new_[48052]_ , \new_[48053]_ , \new_[48056]_ ,
    \new_[48059]_ , \new_[48060]_ , \new_[48063]_ , \new_[48066]_ ,
    \new_[48067]_ , \new_[48068]_ , \new_[48071]_ , \new_[48074]_ ,
    \new_[48075]_ , \new_[48078]_ , \new_[48081]_ , \new_[48082]_ ,
    \new_[48083]_ , \new_[48086]_ , \new_[48089]_ , \new_[48090]_ ,
    \new_[48093]_ , \new_[48096]_ , \new_[48097]_ , \new_[48098]_ ,
    \new_[48101]_ , \new_[48104]_ , \new_[48105]_ , \new_[48108]_ ,
    \new_[48111]_ , \new_[48112]_ , \new_[48113]_ , \new_[48116]_ ,
    \new_[48119]_ , \new_[48120]_ , \new_[48123]_ , \new_[48126]_ ,
    \new_[48127]_ , \new_[48128]_ , \new_[48131]_ , \new_[48134]_ ,
    \new_[48135]_ , \new_[48138]_ , \new_[48141]_ , \new_[48142]_ ,
    \new_[48143]_ , \new_[48146]_ , \new_[48149]_ , \new_[48150]_ ,
    \new_[48153]_ , \new_[48156]_ , \new_[48157]_ , \new_[48158]_ ,
    \new_[48161]_ , \new_[48164]_ , \new_[48165]_ , \new_[48168]_ ,
    \new_[48171]_ , \new_[48172]_ , \new_[48173]_ , \new_[48176]_ ,
    \new_[48179]_ , \new_[48180]_ , \new_[48183]_ , \new_[48186]_ ,
    \new_[48187]_ , \new_[48188]_ , \new_[48191]_ , \new_[48194]_ ,
    \new_[48195]_ , \new_[48198]_ , \new_[48201]_ , \new_[48202]_ ,
    \new_[48203]_ , \new_[48206]_ , \new_[48209]_ , \new_[48210]_ ,
    \new_[48213]_ , \new_[48216]_ , \new_[48217]_ , \new_[48218]_ ,
    \new_[48221]_ , \new_[48224]_ , \new_[48225]_ , \new_[48228]_ ,
    \new_[48231]_ , \new_[48232]_ , \new_[48233]_ , \new_[48236]_ ,
    \new_[48239]_ , \new_[48240]_ , \new_[48243]_ , \new_[48246]_ ,
    \new_[48247]_ , \new_[48248]_ , \new_[48251]_ , \new_[48254]_ ,
    \new_[48255]_ , \new_[48258]_ , \new_[48261]_ , \new_[48262]_ ,
    \new_[48263]_ , \new_[48266]_ , \new_[48269]_ , \new_[48270]_ ,
    \new_[48273]_ , \new_[48276]_ , \new_[48277]_ , \new_[48278]_ ,
    \new_[48281]_ , \new_[48284]_ , \new_[48285]_ , \new_[48288]_ ,
    \new_[48291]_ , \new_[48292]_ , \new_[48293]_ , \new_[48296]_ ,
    \new_[48299]_ , \new_[48300]_ , \new_[48303]_ , \new_[48306]_ ,
    \new_[48307]_ , \new_[48308]_ , \new_[48311]_ , \new_[48314]_ ,
    \new_[48315]_ , \new_[48318]_ , \new_[48321]_ , \new_[48322]_ ,
    \new_[48323]_ , \new_[48326]_ , \new_[48329]_ , \new_[48330]_ ,
    \new_[48333]_ , \new_[48336]_ , \new_[48337]_ , \new_[48338]_ ,
    \new_[48341]_ , \new_[48344]_ , \new_[48345]_ , \new_[48348]_ ,
    \new_[48351]_ , \new_[48352]_ , \new_[48353]_ , \new_[48356]_ ,
    \new_[48359]_ , \new_[48360]_ , \new_[48363]_ , \new_[48366]_ ,
    \new_[48367]_ , \new_[48368]_ , \new_[48371]_ , \new_[48374]_ ,
    \new_[48375]_ , \new_[48378]_ , \new_[48381]_ , \new_[48382]_ ,
    \new_[48383]_ , \new_[48386]_ , \new_[48389]_ , \new_[48390]_ ,
    \new_[48393]_ , \new_[48396]_ , \new_[48397]_ , \new_[48398]_ ,
    \new_[48401]_ , \new_[48404]_ , \new_[48405]_ , \new_[48408]_ ,
    \new_[48411]_ , \new_[48412]_ , \new_[48413]_ , \new_[48416]_ ,
    \new_[48419]_ , \new_[48420]_ , \new_[48423]_ , \new_[48426]_ ,
    \new_[48427]_ , \new_[48428]_ , \new_[48431]_ , \new_[48434]_ ,
    \new_[48435]_ , \new_[48438]_ , \new_[48441]_ , \new_[48442]_ ,
    \new_[48443]_ , \new_[48446]_ , \new_[48449]_ , \new_[48450]_ ,
    \new_[48453]_ , \new_[48456]_ , \new_[48457]_ , \new_[48458]_ ,
    \new_[48461]_ , \new_[48464]_ , \new_[48465]_ , \new_[48468]_ ,
    \new_[48471]_ , \new_[48472]_ , \new_[48473]_ , \new_[48476]_ ,
    \new_[48479]_ , \new_[48480]_ , \new_[48483]_ , \new_[48486]_ ,
    \new_[48487]_ , \new_[48488]_ , \new_[48491]_ , \new_[48494]_ ,
    \new_[48495]_ , \new_[48498]_ , \new_[48501]_ , \new_[48502]_ ,
    \new_[48503]_ , \new_[48506]_ , \new_[48509]_ , \new_[48510]_ ,
    \new_[48513]_ , \new_[48516]_ , \new_[48517]_ , \new_[48518]_ ,
    \new_[48521]_ , \new_[48524]_ , \new_[48525]_ , \new_[48528]_ ,
    \new_[48531]_ , \new_[48532]_ , \new_[48533]_ , \new_[48536]_ ,
    \new_[48539]_ , \new_[48540]_ , \new_[48543]_ , \new_[48546]_ ,
    \new_[48547]_ , \new_[48548]_ , \new_[48551]_ , \new_[48554]_ ,
    \new_[48555]_ , \new_[48558]_ , \new_[48561]_ , \new_[48562]_ ,
    \new_[48563]_ , \new_[48566]_ , \new_[48569]_ , \new_[48570]_ ,
    \new_[48573]_ , \new_[48576]_ , \new_[48577]_ , \new_[48578]_ ,
    \new_[48581]_ , \new_[48584]_ , \new_[48585]_ , \new_[48588]_ ,
    \new_[48591]_ , \new_[48592]_ , \new_[48593]_ , \new_[48596]_ ,
    \new_[48599]_ , \new_[48600]_ , \new_[48603]_ , \new_[48606]_ ,
    \new_[48607]_ , \new_[48608]_ , \new_[48611]_ , \new_[48614]_ ,
    \new_[48615]_ , \new_[48618]_ , \new_[48621]_ , \new_[48622]_ ,
    \new_[48623]_ , \new_[48626]_ , \new_[48629]_ , \new_[48630]_ ,
    \new_[48633]_ , \new_[48636]_ , \new_[48637]_ , \new_[48638]_ ,
    \new_[48641]_ , \new_[48644]_ , \new_[48645]_ , \new_[48648]_ ,
    \new_[48651]_ , \new_[48652]_ , \new_[48653]_ , \new_[48656]_ ,
    \new_[48659]_ , \new_[48660]_ , \new_[48663]_ , \new_[48666]_ ,
    \new_[48667]_ , \new_[48668]_ , \new_[48671]_ , \new_[48674]_ ,
    \new_[48675]_ , \new_[48678]_ , \new_[48681]_ , \new_[48682]_ ,
    \new_[48683]_ , \new_[48686]_ , \new_[48689]_ , \new_[48690]_ ,
    \new_[48693]_ , \new_[48696]_ , \new_[48697]_ , \new_[48698]_ ,
    \new_[48701]_ , \new_[48704]_ , \new_[48705]_ , \new_[48708]_ ,
    \new_[48711]_ , \new_[48712]_ , \new_[48713]_ , \new_[48716]_ ,
    \new_[48719]_ , \new_[48720]_ , \new_[48723]_ , \new_[48726]_ ,
    \new_[48727]_ , \new_[48728]_ , \new_[48731]_ , \new_[48734]_ ,
    \new_[48735]_ , \new_[48738]_ , \new_[48741]_ , \new_[48742]_ ,
    \new_[48743]_ , \new_[48746]_ , \new_[48749]_ , \new_[48750]_ ,
    \new_[48753]_ , \new_[48756]_ , \new_[48757]_ , \new_[48758]_ ,
    \new_[48761]_ , \new_[48764]_ , \new_[48765]_ , \new_[48768]_ ,
    \new_[48771]_ , \new_[48772]_ , \new_[48773]_ , \new_[48776]_ ,
    \new_[48779]_ , \new_[48780]_ , \new_[48783]_ , \new_[48786]_ ,
    \new_[48787]_ , \new_[48788]_ , \new_[48791]_ , \new_[48794]_ ,
    \new_[48795]_ , \new_[48798]_ , \new_[48801]_ , \new_[48802]_ ,
    \new_[48803]_ , \new_[48806]_ , \new_[48809]_ , \new_[48810]_ ,
    \new_[48813]_ , \new_[48816]_ , \new_[48817]_ , \new_[48818]_ ,
    \new_[48821]_ , \new_[48824]_ , \new_[48825]_ , \new_[48828]_ ,
    \new_[48831]_ , \new_[48832]_ , \new_[48833]_ , \new_[48836]_ ,
    \new_[48839]_ , \new_[48840]_ , \new_[48843]_ , \new_[48846]_ ,
    \new_[48847]_ , \new_[48848]_ , \new_[48851]_ , \new_[48854]_ ,
    \new_[48855]_ , \new_[48858]_ , \new_[48861]_ , \new_[48862]_ ,
    \new_[48863]_ , \new_[48866]_ , \new_[48869]_ , \new_[48870]_ ,
    \new_[48873]_ , \new_[48876]_ , \new_[48877]_ , \new_[48878]_ ,
    \new_[48881]_ , \new_[48884]_ , \new_[48885]_ , \new_[48888]_ ,
    \new_[48891]_ , \new_[48892]_ , \new_[48893]_ , \new_[48896]_ ,
    \new_[48899]_ , \new_[48900]_ , \new_[48903]_ , \new_[48906]_ ,
    \new_[48907]_ , \new_[48908]_ , \new_[48911]_ , \new_[48914]_ ,
    \new_[48915]_ , \new_[48918]_ , \new_[48921]_ , \new_[48922]_ ,
    \new_[48923]_ , \new_[48926]_ , \new_[48929]_ , \new_[48930]_ ,
    \new_[48933]_ , \new_[48936]_ , \new_[48937]_ , \new_[48938]_ ,
    \new_[48941]_ , \new_[48944]_ , \new_[48945]_ , \new_[48948]_ ,
    \new_[48951]_ , \new_[48952]_ , \new_[48953]_ , \new_[48956]_ ,
    \new_[48959]_ , \new_[48960]_ , \new_[48963]_ , \new_[48966]_ ,
    \new_[48967]_ , \new_[48968]_ , \new_[48971]_ , \new_[48974]_ ,
    \new_[48975]_ , \new_[48978]_ , \new_[48981]_ , \new_[48982]_ ,
    \new_[48983]_ , \new_[48986]_ , \new_[48989]_ , \new_[48990]_ ,
    \new_[48993]_ , \new_[48996]_ , \new_[48997]_ , \new_[48998]_ ,
    \new_[49001]_ , \new_[49004]_ , \new_[49005]_ , \new_[49008]_ ,
    \new_[49011]_ , \new_[49012]_ , \new_[49013]_ , \new_[49016]_ ,
    \new_[49019]_ , \new_[49020]_ , \new_[49023]_ , \new_[49026]_ ,
    \new_[49027]_ , \new_[49028]_ , \new_[49031]_ , \new_[49034]_ ,
    \new_[49035]_ , \new_[49038]_ , \new_[49041]_ , \new_[49042]_ ,
    \new_[49043]_ , \new_[49046]_ , \new_[49049]_ , \new_[49050]_ ,
    \new_[49053]_ , \new_[49056]_ , \new_[49057]_ , \new_[49058]_ ,
    \new_[49061]_ , \new_[49064]_ , \new_[49065]_ , \new_[49068]_ ,
    \new_[49071]_ , \new_[49072]_ , \new_[49073]_ , \new_[49076]_ ,
    \new_[49079]_ , \new_[49080]_ , \new_[49083]_ , \new_[49086]_ ,
    \new_[49087]_ , \new_[49088]_ , \new_[49091]_ , \new_[49094]_ ,
    \new_[49095]_ , \new_[49098]_ , \new_[49101]_ , \new_[49102]_ ,
    \new_[49103]_ , \new_[49106]_ , \new_[49109]_ , \new_[49110]_ ,
    \new_[49113]_ , \new_[49116]_ , \new_[49117]_ , \new_[49118]_ ,
    \new_[49121]_ , \new_[49124]_ , \new_[49125]_ , \new_[49128]_ ,
    \new_[49131]_ , \new_[49132]_ , \new_[49133]_ , \new_[49136]_ ,
    \new_[49139]_ , \new_[49140]_ , \new_[49143]_ , \new_[49146]_ ,
    \new_[49147]_ , \new_[49148]_ , \new_[49151]_ , \new_[49154]_ ,
    \new_[49155]_ , \new_[49158]_ , \new_[49161]_ , \new_[49162]_ ,
    \new_[49163]_ , \new_[49166]_ , \new_[49169]_ , \new_[49170]_ ,
    \new_[49173]_ , \new_[49176]_ , \new_[49177]_ , \new_[49178]_ ,
    \new_[49181]_ , \new_[49184]_ , \new_[49185]_ , \new_[49188]_ ,
    \new_[49191]_ , \new_[49192]_ , \new_[49193]_ , \new_[49196]_ ,
    \new_[49199]_ , \new_[49200]_ , \new_[49203]_ , \new_[49206]_ ,
    \new_[49207]_ , \new_[49208]_ , \new_[49211]_ , \new_[49214]_ ,
    \new_[49215]_ , \new_[49218]_ , \new_[49221]_ , \new_[49222]_ ,
    \new_[49223]_ , \new_[49226]_ , \new_[49229]_ , \new_[49230]_ ,
    \new_[49233]_ , \new_[49236]_ , \new_[49237]_ , \new_[49238]_ ,
    \new_[49241]_ , \new_[49244]_ , \new_[49245]_ , \new_[49248]_ ,
    \new_[49251]_ , \new_[49252]_ , \new_[49253]_ , \new_[49256]_ ,
    \new_[49259]_ , \new_[49260]_ , \new_[49263]_ , \new_[49266]_ ,
    \new_[49267]_ , \new_[49268]_ , \new_[49271]_ , \new_[49274]_ ,
    \new_[49275]_ , \new_[49278]_ , \new_[49281]_ , \new_[49282]_ ,
    \new_[49283]_ , \new_[49286]_ , \new_[49289]_ , \new_[49290]_ ,
    \new_[49293]_ , \new_[49296]_ , \new_[49297]_ , \new_[49298]_ ,
    \new_[49301]_ , \new_[49304]_ , \new_[49305]_ , \new_[49308]_ ,
    \new_[49311]_ , \new_[49312]_ , \new_[49313]_ , \new_[49316]_ ,
    \new_[49319]_ , \new_[49320]_ , \new_[49323]_ , \new_[49326]_ ,
    \new_[49327]_ , \new_[49328]_ , \new_[49331]_ , \new_[49334]_ ,
    \new_[49335]_ , \new_[49338]_ , \new_[49341]_ , \new_[49342]_ ,
    \new_[49343]_ , \new_[49346]_ , \new_[49349]_ , \new_[49350]_ ,
    \new_[49353]_ , \new_[49356]_ , \new_[49357]_ , \new_[49358]_ ,
    \new_[49361]_ , \new_[49364]_ , \new_[49365]_ , \new_[49368]_ ,
    \new_[49371]_ , \new_[49372]_ , \new_[49373]_ , \new_[49376]_ ,
    \new_[49379]_ , \new_[49380]_ , \new_[49383]_ , \new_[49386]_ ,
    \new_[49387]_ , \new_[49388]_ , \new_[49391]_ , \new_[49394]_ ,
    \new_[49395]_ , \new_[49398]_ , \new_[49401]_ , \new_[49402]_ ,
    \new_[49403]_ , \new_[49406]_ , \new_[49409]_ , \new_[49410]_ ,
    \new_[49413]_ , \new_[49416]_ , \new_[49417]_ , \new_[49418]_ ,
    \new_[49421]_ , \new_[49424]_ , \new_[49425]_ , \new_[49428]_ ,
    \new_[49431]_ , \new_[49432]_ , \new_[49433]_ , \new_[49436]_ ,
    \new_[49439]_ , \new_[49440]_ , \new_[49443]_ , \new_[49446]_ ,
    \new_[49447]_ , \new_[49448]_ , \new_[49451]_ , \new_[49454]_ ,
    \new_[49455]_ , \new_[49458]_ , \new_[49461]_ , \new_[49462]_ ,
    \new_[49463]_ , \new_[49466]_ , \new_[49469]_ , \new_[49470]_ ,
    \new_[49473]_ , \new_[49476]_ , \new_[49477]_ , \new_[49478]_ ,
    \new_[49481]_ , \new_[49484]_ , \new_[49485]_ , \new_[49488]_ ,
    \new_[49491]_ , \new_[49492]_ , \new_[49493]_ , \new_[49496]_ ,
    \new_[49499]_ , \new_[49500]_ , \new_[49503]_ , \new_[49506]_ ,
    \new_[49507]_ , \new_[49508]_ , \new_[49511]_ , \new_[49514]_ ,
    \new_[49515]_ , \new_[49518]_ , \new_[49521]_ , \new_[49522]_ ,
    \new_[49523]_ , \new_[49526]_ , \new_[49529]_ , \new_[49530]_ ,
    \new_[49533]_ , \new_[49536]_ , \new_[49537]_ , \new_[49538]_ ;
  assign A42 = \new_[5254]_  | \new_[3503]_ ;
  assign \new_[1]_  = \new_[49538]_  & \new_[49523]_ ;
  assign \new_[2]_  = \new_[49508]_  & \new_[49493]_ ;
  assign \new_[3]_  = \new_[49478]_  & \new_[49463]_ ;
  assign \new_[4]_  = \new_[49448]_  & \new_[49433]_ ;
  assign \new_[5]_  = \new_[49418]_  & \new_[49403]_ ;
  assign \new_[6]_  = \new_[49388]_  & \new_[49373]_ ;
  assign \new_[7]_  = \new_[49358]_  & \new_[49343]_ ;
  assign \new_[8]_  = \new_[49328]_  & \new_[49313]_ ;
  assign \new_[9]_  = \new_[49298]_  & \new_[49283]_ ;
  assign \new_[10]_  = \new_[49268]_  & \new_[49253]_ ;
  assign \new_[11]_  = \new_[49238]_  & \new_[49223]_ ;
  assign \new_[12]_  = \new_[49208]_  & \new_[49193]_ ;
  assign \new_[13]_  = \new_[49178]_  & \new_[49163]_ ;
  assign \new_[14]_  = \new_[49148]_  & \new_[49133]_ ;
  assign \new_[15]_  = \new_[49118]_  & \new_[49103]_ ;
  assign \new_[16]_  = \new_[49088]_  & \new_[49073]_ ;
  assign \new_[17]_  = \new_[49058]_  & \new_[49043]_ ;
  assign \new_[18]_  = \new_[49028]_  & \new_[49013]_ ;
  assign \new_[19]_  = \new_[48998]_  & \new_[48983]_ ;
  assign \new_[20]_  = \new_[48968]_  & \new_[48953]_ ;
  assign \new_[21]_  = \new_[48938]_  & \new_[48923]_ ;
  assign \new_[22]_  = \new_[48908]_  & \new_[48893]_ ;
  assign \new_[23]_  = \new_[48878]_  & \new_[48863]_ ;
  assign \new_[24]_  = \new_[48848]_  & \new_[48833]_ ;
  assign \new_[25]_  = \new_[48818]_  & \new_[48803]_ ;
  assign \new_[26]_  = \new_[48788]_  & \new_[48773]_ ;
  assign \new_[27]_  = \new_[48758]_  & \new_[48743]_ ;
  assign \new_[28]_  = \new_[48728]_  & \new_[48713]_ ;
  assign \new_[29]_  = \new_[48698]_  & \new_[48683]_ ;
  assign \new_[30]_  = \new_[48668]_  & \new_[48653]_ ;
  assign \new_[31]_  = \new_[48638]_  & \new_[48623]_ ;
  assign \new_[32]_  = \new_[48608]_  & \new_[48593]_ ;
  assign \new_[33]_  = \new_[48578]_  & \new_[48563]_ ;
  assign \new_[34]_  = \new_[48548]_  & \new_[48533]_ ;
  assign \new_[35]_  = \new_[48518]_  & \new_[48503]_ ;
  assign \new_[36]_  = \new_[48488]_  & \new_[48473]_ ;
  assign \new_[37]_  = \new_[48458]_  & \new_[48443]_ ;
  assign \new_[38]_  = \new_[48428]_  & \new_[48413]_ ;
  assign \new_[39]_  = \new_[48398]_  & \new_[48383]_ ;
  assign \new_[40]_  = \new_[48368]_  & \new_[48353]_ ;
  assign \new_[41]_  = \new_[48338]_  & \new_[48323]_ ;
  assign \new_[42]_  = \new_[48308]_  & \new_[48293]_ ;
  assign \new_[43]_  = \new_[48278]_  & \new_[48263]_ ;
  assign \new_[44]_  = \new_[48248]_  & \new_[48233]_ ;
  assign \new_[45]_  = \new_[48218]_  & \new_[48203]_ ;
  assign \new_[46]_  = \new_[48188]_  & \new_[48173]_ ;
  assign \new_[47]_  = \new_[48158]_  & \new_[48143]_ ;
  assign \new_[48]_  = \new_[48128]_  & \new_[48113]_ ;
  assign \new_[49]_  = \new_[48098]_  & \new_[48083]_ ;
  assign \new_[50]_  = \new_[48068]_  & \new_[48053]_ ;
  assign \new_[51]_  = \new_[48038]_  & \new_[48023]_ ;
  assign \new_[52]_  = \new_[48008]_  & \new_[47993]_ ;
  assign \new_[53]_  = \new_[47978]_  & \new_[47963]_ ;
  assign \new_[54]_  = \new_[47948]_  & \new_[47933]_ ;
  assign \new_[55]_  = \new_[47918]_  & \new_[47903]_ ;
  assign \new_[56]_  = \new_[47888]_  & \new_[47873]_ ;
  assign \new_[57]_  = \new_[47858]_  & \new_[47843]_ ;
  assign \new_[58]_  = \new_[47828]_  & \new_[47813]_ ;
  assign \new_[59]_  = \new_[47798]_  & \new_[47783]_ ;
  assign \new_[60]_  = \new_[47768]_  & \new_[47753]_ ;
  assign \new_[61]_  = \new_[47738]_  & \new_[47723]_ ;
  assign \new_[62]_  = \new_[47708]_  & \new_[47693]_ ;
  assign \new_[63]_  = \new_[47678]_  & \new_[47663]_ ;
  assign \new_[64]_  = \new_[47648]_  & \new_[47633]_ ;
  assign \new_[65]_  = \new_[47618]_  & \new_[47603]_ ;
  assign \new_[66]_  = \new_[47588]_  & \new_[47573]_ ;
  assign \new_[67]_  = \new_[47558]_  & \new_[47543]_ ;
  assign \new_[68]_  = \new_[47528]_  & \new_[47513]_ ;
  assign \new_[69]_  = \new_[47498]_  & \new_[47483]_ ;
  assign \new_[70]_  = \new_[47468]_  & \new_[47453]_ ;
  assign \new_[71]_  = \new_[47438]_  & \new_[47423]_ ;
  assign \new_[72]_  = \new_[47408]_  & \new_[47393]_ ;
  assign \new_[73]_  = \new_[47378]_  & \new_[47363]_ ;
  assign \new_[74]_  = \new_[47348]_  & \new_[47333]_ ;
  assign \new_[75]_  = \new_[47318]_  & \new_[47303]_ ;
  assign \new_[76]_  = \new_[47288]_  & \new_[47273]_ ;
  assign \new_[77]_  = \new_[47258]_  & \new_[47243]_ ;
  assign \new_[78]_  = \new_[47228]_  & \new_[47213]_ ;
  assign \new_[79]_  = \new_[47198]_  & \new_[47183]_ ;
  assign \new_[80]_  = \new_[47168]_  & \new_[47153]_ ;
  assign \new_[81]_  = \new_[47138]_  & \new_[47123]_ ;
  assign \new_[82]_  = \new_[47108]_  & \new_[47093]_ ;
  assign \new_[83]_  = \new_[47078]_  & \new_[47063]_ ;
  assign \new_[84]_  = \new_[47048]_  & \new_[47033]_ ;
  assign \new_[85]_  = \new_[47018]_  & \new_[47003]_ ;
  assign \new_[86]_  = \new_[46988]_  & \new_[46973]_ ;
  assign \new_[87]_  = \new_[46958]_  & \new_[46943]_ ;
  assign \new_[88]_  = \new_[46928]_  & \new_[46913]_ ;
  assign \new_[89]_  = \new_[46898]_  & \new_[46883]_ ;
  assign \new_[90]_  = \new_[46868]_  & \new_[46853]_ ;
  assign \new_[91]_  = \new_[46838]_  & \new_[46823]_ ;
  assign \new_[92]_  = \new_[46808]_  & \new_[46793]_ ;
  assign \new_[93]_  = \new_[46778]_  & \new_[46763]_ ;
  assign \new_[94]_  = \new_[46748]_  & \new_[46733]_ ;
  assign \new_[95]_  = \new_[46718]_  & \new_[46703]_ ;
  assign \new_[96]_  = \new_[46688]_  & \new_[46673]_ ;
  assign \new_[97]_  = \new_[46658]_  & \new_[46643]_ ;
  assign \new_[98]_  = \new_[46628]_  & \new_[46613]_ ;
  assign \new_[99]_  = \new_[46598]_  & \new_[46583]_ ;
  assign \new_[100]_  = \new_[46568]_  & \new_[46553]_ ;
  assign \new_[101]_  = \new_[46538]_  & \new_[46523]_ ;
  assign \new_[102]_  = \new_[46508]_  & \new_[46493]_ ;
  assign \new_[103]_  = \new_[46478]_  & \new_[46463]_ ;
  assign \new_[104]_  = \new_[46448]_  & \new_[46433]_ ;
  assign \new_[105]_  = \new_[46418]_  & \new_[46403]_ ;
  assign \new_[106]_  = \new_[46388]_  & \new_[46373]_ ;
  assign \new_[107]_  = \new_[46358]_  & \new_[46343]_ ;
  assign \new_[108]_  = \new_[46328]_  & \new_[46313]_ ;
  assign \new_[109]_  = \new_[46298]_  & \new_[46283]_ ;
  assign \new_[110]_  = \new_[46268]_  & \new_[46253]_ ;
  assign \new_[111]_  = \new_[46238]_  & \new_[46223]_ ;
  assign \new_[112]_  = \new_[46208]_  & \new_[46193]_ ;
  assign \new_[113]_  = \new_[46178]_  & \new_[46163]_ ;
  assign \new_[114]_  = \new_[46148]_  & \new_[46133]_ ;
  assign \new_[115]_  = \new_[46118]_  & \new_[46103]_ ;
  assign \new_[116]_  = \new_[46088]_  & \new_[46073]_ ;
  assign \new_[117]_  = \new_[46058]_  & \new_[46043]_ ;
  assign \new_[118]_  = \new_[46028]_  & \new_[46013]_ ;
  assign \new_[119]_  = \new_[45998]_  & \new_[45983]_ ;
  assign \new_[120]_  = \new_[45968]_  & \new_[45953]_ ;
  assign \new_[121]_  = \new_[45938]_  & \new_[45923]_ ;
  assign \new_[122]_  = \new_[45908]_  & \new_[45893]_ ;
  assign \new_[123]_  = \new_[45878]_  & \new_[45863]_ ;
  assign \new_[124]_  = \new_[45848]_  & \new_[45833]_ ;
  assign \new_[125]_  = \new_[45818]_  & \new_[45803]_ ;
  assign \new_[126]_  = \new_[45788]_  & \new_[45773]_ ;
  assign \new_[127]_  = \new_[45758]_  & \new_[45743]_ ;
  assign \new_[128]_  = \new_[45728]_  & \new_[45713]_ ;
  assign \new_[129]_  = \new_[45698]_  & \new_[45683]_ ;
  assign \new_[130]_  = \new_[45668]_  & \new_[45653]_ ;
  assign \new_[131]_  = \new_[45638]_  & \new_[45623]_ ;
  assign \new_[132]_  = \new_[45608]_  & \new_[45593]_ ;
  assign \new_[133]_  = \new_[45578]_  & \new_[45563]_ ;
  assign \new_[134]_  = \new_[45548]_  & \new_[45533]_ ;
  assign \new_[135]_  = \new_[45518]_  & \new_[45503]_ ;
  assign \new_[136]_  = \new_[45488]_  & \new_[45473]_ ;
  assign \new_[137]_  = \new_[45458]_  & \new_[45443]_ ;
  assign \new_[138]_  = \new_[45428]_  & \new_[45413]_ ;
  assign \new_[139]_  = \new_[45398]_  & \new_[45383]_ ;
  assign \new_[140]_  = \new_[45368]_  & \new_[45353]_ ;
  assign \new_[141]_  = \new_[45338]_  & \new_[45323]_ ;
  assign \new_[142]_  = \new_[45308]_  & \new_[45293]_ ;
  assign \new_[143]_  = \new_[45278]_  & \new_[45263]_ ;
  assign \new_[144]_  = \new_[45248]_  & \new_[45233]_ ;
  assign \new_[145]_  = \new_[45218]_  & \new_[45203]_ ;
  assign \new_[146]_  = \new_[45188]_  & \new_[45173]_ ;
  assign \new_[147]_  = \new_[45158]_  & \new_[45143]_ ;
  assign \new_[148]_  = \new_[45128]_  & \new_[45113]_ ;
  assign \new_[149]_  = \new_[45098]_  & \new_[45083]_ ;
  assign \new_[150]_  = \new_[45068]_  & \new_[45053]_ ;
  assign \new_[151]_  = \new_[45038]_  & \new_[45023]_ ;
  assign \new_[152]_  = \new_[45008]_  & \new_[44993]_ ;
  assign \new_[153]_  = \new_[44978]_  & \new_[44963]_ ;
  assign \new_[154]_  = \new_[44948]_  & \new_[44933]_ ;
  assign \new_[155]_  = \new_[44918]_  & \new_[44903]_ ;
  assign \new_[156]_  = \new_[44888]_  & \new_[44873]_ ;
  assign \new_[157]_  = \new_[44858]_  & \new_[44843]_ ;
  assign \new_[158]_  = \new_[44828]_  & \new_[44813]_ ;
  assign \new_[159]_  = \new_[44798]_  & \new_[44783]_ ;
  assign \new_[160]_  = \new_[44768]_  & \new_[44753]_ ;
  assign \new_[161]_  = \new_[44738]_  & \new_[44723]_ ;
  assign \new_[162]_  = \new_[44708]_  & \new_[44693]_ ;
  assign \new_[163]_  = \new_[44678]_  & \new_[44663]_ ;
  assign \new_[164]_  = \new_[44648]_  & \new_[44633]_ ;
  assign \new_[165]_  = \new_[44618]_  & \new_[44603]_ ;
  assign \new_[166]_  = \new_[44588]_  & \new_[44573]_ ;
  assign \new_[167]_  = \new_[44558]_  & \new_[44543]_ ;
  assign \new_[168]_  = \new_[44528]_  & \new_[44513]_ ;
  assign \new_[169]_  = \new_[44498]_  & \new_[44483]_ ;
  assign \new_[170]_  = \new_[44468]_  & \new_[44453]_ ;
  assign \new_[171]_  = \new_[44438]_  & \new_[44423]_ ;
  assign \new_[172]_  = \new_[44408]_  & \new_[44393]_ ;
  assign \new_[173]_  = \new_[44378]_  & \new_[44363]_ ;
  assign \new_[174]_  = \new_[44348]_  & \new_[44333]_ ;
  assign \new_[175]_  = \new_[44318]_  & \new_[44303]_ ;
  assign \new_[176]_  = \new_[44288]_  & \new_[44273]_ ;
  assign \new_[177]_  = \new_[44258]_  & \new_[44243]_ ;
  assign \new_[178]_  = \new_[44228]_  & \new_[44213]_ ;
  assign \new_[179]_  = \new_[44198]_  & \new_[44183]_ ;
  assign \new_[180]_  = \new_[44168]_  & \new_[44153]_ ;
  assign \new_[181]_  = \new_[44138]_  & \new_[44123]_ ;
  assign \new_[182]_  = \new_[44108]_  & \new_[44093]_ ;
  assign \new_[183]_  = \new_[44078]_  & \new_[44063]_ ;
  assign \new_[184]_  = \new_[44048]_  & \new_[44033]_ ;
  assign \new_[185]_  = \new_[44018]_  & \new_[44003]_ ;
  assign \new_[186]_  = \new_[43988]_  & \new_[43973]_ ;
  assign \new_[187]_  = \new_[43958]_  & \new_[43943]_ ;
  assign \new_[188]_  = \new_[43928]_  & \new_[43913]_ ;
  assign \new_[189]_  = \new_[43898]_  & \new_[43883]_ ;
  assign \new_[190]_  = \new_[43868]_  & \new_[43853]_ ;
  assign \new_[191]_  = \new_[43838]_  & \new_[43823]_ ;
  assign \new_[192]_  = \new_[43808]_  & \new_[43793]_ ;
  assign \new_[193]_  = \new_[43778]_  & \new_[43763]_ ;
  assign \new_[194]_  = \new_[43748]_  & \new_[43733]_ ;
  assign \new_[195]_  = \new_[43718]_  & \new_[43703]_ ;
  assign \new_[196]_  = \new_[43688]_  & \new_[43673]_ ;
  assign \new_[197]_  = \new_[43658]_  & \new_[43643]_ ;
  assign \new_[198]_  = \new_[43628]_  & \new_[43613]_ ;
  assign \new_[199]_  = \new_[43598]_  & \new_[43583]_ ;
  assign \new_[200]_  = \new_[43568]_  & \new_[43553]_ ;
  assign \new_[201]_  = \new_[43538]_  & \new_[43523]_ ;
  assign \new_[202]_  = \new_[43508]_  & \new_[43493]_ ;
  assign \new_[203]_  = \new_[43478]_  & \new_[43463]_ ;
  assign \new_[204]_  = \new_[43448]_  & \new_[43433]_ ;
  assign \new_[205]_  = \new_[43418]_  & \new_[43403]_ ;
  assign \new_[206]_  = \new_[43388]_  & \new_[43373]_ ;
  assign \new_[207]_  = \new_[43358]_  & \new_[43343]_ ;
  assign \new_[208]_  = \new_[43328]_  & \new_[43313]_ ;
  assign \new_[209]_  = \new_[43298]_  & \new_[43283]_ ;
  assign \new_[210]_  = \new_[43268]_  & \new_[43253]_ ;
  assign \new_[211]_  = \new_[43238]_  & \new_[43223]_ ;
  assign \new_[212]_  = \new_[43208]_  & \new_[43193]_ ;
  assign \new_[213]_  = \new_[43178]_  & \new_[43163]_ ;
  assign \new_[214]_  = \new_[43148]_  & \new_[43133]_ ;
  assign \new_[215]_  = \new_[43118]_  & \new_[43103]_ ;
  assign \new_[216]_  = \new_[43088]_  & \new_[43073]_ ;
  assign \new_[217]_  = \new_[43058]_  & \new_[43043]_ ;
  assign \new_[218]_  = \new_[43028]_  & \new_[43013]_ ;
  assign \new_[219]_  = \new_[42998]_  & \new_[42983]_ ;
  assign \new_[220]_  = \new_[42968]_  & \new_[42953]_ ;
  assign \new_[221]_  = \new_[42938]_  & \new_[42923]_ ;
  assign \new_[222]_  = \new_[42908]_  & \new_[42893]_ ;
  assign \new_[223]_  = \new_[42878]_  & \new_[42863]_ ;
  assign \new_[224]_  = \new_[42848]_  & \new_[42833]_ ;
  assign \new_[225]_  = \new_[42818]_  & \new_[42803]_ ;
  assign \new_[226]_  = \new_[42788]_  & \new_[42773]_ ;
  assign \new_[227]_  = \new_[42758]_  & \new_[42743]_ ;
  assign \new_[228]_  = \new_[42728]_  & \new_[42713]_ ;
  assign \new_[229]_  = \new_[42698]_  & \new_[42683]_ ;
  assign \new_[230]_  = \new_[42668]_  & \new_[42653]_ ;
  assign \new_[231]_  = \new_[42638]_  & \new_[42623]_ ;
  assign \new_[232]_  = \new_[42608]_  & \new_[42593]_ ;
  assign \new_[233]_  = \new_[42578]_  & \new_[42563]_ ;
  assign \new_[234]_  = \new_[42548]_  & \new_[42533]_ ;
  assign \new_[235]_  = \new_[42518]_  & \new_[42503]_ ;
  assign \new_[236]_  = \new_[42488]_  & \new_[42473]_ ;
  assign \new_[237]_  = \new_[42458]_  & \new_[42443]_ ;
  assign \new_[238]_  = \new_[42428]_  & \new_[42413]_ ;
  assign \new_[239]_  = \new_[42398]_  & \new_[42383]_ ;
  assign \new_[240]_  = \new_[42368]_  & \new_[42353]_ ;
  assign \new_[241]_  = \new_[42338]_  & \new_[42323]_ ;
  assign \new_[242]_  = \new_[42308]_  & \new_[42293]_ ;
  assign \new_[243]_  = \new_[42278]_  & \new_[42263]_ ;
  assign \new_[244]_  = \new_[42248]_  & \new_[42233]_ ;
  assign \new_[245]_  = \new_[42218]_  & \new_[42203]_ ;
  assign \new_[246]_  = \new_[42188]_  & \new_[42173]_ ;
  assign \new_[247]_  = \new_[42158]_  & \new_[42143]_ ;
  assign \new_[248]_  = \new_[42128]_  & \new_[42113]_ ;
  assign \new_[249]_  = \new_[42098]_  & \new_[42083]_ ;
  assign \new_[250]_  = \new_[42068]_  & \new_[42053]_ ;
  assign \new_[251]_  = \new_[42038]_  & \new_[42023]_ ;
  assign \new_[252]_  = \new_[42008]_  & \new_[41993]_ ;
  assign \new_[253]_  = \new_[41978]_  & \new_[41963]_ ;
  assign \new_[254]_  = \new_[41948]_  & \new_[41933]_ ;
  assign \new_[255]_  = \new_[41918]_  & \new_[41903]_ ;
  assign \new_[256]_  = \new_[41888]_  & \new_[41873]_ ;
  assign \new_[257]_  = \new_[41858]_  & \new_[41843]_ ;
  assign \new_[258]_  = \new_[41828]_  & \new_[41813]_ ;
  assign \new_[259]_  = \new_[41798]_  & \new_[41783]_ ;
  assign \new_[260]_  = \new_[41768]_  & \new_[41753]_ ;
  assign \new_[261]_  = \new_[41738]_  & \new_[41723]_ ;
  assign \new_[262]_  = \new_[41708]_  & \new_[41693]_ ;
  assign \new_[263]_  = \new_[41678]_  & \new_[41663]_ ;
  assign \new_[264]_  = \new_[41648]_  & \new_[41633]_ ;
  assign \new_[265]_  = \new_[41618]_  & \new_[41603]_ ;
  assign \new_[266]_  = \new_[41588]_  & \new_[41573]_ ;
  assign \new_[267]_  = \new_[41558]_  & \new_[41543]_ ;
  assign \new_[268]_  = \new_[41528]_  & \new_[41513]_ ;
  assign \new_[269]_  = \new_[41498]_  & \new_[41483]_ ;
  assign \new_[270]_  = \new_[41468]_  & \new_[41453]_ ;
  assign \new_[271]_  = \new_[41438]_  & \new_[41423]_ ;
  assign \new_[272]_  = \new_[41408]_  & \new_[41393]_ ;
  assign \new_[273]_  = \new_[41378]_  & \new_[41363]_ ;
  assign \new_[274]_  = \new_[41348]_  & \new_[41333]_ ;
  assign \new_[275]_  = \new_[41318]_  & \new_[41303]_ ;
  assign \new_[276]_  = \new_[41288]_  & \new_[41273]_ ;
  assign \new_[277]_  = \new_[41258]_  & \new_[41243]_ ;
  assign \new_[278]_  = \new_[41228]_  & \new_[41213]_ ;
  assign \new_[279]_  = \new_[41198]_  & \new_[41183]_ ;
  assign \new_[280]_  = \new_[41168]_  & \new_[41153]_ ;
  assign \new_[281]_  = \new_[41138]_  & \new_[41123]_ ;
  assign \new_[282]_  = \new_[41108]_  & \new_[41093]_ ;
  assign \new_[283]_  = \new_[41078]_  & \new_[41063]_ ;
  assign \new_[284]_  = \new_[41048]_  & \new_[41033]_ ;
  assign \new_[285]_  = \new_[41018]_  & \new_[41003]_ ;
  assign \new_[286]_  = \new_[40988]_  & \new_[40973]_ ;
  assign \new_[287]_  = \new_[40958]_  & \new_[40943]_ ;
  assign \new_[288]_  = \new_[40928]_  & \new_[40913]_ ;
  assign \new_[289]_  = \new_[40898]_  & \new_[40883]_ ;
  assign \new_[290]_  = \new_[40868]_  & \new_[40853]_ ;
  assign \new_[291]_  = \new_[40838]_  & \new_[40823]_ ;
  assign \new_[292]_  = \new_[40808]_  & \new_[40793]_ ;
  assign \new_[293]_  = \new_[40778]_  & \new_[40763]_ ;
  assign \new_[294]_  = \new_[40748]_  & \new_[40733]_ ;
  assign \new_[295]_  = \new_[40718]_  & \new_[40703]_ ;
  assign \new_[296]_  = \new_[40688]_  & \new_[40673]_ ;
  assign \new_[297]_  = \new_[40658]_  & \new_[40643]_ ;
  assign \new_[298]_  = \new_[40628]_  & \new_[40613]_ ;
  assign \new_[299]_  = \new_[40598]_  & \new_[40583]_ ;
  assign \new_[300]_  = \new_[40568]_  & \new_[40553]_ ;
  assign \new_[301]_  = \new_[40538]_  & \new_[40523]_ ;
  assign \new_[302]_  = \new_[40508]_  & \new_[40493]_ ;
  assign \new_[303]_  = \new_[40478]_  & \new_[40463]_ ;
  assign \new_[304]_  = \new_[40448]_  & \new_[40433]_ ;
  assign \new_[305]_  = \new_[40418]_  & \new_[40403]_ ;
  assign \new_[306]_  = \new_[40388]_  & \new_[40373]_ ;
  assign \new_[307]_  = \new_[40358]_  & \new_[40343]_ ;
  assign \new_[308]_  = \new_[40328]_  & \new_[40313]_ ;
  assign \new_[309]_  = \new_[40298]_  & \new_[40283]_ ;
  assign \new_[310]_  = \new_[40268]_  & \new_[40253]_ ;
  assign \new_[311]_  = \new_[40238]_  & \new_[40223]_ ;
  assign \new_[312]_  = \new_[40208]_  & \new_[40193]_ ;
  assign \new_[313]_  = \new_[40178]_  & \new_[40163]_ ;
  assign \new_[314]_  = \new_[40148]_  & \new_[40133]_ ;
  assign \new_[315]_  = \new_[40118]_  & \new_[40103]_ ;
  assign \new_[316]_  = \new_[40088]_  & \new_[40073]_ ;
  assign \new_[317]_  = \new_[40058]_  & \new_[40043]_ ;
  assign \new_[318]_  = \new_[40028]_  & \new_[40013]_ ;
  assign \new_[319]_  = \new_[39998]_  & \new_[39983]_ ;
  assign \new_[320]_  = \new_[39968]_  & \new_[39953]_ ;
  assign \new_[321]_  = \new_[39938]_  & \new_[39923]_ ;
  assign \new_[322]_  = \new_[39908]_  & \new_[39893]_ ;
  assign \new_[323]_  = \new_[39878]_  & \new_[39863]_ ;
  assign \new_[324]_  = \new_[39848]_  & \new_[39833]_ ;
  assign \new_[325]_  = \new_[39818]_  & \new_[39803]_ ;
  assign \new_[326]_  = \new_[39788]_  & \new_[39773]_ ;
  assign \new_[327]_  = \new_[39758]_  & \new_[39743]_ ;
  assign \new_[328]_  = \new_[39728]_  & \new_[39713]_ ;
  assign \new_[329]_  = \new_[39698]_  & \new_[39683]_ ;
  assign \new_[330]_  = \new_[39668]_  & \new_[39653]_ ;
  assign \new_[331]_  = \new_[39638]_  & \new_[39623]_ ;
  assign \new_[332]_  = \new_[39608]_  & \new_[39593]_ ;
  assign \new_[333]_  = \new_[39578]_  & \new_[39563]_ ;
  assign \new_[334]_  = \new_[39548]_  & \new_[39533]_ ;
  assign \new_[335]_  = \new_[39518]_  & \new_[39503]_ ;
  assign \new_[336]_  = \new_[39488]_  & \new_[39473]_ ;
  assign \new_[337]_  = \new_[39458]_  & \new_[39443]_ ;
  assign \new_[338]_  = \new_[39428]_  & \new_[39413]_ ;
  assign \new_[339]_  = \new_[39398]_  & \new_[39383]_ ;
  assign \new_[340]_  = \new_[39368]_  & \new_[39353]_ ;
  assign \new_[341]_  = \new_[39338]_  & \new_[39323]_ ;
  assign \new_[342]_  = \new_[39308]_  & \new_[39293]_ ;
  assign \new_[343]_  = \new_[39278]_  & \new_[39263]_ ;
  assign \new_[344]_  = \new_[39248]_  & \new_[39233]_ ;
  assign \new_[345]_  = \new_[39218]_  & \new_[39203]_ ;
  assign \new_[346]_  = \new_[39188]_  & \new_[39173]_ ;
  assign \new_[347]_  = \new_[39158]_  & \new_[39143]_ ;
  assign \new_[348]_  = \new_[39128]_  & \new_[39113]_ ;
  assign \new_[349]_  = \new_[39098]_  & \new_[39083]_ ;
  assign \new_[350]_  = \new_[39068]_  & \new_[39053]_ ;
  assign \new_[351]_  = \new_[39038]_  & \new_[39023]_ ;
  assign \new_[352]_  = \new_[39008]_  & \new_[38993]_ ;
  assign \new_[353]_  = \new_[38978]_  & \new_[38963]_ ;
  assign \new_[354]_  = \new_[38948]_  & \new_[38933]_ ;
  assign \new_[355]_  = \new_[38918]_  & \new_[38903]_ ;
  assign \new_[356]_  = \new_[38888]_  & \new_[38873]_ ;
  assign \new_[357]_  = \new_[38858]_  & \new_[38843]_ ;
  assign \new_[358]_  = \new_[38828]_  & \new_[38813]_ ;
  assign \new_[359]_  = \new_[38798]_  & \new_[38783]_ ;
  assign \new_[360]_  = \new_[38768]_  & \new_[38753]_ ;
  assign \new_[361]_  = \new_[38738]_  & \new_[38723]_ ;
  assign \new_[362]_  = \new_[38708]_  & \new_[38693]_ ;
  assign \new_[363]_  = \new_[38678]_  & \new_[38663]_ ;
  assign \new_[364]_  = \new_[38648]_  & \new_[38633]_ ;
  assign \new_[365]_  = \new_[38618]_  & \new_[38603]_ ;
  assign \new_[366]_  = \new_[38588]_  & \new_[38573]_ ;
  assign \new_[367]_  = \new_[38558]_  & \new_[38543]_ ;
  assign \new_[368]_  = \new_[38528]_  & \new_[38513]_ ;
  assign \new_[369]_  = \new_[38498]_  & \new_[38483]_ ;
  assign \new_[370]_  = \new_[38468]_  & \new_[38453]_ ;
  assign \new_[371]_  = \new_[38438]_  & \new_[38423]_ ;
  assign \new_[372]_  = \new_[38408]_  & \new_[38393]_ ;
  assign \new_[373]_  = \new_[38378]_  & \new_[38363]_ ;
  assign \new_[374]_  = \new_[38348]_  & \new_[38333]_ ;
  assign \new_[375]_  = \new_[38318]_  & \new_[38303]_ ;
  assign \new_[376]_  = \new_[38288]_  & \new_[38273]_ ;
  assign \new_[377]_  = \new_[38258]_  & \new_[38243]_ ;
  assign \new_[378]_  = \new_[38228]_  & \new_[38213]_ ;
  assign \new_[379]_  = \new_[38198]_  & \new_[38183]_ ;
  assign \new_[380]_  = \new_[38168]_  & \new_[38153]_ ;
  assign \new_[381]_  = \new_[38138]_  & \new_[38123]_ ;
  assign \new_[382]_  = \new_[38108]_  & \new_[38093]_ ;
  assign \new_[383]_  = \new_[38078]_  & \new_[38063]_ ;
  assign \new_[384]_  = \new_[38048]_  & \new_[38033]_ ;
  assign \new_[385]_  = \new_[38018]_  & \new_[38003]_ ;
  assign \new_[386]_  = \new_[37990]_  & \new_[37975]_ ;
  assign \new_[387]_  = \new_[37962]_  & \new_[37947]_ ;
  assign \new_[388]_  = \new_[37934]_  & \new_[37919]_ ;
  assign \new_[389]_  = \new_[37906]_  & \new_[37891]_ ;
  assign \new_[390]_  = \new_[37878]_  & \new_[37863]_ ;
  assign \new_[391]_  = \new_[37850]_  & \new_[37835]_ ;
  assign \new_[392]_  = \new_[37822]_  & \new_[37807]_ ;
  assign \new_[393]_  = \new_[37794]_  & \new_[37779]_ ;
  assign \new_[394]_  = \new_[37766]_  & \new_[37751]_ ;
  assign \new_[395]_  = \new_[37738]_  & \new_[37723]_ ;
  assign \new_[396]_  = \new_[37710]_  & \new_[37695]_ ;
  assign \new_[397]_  = \new_[37682]_  & \new_[37667]_ ;
  assign \new_[398]_  = \new_[37654]_  & \new_[37639]_ ;
  assign \new_[399]_  = \new_[37626]_  & \new_[37611]_ ;
  assign \new_[400]_  = \new_[37598]_  & \new_[37583]_ ;
  assign \new_[401]_  = \new_[37570]_  & \new_[37555]_ ;
  assign \new_[402]_  = \new_[37542]_  & \new_[37527]_ ;
  assign \new_[403]_  = \new_[37514]_  & \new_[37499]_ ;
  assign \new_[404]_  = \new_[37486]_  & \new_[37471]_ ;
  assign \new_[405]_  = \new_[37458]_  & \new_[37443]_ ;
  assign \new_[406]_  = \new_[37430]_  & \new_[37415]_ ;
  assign \new_[407]_  = \new_[37402]_  & \new_[37387]_ ;
  assign \new_[408]_  = \new_[37374]_  & \new_[37359]_ ;
  assign \new_[409]_  = \new_[37346]_  & \new_[37331]_ ;
  assign \new_[410]_  = \new_[37318]_  & \new_[37303]_ ;
  assign \new_[411]_  = \new_[37290]_  & \new_[37275]_ ;
  assign \new_[412]_  = \new_[37262]_  & \new_[37247]_ ;
  assign \new_[413]_  = \new_[37234]_  & \new_[37219]_ ;
  assign \new_[414]_  = \new_[37206]_  & \new_[37191]_ ;
  assign \new_[415]_  = \new_[37178]_  & \new_[37163]_ ;
  assign \new_[416]_  = \new_[37150]_  & \new_[37135]_ ;
  assign \new_[417]_  = \new_[37122]_  & \new_[37107]_ ;
  assign \new_[418]_  = \new_[37094]_  & \new_[37079]_ ;
  assign \new_[419]_  = \new_[37066]_  & \new_[37051]_ ;
  assign \new_[420]_  = \new_[37038]_  & \new_[37023]_ ;
  assign \new_[421]_  = \new_[37010]_  & \new_[36995]_ ;
  assign \new_[422]_  = \new_[36982]_  & \new_[36967]_ ;
  assign \new_[423]_  = \new_[36954]_  & \new_[36939]_ ;
  assign \new_[424]_  = \new_[36926]_  & \new_[36911]_ ;
  assign \new_[425]_  = \new_[36898]_  & \new_[36883]_ ;
  assign \new_[426]_  = \new_[36870]_  & \new_[36855]_ ;
  assign \new_[427]_  = \new_[36842]_  & \new_[36827]_ ;
  assign \new_[428]_  = \new_[36814]_  & \new_[36799]_ ;
  assign \new_[429]_  = \new_[36786]_  & \new_[36771]_ ;
  assign \new_[430]_  = \new_[36758]_  & \new_[36743]_ ;
  assign \new_[431]_  = \new_[36730]_  & \new_[36715]_ ;
  assign \new_[432]_  = \new_[36702]_  & \new_[36687]_ ;
  assign \new_[433]_  = \new_[36674]_  & \new_[36659]_ ;
  assign \new_[434]_  = \new_[36646]_  & \new_[36631]_ ;
  assign \new_[435]_  = \new_[36618]_  & \new_[36603]_ ;
  assign \new_[436]_  = \new_[36590]_  & \new_[36575]_ ;
  assign \new_[437]_  = \new_[36562]_  & \new_[36547]_ ;
  assign \new_[438]_  = \new_[36534]_  & \new_[36519]_ ;
  assign \new_[439]_  = \new_[36506]_  & \new_[36491]_ ;
  assign \new_[440]_  = \new_[36478]_  & \new_[36463]_ ;
  assign \new_[441]_  = \new_[36450]_  & \new_[36435]_ ;
  assign \new_[442]_  = \new_[36422]_  & \new_[36407]_ ;
  assign \new_[443]_  = \new_[36394]_  & \new_[36379]_ ;
  assign \new_[444]_  = \new_[36366]_  & \new_[36351]_ ;
  assign \new_[445]_  = \new_[36338]_  & \new_[36323]_ ;
  assign \new_[446]_  = \new_[36310]_  & \new_[36295]_ ;
  assign \new_[447]_  = \new_[36282]_  & \new_[36267]_ ;
  assign \new_[448]_  = \new_[36254]_  & \new_[36239]_ ;
  assign \new_[449]_  = \new_[36226]_  & \new_[36211]_ ;
  assign \new_[450]_  = \new_[36198]_  & \new_[36183]_ ;
  assign \new_[451]_  = \new_[36170]_  & \new_[36155]_ ;
  assign \new_[452]_  = \new_[36142]_  & \new_[36127]_ ;
  assign \new_[453]_  = \new_[36114]_  & \new_[36099]_ ;
  assign \new_[454]_  = \new_[36086]_  & \new_[36071]_ ;
  assign \new_[455]_  = \new_[36058]_  & \new_[36043]_ ;
  assign \new_[456]_  = \new_[36030]_  & \new_[36015]_ ;
  assign \new_[457]_  = \new_[36002]_  & \new_[35987]_ ;
  assign \new_[458]_  = \new_[35974]_  & \new_[35959]_ ;
  assign \new_[459]_  = \new_[35946]_  & \new_[35931]_ ;
  assign \new_[460]_  = \new_[35918]_  & \new_[35903]_ ;
  assign \new_[461]_  = \new_[35890]_  & \new_[35875]_ ;
  assign \new_[462]_  = \new_[35862]_  & \new_[35847]_ ;
  assign \new_[463]_  = \new_[35834]_  & \new_[35819]_ ;
  assign \new_[464]_  = \new_[35806]_  & \new_[35791]_ ;
  assign \new_[465]_  = \new_[35778]_  & \new_[35763]_ ;
  assign \new_[466]_  = \new_[35750]_  & \new_[35735]_ ;
  assign \new_[467]_  = \new_[35722]_  & \new_[35707]_ ;
  assign \new_[468]_  = \new_[35694]_  & \new_[35679]_ ;
  assign \new_[469]_  = \new_[35666]_  & \new_[35651]_ ;
  assign \new_[470]_  = \new_[35638]_  & \new_[35623]_ ;
  assign \new_[471]_  = \new_[35610]_  & \new_[35595]_ ;
  assign \new_[472]_  = \new_[35582]_  & \new_[35567]_ ;
  assign \new_[473]_  = \new_[35554]_  & \new_[35539]_ ;
  assign \new_[474]_  = \new_[35526]_  & \new_[35511]_ ;
  assign \new_[475]_  = \new_[35498]_  & \new_[35483]_ ;
  assign \new_[476]_  = \new_[35470]_  & \new_[35455]_ ;
  assign \new_[477]_  = \new_[35442]_  & \new_[35427]_ ;
  assign \new_[478]_  = \new_[35414]_  & \new_[35399]_ ;
  assign \new_[479]_  = \new_[35386]_  & \new_[35371]_ ;
  assign \new_[480]_  = \new_[35358]_  & \new_[35343]_ ;
  assign \new_[481]_  = \new_[35330]_  & \new_[35315]_ ;
  assign \new_[482]_  = \new_[35302]_  & \new_[35287]_ ;
  assign \new_[483]_  = \new_[35274]_  & \new_[35259]_ ;
  assign \new_[484]_  = \new_[35246]_  & \new_[35231]_ ;
  assign \new_[485]_  = \new_[35218]_  & \new_[35203]_ ;
  assign \new_[486]_  = \new_[35190]_  & \new_[35175]_ ;
  assign \new_[487]_  = \new_[35162]_  & \new_[35147]_ ;
  assign \new_[488]_  = \new_[35134]_  & \new_[35119]_ ;
  assign \new_[489]_  = \new_[35106]_  & \new_[35091]_ ;
  assign \new_[490]_  = \new_[35078]_  & \new_[35063]_ ;
  assign \new_[491]_  = \new_[35050]_  & \new_[35035]_ ;
  assign \new_[492]_  = \new_[35022]_  & \new_[35007]_ ;
  assign \new_[493]_  = \new_[34994]_  & \new_[34979]_ ;
  assign \new_[494]_  = \new_[34966]_  & \new_[34951]_ ;
  assign \new_[495]_  = \new_[34938]_  & \new_[34923]_ ;
  assign \new_[496]_  = \new_[34910]_  & \new_[34895]_ ;
  assign \new_[497]_  = \new_[34882]_  & \new_[34867]_ ;
  assign \new_[498]_  = \new_[34854]_  & \new_[34839]_ ;
  assign \new_[499]_  = \new_[34826]_  & \new_[34811]_ ;
  assign \new_[500]_  = \new_[34798]_  & \new_[34783]_ ;
  assign \new_[501]_  = \new_[34770]_  & \new_[34755]_ ;
  assign \new_[502]_  = \new_[34742]_  & \new_[34727]_ ;
  assign \new_[503]_  = \new_[34714]_  & \new_[34699]_ ;
  assign \new_[504]_  = \new_[34686]_  & \new_[34671]_ ;
  assign \new_[505]_  = \new_[34658]_  & \new_[34643]_ ;
  assign \new_[506]_  = \new_[34630]_  & \new_[34615]_ ;
  assign \new_[507]_  = \new_[34602]_  & \new_[34587]_ ;
  assign \new_[508]_  = \new_[34574]_  & \new_[34559]_ ;
  assign \new_[509]_  = \new_[34546]_  & \new_[34531]_ ;
  assign \new_[510]_  = \new_[34518]_  & \new_[34503]_ ;
  assign \new_[511]_  = \new_[34490]_  & \new_[34475]_ ;
  assign \new_[512]_  = \new_[34462]_  & \new_[34447]_ ;
  assign \new_[513]_  = \new_[34434]_  & \new_[34421]_ ;
  assign \new_[514]_  = \new_[34408]_  & \new_[34395]_ ;
  assign \new_[515]_  = \new_[34382]_  & \new_[34369]_ ;
  assign \new_[516]_  = \new_[34356]_  & \new_[34343]_ ;
  assign \new_[517]_  = \new_[34330]_  & \new_[34317]_ ;
  assign \new_[518]_  = \new_[34304]_  & \new_[34291]_ ;
  assign \new_[519]_  = \new_[34278]_  & \new_[34265]_ ;
  assign \new_[520]_  = \new_[34252]_  & \new_[34239]_ ;
  assign \new_[521]_  = \new_[34226]_  & \new_[34213]_ ;
  assign \new_[522]_  = \new_[34200]_  & \new_[34187]_ ;
  assign \new_[523]_  = \new_[34174]_  & \new_[34161]_ ;
  assign \new_[524]_  = \new_[34148]_  & \new_[34135]_ ;
  assign \new_[525]_  = \new_[34122]_  & \new_[34109]_ ;
  assign \new_[526]_  = \new_[34096]_  & \new_[34083]_ ;
  assign \new_[527]_  = \new_[34070]_  & \new_[34057]_ ;
  assign \new_[528]_  = \new_[34044]_  & \new_[34031]_ ;
  assign \new_[529]_  = \new_[34018]_  & \new_[34005]_ ;
  assign \new_[530]_  = \new_[33992]_  & \new_[33979]_ ;
  assign \new_[531]_  = \new_[33966]_  & \new_[33953]_ ;
  assign \new_[532]_  = \new_[33940]_  & \new_[33927]_ ;
  assign \new_[533]_  = \new_[33914]_  & \new_[33901]_ ;
  assign \new_[534]_  = \new_[33888]_  & \new_[33875]_ ;
  assign \new_[535]_  = \new_[33862]_  & \new_[33849]_ ;
  assign \new_[536]_  = \new_[33836]_  & \new_[33823]_ ;
  assign \new_[537]_  = \new_[33810]_  & \new_[33797]_ ;
  assign \new_[538]_  = \new_[33784]_  & \new_[33771]_ ;
  assign \new_[539]_  = \new_[33758]_  & \new_[33745]_ ;
  assign \new_[540]_  = \new_[33732]_  & \new_[33719]_ ;
  assign \new_[541]_  = \new_[33706]_  & \new_[33693]_ ;
  assign \new_[542]_  = \new_[33680]_  & \new_[33667]_ ;
  assign \new_[543]_  = \new_[33654]_  & \new_[33641]_ ;
  assign \new_[544]_  = \new_[33628]_  & \new_[33615]_ ;
  assign \new_[545]_  = \new_[33602]_  & \new_[33589]_ ;
  assign \new_[546]_  = \new_[33576]_  & \new_[33563]_ ;
  assign \new_[547]_  = \new_[33550]_  & \new_[33537]_ ;
  assign \new_[548]_  = \new_[33524]_  & \new_[33511]_ ;
  assign \new_[549]_  = \new_[33498]_  & \new_[33485]_ ;
  assign \new_[550]_  = \new_[33472]_  & \new_[33459]_ ;
  assign \new_[551]_  = \new_[33446]_  & \new_[33433]_ ;
  assign \new_[552]_  = \new_[33420]_  & \new_[33407]_ ;
  assign \new_[553]_  = \new_[33394]_  & \new_[33381]_ ;
  assign \new_[554]_  = \new_[33368]_  & \new_[33355]_ ;
  assign \new_[555]_  = \new_[33342]_  & \new_[33329]_ ;
  assign \new_[556]_  = \new_[33316]_  & \new_[33303]_ ;
  assign \new_[557]_  = \new_[33290]_  & \new_[33277]_ ;
  assign \new_[558]_  = \new_[33264]_  & \new_[33251]_ ;
  assign \new_[559]_  = \new_[33238]_  & \new_[33225]_ ;
  assign \new_[560]_  = \new_[33212]_  & \new_[33199]_ ;
  assign \new_[561]_  = \new_[33186]_  & \new_[33173]_ ;
  assign \new_[562]_  = \new_[33160]_  & \new_[33147]_ ;
  assign \new_[563]_  = \new_[33134]_  & \new_[33121]_ ;
  assign \new_[564]_  = \new_[33108]_  & \new_[33095]_ ;
  assign \new_[565]_  = \new_[33082]_  & \new_[33069]_ ;
  assign \new_[566]_  = \new_[33056]_  & \new_[33043]_ ;
  assign \new_[567]_  = \new_[33030]_  & \new_[33017]_ ;
  assign \new_[568]_  = \new_[33004]_  & \new_[32991]_ ;
  assign \new_[569]_  = \new_[32978]_  & \new_[32965]_ ;
  assign \new_[570]_  = \new_[32952]_  & \new_[32939]_ ;
  assign \new_[571]_  = \new_[32926]_  & \new_[32913]_ ;
  assign \new_[572]_  = \new_[32900]_  & \new_[32887]_ ;
  assign \new_[573]_  = \new_[32874]_  & \new_[32861]_ ;
  assign \new_[574]_  = \new_[32848]_  & \new_[32835]_ ;
  assign \new_[575]_  = \new_[32822]_  & \new_[32809]_ ;
  assign \new_[576]_  = \new_[32796]_  & \new_[32783]_ ;
  assign \new_[577]_  = \new_[32770]_  & \new_[32757]_ ;
  assign \new_[578]_  = \new_[32744]_  & \new_[32731]_ ;
  assign \new_[579]_  = \new_[32718]_  & \new_[32705]_ ;
  assign \new_[580]_  = \new_[32692]_  & \new_[32679]_ ;
  assign \new_[581]_  = \new_[32666]_  & \new_[32653]_ ;
  assign \new_[582]_  = \new_[32640]_  & \new_[32627]_ ;
  assign \new_[583]_  = \new_[32614]_  & \new_[32601]_ ;
  assign \new_[584]_  = \new_[32588]_  & \new_[32575]_ ;
  assign \new_[585]_  = \new_[32562]_  & \new_[32549]_ ;
  assign \new_[586]_  = \new_[32536]_  & \new_[32523]_ ;
  assign \new_[587]_  = \new_[32510]_  & \new_[32497]_ ;
  assign \new_[588]_  = \new_[32484]_  & \new_[32471]_ ;
  assign \new_[589]_  = \new_[32458]_  & \new_[32445]_ ;
  assign \new_[590]_  = \new_[32432]_  & \new_[32419]_ ;
  assign \new_[591]_  = \new_[32406]_  & \new_[32393]_ ;
  assign \new_[592]_  = \new_[32380]_  & \new_[32367]_ ;
  assign \new_[593]_  = \new_[32354]_  & \new_[32341]_ ;
  assign \new_[594]_  = \new_[32328]_  & \new_[32315]_ ;
  assign \new_[595]_  = \new_[32302]_  & \new_[32289]_ ;
  assign \new_[596]_  = \new_[32276]_  & \new_[32263]_ ;
  assign \new_[597]_  = \new_[32250]_  & \new_[32237]_ ;
  assign \new_[598]_  = \new_[32224]_  & \new_[32211]_ ;
  assign \new_[599]_  = \new_[32198]_  & \new_[32185]_ ;
  assign \new_[600]_  = \new_[32172]_  & \new_[32159]_ ;
  assign \new_[601]_  = \new_[32146]_  & \new_[32133]_ ;
  assign \new_[602]_  = \new_[32120]_  & \new_[32107]_ ;
  assign \new_[603]_  = \new_[32094]_  & \new_[32081]_ ;
  assign \new_[604]_  = \new_[32068]_  & \new_[32055]_ ;
  assign \new_[605]_  = \new_[32042]_  & \new_[32029]_ ;
  assign \new_[606]_  = \new_[32016]_  & \new_[32003]_ ;
  assign \new_[607]_  = \new_[31990]_  & \new_[31977]_ ;
  assign \new_[608]_  = \new_[31964]_  & \new_[31951]_ ;
  assign \new_[609]_  = \new_[31938]_  & \new_[31925]_ ;
  assign \new_[610]_  = \new_[31912]_  & \new_[31899]_ ;
  assign \new_[611]_  = \new_[31886]_  & \new_[31873]_ ;
  assign \new_[612]_  = \new_[31860]_  & \new_[31847]_ ;
  assign \new_[613]_  = \new_[31834]_  & \new_[31821]_ ;
  assign \new_[614]_  = \new_[31808]_  & \new_[31795]_ ;
  assign \new_[615]_  = \new_[31782]_  & \new_[31769]_ ;
  assign \new_[616]_  = \new_[31756]_  & \new_[31743]_ ;
  assign \new_[617]_  = \new_[31730]_  & \new_[31717]_ ;
  assign \new_[618]_  = \new_[31704]_  & \new_[31691]_ ;
  assign \new_[619]_  = \new_[31678]_  & \new_[31665]_ ;
  assign \new_[620]_  = \new_[31652]_  & \new_[31639]_ ;
  assign \new_[621]_  = \new_[31626]_  & \new_[31613]_ ;
  assign \new_[622]_  = \new_[31600]_  & \new_[31587]_ ;
  assign \new_[623]_  = \new_[31574]_  & \new_[31561]_ ;
  assign \new_[624]_  = \new_[31548]_  & \new_[31535]_ ;
  assign \new_[625]_  = \new_[31522]_  & \new_[31509]_ ;
  assign \new_[626]_  = \new_[31496]_  & \new_[31483]_ ;
  assign \new_[627]_  = \new_[31470]_  & \new_[31457]_ ;
  assign \new_[628]_  = \new_[31444]_  & \new_[31431]_ ;
  assign \new_[629]_  = \new_[31418]_  & \new_[31405]_ ;
  assign \new_[630]_  = \new_[31392]_  & \new_[31379]_ ;
  assign \new_[631]_  = \new_[31366]_  & \new_[31353]_ ;
  assign \new_[632]_  = \new_[31340]_  & \new_[31327]_ ;
  assign \new_[633]_  = \new_[31314]_  & \new_[31301]_ ;
  assign \new_[634]_  = \new_[31288]_  & \new_[31275]_ ;
  assign \new_[635]_  = \new_[31262]_  & \new_[31249]_ ;
  assign \new_[636]_  = \new_[31236]_  & \new_[31223]_ ;
  assign \new_[637]_  = \new_[31210]_  & \new_[31197]_ ;
  assign \new_[638]_  = \new_[31184]_  & \new_[31171]_ ;
  assign \new_[639]_  = \new_[31158]_  & \new_[31145]_ ;
  assign \new_[640]_  = \new_[31132]_  & \new_[31119]_ ;
  assign \new_[641]_  = \new_[31106]_  & \new_[31093]_ ;
  assign \new_[642]_  = \new_[31080]_  & \new_[31067]_ ;
  assign \new_[643]_  = \new_[31054]_  & \new_[31041]_ ;
  assign \new_[644]_  = \new_[31028]_  & \new_[31015]_ ;
  assign \new_[645]_  = \new_[31002]_  & \new_[30989]_ ;
  assign \new_[646]_  = \new_[30976]_  & \new_[30963]_ ;
  assign \new_[647]_  = \new_[30950]_  & \new_[30937]_ ;
  assign \new_[648]_  = \new_[30924]_  & \new_[30911]_ ;
  assign \new_[649]_  = \new_[30898]_  & \new_[30885]_ ;
  assign \new_[650]_  = \new_[30872]_  & \new_[30859]_ ;
  assign \new_[651]_  = \new_[30846]_  & \new_[30833]_ ;
  assign \new_[652]_  = \new_[30820]_  & \new_[30807]_ ;
  assign \new_[653]_  = \new_[30794]_  & \new_[30781]_ ;
  assign \new_[654]_  = \new_[30768]_  & \new_[30755]_ ;
  assign \new_[655]_  = \new_[30742]_  & \new_[30729]_ ;
  assign \new_[656]_  = \new_[30716]_  & \new_[30703]_ ;
  assign \new_[657]_  = \new_[30690]_  & \new_[30677]_ ;
  assign \new_[658]_  = \new_[30664]_  & \new_[30651]_ ;
  assign \new_[659]_  = \new_[30638]_  & \new_[30625]_ ;
  assign \new_[660]_  = \new_[30612]_  & \new_[30599]_ ;
  assign \new_[661]_  = \new_[30586]_  & \new_[30573]_ ;
  assign \new_[662]_  = \new_[30560]_  & \new_[30547]_ ;
  assign \new_[663]_  = \new_[30534]_  & \new_[30521]_ ;
  assign \new_[664]_  = \new_[30508]_  & \new_[30495]_ ;
  assign \new_[665]_  = \new_[30482]_  & \new_[30469]_ ;
  assign \new_[666]_  = \new_[30456]_  & \new_[30443]_ ;
  assign \new_[667]_  = \new_[30430]_  & \new_[30417]_ ;
  assign \new_[668]_  = \new_[30404]_  & \new_[30391]_ ;
  assign \new_[669]_  = \new_[30378]_  & \new_[30365]_ ;
  assign \new_[670]_  = \new_[30352]_  & \new_[30339]_ ;
  assign \new_[671]_  = \new_[30326]_  & \new_[30313]_ ;
  assign \new_[672]_  = \new_[30300]_  & \new_[30287]_ ;
  assign \new_[673]_  = \new_[30274]_  & \new_[30261]_ ;
  assign \new_[674]_  = \new_[30248]_  & \new_[30235]_ ;
  assign \new_[675]_  = \new_[30222]_  & \new_[30209]_ ;
  assign \new_[676]_  = \new_[30196]_  & \new_[30183]_ ;
  assign \new_[677]_  = \new_[30170]_  & \new_[30157]_ ;
  assign \new_[678]_  = \new_[30144]_  & \new_[30131]_ ;
  assign \new_[679]_  = \new_[30118]_  & \new_[30105]_ ;
  assign \new_[680]_  = \new_[30092]_  & \new_[30079]_ ;
  assign \new_[681]_  = \new_[30066]_  & \new_[30053]_ ;
  assign \new_[682]_  = \new_[30040]_  & \new_[30027]_ ;
  assign \new_[683]_  = \new_[30014]_  & \new_[30001]_ ;
  assign \new_[684]_  = \new_[29988]_  & \new_[29975]_ ;
  assign \new_[685]_  = \new_[29962]_  & \new_[29949]_ ;
  assign \new_[686]_  = \new_[29936]_  & \new_[29923]_ ;
  assign \new_[687]_  = \new_[29910]_  & \new_[29897]_ ;
  assign \new_[688]_  = \new_[29884]_  & \new_[29871]_ ;
  assign \new_[689]_  = \new_[29858]_  & \new_[29845]_ ;
  assign \new_[690]_  = \new_[29832]_  & \new_[29819]_ ;
  assign \new_[691]_  = \new_[29806]_  & \new_[29793]_ ;
  assign \new_[692]_  = \new_[29780]_  & \new_[29767]_ ;
  assign \new_[693]_  = \new_[29754]_  & \new_[29741]_ ;
  assign \new_[694]_  = \new_[29728]_  & \new_[29715]_ ;
  assign \new_[695]_  = \new_[29702]_  & \new_[29689]_ ;
  assign \new_[696]_  = \new_[29676]_  & \new_[29663]_ ;
  assign \new_[697]_  = \new_[29650]_  & \new_[29637]_ ;
  assign \new_[698]_  = \new_[29624]_  & \new_[29611]_ ;
  assign \new_[699]_  = \new_[29598]_  & \new_[29585]_ ;
  assign \new_[700]_  = \new_[29572]_  & \new_[29559]_ ;
  assign \new_[701]_  = \new_[29546]_  & \new_[29533]_ ;
  assign \new_[702]_  = \new_[29520]_  & \new_[29507]_ ;
  assign \new_[703]_  = \new_[29494]_  & \new_[29481]_ ;
  assign \new_[704]_  = \new_[29468]_  & \new_[29455]_ ;
  assign \new_[705]_  = \new_[29442]_  & \new_[29429]_ ;
  assign \new_[706]_  = \new_[29416]_  & \new_[29403]_ ;
  assign \new_[707]_  = \new_[29390]_  & \new_[29377]_ ;
  assign \new_[708]_  = \new_[29364]_  & \new_[29351]_ ;
  assign \new_[709]_  = \new_[29338]_  & \new_[29325]_ ;
  assign \new_[710]_  = \new_[29312]_  & \new_[29299]_ ;
  assign \new_[711]_  = \new_[29286]_  & \new_[29273]_ ;
  assign \new_[712]_  = \new_[29260]_  & \new_[29247]_ ;
  assign \new_[713]_  = \new_[29234]_  & \new_[29221]_ ;
  assign \new_[714]_  = \new_[29208]_  & \new_[29195]_ ;
  assign \new_[715]_  = \new_[29182]_  & \new_[29169]_ ;
  assign \new_[716]_  = \new_[29156]_  & \new_[29143]_ ;
  assign \new_[717]_  = \new_[29130]_  & \new_[29117]_ ;
  assign \new_[718]_  = \new_[29104]_  & \new_[29091]_ ;
  assign \new_[719]_  = \new_[29078]_  & \new_[29065]_ ;
  assign \new_[720]_  = \new_[29052]_  & \new_[29039]_ ;
  assign \new_[721]_  = \new_[29026]_  & \new_[29013]_ ;
  assign \new_[722]_  = \new_[29000]_  & \new_[28987]_ ;
  assign \new_[723]_  = \new_[28974]_  & \new_[28961]_ ;
  assign \new_[724]_  = \new_[28948]_  & \new_[28935]_ ;
  assign \new_[725]_  = \new_[28922]_  & \new_[28909]_ ;
  assign \new_[726]_  = \new_[28896]_  & \new_[28883]_ ;
  assign \new_[727]_  = \new_[28870]_  & \new_[28857]_ ;
  assign \new_[728]_  = \new_[28844]_  & \new_[28831]_ ;
  assign \new_[729]_  = \new_[28818]_  & \new_[28805]_ ;
  assign \new_[730]_  = \new_[28792]_  & \new_[28779]_ ;
  assign \new_[731]_  = \new_[28766]_  & \new_[28753]_ ;
  assign \new_[732]_  = \new_[28740]_  & \new_[28727]_ ;
  assign \new_[733]_  = \new_[28714]_  & \new_[28701]_ ;
  assign \new_[734]_  = \new_[28688]_  & \new_[28675]_ ;
  assign \new_[735]_  = \new_[28662]_  & \new_[28649]_ ;
  assign \new_[736]_  = \new_[28636]_  & \new_[28623]_ ;
  assign \new_[737]_  = \new_[28610]_  & \new_[28597]_ ;
  assign \new_[738]_  = \new_[28584]_  & \new_[28571]_ ;
  assign \new_[739]_  = \new_[28558]_  & \new_[28545]_ ;
  assign \new_[740]_  = \new_[28532]_  & \new_[28519]_ ;
  assign \new_[741]_  = \new_[28506]_  & \new_[28493]_ ;
  assign \new_[742]_  = \new_[28480]_  & \new_[28467]_ ;
  assign \new_[743]_  = \new_[28454]_  & \new_[28441]_ ;
  assign \new_[744]_  = \new_[28428]_  & \new_[28415]_ ;
  assign \new_[745]_  = \new_[28402]_  & \new_[28389]_ ;
  assign \new_[746]_  = \new_[28376]_  & \new_[28363]_ ;
  assign \new_[747]_  = \new_[28350]_  & \new_[28337]_ ;
  assign \new_[748]_  = \new_[28324]_  & \new_[28311]_ ;
  assign \new_[749]_  = \new_[28298]_  & \new_[28285]_ ;
  assign \new_[750]_  = \new_[28272]_  & \new_[28259]_ ;
  assign \new_[751]_  = \new_[28246]_  & \new_[28233]_ ;
  assign \new_[752]_  = \new_[28220]_  & \new_[28207]_ ;
  assign \new_[753]_  = \new_[28194]_  & \new_[28181]_ ;
  assign \new_[754]_  = \new_[28168]_  & \new_[28155]_ ;
  assign \new_[755]_  = \new_[28142]_  & \new_[28129]_ ;
  assign \new_[756]_  = \new_[28116]_  & \new_[28103]_ ;
  assign \new_[757]_  = \new_[28090]_  & \new_[28077]_ ;
  assign \new_[758]_  = \new_[28064]_  & \new_[28051]_ ;
  assign \new_[759]_  = \new_[28038]_  & \new_[28025]_ ;
  assign \new_[760]_  = \new_[28012]_  & \new_[27999]_ ;
  assign \new_[761]_  = \new_[27986]_  & \new_[27973]_ ;
  assign \new_[762]_  = \new_[27960]_  & \new_[27947]_ ;
  assign \new_[763]_  = \new_[27934]_  & \new_[27921]_ ;
  assign \new_[764]_  = \new_[27908]_  & \new_[27895]_ ;
  assign \new_[765]_  = \new_[27882]_  & \new_[27869]_ ;
  assign \new_[766]_  = \new_[27856]_  & \new_[27843]_ ;
  assign \new_[767]_  = \new_[27830]_  & \new_[27817]_ ;
  assign \new_[768]_  = \new_[27804]_  & \new_[27791]_ ;
  assign \new_[769]_  = \new_[27778]_  & \new_[27765]_ ;
  assign \new_[770]_  = \new_[27752]_  & \new_[27739]_ ;
  assign \new_[771]_  = \new_[27726]_  & \new_[27713]_ ;
  assign \new_[772]_  = \new_[27700]_  & \new_[27687]_ ;
  assign \new_[773]_  = \new_[27674]_  & \new_[27661]_ ;
  assign \new_[774]_  = \new_[27648]_  & \new_[27635]_ ;
  assign \new_[775]_  = \new_[27622]_  & \new_[27609]_ ;
  assign \new_[776]_  = \new_[27596]_  & \new_[27583]_ ;
  assign \new_[777]_  = \new_[27570]_  & \new_[27557]_ ;
  assign \new_[778]_  = \new_[27544]_  & \new_[27531]_ ;
  assign \new_[779]_  = \new_[27518]_  & \new_[27505]_ ;
  assign \new_[780]_  = \new_[27492]_  & \new_[27479]_ ;
  assign \new_[781]_  = \new_[27466]_  & \new_[27453]_ ;
  assign \new_[782]_  = \new_[27440]_  & \new_[27427]_ ;
  assign \new_[783]_  = \new_[27414]_  & \new_[27401]_ ;
  assign \new_[784]_  = \new_[27388]_  & \new_[27375]_ ;
  assign \new_[785]_  = \new_[27362]_  & \new_[27349]_ ;
  assign \new_[786]_  = \new_[27336]_  & \new_[27323]_ ;
  assign \new_[787]_  = \new_[27310]_  & \new_[27297]_ ;
  assign \new_[788]_  = \new_[27284]_  & \new_[27271]_ ;
  assign \new_[789]_  = \new_[27258]_  & \new_[27245]_ ;
  assign \new_[790]_  = \new_[27232]_  & \new_[27219]_ ;
  assign \new_[791]_  = \new_[27206]_  & \new_[27193]_ ;
  assign \new_[792]_  = \new_[27180]_  & \new_[27167]_ ;
  assign \new_[793]_  = \new_[27154]_  & \new_[27141]_ ;
  assign \new_[794]_  = \new_[27128]_  & \new_[27115]_ ;
  assign \new_[795]_  = \new_[27102]_  & \new_[27089]_ ;
  assign \new_[796]_  = \new_[27076]_  & \new_[27063]_ ;
  assign \new_[797]_  = \new_[27050]_  & \new_[27037]_ ;
  assign \new_[798]_  = \new_[27024]_  & \new_[27011]_ ;
  assign \new_[799]_  = \new_[26998]_  & \new_[26985]_ ;
  assign \new_[800]_  = \new_[26972]_  & \new_[26959]_ ;
  assign \new_[801]_  = \new_[26946]_  & \new_[26933]_ ;
  assign \new_[802]_  = \new_[26920]_  & \new_[26907]_ ;
  assign \new_[803]_  = \new_[26894]_  & \new_[26881]_ ;
  assign \new_[804]_  = \new_[26868]_  & \new_[26855]_ ;
  assign \new_[805]_  = \new_[26842]_  & \new_[26829]_ ;
  assign \new_[806]_  = \new_[26816]_  & \new_[26803]_ ;
  assign \new_[807]_  = \new_[26790]_  & \new_[26777]_ ;
  assign \new_[808]_  = \new_[26764]_  & \new_[26751]_ ;
  assign \new_[809]_  = \new_[26738]_  & \new_[26725]_ ;
  assign \new_[810]_  = \new_[26712]_  & \new_[26699]_ ;
  assign \new_[811]_  = \new_[26686]_  & \new_[26673]_ ;
  assign \new_[812]_  = \new_[26660]_  & \new_[26647]_ ;
  assign \new_[813]_  = \new_[26634]_  & \new_[26621]_ ;
  assign \new_[814]_  = \new_[26608]_  & \new_[26595]_ ;
  assign \new_[815]_  = \new_[26582]_  & \new_[26569]_ ;
  assign \new_[816]_  = \new_[26556]_  & \new_[26543]_ ;
  assign \new_[817]_  = \new_[26530]_  & \new_[26517]_ ;
  assign \new_[818]_  = \new_[26504]_  & \new_[26491]_ ;
  assign \new_[819]_  = \new_[26478]_  & \new_[26465]_ ;
  assign \new_[820]_  = \new_[26452]_  & \new_[26439]_ ;
  assign \new_[821]_  = \new_[26426]_  & \new_[26413]_ ;
  assign \new_[822]_  = \new_[26400]_  & \new_[26387]_ ;
  assign \new_[823]_  = \new_[26374]_  & \new_[26361]_ ;
  assign \new_[824]_  = \new_[26348]_  & \new_[26335]_ ;
  assign \new_[825]_  = \new_[26322]_  & \new_[26309]_ ;
  assign \new_[826]_  = \new_[26296]_  & \new_[26283]_ ;
  assign \new_[827]_  = \new_[26270]_  & \new_[26257]_ ;
  assign \new_[828]_  = \new_[26244]_  & \new_[26231]_ ;
  assign \new_[829]_  = \new_[26218]_  & \new_[26205]_ ;
  assign \new_[830]_  = \new_[26192]_  & \new_[26179]_ ;
  assign \new_[831]_  = \new_[26166]_  & \new_[26153]_ ;
  assign \new_[832]_  = \new_[26140]_  & \new_[26127]_ ;
  assign \new_[833]_  = \new_[26114]_  & \new_[26101]_ ;
  assign \new_[834]_  = \new_[26088]_  & \new_[26075]_ ;
  assign \new_[835]_  = \new_[26062]_  & \new_[26049]_ ;
  assign \new_[836]_  = \new_[26036]_  & \new_[26023]_ ;
  assign \new_[837]_  = \new_[26010]_  & \new_[25997]_ ;
  assign \new_[838]_  = \new_[25984]_  & \new_[25971]_ ;
  assign \new_[839]_  = \new_[25958]_  & \new_[25945]_ ;
  assign \new_[840]_  = \new_[25932]_  & \new_[25919]_ ;
  assign \new_[841]_  = \new_[25906]_  & \new_[25893]_ ;
  assign \new_[842]_  = \new_[25880]_  & \new_[25867]_ ;
  assign \new_[843]_  = \new_[25854]_  & \new_[25841]_ ;
  assign \new_[844]_  = \new_[25828]_  & \new_[25815]_ ;
  assign \new_[845]_  = \new_[25802]_  & \new_[25789]_ ;
  assign \new_[846]_  = \new_[25776]_  & \new_[25763]_ ;
  assign \new_[847]_  = \new_[25750]_  & \new_[25737]_ ;
  assign \new_[848]_  = \new_[25724]_  & \new_[25711]_ ;
  assign \new_[849]_  = \new_[25698]_  & \new_[25685]_ ;
  assign \new_[850]_  = \new_[25672]_  & \new_[25659]_ ;
  assign \new_[851]_  = \new_[25646]_  & \new_[25633]_ ;
  assign \new_[852]_  = \new_[25620]_  & \new_[25607]_ ;
  assign \new_[853]_  = \new_[25594]_  & \new_[25581]_ ;
  assign \new_[854]_  = \new_[25568]_  & \new_[25555]_ ;
  assign \new_[855]_  = \new_[25542]_  & \new_[25529]_ ;
  assign \new_[856]_  = \new_[25516]_  & \new_[25503]_ ;
  assign \new_[857]_  = \new_[25490]_  & \new_[25477]_ ;
  assign \new_[858]_  = \new_[25464]_  & \new_[25451]_ ;
  assign \new_[859]_  = \new_[25438]_  & \new_[25425]_ ;
  assign \new_[860]_  = \new_[25412]_  & \new_[25399]_ ;
  assign \new_[861]_  = \new_[25386]_  & \new_[25373]_ ;
  assign \new_[862]_  = \new_[25360]_  & \new_[25347]_ ;
  assign \new_[863]_  = \new_[25334]_  & \new_[25321]_ ;
  assign \new_[864]_  = \new_[25308]_  & \new_[25295]_ ;
  assign \new_[865]_  = \new_[25282]_  & \new_[25269]_ ;
  assign \new_[866]_  = \new_[25256]_  & \new_[25243]_ ;
  assign \new_[867]_  = \new_[25230]_  & \new_[25217]_ ;
  assign \new_[868]_  = \new_[25204]_  & \new_[25191]_ ;
  assign \new_[869]_  = \new_[25178]_  & \new_[25165]_ ;
  assign \new_[870]_  = \new_[25152]_  & \new_[25139]_ ;
  assign \new_[871]_  = \new_[25126]_  & \new_[25113]_ ;
  assign \new_[872]_  = \new_[25100]_  & \new_[25087]_ ;
  assign \new_[873]_  = \new_[25074]_  & \new_[25061]_ ;
  assign \new_[874]_  = \new_[25048]_  & \new_[25035]_ ;
  assign \new_[875]_  = \new_[25022]_  & \new_[25009]_ ;
  assign \new_[876]_  = \new_[24996]_  & \new_[24983]_ ;
  assign \new_[877]_  = \new_[24970]_  & \new_[24957]_ ;
  assign \new_[878]_  = \new_[24944]_  & \new_[24931]_ ;
  assign \new_[879]_  = \new_[24918]_  & \new_[24905]_ ;
  assign \new_[880]_  = \new_[24892]_  & \new_[24879]_ ;
  assign \new_[881]_  = \new_[24866]_  & \new_[24853]_ ;
  assign \new_[882]_  = \new_[24840]_  & \new_[24827]_ ;
  assign \new_[883]_  = \new_[24814]_  & \new_[24801]_ ;
  assign \new_[884]_  = \new_[24788]_  & \new_[24775]_ ;
  assign \new_[885]_  = \new_[24762]_  & \new_[24749]_ ;
  assign \new_[886]_  = \new_[24736]_  & \new_[24723]_ ;
  assign \new_[887]_  = \new_[24710]_  & \new_[24697]_ ;
  assign \new_[888]_  = \new_[24684]_  & \new_[24671]_ ;
  assign \new_[889]_  = \new_[24658]_  & \new_[24645]_ ;
  assign \new_[890]_  = \new_[24632]_  & \new_[24619]_ ;
  assign \new_[891]_  = \new_[24606]_  & \new_[24593]_ ;
  assign \new_[892]_  = \new_[24580]_  & \new_[24567]_ ;
  assign \new_[893]_  = \new_[24554]_  & \new_[24541]_ ;
  assign \new_[894]_  = \new_[24528]_  & \new_[24515]_ ;
  assign \new_[895]_  = \new_[24502]_  & \new_[24489]_ ;
  assign \new_[896]_  = \new_[24476]_  & \new_[24463]_ ;
  assign \new_[897]_  = \new_[24450]_  & \new_[24437]_ ;
  assign \new_[898]_  = \new_[24424]_  & \new_[24411]_ ;
  assign \new_[899]_  = \new_[24398]_  & \new_[24385]_ ;
  assign \new_[900]_  = \new_[24372]_  & \new_[24359]_ ;
  assign \new_[901]_  = \new_[24346]_  & \new_[24333]_ ;
  assign \new_[902]_  = \new_[24320]_  & \new_[24307]_ ;
  assign \new_[903]_  = \new_[24294]_  & \new_[24281]_ ;
  assign \new_[904]_  = \new_[24268]_  & \new_[24255]_ ;
  assign \new_[905]_  = \new_[24242]_  & \new_[24229]_ ;
  assign \new_[906]_  = \new_[24216]_  & \new_[24203]_ ;
  assign \new_[907]_  = \new_[24190]_  & \new_[24177]_ ;
  assign \new_[908]_  = \new_[24164]_  & \new_[24151]_ ;
  assign \new_[909]_  = \new_[24138]_  & \new_[24125]_ ;
  assign \new_[910]_  = \new_[24112]_  & \new_[24099]_ ;
  assign \new_[911]_  = \new_[24086]_  & \new_[24073]_ ;
  assign \new_[912]_  = \new_[24060]_  & \new_[24047]_ ;
  assign \new_[913]_  = \new_[24034]_  & \new_[24021]_ ;
  assign \new_[914]_  = \new_[24008]_  & \new_[23995]_ ;
  assign \new_[915]_  = \new_[23982]_  & \new_[23969]_ ;
  assign \new_[916]_  = \new_[23956]_  & \new_[23943]_ ;
  assign \new_[917]_  = \new_[23930]_  & \new_[23917]_ ;
  assign \new_[918]_  = \new_[23904]_  & \new_[23891]_ ;
  assign \new_[919]_  = \new_[23878]_  & \new_[23865]_ ;
  assign \new_[920]_  = \new_[23852]_  & \new_[23839]_ ;
  assign \new_[921]_  = \new_[23826]_  & \new_[23813]_ ;
  assign \new_[922]_  = \new_[23800]_  & \new_[23787]_ ;
  assign \new_[923]_  = \new_[23774]_  & \new_[23761]_ ;
  assign \new_[924]_  = \new_[23748]_  & \new_[23735]_ ;
  assign \new_[925]_  = \new_[23722]_  & \new_[23709]_ ;
  assign \new_[926]_  = \new_[23696]_  & \new_[23683]_ ;
  assign \new_[927]_  = \new_[23670]_  & \new_[23657]_ ;
  assign \new_[928]_  = \new_[23644]_  & \new_[23631]_ ;
  assign \new_[929]_  = \new_[23618]_  & \new_[23605]_ ;
  assign \new_[930]_  = \new_[23592]_  & \new_[23579]_ ;
  assign \new_[931]_  = \new_[23566]_  & \new_[23553]_ ;
  assign \new_[932]_  = \new_[23540]_  & \new_[23527]_ ;
  assign \new_[933]_  = \new_[23514]_  & \new_[23501]_ ;
  assign \new_[934]_  = \new_[23488]_  & \new_[23475]_ ;
  assign \new_[935]_  = \new_[23462]_  & \new_[23449]_ ;
  assign \new_[936]_  = \new_[23436]_  & \new_[23423]_ ;
  assign \new_[937]_  = \new_[23410]_  & \new_[23397]_ ;
  assign \new_[938]_  = \new_[23384]_  & \new_[23371]_ ;
  assign \new_[939]_  = \new_[23358]_  & \new_[23345]_ ;
  assign \new_[940]_  = \new_[23332]_  & \new_[23319]_ ;
  assign \new_[941]_  = \new_[23306]_  & \new_[23293]_ ;
  assign \new_[942]_  = \new_[23280]_  & \new_[23267]_ ;
  assign \new_[943]_  = \new_[23254]_  & \new_[23241]_ ;
  assign \new_[944]_  = \new_[23228]_  & \new_[23215]_ ;
  assign \new_[945]_  = \new_[23202]_  & \new_[23189]_ ;
  assign \new_[946]_  = \new_[23176]_  & \new_[23163]_ ;
  assign \new_[947]_  = \new_[23150]_  & \new_[23137]_ ;
  assign \new_[948]_  = \new_[23124]_  & \new_[23111]_ ;
  assign \new_[949]_  = \new_[23098]_  & \new_[23085]_ ;
  assign \new_[950]_  = \new_[23072]_  & \new_[23059]_ ;
  assign \new_[951]_  = \new_[23046]_  & \new_[23033]_ ;
  assign \new_[952]_  = \new_[23020]_  & \new_[23007]_ ;
  assign \new_[953]_  = \new_[22994]_  & \new_[22981]_ ;
  assign \new_[954]_  = \new_[22968]_  & \new_[22955]_ ;
  assign \new_[955]_  = \new_[22942]_  & \new_[22929]_ ;
  assign \new_[956]_  = \new_[22916]_  & \new_[22903]_ ;
  assign \new_[957]_  = \new_[22890]_  & \new_[22877]_ ;
  assign \new_[958]_  = \new_[22864]_  & \new_[22851]_ ;
  assign \new_[959]_  = \new_[22838]_  & \new_[22825]_ ;
  assign \new_[960]_  = \new_[22812]_  & \new_[22799]_ ;
  assign \new_[961]_  = \new_[22786]_  & \new_[22773]_ ;
  assign \new_[962]_  = \new_[22760]_  & \new_[22747]_ ;
  assign \new_[963]_  = \new_[22734]_  & \new_[22721]_ ;
  assign \new_[964]_  = \new_[22708]_  & \new_[22695]_ ;
  assign \new_[965]_  = \new_[22682]_  & \new_[22669]_ ;
  assign \new_[966]_  = \new_[22656]_  & \new_[22643]_ ;
  assign \new_[967]_  = \new_[22630]_  & \new_[22617]_ ;
  assign \new_[968]_  = \new_[22604]_  & \new_[22591]_ ;
  assign \new_[969]_  = \new_[22578]_  & \new_[22565]_ ;
  assign \new_[970]_  = \new_[22552]_  & \new_[22539]_ ;
  assign \new_[971]_  = \new_[22526]_  & \new_[22513]_ ;
  assign \new_[972]_  = \new_[22500]_  & \new_[22487]_ ;
  assign \new_[973]_  = \new_[22474]_  & \new_[22461]_ ;
  assign \new_[974]_  = \new_[22448]_  & \new_[22435]_ ;
  assign \new_[975]_  = \new_[22422]_  & \new_[22409]_ ;
  assign \new_[976]_  = \new_[22396]_  & \new_[22383]_ ;
  assign \new_[977]_  = \new_[22370]_  & \new_[22357]_ ;
  assign \new_[978]_  = \new_[22344]_  & \new_[22331]_ ;
  assign \new_[979]_  = \new_[22318]_  & \new_[22305]_ ;
  assign \new_[980]_  = \new_[22292]_  & \new_[22279]_ ;
  assign \new_[981]_  = \new_[22266]_  & \new_[22253]_ ;
  assign \new_[982]_  = \new_[22240]_  & \new_[22227]_ ;
  assign \new_[983]_  = \new_[22214]_  & \new_[22201]_ ;
  assign \new_[984]_  = \new_[22188]_  & \new_[22175]_ ;
  assign \new_[985]_  = \new_[22162]_  & \new_[22149]_ ;
  assign \new_[986]_  = \new_[22136]_  & \new_[22123]_ ;
  assign \new_[987]_  = \new_[22110]_  & \new_[22097]_ ;
  assign \new_[988]_  = \new_[22084]_  & \new_[22071]_ ;
  assign \new_[989]_  = \new_[22058]_  & \new_[22045]_ ;
  assign \new_[990]_  = \new_[22032]_  & \new_[22019]_ ;
  assign \new_[991]_  = \new_[22006]_  & \new_[21993]_ ;
  assign \new_[992]_  = \new_[21980]_  & \new_[21967]_ ;
  assign \new_[993]_  = \new_[21954]_  & \new_[21941]_ ;
  assign \new_[994]_  = \new_[21928]_  & \new_[21915]_ ;
  assign \new_[995]_  = \new_[21902]_  & \new_[21889]_ ;
  assign \new_[996]_  = \new_[21876]_  & \new_[21863]_ ;
  assign \new_[997]_  = \new_[21850]_  & \new_[21837]_ ;
  assign \new_[998]_  = \new_[21824]_  & \new_[21811]_ ;
  assign \new_[999]_  = \new_[21798]_  & \new_[21785]_ ;
  assign \new_[1000]_  = \new_[21772]_  & \new_[21759]_ ;
  assign \new_[1001]_  = \new_[21746]_  & \new_[21733]_ ;
  assign \new_[1002]_  = \new_[21720]_  & \new_[21707]_ ;
  assign \new_[1003]_  = \new_[21694]_  & \new_[21681]_ ;
  assign \new_[1004]_  = \new_[21668]_  & \new_[21655]_ ;
  assign \new_[1005]_  = \new_[21642]_  & \new_[21629]_ ;
  assign \new_[1006]_  = \new_[21616]_  & \new_[21603]_ ;
  assign \new_[1007]_  = \new_[21590]_  & \new_[21577]_ ;
  assign \new_[1008]_  = \new_[21564]_  & \new_[21551]_ ;
  assign \new_[1009]_  = \new_[21538]_  & \new_[21525]_ ;
  assign \new_[1010]_  = \new_[21512]_  & \new_[21499]_ ;
  assign \new_[1011]_  = \new_[21486]_  & \new_[21473]_ ;
  assign \new_[1012]_  = \new_[21460]_  & \new_[21447]_ ;
  assign \new_[1013]_  = \new_[21434]_  & \new_[21421]_ ;
  assign \new_[1014]_  = \new_[21408]_  & \new_[21395]_ ;
  assign \new_[1015]_  = \new_[21382]_  & \new_[21369]_ ;
  assign \new_[1016]_  = \new_[21356]_  & \new_[21343]_ ;
  assign \new_[1017]_  = \new_[21330]_  & \new_[21317]_ ;
  assign \new_[1018]_  = \new_[21304]_  & \new_[21291]_ ;
  assign \new_[1019]_  = \new_[21278]_  & \new_[21265]_ ;
  assign \new_[1020]_  = \new_[21252]_  & \new_[21239]_ ;
  assign \new_[1021]_  = \new_[21226]_  & \new_[21213]_ ;
  assign \new_[1022]_  = \new_[21200]_  & \new_[21187]_ ;
  assign \new_[1023]_  = \new_[21174]_  & \new_[21161]_ ;
  assign \new_[1024]_  = \new_[21148]_  & \new_[21135]_ ;
  assign \new_[1025]_  = \new_[21122]_  & \new_[21109]_ ;
  assign \new_[1026]_  = \new_[21096]_  & \new_[21083]_ ;
  assign \new_[1027]_  = \new_[21070]_  & \new_[21057]_ ;
  assign \new_[1028]_  = \new_[21044]_  & \new_[21031]_ ;
  assign \new_[1029]_  = \new_[21018]_  & \new_[21005]_ ;
  assign \new_[1030]_  = \new_[20992]_  & \new_[20979]_ ;
  assign \new_[1031]_  = \new_[20966]_  & \new_[20953]_ ;
  assign \new_[1032]_  = \new_[20940]_  & \new_[20927]_ ;
  assign \new_[1033]_  = \new_[20914]_  & \new_[20901]_ ;
  assign \new_[1034]_  = \new_[20888]_  & \new_[20875]_ ;
  assign \new_[1035]_  = \new_[20862]_  & \new_[20849]_ ;
  assign \new_[1036]_  = \new_[20836]_  & \new_[20823]_ ;
  assign \new_[1037]_  = \new_[20810]_  & \new_[20797]_ ;
  assign \new_[1038]_  = \new_[20784]_  & \new_[20771]_ ;
  assign \new_[1039]_  = \new_[20758]_  & \new_[20745]_ ;
  assign \new_[1040]_  = \new_[20732]_  & \new_[20719]_ ;
  assign \new_[1041]_  = \new_[20706]_  & \new_[20693]_ ;
  assign \new_[1042]_  = \new_[20680]_  & \new_[20667]_ ;
  assign \new_[1043]_  = \new_[20654]_  & \new_[20641]_ ;
  assign \new_[1044]_  = \new_[20628]_  & \new_[20615]_ ;
  assign \new_[1045]_  = \new_[20602]_  & \new_[20589]_ ;
  assign \new_[1046]_  = \new_[20576]_  & \new_[20563]_ ;
  assign \new_[1047]_  = \new_[20550]_  & \new_[20537]_ ;
  assign \new_[1048]_  = \new_[20524]_  & \new_[20511]_ ;
  assign \new_[1049]_  = \new_[20498]_  & \new_[20485]_ ;
  assign \new_[1050]_  = \new_[20472]_  & \new_[20459]_ ;
  assign \new_[1051]_  = \new_[20446]_  & \new_[20433]_ ;
  assign \new_[1052]_  = \new_[20420]_  & \new_[20407]_ ;
  assign \new_[1053]_  = \new_[20394]_  & \new_[20381]_ ;
  assign \new_[1054]_  = \new_[20368]_  & \new_[20355]_ ;
  assign \new_[1055]_  = \new_[20342]_  & \new_[20329]_ ;
  assign \new_[1056]_  = \new_[20316]_  & \new_[20303]_ ;
  assign \new_[1057]_  = \new_[20290]_  & \new_[20277]_ ;
  assign \new_[1058]_  = \new_[20264]_  & \new_[20251]_ ;
  assign \new_[1059]_  = \new_[20238]_  & \new_[20225]_ ;
  assign \new_[1060]_  = \new_[20212]_  & \new_[20199]_ ;
  assign \new_[1061]_  = \new_[20186]_  & \new_[20173]_ ;
  assign \new_[1062]_  = \new_[20160]_  & \new_[20147]_ ;
  assign \new_[1063]_  = \new_[20134]_  & \new_[20121]_ ;
  assign \new_[1064]_  = \new_[20108]_  & \new_[20095]_ ;
  assign \new_[1065]_  = \new_[20082]_  & \new_[20069]_ ;
  assign \new_[1066]_  = \new_[20056]_  & \new_[20043]_ ;
  assign \new_[1067]_  = \new_[20030]_  & \new_[20017]_ ;
  assign \new_[1068]_  = \new_[20004]_  & \new_[19991]_ ;
  assign \new_[1069]_  = \new_[19978]_  & \new_[19965]_ ;
  assign \new_[1070]_  = \new_[19952]_  & \new_[19939]_ ;
  assign \new_[1071]_  = \new_[19926]_  & \new_[19913]_ ;
  assign \new_[1072]_  = \new_[19900]_  & \new_[19887]_ ;
  assign \new_[1073]_  = \new_[19874]_  & \new_[19861]_ ;
  assign \new_[1074]_  = \new_[19848]_  & \new_[19835]_ ;
  assign \new_[1075]_  = \new_[19822]_  & \new_[19809]_ ;
  assign \new_[1076]_  = \new_[19796]_  & \new_[19783]_ ;
  assign \new_[1077]_  = \new_[19770]_  & \new_[19757]_ ;
  assign \new_[1078]_  = \new_[19744]_  & \new_[19731]_ ;
  assign \new_[1079]_  = \new_[19718]_  & \new_[19705]_ ;
  assign \new_[1080]_  = \new_[19692]_  & \new_[19679]_ ;
  assign \new_[1081]_  = \new_[19666]_  & \new_[19653]_ ;
  assign \new_[1082]_  = \new_[19640]_  & \new_[19627]_ ;
  assign \new_[1083]_  = \new_[19614]_  & \new_[19601]_ ;
  assign \new_[1084]_  = \new_[19588]_  & \new_[19575]_ ;
  assign \new_[1085]_  = \new_[19562]_  & \new_[19549]_ ;
  assign \new_[1086]_  = \new_[19536]_  & \new_[19523]_ ;
  assign \new_[1087]_  = \new_[19510]_  & \new_[19497]_ ;
  assign \new_[1088]_  = \new_[19484]_  & \new_[19471]_ ;
  assign \new_[1089]_  = \new_[19458]_  & \new_[19445]_ ;
  assign \new_[1090]_  = \new_[19434]_  & \new_[19421]_ ;
  assign \new_[1091]_  = \new_[19410]_  & \new_[19397]_ ;
  assign \new_[1092]_  = \new_[19386]_  & \new_[19373]_ ;
  assign \new_[1093]_  = \new_[19362]_  & \new_[19349]_ ;
  assign \new_[1094]_  = \new_[19338]_  & \new_[19325]_ ;
  assign \new_[1095]_  = \new_[19314]_  & \new_[19301]_ ;
  assign \new_[1096]_  = \new_[19290]_  & \new_[19277]_ ;
  assign \new_[1097]_  = \new_[19266]_  & \new_[19253]_ ;
  assign \new_[1098]_  = \new_[19242]_  & \new_[19229]_ ;
  assign \new_[1099]_  = \new_[19218]_  & \new_[19205]_ ;
  assign \new_[1100]_  = \new_[19194]_  & \new_[19181]_ ;
  assign \new_[1101]_  = \new_[19170]_  & \new_[19157]_ ;
  assign \new_[1102]_  = \new_[19146]_  & \new_[19133]_ ;
  assign \new_[1103]_  = \new_[19122]_  & \new_[19109]_ ;
  assign \new_[1104]_  = \new_[19098]_  & \new_[19085]_ ;
  assign \new_[1105]_  = \new_[19074]_  & \new_[19061]_ ;
  assign \new_[1106]_  = \new_[19050]_  & \new_[19037]_ ;
  assign \new_[1107]_  = \new_[19026]_  & \new_[19013]_ ;
  assign \new_[1108]_  = \new_[19002]_  & \new_[18989]_ ;
  assign \new_[1109]_  = \new_[18978]_  & \new_[18965]_ ;
  assign \new_[1110]_  = \new_[18954]_  & \new_[18941]_ ;
  assign \new_[1111]_  = \new_[18930]_  & \new_[18917]_ ;
  assign \new_[1112]_  = \new_[18906]_  & \new_[18893]_ ;
  assign \new_[1113]_  = \new_[18882]_  & \new_[18869]_ ;
  assign \new_[1114]_  = \new_[18858]_  & \new_[18845]_ ;
  assign \new_[1115]_  = \new_[18834]_  & \new_[18821]_ ;
  assign \new_[1116]_  = \new_[18810]_  & \new_[18797]_ ;
  assign \new_[1117]_  = \new_[18786]_  & \new_[18773]_ ;
  assign \new_[1118]_  = \new_[18762]_  & \new_[18749]_ ;
  assign \new_[1119]_  = \new_[18738]_  & \new_[18725]_ ;
  assign \new_[1120]_  = \new_[18714]_  & \new_[18701]_ ;
  assign \new_[1121]_  = \new_[18690]_  & \new_[18677]_ ;
  assign \new_[1122]_  = \new_[18666]_  & \new_[18653]_ ;
  assign \new_[1123]_  = \new_[18642]_  & \new_[18629]_ ;
  assign \new_[1124]_  = \new_[18618]_  & \new_[18605]_ ;
  assign \new_[1125]_  = \new_[18594]_  & \new_[18581]_ ;
  assign \new_[1126]_  = \new_[18570]_  & \new_[18557]_ ;
  assign \new_[1127]_  = \new_[18546]_  & \new_[18533]_ ;
  assign \new_[1128]_  = \new_[18522]_  & \new_[18509]_ ;
  assign \new_[1129]_  = \new_[18498]_  & \new_[18485]_ ;
  assign \new_[1130]_  = \new_[18474]_  & \new_[18461]_ ;
  assign \new_[1131]_  = \new_[18450]_  & \new_[18437]_ ;
  assign \new_[1132]_  = \new_[18426]_  & \new_[18413]_ ;
  assign \new_[1133]_  = \new_[18402]_  & \new_[18389]_ ;
  assign \new_[1134]_  = \new_[18378]_  & \new_[18365]_ ;
  assign \new_[1135]_  = \new_[18354]_  & \new_[18341]_ ;
  assign \new_[1136]_  = \new_[18330]_  & \new_[18317]_ ;
  assign \new_[1137]_  = \new_[18306]_  & \new_[18293]_ ;
  assign \new_[1138]_  = \new_[18282]_  & \new_[18269]_ ;
  assign \new_[1139]_  = \new_[18258]_  & \new_[18245]_ ;
  assign \new_[1140]_  = \new_[18234]_  & \new_[18221]_ ;
  assign \new_[1141]_  = \new_[18210]_  & \new_[18197]_ ;
  assign \new_[1142]_  = \new_[18186]_  & \new_[18173]_ ;
  assign \new_[1143]_  = \new_[18162]_  & \new_[18149]_ ;
  assign \new_[1144]_  = \new_[18138]_  & \new_[18125]_ ;
  assign \new_[1145]_  = \new_[18114]_  & \new_[18101]_ ;
  assign \new_[1146]_  = \new_[18090]_  & \new_[18077]_ ;
  assign \new_[1147]_  = \new_[18066]_  & \new_[18053]_ ;
  assign \new_[1148]_  = \new_[18042]_  & \new_[18029]_ ;
  assign \new_[1149]_  = \new_[18018]_  & \new_[18005]_ ;
  assign \new_[1150]_  = \new_[17994]_  & \new_[17981]_ ;
  assign \new_[1151]_  = \new_[17970]_  & \new_[17957]_ ;
  assign \new_[1152]_  = \new_[17946]_  & \new_[17933]_ ;
  assign \new_[1153]_  = \new_[17922]_  & \new_[17909]_ ;
  assign \new_[1154]_  = \new_[17898]_  & \new_[17885]_ ;
  assign \new_[1155]_  = \new_[17874]_  & \new_[17861]_ ;
  assign \new_[1156]_  = \new_[17850]_  & \new_[17837]_ ;
  assign \new_[1157]_  = \new_[17826]_  & \new_[17813]_ ;
  assign \new_[1158]_  = \new_[17802]_  & \new_[17789]_ ;
  assign \new_[1159]_  = \new_[17778]_  & \new_[17765]_ ;
  assign \new_[1160]_  = \new_[17754]_  & \new_[17741]_ ;
  assign \new_[1161]_  = \new_[17730]_  & \new_[17717]_ ;
  assign \new_[1162]_  = \new_[17706]_  & \new_[17693]_ ;
  assign \new_[1163]_  = \new_[17682]_  & \new_[17669]_ ;
  assign \new_[1164]_  = \new_[17658]_  & \new_[17645]_ ;
  assign \new_[1165]_  = \new_[17634]_  & \new_[17621]_ ;
  assign \new_[1166]_  = \new_[17610]_  & \new_[17597]_ ;
  assign \new_[1167]_  = \new_[17586]_  & \new_[17573]_ ;
  assign \new_[1168]_  = \new_[17562]_  & \new_[17549]_ ;
  assign \new_[1169]_  = \new_[17538]_  & \new_[17525]_ ;
  assign \new_[1170]_  = \new_[17514]_  & \new_[17501]_ ;
  assign \new_[1171]_  = \new_[17490]_  & \new_[17477]_ ;
  assign \new_[1172]_  = \new_[17466]_  & \new_[17453]_ ;
  assign \new_[1173]_  = \new_[17442]_  & \new_[17429]_ ;
  assign \new_[1174]_  = \new_[17418]_  & \new_[17405]_ ;
  assign \new_[1175]_  = \new_[17394]_  & \new_[17381]_ ;
  assign \new_[1176]_  = \new_[17370]_  & \new_[17357]_ ;
  assign \new_[1177]_  = \new_[17346]_  & \new_[17333]_ ;
  assign \new_[1178]_  = \new_[17322]_  & \new_[17309]_ ;
  assign \new_[1179]_  = \new_[17298]_  & \new_[17285]_ ;
  assign \new_[1180]_  = \new_[17274]_  & \new_[17261]_ ;
  assign \new_[1181]_  = \new_[17250]_  & \new_[17237]_ ;
  assign \new_[1182]_  = \new_[17226]_  & \new_[17213]_ ;
  assign \new_[1183]_  = \new_[17202]_  & \new_[17189]_ ;
  assign \new_[1184]_  = \new_[17178]_  & \new_[17165]_ ;
  assign \new_[1185]_  = \new_[17154]_  & \new_[17141]_ ;
  assign \new_[1186]_  = \new_[17130]_  & \new_[17117]_ ;
  assign \new_[1187]_  = \new_[17106]_  & \new_[17093]_ ;
  assign \new_[1188]_  = \new_[17082]_  & \new_[17069]_ ;
  assign \new_[1189]_  = \new_[17058]_  & \new_[17045]_ ;
  assign \new_[1190]_  = \new_[17034]_  & \new_[17021]_ ;
  assign \new_[1191]_  = \new_[17010]_  & \new_[16997]_ ;
  assign \new_[1192]_  = \new_[16986]_  & \new_[16973]_ ;
  assign \new_[1193]_  = \new_[16962]_  & \new_[16949]_ ;
  assign \new_[1194]_  = \new_[16938]_  & \new_[16925]_ ;
  assign \new_[1195]_  = \new_[16914]_  & \new_[16901]_ ;
  assign \new_[1196]_  = \new_[16890]_  & \new_[16877]_ ;
  assign \new_[1197]_  = \new_[16866]_  & \new_[16853]_ ;
  assign \new_[1198]_  = \new_[16842]_  & \new_[16829]_ ;
  assign \new_[1199]_  = \new_[16818]_  & \new_[16805]_ ;
  assign \new_[1200]_  = \new_[16794]_  & \new_[16781]_ ;
  assign \new_[1201]_  = \new_[16770]_  & \new_[16757]_ ;
  assign \new_[1202]_  = \new_[16746]_  & \new_[16733]_ ;
  assign \new_[1203]_  = \new_[16722]_  & \new_[16709]_ ;
  assign \new_[1204]_  = \new_[16698]_  & \new_[16685]_ ;
  assign \new_[1205]_  = \new_[16674]_  & \new_[16661]_ ;
  assign \new_[1206]_  = \new_[16650]_  & \new_[16637]_ ;
  assign \new_[1207]_  = \new_[16626]_  & \new_[16613]_ ;
  assign \new_[1208]_  = \new_[16602]_  & \new_[16589]_ ;
  assign \new_[1209]_  = \new_[16578]_  & \new_[16565]_ ;
  assign \new_[1210]_  = \new_[16554]_  & \new_[16541]_ ;
  assign \new_[1211]_  = \new_[16530]_  & \new_[16517]_ ;
  assign \new_[1212]_  = \new_[16506]_  & \new_[16493]_ ;
  assign \new_[1213]_  = \new_[16482]_  & \new_[16469]_ ;
  assign \new_[1214]_  = \new_[16458]_  & \new_[16445]_ ;
  assign \new_[1215]_  = \new_[16434]_  & \new_[16421]_ ;
  assign \new_[1216]_  = \new_[16410]_  & \new_[16397]_ ;
  assign \new_[1217]_  = \new_[16386]_  & \new_[16373]_ ;
  assign \new_[1218]_  = \new_[16362]_  & \new_[16349]_ ;
  assign \new_[1219]_  = \new_[16338]_  & \new_[16325]_ ;
  assign \new_[1220]_  = \new_[16314]_  & \new_[16301]_ ;
  assign \new_[1221]_  = \new_[16290]_  & \new_[16277]_ ;
  assign \new_[1222]_  = \new_[16266]_  & \new_[16253]_ ;
  assign \new_[1223]_  = \new_[16242]_  & \new_[16229]_ ;
  assign \new_[1224]_  = \new_[16218]_  & \new_[16205]_ ;
  assign \new_[1225]_  = \new_[16194]_  & \new_[16181]_ ;
  assign \new_[1226]_  = \new_[16170]_  & \new_[16157]_ ;
  assign \new_[1227]_  = \new_[16146]_  & \new_[16133]_ ;
  assign \new_[1228]_  = \new_[16122]_  & \new_[16109]_ ;
  assign \new_[1229]_  = \new_[16098]_  & \new_[16085]_ ;
  assign \new_[1230]_  = \new_[16074]_  & \new_[16061]_ ;
  assign \new_[1231]_  = \new_[16050]_  & \new_[16037]_ ;
  assign \new_[1232]_  = \new_[16026]_  & \new_[16013]_ ;
  assign \new_[1233]_  = \new_[16002]_  & \new_[15989]_ ;
  assign \new_[1234]_  = \new_[15978]_  & \new_[15965]_ ;
  assign \new_[1235]_  = \new_[15954]_  & \new_[15941]_ ;
  assign \new_[1236]_  = \new_[15930]_  & \new_[15917]_ ;
  assign \new_[1237]_  = \new_[15906]_  & \new_[15893]_ ;
  assign \new_[1238]_  = \new_[15882]_  & \new_[15869]_ ;
  assign \new_[1239]_  = \new_[15858]_  & \new_[15845]_ ;
  assign \new_[1240]_  = \new_[15834]_  & \new_[15821]_ ;
  assign \new_[1241]_  = \new_[15810]_  & \new_[15797]_ ;
  assign \new_[1242]_  = \new_[15786]_  & \new_[15773]_ ;
  assign \new_[1243]_  = \new_[15762]_  & \new_[15749]_ ;
  assign \new_[1244]_  = \new_[15738]_  & \new_[15725]_ ;
  assign \new_[1245]_  = \new_[15714]_  & \new_[15701]_ ;
  assign \new_[1246]_  = \new_[15690]_  & \new_[15677]_ ;
  assign \new_[1247]_  = \new_[15666]_  & \new_[15653]_ ;
  assign \new_[1248]_  = \new_[15642]_  & \new_[15629]_ ;
  assign \new_[1249]_  = \new_[15618]_  & \new_[15605]_ ;
  assign \new_[1250]_  = \new_[15594]_  & \new_[15581]_ ;
  assign \new_[1251]_  = \new_[15570]_  & \new_[15557]_ ;
  assign \new_[1252]_  = \new_[15546]_  & \new_[15533]_ ;
  assign \new_[1253]_  = \new_[15522]_  & \new_[15509]_ ;
  assign \new_[1254]_  = \new_[15498]_  & \new_[15485]_ ;
  assign \new_[1255]_  = \new_[15474]_  & \new_[15461]_ ;
  assign \new_[1256]_  = \new_[15450]_  & \new_[15437]_ ;
  assign \new_[1257]_  = \new_[15426]_  & \new_[15413]_ ;
  assign \new_[1258]_  = \new_[15402]_  & \new_[15389]_ ;
  assign \new_[1259]_  = \new_[15378]_  & \new_[15365]_ ;
  assign \new_[1260]_  = \new_[15354]_  & \new_[15341]_ ;
  assign \new_[1261]_  = \new_[15330]_  & \new_[15317]_ ;
  assign \new_[1262]_  = \new_[15306]_  & \new_[15293]_ ;
  assign \new_[1263]_  = \new_[15282]_  & \new_[15269]_ ;
  assign \new_[1264]_  = \new_[15258]_  & \new_[15245]_ ;
  assign \new_[1265]_  = \new_[15234]_  & \new_[15221]_ ;
  assign \new_[1266]_  = \new_[15210]_  & \new_[15197]_ ;
  assign \new_[1267]_  = \new_[15186]_  & \new_[15173]_ ;
  assign \new_[1268]_  = \new_[15162]_  & \new_[15149]_ ;
  assign \new_[1269]_  = \new_[15138]_  & \new_[15125]_ ;
  assign \new_[1270]_  = \new_[15114]_  & \new_[15101]_ ;
  assign \new_[1271]_  = \new_[15090]_  & \new_[15077]_ ;
  assign \new_[1272]_  = \new_[15066]_  & \new_[15053]_ ;
  assign \new_[1273]_  = \new_[15042]_  & \new_[15029]_ ;
  assign \new_[1274]_  = \new_[15018]_  & \new_[15005]_ ;
  assign \new_[1275]_  = \new_[14994]_  & \new_[14981]_ ;
  assign \new_[1276]_  = \new_[14970]_  & \new_[14957]_ ;
  assign \new_[1277]_  = \new_[14946]_  & \new_[14933]_ ;
  assign \new_[1278]_  = \new_[14922]_  & \new_[14909]_ ;
  assign \new_[1279]_  = \new_[14898]_  & \new_[14885]_ ;
  assign \new_[1280]_  = \new_[14874]_  & \new_[14861]_ ;
  assign \new_[1281]_  = \new_[14850]_  & \new_[14839]_ ;
  assign \new_[1282]_  = \new_[14828]_  & \new_[14817]_ ;
  assign \new_[1283]_  = \new_[14806]_  & \new_[14795]_ ;
  assign \new_[1284]_  = \new_[14784]_  & \new_[14773]_ ;
  assign \new_[1285]_  = \new_[14762]_  & \new_[14751]_ ;
  assign \new_[1286]_  = \new_[14740]_  & \new_[14729]_ ;
  assign \new_[1287]_  = \new_[14718]_  & \new_[14707]_ ;
  assign \new_[1288]_  = \new_[14696]_  & \new_[14685]_ ;
  assign \new_[1289]_  = \new_[14674]_  & \new_[14663]_ ;
  assign \new_[1290]_  = \new_[14652]_  & \new_[14641]_ ;
  assign \new_[1291]_  = \new_[14630]_  & \new_[14619]_ ;
  assign \new_[1292]_  = \new_[14608]_  & \new_[14597]_ ;
  assign \new_[1293]_  = \new_[14586]_  & \new_[14575]_ ;
  assign \new_[1294]_  = \new_[14564]_  & \new_[14553]_ ;
  assign \new_[1295]_  = \new_[14542]_  & \new_[14531]_ ;
  assign \new_[1296]_  = \new_[14520]_  & \new_[14509]_ ;
  assign \new_[1297]_  = \new_[14498]_  & \new_[14487]_ ;
  assign \new_[1298]_  = \new_[14476]_  & \new_[14465]_ ;
  assign \new_[1299]_  = \new_[14454]_  & \new_[14443]_ ;
  assign \new_[1300]_  = \new_[14432]_  & \new_[14421]_ ;
  assign \new_[1301]_  = \new_[14410]_  & \new_[14399]_ ;
  assign \new_[1302]_  = \new_[14388]_  & \new_[14377]_ ;
  assign \new_[1303]_  = \new_[14366]_  & \new_[14355]_ ;
  assign \new_[1304]_  = \new_[14344]_  & \new_[14333]_ ;
  assign \new_[1305]_  = \new_[14322]_  & \new_[14311]_ ;
  assign \new_[1306]_  = \new_[14300]_  & \new_[14289]_ ;
  assign \new_[1307]_  = \new_[14278]_  & \new_[14267]_ ;
  assign \new_[1308]_  = \new_[14256]_  & \new_[14245]_ ;
  assign \new_[1309]_  = \new_[14234]_  & \new_[14223]_ ;
  assign \new_[1310]_  = \new_[14212]_  & \new_[14201]_ ;
  assign \new_[1311]_  = \new_[14190]_  & \new_[14179]_ ;
  assign \new_[1312]_  = \new_[14168]_  & \new_[14157]_ ;
  assign \new_[1313]_  = \new_[14146]_  & \new_[14135]_ ;
  assign \new_[1314]_  = \new_[14124]_  & \new_[14113]_ ;
  assign \new_[1315]_  = \new_[14102]_  & \new_[14091]_ ;
  assign \new_[1316]_  = \new_[14080]_  & \new_[14069]_ ;
  assign \new_[1317]_  = \new_[14058]_  & \new_[14047]_ ;
  assign \new_[1318]_  = \new_[14036]_  & \new_[14025]_ ;
  assign \new_[1319]_  = \new_[14014]_  & \new_[14003]_ ;
  assign \new_[1320]_  = \new_[13992]_  & \new_[13981]_ ;
  assign \new_[1321]_  = \new_[13970]_  & \new_[13959]_ ;
  assign \new_[1322]_  = \new_[13948]_  & \new_[13937]_ ;
  assign \new_[1323]_  = \new_[13926]_  & \new_[13915]_ ;
  assign \new_[1324]_  = \new_[13904]_  & \new_[13893]_ ;
  assign \new_[1325]_  = \new_[13882]_  & \new_[13871]_ ;
  assign \new_[1326]_  = \new_[13860]_  & \new_[13849]_ ;
  assign \new_[1327]_  = \new_[13838]_  & \new_[13827]_ ;
  assign \new_[1328]_  = \new_[13816]_  & \new_[13805]_ ;
  assign \new_[1329]_  = \new_[13794]_  & \new_[13783]_ ;
  assign \new_[1330]_  = \new_[13772]_  & \new_[13761]_ ;
  assign \new_[1331]_  = \new_[13750]_  & \new_[13739]_ ;
  assign \new_[1332]_  = \new_[13728]_  & \new_[13717]_ ;
  assign \new_[1333]_  = \new_[13706]_  & \new_[13695]_ ;
  assign \new_[1334]_  = \new_[13684]_  & \new_[13673]_ ;
  assign \new_[1335]_  = \new_[13662]_  & \new_[13651]_ ;
  assign \new_[1336]_  = \new_[13640]_  & \new_[13629]_ ;
  assign \new_[1337]_  = \new_[13618]_  & \new_[13607]_ ;
  assign \new_[1338]_  = \new_[13596]_  & \new_[13585]_ ;
  assign \new_[1339]_  = \new_[13574]_  & \new_[13563]_ ;
  assign \new_[1340]_  = \new_[13552]_  & \new_[13541]_ ;
  assign \new_[1341]_  = \new_[13530]_  & \new_[13519]_ ;
  assign \new_[1342]_  = \new_[13508]_  & \new_[13497]_ ;
  assign \new_[1343]_  = \new_[13486]_  & \new_[13475]_ ;
  assign \new_[1344]_  = \new_[13464]_  & \new_[13453]_ ;
  assign \new_[1345]_  = \new_[13442]_  & \new_[13431]_ ;
  assign \new_[1346]_  = \new_[13420]_  & \new_[13409]_ ;
  assign \new_[1347]_  = \new_[13398]_  & \new_[13387]_ ;
  assign \new_[1348]_  = \new_[13376]_  & \new_[13365]_ ;
  assign \new_[1349]_  = \new_[13354]_  & \new_[13343]_ ;
  assign \new_[1350]_  = \new_[13332]_  & \new_[13321]_ ;
  assign \new_[1351]_  = \new_[13310]_  & \new_[13299]_ ;
  assign \new_[1352]_  = \new_[13288]_  & \new_[13277]_ ;
  assign \new_[1353]_  = \new_[13266]_  & \new_[13255]_ ;
  assign \new_[1354]_  = \new_[13244]_  & \new_[13233]_ ;
  assign \new_[1355]_  = \new_[13222]_  & \new_[13211]_ ;
  assign \new_[1356]_  = \new_[13200]_  & \new_[13189]_ ;
  assign \new_[1357]_  = \new_[13178]_  & \new_[13167]_ ;
  assign \new_[1358]_  = \new_[13156]_  & \new_[13145]_ ;
  assign \new_[1359]_  = \new_[13134]_  & \new_[13123]_ ;
  assign \new_[1360]_  = \new_[13112]_  & \new_[13101]_ ;
  assign \new_[1361]_  = \new_[13090]_  & \new_[13079]_ ;
  assign \new_[1362]_  = \new_[13068]_  & \new_[13057]_ ;
  assign \new_[1363]_  = \new_[13046]_  & \new_[13035]_ ;
  assign \new_[1364]_  = \new_[13024]_  & \new_[13013]_ ;
  assign \new_[1365]_  = \new_[13002]_  & \new_[12991]_ ;
  assign \new_[1366]_  = \new_[12980]_  & \new_[12969]_ ;
  assign \new_[1367]_  = \new_[12958]_  & \new_[12947]_ ;
  assign \new_[1368]_  = \new_[12936]_  & \new_[12925]_ ;
  assign \new_[1369]_  = \new_[12914]_  & \new_[12903]_ ;
  assign \new_[1370]_  = \new_[12892]_  & \new_[12881]_ ;
  assign \new_[1371]_  = \new_[12870]_  & \new_[12859]_ ;
  assign \new_[1372]_  = \new_[12848]_  & \new_[12837]_ ;
  assign \new_[1373]_  = \new_[12826]_  & \new_[12815]_ ;
  assign \new_[1374]_  = \new_[12804]_  & \new_[12793]_ ;
  assign \new_[1375]_  = \new_[12782]_  & \new_[12771]_ ;
  assign \new_[1376]_  = \new_[12760]_  & \new_[12749]_ ;
  assign \new_[1377]_  = \new_[12738]_  & \new_[12727]_ ;
  assign \new_[1378]_  = \new_[12716]_  & \new_[12705]_ ;
  assign \new_[1379]_  = \new_[12694]_  & \new_[12683]_ ;
  assign \new_[1380]_  = \new_[12672]_  & \new_[12661]_ ;
  assign \new_[1381]_  = \new_[12650]_  & \new_[12639]_ ;
  assign \new_[1382]_  = \new_[12628]_  & \new_[12617]_ ;
  assign \new_[1383]_  = \new_[12606]_  & \new_[12595]_ ;
  assign \new_[1384]_  = \new_[12584]_  & \new_[12573]_ ;
  assign \new_[1385]_  = \new_[12562]_  & \new_[12551]_ ;
  assign \new_[1386]_  = \new_[12540]_  & \new_[12529]_ ;
  assign \new_[1387]_  = \new_[12518]_  & \new_[12507]_ ;
  assign \new_[1388]_  = \new_[12496]_  & \new_[12485]_ ;
  assign \new_[1389]_  = \new_[12474]_  & \new_[12463]_ ;
  assign \new_[1390]_  = \new_[12452]_  & \new_[12441]_ ;
  assign \new_[1391]_  = \new_[12430]_  & \new_[12419]_ ;
  assign \new_[1392]_  = \new_[12408]_  & \new_[12397]_ ;
  assign \new_[1393]_  = \new_[12386]_  & \new_[12375]_ ;
  assign \new_[1394]_  = \new_[12364]_  & \new_[12353]_ ;
  assign \new_[1395]_  = \new_[12342]_  & \new_[12331]_ ;
  assign \new_[1396]_  = \new_[12320]_  & \new_[12309]_ ;
  assign \new_[1397]_  = \new_[12298]_  & \new_[12287]_ ;
  assign \new_[1398]_  = \new_[12276]_  & \new_[12265]_ ;
  assign \new_[1399]_  = \new_[12254]_  & \new_[12243]_ ;
  assign \new_[1400]_  = \new_[12232]_  & \new_[12221]_ ;
  assign \new_[1401]_  = \new_[12210]_  & \new_[12199]_ ;
  assign \new_[1402]_  = \new_[12188]_  & \new_[12177]_ ;
  assign \new_[1403]_  = \new_[12166]_  & \new_[12155]_ ;
  assign \new_[1404]_  = \new_[12144]_  & \new_[12133]_ ;
  assign \new_[1405]_  = \new_[12122]_  & \new_[12111]_ ;
  assign \new_[1406]_  = \new_[12100]_  & \new_[12089]_ ;
  assign \new_[1407]_  = \new_[12078]_  & \new_[12067]_ ;
  assign \new_[1408]_  = \new_[12056]_  & \new_[12045]_ ;
  assign \new_[1409]_  = \new_[12034]_  & \new_[12023]_ ;
  assign \new_[1410]_  = \new_[12012]_  & \new_[12001]_ ;
  assign \new_[1411]_  = \new_[11990]_  & \new_[11979]_ ;
  assign \new_[1412]_  = \new_[11968]_  & \new_[11957]_ ;
  assign \new_[1413]_  = \new_[11946]_  & \new_[11935]_ ;
  assign \new_[1414]_  = \new_[11924]_  & \new_[11913]_ ;
  assign \new_[1415]_  = \new_[11902]_  & \new_[11891]_ ;
  assign \new_[1416]_  = \new_[11880]_  & \new_[11869]_ ;
  assign \new_[1417]_  = \new_[11858]_  & \new_[11847]_ ;
  assign \new_[1418]_  = \new_[11836]_  & \new_[11825]_ ;
  assign \new_[1419]_  = \new_[11814]_  & \new_[11803]_ ;
  assign \new_[1420]_  = \new_[11792]_  & \new_[11781]_ ;
  assign \new_[1421]_  = \new_[11770]_  & \new_[11759]_ ;
  assign \new_[1422]_  = \new_[11748]_  & \new_[11737]_ ;
  assign \new_[1423]_  = \new_[11726]_  & \new_[11715]_ ;
  assign \new_[1424]_  = \new_[11704]_  & \new_[11693]_ ;
  assign \new_[1425]_  = \new_[11682]_  & \new_[11671]_ ;
  assign \new_[1426]_  = \new_[11660]_  & \new_[11649]_ ;
  assign \new_[1427]_  = \new_[11638]_  & \new_[11627]_ ;
  assign \new_[1428]_  = \new_[11616]_  & \new_[11605]_ ;
  assign \new_[1429]_  = \new_[11594]_  & \new_[11583]_ ;
  assign \new_[1430]_  = \new_[11572]_  & \new_[11561]_ ;
  assign \new_[1431]_  = \new_[11550]_  & \new_[11539]_ ;
  assign \new_[1432]_  = \new_[11528]_  & \new_[11517]_ ;
  assign \new_[1433]_  = \new_[11506]_  & \new_[11495]_ ;
  assign \new_[1434]_  = \new_[11484]_  & \new_[11473]_ ;
  assign \new_[1435]_  = \new_[11462]_  & \new_[11451]_ ;
  assign \new_[1436]_  = \new_[11440]_  & \new_[11429]_ ;
  assign \new_[1437]_  = \new_[11418]_  & \new_[11407]_ ;
  assign \new_[1438]_  = \new_[11396]_  & \new_[11385]_ ;
  assign \new_[1439]_  = \new_[11374]_  & \new_[11363]_ ;
  assign \new_[1440]_  = \new_[11352]_  & \new_[11341]_ ;
  assign \new_[1441]_  = \new_[11330]_  & \new_[11319]_ ;
  assign \new_[1442]_  = \new_[11308]_  & \new_[11297]_ ;
  assign \new_[1443]_  = \new_[11286]_  & \new_[11275]_ ;
  assign \new_[1444]_  = \new_[11264]_  & \new_[11253]_ ;
  assign \new_[1445]_  = \new_[11242]_  & \new_[11231]_ ;
  assign \new_[1446]_  = \new_[11220]_  & \new_[11209]_ ;
  assign \new_[1447]_  = \new_[11198]_  & \new_[11187]_ ;
  assign \new_[1448]_  = \new_[11176]_  & \new_[11165]_ ;
  assign \new_[1449]_  = \new_[11154]_  & \new_[11143]_ ;
  assign \new_[1450]_  = \new_[11132]_  & \new_[11121]_ ;
  assign \new_[1451]_  = \new_[11110]_  & \new_[11099]_ ;
  assign \new_[1452]_  = \new_[11088]_  & \new_[11077]_ ;
  assign \new_[1453]_  = \new_[11066]_  & \new_[11055]_ ;
  assign \new_[1454]_  = \new_[11044]_  & \new_[11033]_ ;
  assign \new_[1455]_  = \new_[11022]_  & \new_[11011]_ ;
  assign \new_[1456]_  = \new_[11000]_  & \new_[10989]_ ;
  assign \new_[1457]_  = \new_[10978]_  & \new_[10967]_ ;
  assign \new_[1458]_  = \new_[10956]_  & \new_[10945]_ ;
  assign \new_[1459]_  = \new_[10934]_  & \new_[10923]_ ;
  assign \new_[1460]_  = \new_[10912]_  & \new_[10901]_ ;
  assign \new_[1461]_  = \new_[10890]_  & \new_[10879]_ ;
  assign \new_[1462]_  = \new_[10868]_  & \new_[10857]_ ;
  assign \new_[1463]_  = \new_[10846]_  & \new_[10835]_ ;
  assign \new_[1464]_  = \new_[10824]_  & \new_[10813]_ ;
  assign \new_[1465]_  = \new_[10802]_  & \new_[10791]_ ;
  assign \new_[1466]_  = \new_[10780]_  & \new_[10769]_ ;
  assign \new_[1467]_  = \new_[10758]_  & \new_[10747]_ ;
  assign \new_[1468]_  = \new_[10736]_  & \new_[10725]_ ;
  assign \new_[1469]_  = \new_[10714]_  & \new_[10703]_ ;
  assign \new_[1470]_  = \new_[10692]_  & \new_[10681]_ ;
  assign \new_[1471]_  = \new_[10670]_  & \new_[10659]_ ;
  assign \new_[1472]_  = \new_[10648]_  & \new_[10637]_ ;
  assign \new_[1473]_  = \new_[10626]_  & \new_[10615]_ ;
  assign \new_[1474]_  = \new_[10604]_  & \new_[10593]_ ;
  assign \new_[1475]_  = \new_[10582]_  & \new_[10571]_ ;
  assign \new_[1476]_  = \new_[10560]_  & \new_[10549]_ ;
  assign \new_[1477]_  = \new_[10538]_  & \new_[10527]_ ;
  assign \new_[1478]_  = \new_[10516]_  & \new_[10505]_ ;
  assign \new_[1479]_  = \new_[10494]_  & \new_[10483]_ ;
  assign \new_[1480]_  = \new_[10472]_  & \new_[10461]_ ;
  assign \new_[1481]_  = \new_[10450]_  & \new_[10439]_ ;
  assign \new_[1482]_  = \new_[10428]_  & \new_[10417]_ ;
  assign \new_[1483]_  = \new_[10406]_  & \new_[10395]_ ;
  assign \new_[1484]_  = \new_[10384]_  & \new_[10373]_ ;
  assign \new_[1485]_  = \new_[10362]_  & \new_[10351]_ ;
  assign \new_[1486]_  = \new_[10340]_  & \new_[10329]_ ;
  assign \new_[1487]_  = \new_[10318]_  & \new_[10307]_ ;
  assign \new_[1488]_  = \new_[10296]_  & \new_[10285]_ ;
  assign \new_[1489]_  = \new_[10274]_  & \new_[10263]_ ;
  assign \new_[1490]_  = \new_[10252]_  & \new_[10241]_ ;
  assign \new_[1491]_  = \new_[10230]_  & \new_[10219]_ ;
  assign \new_[1492]_  = \new_[10208]_  & \new_[10197]_ ;
  assign \new_[1493]_  = \new_[10186]_  & \new_[10175]_ ;
  assign \new_[1494]_  = \new_[10164]_  & \new_[10153]_ ;
  assign \new_[1495]_  = \new_[10142]_  & \new_[10131]_ ;
  assign \new_[1496]_  = \new_[10120]_  & \new_[10109]_ ;
  assign \new_[1497]_  = \new_[10098]_  & \new_[10087]_ ;
  assign \new_[1498]_  = \new_[10076]_  & \new_[10065]_ ;
  assign \new_[1499]_  = \new_[10054]_  & \new_[10043]_ ;
  assign \new_[1500]_  = \new_[10032]_  & \new_[10021]_ ;
  assign \new_[1501]_  = \new_[10010]_  & \new_[9999]_ ;
  assign \new_[1502]_  = \new_[9988]_  & \new_[9977]_ ;
  assign \new_[1503]_  = \new_[9966]_  & \new_[9955]_ ;
  assign \new_[1504]_  = \new_[9944]_  & \new_[9933]_ ;
  assign \new_[1505]_  = \new_[9922]_  & \new_[9911]_ ;
  assign \new_[1506]_  = \new_[9900]_  & \new_[9889]_ ;
  assign \new_[1507]_  = \new_[9878]_  & \new_[9867]_ ;
  assign \new_[1508]_  = \new_[9856]_  & \new_[9845]_ ;
  assign \new_[1509]_  = \new_[9834]_  & \new_[9823]_ ;
  assign \new_[1510]_  = \new_[9812]_  & \new_[9801]_ ;
  assign \new_[1511]_  = \new_[9790]_  & \new_[9779]_ ;
  assign \new_[1512]_  = \new_[9768]_  & \new_[9757]_ ;
  assign \new_[1513]_  = \new_[9746]_  & \new_[9735]_ ;
  assign \new_[1514]_  = \new_[9724]_  & \new_[9713]_ ;
  assign \new_[1515]_  = \new_[9702]_  & \new_[9691]_ ;
  assign \new_[1516]_  = \new_[9680]_  & \new_[9669]_ ;
  assign \new_[1517]_  = \new_[9658]_  & \new_[9647]_ ;
  assign \new_[1518]_  = \new_[9636]_  & \new_[9625]_ ;
  assign \new_[1519]_  = \new_[9614]_  & \new_[9603]_ ;
  assign \new_[1520]_  = \new_[9592]_  & \new_[9581]_ ;
  assign \new_[1521]_  = \new_[9570]_  & \new_[9559]_ ;
  assign \new_[1522]_  = \new_[9548]_  & \new_[9537]_ ;
  assign \new_[1523]_  = \new_[9526]_  & \new_[9515]_ ;
  assign \new_[1524]_  = \new_[9504]_  & \new_[9493]_ ;
  assign \new_[1525]_  = \new_[9482]_  & \new_[9471]_ ;
  assign \new_[1526]_  = \new_[9460]_  & \new_[9449]_ ;
  assign \new_[1527]_  = \new_[9438]_  & \new_[9427]_ ;
  assign \new_[1528]_  = \new_[9416]_  & \new_[9405]_ ;
  assign \new_[1529]_  = \new_[9394]_  & \new_[9383]_ ;
  assign \new_[1530]_  = \new_[9372]_  & \new_[9361]_ ;
  assign \new_[1531]_  = \new_[9350]_  & \new_[9339]_ ;
  assign \new_[1532]_  = \new_[9328]_  & \new_[9317]_ ;
  assign \new_[1533]_  = \new_[9306]_  & \new_[9295]_ ;
  assign \new_[1534]_  = \new_[9284]_  & \new_[9273]_ ;
  assign \new_[1535]_  = \new_[9262]_  & \new_[9251]_ ;
  assign \new_[1536]_  = \new_[9240]_  & \new_[9229]_ ;
  assign \new_[1537]_  = \new_[9218]_  & \new_[9207]_ ;
  assign \new_[1538]_  = \new_[9196]_  & \new_[9185]_ ;
  assign \new_[1539]_  = \new_[9174]_  & \new_[9163]_ ;
  assign \new_[1540]_  = \new_[9152]_  & \new_[9141]_ ;
  assign \new_[1541]_  = \new_[9130]_  & \new_[9119]_ ;
  assign \new_[1542]_  = \new_[9108]_  & \new_[9097]_ ;
  assign \new_[1543]_  = \new_[9086]_  & \new_[9075]_ ;
  assign \new_[1544]_  = \new_[9064]_  & \new_[9053]_ ;
  assign \new_[1545]_  = \new_[9042]_  & \new_[9031]_ ;
  assign \new_[1546]_  = \new_[9020]_  & \new_[9009]_ ;
  assign \new_[1547]_  = \new_[8998]_  & \new_[8987]_ ;
  assign \new_[1548]_  = \new_[8976]_  & \new_[8965]_ ;
  assign \new_[1549]_  = \new_[8954]_  & \new_[8943]_ ;
  assign \new_[1550]_  = \new_[8932]_  & \new_[8921]_ ;
  assign \new_[1551]_  = \new_[8910]_  & \new_[8899]_ ;
  assign \new_[1552]_  = \new_[8888]_  & \new_[8877]_ ;
  assign \new_[1553]_  = \new_[8866]_  & \new_[8855]_ ;
  assign \new_[1554]_  = \new_[8844]_  & \new_[8833]_ ;
  assign \new_[1555]_  = \new_[8822]_  & \new_[8811]_ ;
  assign \new_[1556]_  = \new_[8800]_  & \new_[8789]_ ;
  assign \new_[1557]_  = \new_[8778]_  & \new_[8767]_ ;
  assign \new_[1558]_  = \new_[8756]_  & \new_[8745]_ ;
  assign \new_[1559]_  = \new_[8734]_  & \new_[8723]_ ;
  assign \new_[1560]_  = \new_[8712]_  & \new_[8701]_ ;
  assign \new_[1561]_  = \new_[8690]_  & \new_[8679]_ ;
  assign \new_[1562]_  = \new_[8668]_  & \new_[8657]_ ;
  assign \new_[1563]_  = \new_[8646]_  & \new_[8635]_ ;
  assign \new_[1564]_  = \new_[8624]_  & \new_[8613]_ ;
  assign \new_[1565]_  = \new_[8602]_  & \new_[8591]_ ;
  assign \new_[1566]_  = \new_[8580]_  & \new_[8569]_ ;
  assign \new_[1567]_  = \new_[8558]_  & \new_[8547]_ ;
  assign \new_[1568]_  = \new_[8536]_  & \new_[8525]_ ;
  assign \new_[1569]_  = \new_[8514]_  & \new_[8503]_ ;
  assign \new_[1570]_  = \new_[8494]_  & \new_[8483]_ ;
  assign \new_[1571]_  = \new_[8474]_  & \new_[8463]_ ;
  assign \new_[1572]_  = \new_[8454]_  & \new_[8443]_ ;
  assign \new_[1573]_  = \new_[8434]_  & \new_[8423]_ ;
  assign \new_[1574]_  = \new_[8414]_  & \new_[8403]_ ;
  assign \new_[1575]_  = \new_[8394]_  & \new_[8383]_ ;
  assign \new_[1576]_  = \new_[8374]_  & \new_[8363]_ ;
  assign \new_[1577]_  = \new_[8354]_  & \new_[8343]_ ;
  assign \new_[1578]_  = \new_[8334]_  & \new_[8323]_ ;
  assign \new_[1579]_  = \new_[8314]_  & \new_[8303]_ ;
  assign \new_[1580]_  = \new_[8294]_  & \new_[8283]_ ;
  assign \new_[1581]_  = \new_[8274]_  & \new_[8263]_ ;
  assign \new_[1582]_  = \new_[8254]_  & \new_[8243]_ ;
  assign \new_[1583]_  = \new_[8234]_  & \new_[8223]_ ;
  assign \new_[1584]_  = \new_[8214]_  & \new_[8203]_ ;
  assign \new_[1585]_  = \new_[8194]_  & \new_[8183]_ ;
  assign \new_[1586]_  = \new_[8174]_  & \new_[8163]_ ;
  assign \new_[1587]_  = \new_[8154]_  & \new_[8143]_ ;
  assign \new_[1588]_  = \new_[8134]_  & \new_[8123]_ ;
  assign \new_[1589]_  = \new_[8114]_  & \new_[8103]_ ;
  assign \new_[1590]_  = \new_[8094]_  & \new_[8083]_ ;
  assign \new_[1591]_  = \new_[8074]_  & \new_[8063]_ ;
  assign \new_[1592]_  = \new_[8054]_  & \new_[8043]_ ;
  assign \new_[1593]_  = \new_[8034]_  & \new_[8023]_ ;
  assign \new_[1594]_  = \new_[8014]_  & \new_[8003]_ ;
  assign \new_[1595]_  = \new_[7994]_  & \new_[7983]_ ;
  assign \new_[1596]_  = \new_[7974]_  & \new_[7963]_ ;
  assign \new_[1597]_  = \new_[7954]_  & \new_[7943]_ ;
  assign \new_[1598]_  = \new_[7934]_  & \new_[7923]_ ;
  assign \new_[1599]_  = \new_[7914]_  & \new_[7903]_ ;
  assign \new_[1600]_  = \new_[7894]_  & \new_[7883]_ ;
  assign \new_[1601]_  = \new_[7874]_  & \new_[7863]_ ;
  assign \new_[1602]_  = \new_[7854]_  & \new_[7843]_ ;
  assign \new_[1603]_  = \new_[7834]_  & \new_[7823]_ ;
  assign \new_[1604]_  = \new_[7814]_  & \new_[7803]_ ;
  assign \new_[1605]_  = \new_[7794]_  & \new_[7783]_ ;
  assign \new_[1606]_  = \new_[7774]_  & \new_[7763]_ ;
  assign \new_[1607]_  = \new_[7754]_  & \new_[7743]_ ;
  assign \new_[1608]_  = \new_[7734]_  & \new_[7723]_ ;
  assign \new_[1609]_  = \new_[7714]_  & \new_[7703]_ ;
  assign \new_[1610]_  = \new_[7694]_  & \new_[7683]_ ;
  assign \new_[1611]_  = \new_[7674]_  & \new_[7663]_ ;
  assign \new_[1612]_  = \new_[7654]_  & \new_[7643]_ ;
  assign \new_[1613]_  = \new_[7634]_  & \new_[7623]_ ;
  assign \new_[1614]_  = \new_[7614]_  & \new_[7603]_ ;
  assign \new_[1615]_  = \new_[7594]_  & \new_[7583]_ ;
  assign \new_[1616]_  = \new_[7574]_  & \new_[7563]_ ;
  assign \new_[1617]_  = \new_[7554]_  & \new_[7543]_ ;
  assign \new_[1618]_  = \new_[7534]_  & \new_[7523]_ ;
  assign \new_[1619]_  = \new_[7514]_  & \new_[7503]_ ;
  assign \new_[1620]_  = \new_[7494]_  & \new_[7483]_ ;
  assign \new_[1621]_  = \new_[7474]_  & \new_[7463]_ ;
  assign \new_[1622]_  = \new_[7454]_  & \new_[7443]_ ;
  assign \new_[1623]_  = \new_[7434]_  & \new_[7423]_ ;
  assign \new_[1624]_  = \new_[7414]_  & \new_[7403]_ ;
  assign \new_[1625]_  = \new_[7394]_  & \new_[7383]_ ;
  assign \new_[1626]_  = \new_[7374]_  & \new_[7363]_ ;
  assign \new_[1627]_  = \new_[7354]_  & \new_[7343]_ ;
  assign \new_[1628]_  = \new_[7334]_  & \new_[7323]_ ;
  assign \new_[1629]_  = \new_[7314]_  & \new_[7303]_ ;
  assign \new_[1630]_  = \new_[7294]_  & \new_[7283]_ ;
  assign \new_[1631]_  = \new_[7274]_  & \new_[7263]_ ;
  assign \new_[1632]_  = \new_[7254]_  & \new_[7243]_ ;
  assign \new_[1633]_  = \new_[7234]_  & \new_[7223]_ ;
  assign \new_[1634]_  = \new_[7214]_  & \new_[7203]_ ;
  assign \new_[1635]_  = \new_[7194]_  & \new_[7183]_ ;
  assign \new_[1636]_  = \new_[7174]_  & \new_[7163]_ ;
  assign \new_[1637]_  = \new_[7154]_  & \new_[7143]_ ;
  assign \new_[1638]_  = \new_[7134]_  & \new_[7123]_ ;
  assign \new_[1639]_  = \new_[7114]_  & \new_[7103]_ ;
  assign \new_[1640]_  = \new_[7094]_  & \new_[7083]_ ;
  assign \new_[1641]_  = \new_[7074]_  & \new_[7063]_ ;
  assign \new_[1642]_  = \new_[7054]_  & \new_[7043]_ ;
  assign \new_[1643]_  = \new_[7034]_  & \new_[7023]_ ;
  assign \new_[1644]_  = \new_[7014]_  & \new_[7003]_ ;
  assign \new_[1645]_  = \new_[6994]_  & \new_[6983]_ ;
  assign \new_[1646]_  = \new_[6974]_  & \new_[6963]_ ;
  assign \new_[1647]_  = \new_[6954]_  & \new_[6943]_ ;
  assign \new_[1648]_  = \new_[6934]_  & \new_[6923]_ ;
  assign \new_[1649]_  = \new_[6914]_  & \new_[6903]_ ;
  assign \new_[1650]_  = \new_[6894]_  & \new_[6883]_ ;
  assign \new_[1651]_  = \new_[6874]_  & \new_[6863]_ ;
  assign \new_[1652]_  = \new_[6854]_  & \new_[6843]_ ;
  assign \new_[1653]_  = \new_[6834]_  & \new_[6823]_ ;
  assign \new_[1654]_  = \new_[6814]_  & \new_[6803]_ ;
  assign \new_[1655]_  = \new_[6794]_  & \new_[6783]_ ;
  assign \new_[1656]_  = \new_[6774]_  & \new_[6763]_ ;
  assign \new_[1657]_  = \new_[6754]_  & \new_[6743]_ ;
  assign \new_[1658]_  = \new_[6734]_  & \new_[6723]_ ;
  assign \new_[1659]_  = \new_[6714]_  & \new_[6703]_ ;
  assign \new_[1660]_  = \new_[6694]_  & \new_[6683]_ ;
  assign \new_[1661]_  = \new_[6674]_  & \new_[6663]_ ;
  assign \new_[1662]_  = \new_[6654]_  & \new_[6643]_ ;
  assign \new_[1663]_  = \new_[6634]_  & \new_[6623]_ ;
  assign \new_[1664]_  = \new_[6614]_  & \new_[6603]_ ;
  assign \new_[1665]_  = \new_[6594]_  & \new_[6585]_ ;
  assign \new_[1666]_  = \new_[6576]_  & \new_[6567]_ ;
  assign \new_[1667]_  = \new_[6558]_  & \new_[6549]_ ;
  assign \new_[1668]_  = \new_[6540]_  & \new_[6531]_ ;
  assign \new_[1669]_  = \new_[6522]_  & \new_[6513]_ ;
  assign \new_[1670]_  = \new_[6504]_  & \new_[6495]_ ;
  assign \new_[1671]_  = \new_[6486]_  & \new_[6477]_ ;
  assign \new_[1672]_  = \new_[6468]_  & \new_[6459]_ ;
  assign \new_[1673]_  = \new_[6450]_  & \new_[6441]_ ;
  assign \new_[1674]_  = \new_[6432]_  & \new_[6423]_ ;
  assign \new_[1675]_  = \new_[6414]_  & \new_[6405]_ ;
  assign \new_[1676]_  = \new_[6396]_  & \new_[6387]_ ;
  assign \new_[1677]_  = \new_[6378]_  & \new_[6369]_ ;
  assign \new_[1678]_  = \new_[6360]_  & \new_[6351]_ ;
  assign \new_[1679]_  = \new_[6342]_  & \new_[6333]_ ;
  assign \new_[1680]_  = \new_[6324]_  & \new_[6315]_ ;
  assign \new_[1681]_  = \new_[6306]_  & \new_[6297]_ ;
  assign \new_[1682]_  = \new_[6288]_  & \new_[6279]_ ;
  assign \new_[1683]_  = \new_[6270]_  & \new_[6261]_ ;
  assign \new_[1684]_  = \new_[6252]_  & \new_[6243]_ ;
  assign \new_[1685]_  = \new_[6234]_  & \new_[6225]_ ;
  assign \new_[1686]_  = \new_[6216]_  & \new_[6207]_ ;
  assign \new_[1687]_  = \new_[6198]_  & \new_[6189]_ ;
  assign \new_[1688]_  = \new_[6180]_  & \new_[6171]_ ;
  assign \new_[1689]_  = \new_[6162]_  & \new_[6153]_ ;
  assign \new_[1690]_  = \new_[6144]_  & \new_[6135]_ ;
  assign \new_[1691]_  = \new_[6126]_  & \new_[6117]_ ;
  assign \new_[1692]_  = \new_[6108]_  & \new_[6099]_ ;
  assign \new_[1693]_  = \new_[6090]_  & \new_[6081]_ ;
  assign \new_[1694]_  = \new_[6072]_  & \new_[6063]_ ;
  assign \new_[1695]_  = \new_[6054]_  & \new_[6045]_ ;
  assign \new_[1696]_  = \new_[6036]_  & \new_[6027]_ ;
  assign \new_[1697]_  = \new_[6018]_  & \new_[6009]_ ;
  assign \new_[1698]_  = \new_[6000]_  & \new_[5991]_ ;
  assign \new_[1699]_  = \new_[5982]_  & \new_[5973]_ ;
  assign \new_[1700]_  = \new_[5964]_  & \new_[5955]_ ;
  assign \new_[1701]_  = \new_[5946]_  & \new_[5937]_ ;
  assign \new_[1702]_  = \new_[5928]_  & \new_[5919]_ ;
  assign \new_[1703]_  = \new_[5910]_  & \new_[5901]_ ;
  assign \new_[1704]_  = \new_[5892]_  & \new_[5883]_ ;
  assign \new_[1705]_  = \new_[5874]_  & \new_[5865]_ ;
  assign \new_[1706]_  = \new_[5856]_  & \new_[5847]_ ;
  assign \new_[1707]_  = \new_[5838]_  & \new_[5829]_ ;
  assign \new_[1708]_  = \new_[5820]_  & \new_[5811]_ ;
  assign \new_[1709]_  = \new_[5802]_  & \new_[5793]_ ;
  assign \new_[1710]_  = \new_[5784]_  & \new_[5775]_ ;
  assign \new_[1711]_  = \new_[5766]_  & \new_[5757]_ ;
  assign \new_[1712]_  = \new_[5748]_  & \new_[5739]_ ;
  assign \new_[1713]_  = \new_[5730]_  & \new_[5721]_ ;
  assign \new_[1714]_  = \new_[5714]_  & \new_[5705]_ ;
  assign \new_[1715]_  = \new_[5698]_  & \new_[5689]_ ;
  assign \new_[1716]_  = \new_[5682]_  & \new_[5673]_ ;
  assign \new_[1717]_  = \new_[5666]_  & \new_[5657]_ ;
  assign \new_[1718]_  = \new_[5650]_  & \new_[5641]_ ;
  assign \new_[1719]_  = \new_[5634]_  & \new_[5625]_ ;
  assign \new_[1720]_  = \new_[5618]_  & \new_[5609]_ ;
  assign \new_[1721]_  = \new_[5602]_  & \new_[5593]_ ;
  assign \new_[1722]_  = \new_[5586]_  & \new_[5577]_ ;
  assign \new_[1723]_  = \new_[5570]_  & \new_[5561]_ ;
  assign \new_[1724]_  = \new_[5554]_  & \new_[5545]_ ;
  assign \new_[1725]_  = \new_[5538]_  & \new_[5529]_ ;
  assign \new_[1726]_  = \new_[5522]_  & \new_[5513]_ ;
  assign \new_[1727]_  = \new_[5506]_  & \new_[5497]_ ;
  assign \new_[1728]_  = \new_[5490]_  & \new_[5481]_ ;
  assign \new_[1729]_  = \new_[5474]_  & \new_[5467]_ ;
  assign \new_[1730]_  = \new_[5462]_  & \new_[5455]_ ;
  assign \new_[1731]_  = \new_[5450]_  & \new_[5443]_ ;
  assign \new_[1732]_  = \new_[5438]_  & \new_[5431]_ ;
  assign \new_[1733]_  = \new_[5426]_  & \new_[5421]_ ;
  assign \new_[1734]_  = \new_[5416]_  & \new_[5411]_ ;
  assign \new_[1735]_  = \new_[5406]_  & \new_[5401]_ ;
  assign \new_[1736]_  = \new_[5396]_  & \new_[5391]_ ;
  assign \new_[1737]_  = \new_[5386]_  & \new_[5381]_ ;
  assign \new_[1738]_  = \new_[5376]_  & \new_[5371]_ ;
  assign \new_[1739]_  = \new_[5366]_  & \new_[5361]_ ;
  assign \new_[1740]_  = \new_[5356]_  & \new_[5351]_ ;
  assign \new_[1741]_  = \new_[5346]_  & \new_[5341]_ ;
  assign \new_[1742]_  = \new_[5336]_  & \new_[5331]_ ;
  assign \new_[1743]_  = \new_[5326]_  & \new_[5321]_ ;
  assign \new_[1744]_  = \new_[5316]_  & \new_[5311]_ ;
  assign \new_[1745]_  = \new_[5306]_  & \new_[5301]_ ;
  assign \new_[1746]_  = \new_[5298]_  & \new_[5293]_ ;
  assign \new_[1747]_  = \new_[5290]_  & \new_[5287]_ ;
  assign \new_[1748]_  = \new_[5284]_  & \new_[5281]_ ;
  assign \new_[1749]_  = \new_[5278]_  & \new_[5275]_ ;
  assign \new_[1750]_  = \new_[5272]_  & \new_[5269]_ ;
  assign \new_[1751]_  = \new_[5266]_  & \new_[5263]_ ;
  assign \new_[1752]_  = \new_[5260]_  & \new_[5257]_ ;
  assign \new_[1756]_  = \new_[1750]_  | \new_[1751]_ ;
  assign \new_[1757]_  = \new_[1752]_  | \new_[1756]_ ;
  assign \new_[1761]_  = \new_[1747]_  | \new_[1748]_ ;
  assign \new_[1762]_  = \new_[1749]_  | \new_[1761]_ ;
  assign \new_[1763]_  = \new_[1762]_  | \new_[1757]_ ;
  assign \new_[1767]_  = \new_[1744]_  | \new_[1745]_ ;
  assign \new_[1768]_  = \new_[1746]_  | \new_[1767]_ ;
  assign \new_[1771]_  = \new_[1742]_  | \new_[1743]_ ;
  assign \new_[1774]_  = \new_[1740]_  | \new_[1741]_ ;
  assign \new_[1775]_  = \new_[1774]_  | \new_[1771]_ ;
  assign \new_[1776]_  = \new_[1775]_  | \new_[1768]_ ;
  assign \new_[1777]_  = \new_[1776]_  | \new_[1763]_ ;
  assign \new_[1781]_  = \new_[1737]_  | \new_[1738]_ ;
  assign \new_[1782]_  = \new_[1739]_  | \new_[1781]_ ;
  assign \new_[1785]_  = \new_[1735]_  | \new_[1736]_ ;
  assign \new_[1788]_  = \new_[1733]_  | \new_[1734]_ ;
  assign \new_[1789]_  = \new_[1788]_  | \new_[1785]_ ;
  assign \new_[1790]_  = \new_[1789]_  | \new_[1782]_ ;
  assign \new_[1794]_  = \new_[1730]_  | \new_[1731]_ ;
  assign \new_[1795]_  = \new_[1732]_  | \new_[1794]_ ;
  assign \new_[1798]_  = \new_[1728]_  | \new_[1729]_ ;
  assign \new_[1801]_  = \new_[1726]_  | \new_[1727]_ ;
  assign \new_[1802]_  = \new_[1801]_  | \new_[1798]_ ;
  assign \new_[1803]_  = \new_[1802]_  | \new_[1795]_ ;
  assign \new_[1804]_  = \new_[1803]_  | \new_[1790]_ ;
  assign \new_[1805]_  = \new_[1804]_  | \new_[1777]_ ;
  assign \new_[1809]_  = \new_[1723]_  | \new_[1724]_ ;
  assign \new_[1810]_  = \new_[1725]_  | \new_[1809]_ ;
  assign \new_[1814]_  = \new_[1720]_  | \new_[1721]_ ;
  assign \new_[1815]_  = \new_[1722]_  | \new_[1814]_ ;
  assign \new_[1816]_  = \new_[1815]_  | \new_[1810]_ ;
  assign \new_[1820]_  = \new_[1717]_  | \new_[1718]_ ;
  assign \new_[1821]_  = \new_[1719]_  | \new_[1820]_ ;
  assign \new_[1824]_  = \new_[1715]_  | \new_[1716]_ ;
  assign \new_[1827]_  = \new_[1713]_  | \new_[1714]_ ;
  assign \new_[1828]_  = \new_[1827]_  | \new_[1824]_ ;
  assign \new_[1829]_  = \new_[1828]_  | \new_[1821]_ ;
  assign \new_[1830]_  = \new_[1829]_  | \new_[1816]_ ;
  assign \new_[1834]_  = \new_[1710]_  | \new_[1711]_ ;
  assign \new_[1835]_  = \new_[1712]_  | \new_[1834]_ ;
  assign \new_[1838]_  = \new_[1708]_  | \new_[1709]_ ;
  assign \new_[1841]_  = \new_[1706]_  | \new_[1707]_ ;
  assign \new_[1842]_  = \new_[1841]_  | \new_[1838]_ ;
  assign \new_[1843]_  = \new_[1842]_  | \new_[1835]_ ;
  assign \new_[1847]_  = \new_[1703]_  | \new_[1704]_ ;
  assign \new_[1848]_  = \new_[1705]_  | \new_[1847]_ ;
  assign \new_[1851]_  = \new_[1701]_  | \new_[1702]_ ;
  assign \new_[1854]_  = \new_[1699]_  | \new_[1700]_ ;
  assign \new_[1855]_  = \new_[1854]_  | \new_[1851]_ ;
  assign \new_[1856]_  = \new_[1855]_  | \new_[1848]_ ;
  assign \new_[1857]_  = \new_[1856]_  | \new_[1843]_ ;
  assign \new_[1858]_  = \new_[1857]_  | \new_[1830]_ ;
  assign \new_[1859]_  = \new_[1858]_  | \new_[1805]_ ;
  assign \new_[1863]_  = \new_[1696]_  | \new_[1697]_ ;
  assign \new_[1864]_  = \new_[1698]_  | \new_[1863]_ ;
  assign \new_[1868]_  = \new_[1693]_  | \new_[1694]_ ;
  assign \new_[1869]_  = \new_[1695]_  | \new_[1868]_ ;
  assign \new_[1870]_  = \new_[1869]_  | \new_[1864]_ ;
  assign \new_[1874]_  = \new_[1690]_  | \new_[1691]_ ;
  assign \new_[1875]_  = \new_[1692]_  | \new_[1874]_ ;
  assign \new_[1878]_  = \new_[1688]_  | \new_[1689]_ ;
  assign \new_[1881]_  = \new_[1686]_  | \new_[1687]_ ;
  assign \new_[1882]_  = \new_[1881]_  | \new_[1878]_ ;
  assign \new_[1883]_  = \new_[1882]_  | \new_[1875]_ ;
  assign \new_[1884]_  = \new_[1883]_  | \new_[1870]_ ;
  assign \new_[1888]_  = \new_[1683]_  | \new_[1684]_ ;
  assign \new_[1889]_  = \new_[1685]_  | \new_[1888]_ ;
  assign \new_[1892]_  = \new_[1681]_  | \new_[1682]_ ;
  assign \new_[1895]_  = \new_[1679]_  | \new_[1680]_ ;
  assign \new_[1896]_  = \new_[1895]_  | \new_[1892]_ ;
  assign \new_[1897]_  = \new_[1896]_  | \new_[1889]_ ;
  assign \new_[1901]_  = \new_[1676]_  | \new_[1677]_ ;
  assign \new_[1902]_  = \new_[1678]_  | \new_[1901]_ ;
  assign \new_[1905]_  = \new_[1674]_  | \new_[1675]_ ;
  assign \new_[1908]_  = \new_[1672]_  | \new_[1673]_ ;
  assign \new_[1909]_  = \new_[1908]_  | \new_[1905]_ ;
  assign \new_[1910]_  = \new_[1909]_  | \new_[1902]_ ;
  assign \new_[1911]_  = \new_[1910]_  | \new_[1897]_ ;
  assign \new_[1912]_  = \new_[1911]_  | \new_[1884]_ ;
  assign \new_[1916]_  = \new_[1669]_  | \new_[1670]_ ;
  assign \new_[1917]_  = \new_[1671]_  | \new_[1916]_ ;
  assign \new_[1920]_  = \new_[1667]_  | \new_[1668]_ ;
  assign \new_[1923]_  = \new_[1665]_  | \new_[1666]_ ;
  assign \new_[1924]_  = \new_[1923]_  | \new_[1920]_ ;
  assign \new_[1925]_  = \new_[1924]_  | \new_[1917]_ ;
  assign \new_[1929]_  = \new_[1662]_  | \new_[1663]_ ;
  assign \new_[1930]_  = \new_[1664]_  | \new_[1929]_ ;
  assign \new_[1933]_  = \new_[1660]_  | \new_[1661]_ ;
  assign \new_[1936]_  = \new_[1658]_  | \new_[1659]_ ;
  assign \new_[1937]_  = \new_[1936]_  | \new_[1933]_ ;
  assign \new_[1938]_  = \new_[1937]_  | \new_[1930]_ ;
  assign \new_[1939]_  = \new_[1938]_  | \new_[1925]_ ;
  assign \new_[1943]_  = \new_[1655]_  | \new_[1656]_ ;
  assign \new_[1944]_  = \new_[1657]_  | \new_[1943]_ ;
  assign \new_[1947]_  = \new_[1653]_  | \new_[1654]_ ;
  assign \new_[1950]_  = \new_[1651]_  | \new_[1652]_ ;
  assign \new_[1951]_  = \new_[1950]_  | \new_[1947]_ ;
  assign \new_[1952]_  = \new_[1951]_  | \new_[1944]_ ;
  assign \new_[1956]_  = \new_[1648]_  | \new_[1649]_ ;
  assign \new_[1957]_  = \new_[1650]_  | \new_[1956]_ ;
  assign \new_[1960]_  = \new_[1646]_  | \new_[1647]_ ;
  assign \new_[1963]_  = \new_[1644]_  | \new_[1645]_ ;
  assign \new_[1964]_  = \new_[1963]_  | \new_[1960]_ ;
  assign \new_[1965]_  = \new_[1964]_  | \new_[1957]_ ;
  assign \new_[1966]_  = \new_[1965]_  | \new_[1952]_ ;
  assign \new_[1967]_  = \new_[1966]_  | \new_[1939]_ ;
  assign \new_[1968]_  = \new_[1967]_  | \new_[1912]_ ;
  assign \new_[1969]_  = \new_[1968]_  | \new_[1859]_ ;
  assign \new_[1973]_  = \new_[1641]_  | \new_[1642]_ ;
  assign \new_[1974]_  = \new_[1643]_  | \new_[1973]_ ;
  assign \new_[1978]_  = \new_[1638]_  | \new_[1639]_ ;
  assign \new_[1979]_  = \new_[1640]_  | \new_[1978]_ ;
  assign \new_[1980]_  = \new_[1979]_  | \new_[1974]_ ;
  assign \new_[1984]_  = \new_[1635]_  | \new_[1636]_ ;
  assign \new_[1985]_  = \new_[1637]_  | \new_[1984]_ ;
  assign \new_[1988]_  = \new_[1633]_  | \new_[1634]_ ;
  assign \new_[1991]_  = \new_[1631]_  | \new_[1632]_ ;
  assign \new_[1992]_  = \new_[1991]_  | \new_[1988]_ ;
  assign \new_[1993]_  = \new_[1992]_  | \new_[1985]_ ;
  assign \new_[1994]_  = \new_[1993]_  | \new_[1980]_ ;
  assign \new_[1998]_  = \new_[1628]_  | \new_[1629]_ ;
  assign \new_[1999]_  = \new_[1630]_  | \new_[1998]_ ;
  assign \new_[2002]_  = \new_[1626]_  | \new_[1627]_ ;
  assign \new_[2005]_  = \new_[1624]_  | \new_[1625]_ ;
  assign \new_[2006]_  = \new_[2005]_  | \new_[2002]_ ;
  assign \new_[2007]_  = \new_[2006]_  | \new_[1999]_ ;
  assign \new_[2011]_  = \new_[1621]_  | \new_[1622]_ ;
  assign \new_[2012]_  = \new_[1623]_  | \new_[2011]_ ;
  assign \new_[2015]_  = \new_[1619]_  | \new_[1620]_ ;
  assign \new_[2018]_  = \new_[1617]_  | \new_[1618]_ ;
  assign \new_[2019]_  = \new_[2018]_  | \new_[2015]_ ;
  assign \new_[2020]_  = \new_[2019]_  | \new_[2012]_ ;
  assign \new_[2021]_  = \new_[2020]_  | \new_[2007]_ ;
  assign \new_[2022]_  = \new_[2021]_  | \new_[1994]_ ;
  assign \new_[2026]_  = \new_[1614]_  | \new_[1615]_ ;
  assign \new_[2027]_  = \new_[1616]_  | \new_[2026]_ ;
  assign \new_[2030]_  = \new_[1612]_  | \new_[1613]_ ;
  assign \new_[2033]_  = \new_[1610]_  | \new_[1611]_ ;
  assign \new_[2034]_  = \new_[2033]_  | \new_[2030]_ ;
  assign \new_[2035]_  = \new_[2034]_  | \new_[2027]_ ;
  assign \new_[2039]_  = \new_[1607]_  | \new_[1608]_ ;
  assign \new_[2040]_  = \new_[1609]_  | \new_[2039]_ ;
  assign \new_[2043]_  = \new_[1605]_  | \new_[1606]_ ;
  assign \new_[2046]_  = \new_[1603]_  | \new_[1604]_ ;
  assign \new_[2047]_  = \new_[2046]_  | \new_[2043]_ ;
  assign \new_[2048]_  = \new_[2047]_  | \new_[2040]_ ;
  assign \new_[2049]_  = \new_[2048]_  | \new_[2035]_ ;
  assign \new_[2053]_  = \new_[1600]_  | \new_[1601]_ ;
  assign \new_[2054]_  = \new_[1602]_  | \new_[2053]_ ;
  assign \new_[2057]_  = \new_[1598]_  | \new_[1599]_ ;
  assign \new_[2060]_  = \new_[1596]_  | \new_[1597]_ ;
  assign \new_[2061]_  = \new_[2060]_  | \new_[2057]_ ;
  assign \new_[2062]_  = \new_[2061]_  | \new_[2054]_ ;
  assign \new_[2066]_  = \new_[1593]_  | \new_[1594]_ ;
  assign \new_[2067]_  = \new_[1595]_  | \new_[2066]_ ;
  assign \new_[2070]_  = \new_[1591]_  | \new_[1592]_ ;
  assign \new_[2073]_  = \new_[1589]_  | \new_[1590]_ ;
  assign \new_[2074]_  = \new_[2073]_  | \new_[2070]_ ;
  assign \new_[2075]_  = \new_[2074]_  | \new_[2067]_ ;
  assign \new_[2076]_  = \new_[2075]_  | \new_[2062]_ ;
  assign \new_[2077]_  = \new_[2076]_  | \new_[2049]_ ;
  assign \new_[2078]_  = \new_[2077]_  | \new_[2022]_ ;
  assign \new_[2082]_  = \new_[1586]_  | \new_[1587]_ ;
  assign \new_[2083]_  = \new_[1588]_  | \new_[2082]_ ;
  assign \new_[2087]_  = \new_[1583]_  | \new_[1584]_ ;
  assign \new_[2088]_  = \new_[1585]_  | \new_[2087]_ ;
  assign \new_[2089]_  = \new_[2088]_  | \new_[2083]_ ;
  assign \new_[2093]_  = \new_[1580]_  | \new_[1581]_ ;
  assign \new_[2094]_  = \new_[1582]_  | \new_[2093]_ ;
  assign \new_[2097]_  = \new_[1578]_  | \new_[1579]_ ;
  assign \new_[2100]_  = \new_[1576]_  | \new_[1577]_ ;
  assign \new_[2101]_  = \new_[2100]_  | \new_[2097]_ ;
  assign \new_[2102]_  = \new_[2101]_  | \new_[2094]_ ;
  assign \new_[2103]_  = \new_[2102]_  | \new_[2089]_ ;
  assign \new_[2107]_  = \new_[1573]_  | \new_[1574]_ ;
  assign \new_[2108]_  = \new_[1575]_  | \new_[2107]_ ;
  assign \new_[2111]_  = \new_[1571]_  | \new_[1572]_ ;
  assign \new_[2114]_  = \new_[1569]_  | \new_[1570]_ ;
  assign \new_[2115]_  = \new_[2114]_  | \new_[2111]_ ;
  assign \new_[2116]_  = \new_[2115]_  | \new_[2108]_ ;
  assign \new_[2120]_  = \new_[1566]_  | \new_[1567]_ ;
  assign \new_[2121]_  = \new_[1568]_  | \new_[2120]_ ;
  assign \new_[2124]_  = \new_[1564]_  | \new_[1565]_ ;
  assign \new_[2127]_  = \new_[1562]_  | \new_[1563]_ ;
  assign \new_[2128]_  = \new_[2127]_  | \new_[2124]_ ;
  assign \new_[2129]_  = \new_[2128]_  | \new_[2121]_ ;
  assign \new_[2130]_  = \new_[2129]_  | \new_[2116]_ ;
  assign \new_[2131]_  = \new_[2130]_  | \new_[2103]_ ;
  assign \new_[2135]_  = \new_[1559]_  | \new_[1560]_ ;
  assign \new_[2136]_  = \new_[1561]_  | \new_[2135]_ ;
  assign \new_[2139]_  = \new_[1557]_  | \new_[1558]_ ;
  assign \new_[2142]_  = \new_[1555]_  | \new_[1556]_ ;
  assign \new_[2143]_  = \new_[2142]_  | \new_[2139]_ ;
  assign \new_[2144]_  = \new_[2143]_  | \new_[2136]_ ;
  assign \new_[2148]_  = \new_[1552]_  | \new_[1553]_ ;
  assign \new_[2149]_  = \new_[1554]_  | \new_[2148]_ ;
  assign \new_[2152]_  = \new_[1550]_  | \new_[1551]_ ;
  assign \new_[2155]_  = \new_[1548]_  | \new_[1549]_ ;
  assign \new_[2156]_  = \new_[2155]_  | \new_[2152]_ ;
  assign \new_[2157]_  = \new_[2156]_  | \new_[2149]_ ;
  assign \new_[2158]_  = \new_[2157]_  | \new_[2144]_ ;
  assign \new_[2162]_  = \new_[1545]_  | \new_[1546]_ ;
  assign \new_[2163]_  = \new_[1547]_  | \new_[2162]_ ;
  assign \new_[2166]_  = \new_[1543]_  | \new_[1544]_ ;
  assign \new_[2169]_  = \new_[1541]_  | \new_[1542]_ ;
  assign \new_[2170]_  = \new_[2169]_  | \new_[2166]_ ;
  assign \new_[2171]_  = \new_[2170]_  | \new_[2163]_ ;
  assign \new_[2175]_  = \new_[1538]_  | \new_[1539]_ ;
  assign \new_[2176]_  = \new_[1540]_  | \new_[2175]_ ;
  assign \new_[2179]_  = \new_[1536]_  | \new_[1537]_ ;
  assign \new_[2182]_  = \new_[1534]_  | \new_[1535]_ ;
  assign \new_[2183]_  = \new_[2182]_  | \new_[2179]_ ;
  assign \new_[2184]_  = \new_[2183]_  | \new_[2176]_ ;
  assign \new_[2185]_  = \new_[2184]_  | \new_[2171]_ ;
  assign \new_[2186]_  = \new_[2185]_  | \new_[2158]_ ;
  assign \new_[2187]_  = \new_[2186]_  | \new_[2131]_ ;
  assign \new_[2188]_  = \new_[2187]_  | \new_[2078]_ ;
  assign \new_[2189]_  = \new_[2188]_  | \new_[1969]_ ;
  assign \new_[2193]_  = \new_[1531]_  | \new_[1532]_ ;
  assign \new_[2194]_  = \new_[1533]_  | \new_[2193]_ ;
  assign \new_[2198]_  = \new_[1528]_  | \new_[1529]_ ;
  assign \new_[2199]_  = \new_[1530]_  | \new_[2198]_ ;
  assign \new_[2200]_  = \new_[2199]_  | \new_[2194]_ ;
  assign \new_[2204]_  = \new_[1525]_  | \new_[1526]_ ;
  assign \new_[2205]_  = \new_[1527]_  | \new_[2204]_ ;
  assign \new_[2208]_  = \new_[1523]_  | \new_[1524]_ ;
  assign \new_[2211]_  = \new_[1521]_  | \new_[1522]_ ;
  assign \new_[2212]_  = \new_[2211]_  | \new_[2208]_ ;
  assign \new_[2213]_  = \new_[2212]_  | \new_[2205]_ ;
  assign \new_[2214]_  = \new_[2213]_  | \new_[2200]_ ;
  assign \new_[2218]_  = \new_[1518]_  | \new_[1519]_ ;
  assign \new_[2219]_  = \new_[1520]_  | \new_[2218]_ ;
  assign \new_[2222]_  = \new_[1516]_  | \new_[1517]_ ;
  assign \new_[2225]_  = \new_[1514]_  | \new_[1515]_ ;
  assign \new_[2226]_  = \new_[2225]_  | \new_[2222]_ ;
  assign \new_[2227]_  = \new_[2226]_  | \new_[2219]_ ;
  assign \new_[2231]_  = \new_[1511]_  | \new_[1512]_ ;
  assign \new_[2232]_  = \new_[1513]_  | \new_[2231]_ ;
  assign \new_[2235]_  = \new_[1509]_  | \new_[1510]_ ;
  assign \new_[2238]_  = \new_[1507]_  | \new_[1508]_ ;
  assign \new_[2239]_  = \new_[2238]_  | \new_[2235]_ ;
  assign \new_[2240]_  = \new_[2239]_  | \new_[2232]_ ;
  assign \new_[2241]_  = \new_[2240]_  | \new_[2227]_ ;
  assign \new_[2242]_  = \new_[2241]_  | \new_[2214]_ ;
  assign \new_[2246]_  = \new_[1504]_  | \new_[1505]_ ;
  assign \new_[2247]_  = \new_[1506]_  | \new_[2246]_ ;
  assign \new_[2251]_  = \new_[1501]_  | \new_[1502]_ ;
  assign \new_[2252]_  = \new_[1503]_  | \new_[2251]_ ;
  assign \new_[2253]_  = \new_[2252]_  | \new_[2247]_ ;
  assign \new_[2257]_  = \new_[1498]_  | \new_[1499]_ ;
  assign \new_[2258]_  = \new_[1500]_  | \new_[2257]_ ;
  assign \new_[2261]_  = \new_[1496]_  | \new_[1497]_ ;
  assign \new_[2264]_  = \new_[1494]_  | \new_[1495]_ ;
  assign \new_[2265]_  = \new_[2264]_  | \new_[2261]_ ;
  assign \new_[2266]_  = \new_[2265]_  | \new_[2258]_ ;
  assign \new_[2267]_  = \new_[2266]_  | \new_[2253]_ ;
  assign \new_[2271]_  = \new_[1491]_  | \new_[1492]_ ;
  assign \new_[2272]_  = \new_[1493]_  | \new_[2271]_ ;
  assign \new_[2275]_  = \new_[1489]_  | \new_[1490]_ ;
  assign \new_[2278]_  = \new_[1487]_  | \new_[1488]_ ;
  assign \new_[2279]_  = \new_[2278]_  | \new_[2275]_ ;
  assign \new_[2280]_  = \new_[2279]_  | \new_[2272]_ ;
  assign \new_[2284]_  = \new_[1484]_  | \new_[1485]_ ;
  assign \new_[2285]_  = \new_[1486]_  | \new_[2284]_ ;
  assign \new_[2288]_  = \new_[1482]_  | \new_[1483]_ ;
  assign \new_[2291]_  = \new_[1480]_  | \new_[1481]_ ;
  assign \new_[2292]_  = \new_[2291]_  | \new_[2288]_ ;
  assign \new_[2293]_  = \new_[2292]_  | \new_[2285]_ ;
  assign \new_[2294]_  = \new_[2293]_  | \new_[2280]_ ;
  assign \new_[2295]_  = \new_[2294]_  | \new_[2267]_ ;
  assign \new_[2296]_  = \new_[2295]_  | \new_[2242]_ ;
  assign \new_[2300]_  = \new_[1477]_  | \new_[1478]_ ;
  assign \new_[2301]_  = \new_[1479]_  | \new_[2300]_ ;
  assign \new_[2305]_  = \new_[1474]_  | \new_[1475]_ ;
  assign \new_[2306]_  = \new_[1476]_  | \new_[2305]_ ;
  assign \new_[2307]_  = \new_[2306]_  | \new_[2301]_ ;
  assign \new_[2311]_  = \new_[1471]_  | \new_[1472]_ ;
  assign \new_[2312]_  = \new_[1473]_  | \new_[2311]_ ;
  assign \new_[2315]_  = \new_[1469]_  | \new_[1470]_ ;
  assign \new_[2318]_  = \new_[1467]_  | \new_[1468]_ ;
  assign \new_[2319]_  = \new_[2318]_  | \new_[2315]_ ;
  assign \new_[2320]_  = \new_[2319]_  | \new_[2312]_ ;
  assign \new_[2321]_  = \new_[2320]_  | \new_[2307]_ ;
  assign \new_[2325]_  = \new_[1464]_  | \new_[1465]_ ;
  assign \new_[2326]_  = \new_[1466]_  | \new_[2325]_ ;
  assign \new_[2329]_  = \new_[1462]_  | \new_[1463]_ ;
  assign \new_[2332]_  = \new_[1460]_  | \new_[1461]_ ;
  assign \new_[2333]_  = \new_[2332]_  | \new_[2329]_ ;
  assign \new_[2334]_  = \new_[2333]_  | \new_[2326]_ ;
  assign \new_[2338]_  = \new_[1457]_  | \new_[1458]_ ;
  assign \new_[2339]_  = \new_[1459]_  | \new_[2338]_ ;
  assign \new_[2342]_  = \new_[1455]_  | \new_[1456]_ ;
  assign \new_[2345]_  = \new_[1453]_  | \new_[1454]_ ;
  assign \new_[2346]_  = \new_[2345]_  | \new_[2342]_ ;
  assign \new_[2347]_  = \new_[2346]_  | \new_[2339]_ ;
  assign \new_[2348]_  = \new_[2347]_  | \new_[2334]_ ;
  assign \new_[2349]_  = \new_[2348]_  | \new_[2321]_ ;
  assign \new_[2353]_  = \new_[1450]_  | \new_[1451]_ ;
  assign \new_[2354]_  = \new_[1452]_  | \new_[2353]_ ;
  assign \new_[2357]_  = \new_[1448]_  | \new_[1449]_ ;
  assign \new_[2360]_  = \new_[1446]_  | \new_[1447]_ ;
  assign \new_[2361]_  = \new_[2360]_  | \new_[2357]_ ;
  assign \new_[2362]_  = \new_[2361]_  | \new_[2354]_ ;
  assign \new_[2366]_  = \new_[1443]_  | \new_[1444]_ ;
  assign \new_[2367]_  = \new_[1445]_  | \new_[2366]_ ;
  assign \new_[2370]_  = \new_[1441]_  | \new_[1442]_ ;
  assign \new_[2373]_  = \new_[1439]_  | \new_[1440]_ ;
  assign \new_[2374]_  = \new_[2373]_  | \new_[2370]_ ;
  assign \new_[2375]_  = \new_[2374]_  | \new_[2367]_ ;
  assign \new_[2376]_  = \new_[2375]_  | \new_[2362]_ ;
  assign \new_[2380]_  = \new_[1436]_  | \new_[1437]_ ;
  assign \new_[2381]_  = \new_[1438]_  | \new_[2380]_ ;
  assign \new_[2384]_  = \new_[1434]_  | \new_[1435]_ ;
  assign \new_[2387]_  = \new_[1432]_  | \new_[1433]_ ;
  assign \new_[2388]_  = \new_[2387]_  | \new_[2384]_ ;
  assign \new_[2389]_  = \new_[2388]_  | \new_[2381]_ ;
  assign \new_[2393]_  = \new_[1429]_  | \new_[1430]_ ;
  assign \new_[2394]_  = \new_[1431]_  | \new_[2393]_ ;
  assign \new_[2397]_  = \new_[1427]_  | \new_[1428]_ ;
  assign \new_[2400]_  = \new_[1425]_  | \new_[1426]_ ;
  assign \new_[2401]_  = \new_[2400]_  | \new_[2397]_ ;
  assign \new_[2402]_  = \new_[2401]_  | \new_[2394]_ ;
  assign \new_[2403]_  = \new_[2402]_  | \new_[2389]_ ;
  assign \new_[2404]_  = \new_[2403]_  | \new_[2376]_ ;
  assign \new_[2405]_  = \new_[2404]_  | \new_[2349]_ ;
  assign \new_[2406]_  = \new_[2405]_  | \new_[2296]_ ;
  assign \new_[2410]_  = \new_[1422]_  | \new_[1423]_ ;
  assign \new_[2411]_  = \new_[1424]_  | \new_[2410]_ ;
  assign \new_[2415]_  = \new_[1419]_  | \new_[1420]_ ;
  assign \new_[2416]_  = \new_[1421]_  | \new_[2415]_ ;
  assign \new_[2417]_  = \new_[2416]_  | \new_[2411]_ ;
  assign \new_[2421]_  = \new_[1416]_  | \new_[1417]_ ;
  assign \new_[2422]_  = \new_[1418]_  | \new_[2421]_ ;
  assign \new_[2425]_  = \new_[1414]_  | \new_[1415]_ ;
  assign \new_[2428]_  = \new_[1412]_  | \new_[1413]_ ;
  assign \new_[2429]_  = \new_[2428]_  | \new_[2425]_ ;
  assign \new_[2430]_  = \new_[2429]_  | \new_[2422]_ ;
  assign \new_[2431]_  = \new_[2430]_  | \new_[2417]_ ;
  assign \new_[2435]_  = \new_[1409]_  | \new_[1410]_ ;
  assign \new_[2436]_  = \new_[1411]_  | \new_[2435]_ ;
  assign \new_[2439]_  = \new_[1407]_  | \new_[1408]_ ;
  assign \new_[2442]_  = \new_[1405]_  | \new_[1406]_ ;
  assign \new_[2443]_  = \new_[2442]_  | \new_[2439]_ ;
  assign \new_[2444]_  = \new_[2443]_  | \new_[2436]_ ;
  assign \new_[2448]_  = \new_[1402]_  | \new_[1403]_ ;
  assign \new_[2449]_  = \new_[1404]_  | \new_[2448]_ ;
  assign \new_[2452]_  = \new_[1400]_  | \new_[1401]_ ;
  assign \new_[2455]_  = \new_[1398]_  | \new_[1399]_ ;
  assign \new_[2456]_  = \new_[2455]_  | \new_[2452]_ ;
  assign \new_[2457]_  = \new_[2456]_  | \new_[2449]_ ;
  assign \new_[2458]_  = \new_[2457]_  | \new_[2444]_ ;
  assign \new_[2459]_  = \new_[2458]_  | \new_[2431]_ ;
  assign \new_[2463]_  = \new_[1395]_  | \new_[1396]_ ;
  assign \new_[2464]_  = \new_[1397]_  | \new_[2463]_ ;
  assign \new_[2467]_  = \new_[1393]_  | \new_[1394]_ ;
  assign \new_[2470]_  = \new_[1391]_  | \new_[1392]_ ;
  assign \new_[2471]_  = \new_[2470]_  | \new_[2467]_ ;
  assign \new_[2472]_  = \new_[2471]_  | \new_[2464]_ ;
  assign \new_[2476]_  = \new_[1388]_  | \new_[1389]_ ;
  assign \new_[2477]_  = \new_[1390]_  | \new_[2476]_ ;
  assign \new_[2480]_  = \new_[1386]_  | \new_[1387]_ ;
  assign \new_[2483]_  = \new_[1384]_  | \new_[1385]_ ;
  assign \new_[2484]_  = \new_[2483]_  | \new_[2480]_ ;
  assign \new_[2485]_  = \new_[2484]_  | \new_[2477]_ ;
  assign \new_[2486]_  = \new_[2485]_  | \new_[2472]_ ;
  assign \new_[2490]_  = \new_[1381]_  | \new_[1382]_ ;
  assign \new_[2491]_  = \new_[1383]_  | \new_[2490]_ ;
  assign \new_[2494]_  = \new_[1379]_  | \new_[1380]_ ;
  assign \new_[2497]_  = \new_[1377]_  | \new_[1378]_ ;
  assign \new_[2498]_  = \new_[2497]_  | \new_[2494]_ ;
  assign \new_[2499]_  = \new_[2498]_  | \new_[2491]_ ;
  assign \new_[2503]_  = \new_[1374]_  | \new_[1375]_ ;
  assign \new_[2504]_  = \new_[1376]_  | \new_[2503]_ ;
  assign \new_[2507]_  = \new_[1372]_  | \new_[1373]_ ;
  assign \new_[2510]_  = \new_[1370]_  | \new_[1371]_ ;
  assign \new_[2511]_  = \new_[2510]_  | \new_[2507]_ ;
  assign \new_[2512]_  = \new_[2511]_  | \new_[2504]_ ;
  assign \new_[2513]_  = \new_[2512]_  | \new_[2499]_ ;
  assign \new_[2514]_  = \new_[2513]_  | \new_[2486]_ ;
  assign \new_[2515]_  = \new_[2514]_  | \new_[2459]_ ;
  assign \new_[2519]_  = \new_[1367]_  | \new_[1368]_ ;
  assign \new_[2520]_  = \new_[1369]_  | \new_[2519]_ ;
  assign \new_[2524]_  = \new_[1364]_  | \new_[1365]_ ;
  assign \new_[2525]_  = \new_[1366]_  | \new_[2524]_ ;
  assign \new_[2526]_  = \new_[2525]_  | \new_[2520]_ ;
  assign \new_[2530]_  = \new_[1361]_  | \new_[1362]_ ;
  assign \new_[2531]_  = \new_[1363]_  | \new_[2530]_ ;
  assign \new_[2534]_  = \new_[1359]_  | \new_[1360]_ ;
  assign \new_[2537]_  = \new_[1357]_  | \new_[1358]_ ;
  assign \new_[2538]_  = \new_[2537]_  | \new_[2534]_ ;
  assign \new_[2539]_  = \new_[2538]_  | \new_[2531]_ ;
  assign \new_[2540]_  = \new_[2539]_  | \new_[2526]_ ;
  assign \new_[2544]_  = \new_[1354]_  | \new_[1355]_ ;
  assign \new_[2545]_  = \new_[1356]_  | \new_[2544]_ ;
  assign \new_[2548]_  = \new_[1352]_  | \new_[1353]_ ;
  assign \new_[2551]_  = \new_[1350]_  | \new_[1351]_ ;
  assign \new_[2552]_  = \new_[2551]_  | \new_[2548]_ ;
  assign \new_[2553]_  = \new_[2552]_  | \new_[2545]_ ;
  assign \new_[2557]_  = \new_[1347]_  | \new_[1348]_ ;
  assign \new_[2558]_  = \new_[1349]_  | \new_[2557]_ ;
  assign \new_[2561]_  = \new_[1345]_  | \new_[1346]_ ;
  assign \new_[2564]_  = \new_[1343]_  | \new_[1344]_ ;
  assign \new_[2565]_  = \new_[2564]_  | \new_[2561]_ ;
  assign \new_[2566]_  = \new_[2565]_  | \new_[2558]_ ;
  assign \new_[2567]_  = \new_[2566]_  | \new_[2553]_ ;
  assign \new_[2568]_  = \new_[2567]_  | \new_[2540]_ ;
  assign \new_[2572]_  = \new_[1340]_  | \new_[1341]_ ;
  assign \new_[2573]_  = \new_[1342]_  | \new_[2572]_ ;
  assign \new_[2576]_  = \new_[1338]_  | \new_[1339]_ ;
  assign \new_[2579]_  = \new_[1336]_  | \new_[1337]_ ;
  assign \new_[2580]_  = \new_[2579]_  | \new_[2576]_ ;
  assign \new_[2581]_  = \new_[2580]_  | \new_[2573]_ ;
  assign \new_[2585]_  = \new_[1333]_  | \new_[1334]_ ;
  assign \new_[2586]_  = \new_[1335]_  | \new_[2585]_ ;
  assign \new_[2589]_  = \new_[1331]_  | \new_[1332]_ ;
  assign \new_[2592]_  = \new_[1329]_  | \new_[1330]_ ;
  assign \new_[2593]_  = \new_[2592]_  | \new_[2589]_ ;
  assign \new_[2594]_  = \new_[2593]_  | \new_[2586]_ ;
  assign \new_[2595]_  = \new_[2594]_  | \new_[2581]_ ;
  assign \new_[2599]_  = \new_[1326]_  | \new_[1327]_ ;
  assign \new_[2600]_  = \new_[1328]_  | \new_[2599]_ ;
  assign \new_[2603]_  = \new_[1324]_  | \new_[1325]_ ;
  assign \new_[2606]_  = \new_[1322]_  | \new_[1323]_ ;
  assign \new_[2607]_  = \new_[2606]_  | \new_[2603]_ ;
  assign \new_[2608]_  = \new_[2607]_  | \new_[2600]_ ;
  assign \new_[2612]_  = \new_[1319]_  | \new_[1320]_ ;
  assign \new_[2613]_  = \new_[1321]_  | \new_[2612]_ ;
  assign \new_[2616]_  = \new_[1317]_  | \new_[1318]_ ;
  assign \new_[2619]_  = \new_[1315]_  | \new_[1316]_ ;
  assign \new_[2620]_  = \new_[2619]_  | \new_[2616]_ ;
  assign \new_[2621]_  = \new_[2620]_  | \new_[2613]_ ;
  assign \new_[2622]_  = \new_[2621]_  | \new_[2608]_ ;
  assign \new_[2623]_  = \new_[2622]_  | \new_[2595]_ ;
  assign \new_[2624]_  = \new_[2623]_  | \new_[2568]_ ;
  assign \new_[2625]_  = \new_[2624]_  | \new_[2515]_ ;
  assign \new_[2626]_  = \new_[2625]_  | \new_[2406]_ ;
  assign \new_[2627]_  = \new_[2626]_  | \new_[2189]_ ;
  assign \new_[2631]_  = \new_[1312]_  | \new_[1313]_ ;
  assign \new_[2632]_  = \new_[1314]_  | \new_[2631]_ ;
  assign \new_[2636]_  = \new_[1309]_  | \new_[1310]_ ;
  assign \new_[2637]_  = \new_[1311]_  | \new_[2636]_ ;
  assign \new_[2638]_  = \new_[2637]_  | \new_[2632]_ ;
  assign \new_[2642]_  = \new_[1306]_  | \new_[1307]_ ;
  assign \new_[2643]_  = \new_[1308]_  | \new_[2642]_ ;
  assign \new_[2646]_  = \new_[1304]_  | \new_[1305]_ ;
  assign \new_[2649]_  = \new_[1302]_  | \new_[1303]_ ;
  assign \new_[2650]_  = \new_[2649]_  | \new_[2646]_ ;
  assign \new_[2651]_  = \new_[2650]_  | \new_[2643]_ ;
  assign \new_[2652]_  = \new_[2651]_  | \new_[2638]_ ;
  assign \new_[2656]_  = \new_[1299]_  | \new_[1300]_ ;
  assign \new_[2657]_  = \new_[1301]_  | \new_[2656]_ ;
  assign \new_[2660]_  = \new_[1297]_  | \new_[1298]_ ;
  assign \new_[2663]_  = \new_[1295]_  | \new_[1296]_ ;
  assign \new_[2664]_  = \new_[2663]_  | \new_[2660]_ ;
  assign \new_[2665]_  = \new_[2664]_  | \new_[2657]_ ;
  assign \new_[2669]_  = \new_[1292]_  | \new_[1293]_ ;
  assign \new_[2670]_  = \new_[1294]_  | \new_[2669]_ ;
  assign \new_[2673]_  = \new_[1290]_  | \new_[1291]_ ;
  assign \new_[2676]_  = \new_[1288]_  | \new_[1289]_ ;
  assign \new_[2677]_  = \new_[2676]_  | \new_[2673]_ ;
  assign \new_[2678]_  = \new_[2677]_  | \new_[2670]_ ;
  assign \new_[2679]_  = \new_[2678]_  | \new_[2665]_ ;
  assign \new_[2680]_  = \new_[2679]_  | \new_[2652]_ ;
  assign \new_[2684]_  = \new_[1285]_  | \new_[1286]_ ;
  assign \new_[2685]_  = \new_[1287]_  | \new_[2684]_ ;
  assign \new_[2689]_  = \new_[1282]_  | \new_[1283]_ ;
  assign \new_[2690]_  = \new_[1284]_  | \new_[2689]_ ;
  assign \new_[2691]_  = \new_[2690]_  | \new_[2685]_ ;
  assign \new_[2695]_  = \new_[1279]_  | \new_[1280]_ ;
  assign \new_[2696]_  = \new_[1281]_  | \new_[2695]_ ;
  assign \new_[2699]_  = \new_[1277]_  | \new_[1278]_ ;
  assign \new_[2702]_  = \new_[1275]_  | \new_[1276]_ ;
  assign \new_[2703]_  = \new_[2702]_  | \new_[2699]_ ;
  assign \new_[2704]_  = \new_[2703]_  | \new_[2696]_ ;
  assign \new_[2705]_  = \new_[2704]_  | \new_[2691]_ ;
  assign \new_[2709]_  = \new_[1272]_  | \new_[1273]_ ;
  assign \new_[2710]_  = \new_[1274]_  | \new_[2709]_ ;
  assign \new_[2713]_  = \new_[1270]_  | \new_[1271]_ ;
  assign \new_[2716]_  = \new_[1268]_  | \new_[1269]_ ;
  assign \new_[2717]_  = \new_[2716]_  | \new_[2713]_ ;
  assign \new_[2718]_  = \new_[2717]_  | \new_[2710]_ ;
  assign \new_[2722]_  = \new_[1265]_  | \new_[1266]_ ;
  assign \new_[2723]_  = \new_[1267]_  | \new_[2722]_ ;
  assign \new_[2726]_  = \new_[1263]_  | \new_[1264]_ ;
  assign \new_[2729]_  = \new_[1261]_  | \new_[1262]_ ;
  assign \new_[2730]_  = \new_[2729]_  | \new_[2726]_ ;
  assign \new_[2731]_  = \new_[2730]_  | \new_[2723]_ ;
  assign \new_[2732]_  = \new_[2731]_  | \new_[2718]_ ;
  assign \new_[2733]_  = \new_[2732]_  | \new_[2705]_ ;
  assign \new_[2734]_  = \new_[2733]_  | \new_[2680]_ ;
  assign \new_[2738]_  = \new_[1258]_  | \new_[1259]_ ;
  assign \new_[2739]_  = \new_[1260]_  | \new_[2738]_ ;
  assign \new_[2743]_  = \new_[1255]_  | \new_[1256]_ ;
  assign \new_[2744]_  = \new_[1257]_  | \new_[2743]_ ;
  assign \new_[2745]_  = \new_[2744]_  | \new_[2739]_ ;
  assign \new_[2749]_  = \new_[1252]_  | \new_[1253]_ ;
  assign \new_[2750]_  = \new_[1254]_  | \new_[2749]_ ;
  assign \new_[2753]_  = \new_[1250]_  | \new_[1251]_ ;
  assign \new_[2756]_  = \new_[1248]_  | \new_[1249]_ ;
  assign \new_[2757]_  = \new_[2756]_  | \new_[2753]_ ;
  assign \new_[2758]_  = \new_[2757]_  | \new_[2750]_ ;
  assign \new_[2759]_  = \new_[2758]_  | \new_[2745]_ ;
  assign \new_[2763]_  = \new_[1245]_  | \new_[1246]_ ;
  assign \new_[2764]_  = \new_[1247]_  | \new_[2763]_ ;
  assign \new_[2767]_  = \new_[1243]_  | \new_[1244]_ ;
  assign \new_[2770]_  = \new_[1241]_  | \new_[1242]_ ;
  assign \new_[2771]_  = \new_[2770]_  | \new_[2767]_ ;
  assign \new_[2772]_  = \new_[2771]_  | \new_[2764]_ ;
  assign \new_[2776]_  = \new_[1238]_  | \new_[1239]_ ;
  assign \new_[2777]_  = \new_[1240]_  | \new_[2776]_ ;
  assign \new_[2780]_  = \new_[1236]_  | \new_[1237]_ ;
  assign \new_[2783]_  = \new_[1234]_  | \new_[1235]_ ;
  assign \new_[2784]_  = \new_[2783]_  | \new_[2780]_ ;
  assign \new_[2785]_  = \new_[2784]_  | \new_[2777]_ ;
  assign \new_[2786]_  = \new_[2785]_  | \new_[2772]_ ;
  assign \new_[2787]_  = \new_[2786]_  | \new_[2759]_ ;
  assign \new_[2791]_  = \new_[1231]_  | \new_[1232]_ ;
  assign \new_[2792]_  = \new_[1233]_  | \new_[2791]_ ;
  assign \new_[2795]_  = \new_[1229]_  | \new_[1230]_ ;
  assign \new_[2798]_  = \new_[1227]_  | \new_[1228]_ ;
  assign \new_[2799]_  = \new_[2798]_  | \new_[2795]_ ;
  assign \new_[2800]_  = \new_[2799]_  | \new_[2792]_ ;
  assign \new_[2804]_  = \new_[1224]_  | \new_[1225]_ ;
  assign \new_[2805]_  = \new_[1226]_  | \new_[2804]_ ;
  assign \new_[2808]_  = \new_[1222]_  | \new_[1223]_ ;
  assign \new_[2811]_  = \new_[1220]_  | \new_[1221]_ ;
  assign \new_[2812]_  = \new_[2811]_  | \new_[2808]_ ;
  assign \new_[2813]_  = \new_[2812]_  | \new_[2805]_ ;
  assign \new_[2814]_  = \new_[2813]_  | \new_[2800]_ ;
  assign \new_[2818]_  = \new_[1217]_  | \new_[1218]_ ;
  assign \new_[2819]_  = \new_[1219]_  | \new_[2818]_ ;
  assign \new_[2822]_  = \new_[1215]_  | \new_[1216]_ ;
  assign \new_[2825]_  = \new_[1213]_  | \new_[1214]_ ;
  assign \new_[2826]_  = \new_[2825]_  | \new_[2822]_ ;
  assign \new_[2827]_  = \new_[2826]_  | \new_[2819]_ ;
  assign \new_[2831]_  = \new_[1210]_  | \new_[1211]_ ;
  assign \new_[2832]_  = \new_[1212]_  | \new_[2831]_ ;
  assign \new_[2835]_  = \new_[1208]_  | \new_[1209]_ ;
  assign \new_[2838]_  = \new_[1206]_  | \new_[1207]_ ;
  assign \new_[2839]_  = \new_[2838]_  | \new_[2835]_ ;
  assign \new_[2840]_  = \new_[2839]_  | \new_[2832]_ ;
  assign \new_[2841]_  = \new_[2840]_  | \new_[2827]_ ;
  assign \new_[2842]_  = \new_[2841]_  | \new_[2814]_ ;
  assign \new_[2843]_  = \new_[2842]_  | \new_[2787]_ ;
  assign \new_[2844]_  = \new_[2843]_  | \new_[2734]_ ;
  assign \new_[2848]_  = \new_[1203]_  | \new_[1204]_ ;
  assign \new_[2849]_  = \new_[1205]_  | \new_[2848]_ ;
  assign \new_[2853]_  = \new_[1200]_  | \new_[1201]_ ;
  assign \new_[2854]_  = \new_[1202]_  | \new_[2853]_ ;
  assign \new_[2855]_  = \new_[2854]_  | \new_[2849]_ ;
  assign \new_[2859]_  = \new_[1197]_  | \new_[1198]_ ;
  assign \new_[2860]_  = \new_[1199]_  | \new_[2859]_ ;
  assign \new_[2863]_  = \new_[1195]_  | \new_[1196]_ ;
  assign \new_[2866]_  = \new_[1193]_  | \new_[1194]_ ;
  assign \new_[2867]_  = \new_[2866]_  | \new_[2863]_ ;
  assign \new_[2868]_  = \new_[2867]_  | \new_[2860]_ ;
  assign \new_[2869]_  = \new_[2868]_  | \new_[2855]_ ;
  assign \new_[2873]_  = \new_[1190]_  | \new_[1191]_ ;
  assign \new_[2874]_  = \new_[1192]_  | \new_[2873]_ ;
  assign \new_[2877]_  = \new_[1188]_  | \new_[1189]_ ;
  assign \new_[2880]_  = \new_[1186]_  | \new_[1187]_ ;
  assign \new_[2881]_  = \new_[2880]_  | \new_[2877]_ ;
  assign \new_[2882]_  = \new_[2881]_  | \new_[2874]_ ;
  assign \new_[2886]_  = \new_[1183]_  | \new_[1184]_ ;
  assign \new_[2887]_  = \new_[1185]_  | \new_[2886]_ ;
  assign \new_[2890]_  = \new_[1181]_  | \new_[1182]_ ;
  assign \new_[2893]_  = \new_[1179]_  | \new_[1180]_ ;
  assign \new_[2894]_  = \new_[2893]_  | \new_[2890]_ ;
  assign \new_[2895]_  = \new_[2894]_  | \new_[2887]_ ;
  assign \new_[2896]_  = \new_[2895]_  | \new_[2882]_ ;
  assign \new_[2897]_  = \new_[2896]_  | \new_[2869]_ ;
  assign \new_[2901]_  = \new_[1176]_  | \new_[1177]_ ;
  assign \new_[2902]_  = \new_[1178]_  | \new_[2901]_ ;
  assign \new_[2905]_  = \new_[1174]_  | \new_[1175]_ ;
  assign \new_[2908]_  = \new_[1172]_  | \new_[1173]_ ;
  assign \new_[2909]_  = \new_[2908]_  | \new_[2905]_ ;
  assign \new_[2910]_  = \new_[2909]_  | \new_[2902]_ ;
  assign \new_[2914]_  = \new_[1169]_  | \new_[1170]_ ;
  assign \new_[2915]_  = \new_[1171]_  | \new_[2914]_ ;
  assign \new_[2918]_  = \new_[1167]_  | \new_[1168]_ ;
  assign \new_[2921]_  = \new_[1165]_  | \new_[1166]_ ;
  assign \new_[2922]_  = \new_[2921]_  | \new_[2918]_ ;
  assign \new_[2923]_  = \new_[2922]_  | \new_[2915]_ ;
  assign \new_[2924]_  = \new_[2923]_  | \new_[2910]_ ;
  assign \new_[2928]_  = \new_[1162]_  | \new_[1163]_ ;
  assign \new_[2929]_  = \new_[1164]_  | \new_[2928]_ ;
  assign \new_[2932]_  = \new_[1160]_  | \new_[1161]_ ;
  assign \new_[2935]_  = \new_[1158]_  | \new_[1159]_ ;
  assign \new_[2936]_  = \new_[2935]_  | \new_[2932]_ ;
  assign \new_[2937]_  = \new_[2936]_  | \new_[2929]_ ;
  assign \new_[2941]_  = \new_[1155]_  | \new_[1156]_ ;
  assign \new_[2942]_  = \new_[1157]_  | \new_[2941]_ ;
  assign \new_[2945]_  = \new_[1153]_  | \new_[1154]_ ;
  assign \new_[2948]_  = \new_[1151]_  | \new_[1152]_ ;
  assign \new_[2949]_  = \new_[2948]_  | \new_[2945]_ ;
  assign \new_[2950]_  = \new_[2949]_  | \new_[2942]_ ;
  assign \new_[2951]_  = \new_[2950]_  | \new_[2937]_ ;
  assign \new_[2952]_  = \new_[2951]_  | \new_[2924]_ ;
  assign \new_[2953]_  = \new_[2952]_  | \new_[2897]_ ;
  assign \new_[2957]_  = \new_[1148]_  | \new_[1149]_ ;
  assign \new_[2958]_  = \new_[1150]_  | \new_[2957]_ ;
  assign \new_[2962]_  = \new_[1145]_  | \new_[1146]_ ;
  assign \new_[2963]_  = \new_[1147]_  | \new_[2962]_ ;
  assign \new_[2964]_  = \new_[2963]_  | \new_[2958]_ ;
  assign \new_[2968]_  = \new_[1142]_  | \new_[1143]_ ;
  assign \new_[2969]_  = \new_[1144]_  | \new_[2968]_ ;
  assign \new_[2972]_  = \new_[1140]_  | \new_[1141]_ ;
  assign \new_[2975]_  = \new_[1138]_  | \new_[1139]_ ;
  assign \new_[2976]_  = \new_[2975]_  | \new_[2972]_ ;
  assign \new_[2977]_  = \new_[2976]_  | \new_[2969]_ ;
  assign \new_[2978]_  = \new_[2977]_  | \new_[2964]_ ;
  assign \new_[2982]_  = \new_[1135]_  | \new_[1136]_ ;
  assign \new_[2983]_  = \new_[1137]_  | \new_[2982]_ ;
  assign \new_[2986]_  = \new_[1133]_  | \new_[1134]_ ;
  assign \new_[2989]_  = \new_[1131]_  | \new_[1132]_ ;
  assign \new_[2990]_  = \new_[2989]_  | \new_[2986]_ ;
  assign \new_[2991]_  = \new_[2990]_  | \new_[2983]_ ;
  assign \new_[2995]_  = \new_[1128]_  | \new_[1129]_ ;
  assign \new_[2996]_  = \new_[1130]_  | \new_[2995]_ ;
  assign \new_[2999]_  = \new_[1126]_  | \new_[1127]_ ;
  assign \new_[3002]_  = \new_[1124]_  | \new_[1125]_ ;
  assign \new_[3003]_  = \new_[3002]_  | \new_[2999]_ ;
  assign \new_[3004]_  = \new_[3003]_  | \new_[2996]_ ;
  assign \new_[3005]_  = \new_[3004]_  | \new_[2991]_ ;
  assign \new_[3006]_  = \new_[3005]_  | \new_[2978]_ ;
  assign \new_[3010]_  = \new_[1121]_  | \new_[1122]_ ;
  assign \new_[3011]_  = \new_[1123]_  | \new_[3010]_ ;
  assign \new_[3014]_  = \new_[1119]_  | \new_[1120]_ ;
  assign \new_[3017]_  = \new_[1117]_  | \new_[1118]_ ;
  assign \new_[3018]_  = \new_[3017]_  | \new_[3014]_ ;
  assign \new_[3019]_  = \new_[3018]_  | \new_[3011]_ ;
  assign \new_[3023]_  = \new_[1114]_  | \new_[1115]_ ;
  assign \new_[3024]_  = \new_[1116]_  | \new_[3023]_ ;
  assign \new_[3027]_  = \new_[1112]_  | \new_[1113]_ ;
  assign \new_[3030]_  = \new_[1110]_  | \new_[1111]_ ;
  assign \new_[3031]_  = \new_[3030]_  | \new_[3027]_ ;
  assign \new_[3032]_  = \new_[3031]_  | \new_[3024]_ ;
  assign \new_[3033]_  = \new_[3032]_  | \new_[3019]_ ;
  assign \new_[3037]_  = \new_[1107]_  | \new_[1108]_ ;
  assign \new_[3038]_  = \new_[1109]_  | \new_[3037]_ ;
  assign \new_[3041]_  = \new_[1105]_  | \new_[1106]_ ;
  assign \new_[3044]_  = \new_[1103]_  | \new_[1104]_ ;
  assign \new_[3045]_  = \new_[3044]_  | \new_[3041]_ ;
  assign \new_[3046]_  = \new_[3045]_  | \new_[3038]_ ;
  assign \new_[3050]_  = \new_[1100]_  | \new_[1101]_ ;
  assign \new_[3051]_  = \new_[1102]_  | \new_[3050]_ ;
  assign \new_[3054]_  = \new_[1098]_  | \new_[1099]_ ;
  assign \new_[3057]_  = \new_[1096]_  | \new_[1097]_ ;
  assign \new_[3058]_  = \new_[3057]_  | \new_[3054]_ ;
  assign \new_[3059]_  = \new_[3058]_  | \new_[3051]_ ;
  assign \new_[3060]_  = \new_[3059]_  | \new_[3046]_ ;
  assign \new_[3061]_  = \new_[3060]_  | \new_[3033]_ ;
  assign \new_[3062]_  = \new_[3061]_  | \new_[3006]_ ;
  assign \new_[3063]_  = \new_[3062]_  | \new_[2953]_ ;
  assign \new_[3064]_  = \new_[3063]_  | \new_[2844]_ ;
  assign \new_[3068]_  = \new_[1093]_  | \new_[1094]_ ;
  assign \new_[3069]_  = \new_[1095]_  | \new_[3068]_ ;
  assign \new_[3073]_  = \new_[1090]_  | \new_[1091]_ ;
  assign \new_[3074]_  = \new_[1092]_  | \new_[3073]_ ;
  assign \new_[3075]_  = \new_[3074]_  | \new_[3069]_ ;
  assign \new_[3079]_  = \new_[1087]_  | \new_[1088]_ ;
  assign \new_[3080]_  = \new_[1089]_  | \new_[3079]_ ;
  assign \new_[3083]_  = \new_[1085]_  | \new_[1086]_ ;
  assign \new_[3086]_  = \new_[1083]_  | \new_[1084]_ ;
  assign \new_[3087]_  = \new_[3086]_  | \new_[3083]_ ;
  assign \new_[3088]_  = \new_[3087]_  | \new_[3080]_ ;
  assign \new_[3089]_  = \new_[3088]_  | \new_[3075]_ ;
  assign \new_[3093]_  = \new_[1080]_  | \new_[1081]_ ;
  assign \new_[3094]_  = \new_[1082]_  | \new_[3093]_ ;
  assign \new_[3097]_  = \new_[1078]_  | \new_[1079]_ ;
  assign \new_[3100]_  = \new_[1076]_  | \new_[1077]_ ;
  assign \new_[3101]_  = \new_[3100]_  | \new_[3097]_ ;
  assign \new_[3102]_  = \new_[3101]_  | \new_[3094]_ ;
  assign \new_[3106]_  = \new_[1073]_  | \new_[1074]_ ;
  assign \new_[3107]_  = \new_[1075]_  | \new_[3106]_ ;
  assign \new_[3110]_  = \new_[1071]_  | \new_[1072]_ ;
  assign \new_[3113]_  = \new_[1069]_  | \new_[1070]_ ;
  assign \new_[3114]_  = \new_[3113]_  | \new_[3110]_ ;
  assign \new_[3115]_  = \new_[3114]_  | \new_[3107]_ ;
  assign \new_[3116]_  = \new_[3115]_  | \new_[3102]_ ;
  assign \new_[3117]_  = \new_[3116]_  | \new_[3089]_ ;
  assign \new_[3121]_  = \new_[1066]_  | \new_[1067]_ ;
  assign \new_[3122]_  = \new_[1068]_  | \new_[3121]_ ;
  assign \new_[3126]_  = \new_[1063]_  | \new_[1064]_ ;
  assign \new_[3127]_  = \new_[1065]_  | \new_[3126]_ ;
  assign \new_[3128]_  = \new_[3127]_  | \new_[3122]_ ;
  assign \new_[3132]_  = \new_[1060]_  | \new_[1061]_ ;
  assign \new_[3133]_  = \new_[1062]_  | \new_[3132]_ ;
  assign \new_[3136]_  = \new_[1058]_  | \new_[1059]_ ;
  assign \new_[3139]_  = \new_[1056]_  | \new_[1057]_ ;
  assign \new_[3140]_  = \new_[3139]_  | \new_[3136]_ ;
  assign \new_[3141]_  = \new_[3140]_  | \new_[3133]_ ;
  assign \new_[3142]_  = \new_[3141]_  | \new_[3128]_ ;
  assign \new_[3146]_  = \new_[1053]_  | \new_[1054]_ ;
  assign \new_[3147]_  = \new_[1055]_  | \new_[3146]_ ;
  assign \new_[3150]_  = \new_[1051]_  | \new_[1052]_ ;
  assign \new_[3153]_  = \new_[1049]_  | \new_[1050]_ ;
  assign \new_[3154]_  = \new_[3153]_  | \new_[3150]_ ;
  assign \new_[3155]_  = \new_[3154]_  | \new_[3147]_ ;
  assign \new_[3159]_  = \new_[1046]_  | \new_[1047]_ ;
  assign \new_[3160]_  = \new_[1048]_  | \new_[3159]_ ;
  assign \new_[3163]_  = \new_[1044]_  | \new_[1045]_ ;
  assign \new_[3166]_  = \new_[1042]_  | \new_[1043]_ ;
  assign \new_[3167]_  = \new_[3166]_  | \new_[3163]_ ;
  assign \new_[3168]_  = \new_[3167]_  | \new_[3160]_ ;
  assign \new_[3169]_  = \new_[3168]_  | \new_[3155]_ ;
  assign \new_[3170]_  = \new_[3169]_  | \new_[3142]_ ;
  assign \new_[3171]_  = \new_[3170]_  | \new_[3117]_ ;
  assign \new_[3175]_  = \new_[1039]_  | \new_[1040]_ ;
  assign \new_[3176]_  = \new_[1041]_  | \new_[3175]_ ;
  assign \new_[3180]_  = \new_[1036]_  | \new_[1037]_ ;
  assign \new_[3181]_  = \new_[1038]_  | \new_[3180]_ ;
  assign \new_[3182]_  = \new_[3181]_  | \new_[3176]_ ;
  assign \new_[3186]_  = \new_[1033]_  | \new_[1034]_ ;
  assign \new_[3187]_  = \new_[1035]_  | \new_[3186]_ ;
  assign \new_[3190]_  = \new_[1031]_  | \new_[1032]_ ;
  assign \new_[3193]_  = \new_[1029]_  | \new_[1030]_ ;
  assign \new_[3194]_  = \new_[3193]_  | \new_[3190]_ ;
  assign \new_[3195]_  = \new_[3194]_  | \new_[3187]_ ;
  assign \new_[3196]_  = \new_[3195]_  | \new_[3182]_ ;
  assign \new_[3200]_  = \new_[1026]_  | \new_[1027]_ ;
  assign \new_[3201]_  = \new_[1028]_  | \new_[3200]_ ;
  assign \new_[3204]_  = \new_[1024]_  | \new_[1025]_ ;
  assign \new_[3207]_  = \new_[1022]_  | \new_[1023]_ ;
  assign \new_[3208]_  = \new_[3207]_  | \new_[3204]_ ;
  assign \new_[3209]_  = \new_[3208]_  | \new_[3201]_ ;
  assign \new_[3213]_  = \new_[1019]_  | \new_[1020]_ ;
  assign \new_[3214]_  = \new_[1021]_  | \new_[3213]_ ;
  assign \new_[3217]_  = \new_[1017]_  | \new_[1018]_ ;
  assign \new_[3220]_  = \new_[1015]_  | \new_[1016]_ ;
  assign \new_[3221]_  = \new_[3220]_  | \new_[3217]_ ;
  assign \new_[3222]_  = \new_[3221]_  | \new_[3214]_ ;
  assign \new_[3223]_  = \new_[3222]_  | \new_[3209]_ ;
  assign \new_[3224]_  = \new_[3223]_  | \new_[3196]_ ;
  assign \new_[3228]_  = \new_[1012]_  | \new_[1013]_ ;
  assign \new_[3229]_  = \new_[1014]_  | \new_[3228]_ ;
  assign \new_[3232]_  = \new_[1010]_  | \new_[1011]_ ;
  assign \new_[3235]_  = \new_[1008]_  | \new_[1009]_ ;
  assign \new_[3236]_  = \new_[3235]_  | \new_[3232]_ ;
  assign \new_[3237]_  = \new_[3236]_  | \new_[3229]_ ;
  assign \new_[3241]_  = \new_[1005]_  | \new_[1006]_ ;
  assign \new_[3242]_  = \new_[1007]_  | \new_[3241]_ ;
  assign \new_[3245]_  = \new_[1003]_  | \new_[1004]_ ;
  assign \new_[3248]_  = \new_[1001]_  | \new_[1002]_ ;
  assign \new_[3249]_  = \new_[3248]_  | \new_[3245]_ ;
  assign \new_[3250]_  = \new_[3249]_  | \new_[3242]_ ;
  assign \new_[3251]_  = \new_[3250]_  | \new_[3237]_ ;
  assign \new_[3255]_  = \new_[998]_  | \new_[999]_ ;
  assign \new_[3256]_  = \new_[1000]_  | \new_[3255]_ ;
  assign \new_[3259]_  = \new_[996]_  | \new_[997]_ ;
  assign \new_[3262]_  = \new_[994]_  | \new_[995]_ ;
  assign \new_[3263]_  = \new_[3262]_  | \new_[3259]_ ;
  assign \new_[3264]_  = \new_[3263]_  | \new_[3256]_ ;
  assign \new_[3268]_  = \new_[991]_  | \new_[992]_ ;
  assign \new_[3269]_  = \new_[993]_  | \new_[3268]_ ;
  assign \new_[3272]_  = \new_[989]_  | \new_[990]_ ;
  assign \new_[3275]_  = \new_[987]_  | \new_[988]_ ;
  assign \new_[3276]_  = \new_[3275]_  | \new_[3272]_ ;
  assign \new_[3277]_  = \new_[3276]_  | \new_[3269]_ ;
  assign \new_[3278]_  = \new_[3277]_  | \new_[3264]_ ;
  assign \new_[3279]_  = \new_[3278]_  | \new_[3251]_ ;
  assign \new_[3280]_  = \new_[3279]_  | \new_[3224]_ ;
  assign \new_[3281]_  = \new_[3280]_  | \new_[3171]_ ;
  assign \new_[3285]_  = \new_[984]_  | \new_[985]_ ;
  assign \new_[3286]_  = \new_[986]_  | \new_[3285]_ ;
  assign \new_[3290]_  = \new_[981]_  | \new_[982]_ ;
  assign \new_[3291]_  = \new_[983]_  | \new_[3290]_ ;
  assign \new_[3292]_  = \new_[3291]_  | \new_[3286]_ ;
  assign \new_[3296]_  = \new_[978]_  | \new_[979]_ ;
  assign \new_[3297]_  = \new_[980]_  | \new_[3296]_ ;
  assign \new_[3300]_  = \new_[976]_  | \new_[977]_ ;
  assign \new_[3303]_  = \new_[974]_  | \new_[975]_ ;
  assign \new_[3304]_  = \new_[3303]_  | \new_[3300]_ ;
  assign \new_[3305]_  = \new_[3304]_  | \new_[3297]_ ;
  assign \new_[3306]_  = \new_[3305]_  | \new_[3292]_ ;
  assign \new_[3310]_  = \new_[971]_  | \new_[972]_ ;
  assign \new_[3311]_  = \new_[973]_  | \new_[3310]_ ;
  assign \new_[3314]_  = \new_[969]_  | \new_[970]_ ;
  assign \new_[3317]_  = \new_[967]_  | \new_[968]_ ;
  assign \new_[3318]_  = \new_[3317]_  | \new_[3314]_ ;
  assign \new_[3319]_  = \new_[3318]_  | \new_[3311]_ ;
  assign \new_[3323]_  = \new_[964]_  | \new_[965]_ ;
  assign \new_[3324]_  = \new_[966]_  | \new_[3323]_ ;
  assign \new_[3327]_  = \new_[962]_  | \new_[963]_ ;
  assign \new_[3330]_  = \new_[960]_  | \new_[961]_ ;
  assign \new_[3331]_  = \new_[3330]_  | \new_[3327]_ ;
  assign \new_[3332]_  = \new_[3331]_  | \new_[3324]_ ;
  assign \new_[3333]_  = \new_[3332]_  | \new_[3319]_ ;
  assign \new_[3334]_  = \new_[3333]_  | \new_[3306]_ ;
  assign \new_[3338]_  = \new_[957]_  | \new_[958]_ ;
  assign \new_[3339]_  = \new_[959]_  | \new_[3338]_ ;
  assign \new_[3342]_  = \new_[955]_  | \new_[956]_ ;
  assign \new_[3345]_  = \new_[953]_  | \new_[954]_ ;
  assign \new_[3346]_  = \new_[3345]_  | \new_[3342]_ ;
  assign \new_[3347]_  = \new_[3346]_  | \new_[3339]_ ;
  assign \new_[3351]_  = \new_[950]_  | \new_[951]_ ;
  assign \new_[3352]_  = \new_[952]_  | \new_[3351]_ ;
  assign \new_[3355]_  = \new_[948]_  | \new_[949]_ ;
  assign \new_[3358]_  = \new_[946]_  | \new_[947]_ ;
  assign \new_[3359]_  = \new_[3358]_  | \new_[3355]_ ;
  assign \new_[3360]_  = \new_[3359]_  | \new_[3352]_ ;
  assign \new_[3361]_  = \new_[3360]_  | \new_[3347]_ ;
  assign \new_[3365]_  = \new_[943]_  | \new_[944]_ ;
  assign \new_[3366]_  = \new_[945]_  | \new_[3365]_ ;
  assign \new_[3369]_  = \new_[941]_  | \new_[942]_ ;
  assign \new_[3372]_  = \new_[939]_  | \new_[940]_ ;
  assign \new_[3373]_  = \new_[3372]_  | \new_[3369]_ ;
  assign \new_[3374]_  = \new_[3373]_  | \new_[3366]_ ;
  assign \new_[3378]_  = \new_[936]_  | \new_[937]_ ;
  assign \new_[3379]_  = \new_[938]_  | \new_[3378]_ ;
  assign \new_[3382]_  = \new_[934]_  | \new_[935]_ ;
  assign \new_[3385]_  = \new_[932]_  | \new_[933]_ ;
  assign \new_[3386]_  = \new_[3385]_  | \new_[3382]_ ;
  assign \new_[3387]_  = \new_[3386]_  | \new_[3379]_ ;
  assign \new_[3388]_  = \new_[3387]_  | \new_[3374]_ ;
  assign \new_[3389]_  = \new_[3388]_  | \new_[3361]_ ;
  assign \new_[3390]_  = \new_[3389]_  | \new_[3334]_ ;
  assign \new_[3394]_  = \new_[929]_  | \new_[930]_ ;
  assign \new_[3395]_  = \new_[931]_  | \new_[3394]_ ;
  assign \new_[3399]_  = \new_[926]_  | \new_[927]_ ;
  assign \new_[3400]_  = \new_[928]_  | \new_[3399]_ ;
  assign \new_[3401]_  = \new_[3400]_  | \new_[3395]_ ;
  assign \new_[3405]_  = \new_[923]_  | \new_[924]_ ;
  assign \new_[3406]_  = \new_[925]_  | \new_[3405]_ ;
  assign \new_[3409]_  = \new_[921]_  | \new_[922]_ ;
  assign \new_[3412]_  = \new_[919]_  | \new_[920]_ ;
  assign \new_[3413]_  = \new_[3412]_  | \new_[3409]_ ;
  assign \new_[3414]_  = \new_[3413]_  | \new_[3406]_ ;
  assign \new_[3415]_  = \new_[3414]_  | \new_[3401]_ ;
  assign \new_[3419]_  = \new_[916]_  | \new_[917]_ ;
  assign \new_[3420]_  = \new_[918]_  | \new_[3419]_ ;
  assign \new_[3423]_  = \new_[914]_  | \new_[915]_ ;
  assign \new_[3426]_  = \new_[912]_  | \new_[913]_ ;
  assign \new_[3427]_  = \new_[3426]_  | \new_[3423]_ ;
  assign \new_[3428]_  = \new_[3427]_  | \new_[3420]_ ;
  assign \new_[3432]_  = \new_[909]_  | \new_[910]_ ;
  assign \new_[3433]_  = \new_[911]_  | \new_[3432]_ ;
  assign \new_[3436]_  = \new_[907]_  | \new_[908]_ ;
  assign \new_[3439]_  = \new_[905]_  | \new_[906]_ ;
  assign \new_[3440]_  = \new_[3439]_  | \new_[3436]_ ;
  assign \new_[3441]_  = \new_[3440]_  | \new_[3433]_ ;
  assign \new_[3442]_  = \new_[3441]_  | \new_[3428]_ ;
  assign \new_[3443]_  = \new_[3442]_  | \new_[3415]_ ;
  assign \new_[3447]_  = \new_[902]_  | \new_[903]_ ;
  assign \new_[3448]_  = \new_[904]_  | \new_[3447]_ ;
  assign \new_[3451]_  = \new_[900]_  | \new_[901]_ ;
  assign \new_[3454]_  = \new_[898]_  | \new_[899]_ ;
  assign \new_[3455]_  = \new_[3454]_  | \new_[3451]_ ;
  assign \new_[3456]_  = \new_[3455]_  | \new_[3448]_ ;
  assign \new_[3460]_  = \new_[895]_  | \new_[896]_ ;
  assign \new_[3461]_  = \new_[897]_  | \new_[3460]_ ;
  assign \new_[3464]_  = \new_[893]_  | \new_[894]_ ;
  assign \new_[3467]_  = \new_[891]_  | \new_[892]_ ;
  assign \new_[3468]_  = \new_[3467]_  | \new_[3464]_ ;
  assign \new_[3469]_  = \new_[3468]_  | \new_[3461]_ ;
  assign \new_[3470]_  = \new_[3469]_  | \new_[3456]_ ;
  assign \new_[3474]_  = \new_[888]_  | \new_[889]_ ;
  assign \new_[3475]_  = \new_[890]_  | \new_[3474]_ ;
  assign \new_[3478]_  = \new_[886]_  | \new_[887]_ ;
  assign \new_[3481]_  = \new_[884]_  | \new_[885]_ ;
  assign \new_[3482]_  = \new_[3481]_  | \new_[3478]_ ;
  assign \new_[3483]_  = \new_[3482]_  | \new_[3475]_ ;
  assign \new_[3487]_  = \new_[881]_  | \new_[882]_ ;
  assign \new_[3488]_  = \new_[883]_  | \new_[3487]_ ;
  assign \new_[3491]_  = \new_[879]_  | \new_[880]_ ;
  assign \new_[3494]_  = \new_[877]_  | \new_[878]_ ;
  assign \new_[3495]_  = \new_[3494]_  | \new_[3491]_ ;
  assign \new_[3496]_  = \new_[3495]_  | \new_[3488]_ ;
  assign \new_[3497]_  = \new_[3496]_  | \new_[3483]_ ;
  assign \new_[3498]_  = \new_[3497]_  | \new_[3470]_ ;
  assign \new_[3499]_  = \new_[3498]_  | \new_[3443]_ ;
  assign \new_[3500]_  = \new_[3499]_  | \new_[3390]_ ;
  assign \new_[3501]_  = \new_[3500]_  | \new_[3281]_ ;
  assign \new_[3502]_  = \new_[3501]_  | \new_[3064]_ ;
  assign \new_[3503]_  = \new_[3502]_  | \new_[2627]_ ;
  assign \new_[3507]_  = \new_[874]_  | \new_[875]_ ;
  assign \new_[3508]_  = \new_[876]_  | \new_[3507]_ ;
  assign \new_[3512]_  = \new_[871]_  | \new_[872]_ ;
  assign \new_[3513]_  = \new_[873]_  | \new_[3512]_ ;
  assign \new_[3514]_  = \new_[3513]_  | \new_[3508]_ ;
  assign \new_[3518]_  = \new_[868]_  | \new_[869]_ ;
  assign \new_[3519]_  = \new_[870]_  | \new_[3518]_ ;
  assign \new_[3522]_  = \new_[866]_  | \new_[867]_ ;
  assign \new_[3525]_  = \new_[864]_  | \new_[865]_ ;
  assign \new_[3526]_  = \new_[3525]_  | \new_[3522]_ ;
  assign \new_[3527]_  = \new_[3526]_  | \new_[3519]_ ;
  assign \new_[3528]_  = \new_[3527]_  | \new_[3514]_ ;
  assign \new_[3532]_  = \new_[861]_  | \new_[862]_ ;
  assign \new_[3533]_  = \new_[863]_  | \new_[3532]_ ;
  assign \new_[3536]_  = \new_[859]_  | \new_[860]_ ;
  assign \new_[3539]_  = \new_[857]_  | \new_[858]_ ;
  assign \new_[3540]_  = \new_[3539]_  | \new_[3536]_ ;
  assign \new_[3541]_  = \new_[3540]_  | \new_[3533]_ ;
  assign \new_[3545]_  = \new_[854]_  | \new_[855]_ ;
  assign \new_[3546]_  = \new_[856]_  | \new_[3545]_ ;
  assign \new_[3549]_  = \new_[852]_  | \new_[853]_ ;
  assign \new_[3552]_  = \new_[850]_  | \new_[851]_ ;
  assign \new_[3553]_  = \new_[3552]_  | \new_[3549]_ ;
  assign \new_[3554]_  = \new_[3553]_  | \new_[3546]_ ;
  assign \new_[3555]_  = \new_[3554]_  | \new_[3541]_ ;
  assign \new_[3556]_  = \new_[3555]_  | \new_[3528]_ ;
  assign \new_[3560]_  = \new_[847]_  | \new_[848]_ ;
  assign \new_[3561]_  = \new_[849]_  | \new_[3560]_ ;
  assign \new_[3565]_  = \new_[844]_  | \new_[845]_ ;
  assign \new_[3566]_  = \new_[846]_  | \new_[3565]_ ;
  assign \new_[3567]_  = \new_[3566]_  | \new_[3561]_ ;
  assign \new_[3571]_  = \new_[841]_  | \new_[842]_ ;
  assign \new_[3572]_  = \new_[843]_  | \new_[3571]_ ;
  assign \new_[3575]_  = \new_[839]_  | \new_[840]_ ;
  assign \new_[3578]_  = \new_[837]_  | \new_[838]_ ;
  assign \new_[3579]_  = \new_[3578]_  | \new_[3575]_ ;
  assign \new_[3580]_  = \new_[3579]_  | \new_[3572]_ ;
  assign \new_[3581]_  = \new_[3580]_  | \new_[3567]_ ;
  assign \new_[3585]_  = \new_[834]_  | \new_[835]_ ;
  assign \new_[3586]_  = \new_[836]_  | \new_[3585]_ ;
  assign \new_[3589]_  = \new_[832]_  | \new_[833]_ ;
  assign \new_[3592]_  = \new_[830]_  | \new_[831]_ ;
  assign \new_[3593]_  = \new_[3592]_  | \new_[3589]_ ;
  assign \new_[3594]_  = \new_[3593]_  | \new_[3586]_ ;
  assign \new_[3598]_  = \new_[827]_  | \new_[828]_ ;
  assign \new_[3599]_  = \new_[829]_  | \new_[3598]_ ;
  assign \new_[3602]_  = \new_[825]_  | \new_[826]_ ;
  assign \new_[3605]_  = \new_[823]_  | \new_[824]_ ;
  assign \new_[3606]_  = \new_[3605]_  | \new_[3602]_ ;
  assign \new_[3607]_  = \new_[3606]_  | \new_[3599]_ ;
  assign \new_[3608]_  = \new_[3607]_  | \new_[3594]_ ;
  assign \new_[3609]_  = \new_[3608]_  | \new_[3581]_ ;
  assign \new_[3610]_  = \new_[3609]_  | \new_[3556]_ ;
  assign \new_[3614]_  = \new_[820]_  | \new_[821]_ ;
  assign \new_[3615]_  = \new_[822]_  | \new_[3614]_ ;
  assign \new_[3619]_  = \new_[817]_  | \new_[818]_ ;
  assign \new_[3620]_  = \new_[819]_  | \new_[3619]_ ;
  assign \new_[3621]_  = \new_[3620]_  | \new_[3615]_ ;
  assign \new_[3625]_  = \new_[814]_  | \new_[815]_ ;
  assign \new_[3626]_  = \new_[816]_  | \new_[3625]_ ;
  assign \new_[3629]_  = \new_[812]_  | \new_[813]_ ;
  assign \new_[3632]_  = \new_[810]_  | \new_[811]_ ;
  assign \new_[3633]_  = \new_[3632]_  | \new_[3629]_ ;
  assign \new_[3634]_  = \new_[3633]_  | \new_[3626]_ ;
  assign \new_[3635]_  = \new_[3634]_  | \new_[3621]_ ;
  assign \new_[3639]_  = \new_[807]_  | \new_[808]_ ;
  assign \new_[3640]_  = \new_[809]_  | \new_[3639]_ ;
  assign \new_[3643]_  = \new_[805]_  | \new_[806]_ ;
  assign \new_[3646]_  = \new_[803]_  | \new_[804]_ ;
  assign \new_[3647]_  = \new_[3646]_  | \new_[3643]_ ;
  assign \new_[3648]_  = \new_[3647]_  | \new_[3640]_ ;
  assign \new_[3652]_  = \new_[800]_  | \new_[801]_ ;
  assign \new_[3653]_  = \new_[802]_  | \new_[3652]_ ;
  assign \new_[3656]_  = \new_[798]_  | \new_[799]_ ;
  assign \new_[3659]_  = \new_[796]_  | \new_[797]_ ;
  assign \new_[3660]_  = \new_[3659]_  | \new_[3656]_ ;
  assign \new_[3661]_  = \new_[3660]_  | \new_[3653]_ ;
  assign \new_[3662]_  = \new_[3661]_  | \new_[3648]_ ;
  assign \new_[3663]_  = \new_[3662]_  | \new_[3635]_ ;
  assign \new_[3667]_  = \new_[793]_  | \new_[794]_ ;
  assign \new_[3668]_  = \new_[795]_  | \new_[3667]_ ;
  assign \new_[3671]_  = \new_[791]_  | \new_[792]_ ;
  assign \new_[3674]_  = \new_[789]_  | \new_[790]_ ;
  assign \new_[3675]_  = \new_[3674]_  | \new_[3671]_ ;
  assign \new_[3676]_  = \new_[3675]_  | \new_[3668]_ ;
  assign \new_[3680]_  = \new_[786]_  | \new_[787]_ ;
  assign \new_[3681]_  = \new_[788]_  | \new_[3680]_ ;
  assign \new_[3684]_  = \new_[784]_  | \new_[785]_ ;
  assign \new_[3687]_  = \new_[782]_  | \new_[783]_ ;
  assign \new_[3688]_  = \new_[3687]_  | \new_[3684]_ ;
  assign \new_[3689]_  = \new_[3688]_  | \new_[3681]_ ;
  assign \new_[3690]_  = \new_[3689]_  | \new_[3676]_ ;
  assign \new_[3694]_  = \new_[779]_  | \new_[780]_ ;
  assign \new_[3695]_  = \new_[781]_  | \new_[3694]_ ;
  assign \new_[3698]_  = \new_[777]_  | \new_[778]_ ;
  assign \new_[3701]_  = \new_[775]_  | \new_[776]_ ;
  assign \new_[3702]_  = \new_[3701]_  | \new_[3698]_ ;
  assign \new_[3703]_  = \new_[3702]_  | \new_[3695]_ ;
  assign \new_[3707]_  = \new_[772]_  | \new_[773]_ ;
  assign \new_[3708]_  = \new_[774]_  | \new_[3707]_ ;
  assign \new_[3711]_  = \new_[770]_  | \new_[771]_ ;
  assign \new_[3714]_  = \new_[768]_  | \new_[769]_ ;
  assign \new_[3715]_  = \new_[3714]_  | \new_[3711]_ ;
  assign \new_[3716]_  = \new_[3715]_  | \new_[3708]_ ;
  assign \new_[3717]_  = \new_[3716]_  | \new_[3703]_ ;
  assign \new_[3718]_  = \new_[3717]_  | \new_[3690]_ ;
  assign \new_[3719]_  = \new_[3718]_  | \new_[3663]_ ;
  assign \new_[3720]_  = \new_[3719]_  | \new_[3610]_ ;
  assign \new_[3724]_  = \new_[765]_  | \new_[766]_ ;
  assign \new_[3725]_  = \new_[767]_  | \new_[3724]_ ;
  assign \new_[3729]_  = \new_[762]_  | \new_[763]_ ;
  assign \new_[3730]_  = \new_[764]_  | \new_[3729]_ ;
  assign \new_[3731]_  = \new_[3730]_  | \new_[3725]_ ;
  assign \new_[3735]_  = \new_[759]_  | \new_[760]_ ;
  assign \new_[3736]_  = \new_[761]_  | \new_[3735]_ ;
  assign \new_[3739]_  = \new_[757]_  | \new_[758]_ ;
  assign \new_[3742]_  = \new_[755]_  | \new_[756]_ ;
  assign \new_[3743]_  = \new_[3742]_  | \new_[3739]_ ;
  assign \new_[3744]_  = \new_[3743]_  | \new_[3736]_ ;
  assign \new_[3745]_  = \new_[3744]_  | \new_[3731]_ ;
  assign \new_[3749]_  = \new_[752]_  | \new_[753]_ ;
  assign \new_[3750]_  = \new_[754]_  | \new_[3749]_ ;
  assign \new_[3753]_  = \new_[750]_  | \new_[751]_ ;
  assign \new_[3756]_  = \new_[748]_  | \new_[749]_ ;
  assign \new_[3757]_  = \new_[3756]_  | \new_[3753]_ ;
  assign \new_[3758]_  = \new_[3757]_  | \new_[3750]_ ;
  assign \new_[3762]_  = \new_[745]_  | \new_[746]_ ;
  assign \new_[3763]_  = \new_[747]_  | \new_[3762]_ ;
  assign \new_[3766]_  = \new_[743]_  | \new_[744]_ ;
  assign \new_[3769]_  = \new_[741]_  | \new_[742]_ ;
  assign \new_[3770]_  = \new_[3769]_  | \new_[3766]_ ;
  assign \new_[3771]_  = \new_[3770]_  | \new_[3763]_ ;
  assign \new_[3772]_  = \new_[3771]_  | \new_[3758]_ ;
  assign \new_[3773]_  = \new_[3772]_  | \new_[3745]_ ;
  assign \new_[3777]_  = \new_[738]_  | \new_[739]_ ;
  assign \new_[3778]_  = \new_[740]_  | \new_[3777]_ ;
  assign \new_[3781]_  = \new_[736]_  | \new_[737]_ ;
  assign \new_[3784]_  = \new_[734]_  | \new_[735]_ ;
  assign \new_[3785]_  = \new_[3784]_  | \new_[3781]_ ;
  assign \new_[3786]_  = \new_[3785]_  | \new_[3778]_ ;
  assign \new_[3790]_  = \new_[731]_  | \new_[732]_ ;
  assign \new_[3791]_  = \new_[733]_  | \new_[3790]_ ;
  assign \new_[3794]_  = \new_[729]_  | \new_[730]_ ;
  assign \new_[3797]_  = \new_[727]_  | \new_[728]_ ;
  assign \new_[3798]_  = \new_[3797]_  | \new_[3794]_ ;
  assign \new_[3799]_  = \new_[3798]_  | \new_[3791]_ ;
  assign \new_[3800]_  = \new_[3799]_  | \new_[3786]_ ;
  assign \new_[3804]_  = \new_[724]_  | \new_[725]_ ;
  assign \new_[3805]_  = \new_[726]_  | \new_[3804]_ ;
  assign \new_[3808]_  = \new_[722]_  | \new_[723]_ ;
  assign \new_[3811]_  = \new_[720]_  | \new_[721]_ ;
  assign \new_[3812]_  = \new_[3811]_  | \new_[3808]_ ;
  assign \new_[3813]_  = \new_[3812]_  | \new_[3805]_ ;
  assign \new_[3817]_  = \new_[717]_  | \new_[718]_ ;
  assign \new_[3818]_  = \new_[719]_  | \new_[3817]_ ;
  assign \new_[3821]_  = \new_[715]_  | \new_[716]_ ;
  assign \new_[3824]_  = \new_[713]_  | \new_[714]_ ;
  assign \new_[3825]_  = \new_[3824]_  | \new_[3821]_ ;
  assign \new_[3826]_  = \new_[3825]_  | \new_[3818]_ ;
  assign \new_[3827]_  = \new_[3826]_  | \new_[3813]_ ;
  assign \new_[3828]_  = \new_[3827]_  | \new_[3800]_ ;
  assign \new_[3829]_  = \new_[3828]_  | \new_[3773]_ ;
  assign \new_[3833]_  = \new_[710]_  | \new_[711]_ ;
  assign \new_[3834]_  = \new_[712]_  | \new_[3833]_ ;
  assign \new_[3838]_  = \new_[707]_  | \new_[708]_ ;
  assign \new_[3839]_  = \new_[709]_  | \new_[3838]_ ;
  assign \new_[3840]_  = \new_[3839]_  | \new_[3834]_ ;
  assign \new_[3844]_  = \new_[704]_  | \new_[705]_ ;
  assign \new_[3845]_  = \new_[706]_  | \new_[3844]_ ;
  assign \new_[3848]_  = \new_[702]_  | \new_[703]_ ;
  assign \new_[3851]_  = \new_[700]_  | \new_[701]_ ;
  assign \new_[3852]_  = \new_[3851]_  | \new_[3848]_ ;
  assign \new_[3853]_  = \new_[3852]_  | \new_[3845]_ ;
  assign \new_[3854]_  = \new_[3853]_  | \new_[3840]_ ;
  assign \new_[3858]_  = \new_[697]_  | \new_[698]_ ;
  assign \new_[3859]_  = \new_[699]_  | \new_[3858]_ ;
  assign \new_[3862]_  = \new_[695]_  | \new_[696]_ ;
  assign \new_[3865]_  = \new_[693]_  | \new_[694]_ ;
  assign \new_[3866]_  = \new_[3865]_  | \new_[3862]_ ;
  assign \new_[3867]_  = \new_[3866]_  | \new_[3859]_ ;
  assign \new_[3871]_  = \new_[690]_  | \new_[691]_ ;
  assign \new_[3872]_  = \new_[692]_  | \new_[3871]_ ;
  assign \new_[3875]_  = \new_[688]_  | \new_[689]_ ;
  assign \new_[3878]_  = \new_[686]_  | \new_[687]_ ;
  assign \new_[3879]_  = \new_[3878]_  | \new_[3875]_ ;
  assign \new_[3880]_  = \new_[3879]_  | \new_[3872]_ ;
  assign \new_[3881]_  = \new_[3880]_  | \new_[3867]_ ;
  assign \new_[3882]_  = \new_[3881]_  | \new_[3854]_ ;
  assign \new_[3886]_  = \new_[683]_  | \new_[684]_ ;
  assign \new_[3887]_  = \new_[685]_  | \new_[3886]_ ;
  assign \new_[3890]_  = \new_[681]_  | \new_[682]_ ;
  assign \new_[3893]_  = \new_[679]_  | \new_[680]_ ;
  assign \new_[3894]_  = \new_[3893]_  | \new_[3890]_ ;
  assign \new_[3895]_  = \new_[3894]_  | \new_[3887]_ ;
  assign \new_[3899]_  = \new_[676]_  | \new_[677]_ ;
  assign \new_[3900]_  = \new_[678]_  | \new_[3899]_ ;
  assign \new_[3903]_  = \new_[674]_  | \new_[675]_ ;
  assign \new_[3906]_  = \new_[672]_  | \new_[673]_ ;
  assign \new_[3907]_  = \new_[3906]_  | \new_[3903]_ ;
  assign \new_[3908]_  = \new_[3907]_  | \new_[3900]_ ;
  assign \new_[3909]_  = \new_[3908]_  | \new_[3895]_ ;
  assign \new_[3913]_  = \new_[669]_  | \new_[670]_ ;
  assign \new_[3914]_  = \new_[671]_  | \new_[3913]_ ;
  assign \new_[3917]_  = \new_[667]_  | \new_[668]_ ;
  assign \new_[3920]_  = \new_[665]_  | \new_[666]_ ;
  assign \new_[3921]_  = \new_[3920]_  | \new_[3917]_ ;
  assign \new_[3922]_  = \new_[3921]_  | \new_[3914]_ ;
  assign \new_[3926]_  = \new_[662]_  | \new_[663]_ ;
  assign \new_[3927]_  = \new_[664]_  | \new_[3926]_ ;
  assign \new_[3930]_  = \new_[660]_  | \new_[661]_ ;
  assign \new_[3933]_  = \new_[658]_  | \new_[659]_ ;
  assign \new_[3934]_  = \new_[3933]_  | \new_[3930]_ ;
  assign \new_[3935]_  = \new_[3934]_  | \new_[3927]_ ;
  assign \new_[3936]_  = \new_[3935]_  | \new_[3922]_ ;
  assign \new_[3937]_  = \new_[3936]_  | \new_[3909]_ ;
  assign \new_[3938]_  = \new_[3937]_  | \new_[3882]_ ;
  assign \new_[3939]_  = \new_[3938]_  | \new_[3829]_ ;
  assign \new_[3940]_  = \new_[3939]_  | \new_[3720]_ ;
  assign \new_[3944]_  = \new_[655]_  | \new_[656]_ ;
  assign \new_[3945]_  = \new_[657]_  | \new_[3944]_ ;
  assign \new_[3949]_  = \new_[652]_  | \new_[653]_ ;
  assign \new_[3950]_  = \new_[654]_  | \new_[3949]_ ;
  assign \new_[3951]_  = \new_[3950]_  | \new_[3945]_ ;
  assign \new_[3955]_  = \new_[649]_  | \new_[650]_ ;
  assign \new_[3956]_  = \new_[651]_  | \new_[3955]_ ;
  assign \new_[3959]_  = \new_[647]_  | \new_[648]_ ;
  assign \new_[3962]_  = \new_[645]_  | \new_[646]_ ;
  assign \new_[3963]_  = \new_[3962]_  | \new_[3959]_ ;
  assign \new_[3964]_  = \new_[3963]_  | \new_[3956]_ ;
  assign \new_[3965]_  = \new_[3964]_  | \new_[3951]_ ;
  assign \new_[3969]_  = \new_[642]_  | \new_[643]_ ;
  assign \new_[3970]_  = \new_[644]_  | \new_[3969]_ ;
  assign \new_[3973]_  = \new_[640]_  | \new_[641]_ ;
  assign \new_[3976]_  = \new_[638]_  | \new_[639]_ ;
  assign \new_[3977]_  = \new_[3976]_  | \new_[3973]_ ;
  assign \new_[3978]_  = \new_[3977]_  | \new_[3970]_ ;
  assign \new_[3982]_  = \new_[635]_  | \new_[636]_ ;
  assign \new_[3983]_  = \new_[637]_  | \new_[3982]_ ;
  assign \new_[3986]_  = \new_[633]_  | \new_[634]_ ;
  assign \new_[3989]_  = \new_[631]_  | \new_[632]_ ;
  assign \new_[3990]_  = \new_[3989]_  | \new_[3986]_ ;
  assign \new_[3991]_  = \new_[3990]_  | \new_[3983]_ ;
  assign \new_[3992]_  = \new_[3991]_  | \new_[3978]_ ;
  assign \new_[3993]_  = \new_[3992]_  | \new_[3965]_ ;
  assign \new_[3997]_  = \new_[628]_  | \new_[629]_ ;
  assign \new_[3998]_  = \new_[630]_  | \new_[3997]_ ;
  assign \new_[4002]_  = \new_[625]_  | \new_[626]_ ;
  assign \new_[4003]_  = \new_[627]_  | \new_[4002]_ ;
  assign \new_[4004]_  = \new_[4003]_  | \new_[3998]_ ;
  assign \new_[4008]_  = \new_[622]_  | \new_[623]_ ;
  assign \new_[4009]_  = \new_[624]_  | \new_[4008]_ ;
  assign \new_[4012]_  = \new_[620]_  | \new_[621]_ ;
  assign \new_[4015]_  = \new_[618]_  | \new_[619]_ ;
  assign \new_[4016]_  = \new_[4015]_  | \new_[4012]_ ;
  assign \new_[4017]_  = \new_[4016]_  | \new_[4009]_ ;
  assign \new_[4018]_  = \new_[4017]_  | \new_[4004]_ ;
  assign \new_[4022]_  = \new_[615]_  | \new_[616]_ ;
  assign \new_[4023]_  = \new_[617]_  | \new_[4022]_ ;
  assign \new_[4026]_  = \new_[613]_  | \new_[614]_ ;
  assign \new_[4029]_  = \new_[611]_  | \new_[612]_ ;
  assign \new_[4030]_  = \new_[4029]_  | \new_[4026]_ ;
  assign \new_[4031]_  = \new_[4030]_  | \new_[4023]_ ;
  assign \new_[4035]_  = \new_[608]_  | \new_[609]_ ;
  assign \new_[4036]_  = \new_[610]_  | \new_[4035]_ ;
  assign \new_[4039]_  = \new_[606]_  | \new_[607]_ ;
  assign \new_[4042]_  = \new_[604]_  | \new_[605]_ ;
  assign \new_[4043]_  = \new_[4042]_  | \new_[4039]_ ;
  assign \new_[4044]_  = \new_[4043]_  | \new_[4036]_ ;
  assign \new_[4045]_  = \new_[4044]_  | \new_[4031]_ ;
  assign \new_[4046]_  = \new_[4045]_  | \new_[4018]_ ;
  assign \new_[4047]_  = \new_[4046]_  | \new_[3993]_ ;
  assign \new_[4051]_  = \new_[601]_  | \new_[602]_ ;
  assign \new_[4052]_  = \new_[603]_  | \new_[4051]_ ;
  assign \new_[4056]_  = \new_[598]_  | \new_[599]_ ;
  assign \new_[4057]_  = \new_[600]_  | \new_[4056]_ ;
  assign \new_[4058]_  = \new_[4057]_  | \new_[4052]_ ;
  assign \new_[4062]_  = \new_[595]_  | \new_[596]_ ;
  assign \new_[4063]_  = \new_[597]_  | \new_[4062]_ ;
  assign \new_[4066]_  = \new_[593]_  | \new_[594]_ ;
  assign \new_[4069]_  = \new_[591]_  | \new_[592]_ ;
  assign \new_[4070]_  = \new_[4069]_  | \new_[4066]_ ;
  assign \new_[4071]_  = \new_[4070]_  | \new_[4063]_ ;
  assign \new_[4072]_  = \new_[4071]_  | \new_[4058]_ ;
  assign \new_[4076]_  = \new_[588]_  | \new_[589]_ ;
  assign \new_[4077]_  = \new_[590]_  | \new_[4076]_ ;
  assign \new_[4080]_  = \new_[586]_  | \new_[587]_ ;
  assign \new_[4083]_  = \new_[584]_  | \new_[585]_ ;
  assign \new_[4084]_  = \new_[4083]_  | \new_[4080]_ ;
  assign \new_[4085]_  = \new_[4084]_  | \new_[4077]_ ;
  assign \new_[4089]_  = \new_[581]_  | \new_[582]_ ;
  assign \new_[4090]_  = \new_[583]_  | \new_[4089]_ ;
  assign \new_[4093]_  = \new_[579]_  | \new_[580]_ ;
  assign \new_[4096]_  = \new_[577]_  | \new_[578]_ ;
  assign \new_[4097]_  = \new_[4096]_  | \new_[4093]_ ;
  assign \new_[4098]_  = \new_[4097]_  | \new_[4090]_ ;
  assign \new_[4099]_  = \new_[4098]_  | \new_[4085]_ ;
  assign \new_[4100]_  = \new_[4099]_  | \new_[4072]_ ;
  assign \new_[4104]_  = \new_[574]_  | \new_[575]_ ;
  assign \new_[4105]_  = \new_[576]_  | \new_[4104]_ ;
  assign \new_[4108]_  = \new_[572]_  | \new_[573]_ ;
  assign \new_[4111]_  = \new_[570]_  | \new_[571]_ ;
  assign \new_[4112]_  = \new_[4111]_  | \new_[4108]_ ;
  assign \new_[4113]_  = \new_[4112]_  | \new_[4105]_ ;
  assign \new_[4117]_  = \new_[567]_  | \new_[568]_ ;
  assign \new_[4118]_  = \new_[569]_  | \new_[4117]_ ;
  assign \new_[4121]_  = \new_[565]_  | \new_[566]_ ;
  assign \new_[4124]_  = \new_[563]_  | \new_[564]_ ;
  assign \new_[4125]_  = \new_[4124]_  | \new_[4121]_ ;
  assign \new_[4126]_  = \new_[4125]_  | \new_[4118]_ ;
  assign \new_[4127]_  = \new_[4126]_  | \new_[4113]_ ;
  assign \new_[4131]_  = \new_[560]_  | \new_[561]_ ;
  assign \new_[4132]_  = \new_[562]_  | \new_[4131]_ ;
  assign \new_[4135]_  = \new_[558]_  | \new_[559]_ ;
  assign \new_[4138]_  = \new_[556]_  | \new_[557]_ ;
  assign \new_[4139]_  = \new_[4138]_  | \new_[4135]_ ;
  assign \new_[4140]_  = \new_[4139]_  | \new_[4132]_ ;
  assign \new_[4144]_  = \new_[553]_  | \new_[554]_ ;
  assign \new_[4145]_  = \new_[555]_  | \new_[4144]_ ;
  assign \new_[4148]_  = \new_[551]_  | \new_[552]_ ;
  assign \new_[4151]_  = \new_[549]_  | \new_[550]_ ;
  assign \new_[4152]_  = \new_[4151]_  | \new_[4148]_ ;
  assign \new_[4153]_  = \new_[4152]_  | \new_[4145]_ ;
  assign \new_[4154]_  = \new_[4153]_  | \new_[4140]_ ;
  assign \new_[4155]_  = \new_[4154]_  | \new_[4127]_ ;
  assign \new_[4156]_  = \new_[4155]_  | \new_[4100]_ ;
  assign \new_[4157]_  = \new_[4156]_  | \new_[4047]_ ;
  assign \new_[4161]_  = \new_[546]_  | \new_[547]_ ;
  assign \new_[4162]_  = \new_[548]_  | \new_[4161]_ ;
  assign \new_[4166]_  = \new_[543]_  | \new_[544]_ ;
  assign \new_[4167]_  = \new_[545]_  | \new_[4166]_ ;
  assign \new_[4168]_  = \new_[4167]_  | \new_[4162]_ ;
  assign \new_[4172]_  = \new_[540]_  | \new_[541]_ ;
  assign \new_[4173]_  = \new_[542]_  | \new_[4172]_ ;
  assign \new_[4176]_  = \new_[538]_  | \new_[539]_ ;
  assign \new_[4179]_  = \new_[536]_  | \new_[537]_ ;
  assign \new_[4180]_  = \new_[4179]_  | \new_[4176]_ ;
  assign \new_[4181]_  = \new_[4180]_  | \new_[4173]_ ;
  assign \new_[4182]_  = \new_[4181]_  | \new_[4168]_ ;
  assign \new_[4186]_  = \new_[533]_  | \new_[534]_ ;
  assign \new_[4187]_  = \new_[535]_  | \new_[4186]_ ;
  assign \new_[4190]_  = \new_[531]_  | \new_[532]_ ;
  assign \new_[4193]_  = \new_[529]_  | \new_[530]_ ;
  assign \new_[4194]_  = \new_[4193]_  | \new_[4190]_ ;
  assign \new_[4195]_  = \new_[4194]_  | \new_[4187]_ ;
  assign \new_[4199]_  = \new_[526]_  | \new_[527]_ ;
  assign \new_[4200]_  = \new_[528]_  | \new_[4199]_ ;
  assign \new_[4203]_  = \new_[524]_  | \new_[525]_ ;
  assign \new_[4206]_  = \new_[522]_  | \new_[523]_ ;
  assign \new_[4207]_  = \new_[4206]_  | \new_[4203]_ ;
  assign \new_[4208]_  = \new_[4207]_  | \new_[4200]_ ;
  assign \new_[4209]_  = \new_[4208]_  | \new_[4195]_ ;
  assign \new_[4210]_  = \new_[4209]_  | \new_[4182]_ ;
  assign \new_[4214]_  = \new_[519]_  | \new_[520]_ ;
  assign \new_[4215]_  = \new_[521]_  | \new_[4214]_ ;
  assign \new_[4218]_  = \new_[517]_  | \new_[518]_ ;
  assign \new_[4221]_  = \new_[515]_  | \new_[516]_ ;
  assign \new_[4222]_  = \new_[4221]_  | \new_[4218]_ ;
  assign \new_[4223]_  = \new_[4222]_  | \new_[4215]_ ;
  assign \new_[4227]_  = \new_[512]_  | \new_[513]_ ;
  assign \new_[4228]_  = \new_[514]_  | \new_[4227]_ ;
  assign \new_[4231]_  = \new_[510]_  | \new_[511]_ ;
  assign \new_[4234]_  = \new_[508]_  | \new_[509]_ ;
  assign \new_[4235]_  = \new_[4234]_  | \new_[4231]_ ;
  assign \new_[4236]_  = \new_[4235]_  | \new_[4228]_ ;
  assign \new_[4237]_  = \new_[4236]_  | \new_[4223]_ ;
  assign \new_[4241]_  = \new_[505]_  | \new_[506]_ ;
  assign \new_[4242]_  = \new_[507]_  | \new_[4241]_ ;
  assign \new_[4245]_  = \new_[503]_  | \new_[504]_ ;
  assign \new_[4248]_  = \new_[501]_  | \new_[502]_ ;
  assign \new_[4249]_  = \new_[4248]_  | \new_[4245]_ ;
  assign \new_[4250]_  = \new_[4249]_  | \new_[4242]_ ;
  assign \new_[4254]_  = \new_[498]_  | \new_[499]_ ;
  assign \new_[4255]_  = \new_[500]_  | \new_[4254]_ ;
  assign \new_[4258]_  = \new_[496]_  | \new_[497]_ ;
  assign \new_[4261]_  = \new_[494]_  | \new_[495]_ ;
  assign \new_[4262]_  = \new_[4261]_  | \new_[4258]_ ;
  assign \new_[4263]_  = \new_[4262]_  | \new_[4255]_ ;
  assign \new_[4264]_  = \new_[4263]_  | \new_[4250]_ ;
  assign \new_[4265]_  = \new_[4264]_  | \new_[4237]_ ;
  assign \new_[4266]_  = \new_[4265]_  | \new_[4210]_ ;
  assign \new_[4270]_  = \new_[491]_  | \new_[492]_ ;
  assign \new_[4271]_  = \new_[493]_  | \new_[4270]_ ;
  assign \new_[4275]_  = \new_[488]_  | \new_[489]_ ;
  assign \new_[4276]_  = \new_[490]_  | \new_[4275]_ ;
  assign \new_[4277]_  = \new_[4276]_  | \new_[4271]_ ;
  assign \new_[4281]_  = \new_[485]_  | \new_[486]_ ;
  assign \new_[4282]_  = \new_[487]_  | \new_[4281]_ ;
  assign \new_[4285]_  = \new_[483]_  | \new_[484]_ ;
  assign \new_[4288]_  = \new_[481]_  | \new_[482]_ ;
  assign \new_[4289]_  = \new_[4288]_  | \new_[4285]_ ;
  assign \new_[4290]_  = \new_[4289]_  | \new_[4282]_ ;
  assign \new_[4291]_  = \new_[4290]_  | \new_[4277]_ ;
  assign \new_[4295]_  = \new_[478]_  | \new_[479]_ ;
  assign \new_[4296]_  = \new_[480]_  | \new_[4295]_ ;
  assign \new_[4299]_  = \new_[476]_  | \new_[477]_ ;
  assign \new_[4302]_  = \new_[474]_  | \new_[475]_ ;
  assign \new_[4303]_  = \new_[4302]_  | \new_[4299]_ ;
  assign \new_[4304]_  = \new_[4303]_  | \new_[4296]_ ;
  assign \new_[4308]_  = \new_[471]_  | \new_[472]_ ;
  assign \new_[4309]_  = \new_[473]_  | \new_[4308]_ ;
  assign \new_[4312]_  = \new_[469]_  | \new_[470]_ ;
  assign \new_[4315]_  = \new_[467]_  | \new_[468]_ ;
  assign \new_[4316]_  = \new_[4315]_  | \new_[4312]_ ;
  assign \new_[4317]_  = \new_[4316]_  | \new_[4309]_ ;
  assign \new_[4318]_  = \new_[4317]_  | \new_[4304]_ ;
  assign \new_[4319]_  = \new_[4318]_  | \new_[4291]_ ;
  assign \new_[4323]_  = \new_[464]_  | \new_[465]_ ;
  assign \new_[4324]_  = \new_[466]_  | \new_[4323]_ ;
  assign \new_[4327]_  = \new_[462]_  | \new_[463]_ ;
  assign \new_[4330]_  = \new_[460]_  | \new_[461]_ ;
  assign \new_[4331]_  = \new_[4330]_  | \new_[4327]_ ;
  assign \new_[4332]_  = \new_[4331]_  | \new_[4324]_ ;
  assign \new_[4336]_  = \new_[457]_  | \new_[458]_ ;
  assign \new_[4337]_  = \new_[459]_  | \new_[4336]_ ;
  assign \new_[4340]_  = \new_[455]_  | \new_[456]_ ;
  assign \new_[4343]_  = \new_[453]_  | \new_[454]_ ;
  assign \new_[4344]_  = \new_[4343]_  | \new_[4340]_ ;
  assign \new_[4345]_  = \new_[4344]_  | \new_[4337]_ ;
  assign \new_[4346]_  = \new_[4345]_  | \new_[4332]_ ;
  assign \new_[4350]_  = \new_[450]_  | \new_[451]_ ;
  assign \new_[4351]_  = \new_[452]_  | \new_[4350]_ ;
  assign \new_[4354]_  = \new_[448]_  | \new_[449]_ ;
  assign \new_[4357]_  = \new_[446]_  | \new_[447]_ ;
  assign \new_[4358]_  = \new_[4357]_  | \new_[4354]_ ;
  assign \new_[4359]_  = \new_[4358]_  | \new_[4351]_ ;
  assign \new_[4363]_  = \new_[443]_  | \new_[444]_ ;
  assign \new_[4364]_  = \new_[445]_  | \new_[4363]_ ;
  assign \new_[4367]_  = \new_[441]_  | \new_[442]_ ;
  assign \new_[4370]_  = \new_[439]_  | \new_[440]_ ;
  assign \new_[4371]_  = \new_[4370]_  | \new_[4367]_ ;
  assign \new_[4372]_  = \new_[4371]_  | \new_[4364]_ ;
  assign \new_[4373]_  = \new_[4372]_  | \new_[4359]_ ;
  assign \new_[4374]_  = \new_[4373]_  | \new_[4346]_ ;
  assign \new_[4375]_  = \new_[4374]_  | \new_[4319]_ ;
  assign \new_[4376]_  = \new_[4375]_  | \new_[4266]_ ;
  assign \new_[4377]_  = \new_[4376]_  | \new_[4157]_ ;
  assign \new_[4378]_  = \new_[4377]_  | \new_[3940]_ ;
  assign \new_[4382]_  = \new_[436]_  | \new_[437]_ ;
  assign \new_[4383]_  = \new_[438]_  | \new_[4382]_ ;
  assign \new_[4387]_  = \new_[433]_  | \new_[434]_ ;
  assign \new_[4388]_  = \new_[435]_  | \new_[4387]_ ;
  assign \new_[4389]_  = \new_[4388]_  | \new_[4383]_ ;
  assign \new_[4393]_  = \new_[430]_  | \new_[431]_ ;
  assign \new_[4394]_  = \new_[432]_  | \new_[4393]_ ;
  assign \new_[4397]_  = \new_[428]_  | \new_[429]_ ;
  assign \new_[4400]_  = \new_[426]_  | \new_[427]_ ;
  assign \new_[4401]_  = \new_[4400]_  | \new_[4397]_ ;
  assign \new_[4402]_  = \new_[4401]_  | \new_[4394]_ ;
  assign \new_[4403]_  = \new_[4402]_  | \new_[4389]_ ;
  assign \new_[4407]_  = \new_[423]_  | \new_[424]_ ;
  assign \new_[4408]_  = \new_[425]_  | \new_[4407]_ ;
  assign \new_[4411]_  = \new_[421]_  | \new_[422]_ ;
  assign \new_[4414]_  = \new_[419]_  | \new_[420]_ ;
  assign \new_[4415]_  = \new_[4414]_  | \new_[4411]_ ;
  assign \new_[4416]_  = \new_[4415]_  | \new_[4408]_ ;
  assign \new_[4420]_  = \new_[416]_  | \new_[417]_ ;
  assign \new_[4421]_  = \new_[418]_  | \new_[4420]_ ;
  assign \new_[4424]_  = \new_[414]_  | \new_[415]_ ;
  assign \new_[4427]_  = \new_[412]_  | \new_[413]_ ;
  assign \new_[4428]_  = \new_[4427]_  | \new_[4424]_ ;
  assign \new_[4429]_  = \new_[4428]_  | \new_[4421]_ ;
  assign \new_[4430]_  = \new_[4429]_  | \new_[4416]_ ;
  assign \new_[4431]_  = \new_[4430]_  | \new_[4403]_ ;
  assign \new_[4435]_  = \new_[409]_  | \new_[410]_ ;
  assign \new_[4436]_  = \new_[411]_  | \new_[4435]_ ;
  assign \new_[4440]_  = \new_[406]_  | \new_[407]_ ;
  assign \new_[4441]_  = \new_[408]_  | \new_[4440]_ ;
  assign \new_[4442]_  = \new_[4441]_  | \new_[4436]_ ;
  assign \new_[4446]_  = \new_[403]_  | \new_[404]_ ;
  assign \new_[4447]_  = \new_[405]_  | \new_[4446]_ ;
  assign \new_[4450]_  = \new_[401]_  | \new_[402]_ ;
  assign \new_[4453]_  = \new_[399]_  | \new_[400]_ ;
  assign \new_[4454]_  = \new_[4453]_  | \new_[4450]_ ;
  assign \new_[4455]_  = \new_[4454]_  | \new_[4447]_ ;
  assign \new_[4456]_  = \new_[4455]_  | \new_[4442]_ ;
  assign \new_[4460]_  = \new_[396]_  | \new_[397]_ ;
  assign \new_[4461]_  = \new_[398]_  | \new_[4460]_ ;
  assign \new_[4464]_  = \new_[394]_  | \new_[395]_ ;
  assign \new_[4467]_  = \new_[392]_  | \new_[393]_ ;
  assign \new_[4468]_  = \new_[4467]_  | \new_[4464]_ ;
  assign \new_[4469]_  = \new_[4468]_  | \new_[4461]_ ;
  assign \new_[4473]_  = \new_[389]_  | \new_[390]_ ;
  assign \new_[4474]_  = \new_[391]_  | \new_[4473]_ ;
  assign \new_[4477]_  = \new_[387]_  | \new_[388]_ ;
  assign \new_[4480]_  = \new_[385]_  | \new_[386]_ ;
  assign \new_[4481]_  = \new_[4480]_  | \new_[4477]_ ;
  assign \new_[4482]_  = \new_[4481]_  | \new_[4474]_ ;
  assign \new_[4483]_  = \new_[4482]_  | \new_[4469]_ ;
  assign \new_[4484]_  = \new_[4483]_  | \new_[4456]_ ;
  assign \new_[4485]_  = \new_[4484]_  | \new_[4431]_ ;
  assign \new_[4489]_  = \new_[382]_  | \new_[383]_ ;
  assign \new_[4490]_  = \new_[384]_  | \new_[4489]_ ;
  assign \new_[4494]_  = \new_[379]_  | \new_[380]_ ;
  assign \new_[4495]_  = \new_[381]_  | \new_[4494]_ ;
  assign \new_[4496]_  = \new_[4495]_  | \new_[4490]_ ;
  assign \new_[4500]_  = \new_[376]_  | \new_[377]_ ;
  assign \new_[4501]_  = \new_[378]_  | \new_[4500]_ ;
  assign \new_[4504]_  = \new_[374]_  | \new_[375]_ ;
  assign \new_[4507]_  = \new_[372]_  | \new_[373]_ ;
  assign \new_[4508]_  = \new_[4507]_  | \new_[4504]_ ;
  assign \new_[4509]_  = \new_[4508]_  | \new_[4501]_ ;
  assign \new_[4510]_  = \new_[4509]_  | \new_[4496]_ ;
  assign \new_[4514]_  = \new_[369]_  | \new_[370]_ ;
  assign \new_[4515]_  = \new_[371]_  | \new_[4514]_ ;
  assign \new_[4518]_  = \new_[367]_  | \new_[368]_ ;
  assign \new_[4521]_  = \new_[365]_  | \new_[366]_ ;
  assign \new_[4522]_  = \new_[4521]_  | \new_[4518]_ ;
  assign \new_[4523]_  = \new_[4522]_  | \new_[4515]_ ;
  assign \new_[4527]_  = \new_[362]_  | \new_[363]_ ;
  assign \new_[4528]_  = \new_[364]_  | \new_[4527]_ ;
  assign \new_[4531]_  = \new_[360]_  | \new_[361]_ ;
  assign \new_[4534]_  = \new_[358]_  | \new_[359]_ ;
  assign \new_[4535]_  = \new_[4534]_  | \new_[4531]_ ;
  assign \new_[4536]_  = \new_[4535]_  | \new_[4528]_ ;
  assign \new_[4537]_  = \new_[4536]_  | \new_[4523]_ ;
  assign \new_[4538]_  = \new_[4537]_  | \new_[4510]_ ;
  assign \new_[4542]_  = \new_[355]_  | \new_[356]_ ;
  assign \new_[4543]_  = \new_[357]_  | \new_[4542]_ ;
  assign \new_[4546]_  = \new_[353]_  | \new_[354]_ ;
  assign \new_[4549]_  = \new_[351]_  | \new_[352]_ ;
  assign \new_[4550]_  = \new_[4549]_  | \new_[4546]_ ;
  assign \new_[4551]_  = \new_[4550]_  | \new_[4543]_ ;
  assign \new_[4555]_  = \new_[348]_  | \new_[349]_ ;
  assign \new_[4556]_  = \new_[350]_  | \new_[4555]_ ;
  assign \new_[4559]_  = \new_[346]_  | \new_[347]_ ;
  assign \new_[4562]_  = \new_[344]_  | \new_[345]_ ;
  assign \new_[4563]_  = \new_[4562]_  | \new_[4559]_ ;
  assign \new_[4564]_  = \new_[4563]_  | \new_[4556]_ ;
  assign \new_[4565]_  = \new_[4564]_  | \new_[4551]_ ;
  assign \new_[4569]_  = \new_[341]_  | \new_[342]_ ;
  assign \new_[4570]_  = \new_[343]_  | \new_[4569]_ ;
  assign \new_[4573]_  = \new_[339]_  | \new_[340]_ ;
  assign \new_[4576]_  = \new_[337]_  | \new_[338]_ ;
  assign \new_[4577]_  = \new_[4576]_  | \new_[4573]_ ;
  assign \new_[4578]_  = \new_[4577]_  | \new_[4570]_ ;
  assign \new_[4582]_  = \new_[334]_  | \new_[335]_ ;
  assign \new_[4583]_  = \new_[336]_  | \new_[4582]_ ;
  assign \new_[4586]_  = \new_[332]_  | \new_[333]_ ;
  assign \new_[4589]_  = \new_[330]_  | \new_[331]_ ;
  assign \new_[4590]_  = \new_[4589]_  | \new_[4586]_ ;
  assign \new_[4591]_  = \new_[4590]_  | \new_[4583]_ ;
  assign \new_[4592]_  = \new_[4591]_  | \new_[4578]_ ;
  assign \new_[4593]_  = \new_[4592]_  | \new_[4565]_ ;
  assign \new_[4594]_  = \new_[4593]_  | \new_[4538]_ ;
  assign \new_[4595]_  = \new_[4594]_  | \new_[4485]_ ;
  assign \new_[4599]_  = \new_[327]_  | \new_[328]_ ;
  assign \new_[4600]_  = \new_[329]_  | \new_[4599]_ ;
  assign \new_[4604]_  = \new_[324]_  | \new_[325]_ ;
  assign \new_[4605]_  = \new_[326]_  | \new_[4604]_ ;
  assign \new_[4606]_  = \new_[4605]_  | \new_[4600]_ ;
  assign \new_[4610]_  = \new_[321]_  | \new_[322]_ ;
  assign \new_[4611]_  = \new_[323]_  | \new_[4610]_ ;
  assign \new_[4614]_  = \new_[319]_  | \new_[320]_ ;
  assign \new_[4617]_  = \new_[317]_  | \new_[318]_ ;
  assign \new_[4618]_  = \new_[4617]_  | \new_[4614]_ ;
  assign \new_[4619]_  = \new_[4618]_  | \new_[4611]_ ;
  assign \new_[4620]_  = \new_[4619]_  | \new_[4606]_ ;
  assign \new_[4624]_  = \new_[314]_  | \new_[315]_ ;
  assign \new_[4625]_  = \new_[316]_  | \new_[4624]_ ;
  assign \new_[4628]_  = \new_[312]_  | \new_[313]_ ;
  assign \new_[4631]_  = \new_[310]_  | \new_[311]_ ;
  assign \new_[4632]_  = \new_[4631]_  | \new_[4628]_ ;
  assign \new_[4633]_  = \new_[4632]_  | \new_[4625]_ ;
  assign \new_[4637]_  = \new_[307]_  | \new_[308]_ ;
  assign \new_[4638]_  = \new_[309]_  | \new_[4637]_ ;
  assign \new_[4641]_  = \new_[305]_  | \new_[306]_ ;
  assign \new_[4644]_  = \new_[303]_  | \new_[304]_ ;
  assign \new_[4645]_  = \new_[4644]_  | \new_[4641]_ ;
  assign \new_[4646]_  = \new_[4645]_  | \new_[4638]_ ;
  assign \new_[4647]_  = \new_[4646]_  | \new_[4633]_ ;
  assign \new_[4648]_  = \new_[4647]_  | \new_[4620]_ ;
  assign \new_[4652]_  = \new_[300]_  | \new_[301]_ ;
  assign \new_[4653]_  = \new_[302]_  | \new_[4652]_ ;
  assign \new_[4656]_  = \new_[298]_  | \new_[299]_ ;
  assign \new_[4659]_  = \new_[296]_  | \new_[297]_ ;
  assign \new_[4660]_  = \new_[4659]_  | \new_[4656]_ ;
  assign \new_[4661]_  = \new_[4660]_  | \new_[4653]_ ;
  assign \new_[4665]_  = \new_[293]_  | \new_[294]_ ;
  assign \new_[4666]_  = \new_[295]_  | \new_[4665]_ ;
  assign \new_[4669]_  = \new_[291]_  | \new_[292]_ ;
  assign \new_[4672]_  = \new_[289]_  | \new_[290]_ ;
  assign \new_[4673]_  = \new_[4672]_  | \new_[4669]_ ;
  assign \new_[4674]_  = \new_[4673]_  | \new_[4666]_ ;
  assign \new_[4675]_  = \new_[4674]_  | \new_[4661]_ ;
  assign \new_[4679]_  = \new_[286]_  | \new_[287]_ ;
  assign \new_[4680]_  = \new_[288]_  | \new_[4679]_ ;
  assign \new_[4683]_  = \new_[284]_  | \new_[285]_ ;
  assign \new_[4686]_  = \new_[282]_  | \new_[283]_ ;
  assign \new_[4687]_  = \new_[4686]_  | \new_[4683]_ ;
  assign \new_[4688]_  = \new_[4687]_  | \new_[4680]_ ;
  assign \new_[4692]_  = \new_[279]_  | \new_[280]_ ;
  assign \new_[4693]_  = \new_[281]_  | \new_[4692]_ ;
  assign \new_[4696]_  = \new_[277]_  | \new_[278]_ ;
  assign \new_[4699]_  = \new_[275]_  | \new_[276]_ ;
  assign \new_[4700]_  = \new_[4699]_  | \new_[4696]_ ;
  assign \new_[4701]_  = \new_[4700]_  | \new_[4693]_ ;
  assign \new_[4702]_  = \new_[4701]_  | \new_[4688]_ ;
  assign \new_[4703]_  = \new_[4702]_  | \new_[4675]_ ;
  assign \new_[4704]_  = \new_[4703]_  | \new_[4648]_ ;
  assign \new_[4708]_  = \new_[272]_  | \new_[273]_ ;
  assign \new_[4709]_  = \new_[274]_  | \new_[4708]_ ;
  assign \new_[4713]_  = \new_[269]_  | \new_[270]_ ;
  assign \new_[4714]_  = \new_[271]_  | \new_[4713]_ ;
  assign \new_[4715]_  = \new_[4714]_  | \new_[4709]_ ;
  assign \new_[4719]_  = \new_[266]_  | \new_[267]_ ;
  assign \new_[4720]_  = \new_[268]_  | \new_[4719]_ ;
  assign \new_[4723]_  = \new_[264]_  | \new_[265]_ ;
  assign \new_[4726]_  = \new_[262]_  | \new_[263]_ ;
  assign \new_[4727]_  = \new_[4726]_  | \new_[4723]_ ;
  assign \new_[4728]_  = \new_[4727]_  | \new_[4720]_ ;
  assign \new_[4729]_  = \new_[4728]_  | \new_[4715]_ ;
  assign \new_[4733]_  = \new_[259]_  | \new_[260]_ ;
  assign \new_[4734]_  = \new_[261]_  | \new_[4733]_ ;
  assign \new_[4737]_  = \new_[257]_  | \new_[258]_ ;
  assign \new_[4740]_  = \new_[255]_  | \new_[256]_ ;
  assign \new_[4741]_  = \new_[4740]_  | \new_[4737]_ ;
  assign \new_[4742]_  = \new_[4741]_  | \new_[4734]_ ;
  assign \new_[4746]_  = \new_[252]_  | \new_[253]_ ;
  assign \new_[4747]_  = \new_[254]_  | \new_[4746]_ ;
  assign \new_[4750]_  = \new_[250]_  | \new_[251]_ ;
  assign \new_[4753]_  = \new_[248]_  | \new_[249]_ ;
  assign \new_[4754]_  = \new_[4753]_  | \new_[4750]_ ;
  assign \new_[4755]_  = \new_[4754]_  | \new_[4747]_ ;
  assign \new_[4756]_  = \new_[4755]_  | \new_[4742]_ ;
  assign \new_[4757]_  = \new_[4756]_  | \new_[4729]_ ;
  assign \new_[4761]_  = \new_[245]_  | \new_[246]_ ;
  assign \new_[4762]_  = \new_[247]_  | \new_[4761]_ ;
  assign \new_[4765]_  = \new_[243]_  | \new_[244]_ ;
  assign \new_[4768]_  = \new_[241]_  | \new_[242]_ ;
  assign \new_[4769]_  = \new_[4768]_  | \new_[4765]_ ;
  assign \new_[4770]_  = \new_[4769]_  | \new_[4762]_ ;
  assign \new_[4774]_  = \new_[238]_  | \new_[239]_ ;
  assign \new_[4775]_  = \new_[240]_  | \new_[4774]_ ;
  assign \new_[4778]_  = \new_[236]_  | \new_[237]_ ;
  assign \new_[4781]_  = \new_[234]_  | \new_[235]_ ;
  assign \new_[4782]_  = \new_[4781]_  | \new_[4778]_ ;
  assign \new_[4783]_  = \new_[4782]_  | \new_[4775]_ ;
  assign \new_[4784]_  = \new_[4783]_  | \new_[4770]_ ;
  assign \new_[4788]_  = \new_[231]_  | \new_[232]_ ;
  assign \new_[4789]_  = \new_[233]_  | \new_[4788]_ ;
  assign \new_[4792]_  = \new_[229]_  | \new_[230]_ ;
  assign \new_[4795]_  = \new_[227]_  | \new_[228]_ ;
  assign \new_[4796]_  = \new_[4795]_  | \new_[4792]_ ;
  assign \new_[4797]_  = \new_[4796]_  | \new_[4789]_ ;
  assign \new_[4801]_  = \new_[224]_  | \new_[225]_ ;
  assign \new_[4802]_  = \new_[226]_  | \new_[4801]_ ;
  assign \new_[4805]_  = \new_[222]_  | \new_[223]_ ;
  assign \new_[4808]_  = \new_[220]_  | \new_[221]_ ;
  assign \new_[4809]_  = \new_[4808]_  | \new_[4805]_ ;
  assign \new_[4810]_  = \new_[4809]_  | \new_[4802]_ ;
  assign \new_[4811]_  = \new_[4810]_  | \new_[4797]_ ;
  assign \new_[4812]_  = \new_[4811]_  | \new_[4784]_ ;
  assign \new_[4813]_  = \new_[4812]_  | \new_[4757]_ ;
  assign \new_[4814]_  = \new_[4813]_  | \new_[4704]_ ;
  assign \new_[4815]_  = \new_[4814]_  | \new_[4595]_ ;
  assign \new_[4819]_  = \new_[217]_  | \new_[218]_ ;
  assign \new_[4820]_  = \new_[219]_  | \new_[4819]_ ;
  assign \new_[4824]_  = \new_[214]_  | \new_[215]_ ;
  assign \new_[4825]_  = \new_[216]_  | \new_[4824]_ ;
  assign \new_[4826]_  = \new_[4825]_  | \new_[4820]_ ;
  assign \new_[4830]_  = \new_[211]_  | \new_[212]_ ;
  assign \new_[4831]_  = \new_[213]_  | \new_[4830]_ ;
  assign \new_[4834]_  = \new_[209]_  | \new_[210]_ ;
  assign \new_[4837]_  = \new_[207]_  | \new_[208]_ ;
  assign \new_[4838]_  = \new_[4837]_  | \new_[4834]_ ;
  assign \new_[4839]_  = \new_[4838]_  | \new_[4831]_ ;
  assign \new_[4840]_  = \new_[4839]_  | \new_[4826]_ ;
  assign \new_[4844]_  = \new_[204]_  | \new_[205]_ ;
  assign \new_[4845]_  = \new_[206]_  | \new_[4844]_ ;
  assign \new_[4848]_  = \new_[202]_  | \new_[203]_ ;
  assign \new_[4851]_  = \new_[200]_  | \new_[201]_ ;
  assign \new_[4852]_  = \new_[4851]_  | \new_[4848]_ ;
  assign \new_[4853]_  = \new_[4852]_  | \new_[4845]_ ;
  assign \new_[4857]_  = \new_[197]_  | \new_[198]_ ;
  assign \new_[4858]_  = \new_[199]_  | \new_[4857]_ ;
  assign \new_[4861]_  = \new_[195]_  | \new_[196]_ ;
  assign \new_[4864]_  = \new_[193]_  | \new_[194]_ ;
  assign \new_[4865]_  = \new_[4864]_  | \new_[4861]_ ;
  assign \new_[4866]_  = \new_[4865]_  | \new_[4858]_ ;
  assign \new_[4867]_  = \new_[4866]_  | \new_[4853]_ ;
  assign \new_[4868]_  = \new_[4867]_  | \new_[4840]_ ;
  assign \new_[4872]_  = \new_[190]_  | \new_[191]_ ;
  assign \new_[4873]_  = \new_[192]_  | \new_[4872]_ ;
  assign \new_[4877]_  = \new_[187]_  | \new_[188]_ ;
  assign \new_[4878]_  = \new_[189]_  | \new_[4877]_ ;
  assign \new_[4879]_  = \new_[4878]_  | \new_[4873]_ ;
  assign \new_[4883]_  = \new_[184]_  | \new_[185]_ ;
  assign \new_[4884]_  = \new_[186]_  | \new_[4883]_ ;
  assign \new_[4887]_  = \new_[182]_  | \new_[183]_ ;
  assign \new_[4890]_  = \new_[180]_  | \new_[181]_ ;
  assign \new_[4891]_  = \new_[4890]_  | \new_[4887]_ ;
  assign \new_[4892]_  = \new_[4891]_  | \new_[4884]_ ;
  assign \new_[4893]_  = \new_[4892]_  | \new_[4879]_ ;
  assign \new_[4897]_  = \new_[177]_  | \new_[178]_ ;
  assign \new_[4898]_  = \new_[179]_  | \new_[4897]_ ;
  assign \new_[4901]_  = \new_[175]_  | \new_[176]_ ;
  assign \new_[4904]_  = \new_[173]_  | \new_[174]_ ;
  assign \new_[4905]_  = \new_[4904]_  | \new_[4901]_ ;
  assign \new_[4906]_  = \new_[4905]_  | \new_[4898]_ ;
  assign \new_[4910]_  = \new_[170]_  | \new_[171]_ ;
  assign \new_[4911]_  = \new_[172]_  | \new_[4910]_ ;
  assign \new_[4914]_  = \new_[168]_  | \new_[169]_ ;
  assign \new_[4917]_  = \new_[166]_  | \new_[167]_ ;
  assign \new_[4918]_  = \new_[4917]_  | \new_[4914]_ ;
  assign \new_[4919]_  = \new_[4918]_  | \new_[4911]_ ;
  assign \new_[4920]_  = \new_[4919]_  | \new_[4906]_ ;
  assign \new_[4921]_  = \new_[4920]_  | \new_[4893]_ ;
  assign \new_[4922]_  = \new_[4921]_  | \new_[4868]_ ;
  assign \new_[4926]_  = \new_[163]_  | \new_[164]_ ;
  assign \new_[4927]_  = \new_[165]_  | \new_[4926]_ ;
  assign \new_[4931]_  = \new_[160]_  | \new_[161]_ ;
  assign \new_[4932]_  = \new_[162]_  | \new_[4931]_ ;
  assign \new_[4933]_  = \new_[4932]_  | \new_[4927]_ ;
  assign \new_[4937]_  = \new_[157]_  | \new_[158]_ ;
  assign \new_[4938]_  = \new_[159]_  | \new_[4937]_ ;
  assign \new_[4941]_  = \new_[155]_  | \new_[156]_ ;
  assign \new_[4944]_  = \new_[153]_  | \new_[154]_ ;
  assign \new_[4945]_  = \new_[4944]_  | \new_[4941]_ ;
  assign \new_[4946]_  = \new_[4945]_  | \new_[4938]_ ;
  assign \new_[4947]_  = \new_[4946]_  | \new_[4933]_ ;
  assign \new_[4951]_  = \new_[150]_  | \new_[151]_ ;
  assign \new_[4952]_  = \new_[152]_  | \new_[4951]_ ;
  assign \new_[4955]_  = \new_[148]_  | \new_[149]_ ;
  assign \new_[4958]_  = \new_[146]_  | \new_[147]_ ;
  assign \new_[4959]_  = \new_[4958]_  | \new_[4955]_ ;
  assign \new_[4960]_  = \new_[4959]_  | \new_[4952]_ ;
  assign \new_[4964]_  = \new_[143]_  | \new_[144]_ ;
  assign \new_[4965]_  = \new_[145]_  | \new_[4964]_ ;
  assign \new_[4968]_  = \new_[141]_  | \new_[142]_ ;
  assign \new_[4971]_  = \new_[139]_  | \new_[140]_ ;
  assign \new_[4972]_  = \new_[4971]_  | \new_[4968]_ ;
  assign \new_[4973]_  = \new_[4972]_  | \new_[4965]_ ;
  assign \new_[4974]_  = \new_[4973]_  | \new_[4960]_ ;
  assign \new_[4975]_  = \new_[4974]_  | \new_[4947]_ ;
  assign \new_[4979]_  = \new_[136]_  | \new_[137]_ ;
  assign \new_[4980]_  = \new_[138]_  | \new_[4979]_ ;
  assign \new_[4983]_  = \new_[134]_  | \new_[135]_ ;
  assign \new_[4986]_  = \new_[132]_  | \new_[133]_ ;
  assign \new_[4987]_  = \new_[4986]_  | \new_[4983]_ ;
  assign \new_[4988]_  = \new_[4987]_  | \new_[4980]_ ;
  assign \new_[4992]_  = \new_[129]_  | \new_[130]_ ;
  assign \new_[4993]_  = \new_[131]_  | \new_[4992]_ ;
  assign \new_[4996]_  = \new_[127]_  | \new_[128]_ ;
  assign \new_[4999]_  = \new_[125]_  | \new_[126]_ ;
  assign \new_[5000]_  = \new_[4999]_  | \new_[4996]_ ;
  assign \new_[5001]_  = \new_[5000]_  | \new_[4993]_ ;
  assign \new_[5002]_  = \new_[5001]_  | \new_[4988]_ ;
  assign \new_[5006]_  = \new_[122]_  | \new_[123]_ ;
  assign \new_[5007]_  = \new_[124]_  | \new_[5006]_ ;
  assign \new_[5010]_  = \new_[120]_  | \new_[121]_ ;
  assign \new_[5013]_  = \new_[118]_  | \new_[119]_ ;
  assign \new_[5014]_  = \new_[5013]_  | \new_[5010]_ ;
  assign \new_[5015]_  = \new_[5014]_  | \new_[5007]_ ;
  assign \new_[5019]_  = \new_[115]_  | \new_[116]_ ;
  assign \new_[5020]_  = \new_[117]_  | \new_[5019]_ ;
  assign \new_[5023]_  = \new_[113]_  | \new_[114]_ ;
  assign \new_[5026]_  = \new_[111]_  | \new_[112]_ ;
  assign \new_[5027]_  = \new_[5026]_  | \new_[5023]_ ;
  assign \new_[5028]_  = \new_[5027]_  | \new_[5020]_ ;
  assign \new_[5029]_  = \new_[5028]_  | \new_[5015]_ ;
  assign \new_[5030]_  = \new_[5029]_  | \new_[5002]_ ;
  assign \new_[5031]_  = \new_[5030]_  | \new_[4975]_ ;
  assign \new_[5032]_  = \new_[5031]_  | \new_[4922]_ ;
  assign \new_[5036]_  = \new_[108]_  | \new_[109]_ ;
  assign \new_[5037]_  = \new_[110]_  | \new_[5036]_ ;
  assign \new_[5041]_  = \new_[105]_  | \new_[106]_ ;
  assign \new_[5042]_  = \new_[107]_  | \new_[5041]_ ;
  assign \new_[5043]_  = \new_[5042]_  | \new_[5037]_ ;
  assign \new_[5047]_  = \new_[102]_  | \new_[103]_ ;
  assign \new_[5048]_  = \new_[104]_  | \new_[5047]_ ;
  assign \new_[5051]_  = \new_[100]_  | \new_[101]_ ;
  assign \new_[5054]_  = \new_[98]_  | \new_[99]_ ;
  assign \new_[5055]_  = \new_[5054]_  | \new_[5051]_ ;
  assign \new_[5056]_  = \new_[5055]_  | \new_[5048]_ ;
  assign \new_[5057]_  = \new_[5056]_  | \new_[5043]_ ;
  assign \new_[5061]_  = \new_[95]_  | \new_[96]_ ;
  assign \new_[5062]_  = \new_[97]_  | \new_[5061]_ ;
  assign \new_[5065]_  = \new_[93]_  | \new_[94]_ ;
  assign \new_[5068]_  = \new_[91]_  | \new_[92]_ ;
  assign \new_[5069]_  = \new_[5068]_  | \new_[5065]_ ;
  assign \new_[5070]_  = \new_[5069]_  | \new_[5062]_ ;
  assign \new_[5074]_  = \new_[88]_  | \new_[89]_ ;
  assign \new_[5075]_  = \new_[90]_  | \new_[5074]_ ;
  assign \new_[5078]_  = \new_[86]_  | \new_[87]_ ;
  assign \new_[5081]_  = \new_[84]_  | \new_[85]_ ;
  assign \new_[5082]_  = \new_[5081]_  | \new_[5078]_ ;
  assign \new_[5083]_  = \new_[5082]_  | \new_[5075]_ ;
  assign \new_[5084]_  = \new_[5083]_  | \new_[5070]_ ;
  assign \new_[5085]_  = \new_[5084]_  | \new_[5057]_ ;
  assign \new_[5089]_  = \new_[81]_  | \new_[82]_ ;
  assign \new_[5090]_  = \new_[83]_  | \new_[5089]_ ;
  assign \new_[5093]_  = \new_[79]_  | \new_[80]_ ;
  assign \new_[5096]_  = \new_[77]_  | \new_[78]_ ;
  assign \new_[5097]_  = \new_[5096]_  | \new_[5093]_ ;
  assign \new_[5098]_  = \new_[5097]_  | \new_[5090]_ ;
  assign \new_[5102]_  = \new_[74]_  | \new_[75]_ ;
  assign \new_[5103]_  = \new_[76]_  | \new_[5102]_ ;
  assign \new_[5106]_  = \new_[72]_  | \new_[73]_ ;
  assign \new_[5109]_  = \new_[70]_  | \new_[71]_ ;
  assign \new_[5110]_  = \new_[5109]_  | \new_[5106]_ ;
  assign \new_[5111]_  = \new_[5110]_  | \new_[5103]_ ;
  assign \new_[5112]_  = \new_[5111]_  | \new_[5098]_ ;
  assign \new_[5116]_  = \new_[67]_  | \new_[68]_ ;
  assign \new_[5117]_  = \new_[69]_  | \new_[5116]_ ;
  assign \new_[5120]_  = \new_[65]_  | \new_[66]_ ;
  assign \new_[5123]_  = \new_[63]_  | \new_[64]_ ;
  assign \new_[5124]_  = \new_[5123]_  | \new_[5120]_ ;
  assign \new_[5125]_  = \new_[5124]_  | \new_[5117]_ ;
  assign \new_[5129]_  = \new_[60]_  | \new_[61]_ ;
  assign \new_[5130]_  = \new_[62]_  | \new_[5129]_ ;
  assign \new_[5133]_  = \new_[58]_  | \new_[59]_ ;
  assign \new_[5136]_  = \new_[56]_  | \new_[57]_ ;
  assign \new_[5137]_  = \new_[5136]_  | \new_[5133]_ ;
  assign \new_[5138]_  = \new_[5137]_  | \new_[5130]_ ;
  assign \new_[5139]_  = \new_[5138]_  | \new_[5125]_ ;
  assign \new_[5140]_  = \new_[5139]_  | \new_[5112]_ ;
  assign \new_[5141]_  = \new_[5140]_  | \new_[5085]_ ;
  assign \new_[5145]_  = \new_[53]_  | \new_[54]_ ;
  assign \new_[5146]_  = \new_[55]_  | \new_[5145]_ ;
  assign \new_[5150]_  = \new_[50]_  | \new_[51]_ ;
  assign \new_[5151]_  = \new_[52]_  | \new_[5150]_ ;
  assign \new_[5152]_  = \new_[5151]_  | \new_[5146]_ ;
  assign \new_[5156]_  = \new_[47]_  | \new_[48]_ ;
  assign \new_[5157]_  = \new_[49]_  | \new_[5156]_ ;
  assign \new_[5160]_  = \new_[45]_  | \new_[46]_ ;
  assign \new_[5163]_  = \new_[43]_  | \new_[44]_ ;
  assign \new_[5164]_  = \new_[5163]_  | \new_[5160]_ ;
  assign \new_[5165]_  = \new_[5164]_  | \new_[5157]_ ;
  assign \new_[5166]_  = \new_[5165]_  | \new_[5152]_ ;
  assign \new_[5170]_  = \new_[40]_  | \new_[41]_ ;
  assign \new_[5171]_  = \new_[42]_  | \new_[5170]_ ;
  assign \new_[5174]_  = \new_[38]_  | \new_[39]_ ;
  assign \new_[5177]_  = \new_[36]_  | \new_[37]_ ;
  assign \new_[5178]_  = \new_[5177]_  | \new_[5174]_ ;
  assign \new_[5179]_  = \new_[5178]_  | \new_[5171]_ ;
  assign \new_[5183]_  = \new_[33]_  | \new_[34]_ ;
  assign \new_[5184]_  = \new_[35]_  | \new_[5183]_ ;
  assign \new_[5187]_  = \new_[31]_  | \new_[32]_ ;
  assign \new_[5190]_  = \new_[29]_  | \new_[30]_ ;
  assign \new_[5191]_  = \new_[5190]_  | \new_[5187]_ ;
  assign \new_[5192]_  = \new_[5191]_  | \new_[5184]_ ;
  assign \new_[5193]_  = \new_[5192]_  | \new_[5179]_ ;
  assign \new_[5194]_  = \new_[5193]_  | \new_[5166]_ ;
  assign \new_[5198]_  = \new_[26]_  | \new_[27]_ ;
  assign \new_[5199]_  = \new_[28]_  | \new_[5198]_ ;
  assign \new_[5202]_  = \new_[24]_  | \new_[25]_ ;
  assign \new_[5205]_  = \new_[22]_  | \new_[23]_ ;
  assign \new_[5206]_  = \new_[5205]_  | \new_[5202]_ ;
  assign \new_[5207]_  = \new_[5206]_  | \new_[5199]_ ;
  assign \new_[5211]_  = \new_[19]_  | \new_[20]_ ;
  assign \new_[5212]_  = \new_[21]_  | \new_[5211]_ ;
  assign \new_[5215]_  = \new_[17]_  | \new_[18]_ ;
  assign \new_[5218]_  = \new_[15]_  | \new_[16]_ ;
  assign \new_[5219]_  = \new_[5218]_  | \new_[5215]_ ;
  assign \new_[5220]_  = \new_[5219]_  | \new_[5212]_ ;
  assign \new_[5221]_  = \new_[5220]_  | \new_[5207]_ ;
  assign \new_[5225]_  = \new_[12]_  | \new_[13]_ ;
  assign \new_[5226]_  = \new_[14]_  | \new_[5225]_ ;
  assign \new_[5229]_  = \new_[10]_  | \new_[11]_ ;
  assign \new_[5232]_  = \new_[8]_  | \new_[9]_ ;
  assign \new_[5233]_  = \new_[5232]_  | \new_[5229]_ ;
  assign \new_[5234]_  = \new_[5233]_  | \new_[5226]_ ;
  assign \new_[5238]_  = \new_[5]_  | \new_[6]_ ;
  assign \new_[5239]_  = \new_[7]_  | \new_[5238]_ ;
  assign \new_[5242]_  = \new_[3]_  | \new_[4]_ ;
  assign \new_[5245]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[5246]_  = \new_[5245]_  | \new_[5242]_ ;
  assign \new_[5247]_  = \new_[5246]_  | \new_[5239]_ ;
  assign \new_[5248]_  = \new_[5247]_  | \new_[5234]_ ;
  assign \new_[5249]_  = \new_[5248]_  | \new_[5221]_ ;
  assign \new_[5250]_  = \new_[5249]_  | \new_[5194]_ ;
  assign \new_[5251]_  = \new_[5250]_  | \new_[5141]_ ;
  assign \new_[5252]_  = \new_[5251]_  | \new_[5032]_ ;
  assign \new_[5253]_  = \new_[5252]_  | \new_[4815]_ ;
  assign \new_[5254]_  = \new_[5253]_  | \new_[4378]_ ;
  assign \new_[5257]_  = A166 & A167;
  assign \new_[5260]_  = A201 & A199;
  assign \new_[5263]_  = A166 & A167;
  assign \new_[5266]_  = A201 & A200;
  assign \new_[5269]_  = ~A166 & ~A167;
  assign \new_[5272]_  = A201 & A199;
  assign \new_[5275]_  = ~A166 & ~A167;
  assign \new_[5278]_  = A201 & A200;
  assign \new_[5281]_  = ~A167 & ~A168;
  assign \new_[5284]_  = A201 & A199;
  assign \new_[5287]_  = ~A167 & ~A168;
  assign \new_[5290]_  = A201 & A200;
  assign \new_[5293]_  = ~A169 & ~A170;
  assign \new_[5297]_  = A201 & A199;
  assign \new_[5298]_  = ~A167 & \new_[5297]_ ;
  assign \new_[5301]_  = ~A169 & ~A170;
  assign \new_[5305]_  = A201 & A200;
  assign \new_[5306]_  = ~A167 & \new_[5305]_ ;
  assign \new_[5310]_  = A199 & A166;
  assign \new_[5311]_  = A167 & \new_[5310]_ ;
  assign \new_[5315]_  = ~A203 & A202;
  assign \new_[5316]_  = A200 & \new_[5315]_ ;
  assign \new_[5320]_  = ~A199 & A166;
  assign \new_[5321]_  = A167 & \new_[5320]_ ;
  assign \new_[5325]_  = A203 & ~A202;
  assign \new_[5326]_  = A200 & \new_[5325]_ ;
  assign \new_[5330]_  = A199 & A166;
  assign \new_[5331]_  = A167 & \new_[5330]_ ;
  assign \new_[5335]_  = A203 & ~A202;
  assign \new_[5336]_  = ~A200 & \new_[5335]_ ;
  assign \new_[5340]_  = ~A199 & A166;
  assign \new_[5341]_  = A167 & \new_[5340]_ ;
  assign \new_[5345]_  = ~A203 & A202;
  assign \new_[5346]_  = ~A200 & \new_[5345]_ ;
  assign \new_[5350]_  = A199 & ~A166;
  assign \new_[5351]_  = ~A167 & \new_[5350]_ ;
  assign \new_[5355]_  = ~A203 & A202;
  assign \new_[5356]_  = A200 & \new_[5355]_ ;
  assign \new_[5360]_  = ~A199 & ~A166;
  assign \new_[5361]_  = ~A167 & \new_[5360]_ ;
  assign \new_[5365]_  = A203 & ~A202;
  assign \new_[5366]_  = A200 & \new_[5365]_ ;
  assign \new_[5370]_  = A199 & ~A166;
  assign \new_[5371]_  = ~A167 & \new_[5370]_ ;
  assign \new_[5375]_  = A203 & ~A202;
  assign \new_[5376]_  = ~A200 & \new_[5375]_ ;
  assign \new_[5380]_  = ~A199 & ~A166;
  assign \new_[5381]_  = ~A167 & \new_[5380]_ ;
  assign \new_[5385]_  = ~A203 & A202;
  assign \new_[5386]_  = ~A200 & \new_[5385]_ ;
  assign \new_[5390]_  = A199 & ~A167;
  assign \new_[5391]_  = ~A168 & \new_[5390]_ ;
  assign \new_[5395]_  = ~A203 & A202;
  assign \new_[5396]_  = A200 & \new_[5395]_ ;
  assign \new_[5400]_  = ~A199 & ~A167;
  assign \new_[5401]_  = ~A168 & \new_[5400]_ ;
  assign \new_[5405]_  = A203 & ~A202;
  assign \new_[5406]_  = A200 & \new_[5405]_ ;
  assign \new_[5410]_  = A199 & ~A167;
  assign \new_[5411]_  = ~A168 & \new_[5410]_ ;
  assign \new_[5415]_  = A203 & ~A202;
  assign \new_[5416]_  = ~A200 & \new_[5415]_ ;
  assign \new_[5420]_  = ~A199 & ~A167;
  assign \new_[5421]_  = ~A168 & \new_[5420]_ ;
  assign \new_[5425]_  = ~A203 & A202;
  assign \new_[5426]_  = ~A200 & \new_[5425]_ ;
  assign \new_[5430]_  = ~A167 & ~A169;
  assign \new_[5431]_  = ~A170 & \new_[5430]_ ;
  assign \new_[5434]_  = A200 & A199;
  assign \new_[5437]_  = ~A203 & A202;
  assign \new_[5438]_  = \new_[5437]_  & \new_[5434]_ ;
  assign \new_[5442]_  = ~A167 & ~A169;
  assign \new_[5443]_  = ~A170 & \new_[5442]_ ;
  assign \new_[5446]_  = A200 & ~A199;
  assign \new_[5449]_  = A203 & ~A202;
  assign \new_[5450]_  = \new_[5449]_  & \new_[5446]_ ;
  assign \new_[5454]_  = ~A167 & ~A169;
  assign \new_[5455]_  = ~A170 & \new_[5454]_ ;
  assign \new_[5458]_  = ~A200 & A199;
  assign \new_[5461]_  = A203 & ~A202;
  assign \new_[5462]_  = \new_[5461]_  & \new_[5458]_ ;
  assign \new_[5466]_  = ~A167 & ~A169;
  assign \new_[5467]_  = ~A170 & \new_[5466]_ ;
  assign \new_[5470]_  = ~A200 & ~A199;
  assign \new_[5473]_  = ~A203 & A202;
  assign \new_[5474]_  = \new_[5473]_  & \new_[5470]_ ;
  assign \new_[5477]_  = ~A166 & A167;
  assign \new_[5480]_  = ~A200 & ~A199;
  assign \new_[5481]_  = \new_[5480]_  & \new_[5477]_ ;
  assign \new_[5484]_  = A232 & ~A202;
  assign \new_[5488]_  = A300 & A299;
  assign \new_[5489]_  = A234 & \new_[5488]_ ;
  assign \new_[5490]_  = \new_[5489]_  & \new_[5484]_ ;
  assign \new_[5493]_  = ~A166 & A167;
  assign \new_[5496]_  = ~A200 & ~A199;
  assign \new_[5497]_  = \new_[5496]_  & \new_[5493]_ ;
  assign \new_[5500]_  = A232 & ~A202;
  assign \new_[5504]_  = A300 & A298;
  assign \new_[5505]_  = A234 & \new_[5504]_ ;
  assign \new_[5506]_  = \new_[5505]_  & \new_[5500]_ ;
  assign \new_[5509]_  = ~A166 & A167;
  assign \new_[5512]_  = ~A200 & ~A199;
  assign \new_[5513]_  = \new_[5512]_  & \new_[5509]_ ;
  assign \new_[5516]_  = A232 & ~A202;
  assign \new_[5520]_  = A267 & A265;
  assign \new_[5521]_  = A234 & \new_[5520]_ ;
  assign \new_[5522]_  = \new_[5521]_  & \new_[5516]_ ;
  assign \new_[5525]_  = ~A166 & A167;
  assign \new_[5528]_  = ~A200 & ~A199;
  assign \new_[5529]_  = \new_[5528]_  & \new_[5525]_ ;
  assign \new_[5532]_  = A232 & ~A202;
  assign \new_[5536]_  = A267 & A266;
  assign \new_[5537]_  = A234 & \new_[5536]_ ;
  assign \new_[5538]_  = \new_[5537]_  & \new_[5532]_ ;
  assign \new_[5541]_  = ~A166 & A167;
  assign \new_[5544]_  = ~A200 & ~A199;
  assign \new_[5545]_  = \new_[5544]_  & \new_[5541]_ ;
  assign \new_[5548]_  = A233 & ~A202;
  assign \new_[5552]_  = A300 & A299;
  assign \new_[5553]_  = A234 & \new_[5552]_ ;
  assign \new_[5554]_  = \new_[5553]_  & \new_[5548]_ ;
  assign \new_[5557]_  = ~A166 & A167;
  assign \new_[5560]_  = ~A200 & ~A199;
  assign \new_[5561]_  = \new_[5560]_  & \new_[5557]_ ;
  assign \new_[5564]_  = A233 & ~A202;
  assign \new_[5568]_  = A300 & A298;
  assign \new_[5569]_  = A234 & \new_[5568]_ ;
  assign \new_[5570]_  = \new_[5569]_  & \new_[5564]_ ;
  assign \new_[5573]_  = ~A166 & A167;
  assign \new_[5576]_  = ~A200 & ~A199;
  assign \new_[5577]_  = \new_[5576]_  & \new_[5573]_ ;
  assign \new_[5580]_  = A233 & ~A202;
  assign \new_[5584]_  = A267 & A265;
  assign \new_[5585]_  = A234 & \new_[5584]_ ;
  assign \new_[5586]_  = \new_[5585]_  & \new_[5580]_ ;
  assign \new_[5589]_  = ~A166 & A167;
  assign \new_[5592]_  = ~A200 & ~A199;
  assign \new_[5593]_  = \new_[5592]_  & \new_[5589]_ ;
  assign \new_[5596]_  = A233 & ~A202;
  assign \new_[5600]_  = A267 & A266;
  assign \new_[5601]_  = A234 & \new_[5600]_ ;
  assign \new_[5602]_  = \new_[5601]_  & \new_[5596]_ ;
  assign \new_[5605]_  = ~A166 & A167;
  assign \new_[5608]_  = ~A200 & ~A199;
  assign \new_[5609]_  = \new_[5608]_  & \new_[5605]_ ;
  assign \new_[5612]_  = A232 & A203;
  assign \new_[5616]_  = A300 & A299;
  assign \new_[5617]_  = A234 & \new_[5616]_ ;
  assign \new_[5618]_  = \new_[5617]_  & \new_[5612]_ ;
  assign \new_[5621]_  = ~A166 & A167;
  assign \new_[5624]_  = ~A200 & ~A199;
  assign \new_[5625]_  = \new_[5624]_  & \new_[5621]_ ;
  assign \new_[5628]_  = A232 & A203;
  assign \new_[5632]_  = A300 & A298;
  assign \new_[5633]_  = A234 & \new_[5632]_ ;
  assign \new_[5634]_  = \new_[5633]_  & \new_[5628]_ ;
  assign \new_[5637]_  = ~A166 & A167;
  assign \new_[5640]_  = ~A200 & ~A199;
  assign \new_[5641]_  = \new_[5640]_  & \new_[5637]_ ;
  assign \new_[5644]_  = A232 & A203;
  assign \new_[5648]_  = A267 & A265;
  assign \new_[5649]_  = A234 & \new_[5648]_ ;
  assign \new_[5650]_  = \new_[5649]_  & \new_[5644]_ ;
  assign \new_[5653]_  = ~A166 & A167;
  assign \new_[5656]_  = ~A200 & ~A199;
  assign \new_[5657]_  = \new_[5656]_  & \new_[5653]_ ;
  assign \new_[5660]_  = A232 & A203;
  assign \new_[5664]_  = A267 & A266;
  assign \new_[5665]_  = A234 & \new_[5664]_ ;
  assign \new_[5666]_  = \new_[5665]_  & \new_[5660]_ ;
  assign \new_[5669]_  = ~A166 & A167;
  assign \new_[5672]_  = ~A200 & ~A199;
  assign \new_[5673]_  = \new_[5672]_  & \new_[5669]_ ;
  assign \new_[5676]_  = A233 & A203;
  assign \new_[5680]_  = A300 & A299;
  assign \new_[5681]_  = A234 & \new_[5680]_ ;
  assign \new_[5682]_  = \new_[5681]_  & \new_[5676]_ ;
  assign \new_[5685]_  = ~A166 & A167;
  assign \new_[5688]_  = ~A200 & ~A199;
  assign \new_[5689]_  = \new_[5688]_  & \new_[5685]_ ;
  assign \new_[5692]_  = A233 & A203;
  assign \new_[5696]_  = A300 & A298;
  assign \new_[5697]_  = A234 & \new_[5696]_ ;
  assign \new_[5698]_  = \new_[5697]_  & \new_[5692]_ ;
  assign \new_[5701]_  = ~A166 & A167;
  assign \new_[5704]_  = ~A200 & ~A199;
  assign \new_[5705]_  = \new_[5704]_  & \new_[5701]_ ;
  assign \new_[5708]_  = A233 & A203;
  assign \new_[5712]_  = A267 & A265;
  assign \new_[5713]_  = A234 & \new_[5712]_ ;
  assign \new_[5714]_  = \new_[5713]_  & \new_[5708]_ ;
  assign \new_[5717]_  = ~A166 & A167;
  assign \new_[5720]_  = ~A200 & ~A199;
  assign \new_[5721]_  = \new_[5720]_  & \new_[5717]_ ;
  assign \new_[5724]_  = A233 & A203;
  assign \new_[5728]_  = A267 & A266;
  assign \new_[5729]_  = A234 & \new_[5728]_ ;
  assign \new_[5730]_  = \new_[5729]_  & \new_[5724]_ ;
  assign \new_[5733]_  = ~A166 & A167;
  assign \new_[5737]_  = ~A201 & A200;
  assign \new_[5738]_  = A199 & \new_[5737]_ ;
  assign \new_[5739]_  = \new_[5738]_  & \new_[5733]_ ;
  assign \new_[5742]_  = A232 & ~A202;
  assign \new_[5746]_  = A300 & A299;
  assign \new_[5747]_  = A234 & \new_[5746]_ ;
  assign \new_[5748]_  = \new_[5747]_  & \new_[5742]_ ;
  assign \new_[5751]_  = ~A166 & A167;
  assign \new_[5755]_  = ~A201 & A200;
  assign \new_[5756]_  = A199 & \new_[5755]_ ;
  assign \new_[5757]_  = \new_[5756]_  & \new_[5751]_ ;
  assign \new_[5760]_  = A232 & ~A202;
  assign \new_[5764]_  = A300 & A298;
  assign \new_[5765]_  = A234 & \new_[5764]_ ;
  assign \new_[5766]_  = \new_[5765]_  & \new_[5760]_ ;
  assign \new_[5769]_  = ~A166 & A167;
  assign \new_[5773]_  = ~A201 & A200;
  assign \new_[5774]_  = A199 & \new_[5773]_ ;
  assign \new_[5775]_  = \new_[5774]_  & \new_[5769]_ ;
  assign \new_[5778]_  = A232 & ~A202;
  assign \new_[5782]_  = A267 & A265;
  assign \new_[5783]_  = A234 & \new_[5782]_ ;
  assign \new_[5784]_  = \new_[5783]_  & \new_[5778]_ ;
  assign \new_[5787]_  = ~A166 & A167;
  assign \new_[5791]_  = ~A201 & A200;
  assign \new_[5792]_  = A199 & \new_[5791]_ ;
  assign \new_[5793]_  = \new_[5792]_  & \new_[5787]_ ;
  assign \new_[5796]_  = A232 & ~A202;
  assign \new_[5800]_  = A267 & A266;
  assign \new_[5801]_  = A234 & \new_[5800]_ ;
  assign \new_[5802]_  = \new_[5801]_  & \new_[5796]_ ;
  assign \new_[5805]_  = ~A166 & A167;
  assign \new_[5809]_  = ~A201 & A200;
  assign \new_[5810]_  = A199 & \new_[5809]_ ;
  assign \new_[5811]_  = \new_[5810]_  & \new_[5805]_ ;
  assign \new_[5814]_  = A233 & ~A202;
  assign \new_[5818]_  = A300 & A299;
  assign \new_[5819]_  = A234 & \new_[5818]_ ;
  assign \new_[5820]_  = \new_[5819]_  & \new_[5814]_ ;
  assign \new_[5823]_  = ~A166 & A167;
  assign \new_[5827]_  = ~A201 & A200;
  assign \new_[5828]_  = A199 & \new_[5827]_ ;
  assign \new_[5829]_  = \new_[5828]_  & \new_[5823]_ ;
  assign \new_[5832]_  = A233 & ~A202;
  assign \new_[5836]_  = A300 & A298;
  assign \new_[5837]_  = A234 & \new_[5836]_ ;
  assign \new_[5838]_  = \new_[5837]_  & \new_[5832]_ ;
  assign \new_[5841]_  = ~A166 & A167;
  assign \new_[5845]_  = ~A201 & A200;
  assign \new_[5846]_  = A199 & \new_[5845]_ ;
  assign \new_[5847]_  = \new_[5846]_  & \new_[5841]_ ;
  assign \new_[5850]_  = A233 & ~A202;
  assign \new_[5854]_  = A267 & A265;
  assign \new_[5855]_  = A234 & \new_[5854]_ ;
  assign \new_[5856]_  = \new_[5855]_  & \new_[5850]_ ;
  assign \new_[5859]_  = ~A166 & A167;
  assign \new_[5863]_  = ~A201 & A200;
  assign \new_[5864]_  = A199 & \new_[5863]_ ;
  assign \new_[5865]_  = \new_[5864]_  & \new_[5859]_ ;
  assign \new_[5868]_  = A233 & ~A202;
  assign \new_[5872]_  = A267 & A266;
  assign \new_[5873]_  = A234 & \new_[5872]_ ;
  assign \new_[5874]_  = \new_[5873]_  & \new_[5868]_ ;
  assign \new_[5877]_  = ~A166 & A167;
  assign \new_[5881]_  = ~A201 & A200;
  assign \new_[5882]_  = A199 & \new_[5881]_ ;
  assign \new_[5883]_  = \new_[5882]_  & \new_[5877]_ ;
  assign \new_[5886]_  = A232 & A203;
  assign \new_[5890]_  = A300 & A299;
  assign \new_[5891]_  = A234 & \new_[5890]_ ;
  assign \new_[5892]_  = \new_[5891]_  & \new_[5886]_ ;
  assign \new_[5895]_  = ~A166 & A167;
  assign \new_[5899]_  = ~A201 & A200;
  assign \new_[5900]_  = A199 & \new_[5899]_ ;
  assign \new_[5901]_  = \new_[5900]_  & \new_[5895]_ ;
  assign \new_[5904]_  = A232 & A203;
  assign \new_[5908]_  = A300 & A298;
  assign \new_[5909]_  = A234 & \new_[5908]_ ;
  assign \new_[5910]_  = \new_[5909]_  & \new_[5904]_ ;
  assign \new_[5913]_  = ~A166 & A167;
  assign \new_[5917]_  = ~A201 & A200;
  assign \new_[5918]_  = A199 & \new_[5917]_ ;
  assign \new_[5919]_  = \new_[5918]_  & \new_[5913]_ ;
  assign \new_[5922]_  = A232 & A203;
  assign \new_[5926]_  = A267 & A265;
  assign \new_[5927]_  = A234 & \new_[5926]_ ;
  assign \new_[5928]_  = \new_[5927]_  & \new_[5922]_ ;
  assign \new_[5931]_  = ~A166 & A167;
  assign \new_[5935]_  = ~A201 & A200;
  assign \new_[5936]_  = A199 & \new_[5935]_ ;
  assign \new_[5937]_  = \new_[5936]_  & \new_[5931]_ ;
  assign \new_[5940]_  = A232 & A203;
  assign \new_[5944]_  = A267 & A266;
  assign \new_[5945]_  = A234 & \new_[5944]_ ;
  assign \new_[5946]_  = \new_[5945]_  & \new_[5940]_ ;
  assign \new_[5949]_  = ~A166 & A167;
  assign \new_[5953]_  = ~A201 & A200;
  assign \new_[5954]_  = A199 & \new_[5953]_ ;
  assign \new_[5955]_  = \new_[5954]_  & \new_[5949]_ ;
  assign \new_[5958]_  = A233 & A203;
  assign \new_[5962]_  = A300 & A299;
  assign \new_[5963]_  = A234 & \new_[5962]_ ;
  assign \new_[5964]_  = \new_[5963]_  & \new_[5958]_ ;
  assign \new_[5967]_  = ~A166 & A167;
  assign \new_[5971]_  = ~A201 & A200;
  assign \new_[5972]_  = A199 & \new_[5971]_ ;
  assign \new_[5973]_  = \new_[5972]_  & \new_[5967]_ ;
  assign \new_[5976]_  = A233 & A203;
  assign \new_[5980]_  = A300 & A298;
  assign \new_[5981]_  = A234 & \new_[5980]_ ;
  assign \new_[5982]_  = \new_[5981]_  & \new_[5976]_ ;
  assign \new_[5985]_  = ~A166 & A167;
  assign \new_[5989]_  = ~A201 & A200;
  assign \new_[5990]_  = A199 & \new_[5989]_ ;
  assign \new_[5991]_  = \new_[5990]_  & \new_[5985]_ ;
  assign \new_[5994]_  = A233 & A203;
  assign \new_[5998]_  = A267 & A265;
  assign \new_[5999]_  = A234 & \new_[5998]_ ;
  assign \new_[6000]_  = \new_[5999]_  & \new_[5994]_ ;
  assign \new_[6003]_  = ~A166 & A167;
  assign \new_[6007]_  = ~A201 & A200;
  assign \new_[6008]_  = A199 & \new_[6007]_ ;
  assign \new_[6009]_  = \new_[6008]_  & \new_[6003]_ ;
  assign \new_[6012]_  = A233 & A203;
  assign \new_[6016]_  = A267 & A266;
  assign \new_[6017]_  = A234 & \new_[6016]_ ;
  assign \new_[6018]_  = \new_[6017]_  & \new_[6012]_ ;
  assign \new_[6021]_  = ~A166 & A167;
  assign \new_[6025]_  = ~A201 & A200;
  assign \new_[6026]_  = ~A199 & \new_[6025]_ ;
  assign \new_[6027]_  = \new_[6026]_  & \new_[6021]_ ;
  assign \new_[6030]_  = A232 & A202;
  assign \new_[6034]_  = A300 & A299;
  assign \new_[6035]_  = A234 & \new_[6034]_ ;
  assign \new_[6036]_  = \new_[6035]_  & \new_[6030]_ ;
  assign \new_[6039]_  = ~A166 & A167;
  assign \new_[6043]_  = ~A201 & A200;
  assign \new_[6044]_  = ~A199 & \new_[6043]_ ;
  assign \new_[6045]_  = \new_[6044]_  & \new_[6039]_ ;
  assign \new_[6048]_  = A232 & A202;
  assign \new_[6052]_  = A300 & A298;
  assign \new_[6053]_  = A234 & \new_[6052]_ ;
  assign \new_[6054]_  = \new_[6053]_  & \new_[6048]_ ;
  assign \new_[6057]_  = ~A166 & A167;
  assign \new_[6061]_  = ~A201 & A200;
  assign \new_[6062]_  = ~A199 & \new_[6061]_ ;
  assign \new_[6063]_  = \new_[6062]_  & \new_[6057]_ ;
  assign \new_[6066]_  = A232 & A202;
  assign \new_[6070]_  = A267 & A265;
  assign \new_[6071]_  = A234 & \new_[6070]_ ;
  assign \new_[6072]_  = \new_[6071]_  & \new_[6066]_ ;
  assign \new_[6075]_  = ~A166 & A167;
  assign \new_[6079]_  = ~A201 & A200;
  assign \new_[6080]_  = ~A199 & \new_[6079]_ ;
  assign \new_[6081]_  = \new_[6080]_  & \new_[6075]_ ;
  assign \new_[6084]_  = A232 & A202;
  assign \new_[6088]_  = A267 & A266;
  assign \new_[6089]_  = A234 & \new_[6088]_ ;
  assign \new_[6090]_  = \new_[6089]_  & \new_[6084]_ ;
  assign \new_[6093]_  = ~A166 & A167;
  assign \new_[6097]_  = ~A201 & A200;
  assign \new_[6098]_  = ~A199 & \new_[6097]_ ;
  assign \new_[6099]_  = \new_[6098]_  & \new_[6093]_ ;
  assign \new_[6102]_  = A233 & A202;
  assign \new_[6106]_  = A300 & A299;
  assign \new_[6107]_  = A234 & \new_[6106]_ ;
  assign \new_[6108]_  = \new_[6107]_  & \new_[6102]_ ;
  assign \new_[6111]_  = ~A166 & A167;
  assign \new_[6115]_  = ~A201 & A200;
  assign \new_[6116]_  = ~A199 & \new_[6115]_ ;
  assign \new_[6117]_  = \new_[6116]_  & \new_[6111]_ ;
  assign \new_[6120]_  = A233 & A202;
  assign \new_[6124]_  = A300 & A298;
  assign \new_[6125]_  = A234 & \new_[6124]_ ;
  assign \new_[6126]_  = \new_[6125]_  & \new_[6120]_ ;
  assign \new_[6129]_  = ~A166 & A167;
  assign \new_[6133]_  = ~A201 & A200;
  assign \new_[6134]_  = ~A199 & \new_[6133]_ ;
  assign \new_[6135]_  = \new_[6134]_  & \new_[6129]_ ;
  assign \new_[6138]_  = A233 & A202;
  assign \new_[6142]_  = A267 & A265;
  assign \new_[6143]_  = A234 & \new_[6142]_ ;
  assign \new_[6144]_  = \new_[6143]_  & \new_[6138]_ ;
  assign \new_[6147]_  = ~A166 & A167;
  assign \new_[6151]_  = ~A201 & A200;
  assign \new_[6152]_  = ~A199 & \new_[6151]_ ;
  assign \new_[6153]_  = \new_[6152]_  & \new_[6147]_ ;
  assign \new_[6156]_  = A233 & A202;
  assign \new_[6160]_  = A267 & A266;
  assign \new_[6161]_  = A234 & \new_[6160]_ ;
  assign \new_[6162]_  = \new_[6161]_  & \new_[6156]_ ;
  assign \new_[6165]_  = ~A166 & A167;
  assign \new_[6169]_  = ~A201 & A200;
  assign \new_[6170]_  = ~A199 & \new_[6169]_ ;
  assign \new_[6171]_  = \new_[6170]_  & \new_[6165]_ ;
  assign \new_[6174]_  = A232 & ~A203;
  assign \new_[6178]_  = A300 & A299;
  assign \new_[6179]_  = A234 & \new_[6178]_ ;
  assign \new_[6180]_  = \new_[6179]_  & \new_[6174]_ ;
  assign \new_[6183]_  = ~A166 & A167;
  assign \new_[6187]_  = ~A201 & A200;
  assign \new_[6188]_  = ~A199 & \new_[6187]_ ;
  assign \new_[6189]_  = \new_[6188]_  & \new_[6183]_ ;
  assign \new_[6192]_  = A232 & ~A203;
  assign \new_[6196]_  = A300 & A298;
  assign \new_[6197]_  = A234 & \new_[6196]_ ;
  assign \new_[6198]_  = \new_[6197]_  & \new_[6192]_ ;
  assign \new_[6201]_  = ~A166 & A167;
  assign \new_[6205]_  = ~A201 & A200;
  assign \new_[6206]_  = ~A199 & \new_[6205]_ ;
  assign \new_[6207]_  = \new_[6206]_  & \new_[6201]_ ;
  assign \new_[6210]_  = A232 & ~A203;
  assign \new_[6214]_  = A267 & A265;
  assign \new_[6215]_  = A234 & \new_[6214]_ ;
  assign \new_[6216]_  = \new_[6215]_  & \new_[6210]_ ;
  assign \new_[6219]_  = ~A166 & A167;
  assign \new_[6223]_  = ~A201 & A200;
  assign \new_[6224]_  = ~A199 & \new_[6223]_ ;
  assign \new_[6225]_  = \new_[6224]_  & \new_[6219]_ ;
  assign \new_[6228]_  = A232 & ~A203;
  assign \new_[6232]_  = A267 & A266;
  assign \new_[6233]_  = A234 & \new_[6232]_ ;
  assign \new_[6234]_  = \new_[6233]_  & \new_[6228]_ ;
  assign \new_[6237]_  = ~A166 & A167;
  assign \new_[6241]_  = ~A201 & A200;
  assign \new_[6242]_  = ~A199 & \new_[6241]_ ;
  assign \new_[6243]_  = \new_[6242]_  & \new_[6237]_ ;
  assign \new_[6246]_  = A233 & ~A203;
  assign \new_[6250]_  = A300 & A299;
  assign \new_[6251]_  = A234 & \new_[6250]_ ;
  assign \new_[6252]_  = \new_[6251]_  & \new_[6246]_ ;
  assign \new_[6255]_  = ~A166 & A167;
  assign \new_[6259]_  = ~A201 & A200;
  assign \new_[6260]_  = ~A199 & \new_[6259]_ ;
  assign \new_[6261]_  = \new_[6260]_  & \new_[6255]_ ;
  assign \new_[6264]_  = A233 & ~A203;
  assign \new_[6268]_  = A300 & A298;
  assign \new_[6269]_  = A234 & \new_[6268]_ ;
  assign \new_[6270]_  = \new_[6269]_  & \new_[6264]_ ;
  assign \new_[6273]_  = ~A166 & A167;
  assign \new_[6277]_  = ~A201 & A200;
  assign \new_[6278]_  = ~A199 & \new_[6277]_ ;
  assign \new_[6279]_  = \new_[6278]_  & \new_[6273]_ ;
  assign \new_[6282]_  = A233 & ~A203;
  assign \new_[6286]_  = A267 & A265;
  assign \new_[6287]_  = A234 & \new_[6286]_ ;
  assign \new_[6288]_  = \new_[6287]_  & \new_[6282]_ ;
  assign \new_[6291]_  = ~A166 & A167;
  assign \new_[6295]_  = ~A201 & A200;
  assign \new_[6296]_  = ~A199 & \new_[6295]_ ;
  assign \new_[6297]_  = \new_[6296]_  & \new_[6291]_ ;
  assign \new_[6300]_  = A233 & ~A203;
  assign \new_[6304]_  = A267 & A266;
  assign \new_[6305]_  = A234 & \new_[6304]_ ;
  assign \new_[6306]_  = \new_[6305]_  & \new_[6300]_ ;
  assign \new_[6309]_  = ~A166 & A167;
  assign \new_[6313]_  = ~A201 & ~A200;
  assign \new_[6314]_  = A199 & \new_[6313]_ ;
  assign \new_[6315]_  = \new_[6314]_  & \new_[6309]_ ;
  assign \new_[6318]_  = A232 & A202;
  assign \new_[6322]_  = A300 & A299;
  assign \new_[6323]_  = A234 & \new_[6322]_ ;
  assign \new_[6324]_  = \new_[6323]_  & \new_[6318]_ ;
  assign \new_[6327]_  = ~A166 & A167;
  assign \new_[6331]_  = ~A201 & ~A200;
  assign \new_[6332]_  = A199 & \new_[6331]_ ;
  assign \new_[6333]_  = \new_[6332]_  & \new_[6327]_ ;
  assign \new_[6336]_  = A232 & A202;
  assign \new_[6340]_  = A300 & A298;
  assign \new_[6341]_  = A234 & \new_[6340]_ ;
  assign \new_[6342]_  = \new_[6341]_  & \new_[6336]_ ;
  assign \new_[6345]_  = ~A166 & A167;
  assign \new_[6349]_  = ~A201 & ~A200;
  assign \new_[6350]_  = A199 & \new_[6349]_ ;
  assign \new_[6351]_  = \new_[6350]_  & \new_[6345]_ ;
  assign \new_[6354]_  = A232 & A202;
  assign \new_[6358]_  = A267 & A265;
  assign \new_[6359]_  = A234 & \new_[6358]_ ;
  assign \new_[6360]_  = \new_[6359]_  & \new_[6354]_ ;
  assign \new_[6363]_  = ~A166 & A167;
  assign \new_[6367]_  = ~A201 & ~A200;
  assign \new_[6368]_  = A199 & \new_[6367]_ ;
  assign \new_[6369]_  = \new_[6368]_  & \new_[6363]_ ;
  assign \new_[6372]_  = A232 & A202;
  assign \new_[6376]_  = A267 & A266;
  assign \new_[6377]_  = A234 & \new_[6376]_ ;
  assign \new_[6378]_  = \new_[6377]_  & \new_[6372]_ ;
  assign \new_[6381]_  = ~A166 & A167;
  assign \new_[6385]_  = ~A201 & ~A200;
  assign \new_[6386]_  = A199 & \new_[6385]_ ;
  assign \new_[6387]_  = \new_[6386]_  & \new_[6381]_ ;
  assign \new_[6390]_  = A233 & A202;
  assign \new_[6394]_  = A300 & A299;
  assign \new_[6395]_  = A234 & \new_[6394]_ ;
  assign \new_[6396]_  = \new_[6395]_  & \new_[6390]_ ;
  assign \new_[6399]_  = ~A166 & A167;
  assign \new_[6403]_  = ~A201 & ~A200;
  assign \new_[6404]_  = A199 & \new_[6403]_ ;
  assign \new_[6405]_  = \new_[6404]_  & \new_[6399]_ ;
  assign \new_[6408]_  = A233 & A202;
  assign \new_[6412]_  = A300 & A298;
  assign \new_[6413]_  = A234 & \new_[6412]_ ;
  assign \new_[6414]_  = \new_[6413]_  & \new_[6408]_ ;
  assign \new_[6417]_  = ~A166 & A167;
  assign \new_[6421]_  = ~A201 & ~A200;
  assign \new_[6422]_  = A199 & \new_[6421]_ ;
  assign \new_[6423]_  = \new_[6422]_  & \new_[6417]_ ;
  assign \new_[6426]_  = A233 & A202;
  assign \new_[6430]_  = A267 & A265;
  assign \new_[6431]_  = A234 & \new_[6430]_ ;
  assign \new_[6432]_  = \new_[6431]_  & \new_[6426]_ ;
  assign \new_[6435]_  = ~A166 & A167;
  assign \new_[6439]_  = ~A201 & ~A200;
  assign \new_[6440]_  = A199 & \new_[6439]_ ;
  assign \new_[6441]_  = \new_[6440]_  & \new_[6435]_ ;
  assign \new_[6444]_  = A233 & A202;
  assign \new_[6448]_  = A267 & A266;
  assign \new_[6449]_  = A234 & \new_[6448]_ ;
  assign \new_[6450]_  = \new_[6449]_  & \new_[6444]_ ;
  assign \new_[6453]_  = ~A166 & A167;
  assign \new_[6457]_  = ~A201 & ~A200;
  assign \new_[6458]_  = A199 & \new_[6457]_ ;
  assign \new_[6459]_  = \new_[6458]_  & \new_[6453]_ ;
  assign \new_[6462]_  = A232 & ~A203;
  assign \new_[6466]_  = A300 & A299;
  assign \new_[6467]_  = A234 & \new_[6466]_ ;
  assign \new_[6468]_  = \new_[6467]_  & \new_[6462]_ ;
  assign \new_[6471]_  = ~A166 & A167;
  assign \new_[6475]_  = ~A201 & ~A200;
  assign \new_[6476]_  = A199 & \new_[6475]_ ;
  assign \new_[6477]_  = \new_[6476]_  & \new_[6471]_ ;
  assign \new_[6480]_  = A232 & ~A203;
  assign \new_[6484]_  = A300 & A298;
  assign \new_[6485]_  = A234 & \new_[6484]_ ;
  assign \new_[6486]_  = \new_[6485]_  & \new_[6480]_ ;
  assign \new_[6489]_  = ~A166 & A167;
  assign \new_[6493]_  = ~A201 & ~A200;
  assign \new_[6494]_  = A199 & \new_[6493]_ ;
  assign \new_[6495]_  = \new_[6494]_  & \new_[6489]_ ;
  assign \new_[6498]_  = A232 & ~A203;
  assign \new_[6502]_  = A267 & A265;
  assign \new_[6503]_  = A234 & \new_[6502]_ ;
  assign \new_[6504]_  = \new_[6503]_  & \new_[6498]_ ;
  assign \new_[6507]_  = ~A166 & A167;
  assign \new_[6511]_  = ~A201 & ~A200;
  assign \new_[6512]_  = A199 & \new_[6511]_ ;
  assign \new_[6513]_  = \new_[6512]_  & \new_[6507]_ ;
  assign \new_[6516]_  = A232 & ~A203;
  assign \new_[6520]_  = A267 & A266;
  assign \new_[6521]_  = A234 & \new_[6520]_ ;
  assign \new_[6522]_  = \new_[6521]_  & \new_[6516]_ ;
  assign \new_[6525]_  = ~A166 & A167;
  assign \new_[6529]_  = ~A201 & ~A200;
  assign \new_[6530]_  = A199 & \new_[6529]_ ;
  assign \new_[6531]_  = \new_[6530]_  & \new_[6525]_ ;
  assign \new_[6534]_  = A233 & ~A203;
  assign \new_[6538]_  = A300 & A299;
  assign \new_[6539]_  = A234 & \new_[6538]_ ;
  assign \new_[6540]_  = \new_[6539]_  & \new_[6534]_ ;
  assign \new_[6543]_  = ~A166 & A167;
  assign \new_[6547]_  = ~A201 & ~A200;
  assign \new_[6548]_  = A199 & \new_[6547]_ ;
  assign \new_[6549]_  = \new_[6548]_  & \new_[6543]_ ;
  assign \new_[6552]_  = A233 & ~A203;
  assign \new_[6556]_  = A300 & A298;
  assign \new_[6557]_  = A234 & \new_[6556]_ ;
  assign \new_[6558]_  = \new_[6557]_  & \new_[6552]_ ;
  assign \new_[6561]_  = ~A166 & A167;
  assign \new_[6565]_  = ~A201 & ~A200;
  assign \new_[6566]_  = A199 & \new_[6565]_ ;
  assign \new_[6567]_  = \new_[6566]_  & \new_[6561]_ ;
  assign \new_[6570]_  = A233 & ~A203;
  assign \new_[6574]_  = A267 & A265;
  assign \new_[6575]_  = A234 & \new_[6574]_ ;
  assign \new_[6576]_  = \new_[6575]_  & \new_[6570]_ ;
  assign \new_[6579]_  = ~A166 & A167;
  assign \new_[6583]_  = ~A201 & ~A200;
  assign \new_[6584]_  = A199 & \new_[6583]_ ;
  assign \new_[6585]_  = \new_[6584]_  & \new_[6579]_ ;
  assign \new_[6588]_  = A233 & ~A203;
  assign \new_[6592]_  = A267 & A266;
  assign \new_[6593]_  = A234 & \new_[6592]_ ;
  assign \new_[6594]_  = \new_[6593]_  & \new_[6588]_ ;
  assign \new_[6597]_  = ~A166 & A167;
  assign \new_[6601]_  = ~A202 & ~A200;
  assign \new_[6602]_  = ~A199 & \new_[6601]_ ;
  assign \new_[6603]_  = \new_[6602]_  & \new_[6597]_ ;
  assign \new_[6607]_  = A298 & A234;
  assign \new_[6608]_  = A232 & \new_[6607]_ ;
  assign \new_[6612]_  = ~A302 & A301;
  assign \new_[6613]_  = A299 & \new_[6612]_ ;
  assign \new_[6614]_  = \new_[6613]_  & \new_[6608]_ ;
  assign \new_[6617]_  = ~A166 & A167;
  assign \new_[6621]_  = ~A202 & ~A200;
  assign \new_[6622]_  = ~A199 & \new_[6621]_ ;
  assign \new_[6623]_  = \new_[6622]_  & \new_[6617]_ ;
  assign \new_[6627]_  = A298 & A234;
  assign \new_[6628]_  = A232 & \new_[6627]_ ;
  assign \new_[6632]_  = A302 & ~A301;
  assign \new_[6633]_  = ~A299 & \new_[6632]_ ;
  assign \new_[6634]_  = \new_[6633]_  & \new_[6628]_ ;
  assign \new_[6637]_  = ~A166 & A167;
  assign \new_[6641]_  = ~A202 & ~A200;
  assign \new_[6642]_  = ~A199 & \new_[6641]_ ;
  assign \new_[6643]_  = \new_[6642]_  & \new_[6637]_ ;
  assign \new_[6647]_  = ~A298 & A234;
  assign \new_[6648]_  = A232 & \new_[6647]_ ;
  assign \new_[6652]_  = A302 & ~A301;
  assign \new_[6653]_  = A299 & \new_[6652]_ ;
  assign \new_[6654]_  = \new_[6653]_  & \new_[6648]_ ;
  assign \new_[6657]_  = ~A166 & A167;
  assign \new_[6661]_  = ~A202 & ~A200;
  assign \new_[6662]_  = ~A199 & \new_[6661]_ ;
  assign \new_[6663]_  = \new_[6662]_  & \new_[6657]_ ;
  assign \new_[6667]_  = ~A298 & A234;
  assign \new_[6668]_  = A232 & \new_[6667]_ ;
  assign \new_[6672]_  = ~A302 & A301;
  assign \new_[6673]_  = ~A299 & \new_[6672]_ ;
  assign \new_[6674]_  = \new_[6673]_  & \new_[6668]_ ;
  assign \new_[6677]_  = ~A166 & A167;
  assign \new_[6681]_  = ~A202 & ~A200;
  assign \new_[6682]_  = ~A199 & \new_[6681]_ ;
  assign \new_[6683]_  = \new_[6682]_  & \new_[6677]_ ;
  assign \new_[6687]_  = A265 & A234;
  assign \new_[6688]_  = A232 & \new_[6687]_ ;
  assign \new_[6692]_  = ~A269 & A268;
  assign \new_[6693]_  = A266 & \new_[6692]_ ;
  assign \new_[6694]_  = \new_[6693]_  & \new_[6688]_ ;
  assign \new_[6697]_  = ~A166 & A167;
  assign \new_[6701]_  = ~A202 & ~A200;
  assign \new_[6702]_  = ~A199 & \new_[6701]_ ;
  assign \new_[6703]_  = \new_[6702]_  & \new_[6697]_ ;
  assign \new_[6707]_  = ~A265 & A234;
  assign \new_[6708]_  = A232 & \new_[6707]_ ;
  assign \new_[6712]_  = A269 & ~A268;
  assign \new_[6713]_  = A266 & \new_[6712]_ ;
  assign \new_[6714]_  = \new_[6713]_  & \new_[6708]_ ;
  assign \new_[6717]_  = ~A166 & A167;
  assign \new_[6721]_  = ~A202 & ~A200;
  assign \new_[6722]_  = ~A199 & \new_[6721]_ ;
  assign \new_[6723]_  = \new_[6722]_  & \new_[6717]_ ;
  assign \new_[6727]_  = A265 & A234;
  assign \new_[6728]_  = A232 & \new_[6727]_ ;
  assign \new_[6732]_  = A269 & ~A268;
  assign \new_[6733]_  = ~A266 & \new_[6732]_ ;
  assign \new_[6734]_  = \new_[6733]_  & \new_[6728]_ ;
  assign \new_[6737]_  = ~A166 & A167;
  assign \new_[6741]_  = ~A202 & ~A200;
  assign \new_[6742]_  = ~A199 & \new_[6741]_ ;
  assign \new_[6743]_  = \new_[6742]_  & \new_[6737]_ ;
  assign \new_[6747]_  = ~A265 & A234;
  assign \new_[6748]_  = A232 & \new_[6747]_ ;
  assign \new_[6752]_  = ~A269 & A268;
  assign \new_[6753]_  = ~A266 & \new_[6752]_ ;
  assign \new_[6754]_  = \new_[6753]_  & \new_[6748]_ ;
  assign \new_[6757]_  = ~A166 & A167;
  assign \new_[6761]_  = ~A202 & ~A200;
  assign \new_[6762]_  = ~A199 & \new_[6761]_ ;
  assign \new_[6763]_  = \new_[6762]_  & \new_[6757]_ ;
  assign \new_[6767]_  = A298 & A234;
  assign \new_[6768]_  = A233 & \new_[6767]_ ;
  assign \new_[6772]_  = ~A302 & A301;
  assign \new_[6773]_  = A299 & \new_[6772]_ ;
  assign \new_[6774]_  = \new_[6773]_  & \new_[6768]_ ;
  assign \new_[6777]_  = ~A166 & A167;
  assign \new_[6781]_  = ~A202 & ~A200;
  assign \new_[6782]_  = ~A199 & \new_[6781]_ ;
  assign \new_[6783]_  = \new_[6782]_  & \new_[6777]_ ;
  assign \new_[6787]_  = A298 & A234;
  assign \new_[6788]_  = A233 & \new_[6787]_ ;
  assign \new_[6792]_  = A302 & ~A301;
  assign \new_[6793]_  = ~A299 & \new_[6792]_ ;
  assign \new_[6794]_  = \new_[6793]_  & \new_[6788]_ ;
  assign \new_[6797]_  = ~A166 & A167;
  assign \new_[6801]_  = ~A202 & ~A200;
  assign \new_[6802]_  = ~A199 & \new_[6801]_ ;
  assign \new_[6803]_  = \new_[6802]_  & \new_[6797]_ ;
  assign \new_[6807]_  = ~A298 & A234;
  assign \new_[6808]_  = A233 & \new_[6807]_ ;
  assign \new_[6812]_  = A302 & ~A301;
  assign \new_[6813]_  = A299 & \new_[6812]_ ;
  assign \new_[6814]_  = \new_[6813]_  & \new_[6808]_ ;
  assign \new_[6817]_  = ~A166 & A167;
  assign \new_[6821]_  = ~A202 & ~A200;
  assign \new_[6822]_  = ~A199 & \new_[6821]_ ;
  assign \new_[6823]_  = \new_[6822]_  & \new_[6817]_ ;
  assign \new_[6827]_  = ~A298 & A234;
  assign \new_[6828]_  = A233 & \new_[6827]_ ;
  assign \new_[6832]_  = ~A302 & A301;
  assign \new_[6833]_  = ~A299 & \new_[6832]_ ;
  assign \new_[6834]_  = \new_[6833]_  & \new_[6828]_ ;
  assign \new_[6837]_  = ~A166 & A167;
  assign \new_[6841]_  = ~A202 & ~A200;
  assign \new_[6842]_  = ~A199 & \new_[6841]_ ;
  assign \new_[6843]_  = \new_[6842]_  & \new_[6837]_ ;
  assign \new_[6847]_  = A265 & A234;
  assign \new_[6848]_  = A233 & \new_[6847]_ ;
  assign \new_[6852]_  = ~A269 & A268;
  assign \new_[6853]_  = A266 & \new_[6852]_ ;
  assign \new_[6854]_  = \new_[6853]_  & \new_[6848]_ ;
  assign \new_[6857]_  = ~A166 & A167;
  assign \new_[6861]_  = ~A202 & ~A200;
  assign \new_[6862]_  = ~A199 & \new_[6861]_ ;
  assign \new_[6863]_  = \new_[6862]_  & \new_[6857]_ ;
  assign \new_[6867]_  = ~A265 & A234;
  assign \new_[6868]_  = A233 & \new_[6867]_ ;
  assign \new_[6872]_  = A269 & ~A268;
  assign \new_[6873]_  = A266 & \new_[6872]_ ;
  assign \new_[6874]_  = \new_[6873]_  & \new_[6868]_ ;
  assign \new_[6877]_  = ~A166 & A167;
  assign \new_[6881]_  = ~A202 & ~A200;
  assign \new_[6882]_  = ~A199 & \new_[6881]_ ;
  assign \new_[6883]_  = \new_[6882]_  & \new_[6877]_ ;
  assign \new_[6887]_  = A265 & A234;
  assign \new_[6888]_  = A233 & \new_[6887]_ ;
  assign \new_[6892]_  = A269 & ~A268;
  assign \new_[6893]_  = ~A266 & \new_[6892]_ ;
  assign \new_[6894]_  = \new_[6893]_  & \new_[6888]_ ;
  assign \new_[6897]_  = ~A166 & A167;
  assign \new_[6901]_  = ~A202 & ~A200;
  assign \new_[6902]_  = ~A199 & \new_[6901]_ ;
  assign \new_[6903]_  = \new_[6902]_  & \new_[6897]_ ;
  assign \new_[6907]_  = ~A265 & A234;
  assign \new_[6908]_  = A233 & \new_[6907]_ ;
  assign \new_[6912]_  = ~A269 & A268;
  assign \new_[6913]_  = ~A266 & \new_[6912]_ ;
  assign \new_[6914]_  = \new_[6913]_  & \new_[6908]_ ;
  assign \new_[6917]_  = ~A166 & A167;
  assign \new_[6921]_  = ~A202 & ~A200;
  assign \new_[6922]_  = ~A199 & \new_[6921]_ ;
  assign \new_[6923]_  = \new_[6922]_  & \new_[6917]_ ;
  assign \new_[6927]_  = A235 & A233;
  assign \new_[6928]_  = A232 & \new_[6927]_ ;
  assign \new_[6932]_  = A300 & A299;
  assign \new_[6933]_  = ~A236 & \new_[6932]_ ;
  assign \new_[6934]_  = \new_[6933]_  & \new_[6928]_ ;
  assign \new_[6937]_  = ~A166 & A167;
  assign \new_[6941]_  = ~A202 & ~A200;
  assign \new_[6942]_  = ~A199 & \new_[6941]_ ;
  assign \new_[6943]_  = \new_[6942]_  & \new_[6937]_ ;
  assign \new_[6947]_  = A235 & A233;
  assign \new_[6948]_  = A232 & \new_[6947]_ ;
  assign \new_[6952]_  = A300 & A298;
  assign \new_[6953]_  = ~A236 & \new_[6952]_ ;
  assign \new_[6954]_  = \new_[6953]_  & \new_[6948]_ ;
  assign \new_[6957]_  = ~A166 & A167;
  assign \new_[6961]_  = ~A202 & ~A200;
  assign \new_[6962]_  = ~A199 & \new_[6961]_ ;
  assign \new_[6963]_  = \new_[6962]_  & \new_[6957]_ ;
  assign \new_[6967]_  = A235 & A233;
  assign \new_[6968]_  = A232 & \new_[6967]_ ;
  assign \new_[6972]_  = A267 & A265;
  assign \new_[6973]_  = ~A236 & \new_[6972]_ ;
  assign \new_[6974]_  = \new_[6973]_  & \new_[6968]_ ;
  assign \new_[6977]_  = ~A166 & A167;
  assign \new_[6981]_  = ~A202 & ~A200;
  assign \new_[6982]_  = ~A199 & \new_[6981]_ ;
  assign \new_[6983]_  = \new_[6982]_  & \new_[6977]_ ;
  assign \new_[6987]_  = A235 & A233;
  assign \new_[6988]_  = A232 & \new_[6987]_ ;
  assign \new_[6992]_  = A267 & A266;
  assign \new_[6993]_  = ~A236 & \new_[6992]_ ;
  assign \new_[6994]_  = \new_[6993]_  & \new_[6988]_ ;
  assign \new_[6997]_  = ~A166 & A167;
  assign \new_[7001]_  = ~A202 & ~A200;
  assign \new_[7002]_  = ~A199 & \new_[7001]_ ;
  assign \new_[7003]_  = \new_[7002]_  & \new_[6997]_ ;
  assign \new_[7007]_  = ~A235 & A233;
  assign \new_[7008]_  = ~A232 & \new_[7007]_ ;
  assign \new_[7012]_  = A300 & A299;
  assign \new_[7013]_  = A236 & \new_[7012]_ ;
  assign \new_[7014]_  = \new_[7013]_  & \new_[7008]_ ;
  assign \new_[7017]_  = ~A166 & A167;
  assign \new_[7021]_  = ~A202 & ~A200;
  assign \new_[7022]_  = ~A199 & \new_[7021]_ ;
  assign \new_[7023]_  = \new_[7022]_  & \new_[7017]_ ;
  assign \new_[7027]_  = ~A235 & A233;
  assign \new_[7028]_  = ~A232 & \new_[7027]_ ;
  assign \new_[7032]_  = A300 & A298;
  assign \new_[7033]_  = A236 & \new_[7032]_ ;
  assign \new_[7034]_  = \new_[7033]_  & \new_[7028]_ ;
  assign \new_[7037]_  = ~A166 & A167;
  assign \new_[7041]_  = ~A202 & ~A200;
  assign \new_[7042]_  = ~A199 & \new_[7041]_ ;
  assign \new_[7043]_  = \new_[7042]_  & \new_[7037]_ ;
  assign \new_[7047]_  = ~A235 & A233;
  assign \new_[7048]_  = ~A232 & \new_[7047]_ ;
  assign \new_[7052]_  = A267 & A265;
  assign \new_[7053]_  = A236 & \new_[7052]_ ;
  assign \new_[7054]_  = \new_[7053]_  & \new_[7048]_ ;
  assign \new_[7057]_  = ~A166 & A167;
  assign \new_[7061]_  = ~A202 & ~A200;
  assign \new_[7062]_  = ~A199 & \new_[7061]_ ;
  assign \new_[7063]_  = \new_[7062]_  & \new_[7057]_ ;
  assign \new_[7067]_  = ~A235 & A233;
  assign \new_[7068]_  = ~A232 & \new_[7067]_ ;
  assign \new_[7072]_  = A267 & A266;
  assign \new_[7073]_  = A236 & \new_[7072]_ ;
  assign \new_[7074]_  = \new_[7073]_  & \new_[7068]_ ;
  assign \new_[7077]_  = ~A166 & A167;
  assign \new_[7081]_  = ~A202 & ~A200;
  assign \new_[7082]_  = ~A199 & \new_[7081]_ ;
  assign \new_[7083]_  = \new_[7082]_  & \new_[7077]_ ;
  assign \new_[7087]_  = ~A235 & ~A233;
  assign \new_[7088]_  = A232 & \new_[7087]_ ;
  assign \new_[7092]_  = A300 & A299;
  assign \new_[7093]_  = A236 & \new_[7092]_ ;
  assign \new_[7094]_  = \new_[7093]_  & \new_[7088]_ ;
  assign \new_[7097]_  = ~A166 & A167;
  assign \new_[7101]_  = ~A202 & ~A200;
  assign \new_[7102]_  = ~A199 & \new_[7101]_ ;
  assign \new_[7103]_  = \new_[7102]_  & \new_[7097]_ ;
  assign \new_[7107]_  = ~A235 & ~A233;
  assign \new_[7108]_  = A232 & \new_[7107]_ ;
  assign \new_[7112]_  = A300 & A298;
  assign \new_[7113]_  = A236 & \new_[7112]_ ;
  assign \new_[7114]_  = \new_[7113]_  & \new_[7108]_ ;
  assign \new_[7117]_  = ~A166 & A167;
  assign \new_[7121]_  = ~A202 & ~A200;
  assign \new_[7122]_  = ~A199 & \new_[7121]_ ;
  assign \new_[7123]_  = \new_[7122]_  & \new_[7117]_ ;
  assign \new_[7127]_  = ~A235 & ~A233;
  assign \new_[7128]_  = A232 & \new_[7127]_ ;
  assign \new_[7132]_  = A267 & A265;
  assign \new_[7133]_  = A236 & \new_[7132]_ ;
  assign \new_[7134]_  = \new_[7133]_  & \new_[7128]_ ;
  assign \new_[7137]_  = ~A166 & A167;
  assign \new_[7141]_  = ~A202 & ~A200;
  assign \new_[7142]_  = ~A199 & \new_[7141]_ ;
  assign \new_[7143]_  = \new_[7142]_  & \new_[7137]_ ;
  assign \new_[7147]_  = ~A235 & ~A233;
  assign \new_[7148]_  = A232 & \new_[7147]_ ;
  assign \new_[7152]_  = A267 & A266;
  assign \new_[7153]_  = A236 & \new_[7152]_ ;
  assign \new_[7154]_  = \new_[7153]_  & \new_[7148]_ ;
  assign \new_[7157]_  = ~A166 & A167;
  assign \new_[7161]_  = ~A202 & ~A200;
  assign \new_[7162]_  = ~A199 & \new_[7161]_ ;
  assign \new_[7163]_  = \new_[7162]_  & \new_[7157]_ ;
  assign \new_[7167]_  = A235 & ~A233;
  assign \new_[7168]_  = ~A232 & \new_[7167]_ ;
  assign \new_[7172]_  = A300 & A299;
  assign \new_[7173]_  = ~A236 & \new_[7172]_ ;
  assign \new_[7174]_  = \new_[7173]_  & \new_[7168]_ ;
  assign \new_[7177]_  = ~A166 & A167;
  assign \new_[7181]_  = ~A202 & ~A200;
  assign \new_[7182]_  = ~A199 & \new_[7181]_ ;
  assign \new_[7183]_  = \new_[7182]_  & \new_[7177]_ ;
  assign \new_[7187]_  = A235 & ~A233;
  assign \new_[7188]_  = ~A232 & \new_[7187]_ ;
  assign \new_[7192]_  = A300 & A298;
  assign \new_[7193]_  = ~A236 & \new_[7192]_ ;
  assign \new_[7194]_  = \new_[7193]_  & \new_[7188]_ ;
  assign \new_[7197]_  = ~A166 & A167;
  assign \new_[7201]_  = ~A202 & ~A200;
  assign \new_[7202]_  = ~A199 & \new_[7201]_ ;
  assign \new_[7203]_  = \new_[7202]_  & \new_[7197]_ ;
  assign \new_[7207]_  = A235 & ~A233;
  assign \new_[7208]_  = ~A232 & \new_[7207]_ ;
  assign \new_[7212]_  = A267 & A265;
  assign \new_[7213]_  = ~A236 & \new_[7212]_ ;
  assign \new_[7214]_  = \new_[7213]_  & \new_[7208]_ ;
  assign \new_[7217]_  = ~A166 & A167;
  assign \new_[7221]_  = ~A202 & ~A200;
  assign \new_[7222]_  = ~A199 & \new_[7221]_ ;
  assign \new_[7223]_  = \new_[7222]_  & \new_[7217]_ ;
  assign \new_[7227]_  = A235 & ~A233;
  assign \new_[7228]_  = ~A232 & \new_[7227]_ ;
  assign \new_[7232]_  = A267 & A266;
  assign \new_[7233]_  = ~A236 & \new_[7232]_ ;
  assign \new_[7234]_  = \new_[7233]_  & \new_[7228]_ ;
  assign \new_[7237]_  = ~A166 & A167;
  assign \new_[7241]_  = A203 & ~A200;
  assign \new_[7242]_  = ~A199 & \new_[7241]_ ;
  assign \new_[7243]_  = \new_[7242]_  & \new_[7237]_ ;
  assign \new_[7247]_  = A298 & A234;
  assign \new_[7248]_  = A232 & \new_[7247]_ ;
  assign \new_[7252]_  = ~A302 & A301;
  assign \new_[7253]_  = A299 & \new_[7252]_ ;
  assign \new_[7254]_  = \new_[7253]_  & \new_[7248]_ ;
  assign \new_[7257]_  = ~A166 & A167;
  assign \new_[7261]_  = A203 & ~A200;
  assign \new_[7262]_  = ~A199 & \new_[7261]_ ;
  assign \new_[7263]_  = \new_[7262]_  & \new_[7257]_ ;
  assign \new_[7267]_  = A298 & A234;
  assign \new_[7268]_  = A232 & \new_[7267]_ ;
  assign \new_[7272]_  = A302 & ~A301;
  assign \new_[7273]_  = ~A299 & \new_[7272]_ ;
  assign \new_[7274]_  = \new_[7273]_  & \new_[7268]_ ;
  assign \new_[7277]_  = ~A166 & A167;
  assign \new_[7281]_  = A203 & ~A200;
  assign \new_[7282]_  = ~A199 & \new_[7281]_ ;
  assign \new_[7283]_  = \new_[7282]_  & \new_[7277]_ ;
  assign \new_[7287]_  = ~A298 & A234;
  assign \new_[7288]_  = A232 & \new_[7287]_ ;
  assign \new_[7292]_  = A302 & ~A301;
  assign \new_[7293]_  = A299 & \new_[7292]_ ;
  assign \new_[7294]_  = \new_[7293]_  & \new_[7288]_ ;
  assign \new_[7297]_  = ~A166 & A167;
  assign \new_[7301]_  = A203 & ~A200;
  assign \new_[7302]_  = ~A199 & \new_[7301]_ ;
  assign \new_[7303]_  = \new_[7302]_  & \new_[7297]_ ;
  assign \new_[7307]_  = ~A298 & A234;
  assign \new_[7308]_  = A232 & \new_[7307]_ ;
  assign \new_[7312]_  = ~A302 & A301;
  assign \new_[7313]_  = ~A299 & \new_[7312]_ ;
  assign \new_[7314]_  = \new_[7313]_  & \new_[7308]_ ;
  assign \new_[7317]_  = ~A166 & A167;
  assign \new_[7321]_  = A203 & ~A200;
  assign \new_[7322]_  = ~A199 & \new_[7321]_ ;
  assign \new_[7323]_  = \new_[7322]_  & \new_[7317]_ ;
  assign \new_[7327]_  = A265 & A234;
  assign \new_[7328]_  = A232 & \new_[7327]_ ;
  assign \new_[7332]_  = ~A269 & A268;
  assign \new_[7333]_  = A266 & \new_[7332]_ ;
  assign \new_[7334]_  = \new_[7333]_  & \new_[7328]_ ;
  assign \new_[7337]_  = ~A166 & A167;
  assign \new_[7341]_  = A203 & ~A200;
  assign \new_[7342]_  = ~A199 & \new_[7341]_ ;
  assign \new_[7343]_  = \new_[7342]_  & \new_[7337]_ ;
  assign \new_[7347]_  = ~A265 & A234;
  assign \new_[7348]_  = A232 & \new_[7347]_ ;
  assign \new_[7352]_  = A269 & ~A268;
  assign \new_[7353]_  = A266 & \new_[7352]_ ;
  assign \new_[7354]_  = \new_[7353]_  & \new_[7348]_ ;
  assign \new_[7357]_  = ~A166 & A167;
  assign \new_[7361]_  = A203 & ~A200;
  assign \new_[7362]_  = ~A199 & \new_[7361]_ ;
  assign \new_[7363]_  = \new_[7362]_  & \new_[7357]_ ;
  assign \new_[7367]_  = A265 & A234;
  assign \new_[7368]_  = A232 & \new_[7367]_ ;
  assign \new_[7372]_  = A269 & ~A268;
  assign \new_[7373]_  = ~A266 & \new_[7372]_ ;
  assign \new_[7374]_  = \new_[7373]_  & \new_[7368]_ ;
  assign \new_[7377]_  = ~A166 & A167;
  assign \new_[7381]_  = A203 & ~A200;
  assign \new_[7382]_  = ~A199 & \new_[7381]_ ;
  assign \new_[7383]_  = \new_[7382]_  & \new_[7377]_ ;
  assign \new_[7387]_  = ~A265 & A234;
  assign \new_[7388]_  = A232 & \new_[7387]_ ;
  assign \new_[7392]_  = ~A269 & A268;
  assign \new_[7393]_  = ~A266 & \new_[7392]_ ;
  assign \new_[7394]_  = \new_[7393]_  & \new_[7388]_ ;
  assign \new_[7397]_  = ~A166 & A167;
  assign \new_[7401]_  = A203 & ~A200;
  assign \new_[7402]_  = ~A199 & \new_[7401]_ ;
  assign \new_[7403]_  = \new_[7402]_  & \new_[7397]_ ;
  assign \new_[7407]_  = A298 & A234;
  assign \new_[7408]_  = A233 & \new_[7407]_ ;
  assign \new_[7412]_  = ~A302 & A301;
  assign \new_[7413]_  = A299 & \new_[7412]_ ;
  assign \new_[7414]_  = \new_[7413]_  & \new_[7408]_ ;
  assign \new_[7417]_  = ~A166 & A167;
  assign \new_[7421]_  = A203 & ~A200;
  assign \new_[7422]_  = ~A199 & \new_[7421]_ ;
  assign \new_[7423]_  = \new_[7422]_  & \new_[7417]_ ;
  assign \new_[7427]_  = A298 & A234;
  assign \new_[7428]_  = A233 & \new_[7427]_ ;
  assign \new_[7432]_  = A302 & ~A301;
  assign \new_[7433]_  = ~A299 & \new_[7432]_ ;
  assign \new_[7434]_  = \new_[7433]_  & \new_[7428]_ ;
  assign \new_[7437]_  = ~A166 & A167;
  assign \new_[7441]_  = A203 & ~A200;
  assign \new_[7442]_  = ~A199 & \new_[7441]_ ;
  assign \new_[7443]_  = \new_[7442]_  & \new_[7437]_ ;
  assign \new_[7447]_  = ~A298 & A234;
  assign \new_[7448]_  = A233 & \new_[7447]_ ;
  assign \new_[7452]_  = A302 & ~A301;
  assign \new_[7453]_  = A299 & \new_[7452]_ ;
  assign \new_[7454]_  = \new_[7453]_  & \new_[7448]_ ;
  assign \new_[7457]_  = ~A166 & A167;
  assign \new_[7461]_  = A203 & ~A200;
  assign \new_[7462]_  = ~A199 & \new_[7461]_ ;
  assign \new_[7463]_  = \new_[7462]_  & \new_[7457]_ ;
  assign \new_[7467]_  = ~A298 & A234;
  assign \new_[7468]_  = A233 & \new_[7467]_ ;
  assign \new_[7472]_  = ~A302 & A301;
  assign \new_[7473]_  = ~A299 & \new_[7472]_ ;
  assign \new_[7474]_  = \new_[7473]_  & \new_[7468]_ ;
  assign \new_[7477]_  = ~A166 & A167;
  assign \new_[7481]_  = A203 & ~A200;
  assign \new_[7482]_  = ~A199 & \new_[7481]_ ;
  assign \new_[7483]_  = \new_[7482]_  & \new_[7477]_ ;
  assign \new_[7487]_  = A265 & A234;
  assign \new_[7488]_  = A233 & \new_[7487]_ ;
  assign \new_[7492]_  = ~A269 & A268;
  assign \new_[7493]_  = A266 & \new_[7492]_ ;
  assign \new_[7494]_  = \new_[7493]_  & \new_[7488]_ ;
  assign \new_[7497]_  = ~A166 & A167;
  assign \new_[7501]_  = A203 & ~A200;
  assign \new_[7502]_  = ~A199 & \new_[7501]_ ;
  assign \new_[7503]_  = \new_[7502]_  & \new_[7497]_ ;
  assign \new_[7507]_  = ~A265 & A234;
  assign \new_[7508]_  = A233 & \new_[7507]_ ;
  assign \new_[7512]_  = A269 & ~A268;
  assign \new_[7513]_  = A266 & \new_[7512]_ ;
  assign \new_[7514]_  = \new_[7513]_  & \new_[7508]_ ;
  assign \new_[7517]_  = ~A166 & A167;
  assign \new_[7521]_  = A203 & ~A200;
  assign \new_[7522]_  = ~A199 & \new_[7521]_ ;
  assign \new_[7523]_  = \new_[7522]_  & \new_[7517]_ ;
  assign \new_[7527]_  = A265 & A234;
  assign \new_[7528]_  = A233 & \new_[7527]_ ;
  assign \new_[7532]_  = A269 & ~A268;
  assign \new_[7533]_  = ~A266 & \new_[7532]_ ;
  assign \new_[7534]_  = \new_[7533]_  & \new_[7528]_ ;
  assign \new_[7537]_  = ~A166 & A167;
  assign \new_[7541]_  = A203 & ~A200;
  assign \new_[7542]_  = ~A199 & \new_[7541]_ ;
  assign \new_[7543]_  = \new_[7542]_  & \new_[7537]_ ;
  assign \new_[7547]_  = ~A265 & A234;
  assign \new_[7548]_  = A233 & \new_[7547]_ ;
  assign \new_[7552]_  = ~A269 & A268;
  assign \new_[7553]_  = ~A266 & \new_[7552]_ ;
  assign \new_[7554]_  = \new_[7553]_  & \new_[7548]_ ;
  assign \new_[7557]_  = ~A166 & A167;
  assign \new_[7561]_  = A203 & ~A200;
  assign \new_[7562]_  = ~A199 & \new_[7561]_ ;
  assign \new_[7563]_  = \new_[7562]_  & \new_[7557]_ ;
  assign \new_[7567]_  = A235 & A233;
  assign \new_[7568]_  = A232 & \new_[7567]_ ;
  assign \new_[7572]_  = A300 & A299;
  assign \new_[7573]_  = ~A236 & \new_[7572]_ ;
  assign \new_[7574]_  = \new_[7573]_  & \new_[7568]_ ;
  assign \new_[7577]_  = ~A166 & A167;
  assign \new_[7581]_  = A203 & ~A200;
  assign \new_[7582]_  = ~A199 & \new_[7581]_ ;
  assign \new_[7583]_  = \new_[7582]_  & \new_[7577]_ ;
  assign \new_[7587]_  = A235 & A233;
  assign \new_[7588]_  = A232 & \new_[7587]_ ;
  assign \new_[7592]_  = A300 & A298;
  assign \new_[7593]_  = ~A236 & \new_[7592]_ ;
  assign \new_[7594]_  = \new_[7593]_  & \new_[7588]_ ;
  assign \new_[7597]_  = ~A166 & A167;
  assign \new_[7601]_  = A203 & ~A200;
  assign \new_[7602]_  = ~A199 & \new_[7601]_ ;
  assign \new_[7603]_  = \new_[7602]_  & \new_[7597]_ ;
  assign \new_[7607]_  = A235 & A233;
  assign \new_[7608]_  = A232 & \new_[7607]_ ;
  assign \new_[7612]_  = A267 & A265;
  assign \new_[7613]_  = ~A236 & \new_[7612]_ ;
  assign \new_[7614]_  = \new_[7613]_  & \new_[7608]_ ;
  assign \new_[7617]_  = ~A166 & A167;
  assign \new_[7621]_  = A203 & ~A200;
  assign \new_[7622]_  = ~A199 & \new_[7621]_ ;
  assign \new_[7623]_  = \new_[7622]_  & \new_[7617]_ ;
  assign \new_[7627]_  = A235 & A233;
  assign \new_[7628]_  = A232 & \new_[7627]_ ;
  assign \new_[7632]_  = A267 & A266;
  assign \new_[7633]_  = ~A236 & \new_[7632]_ ;
  assign \new_[7634]_  = \new_[7633]_  & \new_[7628]_ ;
  assign \new_[7637]_  = ~A166 & A167;
  assign \new_[7641]_  = A203 & ~A200;
  assign \new_[7642]_  = ~A199 & \new_[7641]_ ;
  assign \new_[7643]_  = \new_[7642]_  & \new_[7637]_ ;
  assign \new_[7647]_  = ~A235 & A233;
  assign \new_[7648]_  = ~A232 & \new_[7647]_ ;
  assign \new_[7652]_  = A300 & A299;
  assign \new_[7653]_  = A236 & \new_[7652]_ ;
  assign \new_[7654]_  = \new_[7653]_  & \new_[7648]_ ;
  assign \new_[7657]_  = ~A166 & A167;
  assign \new_[7661]_  = A203 & ~A200;
  assign \new_[7662]_  = ~A199 & \new_[7661]_ ;
  assign \new_[7663]_  = \new_[7662]_  & \new_[7657]_ ;
  assign \new_[7667]_  = ~A235 & A233;
  assign \new_[7668]_  = ~A232 & \new_[7667]_ ;
  assign \new_[7672]_  = A300 & A298;
  assign \new_[7673]_  = A236 & \new_[7672]_ ;
  assign \new_[7674]_  = \new_[7673]_  & \new_[7668]_ ;
  assign \new_[7677]_  = ~A166 & A167;
  assign \new_[7681]_  = A203 & ~A200;
  assign \new_[7682]_  = ~A199 & \new_[7681]_ ;
  assign \new_[7683]_  = \new_[7682]_  & \new_[7677]_ ;
  assign \new_[7687]_  = ~A235 & A233;
  assign \new_[7688]_  = ~A232 & \new_[7687]_ ;
  assign \new_[7692]_  = A267 & A265;
  assign \new_[7693]_  = A236 & \new_[7692]_ ;
  assign \new_[7694]_  = \new_[7693]_  & \new_[7688]_ ;
  assign \new_[7697]_  = ~A166 & A167;
  assign \new_[7701]_  = A203 & ~A200;
  assign \new_[7702]_  = ~A199 & \new_[7701]_ ;
  assign \new_[7703]_  = \new_[7702]_  & \new_[7697]_ ;
  assign \new_[7707]_  = ~A235 & A233;
  assign \new_[7708]_  = ~A232 & \new_[7707]_ ;
  assign \new_[7712]_  = A267 & A266;
  assign \new_[7713]_  = A236 & \new_[7712]_ ;
  assign \new_[7714]_  = \new_[7713]_  & \new_[7708]_ ;
  assign \new_[7717]_  = ~A166 & A167;
  assign \new_[7721]_  = A203 & ~A200;
  assign \new_[7722]_  = ~A199 & \new_[7721]_ ;
  assign \new_[7723]_  = \new_[7722]_  & \new_[7717]_ ;
  assign \new_[7727]_  = ~A235 & ~A233;
  assign \new_[7728]_  = A232 & \new_[7727]_ ;
  assign \new_[7732]_  = A300 & A299;
  assign \new_[7733]_  = A236 & \new_[7732]_ ;
  assign \new_[7734]_  = \new_[7733]_  & \new_[7728]_ ;
  assign \new_[7737]_  = ~A166 & A167;
  assign \new_[7741]_  = A203 & ~A200;
  assign \new_[7742]_  = ~A199 & \new_[7741]_ ;
  assign \new_[7743]_  = \new_[7742]_  & \new_[7737]_ ;
  assign \new_[7747]_  = ~A235 & ~A233;
  assign \new_[7748]_  = A232 & \new_[7747]_ ;
  assign \new_[7752]_  = A300 & A298;
  assign \new_[7753]_  = A236 & \new_[7752]_ ;
  assign \new_[7754]_  = \new_[7753]_  & \new_[7748]_ ;
  assign \new_[7757]_  = ~A166 & A167;
  assign \new_[7761]_  = A203 & ~A200;
  assign \new_[7762]_  = ~A199 & \new_[7761]_ ;
  assign \new_[7763]_  = \new_[7762]_  & \new_[7757]_ ;
  assign \new_[7767]_  = ~A235 & ~A233;
  assign \new_[7768]_  = A232 & \new_[7767]_ ;
  assign \new_[7772]_  = A267 & A265;
  assign \new_[7773]_  = A236 & \new_[7772]_ ;
  assign \new_[7774]_  = \new_[7773]_  & \new_[7768]_ ;
  assign \new_[7777]_  = ~A166 & A167;
  assign \new_[7781]_  = A203 & ~A200;
  assign \new_[7782]_  = ~A199 & \new_[7781]_ ;
  assign \new_[7783]_  = \new_[7782]_  & \new_[7777]_ ;
  assign \new_[7787]_  = ~A235 & ~A233;
  assign \new_[7788]_  = A232 & \new_[7787]_ ;
  assign \new_[7792]_  = A267 & A266;
  assign \new_[7793]_  = A236 & \new_[7792]_ ;
  assign \new_[7794]_  = \new_[7793]_  & \new_[7788]_ ;
  assign \new_[7797]_  = ~A166 & A167;
  assign \new_[7801]_  = A203 & ~A200;
  assign \new_[7802]_  = ~A199 & \new_[7801]_ ;
  assign \new_[7803]_  = \new_[7802]_  & \new_[7797]_ ;
  assign \new_[7807]_  = A235 & ~A233;
  assign \new_[7808]_  = ~A232 & \new_[7807]_ ;
  assign \new_[7812]_  = A300 & A299;
  assign \new_[7813]_  = ~A236 & \new_[7812]_ ;
  assign \new_[7814]_  = \new_[7813]_  & \new_[7808]_ ;
  assign \new_[7817]_  = ~A166 & A167;
  assign \new_[7821]_  = A203 & ~A200;
  assign \new_[7822]_  = ~A199 & \new_[7821]_ ;
  assign \new_[7823]_  = \new_[7822]_  & \new_[7817]_ ;
  assign \new_[7827]_  = A235 & ~A233;
  assign \new_[7828]_  = ~A232 & \new_[7827]_ ;
  assign \new_[7832]_  = A300 & A298;
  assign \new_[7833]_  = ~A236 & \new_[7832]_ ;
  assign \new_[7834]_  = \new_[7833]_  & \new_[7828]_ ;
  assign \new_[7837]_  = ~A166 & A167;
  assign \new_[7841]_  = A203 & ~A200;
  assign \new_[7842]_  = ~A199 & \new_[7841]_ ;
  assign \new_[7843]_  = \new_[7842]_  & \new_[7837]_ ;
  assign \new_[7847]_  = A235 & ~A233;
  assign \new_[7848]_  = ~A232 & \new_[7847]_ ;
  assign \new_[7852]_  = A267 & A265;
  assign \new_[7853]_  = ~A236 & \new_[7852]_ ;
  assign \new_[7854]_  = \new_[7853]_  & \new_[7848]_ ;
  assign \new_[7857]_  = ~A166 & A167;
  assign \new_[7861]_  = A203 & ~A200;
  assign \new_[7862]_  = ~A199 & \new_[7861]_ ;
  assign \new_[7863]_  = \new_[7862]_  & \new_[7857]_ ;
  assign \new_[7867]_  = A235 & ~A233;
  assign \new_[7868]_  = ~A232 & \new_[7867]_ ;
  assign \new_[7872]_  = A267 & A266;
  assign \new_[7873]_  = ~A236 & \new_[7872]_ ;
  assign \new_[7874]_  = \new_[7873]_  & \new_[7868]_ ;
  assign \new_[7877]_  = A168 & A170;
  assign \new_[7881]_  = ~A199 & A166;
  assign \new_[7882]_  = ~A167 & \new_[7881]_ ;
  assign \new_[7883]_  = \new_[7882]_  & \new_[7877]_ ;
  assign \new_[7887]_  = A232 & ~A202;
  assign \new_[7888]_  = ~A200 & \new_[7887]_ ;
  assign \new_[7892]_  = A300 & A299;
  assign \new_[7893]_  = A234 & \new_[7892]_ ;
  assign \new_[7894]_  = \new_[7893]_  & \new_[7888]_ ;
  assign \new_[7897]_  = A168 & A170;
  assign \new_[7901]_  = ~A199 & A166;
  assign \new_[7902]_  = ~A167 & \new_[7901]_ ;
  assign \new_[7903]_  = \new_[7902]_  & \new_[7897]_ ;
  assign \new_[7907]_  = A232 & ~A202;
  assign \new_[7908]_  = ~A200 & \new_[7907]_ ;
  assign \new_[7912]_  = A300 & A298;
  assign \new_[7913]_  = A234 & \new_[7912]_ ;
  assign \new_[7914]_  = \new_[7913]_  & \new_[7908]_ ;
  assign \new_[7917]_  = A168 & A170;
  assign \new_[7921]_  = ~A199 & A166;
  assign \new_[7922]_  = ~A167 & \new_[7921]_ ;
  assign \new_[7923]_  = \new_[7922]_  & \new_[7917]_ ;
  assign \new_[7927]_  = A232 & ~A202;
  assign \new_[7928]_  = ~A200 & \new_[7927]_ ;
  assign \new_[7932]_  = A267 & A265;
  assign \new_[7933]_  = A234 & \new_[7932]_ ;
  assign \new_[7934]_  = \new_[7933]_  & \new_[7928]_ ;
  assign \new_[7937]_  = A168 & A170;
  assign \new_[7941]_  = ~A199 & A166;
  assign \new_[7942]_  = ~A167 & \new_[7941]_ ;
  assign \new_[7943]_  = \new_[7942]_  & \new_[7937]_ ;
  assign \new_[7947]_  = A232 & ~A202;
  assign \new_[7948]_  = ~A200 & \new_[7947]_ ;
  assign \new_[7952]_  = A267 & A266;
  assign \new_[7953]_  = A234 & \new_[7952]_ ;
  assign \new_[7954]_  = \new_[7953]_  & \new_[7948]_ ;
  assign \new_[7957]_  = A168 & A170;
  assign \new_[7961]_  = ~A199 & A166;
  assign \new_[7962]_  = ~A167 & \new_[7961]_ ;
  assign \new_[7963]_  = \new_[7962]_  & \new_[7957]_ ;
  assign \new_[7967]_  = A233 & ~A202;
  assign \new_[7968]_  = ~A200 & \new_[7967]_ ;
  assign \new_[7972]_  = A300 & A299;
  assign \new_[7973]_  = A234 & \new_[7972]_ ;
  assign \new_[7974]_  = \new_[7973]_  & \new_[7968]_ ;
  assign \new_[7977]_  = A168 & A170;
  assign \new_[7981]_  = ~A199 & A166;
  assign \new_[7982]_  = ~A167 & \new_[7981]_ ;
  assign \new_[7983]_  = \new_[7982]_  & \new_[7977]_ ;
  assign \new_[7987]_  = A233 & ~A202;
  assign \new_[7988]_  = ~A200 & \new_[7987]_ ;
  assign \new_[7992]_  = A300 & A298;
  assign \new_[7993]_  = A234 & \new_[7992]_ ;
  assign \new_[7994]_  = \new_[7993]_  & \new_[7988]_ ;
  assign \new_[7997]_  = A168 & A170;
  assign \new_[8001]_  = ~A199 & A166;
  assign \new_[8002]_  = ~A167 & \new_[8001]_ ;
  assign \new_[8003]_  = \new_[8002]_  & \new_[7997]_ ;
  assign \new_[8007]_  = A233 & ~A202;
  assign \new_[8008]_  = ~A200 & \new_[8007]_ ;
  assign \new_[8012]_  = A267 & A265;
  assign \new_[8013]_  = A234 & \new_[8012]_ ;
  assign \new_[8014]_  = \new_[8013]_  & \new_[8008]_ ;
  assign \new_[8017]_  = A168 & A170;
  assign \new_[8021]_  = ~A199 & A166;
  assign \new_[8022]_  = ~A167 & \new_[8021]_ ;
  assign \new_[8023]_  = \new_[8022]_  & \new_[8017]_ ;
  assign \new_[8027]_  = A233 & ~A202;
  assign \new_[8028]_  = ~A200 & \new_[8027]_ ;
  assign \new_[8032]_  = A267 & A266;
  assign \new_[8033]_  = A234 & \new_[8032]_ ;
  assign \new_[8034]_  = \new_[8033]_  & \new_[8028]_ ;
  assign \new_[8037]_  = A168 & A170;
  assign \new_[8041]_  = ~A199 & A166;
  assign \new_[8042]_  = ~A167 & \new_[8041]_ ;
  assign \new_[8043]_  = \new_[8042]_  & \new_[8037]_ ;
  assign \new_[8047]_  = A232 & A203;
  assign \new_[8048]_  = ~A200 & \new_[8047]_ ;
  assign \new_[8052]_  = A300 & A299;
  assign \new_[8053]_  = A234 & \new_[8052]_ ;
  assign \new_[8054]_  = \new_[8053]_  & \new_[8048]_ ;
  assign \new_[8057]_  = A168 & A170;
  assign \new_[8061]_  = ~A199 & A166;
  assign \new_[8062]_  = ~A167 & \new_[8061]_ ;
  assign \new_[8063]_  = \new_[8062]_  & \new_[8057]_ ;
  assign \new_[8067]_  = A232 & A203;
  assign \new_[8068]_  = ~A200 & \new_[8067]_ ;
  assign \new_[8072]_  = A300 & A298;
  assign \new_[8073]_  = A234 & \new_[8072]_ ;
  assign \new_[8074]_  = \new_[8073]_  & \new_[8068]_ ;
  assign \new_[8077]_  = A168 & A170;
  assign \new_[8081]_  = ~A199 & A166;
  assign \new_[8082]_  = ~A167 & \new_[8081]_ ;
  assign \new_[8083]_  = \new_[8082]_  & \new_[8077]_ ;
  assign \new_[8087]_  = A232 & A203;
  assign \new_[8088]_  = ~A200 & \new_[8087]_ ;
  assign \new_[8092]_  = A267 & A265;
  assign \new_[8093]_  = A234 & \new_[8092]_ ;
  assign \new_[8094]_  = \new_[8093]_  & \new_[8088]_ ;
  assign \new_[8097]_  = A168 & A170;
  assign \new_[8101]_  = ~A199 & A166;
  assign \new_[8102]_  = ~A167 & \new_[8101]_ ;
  assign \new_[8103]_  = \new_[8102]_  & \new_[8097]_ ;
  assign \new_[8107]_  = A232 & A203;
  assign \new_[8108]_  = ~A200 & \new_[8107]_ ;
  assign \new_[8112]_  = A267 & A266;
  assign \new_[8113]_  = A234 & \new_[8112]_ ;
  assign \new_[8114]_  = \new_[8113]_  & \new_[8108]_ ;
  assign \new_[8117]_  = A168 & A170;
  assign \new_[8121]_  = ~A199 & A166;
  assign \new_[8122]_  = ~A167 & \new_[8121]_ ;
  assign \new_[8123]_  = \new_[8122]_  & \new_[8117]_ ;
  assign \new_[8127]_  = A233 & A203;
  assign \new_[8128]_  = ~A200 & \new_[8127]_ ;
  assign \new_[8132]_  = A300 & A299;
  assign \new_[8133]_  = A234 & \new_[8132]_ ;
  assign \new_[8134]_  = \new_[8133]_  & \new_[8128]_ ;
  assign \new_[8137]_  = A168 & A170;
  assign \new_[8141]_  = ~A199 & A166;
  assign \new_[8142]_  = ~A167 & \new_[8141]_ ;
  assign \new_[8143]_  = \new_[8142]_  & \new_[8137]_ ;
  assign \new_[8147]_  = A233 & A203;
  assign \new_[8148]_  = ~A200 & \new_[8147]_ ;
  assign \new_[8152]_  = A300 & A298;
  assign \new_[8153]_  = A234 & \new_[8152]_ ;
  assign \new_[8154]_  = \new_[8153]_  & \new_[8148]_ ;
  assign \new_[8157]_  = A168 & A170;
  assign \new_[8161]_  = ~A199 & A166;
  assign \new_[8162]_  = ~A167 & \new_[8161]_ ;
  assign \new_[8163]_  = \new_[8162]_  & \new_[8157]_ ;
  assign \new_[8167]_  = A233 & A203;
  assign \new_[8168]_  = ~A200 & \new_[8167]_ ;
  assign \new_[8172]_  = A267 & A265;
  assign \new_[8173]_  = A234 & \new_[8172]_ ;
  assign \new_[8174]_  = \new_[8173]_  & \new_[8168]_ ;
  assign \new_[8177]_  = A168 & A170;
  assign \new_[8181]_  = ~A199 & A166;
  assign \new_[8182]_  = ~A167 & \new_[8181]_ ;
  assign \new_[8183]_  = \new_[8182]_  & \new_[8177]_ ;
  assign \new_[8187]_  = A233 & A203;
  assign \new_[8188]_  = ~A200 & \new_[8187]_ ;
  assign \new_[8192]_  = A267 & A266;
  assign \new_[8193]_  = A234 & \new_[8192]_ ;
  assign \new_[8194]_  = \new_[8193]_  & \new_[8188]_ ;
  assign \new_[8197]_  = A168 & A169;
  assign \new_[8201]_  = ~A199 & A166;
  assign \new_[8202]_  = ~A167 & \new_[8201]_ ;
  assign \new_[8203]_  = \new_[8202]_  & \new_[8197]_ ;
  assign \new_[8207]_  = A232 & ~A202;
  assign \new_[8208]_  = ~A200 & \new_[8207]_ ;
  assign \new_[8212]_  = A300 & A299;
  assign \new_[8213]_  = A234 & \new_[8212]_ ;
  assign \new_[8214]_  = \new_[8213]_  & \new_[8208]_ ;
  assign \new_[8217]_  = A168 & A169;
  assign \new_[8221]_  = ~A199 & A166;
  assign \new_[8222]_  = ~A167 & \new_[8221]_ ;
  assign \new_[8223]_  = \new_[8222]_  & \new_[8217]_ ;
  assign \new_[8227]_  = A232 & ~A202;
  assign \new_[8228]_  = ~A200 & \new_[8227]_ ;
  assign \new_[8232]_  = A300 & A298;
  assign \new_[8233]_  = A234 & \new_[8232]_ ;
  assign \new_[8234]_  = \new_[8233]_  & \new_[8228]_ ;
  assign \new_[8237]_  = A168 & A169;
  assign \new_[8241]_  = ~A199 & A166;
  assign \new_[8242]_  = ~A167 & \new_[8241]_ ;
  assign \new_[8243]_  = \new_[8242]_  & \new_[8237]_ ;
  assign \new_[8247]_  = A232 & ~A202;
  assign \new_[8248]_  = ~A200 & \new_[8247]_ ;
  assign \new_[8252]_  = A267 & A265;
  assign \new_[8253]_  = A234 & \new_[8252]_ ;
  assign \new_[8254]_  = \new_[8253]_  & \new_[8248]_ ;
  assign \new_[8257]_  = A168 & A169;
  assign \new_[8261]_  = ~A199 & A166;
  assign \new_[8262]_  = ~A167 & \new_[8261]_ ;
  assign \new_[8263]_  = \new_[8262]_  & \new_[8257]_ ;
  assign \new_[8267]_  = A232 & ~A202;
  assign \new_[8268]_  = ~A200 & \new_[8267]_ ;
  assign \new_[8272]_  = A267 & A266;
  assign \new_[8273]_  = A234 & \new_[8272]_ ;
  assign \new_[8274]_  = \new_[8273]_  & \new_[8268]_ ;
  assign \new_[8277]_  = A168 & A169;
  assign \new_[8281]_  = ~A199 & A166;
  assign \new_[8282]_  = ~A167 & \new_[8281]_ ;
  assign \new_[8283]_  = \new_[8282]_  & \new_[8277]_ ;
  assign \new_[8287]_  = A233 & ~A202;
  assign \new_[8288]_  = ~A200 & \new_[8287]_ ;
  assign \new_[8292]_  = A300 & A299;
  assign \new_[8293]_  = A234 & \new_[8292]_ ;
  assign \new_[8294]_  = \new_[8293]_  & \new_[8288]_ ;
  assign \new_[8297]_  = A168 & A169;
  assign \new_[8301]_  = ~A199 & A166;
  assign \new_[8302]_  = ~A167 & \new_[8301]_ ;
  assign \new_[8303]_  = \new_[8302]_  & \new_[8297]_ ;
  assign \new_[8307]_  = A233 & ~A202;
  assign \new_[8308]_  = ~A200 & \new_[8307]_ ;
  assign \new_[8312]_  = A300 & A298;
  assign \new_[8313]_  = A234 & \new_[8312]_ ;
  assign \new_[8314]_  = \new_[8313]_  & \new_[8308]_ ;
  assign \new_[8317]_  = A168 & A169;
  assign \new_[8321]_  = ~A199 & A166;
  assign \new_[8322]_  = ~A167 & \new_[8321]_ ;
  assign \new_[8323]_  = \new_[8322]_  & \new_[8317]_ ;
  assign \new_[8327]_  = A233 & ~A202;
  assign \new_[8328]_  = ~A200 & \new_[8327]_ ;
  assign \new_[8332]_  = A267 & A265;
  assign \new_[8333]_  = A234 & \new_[8332]_ ;
  assign \new_[8334]_  = \new_[8333]_  & \new_[8328]_ ;
  assign \new_[8337]_  = A168 & A169;
  assign \new_[8341]_  = ~A199 & A166;
  assign \new_[8342]_  = ~A167 & \new_[8341]_ ;
  assign \new_[8343]_  = \new_[8342]_  & \new_[8337]_ ;
  assign \new_[8347]_  = A233 & ~A202;
  assign \new_[8348]_  = ~A200 & \new_[8347]_ ;
  assign \new_[8352]_  = A267 & A266;
  assign \new_[8353]_  = A234 & \new_[8352]_ ;
  assign \new_[8354]_  = \new_[8353]_  & \new_[8348]_ ;
  assign \new_[8357]_  = A168 & A169;
  assign \new_[8361]_  = ~A199 & A166;
  assign \new_[8362]_  = ~A167 & \new_[8361]_ ;
  assign \new_[8363]_  = \new_[8362]_  & \new_[8357]_ ;
  assign \new_[8367]_  = A232 & A203;
  assign \new_[8368]_  = ~A200 & \new_[8367]_ ;
  assign \new_[8372]_  = A300 & A299;
  assign \new_[8373]_  = A234 & \new_[8372]_ ;
  assign \new_[8374]_  = \new_[8373]_  & \new_[8368]_ ;
  assign \new_[8377]_  = A168 & A169;
  assign \new_[8381]_  = ~A199 & A166;
  assign \new_[8382]_  = ~A167 & \new_[8381]_ ;
  assign \new_[8383]_  = \new_[8382]_  & \new_[8377]_ ;
  assign \new_[8387]_  = A232 & A203;
  assign \new_[8388]_  = ~A200 & \new_[8387]_ ;
  assign \new_[8392]_  = A300 & A298;
  assign \new_[8393]_  = A234 & \new_[8392]_ ;
  assign \new_[8394]_  = \new_[8393]_  & \new_[8388]_ ;
  assign \new_[8397]_  = A168 & A169;
  assign \new_[8401]_  = ~A199 & A166;
  assign \new_[8402]_  = ~A167 & \new_[8401]_ ;
  assign \new_[8403]_  = \new_[8402]_  & \new_[8397]_ ;
  assign \new_[8407]_  = A232 & A203;
  assign \new_[8408]_  = ~A200 & \new_[8407]_ ;
  assign \new_[8412]_  = A267 & A265;
  assign \new_[8413]_  = A234 & \new_[8412]_ ;
  assign \new_[8414]_  = \new_[8413]_  & \new_[8408]_ ;
  assign \new_[8417]_  = A168 & A169;
  assign \new_[8421]_  = ~A199 & A166;
  assign \new_[8422]_  = ~A167 & \new_[8421]_ ;
  assign \new_[8423]_  = \new_[8422]_  & \new_[8417]_ ;
  assign \new_[8427]_  = A232 & A203;
  assign \new_[8428]_  = ~A200 & \new_[8427]_ ;
  assign \new_[8432]_  = A267 & A266;
  assign \new_[8433]_  = A234 & \new_[8432]_ ;
  assign \new_[8434]_  = \new_[8433]_  & \new_[8428]_ ;
  assign \new_[8437]_  = A168 & A169;
  assign \new_[8441]_  = ~A199 & A166;
  assign \new_[8442]_  = ~A167 & \new_[8441]_ ;
  assign \new_[8443]_  = \new_[8442]_  & \new_[8437]_ ;
  assign \new_[8447]_  = A233 & A203;
  assign \new_[8448]_  = ~A200 & \new_[8447]_ ;
  assign \new_[8452]_  = A300 & A299;
  assign \new_[8453]_  = A234 & \new_[8452]_ ;
  assign \new_[8454]_  = \new_[8453]_  & \new_[8448]_ ;
  assign \new_[8457]_  = A168 & A169;
  assign \new_[8461]_  = ~A199 & A166;
  assign \new_[8462]_  = ~A167 & \new_[8461]_ ;
  assign \new_[8463]_  = \new_[8462]_  & \new_[8457]_ ;
  assign \new_[8467]_  = A233 & A203;
  assign \new_[8468]_  = ~A200 & \new_[8467]_ ;
  assign \new_[8472]_  = A300 & A298;
  assign \new_[8473]_  = A234 & \new_[8472]_ ;
  assign \new_[8474]_  = \new_[8473]_  & \new_[8468]_ ;
  assign \new_[8477]_  = A168 & A169;
  assign \new_[8481]_  = ~A199 & A166;
  assign \new_[8482]_  = ~A167 & \new_[8481]_ ;
  assign \new_[8483]_  = \new_[8482]_  & \new_[8477]_ ;
  assign \new_[8487]_  = A233 & A203;
  assign \new_[8488]_  = ~A200 & \new_[8487]_ ;
  assign \new_[8492]_  = A267 & A265;
  assign \new_[8493]_  = A234 & \new_[8492]_ ;
  assign \new_[8494]_  = \new_[8493]_  & \new_[8488]_ ;
  assign \new_[8497]_  = A168 & A169;
  assign \new_[8501]_  = ~A199 & A166;
  assign \new_[8502]_  = ~A167 & \new_[8501]_ ;
  assign \new_[8503]_  = \new_[8502]_  & \new_[8497]_ ;
  assign \new_[8507]_  = A233 & A203;
  assign \new_[8508]_  = ~A200 & \new_[8507]_ ;
  assign \new_[8512]_  = A267 & A266;
  assign \new_[8513]_  = A234 & \new_[8512]_ ;
  assign \new_[8514]_  = \new_[8513]_  & \new_[8508]_ ;
  assign \new_[8518]_  = A199 & ~A166;
  assign \new_[8519]_  = A167 & \new_[8518]_ ;
  assign \new_[8523]_  = ~A202 & ~A201;
  assign \new_[8524]_  = A200 & \new_[8523]_ ;
  assign \new_[8525]_  = \new_[8524]_  & \new_[8519]_ ;
  assign \new_[8529]_  = A298 & A234;
  assign \new_[8530]_  = A232 & \new_[8529]_ ;
  assign \new_[8534]_  = ~A302 & A301;
  assign \new_[8535]_  = A299 & \new_[8534]_ ;
  assign \new_[8536]_  = \new_[8535]_  & \new_[8530]_ ;
  assign \new_[8540]_  = A199 & ~A166;
  assign \new_[8541]_  = A167 & \new_[8540]_ ;
  assign \new_[8545]_  = ~A202 & ~A201;
  assign \new_[8546]_  = A200 & \new_[8545]_ ;
  assign \new_[8547]_  = \new_[8546]_  & \new_[8541]_ ;
  assign \new_[8551]_  = A298 & A234;
  assign \new_[8552]_  = A232 & \new_[8551]_ ;
  assign \new_[8556]_  = A302 & ~A301;
  assign \new_[8557]_  = ~A299 & \new_[8556]_ ;
  assign \new_[8558]_  = \new_[8557]_  & \new_[8552]_ ;
  assign \new_[8562]_  = A199 & ~A166;
  assign \new_[8563]_  = A167 & \new_[8562]_ ;
  assign \new_[8567]_  = ~A202 & ~A201;
  assign \new_[8568]_  = A200 & \new_[8567]_ ;
  assign \new_[8569]_  = \new_[8568]_  & \new_[8563]_ ;
  assign \new_[8573]_  = ~A298 & A234;
  assign \new_[8574]_  = A232 & \new_[8573]_ ;
  assign \new_[8578]_  = A302 & ~A301;
  assign \new_[8579]_  = A299 & \new_[8578]_ ;
  assign \new_[8580]_  = \new_[8579]_  & \new_[8574]_ ;
  assign \new_[8584]_  = A199 & ~A166;
  assign \new_[8585]_  = A167 & \new_[8584]_ ;
  assign \new_[8589]_  = ~A202 & ~A201;
  assign \new_[8590]_  = A200 & \new_[8589]_ ;
  assign \new_[8591]_  = \new_[8590]_  & \new_[8585]_ ;
  assign \new_[8595]_  = ~A298 & A234;
  assign \new_[8596]_  = A232 & \new_[8595]_ ;
  assign \new_[8600]_  = ~A302 & A301;
  assign \new_[8601]_  = ~A299 & \new_[8600]_ ;
  assign \new_[8602]_  = \new_[8601]_  & \new_[8596]_ ;
  assign \new_[8606]_  = A199 & ~A166;
  assign \new_[8607]_  = A167 & \new_[8606]_ ;
  assign \new_[8611]_  = ~A202 & ~A201;
  assign \new_[8612]_  = A200 & \new_[8611]_ ;
  assign \new_[8613]_  = \new_[8612]_  & \new_[8607]_ ;
  assign \new_[8617]_  = A265 & A234;
  assign \new_[8618]_  = A232 & \new_[8617]_ ;
  assign \new_[8622]_  = ~A269 & A268;
  assign \new_[8623]_  = A266 & \new_[8622]_ ;
  assign \new_[8624]_  = \new_[8623]_  & \new_[8618]_ ;
  assign \new_[8628]_  = A199 & ~A166;
  assign \new_[8629]_  = A167 & \new_[8628]_ ;
  assign \new_[8633]_  = ~A202 & ~A201;
  assign \new_[8634]_  = A200 & \new_[8633]_ ;
  assign \new_[8635]_  = \new_[8634]_  & \new_[8629]_ ;
  assign \new_[8639]_  = ~A265 & A234;
  assign \new_[8640]_  = A232 & \new_[8639]_ ;
  assign \new_[8644]_  = A269 & ~A268;
  assign \new_[8645]_  = A266 & \new_[8644]_ ;
  assign \new_[8646]_  = \new_[8645]_  & \new_[8640]_ ;
  assign \new_[8650]_  = A199 & ~A166;
  assign \new_[8651]_  = A167 & \new_[8650]_ ;
  assign \new_[8655]_  = ~A202 & ~A201;
  assign \new_[8656]_  = A200 & \new_[8655]_ ;
  assign \new_[8657]_  = \new_[8656]_  & \new_[8651]_ ;
  assign \new_[8661]_  = A265 & A234;
  assign \new_[8662]_  = A232 & \new_[8661]_ ;
  assign \new_[8666]_  = A269 & ~A268;
  assign \new_[8667]_  = ~A266 & \new_[8666]_ ;
  assign \new_[8668]_  = \new_[8667]_  & \new_[8662]_ ;
  assign \new_[8672]_  = A199 & ~A166;
  assign \new_[8673]_  = A167 & \new_[8672]_ ;
  assign \new_[8677]_  = ~A202 & ~A201;
  assign \new_[8678]_  = A200 & \new_[8677]_ ;
  assign \new_[8679]_  = \new_[8678]_  & \new_[8673]_ ;
  assign \new_[8683]_  = ~A265 & A234;
  assign \new_[8684]_  = A232 & \new_[8683]_ ;
  assign \new_[8688]_  = ~A269 & A268;
  assign \new_[8689]_  = ~A266 & \new_[8688]_ ;
  assign \new_[8690]_  = \new_[8689]_  & \new_[8684]_ ;
  assign \new_[8694]_  = A199 & ~A166;
  assign \new_[8695]_  = A167 & \new_[8694]_ ;
  assign \new_[8699]_  = ~A202 & ~A201;
  assign \new_[8700]_  = A200 & \new_[8699]_ ;
  assign \new_[8701]_  = \new_[8700]_  & \new_[8695]_ ;
  assign \new_[8705]_  = A298 & A234;
  assign \new_[8706]_  = A233 & \new_[8705]_ ;
  assign \new_[8710]_  = ~A302 & A301;
  assign \new_[8711]_  = A299 & \new_[8710]_ ;
  assign \new_[8712]_  = \new_[8711]_  & \new_[8706]_ ;
  assign \new_[8716]_  = A199 & ~A166;
  assign \new_[8717]_  = A167 & \new_[8716]_ ;
  assign \new_[8721]_  = ~A202 & ~A201;
  assign \new_[8722]_  = A200 & \new_[8721]_ ;
  assign \new_[8723]_  = \new_[8722]_  & \new_[8717]_ ;
  assign \new_[8727]_  = A298 & A234;
  assign \new_[8728]_  = A233 & \new_[8727]_ ;
  assign \new_[8732]_  = A302 & ~A301;
  assign \new_[8733]_  = ~A299 & \new_[8732]_ ;
  assign \new_[8734]_  = \new_[8733]_  & \new_[8728]_ ;
  assign \new_[8738]_  = A199 & ~A166;
  assign \new_[8739]_  = A167 & \new_[8738]_ ;
  assign \new_[8743]_  = ~A202 & ~A201;
  assign \new_[8744]_  = A200 & \new_[8743]_ ;
  assign \new_[8745]_  = \new_[8744]_  & \new_[8739]_ ;
  assign \new_[8749]_  = ~A298 & A234;
  assign \new_[8750]_  = A233 & \new_[8749]_ ;
  assign \new_[8754]_  = A302 & ~A301;
  assign \new_[8755]_  = A299 & \new_[8754]_ ;
  assign \new_[8756]_  = \new_[8755]_  & \new_[8750]_ ;
  assign \new_[8760]_  = A199 & ~A166;
  assign \new_[8761]_  = A167 & \new_[8760]_ ;
  assign \new_[8765]_  = ~A202 & ~A201;
  assign \new_[8766]_  = A200 & \new_[8765]_ ;
  assign \new_[8767]_  = \new_[8766]_  & \new_[8761]_ ;
  assign \new_[8771]_  = ~A298 & A234;
  assign \new_[8772]_  = A233 & \new_[8771]_ ;
  assign \new_[8776]_  = ~A302 & A301;
  assign \new_[8777]_  = ~A299 & \new_[8776]_ ;
  assign \new_[8778]_  = \new_[8777]_  & \new_[8772]_ ;
  assign \new_[8782]_  = A199 & ~A166;
  assign \new_[8783]_  = A167 & \new_[8782]_ ;
  assign \new_[8787]_  = ~A202 & ~A201;
  assign \new_[8788]_  = A200 & \new_[8787]_ ;
  assign \new_[8789]_  = \new_[8788]_  & \new_[8783]_ ;
  assign \new_[8793]_  = A265 & A234;
  assign \new_[8794]_  = A233 & \new_[8793]_ ;
  assign \new_[8798]_  = ~A269 & A268;
  assign \new_[8799]_  = A266 & \new_[8798]_ ;
  assign \new_[8800]_  = \new_[8799]_  & \new_[8794]_ ;
  assign \new_[8804]_  = A199 & ~A166;
  assign \new_[8805]_  = A167 & \new_[8804]_ ;
  assign \new_[8809]_  = ~A202 & ~A201;
  assign \new_[8810]_  = A200 & \new_[8809]_ ;
  assign \new_[8811]_  = \new_[8810]_  & \new_[8805]_ ;
  assign \new_[8815]_  = ~A265 & A234;
  assign \new_[8816]_  = A233 & \new_[8815]_ ;
  assign \new_[8820]_  = A269 & ~A268;
  assign \new_[8821]_  = A266 & \new_[8820]_ ;
  assign \new_[8822]_  = \new_[8821]_  & \new_[8816]_ ;
  assign \new_[8826]_  = A199 & ~A166;
  assign \new_[8827]_  = A167 & \new_[8826]_ ;
  assign \new_[8831]_  = ~A202 & ~A201;
  assign \new_[8832]_  = A200 & \new_[8831]_ ;
  assign \new_[8833]_  = \new_[8832]_  & \new_[8827]_ ;
  assign \new_[8837]_  = A265 & A234;
  assign \new_[8838]_  = A233 & \new_[8837]_ ;
  assign \new_[8842]_  = A269 & ~A268;
  assign \new_[8843]_  = ~A266 & \new_[8842]_ ;
  assign \new_[8844]_  = \new_[8843]_  & \new_[8838]_ ;
  assign \new_[8848]_  = A199 & ~A166;
  assign \new_[8849]_  = A167 & \new_[8848]_ ;
  assign \new_[8853]_  = ~A202 & ~A201;
  assign \new_[8854]_  = A200 & \new_[8853]_ ;
  assign \new_[8855]_  = \new_[8854]_  & \new_[8849]_ ;
  assign \new_[8859]_  = ~A265 & A234;
  assign \new_[8860]_  = A233 & \new_[8859]_ ;
  assign \new_[8864]_  = ~A269 & A268;
  assign \new_[8865]_  = ~A266 & \new_[8864]_ ;
  assign \new_[8866]_  = \new_[8865]_  & \new_[8860]_ ;
  assign \new_[8870]_  = A199 & ~A166;
  assign \new_[8871]_  = A167 & \new_[8870]_ ;
  assign \new_[8875]_  = ~A202 & ~A201;
  assign \new_[8876]_  = A200 & \new_[8875]_ ;
  assign \new_[8877]_  = \new_[8876]_  & \new_[8871]_ ;
  assign \new_[8881]_  = A235 & A233;
  assign \new_[8882]_  = A232 & \new_[8881]_ ;
  assign \new_[8886]_  = A300 & A299;
  assign \new_[8887]_  = ~A236 & \new_[8886]_ ;
  assign \new_[8888]_  = \new_[8887]_  & \new_[8882]_ ;
  assign \new_[8892]_  = A199 & ~A166;
  assign \new_[8893]_  = A167 & \new_[8892]_ ;
  assign \new_[8897]_  = ~A202 & ~A201;
  assign \new_[8898]_  = A200 & \new_[8897]_ ;
  assign \new_[8899]_  = \new_[8898]_  & \new_[8893]_ ;
  assign \new_[8903]_  = A235 & A233;
  assign \new_[8904]_  = A232 & \new_[8903]_ ;
  assign \new_[8908]_  = A300 & A298;
  assign \new_[8909]_  = ~A236 & \new_[8908]_ ;
  assign \new_[8910]_  = \new_[8909]_  & \new_[8904]_ ;
  assign \new_[8914]_  = A199 & ~A166;
  assign \new_[8915]_  = A167 & \new_[8914]_ ;
  assign \new_[8919]_  = ~A202 & ~A201;
  assign \new_[8920]_  = A200 & \new_[8919]_ ;
  assign \new_[8921]_  = \new_[8920]_  & \new_[8915]_ ;
  assign \new_[8925]_  = A235 & A233;
  assign \new_[8926]_  = A232 & \new_[8925]_ ;
  assign \new_[8930]_  = A267 & A265;
  assign \new_[8931]_  = ~A236 & \new_[8930]_ ;
  assign \new_[8932]_  = \new_[8931]_  & \new_[8926]_ ;
  assign \new_[8936]_  = A199 & ~A166;
  assign \new_[8937]_  = A167 & \new_[8936]_ ;
  assign \new_[8941]_  = ~A202 & ~A201;
  assign \new_[8942]_  = A200 & \new_[8941]_ ;
  assign \new_[8943]_  = \new_[8942]_  & \new_[8937]_ ;
  assign \new_[8947]_  = A235 & A233;
  assign \new_[8948]_  = A232 & \new_[8947]_ ;
  assign \new_[8952]_  = A267 & A266;
  assign \new_[8953]_  = ~A236 & \new_[8952]_ ;
  assign \new_[8954]_  = \new_[8953]_  & \new_[8948]_ ;
  assign \new_[8958]_  = A199 & ~A166;
  assign \new_[8959]_  = A167 & \new_[8958]_ ;
  assign \new_[8963]_  = ~A202 & ~A201;
  assign \new_[8964]_  = A200 & \new_[8963]_ ;
  assign \new_[8965]_  = \new_[8964]_  & \new_[8959]_ ;
  assign \new_[8969]_  = ~A235 & A233;
  assign \new_[8970]_  = ~A232 & \new_[8969]_ ;
  assign \new_[8974]_  = A300 & A299;
  assign \new_[8975]_  = A236 & \new_[8974]_ ;
  assign \new_[8976]_  = \new_[8975]_  & \new_[8970]_ ;
  assign \new_[8980]_  = A199 & ~A166;
  assign \new_[8981]_  = A167 & \new_[8980]_ ;
  assign \new_[8985]_  = ~A202 & ~A201;
  assign \new_[8986]_  = A200 & \new_[8985]_ ;
  assign \new_[8987]_  = \new_[8986]_  & \new_[8981]_ ;
  assign \new_[8991]_  = ~A235 & A233;
  assign \new_[8992]_  = ~A232 & \new_[8991]_ ;
  assign \new_[8996]_  = A300 & A298;
  assign \new_[8997]_  = A236 & \new_[8996]_ ;
  assign \new_[8998]_  = \new_[8997]_  & \new_[8992]_ ;
  assign \new_[9002]_  = A199 & ~A166;
  assign \new_[9003]_  = A167 & \new_[9002]_ ;
  assign \new_[9007]_  = ~A202 & ~A201;
  assign \new_[9008]_  = A200 & \new_[9007]_ ;
  assign \new_[9009]_  = \new_[9008]_  & \new_[9003]_ ;
  assign \new_[9013]_  = ~A235 & A233;
  assign \new_[9014]_  = ~A232 & \new_[9013]_ ;
  assign \new_[9018]_  = A267 & A265;
  assign \new_[9019]_  = A236 & \new_[9018]_ ;
  assign \new_[9020]_  = \new_[9019]_  & \new_[9014]_ ;
  assign \new_[9024]_  = A199 & ~A166;
  assign \new_[9025]_  = A167 & \new_[9024]_ ;
  assign \new_[9029]_  = ~A202 & ~A201;
  assign \new_[9030]_  = A200 & \new_[9029]_ ;
  assign \new_[9031]_  = \new_[9030]_  & \new_[9025]_ ;
  assign \new_[9035]_  = ~A235 & A233;
  assign \new_[9036]_  = ~A232 & \new_[9035]_ ;
  assign \new_[9040]_  = A267 & A266;
  assign \new_[9041]_  = A236 & \new_[9040]_ ;
  assign \new_[9042]_  = \new_[9041]_  & \new_[9036]_ ;
  assign \new_[9046]_  = A199 & ~A166;
  assign \new_[9047]_  = A167 & \new_[9046]_ ;
  assign \new_[9051]_  = ~A202 & ~A201;
  assign \new_[9052]_  = A200 & \new_[9051]_ ;
  assign \new_[9053]_  = \new_[9052]_  & \new_[9047]_ ;
  assign \new_[9057]_  = ~A235 & ~A233;
  assign \new_[9058]_  = A232 & \new_[9057]_ ;
  assign \new_[9062]_  = A300 & A299;
  assign \new_[9063]_  = A236 & \new_[9062]_ ;
  assign \new_[9064]_  = \new_[9063]_  & \new_[9058]_ ;
  assign \new_[9068]_  = A199 & ~A166;
  assign \new_[9069]_  = A167 & \new_[9068]_ ;
  assign \new_[9073]_  = ~A202 & ~A201;
  assign \new_[9074]_  = A200 & \new_[9073]_ ;
  assign \new_[9075]_  = \new_[9074]_  & \new_[9069]_ ;
  assign \new_[9079]_  = ~A235 & ~A233;
  assign \new_[9080]_  = A232 & \new_[9079]_ ;
  assign \new_[9084]_  = A300 & A298;
  assign \new_[9085]_  = A236 & \new_[9084]_ ;
  assign \new_[9086]_  = \new_[9085]_  & \new_[9080]_ ;
  assign \new_[9090]_  = A199 & ~A166;
  assign \new_[9091]_  = A167 & \new_[9090]_ ;
  assign \new_[9095]_  = ~A202 & ~A201;
  assign \new_[9096]_  = A200 & \new_[9095]_ ;
  assign \new_[9097]_  = \new_[9096]_  & \new_[9091]_ ;
  assign \new_[9101]_  = ~A235 & ~A233;
  assign \new_[9102]_  = A232 & \new_[9101]_ ;
  assign \new_[9106]_  = A267 & A265;
  assign \new_[9107]_  = A236 & \new_[9106]_ ;
  assign \new_[9108]_  = \new_[9107]_  & \new_[9102]_ ;
  assign \new_[9112]_  = A199 & ~A166;
  assign \new_[9113]_  = A167 & \new_[9112]_ ;
  assign \new_[9117]_  = ~A202 & ~A201;
  assign \new_[9118]_  = A200 & \new_[9117]_ ;
  assign \new_[9119]_  = \new_[9118]_  & \new_[9113]_ ;
  assign \new_[9123]_  = ~A235 & ~A233;
  assign \new_[9124]_  = A232 & \new_[9123]_ ;
  assign \new_[9128]_  = A267 & A266;
  assign \new_[9129]_  = A236 & \new_[9128]_ ;
  assign \new_[9130]_  = \new_[9129]_  & \new_[9124]_ ;
  assign \new_[9134]_  = A199 & ~A166;
  assign \new_[9135]_  = A167 & \new_[9134]_ ;
  assign \new_[9139]_  = ~A202 & ~A201;
  assign \new_[9140]_  = A200 & \new_[9139]_ ;
  assign \new_[9141]_  = \new_[9140]_  & \new_[9135]_ ;
  assign \new_[9145]_  = A235 & ~A233;
  assign \new_[9146]_  = ~A232 & \new_[9145]_ ;
  assign \new_[9150]_  = A300 & A299;
  assign \new_[9151]_  = ~A236 & \new_[9150]_ ;
  assign \new_[9152]_  = \new_[9151]_  & \new_[9146]_ ;
  assign \new_[9156]_  = A199 & ~A166;
  assign \new_[9157]_  = A167 & \new_[9156]_ ;
  assign \new_[9161]_  = ~A202 & ~A201;
  assign \new_[9162]_  = A200 & \new_[9161]_ ;
  assign \new_[9163]_  = \new_[9162]_  & \new_[9157]_ ;
  assign \new_[9167]_  = A235 & ~A233;
  assign \new_[9168]_  = ~A232 & \new_[9167]_ ;
  assign \new_[9172]_  = A300 & A298;
  assign \new_[9173]_  = ~A236 & \new_[9172]_ ;
  assign \new_[9174]_  = \new_[9173]_  & \new_[9168]_ ;
  assign \new_[9178]_  = A199 & ~A166;
  assign \new_[9179]_  = A167 & \new_[9178]_ ;
  assign \new_[9183]_  = ~A202 & ~A201;
  assign \new_[9184]_  = A200 & \new_[9183]_ ;
  assign \new_[9185]_  = \new_[9184]_  & \new_[9179]_ ;
  assign \new_[9189]_  = A235 & ~A233;
  assign \new_[9190]_  = ~A232 & \new_[9189]_ ;
  assign \new_[9194]_  = A267 & A265;
  assign \new_[9195]_  = ~A236 & \new_[9194]_ ;
  assign \new_[9196]_  = \new_[9195]_  & \new_[9190]_ ;
  assign \new_[9200]_  = A199 & ~A166;
  assign \new_[9201]_  = A167 & \new_[9200]_ ;
  assign \new_[9205]_  = ~A202 & ~A201;
  assign \new_[9206]_  = A200 & \new_[9205]_ ;
  assign \new_[9207]_  = \new_[9206]_  & \new_[9201]_ ;
  assign \new_[9211]_  = A235 & ~A233;
  assign \new_[9212]_  = ~A232 & \new_[9211]_ ;
  assign \new_[9216]_  = A267 & A266;
  assign \new_[9217]_  = ~A236 & \new_[9216]_ ;
  assign \new_[9218]_  = \new_[9217]_  & \new_[9212]_ ;
  assign \new_[9222]_  = A199 & ~A166;
  assign \new_[9223]_  = A167 & \new_[9222]_ ;
  assign \new_[9227]_  = A203 & ~A201;
  assign \new_[9228]_  = A200 & \new_[9227]_ ;
  assign \new_[9229]_  = \new_[9228]_  & \new_[9223]_ ;
  assign \new_[9233]_  = A298 & A234;
  assign \new_[9234]_  = A232 & \new_[9233]_ ;
  assign \new_[9238]_  = ~A302 & A301;
  assign \new_[9239]_  = A299 & \new_[9238]_ ;
  assign \new_[9240]_  = \new_[9239]_  & \new_[9234]_ ;
  assign \new_[9244]_  = A199 & ~A166;
  assign \new_[9245]_  = A167 & \new_[9244]_ ;
  assign \new_[9249]_  = A203 & ~A201;
  assign \new_[9250]_  = A200 & \new_[9249]_ ;
  assign \new_[9251]_  = \new_[9250]_  & \new_[9245]_ ;
  assign \new_[9255]_  = A298 & A234;
  assign \new_[9256]_  = A232 & \new_[9255]_ ;
  assign \new_[9260]_  = A302 & ~A301;
  assign \new_[9261]_  = ~A299 & \new_[9260]_ ;
  assign \new_[9262]_  = \new_[9261]_  & \new_[9256]_ ;
  assign \new_[9266]_  = A199 & ~A166;
  assign \new_[9267]_  = A167 & \new_[9266]_ ;
  assign \new_[9271]_  = A203 & ~A201;
  assign \new_[9272]_  = A200 & \new_[9271]_ ;
  assign \new_[9273]_  = \new_[9272]_  & \new_[9267]_ ;
  assign \new_[9277]_  = ~A298 & A234;
  assign \new_[9278]_  = A232 & \new_[9277]_ ;
  assign \new_[9282]_  = A302 & ~A301;
  assign \new_[9283]_  = A299 & \new_[9282]_ ;
  assign \new_[9284]_  = \new_[9283]_  & \new_[9278]_ ;
  assign \new_[9288]_  = A199 & ~A166;
  assign \new_[9289]_  = A167 & \new_[9288]_ ;
  assign \new_[9293]_  = A203 & ~A201;
  assign \new_[9294]_  = A200 & \new_[9293]_ ;
  assign \new_[9295]_  = \new_[9294]_  & \new_[9289]_ ;
  assign \new_[9299]_  = ~A298 & A234;
  assign \new_[9300]_  = A232 & \new_[9299]_ ;
  assign \new_[9304]_  = ~A302 & A301;
  assign \new_[9305]_  = ~A299 & \new_[9304]_ ;
  assign \new_[9306]_  = \new_[9305]_  & \new_[9300]_ ;
  assign \new_[9310]_  = A199 & ~A166;
  assign \new_[9311]_  = A167 & \new_[9310]_ ;
  assign \new_[9315]_  = A203 & ~A201;
  assign \new_[9316]_  = A200 & \new_[9315]_ ;
  assign \new_[9317]_  = \new_[9316]_  & \new_[9311]_ ;
  assign \new_[9321]_  = A265 & A234;
  assign \new_[9322]_  = A232 & \new_[9321]_ ;
  assign \new_[9326]_  = ~A269 & A268;
  assign \new_[9327]_  = A266 & \new_[9326]_ ;
  assign \new_[9328]_  = \new_[9327]_  & \new_[9322]_ ;
  assign \new_[9332]_  = A199 & ~A166;
  assign \new_[9333]_  = A167 & \new_[9332]_ ;
  assign \new_[9337]_  = A203 & ~A201;
  assign \new_[9338]_  = A200 & \new_[9337]_ ;
  assign \new_[9339]_  = \new_[9338]_  & \new_[9333]_ ;
  assign \new_[9343]_  = ~A265 & A234;
  assign \new_[9344]_  = A232 & \new_[9343]_ ;
  assign \new_[9348]_  = A269 & ~A268;
  assign \new_[9349]_  = A266 & \new_[9348]_ ;
  assign \new_[9350]_  = \new_[9349]_  & \new_[9344]_ ;
  assign \new_[9354]_  = A199 & ~A166;
  assign \new_[9355]_  = A167 & \new_[9354]_ ;
  assign \new_[9359]_  = A203 & ~A201;
  assign \new_[9360]_  = A200 & \new_[9359]_ ;
  assign \new_[9361]_  = \new_[9360]_  & \new_[9355]_ ;
  assign \new_[9365]_  = A265 & A234;
  assign \new_[9366]_  = A232 & \new_[9365]_ ;
  assign \new_[9370]_  = A269 & ~A268;
  assign \new_[9371]_  = ~A266 & \new_[9370]_ ;
  assign \new_[9372]_  = \new_[9371]_  & \new_[9366]_ ;
  assign \new_[9376]_  = A199 & ~A166;
  assign \new_[9377]_  = A167 & \new_[9376]_ ;
  assign \new_[9381]_  = A203 & ~A201;
  assign \new_[9382]_  = A200 & \new_[9381]_ ;
  assign \new_[9383]_  = \new_[9382]_  & \new_[9377]_ ;
  assign \new_[9387]_  = ~A265 & A234;
  assign \new_[9388]_  = A232 & \new_[9387]_ ;
  assign \new_[9392]_  = ~A269 & A268;
  assign \new_[9393]_  = ~A266 & \new_[9392]_ ;
  assign \new_[9394]_  = \new_[9393]_  & \new_[9388]_ ;
  assign \new_[9398]_  = A199 & ~A166;
  assign \new_[9399]_  = A167 & \new_[9398]_ ;
  assign \new_[9403]_  = A203 & ~A201;
  assign \new_[9404]_  = A200 & \new_[9403]_ ;
  assign \new_[9405]_  = \new_[9404]_  & \new_[9399]_ ;
  assign \new_[9409]_  = A298 & A234;
  assign \new_[9410]_  = A233 & \new_[9409]_ ;
  assign \new_[9414]_  = ~A302 & A301;
  assign \new_[9415]_  = A299 & \new_[9414]_ ;
  assign \new_[9416]_  = \new_[9415]_  & \new_[9410]_ ;
  assign \new_[9420]_  = A199 & ~A166;
  assign \new_[9421]_  = A167 & \new_[9420]_ ;
  assign \new_[9425]_  = A203 & ~A201;
  assign \new_[9426]_  = A200 & \new_[9425]_ ;
  assign \new_[9427]_  = \new_[9426]_  & \new_[9421]_ ;
  assign \new_[9431]_  = A298 & A234;
  assign \new_[9432]_  = A233 & \new_[9431]_ ;
  assign \new_[9436]_  = A302 & ~A301;
  assign \new_[9437]_  = ~A299 & \new_[9436]_ ;
  assign \new_[9438]_  = \new_[9437]_  & \new_[9432]_ ;
  assign \new_[9442]_  = A199 & ~A166;
  assign \new_[9443]_  = A167 & \new_[9442]_ ;
  assign \new_[9447]_  = A203 & ~A201;
  assign \new_[9448]_  = A200 & \new_[9447]_ ;
  assign \new_[9449]_  = \new_[9448]_  & \new_[9443]_ ;
  assign \new_[9453]_  = ~A298 & A234;
  assign \new_[9454]_  = A233 & \new_[9453]_ ;
  assign \new_[9458]_  = A302 & ~A301;
  assign \new_[9459]_  = A299 & \new_[9458]_ ;
  assign \new_[9460]_  = \new_[9459]_  & \new_[9454]_ ;
  assign \new_[9464]_  = A199 & ~A166;
  assign \new_[9465]_  = A167 & \new_[9464]_ ;
  assign \new_[9469]_  = A203 & ~A201;
  assign \new_[9470]_  = A200 & \new_[9469]_ ;
  assign \new_[9471]_  = \new_[9470]_  & \new_[9465]_ ;
  assign \new_[9475]_  = ~A298 & A234;
  assign \new_[9476]_  = A233 & \new_[9475]_ ;
  assign \new_[9480]_  = ~A302 & A301;
  assign \new_[9481]_  = ~A299 & \new_[9480]_ ;
  assign \new_[9482]_  = \new_[9481]_  & \new_[9476]_ ;
  assign \new_[9486]_  = A199 & ~A166;
  assign \new_[9487]_  = A167 & \new_[9486]_ ;
  assign \new_[9491]_  = A203 & ~A201;
  assign \new_[9492]_  = A200 & \new_[9491]_ ;
  assign \new_[9493]_  = \new_[9492]_  & \new_[9487]_ ;
  assign \new_[9497]_  = A265 & A234;
  assign \new_[9498]_  = A233 & \new_[9497]_ ;
  assign \new_[9502]_  = ~A269 & A268;
  assign \new_[9503]_  = A266 & \new_[9502]_ ;
  assign \new_[9504]_  = \new_[9503]_  & \new_[9498]_ ;
  assign \new_[9508]_  = A199 & ~A166;
  assign \new_[9509]_  = A167 & \new_[9508]_ ;
  assign \new_[9513]_  = A203 & ~A201;
  assign \new_[9514]_  = A200 & \new_[9513]_ ;
  assign \new_[9515]_  = \new_[9514]_  & \new_[9509]_ ;
  assign \new_[9519]_  = ~A265 & A234;
  assign \new_[9520]_  = A233 & \new_[9519]_ ;
  assign \new_[9524]_  = A269 & ~A268;
  assign \new_[9525]_  = A266 & \new_[9524]_ ;
  assign \new_[9526]_  = \new_[9525]_  & \new_[9520]_ ;
  assign \new_[9530]_  = A199 & ~A166;
  assign \new_[9531]_  = A167 & \new_[9530]_ ;
  assign \new_[9535]_  = A203 & ~A201;
  assign \new_[9536]_  = A200 & \new_[9535]_ ;
  assign \new_[9537]_  = \new_[9536]_  & \new_[9531]_ ;
  assign \new_[9541]_  = A265 & A234;
  assign \new_[9542]_  = A233 & \new_[9541]_ ;
  assign \new_[9546]_  = A269 & ~A268;
  assign \new_[9547]_  = ~A266 & \new_[9546]_ ;
  assign \new_[9548]_  = \new_[9547]_  & \new_[9542]_ ;
  assign \new_[9552]_  = A199 & ~A166;
  assign \new_[9553]_  = A167 & \new_[9552]_ ;
  assign \new_[9557]_  = A203 & ~A201;
  assign \new_[9558]_  = A200 & \new_[9557]_ ;
  assign \new_[9559]_  = \new_[9558]_  & \new_[9553]_ ;
  assign \new_[9563]_  = ~A265 & A234;
  assign \new_[9564]_  = A233 & \new_[9563]_ ;
  assign \new_[9568]_  = ~A269 & A268;
  assign \new_[9569]_  = ~A266 & \new_[9568]_ ;
  assign \new_[9570]_  = \new_[9569]_  & \new_[9564]_ ;
  assign \new_[9574]_  = A199 & ~A166;
  assign \new_[9575]_  = A167 & \new_[9574]_ ;
  assign \new_[9579]_  = A203 & ~A201;
  assign \new_[9580]_  = A200 & \new_[9579]_ ;
  assign \new_[9581]_  = \new_[9580]_  & \new_[9575]_ ;
  assign \new_[9585]_  = A235 & A233;
  assign \new_[9586]_  = A232 & \new_[9585]_ ;
  assign \new_[9590]_  = A300 & A299;
  assign \new_[9591]_  = ~A236 & \new_[9590]_ ;
  assign \new_[9592]_  = \new_[9591]_  & \new_[9586]_ ;
  assign \new_[9596]_  = A199 & ~A166;
  assign \new_[9597]_  = A167 & \new_[9596]_ ;
  assign \new_[9601]_  = A203 & ~A201;
  assign \new_[9602]_  = A200 & \new_[9601]_ ;
  assign \new_[9603]_  = \new_[9602]_  & \new_[9597]_ ;
  assign \new_[9607]_  = A235 & A233;
  assign \new_[9608]_  = A232 & \new_[9607]_ ;
  assign \new_[9612]_  = A300 & A298;
  assign \new_[9613]_  = ~A236 & \new_[9612]_ ;
  assign \new_[9614]_  = \new_[9613]_  & \new_[9608]_ ;
  assign \new_[9618]_  = A199 & ~A166;
  assign \new_[9619]_  = A167 & \new_[9618]_ ;
  assign \new_[9623]_  = A203 & ~A201;
  assign \new_[9624]_  = A200 & \new_[9623]_ ;
  assign \new_[9625]_  = \new_[9624]_  & \new_[9619]_ ;
  assign \new_[9629]_  = A235 & A233;
  assign \new_[9630]_  = A232 & \new_[9629]_ ;
  assign \new_[9634]_  = A267 & A265;
  assign \new_[9635]_  = ~A236 & \new_[9634]_ ;
  assign \new_[9636]_  = \new_[9635]_  & \new_[9630]_ ;
  assign \new_[9640]_  = A199 & ~A166;
  assign \new_[9641]_  = A167 & \new_[9640]_ ;
  assign \new_[9645]_  = A203 & ~A201;
  assign \new_[9646]_  = A200 & \new_[9645]_ ;
  assign \new_[9647]_  = \new_[9646]_  & \new_[9641]_ ;
  assign \new_[9651]_  = A235 & A233;
  assign \new_[9652]_  = A232 & \new_[9651]_ ;
  assign \new_[9656]_  = A267 & A266;
  assign \new_[9657]_  = ~A236 & \new_[9656]_ ;
  assign \new_[9658]_  = \new_[9657]_  & \new_[9652]_ ;
  assign \new_[9662]_  = A199 & ~A166;
  assign \new_[9663]_  = A167 & \new_[9662]_ ;
  assign \new_[9667]_  = A203 & ~A201;
  assign \new_[9668]_  = A200 & \new_[9667]_ ;
  assign \new_[9669]_  = \new_[9668]_  & \new_[9663]_ ;
  assign \new_[9673]_  = ~A235 & A233;
  assign \new_[9674]_  = ~A232 & \new_[9673]_ ;
  assign \new_[9678]_  = A300 & A299;
  assign \new_[9679]_  = A236 & \new_[9678]_ ;
  assign \new_[9680]_  = \new_[9679]_  & \new_[9674]_ ;
  assign \new_[9684]_  = A199 & ~A166;
  assign \new_[9685]_  = A167 & \new_[9684]_ ;
  assign \new_[9689]_  = A203 & ~A201;
  assign \new_[9690]_  = A200 & \new_[9689]_ ;
  assign \new_[9691]_  = \new_[9690]_  & \new_[9685]_ ;
  assign \new_[9695]_  = ~A235 & A233;
  assign \new_[9696]_  = ~A232 & \new_[9695]_ ;
  assign \new_[9700]_  = A300 & A298;
  assign \new_[9701]_  = A236 & \new_[9700]_ ;
  assign \new_[9702]_  = \new_[9701]_  & \new_[9696]_ ;
  assign \new_[9706]_  = A199 & ~A166;
  assign \new_[9707]_  = A167 & \new_[9706]_ ;
  assign \new_[9711]_  = A203 & ~A201;
  assign \new_[9712]_  = A200 & \new_[9711]_ ;
  assign \new_[9713]_  = \new_[9712]_  & \new_[9707]_ ;
  assign \new_[9717]_  = ~A235 & A233;
  assign \new_[9718]_  = ~A232 & \new_[9717]_ ;
  assign \new_[9722]_  = A267 & A265;
  assign \new_[9723]_  = A236 & \new_[9722]_ ;
  assign \new_[9724]_  = \new_[9723]_  & \new_[9718]_ ;
  assign \new_[9728]_  = A199 & ~A166;
  assign \new_[9729]_  = A167 & \new_[9728]_ ;
  assign \new_[9733]_  = A203 & ~A201;
  assign \new_[9734]_  = A200 & \new_[9733]_ ;
  assign \new_[9735]_  = \new_[9734]_  & \new_[9729]_ ;
  assign \new_[9739]_  = ~A235 & A233;
  assign \new_[9740]_  = ~A232 & \new_[9739]_ ;
  assign \new_[9744]_  = A267 & A266;
  assign \new_[9745]_  = A236 & \new_[9744]_ ;
  assign \new_[9746]_  = \new_[9745]_  & \new_[9740]_ ;
  assign \new_[9750]_  = A199 & ~A166;
  assign \new_[9751]_  = A167 & \new_[9750]_ ;
  assign \new_[9755]_  = A203 & ~A201;
  assign \new_[9756]_  = A200 & \new_[9755]_ ;
  assign \new_[9757]_  = \new_[9756]_  & \new_[9751]_ ;
  assign \new_[9761]_  = ~A235 & ~A233;
  assign \new_[9762]_  = A232 & \new_[9761]_ ;
  assign \new_[9766]_  = A300 & A299;
  assign \new_[9767]_  = A236 & \new_[9766]_ ;
  assign \new_[9768]_  = \new_[9767]_  & \new_[9762]_ ;
  assign \new_[9772]_  = A199 & ~A166;
  assign \new_[9773]_  = A167 & \new_[9772]_ ;
  assign \new_[9777]_  = A203 & ~A201;
  assign \new_[9778]_  = A200 & \new_[9777]_ ;
  assign \new_[9779]_  = \new_[9778]_  & \new_[9773]_ ;
  assign \new_[9783]_  = ~A235 & ~A233;
  assign \new_[9784]_  = A232 & \new_[9783]_ ;
  assign \new_[9788]_  = A300 & A298;
  assign \new_[9789]_  = A236 & \new_[9788]_ ;
  assign \new_[9790]_  = \new_[9789]_  & \new_[9784]_ ;
  assign \new_[9794]_  = A199 & ~A166;
  assign \new_[9795]_  = A167 & \new_[9794]_ ;
  assign \new_[9799]_  = A203 & ~A201;
  assign \new_[9800]_  = A200 & \new_[9799]_ ;
  assign \new_[9801]_  = \new_[9800]_  & \new_[9795]_ ;
  assign \new_[9805]_  = ~A235 & ~A233;
  assign \new_[9806]_  = A232 & \new_[9805]_ ;
  assign \new_[9810]_  = A267 & A265;
  assign \new_[9811]_  = A236 & \new_[9810]_ ;
  assign \new_[9812]_  = \new_[9811]_  & \new_[9806]_ ;
  assign \new_[9816]_  = A199 & ~A166;
  assign \new_[9817]_  = A167 & \new_[9816]_ ;
  assign \new_[9821]_  = A203 & ~A201;
  assign \new_[9822]_  = A200 & \new_[9821]_ ;
  assign \new_[9823]_  = \new_[9822]_  & \new_[9817]_ ;
  assign \new_[9827]_  = ~A235 & ~A233;
  assign \new_[9828]_  = A232 & \new_[9827]_ ;
  assign \new_[9832]_  = A267 & A266;
  assign \new_[9833]_  = A236 & \new_[9832]_ ;
  assign \new_[9834]_  = \new_[9833]_  & \new_[9828]_ ;
  assign \new_[9838]_  = A199 & ~A166;
  assign \new_[9839]_  = A167 & \new_[9838]_ ;
  assign \new_[9843]_  = A203 & ~A201;
  assign \new_[9844]_  = A200 & \new_[9843]_ ;
  assign \new_[9845]_  = \new_[9844]_  & \new_[9839]_ ;
  assign \new_[9849]_  = A235 & ~A233;
  assign \new_[9850]_  = ~A232 & \new_[9849]_ ;
  assign \new_[9854]_  = A300 & A299;
  assign \new_[9855]_  = ~A236 & \new_[9854]_ ;
  assign \new_[9856]_  = \new_[9855]_  & \new_[9850]_ ;
  assign \new_[9860]_  = A199 & ~A166;
  assign \new_[9861]_  = A167 & \new_[9860]_ ;
  assign \new_[9865]_  = A203 & ~A201;
  assign \new_[9866]_  = A200 & \new_[9865]_ ;
  assign \new_[9867]_  = \new_[9866]_  & \new_[9861]_ ;
  assign \new_[9871]_  = A235 & ~A233;
  assign \new_[9872]_  = ~A232 & \new_[9871]_ ;
  assign \new_[9876]_  = A300 & A298;
  assign \new_[9877]_  = ~A236 & \new_[9876]_ ;
  assign \new_[9878]_  = \new_[9877]_  & \new_[9872]_ ;
  assign \new_[9882]_  = A199 & ~A166;
  assign \new_[9883]_  = A167 & \new_[9882]_ ;
  assign \new_[9887]_  = A203 & ~A201;
  assign \new_[9888]_  = A200 & \new_[9887]_ ;
  assign \new_[9889]_  = \new_[9888]_  & \new_[9883]_ ;
  assign \new_[9893]_  = A235 & ~A233;
  assign \new_[9894]_  = ~A232 & \new_[9893]_ ;
  assign \new_[9898]_  = A267 & A265;
  assign \new_[9899]_  = ~A236 & \new_[9898]_ ;
  assign \new_[9900]_  = \new_[9899]_  & \new_[9894]_ ;
  assign \new_[9904]_  = A199 & ~A166;
  assign \new_[9905]_  = A167 & \new_[9904]_ ;
  assign \new_[9909]_  = A203 & ~A201;
  assign \new_[9910]_  = A200 & \new_[9909]_ ;
  assign \new_[9911]_  = \new_[9910]_  & \new_[9905]_ ;
  assign \new_[9915]_  = A235 & ~A233;
  assign \new_[9916]_  = ~A232 & \new_[9915]_ ;
  assign \new_[9920]_  = A267 & A266;
  assign \new_[9921]_  = ~A236 & \new_[9920]_ ;
  assign \new_[9922]_  = \new_[9921]_  & \new_[9916]_ ;
  assign \new_[9926]_  = ~A199 & ~A166;
  assign \new_[9927]_  = A167 & \new_[9926]_ ;
  assign \new_[9931]_  = A202 & ~A201;
  assign \new_[9932]_  = A200 & \new_[9931]_ ;
  assign \new_[9933]_  = \new_[9932]_  & \new_[9927]_ ;
  assign \new_[9937]_  = A298 & A234;
  assign \new_[9938]_  = A232 & \new_[9937]_ ;
  assign \new_[9942]_  = ~A302 & A301;
  assign \new_[9943]_  = A299 & \new_[9942]_ ;
  assign \new_[9944]_  = \new_[9943]_  & \new_[9938]_ ;
  assign \new_[9948]_  = ~A199 & ~A166;
  assign \new_[9949]_  = A167 & \new_[9948]_ ;
  assign \new_[9953]_  = A202 & ~A201;
  assign \new_[9954]_  = A200 & \new_[9953]_ ;
  assign \new_[9955]_  = \new_[9954]_  & \new_[9949]_ ;
  assign \new_[9959]_  = A298 & A234;
  assign \new_[9960]_  = A232 & \new_[9959]_ ;
  assign \new_[9964]_  = A302 & ~A301;
  assign \new_[9965]_  = ~A299 & \new_[9964]_ ;
  assign \new_[9966]_  = \new_[9965]_  & \new_[9960]_ ;
  assign \new_[9970]_  = ~A199 & ~A166;
  assign \new_[9971]_  = A167 & \new_[9970]_ ;
  assign \new_[9975]_  = A202 & ~A201;
  assign \new_[9976]_  = A200 & \new_[9975]_ ;
  assign \new_[9977]_  = \new_[9976]_  & \new_[9971]_ ;
  assign \new_[9981]_  = ~A298 & A234;
  assign \new_[9982]_  = A232 & \new_[9981]_ ;
  assign \new_[9986]_  = A302 & ~A301;
  assign \new_[9987]_  = A299 & \new_[9986]_ ;
  assign \new_[9988]_  = \new_[9987]_  & \new_[9982]_ ;
  assign \new_[9992]_  = ~A199 & ~A166;
  assign \new_[9993]_  = A167 & \new_[9992]_ ;
  assign \new_[9997]_  = A202 & ~A201;
  assign \new_[9998]_  = A200 & \new_[9997]_ ;
  assign \new_[9999]_  = \new_[9998]_  & \new_[9993]_ ;
  assign \new_[10003]_  = ~A298 & A234;
  assign \new_[10004]_  = A232 & \new_[10003]_ ;
  assign \new_[10008]_  = ~A302 & A301;
  assign \new_[10009]_  = ~A299 & \new_[10008]_ ;
  assign \new_[10010]_  = \new_[10009]_  & \new_[10004]_ ;
  assign \new_[10014]_  = ~A199 & ~A166;
  assign \new_[10015]_  = A167 & \new_[10014]_ ;
  assign \new_[10019]_  = A202 & ~A201;
  assign \new_[10020]_  = A200 & \new_[10019]_ ;
  assign \new_[10021]_  = \new_[10020]_  & \new_[10015]_ ;
  assign \new_[10025]_  = A265 & A234;
  assign \new_[10026]_  = A232 & \new_[10025]_ ;
  assign \new_[10030]_  = ~A269 & A268;
  assign \new_[10031]_  = A266 & \new_[10030]_ ;
  assign \new_[10032]_  = \new_[10031]_  & \new_[10026]_ ;
  assign \new_[10036]_  = ~A199 & ~A166;
  assign \new_[10037]_  = A167 & \new_[10036]_ ;
  assign \new_[10041]_  = A202 & ~A201;
  assign \new_[10042]_  = A200 & \new_[10041]_ ;
  assign \new_[10043]_  = \new_[10042]_  & \new_[10037]_ ;
  assign \new_[10047]_  = ~A265 & A234;
  assign \new_[10048]_  = A232 & \new_[10047]_ ;
  assign \new_[10052]_  = A269 & ~A268;
  assign \new_[10053]_  = A266 & \new_[10052]_ ;
  assign \new_[10054]_  = \new_[10053]_  & \new_[10048]_ ;
  assign \new_[10058]_  = ~A199 & ~A166;
  assign \new_[10059]_  = A167 & \new_[10058]_ ;
  assign \new_[10063]_  = A202 & ~A201;
  assign \new_[10064]_  = A200 & \new_[10063]_ ;
  assign \new_[10065]_  = \new_[10064]_  & \new_[10059]_ ;
  assign \new_[10069]_  = A265 & A234;
  assign \new_[10070]_  = A232 & \new_[10069]_ ;
  assign \new_[10074]_  = A269 & ~A268;
  assign \new_[10075]_  = ~A266 & \new_[10074]_ ;
  assign \new_[10076]_  = \new_[10075]_  & \new_[10070]_ ;
  assign \new_[10080]_  = ~A199 & ~A166;
  assign \new_[10081]_  = A167 & \new_[10080]_ ;
  assign \new_[10085]_  = A202 & ~A201;
  assign \new_[10086]_  = A200 & \new_[10085]_ ;
  assign \new_[10087]_  = \new_[10086]_  & \new_[10081]_ ;
  assign \new_[10091]_  = ~A265 & A234;
  assign \new_[10092]_  = A232 & \new_[10091]_ ;
  assign \new_[10096]_  = ~A269 & A268;
  assign \new_[10097]_  = ~A266 & \new_[10096]_ ;
  assign \new_[10098]_  = \new_[10097]_  & \new_[10092]_ ;
  assign \new_[10102]_  = ~A199 & ~A166;
  assign \new_[10103]_  = A167 & \new_[10102]_ ;
  assign \new_[10107]_  = A202 & ~A201;
  assign \new_[10108]_  = A200 & \new_[10107]_ ;
  assign \new_[10109]_  = \new_[10108]_  & \new_[10103]_ ;
  assign \new_[10113]_  = A298 & A234;
  assign \new_[10114]_  = A233 & \new_[10113]_ ;
  assign \new_[10118]_  = ~A302 & A301;
  assign \new_[10119]_  = A299 & \new_[10118]_ ;
  assign \new_[10120]_  = \new_[10119]_  & \new_[10114]_ ;
  assign \new_[10124]_  = ~A199 & ~A166;
  assign \new_[10125]_  = A167 & \new_[10124]_ ;
  assign \new_[10129]_  = A202 & ~A201;
  assign \new_[10130]_  = A200 & \new_[10129]_ ;
  assign \new_[10131]_  = \new_[10130]_  & \new_[10125]_ ;
  assign \new_[10135]_  = A298 & A234;
  assign \new_[10136]_  = A233 & \new_[10135]_ ;
  assign \new_[10140]_  = A302 & ~A301;
  assign \new_[10141]_  = ~A299 & \new_[10140]_ ;
  assign \new_[10142]_  = \new_[10141]_  & \new_[10136]_ ;
  assign \new_[10146]_  = ~A199 & ~A166;
  assign \new_[10147]_  = A167 & \new_[10146]_ ;
  assign \new_[10151]_  = A202 & ~A201;
  assign \new_[10152]_  = A200 & \new_[10151]_ ;
  assign \new_[10153]_  = \new_[10152]_  & \new_[10147]_ ;
  assign \new_[10157]_  = ~A298 & A234;
  assign \new_[10158]_  = A233 & \new_[10157]_ ;
  assign \new_[10162]_  = A302 & ~A301;
  assign \new_[10163]_  = A299 & \new_[10162]_ ;
  assign \new_[10164]_  = \new_[10163]_  & \new_[10158]_ ;
  assign \new_[10168]_  = ~A199 & ~A166;
  assign \new_[10169]_  = A167 & \new_[10168]_ ;
  assign \new_[10173]_  = A202 & ~A201;
  assign \new_[10174]_  = A200 & \new_[10173]_ ;
  assign \new_[10175]_  = \new_[10174]_  & \new_[10169]_ ;
  assign \new_[10179]_  = ~A298 & A234;
  assign \new_[10180]_  = A233 & \new_[10179]_ ;
  assign \new_[10184]_  = ~A302 & A301;
  assign \new_[10185]_  = ~A299 & \new_[10184]_ ;
  assign \new_[10186]_  = \new_[10185]_  & \new_[10180]_ ;
  assign \new_[10190]_  = ~A199 & ~A166;
  assign \new_[10191]_  = A167 & \new_[10190]_ ;
  assign \new_[10195]_  = A202 & ~A201;
  assign \new_[10196]_  = A200 & \new_[10195]_ ;
  assign \new_[10197]_  = \new_[10196]_  & \new_[10191]_ ;
  assign \new_[10201]_  = A265 & A234;
  assign \new_[10202]_  = A233 & \new_[10201]_ ;
  assign \new_[10206]_  = ~A269 & A268;
  assign \new_[10207]_  = A266 & \new_[10206]_ ;
  assign \new_[10208]_  = \new_[10207]_  & \new_[10202]_ ;
  assign \new_[10212]_  = ~A199 & ~A166;
  assign \new_[10213]_  = A167 & \new_[10212]_ ;
  assign \new_[10217]_  = A202 & ~A201;
  assign \new_[10218]_  = A200 & \new_[10217]_ ;
  assign \new_[10219]_  = \new_[10218]_  & \new_[10213]_ ;
  assign \new_[10223]_  = ~A265 & A234;
  assign \new_[10224]_  = A233 & \new_[10223]_ ;
  assign \new_[10228]_  = A269 & ~A268;
  assign \new_[10229]_  = A266 & \new_[10228]_ ;
  assign \new_[10230]_  = \new_[10229]_  & \new_[10224]_ ;
  assign \new_[10234]_  = ~A199 & ~A166;
  assign \new_[10235]_  = A167 & \new_[10234]_ ;
  assign \new_[10239]_  = A202 & ~A201;
  assign \new_[10240]_  = A200 & \new_[10239]_ ;
  assign \new_[10241]_  = \new_[10240]_  & \new_[10235]_ ;
  assign \new_[10245]_  = A265 & A234;
  assign \new_[10246]_  = A233 & \new_[10245]_ ;
  assign \new_[10250]_  = A269 & ~A268;
  assign \new_[10251]_  = ~A266 & \new_[10250]_ ;
  assign \new_[10252]_  = \new_[10251]_  & \new_[10246]_ ;
  assign \new_[10256]_  = ~A199 & ~A166;
  assign \new_[10257]_  = A167 & \new_[10256]_ ;
  assign \new_[10261]_  = A202 & ~A201;
  assign \new_[10262]_  = A200 & \new_[10261]_ ;
  assign \new_[10263]_  = \new_[10262]_  & \new_[10257]_ ;
  assign \new_[10267]_  = ~A265 & A234;
  assign \new_[10268]_  = A233 & \new_[10267]_ ;
  assign \new_[10272]_  = ~A269 & A268;
  assign \new_[10273]_  = ~A266 & \new_[10272]_ ;
  assign \new_[10274]_  = \new_[10273]_  & \new_[10268]_ ;
  assign \new_[10278]_  = ~A199 & ~A166;
  assign \new_[10279]_  = A167 & \new_[10278]_ ;
  assign \new_[10283]_  = A202 & ~A201;
  assign \new_[10284]_  = A200 & \new_[10283]_ ;
  assign \new_[10285]_  = \new_[10284]_  & \new_[10279]_ ;
  assign \new_[10289]_  = A235 & A233;
  assign \new_[10290]_  = A232 & \new_[10289]_ ;
  assign \new_[10294]_  = A300 & A299;
  assign \new_[10295]_  = ~A236 & \new_[10294]_ ;
  assign \new_[10296]_  = \new_[10295]_  & \new_[10290]_ ;
  assign \new_[10300]_  = ~A199 & ~A166;
  assign \new_[10301]_  = A167 & \new_[10300]_ ;
  assign \new_[10305]_  = A202 & ~A201;
  assign \new_[10306]_  = A200 & \new_[10305]_ ;
  assign \new_[10307]_  = \new_[10306]_  & \new_[10301]_ ;
  assign \new_[10311]_  = A235 & A233;
  assign \new_[10312]_  = A232 & \new_[10311]_ ;
  assign \new_[10316]_  = A300 & A298;
  assign \new_[10317]_  = ~A236 & \new_[10316]_ ;
  assign \new_[10318]_  = \new_[10317]_  & \new_[10312]_ ;
  assign \new_[10322]_  = ~A199 & ~A166;
  assign \new_[10323]_  = A167 & \new_[10322]_ ;
  assign \new_[10327]_  = A202 & ~A201;
  assign \new_[10328]_  = A200 & \new_[10327]_ ;
  assign \new_[10329]_  = \new_[10328]_  & \new_[10323]_ ;
  assign \new_[10333]_  = A235 & A233;
  assign \new_[10334]_  = A232 & \new_[10333]_ ;
  assign \new_[10338]_  = A267 & A265;
  assign \new_[10339]_  = ~A236 & \new_[10338]_ ;
  assign \new_[10340]_  = \new_[10339]_  & \new_[10334]_ ;
  assign \new_[10344]_  = ~A199 & ~A166;
  assign \new_[10345]_  = A167 & \new_[10344]_ ;
  assign \new_[10349]_  = A202 & ~A201;
  assign \new_[10350]_  = A200 & \new_[10349]_ ;
  assign \new_[10351]_  = \new_[10350]_  & \new_[10345]_ ;
  assign \new_[10355]_  = A235 & A233;
  assign \new_[10356]_  = A232 & \new_[10355]_ ;
  assign \new_[10360]_  = A267 & A266;
  assign \new_[10361]_  = ~A236 & \new_[10360]_ ;
  assign \new_[10362]_  = \new_[10361]_  & \new_[10356]_ ;
  assign \new_[10366]_  = ~A199 & ~A166;
  assign \new_[10367]_  = A167 & \new_[10366]_ ;
  assign \new_[10371]_  = A202 & ~A201;
  assign \new_[10372]_  = A200 & \new_[10371]_ ;
  assign \new_[10373]_  = \new_[10372]_  & \new_[10367]_ ;
  assign \new_[10377]_  = ~A235 & A233;
  assign \new_[10378]_  = ~A232 & \new_[10377]_ ;
  assign \new_[10382]_  = A300 & A299;
  assign \new_[10383]_  = A236 & \new_[10382]_ ;
  assign \new_[10384]_  = \new_[10383]_  & \new_[10378]_ ;
  assign \new_[10388]_  = ~A199 & ~A166;
  assign \new_[10389]_  = A167 & \new_[10388]_ ;
  assign \new_[10393]_  = A202 & ~A201;
  assign \new_[10394]_  = A200 & \new_[10393]_ ;
  assign \new_[10395]_  = \new_[10394]_  & \new_[10389]_ ;
  assign \new_[10399]_  = ~A235 & A233;
  assign \new_[10400]_  = ~A232 & \new_[10399]_ ;
  assign \new_[10404]_  = A300 & A298;
  assign \new_[10405]_  = A236 & \new_[10404]_ ;
  assign \new_[10406]_  = \new_[10405]_  & \new_[10400]_ ;
  assign \new_[10410]_  = ~A199 & ~A166;
  assign \new_[10411]_  = A167 & \new_[10410]_ ;
  assign \new_[10415]_  = A202 & ~A201;
  assign \new_[10416]_  = A200 & \new_[10415]_ ;
  assign \new_[10417]_  = \new_[10416]_  & \new_[10411]_ ;
  assign \new_[10421]_  = ~A235 & A233;
  assign \new_[10422]_  = ~A232 & \new_[10421]_ ;
  assign \new_[10426]_  = A267 & A265;
  assign \new_[10427]_  = A236 & \new_[10426]_ ;
  assign \new_[10428]_  = \new_[10427]_  & \new_[10422]_ ;
  assign \new_[10432]_  = ~A199 & ~A166;
  assign \new_[10433]_  = A167 & \new_[10432]_ ;
  assign \new_[10437]_  = A202 & ~A201;
  assign \new_[10438]_  = A200 & \new_[10437]_ ;
  assign \new_[10439]_  = \new_[10438]_  & \new_[10433]_ ;
  assign \new_[10443]_  = ~A235 & A233;
  assign \new_[10444]_  = ~A232 & \new_[10443]_ ;
  assign \new_[10448]_  = A267 & A266;
  assign \new_[10449]_  = A236 & \new_[10448]_ ;
  assign \new_[10450]_  = \new_[10449]_  & \new_[10444]_ ;
  assign \new_[10454]_  = ~A199 & ~A166;
  assign \new_[10455]_  = A167 & \new_[10454]_ ;
  assign \new_[10459]_  = A202 & ~A201;
  assign \new_[10460]_  = A200 & \new_[10459]_ ;
  assign \new_[10461]_  = \new_[10460]_  & \new_[10455]_ ;
  assign \new_[10465]_  = ~A235 & ~A233;
  assign \new_[10466]_  = A232 & \new_[10465]_ ;
  assign \new_[10470]_  = A300 & A299;
  assign \new_[10471]_  = A236 & \new_[10470]_ ;
  assign \new_[10472]_  = \new_[10471]_  & \new_[10466]_ ;
  assign \new_[10476]_  = ~A199 & ~A166;
  assign \new_[10477]_  = A167 & \new_[10476]_ ;
  assign \new_[10481]_  = A202 & ~A201;
  assign \new_[10482]_  = A200 & \new_[10481]_ ;
  assign \new_[10483]_  = \new_[10482]_  & \new_[10477]_ ;
  assign \new_[10487]_  = ~A235 & ~A233;
  assign \new_[10488]_  = A232 & \new_[10487]_ ;
  assign \new_[10492]_  = A300 & A298;
  assign \new_[10493]_  = A236 & \new_[10492]_ ;
  assign \new_[10494]_  = \new_[10493]_  & \new_[10488]_ ;
  assign \new_[10498]_  = ~A199 & ~A166;
  assign \new_[10499]_  = A167 & \new_[10498]_ ;
  assign \new_[10503]_  = A202 & ~A201;
  assign \new_[10504]_  = A200 & \new_[10503]_ ;
  assign \new_[10505]_  = \new_[10504]_  & \new_[10499]_ ;
  assign \new_[10509]_  = ~A235 & ~A233;
  assign \new_[10510]_  = A232 & \new_[10509]_ ;
  assign \new_[10514]_  = A267 & A265;
  assign \new_[10515]_  = A236 & \new_[10514]_ ;
  assign \new_[10516]_  = \new_[10515]_  & \new_[10510]_ ;
  assign \new_[10520]_  = ~A199 & ~A166;
  assign \new_[10521]_  = A167 & \new_[10520]_ ;
  assign \new_[10525]_  = A202 & ~A201;
  assign \new_[10526]_  = A200 & \new_[10525]_ ;
  assign \new_[10527]_  = \new_[10526]_  & \new_[10521]_ ;
  assign \new_[10531]_  = ~A235 & ~A233;
  assign \new_[10532]_  = A232 & \new_[10531]_ ;
  assign \new_[10536]_  = A267 & A266;
  assign \new_[10537]_  = A236 & \new_[10536]_ ;
  assign \new_[10538]_  = \new_[10537]_  & \new_[10532]_ ;
  assign \new_[10542]_  = ~A199 & ~A166;
  assign \new_[10543]_  = A167 & \new_[10542]_ ;
  assign \new_[10547]_  = A202 & ~A201;
  assign \new_[10548]_  = A200 & \new_[10547]_ ;
  assign \new_[10549]_  = \new_[10548]_  & \new_[10543]_ ;
  assign \new_[10553]_  = A235 & ~A233;
  assign \new_[10554]_  = ~A232 & \new_[10553]_ ;
  assign \new_[10558]_  = A300 & A299;
  assign \new_[10559]_  = ~A236 & \new_[10558]_ ;
  assign \new_[10560]_  = \new_[10559]_  & \new_[10554]_ ;
  assign \new_[10564]_  = ~A199 & ~A166;
  assign \new_[10565]_  = A167 & \new_[10564]_ ;
  assign \new_[10569]_  = A202 & ~A201;
  assign \new_[10570]_  = A200 & \new_[10569]_ ;
  assign \new_[10571]_  = \new_[10570]_  & \new_[10565]_ ;
  assign \new_[10575]_  = A235 & ~A233;
  assign \new_[10576]_  = ~A232 & \new_[10575]_ ;
  assign \new_[10580]_  = A300 & A298;
  assign \new_[10581]_  = ~A236 & \new_[10580]_ ;
  assign \new_[10582]_  = \new_[10581]_  & \new_[10576]_ ;
  assign \new_[10586]_  = ~A199 & ~A166;
  assign \new_[10587]_  = A167 & \new_[10586]_ ;
  assign \new_[10591]_  = A202 & ~A201;
  assign \new_[10592]_  = A200 & \new_[10591]_ ;
  assign \new_[10593]_  = \new_[10592]_  & \new_[10587]_ ;
  assign \new_[10597]_  = A235 & ~A233;
  assign \new_[10598]_  = ~A232 & \new_[10597]_ ;
  assign \new_[10602]_  = A267 & A265;
  assign \new_[10603]_  = ~A236 & \new_[10602]_ ;
  assign \new_[10604]_  = \new_[10603]_  & \new_[10598]_ ;
  assign \new_[10608]_  = ~A199 & ~A166;
  assign \new_[10609]_  = A167 & \new_[10608]_ ;
  assign \new_[10613]_  = A202 & ~A201;
  assign \new_[10614]_  = A200 & \new_[10613]_ ;
  assign \new_[10615]_  = \new_[10614]_  & \new_[10609]_ ;
  assign \new_[10619]_  = A235 & ~A233;
  assign \new_[10620]_  = ~A232 & \new_[10619]_ ;
  assign \new_[10624]_  = A267 & A266;
  assign \new_[10625]_  = ~A236 & \new_[10624]_ ;
  assign \new_[10626]_  = \new_[10625]_  & \new_[10620]_ ;
  assign \new_[10630]_  = ~A199 & ~A166;
  assign \new_[10631]_  = A167 & \new_[10630]_ ;
  assign \new_[10635]_  = ~A203 & ~A201;
  assign \new_[10636]_  = A200 & \new_[10635]_ ;
  assign \new_[10637]_  = \new_[10636]_  & \new_[10631]_ ;
  assign \new_[10641]_  = A298 & A234;
  assign \new_[10642]_  = A232 & \new_[10641]_ ;
  assign \new_[10646]_  = ~A302 & A301;
  assign \new_[10647]_  = A299 & \new_[10646]_ ;
  assign \new_[10648]_  = \new_[10647]_  & \new_[10642]_ ;
  assign \new_[10652]_  = ~A199 & ~A166;
  assign \new_[10653]_  = A167 & \new_[10652]_ ;
  assign \new_[10657]_  = ~A203 & ~A201;
  assign \new_[10658]_  = A200 & \new_[10657]_ ;
  assign \new_[10659]_  = \new_[10658]_  & \new_[10653]_ ;
  assign \new_[10663]_  = A298 & A234;
  assign \new_[10664]_  = A232 & \new_[10663]_ ;
  assign \new_[10668]_  = A302 & ~A301;
  assign \new_[10669]_  = ~A299 & \new_[10668]_ ;
  assign \new_[10670]_  = \new_[10669]_  & \new_[10664]_ ;
  assign \new_[10674]_  = ~A199 & ~A166;
  assign \new_[10675]_  = A167 & \new_[10674]_ ;
  assign \new_[10679]_  = ~A203 & ~A201;
  assign \new_[10680]_  = A200 & \new_[10679]_ ;
  assign \new_[10681]_  = \new_[10680]_  & \new_[10675]_ ;
  assign \new_[10685]_  = ~A298 & A234;
  assign \new_[10686]_  = A232 & \new_[10685]_ ;
  assign \new_[10690]_  = A302 & ~A301;
  assign \new_[10691]_  = A299 & \new_[10690]_ ;
  assign \new_[10692]_  = \new_[10691]_  & \new_[10686]_ ;
  assign \new_[10696]_  = ~A199 & ~A166;
  assign \new_[10697]_  = A167 & \new_[10696]_ ;
  assign \new_[10701]_  = ~A203 & ~A201;
  assign \new_[10702]_  = A200 & \new_[10701]_ ;
  assign \new_[10703]_  = \new_[10702]_  & \new_[10697]_ ;
  assign \new_[10707]_  = ~A298 & A234;
  assign \new_[10708]_  = A232 & \new_[10707]_ ;
  assign \new_[10712]_  = ~A302 & A301;
  assign \new_[10713]_  = ~A299 & \new_[10712]_ ;
  assign \new_[10714]_  = \new_[10713]_  & \new_[10708]_ ;
  assign \new_[10718]_  = ~A199 & ~A166;
  assign \new_[10719]_  = A167 & \new_[10718]_ ;
  assign \new_[10723]_  = ~A203 & ~A201;
  assign \new_[10724]_  = A200 & \new_[10723]_ ;
  assign \new_[10725]_  = \new_[10724]_  & \new_[10719]_ ;
  assign \new_[10729]_  = A265 & A234;
  assign \new_[10730]_  = A232 & \new_[10729]_ ;
  assign \new_[10734]_  = ~A269 & A268;
  assign \new_[10735]_  = A266 & \new_[10734]_ ;
  assign \new_[10736]_  = \new_[10735]_  & \new_[10730]_ ;
  assign \new_[10740]_  = ~A199 & ~A166;
  assign \new_[10741]_  = A167 & \new_[10740]_ ;
  assign \new_[10745]_  = ~A203 & ~A201;
  assign \new_[10746]_  = A200 & \new_[10745]_ ;
  assign \new_[10747]_  = \new_[10746]_  & \new_[10741]_ ;
  assign \new_[10751]_  = ~A265 & A234;
  assign \new_[10752]_  = A232 & \new_[10751]_ ;
  assign \new_[10756]_  = A269 & ~A268;
  assign \new_[10757]_  = A266 & \new_[10756]_ ;
  assign \new_[10758]_  = \new_[10757]_  & \new_[10752]_ ;
  assign \new_[10762]_  = ~A199 & ~A166;
  assign \new_[10763]_  = A167 & \new_[10762]_ ;
  assign \new_[10767]_  = ~A203 & ~A201;
  assign \new_[10768]_  = A200 & \new_[10767]_ ;
  assign \new_[10769]_  = \new_[10768]_  & \new_[10763]_ ;
  assign \new_[10773]_  = A265 & A234;
  assign \new_[10774]_  = A232 & \new_[10773]_ ;
  assign \new_[10778]_  = A269 & ~A268;
  assign \new_[10779]_  = ~A266 & \new_[10778]_ ;
  assign \new_[10780]_  = \new_[10779]_  & \new_[10774]_ ;
  assign \new_[10784]_  = ~A199 & ~A166;
  assign \new_[10785]_  = A167 & \new_[10784]_ ;
  assign \new_[10789]_  = ~A203 & ~A201;
  assign \new_[10790]_  = A200 & \new_[10789]_ ;
  assign \new_[10791]_  = \new_[10790]_  & \new_[10785]_ ;
  assign \new_[10795]_  = ~A265 & A234;
  assign \new_[10796]_  = A232 & \new_[10795]_ ;
  assign \new_[10800]_  = ~A269 & A268;
  assign \new_[10801]_  = ~A266 & \new_[10800]_ ;
  assign \new_[10802]_  = \new_[10801]_  & \new_[10796]_ ;
  assign \new_[10806]_  = ~A199 & ~A166;
  assign \new_[10807]_  = A167 & \new_[10806]_ ;
  assign \new_[10811]_  = ~A203 & ~A201;
  assign \new_[10812]_  = A200 & \new_[10811]_ ;
  assign \new_[10813]_  = \new_[10812]_  & \new_[10807]_ ;
  assign \new_[10817]_  = A298 & A234;
  assign \new_[10818]_  = A233 & \new_[10817]_ ;
  assign \new_[10822]_  = ~A302 & A301;
  assign \new_[10823]_  = A299 & \new_[10822]_ ;
  assign \new_[10824]_  = \new_[10823]_  & \new_[10818]_ ;
  assign \new_[10828]_  = ~A199 & ~A166;
  assign \new_[10829]_  = A167 & \new_[10828]_ ;
  assign \new_[10833]_  = ~A203 & ~A201;
  assign \new_[10834]_  = A200 & \new_[10833]_ ;
  assign \new_[10835]_  = \new_[10834]_  & \new_[10829]_ ;
  assign \new_[10839]_  = A298 & A234;
  assign \new_[10840]_  = A233 & \new_[10839]_ ;
  assign \new_[10844]_  = A302 & ~A301;
  assign \new_[10845]_  = ~A299 & \new_[10844]_ ;
  assign \new_[10846]_  = \new_[10845]_  & \new_[10840]_ ;
  assign \new_[10850]_  = ~A199 & ~A166;
  assign \new_[10851]_  = A167 & \new_[10850]_ ;
  assign \new_[10855]_  = ~A203 & ~A201;
  assign \new_[10856]_  = A200 & \new_[10855]_ ;
  assign \new_[10857]_  = \new_[10856]_  & \new_[10851]_ ;
  assign \new_[10861]_  = ~A298 & A234;
  assign \new_[10862]_  = A233 & \new_[10861]_ ;
  assign \new_[10866]_  = A302 & ~A301;
  assign \new_[10867]_  = A299 & \new_[10866]_ ;
  assign \new_[10868]_  = \new_[10867]_  & \new_[10862]_ ;
  assign \new_[10872]_  = ~A199 & ~A166;
  assign \new_[10873]_  = A167 & \new_[10872]_ ;
  assign \new_[10877]_  = ~A203 & ~A201;
  assign \new_[10878]_  = A200 & \new_[10877]_ ;
  assign \new_[10879]_  = \new_[10878]_  & \new_[10873]_ ;
  assign \new_[10883]_  = ~A298 & A234;
  assign \new_[10884]_  = A233 & \new_[10883]_ ;
  assign \new_[10888]_  = ~A302 & A301;
  assign \new_[10889]_  = ~A299 & \new_[10888]_ ;
  assign \new_[10890]_  = \new_[10889]_  & \new_[10884]_ ;
  assign \new_[10894]_  = ~A199 & ~A166;
  assign \new_[10895]_  = A167 & \new_[10894]_ ;
  assign \new_[10899]_  = ~A203 & ~A201;
  assign \new_[10900]_  = A200 & \new_[10899]_ ;
  assign \new_[10901]_  = \new_[10900]_  & \new_[10895]_ ;
  assign \new_[10905]_  = A265 & A234;
  assign \new_[10906]_  = A233 & \new_[10905]_ ;
  assign \new_[10910]_  = ~A269 & A268;
  assign \new_[10911]_  = A266 & \new_[10910]_ ;
  assign \new_[10912]_  = \new_[10911]_  & \new_[10906]_ ;
  assign \new_[10916]_  = ~A199 & ~A166;
  assign \new_[10917]_  = A167 & \new_[10916]_ ;
  assign \new_[10921]_  = ~A203 & ~A201;
  assign \new_[10922]_  = A200 & \new_[10921]_ ;
  assign \new_[10923]_  = \new_[10922]_  & \new_[10917]_ ;
  assign \new_[10927]_  = ~A265 & A234;
  assign \new_[10928]_  = A233 & \new_[10927]_ ;
  assign \new_[10932]_  = A269 & ~A268;
  assign \new_[10933]_  = A266 & \new_[10932]_ ;
  assign \new_[10934]_  = \new_[10933]_  & \new_[10928]_ ;
  assign \new_[10938]_  = ~A199 & ~A166;
  assign \new_[10939]_  = A167 & \new_[10938]_ ;
  assign \new_[10943]_  = ~A203 & ~A201;
  assign \new_[10944]_  = A200 & \new_[10943]_ ;
  assign \new_[10945]_  = \new_[10944]_  & \new_[10939]_ ;
  assign \new_[10949]_  = A265 & A234;
  assign \new_[10950]_  = A233 & \new_[10949]_ ;
  assign \new_[10954]_  = A269 & ~A268;
  assign \new_[10955]_  = ~A266 & \new_[10954]_ ;
  assign \new_[10956]_  = \new_[10955]_  & \new_[10950]_ ;
  assign \new_[10960]_  = ~A199 & ~A166;
  assign \new_[10961]_  = A167 & \new_[10960]_ ;
  assign \new_[10965]_  = ~A203 & ~A201;
  assign \new_[10966]_  = A200 & \new_[10965]_ ;
  assign \new_[10967]_  = \new_[10966]_  & \new_[10961]_ ;
  assign \new_[10971]_  = ~A265 & A234;
  assign \new_[10972]_  = A233 & \new_[10971]_ ;
  assign \new_[10976]_  = ~A269 & A268;
  assign \new_[10977]_  = ~A266 & \new_[10976]_ ;
  assign \new_[10978]_  = \new_[10977]_  & \new_[10972]_ ;
  assign \new_[10982]_  = ~A199 & ~A166;
  assign \new_[10983]_  = A167 & \new_[10982]_ ;
  assign \new_[10987]_  = ~A203 & ~A201;
  assign \new_[10988]_  = A200 & \new_[10987]_ ;
  assign \new_[10989]_  = \new_[10988]_  & \new_[10983]_ ;
  assign \new_[10993]_  = A235 & A233;
  assign \new_[10994]_  = A232 & \new_[10993]_ ;
  assign \new_[10998]_  = A300 & A299;
  assign \new_[10999]_  = ~A236 & \new_[10998]_ ;
  assign \new_[11000]_  = \new_[10999]_  & \new_[10994]_ ;
  assign \new_[11004]_  = ~A199 & ~A166;
  assign \new_[11005]_  = A167 & \new_[11004]_ ;
  assign \new_[11009]_  = ~A203 & ~A201;
  assign \new_[11010]_  = A200 & \new_[11009]_ ;
  assign \new_[11011]_  = \new_[11010]_  & \new_[11005]_ ;
  assign \new_[11015]_  = A235 & A233;
  assign \new_[11016]_  = A232 & \new_[11015]_ ;
  assign \new_[11020]_  = A300 & A298;
  assign \new_[11021]_  = ~A236 & \new_[11020]_ ;
  assign \new_[11022]_  = \new_[11021]_  & \new_[11016]_ ;
  assign \new_[11026]_  = ~A199 & ~A166;
  assign \new_[11027]_  = A167 & \new_[11026]_ ;
  assign \new_[11031]_  = ~A203 & ~A201;
  assign \new_[11032]_  = A200 & \new_[11031]_ ;
  assign \new_[11033]_  = \new_[11032]_  & \new_[11027]_ ;
  assign \new_[11037]_  = A235 & A233;
  assign \new_[11038]_  = A232 & \new_[11037]_ ;
  assign \new_[11042]_  = A267 & A265;
  assign \new_[11043]_  = ~A236 & \new_[11042]_ ;
  assign \new_[11044]_  = \new_[11043]_  & \new_[11038]_ ;
  assign \new_[11048]_  = ~A199 & ~A166;
  assign \new_[11049]_  = A167 & \new_[11048]_ ;
  assign \new_[11053]_  = ~A203 & ~A201;
  assign \new_[11054]_  = A200 & \new_[11053]_ ;
  assign \new_[11055]_  = \new_[11054]_  & \new_[11049]_ ;
  assign \new_[11059]_  = A235 & A233;
  assign \new_[11060]_  = A232 & \new_[11059]_ ;
  assign \new_[11064]_  = A267 & A266;
  assign \new_[11065]_  = ~A236 & \new_[11064]_ ;
  assign \new_[11066]_  = \new_[11065]_  & \new_[11060]_ ;
  assign \new_[11070]_  = ~A199 & ~A166;
  assign \new_[11071]_  = A167 & \new_[11070]_ ;
  assign \new_[11075]_  = ~A203 & ~A201;
  assign \new_[11076]_  = A200 & \new_[11075]_ ;
  assign \new_[11077]_  = \new_[11076]_  & \new_[11071]_ ;
  assign \new_[11081]_  = ~A235 & A233;
  assign \new_[11082]_  = ~A232 & \new_[11081]_ ;
  assign \new_[11086]_  = A300 & A299;
  assign \new_[11087]_  = A236 & \new_[11086]_ ;
  assign \new_[11088]_  = \new_[11087]_  & \new_[11082]_ ;
  assign \new_[11092]_  = ~A199 & ~A166;
  assign \new_[11093]_  = A167 & \new_[11092]_ ;
  assign \new_[11097]_  = ~A203 & ~A201;
  assign \new_[11098]_  = A200 & \new_[11097]_ ;
  assign \new_[11099]_  = \new_[11098]_  & \new_[11093]_ ;
  assign \new_[11103]_  = ~A235 & A233;
  assign \new_[11104]_  = ~A232 & \new_[11103]_ ;
  assign \new_[11108]_  = A300 & A298;
  assign \new_[11109]_  = A236 & \new_[11108]_ ;
  assign \new_[11110]_  = \new_[11109]_  & \new_[11104]_ ;
  assign \new_[11114]_  = ~A199 & ~A166;
  assign \new_[11115]_  = A167 & \new_[11114]_ ;
  assign \new_[11119]_  = ~A203 & ~A201;
  assign \new_[11120]_  = A200 & \new_[11119]_ ;
  assign \new_[11121]_  = \new_[11120]_  & \new_[11115]_ ;
  assign \new_[11125]_  = ~A235 & A233;
  assign \new_[11126]_  = ~A232 & \new_[11125]_ ;
  assign \new_[11130]_  = A267 & A265;
  assign \new_[11131]_  = A236 & \new_[11130]_ ;
  assign \new_[11132]_  = \new_[11131]_  & \new_[11126]_ ;
  assign \new_[11136]_  = ~A199 & ~A166;
  assign \new_[11137]_  = A167 & \new_[11136]_ ;
  assign \new_[11141]_  = ~A203 & ~A201;
  assign \new_[11142]_  = A200 & \new_[11141]_ ;
  assign \new_[11143]_  = \new_[11142]_  & \new_[11137]_ ;
  assign \new_[11147]_  = ~A235 & A233;
  assign \new_[11148]_  = ~A232 & \new_[11147]_ ;
  assign \new_[11152]_  = A267 & A266;
  assign \new_[11153]_  = A236 & \new_[11152]_ ;
  assign \new_[11154]_  = \new_[11153]_  & \new_[11148]_ ;
  assign \new_[11158]_  = ~A199 & ~A166;
  assign \new_[11159]_  = A167 & \new_[11158]_ ;
  assign \new_[11163]_  = ~A203 & ~A201;
  assign \new_[11164]_  = A200 & \new_[11163]_ ;
  assign \new_[11165]_  = \new_[11164]_  & \new_[11159]_ ;
  assign \new_[11169]_  = ~A235 & ~A233;
  assign \new_[11170]_  = A232 & \new_[11169]_ ;
  assign \new_[11174]_  = A300 & A299;
  assign \new_[11175]_  = A236 & \new_[11174]_ ;
  assign \new_[11176]_  = \new_[11175]_  & \new_[11170]_ ;
  assign \new_[11180]_  = ~A199 & ~A166;
  assign \new_[11181]_  = A167 & \new_[11180]_ ;
  assign \new_[11185]_  = ~A203 & ~A201;
  assign \new_[11186]_  = A200 & \new_[11185]_ ;
  assign \new_[11187]_  = \new_[11186]_  & \new_[11181]_ ;
  assign \new_[11191]_  = ~A235 & ~A233;
  assign \new_[11192]_  = A232 & \new_[11191]_ ;
  assign \new_[11196]_  = A300 & A298;
  assign \new_[11197]_  = A236 & \new_[11196]_ ;
  assign \new_[11198]_  = \new_[11197]_  & \new_[11192]_ ;
  assign \new_[11202]_  = ~A199 & ~A166;
  assign \new_[11203]_  = A167 & \new_[11202]_ ;
  assign \new_[11207]_  = ~A203 & ~A201;
  assign \new_[11208]_  = A200 & \new_[11207]_ ;
  assign \new_[11209]_  = \new_[11208]_  & \new_[11203]_ ;
  assign \new_[11213]_  = ~A235 & ~A233;
  assign \new_[11214]_  = A232 & \new_[11213]_ ;
  assign \new_[11218]_  = A267 & A265;
  assign \new_[11219]_  = A236 & \new_[11218]_ ;
  assign \new_[11220]_  = \new_[11219]_  & \new_[11214]_ ;
  assign \new_[11224]_  = ~A199 & ~A166;
  assign \new_[11225]_  = A167 & \new_[11224]_ ;
  assign \new_[11229]_  = ~A203 & ~A201;
  assign \new_[11230]_  = A200 & \new_[11229]_ ;
  assign \new_[11231]_  = \new_[11230]_  & \new_[11225]_ ;
  assign \new_[11235]_  = ~A235 & ~A233;
  assign \new_[11236]_  = A232 & \new_[11235]_ ;
  assign \new_[11240]_  = A267 & A266;
  assign \new_[11241]_  = A236 & \new_[11240]_ ;
  assign \new_[11242]_  = \new_[11241]_  & \new_[11236]_ ;
  assign \new_[11246]_  = ~A199 & ~A166;
  assign \new_[11247]_  = A167 & \new_[11246]_ ;
  assign \new_[11251]_  = ~A203 & ~A201;
  assign \new_[11252]_  = A200 & \new_[11251]_ ;
  assign \new_[11253]_  = \new_[11252]_  & \new_[11247]_ ;
  assign \new_[11257]_  = A235 & ~A233;
  assign \new_[11258]_  = ~A232 & \new_[11257]_ ;
  assign \new_[11262]_  = A300 & A299;
  assign \new_[11263]_  = ~A236 & \new_[11262]_ ;
  assign \new_[11264]_  = \new_[11263]_  & \new_[11258]_ ;
  assign \new_[11268]_  = ~A199 & ~A166;
  assign \new_[11269]_  = A167 & \new_[11268]_ ;
  assign \new_[11273]_  = ~A203 & ~A201;
  assign \new_[11274]_  = A200 & \new_[11273]_ ;
  assign \new_[11275]_  = \new_[11274]_  & \new_[11269]_ ;
  assign \new_[11279]_  = A235 & ~A233;
  assign \new_[11280]_  = ~A232 & \new_[11279]_ ;
  assign \new_[11284]_  = A300 & A298;
  assign \new_[11285]_  = ~A236 & \new_[11284]_ ;
  assign \new_[11286]_  = \new_[11285]_  & \new_[11280]_ ;
  assign \new_[11290]_  = ~A199 & ~A166;
  assign \new_[11291]_  = A167 & \new_[11290]_ ;
  assign \new_[11295]_  = ~A203 & ~A201;
  assign \new_[11296]_  = A200 & \new_[11295]_ ;
  assign \new_[11297]_  = \new_[11296]_  & \new_[11291]_ ;
  assign \new_[11301]_  = A235 & ~A233;
  assign \new_[11302]_  = ~A232 & \new_[11301]_ ;
  assign \new_[11306]_  = A267 & A265;
  assign \new_[11307]_  = ~A236 & \new_[11306]_ ;
  assign \new_[11308]_  = \new_[11307]_  & \new_[11302]_ ;
  assign \new_[11312]_  = ~A199 & ~A166;
  assign \new_[11313]_  = A167 & \new_[11312]_ ;
  assign \new_[11317]_  = ~A203 & ~A201;
  assign \new_[11318]_  = A200 & \new_[11317]_ ;
  assign \new_[11319]_  = \new_[11318]_  & \new_[11313]_ ;
  assign \new_[11323]_  = A235 & ~A233;
  assign \new_[11324]_  = ~A232 & \new_[11323]_ ;
  assign \new_[11328]_  = A267 & A266;
  assign \new_[11329]_  = ~A236 & \new_[11328]_ ;
  assign \new_[11330]_  = \new_[11329]_  & \new_[11324]_ ;
  assign \new_[11334]_  = A199 & ~A166;
  assign \new_[11335]_  = A167 & \new_[11334]_ ;
  assign \new_[11339]_  = A202 & ~A201;
  assign \new_[11340]_  = ~A200 & \new_[11339]_ ;
  assign \new_[11341]_  = \new_[11340]_  & \new_[11335]_ ;
  assign \new_[11345]_  = A298 & A234;
  assign \new_[11346]_  = A232 & \new_[11345]_ ;
  assign \new_[11350]_  = ~A302 & A301;
  assign \new_[11351]_  = A299 & \new_[11350]_ ;
  assign \new_[11352]_  = \new_[11351]_  & \new_[11346]_ ;
  assign \new_[11356]_  = A199 & ~A166;
  assign \new_[11357]_  = A167 & \new_[11356]_ ;
  assign \new_[11361]_  = A202 & ~A201;
  assign \new_[11362]_  = ~A200 & \new_[11361]_ ;
  assign \new_[11363]_  = \new_[11362]_  & \new_[11357]_ ;
  assign \new_[11367]_  = A298 & A234;
  assign \new_[11368]_  = A232 & \new_[11367]_ ;
  assign \new_[11372]_  = A302 & ~A301;
  assign \new_[11373]_  = ~A299 & \new_[11372]_ ;
  assign \new_[11374]_  = \new_[11373]_  & \new_[11368]_ ;
  assign \new_[11378]_  = A199 & ~A166;
  assign \new_[11379]_  = A167 & \new_[11378]_ ;
  assign \new_[11383]_  = A202 & ~A201;
  assign \new_[11384]_  = ~A200 & \new_[11383]_ ;
  assign \new_[11385]_  = \new_[11384]_  & \new_[11379]_ ;
  assign \new_[11389]_  = ~A298 & A234;
  assign \new_[11390]_  = A232 & \new_[11389]_ ;
  assign \new_[11394]_  = A302 & ~A301;
  assign \new_[11395]_  = A299 & \new_[11394]_ ;
  assign \new_[11396]_  = \new_[11395]_  & \new_[11390]_ ;
  assign \new_[11400]_  = A199 & ~A166;
  assign \new_[11401]_  = A167 & \new_[11400]_ ;
  assign \new_[11405]_  = A202 & ~A201;
  assign \new_[11406]_  = ~A200 & \new_[11405]_ ;
  assign \new_[11407]_  = \new_[11406]_  & \new_[11401]_ ;
  assign \new_[11411]_  = ~A298 & A234;
  assign \new_[11412]_  = A232 & \new_[11411]_ ;
  assign \new_[11416]_  = ~A302 & A301;
  assign \new_[11417]_  = ~A299 & \new_[11416]_ ;
  assign \new_[11418]_  = \new_[11417]_  & \new_[11412]_ ;
  assign \new_[11422]_  = A199 & ~A166;
  assign \new_[11423]_  = A167 & \new_[11422]_ ;
  assign \new_[11427]_  = A202 & ~A201;
  assign \new_[11428]_  = ~A200 & \new_[11427]_ ;
  assign \new_[11429]_  = \new_[11428]_  & \new_[11423]_ ;
  assign \new_[11433]_  = A265 & A234;
  assign \new_[11434]_  = A232 & \new_[11433]_ ;
  assign \new_[11438]_  = ~A269 & A268;
  assign \new_[11439]_  = A266 & \new_[11438]_ ;
  assign \new_[11440]_  = \new_[11439]_  & \new_[11434]_ ;
  assign \new_[11444]_  = A199 & ~A166;
  assign \new_[11445]_  = A167 & \new_[11444]_ ;
  assign \new_[11449]_  = A202 & ~A201;
  assign \new_[11450]_  = ~A200 & \new_[11449]_ ;
  assign \new_[11451]_  = \new_[11450]_  & \new_[11445]_ ;
  assign \new_[11455]_  = ~A265 & A234;
  assign \new_[11456]_  = A232 & \new_[11455]_ ;
  assign \new_[11460]_  = A269 & ~A268;
  assign \new_[11461]_  = A266 & \new_[11460]_ ;
  assign \new_[11462]_  = \new_[11461]_  & \new_[11456]_ ;
  assign \new_[11466]_  = A199 & ~A166;
  assign \new_[11467]_  = A167 & \new_[11466]_ ;
  assign \new_[11471]_  = A202 & ~A201;
  assign \new_[11472]_  = ~A200 & \new_[11471]_ ;
  assign \new_[11473]_  = \new_[11472]_  & \new_[11467]_ ;
  assign \new_[11477]_  = A265 & A234;
  assign \new_[11478]_  = A232 & \new_[11477]_ ;
  assign \new_[11482]_  = A269 & ~A268;
  assign \new_[11483]_  = ~A266 & \new_[11482]_ ;
  assign \new_[11484]_  = \new_[11483]_  & \new_[11478]_ ;
  assign \new_[11488]_  = A199 & ~A166;
  assign \new_[11489]_  = A167 & \new_[11488]_ ;
  assign \new_[11493]_  = A202 & ~A201;
  assign \new_[11494]_  = ~A200 & \new_[11493]_ ;
  assign \new_[11495]_  = \new_[11494]_  & \new_[11489]_ ;
  assign \new_[11499]_  = ~A265 & A234;
  assign \new_[11500]_  = A232 & \new_[11499]_ ;
  assign \new_[11504]_  = ~A269 & A268;
  assign \new_[11505]_  = ~A266 & \new_[11504]_ ;
  assign \new_[11506]_  = \new_[11505]_  & \new_[11500]_ ;
  assign \new_[11510]_  = A199 & ~A166;
  assign \new_[11511]_  = A167 & \new_[11510]_ ;
  assign \new_[11515]_  = A202 & ~A201;
  assign \new_[11516]_  = ~A200 & \new_[11515]_ ;
  assign \new_[11517]_  = \new_[11516]_  & \new_[11511]_ ;
  assign \new_[11521]_  = A298 & A234;
  assign \new_[11522]_  = A233 & \new_[11521]_ ;
  assign \new_[11526]_  = ~A302 & A301;
  assign \new_[11527]_  = A299 & \new_[11526]_ ;
  assign \new_[11528]_  = \new_[11527]_  & \new_[11522]_ ;
  assign \new_[11532]_  = A199 & ~A166;
  assign \new_[11533]_  = A167 & \new_[11532]_ ;
  assign \new_[11537]_  = A202 & ~A201;
  assign \new_[11538]_  = ~A200 & \new_[11537]_ ;
  assign \new_[11539]_  = \new_[11538]_  & \new_[11533]_ ;
  assign \new_[11543]_  = A298 & A234;
  assign \new_[11544]_  = A233 & \new_[11543]_ ;
  assign \new_[11548]_  = A302 & ~A301;
  assign \new_[11549]_  = ~A299 & \new_[11548]_ ;
  assign \new_[11550]_  = \new_[11549]_  & \new_[11544]_ ;
  assign \new_[11554]_  = A199 & ~A166;
  assign \new_[11555]_  = A167 & \new_[11554]_ ;
  assign \new_[11559]_  = A202 & ~A201;
  assign \new_[11560]_  = ~A200 & \new_[11559]_ ;
  assign \new_[11561]_  = \new_[11560]_  & \new_[11555]_ ;
  assign \new_[11565]_  = ~A298 & A234;
  assign \new_[11566]_  = A233 & \new_[11565]_ ;
  assign \new_[11570]_  = A302 & ~A301;
  assign \new_[11571]_  = A299 & \new_[11570]_ ;
  assign \new_[11572]_  = \new_[11571]_  & \new_[11566]_ ;
  assign \new_[11576]_  = A199 & ~A166;
  assign \new_[11577]_  = A167 & \new_[11576]_ ;
  assign \new_[11581]_  = A202 & ~A201;
  assign \new_[11582]_  = ~A200 & \new_[11581]_ ;
  assign \new_[11583]_  = \new_[11582]_  & \new_[11577]_ ;
  assign \new_[11587]_  = ~A298 & A234;
  assign \new_[11588]_  = A233 & \new_[11587]_ ;
  assign \new_[11592]_  = ~A302 & A301;
  assign \new_[11593]_  = ~A299 & \new_[11592]_ ;
  assign \new_[11594]_  = \new_[11593]_  & \new_[11588]_ ;
  assign \new_[11598]_  = A199 & ~A166;
  assign \new_[11599]_  = A167 & \new_[11598]_ ;
  assign \new_[11603]_  = A202 & ~A201;
  assign \new_[11604]_  = ~A200 & \new_[11603]_ ;
  assign \new_[11605]_  = \new_[11604]_  & \new_[11599]_ ;
  assign \new_[11609]_  = A265 & A234;
  assign \new_[11610]_  = A233 & \new_[11609]_ ;
  assign \new_[11614]_  = ~A269 & A268;
  assign \new_[11615]_  = A266 & \new_[11614]_ ;
  assign \new_[11616]_  = \new_[11615]_  & \new_[11610]_ ;
  assign \new_[11620]_  = A199 & ~A166;
  assign \new_[11621]_  = A167 & \new_[11620]_ ;
  assign \new_[11625]_  = A202 & ~A201;
  assign \new_[11626]_  = ~A200 & \new_[11625]_ ;
  assign \new_[11627]_  = \new_[11626]_  & \new_[11621]_ ;
  assign \new_[11631]_  = ~A265 & A234;
  assign \new_[11632]_  = A233 & \new_[11631]_ ;
  assign \new_[11636]_  = A269 & ~A268;
  assign \new_[11637]_  = A266 & \new_[11636]_ ;
  assign \new_[11638]_  = \new_[11637]_  & \new_[11632]_ ;
  assign \new_[11642]_  = A199 & ~A166;
  assign \new_[11643]_  = A167 & \new_[11642]_ ;
  assign \new_[11647]_  = A202 & ~A201;
  assign \new_[11648]_  = ~A200 & \new_[11647]_ ;
  assign \new_[11649]_  = \new_[11648]_  & \new_[11643]_ ;
  assign \new_[11653]_  = A265 & A234;
  assign \new_[11654]_  = A233 & \new_[11653]_ ;
  assign \new_[11658]_  = A269 & ~A268;
  assign \new_[11659]_  = ~A266 & \new_[11658]_ ;
  assign \new_[11660]_  = \new_[11659]_  & \new_[11654]_ ;
  assign \new_[11664]_  = A199 & ~A166;
  assign \new_[11665]_  = A167 & \new_[11664]_ ;
  assign \new_[11669]_  = A202 & ~A201;
  assign \new_[11670]_  = ~A200 & \new_[11669]_ ;
  assign \new_[11671]_  = \new_[11670]_  & \new_[11665]_ ;
  assign \new_[11675]_  = ~A265 & A234;
  assign \new_[11676]_  = A233 & \new_[11675]_ ;
  assign \new_[11680]_  = ~A269 & A268;
  assign \new_[11681]_  = ~A266 & \new_[11680]_ ;
  assign \new_[11682]_  = \new_[11681]_  & \new_[11676]_ ;
  assign \new_[11686]_  = A199 & ~A166;
  assign \new_[11687]_  = A167 & \new_[11686]_ ;
  assign \new_[11691]_  = A202 & ~A201;
  assign \new_[11692]_  = ~A200 & \new_[11691]_ ;
  assign \new_[11693]_  = \new_[11692]_  & \new_[11687]_ ;
  assign \new_[11697]_  = A235 & A233;
  assign \new_[11698]_  = A232 & \new_[11697]_ ;
  assign \new_[11702]_  = A300 & A299;
  assign \new_[11703]_  = ~A236 & \new_[11702]_ ;
  assign \new_[11704]_  = \new_[11703]_  & \new_[11698]_ ;
  assign \new_[11708]_  = A199 & ~A166;
  assign \new_[11709]_  = A167 & \new_[11708]_ ;
  assign \new_[11713]_  = A202 & ~A201;
  assign \new_[11714]_  = ~A200 & \new_[11713]_ ;
  assign \new_[11715]_  = \new_[11714]_  & \new_[11709]_ ;
  assign \new_[11719]_  = A235 & A233;
  assign \new_[11720]_  = A232 & \new_[11719]_ ;
  assign \new_[11724]_  = A300 & A298;
  assign \new_[11725]_  = ~A236 & \new_[11724]_ ;
  assign \new_[11726]_  = \new_[11725]_  & \new_[11720]_ ;
  assign \new_[11730]_  = A199 & ~A166;
  assign \new_[11731]_  = A167 & \new_[11730]_ ;
  assign \new_[11735]_  = A202 & ~A201;
  assign \new_[11736]_  = ~A200 & \new_[11735]_ ;
  assign \new_[11737]_  = \new_[11736]_  & \new_[11731]_ ;
  assign \new_[11741]_  = A235 & A233;
  assign \new_[11742]_  = A232 & \new_[11741]_ ;
  assign \new_[11746]_  = A267 & A265;
  assign \new_[11747]_  = ~A236 & \new_[11746]_ ;
  assign \new_[11748]_  = \new_[11747]_  & \new_[11742]_ ;
  assign \new_[11752]_  = A199 & ~A166;
  assign \new_[11753]_  = A167 & \new_[11752]_ ;
  assign \new_[11757]_  = A202 & ~A201;
  assign \new_[11758]_  = ~A200 & \new_[11757]_ ;
  assign \new_[11759]_  = \new_[11758]_  & \new_[11753]_ ;
  assign \new_[11763]_  = A235 & A233;
  assign \new_[11764]_  = A232 & \new_[11763]_ ;
  assign \new_[11768]_  = A267 & A266;
  assign \new_[11769]_  = ~A236 & \new_[11768]_ ;
  assign \new_[11770]_  = \new_[11769]_  & \new_[11764]_ ;
  assign \new_[11774]_  = A199 & ~A166;
  assign \new_[11775]_  = A167 & \new_[11774]_ ;
  assign \new_[11779]_  = A202 & ~A201;
  assign \new_[11780]_  = ~A200 & \new_[11779]_ ;
  assign \new_[11781]_  = \new_[11780]_  & \new_[11775]_ ;
  assign \new_[11785]_  = ~A235 & A233;
  assign \new_[11786]_  = ~A232 & \new_[11785]_ ;
  assign \new_[11790]_  = A300 & A299;
  assign \new_[11791]_  = A236 & \new_[11790]_ ;
  assign \new_[11792]_  = \new_[11791]_  & \new_[11786]_ ;
  assign \new_[11796]_  = A199 & ~A166;
  assign \new_[11797]_  = A167 & \new_[11796]_ ;
  assign \new_[11801]_  = A202 & ~A201;
  assign \new_[11802]_  = ~A200 & \new_[11801]_ ;
  assign \new_[11803]_  = \new_[11802]_  & \new_[11797]_ ;
  assign \new_[11807]_  = ~A235 & A233;
  assign \new_[11808]_  = ~A232 & \new_[11807]_ ;
  assign \new_[11812]_  = A300 & A298;
  assign \new_[11813]_  = A236 & \new_[11812]_ ;
  assign \new_[11814]_  = \new_[11813]_  & \new_[11808]_ ;
  assign \new_[11818]_  = A199 & ~A166;
  assign \new_[11819]_  = A167 & \new_[11818]_ ;
  assign \new_[11823]_  = A202 & ~A201;
  assign \new_[11824]_  = ~A200 & \new_[11823]_ ;
  assign \new_[11825]_  = \new_[11824]_  & \new_[11819]_ ;
  assign \new_[11829]_  = ~A235 & A233;
  assign \new_[11830]_  = ~A232 & \new_[11829]_ ;
  assign \new_[11834]_  = A267 & A265;
  assign \new_[11835]_  = A236 & \new_[11834]_ ;
  assign \new_[11836]_  = \new_[11835]_  & \new_[11830]_ ;
  assign \new_[11840]_  = A199 & ~A166;
  assign \new_[11841]_  = A167 & \new_[11840]_ ;
  assign \new_[11845]_  = A202 & ~A201;
  assign \new_[11846]_  = ~A200 & \new_[11845]_ ;
  assign \new_[11847]_  = \new_[11846]_  & \new_[11841]_ ;
  assign \new_[11851]_  = ~A235 & A233;
  assign \new_[11852]_  = ~A232 & \new_[11851]_ ;
  assign \new_[11856]_  = A267 & A266;
  assign \new_[11857]_  = A236 & \new_[11856]_ ;
  assign \new_[11858]_  = \new_[11857]_  & \new_[11852]_ ;
  assign \new_[11862]_  = A199 & ~A166;
  assign \new_[11863]_  = A167 & \new_[11862]_ ;
  assign \new_[11867]_  = A202 & ~A201;
  assign \new_[11868]_  = ~A200 & \new_[11867]_ ;
  assign \new_[11869]_  = \new_[11868]_  & \new_[11863]_ ;
  assign \new_[11873]_  = ~A235 & ~A233;
  assign \new_[11874]_  = A232 & \new_[11873]_ ;
  assign \new_[11878]_  = A300 & A299;
  assign \new_[11879]_  = A236 & \new_[11878]_ ;
  assign \new_[11880]_  = \new_[11879]_  & \new_[11874]_ ;
  assign \new_[11884]_  = A199 & ~A166;
  assign \new_[11885]_  = A167 & \new_[11884]_ ;
  assign \new_[11889]_  = A202 & ~A201;
  assign \new_[11890]_  = ~A200 & \new_[11889]_ ;
  assign \new_[11891]_  = \new_[11890]_  & \new_[11885]_ ;
  assign \new_[11895]_  = ~A235 & ~A233;
  assign \new_[11896]_  = A232 & \new_[11895]_ ;
  assign \new_[11900]_  = A300 & A298;
  assign \new_[11901]_  = A236 & \new_[11900]_ ;
  assign \new_[11902]_  = \new_[11901]_  & \new_[11896]_ ;
  assign \new_[11906]_  = A199 & ~A166;
  assign \new_[11907]_  = A167 & \new_[11906]_ ;
  assign \new_[11911]_  = A202 & ~A201;
  assign \new_[11912]_  = ~A200 & \new_[11911]_ ;
  assign \new_[11913]_  = \new_[11912]_  & \new_[11907]_ ;
  assign \new_[11917]_  = ~A235 & ~A233;
  assign \new_[11918]_  = A232 & \new_[11917]_ ;
  assign \new_[11922]_  = A267 & A265;
  assign \new_[11923]_  = A236 & \new_[11922]_ ;
  assign \new_[11924]_  = \new_[11923]_  & \new_[11918]_ ;
  assign \new_[11928]_  = A199 & ~A166;
  assign \new_[11929]_  = A167 & \new_[11928]_ ;
  assign \new_[11933]_  = A202 & ~A201;
  assign \new_[11934]_  = ~A200 & \new_[11933]_ ;
  assign \new_[11935]_  = \new_[11934]_  & \new_[11929]_ ;
  assign \new_[11939]_  = ~A235 & ~A233;
  assign \new_[11940]_  = A232 & \new_[11939]_ ;
  assign \new_[11944]_  = A267 & A266;
  assign \new_[11945]_  = A236 & \new_[11944]_ ;
  assign \new_[11946]_  = \new_[11945]_  & \new_[11940]_ ;
  assign \new_[11950]_  = A199 & ~A166;
  assign \new_[11951]_  = A167 & \new_[11950]_ ;
  assign \new_[11955]_  = A202 & ~A201;
  assign \new_[11956]_  = ~A200 & \new_[11955]_ ;
  assign \new_[11957]_  = \new_[11956]_  & \new_[11951]_ ;
  assign \new_[11961]_  = A235 & ~A233;
  assign \new_[11962]_  = ~A232 & \new_[11961]_ ;
  assign \new_[11966]_  = A300 & A299;
  assign \new_[11967]_  = ~A236 & \new_[11966]_ ;
  assign \new_[11968]_  = \new_[11967]_  & \new_[11962]_ ;
  assign \new_[11972]_  = A199 & ~A166;
  assign \new_[11973]_  = A167 & \new_[11972]_ ;
  assign \new_[11977]_  = A202 & ~A201;
  assign \new_[11978]_  = ~A200 & \new_[11977]_ ;
  assign \new_[11979]_  = \new_[11978]_  & \new_[11973]_ ;
  assign \new_[11983]_  = A235 & ~A233;
  assign \new_[11984]_  = ~A232 & \new_[11983]_ ;
  assign \new_[11988]_  = A300 & A298;
  assign \new_[11989]_  = ~A236 & \new_[11988]_ ;
  assign \new_[11990]_  = \new_[11989]_  & \new_[11984]_ ;
  assign \new_[11994]_  = A199 & ~A166;
  assign \new_[11995]_  = A167 & \new_[11994]_ ;
  assign \new_[11999]_  = A202 & ~A201;
  assign \new_[12000]_  = ~A200 & \new_[11999]_ ;
  assign \new_[12001]_  = \new_[12000]_  & \new_[11995]_ ;
  assign \new_[12005]_  = A235 & ~A233;
  assign \new_[12006]_  = ~A232 & \new_[12005]_ ;
  assign \new_[12010]_  = A267 & A265;
  assign \new_[12011]_  = ~A236 & \new_[12010]_ ;
  assign \new_[12012]_  = \new_[12011]_  & \new_[12006]_ ;
  assign \new_[12016]_  = A199 & ~A166;
  assign \new_[12017]_  = A167 & \new_[12016]_ ;
  assign \new_[12021]_  = A202 & ~A201;
  assign \new_[12022]_  = ~A200 & \new_[12021]_ ;
  assign \new_[12023]_  = \new_[12022]_  & \new_[12017]_ ;
  assign \new_[12027]_  = A235 & ~A233;
  assign \new_[12028]_  = ~A232 & \new_[12027]_ ;
  assign \new_[12032]_  = A267 & A266;
  assign \new_[12033]_  = ~A236 & \new_[12032]_ ;
  assign \new_[12034]_  = \new_[12033]_  & \new_[12028]_ ;
  assign \new_[12038]_  = A199 & ~A166;
  assign \new_[12039]_  = A167 & \new_[12038]_ ;
  assign \new_[12043]_  = ~A203 & ~A201;
  assign \new_[12044]_  = ~A200 & \new_[12043]_ ;
  assign \new_[12045]_  = \new_[12044]_  & \new_[12039]_ ;
  assign \new_[12049]_  = A298 & A234;
  assign \new_[12050]_  = A232 & \new_[12049]_ ;
  assign \new_[12054]_  = ~A302 & A301;
  assign \new_[12055]_  = A299 & \new_[12054]_ ;
  assign \new_[12056]_  = \new_[12055]_  & \new_[12050]_ ;
  assign \new_[12060]_  = A199 & ~A166;
  assign \new_[12061]_  = A167 & \new_[12060]_ ;
  assign \new_[12065]_  = ~A203 & ~A201;
  assign \new_[12066]_  = ~A200 & \new_[12065]_ ;
  assign \new_[12067]_  = \new_[12066]_  & \new_[12061]_ ;
  assign \new_[12071]_  = A298 & A234;
  assign \new_[12072]_  = A232 & \new_[12071]_ ;
  assign \new_[12076]_  = A302 & ~A301;
  assign \new_[12077]_  = ~A299 & \new_[12076]_ ;
  assign \new_[12078]_  = \new_[12077]_  & \new_[12072]_ ;
  assign \new_[12082]_  = A199 & ~A166;
  assign \new_[12083]_  = A167 & \new_[12082]_ ;
  assign \new_[12087]_  = ~A203 & ~A201;
  assign \new_[12088]_  = ~A200 & \new_[12087]_ ;
  assign \new_[12089]_  = \new_[12088]_  & \new_[12083]_ ;
  assign \new_[12093]_  = ~A298 & A234;
  assign \new_[12094]_  = A232 & \new_[12093]_ ;
  assign \new_[12098]_  = A302 & ~A301;
  assign \new_[12099]_  = A299 & \new_[12098]_ ;
  assign \new_[12100]_  = \new_[12099]_  & \new_[12094]_ ;
  assign \new_[12104]_  = A199 & ~A166;
  assign \new_[12105]_  = A167 & \new_[12104]_ ;
  assign \new_[12109]_  = ~A203 & ~A201;
  assign \new_[12110]_  = ~A200 & \new_[12109]_ ;
  assign \new_[12111]_  = \new_[12110]_  & \new_[12105]_ ;
  assign \new_[12115]_  = ~A298 & A234;
  assign \new_[12116]_  = A232 & \new_[12115]_ ;
  assign \new_[12120]_  = ~A302 & A301;
  assign \new_[12121]_  = ~A299 & \new_[12120]_ ;
  assign \new_[12122]_  = \new_[12121]_  & \new_[12116]_ ;
  assign \new_[12126]_  = A199 & ~A166;
  assign \new_[12127]_  = A167 & \new_[12126]_ ;
  assign \new_[12131]_  = ~A203 & ~A201;
  assign \new_[12132]_  = ~A200 & \new_[12131]_ ;
  assign \new_[12133]_  = \new_[12132]_  & \new_[12127]_ ;
  assign \new_[12137]_  = A265 & A234;
  assign \new_[12138]_  = A232 & \new_[12137]_ ;
  assign \new_[12142]_  = ~A269 & A268;
  assign \new_[12143]_  = A266 & \new_[12142]_ ;
  assign \new_[12144]_  = \new_[12143]_  & \new_[12138]_ ;
  assign \new_[12148]_  = A199 & ~A166;
  assign \new_[12149]_  = A167 & \new_[12148]_ ;
  assign \new_[12153]_  = ~A203 & ~A201;
  assign \new_[12154]_  = ~A200 & \new_[12153]_ ;
  assign \new_[12155]_  = \new_[12154]_  & \new_[12149]_ ;
  assign \new_[12159]_  = ~A265 & A234;
  assign \new_[12160]_  = A232 & \new_[12159]_ ;
  assign \new_[12164]_  = A269 & ~A268;
  assign \new_[12165]_  = A266 & \new_[12164]_ ;
  assign \new_[12166]_  = \new_[12165]_  & \new_[12160]_ ;
  assign \new_[12170]_  = A199 & ~A166;
  assign \new_[12171]_  = A167 & \new_[12170]_ ;
  assign \new_[12175]_  = ~A203 & ~A201;
  assign \new_[12176]_  = ~A200 & \new_[12175]_ ;
  assign \new_[12177]_  = \new_[12176]_  & \new_[12171]_ ;
  assign \new_[12181]_  = A265 & A234;
  assign \new_[12182]_  = A232 & \new_[12181]_ ;
  assign \new_[12186]_  = A269 & ~A268;
  assign \new_[12187]_  = ~A266 & \new_[12186]_ ;
  assign \new_[12188]_  = \new_[12187]_  & \new_[12182]_ ;
  assign \new_[12192]_  = A199 & ~A166;
  assign \new_[12193]_  = A167 & \new_[12192]_ ;
  assign \new_[12197]_  = ~A203 & ~A201;
  assign \new_[12198]_  = ~A200 & \new_[12197]_ ;
  assign \new_[12199]_  = \new_[12198]_  & \new_[12193]_ ;
  assign \new_[12203]_  = ~A265 & A234;
  assign \new_[12204]_  = A232 & \new_[12203]_ ;
  assign \new_[12208]_  = ~A269 & A268;
  assign \new_[12209]_  = ~A266 & \new_[12208]_ ;
  assign \new_[12210]_  = \new_[12209]_  & \new_[12204]_ ;
  assign \new_[12214]_  = A199 & ~A166;
  assign \new_[12215]_  = A167 & \new_[12214]_ ;
  assign \new_[12219]_  = ~A203 & ~A201;
  assign \new_[12220]_  = ~A200 & \new_[12219]_ ;
  assign \new_[12221]_  = \new_[12220]_  & \new_[12215]_ ;
  assign \new_[12225]_  = A298 & A234;
  assign \new_[12226]_  = A233 & \new_[12225]_ ;
  assign \new_[12230]_  = ~A302 & A301;
  assign \new_[12231]_  = A299 & \new_[12230]_ ;
  assign \new_[12232]_  = \new_[12231]_  & \new_[12226]_ ;
  assign \new_[12236]_  = A199 & ~A166;
  assign \new_[12237]_  = A167 & \new_[12236]_ ;
  assign \new_[12241]_  = ~A203 & ~A201;
  assign \new_[12242]_  = ~A200 & \new_[12241]_ ;
  assign \new_[12243]_  = \new_[12242]_  & \new_[12237]_ ;
  assign \new_[12247]_  = A298 & A234;
  assign \new_[12248]_  = A233 & \new_[12247]_ ;
  assign \new_[12252]_  = A302 & ~A301;
  assign \new_[12253]_  = ~A299 & \new_[12252]_ ;
  assign \new_[12254]_  = \new_[12253]_  & \new_[12248]_ ;
  assign \new_[12258]_  = A199 & ~A166;
  assign \new_[12259]_  = A167 & \new_[12258]_ ;
  assign \new_[12263]_  = ~A203 & ~A201;
  assign \new_[12264]_  = ~A200 & \new_[12263]_ ;
  assign \new_[12265]_  = \new_[12264]_  & \new_[12259]_ ;
  assign \new_[12269]_  = ~A298 & A234;
  assign \new_[12270]_  = A233 & \new_[12269]_ ;
  assign \new_[12274]_  = A302 & ~A301;
  assign \new_[12275]_  = A299 & \new_[12274]_ ;
  assign \new_[12276]_  = \new_[12275]_  & \new_[12270]_ ;
  assign \new_[12280]_  = A199 & ~A166;
  assign \new_[12281]_  = A167 & \new_[12280]_ ;
  assign \new_[12285]_  = ~A203 & ~A201;
  assign \new_[12286]_  = ~A200 & \new_[12285]_ ;
  assign \new_[12287]_  = \new_[12286]_  & \new_[12281]_ ;
  assign \new_[12291]_  = ~A298 & A234;
  assign \new_[12292]_  = A233 & \new_[12291]_ ;
  assign \new_[12296]_  = ~A302 & A301;
  assign \new_[12297]_  = ~A299 & \new_[12296]_ ;
  assign \new_[12298]_  = \new_[12297]_  & \new_[12292]_ ;
  assign \new_[12302]_  = A199 & ~A166;
  assign \new_[12303]_  = A167 & \new_[12302]_ ;
  assign \new_[12307]_  = ~A203 & ~A201;
  assign \new_[12308]_  = ~A200 & \new_[12307]_ ;
  assign \new_[12309]_  = \new_[12308]_  & \new_[12303]_ ;
  assign \new_[12313]_  = A265 & A234;
  assign \new_[12314]_  = A233 & \new_[12313]_ ;
  assign \new_[12318]_  = ~A269 & A268;
  assign \new_[12319]_  = A266 & \new_[12318]_ ;
  assign \new_[12320]_  = \new_[12319]_  & \new_[12314]_ ;
  assign \new_[12324]_  = A199 & ~A166;
  assign \new_[12325]_  = A167 & \new_[12324]_ ;
  assign \new_[12329]_  = ~A203 & ~A201;
  assign \new_[12330]_  = ~A200 & \new_[12329]_ ;
  assign \new_[12331]_  = \new_[12330]_  & \new_[12325]_ ;
  assign \new_[12335]_  = ~A265 & A234;
  assign \new_[12336]_  = A233 & \new_[12335]_ ;
  assign \new_[12340]_  = A269 & ~A268;
  assign \new_[12341]_  = A266 & \new_[12340]_ ;
  assign \new_[12342]_  = \new_[12341]_  & \new_[12336]_ ;
  assign \new_[12346]_  = A199 & ~A166;
  assign \new_[12347]_  = A167 & \new_[12346]_ ;
  assign \new_[12351]_  = ~A203 & ~A201;
  assign \new_[12352]_  = ~A200 & \new_[12351]_ ;
  assign \new_[12353]_  = \new_[12352]_  & \new_[12347]_ ;
  assign \new_[12357]_  = A265 & A234;
  assign \new_[12358]_  = A233 & \new_[12357]_ ;
  assign \new_[12362]_  = A269 & ~A268;
  assign \new_[12363]_  = ~A266 & \new_[12362]_ ;
  assign \new_[12364]_  = \new_[12363]_  & \new_[12358]_ ;
  assign \new_[12368]_  = A199 & ~A166;
  assign \new_[12369]_  = A167 & \new_[12368]_ ;
  assign \new_[12373]_  = ~A203 & ~A201;
  assign \new_[12374]_  = ~A200 & \new_[12373]_ ;
  assign \new_[12375]_  = \new_[12374]_  & \new_[12369]_ ;
  assign \new_[12379]_  = ~A265 & A234;
  assign \new_[12380]_  = A233 & \new_[12379]_ ;
  assign \new_[12384]_  = ~A269 & A268;
  assign \new_[12385]_  = ~A266 & \new_[12384]_ ;
  assign \new_[12386]_  = \new_[12385]_  & \new_[12380]_ ;
  assign \new_[12390]_  = A199 & ~A166;
  assign \new_[12391]_  = A167 & \new_[12390]_ ;
  assign \new_[12395]_  = ~A203 & ~A201;
  assign \new_[12396]_  = ~A200 & \new_[12395]_ ;
  assign \new_[12397]_  = \new_[12396]_  & \new_[12391]_ ;
  assign \new_[12401]_  = A235 & A233;
  assign \new_[12402]_  = A232 & \new_[12401]_ ;
  assign \new_[12406]_  = A300 & A299;
  assign \new_[12407]_  = ~A236 & \new_[12406]_ ;
  assign \new_[12408]_  = \new_[12407]_  & \new_[12402]_ ;
  assign \new_[12412]_  = A199 & ~A166;
  assign \new_[12413]_  = A167 & \new_[12412]_ ;
  assign \new_[12417]_  = ~A203 & ~A201;
  assign \new_[12418]_  = ~A200 & \new_[12417]_ ;
  assign \new_[12419]_  = \new_[12418]_  & \new_[12413]_ ;
  assign \new_[12423]_  = A235 & A233;
  assign \new_[12424]_  = A232 & \new_[12423]_ ;
  assign \new_[12428]_  = A300 & A298;
  assign \new_[12429]_  = ~A236 & \new_[12428]_ ;
  assign \new_[12430]_  = \new_[12429]_  & \new_[12424]_ ;
  assign \new_[12434]_  = A199 & ~A166;
  assign \new_[12435]_  = A167 & \new_[12434]_ ;
  assign \new_[12439]_  = ~A203 & ~A201;
  assign \new_[12440]_  = ~A200 & \new_[12439]_ ;
  assign \new_[12441]_  = \new_[12440]_  & \new_[12435]_ ;
  assign \new_[12445]_  = A235 & A233;
  assign \new_[12446]_  = A232 & \new_[12445]_ ;
  assign \new_[12450]_  = A267 & A265;
  assign \new_[12451]_  = ~A236 & \new_[12450]_ ;
  assign \new_[12452]_  = \new_[12451]_  & \new_[12446]_ ;
  assign \new_[12456]_  = A199 & ~A166;
  assign \new_[12457]_  = A167 & \new_[12456]_ ;
  assign \new_[12461]_  = ~A203 & ~A201;
  assign \new_[12462]_  = ~A200 & \new_[12461]_ ;
  assign \new_[12463]_  = \new_[12462]_  & \new_[12457]_ ;
  assign \new_[12467]_  = A235 & A233;
  assign \new_[12468]_  = A232 & \new_[12467]_ ;
  assign \new_[12472]_  = A267 & A266;
  assign \new_[12473]_  = ~A236 & \new_[12472]_ ;
  assign \new_[12474]_  = \new_[12473]_  & \new_[12468]_ ;
  assign \new_[12478]_  = A199 & ~A166;
  assign \new_[12479]_  = A167 & \new_[12478]_ ;
  assign \new_[12483]_  = ~A203 & ~A201;
  assign \new_[12484]_  = ~A200 & \new_[12483]_ ;
  assign \new_[12485]_  = \new_[12484]_  & \new_[12479]_ ;
  assign \new_[12489]_  = ~A235 & A233;
  assign \new_[12490]_  = ~A232 & \new_[12489]_ ;
  assign \new_[12494]_  = A300 & A299;
  assign \new_[12495]_  = A236 & \new_[12494]_ ;
  assign \new_[12496]_  = \new_[12495]_  & \new_[12490]_ ;
  assign \new_[12500]_  = A199 & ~A166;
  assign \new_[12501]_  = A167 & \new_[12500]_ ;
  assign \new_[12505]_  = ~A203 & ~A201;
  assign \new_[12506]_  = ~A200 & \new_[12505]_ ;
  assign \new_[12507]_  = \new_[12506]_  & \new_[12501]_ ;
  assign \new_[12511]_  = ~A235 & A233;
  assign \new_[12512]_  = ~A232 & \new_[12511]_ ;
  assign \new_[12516]_  = A300 & A298;
  assign \new_[12517]_  = A236 & \new_[12516]_ ;
  assign \new_[12518]_  = \new_[12517]_  & \new_[12512]_ ;
  assign \new_[12522]_  = A199 & ~A166;
  assign \new_[12523]_  = A167 & \new_[12522]_ ;
  assign \new_[12527]_  = ~A203 & ~A201;
  assign \new_[12528]_  = ~A200 & \new_[12527]_ ;
  assign \new_[12529]_  = \new_[12528]_  & \new_[12523]_ ;
  assign \new_[12533]_  = ~A235 & A233;
  assign \new_[12534]_  = ~A232 & \new_[12533]_ ;
  assign \new_[12538]_  = A267 & A265;
  assign \new_[12539]_  = A236 & \new_[12538]_ ;
  assign \new_[12540]_  = \new_[12539]_  & \new_[12534]_ ;
  assign \new_[12544]_  = A199 & ~A166;
  assign \new_[12545]_  = A167 & \new_[12544]_ ;
  assign \new_[12549]_  = ~A203 & ~A201;
  assign \new_[12550]_  = ~A200 & \new_[12549]_ ;
  assign \new_[12551]_  = \new_[12550]_  & \new_[12545]_ ;
  assign \new_[12555]_  = ~A235 & A233;
  assign \new_[12556]_  = ~A232 & \new_[12555]_ ;
  assign \new_[12560]_  = A267 & A266;
  assign \new_[12561]_  = A236 & \new_[12560]_ ;
  assign \new_[12562]_  = \new_[12561]_  & \new_[12556]_ ;
  assign \new_[12566]_  = A199 & ~A166;
  assign \new_[12567]_  = A167 & \new_[12566]_ ;
  assign \new_[12571]_  = ~A203 & ~A201;
  assign \new_[12572]_  = ~A200 & \new_[12571]_ ;
  assign \new_[12573]_  = \new_[12572]_  & \new_[12567]_ ;
  assign \new_[12577]_  = ~A235 & ~A233;
  assign \new_[12578]_  = A232 & \new_[12577]_ ;
  assign \new_[12582]_  = A300 & A299;
  assign \new_[12583]_  = A236 & \new_[12582]_ ;
  assign \new_[12584]_  = \new_[12583]_  & \new_[12578]_ ;
  assign \new_[12588]_  = A199 & ~A166;
  assign \new_[12589]_  = A167 & \new_[12588]_ ;
  assign \new_[12593]_  = ~A203 & ~A201;
  assign \new_[12594]_  = ~A200 & \new_[12593]_ ;
  assign \new_[12595]_  = \new_[12594]_  & \new_[12589]_ ;
  assign \new_[12599]_  = ~A235 & ~A233;
  assign \new_[12600]_  = A232 & \new_[12599]_ ;
  assign \new_[12604]_  = A300 & A298;
  assign \new_[12605]_  = A236 & \new_[12604]_ ;
  assign \new_[12606]_  = \new_[12605]_  & \new_[12600]_ ;
  assign \new_[12610]_  = A199 & ~A166;
  assign \new_[12611]_  = A167 & \new_[12610]_ ;
  assign \new_[12615]_  = ~A203 & ~A201;
  assign \new_[12616]_  = ~A200 & \new_[12615]_ ;
  assign \new_[12617]_  = \new_[12616]_  & \new_[12611]_ ;
  assign \new_[12621]_  = ~A235 & ~A233;
  assign \new_[12622]_  = A232 & \new_[12621]_ ;
  assign \new_[12626]_  = A267 & A265;
  assign \new_[12627]_  = A236 & \new_[12626]_ ;
  assign \new_[12628]_  = \new_[12627]_  & \new_[12622]_ ;
  assign \new_[12632]_  = A199 & ~A166;
  assign \new_[12633]_  = A167 & \new_[12632]_ ;
  assign \new_[12637]_  = ~A203 & ~A201;
  assign \new_[12638]_  = ~A200 & \new_[12637]_ ;
  assign \new_[12639]_  = \new_[12638]_  & \new_[12633]_ ;
  assign \new_[12643]_  = ~A235 & ~A233;
  assign \new_[12644]_  = A232 & \new_[12643]_ ;
  assign \new_[12648]_  = A267 & A266;
  assign \new_[12649]_  = A236 & \new_[12648]_ ;
  assign \new_[12650]_  = \new_[12649]_  & \new_[12644]_ ;
  assign \new_[12654]_  = A199 & ~A166;
  assign \new_[12655]_  = A167 & \new_[12654]_ ;
  assign \new_[12659]_  = ~A203 & ~A201;
  assign \new_[12660]_  = ~A200 & \new_[12659]_ ;
  assign \new_[12661]_  = \new_[12660]_  & \new_[12655]_ ;
  assign \new_[12665]_  = A235 & ~A233;
  assign \new_[12666]_  = ~A232 & \new_[12665]_ ;
  assign \new_[12670]_  = A300 & A299;
  assign \new_[12671]_  = ~A236 & \new_[12670]_ ;
  assign \new_[12672]_  = \new_[12671]_  & \new_[12666]_ ;
  assign \new_[12676]_  = A199 & ~A166;
  assign \new_[12677]_  = A167 & \new_[12676]_ ;
  assign \new_[12681]_  = ~A203 & ~A201;
  assign \new_[12682]_  = ~A200 & \new_[12681]_ ;
  assign \new_[12683]_  = \new_[12682]_  & \new_[12677]_ ;
  assign \new_[12687]_  = A235 & ~A233;
  assign \new_[12688]_  = ~A232 & \new_[12687]_ ;
  assign \new_[12692]_  = A300 & A298;
  assign \new_[12693]_  = ~A236 & \new_[12692]_ ;
  assign \new_[12694]_  = \new_[12693]_  & \new_[12688]_ ;
  assign \new_[12698]_  = A199 & ~A166;
  assign \new_[12699]_  = A167 & \new_[12698]_ ;
  assign \new_[12703]_  = ~A203 & ~A201;
  assign \new_[12704]_  = ~A200 & \new_[12703]_ ;
  assign \new_[12705]_  = \new_[12704]_  & \new_[12699]_ ;
  assign \new_[12709]_  = A235 & ~A233;
  assign \new_[12710]_  = ~A232 & \new_[12709]_ ;
  assign \new_[12714]_  = A267 & A265;
  assign \new_[12715]_  = ~A236 & \new_[12714]_ ;
  assign \new_[12716]_  = \new_[12715]_  & \new_[12710]_ ;
  assign \new_[12720]_  = A199 & ~A166;
  assign \new_[12721]_  = A167 & \new_[12720]_ ;
  assign \new_[12725]_  = ~A203 & ~A201;
  assign \new_[12726]_  = ~A200 & \new_[12725]_ ;
  assign \new_[12727]_  = \new_[12726]_  & \new_[12721]_ ;
  assign \new_[12731]_  = A235 & ~A233;
  assign \new_[12732]_  = ~A232 & \new_[12731]_ ;
  assign \new_[12736]_  = A267 & A266;
  assign \new_[12737]_  = ~A236 & \new_[12736]_ ;
  assign \new_[12738]_  = \new_[12737]_  & \new_[12732]_ ;
  assign \new_[12742]_  = ~A167 & A168;
  assign \new_[12743]_  = A170 & \new_[12742]_ ;
  assign \new_[12747]_  = A200 & A199;
  assign \new_[12748]_  = A166 & \new_[12747]_ ;
  assign \new_[12749]_  = \new_[12748]_  & \new_[12743]_ ;
  assign \new_[12753]_  = A232 & ~A202;
  assign \new_[12754]_  = ~A201 & \new_[12753]_ ;
  assign \new_[12758]_  = A300 & A299;
  assign \new_[12759]_  = A234 & \new_[12758]_ ;
  assign \new_[12760]_  = \new_[12759]_  & \new_[12754]_ ;
  assign \new_[12764]_  = ~A167 & A168;
  assign \new_[12765]_  = A170 & \new_[12764]_ ;
  assign \new_[12769]_  = A200 & A199;
  assign \new_[12770]_  = A166 & \new_[12769]_ ;
  assign \new_[12771]_  = \new_[12770]_  & \new_[12765]_ ;
  assign \new_[12775]_  = A232 & ~A202;
  assign \new_[12776]_  = ~A201 & \new_[12775]_ ;
  assign \new_[12780]_  = A300 & A298;
  assign \new_[12781]_  = A234 & \new_[12780]_ ;
  assign \new_[12782]_  = \new_[12781]_  & \new_[12776]_ ;
  assign \new_[12786]_  = ~A167 & A168;
  assign \new_[12787]_  = A170 & \new_[12786]_ ;
  assign \new_[12791]_  = A200 & A199;
  assign \new_[12792]_  = A166 & \new_[12791]_ ;
  assign \new_[12793]_  = \new_[12792]_  & \new_[12787]_ ;
  assign \new_[12797]_  = A232 & ~A202;
  assign \new_[12798]_  = ~A201 & \new_[12797]_ ;
  assign \new_[12802]_  = A267 & A265;
  assign \new_[12803]_  = A234 & \new_[12802]_ ;
  assign \new_[12804]_  = \new_[12803]_  & \new_[12798]_ ;
  assign \new_[12808]_  = ~A167 & A168;
  assign \new_[12809]_  = A170 & \new_[12808]_ ;
  assign \new_[12813]_  = A200 & A199;
  assign \new_[12814]_  = A166 & \new_[12813]_ ;
  assign \new_[12815]_  = \new_[12814]_  & \new_[12809]_ ;
  assign \new_[12819]_  = A232 & ~A202;
  assign \new_[12820]_  = ~A201 & \new_[12819]_ ;
  assign \new_[12824]_  = A267 & A266;
  assign \new_[12825]_  = A234 & \new_[12824]_ ;
  assign \new_[12826]_  = \new_[12825]_  & \new_[12820]_ ;
  assign \new_[12830]_  = ~A167 & A168;
  assign \new_[12831]_  = A170 & \new_[12830]_ ;
  assign \new_[12835]_  = A200 & A199;
  assign \new_[12836]_  = A166 & \new_[12835]_ ;
  assign \new_[12837]_  = \new_[12836]_  & \new_[12831]_ ;
  assign \new_[12841]_  = A233 & ~A202;
  assign \new_[12842]_  = ~A201 & \new_[12841]_ ;
  assign \new_[12846]_  = A300 & A299;
  assign \new_[12847]_  = A234 & \new_[12846]_ ;
  assign \new_[12848]_  = \new_[12847]_  & \new_[12842]_ ;
  assign \new_[12852]_  = ~A167 & A168;
  assign \new_[12853]_  = A170 & \new_[12852]_ ;
  assign \new_[12857]_  = A200 & A199;
  assign \new_[12858]_  = A166 & \new_[12857]_ ;
  assign \new_[12859]_  = \new_[12858]_  & \new_[12853]_ ;
  assign \new_[12863]_  = A233 & ~A202;
  assign \new_[12864]_  = ~A201 & \new_[12863]_ ;
  assign \new_[12868]_  = A300 & A298;
  assign \new_[12869]_  = A234 & \new_[12868]_ ;
  assign \new_[12870]_  = \new_[12869]_  & \new_[12864]_ ;
  assign \new_[12874]_  = ~A167 & A168;
  assign \new_[12875]_  = A170 & \new_[12874]_ ;
  assign \new_[12879]_  = A200 & A199;
  assign \new_[12880]_  = A166 & \new_[12879]_ ;
  assign \new_[12881]_  = \new_[12880]_  & \new_[12875]_ ;
  assign \new_[12885]_  = A233 & ~A202;
  assign \new_[12886]_  = ~A201 & \new_[12885]_ ;
  assign \new_[12890]_  = A267 & A265;
  assign \new_[12891]_  = A234 & \new_[12890]_ ;
  assign \new_[12892]_  = \new_[12891]_  & \new_[12886]_ ;
  assign \new_[12896]_  = ~A167 & A168;
  assign \new_[12897]_  = A170 & \new_[12896]_ ;
  assign \new_[12901]_  = A200 & A199;
  assign \new_[12902]_  = A166 & \new_[12901]_ ;
  assign \new_[12903]_  = \new_[12902]_  & \new_[12897]_ ;
  assign \new_[12907]_  = A233 & ~A202;
  assign \new_[12908]_  = ~A201 & \new_[12907]_ ;
  assign \new_[12912]_  = A267 & A266;
  assign \new_[12913]_  = A234 & \new_[12912]_ ;
  assign \new_[12914]_  = \new_[12913]_  & \new_[12908]_ ;
  assign \new_[12918]_  = ~A167 & A168;
  assign \new_[12919]_  = A170 & \new_[12918]_ ;
  assign \new_[12923]_  = A200 & A199;
  assign \new_[12924]_  = A166 & \new_[12923]_ ;
  assign \new_[12925]_  = \new_[12924]_  & \new_[12919]_ ;
  assign \new_[12929]_  = A232 & A203;
  assign \new_[12930]_  = ~A201 & \new_[12929]_ ;
  assign \new_[12934]_  = A300 & A299;
  assign \new_[12935]_  = A234 & \new_[12934]_ ;
  assign \new_[12936]_  = \new_[12935]_  & \new_[12930]_ ;
  assign \new_[12940]_  = ~A167 & A168;
  assign \new_[12941]_  = A170 & \new_[12940]_ ;
  assign \new_[12945]_  = A200 & A199;
  assign \new_[12946]_  = A166 & \new_[12945]_ ;
  assign \new_[12947]_  = \new_[12946]_  & \new_[12941]_ ;
  assign \new_[12951]_  = A232 & A203;
  assign \new_[12952]_  = ~A201 & \new_[12951]_ ;
  assign \new_[12956]_  = A300 & A298;
  assign \new_[12957]_  = A234 & \new_[12956]_ ;
  assign \new_[12958]_  = \new_[12957]_  & \new_[12952]_ ;
  assign \new_[12962]_  = ~A167 & A168;
  assign \new_[12963]_  = A170 & \new_[12962]_ ;
  assign \new_[12967]_  = A200 & A199;
  assign \new_[12968]_  = A166 & \new_[12967]_ ;
  assign \new_[12969]_  = \new_[12968]_  & \new_[12963]_ ;
  assign \new_[12973]_  = A232 & A203;
  assign \new_[12974]_  = ~A201 & \new_[12973]_ ;
  assign \new_[12978]_  = A267 & A265;
  assign \new_[12979]_  = A234 & \new_[12978]_ ;
  assign \new_[12980]_  = \new_[12979]_  & \new_[12974]_ ;
  assign \new_[12984]_  = ~A167 & A168;
  assign \new_[12985]_  = A170 & \new_[12984]_ ;
  assign \new_[12989]_  = A200 & A199;
  assign \new_[12990]_  = A166 & \new_[12989]_ ;
  assign \new_[12991]_  = \new_[12990]_  & \new_[12985]_ ;
  assign \new_[12995]_  = A232 & A203;
  assign \new_[12996]_  = ~A201 & \new_[12995]_ ;
  assign \new_[13000]_  = A267 & A266;
  assign \new_[13001]_  = A234 & \new_[13000]_ ;
  assign \new_[13002]_  = \new_[13001]_  & \new_[12996]_ ;
  assign \new_[13006]_  = ~A167 & A168;
  assign \new_[13007]_  = A170 & \new_[13006]_ ;
  assign \new_[13011]_  = A200 & A199;
  assign \new_[13012]_  = A166 & \new_[13011]_ ;
  assign \new_[13013]_  = \new_[13012]_  & \new_[13007]_ ;
  assign \new_[13017]_  = A233 & A203;
  assign \new_[13018]_  = ~A201 & \new_[13017]_ ;
  assign \new_[13022]_  = A300 & A299;
  assign \new_[13023]_  = A234 & \new_[13022]_ ;
  assign \new_[13024]_  = \new_[13023]_  & \new_[13018]_ ;
  assign \new_[13028]_  = ~A167 & A168;
  assign \new_[13029]_  = A170 & \new_[13028]_ ;
  assign \new_[13033]_  = A200 & A199;
  assign \new_[13034]_  = A166 & \new_[13033]_ ;
  assign \new_[13035]_  = \new_[13034]_  & \new_[13029]_ ;
  assign \new_[13039]_  = A233 & A203;
  assign \new_[13040]_  = ~A201 & \new_[13039]_ ;
  assign \new_[13044]_  = A300 & A298;
  assign \new_[13045]_  = A234 & \new_[13044]_ ;
  assign \new_[13046]_  = \new_[13045]_  & \new_[13040]_ ;
  assign \new_[13050]_  = ~A167 & A168;
  assign \new_[13051]_  = A170 & \new_[13050]_ ;
  assign \new_[13055]_  = A200 & A199;
  assign \new_[13056]_  = A166 & \new_[13055]_ ;
  assign \new_[13057]_  = \new_[13056]_  & \new_[13051]_ ;
  assign \new_[13061]_  = A233 & A203;
  assign \new_[13062]_  = ~A201 & \new_[13061]_ ;
  assign \new_[13066]_  = A267 & A265;
  assign \new_[13067]_  = A234 & \new_[13066]_ ;
  assign \new_[13068]_  = \new_[13067]_  & \new_[13062]_ ;
  assign \new_[13072]_  = ~A167 & A168;
  assign \new_[13073]_  = A170 & \new_[13072]_ ;
  assign \new_[13077]_  = A200 & A199;
  assign \new_[13078]_  = A166 & \new_[13077]_ ;
  assign \new_[13079]_  = \new_[13078]_  & \new_[13073]_ ;
  assign \new_[13083]_  = A233 & A203;
  assign \new_[13084]_  = ~A201 & \new_[13083]_ ;
  assign \new_[13088]_  = A267 & A266;
  assign \new_[13089]_  = A234 & \new_[13088]_ ;
  assign \new_[13090]_  = \new_[13089]_  & \new_[13084]_ ;
  assign \new_[13094]_  = ~A167 & A168;
  assign \new_[13095]_  = A170 & \new_[13094]_ ;
  assign \new_[13099]_  = A200 & ~A199;
  assign \new_[13100]_  = A166 & \new_[13099]_ ;
  assign \new_[13101]_  = \new_[13100]_  & \new_[13095]_ ;
  assign \new_[13105]_  = A232 & A202;
  assign \new_[13106]_  = ~A201 & \new_[13105]_ ;
  assign \new_[13110]_  = A300 & A299;
  assign \new_[13111]_  = A234 & \new_[13110]_ ;
  assign \new_[13112]_  = \new_[13111]_  & \new_[13106]_ ;
  assign \new_[13116]_  = ~A167 & A168;
  assign \new_[13117]_  = A170 & \new_[13116]_ ;
  assign \new_[13121]_  = A200 & ~A199;
  assign \new_[13122]_  = A166 & \new_[13121]_ ;
  assign \new_[13123]_  = \new_[13122]_  & \new_[13117]_ ;
  assign \new_[13127]_  = A232 & A202;
  assign \new_[13128]_  = ~A201 & \new_[13127]_ ;
  assign \new_[13132]_  = A300 & A298;
  assign \new_[13133]_  = A234 & \new_[13132]_ ;
  assign \new_[13134]_  = \new_[13133]_  & \new_[13128]_ ;
  assign \new_[13138]_  = ~A167 & A168;
  assign \new_[13139]_  = A170 & \new_[13138]_ ;
  assign \new_[13143]_  = A200 & ~A199;
  assign \new_[13144]_  = A166 & \new_[13143]_ ;
  assign \new_[13145]_  = \new_[13144]_  & \new_[13139]_ ;
  assign \new_[13149]_  = A232 & A202;
  assign \new_[13150]_  = ~A201 & \new_[13149]_ ;
  assign \new_[13154]_  = A267 & A265;
  assign \new_[13155]_  = A234 & \new_[13154]_ ;
  assign \new_[13156]_  = \new_[13155]_  & \new_[13150]_ ;
  assign \new_[13160]_  = ~A167 & A168;
  assign \new_[13161]_  = A170 & \new_[13160]_ ;
  assign \new_[13165]_  = A200 & ~A199;
  assign \new_[13166]_  = A166 & \new_[13165]_ ;
  assign \new_[13167]_  = \new_[13166]_  & \new_[13161]_ ;
  assign \new_[13171]_  = A232 & A202;
  assign \new_[13172]_  = ~A201 & \new_[13171]_ ;
  assign \new_[13176]_  = A267 & A266;
  assign \new_[13177]_  = A234 & \new_[13176]_ ;
  assign \new_[13178]_  = \new_[13177]_  & \new_[13172]_ ;
  assign \new_[13182]_  = ~A167 & A168;
  assign \new_[13183]_  = A170 & \new_[13182]_ ;
  assign \new_[13187]_  = A200 & ~A199;
  assign \new_[13188]_  = A166 & \new_[13187]_ ;
  assign \new_[13189]_  = \new_[13188]_  & \new_[13183]_ ;
  assign \new_[13193]_  = A233 & A202;
  assign \new_[13194]_  = ~A201 & \new_[13193]_ ;
  assign \new_[13198]_  = A300 & A299;
  assign \new_[13199]_  = A234 & \new_[13198]_ ;
  assign \new_[13200]_  = \new_[13199]_  & \new_[13194]_ ;
  assign \new_[13204]_  = ~A167 & A168;
  assign \new_[13205]_  = A170 & \new_[13204]_ ;
  assign \new_[13209]_  = A200 & ~A199;
  assign \new_[13210]_  = A166 & \new_[13209]_ ;
  assign \new_[13211]_  = \new_[13210]_  & \new_[13205]_ ;
  assign \new_[13215]_  = A233 & A202;
  assign \new_[13216]_  = ~A201 & \new_[13215]_ ;
  assign \new_[13220]_  = A300 & A298;
  assign \new_[13221]_  = A234 & \new_[13220]_ ;
  assign \new_[13222]_  = \new_[13221]_  & \new_[13216]_ ;
  assign \new_[13226]_  = ~A167 & A168;
  assign \new_[13227]_  = A170 & \new_[13226]_ ;
  assign \new_[13231]_  = A200 & ~A199;
  assign \new_[13232]_  = A166 & \new_[13231]_ ;
  assign \new_[13233]_  = \new_[13232]_  & \new_[13227]_ ;
  assign \new_[13237]_  = A233 & A202;
  assign \new_[13238]_  = ~A201 & \new_[13237]_ ;
  assign \new_[13242]_  = A267 & A265;
  assign \new_[13243]_  = A234 & \new_[13242]_ ;
  assign \new_[13244]_  = \new_[13243]_  & \new_[13238]_ ;
  assign \new_[13248]_  = ~A167 & A168;
  assign \new_[13249]_  = A170 & \new_[13248]_ ;
  assign \new_[13253]_  = A200 & ~A199;
  assign \new_[13254]_  = A166 & \new_[13253]_ ;
  assign \new_[13255]_  = \new_[13254]_  & \new_[13249]_ ;
  assign \new_[13259]_  = A233 & A202;
  assign \new_[13260]_  = ~A201 & \new_[13259]_ ;
  assign \new_[13264]_  = A267 & A266;
  assign \new_[13265]_  = A234 & \new_[13264]_ ;
  assign \new_[13266]_  = \new_[13265]_  & \new_[13260]_ ;
  assign \new_[13270]_  = ~A167 & A168;
  assign \new_[13271]_  = A170 & \new_[13270]_ ;
  assign \new_[13275]_  = A200 & ~A199;
  assign \new_[13276]_  = A166 & \new_[13275]_ ;
  assign \new_[13277]_  = \new_[13276]_  & \new_[13271]_ ;
  assign \new_[13281]_  = A232 & ~A203;
  assign \new_[13282]_  = ~A201 & \new_[13281]_ ;
  assign \new_[13286]_  = A300 & A299;
  assign \new_[13287]_  = A234 & \new_[13286]_ ;
  assign \new_[13288]_  = \new_[13287]_  & \new_[13282]_ ;
  assign \new_[13292]_  = ~A167 & A168;
  assign \new_[13293]_  = A170 & \new_[13292]_ ;
  assign \new_[13297]_  = A200 & ~A199;
  assign \new_[13298]_  = A166 & \new_[13297]_ ;
  assign \new_[13299]_  = \new_[13298]_  & \new_[13293]_ ;
  assign \new_[13303]_  = A232 & ~A203;
  assign \new_[13304]_  = ~A201 & \new_[13303]_ ;
  assign \new_[13308]_  = A300 & A298;
  assign \new_[13309]_  = A234 & \new_[13308]_ ;
  assign \new_[13310]_  = \new_[13309]_  & \new_[13304]_ ;
  assign \new_[13314]_  = ~A167 & A168;
  assign \new_[13315]_  = A170 & \new_[13314]_ ;
  assign \new_[13319]_  = A200 & ~A199;
  assign \new_[13320]_  = A166 & \new_[13319]_ ;
  assign \new_[13321]_  = \new_[13320]_  & \new_[13315]_ ;
  assign \new_[13325]_  = A232 & ~A203;
  assign \new_[13326]_  = ~A201 & \new_[13325]_ ;
  assign \new_[13330]_  = A267 & A265;
  assign \new_[13331]_  = A234 & \new_[13330]_ ;
  assign \new_[13332]_  = \new_[13331]_  & \new_[13326]_ ;
  assign \new_[13336]_  = ~A167 & A168;
  assign \new_[13337]_  = A170 & \new_[13336]_ ;
  assign \new_[13341]_  = A200 & ~A199;
  assign \new_[13342]_  = A166 & \new_[13341]_ ;
  assign \new_[13343]_  = \new_[13342]_  & \new_[13337]_ ;
  assign \new_[13347]_  = A232 & ~A203;
  assign \new_[13348]_  = ~A201 & \new_[13347]_ ;
  assign \new_[13352]_  = A267 & A266;
  assign \new_[13353]_  = A234 & \new_[13352]_ ;
  assign \new_[13354]_  = \new_[13353]_  & \new_[13348]_ ;
  assign \new_[13358]_  = ~A167 & A168;
  assign \new_[13359]_  = A170 & \new_[13358]_ ;
  assign \new_[13363]_  = A200 & ~A199;
  assign \new_[13364]_  = A166 & \new_[13363]_ ;
  assign \new_[13365]_  = \new_[13364]_  & \new_[13359]_ ;
  assign \new_[13369]_  = A233 & ~A203;
  assign \new_[13370]_  = ~A201 & \new_[13369]_ ;
  assign \new_[13374]_  = A300 & A299;
  assign \new_[13375]_  = A234 & \new_[13374]_ ;
  assign \new_[13376]_  = \new_[13375]_  & \new_[13370]_ ;
  assign \new_[13380]_  = ~A167 & A168;
  assign \new_[13381]_  = A170 & \new_[13380]_ ;
  assign \new_[13385]_  = A200 & ~A199;
  assign \new_[13386]_  = A166 & \new_[13385]_ ;
  assign \new_[13387]_  = \new_[13386]_  & \new_[13381]_ ;
  assign \new_[13391]_  = A233 & ~A203;
  assign \new_[13392]_  = ~A201 & \new_[13391]_ ;
  assign \new_[13396]_  = A300 & A298;
  assign \new_[13397]_  = A234 & \new_[13396]_ ;
  assign \new_[13398]_  = \new_[13397]_  & \new_[13392]_ ;
  assign \new_[13402]_  = ~A167 & A168;
  assign \new_[13403]_  = A170 & \new_[13402]_ ;
  assign \new_[13407]_  = A200 & ~A199;
  assign \new_[13408]_  = A166 & \new_[13407]_ ;
  assign \new_[13409]_  = \new_[13408]_  & \new_[13403]_ ;
  assign \new_[13413]_  = A233 & ~A203;
  assign \new_[13414]_  = ~A201 & \new_[13413]_ ;
  assign \new_[13418]_  = A267 & A265;
  assign \new_[13419]_  = A234 & \new_[13418]_ ;
  assign \new_[13420]_  = \new_[13419]_  & \new_[13414]_ ;
  assign \new_[13424]_  = ~A167 & A168;
  assign \new_[13425]_  = A170 & \new_[13424]_ ;
  assign \new_[13429]_  = A200 & ~A199;
  assign \new_[13430]_  = A166 & \new_[13429]_ ;
  assign \new_[13431]_  = \new_[13430]_  & \new_[13425]_ ;
  assign \new_[13435]_  = A233 & ~A203;
  assign \new_[13436]_  = ~A201 & \new_[13435]_ ;
  assign \new_[13440]_  = A267 & A266;
  assign \new_[13441]_  = A234 & \new_[13440]_ ;
  assign \new_[13442]_  = \new_[13441]_  & \new_[13436]_ ;
  assign \new_[13446]_  = ~A167 & A168;
  assign \new_[13447]_  = A170 & \new_[13446]_ ;
  assign \new_[13451]_  = ~A200 & A199;
  assign \new_[13452]_  = A166 & \new_[13451]_ ;
  assign \new_[13453]_  = \new_[13452]_  & \new_[13447]_ ;
  assign \new_[13457]_  = A232 & A202;
  assign \new_[13458]_  = ~A201 & \new_[13457]_ ;
  assign \new_[13462]_  = A300 & A299;
  assign \new_[13463]_  = A234 & \new_[13462]_ ;
  assign \new_[13464]_  = \new_[13463]_  & \new_[13458]_ ;
  assign \new_[13468]_  = ~A167 & A168;
  assign \new_[13469]_  = A170 & \new_[13468]_ ;
  assign \new_[13473]_  = ~A200 & A199;
  assign \new_[13474]_  = A166 & \new_[13473]_ ;
  assign \new_[13475]_  = \new_[13474]_  & \new_[13469]_ ;
  assign \new_[13479]_  = A232 & A202;
  assign \new_[13480]_  = ~A201 & \new_[13479]_ ;
  assign \new_[13484]_  = A300 & A298;
  assign \new_[13485]_  = A234 & \new_[13484]_ ;
  assign \new_[13486]_  = \new_[13485]_  & \new_[13480]_ ;
  assign \new_[13490]_  = ~A167 & A168;
  assign \new_[13491]_  = A170 & \new_[13490]_ ;
  assign \new_[13495]_  = ~A200 & A199;
  assign \new_[13496]_  = A166 & \new_[13495]_ ;
  assign \new_[13497]_  = \new_[13496]_  & \new_[13491]_ ;
  assign \new_[13501]_  = A232 & A202;
  assign \new_[13502]_  = ~A201 & \new_[13501]_ ;
  assign \new_[13506]_  = A267 & A265;
  assign \new_[13507]_  = A234 & \new_[13506]_ ;
  assign \new_[13508]_  = \new_[13507]_  & \new_[13502]_ ;
  assign \new_[13512]_  = ~A167 & A168;
  assign \new_[13513]_  = A170 & \new_[13512]_ ;
  assign \new_[13517]_  = ~A200 & A199;
  assign \new_[13518]_  = A166 & \new_[13517]_ ;
  assign \new_[13519]_  = \new_[13518]_  & \new_[13513]_ ;
  assign \new_[13523]_  = A232 & A202;
  assign \new_[13524]_  = ~A201 & \new_[13523]_ ;
  assign \new_[13528]_  = A267 & A266;
  assign \new_[13529]_  = A234 & \new_[13528]_ ;
  assign \new_[13530]_  = \new_[13529]_  & \new_[13524]_ ;
  assign \new_[13534]_  = ~A167 & A168;
  assign \new_[13535]_  = A170 & \new_[13534]_ ;
  assign \new_[13539]_  = ~A200 & A199;
  assign \new_[13540]_  = A166 & \new_[13539]_ ;
  assign \new_[13541]_  = \new_[13540]_  & \new_[13535]_ ;
  assign \new_[13545]_  = A233 & A202;
  assign \new_[13546]_  = ~A201 & \new_[13545]_ ;
  assign \new_[13550]_  = A300 & A299;
  assign \new_[13551]_  = A234 & \new_[13550]_ ;
  assign \new_[13552]_  = \new_[13551]_  & \new_[13546]_ ;
  assign \new_[13556]_  = ~A167 & A168;
  assign \new_[13557]_  = A170 & \new_[13556]_ ;
  assign \new_[13561]_  = ~A200 & A199;
  assign \new_[13562]_  = A166 & \new_[13561]_ ;
  assign \new_[13563]_  = \new_[13562]_  & \new_[13557]_ ;
  assign \new_[13567]_  = A233 & A202;
  assign \new_[13568]_  = ~A201 & \new_[13567]_ ;
  assign \new_[13572]_  = A300 & A298;
  assign \new_[13573]_  = A234 & \new_[13572]_ ;
  assign \new_[13574]_  = \new_[13573]_  & \new_[13568]_ ;
  assign \new_[13578]_  = ~A167 & A168;
  assign \new_[13579]_  = A170 & \new_[13578]_ ;
  assign \new_[13583]_  = ~A200 & A199;
  assign \new_[13584]_  = A166 & \new_[13583]_ ;
  assign \new_[13585]_  = \new_[13584]_  & \new_[13579]_ ;
  assign \new_[13589]_  = A233 & A202;
  assign \new_[13590]_  = ~A201 & \new_[13589]_ ;
  assign \new_[13594]_  = A267 & A265;
  assign \new_[13595]_  = A234 & \new_[13594]_ ;
  assign \new_[13596]_  = \new_[13595]_  & \new_[13590]_ ;
  assign \new_[13600]_  = ~A167 & A168;
  assign \new_[13601]_  = A170 & \new_[13600]_ ;
  assign \new_[13605]_  = ~A200 & A199;
  assign \new_[13606]_  = A166 & \new_[13605]_ ;
  assign \new_[13607]_  = \new_[13606]_  & \new_[13601]_ ;
  assign \new_[13611]_  = A233 & A202;
  assign \new_[13612]_  = ~A201 & \new_[13611]_ ;
  assign \new_[13616]_  = A267 & A266;
  assign \new_[13617]_  = A234 & \new_[13616]_ ;
  assign \new_[13618]_  = \new_[13617]_  & \new_[13612]_ ;
  assign \new_[13622]_  = ~A167 & A168;
  assign \new_[13623]_  = A170 & \new_[13622]_ ;
  assign \new_[13627]_  = ~A200 & A199;
  assign \new_[13628]_  = A166 & \new_[13627]_ ;
  assign \new_[13629]_  = \new_[13628]_  & \new_[13623]_ ;
  assign \new_[13633]_  = A232 & ~A203;
  assign \new_[13634]_  = ~A201 & \new_[13633]_ ;
  assign \new_[13638]_  = A300 & A299;
  assign \new_[13639]_  = A234 & \new_[13638]_ ;
  assign \new_[13640]_  = \new_[13639]_  & \new_[13634]_ ;
  assign \new_[13644]_  = ~A167 & A168;
  assign \new_[13645]_  = A170 & \new_[13644]_ ;
  assign \new_[13649]_  = ~A200 & A199;
  assign \new_[13650]_  = A166 & \new_[13649]_ ;
  assign \new_[13651]_  = \new_[13650]_  & \new_[13645]_ ;
  assign \new_[13655]_  = A232 & ~A203;
  assign \new_[13656]_  = ~A201 & \new_[13655]_ ;
  assign \new_[13660]_  = A300 & A298;
  assign \new_[13661]_  = A234 & \new_[13660]_ ;
  assign \new_[13662]_  = \new_[13661]_  & \new_[13656]_ ;
  assign \new_[13666]_  = ~A167 & A168;
  assign \new_[13667]_  = A170 & \new_[13666]_ ;
  assign \new_[13671]_  = ~A200 & A199;
  assign \new_[13672]_  = A166 & \new_[13671]_ ;
  assign \new_[13673]_  = \new_[13672]_  & \new_[13667]_ ;
  assign \new_[13677]_  = A232 & ~A203;
  assign \new_[13678]_  = ~A201 & \new_[13677]_ ;
  assign \new_[13682]_  = A267 & A265;
  assign \new_[13683]_  = A234 & \new_[13682]_ ;
  assign \new_[13684]_  = \new_[13683]_  & \new_[13678]_ ;
  assign \new_[13688]_  = ~A167 & A168;
  assign \new_[13689]_  = A170 & \new_[13688]_ ;
  assign \new_[13693]_  = ~A200 & A199;
  assign \new_[13694]_  = A166 & \new_[13693]_ ;
  assign \new_[13695]_  = \new_[13694]_  & \new_[13689]_ ;
  assign \new_[13699]_  = A232 & ~A203;
  assign \new_[13700]_  = ~A201 & \new_[13699]_ ;
  assign \new_[13704]_  = A267 & A266;
  assign \new_[13705]_  = A234 & \new_[13704]_ ;
  assign \new_[13706]_  = \new_[13705]_  & \new_[13700]_ ;
  assign \new_[13710]_  = ~A167 & A168;
  assign \new_[13711]_  = A170 & \new_[13710]_ ;
  assign \new_[13715]_  = ~A200 & A199;
  assign \new_[13716]_  = A166 & \new_[13715]_ ;
  assign \new_[13717]_  = \new_[13716]_  & \new_[13711]_ ;
  assign \new_[13721]_  = A233 & ~A203;
  assign \new_[13722]_  = ~A201 & \new_[13721]_ ;
  assign \new_[13726]_  = A300 & A299;
  assign \new_[13727]_  = A234 & \new_[13726]_ ;
  assign \new_[13728]_  = \new_[13727]_  & \new_[13722]_ ;
  assign \new_[13732]_  = ~A167 & A168;
  assign \new_[13733]_  = A170 & \new_[13732]_ ;
  assign \new_[13737]_  = ~A200 & A199;
  assign \new_[13738]_  = A166 & \new_[13737]_ ;
  assign \new_[13739]_  = \new_[13738]_  & \new_[13733]_ ;
  assign \new_[13743]_  = A233 & ~A203;
  assign \new_[13744]_  = ~A201 & \new_[13743]_ ;
  assign \new_[13748]_  = A300 & A298;
  assign \new_[13749]_  = A234 & \new_[13748]_ ;
  assign \new_[13750]_  = \new_[13749]_  & \new_[13744]_ ;
  assign \new_[13754]_  = ~A167 & A168;
  assign \new_[13755]_  = A170 & \new_[13754]_ ;
  assign \new_[13759]_  = ~A200 & A199;
  assign \new_[13760]_  = A166 & \new_[13759]_ ;
  assign \new_[13761]_  = \new_[13760]_  & \new_[13755]_ ;
  assign \new_[13765]_  = A233 & ~A203;
  assign \new_[13766]_  = ~A201 & \new_[13765]_ ;
  assign \new_[13770]_  = A267 & A265;
  assign \new_[13771]_  = A234 & \new_[13770]_ ;
  assign \new_[13772]_  = \new_[13771]_  & \new_[13766]_ ;
  assign \new_[13776]_  = ~A167 & A168;
  assign \new_[13777]_  = A170 & \new_[13776]_ ;
  assign \new_[13781]_  = ~A200 & A199;
  assign \new_[13782]_  = A166 & \new_[13781]_ ;
  assign \new_[13783]_  = \new_[13782]_  & \new_[13777]_ ;
  assign \new_[13787]_  = A233 & ~A203;
  assign \new_[13788]_  = ~A201 & \new_[13787]_ ;
  assign \new_[13792]_  = A267 & A266;
  assign \new_[13793]_  = A234 & \new_[13792]_ ;
  assign \new_[13794]_  = \new_[13793]_  & \new_[13788]_ ;
  assign \new_[13798]_  = ~A167 & A168;
  assign \new_[13799]_  = A169 & \new_[13798]_ ;
  assign \new_[13803]_  = A200 & A199;
  assign \new_[13804]_  = A166 & \new_[13803]_ ;
  assign \new_[13805]_  = \new_[13804]_  & \new_[13799]_ ;
  assign \new_[13809]_  = A232 & ~A202;
  assign \new_[13810]_  = ~A201 & \new_[13809]_ ;
  assign \new_[13814]_  = A300 & A299;
  assign \new_[13815]_  = A234 & \new_[13814]_ ;
  assign \new_[13816]_  = \new_[13815]_  & \new_[13810]_ ;
  assign \new_[13820]_  = ~A167 & A168;
  assign \new_[13821]_  = A169 & \new_[13820]_ ;
  assign \new_[13825]_  = A200 & A199;
  assign \new_[13826]_  = A166 & \new_[13825]_ ;
  assign \new_[13827]_  = \new_[13826]_  & \new_[13821]_ ;
  assign \new_[13831]_  = A232 & ~A202;
  assign \new_[13832]_  = ~A201 & \new_[13831]_ ;
  assign \new_[13836]_  = A300 & A298;
  assign \new_[13837]_  = A234 & \new_[13836]_ ;
  assign \new_[13838]_  = \new_[13837]_  & \new_[13832]_ ;
  assign \new_[13842]_  = ~A167 & A168;
  assign \new_[13843]_  = A169 & \new_[13842]_ ;
  assign \new_[13847]_  = A200 & A199;
  assign \new_[13848]_  = A166 & \new_[13847]_ ;
  assign \new_[13849]_  = \new_[13848]_  & \new_[13843]_ ;
  assign \new_[13853]_  = A232 & ~A202;
  assign \new_[13854]_  = ~A201 & \new_[13853]_ ;
  assign \new_[13858]_  = A267 & A265;
  assign \new_[13859]_  = A234 & \new_[13858]_ ;
  assign \new_[13860]_  = \new_[13859]_  & \new_[13854]_ ;
  assign \new_[13864]_  = ~A167 & A168;
  assign \new_[13865]_  = A169 & \new_[13864]_ ;
  assign \new_[13869]_  = A200 & A199;
  assign \new_[13870]_  = A166 & \new_[13869]_ ;
  assign \new_[13871]_  = \new_[13870]_  & \new_[13865]_ ;
  assign \new_[13875]_  = A232 & ~A202;
  assign \new_[13876]_  = ~A201 & \new_[13875]_ ;
  assign \new_[13880]_  = A267 & A266;
  assign \new_[13881]_  = A234 & \new_[13880]_ ;
  assign \new_[13882]_  = \new_[13881]_  & \new_[13876]_ ;
  assign \new_[13886]_  = ~A167 & A168;
  assign \new_[13887]_  = A169 & \new_[13886]_ ;
  assign \new_[13891]_  = A200 & A199;
  assign \new_[13892]_  = A166 & \new_[13891]_ ;
  assign \new_[13893]_  = \new_[13892]_  & \new_[13887]_ ;
  assign \new_[13897]_  = A233 & ~A202;
  assign \new_[13898]_  = ~A201 & \new_[13897]_ ;
  assign \new_[13902]_  = A300 & A299;
  assign \new_[13903]_  = A234 & \new_[13902]_ ;
  assign \new_[13904]_  = \new_[13903]_  & \new_[13898]_ ;
  assign \new_[13908]_  = ~A167 & A168;
  assign \new_[13909]_  = A169 & \new_[13908]_ ;
  assign \new_[13913]_  = A200 & A199;
  assign \new_[13914]_  = A166 & \new_[13913]_ ;
  assign \new_[13915]_  = \new_[13914]_  & \new_[13909]_ ;
  assign \new_[13919]_  = A233 & ~A202;
  assign \new_[13920]_  = ~A201 & \new_[13919]_ ;
  assign \new_[13924]_  = A300 & A298;
  assign \new_[13925]_  = A234 & \new_[13924]_ ;
  assign \new_[13926]_  = \new_[13925]_  & \new_[13920]_ ;
  assign \new_[13930]_  = ~A167 & A168;
  assign \new_[13931]_  = A169 & \new_[13930]_ ;
  assign \new_[13935]_  = A200 & A199;
  assign \new_[13936]_  = A166 & \new_[13935]_ ;
  assign \new_[13937]_  = \new_[13936]_  & \new_[13931]_ ;
  assign \new_[13941]_  = A233 & ~A202;
  assign \new_[13942]_  = ~A201 & \new_[13941]_ ;
  assign \new_[13946]_  = A267 & A265;
  assign \new_[13947]_  = A234 & \new_[13946]_ ;
  assign \new_[13948]_  = \new_[13947]_  & \new_[13942]_ ;
  assign \new_[13952]_  = ~A167 & A168;
  assign \new_[13953]_  = A169 & \new_[13952]_ ;
  assign \new_[13957]_  = A200 & A199;
  assign \new_[13958]_  = A166 & \new_[13957]_ ;
  assign \new_[13959]_  = \new_[13958]_  & \new_[13953]_ ;
  assign \new_[13963]_  = A233 & ~A202;
  assign \new_[13964]_  = ~A201 & \new_[13963]_ ;
  assign \new_[13968]_  = A267 & A266;
  assign \new_[13969]_  = A234 & \new_[13968]_ ;
  assign \new_[13970]_  = \new_[13969]_  & \new_[13964]_ ;
  assign \new_[13974]_  = ~A167 & A168;
  assign \new_[13975]_  = A169 & \new_[13974]_ ;
  assign \new_[13979]_  = A200 & A199;
  assign \new_[13980]_  = A166 & \new_[13979]_ ;
  assign \new_[13981]_  = \new_[13980]_  & \new_[13975]_ ;
  assign \new_[13985]_  = A232 & A203;
  assign \new_[13986]_  = ~A201 & \new_[13985]_ ;
  assign \new_[13990]_  = A300 & A299;
  assign \new_[13991]_  = A234 & \new_[13990]_ ;
  assign \new_[13992]_  = \new_[13991]_  & \new_[13986]_ ;
  assign \new_[13996]_  = ~A167 & A168;
  assign \new_[13997]_  = A169 & \new_[13996]_ ;
  assign \new_[14001]_  = A200 & A199;
  assign \new_[14002]_  = A166 & \new_[14001]_ ;
  assign \new_[14003]_  = \new_[14002]_  & \new_[13997]_ ;
  assign \new_[14007]_  = A232 & A203;
  assign \new_[14008]_  = ~A201 & \new_[14007]_ ;
  assign \new_[14012]_  = A300 & A298;
  assign \new_[14013]_  = A234 & \new_[14012]_ ;
  assign \new_[14014]_  = \new_[14013]_  & \new_[14008]_ ;
  assign \new_[14018]_  = ~A167 & A168;
  assign \new_[14019]_  = A169 & \new_[14018]_ ;
  assign \new_[14023]_  = A200 & A199;
  assign \new_[14024]_  = A166 & \new_[14023]_ ;
  assign \new_[14025]_  = \new_[14024]_  & \new_[14019]_ ;
  assign \new_[14029]_  = A232 & A203;
  assign \new_[14030]_  = ~A201 & \new_[14029]_ ;
  assign \new_[14034]_  = A267 & A265;
  assign \new_[14035]_  = A234 & \new_[14034]_ ;
  assign \new_[14036]_  = \new_[14035]_  & \new_[14030]_ ;
  assign \new_[14040]_  = ~A167 & A168;
  assign \new_[14041]_  = A169 & \new_[14040]_ ;
  assign \new_[14045]_  = A200 & A199;
  assign \new_[14046]_  = A166 & \new_[14045]_ ;
  assign \new_[14047]_  = \new_[14046]_  & \new_[14041]_ ;
  assign \new_[14051]_  = A232 & A203;
  assign \new_[14052]_  = ~A201 & \new_[14051]_ ;
  assign \new_[14056]_  = A267 & A266;
  assign \new_[14057]_  = A234 & \new_[14056]_ ;
  assign \new_[14058]_  = \new_[14057]_  & \new_[14052]_ ;
  assign \new_[14062]_  = ~A167 & A168;
  assign \new_[14063]_  = A169 & \new_[14062]_ ;
  assign \new_[14067]_  = A200 & A199;
  assign \new_[14068]_  = A166 & \new_[14067]_ ;
  assign \new_[14069]_  = \new_[14068]_  & \new_[14063]_ ;
  assign \new_[14073]_  = A233 & A203;
  assign \new_[14074]_  = ~A201 & \new_[14073]_ ;
  assign \new_[14078]_  = A300 & A299;
  assign \new_[14079]_  = A234 & \new_[14078]_ ;
  assign \new_[14080]_  = \new_[14079]_  & \new_[14074]_ ;
  assign \new_[14084]_  = ~A167 & A168;
  assign \new_[14085]_  = A169 & \new_[14084]_ ;
  assign \new_[14089]_  = A200 & A199;
  assign \new_[14090]_  = A166 & \new_[14089]_ ;
  assign \new_[14091]_  = \new_[14090]_  & \new_[14085]_ ;
  assign \new_[14095]_  = A233 & A203;
  assign \new_[14096]_  = ~A201 & \new_[14095]_ ;
  assign \new_[14100]_  = A300 & A298;
  assign \new_[14101]_  = A234 & \new_[14100]_ ;
  assign \new_[14102]_  = \new_[14101]_  & \new_[14096]_ ;
  assign \new_[14106]_  = ~A167 & A168;
  assign \new_[14107]_  = A169 & \new_[14106]_ ;
  assign \new_[14111]_  = A200 & A199;
  assign \new_[14112]_  = A166 & \new_[14111]_ ;
  assign \new_[14113]_  = \new_[14112]_  & \new_[14107]_ ;
  assign \new_[14117]_  = A233 & A203;
  assign \new_[14118]_  = ~A201 & \new_[14117]_ ;
  assign \new_[14122]_  = A267 & A265;
  assign \new_[14123]_  = A234 & \new_[14122]_ ;
  assign \new_[14124]_  = \new_[14123]_  & \new_[14118]_ ;
  assign \new_[14128]_  = ~A167 & A168;
  assign \new_[14129]_  = A169 & \new_[14128]_ ;
  assign \new_[14133]_  = A200 & A199;
  assign \new_[14134]_  = A166 & \new_[14133]_ ;
  assign \new_[14135]_  = \new_[14134]_  & \new_[14129]_ ;
  assign \new_[14139]_  = A233 & A203;
  assign \new_[14140]_  = ~A201 & \new_[14139]_ ;
  assign \new_[14144]_  = A267 & A266;
  assign \new_[14145]_  = A234 & \new_[14144]_ ;
  assign \new_[14146]_  = \new_[14145]_  & \new_[14140]_ ;
  assign \new_[14150]_  = ~A167 & A168;
  assign \new_[14151]_  = A169 & \new_[14150]_ ;
  assign \new_[14155]_  = A200 & ~A199;
  assign \new_[14156]_  = A166 & \new_[14155]_ ;
  assign \new_[14157]_  = \new_[14156]_  & \new_[14151]_ ;
  assign \new_[14161]_  = A232 & A202;
  assign \new_[14162]_  = ~A201 & \new_[14161]_ ;
  assign \new_[14166]_  = A300 & A299;
  assign \new_[14167]_  = A234 & \new_[14166]_ ;
  assign \new_[14168]_  = \new_[14167]_  & \new_[14162]_ ;
  assign \new_[14172]_  = ~A167 & A168;
  assign \new_[14173]_  = A169 & \new_[14172]_ ;
  assign \new_[14177]_  = A200 & ~A199;
  assign \new_[14178]_  = A166 & \new_[14177]_ ;
  assign \new_[14179]_  = \new_[14178]_  & \new_[14173]_ ;
  assign \new_[14183]_  = A232 & A202;
  assign \new_[14184]_  = ~A201 & \new_[14183]_ ;
  assign \new_[14188]_  = A300 & A298;
  assign \new_[14189]_  = A234 & \new_[14188]_ ;
  assign \new_[14190]_  = \new_[14189]_  & \new_[14184]_ ;
  assign \new_[14194]_  = ~A167 & A168;
  assign \new_[14195]_  = A169 & \new_[14194]_ ;
  assign \new_[14199]_  = A200 & ~A199;
  assign \new_[14200]_  = A166 & \new_[14199]_ ;
  assign \new_[14201]_  = \new_[14200]_  & \new_[14195]_ ;
  assign \new_[14205]_  = A232 & A202;
  assign \new_[14206]_  = ~A201 & \new_[14205]_ ;
  assign \new_[14210]_  = A267 & A265;
  assign \new_[14211]_  = A234 & \new_[14210]_ ;
  assign \new_[14212]_  = \new_[14211]_  & \new_[14206]_ ;
  assign \new_[14216]_  = ~A167 & A168;
  assign \new_[14217]_  = A169 & \new_[14216]_ ;
  assign \new_[14221]_  = A200 & ~A199;
  assign \new_[14222]_  = A166 & \new_[14221]_ ;
  assign \new_[14223]_  = \new_[14222]_  & \new_[14217]_ ;
  assign \new_[14227]_  = A232 & A202;
  assign \new_[14228]_  = ~A201 & \new_[14227]_ ;
  assign \new_[14232]_  = A267 & A266;
  assign \new_[14233]_  = A234 & \new_[14232]_ ;
  assign \new_[14234]_  = \new_[14233]_  & \new_[14228]_ ;
  assign \new_[14238]_  = ~A167 & A168;
  assign \new_[14239]_  = A169 & \new_[14238]_ ;
  assign \new_[14243]_  = A200 & ~A199;
  assign \new_[14244]_  = A166 & \new_[14243]_ ;
  assign \new_[14245]_  = \new_[14244]_  & \new_[14239]_ ;
  assign \new_[14249]_  = A233 & A202;
  assign \new_[14250]_  = ~A201 & \new_[14249]_ ;
  assign \new_[14254]_  = A300 & A299;
  assign \new_[14255]_  = A234 & \new_[14254]_ ;
  assign \new_[14256]_  = \new_[14255]_  & \new_[14250]_ ;
  assign \new_[14260]_  = ~A167 & A168;
  assign \new_[14261]_  = A169 & \new_[14260]_ ;
  assign \new_[14265]_  = A200 & ~A199;
  assign \new_[14266]_  = A166 & \new_[14265]_ ;
  assign \new_[14267]_  = \new_[14266]_  & \new_[14261]_ ;
  assign \new_[14271]_  = A233 & A202;
  assign \new_[14272]_  = ~A201 & \new_[14271]_ ;
  assign \new_[14276]_  = A300 & A298;
  assign \new_[14277]_  = A234 & \new_[14276]_ ;
  assign \new_[14278]_  = \new_[14277]_  & \new_[14272]_ ;
  assign \new_[14282]_  = ~A167 & A168;
  assign \new_[14283]_  = A169 & \new_[14282]_ ;
  assign \new_[14287]_  = A200 & ~A199;
  assign \new_[14288]_  = A166 & \new_[14287]_ ;
  assign \new_[14289]_  = \new_[14288]_  & \new_[14283]_ ;
  assign \new_[14293]_  = A233 & A202;
  assign \new_[14294]_  = ~A201 & \new_[14293]_ ;
  assign \new_[14298]_  = A267 & A265;
  assign \new_[14299]_  = A234 & \new_[14298]_ ;
  assign \new_[14300]_  = \new_[14299]_  & \new_[14294]_ ;
  assign \new_[14304]_  = ~A167 & A168;
  assign \new_[14305]_  = A169 & \new_[14304]_ ;
  assign \new_[14309]_  = A200 & ~A199;
  assign \new_[14310]_  = A166 & \new_[14309]_ ;
  assign \new_[14311]_  = \new_[14310]_  & \new_[14305]_ ;
  assign \new_[14315]_  = A233 & A202;
  assign \new_[14316]_  = ~A201 & \new_[14315]_ ;
  assign \new_[14320]_  = A267 & A266;
  assign \new_[14321]_  = A234 & \new_[14320]_ ;
  assign \new_[14322]_  = \new_[14321]_  & \new_[14316]_ ;
  assign \new_[14326]_  = ~A167 & A168;
  assign \new_[14327]_  = A169 & \new_[14326]_ ;
  assign \new_[14331]_  = A200 & ~A199;
  assign \new_[14332]_  = A166 & \new_[14331]_ ;
  assign \new_[14333]_  = \new_[14332]_  & \new_[14327]_ ;
  assign \new_[14337]_  = A232 & ~A203;
  assign \new_[14338]_  = ~A201 & \new_[14337]_ ;
  assign \new_[14342]_  = A300 & A299;
  assign \new_[14343]_  = A234 & \new_[14342]_ ;
  assign \new_[14344]_  = \new_[14343]_  & \new_[14338]_ ;
  assign \new_[14348]_  = ~A167 & A168;
  assign \new_[14349]_  = A169 & \new_[14348]_ ;
  assign \new_[14353]_  = A200 & ~A199;
  assign \new_[14354]_  = A166 & \new_[14353]_ ;
  assign \new_[14355]_  = \new_[14354]_  & \new_[14349]_ ;
  assign \new_[14359]_  = A232 & ~A203;
  assign \new_[14360]_  = ~A201 & \new_[14359]_ ;
  assign \new_[14364]_  = A300 & A298;
  assign \new_[14365]_  = A234 & \new_[14364]_ ;
  assign \new_[14366]_  = \new_[14365]_  & \new_[14360]_ ;
  assign \new_[14370]_  = ~A167 & A168;
  assign \new_[14371]_  = A169 & \new_[14370]_ ;
  assign \new_[14375]_  = A200 & ~A199;
  assign \new_[14376]_  = A166 & \new_[14375]_ ;
  assign \new_[14377]_  = \new_[14376]_  & \new_[14371]_ ;
  assign \new_[14381]_  = A232 & ~A203;
  assign \new_[14382]_  = ~A201 & \new_[14381]_ ;
  assign \new_[14386]_  = A267 & A265;
  assign \new_[14387]_  = A234 & \new_[14386]_ ;
  assign \new_[14388]_  = \new_[14387]_  & \new_[14382]_ ;
  assign \new_[14392]_  = ~A167 & A168;
  assign \new_[14393]_  = A169 & \new_[14392]_ ;
  assign \new_[14397]_  = A200 & ~A199;
  assign \new_[14398]_  = A166 & \new_[14397]_ ;
  assign \new_[14399]_  = \new_[14398]_  & \new_[14393]_ ;
  assign \new_[14403]_  = A232 & ~A203;
  assign \new_[14404]_  = ~A201 & \new_[14403]_ ;
  assign \new_[14408]_  = A267 & A266;
  assign \new_[14409]_  = A234 & \new_[14408]_ ;
  assign \new_[14410]_  = \new_[14409]_  & \new_[14404]_ ;
  assign \new_[14414]_  = ~A167 & A168;
  assign \new_[14415]_  = A169 & \new_[14414]_ ;
  assign \new_[14419]_  = A200 & ~A199;
  assign \new_[14420]_  = A166 & \new_[14419]_ ;
  assign \new_[14421]_  = \new_[14420]_  & \new_[14415]_ ;
  assign \new_[14425]_  = A233 & ~A203;
  assign \new_[14426]_  = ~A201 & \new_[14425]_ ;
  assign \new_[14430]_  = A300 & A299;
  assign \new_[14431]_  = A234 & \new_[14430]_ ;
  assign \new_[14432]_  = \new_[14431]_  & \new_[14426]_ ;
  assign \new_[14436]_  = ~A167 & A168;
  assign \new_[14437]_  = A169 & \new_[14436]_ ;
  assign \new_[14441]_  = A200 & ~A199;
  assign \new_[14442]_  = A166 & \new_[14441]_ ;
  assign \new_[14443]_  = \new_[14442]_  & \new_[14437]_ ;
  assign \new_[14447]_  = A233 & ~A203;
  assign \new_[14448]_  = ~A201 & \new_[14447]_ ;
  assign \new_[14452]_  = A300 & A298;
  assign \new_[14453]_  = A234 & \new_[14452]_ ;
  assign \new_[14454]_  = \new_[14453]_  & \new_[14448]_ ;
  assign \new_[14458]_  = ~A167 & A168;
  assign \new_[14459]_  = A169 & \new_[14458]_ ;
  assign \new_[14463]_  = A200 & ~A199;
  assign \new_[14464]_  = A166 & \new_[14463]_ ;
  assign \new_[14465]_  = \new_[14464]_  & \new_[14459]_ ;
  assign \new_[14469]_  = A233 & ~A203;
  assign \new_[14470]_  = ~A201 & \new_[14469]_ ;
  assign \new_[14474]_  = A267 & A265;
  assign \new_[14475]_  = A234 & \new_[14474]_ ;
  assign \new_[14476]_  = \new_[14475]_  & \new_[14470]_ ;
  assign \new_[14480]_  = ~A167 & A168;
  assign \new_[14481]_  = A169 & \new_[14480]_ ;
  assign \new_[14485]_  = A200 & ~A199;
  assign \new_[14486]_  = A166 & \new_[14485]_ ;
  assign \new_[14487]_  = \new_[14486]_  & \new_[14481]_ ;
  assign \new_[14491]_  = A233 & ~A203;
  assign \new_[14492]_  = ~A201 & \new_[14491]_ ;
  assign \new_[14496]_  = A267 & A266;
  assign \new_[14497]_  = A234 & \new_[14496]_ ;
  assign \new_[14498]_  = \new_[14497]_  & \new_[14492]_ ;
  assign \new_[14502]_  = ~A167 & A168;
  assign \new_[14503]_  = A169 & \new_[14502]_ ;
  assign \new_[14507]_  = ~A200 & A199;
  assign \new_[14508]_  = A166 & \new_[14507]_ ;
  assign \new_[14509]_  = \new_[14508]_  & \new_[14503]_ ;
  assign \new_[14513]_  = A232 & A202;
  assign \new_[14514]_  = ~A201 & \new_[14513]_ ;
  assign \new_[14518]_  = A300 & A299;
  assign \new_[14519]_  = A234 & \new_[14518]_ ;
  assign \new_[14520]_  = \new_[14519]_  & \new_[14514]_ ;
  assign \new_[14524]_  = ~A167 & A168;
  assign \new_[14525]_  = A169 & \new_[14524]_ ;
  assign \new_[14529]_  = ~A200 & A199;
  assign \new_[14530]_  = A166 & \new_[14529]_ ;
  assign \new_[14531]_  = \new_[14530]_  & \new_[14525]_ ;
  assign \new_[14535]_  = A232 & A202;
  assign \new_[14536]_  = ~A201 & \new_[14535]_ ;
  assign \new_[14540]_  = A300 & A298;
  assign \new_[14541]_  = A234 & \new_[14540]_ ;
  assign \new_[14542]_  = \new_[14541]_  & \new_[14536]_ ;
  assign \new_[14546]_  = ~A167 & A168;
  assign \new_[14547]_  = A169 & \new_[14546]_ ;
  assign \new_[14551]_  = ~A200 & A199;
  assign \new_[14552]_  = A166 & \new_[14551]_ ;
  assign \new_[14553]_  = \new_[14552]_  & \new_[14547]_ ;
  assign \new_[14557]_  = A232 & A202;
  assign \new_[14558]_  = ~A201 & \new_[14557]_ ;
  assign \new_[14562]_  = A267 & A265;
  assign \new_[14563]_  = A234 & \new_[14562]_ ;
  assign \new_[14564]_  = \new_[14563]_  & \new_[14558]_ ;
  assign \new_[14568]_  = ~A167 & A168;
  assign \new_[14569]_  = A169 & \new_[14568]_ ;
  assign \new_[14573]_  = ~A200 & A199;
  assign \new_[14574]_  = A166 & \new_[14573]_ ;
  assign \new_[14575]_  = \new_[14574]_  & \new_[14569]_ ;
  assign \new_[14579]_  = A232 & A202;
  assign \new_[14580]_  = ~A201 & \new_[14579]_ ;
  assign \new_[14584]_  = A267 & A266;
  assign \new_[14585]_  = A234 & \new_[14584]_ ;
  assign \new_[14586]_  = \new_[14585]_  & \new_[14580]_ ;
  assign \new_[14590]_  = ~A167 & A168;
  assign \new_[14591]_  = A169 & \new_[14590]_ ;
  assign \new_[14595]_  = ~A200 & A199;
  assign \new_[14596]_  = A166 & \new_[14595]_ ;
  assign \new_[14597]_  = \new_[14596]_  & \new_[14591]_ ;
  assign \new_[14601]_  = A233 & A202;
  assign \new_[14602]_  = ~A201 & \new_[14601]_ ;
  assign \new_[14606]_  = A300 & A299;
  assign \new_[14607]_  = A234 & \new_[14606]_ ;
  assign \new_[14608]_  = \new_[14607]_  & \new_[14602]_ ;
  assign \new_[14612]_  = ~A167 & A168;
  assign \new_[14613]_  = A169 & \new_[14612]_ ;
  assign \new_[14617]_  = ~A200 & A199;
  assign \new_[14618]_  = A166 & \new_[14617]_ ;
  assign \new_[14619]_  = \new_[14618]_  & \new_[14613]_ ;
  assign \new_[14623]_  = A233 & A202;
  assign \new_[14624]_  = ~A201 & \new_[14623]_ ;
  assign \new_[14628]_  = A300 & A298;
  assign \new_[14629]_  = A234 & \new_[14628]_ ;
  assign \new_[14630]_  = \new_[14629]_  & \new_[14624]_ ;
  assign \new_[14634]_  = ~A167 & A168;
  assign \new_[14635]_  = A169 & \new_[14634]_ ;
  assign \new_[14639]_  = ~A200 & A199;
  assign \new_[14640]_  = A166 & \new_[14639]_ ;
  assign \new_[14641]_  = \new_[14640]_  & \new_[14635]_ ;
  assign \new_[14645]_  = A233 & A202;
  assign \new_[14646]_  = ~A201 & \new_[14645]_ ;
  assign \new_[14650]_  = A267 & A265;
  assign \new_[14651]_  = A234 & \new_[14650]_ ;
  assign \new_[14652]_  = \new_[14651]_  & \new_[14646]_ ;
  assign \new_[14656]_  = ~A167 & A168;
  assign \new_[14657]_  = A169 & \new_[14656]_ ;
  assign \new_[14661]_  = ~A200 & A199;
  assign \new_[14662]_  = A166 & \new_[14661]_ ;
  assign \new_[14663]_  = \new_[14662]_  & \new_[14657]_ ;
  assign \new_[14667]_  = A233 & A202;
  assign \new_[14668]_  = ~A201 & \new_[14667]_ ;
  assign \new_[14672]_  = A267 & A266;
  assign \new_[14673]_  = A234 & \new_[14672]_ ;
  assign \new_[14674]_  = \new_[14673]_  & \new_[14668]_ ;
  assign \new_[14678]_  = ~A167 & A168;
  assign \new_[14679]_  = A169 & \new_[14678]_ ;
  assign \new_[14683]_  = ~A200 & A199;
  assign \new_[14684]_  = A166 & \new_[14683]_ ;
  assign \new_[14685]_  = \new_[14684]_  & \new_[14679]_ ;
  assign \new_[14689]_  = A232 & ~A203;
  assign \new_[14690]_  = ~A201 & \new_[14689]_ ;
  assign \new_[14694]_  = A300 & A299;
  assign \new_[14695]_  = A234 & \new_[14694]_ ;
  assign \new_[14696]_  = \new_[14695]_  & \new_[14690]_ ;
  assign \new_[14700]_  = ~A167 & A168;
  assign \new_[14701]_  = A169 & \new_[14700]_ ;
  assign \new_[14705]_  = ~A200 & A199;
  assign \new_[14706]_  = A166 & \new_[14705]_ ;
  assign \new_[14707]_  = \new_[14706]_  & \new_[14701]_ ;
  assign \new_[14711]_  = A232 & ~A203;
  assign \new_[14712]_  = ~A201 & \new_[14711]_ ;
  assign \new_[14716]_  = A300 & A298;
  assign \new_[14717]_  = A234 & \new_[14716]_ ;
  assign \new_[14718]_  = \new_[14717]_  & \new_[14712]_ ;
  assign \new_[14722]_  = ~A167 & A168;
  assign \new_[14723]_  = A169 & \new_[14722]_ ;
  assign \new_[14727]_  = ~A200 & A199;
  assign \new_[14728]_  = A166 & \new_[14727]_ ;
  assign \new_[14729]_  = \new_[14728]_  & \new_[14723]_ ;
  assign \new_[14733]_  = A232 & ~A203;
  assign \new_[14734]_  = ~A201 & \new_[14733]_ ;
  assign \new_[14738]_  = A267 & A265;
  assign \new_[14739]_  = A234 & \new_[14738]_ ;
  assign \new_[14740]_  = \new_[14739]_  & \new_[14734]_ ;
  assign \new_[14744]_  = ~A167 & A168;
  assign \new_[14745]_  = A169 & \new_[14744]_ ;
  assign \new_[14749]_  = ~A200 & A199;
  assign \new_[14750]_  = A166 & \new_[14749]_ ;
  assign \new_[14751]_  = \new_[14750]_  & \new_[14745]_ ;
  assign \new_[14755]_  = A232 & ~A203;
  assign \new_[14756]_  = ~A201 & \new_[14755]_ ;
  assign \new_[14760]_  = A267 & A266;
  assign \new_[14761]_  = A234 & \new_[14760]_ ;
  assign \new_[14762]_  = \new_[14761]_  & \new_[14756]_ ;
  assign \new_[14766]_  = ~A167 & A168;
  assign \new_[14767]_  = A169 & \new_[14766]_ ;
  assign \new_[14771]_  = ~A200 & A199;
  assign \new_[14772]_  = A166 & \new_[14771]_ ;
  assign \new_[14773]_  = \new_[14772]_  & \new_[14767]_ ;
  assign \new_[14777]_  = A233 & ~A203;
  assign \new_[14778]_  = ~A201 & \new_[14777]_ ;
  assign \new_[14782]_  = A300 & A299;
  assign \new_[14783]_  = A234 & \new_[14782]_ ;
  assign \new_[14784]_  = \new_[14783]_  & \new_[14778]_ ;
  assign \new_[14788]_  = ~A167 & A168;
  assign \new_[14789]_  = A169 & \new_[14788]_ ;
  assign \new_[14793]_  = ~A200 & A199;
  assign \new_[14794]_  = A166 & \new_[14793]_ ;
  assign \new_[14795]_  = \new_[14794]_  & \new_[14789]_ ;
  assign \new_[14799]_  = A233 & ~A203;
  assign \new_[14800]_  = ~A201 & \new_[14799]_ ;
  assign \new_[14804]_  = A300 & A298;
  assign \new_[14805]_  = A234 & \new_[14804]_ ;
  assign \new_[14806]_  = \new_[14805]_  & \new_[14800]_ ;
  assign \new_[14810]_  = ~A167 & A168;
  assign \new_[14811]_  = A169 & \new_[14810]_ ;
  assign \new_[14815]_  = ~A200 & A199;
  assign \new_[14816]_  = A166 & \new_[14815]_ ;
  assign \new_[14817]_  = \new_[14816]_  & \new_[14811]_ ;
  assign \new_[14821]_  = A233 & ~A203;
  assign \new_[14822]_  = ~A201 & \new_[14821]_ ;
  assign \new_[14826]_  = A267 & A265;
  assign \new_[14827]_  = A234 & \new_[14826]_ ;
  assign \new_[14828]_  = \new_[14827]_  & \new_[14822]_ ;
  assign \new_[14832]_  = ~A167 & A168;
  assign \new_[14833]_  = A169 & \new_[14832]_ ;
  assign \new_[14837]_  = ~A200 & A199;
  assign \new_[14838]_  = A166 & \new_[14837]_ ;
  assign \new_[14839]_  = \new_[14838]_  & \new_[14833]_ ;
  assign \new_[14843]_  = A233 & ~A203;
  assign \new_[14844]_  = ~A201 & \new_[14843]_ ;
  assign \new_[14848]_  = A267 & A266;
  assign \new_[14849]_  = A234 & \new_[14848]_ ;
  assign \new_[14850]_  = \new_[14849]_  & \new_[14844]_ ;
  assign \new_[14854]_  = ~A199 & ~A166;
  assign \new_[14855]_  = A167 & \new_[14854]_ ;
  assign \new_[14859]_  = A232 & ~A202;
  assign \new_[14860]_  = ~A200 & \new_[14859]_ ;
  assign \new_[14861]_  = \new_[14860]_  & \new_[14855]_ ;
  assign \new_[14865]_  = ~A236 & A235;
  assign \new_[14866]_  = A233 & \new_[14865]_ ;
  assign \new_[14869]_  = A299 & A298;
  assign \new_[14872]_  = ~A302 & A301;
  assign \new_[14873]_  = \new_[14872]_  & \new_[14869]_ ;
  assign \new_[14874]_  = \new_[14873]_  & \new_[14866]_ ;
  assign \new_[14878]_  = ~A199 & ~A166;
  assign \new_[14879]_  = A167 & \new_[14878]_ ;
  assign \new_[14883]_  = A232 & ~A202;
  assign \new_[14884]_  = ~A200 & \new_[14883]_ ;
  assign \new_[14885]_  = \new_[14884]_  & \new_[14879]_ ;
  assign \new_[14889]_  = ~A236 & A235;
  assign \new_[14890]_  = A233 & \new_[14889]_ ;
  assign \new_[14893]_  = ~A299 & A298;
  assign \new_[14896]_  = A302 & ~A301;
  assign \new_[14897]_  = \new_[14896]_  & \new_[14893]_ ;
  assign \new_[14898]_  = \new_[14897]_  & \new_[14890]_ ;
  assign \new_[14902]_  = ~A199 & ~A166;
  assign \new_[14903]_  = A167 & \new_[14902]_ ;
  assign \new_[14907]_  = A232 & ~A202;
  assign \new_[14908]_  = ~A200 & \new_[14907]_ ;
  assign \new_[14909]_  = \new_[14908]_  & \new_[14903]_ ;
  assign \new_[14913]_  = ~A236 & A235;
  assign \new_[14914]_  = A233 & \new_[14913]_ ;
  assign \new_[14917]_  = A299 & ~A298;
  assign \new_[14920]_  = A302 & ~A301;
  assign \new_[14921]_  = \new_[14920]_  & \new_[14917]_ ;
  assign \new_[14922]_  = \new_[14921]_  & \new_[14914]_ ;
  assign \new_[14926]_  = ~A199 & ~A166;
  assign \new_[14927]_  = A167 & \new_[14926]_ ;
  assign \new_[14931]_  = A232 & ~A202;
  assign \new_[14932]_  = ~A200 & \new_[14931]_ ;
  assign \new_[14933]_  = \new_[14932]_  & \new_[14927]_ ;
  assign \new_[14937]_  = ~A236 & A235;
  assign \new_[14938]_  = A233 & \new_[14937]_ ;
  assign \new_[14941]_  = ~A299 & ~A298;
  assign \new_[14944]_  = ~A302 & A301;
  assign \new_[14945]_  = \new_[14944]_  & \new_[14941]_ ;
  assign \new_[14946]_  = \new_[14945]_  & \new_[14938]_ ;
  assign \new_[14950]_  = ~A199 & ~A166;
  assign \new_[14951]_  = A167 & \new_[14950]_ ;
  assign \new_[14955]_  = A232 & ~A202;
  assign \new_[14956]_  = ~A200 & \new_[14955]_ ;
  assign \new_[14957]_  = \new_[14956]_  & \new_[14951]_ ;
  assign \new_[14961]_  = ~A236 & A235;
  assign \new_[14962]_  = A233 & \new_[14961]_ ;
  assign \new_[14965]_  = A266 & A265;
  assign \new_[14968]_  = ~A269 & A268;
  assign \new_[14969]_  = \new_[14968]_  & \new_[14965]_ ;
  assign \new_[14970]_  = \new_[14969]_  & \new_[14962]_ ;
  assign \new_[14974]_  = ~A199 & ~A166;
  assign \new_[14975]_  = A167 & \new_[14974]_ ;
  assign \new_[14979]_  = A232 & ~A202;
  assign \new_[14980]_  = ~A200 & \new_[14979]_ ;
  assign \new_[14981]_  = \new_[14980]_  & \new_[14975]_ ;
  assign \new_[14985]_  = ~A236 & A235;
  assign \new_[14986]_  = A233 & \new_[14985]_ ;
  assign \new_[14989]_  = A266 & ~A265;
  assign \new_[14992]_  = A269 & ~A268;
  assign \new_[14993]_  = \new_[14992]_  & \new_[14989]_ ;
  assign \new_[14994]_  = \new_[14993]_  & \new_[14986]_ ;
  assign \new_[14998]_  = ~A199 & ~A166;
  assign \new_[14999]_  = A167 & \new_[14998]_ ;
  assign \new_[15003]_  = A232 & ~A202;
  assign \new_[15004]_  = ~A200 & \new_[15003]_ ;
  assign \new_[15005]_  = \new_[15004]_  & \new_[14999]_ ;
  assign \new_[15009]_  = ~A236 & A235;
  assign \new_[15010]_  = A233 & \new_[15009]_ ;
  assign \new_[15013]_  = ~A266 & A265;
  assign \new_[15016]_  = A269 & ~A268;
  assign \new_[15017]_  = \new_[15016]_  & \new_[15013]_ ;
  assign \new_[15018]_  = \new_[15017]_  & \new_[15010]_ ;
  assign \new_[15022]_  = ~A199 & ~A166;
  assign \new_[15023]_  = A167 & \new_[15022]_ ;
  assign \new_[15027]_  = A232 & ~A202;
  assign \new_[15028]_  = ~A200 & \new_[15027]_ ;
  assign \new_[15029]_  = \new_[15028]_  & \new_[15023]_ ;
  assign \new_[15033]_  = ~A236 & A235;
  assign \new_[15034]_  = A233 & \new_[15033]_ ;
  assign \new_[15037]_  = ~A266 & ~A265;
  assign \new_[15040]_  = ~A269 & A268;
  assign \new_[15041]_  = \new_[15040]_  & \new_[15037]_ ;
  assign \new_[15042]_  = \new_[15041]_  & \new_[15034]_ ;
  assign \new_[15046]_  = ~A199 & ~A166;
  assign \new_[15047]_  = A167 & \new_[15046]_ ;
  assign \new_[15051]_  = ~A232 & ~A202;
  assign \new_[15052]_  = ~A200 & \new_[15051]_ ;
  assign \new_[15053]_  = \new_[15052]_  & \new_[15047]_ ;
  assign \new_[15057]_  = A236 & ~A235;
  assign \new_[15058]_  = A233 & \new_[15057]_ ;
  assign \new_[15061]_  = A299 & A298;
  assign \new_[15064]_  = ~A302 & A301;
  assign \new_[15065]_  = \new_[15064]_  & \new_[15061]_ ;
  assign \new_[15066]_  = \new_[15065]_  & \new_[15058]_ ;
  assign \new_[15070]_  = ~A199 & ~A166;
  assign \new_[15071]_  = A167 & \new_[15070]_ ;
  assign \new_[15075]_  = ~A232 & ~A202;
  assign \new_[15076]_  = ~A200 & \new_[15075]_ ;
  assign \new_[15077]_  = \new_[15076]_  & \new_[15071]_ ;
  assign \new_[15081]_  = A236 & ~A235;
  assign \new_[15082]_  = A233 & \new_[15081]_ ;
  assign \new_[15085]_  = ~A299 & A298;
  assign \new_[15088]_  = A302 & ~A301;
  assign \new_[15089]_  = \new_[15088]_  & \new_[15085]_ ;
  assign \new_[15090]_  = \new_[15089]_  & \new_[15082]_ ;
  assign \new_[15094]_  = ~A199 & ~A166;
  assign \new_[15095]_  = A167 & \new_[15094]_ ;
  assign \new_[15099]_  = ~A232 & ~A202;
  assign \new_[15100]_  = ~A200 & \new_[15099]_ ;
  assign \new_[15101]_  = \new_[15100]_  & \new_[15095]_ ;
  assign \new_[15105]_  = A236 & ~A235;
  assign \new_[15106]_  = A233 & \new_[15105]_ ;
  assign \new_[15109]_  = A299 & ~A298;
  assign \new_[15112]_  = A302 & ~A301;
  assign \new_[15113]_  = \new_[15112]_  & \new_[15109]_ ;
  assign \new_[15114]_  = \new_[15113]_  & \new_[15106]_ ;
  assign \new_[15118]_  = ~A199 & ~A166;
  assign \new_[15119]_  = A167 & \new_[15118]_ ;
  assign \new_[15123]_  = ~A232 & ~A202;
  assign \new_[15124]_  = ~A200 & \new_[15123]_ ;
  assign \new_[15125]_  = \new_[15124]_  & \new_[15119]_ ;
  assign \new_[15129]_  = A236 & ~A235;
  assign \new_[15130]_  = A233 & \new_[15129]_ ;
  assign \new_[15133]_  = ~A299 & ~A298;
  assign \new_[15136]_  = ~A302 & A301;
  assign \new_[15137]_  = \new_[15136]_  & \new_[15133]_ ;
  assign \new_[15138]_  = \new_[15137]_  & \new_[15130]_ ;
  assign \new_[15142]_  = ~A199 & ~A166;
  assign \new_[15143]_  = A167 & \new_[15142]_ ;
  assign \new_[15147]_  = ~A232 & ~A202;
  assign \new_[15148]_  = ~A200 & \new_[15147]_ ;
  assign \new_[15149]_  = \new_[15148]_  & \new_[15143]_ ;
  assign \new_[15153]_  = A236 & ~A235;
  assign \new_[15154]_  = A233 & \new_[15153]_ ;
  assign \new_[15157]_  = A266 & A265;
  assign \new_[15160]_  = ~A269 & A268;
  assign \new_[15161]_  = \new_[15160]_  & \new_[15157]_ ;
  assign \new_[15162]_  = \new_[15161]_  & \new_[15154]_ ;
  assign \new_[15166]_  = ~A199 & ~A166;
  assign \new_[15167]_  = A167 & \new_[15166]_ ;
  assign \new_[15171]_  = ~A232 & ~A202;
  assign \new_[15172]_  = ~A200 & \new_[15171]_ ;
  assign \new_[15173]_  = \new_[15172]_  & \new_[15167]_ ;
  assign \new_[15177]_  = A236 & ~A235;
  assign \new_[15178]_  = A233 & \new_[15177]_ ;
  assign \new_[15181]_  = A266 & ~A265;
  assign \new_[15184]_  = A269 & ~A268;
  assign \new_[15185]_  = \new_[15184]_  & \new_[15181]_ ;
  assign \new_[15186]_  = \new_[15185]_  & \new_[15178]_ ;
  assign \new_[15190]_  = ~A199 & ~A166;
  assign \new_[15191]_  = A167 & \new_[15190]_ ;
  assign \new_[15195]_  = ~A232 & ~A202;
  assign \new_[15196]_  = ~A200 & \new_[15195]_ ;
  assign \new_[15197]_  = \new_[15196]_  & \new_[15191]_ ;
  assign \new_[15201]_  = A236 & ~A235;
  assign \new_[15202]_  = A233 & \new_[15201]_ ;
  assign \new_[15205]_  = ~A266 & A265;
  assign \new_[15208]_  = A269 & ~A268;
  assign \new_[15209]_  = \new_[15208]_  & \new_[15205]_ ;
  assign \new_[15210]_  = \new_[15209]_  & \new_[15202]_ ;
  assign \new_[15214]_  = ~A199 & ~A166;
  assign \new_[15215]_  = A167 & \new_[15214]_ ;
  assign \new_[15219]_  = ~A232 & ~A202;
  assign \new_[15220]_  = ~A200 & \new_[15219]_ ;
  assign \new_[15221]_  = \new_[15220]_  & \new_[15215]_ ;
  assign \new_[15225]_  = A236 & ~A235;
  assign \new_[15226]_  = A233 & \new_[15225]_ ;
  assign \new_[15229]_  = ~A266 & ~A265;
  assign \new_[15232]_  = ~A269 & A268;
  assign \new_[15233]_  = \new_[15232]_  & \new_[15229]_ ;
  assign \new_[15234]_  = \new_[15233]_  & \new_[15226]_ ;
  assign \new_[15238]_  = ~A199 & ~A166;
  assign \new_[15239]_  = A167 & \new_[15238]_ ;
  assign \new_[15243]_  = A232 & ~A202;
  assign \new_[15244]_  = ~A200 & \new_[15243]_ ;
  assign \new_[15245]_  = \new_[15244]_  & \new_[15239]_ ;
  assign \new_[15249]_  = A236 & ~A235;
  assign \new_[15250]_  = ~A233 & \new_[15249]_ ;
  assign \new_[15253]_  = A299 & A298;
  assign \new_[15256]_  = ~A302 & A301;
  assign \new_[15257]_  = \new_[15256]_  & \new_[15253]_ ;
  assign \new_[15258]_  = \new_[15257]_  & \new_[15250]_ ;
  assign \new_[15262]_  = ~A199 & ~A166;
  assign \new_[15263]_  = A167 & \new_[15262]_ ;
  assign \new_[15267]_  = A232 & ~A202;
  assign \new_[15268]_  = ~A200 & \new_[15267]_ ;
  assign \new_[15269]_  = \new_[15268]_  & \new_[15263]_ ;
  assign \new_[15273]_  = A236 & ~A235;
  assign \new_[15274]_  = ~A233 & \new_[15273]_ ;
  assign \new_[15277]_  = ~A299 & A298;
  assign \new_[15280]_  = A302 & ~A301;
  assign \new_[15281]_  = \new_[15280]_  & \new_[15277]_ ;
  assign \new_[15282]_  = \new_[15281]_  & \new_[15274]_ ;
  assign \new_[15286]_  = ~A199 & ~A166;
  assign \new_[15287]_  = A167 & \new_[15286]_ ;
  assign \new_[15291]_  = A232 & ~A202;
  assign \new_[15292]_  = ~A200 & \new_[15291]_ ;
  assign \new_[15293]_  = \new_[15292]_  & \new_[15287]_ ;
  assign \new_[15297]_  = A236 & ~A235;
  assign \new_[15298]_  = ~A233 & \new_[15297]_ ;
  assign \new_[15301]_  = A299 & ~A298;
  assign \new_[15304]_  = A302 & ~A301;
  assign \new_[15305]_  = \new_[15304]_  & \new_[15301]_ ;
  assign \new_[15306]_  = \new_[15305]_  & \new_[15298]_ ;
  assign \new_[15310]_  = ~A199 & ~A166;
  assign \new_[15311]_  = A167 & \new_[15310]_ ;
  assign \new_[15315]_  = A232 & ~A202;
  assign \new_[15316]_  = ~A200 & \new_[15315]_ ;
  assign \new_[15317]_  = \new_[15316]_  & \new_[15311]_ ;
  assign \new_[15321]_  = A236 & ~A235;
  assign \new_[15322]_  = ~A233 & \new_[15321]_ ;
  assign \new_[15325]_  = ~A299 & ~A298;
  assign \new_[15328]_  = ~A302 & A301;
  assign \new_[15329]_  = \new_[15328]_  & \new_[15325]_ ;
  assign \new_[15330]_  = \new_[15329]_  & \new_[15322]_ ;
  assign \new_[15334]_  = ~A199 & ~A166;
  assign \new_[15335]_  = A167 & \new_[15334]_ ;
  assign \new_[15339]_  = A232 & ~A202;
  assign \new_[15340]_  = ~A200 & \new_[15339]_ ;
  assign \new_[15341]_  = \new_[15340]_  & \new_[15335]_ ;
  assign \new_[15345]_  = A236 & ~A235;
  assign \new_[15346]_  = ~A233 & \new_[15345]_ ;
  assign \new_[15349]_  = A266 & A265;
  assign \new_[15352]_  = ~A269 & A268;
  assign \new_[15353]_  = \new_[15352]_  & \new_[15349]_ ;
  assign \new_[15354]_  = \new_[15353]_  & \new_[15346]_ ;
  assign \new_[15358]_  = ~A199 & ~A166;
  assign \new_[15359]_  = A167 & \new_[15358]_ ;
  assign \new_[15363]_  = A232 & ~A202;
  assign \new_[15364]_  = ~A200 & \new_[15363]_ ;
  assign \new_[15365]_  = \new_[15364]_  & \new_[15359]_ ;
  assign \new_[15369]_  = A236 & ~A235;
  assign \new_[15370]_  = ~A233 & \new_[15369]_ ;
  assign \new_[15373]_  = A266 & ~A265;
  assign \new_[15376]_  = A269 & ~A268;
  assign \new_[15377]_  = \new_[15376]_  & \new_[15373]_ ;
  assign \new_[15378]_  = \new_[15377]_  & \new_[15370]_ ;
  assign \new_[15382]_  = ~A199 & ~A166;
  assign \new_[15383]_  = A167 & \new_[15382]_ ;
  assign \new_[15387]_  = A232 & ~A202;
  assign \new_[15388]_  = ~A200 & \new_[15387]_ ;
  assign \new_[15389]_  = \new_[15388]_  & \new_[15383]_ ;
  assign \new_[15393]_  = A236 & ~A235;
  assign \new_[15394]_  = ~A233 & \new_[15393]_ ;
  assign \new_[15397]_  = ~A266 & A265;
  assign \new_[15400]_  = A269 & ~A268;
  assign \new_[15401]_  = \new_[15400]_  & \new_[15397]_ ;
  assign \new_[15402]_  = \new_[15401]_  & \new_[15394]_ ;
  assign \new_[15406]_  = ~A199 & ~A166;
  assign \new_[15407]_  = A167 & \new_[15406]_ ;
  assign \new_[15411]_  = A232 & ~A202;
  assign \new_[15412]_  = ~A200 & \new_[15411]_ ;
  assign \new_[15413]_  = \new_[15412]_  & \new_[15407]_ ;
  assign \new_[15417]_  = A236 & ~A235;
  assign \new_[15418]_  = ~A233 & \new_[15417]_ ;
  assign \new_[15421]_  = ~A266 & ~A265;
  assign \new_[15424]_  = ~A269 & A268;
  assign \new_[15425]_  = \new_[15424]_  & \new_[15421]_ ;
  assign \new_[15426]_  = \new_[15425]_  & \new_[15418]_ ;
  assign \new_[15430]_  = ~A199 & ~A166;
  assign \new_[15431]_  = A167 & \new_[15430]_ ;
  assign \new_[15435]_  = ~A232 & ~A202;
  assign \new_[15436]_  = ~A200 & \new_[15435]_ ;
  assign \new_[15437]_  = \new_[15436]_  & \new_[15431]_ ;
  assign \new_[15441]_  = ~A236 & A235;
  assign \new_[15442]_  = ~A233 & \new_[15441]_ ;
  assign \new_[15445]_  = A299 & A298;
  assign \new_[15448]_  = ~A302 & A301;
  assign \new_[15449]_  = \new_[15448]_  & \new_[15445]_ ;
  assign \new_[15450]_  = \new_[15449]_  & \new_[15442]_ ;
  assign \new_[15454]_  = ~A199 & ~A166;
  assign \new_[15455]_  = A167 & \new_[15454]_ ;
  assign \new_[15459]_  = ~A232 & ~A202;
  assign \new_[15460]_  = ~A200 & \new_[15459]_ ;
  assign \new_[15461]_  = \new_[15460]_  & \new_[15455]_ ;
  assign \new_[15465]_  = ~A236 & A235;
  assign \new_[15466]_  = ~A233 & \new_[15465]_ ;
  assign \new_[15469]_  = ~A299 & A298;
  assign \new_[15472]_  = A302 & ~A301;
  assign \new_[15473]_  = \new_[15472]_  & \new_[15469]_ ;
  assign \new_[15474]_  = \new_[15473]_  & \new_[15466]_ ;
  assign \new_[15478]_  = ~A199 & ~A166;
  assign \new_[15479]_  = A167 & \new_[15478]_ ;
  assign \new_[15483]_  = ~A232 & ~A202;
  assign \new_[15484]_  = ~A200 & \new_[15483]_ ;
  assign \new_[15485]_  = \new_[15484]_  & \new_[15479]_ ;
  assign \new_[15489]_  = ~A236 & A235;
  assign \new_[15490]_  = ~A233 & \new_[15489]_ ;
  assign \new_[15493]_  = A299 & ~A298;
  assign \new_[15496]_  = A302 & ~A301;
  assign \new_[15497]_  = \new_[15496]_  & \new_[15493]_ ;
  assign \new_[15498]_  = \new_[15497]_  & \new_[15490]_ ;
  assign \new_[15502]_  = ~A199 & ~A166;
  assign \new_[15503]_  = A167 & \new_[15502]_ ;
  assign \new_[15507]_  = ~A232 & ~A202;
  assign \new_[15508]_  = ~A200 & \new_[15507]_ ;
  assign \new_[15509]_  = \new_[15508]_  & \new_[15503]_ ;
  assign \new_[15513]_  = ~A236 & A235;
  assign \new_[15514]_  = ~A233 & \new_[15513]_ ;
  assign \new_[15517]_  = ~A299 & ~A298;
  assign \new_[15520]_  = ~A302 & A301;
  assign \new_[15521]_  = \new_[15520]_  & \new_[15517]_ ;
  assign \new_[15522]_  = \new_[15521]_  & \new_[15514]_ ;
  assign \new_[15526]_  = ~A199 & ~A166;
  assign \new_[15527]_  = A167 & \new_[15526]_ ;
  assign \new_[15531]_  = ~A232 & ~A202;
  assign \new_[15532]_  = ~A200 & \new_[15531]_ ;
  assign \new_[15533]_  = \new_[15532]_  & \new_[15527]_ ;
  assign \new_[15537]_  = ~A236 & A235;
  assign \new_[15538]_  = ~A233 & \new_[15537]_ ;
  assign \new_[15541]_  = A266 & A265;
  assign \new_[15544]_  = ~A269 & A268;
  assign \new_[15545]_  = \new_[15544]_  & \new_[15541]_ ;
  assign \new_[15546]_  = \new_[15545]_  & \new_[15538]_ ;
  assign \new_[15550]_  = ~A199 & ~A166;
  assign \new_[15551]_  = A167 & \new_[15550]_ ;
  assign \new_[15555]_  = ~A232 & ~A202;
  assign \new_[15556]_  = ~A200 & \new_[15555]_ ;
  assign \new_[15557]_  = \new_[15556]_  & \new_[15551]_ ;
  assign \new_[15561]_  = ~A236 & A235;
  assign \new_[15562]_  = ~A233 & \new_[15561]_ ;
  assign \new_[15565]_  = A266 & ~A265;
  assign \new_[15568]_  = A269 & ~A268;
  assign \new_[15569]_  = \new_[15568]_  & \new_[15565]_ ;
  assign \new_[15570]_  = \new_[15569]_  & \new_[15562]_ ;
  assign \new_[15574]_  = ~A199 & ~A166;
  assign \new_[15575]_  = A167 & \new_[15574]_ ;
  assign \new_[15579]_  = ~A232 & ~A202;
  assign \new_[15580]_  = ~A200 & \new_[15579]_ ;
  assign \new_[15581]_  = \new_[15580]_  & \new_[15575]_ ;
  assign \new_[15585]_  = ~A236 & A235;
  assign \new_[15586]_  = ~A233 & \new_[15585]_ ;
  assign \new_[15589]_  = ~A266 & A265;
  assign \new_[15592]_  = A269 & ~A268;
  assign \new_[15593]_  = \new_[15592]_  & \new_[15589]_ ;
  assign \new_[15594]_  = \new_[15593]_  & \new_[15586]_ ;
  assign \new_[15598]_  = ~A199 & ~A166;
  assign \new_[15599]_  = A167 & \new_[15598]_ ;
  assign \new_[15603]_  = ~A232 & ~A202;
  assign \new_[15604]_  = ~A200 & \new_[15603]_ ;
  assign \new_[15605]_  = \new_[15604]_  & \new_[15599]_ ;
  assign \new_[15609]_  = ~A236 & A235;
  assign \new_[15610]_  = ~A233 & \new_[15609]_ ;
  assign \new_[15613]_  = ~A266 & ~A265;
  assign \new_[15616]_  = ~A269 & A268;
  assign \new_[15617]_  = \new_[15616]_  & \new_[15613]_ ;
  assign \new_[15618]_  = \new_[15617]_  & \new_[15610]_ ;
  assign \new_[15622]_  = ~A199 & ~A166;
  assign \new_[15623]_  = A167 & \new_[15622]_ ;
  assign \new_[15627]_  = A232 & A203;
  assign \new_[15628]_  = ~A200 & \new_[15627]_ ;
  assign \new_[15629]_  = \new_[15628]_  & \new_[15623]_ ;
  assign \new_[15633]_  = ~A236 & A235;
  assign \new_[15634]_  = A233 & \new_[15633]_ ;
  assign \new_[15637]_  = A299 & A298;
  assign \new_[15640]_  = ~A302 & A301;
  assign \new_[15641]_  = \new_[15640]_  & \new_[15637]_ ;
  assign \new_[15642]_  = \new_[15641]_  & \new_[15634]_ ;
  assign \new_[15646]_  = ~A199 & ~A166;
  assign \new_[15647]_  = A167 & \new_[15646]_ ;
  assign \new_[15651]_  = A232 & A203;
  assign \new_[15652]_  = ~A200 & \new_[15651]_ ;
  assign \new_[15653]_  = \new_[15652]_  & \new_[15647]_ ;
  assign \new_[15657]_  = ~A236 & A235;
  assign \new_[15658]_  = A233 & \new_[15657]_ ;
  assign \new_[15661]_  = ~A299 & A298;
  assign \new_[15664]_  = A302 & ~A301;
  assign \new_[15665]_  = \new_[15664]_  & \new_[15661]_ ;
  assign \new_[15666]_  = \new_[15665]_  & \new_[15658]_ ;
  assign \new_[15670]_  = ~A199 & ~A166;
  assign \new_[15671]_  = A167 & \new_[15670]_ ;
  assign \new_[15675]_  = A232 & A203;
  assign \new_[15676]_  = ~A200 & \new_[15675]_ ;
  assign \new_[15677]_  = \new_[15676]_  & \new_[15671]_ ;
  assign \new_[15681]_  = ~A236 & A235;
  assign \new_[15682]_  = A233 & \new_[15681]_ ;
  assign \new_[15685]_  = A299 & ~A298;
  assign \new_[15688]_  = A302 & ~A301;
  assign \new_[15689]_  = \new_[15688]_  & \new_[15685]_ ;
  assign \new_[15690]_  = \new_[15689]_  & \new_[15682]_ ;
  assign \new_[15694]_  = ~A199 & ~A166;
  assign \new_[15695]_  = A167 & \new_[15694]_ ;
  assign \new_[15699]_  = A232 & A203;
  assign \new_[15700]_  = ~A200 & \new_[15699]_ ;
  assign \new_[15701]_  = \new_[15700]_  & \new_[15695]_ ;
  assign \new_[15705]_  = ~A236 & A235;
  assign \new_[15706]_  = A233 & \new_[15705]_ ;
  assign \new_[15709]_  = ~A299 & ~A298;
  assign \new_[15712]_  = ~A302 & A301;
  assign \new_[15713]_  = \new_[15712]_  & \new_[15709]_ ;
  assign \new_[15714]_  = \new_[15713]_  & \new_[15706]_ ;
  assign \new_[15718]_  = ~A199 & ~A166;
  assign \new_[15719]_  = A167 & \new_[15718]_ ;
  assign \new_[15723]_  = A232 & A203;
  assign \new_[15724]_  = ~A200 & \new_[15723]_ ;
  assign \new_[15725]_  = \new_[15724]_  & \new_[15719]_ ;
  assign \new_[15729]_  = ~A236 & A235;
  assign \new_[15730]_  = A233 & \new_[15729]_ ;
  assign \new_[15733]_  = A266 & A265;
  assign \new_[15736]_  = ~A269 & A268;
  assign \new_[15737]_  = \new_[15736]_  & \new_[15733]_ ;
  assign \new_[15738]_  = \new_[15737]_  & \new_[15730]_ ;
  assign \new_[15742]_  = ~A199 & ~A166;
  assign \new_[15743]_  = A167 & \new_[15742]_ ;
  assign \new_[15747]_  = A232 & A203;
  assign \new_[15748]_  = ~A200 & \new_[15747]_ ;
  assign \new_[15749]_  = \new_[15748]_  & \new_[15743]_ ;
  assign \new_[15753]_  = ~A236 & A235;
  assign \new_[15754]_  = A233 & \new_[15753]_ ;
  assign \new_[15757]_  = A266 & ~A265;
  assign \new_[15760]_  = A269 & ~A268;
  assign \new_[15761]_  = \new_[15760]_  & \new_[15757]_ ;
  assign \new_[15762]_  = \new_[15761]_  & \new_[15754]_ ;
  assign \new_[15766]_  = ~A199 & ~A166;
  assign \new_[15767]_  = A167 & \new_[15766]_ ;
  assign \new_[15771]_  = A232 & A203;
  assign \new_[15772]_  = ~A200 & \new_[15771]_ ;
  assign \new_[15773]_  = \new_[15772]_  & \new_[15767]_ ;
  assign \new_[15777]_  = ~A236 & A235;
  assign \new_[15778]_  = A233 & \new_[15777]_ ;
  assign \new_[15781]_  = ~A266 & A265;
  assign \new_[15784]_  = A269 & ~A268;
  assign \new_[15785]_  = \new_[15784]_  & \new_[15781]_ ;
  assign \new_[15786]_  = \new_[15785]_  & \new_[15778]_ ;
  assign \new_[15790]_  = ~A199 & ~A166;
  assign \new_[15791]_  = A167 & \new_[15790]_ ;
  assign \new_[15795]_  = A232 & A203;
  assign \new_[15796]_  = ~A200 & \new_[15795]_ ;
  assign \new_[15797]_  = \new_[15796]_  & \new_[15791]_ ;
  assign \new_[15801]_  = ~A236 & A235;
  assign \new_[15802]_  = A233 & \new_[15801]_ ;
  assign \new_[15805]_  = ~A266 & ~A265;
  assign \new_[15808]_  = ~A269 & A268;
  assign \new_[15809]_  = \new_[15808]_  & \new_[15805]_ ;
  assign \new_[15810]_  = \new_[15809]_  & \new_[15802]_ ;
  assign \new_[15814]_  = ~A199 & ~A166;
  assign \new_[15815]_  = A167 & \new_[15814]_ ;
  assign \new_[15819]_  = ~A232 & A203;
  assign \new_[15820]_  = ~A200 & \new_[15819]_ ;
  assign \new_[15821]_  = \new_[15820]_  & \new_[15815]_ ;
  assign \new_[15825]_  = A236 & ~A235;
  assign \new_[15826]_  = A233 & \new_[15825]_ ;
  assign \new_[15829]_  = A299 & A298;
  assign \new_[15832]_  = ~A302 & A301;
  assign \new_[15833]_  = \new_[15832]_  & \new_[15829]_ ;
  assign \new_[15834]_  = \new_[15833]_  & \new_[15826]_ ;
  assign \new_[15838]_  = ~A199 & ~A166;
  assign \new_[15839]_  = A167 & \new_[15838]_ ;
  assign \new_[15843]_  = ~A232 & A203;
  assign \new_[15844]_  = ~A200 & \new_[15843]_ ;
  assign \new_[15845]_  = \new_[15844]_  & \new_[15839]_ ;
  assign \new_[15849]_  = A236 & ~A235;
  assign \new_[15850]_  = A233 & \new_[15849]_ ;
  assign \new_[15853]_  = ~A299 & A298;
  assign \new_[15856]_  = A302 & ~A301;
  assign \new_[15857]_  = \new_[15856]_  & \new_[15853]_ ;
  assign \new_[15858]_  = \new_[15857]_  & \new_[15850]_ ;
  assign \new_[15862]_  = ~A199 & ~A166;
  assign \new_[15863]_  = A167 & \new_[15862]_ ;
  assign \new_[15867]_  = ~A232 & A203;
  assign \new_[15868]_  = ~A200 & \new_[15867]_ ;
  assign \new_[15869]_  = \new_[15868]_  & \new_[15863]_ ;
  assign \new_[15873]_  = A236 & ~A235;
  assign \new_[15874]_  = A233 & \new_[15873]_ ;
  assign \new_[15877]_  = A299 & ~A298;
  assign \new_[15880]_  = A302 & ~A301;
  assign \new_[15881]_  = \new_[15880]_  & \new_[15877]_ ;
  assign \new_[15882]_  = \new_[15881]_  & \new_[15874]_ ;
  assign \new_[15886]_  = ~A199 & ~A166;
  assign \new_[15887]_  = A167 & \new_[15886]_ ;
  assign \new_[15891]_  = ~A232 & A203;
  assign \new_[15892]_  = ~A200 & \new_[15891]_ ;
  assign \new_[15893]_  = \new_[15892]_  & \new_[15887]_ ;
  assign \new_[15897]_  = A236 & ~A235;
  assign \new_[15898]_  = A233 & \new_[15897]_ ;
  assign \new_[15901]_  = ~A299 & ~A298;
  assign \new_[15904]_  = ~A302 & A301;
  assign \new_[15905]_  = \new_[15904]_  & \new_[15901]_ ;
  assign \new_[15906]_  = \new_[15905]_  & \new_[15898]_ ;
  assign \new_[15910]_  = ~A199 & ~A166;
  assign \new_[15911]_  = A167 & \new_[15910]_ ;
  assign \new_[15915]_  = ~A232 & A203;
  assign \new_[15916]_  = ~A200 & \new_[15915]_ ;
  assign \new_[15917]_  = \new_[15916]_  & \new_[15911]_ ;
  assign \new_[15921]_  = A236 & ~A235;
  assign \new_[15922]_  = A233 & \new_[15921]_ ;
  assign \new_[15925]_  = A266 & A265;
  assign \new_[15928]_  = ~A269 & A268;
  assign \new_[15929]_  = \new_[15928]_  & \new_[15925]_ ;
  assign \new_[15930]_  = \new_[15929]_  & \new_[15922]_ ;
  assign \new_[15934]_  = ~A199 & ~A166;
  assign \new_[15935]_  = A167 & \new_[15934]_ ;
  assign \new_[15939]_  = ~A232 & A203;
  assign \new_[15940]_  = ~A200 & \new_[15939]_ ;
  assign \new_[15941]_  = \new_[15940]_  & \new_[15935]_ ;
  assign \new_[15945]_  = A236 & ~A235;
  assign \new_[15946]_  = A233 & \new_[15945]_ ;
  assign \new_[15949]_  = A266 & ~A265;
  assign \new_[15952]_  = A269 & ~A268;
  assign \new_[15953]_  = \new_[15952]_  & \new_[15949]_ ;
  assign \new_[15954]_  = \new_[15953]_  & \new_[15946]_ ;
  assign \new_[15958]_  = ~A199 & ~A166;
  assign \new_[15959]_  = A167 & \new_[15958]_ ;
  assign \new_[15963]_  = ~A232 & A203;
  assign \new_[15964]_  = ~A200 & \new_[15963]_ ;
  assign \new_[15965]_  = \new_[15964]_  & \new_[15959]_ ;
  assign \new_[15969]_  = A236 & ~A235;
  assign \new_[15970]_  = A233 & \new_[15969]_ ;
  assign \new_[15973]_  = ~A266 & A265;
  assign \new_[15976]_  = A269 & ~A268;
  assign \new_[15977]_  = \new_[15976]_  & \new_[15973]_ ;
  assign \new_[15978]_  = \new_[15977]_  & \new_[15970]_ ;
  assign \new_[15982]_  = ~A199 & ~A166;
  assign \new_[15983]_  = A167 & \new_[15982]_ ;
  assign \new_[15987]_  = ~A232 & A203;
  assign \new_[15988]_  = ~A200 & \new_[15987]_ ;
  assign \new_[15989]_  = \new_[15988]_  & \new_[15983]_ ;
  assign \new_[15993]_  = A236 & ~A235;
  assign \new_[15994]_  = A233 & \new_[15993]_ ;
  assign \new_[15997]_  = ~A266 & ~A265;
  assign \new_[16000]_  = ~A269 & A268;
  assign \new_[16001]_  = \new_[16000]_  & \new_[15997]_ ;
  assign \new_[16002]_  = \new_[16001]_  & \new_[15994]_ ;
  assign \new_[16006]_  = ~A199 & ~A166;
  assign \new_[16007]_  = A167 & \new_[16006]_ ;
  assign \new_[16011]_  = A232 & A203;
  assign \new_[16012]_  = ~A200 & \new_[16011]_ ;
  assign \new_[16013]_  = \new_[16012]_  & \new_[16007]_ ;
  assign \new_[16017]_  = A236 & ~A235;
  assign \new_[16018]_  = ~A233 & \new_[16017]_ ;
  assign \new_[16021]_  = A299 & A298;
  assign \new_[16024]_  = ~A302 & A301;
  assign \new_[16025]_  = \new_[16024]_  & \new_[16021]_ ;
  assign \new_[16026]_  = \new_[16025]_  & \new_[16018]_ ;
  assign \new_[16030]_  = ~A199 & ~A166;
  assign \new_[16031]_  = A167 & \new_[16030]_ ;
  assign \new_[16035]_  = A232 & A203;
  assign \new_[16036]_  = ~A200 & \new_[16035]_ ;
  assign \new_[16037]_  = \new_[16036]_  & \new_[16031]_ ;
  assign \new_[16041]_  = A236 & ~A235;
  assign \new_[16042]_  = ~A233 & \new_[16041]_ ;
  assign \new_[16045]_  = ~A299 & A298;
  assign \new_[16048]_  = A302 & ~A301;
  assign \new_[16049]_  = \new_[16048]_  & \new_[16045]_ ;
  assign \new_[16050]_  = \new_[16049]_  & \new_[16042]_ ;
  assign \new_[16054]_  = ~A199 & ~A166;
  assign \new_[16055]_  = A167 & \new_[16054]_ ;
  assign \new_[16059]_  = A232 & A203;
  assign \new_[16060]_  = ~A200 & \new_[16059]_ ;
  assign \new_[16061]_  = \new_[16060]_  & \new_[16055]_ ;
  assign \new_[16065]_  = A236 & ~A235;
  assign \new_[16066]_  = ~A233 & \new_[16065]_ ;
  assign \new_[16069]_  = A299 & ~A298;
  assign \new_[16072]_  = A302 & ~A301;
  assign \new_[16073]_  = \new_[16072]_  & \new_[16069]_ ;
  assign \new_[16074]_  = \new_[16073]_  & \new_[16066]_ ;
  assign \new_[16078]_  = ~A199 & ~A166;
  assign \new_[16079]_  = A167 & \new_[16078]_ ;
  assign \new_[16083]_  = A232 & A203;
  assign \new_[16084]_  = ~A200 & \new_[16083]_ ;
  assign \new_[16085]_  = \new_[16084]_  & \new_[16079]_ ;
  assign \new_[16089]_  = A236 & ~A235;
  assign \new_[16090]_  = ~A233 & \new_[16089]_ ;
  assign \new_[16093]_  = ~A299 & ~A298;
  assign \new_[16096]_  = ~A302 & A301;
  assign \new_[16097]_  = \new_[16096]_  & \new_[16093]_ ;
  assign \new_[16098]_  = \new_[16097]_  & \new_[16090]_ ;
  assign \new_[16102]_  = ~A199 & ~A166;
  assign \new_[16103]_  = A167 & \new_[16102]_ ;
  assign \new_[16107]_  = A232 & A203;
  assign \new_[16108]_  = ~A200 & \new_[16107]_ ;
  assign \new_[16109]_  = \new_[16108]_  & \new_[16103]_ ;
  assign \new_[16113]_  = A236 & ~A235;
  assign \new_[16114]_  = ~A233 & \new_[16113]_ ;
  assign \new_[16117]_  = A266 & A265;
  assign \new_[16120]_  = ~A269 & A268;
  assign \new_[16121]_  = \new_[16120]_  & \new_[16117]_ ;
  assign \new_[16122]_  = \new_[16121]_  & \new_[16114]_ ;
  assign \new_[16126]_  = ~A199 & ~A166;
  assign \new_[16127]_  = A167 & \new_[16126]_ ;
  assign \new_[16131]_  = A232 & A203;
  assign \new_[16132]_  = ~A200 & \new_[16131]_ ;
  assign \new_[16133]_  = \new_[16132]_  & \new_[16127]_ ;
  assign \new_[16137]_  = A236 & ~A235;
  assign \new_[16138]_  = ~A233 & \new_[16137]_ ;
  assign \new_[16141]_  = A266 & ~A265;
  assign \new_[16144]_  = A269 & ~A268;
  assign \new_[16145]_  = \new_[16144]_  & \new_[16141]_ ;
  assign \new_[16146]_  = \new_[16145]_  & \new_[16138]_ ;
  assign \new_[16150]_  = ~A199 & ~A166;
  assign \new_[16151]_  = A167 & \new_[16150]_ ;
  assign \new_[16155]_  = A232 & A203;
  assign \new_[16156]_  = ~A200 & \new_[16155]_ ;
  assign \new_[16157]_  = \new_[16156]_  & \new_[16151]_ ;
  assign \new_[16161]_  = A236 & ~A235;
  assign \new_[16162]_  = ~A233 & \new_[16161]_ ;
  assign \new_[16165]_  = ~A266 & A265;
  assign \new_[16168]_  = A269 & ~A268;
  assign \new_[16169]_  = \new_[16168]_  & \new_[16165]_ ;
  assign \new_[16170]_  = \new_[16169]_  & \new_[16162]_ ;
  assign \new_[16174]_  = ~A199 & ~A166;
  assign \new_[16175]_  = A167 & \new_[16174]_ ;
  assign \new_[16179]_  = A232 & A203;
  assign \new_[16180]_  = ~A200 & \new_[16179]_ ;
  assign \new_[16181]_  = \new_[16180]_  & \new_[16175]_ ;
  assign \new_[16185]_  = A236 & ~A235;
  assign \new_[16186]_  = ~A233 & \new_[16185]_ ;
  assign \new_[16189]_  = ~A266 & ~A265;
  assign \new_[16192]_  = ~A269 & A268;
  assign \new_[16193]_  = \new_[16192]_  & \new_[16189]_ ;
  assign \new_[16194]_  = \new_[16193]_  & \new_[16186]_ ;
  assign \new_[16198]_  = ~A199 & ~A166;
  assign \new_[16199]_  = A167 & \new_[16198]_ ;
  assign \new_[16203]_  = ~A232 & A203;
  assign \new_[16204]_  = ~A200 & \new_[16203]_ ;
  assign \new_[16205]_  = \new_[16204]_  & \new_[16199]_ ;
  assign \new_[16209]_  = ~A236 & A235;
  assign \new_[16210]_  = ~A233 & \new_[16209]_ ;
  assign \new_[16213]_  = A299 & A298;
  assign \new_[16216]_  = ~A302 & A301;
  assign \new_[16217]_  = \new_[16216]_  & \new_[16213]_ ;
  assign \new_[16218]_  = \new_[16217]_  & \new_[16210]_ ;
  assign \new_[16222]_  = ~A199 & ~A166;
  assign \new_[16223]_  = A167 & \new_[16222]_ ;
  assign \new_[16227]_  = ~A232 & A203;
  assign \new_[16228]_  = ~A200 & \new_[16227]_ ;
  assign \new_[16229]_  = \new_[16228]_  & \new_[16223]_ ;
  assign \new_[16233]_  = ~A236 & A235;
  assign \new_[16234]_  = ~A233 & \new_[16233]_ ;
  assign \new_[16237]_  = ~A299 & A298;
  assign \new_[16240]_  = A302 & ~A301;
  assign \new_[16241]_  = \new_[16240]_  & \new_[16237]_ ;
  assign \new_[16242]_  = \new_[16241]_  & \new_[16234]_ ;
  assign \new_[16246]_  = ~A199 & ~A166;
  assign \new_[16247]_  = A167 & \new_[16246]_ ;
  assign \new_[16251]_  = ~A232 & A203;
  assign \new_[16252]_  = ~A200 & \new_[16251]_ ;
  assign \new_[16253]_  = \new_[16252]_  & \new_[16247]_ ;
  assign \new_[16257]_  = ~A236 & A235;
  assign \new_[16258]_  = ~A233 & \new_[16257]_ ;
  assign \new_[16261]_  = A299 & ~A298;
  assign \new_[16264]_  = A302 & ~A301;
  assign \new_[16265]_  = \new_[16264]_  & \new_[16261]_ ;
  assign \new_[16266]_  = \new_[16265]_  & \new_[16258]_ ;
  assign \new_[16270]_  = ~A199 & ~A166;
  assign \new_[16271]_  = A167 & \new_[16270]_ ;
  assign \new_[16275]_  = ~A232 & A203;
  assign \new_[16276]_  = ~A200 & \new_[16275]_ ;
  assign \new_[16277]_  = \new_[16276]_  & \new_[16271]_ ;
  assign \new_[16281]_  = ~A236 & A235;
  assign \new_[16282]_  = ~A233 & \new_[16281]_ ;
  assign \new_[16285]_  = ~A299 & ~A298;
  assign \new_[16288]_  = ~A302 & A301;
  assign \new_[16289]_  = \new_[16288]_  & \new_[16285]_ ;
  assign \new_[16290]_  = \new_[16289]_  & \new_[16282]_ ;
  assign \new_[16294]_  = ~A199 & ~A166;
  assign \new_[16295]_  = A167 & \new_[16294]_ ;
  assign \new_[16299]_  = ~A232 & A203;
  assign \new_[16300]_  = ~A200 & \new_[16299]_ ;
  assign \new_[16301]_  = \new_[16300]_  & \new_[16295]_ ;
  assign \new_[16305]_  = ~A236 & A235;
  assign \new_[16306]_  = ~A233 & \new_[16305]_ ;
  assign \new_[16309]_  = A266 & A265;
  assign \new_[16312]_  = ~A269 & A268;
  assign \new_[16313]_  = \new_[16312]_  & \new_[16309]_ ;
  assign \new_[16314]_  = \new_[16313]_  & \new_[16306]_ ;
  assign \new_[16318]_  = ~A199 & ~A166;
  assign \new_[16319]_  = A167 & \new_[16318]_ ;
  assign \new_[16323]_  = ~A232 & A203;
  assign \new_[16324]_  = ~A200 & \new_[16323]_ ;
  assign \new_[16325]_  = \new_[16324]_  & \new_[16319]_ ;
  assign \new_[16329]_  = ~A236 & A235;
  assign \new_[16330]_  = ~A233 & \new_[16329]_ ;
  assign \new_[16333]_  = A266 & ~A265;
  assign \new_[16336]_  = A269 & ~A268;
  assign \new_[16337]_  = \new_[16336]_  & \new_[16333]_ ;
  assign \new_[16338]_  = \new_[16337]_  & \new_[16330]_ ;
  assign \new_[16342]_  = ~A199 & ~A166;
  assign \new_[16343]_  = A167 & \new_[16342]_ ;
  assign \new_[16347]_  = ~A232 & A203;
  assign \new_[16348]_  = ~A200 & \new_[16347]_ ;
  assign \new_[16349]_  = \new_[16348]_  & \new_[16343]_ ;
  assign \new_[16353]_  = ~A236 & A235;
  assign \new_[16354]_  = ~A233 & \new_[16353]_ ;
  assign \new_[16357]_  = ~A266 & A265;
  assign \new_[16360]_  = A269 & ~A268;
  assign \new_[16361]_  = \new_[16360]_  & \new_[16357]_ ;
  assign \new_[16362]_  = \new_[16361]_  & \new_[16354]_ ;
  assign \new_[16366]_  = ~A199 & ~A166;
  assign \new_[16367]_  = A167 & \new_[16366]_ ;
  assign \new_[16371]_  = ~A232 & A203;
  assign \new_[16372]_  = ~A200 & \new_[16371]_ ;
  assign \new_[16373]_  = \new_[16372]_  & \new_[16367]_ ;
  assign \new_[16377]_  = ~A236 & A235;
  assign \new_[16378]_  = ~A233 & \new_[16377]_ ;
  assign \new_[16381]_  = ~A266 & ~A265;
  assign \new_[16384]_  = ~A269 & A268;
  assign \new_[16385]_  = \new_[16384]_  & \new_[16381]_ ;
  assign \new_[16386]_  = \new_[16385]_  & \new_[16378]_ ;
  assign \new_[16390]_  = ~A167 & A168;
  assign \new_[16391]_  = A170 & \new_[16390]_ ;
  assign \new_[16395]_  = ~A200 & ~A199;
  assign \new_[16396]_  = A166 & \new_[16395]_ ;
  assign \new_[16397]_  = \new_[16396]_  & \new_[16391]_ ;
  assign \new_[16401]_  = A234 & A232;
  assign \new_[16402]_  = ~A202 & \new_[16401]_ ;
  assign \new_[16405]_  = A299 & A298;
  assign \new_[16408]_  = ~A302 & A301;
  assign \new_[16409]_  = \new_[16408]_  & \new_[16405]_ ;
  assign \new_[16410]_  = \new_[16409]_  & \new_[16402]_ ;
  assign \new_[16414]_  = ~A167 & A168;
  assign \new_[16415]_  = A170 & \new_[16414]_ ;
  assign \new_[16419]_  = ~A200 & ~A199;
  assign \new_[16420]_  = A166 & \new_[16419]_ ;
  assign \new_[16421]_  = \new_[16420]_  & \new_[16415]_ ;
  assign \new_[16425]_  = A234 & A232;
  assign \new_[16426]_  = ~A202 & \new_[16425]_ ;
  assign \new_[16429]_  = ~A299 & A298;
  assign \new_[16432]_  = A302 & ~A301;
  assign \new_[16433]_  = \new_[16432]_  & \new_[16429]_ ;
  assign \new_[16434]_  = \new_[16433]_  & \new_[16426]_ ;
  assign \new_[16438]_  = ~A167 & A168;
  assign \new_[16439]_  = A170 & \new_[16438]_ ;
  assign \new_[16443]_  = ~A200 & ~A199;
  assign \new_[16444]_  = A166 & \new_[16443]_ ;
  assign \new_[16445]_  = \new_[16444]_  & \new_[16439]_ ;
  assign \new_[16449]_  = A234 & A232;
  assign \new_[16450]_  = ~A202 & \new_[16449]_ ;
  assign \new_[16453]_  = A299 & ~A298;
  assign \new_[16456]_  = A302 & ~A301;
  assign \new_[16457]_  = \new_[16456]_  & \new_[16453]_ ;
  assign \new_[16458]_  = \new_[16457]_  & \new_[16450]_ ;
  assign \new_[16462]_  = ~A167 & A168;
  assign \new_[16463]_  = A170 & \new_[16462]_ ;
  assign \new_[16467]_  = ~A200 & ~A199;
  assign \new_[16468]_  = A166 & \new_[16467]_ ;
  assign \new_[16469]_  = \new_[16468]_  & \new_[16463]_ ;
  assign \new_[16473]_  = A234 & A232;
  assign \new_[16474]_  = ~A202 & \new_[16473]_ ;
  assign \new_[16477]_  = ~A299 & ~A298;
  assign \new_[16480]_  = ~A302 & A301;
  assign \new_[16481]_  = \new_[16480]_  & \new_[16477]_ ;
  assign \new_[16482]_  = \new_[16481]_  & \new_[16474]_ ;
  assign \new_[16486]_  = ~A167 & A168;
  assign \new_[16487]_  = A170 & \new_[16486]_ ;
  assign \new_[16491]_  = ~A200 & ~A199;
  assign \new_[16492]_  = A166 & \new_[16491]_ ;
  assign \new_[16493]_  = \new_[16492]_  & \new_[16487]_ ;
  assign \new_[16497]_  = A234 & A232;
  assign \new_[16498]_  = ~A202 & \new_[16497]_ ;
  assign \new_[16501]_  = A266 & A265;
  assign \new_[16504]_  = ~A269 & A268;
  assign \new_[16505]_  = \new_[16504]_  & \new_[16501]_ ;
  assign \new_[16506]_  = \new_[16505]_  & \new_[16498]_ ;
  assign \new_[16510]_  = ~A167 & A168;
  assign \new_[16511]_  = A170 & \new_[16510]_ ;
  assign \new_[16515]_  = ~A200 & ~A199;
  assign \new_[16516]_  = A166 & \new_[16515]_ ;
  assign \new_[16517]_  = \new_[16516]_  & \new_[16511]_ ;
  assign \new_[16521]_  = A234 & A232;
  assign \new_[16522]_  = ~A202 & \new_[16521]_ ;
  assign \new_[16525]_  = A266 & ~A265;
  assign \new_[16528]_  = A269 & ~A268;
  assign \new_[16529]_  = \new_[16528]_  & \new_[16525]_ ;
  assign \new_[16530]_  = \new_[16529]_  & \new_[16522]_ ;
  assign \new_[16534]_  = ~A167 & A168;
  assign \new_[16535]_  = A170 & \new_[16534]_ ;
  assign \new_[16539]_  = ~A200 & ~A199;
  assign \new_[16540]_  = A166 & \new_[16539]_ ;
  assign \new_[16541]_  = \new_[16540]_  & \new_[16535]_ ;
  assign \new_[16545]_  = A234 & A232;
  assign \new_[16546]_  = ~A202 & \new_[16545]_ ;
  assign \new_[16549]_  = ~A266 & A265;
  assign \new_[16552]_  = A269 & ~A268;
  assign \new_[16553]_  = \new_[16552]_  & \new_[16549]_ ;
  assign \new_[16554]_  = \new_[16553]_  & \new_[16546]_ ;
  assign \new_[16558]_  = ~A167 & A168;
  assign \new_[16559]_  = A170 & \new_[16558]_ ;
  assign \new_[16563]_  = ~A200 & ~A199;
  assign \new_[16564]_  = A166 & \new_[16563]_ ;
  assign \new_[16565]_  = \new_[16564]_  & \new_[16559]_ ;
  assign \new_[16569]_  = A234 & A232;
  assign \new_[16570]_  = ~A202 & \new_[16569]_ ;
  assign \new_[16573]_  = ~A266 & ~A265;
  assign \new_[16576]_  = ~A269 & A268;
  assign \new_[16577]_  = \new_[16576]_  & \new_[16573]_ ;
  assign \new_[16578]_  = \new_[16577]_  & \new_[16570]_ ;
  assign \new_[16582]_  = ~A167 & A168;
  assign \new_[16583]_  = A170 & \new_[16582]_ ;
  assign \new_[16587]_  = ~A200 & ~A199;
  assign \new_[16588]_  = A166 & \new_[16587]_ ;
  assign \new_[16589]_  = \new_[16588]_  & \new_[16583]_ ;
  assign \new_[16593]_  = A234 & A233;
  assign \new_[16594]_  = ~A202 & \new_[16593]_ ;
  assign \new_[16597]_  = A299 & A298;
  assign \new_[16600]_  = ~A302 & A301;
  assign \new_[16601]_  = \new_[16600]_  & \new_[16597]_ ;
  assign \new_[16602]_  = \new_[16601]_  & \new_[16594]_ ;
  assign \new_[16606]_  = ~A167 & A168;
  assign \new_[16607]_  = A170 & \new_[16606]_ ;
  assign \new_[16611]_  = ~A200 & ~A199;
  assign \new_[16612]_  = A166 & \new_[16611]_ ;
  assign \new_[16613]_  = \new_[16612]_  & \new_[16607]_ ;
  assign \new_[16617]_  = A234 & A233;
  assign \new_[16618]_  = ~A202 & \new_[16617]_ ;
  assign \new_[16621]_  = ~A299 & A298;
  assign \new_[16624]_  = A302 & ~A301;
  assign \new_[16625]_  = \new_[16624]_  & \new_[16621]_ ;
  assign \new_[16626]_  = \new_[16625]_  & \new_[16618]_ ;
  assign \new_[16630]_  = ~A167 & A168;
  assign \new_[16631]_  = A170 & \new_[16630]_ ;
  assign \new_[16635]_  = ~A200 & ~A199;
  assign \new_[16636]_  = A166 & \new_[16635]_ ;
  assign \new_[16637]_  = \new_[16636]_  & \new_[16631]_ ;
  assign \new_[16641]_  = A234 & A233;
  assign \new_[16642]_  = ~A202 & \new_[16641]_ ;
  assign \new_[16645]_  = A299 & ~A298;
  assign \new_[16648]_  = A302 & ~A301;
  assign \new_[16649]_  = \new_[16648]_  & \new_[16645]_ ;
  assign \new_[16650]_  = \new_[16649]_  & \new_[16642]_ ;
  assign \new_[16654]_  = ~A167 & A168;
  assign \new_[16655]_  = A170 & \new_[16654]_ ;
  assign \new_[16659]_  = ~A200 & ~A199;
  assign \new_[16660]_  = A166 & \new_[16659]_ ;
  assign \new_[16661]_  = \new_[16660]_  & \new_[16655]_ ;
  assign \new_[16665]_  = A234 & A233;
  assign \new_[16666]_  = ~A202 & \new_[16665]_ ;
  assign \new_[16669]_  = ~A299 & ~A298;
  assign \new_[16672]_  = ~A302 & A301;
  assign \new_[16673]_  = \new_[16672]_  & \new_[16669]_ ;
  assign \new_[16674]_  = \new_[16673]_  & \new_[16666]_ ;
  assign \new_[16678]_  = ~A167 & A168;
  assign \new_[16679]_  = A170 & \new_[16678]_ ;
  assign \new_[16683]_  = ~A200 & ~A199;
  assign \new_[16684]_  = A166 & \new_[16683]_ ;
  assign \new_[16685]_  = \new_[16684]_  & \new_[16679]_ ;
  assign \new_[16689]_  = A234 & A233;
  assign \new_[16690]_  = ~A202 & \new_[16689]_ ;
  assign \new_[16693]_  = A266 & A265;
  assign \new_[16696]_  = ~A269 & A268;
  assign \new_[16697]_  = \new_[16696]_  & \new_[16693]_ ;
  assign \new_[16698]_  = \new_[16697]_  & \new_[16690]_ ;
  assign \new_[16702]_  = ~A167 & A168;
  assign \new_[16703]_  = A170 & \new_[16702]_ ;
  assign \new_[16707]_  = ~A200 & ~A199;
  assign \new_[16708]_  = A166 & \new_[16707]_ ;
  assign \new_[16709]_  = \new_[16708]_  & \new_[16703]_ ;
  assign \new_[16713]_  = A234 & A233;
  assign \new_[16714]_  = ~A202 & \new_[16713]_ ;
  assign \new_[16717]_  = A266 & ~A265;
  assign \new_[16720]_  = A269 & ~A268;
  assign \new_[16721]_  = \new_[16720]_  & \new_[16717]_ ;
  assign \new_[16722]_  = \new_[16721]_  & \new_[16714]_ ;
  assign \new_[16726]_  = ~A167 & A168;
  assign \new_[16727]_  = A170 & \new_[16726]_ ;
  assign \new_[16731]_  = ~A200 & ~A199;
  assign \new_[16732]_  = A166 & \new_[16731]_ ;
  assign \new_[16733]_  = \new_[16732]_  & \new_[16727]_ ;
  assign \new_[16737]_  = A234 & A233;
  assign \new_[16738]_  = ~A202 & \new_[16737]_ ;
  assign \new_[16741]_  = ~A266 & A265;
  assign \new_[16744]_  = A269 & ~A268;
  assign \new_[16745]_  = \new_[16744]_  & \new_[16741]_ ;
  assign \new_[16746]_  = \new_[16745]_  & \new_[16738]_ ;
  assign \new_[16750]_  = ~A167 & A168;
  assign \new_[16751]_  = A170 & \new_[16750]_ ;
  assign \new_[16755]_  = ~A200 & ~A199;
  assign \new_[16756]_  = A166 & \new_[16755]_ ;
  assign \new_[16757]_  = \new_[16756]_  & \new_[16751]_ ;
  assign \new_[16761]_  = A234 & A233;
  assign \new_[16762]_  = ~A202 & \new_[16761]_ ;
  assign \new_[16765]_  = ~A266 & ~A265;
  assign \new_[16768]_  = ~A269 & A268;
  assign \new_[16769]_  = \new_[16768]_  & \new_[16765]_ ;
  assign \new_[16770]_  = \new_[16769]_  & \new_[16762]_ ;
  assign \new_[16774]_  = ~A167 & A168;
  assign \new_[16775]_  = A170 & \new_[16774]_ ;
  assign \new_[16779]_  = ~A200 & ~A199;
  assign \new_[16780]_  = A166 & \new_[16779]_ ;
  assign \new_[16781]_  = \new_[16780]_  & \new_[16775]_ ;
  assign \new_[16785]_  = A233 & A232;
  assign \new_[16786]_  = ~A202 & \new_[16785]_ ;
  assign \new_[16789]_  = ~A236 & A235;
  assign \new_[16792]_  = A300 & A299;
  assign \new_[16793]_  = \new_[16792]_  & \new_[16789]_ ;
  assign \new_[16794]_  = \new_[16793]_  & \new_[16786]_ ;
  assign \new_[16798]_  = ~A167 & A168;
  assign \new_[16799]_  = A170 & \new_[16798]_ ;
  assign \new_[16803]_  = ~A200 & ~A199;
  assign \new_[16804]_  = A166 & \new_[16803]_ ;
  assign \new_[16805]_  = \new_[16804]_  & \new_[16799]_ ;
  assign \new_[16809]_  = A233 & A232;
  assign \new_[16810]_  = ~A202 & \new_[16809]_ ;
  assign \new_[16813]_  = ~A236 & A235;
  assign \new_[16816]_  = A300 & A298;
  assign \new_[16817]_  = \new_[16816]_  & \new_[16813]_ ;
  assign \new_[16818]_  = \new_[16817]_  & \new_[16810]_ ;
  assign \new_[16822]_  = ~A167 & A168;
  assign \new_[16823]_  = A170 & \new_[16822]_ ;
  assign \new_[16827]_  = ~A200 & ~A199;
  assign \new_[16828]_  = A166 & \new_[16827]_ ;
  assign \new_[16829]_  = \new_[16828]_  & \new_[16823]_ ;
  assign \new_[16833]_  = A233 & A232;
  assign \new_[16834]_  = ~A202 & \new_[16833]_ ;
  assign \new_[16837]_  = ~A236 & A235;
  assign \new_[16840]_  = A267 & A265;
  assign \new_[16841]_  = \new_[16840]_  & \new_[16837]_ ;
  assign \new_[16842]_  = \new_[16841]_  & \new_[16834]_ ;
  assign \new_[16846]_  = ~A167 & A168;
  assign \new_[16847]_  = A170 & \new_[16846]_ ;
  assign \new_[16851]_  = ~A200 & ~A199;
  assign \new_[16852]_  = A166 & \new_[16851]_ ;
  assign \new_[16853]_  = \new_[16852]_  & \new_[16847]_ ;
  assign \new_[16857]_  = A233 & A232;
  assign \new_[16858]_  = ~A202 & \new_[16857]_ ;
  assign \new_[16861]_  = ~A236 & A235;
  assign \new_[16864]_  = A267 & A266;
  assign \new_[16865]_  = \new_[16864]_  & \new_[16861]_ ;
  assign \new_[16866]_  = \new_[16865]_  & \new_[16858]_ ;
  assign \new_[16870]_  = ~A167 & A168;
  assign \new_[16871]_  = A170 & \new_[16870]_ ;
  assign \new_[16875]_  = ~A200 & ~A199;
  assign \new_[16876]_  = A166 & \new_[16875]_ ;
  assign \new_[16877]_  = \new_[16876]_  & \new_[16871]_ ;
  assign \new_[16881]_  = A233 & ~A232;
  assign \new_[16882]_  = ~A202 & \new_[16881]_ ;
  assign \new_[16885]_  = A236 & ~A235;
  assign \new_[16888]_  = A300 & A299;
  assign \new_[16889]_  = \new_[16888]_  & \new_[16885]_ ;
  assign \new_[16890]_  = \new_[16889]_  & \new_[16882]_ ;
  assign \new_[16894]_  = ~A167 & A168;
  assign \new_[16895]_  = A170 & \new_[16894]_ ;
  assign \new_[16899]_  = ~A200 & ~A199;
  assign \new_[16900]_  = A166 & \new_[16899]_ ;
  assign \new_[16901]_  = \new_[16900]_  & \new_[16895]_ ;
  assign \new_[16905]_  = A233 & ~A232;
  assign \new_[16906]_  = ~A202 & \new_[16905]_ ;
  assign \new_[16909]_  = A236 & ~A235;
  assign \new_[16912]_  = A300 & A298;
  assign \new_[16913]_  = \new_[16912]_  & \new_[16909]_ ;
  assign \new_[16914]_  = \new_[16913]_  & \new_[16906]_ ;
  assign \new_[16918]_  = ~A167 & A168;
  assign \new_[16919]_  = A170 & \new_[16918]_ ;
  assign \new_[16923]_  = ~A200 & ~A199;
  assign \new_[16924]_  = A166 & \new_[16923]_ ;
  assign \new_[16925]_  = \new_[16924]_  & \new_[16919]_ ;
  assign \new_[16929]_  = A233 & ~A232;
  assign \new_[16930]_  = ~A202 & \new_[16929]_ ;
  assign \new_[16933]_  = A236 & ~A235;
  assign \new_[16936]_  = A267 & A265;
  assign \new_[16937]_  = \new_[16936]_  & \new_[16933]_ ;
  assign \new_[16938]_  = \new_[16937]_  & \new_[16930]_ ;
  assign \new_[16942]_  = ~A167 & A168;
  assign \new_[16943]_  = A170 & \new_[16942]_ ;
  assign \new_[16947]_  = ~A200 & ~A199;
  assign \new_[16948]_  = A166 & \new_[16947]_ ;
  assign \new_[16949]_  = \new_[16948]_  & \new_[16943]_ ;
  assign \new_[16953]_  = A233 & ~A232;
  assign \new_[16954]_  = ~A202 & \new_[16953]_ ;
  assign \new_[16957]_  = A236 & ~A235;
  assign \new_[16960]_  = A267 & A266;
  assign \new_[16961]_  = \new_[16960]_  & \new_[16957]_ ;
  assign \new_[16962]_  = \new_[16961]_  & \new_[16954]_ ;
  assign \new_[16966]_  = ~A167 & A168;
  assign \new_[16967]_  = A170 & \new_[16966]_ ;
  assign \new_[16971]_  = ~A200 & ~A199;
  assign \new_[16972]_  = A166 & \new_[16971]_ ;
  assign \new_[16973]_  = \new_[16972]_  & \new_[16967]_ ;
  assign \new_[16977]_  = ~A233 & A232;
  assign \new_[16978]_  = ~A202 & \new_[16977]_ ;
  assign \new_[16981]_  = A236 & ~A235;
  assign \new_[16984]_  = A300 & A299;
  assign \new_[16985]_  = \new_[16984]_  & \new_[16981]_ ;
  assign \new_[16986]_  = \new_[16985]_  & \new_[16978]_ ;
  assign \new_[16990]_  = ~A167 & A168;
  assign \new_[16991]_  = A170 & \new_[16990]_ ;
  assign \new_[16995]_  = ~A200 & ~A199;
  assign \new_[16996]_  = A166 & \new_[16995]_ ;
  assign \new_[16997]_  = \new_[16996]_  & \new_[16991]_ ;
  assign \new_[17001]_  = ~A233 & A232;
  assign \new_[17002]_  = ~A202 & \new_[17001]_ ;
  assign \new_[17005]_  = A236 & ~A235;
  assign \new_[17008]_  = A300 & A298;
  assign \new_[17009]_  = \new_[17008]_  & \new_[17005]_ ;
  assign \new_[17010]_  = \new_[17009]_  & \new_[17002]_ ;
  assign \new_[17014]_  = ~A167 & A168;
  assign \new_[17015]_  = A170 & \new_[17014]_ ;
  assign \new_[17019]_  = ~A200 & ~A199;
  assign \new_[17020]_  = A166 & \new_[17019]_ ;
  assign \new_[17021]_  = \new_[17020]_  & \new_[17015]_ ;
  assign \new_[17025]_  = ~A233 & A232;
  assign \new_[17026]_  = ~A202 & \new_[17025]_ ;
  assign \new_[17029]_  = A236 & ~A235;
  assign \new_[17032]_  = A267 & A265;
  assign \new_[17033]_  = \new_[17032]_  & \new_[17029]_ ;
  assign \new_[17034]_  = \new_[17033]_  & \new_[17026]_ ;
  assign \new_[17038]_  = ~A167 & A168;
  assign \new_[17039]_  = A170 & \new_[17038]_ ;
  assign \new_[17043]_  = ~A200 & ~A199;
  assign \new_[17044]_  = A166 & \new_[17043]_ ;
  assign \new_[17045]_  = \new_[17044]_  & \new_[17039]_ ;
  assign \new_[17049]_  = ~A233 & A232;
  assign \new_[17050]_  = ~A202 & \new_[17049]_ ;
  assign \new_[17053]_  = A236 & ~A235;
  assign \new_[17056]_  = A267 & A266;
  assign \new_[17057]_  = \new_[17056]_  & \new_[17053]_ ;
  assign \new_[17058]_  = \new_[17057]_  & \new_[17050]_ ;
  assign \new_[17062]_  = ~A167 & A168;
  assign \new_[17063]_  = A170 & \new_[17062]_ ;
  assign \new_[17067]_  = ~A200 & ~A199;
  assign \new_[17068]_  = A166 & \new_[17067]_ ;
  assign \new_[17069]_  = \new_[17068]_  & \new_[17063]_ ;
  assign \new_[17073]_  = ~A233 & ~A232;
  assign \new_[17074]_  = ~A202 & \new_[17073]_ ;
  assign \new_[17077]_  = ~A236 & A235;
  assign \new_[17080]_  = A300 & A299;
  assign \new_[17081]_  = \new_[17080]_  & \new_[17077]_ ;
  assign \new_[17082]_  = \new_[17081]_  & \new_[17074]_ ;
  assign \new_[17086]_  = ~A167 & A168;
  assign \new_[17087]_  = A170 & \new_[17086]_ ;
  assign \new_[17091]_  = ~A200 & ~A199;
  assign \new_[17092]_  = A166 & \new_[17091]_ ;
  assign \new_[17093]_  = \new_[17092]_  & \new_[17087]_ ;
  assign \new_[17097]_  = ~A233 & ~A232;
  assign \new_[17098]_  = ~A202 & \new_[17097]_ ;
  assign \new_[17101]_  = ~A236 & A235;
  assign \new_[17104]_  = A300 & A298;
  assign \new_[17105]_  = \new_[17104]_  & \new_[17101]_ ;
  assign \new_[17106]_  = \new_[17105]_  & \new_[17098]_ ;
  assign \new_[17110]_  = ~A167 & A168;
  assign \new_[17111]_  = A170 & \new_[17110]_ ;
  assign \new_[17115]_  = ~A200 & ~A199;
  assign \new_[17116]_  = A166 & \new_[17115]_ ;
  assign \new_[17117]_  = \new_[17116]_  & \new_[17111]_ ;
  assign \new_[17121]_  = ~A233 & ~A232;
  assign \new_[17122]_  = ~A202 & \new_[17121]_ ;
  assign \new_[17125]_  = ~A236 & A235;
  assign \new_[17128]_  = A267 & A265;
  assign \new_[17129]_  = \new_[17128]_  & \new_[17125]_ ;
  assign \new_[17130]_  = \new_[17129]_  & \new_[17122]_ ;
  assign \new_[17134]_  = ~A167 & A168;
  assign \new_[17135]_  = A170 & \new_[17134]_ ;
  assign \new_[17139]_  = ~A200 & ~A199;
  assign \new_[17140]_  = A166 & \new_[17139]_ ;
  assign \new_[17141]_  = \new_[17140]_  & \new_[17135]_ ;
  assign \new_[17145]_  = ~A233 & ~A232;
  assign \new_[17146]_  = ~A202 & \new_[17145]_ ;
  assign \new_[17149]_  = ~A236 & A235;
  assign \new_[17152]_  = A267 & A266;
  assign \new_[17153]_  = \new_[17152]_  & \new_[17149]_ ;
  assign \new_[17154]_  = \new_[17153]_  & \new_[17146]_ ;
  assign \new_[17158]_  = ~A167 & A168;
  assign \new_[17159]_  = A170 & \new_[17158]_ ;
  assign \new_[17163]_  = ~A200 & ~A199;
  assign \new_[17164]_  = A166 & \new_[17163]_ ;
  assign \new_[17165]_  = \new_[17164]_  & \new_[17159]_ ;
  assign \new_[17169]_  = A234 & A232;
  assign \new_[17170]_  = A203 & \new_[17169]_ ;
  assign \new_[17173]_  = A299 & A298;
  assign \new_[17176]_  = ~A302 & A301;
  assign \new_[17177]_  = \new_[17176]_  & \new_[17173]_ ;
  assign \new_[17178]_  = \new_[17177]_  & \new_[17170]_ ;
  assign \new_[17182]_  = ~A167 & A168;
  assign \new_[17183]_  = A170 & \new_[17182]_ ;
  assign \new_[17187]_  = ~A200 & ~A199;
  assign \new_[17188]_  = A166 & \new_[17187]_ ;
  assign \new_[17189]_  = \new_[17188]_  & \new_[17183]_ ;
  assign \new_[17193]_  = A234 & A232;
  assign \new_[17194]_  = A203 & \new_[17193]_ ;
  assign \new_[17197]_  = ~A299 & A298;
  assign \new_[17200]_  = A302 & ~A301;
  assign \new_[17201]_  = \new_[17200]_  & \new_[17197]_ ;
  assign \new_[17202]_  = \new_[17201]_  & \new_[17194]_ ;
  assign \new_[17206]_  = ~A167 & A168;
  assign \new_[17207]_  = A170 & \new_[17206]_ ;
  assign \new_[17211]_  = ~A200 & ~A199;
  assign \new_[17212]_  = A166 & \new_[17211]_ ;
  assign \new_[17213]_  = \new_[17212]_  & \new_[17207]_ ;
  assign \new_[17217]_  = A234 & A232;
  assign \new_[17218]_  = A203 & \new_[17217]_ ;
  assign \new_[17221]_  = A299 & ~A298;
  assign \new_[17224]_  = A302 & ~A301;
  assign \new_[17225]_  = \new_[17224]_  & \new_[17221]_ ;
  assign \new_[17226]_  = \new_[17225]_  & \new_[17218]_ ;
  assign \new_[17230]_  = ~A167 & A168;
  assign \new_[17231]_  = A170 & \new_[17230]_ ;
  assign \new_[17235]_  = ~A200 & ~A199;
  assign \new_[17236]_  = A166 & \new_[17235]_ ;
  assign \new_[17237]_  = \new_[17236]_  & \new_[17231]_ ;
  assign \new_[17241]_  = A234 & A232;
  assign \new_[17242]_  = A203 & \new_[17241]_ ;
  assign \new_[17245]_  = ~A299 & ~A298;
  assign \new_[17248]_  = ~A302 & A301;
  assign \new_[17249]_  = \new_[17248]_  & \new_[17245]_ ;
  assign \new_[17250]_  = \new_[17249]_  & \new_[17242]_ ;
  assign \new_[17254]_  = ~A167 & A168;
  assign \new_[17255]_  = A170 & \new_[17254]_ ;
  assign \new_[17259]_  = ~A200 & ~A199;
  assign \new_[17260]_  = A166 & \new_[17259]_ ;
  assign \new_[17261]_  = \new_[17260]_  & \new_[17255]_ ;
  assign \new_[17265]_  = A234 & A232;
  assign \new_[17266]_  = A203 & \new_[17265]_ ;
  assign \new_[17269]_  = A266 & A265;
  assign \new_[17272]_  = ~A269 & A268;
  assign \new_[17273]_  = \new_[17272]_  & \new_[17269]_ ;
  assign \new_[17274]_  = \new_[17273]_  & \new_[17266]_ ;
  assign \new_[17278]_  = ~A167 & A168;
  assign \new_[17279]_  = A170 & \new_[17278]_ ;
  assign \new_[17283]_  = ~A200 & ~A199;
  assign \new_[17284]_  = A166 & \new_[17283]_ ;
  assign \new_[17285]_  = \new_[17284]_  & \new_[17279]_ ;
  assign \new_[17289]_  = A234 & A232;
  assign \new_[17290]_  = A203 & \new_[17289]_ ;
  assign \new_[17293]_  = A266 & ~A265;
  assign \new_[17296]_  = A269 & ~A268;
  assign \new_[17297]_  = \new_[17296]_  & \new_[17293]_ ;
  assign \new_[17298]_  = \new_[17297]_  & \new_[17290]_ ;
  assign \new_[17302]_  = ~A167 & A168;
  assign \new_[17303]_  = A170 & \new_[17302]_ ;
  assign \new_[17307]_  = ~A200 & ~A199;
  assign \new_[17308]_  = A166 & \new_[17307]_ ;
  assign \new_[17309]_  = \new_[17308]_  & \new_[17303]_ ;
  assign \new_[17313]_  = A234 & A232;
  assign \new_[17314]_  = A203 & \new_[17313]_ ;
  assign \new_[17317]_  = ~A266 & A265;
  assign \new_[17320]_  = A269 & ~A268;
  assign \new_[17321]_  = \new_[17320]_  & \new_[17317]_ ;
  assign \new_[17322]_  = \new_[17321]_  & \new_[17314]_ ;
  assign \new_[17326]_  = ~A167 & A168;
  assign \new_[17327]_  = A170 & \new_[17326]_ ;
  assign \new_[17331]_  = ~A200 & ~A199;
  assign \new_[17332]_  = A166 & \new_[17331]_ ;
  assign \new_[17333]_  = \new_[17332]_  & \new_[17327]_ ;
  assign \new_[17337]_  = A234 & A232;
  assign \new_[17338]_  = A203 & \new_[17337]_ ;
  assign \new_[17341]_  = ~A266 & ~A265;
  assign \new_[17344]_  = ~A269 & A268;
  assign \new_[17345]_  = \new_[17344]_  & \new_[17341]_ ;
  assign \new_[17346]_  = \new_[17345]_  & \new_[17338]_ ;
  assign \new_[17350]_  = ~A167 & A168;
  assign \new_[17351]_  = A170 & \new_[17350]_ ;
  assign \new_[17355]_  = ~A200 & ~A199;
  assign \new_[17356]_  = A166 & \new_[17355]_ ;
  assign \new_[17357]_  = \new_[17356]_  & \new_[17351]_ ;
  assign \new_[17361]_  = A234 & A233;
  assign \new_[17362]_  = A203 & \new_[17361]_ ;
  assign \new_[17365]_  = A299 & A298;
  assign \new_[17368]_  = ~A302 & A301;
  assign \new_[17369]_  = \new_[17368]_  & \new_[17365]_ ;
  assign \new_[17370]_  = \new_[17369]_  & \new_[17362]_ ;
  assign \new_[17374]_  = ~A167 & A168;
  assign \new_[17375]_  = A170 & \new_[17374]_ ;
  assign \new_[17379]_  = ~A200 & ~A199;
  assign \new_[17380]_  = A166 & \new_[17379]_ ;
  assign \new_[17381]_  = \new_[17380]_  & \new_[17375]_ ;
  assign \new_[17385]_  = A234 & A233;
  assign \new_[17386]_  = A203 & \new_[17385]_ ;
  assign \new_[17389]_  = ~A299 & A298;
  assign \new_[17392]_  = A302 & ~A301;
  assign \new_[17393]_  = \new_[17392]_  & \new_[17389]_ ;
  assign \new_[17394]_  = \new_[17393]_  & \new_[17386]_ ;
  assign \new_[17398]_  = ~A167 & A168;
  assign \new_[17399]_  = A170 & \new_[17398]_ ;
  assign \new_[17403]_  = ~A200 & ~A199;
  assign \new_[17404]_  = A166 & \new_[17403]_ ;
  assign \new_[17405]_  = \new_[17404]_  & \new_[17399]_ ;
  assign \new_[17409]_  = A234 & A233;
  assign \new_[17410]_  = A203 & \new_[17409]_ ;
  assign \new_[17413]_  = A299 & ~A298;
  assign \new_[17416]_  = A302 & ~A301;
  assign \new_[17417]_  = \new_[17416]_  & \new_[17413]_ ;
  assign \new_[17418]_  = \new_[17417]_  & \new_[17410]_ ;
  assign \new_[17422]_  = ~A167 & A168;
  assign \new_[17423]_  = A170 & \new_[17422]_ ;
  assign \new_[17427]_  = ~A200 & ~A199;
  assign \new_[17428]_  = A166 & \new_[17427]_ ;
  assign \new_[17429]_  = \new_[17428]_  & \new_[17423]_ ;
  assign \new_[17433]_  = A234 & A233;
  assign \new_[17434]_  = A203 & \new_[17433]_ ;
  assign \new_[17437]_  = ~A299 & ~A298;
  assign \new_[17440]_  = ~A302 & A301;
  assign \new_[17441]_  = \new_[17440]_  & \new_[17437]_ ;
  assign \new_[17442]_  = \new_[17441]_  & \new_[17434]_ ;
  assign \new_[17446]_  = ~A167 & A168;
  assign \new_[17447]_  = A170 & \new_[17446]_ ;
  assign \new_[17451]_  = ~A200 & ~A199;
  assign \new_[17452]_  = A166 & \new_[17451]_ ;
  assign \new_[17453]_  = \new_[17452]_  & \new_[17447]_ ;
  assign \new_[17457]_  = A234 & A233;
  assign \new_[17458]_  = A203 & \new_[17457]_ ;
  assign \new_[17461]_  = A266 & A265;
  assign \new_[17464]_  = ~A269 & A268;
  assign \new_[17465]_  = \new_[17464]_  & \new_[17461]_ ;
  assign \new_[17466]_  = \new_[17465]_  & \new_[17458]_ ;
  assign \new_[17470]_  = ~A167 & A168;
  assign \new_[17471]_  = A170 & \new_[17470]_ ;
  assign \new_[17475]_  = ~A200 & ~A199;
  assign \new_[17476]_  = A166 & \new_[17475]_ ;
  assign \new_[17477]_  = \new_[17476]_  & \new_[17471]_ ;
  assign \new_[17481]_  = A234 & A233;
  assign \new_[17482]_  = A203 & \new_[17481]_ ;
  assign \new_[17485]_  = A266 & ~A265;
  assign \new_[17488]_  = A269 & ~A268;
  assign \new_[17489]_  = \new_[17488]_  & \new_[17485]_ ;
  assign \new_[17490]_  = \new_[17489]_  & \new_[17482]_ ;
  assign \new_[17494]_  = ~A167 & A168;
  assign \new_[17495]_  = A170 & \new_[17494]_ ;
  assign \new_[17499]_  = ~A200 & ~A199;
  assign \new_[17500]_  = A166 & \new_[17499]_ ;
  assign \new_[17501]_  = \new_[17500]_  & \new_[17495]_ ;
  assign \new_[17505]_  = A234 & A233;
  assign \new_[17506]_  = A203 & \new_[17505]_ ;
  assign \new_[17509]_  = ~A266 & A265;
  assign \new_[17512]_  = A269 & ~A268;
  assign \new_[17513]_  = \new_[17512]_  & \new_[17509]_ ;
  assign \new_[17514]_  = \new_[17513]_  & \new_[17506]_ ;
  assign \new_[17518]_  = ~A167 & A168;
  assign \new_[17519]_  = A170 & \new_[17518]_ ;
  assign \new_[17523]_  = ~A200 & ~A199;
  assign \new_[17524]_  = A166 & \new_[17523]_ ;
  assign \new_[17525]_  = \new_[17524]_  & \new_[17519]_ ;
  assign \new_[17529]_  = A234 & A233;
  assign \new_[17530]_  = A203 & \new_[17529]_ ;
  assign \new_[17533]_  = ~A266 & ~A265;
  assign \new_[17536]_  = ~A269 & A268;
  assign \new_[17537]_  = \new_[17536]_  & \new_[17533]_ ;
  assign \new_[17538]_  = \new_[17537]_  & \new_[17530]_ ;
  assign \new_[17542]_  = ~A167 & A168;
  assign \new_[17543]_  = A170 & \new_[17542]_ ;
  assign \new_[17547]_  = ~A200 & ~A199;
  assign \new_[17548]_  = A166 & \new_[17547]_ ;
  assign \new_[17549]_  = \new_[17548]_  & \new_[17543]_ ;
  assign \new_[17553]_  = A233 & A232;
  assign \new_[17554]_  = A203 & \new_[17553]_ ;
  assign \new_[17557]_  = ~A236 & A235;
  assign \new_[17560]_  = A300 & A299;
  assign \new_[17561]_  = \new_[17560]_  & \new_[17557]_ ;
  assign \new_[17562]_  = \new_[17561]_  & \new_[17554]_ ;
  assign \new_[17566]_  = ~A167 & A168;
  assign \new_[17567]_  = A170 & \new_[17566]_ ;
  assign \new_[17571]_  = ~A200 & ~A199;
  assign \new_[17572]_  = A166 & \new_[17571]_ ;
  assign \new_[17573]_  = \new_[17572]_  & \new_[17567]_ ;
  assign \new_[17577]_  = A233 & A232;
  assign \new_[17578]_  = A203 & \new_[17577]_ ;
  assign \new_[17581]_  = ~A236 & A235;
  assign \new_[17584]_  = A300 & A298;
  assign \new_[17585]_  = \new_[17584]_  & \new_[17581]_ ;
  assign \new_[17586]_  = \new_[17585]_  & \new_[17578]_ ;
  assign \new_[17590]_  = ~A167 & A168;
  assign \new_[17591]_  = A170 & \new_[17590]_ ;
  assign \new_[17595]_  = ~A200 & ~A199;
  assign \new_[17596]_  = A166 & \new_[17595]_ ;
  assign \new_[17597]_  = \new_[17596]_  & \new_[17591]_ ;
  assign \new_[17601]_  = A233 & A232;
  assign \new_[17602]_  = A203 & \new_[17601]_ ;
  assign \new_[17605]_  = ~A236 & A235;
  assign \new_[17608]_  = A267 & A265;
  assign \new_[17609]_  = \new_[17608]_  & \new_[17605]_ ;
  assign \new_[17610]_  = \new_[17609]_  & \new_[17602]_ ;
  assign \new_[17614]_  = ~A167 & A168;
  assign \new_[17615]_  = A170 & \new_[17614]_ ;
  assign \new_[17619]_  = ~A200 & ~A199;
  assign \new_[17620]_  = A166 & \new_[17619]_ ;
  assign \new_[17621]_  = \new_[17620]_  & \new_[17615]_ ;
  assign \new_[17625]_  = A233 & A232;
  assign \new_[17626]_  = A203 & \new_[17625]_ ;
  assign \new_[17629]_  = ~A236 & A235;
  assign \new_[17632]_  = A267 & A266;
  assign \new_[17633]_  = \new_[17632]_  & \new_[17629]_ ;
  assign \new_[17634]_  = \new_[17633]_  & \new_[17626]_ ;
  assign \new_[17638]_  = ~A167 & A168;
  assign \new_[17639]_  = A170 & \new_[17638]_ ;
  assign \new_[17643]_  = ~A200 & ~A199;
  assign \new_[17644]_  = A166 & \new_[17643]_ ;
  assign \new_[17645]_  = \new_[17644]_  & \new_[17639]_ ;
  assign \new_[17649]_  = A233 & ~A232;
  assign \new_[17650]_  = A203 & \new_[17649]_ ;
  assign \new_[17653]_  = A236 & ~A235;
  assign \new_[17656]_  = A300 & A299;
  assign \new_[17657]_  = \new_[17656]_  & \new_[17653]_ ;
  assign \new_[17658]_  = \new_[17657]_  & \new_[17650]_ ;
  assign \new_[17662]_  = ~A167 & A168;
  assign \new_[17663]_  = A170 & \new_[17662]_ ;
  assign \new_[17667]_  = ~A200 & ~A199;
  assign \new_[17668]_  = A166 & \new_[17667]_ ;
  assign \new_[17669]_  = \new_[17668]_  & \new_[17663]_ ;
  assign \new_[17673]_  = A233 & ~A232;
  assign \new_[17674]_  = A203 & \new_[17673]_ ;
  assign \new_[17677]_  = A236 & ~A235;
  assign \new_[17680]_  = A300 & A298;
  assign \new_[17681]_  = \new_[17680]_  & \new_[17677]_ ;
  assign \new_[17682]_  = \new_[17681]_  & \new_[17674]_ ;
  assign \new_[17686]_  = ~A167 & A168;
  assign \new_[17687]_  = A170 & \new_[17686]_ ;
  assign \new_[17691]_  = ~A200 & ~A199;
  assign \new_[17692]_  = A166 & \new_[17691]_ ;
  assign \new_[17693]_  = \new_[17692]_  & \new_[17687]_ ;
  assign \new_[17697]_  = A233 & ~A232;
  assign \new_[17698]_  = A203 & \new_[17697]_ ;
  assign \new_[17701]_  = A236 & ~A235;
  assign \new_[17704]_  = A267 & A265;
  assign \new_[17705]_  = \new_[17704]_  & \new_[17701]_ ;
  assign \new_[17706]_  = \new_[17705]_  & \new_[17698]_ ;
  assign \new_[17710]_  = ~A167 & A168;
  assign \new_[17711]_  = A170 & \new_[17710]_ ;
  assign \new_[17715]_  = ~A200 & ~A199;
  assign \new_[17716]_  = A166 & \new_[17715]_ ;
  assign \new_[17717]_  = \new_[17716]_  & \new_[17711]_ ;
  assign \new_[17721]_  = A233 & ~A232;
  assign \new_[17722]_  = A203 & \new_[17721]_ ;
  assign \new_[17725]_  = A236 & ~A235;
  assign \new_[17728]_  = A267 & A266;
  assign \new_[17729]_  = \new_[17728]_  & \new_[17725]_ ;
  assign \new_[17730]_  = \new_[17729]_  & \new_[17722]_ ;
  assign \new_[17734]_  = ~A167 & A168;
  assign \new_[17735]_  = A170 & \new_[17734]_ ;
  assign \new_[17739]_  = ~A200 & ~A199;
  assign \new_[17740]_  = A166 & \new_[17739]_ ;
  assign \new_[17741]_  = \new_[17740]_  & \new_[17735]_ ;
  assign \new_[17745]_  = ~A233 & A232;
  assign \new_[17746]_  = A203 & \new_[17745]_ ;
  assign \new_[17749]_  = A236 & ~A235;
  assign \new_[17752]_  = A300 & A299;
  assign \new_[17753]_  = \new_[17752]_  & \new_[17749]_ ;
  assign \new_[17754]_  = \new_[17753]_  & \new_[17746]_ ;
  assign \new_[17758]_  = ~A167 & A168;
  assign \new_[17759]_  = A170 & \new_[17758]_ ;
  assign \new_[17763]_  = ~A200 & ~A199;
  assign \new_[17764]_  = A166 & \new_[17763]_ ;
  assign \new_[17765]_  = \new_[17764]_  & \new_[17759]_ ;
  assign \new_[17769]_  = ~A233 & A232;
  assign \new_[17770]_  = A203 & \new_[17769]_ ;
  assign \new_[17773]_  = A236 & ~A235;
  assign \new_[17776]_  = A300 & A298;
  assign \new_[17777]_  = \new_[17776]_  & \new_[17773]_ ;
  assign \new_[17778]_  = \new_[17777]_  & \new_[17770]_ ;
  assign \new_[17782]_  = ~A167 & A168;
  assign \new_[17783]_  = A170 & \new_[17782]_ ;
  assign \new_[17787]_  = ~A200 & ~A199;
  assign \new_[17788]_  = A166 & \new_[17787]_ ;
  assign \new_[17789]_  = \new_[17788]_  & \new_[17783]_ ;
  assign \new_[17793]_  = ~A233 & A232;
  assign \new_[17794]_  = A203 & \new_[17793]_ ;
  assign \new_[17797]_  = A236 & ~A235;
  assign \new_[17800]_  = A267 & A265;
  assign \new_[17801]_  = \new_[17800]_  & \new_[17797]_ ;
  assign \new_[17802]_  = \new_[17801]_  & \new_[17794]_ ;
  assign \new_[17806]_  = ~A167 & A168;
  assign \new_[17807]_  = A170 & \new_[17806]_ ;
  assign \new_[17811]_  = ~A200 & ~A199;
  assign \new_[17812]_  = A166 & \new_[17811]_ ;
  assign \new_[17813]_  = \new_[17812]_  & \new_[17807]_ ;
  assign \new_[17817]_  = ~A233 & A232;
  assign \new_[17818]_  = A203 & \new_[17817]_ ;
  assign \new_[17821]_  = A236 & ~A235;
  assign \new_[17824]_  = A267 & A266;
  assign \new_[17825]_  = \new_[17824]_  & \new_[17821]_ ;
  assign \new_[17826]_  = \new_[17825]_  & \new_[17818]_ ;
  assign \new_[17830]_  = ~A167 & A168;
  assign \new_[17831]_  = A170 & \new_[17830]_ ;
  assign \new_[17835]_  = ~A200 & ~A199;
  assign \new_[17836]_  = A166 & \new_[17835]_ ;
  assign \new_[17837]_  = \new_[17836]_  & \new_[17831]_ ;
  assign \new_[17841]_  = ~A233 & ~A232;
  assign \new_[17842]_  = A203 & \new_[17841]_ ;
  assign \new_[17845]_  = ~A236 & A235;
  assign \new_[17848]_  = A300 & A299;
  assign \new_[17849]_  = \new_[17848]_  & \new_[17845]_ ;
  assign \new_[17850]_  = \new_[17849]_  & \new_[17842]_ ;
  assign \new_[17854]_  = ~A167 & A168;
  assign \new_[17855]_  = A170 & \new_[17854]_ ;
  assign \new_[17859]_  = ~A200 & ~A199;
  assign \new_[17860]_  = A166 & \new_[17859]_ ;
  assign \new_[17861]_  = \new_[17860]_  & \new_[17855]_ ;
  assign \new_[17865]_  = ~A233 & ~A232;
  assign \new_[17866]_  = A203 & \new_[17865]_ ;
  assign \new_[17869]_  = ~A236 & A235;
  assign \new_[17872]_  = A300 & A298;
  assign \new_[17873]_  = \new_[17872]_  & \new_[17869]_ ;
  assign \new_[17874]_  = \new_[17873]_  & \new_[17866]_ ;
  assign \new_[17878]_  = ~A167 & A168;
  assign \new_[17879]_  = A170 & \new_[17878]_ ;
  assign \new_[17883]_  = ~A200 & ~A199;
  assign \new_[17884]_  = A166 & \new_[17883]_ ;
  assign \new_[17885]_  = \new_[17884]_  & \new_[17879]_ ;
  assign \new_[17889]_  = ~A233 & ~A232;
  assign \new_[17890]_  = A203 & \new_[17889]_ ;
  assign \new_[17893]_  = ~A236 & A235;
  assign \new_[17896]_  = A267 & A265;
  assign \new_[17897]_  = \new_[17896]_  & \new_[17893]_ ;
  assign \new_[17898]_  = \new_[17897]_  & \new_[17890]_ ;
  assign \new_[17902]_  = ~A167 & A168;
  assign \new_[17903]_  = A170 & \new_[17902]_ ;
  assign \new_[17907]_  = ~A200 & ~A199;
  assign \new_[17908]_  = A166 & \new_[17907]_ ;
  assign \new_[17909]_  = \new_[17908]_  & \new_[17903]_ ;
  assign \new_[17913]_  = ~A233 & ~A232;
  assign \new_[17914]_  = A203 & \new_[17913]_ ;
  assign \new_[17917]_  = ~A236 & A235;
  assign \new_[17920]_  = A267 & A266;
  assign \new_[17921]_  = \new_[17920]_  & \new_[17917]_ ;
  assign \new_[17922]_  = \new_[17921]_  & \new_[17914]_ ;
  assign \new_[17926]_  = ~A167 & A168;
  assign \new_[17927]_  = A169 & \new_[17926]_ ;
  assign \new_[17931]_  = ~A200 & ~A199;
  assign \new_[17932]_  = A166 & \new_[17931]_ ;
  assign \new_[17933]_  = \new_[17932]_  & \new_[17927]_ ;
  assign \new_[17937]_  = A234 & A232;
  assign \new_[17938]_  = ~A202 & \new_[17937]_ ;
  assign \new_[17941]_  = A299 & A298;
  assign \new_[17944]_  = ~A302 & A301;
  assign \new_[17945]_  = \new_[17944]_  & \new_[17941]_ ;
  assign \new_[17946]_  = \new_[17945]_  & \new_[17938]_ ;
  assign \new_[17950]_  = ~A167 & A168;
  assign \new_[17951]_  = A169 & \new_[17950]_ ;
  assign \new_[17955]_  = ~A200 & ~A199;
  assign \new_[17956]_  = A166 & \new_[17955]_ ;
  assign \new_[17957]_  = \new_[17956]_  & \new_[17951]_ ;
  assign \new_[17961]_  = A234 & A232;
  assign \new_[17962]_  = ~A202 & \new_[17961]_ ;
  assign \new_[17965]_  = ~A299 & A298;
  assign \new_[17968]_  = A302 & ~A301;
  assign \new_[17969]_  = \new_[17968]_  & \new_[17965]_ ;
  assign \new_[17970]_  = \new_[17969]_  & \new_[17962]_ ;
  assign \new_[17974]_  = ~A167 & A168;
  assign \new_[17975]_  = A169 & \new_[17974]_ ;
  assign \new_[17979]_  = ~A200 & ~A199;
  assign \new_[17980]_  = A166 & \new_[17979]_ ;
  assign \new_[17981]_  = \new_[17980]_  & \new_[17975]_ ;
  assign \new_[17985]_  = A234 & A232;
  assign \new_[17986]_  = ~A202 & \new_[17985]_ ;
  assign \new_[17989]_  = A299 & ~A298;
  assign \new_[17992]_  = A302 & ~A301;
  assign \new_[17993]_  = \new_[17992]_  & \new_[17989]_ ;
  assign \new_[17994]_  = \new_[17993]_  & \new_[17986]_ ;
  assign \new_[17998]_  = ~A167 & A168;
  assign \new_[17999]_  = A169 & \new_[17998]_ ;
  assign \new_[18003]_  = ~A200 & ~A199;
  assign \new_[18004]_  = A166 & \new_[18003]_ ;
  assign \new_[18005]_  = \new_[18004]_  & \new_[17999]_ ;
  assign \new_[18009]_  = A234 & A232;
  assign \new_[18010]_  = ~A202 & \new_[18009]_ ;
  assign \new_[18013]_  = ~A299 & ~A298;
  assign \new_[18016]_  = ~A302 & A301;
  assign \new_[18017]_  = \new_[18016]_  & \new_[18013]_ ;
  assign \new_[18018]_  = \new_[18017]_  & \new_[18010]_ ;
  assign \new_[18022]_  = ~A167 & A168;
  assign \new_[18023]_  = A169 & \new_[18022]_ ;
  assign \new_[18027]_  = ~A200 & ~A199;
  assign \new_[18028]_  = A166 & \new_[18027]_ ;
  assign \new_[18029]_  = \new_[18028]_  & \new_[18023]_ ;
  assign \new_[18033]_  = A234 & A232;
  assign \new_[18034]_  = ~A202 & \new_[18033]_ ;
  assign \new_[18037]_  = A266 & A265;
  assign \new_[18040]_  = ~A269 & A268;
  assign \new_[18041]_  = \new_[18040]_  & \new_[18037]_ ;
  assign \new_[18042]_  = \new_[18041]_  & \new_[18034]_ ;
  assign \new_[18046]_  = ~A167 & A168;
  assign \new_[18047]_  = A169 & \new_[18046]_ ;
  assign \new_[18051]_  = ~A200 & ~A199;
  assign \new_[18052]_  = A166 & \new_[18051]_ ;
  assign \new_[18053]_  = \new_[18052]_  & \new_[18047]_ ;
  assign \new_[18057]_  = A234 & A232;
  assign \new_[18058]_  = ~A202 & \new_[18057]_ ;
  assign \new_[18061]_  = A266 & ~A265;
  assign \new_[18064]_  = A269 & ~A268;
  assign \new_[18065]_  = \new_[18064]_  & \new_[18061]_ ;
  assign \new_[18066]_  = \new_[18065]_  & \new_[18058]_ ;
  assign \new_[18070]_  = ~A167 & A168;
  assign \new_[18071]_  = A169 & \new_[18070]_ ;
  assign \new_[18075]_  = ~A200 & ~A199;
  assign \new_[18076]_  = A166 & \new_[18075]_ ;
  assign \new_[18077]_  = \new_[18076]_  & \new_[18071]_ ;
  assign \new_[18081]_  = A234 & A232;
  assign \new_[18082]_  = ~A202 & \new_[18081]_ ;
  assign \new_[18085]_  = ~A266 & A265;
  assign \new_[18088]_  = A269 & ~A268;
  assign \new_[18089]_  = \new_[18088]_  & \new_[18085]_ ;
  assign \new_[18090]_  = \new_[18089]_  & \new_[18082]_ ;
  assign \new_[18094]_  = ~A167 & A168;
  assign \new_[18095]_  = A169 & \new_[18094]_ ;
  assign \new_[18099]_  = ~A200 & ~A199;
  assign \new_[18100]_  = A166 & \new_[18099]_ ;
  assign \new_[18101]_  = \new_[18100]_  & \new_[18095]_ ;
  assign \new_[18105]_  = A234 & A232;
  assign \new_[18106]_  = ~A202 & \new_[18105]_ ;
  assign \new_[18109]_  = ~A266 & ~A265;
  assign \new_[18112]_  = ~A269 & A268;
  assign \new_[18113]_  = \new_[18112]_  & \new_[18109]_ ;
  assign \new_[18114]_  = \new_[18113]_  & \new_[18106]_ ;
  assign \new_[18118]_  = ~A167 & A168;
  assign \new_[18119]_  = A169 & \new_[18118]_ ;
  assign \new_[18123]_  = ~A200 & ~A199;
  assign \new_[18124]_  = A166 & \new_[18123]_ ;
  assign \new_[18125]_  = \new_[18124]_  & \new_[18119]_ ;
  assign \new_[18129]_  = A234 & A233;
  assign \new_[18130]_  = ~A202 & \new_[18129]_ ;
  assign \new_[18133]_  = A299 & A298;
  assign \new_[18136]_  = ~A302 & A301;
  assign \new_[18137]_  = \new_[18136]_  & \new_[18133]_ ;
  assign \new_[18138]_  = \new_[18137]_  & \new_[18130]_ ;
  assign \new_[18142]_  = ~A167 & A168;
  assign \new_[18143]_  = A169 & \new_[18142]_ ;
  assign \new_[18147]_  = ~A200 & ~A199;
  assign \new_[18148]_  = A166 & \new_[18147]_ ;
  assign \new_[18149]_  = \new_[18148]_  & \new_[18143]_ ;
  assign \new_[18153]_  = A234 & A233;
  assign \new_[18154]_  = ~A202 & \new_[18153]_ ;
  assign \new_[18157]_  = ~A299 & A298;
  assign \new_[18160]_  = A302 & ~A301;
  assign \new_[18161]_  = \new_[18160]_  & \new_[18157]_ ;
  assign \new_[18162]_  = \new_[18161]_  & \new_[18154]_ ;
  assign \new_[18166]_  = ~A167 & A168;
  assign \new_[18167]_  = A169 & \new_[18166]_ ;
  assign \new_[18171]_  = ~A200 & ~A199;
  assign \new_[18172]_  = A166 & \new_[18171]_ ;
  assign \new_[18173]_  = \new_[18172]_  & \new_[18167]_ ;
  assign \new_[18177]_  = A234 & A233;
  assign \new_[18178]_  = ~A202 & \new_[18177]_ ;
  assign \new_[18181]_  = A299 & ~A298;
  assign \new_[18184]_  = A302 & ~A301;
  assign \new_[18185]_  = \new_[18184]_  & \new_[18181]_ ;
  assign \new_[18186]_  = \new_[18185]_  & \new_[18178]_ ;
  assign \new_[18190]_  = ~A167 & A168;
  assign \new_[18191]_  = A169 & \new_[18190]_ ;
  assign \new_[18195]_  = ~A200 & ~A199;
  assign \new_[18196]_  = A166 & \new_[18195]_ ;
  assign \new_[18197]_  = \new_[18196]_  & \new_[18191]_ ;
  assign \new_[18201]_  = A234 & A233;
  assign \new_[18202]_  = ~A202 & \new_[18201]_ ;
  assign \new_[18205]_  = ~A299 & ~A298;
  assign \new_[18208]_  = ~A302 & A301;
  assign \new_[18209]_  = \new_[18208]_  & \new_[18205]_ ;
  assign \new_[18210]_  = \new_[18209]_  & \new_[18202]_ ;
  assign \new_[18214]_  = ~A167 & A168;
  assign \new_[18215]_  = A169 & \new_[18214]_ ;
  assign \new_[18219]_  = ~A200 & ~A199;
  assign \new_[18220]_  = A166 & \new_[18219]_ ;
  assign \new_[18221]_  = \new_[18220]_  & \new_[18215]_ ;
  assign \new_[18225]_  = A234 & A233;
  assign \new_[18226]_  = ~A202 & \new_[18225]_ ;
  assign \new_[18229]_  = A266 & A265;
  assign \new_[18232]_  = ~A269 & A268;
  assign \new_[18233]_  = \new_[18232]_  & \new_[18229]_ ;
  assign \new_[18234]_  = \new_[18233]_  & \new_[18226]_ ;
  assign \new_[18238]_  = ~A167 & A168;
  assign \new_[18239]_  = A169 & \new_[18238]_ ;
  assign \new_[18243]_  = ~A200 & ~A199;
  assign \new_[18244]_  = A166 & \new_[18243]_ ;
  assign \new_[18245]_  = \new_[18244]_  & \new_[18239]_ ;
  assign \new_[18249]_  = A234 & A233;
  assign \new_[18250]_  = ~A202 & \new_[18249]_ ;
  assign \new_[18253]_  = A266 & ~A265;
  assign \new_[18256]_  = A269 & ~A268;
  assign \new_[18257]_  = \new_[18256]_  & \new_[18253]_ ;
  assign \new_[18258]_  = \new_[18257]_  & \new_[18250]_ ;
  assign \new_[18262]_  = ~A167 & A168;
  assign \new_[18263]_  = A169 & \new_[18262]_ ;
  assign \new_[18267]_  = ~A200 & ~A199;
  assign \new_[18268]_  = A166 & \new_[18267]_ ;
  assign \new_[18269]_  = \new_[18268]_  & \new_[18263]_ ;
  assign \new_[18273]_  = A234 & A233;
  assign \new_[18274]_  = ~A202 & \new_[18273]_ ;
  assign \new_[18277]_  = ~A266 & A265;
  assign \new_[18280]_  = A269 & ~A268;
  assign \new_[18281]_  = \new_[18280]_  & \new_[18277]_ ;
  assign \new_[18282]_  = \new_[18281]_  & \new_[18274]_ ;
  assign \new_[18286]_  = ~A167 & A168;
  assign \new_[18287]_  = A169 & \new_[18286]_ ;
  assign \new_[18291]_  = ~A200 & ~A199;
  assign \new_[18292]_  = A166 & \new_[18291]_ ;
  assign \new_[18293]_  = \new_[18292]_  & \new_[18287]_ ;
  assign \new_[18297]_  = A234 & A233;
  assign \new_[18298]_  = ~A202 & \new_[18297]_ ;
  assign \new_[18301]_  = ~A266 & ~A265;
  assign \new_[18304]_  = ~A269 & A268;
  assign \new_[18305]_  = \new_[18304]_  & \new_[18301]_ ;
  assign \new_[18306]_  = \new_[18305]_  & \new_[18298]_ ;
  assign \new_[18310]_  = ~A167 & A168;
  assign \new_[18311]_  = A169 & \new_[18310]_ ;
  assign \new_[18315]_  = ~A200 & ~A199;
  assign \new_[18316]_  = A166 & \new_[18315]_ ;
  assign \new_[18317]_  = \new_[18316]_  & \new_[18311]_ ;
  assign \new_[18321]_  = A233 & A232;
  assign \new_[18322]_  = ~A202 & \new_[18321]_ ;
  assign \new_[18325]_  = ~A236 & A235;
  assign \new_[18328]_  = A300 & A299;
  assign \new_[18329]_  = \new_[18328]_  & \new_[18325]_ ;
  assign \new_[18330]_  = \new_[18329]_  & \new_[18322]_ ;
  assign \new_[18334]_  = ~A167 & A168;
  assign \new_[18335]_  = A169 & \new_[18334]_ ;
  assign \new_[18339]_  = ~A200 & ~A199;
  assign \new_[18340]_  = A166 & \new_[18339]_ ;
  assign \new_[18341]_  = \new_[18340]_  & \new_[18335]_ ;
  assign \new_[18345]_  = A233 & A232;
  assign \new_[18346]_  = ~A202 & \new_[18345]_ ;
  assign \new_[18349]_  = ~A236 & A235;
  assign \new_[18352]_  = A300 & A298;
  assign \new_[18353]_  = \new_[18352]_  & \new_[18349]_ ;
  assign \new_[18354]_  = \new_[18353]_  & \new_[18346]_ ;
  assign \new_[18358]_  = ~A167 & A168;
  assign \new_[18359]_  = A169 & \new_[18358]_ ;
  assign \new_[18363]_  = ~A200 & ~A199;
  assign \new_[18364]_  = A166 & \new_[18363]_ ;
  assign \new_[18365]_  = \new_[18364]_  & \new_[18359]_ ;
  assign \new_[18369]_  = A233 & A232;
  assign \new_[18370]_  = ~A202 & \new_[18369]_ ;
  assign \new_[18373]_  = ~A236 & A235;
  assign \new_[18376]_  = A267 & A265;
  assign \new_[18377]_  = \new_[18376]_  & \new_[18373]_ ;
  assign \new_[18378]_  = \new_[18377]_  & \new_[18370]_ ;
  assign \new_[18382]_  = ~A167 & A168;
  assign \new_[18383]_  = A169 & \new_[18382]_ ;
  assign \new_[18387]_  = ~A200 & ~A199;
  assign \new_[18388]_  = A166 & \new_[18387]_ ;
  assign \new_[18389]_  = \new_[18388]_  & \new_[18383]_ ;
  assign \new_[18393]_  = A233 & A232;
  assign \new_[18394]_  = ~A202 & \new_[18393]_ ;
  assign \new_[18397]_  = ~A236 & A235;
  assign \new_[18400]_  = A267 & A266;
  assign \new_[18401]_  = \new_[18400]_  & \new_[18397]_ ;
  assign \new_[18402]_  = \new_[18401]_  & \new_[18394]_ ;
  assign \new_[18406]_  = ~A167 & A168;
  assign \new_[18407]_  = A169 & \new_[18406]_ ;
  assign \new_[18411]_  = ~A200 & ~A199;
  assign \new_[18412]_  = A166 & \new_[18411]_ ;
  assign \new_[18413]_  = \new_[18412]_  & \new_[18407]_ ;
  assign \new_[18417]_  = A233 & ~A232;
  assign \new_[18418]_  = ~A202 & \new_[18417]_ ;
  assign \new_[18421]_  = A236 & ~A235;
  assign \new_[18424]_  = A300 & A299;
  assign \new_[18425]_  = \new_[18424]_  & \new_[18421]_ ;
  assign \new_[18426]_  = \new_[18425]_  & \new_[18418]_ ;
  assign \new_[18430]_  = ~A167 & A168;
  assign \new_[18431]_  = A169 & \new_[18430]_ ;
  assign \new_[18435]_  = ~A200 & ~A199;
  assign \new_[18436]_  = A166 & \new_[18435]_ ;
  assign \new_[18437]_  = \new_[18436]_  & \new_[18431]_ ;
  assign \new_[18441]_  = A233 & ~A232;
  assign \new_[18442]_  = ~A202 & \new_[18441]_ ;
  assign \new_[18445]_  = A236 & ~A235;
  assign \new_[18448]_  = A300 & A298;
  assign \new_[18449]_  = \new_[18448]_  & \new_[18445]_ ;
  assign \new_[18450]_  = \new_[18449]_  & \new_[18442]_ ;
  assign \new_[18454]_  = ~A167 & A168;
  assign \new_[18455]_  = A169 & \new_[18454]_ ;
  assign \new_[18459]_  = ~A200 & ~A199;
  assign \new_[18460]_  = A166 & \new_[18459]_ ;
  assign \new_[18461]_  = \new_[18460]_  & \new_[18455]_ ;
  assign \new_[18465]_  = A233 & ~A232;
  assign \new_[18466]_  = ~A202 & \new_[18465]_ ;
  assign \new_[18469]_  = A236 & ~A235;
  assign \new_[18472]_  = A267 & A265;
  assign \new_[18473]_  = \new_[18472]_  & \new_[18469]_ ;
  assign \new_[18474]_  = \new_[18473]_  & \new_[18466]_ ;
  assign \new_[18478]_  = ~A167 & A168;
  assign \new_[18479]_  = A169 & \new_[18478]_ ;
  assign \new_[18483]_  = ~A200 & ~A199;
  assign \new_[18484]_  = A166 & \new_[18483]_ ;
  assign \new_[18485]_  = \new_[18484]_  & \new_[18479]_ ;
  assign \new_[18489]_  = A233 & ~A232;
  assign \new_[18490]_  = ~A202 & \new_[18489]_ ;
  assign \new_[18493]_  = A236 & ~A235;
  assign \new_[18496]_  = A267 & A266;
  assign \new_[18497]_  = \new_[18496]_  & \new_[18493]_ ;
  assign \new_[18498]_  = \new_[18497]_  & \new_[18490]_ ;
  assign \new_[18502]_  = ~A167 & A168;
  assign \new_[18503]_  = A169 & \new_[18502]_ ;
  assign \new_[18507]_  = ~A200 & ~A199;
  assign \new_[18508]_  = A166 & \new_[18507]_ ;
  assign \new_[18509]_  = \new_[18508]_  & \new_[18503]_ ;
  assign \new_[18513]_  = ~A233 & A232;
  assign \new_[18514]_  = ~A202 & \new_[18513]_ ;
  assign \new_[18517]_  = A236 & ~A235;
  assign \new_[18520]_  = A300 & A299;
  assign \new_[18521]_  = \new_[18520]_  & \new_[18517]_ ;
  assign \new_[18522]_  = \new_[18521]_  & \new_[18514]_ ;
  assign \new_[18526]_  = ~A167 & A168;
  assign \new_[18527]_  = A169 & \new_[18526]_ ;
  assign \new_[18531]_  = ~A200 & ~A199;
  assign \new_[18532]_  = A166 & \new_[18531]_ ;
  assign \new_[18533]_  = \new_[18532]_  & \new_[18527]_ ;
  assign \new_[18537]_  = ~A233 & A232;
  assign \new_[18538]_  = ~A202 & \new_[18537]_ ;
  assign \new_[18541]_  = A236 & ~A235;
  assign \new_[18544]_  = A300 & A298;
  assign \new_[18545]_  = \new_[18544]_  & \new_[18541]_ ;
  assign \new_[18546]_  = \new_[18545]_  & \new_[18538]_ ;
  assign \new_[18550]_  = ~A167 & A168;
  assign \new_[18551]_  = A169 & \new_[18550]_ ;
  assign \new_[18555]_  = ~A200 & ~A199;
  assign \new_[18556]_  = A166 & \new_[18555]_ ;
  assign \new_[18557]_  = \new_[18556]_  & \new_[18551]_ ;
  assign \new_[18561]_  = ~A233 & A232;
  assign \new_[18562]_  = ~A202 & \new_[18561]_ ;
  assign \new_[18565]_  = A236 & ~A235;
  assign \new_[18568]_  = A267 & A265;
  assign \new_[18569]_  = \new_[18568]_  & \new_[18565]_ ;
  assign \new_[18570]_  = \new_[18569]_  & \new_[18562]_ ;
  assign \new_[18574]_  = ~A167 & A168;
  assign \new_[18575]_  = A169 & \new_[18574]_ ;
  assign \new_[18579]_  = ~A200 & ~A199;
  assign \new_[18580]_  = A166 & \new_[18579]_ ;
  assign \new_[18581]_  = \new_[18580]_  & \new_[18575]_ ;
  assign \new_[18585]_  = ~A233 & A232;
  assign \new_[18586]_  = ~A202 & \new_[18585]_ ;
  assign \new_[18589]_  = A236 & ~A235;
  assign \new_[18592]_  = A267 & A266;
  assign \new_[18593]_  = \new_[18592]_  & \new_[18589]_ ;
  assign \new_[18594]_  = \new_[18593]_  & \new_[18586]_ ;
  assign \new_[18598]_  = ~A167 & A168;
  assign \new_[18599]_  = A169 & \new_[18598]_ ;
  assign \new_[18603]_  = ~A200 & ~A199;
  assign \new_[18604]_  = A166 & \new_[18603]_ ;
  assign \new_[18605]_  = \new_[18604]_  & \new_[18599]_ ;
  assign \new_[18609]_  = ~A233 & ~A232;
  assign \new_[18610]_  = ~A202 & \new_[18609]_ ;
  assign \new_[18613]_  = ~A236 & A235;
  assign \new_[18616]_  = A300 & A299;
  assign \new_[18617]_  = \new_[18616]_  & \new_[18613]_ ;
  assign \new_[18618]_  = \new_[18617]_  & \new_[18610]_ ;
  assign \new_[18622]_  = ~A167 & A168;
  assign \new_[18623]_  = A169 & \new_[18622]_ ;
  assign \new_[18627]_  = ~A200 & ~A199;
  assign \new_[18628]_  = A166 & \new_[18627]_ ;
  assign \new_[18629]_  = \new_[18628]_  & \new_[18623]_ ;
  assign \new_[18633]_  = ~A233 & ~A232;
  assign \new_[18634]_  = ~A202 & \new_[18633]_ ;
  assign \new_[18637]_  = ~A236 & A235;
  assign \new_[18640]_  = A300 & A298;
  assign \new_[18641]_  = \new_[18640]_  & \new_[18637]_ ;
  assign \new_[18642]_  = \new_[18641]_  & \new_[18634]_ ;
  assign \new_[18646]_  = ~A167 & A168;
  assign \new_[18647]_  = A169 & \new_[18646]_ ;
  assign \new_[18651]_  = ~A200 & ~A199;
  assign \new_[18652]_  = A166 & \new_[18651]_ ;
  assign \new_[18653]_  = \new_[18652]_  & \new_[18647]_ ;
  assign \new_[18657]_  = ~A233 & ~A232;
  assign \new_[18658]_  = ~A202 & \new_[18657]_ ;
  assign \new_[18661]_  = ~A236 & A235;
  assign \new_[18664]_  = A267 & A265;
  assign \new_[18665]_  = \new_[18664]_  & \new_[18661]_ ;
  assign \new_[18666]_  = \new_[18665]_  & \new_[18658]_ ;
  assign \new_[18670]_  = ~A167 & A168;
  assign \new_[18671]_  = A169 & \new_[18670]_ ;
  assign \new_[18675]_  = ~A200 & ~A199;
  assign \new_[18676]_  = A166 & \new_[18675]_ ;
  assign \new_[18677]_  = \new_[18676]_  & \new_[18671]_ ;
  assign \new_[18681]_  = ~A233 & ~A232;
  assign \new_[18682]_  = ~A202 & \new_[18681]_ ;
  assign \new_[18685]_  = ~A236 & A235;
  assign \new_[18688]_  = A267 & A266;
  assign \new_[18689]_  = \new_[18688]_  & \new_[18685]_ ;
  assign \new_[18690]_  = \new_[18689]_  & \new_[18682]_ ;
  assign \new_[18694]_  = ~A167 & A168;
  assign \new_[18695]_  = A169 & \new_[18694]_ ;
  assign \new_[18699]_  = ~A200 & ~A199;
  assign \new_[18700]_  = A166 & \new_[18699]_ ;
  assign \new_[18701]_  = \new_[18700]_  & \new_[18695]_ ;
  assign \new_[18705]_  = A234 & A232;
  assign \new_[18706]_  = A203 & \new_[18705]_ ;
  assign \new_[18709]_  = A299 & A298;
  assign \new_[18712]_  = ~A302 & A301;
  assign \new_[18713]_  = \new_[18712]_  & \new_[18709]_ ;
  assign \new_[18714]_  = \new_[18713]_  & \new_[18706]_ ;
  assign \new_[18718]_  = ~A167 & A168;
  assign \new_[18719]_  = A169 & \new_[18718]_ ;
  assign \new_[18723]_  = ~A200 & ~A199;
  assign \new_[18724]_  = A166 & \new_[18723]_ ;
  assign \new_[18725]_  = \new_[18724]_  & \new_[18719]_ ;
  assign \new_[18729]_  = A234 & A232;
  assign \new_[18730]_  = A203 & \new_[18729]_ ;
  assign \new_[18733]_  = ~A299 & A298;
  assign \new_[18736]_  = A302 & ~A301;
  assign \new_[18737]_  = \new_[18736]_  & \new_[18733]_ ;
  assign \new_[18738]_  = \new_[18737]_  & \new_[18730]_ ;
  assign \new_[18742]_  = ~A167 & A168;
  assign \new_[18743]_  = A169 & \new_[18742]_ ;
  assign \new_[18747]_  = ~A200 & ~A199;
  assign \new_[18748]_  = A166 & \new_[18747]_ ;
  assign \new_[18749]_  = \new_[18748]_  & \new_[18743]_ ;
  assign \new_[18753]_  = A234 & A232;
  assign \new_[18754]_  = A203 & \new_[18753]_ ;
  assign \new_[18757]_  = A299 & ~A298;
  assign \new_[18760]_  = A302 & ~A301;
  assign \new_[18761]_  = \new_[18760]_  & \new_[18757]_ ;
  assign \new_[18762]_  = \new_[18761]_  & \new_[18754]_ ;
  assign \new_[18766]_  = ~A167 & A168;
  assign \new_[18767]_  = A169 & \new_[18766]_ ;
  assign \new_[18771]_  = ~A200 & ~A199;
  assign \new_[18772]_  = A166 & \new_[18771]_ ;
  assign \new_[18773]_  = \new_[18772]_  & \new_[18767]_ ;
  assign \new_[18777]_  = A234 & A232;
  assign \new_[18778]_  = A203 & \new_[18777]_ ;
  assign \new_[18781]_  = ~A299 & ~A298;
  assign \new_[18784]_  = ~A302 & A301;
  assign \new_[18785]_  = \new_[18784]_  & \new_[18781]_ ;
  assign \new_[18786]_  = \new_[18785]_  & \new_[18778]_ ;
  assign \new_[18790]_  = ~A167 & A168;
  assign \new_[18791]_  = A169 & \new_[18790]_ ;
  assign \new_[18795]_  = ~A200 & ~A199;
  assign \new_[18796]_  = A166 & \new_[18795]_ ;
  assign \new_[18797]_  = \new_[18796]_  & \new_[18791]_ ;
  assign \new_[18801]_  = A234 & A232;
  assign \new_[18802]_  = A203 & \new_[18801]_ ;
  assign \new_[18805]_  = A266 & A265;
  assign \new_[18808]_  = ~A269 & A268;
  assign \new_[18809]_  = \new_[18808]_  & \new_[18805]_ ;
  assign \new_[18810]_  = \new_[18809]_  & \new_[18802]_ ;
  assign \new_[18814]_  = ~A167 & A168;
  assign \new_[18815]_  = A169 & \new_[18814]_ ;
  assign \new_[18819]_  = ~A200 & ~A199;
  assign \new_[18820]_  = A166 & \new_[18819]_ ;
  assign \new_[18821]_  = \new_[18820]_  & \new_[18815]_ ;
  assign \new_[18825]_  = A234 & A232;
  assign \new_[18826]_  = A203 & \new_[18825]_ ;
  assign \new_[18829]_  = A266 & ~A265;
  assign \new_[18832]_  = A269 & ~A268;
  assign \new_[18833]_  = \new_[18832]_  & \new_[18829]_ ;
  assign \new_[18834]_  = \new_[18833]_  & \new_[18826]_ ;
  assign \new_[18838]_  = ~A167 & A168;
  assign \new_[18839]_  = A169 & \new_[18838]_ ;
  assign \new_[18843]_  = ~A200 & ~A199;
  assign \new_[18844]_  = A166 & \new_[18843]_ ;
  assign \new_[18845]_  = \new_[18844]_  & \new_[18839]_ ;
  assign \new_[18849]_  = A234 & A232;
  assign \new_[18850]_  = A203 & \new_[18849]_ ;
  assign \new_[18853]_  = ~A266 & A265;
  assign \new_[18856]_  = A269 & ~A268;
  assign \new_[18857]_  = \new_[18856]_  & \new_[18853]_ ;
  assign \new_[18858]_  = \new_[18857]_  & \new_[18850]_ ;
  assign \new_[18862]_  = ~A167 & A168;
  assign \new_[18863]_  = A169 & \new_[18862]_ ;
  assign \new_[18867]_  = ~A200 & ~A199;
  assign \new_[18868]_  = A166 & \new_[18867]_ ;
  assign \new_[18869]_  = \new_[18868]_  & \new_[18863]_ ;
  assign \new_[18873]_  = A234 & A232;
  assign \new_[18874]_  = A203 & \new_[18873]_ ;
  assign \new_[18877]_  = ~A266 & ~A265;
  assign \new_[18880]_  = ~A269 & A268;
  assign \new_[18881]_  = \new_[18880]_  & \new_[18877]_ ;
  assign \new_[18882]_  = \new_[18881]_  & \new_[18874]_ ;
  assign \new_[18886]_  = ~A167 & A168;
  assign \new_[18887]_  = A169 & \new_[18886]_ ;
  assign \new_[18891]_  = ~A200 & ~A199;
  assign \new_[18892]_  = A166 & \new_[18891]_ ;
  assign \new_[18893]_  = \new_[18892]_  & \new_[18887]_ ;
  assign \new_[18897]_  = A234 & A233;
  assign \new_[18898]_  = A203 & \new_[18897]_ ;
  assign \new_[18901]_  = A299 & A298;
  assign \new_[18904]_  = ~A302 & A301;
  assign \new_[18905]_  = \new_[18904]_  & \new_[18901]_ ;
  assign \new_[18906]_  = \new_[18905]_  & \new_[18898]_ ;
  assign \new_[18910]_  = ~A167 & A168;
  assign \new_[18911]_  = A169 & \new_[18910]_ ;
  assign \new_[18915]_  = ~A200 & ~A199;
  assign \new_[18916]_  = A166 & \new_[18915]_ ;
  assign \new_[18917]_  = \new_[18916]_  & \new_[18911]_ ;
  assign \new_[18921]_  = A234 & A233;
  assign \new_[18922]_  = A203 & \new_[18921]_ ;
  assign \new_[18925]_  = ~A299 & A298;
  assign \new_[18928]_  = A302 & ~A301;
  assign \new_[18929]_  = \new_[18928]_  & \new_[18925]_ ;
  assign \new_[18930]_  = \new_[18929]_  & \new_[18922]_ ;
  assign \new_[18934]_  = ~A167 & A168;
  assign \new_[18935]_  = A169 & \new_[18934]_ ;
  assign \new_[18939]_  = ~A200 & ~A199;
  assign \new_[18940]_  = A166 & \new_[18939]_ ;
  assign \new_[18941]_  = \new_[18940]_  & \new_[18935]_ ;
  assign \new_[18945]_  = A234 & A233;
  assign \new_[18946]_  = A203 & \new_[18945]_ ;
  assign \new_[18949]_  = A299 & ~A298;
  assign \new_[18952]_  = A302 & ~A301;
  assign \new_[18953]_  = \new_[18952]_  & \new_[18949]_ ;
  assign \new_[18954]_  = \new_[18953]_  & \new_[18946]_ ;
  assign \new_[18958]_  = ~A167 & A168;
  assign \new_[18959]_  = A169 & \new_[18958]_ ;
  assign \new_[18963]_  = ~A200 & ~A199;
  assign \new_[18964]_  = A166 & \new_[18963]_ ;
  assign \new_[18965]_  = \new_[18964]_  & \new_[18959]_ ;
  assign \new_[18969]_  = A234 & A233;
  assign \new_[18970]_  = A203 & \new_[18969]_ ;
  assign \new_[18973]_  = ~A299 & ~A298;
  assign \new_[18976]_  = ~A302 & A301;
  assign \new_[18977]_  = \new_[18976]_  & \new_[18973]_ ;
  assign \new_[18978]_  = \new_[18977]_  & \new_[18970]_ ;
  assign \new_[18982]_  = ~A167 & A168;
  assign \new_[18983]_  = A169 & \new_[18982]_ ;
  assign \new_[18987]_  = ~A200 & ~A199;
  assign \new_[18988]_  = A166 & \new_[18987]_ ;
  assign \new_[18989]_  = \new_[18988]_  & \new_[18983]_ ;
  assign \new_[18993]_  = A234 & A233;
  assign \new_[18994]_  = A203 & \new_[18993]_ ;
  assign \new_[18997]_  = A266 & A265;
  assign \new_[19000]_  = ~A269 & A268;
  assign \new_[19001]_  = \new_[19000]_  & \new_[18997]_ ;
  assign \new_[19002]_  = \new_[19001]_  & \new_[18994]_ ;
  assign \new_[19006]_  = ~A167 & A168;
  assign \new_[19007]_  = A169 & \new_[19006]_ ;
  assign \new_[19011]_  = ~A200 & ~A199;
  assign \new_[19012]_  = A166 & \new_[19011]_ ;
  assign \new_[19013]_  = \new_[19012]_  & \new_[19007]_ ;
  assign \new_[19017]_  = A234 & A233;
  assign \new_[19018]_  = A203 & \new_[19017]_ ;
  assign \new_[19021]_  = A266 & ~A265;
  assign \new_[19024]_  = A269 & ~A268;
  assign \new_[19025]_  = \new_[19024]_  & \new_[19021]_ ;
  assign \new_[19026]_  = \new_[19025]_  & \new_[19018]_ ;
  assign \new_[19030]_  = ~A167 & A168;
  assign \new_[19031]_  = A169 & \new_[19030]_ ;
  assign \new_[19035]_  = ~A200 & ~A199;
  assign \new_[19036]_  = A166 & \new_[19035]_ ;
  assign \new_[19037]_  = \new_[19036]_  & \new_[19031]_ ;
  assign \new_[19041]_  = A234 & A233;
  assign \new_[19042]_  = A203 & \new_[19041]_ ;
  assign \new_[19045]_  = ~A266 & A265;
  assign \new_[19048]_  = A269 & ~A268;
  assign \new_[19049]_  = \new_[19048]_  & \new_[19045]_ ;
  assign \new_[19050]_  = \new_[19049]_  & \new_[19042]_ ;
  assign \new_[19054]_  = ~A167 & A168;
  assign \new_[19055]_  = A169 & \new_[19054]_ ;
  assign \new_[19059]_  = ~A200 & ~A199;
  assign \new_[19060]_  = A166 & \new_[19059]_ ;
  assign \new_[19061]_  = \new_[19060]_  & \new_[19055]_ ;
  assign \new_[19065]_  = A234 & A233;
  assign \new_[19066]_  = A203 & \new_[19065]_ ;
  assign \new_[19069]_  = ~A266 & ~A265;
  assign \new_[19072]_  = ~A269 & A268;
  assign \new_[19073]_  = \new_[19072]_  & \new_[19069]_ ;
  assign \new_[19074]_  = \new_[19073]_  & \new_[19066]_ ;
  assign \new_[19078]_  = ~A167 & A168;
  assign \new_[19079]_  = A169 & \new_[19078]_ ;
  assign \new_[19083]_  = ~A200 & ~A199;
  assign \new_[19084]_  = A166 & \new_[19083]_ ;
  assign \new_[19085]_  = \new_[19084]_  & \new_[19079]_ ;
  assign \new_[19089]_  = A233 & A232;
  assign \new_[19090]_  = A203 & \new_[19089]_ ;
  assign \new_[19093]_  = ~A236 & A235;
  assign \new_[19096]_  = A300 & A299;
  assign \new_[19097]_  = \new_[19096]_  & \new_[19093]_ ;
  assign \new_[19098]_  = \new_[19097]_  & \new_[19090]_ ;
  assign \new_[19102]_  = ~A167 & A168;
  assign \new_[19103]_  = A169 & \new_[19102]_ ;
  assign \new_[19107]_  = ~A200 & ~A199;
  assign \new_[19108]_  = A166 & \new_[19107]_ ;
  assign \new_[19109]_  = \new_[19108]_  & \new_[19103]_ ;
  assign \new_[19113]_  = A233 & A232;
  assign \new_[19114]_  = A203 & \new_[19113]_ ;
  assign \new_[19117]_  = ~A236 & A235;
  assign \new_[19120]_  = A300 & A298;
  assign \new_[19121]_  = \new_[19120]_  & \new_[19117]_ ;
  assign \new_[19122]_  = \new_[19121]_  & \new_[19114]_ ;
  assign \new_[19126]_  = ~A167 & A168;
  assign \new_[19127]_  = A169 & \new_[19126]_ ;
  assign \new_[19131]_  = ~A200 & ~A199;
  assign \new_[19132]_  = A166 & \new_[19131]_ ;
  assign \new_[19133]_  = \new_[19132]_  & \new_[19127]_ ;
  assign \new_[19137]_  = A233 & A232;
  assign \new_[19138]_  = A203 & \new_[19137]_ ;
  assign \new_[19141]_  = ~A236 & A235;
  assign \new_[19144]_  = A267 & A265;
  assign \new_[19145]_  = \new_[19144]_  & \new_[19141]_ ;
  assign \new_[19146]_  = \new_[19145]_  & \new_[19138]_ ;
  assign \new_[19150]_  = ~A167 & A168;
  assign \new_[19151]_  = A169 & \new_[19150]_ ;
  assign \new_[19155]_  = ~A200 & ~A199;
  assign \new_[19156]_  = A166 & \new_[19155]_ ;
  assign \new_[19157]_  = \new_[19156]_  & \new_[19151]_ ;
  assign \new_[19161]_  = A233 & A232;
  assign \new_[19162]_  = A203 & \new_[19161]_ ;
  assign \new_[19165]_  = ~A236 & A235;
  assign \new_[19168]_  = A267 & A266;
  assign \new_[19169]_  = \new_[19168]_  & \new_[19165]_ ;
  assign \new_[19170]_  = \new_[19169]_  & \new_[19162]_ ;
  assign \new_[19174]_  = ~A167 & A168;
  assign \new_[19175]_  = A169 & \new_[19174]_ ;
  assign \new_[19179]_  = ~A200 & ~A199;
  assign \new_[19180]_  = A166 & \new_[19179]_ ;
  assign \new_[19181]_  = \new_[19180]_  & \new_[19175]_ ;
  assign \new_[19185]_  = A233 & ~A232;
  assign \new_[19186]_  = A203 & \new_[19185]_ ;
  assign \new_[19189]_  = A236 & ~A235;
  assign \new_[19192]_  = A300 & A299;
  assign \new_[19193]_  = \new_[19192]_  & \new_[19189]_ ;
  assign \new_[19194]_  = \new_[19193]_  & \new_[19186]_ ;
  assign \new_[19198]_  = ~A167 & A168;
  assign \new_[19199]_  = A169 & \new_[19198]_ ;
  assign \new_[19203]_  = ~A200 & ~A199;
  assign \new_[19204]_  = A166 & \new_[19203]_ ;
  assign \new_[19205]_  = \new_[19204]_  & \new_[19199]_ ;
  assign \new_[19209]_  = A233 & ~A232;
  assign \new_[19210]_  = A203 & \new_[19209]_ ;
  assign \new_[19213]_  = A236 & ~A235;
  assign \new_[19216]_  = A300 & A298;
  assign \new_[19217]_  = \new_[19216]_  & \new_[19213]_ ;
  assign \new_[19218]_  = \new_[19217]_  & \new_[19210]_ ;
  assign \new_[19222]_  = ~A167 & A168;
  assign \new_[19223]_  = A169 & \new_[19222]_ ;
  assign \new_[19227]_  = ~A200 & ~A199;
  assign \new_[19228]_  = A166 & \new_[19227]_ ;
  assign \new_[19229]_  = \new_[19228]_  & \new_[19223]_ ;
  assign \new_[19233]_  = A233 & ~A232;
  assign \new_[19234]_  = A203 & \new_[19233]_ ;
  assign \new_[19237]_  = A236 & ~A235;
  assign \new_[19240]_  = A267 & A265;
  assign \new_[19241]_  = \new_[19240]_  & \new_[19237]_ ;
  assign \new_[19242]_  = \new_[19241]_  & \new_[19234]_ ;
  assign \new_[19246]_  = ~A167 & A168;
  assign \new_[19247]_  = A169 & \new_[19246]_ ;
  assign \new_[19251]_  = ~A200 & ~A199;
  assign \new_[19252]_  = A166 & \new_[19251]_ ;
  assign \new_[19253]_  = \new_[19252]_  & \new_[19247]_ ;
  assign \new_[19257]_  = A233 & ~A232;
  assign \new_[19258]_  = A203 & \new_[19257]_ ;
  assign \new_[19261]_  = A236 & ~A235;
  assign \new_[19264]_  = A267 & A266;
  assign \new_[19265]_  = \new_[19264]_  & \new_[19261]_ ;
  assign \new_[19266]_  = \new_[19265]_  & \new_[19258]_ ;
  assign \new_[19270]_  = ~A167 & A168;
  assign \new_[19271]_  = A169 & \new_[19270]_ ;
  assign \new_[19275]_  = ~A200 & ~A199;
  assign \new_[19276]_  = A166 & \new_[19275]_ ;
  assign \new_[19277]_  = \new_[19276]_  & \new_[19271]_ ;
  assign \new_[19281]_  = ~A233 & A232;
  assign \new_[19282]_  = A203 & \new_[19281]_ ;
  assign \new_[19285]_  = A236 & ~A235;
  assign \new_[19288]_  = A300 & A299;
  assign \new_[19289]_  = \new_[19288]_  & \new_[19285]_ ;
  assign \new_[19290]_  = \new_[19289]_  & \new_[19282]_ ;
  assign \new_[19294]_  = ~A167 & A168;
  assign \new_[19295]_  = A169 & \new_[19294]_ ;
  assign \new_[19299]_  = ~A200 & ~A199;
  assign \new_[19300]_  = A166 & \new_[19299]_ ;
  assign \new_[19301]_  = \new_[19300]_  & \new_[19295]_ ;
  assign \new_[19305]_  = ~A233 & A232;
  assign \new_[19306]_  = A203 & \new_[19305]_ ;
  assign \new_[19309]_  = A236 & ~A235;
  assign \new_[19312]_  = A300 & A298;
  assign \new_[19313]_  = \new_[19312]_  & \new_[19309]_ ;
  assign \new_[19314]_  = \new_[19313]_  & \new_[19306]_ ;
  assign \new_[19318]_  = ~A167 & A168;
  assign \new_[19319]_  = A169 & \new_[19318]_ ;
  assign \new_[19323]_  = ~A200 & ~A199;
  assign \new_[19324]_  = A166 & \new_[19323]_ ;
  assign \new_[19325]_  = \new_[19324]_  & \new_[19319]_ ;
  assign \new_[19329]_  = ~A233 & A232;
  assign \new_[19330]_  = A203 & \new_[19329]_ ;
  assign \new_[19333]_  = A236 & ~A235;
  assign \new_[19336]_  = A267 & A265;
  assign \new_[19337]_  = \new_[19336]_  & \new_[19333]_ ;
  assign \new_[19338]_  = \new_[19337]_  & \new_[19330]_ ;
  assign \new_[19342]_  = ~A167 & A168;
  assign \new_[19343]_  = A169 & \new_[19342]_ ;
  assign \new_[19347]_  = ~A200 & ~A199;
  assign \new_[19348]_  = A166 & \new_[19347]_ ;
  assign \new_[19349]_  = \new_[19348]_  & \new_[19343]_ ;
  assign \new_[19353]_  = ~A233 & A232;
  assign \new_[19354]_  = A203 & \new_[19353]_ ;
  assign \new_[19357]_  = A236 & ~A235;
  assign \new_[19360]_  = A267 & A266;
  assign \new_[19361]_  = \new_[19360]_  & \new_[19357]_ ;
  assign \new_[19362]_  = \new_[19361]_  & \new_[19354]_ ;
  assign \new_[19366]_  = ~A167 & A168;
  assign \new_[19367]_  = A169 & \new_[19366]_ ;
  assign \new_[19371]_  = ~A200 & ~A199;
  assign \new_[19372]_  = A166 & \new_[19371]_ ;
  assign \new_[19373]_  = \new_[19372]_  & \new_[19367]_ ;
  assign \new_[19377]_  = ~A233 & ~A232;
  assign \new_[19378]_  = A203 & \new_[19377]_ ;
  assign \new_[19381]_  = ~A236 & A235;
  assign \new_[19384]_  = A300 & A299;
  assign \new_[19385]_  = \new_[19384]_  & \new_[19381]_ ;
  assign \new_[19386]_  = \new_[19385]_  & \new_[19378]_ ;
  assign \new_[19390]_  = ~A167 & A168;
  assign \new_[19391]_  = A169 & \new_[19390]_ ;
  assign \new_[19395]_  = ~A200 & ~A199;
  assign \new_[19396]_  = A166 & \new_[19395]_ ;
  assign \new_[19397]_  = \new_[19396]_  & \new_[19391]_ ;
  assign \new_[19401]_  = ~A233 & ~A232;
  assign \new_[19402]_  = A203 & \new_[19401]_ ;
  assign \new_[19405]_  = ~A236 & A235;
  assign \new_[19408]_  = A300 & A298;
  assign \new_[19409]_  = \new_[19408]_  & \new_[19405]_ ;
  assign \new_[19410]_  = \new_[19409]_  & \new_[19402]_ ;
  assign \new_[19414]_  = ~A167 & A168;
  assign \new_[19415]_  = A169 & \new_[19414]_ ;
  assign \new_[19419]_  = ~A200 & ~A199;
  assign \new_[19420]_  = A166 & \new_[19419]_ ;
  assign \new_[19421]_  = \new_[19420]_  & \new_[19415]_ ;
  assign \new_[19425]_  = ~A233 & ~A232;
  assign \new_[19426]_  = A203 & \new_[19425]_ ;
  assign \new_[19429]_  = ~A236 & A235;
  assign \new_[19432]_  = A267 & A265;
  assign \new_[19433]_  = \new_[19432]_  & \new_[19429]_ ;
  assign \new_[19434]_  = \new_[19433]_  & \new_[19426]_ ;
  assign \new_[19438]_  = ~A167 & A168;
  assign \new_[19439]_  = A169 & \new_[19438]_ ;
  assign \new_[19443]_  = ~A200 & ~A199;
  assign \new_[19444]_  = A166 & \new_[19443]_ ;
  assign \new_[19445]_  = \new_[19444]_  & \new_[19439]_ ;
  assign \new_[19449]_  = ~A233 & ~A232;
  assign \new_[19450]_  = A203 & \new_[19449]_ ;
  assign \new_[19453]_  = ~A236 & A235;
  assign \new_[19456]_  = A267 & A266;
  assign \new_[19457]_  = \new_[19456]_  & \new_[19453]_ ;
  assign \new_[19458]_  = \new_[19457]_  & \new_[19450]_ ;
  assign \new_[19462]_  = A199 & ~A166;
  assign \new_[19463]_  = A167 & \new_[19462]_ ;
  assign \new_[19466]_  = ~A201 & A200;
  assign \new_[19469]_  = A232 & ~A202;
  assign \new_[19470]_  = \new_[19469]_  & \new_[19466]_ ;
  assign \new_[19471]_  = \new_[19470]_  & \new_[19463]_ ;
  assign \new_[19475]_  = ~A236 & A235;
  assign \new_[19476]_  = A233 & \new_[19475]_ ;
  assign \new_[19479]_  = A299 & A298;
  assign \new_[19482]_  = ~A302 & A301;
  assign \new_[19483]_  = \new_[19482]_  & \new_[19479]_ ;
  assign \new_[19484]_  = \new_[19483]_  & \new_[19476]_ ;
  assign \new_[19488]_  = A199 & ~A166;
  assign \new_[19489]_  = A167 & \new_[19488]_ ;
  assign \new_[19492]_  = ~A201 & A200;
  assign \new_[19495]_  = A232 & ~A202;
  assign \new_[19496]_  = \new_[19495]_  & \new_[19492]_ ;
  assign \new_[19497]_  = \new_[19496]_  & \new_[19489]_ ;
  assign \new_[19501]_  = ~A236 & A235;
  assign \new_[19502]_  = A233 & \new_[19501]_ ;
  assign \new_[19505]_  = ~A299 & A298;
  assign \new_[19508]_  = A302 & ~A301;
  assign \new_[19509]_  = \new_[19508]_  & \new_[19505]_ ;
  assign \new_[19510]_  = \new_[19509]_  & \new_[19502]_ ;
  assign \new_[19514]_  = A199 & ~A166;
  assign \new_[19515]_  = A167 & \new_[19514]_ ;
  assign \new_[19518]_  = ~A201 & A200;
  assign \new_[19521]_  = A232 & ~A202;
  assign \new_[19522]_  = \new_[19521]_  & \new_[19518]_ ;
  assign \new_[19523]_  = \new_[19522]_  & \new_[19515]_ ;
  assign \new_[19527]_  = ~A236 & A235;
  assign \new_[19528]_  = A233 & \new_[19527]_ ;
  assign \new_[19531]_  = A299 & ~A298;
  assign \new_[19534]_  = A302 & ~A301;
  assign \new_[19535]_  = \new_[19534]_  & \new_[19531]_ ;
  assign \new_[19536]_  = \new_[19535]_  & \new_[19528]_ ;
  assign \new_[19540]_  = A199 & ~A166;
  assign \new_[19541]_  = A167 & \new_[19540]_ ;
  assign \new_[19544]_  = ~A201 & A200;
  assign \new_[19547]_  = A232 & ~A202;
  assign \new_[19548]_  = \new_[19547]_  & \new_[19544]_ ;
  assign \new_[19549]_  = \new_[19548]_  & \new_[19541]_ ;
  assign \new_[19553]_  = ~A236 & A235;
  assign \new_[19554]_  = A233 & \new_[19553]_ ;
  assign \new_[19557]_  = ~A299 & ~A298;
  assign \new_[19560]_  = ~A302 & A301;
  assign \new_[19561]_  = \new_[19560]_  & \new_[19557]_ ;
  assign \new_[19562]_  = \new_[19561]_  & \new_[19554]_ ;
  assign \new_[19566]_  = A199 & ~A166;
  assign \new_[19567]_  = A167 & \new_[19566]_ ;
  assign \new_[19570]_  = ~A201 & A200;
  assign \new_[19573]_  = A232 & ~A202;
  assign \new_[19574]_  = \new_[19573]_  & \new_[19570]_ ;
  assign \new_[19575]_  = \new_[19574]_  & \new_[19567]_ ;
  assign \new_[19579]_  = ~A236 & A235;
  assign \new_[19580]_  = A233 & \new_[19579]_ ;
  assign \new_[19583]_  = A266 & A265;
  assign \new_[19586]_  = ~A269 & A268;
  assign \new_[19587]_  = \new_[19586]_  & \new_[19583]_ ;
  assign \new_[19588]_  = \new_[19587]_  & \new_[19580]_ ;
  assign \new_[19592]_  = A199 & ~A166;
  assign \new_[19593]_  = A167 & \new_[19592]_ ;
  assign \new_[19596]_  = ~A201 & A200;
  assign \new_[19599]_  = A232 & ~A202;
  assign \new_[19600]_  = \new_[19599]_  & \new_[19596]_ ;
  assign \new_[19601]_  = \new_[19600]_  & \new_[19593]_ ;
  assign \new_[19605]_  = ~A236 & A235;
  assign \new_[19606]_  = A233 & \new_[19605]_ ;
  assign \new_[19609]_  = A266 & ~A265;
  assign \new_[19612]_  = A269 & ~A268;
  assign \new_[19613]_  = \new_[19612]_  & \new_[19609]_ ;
  assign \new_[19614]_  = \new_[19613]_  & \new_[19606]_ ;
  assign \new_[19618]_  = A199 & ~A166;
  assign \new_[19619]_  = A167 & \new_[19618]_ ;
  assign \new_[19622]_  = ~A201 & A200;
  assign \new_[19625]_  = A232 & ~A202;
  assign \new_[19626]_  = \new_[19625]_  & \new_[19622]_ ;
  assign \new_[19627]_  = \new_[19626]_  & \new_[19619]_ ;
  assign \new_[19631]_  = ~A236 & A235;
  assign \new_[19632]_  = A233 & \new_[19631]_ ;
  assign \new_[19635]_  = ~A266 & A265;
  assign \new_[19638]_  = A269 & ~A268;
  assign \new_[19639]_  = \new_[19638]_  & \new_[19635]_ ;
  assign \new_[19640]_  = \new_[19639]_  & \new_[19632]_ ;
  assign \new_[19644]_  = A199 & ~A166;
  assign \new_[19645]_  = A167 & \new_[19644]_ ;
  assign \new_[19648]_  = ~A201 & A200;
  assign \new_[19651]_  = A232 & ~A202;
  assign \new_[19652]_  = \new_[19651]_  & \new_[19648]_ ;
  assign \new_[19653]_  = \new_[19652]_  & \new_[19645]_ ;
  assign \new_[19657]_  = ~A236 & A235;
  assign \new_[19658]_  = A233 & \new_[19657]_ ;
  assign \new_[19661]_  = ~A266 & ~A265;
  assign \new_[19664]_  = ~A269 & A268;
  assign \new_[19665]_  = \new_[19664]_  & \new_[19661]_ ;
  assign \new_[19666]_  = \new_[19665]_  & \new_[19658]_ ;
  assign \new_[19670]_  = A199 & ~A166;
  assign \new_[19671]_  = A167 & \new_[19670]_ ;
  assign \new_[19674]_  = ~A201 & A200;
  assign \new_[19677]_  = ~A232 & ~A202;
  assign \new_[19678]_  = \new_[19677]_  & \new_[19674]_ ;
  assign \new_[19679]_  = \new_[19678]_  & \new_[19671]_ ;
  assign \new_[19683]_  = A236 & ~A235;
  assign \new_[19684]_  = A233 & \new_[19683]_ ;
  assign \new_[19687]_  = A299 & A298;
  assign \new_[19690]_  = ~A302 & A301;
  assign \new_[19691]_  = \new_[19690]_  & \new_[19687]_ ;
  assign \new_[19692]_  = \new_[19691]_  & \new_[19684]_ ;
  assign \new_[19696]_  = A199 & ~A166;
  assign \new_[19697]_  = A167 & \new_[19696]_ ;
  assign \new_[19700]_  = ~A201 & A200;
  assign \new_[19703]_  = ~A232 & ~A202;
  assign \new_[19704]_  = \new_[19703]_  & \new_[19700]_ ;
  assign \new_[19705]_  = \new_[19704]_  & \new_[19697]_ ;
  assign \new_[19709]_  = A236 & ~A235;
  assign \new_[19710]_  = A233 & \new_[19709]_ ;
  assign \new_[19713]_  = ~A299 & A298;
  assign \new_[19716]_  = A302 & ~A301;
  assign \new_[19717]_  = \new_[19716]_  & \new_[19713]_ ;
  assign \new_[19718]_  = \new_[19717]_  & \new_[19710]_ ;
  assign \new_[19722]_  = A199 & ~A166;
  assign \new_[19723]_  = A167 & \new_[19722]_ ;
  assign \new_[19726]_  = ~A201 & A200;
  assign \new_[19729]_  = ~A232 & ~A202;
  assign \new_[19730]_  = \new_[19729]_  & \new_[19726]_ ;
  assign \new_[19731]_  = \new_[19730]_  & \new_[19723]_ ;
  assign \new_[19735]_  = A236 & ~A235;
  assign \new_[19736]_  = A233 & \new_[19735]_ ;
  assign \new_[19739]_  = A299 & ~A298;
  assign \new_[19742]_  = A302 & ~A301;
  assign \new_[19743]_  = \new_[19742]_  & \new_[19739]_ ;
  assign \new_[19744]_  = \new_[19743]_  & \new_[19736]_ ;
  assign \new_[19748]_  = A199 & ~A166;
  assign \new_[19749]_  = A167 & \new_[19748]_ ;
  assign \new_[19752]_  = ~A201 & A200;
  assign \new_[19755]_  = ~A232 & ~A202;
  assign \new_[19756]_  = \new_[19755]_  & \new_[19752]_ ;
  assign \new_[19757]_  = \new_[19756]_  & \new_[19749]_ ;
  assign \new_[19761]_  = A236 & ~A235;
  assign \new_[19762]_  = A233 & \new_[19761]_ ;
  assign \new_[19765]_  = ~A299 & ~A298;
  assign \new_[19768]_  = ~A302 & A301;
  assign \new_[19769]_  = \new_[19768]_  & \new_[19765]_ ;
  assign \new_[19770]_  = \new_[19769]_  & \new_[19762]_ ;
  assign \new_[19774]_  = A199 & ~A166;
  assign \new_[19775]_  = A167 & \new_[19774]_ ;
  assign \new_[19778]_  = ~A201 & A200;
  assign \new_[19781]_  = ~A232 & ~A202;
  assign \new_[19782]_  = \new_[19781]_  & \new_[19778]_ ;
  assign \new_[19783]_  = \new_[19782]_  & \new_[19775]_ ;
  assign \new_[19787]_  = A236 & ~A235;
  assign \new_[19788]_  = A233 & \new_[19787]_ ;
  assign \new_[19791]_  = A266 & A265;
  assign \new_[19794]_  = ~A269 & A268;
  assign \new_[19795]_  = \new_[19794]_  & \new_[19791]_ ;
  assign \new_[19796]_  = \new_[19795]_  & \new_[19788]_ ;
  assign \new_[19800]_  = A199 & ~A166;
  assign \new_[19801]_  = A167 & \new_[19800]_ ;
  assign \new_[19804]_  = ~A201 & A200;
  assign \new_[19807]_  = ~A232 & ~A202;
  assign \new_[19808]_  = \new_[19807]_  & \new_[19804]_ ;
  assign \new_[19809]_  = \new_[19808]_  & \new_[19801]_ ;
  assign \new_[19813]_  = A236 & ~A235;
  assign \new_[19814]_  = A233 & \new_[19813]_ ;
  assign \new_[19817]_  = A266 & ~A265;
  assign \new_[19820]_  = A269 & ~A268;
  assign \new_[19821]_  = \new_[19820]_  & \new_[19817]_ ;
  assign \new_[19822]_  = \new_[19821]_  & \new_[19814]_ ;
  assign \new_[19826]_  = A199 & ~A166;
  assign \new_[19827]_  = A167 & \new_[19826]_ ;
  assign \new_[19830]_  = ~A201 & A200;
  assign \new_[19833]_  = ~A232 & ~A202;
  assign \new_[19834]_  = \new_[19833]_  & \new_[19830]_ ;
  assign \new_[19835]_  = \new_[19834]_  & \new_[19827]_ ;
  assign \new_[19839]_  = A236 & ~A235;
  assign \new_[19840]_  = A233 & \new_[19839]_ ;
  assign \new_[19843]_  = ~A266 & A265;
  assign \new_[19846]_  = A269 & ~A268;
  assign \new_[19847]_  = \new_[19846]_  & \new_[19843]_ ;
  assign \new_[19848]_  = \new_[19847]_  & \new_[19840]_ ;
  assign \new_[19852]_  = A199 & ~A166;
  assign \new_[19853]_  = A167 & \new_[19852]_ ;
  assign \new_[19856]_  = ~A201 & A200;
  assign \new_[19859]_  = ~A232 & ~A202;
  assign \new_[19860]_  = \new_[19859]_  & \new_[19856]_ ;
  assign \new_[19861]_  = \new_[19860]_  & \new_[19853]_ ;
  assign \new_[19865]_  = A236 & ~A235;
  assign \new_[19866]_  = A233 & \new_[19865]_ ;
  assign \new_[19869]_  = ~A266 & ~A265;
  assign \new_[19872]_  = ~A269 & A268;
  assign \new_[19873]_  = \new_[19872]_  & \new_[19869]_ ;
  assign \new_[19874]_  = \new_[19873]_  & \new_[19866]_ ;
  assign \new_[19878]_  = A199 & ~A166;
  assign \new_[19879]_  = A167 & \new_[19878]_ ;
  assign \new_[19882]_  = ~A201 & A200;
  assign \new_[19885]_  = A232 & ~A202;
  assign \new_[19886]_  = \new_[19885]_  & \new_[19882]_ ;
  assign \new_[19887]_  = \new_[19886]_  & \new_[19879]_ ;
  assign \new_[19891]_  = A236 & ~A235;
  assign \new_[19892]_  = ~A233 & \new_[19891]_ ;
  assign \new_[19895]_  = A299 & A298;
  assign \new_[19898]_  = ~A302 & A301;
  assign \new_[19899]_  = \new_[19898]_  & \new_[19895]_ ;
  assign \new_[19900]_  = \new_[19899]_  & \new_[19892]_ ;
  assign \new_[19904]_  = A199 & ~A166;
  assign \new_[19905]_  = A167 & \new_[19904]_ ;
  assign \new_[19908]_  = ~A201 & A200;
  assign \new_[19911]_  = A232 & ~A202;
  assign \new_[19912]_  = \new_[19911]_  & \new_[19908]_ ;
  assign \new_[19913]_  = \new_[19912]_  & \new_[19905]_ ;
  assign \new_[19917]_  = A236 & ~A235;
  assign \new_[19918]_  = ~A233 & \new_[19917]_ ;
  assign \new_[19921]_  = ~A299 & A298;
  assign \new_[19924]_  = A302 & ~A301;
  assign \new_[19925]_  = \new_[19924]_  & \new_[19921]_ ;
  assign \new_[19926]_  = \new_[19925]_  & \new_[19918]_ ;
  assign \new_[19930]_  = A199 & ~A166;
  assign \new_[19931]_  = A167 & \new_[19930]_ ;
  assign \new_[19934]_  = ~A201 & A200;
  assign \new_[19937]_  = A232 & ~A202;
  assign \new_[19938]_  = \new_[19937]_  & \new_[19934]_ ;
  assign \new_[19939]_  = \new_[19938]_  & \new_[19931]_ ;
  assign \new_[19943]_  = A236 & ~A235;
  assign \new_[19944]_  = ~A233 & \new_[19943]_ ;
  assign \new_[19947]_  = A299 & ~A298;
  assign \new_[19950]_  = A302 & ~A301;
  assign \new_[19951]_  = \new_[19950]_  & \new_[19947]_ ;
  assign \new_[19952]_  = \new_[19951]_  & \new_[19944]_ ;
  assign \new_[19956]_  = A199 & ~A166;
  assign \new_[19957]_  = A167 & \new_[19956]_ ;
  assign \new_[19960]_  = ~A201 & A200;
  assign \new_[19963]_  = A232 & ~A202;
  assign \new_[19964]_  = \new_[19963]_  & \new_[19960]_ ;
  assign \new_[19965]_  = \new_[19964]_  & \new_[19957]_ ;
  assign \new_[19969]_  = A236 & ~A235;
  assign \new_[19970]_  = ~A233 & \new_[19969]_ ;
  assign \new_[19973]_  = ~A299 & ~A298;
  assign \new_[19976]_  = ~A302 & A301;
  assign \new_[19977]_  = \new_[19976]_  & \new_[19973]_ ;
  assign \new_[19978]_  = \new_[19977]_  & \new_[19970]_ ;
  assign \new_[19982]_  = A199 & ~A166;
  assign \new_[19983]_  = A167 & \new_[19982]_ ;
  assign \new_[19986]_  = ~A201 & A200;
  assign \new_[19989]_  = A232 & ~A202;
  assign \new_[19990]_  = \new_[19989]_  & \new_[19986]_ ;
  assign \new_[19991]_  = \new_[19990]_  & \new_[19983]_ ;
  assign \new_[19995]_  = A236 & ~A235;
  assign \new_[19996]_  = ~A233 & \new_[19995]_ ;
  assign \new_[19999]_  = A266 & A265;
  assign \new_[20002]_  = ~A269 & A268;
  assign \new_[20003]_  = \new_[20002]_  & \new_[19999]_ ;
  assign \new_[20004]_  = \new_[20003]_  & \new_[19996]_ ;
  assign \new_[20008]_  = A199 & ~A166;
  assign \new_[20009]_  = A167 & \new_[20008]_ ;
  assign \new_[20012]_  = ~A201 & A200;
  assign \new_[20015]_  = A232 & ~A202;
  assign \new_[20016]_  = \new_[20015]_  & \new_[20012]_ ;
  assign \new_[20017]_  = \new_[20016]_  & \new_[20009]_ ;
  assign \new_[20021]_  = A236 & ~A235;
  assign \new_[20022]_  = ~A233 & \new_[20021]_ ;
  assign \new_[20025]_  = A266 & ~A265;
  assign \new_[20028]_  = A269 & ~A268;
  assign \new_[20029]_  = \new_[20028]_  & \new_[20025]_ ;
  assign \new_[20030]_  = \new_[20029]_  & \new_[20022]_ ;
  assign \new_[20034]_  = A199 & ~A166;
  assign \new_[20035]_  = A167 & \new_[20034]_ ;
  assign \new_[20038]_  = ~A201 & A200;
  assign \new_[20041]_  = A232 & ~A202;
  assign \new_[20042]_  = \new_[20041]_  & \new_[20038]_ ;
  assign \new_[20043]_  = \new_[20042]_  & \new_[20035]_ ;
  assign \new_[20047]_  = A236 & ~A235;
  assign \new_[20048]_  = ~A233 & \new_[20047]_ ;
  assign \new_[20051]_  = ~A266 & A265;
  assign \new_[20054]_  = A269 & ~A268;
  assign \new_[20055]_  = \new_[20054]_  & \new_[20051]_ ;
  assign \new_[20056]_  = \new_[20055]_  & \new_[20048]_ ;
  assign \new_[20060]_  = A199 & ~A166;
  assign \new_[20061]_  = A167 & \new_[20060]_ ;
  assign \new_[20064]_  = ~A201 & A200;
  assign \new_[20067]_  = A232 & ~A202;
  assign \new_[20068]_  = \new_[20067]_  & \new_[20064]_ ;
  assign \new_[20069]_  = \new_[20068]_  & \new_[20061]_ ;
  assign \new_[20073]_  = A236 & ~A235;
  assign \new_[20074]_  = ~A233 & \new_[20073]_ ;
  assign \new_[20077]_  = ~A266 & ~A265;
  assign \new_[20080]_  = ~A269 & A268;
  assign \new_[20081]_  = \new_[20080]_  & \new_[20077]_ ;
  assign \new_[20082]_  = \new_[20081]_  & \new_[20074]_ ;
  assign \new_[20086]_  = A199 & ~A166;
  assign \new_[20087]_  = A167 & \new_[20086]_ ;
  assign \new_[20090]_  = ~A201 & A200;
  assign \new_[20093]_  = ~A232 & ~A202;
  assign \new_[20094]_  = \new_[20093]_  & \new_[20090]_ ;
  assign \new_[20095]_  = \new_[20094]_  & \new_[20087]_ ;
  assign \new_[20099]_  = ~A236 & A235;
  assign \new_[20100]_  = ~A233 & \new_[20099]_ ;
  assign \new_[20103]_  = A299 & A298;
  assign \new_[20106]_  = ~A302 & A301;
  assign \new_[20107]_  = \new_[20106]_  & \new_[20103]_ ;
  assign \new_[20108]_  = \new_[20107]_  & \new_[20100]_ ;
  assign \new_[20112]_  = A199 & ~A166;
  assign \new_[20113]_  = A167 & \new_[20112]_ ;
  assign \new_[20116]_  = ~A201 & A200;
  assign \new_[20119]_  = ~A232 & ~A202;
  assign \new_[20120]_  = \new_[20119]_  & \new_[20116]_ ;
  assign \new_[20121]_  = \new_[20120]_  & \new_[20113]_ ;
  assign \new_[20125]_  = ~A236 & A235;
  assign \new_[20126]_  = ~A233 & \new_[20125]_ ;
  assign \new_[20129]_  = ~A299 & A298;
  assign \new_[20132]_  = A302 & ~A301;
  assign \new_[20133]_  = \new_[20132]_  & \new_[20129]_ ;
  assign \new_[20134]_  = \new_[20133]_  & \new_[20126]_ ;
  assign \new_[20138]_  = A199 & ~A166;
  assign \new_[20139]_  = A167 & \new_[20138]_ ;
  assign \new_[20142]_  = ~A201 & A200;
  assign \new_[20145]_  = ~A232 & ~A202;
  assign \new_[20146]_  = \new_[20145]_  & \new_[20142]_ ;
  assign \new_[20147]_  = \new_[20146]_  & \new_[20139]_ ;
  assign \new_[20151]_  = ~A236 & A235;
  assign \new_[20152]_  = ~A233 & \new_[20151]_ ;
  assign \new_[20155]_  = A299 & ~A298;
  assign \new_[20158]_  = A302 & ~A301;
  assign \new_[20159]_  = \new_[20158]_  & \new_[20155]_ ;
  assign \new_[20160]_  = \new_[20159]_  & \new_[20152]_ ;
  assign \new_[20164]_  = A199 & ~A166;
  assign \new_[20165]_  = A167 & \new_[20164]_ ;
  assign \new_[20168]_  = ~A201 & A200;
  assign \new_[20171]_  = ~A232 & ~A202;
  assign \new_[20172]_  = \new_[20171]_  & \new_[20168]_ ;
  assign \new_[20173]_  = \new_[20172]_  & \new_[20165]_ ;
  assign \new_[20177]_  = ~A236 & A235;
  assign \new_[20178]_  = ~A233 & \new_[20177]_ ;
  assign \new_[20181]_  = ~A299 & ~A298;
  assign \new_[20184]_  = ~A302 & A301;
  assign \new_[20185]_  = \new_[20184]_  & \new_[20181]_ ;
  assign \new_[20186]_  = \new_[20185]_  & \new_[20178]_ ;
  assign \new_[20190]_  = A199 & ~A166;
  assign \new_[20191]_  = A167 & \new_[20190]_ ;
  assign \new_[20194]_  = ~A201 & A200;
  assign \new_[20197]_  = ~A232 & ~A202;
  assign \new_[20198]_  = \new_[20197]_  & \new_[20194]_ ;
  assign \new_[20199]_  = \new_[20198]_  & \new_[20191]_ ;
  assign \new_[20203]_  = ~A236 & A235;
  assign \new_[20204]_  = ~A233 & \new_[20203]_ ;
  assign \new_[20207]_  = A266 & A265;
  assign \new_[20210]_  = ~A269 & A268;
  assign \new_[20211]_  = \new_[20210]_  & \new_[20207]_ ;
  assign \new_[20212]_  = \new_[20211]_  & \new_[20204]_ ;
  assign \new_[20216]_  = A199 & ~A166;
  assign \new_[20217]_  = A167 & \new_[20216]_ ;
  assign \new_[20220]_  = ~A201 & A200;
  assign \new_[20223]_  = ~A232 & ~A202;
  assign \new_[20224]_  = \new_[20223]_  & \new_[20220]_ ;
  assign \new_[20225]_  = \new_[20224]_  & \new_[20217]_ ;
  assign \new_[20229]_  = ~A236 & A235;
  assign \new_[20230]_  = ~A233 & \new_[20229]_ ;
  assign \new_[20233]_  = A266 & ~A265;
  assign \new_[20236]_  = A269 & ~A268;
  assign \new_[20237]_  = \new_[20236]_  & \new_[20233]_ ;
  assign \new_[20238]_  = \new_[20237]_  & \new_[20230]_ ;
  assign \new_[20242]_  = A199 & ~A166;
  assign \new_[20243]_  = A167 & \new_[20242]_ ;
  assign \new_[20246]_  = ~A201 & A200;
  assign \new_[20249]_  = ~A232 & ~A202;
  assign \new_[20250]_  = \new_[20249]_  & \new_[20246]_ ;
  assign \new_[20251]_  = \new_[20250]_  & \new_[20243]_ ;
  assign \new_[20255]_  = ~A236 & A235;
  assign \new_[20256]_  = ~A233 & \new_[20255]_ ;
  assign \new_[20259]_  = ~A266 & A265;
  assign \new_[20262]_  = A269 & ~A268;
  assign \new_[20263]_  = \new_[20262]_  & \new_[20259]_ ;
  assign \new_[20264]_  = \new_[20263]_  & \new_[20256]_ ;
  assign \new_[20268]_  = A199 & ~A166;
  assign \new_[20269]_  = A167 & \new_[20268]_ ;
  assign \new_[20272]_  = ~A201 & A200;
  assign \new_[20275]_  = ~A232 & ~A202;
  assign \new_[20276]_  = \new_[20275]_  & \new_[20272]_ ;
  assign \new_[20277]_  = \new_[20276]_  & \new_[20269]_ ;
  assign \new_[20281]_  = ~A236 & A235;
  assign \new_[20282]_  = ~A233 & \new_[20281]_ ;
  assign \new_[20285]_  = ~A266 & ~A265;
  assign \new_[20288]_  = ~A269 & A268;
  assign \new_[20289]_  = \new_[20288]_  & \new_[20285]_ ;
  assign \new_[20290]_  = \new_[20289]_  & \new_[20282]_ ;
  assign \new_[20294]_  = A199 & ~A166;
  assign \new_[20295]_  = A167 & \new_[20294]_ ;
  assign \new_[20298]_  = ~A201 & A200;
  assign \new_[20301]_  = A232 & A203;
  assign \new_[20302]_  = \new_[20301]_  & \new_[20298]_ ;
  assign \new_[20303]_  = \new_[20302]_  & \new_[20295]_ ;
  assign \new_[20307]_  = ~A236 & A235;
  assign \new_[20308]_  = A233 & \new_[20307]_ ;
  assign \new_[20311]_  = A299 & A298;
  assign \new_[20314]_  = ~A302 & A301;
  assign \new_[20315]_  = \new_[20314]_  & \new_[20311]_ ;
  assign \new_[20316]_  = \new_[20315]_  & \new_[20308]_ ;
  assign \new_[20320]_  = A199 & ~A166;
  assign \new_[20321]_  = A167 & \new_[20320]_ ;
  assign \new_[20324]_  = ~A201 & A200;
  assign \new_[20327]_  = A232 & A203;
  assign \new_[20328]_  = \new_[20327]_  & \new_[20324]_ ;
  assign \new_[20329]_  = \new_[20328]_  & \new_[20321]_ ;
  assign \new_[20333]_  = ~A236 & A235;
  assign \new_[20334]_  = A233 & \new_[20333]_ ;
  assign \new_[20337]_  = ~A299 & A298;
  assign \new_[20340]_  = A302 & ~A301;
  assign \new_[20341]_  = \new_[20340]_  & \new_[20337]_ ;
  assign \new_[20342]_  = \new_[20341]_  & \new_[20334]_ ;
  assign \new_[20346]_  = A199 & ~A166;
  assign \new_[20347]_  = A167 & \new_[20346]_ ;
  assign \new_[20350]_  = ~A201 & A200;
  assign \new_[20353]_  = A232 & A203;
  assign \new_[20354]_  = \new_[20353]_  & \new_[20350]_ ;
  assign \new_[20355]_  = \new_[20354]_  & \new_[20347]_ ;
  assign \new_[20359]_  = ~A236 & A235;
  assign \new_[20360]_  = A233 & \new_[20359]_ ;
  assign \new_[20363]_  = A299 & ~A298;
  assign \new_[20366]_  = A302 & ~A301;
  assign \new_[20367]_  = \new_[20366]_  & \new_[20363]_ ;
  assign \new_[20368]_  = \new_[20367]_  & \new_[20360]_ ;
  assign \new_[20372]_  = A199 & ~A166;
  assign \new_[20373]_  = A167 & \new_[20372]_ ;
  assign \new_[20376]_  = ~A201 & A200;
  assign \new_[20379]_  = A232 & A203;
  assign \new_[20380]_  = \new_[20379]_  & \new_[20376]_ ;
  assign \new_[20381]_  = \new_[20380]_  & \new_[20373]_ ;
  assign \new_[20385]_  = ~A236 & A235;
  assign \new_[20386]_  = A233 & \new_[20385]_ ;
  assign \new_[20389]_  = ~A299 & ~A298;
  assign \new_[20392]_  = ~A302 & A301;
  assign \new_[20393]_  = \new_[20392]_  & \new_[20389]_ ;
  assign \new_[20394]_  = \new_[20393]_  & \new_[20386]_ ;
  assign \new_[20398]_  = A199 & ~A166;
  assign \new_[20399]_  = A167 & \new_[20398]_ ;
  assign \new_[20402]_  = ~A201 & A200;
  assign \new_[20405]_  = A232 & A203;
  assign \new_[20406]_  = \new_[20405]_  & \new_[20402]_ ;
  assign \new_[20407]_  = \new_[20406]_  & \new_[20399]_ ;
  assign \new_[20411]_  = ~A236 & A235;
  assign \new_[20412]_  = A233 & \new_[20411]_ ;
  assign \new_[20415]_  = A266 & A265;
  assign \new_[20418]_  = ~A269 & A268;
  assign \new_[20419]_  = \new_[20418]_  & \new_[20415]_ ;
  assign \new_[20420]_  = \new_[20419]_  & \new_[20412]_ ;
  assign \new_[20424]_  = A199 & ~A166;
  assign \new_[20425]_  = A167 & \new_[20424]_ ;
  assign \new_[20428]_  = ~A201 & A200;
  assign \new_[20431]_  = A232 & A203;
  assign \new_[20432]_  = \new_[20431]_  & \new_[20428]_ ;
  assign \new_[20433]_  = \new_[20432]_  & \new_[20425]_ ;
  assign \new_[20437]_  = ~A236 & A235;
  assign \new_[20438]_  = A233 & \new_[20437]_ ;
  assign \new_[20441]_  = A266 & ~A265;
  assign \new_[20444]_  = A269 & ~A268;
  assign \new_[20445]_  = \new_[20444]_  & \new_[20441]_ ;
  assign \new_[20446]_  = \new_[20445]_  & \new_[20438]_ ;
  assign \new_[20450]_  = A199 & ~A166;
  assign \new_[20451]_  = A167 & \new_[20450]_ ;
  assign \new_[20454]_  = ~A201 & A200;
  assign \new_[20457]_  = A232 & A203;
  assign \new_[20458]_  = \new_[20457]_  & \new_[20454]_ ;
  assign \new_[20459]_  = \new_[20458]_  & \new_[20451]_ ;
  assign \new_[20463]_  = ~A236 & A235;
  assign \new_[20464]_  = A233 & \new_[20463]_ ;
  assign \new_[20467]_  = ~A266 & A265;
  assign \new_[20470]_  = A269 & ~A268;
  assign \new_[20471]_  = \new_[20470]_  & \new_[20467]_ ;
  assign \new_[20472]_  = \new_[20471]_  & \new_[20464]_ ;
  assign \new_[20476]_  = A199 & ~A166;
  assign \new_[20477]_  = A167 & \new_[20476]_ ;
  assign \new_[20480]_  = ~A201 & A200;
  assign \new_[20483]_  = A232 & A203;
  assign \new_[20484]_  = \new_[20483]_  & \new_[20480]_ ;
  assign \new_[20485]_  = \new_[20484]_  & \new_[20477]_ ;
  assign \new_[20489]_  = ~A236 & A235;
  assign \new_[20490]_  = A233 & \new_[20489]_ ;
  assign \new_[20493]_  = ~A266 & ~A265;
  assign \new_[20496]_  = ~A269 & A268;
  assign \new_[20497]_  = \new_[20496]_  & \new_[20493]_ ;
  assign \new_[20498]_  = \new_[20497]_  & \new_[20490]_ ;
  assign \new_[20502]_  = A199 & ~A166;
  assign \new_[20503]_  = A167 & \new_[20502]_ ;
  assign \new_[20506]_  = ~A201 & A200;
  assign \new_[20509]_  = ~A232 & A203;
  assign \new_[20510]_  = \new_[20509]_  & \new_[20506]_ ;
  assign \new_[20511]_  = \new_[20510]_  & \new_[20503]_ ;
  assign \new_[20515]_  = A236 & ~A235;
  assign \new_[20516]_  = A233 & \new_[20515]_ ;
  assign \new_[20519]_  = A299 & A298;
  assign \new_[20522]_  = ~A302 & A301;
  assign \new_[20523]_  = \new_[20522]_  & \new_[20519]_ ;
  assign \new_[20524]_  = \new_[20523]_  & \new_[20516]_ ;
  assign \new_[20528]_  = A199 & ~A166;
  assign \new_[20529]_  = A167 & \new_[20528]_ ;
  assign \new_[20532]_  = ~A201 & A200;
  assign \new_[20535]_  = ~A232 & A203;
  assign \new_[20536]_  = \new_[20535]_  & \new_[20532]_ ;
  assign \new_[20537]_  = \new_[20536]_  & \new_[20529]_ ;
  assign \new_[20541]_  = A236 & ~A235;
  assign \new_[20542]_  = A233 & \new_[20541]_ ;
  assign \new_[20545]_  = ~A299 & A298;
  assign \new_[20548]_  = A302 & ~A301;
  assign \new_[20549]_  = \new_[20548]_  & \new_[20545]_ ;
  assign \new_[20550]_  = \new_[20549]_  & \new_[20542]_ ;
  assign \new_[20554]_  = A199 & ~A166;
  assign \new_[20555]_  = A167 & \new_[20554]_ ;
  assign \new_[20558]_  = ~A201 & A200;
  assign \new_[20561]_  = ~A232 & A203;
  assign \new_[20562]_  = \new_[20561]_  & \new_[20558]_ ;
  assign \new_[20563]_  = \new_[20562]_  & \new_[20555]_ ;
  assign \new_[20567]_  = A236 & ~A235;
  assign \new_[20568]_  = A233 & \new_[20567]_ ;
  assign \new_[20571]_  = A299 & ~A298;
  assign \new_[20574]_  = A302 & ~A301;
  assign \new_[20575]_  = \new_[20574]_  & \new_[20571]_ ;
  assign \new_[20576]_  = \new_[20575]_  & \new_[20568]_ ;
  assign \new_[20580]_  = A199 & ~A166;
  assign \new_[20581]_  = A167 & \new_[20580]_ ;
  assign \new_[20584]_  = ~A201 & A200;
  assign \new_[20587]_  = ~A232 & A203;
  assign \new_[20588]_  = \new_[20587]_  & \new_[20584]_ ;
  assign \new_[20589]_  = \new_[20588]_  & \new_[20581]_ ;
  assign \new_[20593]_  = A236 & ~A235;
  assign \new_[20594]_  = A233 & \new_[20593]_ ;
  assign \new_[20597]_  = ~A299 & ~A298;
  assign \new_[20600]_  = ~A302 & A301;
  assign \new_[20601]_  = \new_[20600]_  & \new_[20597]_ ;
  assign \new_[20602]_  = \new_[20601]_  & \new_[20594]_ ;
  assign \new_[20606]_  = A199 & ~A166;
  assign \new_[20607]_  = A167 & \new_[20606]_ ;
  assign \new_[20610]_  = ~A201 & A200;
  assign \new_[20613]_  = ~A232 & A203;
  assign \new_[20614]_  = \new_[20613]_  & \new_[20610]_ ;
  assign \new_[20615]_  = \new_[20614]_  & \new_[20607]_ ;
  assign \new_[20619]_  = A236 & ~A235;
  assign \new_[20620]_  = A233 & \new_[20619]_ ;
  assign \new_[20623]_  = A266 & A265;
  assign \new_[20626]_  = ~A269 & A268;
  assign \new_[20627]_  = \new_[20626]_  & \new_[20623]_ ;
  assign \new_[20628]_  = \new_[20627]_  & \new_[20620]_ ;
  assign \new_[20632]_  = A199 & ~A166;
  assign \new_[20633]_  = A167 & \new_[20632]_ ;
  assign \new_[20636]_  = ~A201 & A200;
  assign \new_[20639]_  = ~A232 & A203;
  assign \new_[20640]_  = \new_[20639]_  & \new_[20636]_ ;
  assign \new_[20641]_  = \new_[20640]_  & \new_[20633]_ ;
  assign \new_[20645]_  = A236 & ~A235;
  assign \new_[20646]_  = A233 & \new_[20645]_ ;
  assign \new_[20649]_  = A266 & ~A265;
  assign \new_[20652]_  = A269 & ~A268;
  assign \new_[20653]_  = \new_[20652]_  & \new_[20649]_ ;
  assign \new_[20654]_  = \new_[20653]_  & \new_[20646]_ ;
  assign \new_[20658]_  = A199 & ~A166;
  assign \new_[20659]_  = A167 & \new_[20658]_ ;
  assign \new_[20662]_  = ~A201 & A200;
  assign \new_[20665]_  = ~A232 & A203;
  assign \new_[20666]_  = \new_[20665]_  & \new_[20662]_ ;
  assign \new_[20667]_  = \new_[20666]_  & \new_[20659]_ ;
  assign \new_[20671]_  = A236 & ~A235;
  assign \new_[20672]_  = A233 & \new_[20671]_ ;
  assign \new_[20675]_  = ~A266 & A265;
  assign \new_[20678]_  = A269 & ~A268;
  assign \new_[20679]_  = \new_[20678]_  & \new_[20675]_ ;
  assign \new_[20680]_  = \new_[20679]_  & \new_[20672]_ ;
  assign \new_[20684]_  = A199 & ~A166;
  assign \new_[20685]_  = A167 & \new_[20684]_ ;
  assign \new_[20688]_  = ~A201 & A200;
  assign \new_[20691]_  = ~A232 & A203;
  assign \new_[20692]_  = \new_[20691]_  & \new_[20688]_ ;
  assign \new_[20693]_  = \new_[20692]_  & \new_[20685]_ ;
  assign \new_[20697]_  = A236 & ~A235;
  assign \new_[20698]_  = A233 & \new_[20697]_ ;
  assign \new_[20701]_  = ~A266 & ~A265;
  assign \new_[20704]_  = ~A269 & A268;
  assign \new_[20705]_  = \new_[20704]_  & \new_[20701]_ ;
  assign \new_[20706]_  = \new_[20705]_  & \new_[20698]_ ;
  assign \new_[20710]_  = A199 & ~A166;
  assign \new_[20711]_  = A167 & \new_[20710]_ ;
  assign \new_[20714]_  = ~A201 & A200;
  assign \new_[20717]_  = A232 & A203;
  assign \new_[20718]_  = \new_[20717]_  & \new_[20714]_ ;
  assign \new_[20719]_  = \new_[20718]_  & \new_[20711]_ ;
  assign \new_[20723]_  = A236 & ~A235;
  assign \new_[20724]_  = ~A233 & \new_[20723]_ ;
  assign \new_[20727]_  = A299 & A298;
  assign \new_[20730]_  = ~A302 & A301;
  assign \new_[20731]_  = \new_[20730]_  & \new_[20727]_ ;
  assign \new_[20732]_  = \new_[20731]_  & \new_[20724]_ ;
  assign \new_[20736]_  = A199 & ~A166;
  assign \new_[20737]_  = A167 & \new_[20736]_ ;
  assign \new_[20740]_  = ~A201 & A200;
  assign \new_[20743]_  = A232 & A203;
  assign \new_[20744]_  = \new_[20743]_  & \new_[20740]_ ;
  assign \new_[20745]_  = \new_[20744]_  & \new_[20737]_ ;
  assign \new_[20749]_  = A236 & ~A235;
  assign \new_[20750]_  = ~A233 & \new_[20749]_ ;
  assign \new_[20753]_  = ~A299 & A298;
  assign \new_[20756]_  = A302 & ~A301;
  assign \new_[20757]_  = \new_[20756]_  & \new_[20753]_ ;
  assign \new_[20758]_  = \new_[20757]_  & \new_[20750]_ ;
  assign \new_[20762]_  = A199 & ~A166;
  assign \new_[20763]_  = A167 & \new_[20762]_ ;
  assign \new_[20766]_  = ~A201 & A200;
  assign \new_[20769]_  = A232 & A203;
  assign \new_[20770]_  = \new_[20769]_  & \new_[20766]_ ;
  assign \new_[20771]_  = \new_[20770]_  & \new_[20763]_ ;
  assign \new_[20775]_  = A236 & ~A235;
  assign \new_[20776]_  = ~A233 & \new_[20775]_ ;
  assign \new_[20779]_  = A299 & ~A298;
  assign \new_[20782]_  = A302 & ~A301;
  assign \new_[20783]_  = \new_[20782]_  & \new_[20779]_ ;
  assign \new_[20784]_  = \new_[20783]_  & \new_[20776]_ ;
  assign \new_[20788]_  = A199 & ~A166;
  assign \new_[20789]_  = A167 & \new_[20788]_ ;
  assign \new_[20792]_  = ~A201 & A200;
  assign \new_[20795]_  = A232 & A203;
  assign \new_[20796]_  = \new_[20795]_  & \new_[20792]_ ;
  assign \new_[20797]_  = \new_[20796]_  & \new_[20789]_ ;
  assign \new_[20801]_  = A236 & ~A235;
  assign \new_[20802]_  = ~A233 & \new_[20801]_ ;
  assign \new_[20805]_  = ~A299 & ~A298;
  assign \new_[20808]_  = ~A302 & A301;
  assign \new_[20809]_  = \new_[20808]_  & \new_[20805]_ ;
  assign \new_[20810]_  = \new_[20809]_  & \new_[20802]_ ;
  assign \new_[20814]_  = A199 & ~A166;
  assign \new_[20815]_  = A167 & \new_[20814]_ ;
  assign \new_[20818]_  = ~A201 & A200;
  assign \new_[20821]_  = A232 & A203;
  assign \new_[20822]_  = \new_[20821]_  & \new_[20818]_ ;
  assign \new_[20823]_  = \new_[20822]_  & \new_[20815]_ ;
  assign \new_[20827]_  = A236 & ~A235;
  assign \new_[20828]_  = ~A233 & \new_[20827]_ ;
  assign \new_[20831]_  = A266 & A265;
  assign \new_[20834]_  = ~A269 & A268;
  assign \new_[20835]_  = \new_[20834]_  & \new_[20831]_ ;
  assign \new_[20836]_  = \new_[20835]_  & \new_[20828]_ ;
  assign \new_[20840]_  = A199 & ~A166;
  assign \new_[20841]_  = A167 & \new_[20840]_ ;
  assign \new_[20844]_  = ~A201 & A200;
  assign \new_[20847]_  = A232 & A203;
  assign \new_[20848]_  = \new_[20847]_  & \new_[20844]_ ;
  assign \new_[20849]_  = \new_[20848]_  & \new_[20841]_ ;
  assign \new_[20853]_  = A236 & ~A235;
  assign \new_[20854]_  = ~A233 & \new_[20853]_ ;
  assign \new_[20857]_  = A266 & ~A265;
  assign \new_[20860]_  = A269 & ~A268;
  assign \new_[20861]_  = \new_[20860]_  & \new_[20857]_ ;
  assign \new_[20862]_  = \new_[20861]_  & \new_[20854]_ ;
  assign \new_[20866]_  = A199 & ~A166;
  assign \new_[20867]_  = A167 & \new_[20866]_ ;
  assign \new_[20870]_  = ~A201 & A200;
  assign \new_[20873]_  = A232 & A203;
  assign \new_[20874]_  = \new_[20873]_  & \new_[20870]_ ;
  assign \new_[20875]_  = \new_[20874]_  & \new_[20867]_ ;
  assign \new_[20879]_  = A236 & ~A235;
  assign \new_[20880]_  = ~A233 & \new_[20879]_ ;
  assign \new_[20883]_  = ~A266 & A265;
  assign \new_[20886]_  = A269 & ~A268;
  assign \new_[20887]_  = \new_[20886]_  & \new_[20883]_ ;
  assign \new_[20888]_  = \new_[20887]_  & \new_[20880]_ ;
  assign \new_[20892]_  = A199 & ~A166;
  assign \new_[20893]_  = A167 & \new_[20892]_ ;
  assign \new_[20896]_  = ~A201 & A200;
  assign \new_[20899]_  = A232 & A203;
  assign \new_[20900]_  = \new_[20899]_  & \new_[20896]_ ;
  assign \new_[20901]_  = \new_[20900]_  & \new_[20893]_ ;
  assign \new_[20905]_  = A236 & ~A235;
  assign \new_[20906]_  = ~A233 & \new_[20905]_ ;
  assign \new_[20909]_  = ~A266 & ~A265;
  assign \new_[20912]_  = ~A269 & A268;
  assign \new_[20913]_  = \new_[20912]_  & \new_[20909]_ ;
  assign \new_[20914]_  = \new_[20913]_  & \new_[20906]_ ;
  assign \new_[20918]_  = A199 & ~A166;
  assign \new_[20919]_  = A167 & \new_[20918]_ ;
  assign \new_[20922]_  = ~A201 & A200;
  assign \new_[20925]_  = ~A232 & A203;
  assign \new_[20926]_  = \new_[20925]_  & \new_[20922]_ ;
  assign \new_[20927]_  = \new_[20926]_  & \new_[20919]_ ;
  assign \new_[20931]_  = ~A236 & A235;
  assign \new_[20932]_  = ~A233 & \new_[20931]_ ;
  assign \new_[20935]_  = A299 & A298;
  assign \new_[20938]_  = ~A302 & A301;
  assign \new_[20939]_  = \new_[20938]_  & \new_[20935]_ ;
  assign \new_[20940]_  = \new_[20939]_  & \new_[20932]_ ;
  assign \new_[20944]_  = A199 & ~A166;
  assign \new_[20945]_  = A167 & \new_[20944]_ ;
  assign \new_[20948]_  = ~A201 & A200;
  assign \new_[20951]_  = ~A232 & A203;
  assign \new_[20952]_  = \new_[20951]_  & \new_[20948]_ ;
  assign \new_[20953]_  = \new_[20952]_  & \new_[20945]_ ;
  assign \new_[20957]_  = ~A236 & A235;
  assign \new_[20958]_  = ~A233 & \new_[20957]_ ;
  assign \new_[20961]_  = ~A299 & A298;
  assign \new_[20964]_  = A302 & ~A301;
  assign \new_[20965]_  = \new_[20964]_  & \new_[20961]_ ;
  assign \new_[20966]_  = \new_[20965]_  & \new_[20958]_ ;
  assign \new_[20970]_  = A199 & ~A166;
  assign \new_[20971]_  = A167 & \new_[20970]_ ;
  assign \new_[20974]_  = ~A201 & A200;
  assign \new_[20977]_  = ~A232 & A203;
  assign \new_[20978]_  = \new_[20977]_  & \new_[20974]_ ;
  assign \new_[20979]_  = \new_[20978]_  & \new_[20971]_ ;
  assign \new_[20983]_  = ~A236 & A235;
  assign \new_[20984]_  = ~A233 & \new_[20983]_ ;
  assign \new_[20987]_  = A299 & ~A298;
  assign \new_[20990]_  = A302 & ~A301;
  assign \new_[20991]_  = \new_[20990]_  & \new_[20987]_ ;
  assign \new_[20992]_  = \new_[20991]_  & \new_[20984]_ ;
  assign \new_[20996]_  = A199 & ~A166;
  assign \new_[20997]_  = A167 & \new_[20996]_ ;
  assign \new_[21000]_  = ~A201 & A200;
  assign \new_[21003]_  = ~A232 & A203;
  assign \new_[21004]_  = \new_[21003]_  & \new_[21000]_ ;
  assign \new_[21005]_  = \new_[21004]_  & \new_[20997]_ ;
  assign \new_[21009]_  = ~A236 & A235;
  assign \new_[21010]_  = ~A233 & \new_[21009]_ ;
  assign \new_[21013]_  = ~A299 & ~A298;
  assign \new_[21016]_  = ~A302 & A301;
  assign \new_[21017]_  = \new_[21016]_  & \new_[21013]_ ;
  assign \new_[21018]_  = \new_[21017]_  & \new_[21010]_ ;
  assign \new_[21022]_  = A199 & ~A166;
  assign \new_[21023]_  = A167 & \new_[21022]_ ;
  assign \new_[21026]_  = ~A201 & A200;
  assign \new_[21029]_  = ~A232 & A203;
  assign \new_[21030]_  = \new_[21029]_  & \new_[21026]_ ;
  assign \new_[21031]_  = \new_[21030]_  & \new_[21023]_ ;
  assign \new_[21035]_  = ~A236 & A235;
  assign \new_[21036]_  = ~A233 & \new_[21035]_ ;
  assign \new_[21039]_  = A266 & A265;
  assign \new_[21042]_  = ~A269 & A268;
  assign \new_[21043]_  = \new_[21042]_  & \new_[21039]_ ;
  assign \new_[21044]_  = \new_[21043]_  & \new_[21036]_ ;
  assign \new_[21048]_  = A199 & ~A166;
  assign \new_[21049]_  = A167 & \new_[21048]_ ;
  assign \new_[21052]_  = ~A201 & A200;
  assign \new_[21055]_  = ~A232 & A203;
  assign \new_[21056]_  = \new_[21055]_  & \new_[21052]_ ;
  assign \new_[21057]_  = \new_[21056]_  & \new_[21049]_ ;
  assign \new_[21061]_  = ~A236 & A235;
  assign \new_[21062]_  = ~A233 & \new_[21061]_ ;
  assign \new_[21065]_  = A266 & ~A265;
  assign \new_[21068]_  = A269 & ~A268;
  assign \new_[21069]_  = \new_[21068]_  & \new_[21065]_ ;
  assign \new_[21070]_  = \new_[21069]_  & \new_[21062]_ ;
  assign \new_[21074]_  = A199 & ~A166;
  assign \new_[21075]_  = A167 & \new_[21074]_ ;
  assign \new_[21078]_  = ~A201 & A200;
  assign \new_[21081]_  = ~A232 & A203;
  assign \new_[21082]_  = \new_[21081]_  & \new_[21078]_ ;
  assign \new_[21083]_  = \new_[21082]_  & \new_[21075]_ ;
  assign \new_[21087]_  = ~A236 & A235;
  assign \new_[21088]_  = ~A233 & \new_[21087]_ ;
  assign \new_[21091]_  = ~A266 & A265;
  assign \new_[21094]_  = A269 & ~A268;
  assign \new_[21095]_  = \new_[21094]_  & \new_[21091]_ ;
  assign \new_[21096]_  = \new_[21095]_  & \new_[21088]_ ;
  assign \new_[21100]_  = A199 & ~A166;
  assign \new_[21101]_  = A167 & \new_[21100]_ ;
  assign \new_[21104]_  = ~A201 & A200;
  assign \new_[21107]_  = ~A232 & A203;
  assign \new_[21108]_  = \new_[21107]_  & \new_[21104]_ ;
  assign \new_[21109]_  = \new_[21108]_  & \new_[21101]_ ;
  assign \new_[21113]_  = ~A236 & A235;
  assign \new_[21114]_  = ~A233 & \new_[21113]_ ;
  assign \new_[21117]_  = ~A266 & ~A265;
  assign \new_[21120]_  = ~A269 & A268;
  assign \new_[21121]_  = \new_[21120]_  & \new_[21117]_ ;
  assign \new_[21122]_  = \new_[21121]_  & \new_[21114]_ ;
  assign \new_[21126]_  = ~A199 & ~A166;
  assign \new_[21127]_  = A167 & \new_[21126]_ ;
  assign \new_[21130]_  = ~A201 & A200;
  assign \new_[21133]_  = A232 & A202;
  assign \new_[21134]_  = \new_[21133]_  & \new_[21130]_ ;
  assign \new_[21135]_  = \new_[21134]_  & \new_[21127]_ ;
  assign \new_[21139]_  = ~A236 & A235;
  assign \new_[21140]_  = A233 & \new_[21139]_ ;
  assign \new_[21143]_  = A299 & A298;
  assign \new_[21146]_  = ~A302 & A301;
  assign \new_[21147]_  = \new_[21146]_  & \new_[21143]_ ;
  assign \new_[21148]_  = \new_[21147]_  & \new_[21140]_ ;
  assign \new_[21152]_  = ~A199 & ~A166;
  assign \new_[21153]_  = A167 & \new_[21152]_ ;
  assign \new_[21156]_  = ~A201 & A200;
  assign \new_[21159]_  = A232 & A202;
  assign \new_[21160]_  = \new_[21159]_  & \new_[21156]_ ;
  assign \new_[21161]_  = \new_[21160]_  & \new_[21153]_ ;
  assign \new_[21165]_  = ~A236 & A235;
  assign \new_[21166]_  = A233 & \new_[21165]_ ;
  assign \new_[21169]_  = ~A299 & A298;
  assign \new_[21172]_  = A302 & ~A301;
  assign \new_[21173]_  = \new_[21172]_  & \new_[21169]_ ;
  assign \new_[21174]_  = \new_[21173]_  & \new_[21166]_ ;
  assign \new_[21178]_  = ~A199 & ~A166;
  assign \new_[21179]_  = A167 & \new_[21178]_ ;
  assign \new_[21182]_  = ~A201 & A200;
  assign \new_[21185]_  = A232 & A202;
  assign \new_[21186]_  = \new_[21185]_  & \new_[21182]_ ;
  assign \new_[21187]_  = \new_[21186]_  & \new_[21179]_ ;
  assign \new_[21191]_  = ~A236 & A235;
  assign \new_[21192]_  = A233 & \new_[21191]_ ;
  assign \new_[21195]_  = A299 & ~A298;
  assign \new_[21198]_  = A302 & ~A301;
  assign \new_[21199]_  = \new_[21198]_  & \new_[21195]_ ;
  assign \new_[21200]_  = \new_[21199]_  & \new_[21192]_ ;
  assign \new_[21204]_  = ~A199 & ~A166;
  assign \new_[21205]_  = A167 & \new_[21204]_ ;
  assign \new_[21208]_  = ~A201 & A200;
  assign \new_[21211]_  = A232 & A202;
  assign \new_[21212]_  = \new_[21211]_  & \new_[21208]_ ;
  assign \new_[21213]_  = \new_[21212]_  & \new_[21205]_ ;
  assign \new_[21217]_  = ~A236 & A235;
  assign \new_[21218]_  = A233 & \new_[21217]_ ;
  assign \new_[21221]_  = ~A299 & ~A298;
  assign \new_[21224]_  = ~A302 & A301;
  assign \new_[21225]_  = \new_[21224]_  & \new_[21221]_ ;
  assign \new_[21226]_  = \new_[21225]_  & \new_[21218]_ ;
  assign \new_[21230]_  = ~A199 & ~A166;
  assign \new_[21231]_  = A167 & \new_[21230]_ ;
  assign \new_[21234]_  = ~A201 & A200;
  assign \new_[21237]_  = A232 & A202;
  assign \new_[21238]_  = \new_[21237]_  & \new_[21234]_ ;
  assign \new_[21239]_  = \new_[21238]_  & \new_[21231]_ ;
  assign \new_[21243]_  = ~A236 & A235;
  assign \new_[21244]_  = A233 & \new_[21243]_ ;
  assign \new_[21247]_  = A266 & A265;
  assign \new_[21250]_  = ~A269 & A268;
  assign \new_[21251]_  = \new_[21250]_  & \new_[21247]_ ;
  assign \new_[21252]_  = \new_[21251]_  & \new_[21244]_ ;
  assign \new_[21256]_  = ~A199 & ~A166;
  assign \new_[21257]_  = A167 & \new_[21256]_ ;
  assign \new_[21260]_  = ~A201 & A200;
  assign \new_[21263]_  = A232 & A202;
  assign \new_[21264]_  = \new_[21263]_  & \new_[21260]_ ;
  assign \new_[21265]_  = \new_[21264]_  & \new_[21257]_ ;
  assign \new_[21269]_  = ~A236 & A235;
  assign \new_[21270]_  = A233 & \new_[21269]_ ;
  assign \new_[21273]_  = A266 & ~A265;
  assign \new_[21276]_  = A269 & ~A268;
  assign \new_[21277]_  = \new_[21276]_  & \new_[21273]_ ;
  assign \new_[21278]_  = \new_[21277]_  & \new_[21270]_ ;
  assign \new_[21282]_  = ~A199 & ~A166;
  assign \new_[21283]_  = A167 & \new_[21282]_ ;
  assign \new_[21286]_  = ~A201 & A200;
  assign \new_[21289]_  = A232 & A202;
  assign \new_[21290]_  = \new_[21289]_  & \new_[21286]_ ;
  assign \new_[21291]_  = \new_[21290]_  & \new_[21283]_ ;
  assign \new_[21295]_  = ~A236 & A235;
  assign \new_[21296]_  = A233 & \new_[21295]_ ;
  assign \new_[21299]_  = ~A266 & A265;
  assign \new_[21302]_  = A269 & ~A268;
  assign \new_[21303]_  = \new_[21302]_  & \new_[21299]_ ;
  assign \new_[21304]_  = \new_[21303]_  & \new_[21296]_ ;
  assign \new_[21308]_  = ~A199 & ~A166;
  assign \new_[21309]_  = A167 & \new_[21308]_ ;
  assign \new_[21312]_  = ~A201 & A200;
  assign \new_[21315]_  = A232 & A202;
  assign \new_[21316]_  = \new_[21315]_  & \new_[21312]_ ;
  assign \new_[21317]_  = \new_[21316]_  & \new_[21309]_ ;
  assign \new_[21321]_  = ~A236 & A235;
  assign \new_[21322]_  = A233 & \new_[21321]_ ;
  assign \new_[21325]_  = ~A266 & ~A265;
  assign \new_[21328]_  = ~A269 & A268;
  assign \new_[21329]_  = \new_[21328]_  & \new_[21325]_ ;
  assign \new_[21330]_  = \new_[21329]_  & \new_[21322]_ ;
  assign \new_[21334]_  = ~A199 & ~A166;
  assign \new_[21335]_  = A167 & \new_[21334]_ ;
  assign \new_[21338]_  = ~A201 & A200;
  assign \new_[21341]_  = ~A232 & A202;
  assign \new_[21342]_  = \new_[21341]_  & \new_[21338]_ ;
  assign \new_[21343]_  = \new_[21342]_  & \new_[21335]_ ;
  assign \new_[21347]_  = A236 & ~A235;
  assign \new_[21348]_  = A233 & \new_[21347]_ ;
  assign \new_[21351]_  = A299 & A298;
  assign \new_[21354]_  = ~A302 & A301;
  assign \new_[21355]_  = \new_[21354]_  & \new_[21351]_ ;
  assign \new_[21356]_  = \new_[21355]_  & \new_[21348]_ ;
  assign \new_[21360]_  = ~A199 & ~A166;
  assign \new_[21361]_  = A167 & \new_[21360]_ ;
  assign \new_[21364]_  = ~A201 & A200;
  assign \new_[21367]_  = ~A232 & A202;
  assign \new_[21368]_  = \new_[21367]_  & \new_[21364]_ ;
  assign \new_[21369]_  = \new_[21368]_  & \new_[21361]_ ;
  assign \new_[21373]_  = A236 & ~A235;
  assign \new_[21374]_  = A233 & \new_[21373]_ ;
  assign \new_[21377]_  = ~A299 & A298;
  assign \new_[21380]_  = A302 & ~A301;
  assign \new_[21381]_  = \new_[21380]_  & \new_[21377]_ ;
  assign \new_[21382]_  = \new_[21381]_  & \new_[21374]_ ;
  assign \new_[21386]_  = ~A199 & ~A166;
  assign \new_[21387]_  = A167 & \new_[21386]_ ;
  assign \new_[21390]_  = ~A201 & A200;
  assign \new_[21393]_  = ~A232 & A202;
  assign \new_[21394]_  = \new_[21393]_  & \new_[21390]_ ;
  assign \new_[21395]_  = \new_[21394]_  & \new_[21387]_ ;
  assign \new_[21399]_  = A236 & ~A235;
  assign \new_[21400]_  = A233 & \new_[21399]_ ;
  assign \new_[21403]_  = A299 & ~A298;
  assign \new_[21406]_  = A302 & ~A301;
  assign \new_[21407]_  = \new_[21406]_  & \new_[21403]_ ;
  assign \new_[21408]_  = \new_[21407]_  & \new_[21400]_ ;
  assign \new_[21412]_  = ~A199 & ~A166;
  assign \new_[21413]_  = A167 & \new_[21412]_ ;
  assign \new_[21416]_  = ~A201 & A200;
  assign \new_[21419]_  = ~A232 & A202;
  assign \new_[21420]_  = \new_[21419]_  & \new_[21416]_ ;
  assign \new_[21421]_  = \new_[21420]_  & \new_[21413]_ ;
  assign \new_[21425]_  = A236 & ~A235;
  assign \new_[21426]_  = A233 & \new_[21425]_ ;
  assign \new_[21429]_  = ~A299 & ~A298;
  assign \new_[21432]_  = ~A302 & A301;
  assign \new_[21433]_  = \new_[21432]_  & \new_[21429]_ ;
  assign \new_[21434]_  = \new_[21433]_  & \new_[21426]_ ;
  assign \new_[21438]_  = ~A199 & ~A166;
  assign \new_[21439]_  = A167 & \new_[21438]_ ;
  assign \new_[21442]_  = ~A201 & A200;
  assign \new_[21445]_  = ~A232 & A202;
  assign \new_[21446]_  = \new_[21445]_  & \new_[21442]_ ;
  assign \new_[21447]_  = \new_[21446]_  & \new_[21439]_ ;
  assign \new_[21451]_  = A236 & ~A235;
  assign \new_[21452]_  = A233 & \new_[21451]_ ;
  assign \new_[21455]_  = A266 & A265;
  assign \new_[21458]_  = ~A269 & A268;
  assign \new_[21459]_  = \new_[21458]_  & \new_[21455]_ ;
  assign \new_[21460]_  = \new_[21459]_  & \new_[21452]_ ;
  assign \new_[21464]_  = ~A199 & ~A166;
  assign \new_[21465]_  = A167 & \new_[21464]_ ;
  assign \new_[21468]_  = ~A201 & A200;
  assign \new_[21471]_  = ~A232 & A202;
  assign \new_[21472]_  = \new_[21471]_  & \new_[21468]_ ;
  assign \new_[21473]_  = \new_[21472]_  & \new_[21465]_ ;
  assign \new_[21477]_  = A236 & ~A235;
  assign \new_[21478]_  = A233 & \new_[21477]_ ;
  assign \new_[21481]_  = A266 & ~A265;
  assign \new_[21484]_  = A269 & ~A268;
  assign \new_[21485]_  = \new_[21484]_  & \new_[21481]_ ;
  assign \new_[21486]_  = \new_[21485]_  & \new_[21478]_ ;
  assign \new_[21490]_  = ~A199 & ~A166;
  assign \new_[21491]_  = A167 & \new_[21490]_ ;
  assign \new_[21494]_  = ~A201 & A200;
  assign \new_[21497]_  = ~A232 & A202;
  assign \new_[21498]_  = \new_[21497]_  & \new_[21494]_ ;
  assign \new_[21499]_  = \new_[21498]_  & \new_[21491]_ ;
  assign \new_[21503]_  = A236 & ~A235;
  assign \new_[21504]_  = A233 & \new_[21503]_ ;
  assign \new_[21507]_  = ~A266 & A265;
  assign \new_[21510]_  = A269 & ~A268;
  assign \new_[21511]_  = \new_[21510]_  & \new_[21507]_ ;
  assign \new_[21512]_  = \new_[21511]_  & \new_[21504]_ ;
  assign \new_[21516]_  = ~A199 & ~A166;
  assign \new_[21517]_  = A167 & \new_[21516]_ ;
  assign \new_[21520]_  = ~A201 & A200;
  assign \new_[21523]_  = ~A232 & A202;
  assign \new_[21524]_  = \new_[21523]_  & \new_[21520]_ ;
  assign \new_[21525]_  = \new_[21524]_  & \new_[21517]_ ;
  assign \new_[21529]_  = A236 & ~A235;
  assign \new_[21530]_  = A233 & \new_[21529]_ ;
  assign \new_[21533]_  = ~A266 & ~A265;
  assign \new_[21536]_  = ~A269 & A268;
  assign \new_[21537]_  = \new_[21536]_  & \new_[21533]_ ;
  assign \new_[21538]_  = \new_[21537]_  & \new_[21530]_ ;
  assign \new_[21542]_  = ~A199 & ~A166;
  assign \new_[21543]_  = A167 & \new_[21542]_ ;
  assign \new_[21546]_  = ~A201 & A200;
  assign \new_[21549]_  = A232 & A202;
  assign \new_[21550]_  = \new_[21549]_  & \new_[21546]_ ;
  assign \new_[21551]_  = \new_[21550]_  & \new_[21543]_ ;
  assign \new_[21555]_  = A236 & ~A235;
  assign \new_[21556]_  = ~A233 & \new_[21555]_ ;
  assign \new_[21559]_  = A299 & A298;
  assign \new_[21562]_  = ~A302 & A301;
  assign \new_[21563]_  = \new_[21562]_  & \new_[21559]_ ;
  assign \new_[21564]_  = \new_[21563]_  & \new_[21556]_ ;
  assign \new_[21568]_  = ~A199 & ~A166;
  assign \new_[21569]_  = A167 & \new_[21568]_ ;
  assign \new_[21572]_  = ~A201 & A200;
  assign \new_[21575]_  = A232 & A202;
  assign \new_[21576]_  = \new_[21575]_  & \new_[21572]_ ;
  assign \new_[21577]_  = \new_[21576]_  & \new_[21569]_ ;
  assign \new_[21581]_  = A236 & ~A235;
  assign \new_[21582]_  = ~A233 & \new_[21581]_ ;
  assign \new_[21585]_  = ~A299 & A298;
  assign \new_[21588]_  = A302 & ~A301;
  assign \new_[21589]_  = \new_[21588]_  & \new_[21585]_ ;
  assign \new_[21590]_  = \new_[21589]_  & \new_[21582]_ ;
  assign \new_[21594]_  = ~A199 & ~A166;
  assign \new_[21595]_  = A167 & \new_[21594]_ ;
  assign \new_[21598]_  = ~A201 & A200;
  assign \new_[21601]_  = A232 & A202;
  assign \new_[21602]_  = \new_[21601]_  & \new_[21598]_ ;
  assign \new_[21603]_  = \new_[21602]_  & \new_[21595]_ ;
  assign \new_[21607]_  = A236 & ~A235;
  assign \new_[21608]_  = ~A233 & \new_[21607]_ ;
  assign \new_[21611]_  = A299 & ~A298;
  assign \new_[21614]_  = A302 & ~A301;
  assign \new_[21615]_  = \new_[21614]_  & \new_[21611]_ ;
  assign \new_[21616]_  = \new_[21615]_  & \new_[21608]_ ;
  assign \new_[21620]_  = ~A199 & ~A166;
  assign \new_[21621]_  = A167 & \new_[21620]_ ;
  assign \new_[21624]_  = ~A201 & A200;
  assign \new_[21627]_  = A232 & A202;
  assign \new_[21628]_  = \new_[21627]_  & \new_[21624]_ ;
  assign \new_[21629]_  = \new_[21628]_  & \new_[21621]_ ;
  assign \new_[21633]_  = A236 & ~A235;
  assign \new_[21634]_  = ~A233 & \new_[21633]_ ;
  assign \new_[21637]_  = ~A299 & ~A298;
  assign \new_[21640]_  = ~A302 & A301;
  assign \new_[21641]_  = \new_[21640]_  & \new_[21637]_ ;
  assign \new_[21642]_  = \new_[21641]_  & \new_[21634]_ ;
  assign \new_[21646]_  = ~A199 & ~A166;
  assign \new_[21647]_  = A167 & \new_[21646]_ ;
  assign \new_[21650]_  = ~A201 & A200;
  assign \new_[21653]_  = A232 & A202;
  assign \new_[21654]_  = \new_[21653]_  & \new_[21650]_ ;
  assign \new_[21655]_  = \new_[21654]_  & \new_[21647]_ ;
  assign \new_[21659]_  = A236 & ~A235;
  assign \new_[21660]_  = ~A233 & \new_[21659]_ ;
  assign \new_[21663]_  = A266 & A265;
  assign \new_[21666]_  = ~A269 & A268;
  assign \new_[21667]_  = \new_[21666]_  & \new_[21663]_ ;
  assign \new_[21668]_  = \new_[21667]_  & \new_[21660]_ ;
  assign \new_[21672]_  = ~A199 & ~A166;
  assign \new_[21673]_  = A167 & \new_[21672]_ ;
  assign \new_[21676]_  = ~A201 & A200;
  assign \new_[21679]_  = A232 & A202;
  assign \new_[21680]_  = \new_[21679]_  & \new_[21676]_ ;
  assign \new_[21681]_  = \new_[21680]_  & \new_[21673]_ ;
  assign \new_[21685]_  = A236 & ~A235;
  assign \new_[21686]_  = ~A233 & \new_[21685]_ ;
  assign \new_[21689]_  = A266 & ~A265;
  assign \new_[21692]_  = A269 & ~A268;
  assign \new_[21693]_  = \new_[21692]_  & \new_[21689]_ ;
  assign \new_[21694]_  = \new_[21693]_  & \new_[21686]_ ;
  assign \new_[21698]_  = ~A199 & ~A166;
  assign \new_[21699]_  = A167 & \new_[21698]_ ;
  assign \new_[21702]_  = ~A201 & A200;
  assign \new_[21705]_  = A232 & A202;
  assign \new_[21706]_  = \new_[21705]_  & \new_[21702]_ ;
  assign \new_[21707]_  = \new_[21706]_  & \new_[21699]_ ;
  assign \new_[21711]_  = A236 & ~A235;
  assign \new_[21712]_  = ~A233 & \new_[21711]_ ;
  assign \new_[21715]_  = ~A266 & A265;
  assign \new_[21718]_  = A269 & ~A268;
  assign \new_[21719]_  = \new_[21718]_  & \new_[21715]_ ;
  assign \new_[21720]_  = \new_[21719]_  & \new_[21712]_ ;
  assign \new_[21724]_  = ~A199 & ~A166;
  assign \new_[21725]_  = A167 & \new_[21724]_ ;
  assign \new_[21728]_  = ~A201 & A200;
  assign \new_[21731]_  = A232 & A202;
  assign \new_[21732]_  = \new_[21731]_  & \new_[21728]_ ;
  assign \new_[21733]_  = \new_[21732]_  & \new_[21725]_ ;
  assign \new_[21737]_  = A236 & ~A235;
  assign \new_[21738]_  = ~A233 & \new_[21737]_ ;
  assign \new_[21741]_  = ~A266 & ~A265;
  assign \new_[21744]_  = ~A269 & A268;
  assign \new_[21745]_  = \new_[21744]_  & \new_[21741]_ ;
  assign \new_[21746]_  = \new_[21745]_  & \new_[21738]_ ;
  assign \new_[21750]_  = ~A199 & ~A166;
  assign \new_[21751]_  = A167 & \new_[21750]_ ;
  assign \new_[21754]_  = ~A201 & A200;
  assign \new_[21757]_  = ~A232 & A202;
  assign \new_[21758]_  = \new_[21757]_  & \new_[21754]_ ;
  assign \new_[21759]_  = \new_[21758]_  & \new_[21751]_ ;
  assign \new_[21763]_  = ~A236 & A235;
  assign \new_[21764]_  = ~A233 & \new_[21763]_ ;
  assign \new_[21767]_  = A299 & A298;
  assign \new_[21770]_  = ~A302 & A301;
  assign \new_[21771]_  = \new_[21770]_  & \new_[21767]_ ;
  assign \new_[21772]_  = \new_[21771]_  & \new_[21764]_ ;
  assign \new_[21776]_  = ~A199 & ~A166;
  assign \new_[21777]_  = A167 & \new_[21776]_ ;
  assign \new_[21780]_  = ~A201 & A200;
  assign \new_[21783]_  = ~A232 & A202;
  assign \new_[21784]_  = \new_[21783]_  & \new_[21780]_ ;
  assign \new_[21785]_  = \new_[21784]_  & \new_[21777]_ ;
  assign \new_[21789]_  = ~A236 & A235;
  assign \new_[21790]_  = ~A233 & \new_[21789]_ ;
  assign \new_[21793]_  = ~A299 & A298;
  assign \new_[21796]_  = A302 & ~A301;
  assign \new_[21797]_  = \new_[21796]_  & \new_[21793]_ ;
  assign \new_[21798]_  = \new_[21797]_  & \new_[21790]_ ;
  assign \new_[21802]_  = ~A199 & ~A166;
  assign \new_[21803]_  = A167 & \new_[21802]_ ;
  assign \new_[21806]_  = ~A201 & A200;
  assign \new_[21809]_  = ~A232 & A202;
  assign \new_[21810]_  = \new_[21809]_  & \new_[21806]_ ;
  assign \new_[21811]_  = \new_[21810]_  & \new_[21803]_ ;
  assign \new_[21815]_  = ~A236 & A235;
  assign \new_[21816]_  = ~A233 & \new_[21815]_ ;
  assign \new_[21819]_  = A299 & ~A298;
  assign \new_[21822]_  = A302 & ~A301;
  assign \new_[21823]_  = \new_[21822]_  & \new_[21819]_ ;
  assign \new_[21824]_  = \new_[21823]_  & \new_[21816]_ ;
  assign \new_[21828]_  = ~A199 & ~A166;
  assign \new_[21829]_  = A167 & \new_[21828]_ ;
  assign \new_[21832]_  = ~A201 & A200;
  assign \new_[21835]_  = ~A232 & A202;
  assign \new_[21836]_  = \new_[21835]_  & \new_[21832]_ ;
  assign \new_[21837]_  = \new_[21836]_  & \new_[21829]_ ;
  assign \new_[21841]_  = ~A236 & A235;
  assign \new_[21842]_  = ~A233 & \new_[21841]_ ;
  assign \new_[21845]_  = ~A299 & ~A298;
  assign \new_[21848]_  = ~A302 & A301;
  assign \new_[21849]_  = \new_[21848]_  & \new_[21845]_ ;
  assign \new_[21850]_  = \new_[21849]_  & \new_[21842]_ ;
  assign \new_[21854]_  = ~A199 & ~A166;
  assign \new_[21855]_  = A167 & \new_[21854]_ ;
  assign \new_[21858]_  = ~A201 & A200;
  assign \new_[21861]_  = ~A232 & A202;
  assign \new_[21862]_  = \new_[21861]_  & \new_[21858]_ ;
  assign \new_[21863]_  = \new_[21862]_  & \new_[21855]_ ;
  assign \new_[21867]_  = ~A236 & A235;
  assign \new_[21868]_  = ~A233 & \new_[21867]_ ;
  assign \new_[21871]_  = A266 & A265;
  assign \new_[21874]_  = ~A269 & A268;
  assign \new_[21875]_  = \new_[21874]_  & \new_[21871]_ ;
  assign \new_[21876]_  = \new_[21875]_  & \new_[21868]_ ;
  assign \new_[21880]_  = ~A199 & ~A166;
  assign \new_[21881]_  = A167 & \new_[21880]_ ;
  assign \new_[21884]_  = ~A201 & A200;
  assign \new_[21887]_  = ~A232 & A202;
  assign \new_[21888]_  = \new_[21887]_  & \new_[21884]_ ;
  assign \new_[21889]_  = \new_[21888]_  & \new_[21881]_ ;
  assign \new_[21893]_  = ~A236 & A235;
  assign \new_[21894]_  = ~A233 & \new_[21893]_ ;
  assign \new_[21897]_  = A266 & ~A265;
  assign \new_[21900]_  = A269 & ~A268;
  assign \new_[21901]_  = \new_[21900]_  & \new_[21897]_ ;
  assign \new_[21902]_  = \new_[21901]_  & \new_[21894]_ ;
  assign \new_[21906]_  = ~A199 & ~A166;
  assign \new_[21907]_  = A167 & \new_[21906]_ ;
  assign \new_[21910]_  = ~A201 & A200;
  assign \new_[21913]_  = ~A232 & A202;
  assign \new_[21914]_  = \new_[21913]_  & \new_[21910]_ ;
  assign \new_[21915]_  = \new_[21914]_  & \new_[21907]_ ;
  assign \new_[21919]_  = ~A236 & A235;
  assign \new_[21920]_  = ~A233 & \new_[21919]_ ;
  assign \new_[21923]_  = ~A266 & A265;
  assign \new_[21926]_  = A269 & ~A268;
  assign \new_[21927]_  = \new_[21926]_  & \new_[21923]_ ;
  assign \new_[21928]_  = \new_[21927]_  & \new_[21920]_ ;
  assign \new_[21932]_  = ~A199 & ~A166;
  assign \new_[21933]_  = A167 & \new_[21932]_ ;
  assign \new_[21936]_  = ~A201 & A200;
  assign \new_[21939]_  = ~A232 & A202;
  assign \new_[21940]_  = \new_[21939]_  & \new_[21936]_ ;
  assign \new_[21941]_  = \new_[21940]_  & \new_[21933]_ ;
  assign \new_[21945]_  = ~A236 & A235;
  assign \new_[21946]_  = ~A233 & \new_[21945]_ ;
  assign \new_[21949]_  = ~A266 & ~A265;
  assign \new_[21952]_  = ~A269 & A268;
  assign \new_[21953]_  = \new_[21952]_  & \new_[21949]_ ;
  assign \new_[21954]_  = \new_[21953]_  & \new_[21946]_ ;
  assign \new_[21958]_  = ~A199 & ~A166;
  assign \new_[21959]_  = A167 & \new_[21958]_ ;
  assign \new_[21962]_  = ~A201 & A200;
  assign \new_[21965]_  = A232 & ~A203;
  assign \new_[21966]_  = \new_[21965]_  & \new_[21962]_ ;
  assign \new_[21967]_  = \new_[21966]_  & \new_[21959]_ ;
  assign \new_[21971]_  = ~A236 & A235;
  assign \new_[21972]_  = A233 & \new_[21971]_ ;
  assign \new_[21975]_  = A299 & A298;
  assign \new_[21978]_  = ~A302 & A301;
  assign \new_[21979]_  = \new_[21978]_  & \new_[21975]_ ;
  assign \new_[21980]_  = \new_[21979]_  & \new_[21972]_ ;
  assign \new_[21984]_  = ~A199 & ~A166;
  assign \new_[21985]_  = A167 & \new_[21984]_ ;
  assign \new_[21988]_  = ~A201 & A200;
  assign \new_[21991]_  = A232 & ~A203;
  assign \new_[21992]_  = \new_[21991]_  & \new_[21988]_ ;
  assign \new_[21993]_  = \new_[21992]_  & \new_[21985]_ ;
  assign \new_[21997]_  = ~A236 & A235;
  assign \new_[21998]_  = A233 & \new_[21997]_ ;
  assign \new_[22001]_  = ~A299 & A298;
  assign \new_[22004]_  = A302 & ~A301;
  assign \new_[22005]_  = \new_[22004]_  & \new_[22001]_ ;
  assign \new_[22006]_  = \new_[22005]_  & \new_[21998]_ ;
  assign \new_[22010]_  = ~A199 & ~A166;
  assign \new_[22011]_  = A167 & \new_[22010]_ ;
  assign \new_[22014]_  = ~A201 & A200;
  assign \new_[22017]_  = A232 & ~A203;
  assign \new_[22018]_  = \new_[22017]_  & \new_[22014]_ ;
  assign \new_[22019]_  = \new_[22018]_  & \new_[22011]_ ;
  assign \new_[22023]_  = ~A236 & A235;
  assign \new_[22024]_  = A233 & \new_[22023]_ ;
  assign \new_[22027]_  = A299 & ~A298;
  assign \new_[22030]_  = A302 & ~A301;
  assign \new_[22031]_  = \new_[22030]_  & \new_[22027]_ ;
  assign \new_[22032]_  = \new_[22031]_  & \new_[22024]_ ;
  assign \new_[22036]_  = ~A199 & ~A166;
  assign \new_[22037]_  = A167 & \new_[22036]_ ;
  assign \new_[22040]_  = ~A201 & A200;
  assign \new_[22043]_  = A232 & ~A203;
  assign \new_[22044]_  = \new_[22043]_  & \new_[22040]_ ;
  assign \new_[22045]_  = \new_[22044]_  & \new_[22037]_ ;
  assign \new_[22049]_  = ~A236 & A235;
  assign \new_[22050]_  = A233 & \new_[22049]_ ;
  assign \new_[22053]_  = ~A299 & ~A298;
  assign \new_[22056]_  = ~A302 & A301;
  assign \new_[22057]_  = \new_[22056]_  & \new_[22053]_ ;
  assign \new_[22058]_  = \new_[22057]_  & \new_[22050]_ ;
  assign \new_[22062]_  = ~A199 & ~A166;
  assign \new_[22063]_  = A167 & \new_[22062]_ ;
  assign \new_[22066]_  = ~A201 & A200;
  assign \new_[22069]_  = A232 & ~A203;
  assign \new_[22070]_  = \new_[22069]_  & \new_[22066]_ ;
  assign \new_[22071]_  = \new_[22070]_  & \new_[22063]_ ;
  assign \new_[22075]_  = ~A236 & A235;
  assign \new_[22076]_  = A233 & \new_[22075]_ ;
  assign \new_[22079]_  = A266 & A265;
  assign \new_[22082]_  = ~A269 & A268;
  assign \new_[22083]_  = \new_[22082]_  & \new_[22079]_ ;
  assign \new_[22084]_  = \new_[22083]_  & \new_[22076]_ ;
  assign \new_[22088]_  = ~A199 & ~A166;
  assign \new_[22089]_  = A167 & \new_[22088]_ ;
  assign \new_[22092]_  = ~A201 & A200;
  assign \new_[22095]_  = A232 & ~A203;
  assign \new_[22096]_  = \new_[22095]_  & \new_[22092]_ ;
  assign \new_[22097]_  = \new_[22096]_  & \new_[22089]_ ;
  assign \new_[22101]_  = ~A236 & A235;
  assign \new_[22102]_  = A233 & \new_[22101]_ ;
  assign \new_[22105]_  = A266 & ~A265;
  assign \new_[22108]_  = A269 & ~A268;
  assign \new_[22109]_  = \new_[22108]_  & \new_[22105]_ ;
  assign \new_[22110]_  = \new_[22109]_  & \new_[22102]_ ;
  assign \new_[22114]_  = ~A199 & ~A166;
  assign \new_[22115]_  = A167 & \new_[22114]_ ;
  assign \new_[22118]_  = ~A201 & A200;
  assign \new_[22121]_  = A232 & ~A203;
  assign \new_[22122]_  = \new_[22121]_  & \new_[22118]_ ;
  assign \new_[22123]_  = \new_[22122]_  & \new_[22115]_ ;
  assign \new_[22127]_  = ~A236 & A235;
  assign \new_[22128]_  = A233 & \new_[22127]_ ;
  assign \new_[22131]_  = ~A266 & A265;
  assign \new_[22134]_  = A269 & ~A268;
  assign \new_[22135]_  = \new_[22134]_  & \new_[22131]_ ;
  assign \new_[22136]_  = \new_[22135]_  & \new_[22128]_ ;
  assign \new_[22140]_  = ~A199 & ~A166;
  assign \new_[22141]_  = A167 & \new_[22140]_ ;
  assign \new_[22144]_  = ~A201 & A200;
  assign \new_[22147]_  = A232 & ~A203;
  assign \new_[22148]_  = \new_[22147]_  & \new_[22144]_ ;
  assign \new_[22149]_  = \new_[22148]_  & \new_[22141]_ ;
  assign \new_[22153]_  = ~A236 & A235;
  assign \new_[22154]_  = A233 & \new_[22153]_ ;
  assign \new_[22157]_  = ~A266 & ~A265;
  assign \new_[22160]_  = ~A269 & A268;
  assign \new_[22161]_  = \new_[22160]_  & \new_[22157]_ ;
  assign \new_[22162]_  = \new_[22161]_  & \new_[22154]_ ;
  assign \new_[22166]_  = ~A199 & ~A166;
  assign \new_[22167]_  = A167 & \new_[22166]_ ;
  assign \new_[22170]_  = ~A201 & A200;
  assign \new_[22173]_  = ~A232 & ~A203;
  assign \new_[22174]_  = \new_[22173]_  & \new_[22170]_ ;
  assign \new_[22175]_  = \new_[22174]_  & \new_[22167]_ ;
  assign \new_[22179]_  = A236 & ~A235;
  assign \new_[22180]_  = A233 & \new_[22179]_ ;
  assign \new_[22183]_  = A299 & A298;
  assign \new_[22186]_  = ~A302 & A301;
  assign \new_[22187]_  = \new_[22186]_  & \new_[22183]_ ;
  assign \new_[22188]_  = \new_[22187]_  & \new_[22180]_ ;
  assign \new_[22192]_  = ~A199 & ~A166;
  assign \new_[22193]_  = A167 & \new_[22192]_ ;
  assign \new_[22196]_  = ~A201 & A200;
  assign \new_[22199]_  = ~A232 & ~A203;
  assign \new_[22200]_  = \new_[22199]_  & \new_[22196]_ ;
  assign \new_[22201]_  = \new_[22200]_  & \new_[22193]_ ;
  assign \new_[22205]_  = A236 & ~A235;
  assign \new_[22206]_  = A233 & \new_[22205]_ ;
  assign \new_[22209]_  = ~A299 & A298;
  assign \new_[22212]_  = A302 & ~A301;
  assign \new_[22213]_  = \new_[22212]_  & \new_[22209]_ ;
  assign \new_[22214]_  = \new_[22213]_  & \new_[22206]_ ;
  assign \new_[22218]_  = ~A199 & ~A166;
  assign \new_[22219]_  = A167 & \new_[22218]_ ;
  assign \new_[22222]_  = ~A201 & A200;
  assign \new_[22225]_  = ~A232 & ~A203;
  assign \new_[22226]_  = \new_[22225]_  & \new_[22222]_ ;
  assign \new_[22227]_  = \new_[22226]_  & \new_[22219]_ ;
  assign \new_[22231]_  = A236 & ~A235;
  assign \new_[22232]_  = A233 & \new_[22231]_ ;
  assign \new_[22235]_  = A299 & ~A298;
  assign \new_[22238]_  = A302 & ~A301;
  assign \new_[22239]_  = \new_[22238]_  & \new_[22235]_ ;
  assign \new_[22240]_  = \new_[22239]_  & \new_[22232]_ ;
  assign \new_[22244]_  = ~A199 & ~A166;
  assign \new_[22245]_  = A167 & \new_[22244]_ ;
  assign \new_[22248]_  = ~A201 & A200;
  assign \new_[22251]_  = ~A232 & ~A203;
  assign \new_[22252]_  = \new_[22251]_  & \new_[22248]_ ;
  assign \new_[22253]_  = \new_[22252]_  & \new_[22245]_ ;
  assign \new_[22257]_  = A236 & ~A235;
  assign \new_[22258]_  = A233 & \new_[22257]_ ;
  assign \new_[22261]_  = ~A299 & ~A298;
  assign \new_[22264]_  = ~A302 & A301;
  assign \new_[22265]_  = \new_[22264]_  & \new_[22261]_ ;
  assign \new_[22266]_  = \new_[22265]_  & \new_[22258]_ ;
  assign \new_[22270]_  = ~A199 & ~A166;
  assign \new_[22271]_  = A167 & \new_[22270]_ ;
  assign \new_[22274]_  = ~A201 & A200;
  assign \new_[22277]_  = ~A232 & ~A203;
  assign \new_[22278]_  = \new_[22277]_  & \new_[22274]_ ;
  assign \new_[22279]_  = \new_[22278]_  & \new_[22271]_ ;
  assign \new_[22283]_  = A236 & ~A235;
  assign \new_[22284]_  = A233 & \new_[22283]_ ;
  assign \new_[22287]_  = A266 & A265;
  assign \new_[22290]_  = ~A269 & A268;
  assign \new_[22291]_  = \new_[22290]_  & \new_[22287]_ ;
  assign \new_[22292]_  = \new_[22291]_  & \new_[22284]_ ;
  assign \new_[22296]_  = ~A199 & ~A166;
  assign \new_[22297]_  = A167 & \new_[22296]_ ;
  assign \new_[22300]_  = ~A201 & A200;
  assign \new_[22303]_  = ~A232 & ~A203;
  assign \new_[22304]_  = \new_[22303]_  & \new_[22300]_ ;
  assign \new_[22305]_  = \new_[22304]_  & \new_[22297]_ ;
  assign \new_[22309]_  = A236 & ~A235;
  assign \new_[22310]_  = A233 & \new_[22309]_ ;
  assign \new_[22313]_  = A266 & ~A265;
  assign \new_[22316]_  = A269 & ~A268;
  assign \new_[22317]_  = \new_[22316]_  & \new_[22313]_ ;
  assign \new_[22318]_  = \new_[22317]_  & \new_[22310]_ ;
  assign \new_[22322]_  = ~A199 & ~A166;
  assign \new_[22323]_  = A167 & \new_[22322]_ ;
  assign \new_[22326]_  = ~A201 & A200;
  assign \new_[22329]_  = ~A232 & ~A203;
  assign \new_[22330]_  = \new_[22329]_  & \new_[22326]_ ;
  assign \new_[22331]_  = \new_[22330]_  & \new_[22323]_ ;
  assign \new_[22335]_  = A236 & ~A235;
  assign \new_[22336]_  = A233 & \new_[22335]_ ;
  assign \new_[22339]_  = ~A266 & A265;
  assign \new_[22342]_  = A269 & ~A268;
  assign \new_[22343]_  = \new_[22342]_  & \new_[22339]_ ;
  assign \new_[22344]_  = \new_[22343]_  & \new_[22336]_ ;
  assign \new_[22348]_  = ~A199 & ~A166;
  assign \new_[22349]_  = A167 & \new_[22348]_ ;
  assign \new_[22352]_  = ~A201 & A200;
  assign \new_[22355]_  = ~A232 & ~A203;
  assign \new_[22356]_  = \new_[22355]_  & \new_[22352]_ ;
  assign \new_[22357]_  = \new_[22356]_  & \new_[22349]_ ;
  assign \new_[22361]_  = A236 & ~A235;
  assign \new_[22362]_  = A233 & \new_[22361]_ ;
  assign \new_[22365]_  = ~A266 & ~A265;
  assign \new_[22368]_  = ~A269 & A268;
  assign \new_[22369]_  = \new_[22368]_  & \new_[22365]_ ;
  assign \new_[22370]_  = \new_[22369]_  & \new_[22362]_ ;
  assign \new_[22374]_  = ~A199 & ~A166;
  assign \new_[22375]_  = A167 & \new_[22374]_ ;
  assign \new_[22378]_  = ~A201 & A200;
  assign \new_[22381]_  = A232 & ~A203;
  assign \new_[22382]_  = \new_[22381]_  & \new_[22378]_ ;
  assign \new_[22383]_  = \new_[22382]_  & \new_[22375]_ ;
  assign \new_[22387]_  = A236 & ~A235;
  assign \new_[22388]_  = ~A233 & \new_[22387]_ ;
  assign \new_[22391]_  = A299 & A298;
  assign \new_[22394]_  = ~A302 & A301;
  assign \new_[22395]_  = \new_[22394]_  & \new_[22391]_ ;
  assign \new_[22396]_  = \new_[22395]_  & \new_[22388]_ ;
  assign \new_[22400]_  = ~A199 & ~A166;
  assign \new_[22401]_  = A167 & \new_[22400]_ ;
  assign \new_[22404]_  = ~A201 & A200;
  assign \new_[22407]_  = A232 & ~A203;
  assign \new_[22408]_  = \new_[22407]_  & \new_[22404]_ ;
  assign \new_[22409]_  = \new_[22408]_  & \new_[22401]_ ;
  assign \new_[22413]_  = A236 & ~A235;
  assign \new_[22414]_  = ~A233 & \new_[22413]_ ;
  assign \new_[22417]_  = ~A299 & A298;
  assign \new_[22420]_  = A302 & ~A301;
  assign \new_[22421]_  = \new_[22420]_  & \new_[22417]_ ;
  assign \new_[22422]_  = \new_[22421]_  & \new_[22414]_ ;
  assign \new_[22426]_  = ~A199 & ~A166;
  assign \new_[22427]_  = A167 & \new_[22426]_ ;
  assign \new_[22430]_  = ~A201 & A200;
  assign \new_[22433]_  = A232 & ~A203;
  assign \new_[22434]_  = \new_[22433]_  & \new_[22430]_ ;
  assign \new_[22435]_  = \new_[22434]_  & \new_[22427]_ ;
  assign \new_[22439]_  = A236 & ~A235;
  assign \new_[22440]_  = ~A233 & \new_[22439]_ ;
  assign \new_[22443]_  = A299 & ~A298;
  assign \new_[22446]_  = A302 & ~A301;
  assign \new_[22447]_  = \new_[22446]_  & \new_[22443]_ ;
  assign \new_[22448]_  = \new_[22447]_  & \new_[22440]_ ;
  assign \new_[22452]_  = ~A199 & ~A166;
  assign \new_[22453]_  = A167 & \new_[22452]_ ;
  assign \new_[22456]_  = ~A201 & A200;
  assign \new_[22459]_  = A232 & ~A203;
  assign \new_[22460]_  = \new_[22459]_  & \new_[22456]_ ;
  assign \new_[22461]_  = \new_[22460]_  & \new_[22453]_ ;
  assign \new_[22465]_  = A236 & ~A235;
  assign \new_[22466]_  = ~A233 & \new_[22465]_ ;
  assign \new_[22469]_  = ~A299 & ~A298;
  assign \new_[22472]_  = ~A302 & A301;
  assign \new_[22473]_  = \new_[22472]_  & \new_[22469]_ ;
  assign \new_[22474]_  = \new_[22473]_  & \new_[22466]_ ;
  assign \new_[22478]_  = ~A199 & ~A166;
  assign \new_[22479]_  = A167 & \new_[22478]_ ;
  assign \new_[22482]_  = ~A201 & A200;
  assign \new_[22485]_  = A232 & ~A203;
  assign \new_[22486]_  = \new_[22485]_  & \new_[22482]_ ;
  assign \new_[22487]_  = \new_[22486]_  & \new_[22479]_ ;
  assign \new_[22491]_  = A236 & ~A235;
  assign \new_[22492]_  = ~A233 & \new_[22491]_ ;
  assign \new_[22495]_  = A266 & A265;
  assign \new_[22498]_  = ~A269 & A268;
  assign \new_[22499]_  = \new_[22498]_  & \new_[22495]_ ;
  assign \new_[22500]_  = \new_[22499]_  & \new_[22492]_ ;
  assign \new_[22504]_  = ~A199 & ~A166;
  assign \new_[22505]_  = A167 & \new_[22504]_ ;
  assign \new_[22508]_  = ~A201 & A200;
  assign \new_[22511]_  = A232 & ~A203;
  assign \new_[22512]_  = \new_[22511]_  & \new_[22508]_ ;
  assign \new_[22513]_  = \new_[22512]_  & \new_[22505]_ ;
  assign \new_[22517]_  = A236 & ~A235;
  assign \new_[22518]_  = ~A233 & \new_[22517]_ ;
  assign \new_[22521]_  = A266 & ~A265;
  assign \new_[22524]_  = A269 & ~A268;
  assign \new_[22525]_  = \new_[22524]_  & \new_[22521]_ ;
  assign \new_[22526]_  = \new_[22525]_  & \new_[22518]_ ;
  assign \new_[22530]_  = ~A199 & ~A166;
  assign \new_[22531]_  = A167 & \new_[22530]_ ;
  assign \new_[22534]_  = ~A201 & A200;
  assign \new_[22537]_  = A232 & ~A203;
  assign \new_[22538]_  = \new_[22537]_  & \new_[22534]_ ;
  assign \new_[22539]_  = \new_[22538]_  & \new_[22531]_ ;
  assign \new_[22543]_  = A236 & ~A235;
  assign \new_[22544]_  = ~A233 & \new_[22543]_ ;
  assign \new_[22547]_  = ~A266 & A265;
  assign \new_[22550]_  = A269 & ~A268;
  assign \new_[22551]_  = \new_[22550]_  & \new_[22547]_ ;
  assign \new_[22552]_  = \new_[22551]_  & \new_[22544]_ ;
  assign \new_[22556]_  = ~A199 & ~A166;
  assign \new_[22557]_  = A167 & \new_[22556]_ ;
  assign \new_[22560]_  = ~A201 & A200;
  assign \new_[22563]_  = A232 & ~A203;
  assign \new_[22564]_  = \new_[22563]_  & \new_[22560]_ ;
  assign \new_[22565]_  = \new_[22564]_  & \new_[22557]_ ;
  assign \new_[22569]_  = A236 & ~A235;
  assign \new_[22570]_  = ~A233 & \new_[22569]_ ;
  assign \new_[22573]_  = ~A266 & ~A265;
  assign \new_[22576]_  = ~A269 & A268;
  assign \new_[22577]_  = \new_[22576]_  & \new_[22573]_ ;
  assign \new_[22578]_  = \new_[22577]_  & \new_[22570]_ ;
  assign \new_[22582]_  = ~A199 & ~A166;
  assign \new_[22583]_  = A167 & \new_[22582]_ ;
  assign \new_[22586]_  = ~A201 & A200;
  assign \new_[22589]_  = ~A232 & ~A203;
  assign \new_[22590]_  = \new_[22589]_  & \new_[22586]_ ;
  assign \new_[22591]_  = \new_[22590]_  & \new_[22583]_ ;
  assign \new_[22595]_  = ~A236 & A235;
  assign \new_[22596]_  = ~A233 & \new_[22595]_ ;
  assign \new_[22599]_  = A299 & A298;
  assign \new_[22602]_  = ~A302 & A301;
  assign \new_[22603]_  = \new_[22602]_  & \new_[22599]_ ;
  assign \new_[22604]_  = \new_[22603]_  & \new_[22596]_ ;
  assign \new_[22608]_  = ~A199 & ~A166;
  assign \new_[22609]_  = A167 & \new_[22608]_ ;
  assign \new_[22612]_  = ~A201 & A200;
  assign \new_[22615]_  = ~A232 & ~A203;
  assign \new_[22616]_  = \new_[22615]_  & \new_[22612]_ ;
  assign \new_[22617]_  = \new_[22616]_  & \new_[22609]_ ;
  assign \new_[22621]_  = ~A236 & A235;
  assign \new_[22622]_  = ~A233 & \new_[22621]_ ;
  assign \new_[22625]_  = ~A299 & A298;
  assign \new_[22628]_  = A302 & ~A301;
  assign \new_[22629]_  = \new_[22628]_  & \new_[22625]_ ;
  assign \new_[22630]_  = \new_[22629]_  & \new_[22622]_ ;
  assign \new_[22634]_  = ~A199 & ~A166;
  assign \new_[22635]_  = A167 & \new_[22634]_ ;
  assign \new_[22638]_  = ~A201 & A200;
  assign \new_[22641]_  = ~A232 & ~A203;
  assign \new_[22642]_  = \new_[22641]_  & \new_[22638]_ ;
  assign \new_[22643]_  = \new_[22642]_  & \new_[22635]_ ;
  assign \new_[22647]_  = ~A236 & A235;
  assign \new_[22648]_  = ~A233 & \new_[22647]_ ;
  assign \new_[22651]_  = A299 & ~A298;
  assign \new_[22654]_  = A302 & ~A301;
  assign \new_[22655]_  = \new_[22654]_  & \new_[22651]_ ;
  assign \new_[22656]_  = \new_[22655]_  & \new_[22648]_ ;
  assign \new_[22660]_  = ~A199 & ~A166;
  assign \new_[22661]_  = A167 & \new_[22660]_ ;
  assign \new_[22664]_  = ~A201 & A200;
  assign \new_[22667]_  = ~A232 & ~A203;
  assign \new_[22668]_  = \new_[22667]_  & \new_[22664]_ ;
  assign \new_[22669]_  = \new_[22668]_  & \new_[22661]_ ;
  assign \new_[22673]_  = ~A236 & A235;
  assign \new_[22674]_  = ~A233 & \new_[22673]_ ;
  assign \new_[22677]_  = ~A299 & ~A298;
  assign \new_[22680]_  = ~A302 & A301;
  assign \new_[22681]_  = \new_[22680]_  & \new_[22677]_ ;
  assign \new_[22682]_  = \new_[22681]_  & \new_[22674]_ ;
  assign \new_[22686]_  = ~A199 & ~A166;
  assign \new_[22687]_  = A167 & \new_[22686]_ ;
  assign \new_[22690]_  = ~A201 & A200;
  assign \new_[22693]_  = ~A232 & ~A203;
  assign \new_[22694]_  = \new_[22693]_  & \new_[22690]_ ;
  assign \new_[22695]_  = \new_[22694]_  & \new_[22687]_ ;
  assign \new_[22699]_  = ~A236 & A235;
  assign \new_[22700]_  = ~A233 & \new_[22699]_ ;
  assign \new_[22703]_  = A266 & A265;
  assign \new_[22706]_  = ~A269 & A268;
  assign \new_[22707]_  = \new_[22706]_  & \new_[22703]_ ;
  assign \new_[22708]_  = \new_[22707]_  & \new_[22700]_ ;
  assign \new_[22712]_  = ~A199 & ~A166;
  assign \new_[22713]_  = A167 & \new_[22712]_ ;
  assign \new_[22716]_  = ~A201 & A200;
  assign \new_[22719]_  = ~A232 & ~A203;
  assign \new_[22720]_  = \new_[22719]_  & \new_[22716]_ ;
  assign \new_[22721]_  = \new_[22720]_  & \new_[22713]_ ;
  assign \new_[22725]_  = ~A236 & A235;
  assign \new_[22726]_  = ~A233 & \new_[22725]_ ;
  assign \new_[22729]_  = A266 & ~A265;
  assign \new_[22732]_  = A269 & ~A268;
  assign \new_[22733]_  = \new_[22732]_  & \new_[22729]_ ;
  assign \new_[22734]_  = \new_[22733]_  & \new_[22726]_ ;
  assign \new_[22738]_  = ~A199 & ~A166;
  assign \new_[22739]_  = A167 & \new_[22738]_ ;
  assign \new_[22742]_  = ~A201 & A200;
  assign \new_[22745]_  = ~A232 & ~A203;
  assign \new_[22746]_  = \new_[22745]_  & \new_[22742]_ ;
  assign \new_[22747]_  = \new_[22746]_  & \new_[22739]_ ;
  assign \new_[22751]_  = ~A236 & A235;
  assign \new_[22752]_  = ~A233 & \new_[22751]_ ;
  assign \new_[22755]_  = ~A266 & A265;
  assign \new_[22758]_  = A269 & ~A268;
  assign \new_[22759]_  = \new_[22758]_  & \new_[22755]_ ;
  assign \new_[22760]_  = \new_[22759]_  & \new_[22752]_ ;
  assign \new_[22764]_  = ~A199 & ~A166;
  assign \new_[22765]_  = A167 & \new_[22764]_ ;
  assign \new_[22768]_  = ~A201 & A200;
  assign \new_[22771]_  = ~A232 & ~A203;
  assign \new_[22772]_  = \new_[22771]_  & \new_[22768]_ ;
  assign \new_[22773]_  = \new_[22772]_  & \new_[22765]_ ;
  assign \new_[22777]_  = ~A236 & A235;
  assign \new_[22778]_  = ~A233 & \new_[22777]_ ;
  assign \new_[22781]_  = ~A266 & ~A265;
  assign \new_[22784]_  = ~A269 & A268;
  assign \new_[22785]_  = \new_[22784]_  & \new_[22781]_ ;
  assign \new_[22786]_  = \new_[22785]_  & \new_[22778]_ ;
  assign \new_[22790]_  = A199 & ~A166;
  assign \new_[22791]_  = A167 & \new_[22790]_ ;
  assign \new_[22794]_  = ~A201 & ~A200;
  assign \new_[22797]_  = A232 & A202;
  assign \new_[22798]_  = \new_[22797]_  & \new_[22794]_ ;
  assign \new_[22799]_  = \new_[22798]_  & \new_[22791]_ ;
  assign \new_[22803]_  = ~A236 & A235;
  assign \new_[22804]_  = A233 & \new_[22803]_ ;
  assign \new_[22807]_  = A299 & A298;
  assign \new_[22810]_  = ~A302 & A301;
  assign \new_[22811]_  = \new_[22810]_  & \new_[22807]_ ;
  assign \new_[22812]_  = \new_[22811]_  & \new_[22804]_ ;
  assign \new_[22816]_  = A199 & ~A166;
  assign \new_[22817]_  = A167 & \new_[22816]_ ;
  assign \new_[22820]_  = ~A201 & ~A200;
  assign \new_[22823]_  = A232 & A202;
  assign \new_[22824]_  = \new_[22823]_  & \new_[22820]_ ;
  assign \new_[22825]_  = \new_[22824]_  & \new_[22817]_ ;
  assign \new_[22829]_  = ~A236 & A235;
  assign \new_[22830]_  = A233 & \new_[22829]_ ;
  assign \new_[22833]_  = ~A299 & A298;
  assign \new_[22836]_  = A302 & ~A301;
  assign \new_[22837]_  = \new_[22836]_  & \new_[22833]_ ;
  assign \new_[22838]_  = \new_[22837]_  & \new_[22830]_ ;
  assign \new_[22842]_  = A199 & ~A166;
  assign \new_[22843]_  = A167 & \new_[22842]_ ;
  assign \new_[22846]_  = ~A201 & ~A200;
  assign \new_[22849]_  = A232 & A202;
  assign \new_[22850]_  = \new_[22849]_  & \new_[22846]_ ;
  assign \new_[22851]_  = \new_[22850]_  & \new_[22843]_ ;
  assign \new_[22855]_  = ~A236 & A235;
  assign \new_[22856]_  = A233 & \new_[22855]_ ;
  assign \new_[22859]_  = A299 & ~A298;
  assign \new_[22862]_  = A302 & ~A301;
  assign \new_[22863]_  = \new_[22862]_  & \new_[22859]_ ;
  assign \new_[22864]_  = \new_[22863]_  & \new_[22856]_ ;
  assign \new_[22868]_  = A199 & ~A166;
  assign \new_[22869]_  = A167 & \new_[22868]_ ;
  assign \new_[22872]_  = ~A201 & ~A200;
  assign \new_[22875]_  = A232 & A202;
  assign \new_[22876]_  = \new_[22875]_  & \new_[22872]_ ;
  assign \new_[22877]_  = \new_[22876]_  & \new_[22869]_ ;
  assign \new_[22881]_  = ~A236 & A235;
  assign \new_[22882]_  = A233 & \new_[22881]_ ;
  assign \new_[22885]_  = ~A299 & ~A298;
  assign \new_[22888]_  = ~A302 & A301;
  assign \new_[22889]_  = \new_[22888]_  & \new_[22885]_ ;
  assign \new_[22890]_  = \new_[22889]_  & \new_[22882]_ ;
  assign \new_[22894]_  = A199 & ~A166;
  assign \new_[22895]_  = A167 & \new_[22894]_ ;
  assign \new_[22898]_  = ~A201 & ~A200;
  assign \new_[22901]_  = A232 & A202;
  assign \new_[22902]_  = \new_[22901]_  & \new_[22898]_ ;
  assign \new_[22903]_  = \new_[22902]_  & \new_[22895]_ ;
  assign \new_[22907]_  = ~A236 & A235;
  assign \new_[22908]_  = A233 & \new_[22907]_ ;
  assign \new_[22911]_  = A266 & A265;
  assign \new_[22914]_  = ~A269 & A268;
  assign \new_[22915]_  = \new_[22914]_  & \new_[22911]_ ;
  assign \new_[22916]_  = \new_[22915]_  & \new_[22908]_ ;
  assign \new_[22920]_  = A199 & ~A166;
  assign \new_[22921]_  = A167 & \new_[22920]_ ;
  assign \new_[22924]_  = ~A201 & ~A200;
  assign \new_[22927]_  = A232 & A202;
  assign \new_[22928]_  = \new_[22927]_  & \new_[22924]_ ;
  assign \new_[22929]_  = \new_[22928]_  & \new_[22921]_ ;
  assign \new_[22933]_  = ~A236 & A235;
  assign \new_[22934]_  = A233 & \new_[22933]_ ;
  assign \new_[22937]_  = A266 & ~A265;
  assign \new_[22940]_  = A269 & ~A268;
  assign \new_[22941]_  = \new_[22940]_  & \new_[22937]_ ;
  assign \new_[22942]_  = \new_[22941]_  & \new_[22934]_ ;
  assign \new_[22946]_  = A199 & ~A166;
  assign \new_[22947]_  = A167 & \new_[22946]_ ;
  assign \new_[22950]_  = ~A201 & ~A200;
  assign \new_[22953]_  = A232 & A202;
  assign \new_[22954]_  = \new_[22953]_  & \new_[22950]_ ;
  assign \new_[22955]_  = \new_[22954]_  & \new_[22947]_ ;
  assign \new_[22959]_  = ~A236 & A235;
  assign \new_[22960]_  = A233 & \new_[22959]_ ;
  assign \new_[22963]_  = ~A266 & A265;
  assign \new_[22966]_  = A269 & ~A268;
  assign \new_[22967]_  = \new_[22966]_  & \new_[22963]_ ;
  assign \new_[22968]_  = \new_[22967]_  & \new_[22960]_ ;
  assign \new_[22972]_  = A199 & ~A166;
  assign \new_[22973]_  = A167 & \new_[22972]_ ;
  assign \new_[22976]_  = ~A201 & ~A200;
  assign \new_[22979]_  = A232 & A202;
  assign \new_[22980]_  = \new_[22979]_  & \new_[22976]_ ;
  assign \new_[22981]_  = \new_[22980]_  & \new_[22973]_ ;
  assign \new_[22985]_  = ~A236 & A235;
  assign \new_[22986]_  = A233 & \new_[22985]_ ;
  assign \new_[22989]_  = ~A266 & ~A265;
  assign \new_[22992]_  = ~A269 & A268;
  assign \new_[22993]_  = \new_[22992]_  & \new_[22989]_ ;
  assign \new_[22994]_  = \new_[22993]_  & \new_[22986]_ ;
  assign \new_[22998]_  = A199 & ~A166;
  assign \new_[22999]_  = A167 & \new_[22998]_ ;
  assign \new_[23002]_  = ~A201 & ~A200;
  assign \new_[23005]_  = ~A232 & A202;
  assign \new_[23006]_  = \new_[23005]_  & \new_[23002]_ ;
  assign \new_[23007]_  = \new_[23006]_  & \new_[22999]_ ;
  assign \new_[23011]_  = A236 & ~A235;
  assign \new_[23012]_  = A233 & \new_[23011]_ ;
  assign \new_[23015]_  = A299 & A298;
  assign \new_[23018]_  = ~A302 & A301;
  assign \new_[23019]_  = \new_[23018]_  & \new_[23015]_ ;
  assign \new_[23020]_  = \new_[23019]_  & \new_[23012]_ ;
  assign \new_[23024]_  = A199 & ~A166;
  assign \new_[23025]_  = A167 & \new_[23024]_ ;
  assign \new_[23028]_  = ~A201 & ~A200;
  assign \new_[23031]_  = ~A232 & A202;
  assign \new_[23032]_  = \new_[23031]_  & \new_[23028]_ ;
  assign \new_[23033]_  = \new_[23032]_  & \new_[23025]_ ;
  assign \new_[23037]_  = A236 & ~A235;
  assign \new_[23038]_  = A233 & \new_[23037]_ ;
  assign \new_[23041]_  = ~A299 & A298;
  assign \new_[23044]_  = A302 & ~A301;
  assign \new_[23045]_  = \new_[23044]_  & \new_[23041]_ ;
  assign \new_[23046]_  = \new_[23045]_  & \new_[23038]_ ;
  assign \new_[23050]_  = A199 & ~A166;
  assign \new_[23051]_  = A167 & \new_[23050]_ ;
  assign \new_[23054]_  = ~A201 & ~A200;
  assign \new_[23057]_  = ~A232 & A202;
  assign \new_[23058]_  = \new_[23057]_  & \new_[23054]_ ;
  assign \new_[23059]_  = \new_[23058]_  & \new_[23051]_ ;
  assign \new_[23063]_  = A236 & ~A235;
  assign \new_[23064]_  = A233 & \new_[23063]_ ;
  assign \new_[23067]_  = A299 & ~A298;
  assign \new_[23070]_  = A302 & ~A301;
  assign \new_[23071]_  = \new_[23070]_  & \new_[23067]_ ;
  assign \new_[23072]_  = \new_[23071]_  & \new_[23064]_ ;
  assign \new_[23076]_  = A199 & ~A166;
  assign \new_[23077]_  = A167 & \new_[23076]_ ;
  assign \new_[23080]_  = ~A201 & ~A200;
  assign \new_[23083]_  = ~A232 & A202;
  assign \new_[23084]_  = \new_[23083]_  & \new_[23080]_ ;
  assign \new_[23085]_  = \new_[23084]_  & \new_[23077]_ ;
  assign \new_[23089]_  = A236 & ~A235;
  assign \new_[23090]_  = A233 & \new_[23089]_ ;
  assign \new_[23093]_  = ~A299 & ~A298;
  assign \new_[23096]_  = ~A302 & A301;
  assign \new_[23097]_  = \new_[23096]_  & \new_[23093]_ ;
  assign \new_[23098]_  = \new_[23097]_  & \new_[23090]_ ;
  assign \new_[23102]_  = A199 & ~A166;
  assign \new_[23103]_  = A167 & \new_[23102]_ ;
  assign \new_[23106]_  = ~A201 & ~A200;
  assign \new_[23109]_  = ~A232 & A202;
  assign \new_[23110]_  = \new_[23109]_  & \new_[23106]_ ;
  assign \new_[23111]_  = \new_[23110]_  & \new_[23103]_ ;
  assign \new_[23115]_  = A236 & ~A235;
  assign \new_[23116]_  = A233 & \new_[23115]_ ;
  assign \new_[23119]_  = A266 & A265;
  assign \new_[23122]_  = ~A269 & A268;
  assign \new_[23123]_  = \new_[23122]_  & \new_[23119]_ ;
  assign \new_[23124]_  = \new_[23123]_  & \new_[23116]_ ;
  assign \new_[23128]_  = A199 & ~A166;
  assign \new_[23129]_  = A167 & \new_[23128]_ ;
  assign \new_[23132]_  = ~A201 & ~A200;
  assign \new_[23135]_  = ~A232 & A202;
  assign \new_[23136]_  = \new_[23135]_  & \new_[23132]_ ;
  assign \new_[23137]_  = \new_[23136]_  & \new_[23129]_ ;
  assign \new_[23141]_  = A236 & ~A235;
  assign \new_[23142]_  = A233 & \new_[23141]_ ;
  assign \new_[23145]_  = A266 & ~A265;
  assign \new_[23148]_  = A269 & ~A268;
  assign \new_[23149]_  = \new_[23148]_  & \new_[23145]_ ;
  assign \new_[23150]_  = \new_[23149]_  & \new_[23142]_ ;
  assign \new_[23154]_  = A199 & ~A166;
  assign \new_[23155]_  = A167 & \new_[23154]_ ;
  assign \new_[23158]_  = ~A201 & ~A200;
  assign \new_[23161]_  = ~A232 & A202;
  assign \new_[23162]_  = \new_[23161]_  & \new_[23158]_ ;
  assign \new_[23163]_  = \new_[23162]_  & \new_[23155]_ ;
  assign \new_[23167]_  = A236 & ~A235;
  assign \new_[23168]_  = A233 & \new_[23167]_ ;
  assign \new_[23171]_  = ~A266 & A265;
  assign \new_[23174]_  = A269 & ~A268;
  assign \new_[23175]_  = \new_[23174]_  & \new_[23171]_ ;
  assign \new_[23176]_  = \new_[23175]_  & \new_[23168]_ ;
  assign \new_[23180]_  = A199 & ~A166;
  assign \new_[23181]_  = A167 & \new_[23180]_ ;
  assign \new_[23184]_  = ~A201 & ~A200;
  assign \new_[23187]_  = ~A232 & A202;
  assign \new_[23188]_  = \new_[23187]_  & \new_[23184]_ ;
  assign \new_[23189]_  = \new_[23188]_  & \new_[23181]_ ;
  assign \new_[23193]_  = A236 & ~A235;
  assign \new_[23194]_  = A233 & \new_[23193]_ ;
  assign \new_[23197]_  = ~A266 & ~A265;
  assign \new_[23200]_  = ~A269 & A268;
  assign \new_[23201]_  = \new_[23200]_  & \new_[23197]_ ;
  assign \new_[23202]_  = \new_[23201]_  & \new_[23194]_ ;
  assign \new_[23206]_  = A199 & ~A166;
  assign \new_[23207]_  = A167 & \new_[23206]_ ;
  assign \new_[23210]_  = ~A201 & ~A200;
  assign \new_[23213]_  = A232 & A202;
  assign \new_[23214]_  = \new_[23213]_  & \new_[23210]_ ;
  assign \new_[23215]_  = \new_[23214]_  & \new_[23207]_ ;
  assign \new_[23219]_  = A236 & ~A235;
  assign \new_[23220]_  = ~A233 & \new_[23219]_ ;
  assign \new_[23223]_  = A299 & A298;
  assign \new_[23226]_  = ~A302 & A301;
  assign \new_[23227]_  = \new_[23226]_  & \new_[23223]_ ;
  assign \new_[23228]_  = \new_[23227]_  & \new_[23220]_ ;
  assign \new_[23232]_  = A199 & ~A166;
  assign \new_[23233]_  = A167 & \new_[23232]_ ;
  assign \new_[23236]_  = ~A201 & ~A200;
  assign \new_[23239]_  = A232 & A202;
  assign \new_[23240]_  = \new_[23239]_  & \new_[23236]_ ;
  assign \new_[23241]_  = \new_[23240]_  & \new_[23233]_ ;
  assign \new_[23245]_  = A236 & ~A235;
  assign \new_[23246]_  = ~A233 & \new_[23245]_ ;
  assign \new_[23249]_  = ~A299 & A298;
  assign \new_[23252]_  = A302 & ~A301;
  assign \new_[23253]_  = \new_[23252]_  & \new_[23249]_ ;
  assign \new_[23254]_  = \new_[23253]_  & \new_[23246]_ ;
  assign \new_[23258]_  = A199 & ~A166;
  assign \new_[23259]_  = A167 & \new_[23258]_ ;
  assign \new_[23262]_  = ~A201 & ~A200;
  assign \new_[23265]_  = A232 & A202;
  assign \new_[23266]_  = \new_[23265]_  & \new_[23262]_ ;
  assign \new_[23267]_  = \new_[23266]_  & \new_[23259]_ ;
  assign \new_[23271]_  = A236 & ~A235;
  assign \new_[23272]_  = ~A233 & \new_[23271]_ ;
  assign \new_[23275]_  = A299 & ~A298;
  assign \new_[23278]_  = A302 & ~A301;
  assign \new_[23279]_  = \new_[23278]_  & \new_[23275]_ ;
  assign \new_[23280]_  = \new_[23279]_  & \new_[23272]_ ;
  assign \new_[23284]_  = A199 & ~A166;
  assign \new_[23285]_  = A167 & \new_[23284]_ ;
  assign \new_[23288]_  = ~A201 & ~A200;
  assign \new_[23291]_  = A232 & A202;
  assign \new_[23292]_  = \new_[23291]_  & \new_[23288]_ ;
  assign \new_[23293]_  = \new_[23292]_  & \new_[23285]_ ;
  assign \new_[23297]_  = A236 & ~A235;
  assign \new_[23298]_  = ~A233 & \new_[23297]_ ;
  assign \new_[23301]_  = ~A299 & ~A298;
  assign \new_[23304]_  = ~A302 & A301;
  assign \new_[23305]_  = \new_[23304]_  & \new_[23301]_ ;
  assign \new_[23306]_  = \new_[23305]_  & \new_[23298]_ ;
  assign \new_[23310]_  = A199 & ~A166;
  assign \new_[23311]_  = A167 & \new_[23310]_ ;
  assign \new_[23314]_  = ~A201 & ~A200;
  assign \new_[23317]_  = A232 & A202;
  assign \new_[23318]_  = \new_[23317]_  & \new_[23314]_ ;
  assign \new_[23319]_  = \new_[23318]_  & \new_[23311]_ ;
  assign \new_[23323]_  = A236 & ~A235;
  assign \new_[23324]_  = ~A233 & \new_[23323]_ ;
  assign \new_[23327]_  = A266 & A265;
  assign \new_[23330]_  = ~A269 & A268;
  assign \new_[23331]_  = \new_[23330]_  & \new_[23327]_ ;
  assign \new_[23332]_  = \new_[23331]_  & \new_[23324]_ ;
  assign \new_[23336]_  = A199 & ~A166;
  assign \new_[23337]_  = A167 & \new_[23336]_ ;
  assign \new_[23340]_  = ~A201 & ~A200;
  assign \new_[23343]_  = A232 & A202;
  assign \new_[23344]_  = \new_[23343]_  & \new_[23340]_ ;
  assign \new_[23345]_  = \new_[23344]_  & \new_[23337]_ ;
  assign \new_[23349]_  = A236 & ~A235;
  assign \new_[23350]_  = ~A233 & \new_[23349]_ ;
  assign \new_[23353]_  = A266 & ~A265;
  assign \new_[23356]_  = A269 & ~A268;
  assign \new_[23357]_  = \new_[23356]_  & \new_[23353]_ ;
  assign \new_[23358]_  = \new_[23357]_  & \new_[23350]_ ;
  assign \new_[23362]_  = A199 & ~A166;
  assign \new_[23363]_  = A167 & \new_[23362]_ ;
  assign \new_[23366]_  = ~A201 & ~A200;
  assign \new_[23369]_  = A232 & A202;
  assign \new_[23370]_  = \new_[23369]_  & \new_[23366]_ ;
  assign \new_[23371]_  = \new_[23370]_  & \new_[23363]_ ;
  assign \new_[23375]_  = A236 & ~A235;
  assign \new_[23376]_  = ~A233 & \new_[23375]_ ;
  assign \new_[23379]_  = ~A266 & A265;
  assign \new_[23382]_  = A269 & ~A268;
  assign \new_[23383]_  = \new_[23382]_  & \new_[23379]_ ;
  assign \new_[23384]_  = \new_[23383]_  & \new_[23376]_ ;
  assign \new_[23388]_  = A199 & ~A166;
  assign \new_[23389]_  = A167 & \new_[23388]_ ;
  assign \new_[23392]_  = ~A201 & ~A200;
  assign \new_[23395]_  = A232 & A202;
  assign \new_[23396]_  = \new_[23395]_  & \new_[23392]_ ;
  assign \new_[23397]_  = \new_[23396]_  & \new_[23389]_ ;
  assign \new_[23401]_  = A236 & ~A235;
  assign \new_[23402]_  = ~A233 & \new_[23401]_ ;
  assign \new_[23405]_  = ~A266 & ~A265;
  assign \new_[23408]_  = ~A269 & A268;
  assign \new_[23409]_  = \new_[23408]_  & \new_[23405]_ ;
  assign \new_[23410]_  = \new_[23409]_  & \new_[23402]_ ;
  assign \new_[23414]_  = A199 & ~A166;
  assign \new_[23415]_  = A167 & \new_[23414]_ ;
  assign \new_[23418]_  = ~A201 & ~A200;
  assign \new_[23421]_  = ~A232 & A202;
  assign \new_[23422]_  = \new_[23421]_  & \new_[23418]_ ;
  assign \new_[23423]_  = \new_[23422]_  & \new_[23415]_ ;
  assign \new_[23427]_  = ~A236 & A235;
  assign \new_[23428]_  = ~A233 & \new_[23427]_ ;
  assign \new_[23431]_  = A299 & A298;
  assign \new_[23434]_  = ~A302 & A301;
  assign \new_[23435]_  = \new_[23434]_  & \new_[23431]_ ;
  assign \new_[23436]_  = \new_[23435]_  & \new_[23428]_ ;
  assign \new_[23440]_  = A199 & ~A166;
  assign \new_[23441]_  = A167 & \new_[23440]_ ;
  assign \new_[23444]_  = ~A201 & ~A200;
  assign \new_[23447]_  = ~A232 & A202;
  assign \new_[23448]_  = \new_[23447]_  & \new_[23444]_ ;
  assign \new_[23449]_  = \new_[23448]_  & \new_[23441]_ ;
  assign \new_[23453]_  = ~A236 & A235;
  assign \new_[23454]_  = ~A233 & \new_[23453]_ ;
  assign \new_[23457]_  = ~A299 & A298;
  assign \new_[23460]_  = A302 & ~A301;
  assign \new_[23461]_  = \new_[23460]_  & \new_[23457]_ ;
  assign \new_[23462]_  = \new_[23461]_  & \new_[23454]_ ;
  assign \new_[23466]_  = A199 & ~A166;
  assign \new_[23467]_  = A167 & \new_[23466]_ ;
  assign \new_[23470]_  = ~A201 & ~A200;
  assign \new_[23473]_  = ~A232 & A202;
  assign \new_[23474]_  = \new_[23473]_  & \new_[23470]_ ;
  assign \new_[23475]_  = \new_[23474]_  & \new_[23467]_ ;
  assign \new_[23479]_  = ~A236 & A235;
  assign \new_[23480]_  = ~A233 & \new_[23479]_ ;
  assign \new_[23483]_  = A299 & ~A298;
  assign \new_[23486]_  = A302 & ~A301;
  assign \new_[23487]_  = \new_[23486]_  & \new_[23483]_ ;
  assign \new_[23488]_  = \new_[23487]_  & \new_[23480]_ ;
  assign \new_[23492]_  = A199 & ~A166;
  assign \new_[23493]_  = A167 & \new_[23492]_ ;
  assign \new_[23496]_  = ~A201 & ~A200;
  assign \new_[23499]_  = ~A232 & A202;
  assign \new_[23500]_  = \new_[23499]_  & \new_[23496]_ ;
  assign \new_[23501]_  = \new_[23500]_  & \new_[23493]_ ;
  assign \new_[23505]_  = ~A236 & A235;
  assign \new_[23506]_  = ~A233 & \new_[23505]_ ;
  assign \new_[23509]_  = ~A299 & ~A298;
  assign \new_[23512]_  = ~A302 & A301;
  assign \new_[23513]_  = \new_[23512]_  & \new_[23509]_ ;
  assign \new_[23514]_  = \new_[23513]_  & \new_[23506]_ ;
  assign \new_[23518]_  = A199 & ~A166;
  assign \new_[23519]_  = A167 & \new_[23518]_ ;
  assign \new_[23522]_  = ~A201 & ~A200;
  assign \new_[23525]_  = ~A232 & A202;
  assign \new_[23526]_  = \new_[23525]_  & \new_[23522]_ ;
  assign \new_[23527]_  = \new_[23526]_  & \new_[23519]_ ;
  assign \new_[23531]_  = ~A236 & A235;
  assign \new_[23532]_  = ~A233 & \new_[23531]_ ;
  assign \new_[23535]_  = A266 & A265;
  assign \new_[23538]_  = ~A269 & A268;
  assign \new_[23539]_  = \new_[23538]_  & \new_[23535]_ ;
  assign \new_[23540]_  = \new_[23539]_  & \new_[23532]_ ;
  assign \new_[23544]_  = A199 & ~A166;
  assign \new_[23545]_  = A167 & \new_[23544]_ ;
  assign \new_[23548]_  = ~A201 & ~A200;
  assign \new_[23551]_  = ~A232 & A202;
  assign \new_[23552]_  = \new_[23551]_  & \new_[23548]_ ;
  assign \new_[23553]_  = \new_[23552]_  & \new_[23545]_ ;
  assign \new_[23557]_  = ~A236 & A235;
  assign \new_[23558]_  = ~A233 & \new_[23557]_ ;
  assign \new_[23561]_  = A266 & ~A265;
  assign \new_[23564]_  = A269 & ~A268;
  assign \new_[23565]_  = \new_[23564]_  & \new_[23561]_ ;
  assign \new_[23566]_  = \new_[23565]_  & \new_[23558]_ ;
  assign \new_[23570]_  = A199 & ~A166;
  assign \new_[23571]_  = A167 & \new_[23570]_ ;
  assign \new_[23574]_  = ~A201 & ~A200;
  assign \new_[23577]_  = ~A232 & A202;
  assign \new_[23578]_  = \new_[23577]_  & \new_[23574]_ ;
  assign \new_[23579]_  = \new_[23578]_  & \new_[23571]_ ;
  assign \new_[23583]_  = ~A236 & A235;
  assign \new_[23584]_  = ~A233 & \new_[23583]_ ;
  assign \new_[23587]_  = ~A266 & A265;
  assign \new_[23590]_  = A269 & ~A268;
  assign \new_[23591]_  = \new_[23590]_  & \new_[23587]_ ;
  assign \new_[23592]_  = \new_[23591]_  & \new_[23584]_ ;
  assign \new_[23596]_  = A199 & ~A166;
  assign \new_[23597]_  = A167 & \new_[23596]_ ;
  assign \new_[23600]_  = ~A201 & ~A200;
  assign \new_[23603]_  = ~A232 & A202;
  assign \new_[23604]_  = \new_[23603]_  & \new_[23600]_ ;
  assign \new_[23605]_  = \new_[23604]_  & \new_[23597]_ ;
  assign \new_[23609]_  = ~A236 & A235;
  assign \new_[23610]_  = ~A233 & \new_[23609]_ ;
  assign \new_[23613]_  = ~A266 & ~A265;
  assign \new_[23616]_  = ~A269 & A268;
  assign \new_[23617]_  = \new_[23616]_  & \new_[23613]_ ;
  assign \new_[23618]_  = \new_[23617]_  & \new_[23610]_ ;
  assign \new_[23622]_  = A199 & ~A166;
  assign \new_[23623]_  = A167 & \new_[23622]_ ;
  assign \new_[23626]_  = ~A201 & ~A200;
  assign \new_[23629]_  = A232 & ~A203;
  assign \new_[23630]_  = \new_[23629]_  & \new_[23626]_ ;
  assign \new_[23631]_  = \new_[23630]_  & \new_[23623]_ ;
  assign \new_[23635]_  = ~A236 & A235;
  assign \new_[23636]_  = A233 & \new_[23635]_ ;
  assign \new_[23639]_  = A299 & A298;
  assign \new_[23642]_  = ~A302 & A301;
  assign \new_[23643]_  = \new_[23642]_  & \new_[23639]_ ;
  assign \new_[23644]_  = \new_[23643]_  & \new_[23636]_ ;
  assign \new_[23648]_  = A199 & ~A166;
  assign \new_[23649]_  = A167 & \new_[23648]_ ;
  assign \new_[23652]_  = ~A201 & ~A200;
  assign \new_[23655]_  = A232 & ~A203;
  assign \new_[23656]_  = \new_[23655]_  & \new_[23652]_ ;
  assign \new_[23657]_  = \new_[23656]_  & \new_[23649]_ ;
  assign \new_[23661]_  = ~A236 & A235;
  assign \new_[23662]_  = A233 & \new_[23661]_ ;
  assign \new_[23665]_  = ~A299 & A298;
  assign \new_[23668]_  = A302 & ~A301;
  assign \new_[23669]_  = \new_[23668]_  & \new_[23665]_ ;
  assign \new_[23670]_  = \new_[23669]_  & \new_[23662]_ ;
  assign \new_[23674]_  = A199 & ~A166;
  assign \new_[23675]_  = A167 & \new_[23674]_ ;
  assign \new_[23678]_  = ~A201 & ~A200;
  assign \new_[23681]_  = A232 & ~A203;
  assign \new_[23682]_  = \new_[23681]_  & \new_[23678]_ ;
  assign \new_[23683]_  = \new_[23682]_  & \new_[23675]_ ;
  assign \new_[23687]_  = ~A236 & A235;
  assign \new_[23688]_  = A233 & \new_[23687]_ ;
  assign \new_[23691]_  = A299 & ~A298;
  assign \new_[23694]_  = A302 & ~A301;
  assign \new_[23695]_  = \new_[23694]_  & \new_[23691]_ ;
  assign \new_[23696]_  = \new_[23695]_  & \new_[23688]_ ;
  assign \new_[23700]_  = A199 & ~A166;
  assign \new_[23701]_  = A167 & \new_[23700]_ ;
  assign \new_[23704]_  = ~A201 & ~A200;
  assign \new_[23707]_  = A232 & ~A203;
  assign \new_[23708]_  = \new_[23707]_  & \new_[23704]_ ;
  assign \new_[23709]_  = \new_[23708]_  & \new_[23701]_ ;
  assign \new_[23713]_  = ~A236 & A235;
  assign \new_[23714]_  = A233 & \new_[23713]_ ;
  assign \new_[23717]_  = ~A299 & ~A298;
  assign \new_[23720]_  = ~A302 & A301;
  assign \new_[23721]_  = \new_[23720]_  & \new_[23717]_ ;
  assign \new_[23722]_  = \new_[23721]_  & \new_[23714]_ ;
  assign \new_[23726]_  = A199 & ~A166;
  assign \new_[23727]_  = A167 & \new_[23726]_ ;
  assign \new_[23730]_  = ~A201 & ~A200;
  assign \new_[23733]_  = A232 & ~A203;
  assign \new_[23734]_  = \new_[23733]_  & \new_[23730]_ ;
  assign \new_[23735]_  = \new_[23734]_  & \new_[23727]_ ;
  assign \new_[23739]_  = ~A236 & A235;
  assign \new_[23740]_  = A233 & \new_[23739]_ ;
  assign \new_[23743]_  = A266 & A265;
  assign \new_[23746]_  = ~A269 & A268;
  assign \new_[23747]_  = \new_[23746]_  & \new_[23743]_ ;
  assign \new_[23748]_  = \new_[23747]_  & \new_[23740]_ ;
  assign \new_[23752]_  = A199 & ~A166;
  assign \new_[23753]_  = A167 & \new_[23752]_ ;
  assign \new_[23756]_  = ~A201 & ~A200;
  assign \new_[23759]_  = A232 & ~A203;
  assign \new_[23760]_  = \new_[23759]_  & \new_[23756]_ ;
  assign \new_[23761]_  = \new_[23760]_  & \new_[23753]_ ;
  assign \new_[23765]_  = ~A236 & A235;
  assign \new_[23766]_  = A233 & \new_[23765]_ ;
  assign \new_[23769]_  = A266 & ~A265;
  assign \new_[23772]_  = A269 & ~A268;
  assign \new_[23773]_  = \new_[23772]_  & \new_[23769]_ ;
  assign \new_[23774]_  = \new_[23773]_  & \new_[23766]_ ;
  assign \new_[23778]_  = A199 & ~A166;
  assign \new_[23779]_  = A167 & \new_[23778]_ ;
  assign \new_[23782]_  = ~A201 & ~A200;
  assign \new_[23785]_  = A232 & ~A203;
  assign \new_[23786]_  = \new_[23785]_  & \new_[23782]_ ;
  assign \new_[23787]_  = \new_[23786]_  & \new_[23779]_ ;
  assign \new_[23791]_  = ~A236 & A235;
  assign \new_[23792]_  = A233 & \new_[23791]_ ;
  assign \new_[23795]_  = ~A266 & A265;
  assign \new_[23798]_  = A269 & ~A268;
  assign \new_[23799]_  = \new_[23798]_  & \new_[23795]_ ;
  assign \new_[23800]_  = \new_[23799]_  & \new_[23792]_ ;
  assign \new_[23804]_  = A199 & ~A166;
  assign \new_[23805]_  = A167 & \new_[23804]_ ;
  assign \new_[23808]_  = ~A201 & ~A200;
  assign \new_[23811]_  = A232 & ~A203;
  assign \new_[23812]_  = \new_[23811]_  & \new_[23808]_ ;
  assign \new_[23813]_  = \new_[23812]_  & \new_[23805]_ ;
  assign \new_[23817]_  = ~A236 & A235;
  assign \new_[23818]_  = A233 & \new_[23817]_ ;
  assign \new_[23821]_  = ~A266 & ~A265;
  assign \new_[23824]_  = ~A269 & A268;
  assign \new_[23825]_  = \new_[23824]_  & \new_[23821]_ ;
  assign \new_[23826]_  = \new_[23825]_  & \new_[23818]_ ;
  assign \new_[23830]_  = A199 & ~A166;
  assign \new_[23831]_  = A167 & \new_[23830]_ ;
  assign \new_[23834]_  = ~A201 & ~A200;
  assign \new_[23837]_  = ~A232 & ~A203;
  assign \new_[23838]_  = \new_[23837]_  & \new_[23834]_ ;
  assign \new_[23839]_  = \new_[23838]_  & \new_[23831]_ ;
  assign \new_[23843]_  = A236 & ~A235;
  assign \new_[23844]_  = A233 & \new_[23843]_ ;
  assign \new_[23847]_  = A299 & A298;
  assign \new_[23850]_  = ~A302 & A301;
  assign \new_[23851]_  = \new_[23850]_  & \new_[23847]_ ;
  assign \new_[23852]_  = \new_[23851]_  & \new_[23844]_ ;
  assign \new_[23856]_  = A199 & ~A166;
  assign \new_[23857]_  = A167 & \new_[23856]_ ;
  assign \new_[23860]_  = ~A201 & ~A200;
  assign \new_[23863]_  = ~A232 & ~A203;
  assign \new_[23864]_  = \new_[23863]_  & \new_[23860]_ ;
  assign \new_[23865]_  = \new_[23864]_  & \new_[23857]_ ;
  assign \new_[23869]_  = A236 & ~A235;
  assign \new_[23870]_  = A233 & \new_[23869]_ ;
  assign \new_[23873]_  = ~A299 & A298;
  assign \new_[23876]_  = A302 & ~A301;
  assign \new_[23877]_  = \new_[23876]_  & \new_[23873]_ ;
  assign \new_[23878]_  = \new_[23877]_  & \new_[23870]_ ;
  assign \new_[23882]_  = A199 & ~A166;
  assign \new_[23883]_  = A167 & \new_[23882]_ ;
  assign \new_[23886]_  = ~A201 & ~A200;
  assign \new_[23889]_  = ~A232 & ~A203;
  assign \new_[23890]_  = \new_[23889]_  & \new_[23886]_ ;
  assign \new_[23891]_  = \new_[23890]_  & \new_[23883]_ ;
  assign \new_[23895]_  = A236 & ~A235;
  assign \new_[23896]_  = A233 & \new_[23895]_ ;
  assign \new_[23899]_  = A299 & ~A298;
  assign \new_[23902]_  = A302 & ~A301;
  assign \new_[23903]_  = \new_[23902]_  & \new_[23899]_ ;
  assign \new_[23904]_  = \new_[23903]_  & \new_[23896]_ ;
  assign \new_[23908]_  = A199 & ~A166;
  assign \new_[23909]_  = A167 & \new_[23908]_ ;
  assign \new_[23912]_  = ~A201 & ~A200;
  assign \new_[23915]_  = ~A232 & ~A203;
  assign \new_[23916]_  = \new_[23915]_  & \new_[23912]_ ;
  assign \new_[23917]_  = \new_[23916]_  & \new_[23909]_ ;
  assign \new_[23921]_  = A236 & ~A235;
  assign \new_[23922]_  = A233 & \new_[23921]_ ;
  assign \new_[23925]_  = ~A299 & ~A298;
  assign \new_[23928]_  = ~A302 & A301;
  assign \new_[23929]_  = \new_[23928]_  & \new_[23925]_ ;
  assign \new_[23930]_  = \new_[23929]_  & \new_[23922]_ ;
  assign \new_[23934]_  = A199 & ~A166;
  assign \new_[23935]_  = A167 & \new_[23934]_ ;
  assign \new_[23938]_  = ~A201 & ~A200;
  assign \new_[23941]_  = ~A232 & ~A203;
  assign \new_[23942]_  = \new_[23941]_  & \new_[23938]_ ;
  assign \new_[23943]_  = \new_[23942]_  & \new_[23935]_ ;
  assign \new_[23947]_  = A236 & ~A235;
  assign \new_[23948]_  = A233 & \new_[23947]_ ;
  assign \new_[23951]_  = A266 & A265;
  assign \new_[23954]_  = ~A269 & A268;
  assign \new_[23955]_  = \new_[23954]_  & \new_[23951]_ ;
  assign \new_[23956]_  = \new_[23955]_  & \new_[23948]_ ;
  assign \new_[23960]_  = A199 & ~A166;
  assign \new_[23961]_  = A167 & \new_[23960]_ ;
  assign \new_[23964]_  = ~A201 & ~A200;
  assign \new_[23967]_  = ~A232 & ~A203;
  assign \new_[23968]_  = \new_[23967]_  & \new_[23964]_ ;
  assign \new_[23969]_  = \new_[23968]_  & \new_[23961]_ ;
  assign \new_[23973]_  = A236 & ~A235;
  assign \new_[23974]_  = A233 & \new_[23973]_ ;
  assign \new_[23977]_  = A266 & ~A265;
  assign \new_[23980]_  = A269 & ~A268;
  assign \new_[23981]_  = \new_[23980]_  & \new_[23977]_ ;
  assign \new_[23982]_  = \new_[23981]_  & \new_[23974]_ ;
  assign \new_[23986]_  = A199 & ~A166;
  assign \new_[23987]_  = A167 & \new_[23986]_ ;
  assign \new_[23990]_  = ~A201 & ~A200;
  assign \new_[23993]_  = ~A232 & ~A203;
  assign \new_[23994]_  = \new_[23993]_  & \new_[23990]_ ;
  assign \new_[23995]_  = \new_[23994]_  & \new_[23987]_ ;
  assign \new_[23999]_  = A236 & ~A235;
  assign \new_[24000]_  = A233 & \new_[23999]_ ;
  assign \new_[24003]_  = ~A266 & A265;
  assign \new_[24006]_  = A269 & ~A268;
  assign \new_[24007]_  = \new_[24006]_  & \new_[24003]_ ;
  assign \new_[24008]_  = \new_[24007]_  & \new_[24000]_ ;
  assign \new_[24012]_  = A199 & ~A166;
  assign \new_[24013]_  = A167 & \new_[24012]_ ;
  assign \new_[24016]_  = ~A201 & ~A200;
  assign \new_[24019]_  = ~A232 & ~A203;
  assign \new_[24020]_  = \new_[24019]_  & \new_[24016]_ ;
  assign \new_[24021]_  = \new_[24020]_  & \new_[24013]_ ;
  assign \new_[24025]_  = A236 & ~A235;
  assign \new_[24026]_  = A233 & \new_[24025]_ ;
  assign \new_[24029]_  = ~A266 & ~A265;
  assign \new_[24032]_  = ~A269 & A268;
  assign \new_[24033]_  = \new_[24032]_  & \new_[24029]_ ;
  assign \new_[24034]_  = \new_[24033]_  & \new_[24026]_ ;
  assign \new_[24038]_  = A199 & ~A166;
  assign \new_[24039]_  = A167 & \new_[24038]_ ;
  assign \new_[24042]_  = ~A201 & ~A200;
  assign \new_[24045]_  = A232 & ~A203;
  assign \new_[24046]_  = \new_[24045]_  & \new_[24042]_ ;
  assign \new_[24047]_  = \new_[24046]_  & \new_[24039]_ ;
  assign \new_[24051]_  = A236 & ~A235;
  assign \new_[24052]_  = ~A233 & \new_[24051]_ ;
  assign \new_[24055]_  = A299 & A298;
  assign \new_[24058]_  = ~A302 & A301;
  assign \new_[24059]_  = \new_[24058]_  & \new_[24055]_ ;
  assign \new_[24060]_  = \new_[24059]_  & \new_[24052]_ ;
  assign \new_[24064]_  = A199 & ~A166;
  assign \new_[24065]_  = A167 & \new_[24064]_ ;
  assign \new_[24068]_  = ~A201 & ~A200;
  assign \new_[24071]_  = A232 & ~A203;
  assign \new_[24072]_  = \new_[24071]_  & \new_[24068]_ ;
  assign \new_[24073]_  = \new_[24072]_  & \new_[24065]_ ;
  assign \new_[24077]_  = A236 & ~A235;
  assign \new_[24078]_  = ~A233 & \new_[24077]_ ;
  assign \new_[24081]_  = ~A299 & A298;
  assign \new_[24084]_  = A302 & ~A301;
  assign \new_[24085]_  = \new_[24084]_  & \new_[24081]_ ;
  assign \new_[24086]_  = \new_[24085]_  & \new_[24078]_ ;
  assign \new_[24090]_  = A199 & ~A166;
  assign \new_[24091]_  = A167 & \new_[24090]_ ;
  assign \new_[24094]_  = ~A201 & ~A200;
  assign \new_[24097]_  = A232 & ~A203;
  assign \new_[24098]_  = \new_[24097]_  & \new_[24094]_ ;
  assign \new_[24099]_  = \new_[24098]_  & \new_[24091]_ ;
  assign \new_[24103]_  = A236 & ~A235;
  assign \new_[24104]_  = ~A233 & \new_[24103]_ ;
  assign \new_[24107]_  = A299 & ~A298;
  assign \new_[24110]_  = A302 & ~A301;
  assign \new_[24111]_  = \new_[24110]_  & \new_[24107]_ ;
  assign \new_[24112]_  = \new_[24111]_  & \new_[24104]_ ;
  assign \new_[24116]_  = A199 & ~A166;
  assign \new_[24117]_  = A167 & \new_[24116]_ ;
  assign \new_[24120]_  = ~A201 & ~A200;
  assign \new_[24123]_  = A232 & ~A203;
  assign \new_[24124]_  = \new_[24123]_  & \new_[24120]_ ;
  assign \new_[24125]_  = \new_[24124]_  & \new_[24117]_ ;
  assign \new_[24129]_  = A236 & ~A235;
  assign \new_[24130]_  = ~A233 & \new_[24129]_ ;
  assign \new_[24133]_  = ~A299 & ~A298;
  assign \new_[24136]_  = ~A302 & A301;
  assign \new_[24137]_  = \new_[24136]_  & \new_[24133]_ ;
  assign \new_[24138]_  = \new_[24137]_  & \new_[24130]_ ;
  assign \new_[24142]_  = A199 & ~A166;
  assign \new_[24143]_  = A167 & \new_[24142]_ ;
  assign \new_[24146]_  = ~A201 & ~A200;
  assign \new_[24149]_  = A232 & ~A203;
  assign \new_[24150]_  = \new_[24149]_  & \new_[24146]_ ;
  assign \new_[24151]_  = \new_[24150]_  & \new_[24143]_ ;
  assign \new_[24155]_  = A236 & ~A235;
  assign \new_[24156]_  = ~A233 & \new_[24155]_ ;
  assign \new_[24159]_  = A266 & A265;
  assign \new_[24162]_  = ~A269 & A268;
  assign \new_[24163]_  = \new_[24162]_  & \new_[24159]_ ;
  assign \new_[24164]_  = \new_[24163]_  & \new_[24156]_ ;
  assign \new_[24168]_  = A199 & ~A166;
  assign \new_[24169]_  = A167 & \new_[24168]_ ;
  assign \new_[24172]_  = ~A201 & ~A200;
  assign \new_[24175]_  = A232 & ~A203;
  assign \new_[24176]_  = \new_[24175]_  & \new_[24172]_ ;
  assign \new_[24177]_  = \new_[24176]_  & \new_[24169]_ ;
  assign \new_[24181]_  = A236 & ~A235;
  assign \new_[24182]_  = ~A233 & \new_[24181]_ ;
  assign \new_[24185]_  = A266 & ~A265;
  assign \new_[24188]_  = A269 & ~A268;
  assign \new_[24189]_  = \new_[24188]_  & \new_[24185]_ ;
  assign \new_[24190]_  = \new_[24189]_  & \new_[24182]_ ;
  assign \new_[24194]_  = A199 & ~A166;
  assign \new_[24195]_  = A167 & \new_[24194]_ ;
  assign \new_[24198]_  = ~A201 & ~A200;
  assign \new_[24201]_  = A232 & ~A203;
  assign \new_[24202]_  = \new_[24201]_  & \new_[24198]_ ;
  assign \new_[24203]_  = \new_[24202]_  & \new_[24195]_ ;
  assign \new_[24207]_  = A236 & ~A235;
  assign \new_[24208]_  = ~A233 & \new_[24207]_ ;
  assign \new_[24211]_  = ~A266 & A265;
  assign \new_[24214]_  = A269 & ~A268;
  assign \new_[24215]_  = \new_[24214]_  & \new_[24211]_ ;
  assign \new_[24216]_  = \new_[24215]_  & \new_[24208]_ ;
  assign \new_[24220]_  = A199 & ~A166;
  assign \new_[24221]_  = A167 & \new_[24220]_ ;
  assign \new_[24224]_  = ~A201 & ~A200;
  assign \new_[24227]_  = A232 & ~A203;
  assign \new_[24228]_  = \new_[24227]_  & \new_[24224]_ ;
  assign \new_[24229]_  = \new_[24228]_  & \new_[24221]_ ;
  assign \new_[24233]_  = A236 & ~A235;
  assign \new_[24234]_  = ~A233 & \new_[24233]_ ;
  assign \new_[24237]_  = ~A266 & ~A265;
  assign \new_[24240]_  = ~A269 & A268;
  assign \new_[24241]_  = \new_[24240]_  & \new_[24237]_ ;
  assign \new_[24242]_  = \new_[24241]_  & \new_[24234]_ ;
  assign \new_[24246]_  = A199 & ~A166;
  assign \new_[24247]_  = A167 & \new_[24246]_ ;
  assign \new_[24250]_  = ~A201 & ~A200;
  assign \new_[24253]_  = ~A232 & ~A203;
  assign \new_[24254]_  = \new_[24253]_  & \new_[24250]_ ;
  assign \new_[24255]_  = \new_[24254]_  & \new_[24247]_ ;
  assign \new_[24259]_  = ~A236 & A235;
  assign \new_[24260]_  = ~A233 & \new_[24259]_ ;
  assign \new_[24263]_  = A299 & A298;
  assign \new_[24266]_  = ~A302 & A301;
  assign \new_[24267]_  = \new_[24266]_  & \new_[24263]_ ;
  assign \new_[24268]_  = \new_[24267]_  & \new_[24260]_ ;
  assign \new_[24272]_  = A199 & ~A166;
  assign \new_[24273]_  = A167 & \new_[24272]_ ;
  assign \new_[24276]_  = ~A201 & ~A200;
  assign \new_[24279]_  = ~A232 & ~A203;
  assign \new_[24280]_  = \new_[24279]_  & \new_[24276]_ ;
  assign \new_[24281]_  = \new_[24280]_  & \new_[24273]_ ;
  assign \new_[24285]_  = ~A236 & A235;
  assign \new_[24286]_  = ~A233 & \new_[24285]_ ;
  assign \new_[24289]_  = ~A299 & A298;
  assign \new_[24292]_  = A302 & ~A301;
  assign \new_[24293]_  = \new_[24292]_  & \new_[24289]_ ;
  assign \new_[24294]_  = \new_[24293]_  & \new_[24286]_ ;
  assign \new_[24298]_  = A199 & ~A166;
  assign \new_[24299]_  = A167 & \new_[24298]_ ;
  assign \new_[24302]_  = ~A201 & ~A200;
  assign \new_[24305]_  = ~A232 & ~A203;
  assign \new_[24306]_  = \new_[24305]_  & \new_[24302]_ ;
  assign \new_[24307]_  = \new_[24306]_  & \new_[24299]_ ;
  assign \new_[24311]_  = ~A236 & A235;
  assign \new_[24312]_  = ~A233 & \new_[24311]_ ;
  assign \new_[24315]_  = A299 & ~A298;
  assign \new_[24318]_  = A302 & ~A301;
  assign \new_[24319]_  = \new_[24318]_  & \new_[24315]_ ;
  assign \new_[24320]_  = \new_[24319]_  & \new_[24312]_ ;
  assign \new_[24324]_  = A199 & ~A166;
  assign \new_[24325]_  = A167 & \new_[24324]_ ;
  assign \new_[24328]_  = ~A201 & ~A200;
  assign \new_[24331]_  = ~A232 & ~A203;
  assign \new_[24332]_  = \new_[24331]_  & \new_[24328]_ ;
  assign \new_[24333]_  = \new_[24332]_  & \new_[24325]_ ;
  assign \new_[24337]_  = ~A236 & A235;
  assign \new_[24338]_  = ~A233 & \new_[24337]_ ;
  assign \new_[24341]_  = ~A299 & ~A298;
  assign \new_[24344]_  = ~A302 & A301;
  assign \new_[24345]_  = \new_[24344]_  & \new_[24341]_ ;
  assign \new_[24346]_  = \new_[24345]_  & \new_[24338]_ ;
  assign \new_[24350]_  = A199 & ~A166;
  assign \new_[24351]_  = A167 & \new_[24350]_ ;
  assign \new_[24354]_  = ~A201 & ~A200;
  assign \new_[24357]_  = ~A232 & ~A203;
  assign \new_[24358]_  = \new_[24357]_  & \new_[24354]_ ;
  assign \new_[24359]_  = \new_[24358]_  & \new_[24351]_ ;
  assign \new_[24363]_  = ~A236 & A235;
  assign \new_[24364]_  = ~A233 & \new_[24363]_ ;
  assign \new_[24367]_  = A266 & A265;
  assign \new_[24370]_  = ~A269 & A268;
  assign \new_[24371]_  = \new_[24370]_  & \new_[24367]_ ;
  assign \new_[24372]_  = \new_[24371]_  & \new_[24364]_ ;
  assign \new_[24376]_  = A199 & ~A166;
  assign \new_[24377]_  = A167 & \new_[24376]_ ;
  assign \new_[24380]_  = ~A201 & ~A200;
  assign \new_[24383]_  = ~A232 & ~A203;
  assign \new_[24384]_  = \new_[24383]_  & \new_[24380]_ ;
  assign \new_[24385]_  = \new_[24384]_  & \new_[24377]_ ;
  assign \new_[24389]_  = ~A236 & A235;
  assign \new_[24390]_  = ~A233 & \new_[24389]_ ;
  assign \new_[24393]_  = A266 & ~A265;
  assign \new_[24396]_  = A269 & ~A268;
  assign \new_[24397]_  = \new_[24396]_  & \new_[24393]_ ;
  assign \new_[24398]_  = \new_[24397]_  & \new_[24390]_ ;
  assign \new_[24402]_  = A199 & ~A166;
  assign \new_[24403]_  = A167 & \new_[24402]_ ;
  assign \new_[24406]_  = ~A201 & ~A200;
  assign \new_[24409]_  = ~A232 & ~A203;
  assign \new_[24410]_  = \new_[24409]_  & \new_[24406]_ ;
  assign \new_[24411]_  = \new_[24410]_  & \new_[24403]_ ;
  assign \new_[24415]_  = ~A236 & A235;
  assign \new_[24416]_  = ~A233 & \new_[24415]_ ;
  assign \new_[24419]_  = ~A266 & A265;
  assign \new_[24422]_  = A269 & ~A268;
  assign \new_[24423]_  = \new_[24422]_  & \new_[24419]_ ;
  assign \new_[24424]_  = \new_[24423]_  & \new_[24416]_ ;
  assign \new_[24428]_  = A199 & ~A166;
  assign \new_[24429]_  = A167 & \new_[24428]_ ;
  assign \new_[24432]_  = ~A201 & ~A200;
  assign \new_[24435]_  = ~A232 & ~A203;
  assign \new_[24436]_  = \new_[24435]_  & \new_[24432]_ ;
  assign \new_[24437]_  = \new_[24436]_  & \new_[24429]_ ;
  assign \new_[24441]_  = ~A236 & A235;
  assign \new_[24442]_  = ~A233 & \new_[24441]_ ;
  assign \new_[24445]_  = ~A266 & ~A265;
  assign \new_[24448]_  = ~A269 & A268;
  assign \new_[24449]_  = \new_[24448]_  & \new_[24445]_ ;
  assign \new_[24450]_  = \new_[24449]_  & \new_[24442]_ ;
  assign \new_[24454]_  = ~A167 & A168;
  assign \new_[24455]_  = A170 & \new_[24454]_ ;
  assign \new_[24458]_  = A199 & A166;
  assign \new_[24461]_  = ~A201 & A200;
  assign \new_[24462]_  = \new_[24461]_  & \new_[24458]_ ;
  assign \new_[24463]_  = \new_[24462]_  & \new_[24455]_ ;
  assign \new_[24467]_  = A234 & A232;
  assign \new_[24468]_  = ~A202 & \new_[24467]_ ;
  assign \new_[24471]_  = A299 & A298;
  assign \new_[24474]_  = ~A302 & A301;
  assign \new_[24475]_  = \new_[24474]_  & \new_[24471]_ ;
  assign \new_[24476]_  = \new_[24475]_  & \new_[24468]_ ;
  assign \new_[24480]_  = ~A167 & A168;
  assign \new_[24481]_  = A170 & \new_[24480]_ ;
  assign \new_[24484]_  = A199 & A166;
  assign \new_[24487]_  = ~A201 & A200;
  assign \new_[24488]_  = \new_[24487]_  & \new_[24484]_ ;
  assign \new_[24489]_  = \new_[24488]_  & \new_[24481]_ ;
  assign \new_[24493]_  = A234 & A232;
  assign \new_[24494]_  = ~A202 & \new_[24493]_ ;
  assign \new_[24497]_  = ~A299 & A298;
  assign \new_[24500]_  = A302 & ~A301;
  assign \new_[24501]_  = \new_[24500]_  & \new_[24497]_ ;
  assign \new_[24502]_  = \new_[24501]_  & \new_[24494]_ ;
  assign \new_[24506]_  = ~A167 & A168;
  assign \new_[24507]_  = A170 & \new_[24506]_ ;
  assign \new_[24510]_  = A199 & A166;
  assign \new_[24513]_  = ~A201 & A200;
  assign \new_[24514]_  = \new_[24513]_  & \new_[24510]_ ;
  assign \new_[24515]_  = \new_[24514]_  & \new_[24507]_ ;
  assign \new_[24519]_  = A234 & A232;
  assign \new_[24520]_  = ~A202 & \new_[24519]_ ;
  assign \new_[24523]_  = A299 & ~A298;
  assign \new_[24526]_  = A302 & ~A301;
  assign \new_[24527]_  = \new_[24526]_  & \new_[24523]_ ;
  assign \new_[24528]_  = \new_[24527]_  & \new_[24520]_ ;
  assign \new_[24532]_  = ~A167 & A168;
  assign \new_[24533]_  = A170 & \new_[24532]_ ;
  assign \new_[24536]_  = A199 & A166;
  assign \new_[24539]_  = ~A201 & A200;
  assign \new_[24540]_  = \new_[24539]_  & \new_[24536]_ ;
  assign \new_[24541]_  = \new_[24540]_  & \new_[24533]_ ;
  assign \new_[24545]_  = A234 & A232;
  assign \new_[24546]_  = ~A202 & \new_[24545]_ ;
  assign \new_[24549]_  = ~A299 & ~A298;
  assign \new_[24552]_  = ~A302 & A301;
  assign \new_[24553]_  = \new_[24552]_  & \new_[24549]_ ;
  assign \new_[24554]_  = \new_[24553]_  & \new_[24546]_ ;
  assign \new_[24558]_  = ~A167 & A168;
  assign \new_[24559]_  = A170 & \new_[24558]_ ;
  assign \new_[24562]_  = A199 & A166;
  assign \new_[24565]_  = ~A201 & A200;
  assign \new_[24566]_  = \new_[24565]_  & \new_[24562]_ ;
  assign \new_[24567]_  = \new_[24566]_  & \new_[24559]_ ;
  assign \new_[24571]_  = A234 & A232;
  assign \new_[24572]_  = ~A202 & \new_[24571]_ ;
  assign \new_[24575]_  = A266 & A265;
  assign \new_[24578]_  = ~A269 & A268;
  assign \new_[24579]_  = \new_[24578]_  & \new_[24575]_ ;
  assign \new_[24580]_  = \new_[24579]_  & \new_[24572]_ ;
  assign \new_[24584]_  = ~A167 & A168;
  assign \new_[24585]_  = A170 & \new_[24584]_ ;
  assign \new_[24588]_  = A199 & A166;
  assign \new_[24591]_  = ~A201 & A200;
  assign \new_[24592]_  = \new_[24591]_  & \new_[24588]_ ;
  assign \new_[24593]_  = \new_[24592]_  & \new_[24585]_ ;
  assign \new_[24597]_  = A234 & A232;
  assign \new_[24598]_  = ~A202 & \new_[24597]_ ;
  assign \new_[24601]_  = A266 & ~A265;
  assign \new_[24604]_  = A269 & ~A268;
  assign \new_[24605]_  = \new_[24604]_  & \new_[24601]_ ;
  assign \new_[24606]_  = \new_[24605]_  & \new_[24598]_ ;
  assign \new_[24610]_  = ~A167 & A168;
  assign \new_[24611]_  = A170 & \new_[24610]_ ;
  assign \new_[24614]_  = A199 & A166;
  assign \new_[24617]_  = ~A201 & A200;
  assign \new_[24618]_  = \new_[24617]_  & \new_[24614]_ ;
  assign \new_[24619]_  = \new_[24618]_  & \new_[24611]_ ;
  assign \new_[24623]_  = A234 & A232;
  assign \new_[24624]_  = ~A202 & \new_[24623]_ ;
  assign \new_[24627]_  = ~A266 & A265;
  assign \new_[24630]_  = A269 & ~A268;
  assign \new_[24631]_  = \new_[24630]_  & \new_[24627]_ ;
  assign \new_[24632]_  = \new_[24631]_  & \new_[24624]_ ;
  assign \new_[24636]_  = ~A167 & A168;
  assign \new_[24637]_  = A170 & \new_[24636]_ ;
  assign \new_[24640]_  = A199 & A166;
  assign \new_[24643]_  = ~A201 & A200;
  assign \new_[24644]_  = \new_[24643]_  & \new_[24640]_ ;
  assign \new_[24645]_  = \new_[24644]_  & \new_[24637]_ ;
  assign \new_[24649]_  = A234 & A232;
  assign \new_[24650]_  = ~A202 & \new_[24649]_ ;
  assign \new_[24653]_  = ~A266 & ~A265;
  assign \new_[24656]_  = ~A269 & A268;
  assign \new_[24657]_  = \new_[24656]_  & \new_[24653]_ ;
  assign \new_[24658]_  = \new_[24657]_  & \new_[24650]_ ;
  assign \new_[24662]_  = ~A167 & A168;
  assign \new_[24663]_  = A170 & \new_[24662]_ ;
  assign \new_[24666]_  = A199 & A166;
  assign \new_[24669]_  = ~A201 & A200;
  assign \new_[24670]_  = \new_[24669]_  & \new_[24666]_ ;
  assign \new_[24671]_  = \new_[24670]_  & \new_[24663]_ ;
  assign \new_[24675]_  = A234 & A233;
  assign \new_[24676]_  = ~A202 & \new_[24675]_ ;
  assign \new_[24679]_  = A299 & A298;
  assign \new_[24682]_  = ~A302 & A301;
  assign \new_[24683]_  = \new_[24682]_  & \new_[24679]_ ;
  assign \new_[24684]_  = \new_[24683]_  & \new_[24676]_ ;
  assign \new_[24688]_  = ~A167 & A168;
  assign \new_[24689]_  = A170 & \new_[24688]_ ;
  assign \new_[24692]_  = A199 & A166;
  assign \new_[24695]_  = ~A201 & A200;
  assign \new_[24696]_  = \new_[24695]_  & \new_[24692]_ ;
  assign \new_[24697]_  = \new_[24696]_  & \new_[24689]_ ;
  assign \new_[24701]_  = A234 & A233;
  assign \new_[24702]_  = ~A202 & \new_[24701]_ ;
  assign \new_[24705]_  = ~A299 & A298;
  assign \new_[24708]_  = A302 & ~A301;
  assign \new_[24709]_  = \new_[24708]_  & \new_[24705]_ ;
  assign \new_[24710]_  = \new_[24709]_  & \new_[24702]_ ;
  assign \new_[24714]_  = ~A167 & A168;
  assign \new_[24715]_  = A170 & \new_[24714]_ ;
  assign \new_[24718]_  = A199 & A166;
  assign \new_[24721]_  = ~A201 & A200;
  assign \new_[24722]_  = \new_[24721]_  & \new_[24718]_ ;
  assign \new_[24723]_  = \new_[24722]_  & \new_[24715]_ ;
  assign \new_[24727]_  = A234 & A233;
  assign \new_[24728]_  = ~A202 & \new_[24727]_ ;
  assign \new_[24731]_  = A299 & ~A298;
  assign \new_[24734]_  = A302 & ~A301;
  assign \new_[24735]_  = \new_[24734]_  & \new_[24731]_ ;
  assign \new_[24736]_  = \new_[24735]_  & \new_[24728]_ ;
  assign \new_[24740]_  = ~A167 & A168;
  assign \new_[24741]_  = A170 & \new_[24740]_ ;
  assign \new_[24744]_  = A199 & A166;
  assign \new_[24747]_  = ~A201 & A200;
  assign \new_[24748]_  = \new_[24747]_  & \new_[24744]_ ;
  assign \new_[24749]_  = \new_[24748]_  & \new_[24741]_ ;
  assign \new_[24753]_  = A234 & A233;
  assign \new_[24754]_  = ~A202 & \new_[24753]_ ;
  assign \new_[24757]_  = ~A299 & ~A298;
  assign \new_[24760]_  = ~A302 & A301;
  assign \new_[24761]_  = \new_[24760]_  & \new_[24757]_ ;
  assign \new_[24762]_  = \new_[24761]_  & \new_[24754]_ ;
  assign \new_[24766]_  = ~A167 & A168;
  assign \new_[24767]_  = A170 & \new_[24766]_ ;
  assign \new_[24770]_  = A199 & A166;
  assign \new_[24773]_  = ~A201 & A200;
  assign \new_[24774]_  = \new_[24773]_  & \new_[24770]_ ;
  assign \new_[24775]_  = \new_[24774]_  & \new_[24767]_ ;
  assign \new_[24779]_  = A234 & A233;
  assign \new_[24780]_  = ~A202 & \new_[24779]_ ;
  assign \new_[24783]_  = A266 & A265;
  assign \new_[24786]_  = ~A269 & A268;
  assign \new_[24787]_  = \new_[24786]_  & \new_[24783]_ ;
  assign \new_[24788]_  = \new_[24787]_  & \new_[24780]_ ;
  assign \new_[24792]_  = ~A167 & A168;
  assign \new_[24793]_  = A170 & \new_[24792]_ ;
  assign \new_[24796]_  = A199 & A166;
  assign \new_[24799]_  = ~A201 & A200;
  assign \new_[24800]_  = \new_[24799]_  & \new_[24796]_ ;
  assign \new_[24801]_  = \new_[24800]_  & \new_[24793]_ ;
  assign \new_[24805]_  = A234 & A233;
  assign \new_[24806]_  = ~A202 & \new_[24805]_ ;
  assign \new_[24809]_  = A266 & ~A265;
  assign \new_[24812]_  = A269 & ~A268;
  assign \new_[24813]_  = \new_[24812]_  & \new_[24809]_ ;
  assign \new_[24814]_  = \new_[24813]_  & \new_[24806]_ ;
  assign \new_[24818]_  = ~A167 & A168;
  assign \new_[24819]_  = A170 & \new_[24818]_ ;
  assign \new_[24822]_  = A199 & A166;
  assign \new_[24825]_  = ~A201 & A200;
  assign \new_[24826]_  = \new_[24825]_  & \new_[24822]_ ;
  assign \new_[24827]_  = \new_[24826]_  & \new_[24819]_ ;
  assign \new_[24831]_  = A234 & A233;
  assign \new_[24832]_  = ~A202 & \new_[24831]_ ;
  assign \new_[24835]_  = ~A266 & A265;
  assign \new_[24838]_  = A269 & ~A268;
  assign \new_[24839]_  = \new_[24838]_  & \new_[24835]_ ;
  assign \new_[24840]_  = \new_[24839]_  & \new_[24832]_ ;
  assign \new_[24844]_  = ~A167 & A168;
  assign \new_[24845]_  = A170 & \new_[24844]_ ;
  assign \new_[24848]_  = A199 & A166;
  assign \new_[24851]_  = ~A201 & A200;
  assign \new_[24852]_  = \new_[24851]_  & \new_[24848]_ ;
  assign \new_[24853]_  = \new_[24852]_  & \new_[24845]_ ;
  assign \new_[24857]_  = A234 & A233;
  assign \new_[24858]_  = ~A202 & \new_[24857]_ ;
  assign \new_[24861]_  = ~A266 & ~A265;
  assign \new_[24864]_  = ~A269 & A268;
  assign \new_[24865]_  = \new_[24864]_  & \new_[24861]_ ;
  assign \new_[24866]_  = \new_[24865]_  & \new_[24858]_ ;
  assign \new_[24870]_  = ~A167 & A168;
  assign \new_[24871]_  = A170 & \new_[24870]_ ;
  assign \new_[24874]_  = A199 & A166;
  assign \new_[24877]_  = ~A201 & A200;
  assign \new_[24878]_  = \new_[24877]_  & \new_[24874]_ ;
  assign \new_[24879]_  = \new_[24878]_  & \new_[24871]_ ;
  assign \new_[24883]_  = A233 & A232;
  assign \new_[24884]_  = ~A202 & \new_[24883]_ ;
  assign \new_[24887]_  = ~A236 & A235;
  assign \new_[24890]_  = A300 & A299;
  assign \new_[24891]_  = \new_[24890]_  & \new_[24887]_ ;
  assign \new_[24892]_  = \new_[24891]_  & \new_[24884]_ ;
  assign \new_[24896]_  = ~A167 & A168;
  assign \new_[24897]_  = A170 & \new_[24896]_ ;
  assign \new_[24900]_  = A199 & A166;
  assign \new_[24903]_  = ~A201 & A200;
  assign \new_[24904]_  = \new_[24903]_  & \new_[24900]_ ;
  assign \new_[24905]_  = \new_[24904]_  & \new_[24897]_ ;
  assign \new_[24909]_  = A233 & A232;
  assign \new_[24910]_  = ~A202 & \new_[24909]_ ;
  assign \new_[24913]_  = ~A236 & A235;
  assign \new_[24916]_  = A300 & A298;
  assign \new_[24917]_  = \new_[24916]_  & \new_[24913]_ ;
  assign \new_[24918]_  = \new_[24917]_  & \new_[24910]_ ;
  assign \new_[24922]_  = ~A167 & A168;
  assign \new_[24923]_  = A170 & \new_[24922]_ ;
  assign \new_[24926]_  = A199 & A166;
  assign \new_[24929]_  = ~A201 & A200;
  assign \new_[24930]_  = \new_[24929]_  & \new_[24926]_ ;
  assign \new_[24931]_  = \new_[24930]_  & \new_[24923]_ ;
  assign \new_[24935]_  = A233 & A232;
  assign \new_[24936]_  = ~A202 & \new_[24935]_ ;
  assign \new_[24939]_  = ~A236 & A235;
  assign \new_[24942]_  = A267 & A265;
  assign \new_[24943]_  = \new_[24942]_  & \new_[24939]_ ;
  assign \new_[24944]_  = \new_[24943]_  & \new_[24936]_ ;
  assign \new_[24948]_  = ~A167 & A168;
  assign \new_[24949]_  = A170 & \new_[24948]_ ;
  assign \new_[24952]_  = A199 & A166;
  assign \new_[24955]_  = ~A201 & A200;
  assign \new_[24956]_  = \new_[24955]_  & \new_[24952]_ ;
  assign \new_[24957]_  = \new_[24956]_  & \new_[24949]_ ;
  assign \new_[24961]_  = A233 & A232;
  assign \new_[24962]_  = ~A202 & \new_[24961]_ ;
  assign \new_[24965]_  = ~A236 & A235;
  assign \new_[24968]_  = A267 & A266;
  assign \new_[24969]_  = \new_[24968]_  & \new_[24965]_ ;
  assign \new_[24970]_  = \new_[24969]_  & \new_[24962]_ ;
  assign \new_[24974]_  = ~A167 & A168;
  assign \new_[24975]_  = A170 & \new_[24974]_ ;
  assign \new_[24978]_  = A199 & A166;
  assign \new_[24981]_  = ~A201 & A200;
  assign \new_[24982]_  = \new_[24981]_  & \new_[24978]_ ;
  assign \new_[24983]_  = \new_[24982]_  & \new_[24975]_ ;
  assign \new_[24987]_  = A233 & ~A232;
  assign \new_[24988]_  = ~A202 & \new_[24987]_ ;
  assign \new_[24991]_  = A236 & ~A235;
  assign \new_[24994]_  = A300 & A299;
  assign \new_[24995]_  = \new_[24994]_  & \new_[24991]_ ;
  assign \new_[24996]_  = \new_[24995]_  & \new_[24988]_ ;
  assign \new_[25000]_  = ~A167 & A168;
  assign \new_[25001]_  = A170 & \new_[25000]_ ;
  assign \new_[25004]_  = A199 & A166;
  assign \new_[25007]_  = ~A201 & A200;
  assign \new_[25008]_  = \new_[25007]_  & \new_[25004]_ ;
  assign \new_[25009]_  = \new_[25008]_  & \new_[25001]_ ;
  assign \new_[25013]_  = A233 & ~A232;
  assign \new_[25014]_  = ~A202 & \new_[25013]_ ;
  assign \new_[25017]_  = A236 & ~A235;
  assign \new_[25020]_  = A300 & A298;
  assign \new_[25021]_  = \new_[25020]_  & \new_[25017]_ ;
  assign \new_[25022]_  = \new_[25021]_  & \new_[25014]_ ;
  assign \new_[25026]_  = ~A167 & A168;
  assign \new_[25027]_  = A170 & \new_[25026]_ ;
  assign \new_[25030]_  = A199 & A166;
  assign \new_[25033]_  = ~A201 & A200;
  assign \new_[25034]_  = \new_[25033]_  & \new_[25030]_ ;
  assign \new_[25035]_  = \new_[25034]_  & \new_[25027]_ ;
  assign \new_[25039]_  = A233 & ~A232;
  assign \new_[25040]_  = ~A202 & \new_[25039]_ ;
  assign \new_[25043]_  = A236 & ~A235;
  assign \new_[25046]_  = A267 & A265;
  assign \new_[25047]_  = \new_[25046]_  & \new_[25043]_ ;
  assign \new_[25048]_  = \new_[25047]_  & \new_[25040]_ ;
  assign \new_[25052]_  = ~A167 & A168;
  assign \new_[25053]_  = A170 & \new_[25052]_ ;
  assign \new_[25056]_  = A199 & A166;
  assign \new_[25059]_  = ~A201 & A200;
  assign \new_[25060]_  = \new_[25059]_  & \new_[25056]_ ;
  assign \new_[25061]_  = \new_[25060]_  & \new_[25053]_ ;
  assign \new_[25065]_  = A233 & ~A232;
  assign \new_[25066]_  = ~A202 & \new_[25065]_ ;
  assign \new_[25069]_  = A236 & ~A235;
  assign \new_[25072]_  = A267 & A266;
  assign \new_[25073]_  = \new_[25072]_  & \new_[25069]_ ;
  assign \new_[25074]_  = \new_[25073]_  & \new_[25066]_ ;
  assign \new_[25078]_  = ~A167 & A168;
  assign \new_[25079]_  = A170 & \new_[25078]_ ;
  assign \new_[25082]_  = A199 & A166;
  assign \new_[25085]_  = ~A201 & A200;
  assign \new_[25086]_  = \new_[25085]_  & \new_[25082]_ ;
  assign \new_[25087]_  = \new_[25086]_  & \new_[25079]_ ;
  assign \new_[25091]_  = ~A233 & A232;
  assign \new_[25092]_  = ~A202 & \new_[25091]_ ;
  assign \new_[25095]_  = A236 & ~A235;
  assign \new_[25098]_  = A300 & A299;
  assign \new_[25099]_  = \new_[25098]_  & \new_[25095]_ ;
  assign \new_[25100]_  = \new_[25099]_  & \new_[25092]_ ;
  assign \new_[25104]_  = ~A167 & A168;
  assign \new_[25105]_  = A170 & \new_[25104]_ ;
  assign \new_[25108]_  = A199 & A166;
  assign \new_[25111]_  = ~A201 & A200;
  assign \new_[25112]_  = \new_[25111]_  & \new_[25108]_ ;
  assign \new_[25113]_  = \new_[25112]_  & \new_[25105]_ ;
  assign \new_[25117]_  = ~A233 & A232;
  assign \new_[25118]_  = ~A202 & \new_[25117]_ ;
  assign \new_[25121]_  = A236 & ~A235;
  assign \new_[25124]_  = A300 & A298;
  assign \new_[25125]_  = \new_[25124]_  & \new_[25121]_ ;
  assign \new_[25126]_  = \new_[25125]_  & \new_[25118]_ ;
  assign \new_[25130]_  = ~A167 & A168;
  assign \new_[25131]_  = A170 & \new_[25130]_ ;
  assign \new_[25134]_  = A199 & A166;
  assign \new_[25137]_  = ~A201 & A200;
  assign \new_[25138]_  = \new_[25137]_  & \new_[25134]_ ;
  assign \new_[25139]_  = \new_[25138]_  & \new_[25131]_ ;
  assign \new_[25143]_  = ~A233 & A232;
  assign \new_[25144]_  = ~A202 & \new_[25143]_ ;
  assign \new_[25147]_  = A236 & ~A235;
  assign \new_[25150]_  = A267 & A265;
  assign \new_[25151]_  = \new_[25150]_  & \new_[25147]_ ;
  assign \new_[25152]_  = \new_[25151]_  & \new_[25144]_ ;
  assign \new_[25156]_  = ~A167 & A168;
  assign \new_[25157]_  = A170 & \new_[25156]_ ;
  assign \new_[25160]_  = A199 & A166;
  assign \new_[25163]_  = ~A201 & A200;
  assign \new_[25164]_  = \new_[25163]_  & \new_[25160]_ ;
  assign \new_[25165]_  = \new_[25164]_  & \new_[25157]_ ;
  assign \new_[25169]_  = ~A233 & A232;
  assign \new_[25170]_  = ~A202 & \new_[25169]_ ;
  assign \new_[25173]_  = A236 & ~A235;
  assign \new_[25176]_  = A267 & A266;
  assign \new_[25177]_  = \new_[25176]_  & \new_[25173]_ ;
  assign \new_[25178]_  = \new_[25177]_  & \new_[25170]_ ;
  assign \new_[25182]_  = ~A167 & A168;
  assign \new_[25183]_  = A170 & \new_[25182]_ ;
  assign \new_[25186]_  = A199 & A166;
  assign \new_[25189]_  = ~A201 & A200;
  assign \new_[25190]_  = \new_[25189]_  & \new_[25186]_ ;
  assign \new_[25191]_  = \new_[25190]_  & \new_[25183]_ ;
  assign \new_[25195]_  = ~A233 & ~A232;
  assign \new_[25196]_  = ~A202 & \new_[25195]_ ;
  assign \new_[25199]_  = ~A236 & A235;
  assign \new_[25202]_  = A300 & A299;
  assign \new_[25203]_  = \new_[25202]_  & \new_[25199]_ ;
  assign \new_[25204]_  = \new_[25203]_  & \new_[25196]_ ;
  assign \new_[25208]_  = ~A167 & A168;
  assign \new_[25209]_  = A170 & \new_[25208]_ ;
  assign \new_[25212]_  = A199 & A166;
  assign \new_[25215]_  = ~A201 & A200;
  assign \new_[25216]_  = \new_[25215]_  & \new_[25212]_ ;
  assign \new_[25217]_  = \new_[25216]_  & \new_[25209]_ ;
  assign \new_[25221]_  = ~A233 & ~A232;
  assign \new_[25222]_  = ~A202 & \new_[25221]_ ;
  assign \new_[25225]_  = ~A236 & A235;
  assign \new_[25228]_  = A300 & A298;
  assign \new_[25229]_  = \new_[25228]_  & \new_[25225]_ ;
  assign \new_[25230]_  = \new_[25229]_  & \new_[25222]_ ;
  assign \new_[25234]_  = ~A167 & A168;
  assign \new_[25235]_  = A170 & \new_[25234]_ ;
  assign \new_[25238]_  = A199 & A166;
  assign \new_[25241]_  = ~A201 & A200;
  assign \new_[25242]_  = \new_[25241]_  & \new_[25238]_ ;
  assign \new_[25243]_  = \new_[25242]_  & \new_[25235]_ ;
  assign \new_[25247]_  = ~A233 & ~A232;
  assign \new_[25248]_  = ~A202 & \new_[25247]_ ;
  assign \new_[25251]_  = ~A236 & A235;
  assign \new_[25254]_  = A267 & A265;
  assign \new_[25255]_  = \new_[25254]_  & \new_[25251]_ ;
  assign \new_[25256]_  = \new_[25255]_  & \new_[25248]_ ;
  assign \new_[25260]_  = ~A167 & A168;
  assign \new_[25261]_  = A170 & \new_[25260]_ ;
  assign \new_[25264]_  = A199 & A166;
  assign \new_[25267]_  = ~A201 & A200;
  assign \new_[25268]_  = \new_[25267]_  & \new_[25264]_ ;
  assign \new_[25269]_  = \new_[25268]_  & \new_[25261]_ ;
  assign \new_[25273]_  = ~A233 & ~A232;
  assign \new_[25274]_  = ~A202 & \new_[25273]_ ;
  assign \new_[25277]_  = ~A236 & A235;
  assign \new_[25280]_  = A267 & A266;
  assign \new_[25281]_  = \new_[25280]_  & \new_[25277]_ ;
  assign \new_[25282]_  = \new_[25281]_  & \new_[25274]_ ;
  assign \new_[25286]_  = ~A167 & A168;
  assign \new_[25287]_  = A170 & \new_[25286]_ ;
  assign \new_[25290]_  = A199 & A166;
  assign \new_[25293]_  = ~A201 & A200;
  assign \new_[25294]_  = \new_[25293]_  & \new_[25290]_ ;
  assign \new_[25295]_  = \new_[25294]_  & \new_[25287]_ ;
  assign \new_[25299]_  = A234 & A232;
  assign \new_[25300]_  = A203 & \new_[25299]_ ;
  assign \new_[25303]_  = A299 & A298;
  assign \new_[25306]_  = ~A302 & A301;
  assign \new_[25307]_  = \new_[25306]_  & \new_[25303]_ ;
  assign \new_[25308]_  = \new_[25307]_  & \new_[25300]_ ;
  assign \new_[25312]_  = ~A167 & A168;
  assign \new_[25313]_  = A170 & \new_[25312]_ ;
  assign \new_[25316]_  = A199 & A166;
  assign \new_[25319]_  = ~A201 & A200;
  assign \new_[25320]_  = \new_[25319]_  & \new_[25316]_ ;
  assign \new_[25321]_  = \new_[25320]_  & \new_[25313]_ ;
  assign \new_[25325]_  = A234 & A232;
  assign \new_[25326]_  = A203 & \new_[25325]_ ;
  assign \new_[25329]_  = ~A299 & A298;
  assign \new_[25332]_  = A302 & ~A301;
  assign \new_[25333]_  = \new_[25332]_  & \new_[25329]_ ;
  assign \new_[25334]_  = \new_[25333]_  & \new_[25326]_ ;
  assign \new_[25338]_  = ~A167 & A168;
  assign \new_[25339]_  = A170 & \new_[25338]_ ;
  assign \new_[25342]_  = A199 & A166;
  assign \new_[25345]_  = ~A201 & A200;
  assign \new_[25346]_  = \new_[25345]_  & \new_[25342]_ ;
  assign \new_[25347]_  = \new_[25346]_  & \new_[25339]_ ;
  assign \new_[25351]_  = A234 & A232;
  assign \new_[25352]_  = A203 & \new_[25351]_ ;
  assign \new_[25355]_  = A299 & ~A298;
  assign \new_[25358]_  = A302 & ~A301;
  assign \new_[25359]_  = \new_[25358]_  & \new_[25355]_ ;
  assign \new_[25360]_  = \new_[25359]_  & \new_[25352]_ ;
  assign \new_[25364]_  = ~A167 & A168;
  assign \new_[25365]_  = A170 & \new_[25364]_ ;
  assign \new_[25368]_  = A199 & A166;
  assign \new_[25371]_  = ~A201 & A200;
  assign \new_[25372]_  = \new_[25371]_  & \new_[25368]_ ;
  assign \new_[25373]_  = \new_[25372]_  & \new_[25365]_ ;
  assign \new_[25377]_  = A234 & A232;
  assign \new_[25378]_  = A203 & \new_[25377]_ ;
  assign \new_[25381]_  = ~A299 & ~A298;
  assign \new_[25384]_  = ~A302 & A301;
  assign \new_[25385]_  = \new_[25384]_  & \new_[25381]_ ;
  assign \new_[25386]_  = \new_[25385]_  & \new_[25378]_ ;
  assign \new_[25390]_  = ~A167 & A168;
  assign \new_[25391]_  = A170 & \new_[25390]_ ;
  assign \new_[25394]_  = A199 & A166;
  assign \new_[25397]_  = ~A201 & A200;
  assign \new_[25398]_  = \new_[25397]_  & \new_[25394]_ ;
  assign \new_[25399]_  = \new_[25398]_  & \new_[25391]_ ;
  assign \new_[25403]_  = A234 & A232;
  assign \new_[25404]_  = A203 & \new_[25403]_ ;
  assign \new_[25407]_  = A266 & A265;
  assign \new_[25410]_  = ~A269 & A268;
  assign \new_[25411]_  = \new_[25410]_  & \new_[25407]_ ;
  assign \new_[25412]_  = \new_[25411]_  & \new_[25404]_ ;
  assign \new_[25416]_  = ~A167 & A168;
  assign \new_[25417]_  = A170 & \new_[25416]_ ;
  assign \new_[25420]_  = A199 & A166;
  assign \new_[25423]_  = ~A201 & A200;
  assign \new_[25424]_  = \new_[25423]_  & \new_[25420]_ ;
  assign \new_[25425]_  = \new_[25424]_  & \new_[25417]_ ;
  assign \new_[25429]_  = A234 & A232;
  assign \new_[25430]_  = A203 & \new_[25429]_ ;
  assign \new_[25433]_  = A266 & ~A265;
  assign \new_[25436]_  = A269 & ~A268;
  assign \new_[25437]_  = \new_[25436]_  & \new_[25433]_ ;
  assign \new_[25438]_  = \new_[25437]_  & \new_[25430]_ ;
  assign \new_[25442]_  = ~A167 & A168;
  assign \new_[25443]_  = A170 & \new_[25442]_ ;
  assign \new_[25446]_  = A199 & A166;
  assign \new_[25449]_  = ~A201 & A200;
  assign \new_[25450]_  = \new_[25449]_  & \new_[25446]_ ;
  assign \new_[25451]_  = \new_[25450]_  & \new_[25443]_ ;
  assign \new_[25455]_  = A234 & A232;
  assign \new_[25456]_  = A203 & \new_[25455]_ ;
  assign \new_[25459]_  = ~A266 & A265;
  assign \new_[25462]_  = A269 & ~A268;
  assign \new_[25463]_  = \new_[25462]_  & \new_[25459]_ ;
  assign \new_[25464]_  = \new_[25463]_  & \new_[25456]_ ;
  assign \new_[25468]_  = ~A167 & A168;
  assign \new_[25469]_  = A170 & \new_[25468]_ ;
  assign \new_[25472]_  = A199 & A166;
  assign \new_[25475]_  = ~A201 & A200;
  assign \new_[25476]_  = \new_[25475]_  & \new_[25472]_ ;
  assign \new_[25477]_  = \new_[25476]_  & \new_[25469]_ ;
  assign \new_[25481]_  = A234 & A232;
  assign \new_[25482]_  = A203 & \new_[25481]_ ;
  assign \new_[25485]_  = ~A266 & ~A265;
  assign \new_[25488]_  = ~A269 & A268;
  assign \new_[25489]_  = \new_[25488]_  & \new_[25485]_ ;
  assign \new_[25490]_  = \new_[25489]_  & \new_[25482]_ ;
  assign \new_[25494]_  = ~A167 & A168;
  assign \new_[25495]_  = A170 & \new_[25494]_ ;
  assign \new_[25498]_  = A199 & A166;
  assign \new_[25501]_  = ~A201 & A200;
  assign \new_[25502]_  = \new_[25501]_  & \new_[25498]_ ;
  assign \new_[25503]_  = \new_[25502]_  & \new_[25495]_ ;
  assign \new_[25507]_  = A234 & A233;
  assign \new_[25508]_  = A203 & \new_[25507]_ ;
  assign \new_[25511]_  = A299 & A298;
  assign \new_[25514]_  = ~A302 & A301;
  assign \new_[25515]_  = \new_[25514]_  & \new_[25511]_ ;
  assign \new_[25516]_  = \new_[25515]_  & \new_[25508]_ ;
  assign \new_[25520]_  = ~A167 & A168;
  assign \new_[25521]_  = A170 & \new_[25520]_ ;
  assign \new_[25524]_  = A199 & A166;
  assign \new_[25527]_  = ~A201 & A200;
  assign \new_[25528]_  = \new_[25527]_  & \new_[25524]_ ;
  assign \new_[25529]_  = \new_[25528]_  & \new_[25521]_ ;
  assign \new_[25533]_  = A234 & A233;
  assign \new_[25534]_  = A203 & \new_[25533]_ ;
  assign \new_[25537]_  = ~A299 & A298;
  assign \new_[25540]_  = A302 & ~A301;
  assign \new_[25541]_  = \new_[25540]_  & \new_[25537]_ ;
  assign \new_[25542]_  = \new_[25541]_  & \new_[25534]_ ;
  assign \new_[25546]_  = ~A167 & A168;
  assign \new_[25547]_  = A170 & \new_[25546]_ ;
  assign \new_[25550]_  = A199 & A166;
  assign \new_[25553]_  = ~A201 & A200;
  assign \new_[25554]_  = \new_[25553]_  & \new_[25550]_ ;
  assign \new_[25555]_  = \new_[25554]_  & \new_[25547]_ ;
  assign \new_[25559]_  = A234 & A233;
  assign \new_[25560]_  = A203 & \new_[25559]_ ;
  assign \new_[25563]_  = A299 & ~A298;
  assign \new_[25566]_  = A302 & ~A301;
  assign \new_[25567]_  = \new_[25566]_  & \new_[25563]_ ;
  assign \new_[25568]_  = \new_[25567]_  & \new_[25560]_ ;
  assign \new_[25572]_  = ~A167 & A168;
  assign \new_[25573]_  = A170 & \new_[25572]_ ;
  assign \new_[25576]_  = A199 & A166;
  assign \new_[25579]_  = ~A201 & A200;
  assign \new_[25580]_  = \new_[25579]_  & \new_[25576]_ ;
  assign \new_[25581]_  = \new_[25580]_  & \new_[25573]_ ;
  assign \new_[25585]_  = A234 & A233;
  assign \new_[25586]_  = A203 & \new_[25585]_ ;
  assign \new_[25589]_  = ~A299 & ~A298;
  assign \new_[25592]_  = ~A302 & A301;
  assign \new_[25593]_  = \new_[25592]_  & \new_[25589]_ ;
  assign \new_[25594]_  = \new_[25593]_  & \new_[25586]_ ;
  assign \new_[25598]_  = ~A167 & A168;
  assign \new_[25599]_  = A170 & \new_[25598]_ ;
  assign \new_[25602]_  = A199 & A166;
  assign \new_[25605]_  = ~A201 & A200;
  assign \new_[25606]_  = \new_[25605]_  & \new_[25602]_ ;
  assign \new_[25607]_  = \new_[25606]_  & \new_[25599]_ ;
  assign \new_[25611]_  = A234 & A233;
  assign \new_[25612]_  = A203 & \new_[25611]_ ;
  assign \new_[25615]_  = A266 & A265;
  assign \new_[25618]_  = ~A269 & A268;
  assign \new_[25619]_  = \new_[25618]_  & \new_[25615]_ ;
  assign \new_[25620]_  = \new_[25619]_  & \new_[25612]_ ;
  assign \new_[25624]_  = ~A167 & A168;
  assign \new_[25625]_  = A170 & \new_[25624]_ ;
  assign \new_[25628]_  = A199 & A166;
  assign \new_[25631]_  = ~A201 & A200;
  assign \new_[25632]_  = \new_[25631]_  & \new_[25628]_ ;
  assign \new_[25633]_  = \new_[25632]_  & \new_[25625]_ ;
  assign \new_[25637]_  = A234 & A233;
  assign \new_[25638]_  = A203 & \new_[25637]_ ;
  assign \new_[25641]_  = A266 & ~A265;
  assign \new_[25644]_  = A269 & ~A268;
  assign \new_[25645]_  = \new_[25644]_  & \new_[25641]_ ;
  assign \new_[25646]_  = \new_[25645]_  & \new_[25638]_ ;
  assign \new_[25650]_  = ~A167 & A168;
  assign \new_[25651]_  = A170 & \new_[25650]_ ;
  assign \new_[25654]_  = A199 & A166;
  assign \new_[25657]_  = ~A201 & A200;
  assign \new_[25658]_  = \new_[25657]_  & \new_[25654]_ ;
  assign \new_[25659]_  = \new_[25658]_  & \new_[25651]_ ;
  assign \new_[25663]_  = A234 & A233;
  assign \new_[25664]_  = A203 & \new_[25663]_ ;
  assign \new_[25667]_  = ~A266 & A265;
  assign \new_[25670]_  = A269 & ~A268;
  assign \new_[25671]_  = \new_[25670]_  & \new_[25667]_ ;
  assign \new_[25672]_  = \new_[25671]_  & \new_[25664]_ ;
  assign \new_[25676]_  = ~A167 & A168;
  assign \new_[25677]_  = A170 & \new_[25676]_ ;
  assign \new_[25680]_  = A199 & A166;
  assign \new_[25683]_  = ~A201 & A200;
  assign \new_[25684]_  = \new_[25683]_  & \new_[25680]_ ;
  assign \new_[25685]_  = \new_[25684]_  & \new_[25677]_ ;
  assign \new_[25689]_  = A234 & A233;
  assign \new_[25690]_  = A203 & \new_[25689]_ ;
  assign \new_[25693]_  = ~A266 & ~A265;
  assign \new_[25696]_  = ~A269 & A268;
  assign \new_[25697]_  = \new_[25696]_  & \new_[25693]_ ;
  assign \new_[25698]_  = \new_[25697]_  & \new_[25690]_ ;
  assign \new_[25702]_  = ~A167 & A168;
  assign \new_[25703]_  = A170 & \new_[25702]_ ;
  assign \new_[25706]_  = A199 & A166;
  assign \new_[25709]_  = ~A201 & A200;
  assign \new_[25710]_  = \new_[25709]_  & \new_[25706]_ ;
  assign \new_[25711]_  = \new_[25710]_  & \new_[25703]_ ;
  assign \new_[25715]_  = A233 & A232;
  assign \new_[25716]_  = A203 & \new_[25715]_ ;
  assign \new_[25719]_  = ~A236 & A235;
  assign \new_[25722]_  = A300 & A299;
  assign \new_[25723]_  = \new_[25722]_  & \new_[25719]_ ;
  assign \new_[25724]_  = \new_[25723]_  & \new_[25716]_ ;
  assign \new_[25728]_  = ~A167 & A168;
  assign \new_[25729]_  = A170 & \new_[25728]_ ;
  assign \new_[25732]_  = A199 & A166;
  assign \new_[25735]_  = ~A201 & A200;
  assign \new_[25736]_  = \new_[25735]_  & \new_[25732]_ ;
  assign \new_[25737]_  = \new_[25736]_  & \new_[25729]_ ;
  assign \new_[25741]_  = A233 & A232;
  assign \new_[25742]_  = A203 & \new_[25741]_ ;
  assign \new_[25745]_  = ~A236 & A235;
  assign \new_[25748]_  = A300 & A298;
  assign \new_[25749]_  = \new_[25748]_  & \new_[25745]_ ;
  assign \new_[25750]_  = \new_[25749]_  & \new_[25742]_ ;
  assign \new_[25754]_  = ~A167 & A168;
  assign \new_[25755]_  = A170 & \new_[25754]_ ;
  assign \new_[25758]_  = A199 & A166;
  assign \new_[25761]_  = ~A201 & A200;
  assign \new_[25762]_  = \new_[25761]_  & \new_[25758]_ ;
  assign \new_[25763]_  = \new_[25762]_  & \new_[25755]_ ;
  assign \new_[25767]_  = A233 & A232;
  assign \new_[25768]_  = A203 & \new_[25767]_ ;
  assign \new_[25771]_  = ~A236 & A235;
  assign \new_[25774]_  = A267 & A265;
  assign \new_[25775]_  = \new_[25774]_  & \new_[25771]_ ;
  assign \new_[25776]_  = \new_[25775]_  & \new_[25768]_ ;
  assign \new_[25780]_  = ~A167 & A168;
  assign \new_[25781]_  = A170 & \new_[25780]_ ;
  assign \new_[25784]_  = A199 & A166;
  assign \new_[25787]_  = ~A201 & A200;
  assign \new_[25788]_  = \new_[25787]_  & \new_[25784]_ ;
  assign \new_[25789]_  = \new_[25788]_  & \new_[25781]_ ;
  assign \new_[25793]_  = A233 & A232;
  assign \new_[25794]_  = A203 & \new_[25793]_ ;
  assign \new_[25797]_  = ~A236 & A235;
  assign \new_[25800]_  = A267 & A266;
  assign \new_[25801]_  = \new_[25800]_  & \new_[25797]_ ;
  assign \new_[25802]_  = \new_[25801]_  & \new_[25794]_ ;
  assign \new_[25806]_  = ~A167 & A168;
  assign \new_[25807]_  = A170 & \new_[25806]_ ;
  assign \new_[25810]_  = A199 & A166;
  assign \new_[25813]_  = ~A201 & A200;
  assign \new_[25814]_  = \new_[25813]_  & \new_[25810]_ ;
  assign \new_[25815]_  = \new_[25814]_  & \new_[25807]_ ;
  assign \new_[25819]_  = A233 & ~A232;
  assign \new_[25820]_  = A203 & \new_[25819]_ ;
  assign \new_[25823]_  = A236 & ~A235;
  assign \new_[25826]_  = A300 & A299;
  assign \new_[25827]_  = \new_[25826]_  & \new_[25823]_ ;
  assign \new_[25828]_  = \new_[25827]_  & \new_[25820]_ ;
  assign \new_[25832]_  = ~A167 & A168;
  assign \new_[25833]_  = A170 & \new_[25832]_ ;
  assign \new_[25836]_  = A199 & A166;
  assign \new_[25839]_  = ~A201 & A200;
  assign \new_[25840]_  = \new_[25839]_  & \new_[25836]_ ;
  assign \new_[25841]_  = \new_[25840]_  & \new_[25833]_ ;
  assign \new_[25845]_  = A233 & ~A232;
  assign \new_[25846]_  = A203 & \new_[25845]_ ;
  assign \new_[25849]_  = A236 & ~A235;
  assign \new_[25852]_  = A300 & A298;
  assign \new_[25853]_  = \new_[25852]_  & \new_[25849]_ ;
  assign \new_[25854]_  = \new_[25853]_  & \new_[25846]_ ;
  assign \new_[25858]_  = ~A167 & A168;
  assign \new_[25859]_  = A170 & \new_[25858]_ ;
  assign \new_[25862]_  = A199 & A166;
  assign \new_[25865]_  = ~A201 & A200;
  assign \new_[25866]_  = \new_[25865]_  & \new_[25862]_ ;
  assign \new_[25867]_  = \new_[25866]_  & \new_[25859]_ ;
  assign \new_[25871]_  = A233 & ~A232;
  assign \new_[25872]_  = A203 & \new_[25871]_ ;
  assign \new_[25875]_  = A236 & ~A235;
  assign \new_[25878]_  = A267 & A265;
  assign \new_[25879]_  = \new_[25878]_  & \new_[25875]_ ;
  assign \new_[25880]_  = \new_[25879]_  & \new_[25872]_ ;
  assign \new_[25884]_  = ~A167 & A168;
  assign \new_[25885]_  = A170 & \new_[25884]_ ;
  assign \new_[25888]_  = A199 & A166;
  assign \new_[25891]_  = ~A201 & A200;
  assign \new_[25892]_  = \new_[25891]_  & \new_[25888]_ ;
  assign \new_[25893]_  = \new_[25892]_  & \new_[25885]_ ;
  assign \new_[25897]_  = A233 & ~A232;
  assign \new_[25898]_  = A203 & \new_[25897]_ ;
  assign \new_[25901]_  = A236 & ~A235;
  assign \new_[25904]_  = A267 & A266;
  assign \new_[25905]_  = \new_[25904]_  & \new_[25901]_ ;
  assign \new_[25906]_  = \new_[25905]_  & \new_[25898]_ ;
  assign \new_[25910]_  = ~A167 & A168;
  assign \new_[25911]_  = A170 & \new_[25910]_ ;
  assign \new_[25914]_  = A199 & A166;
  assign \new_[25917]_  = ~A201 & A200;
  assign \new_[25918]_  = \new_[25917]_  & \new_[25914]_ ;
  assign \new_[25919]_  = \new_[25918]_  & \new_[25911]_ ;
  assign \new_[25923]_  = ~A233 & A232;
  assign \new_[25924]_  = A203 & \new_[25923]_ ;
  assign \new_[25927]_  = A236 & ~A235;
  assign \new_[25930]_  = A300 & A299;
  assign \new_[25931]_  = \new_[25930]_  & \new_[25927]_ ;
  assign \new_[25932]_  = \new_[25931]_  & \new_[25924]_ ;
  assign \new_[25936]_  = ~A167 & A168;
  assign \new_[25937]_  = A170 & \new_[25936]_ ;
  assign \new_[25940]_  = A199 & A166;
  assign \new_[25943]_  = ~A201 & A200;
  assign \new_[25944]_  = \new_[25943]_  & \new_[25940]_ ;
  assign \new_[25945]_  = \new_[25944]_  & \new_[25937]_ ;
  assign \new_[25949]_  = ~A233 & A232;
  assign \new_[25950]_  = A203 & \new_[25949]_ ;
  assign \new_[25953]_  = A236 & ~A235;
  assign \new_[25956]_  = A300 & A298;
  assign \new_[25957]_  = \new_[25956]_  & \new_[25953]_ ;
  assign \new_[25958]_  = \new_[25957]_  & \new_[25950]_ ;
  assign \new_[25962]_  = ~A167 & A168;
  assign \new_[25963]_  = A170 & \new_[25962]_ ;
  assign \new_[25966]_  = A199 & A166;
  assign \new_[25969]_  = ~A201 & A200;
  assign \new_[25970]_  = \new_[25969]_  & \new_[25966]_ ;
  assign \new_[25971]_  = \new_[25970]_  & \new_[25963]_ ;
  assign \new_[25975]_  = ~A233 & A232;
  assign \new_[25976]_  = A203 & \new_[25975]_ ;
  assign \new_[25979]_  = A236 & ~A235;
  assign \new_[25982]_  = A267 & A265;
  assign \new_[25983]_  = \new_[25982]_  & \new_[25979]_ ;
  assign \new_[25984]_  = \new_[25983]_  & \new_[25976]_ ;
  assign \new_[25988]_  = ~A167 & A168;
  assign \new_[25989]_  = A170 & \new_[25988]_ ;
  assign \new_[25992]_  = A199 & A166;
  assign \new_[25995]_  = ~A201 & A200;
  assign \new_[25996]_  = \new_[25995]_  & \new_[25992]_ ;
  assign \new_[25997]_  = \new_[25996]_  & \new_[25989]_ ;
  assign \new_[26001]_  = ~A233 & A232;
  assign \new_[26002]_  = A203 & \new_[26001]_ ;
  assign \new_[26005]_  = A236 & ~A235;
  assign \new_[26008]_  = A267 & A266;
  assign \new_[26009]_  = \new_[26008]_  & \new_[26005]_ ;
  assign \new_[26010]_  = \new_[26009]_  & \new_[26002]_ ;
  assign \new_[26014]_  = ~A167 & A168;
  assign \new_[26015]_  = A170 & \new_[26014]_ ;
  assign \new_[26018]_  = A199 & A166;
  assign \new_[26021]_  = ~A201 & A200;
  assign \new_[26022]_  = \new_[26021]_  & \new_[26018]_ ;
  assign \new_[26023]_  = \new_[26022]_  & \new_[26015]_ ;
  assign \new_[26027]_  = ~A233 & ~A232;
  assign \new_[26028]_  = A203 & \new_[26027]_ ;
  assign \new_[26031]_  = ~A236 & A235;
  assign \new_[26034]_  = A300 & A299;
  assign \new_[26035]_  = \new_[26034]_  & \new_[26031]_ ;
  assign \new_[26036]_  = \new_[26035]_  & \new_[26028]_ ;
  assign \new_[26040]_  = ~A167 & A168;
  assign \new_[26041]_  = A170 & \new_[26040]_ ;
  assign \new_[26044]_  = A199 & A166;
  assign \new_[26047]_  = ~A201 & A200;
  assign \new_[26048]_  = \new_[26047]_  & \new_[26044]_ ;
  assign \new_[26049]_  = \new_[26048]_  & \new_[26041]_ ;
  assign \new_[26053]_  = ~A233 & ~A232;
  assign \new_[26054]_  = A203 & \new_[26053]_ ;
  assign \new_[26057]_  = ~A236 & A235;
  assign \new_[26060]_  = A300 & A298;
  assign \new_[26061]_  = \new_[26060]_  & \new_[26057]_ ;
  assign \new_[26062]_  = \new_[26061]_  & \new_[26054]_ ;
  assign \new_[26066]_  = ~A167 & A168;
  assign \new_[26067]_  = A170 & \new_[26066]_ ;
  assign \new_[26070]_  = A199 & A166;
  assign \new_[26073]_  = ~A201 & A200;
  assign \new_[26074]_  = \new_[26073]_  & \new_[26070]_ ;
  assign \new_[26075]_  = \new_[26074]_  & \new_[26067]_ ;
  assign \new_[26079]_  = ~A233 & ~A232;
  assign \new_[26080]_  = A203 & \new_[26079]_ ;
  assign \new_[26083]_  = ~A236 & A235;
  assign \new_[26086]_  = A267 & A265;
  assign \new_[26087]_  = \new_[26086]_  & \new_[26083]_ ;
  assign \new_[26088]_  = \new_[26087]_  & \new_[26080]_ ;
  assign \new_[26092]_  = ~A167 & A168;
  assign \new_[26093]_  = A170 & \new_[26092]_ ;
  assign \new_[26096]_  = A199 & A166;
  assign \new_[26099]_  = ~A201 & A200;
  assign \new_[26100]_  = \new_[26099]_  & \new_[26096]_ ;
  assign \new_[26101]_  = \new_[26100]_  & \new_[26093]_ ;
  assign \new_[26105]_  = ~A233 & ~A232;
  assign \new_[26106]_  = A203 & \new_[26105]_ ;
  assign \new_[26109]_  = ~A236 & A235;
  assign \new_[26112]_  = A267 & A266;
  assign \new_[26113]_  = \new_[26112]_  & \new_[26109]_ ;
  assign \new_[26114]_  = \new_[26113]_  & \new_[26106]_ ;
  assign \new_[26118]_  = ~A167 & A168;
  assign \new_[26119]_  = A170 & \new_[26118]_ ;
  assign \new_[26122]_  = ~A199 & A166;
  assign \new_[26125]_  = ~A201 & A200;
  assign \new_[26126]_  = \new_[26125]_  & \new_[26122]_ ;
  assign \new_[26127]_  = \new_[26126]_  & \new_[26119]_ ;
  assign \new_[26131]_  = A234 & A232;
  assign \new_[26132]_  = A202 & \new_[26131]_ ;
  assign \new_[26135]_  = A299 & A298;
  assign \new_[26138]_  = ~A302 & A301;
  assign \new_[26139]_  = \new_[26138]_  & \new_[26135]_ ;
  assign \new_[26140]_  = \new_[26139]_  & \new_[26132]_ ;
  assign \new_[26144]_  = ~A167 & A168;
  assign \new_[26145]_  = A170 & \new_[26144]_ ;
  assign \new_[26148]_  = ~A199 & A166;
  assign \new_[26151]_  = ~A201 & A200;
  assign \new_[26152]_  = \new_[26151]_  & \new_[26148]_ ;
  assign \new_[26153]_  = \new_[26152]_  & \new_[26145]_ ;
  assign \new_[26157]_  = A234 & A232;
  assign \new_[26158]_  = A202 & \new_[26157]_ ;
  assign \new_[26161]_  = ~A299 & A298;
  assign \new_[26164]_  = A302 & ~A301;
  assign \new_[26165]_  = \new_[26164]_  & \new_[26161]_ ;
  assign \new_[26166]_  = \new_[26165]_  & \new_[26158]_ ;
  assign \new_[26170]_  = ~A167 & A168;
  assign \new_[26171]_  = A170 & \new_[26170]_ ;
  assign \new_[26174]_  = ~A199 & A166;
  assign \new_[26177]_  = ~A201 & A200;
  assign \new_[26178]_  = \new_[26177]_  & \new_[26174]_ ;
  assign \new_[26179]_  = \new_[26178]_  & \new_[26171]_ ;
  assign \new_[26183]_  = A234 & A232;
  assign \new_[26184]_  = A202 & \new_[26183]_ ;
  assign \new_[26187]_  = A299 & ~A298;
  assign \new_[26190]_  = A302 & ~A301;
  assign \new_[26191]_  = \new_[26190]_  & \new_[26187]_ ;
  assign \new_[26192]_  = \new_[26191]_  & \new_[26184]_ ;
  assign \new_[26196]_  = ~A167 & A168;
  assign \new_[26197]_  = A170 & \new_[26196]_ ;
  assign \new_[26200]_  = ~A199 & A166;
  assign \new_[26203]_  = ~A201 & A200;
  assign \new_[26204]_  = \new_[26203]_  & \new_[26200]_ ;
  assign \new_[26205]_  = \new_[26204]_  & \new_[26197]_ ;
  assign \new_[26209]_  = A234 & A232;
  assign \new_[26210]_  = A202 & \new_[26209]_ ;
  assign \new_[26213]_  = ~A299 & ~A298;
  assign \new_[26216]_  = ~A302 & A301;
  assign \new_[26217]_  = \new_[26216]_  & \new_[26213]_ ;
  assign \new_[26218]_  = \new_[26217]_  & \new_[26210]_ ;
  assign \new_[26222]_  = ~A167 & A168;
  assign \new_[26223]_  = A170 & \new_[26222]_ ;
  assign \new_[26226]_  = ~A199 & A166;
  assign \new_[26229]_  = ~A201 & A200;
  assign \new_[26230]_  = \new_[26229]_  & \new_[26226]_ ;
  assign \new_[26231]_  = \new_[26230]_  & \new_[26223]_ ;
  assign \new_[26235]_  = A234 & A232;
  assign \new_[26236]_  = A202 & \new_[26235]_ ;
  assign \new_[26239]_  = A266 & A265;
  assign \new_[26242]_  = ~A269 & A268;
  assign \new_[26243]_  = \new_[26242]_  & \new_[26239]_ ;
  assign \new_[26244]_  = \new_[26243]_  & \new_[26236]_ ;
  assign \new_[26248]_  = ~A167 & A168;
  assign \new_[26249]_  = A170 & \new_[26248]_ ;
  assign \new_[26252]_  = ~A199 & A166;
  assign \new_[26255]_  = ~A201 & A200;
  assign \new_[26256]_  = \new_[26255]_  & \new_[26252]_ ;
  assign \new_[26257]_  = \new_[26256]_  & \new_[26249]_ ;
  assign \new_[26261]_  = A234 & A232;
  assign \new_[26262]_  = A202 & \new_[26261]_ ;
  assign \new_[26265]_  = A266 & ~A265;
  assign \new_[26268]_  = A269 & ~A268;
  assign \new_[26269]_  = \new_[26268]_  & \new_[26265]_ ;
  assign \new_[26270]_  = \new_[26269]_  & \new_[26262]_ ;
  assign \new_[26274]_  = ~A167 & A168;
  assign \new_[26275]_  = A170 & \new_[26274]_ ;
  assign \new_[26278]_  = ~A199 & A166;
  assign \new_[26281]_  = ~A201 & A200;
  assign \new_[26282]_  = \new_[26281]_  & \new_[26278]_ ;
  assign \new_[26283]_  = \new_[26282]_  & \new_[26275]_ ;
  assign \new_[26287]_  = A234 & A232;
  assign \new_[26288]_  = A202 & \new_[26287]_ ;
  assign \new_[26291]_  = ~A266 & A265;
  assign \new_[26294]_  = A269 & ~A268;
  assign \new_[26295]_  = \new_[26294]_  & \new_[26291]_ ;
  assign \new_[26296]_  = \new_[26295]_  & \new_[26288]_ ;
  assign \new_[26300]_  = ~A167 & A168;
  assign \new_[26301]_  = A170 & \new_[26300]_ ;
  assign \new_[26304]_  = ~A199 & A166;
  assign \new_[26307]_  = ~A201 & A200;
  assign \new_[26308]_  = \new_[26307]_  & \new_[26304]_ ;
  assign \new_[26309]_  = \new_[26308]_  & \new_[26301]_ ;
  assign \new_[26313]_  = A234 & A232;
  assign \new_[26314]_  = A202 & \new_[26313]_ ;
  assign \new_[26317]_  = ~A266 & ~A265;
  assign \new_[26320]_  = ~A269 & A268;
  assign \new_[26321]_  = \new_[26320]_  & \new_[26317]_ ;
  assign \new_[26322]_  = \new_[26321]_  & \new_[26314]_ ;
  assign \new_[26326]_  = ~A167 & A168;
  assign \new_[26327]_  = A170 & \new_[26326]_ ;
  assign \new_[26330]_  = ~A199 & A166;
  assign \new_[26333]_  = ~A201 & A200;
  assign \new_[26334]_  = \new_[26333]_  & \new_[26330]_ ;
  assign \new_[26335]_  = \new_[26334]_  & \new_[26327]_ ;
  assign \new_[26339]_  = A234 & A233;
  assign \new_[26340]_  = A202 & \new_[26339]_ ;
  assign \new_[26343]_  = A299 & A298;
  assign \new_[26346]_  = ~A302 & A301;
  assign \new_[26347]_  = \new_[26346]_  & \new_[26343]_ ;
  assign \new_[26348]_  = \new_[26347]_  & \new_[26340]_ ;
  assign \new_[26352]_  = ~A167 & A168;
  assign \new_[26353]_  = A170 & \new_[26352]_ ;
  assign \new_[26356]_  = ~A199 & A166;
  assign \new_[26359]_  = ~A201 & A200;
  assign \new_[26360]_  = \new_[26359]_  & \new_[26356]_ ;
  assign \new_[26361]_  = \new_[26360]_  & \new_[26353]_ ;
  assign \new_[26365]_  = A234 & A233;
  assign \new_[26366]_  = A202 & \new_[26365]_ ;
  assign \new_[26369]_  = ~A299 & A298;
  assign \new_[26372]_  = A302 & ~A301;
  assign \new_[26373]_  = \new_[26372]_  & \new_[26369]_ ;
  assign \new_[26374]_  = \new_[26373]_  & \new_[26366]_ ;
  assign \new_[26378]_  = ~A167 & A168;
  assign \new_[26379]_  = A170 & \new_[26378]_ ;
  assign \new_[26382]_  = ~A199 & A166;
  assign \new_[26385]_  = ~A201 & A200;
  assign \new_[26386]_  = \new_[26385]_  & \new_[26382]_ ;
  assign \new_[26387]_  = \new_[26386]_  & \new_[26379]_ ;
  assign \new_[26391]_  = A234 & A233;
  assign \new_[26392]_  = A202 & \new_[26391]_ ;
  assign \new_[26395]_  = A299 & ~A298;
  assign \new_[26398]_  = A302 & ~A301;
  assign \new_[26399]_  = \new_[26398]_  & \new_[26395]_ ;
  assign \new_[26400]_  = \new_[26399]_  & \new_[26392]_ ;
  assign \new_[26404]_  = ~A167 & A168;
  assign \new_[26405]_  = A170 & \new_[26404]_ ;
  assign \new_[26408]_  = ~A199 & A166;
  assign \new_[26411]_  = ~A201 & A200;
  assign \new_[26412]_  = \new_[26411]_  & \new_[26408]_ ;
  assign \new_[26413]_  = \new_[26412]_  & \new_[26405]_ ;
  assign \new_[26417]_  = A234 & A233;
  assign \new_[26418]_  = A202 & \new_[26417]_ ;
  assign \new_[26421]_  = ~A299 & ~A298;
  assign \new_[26424]_  = ~A302 & A301;
  assign \new_[26425]_  = \new_[26424]_  & \new_[26421]_ ;
  assign \new_[26426]_  = \new_[26425]_  & \new_[26418]_ ;
  assign \new_[26430]_  = ~A167 & A168;
  assign \new_[26431]_  = A170 & \new_[26430]_ ;
  assign \new_[26434]_  = ~A199 & A166;
  assign \new_[26437]_  = ~A201 & A200;
  assign \new_[26438]_  = \new_[26437]_  & \new_[26434]_ ;
  assign \new_[26439]_  = \new_[26438]_  & \new_[26431]_ ;
  assign \new_[26443]_  = A234 & A233;
  assign \new_[26444]_  = A202 & \new_[26443]_ ;
  assign \new_[26447]_  = A266 & A265;
  assign \new_[26450]_  = ~A269 & A268;
  assign \new_[26451]_  = \new_[26450]_  & \new_[26447]_ ;
  assign \new_[26452]_  = \new_[26451]_  & \new_[26444]_ ;
  assign \new_[26456]_  = ~A167 & A168;
  assign \new_[26457]_  = A170 & \new_[26456]_ ;
  assign \new_[26460]_  = ~A199 & A166;
  assign \new_[26463]_  = ~A201 & A200;
  assign \new_[26464]_  = \new_[26463]_  & \new_[26460]_ ;
  assign \new_[26465]_  = \new_[26464]_  & \new_[26457]_ ;
  assign \new_[26469]_  = A234 & A233;
  assign \new_[26470]_  = A202 & \new_[26469]_ ;
  assign \new_[26473]_  = A266 & ~A265;
  assign \new_[26476]_  = A269 & ~A268;
  assign \new_[26477]_  = \new_[26476]_  & \new_[26473]_ ;
  assign \new_[26478]_  = \new_[26477]_  & \new_[26470]_ ;
  assign \new_[26482]_  = ~A167 & A168;
  assign \new_[26483]_  = A170 & \new_[26482]_ ;
  assign \new_[26486]_  = ~A199 & A166;
  assign \new_[26489]_  = ~A201 & A200;
  assign \new_[26490]_  = \new_[26489]_  & \new_[26486]_ ;
  assign \new_[26491]_  = \new_[26490]_  & \new_[26483]_ ;
  assign \new_[26495]_  = A234 & A233;
  assign \new_[26496]_  = A202 & \new_[26495]_ ;
  assign \new_[26499]_  = ~A266 & A265;
  assign \new_[26502]_  = A269 & ~A268;
  assign \new_[26503]_  = \new_[26502]_  & \new_[26499]_ ;
  assign \new_[26504]_  = \new_[26503]_  & \new_[26496]_ ;
  assign \new_[26508]_  = ~A167 & A168;
  assign \new_[26509]_  = A170 & \new_[26508]_ ;
  assign \new_[26512]_  = ~A199 & A166;
  assign \new_[26515]_  = ~A201 & A200;
  assign \new_[26516]_  = \new_[26515]_  & \new_[26512]_ ;
  assign \new_[26517]_  = \new_[26516]_  & \new_[26509]_ ;
  assign \new_[26521]_  = A234 & A233;
  assign \new_[26522]_  = A202 & \new_[26521]_ ;
  assign \new_[26525]_  = ~A266 & ~A265;
  assign \new_[26528]_  = ~A269 & A268;
  assign \new_[26529]_  = \new_[26528]_  & \new_[26525]_ ;
  assign \new_[26530]_  = \new_[26529]_  & \new_[26522]_ ;
  assign \new_[26534]_  = ~A167 & A168;
  assign \new_[26535]_  = A170 & \new_[26534]_ ;
  assign \new_[26538]_  = ~A199 & A166;
  assign \new_[26541]_  = ~A201 & A200;
  assign \new_[26542]_  = \new_[26541]_  & \new_[26538]_ ;
  assign \new_[26543]_  = \new_[26542]_  & \new_[26535]_ ;
  assign \new_[26547]_  = A233 & A232;
  assign \new_[26548]_  = A202 & \new_[26547]_ ;
  assign \new_[26551]_  = ~A236 & A235;
  assign \new_[26554]_  = A300 & A299;
  assign \new_[26555]_  = \new_[26554]_  & \new_[26551]_ ;
  assign \new_[26556]_  = \new_[26555]_  & \new_[26548]_ ;
  assign \new_[26560]_  = ~A167 & A168;
  assign \new_[26561]_  = A170 & \new_[26560]_ ;
  assign \new_[26564]_  = ~A199 & A166;
  assign \new_[26567]_  = ~A201 & A200;
  assign \new_[26568]_  = \new_[26567]_  & \new_[26564]_ ;
  assign \new_[26569]_  = \new_[26568]_  & \new_[26561]_ ;
  assign \new_[26573]_  = A233 & A232;
  assign \new_[26574]_  = A202 & \new_[26573]_ ;
  assign \new_[26577]_  = ~A236 & A235;
  assign \new_[26580]_  = A300 & A298;
  assign \new_[26581]_  = \new_[26580]_  & \new_[26577]_ ;
  assign \new_[26582]_  = \new_[26581]_  & \new_[26574]_ ;
  assign \new_[26586]_  = ~A167 & A168;
  assign \new_[26587]_  = A170 & \new_[26586]_ ;
  assign \new_[26590]_  = ~A199 & A166;
  assign \new_[26593]_  = ~A201 & A200;
  assign \new_[26594]_  = \new_[26593]_  & \new_[26590]_ ;
  assign \new_[26595]_  = \new_[26594]_  & \new_[26587]_ ;
  assign \new_[26599]_  = A233 & A232;
  assign \new_[26600]_  = A202 & \new_[26599]_ ;
  assign \new_[26603]_  = ~A236 & A235;
  assign \new_[26606]_  = A267 & A265;
  assign \new_[26607]_  = \new_[26606]_  & \new_[26603]_ ;
  assign \new_[26608]_  = \new_[26607]_  & \new_[26600]_ ;
  assign \new_[26612]_  = ~A167 & A168;
  assign \new_[26613]_  = A170 & \new_[26612]_ ;
  assign \new_[26616]_  = ~A199 & A166;
  assign \new_[26619]_  = ~A201 & A200;
  assign \new_[26620]_  = \new_[26619]_  & \new_[26616]_ ;
  assign \new_[26621]_  = \new_[26620]_  & \new_[26613]_ ;
  assign \new_[26625]_  = A233 & A232;
  assign \new_[26626]_  = A202 & \new_[26625]_ ;
  assign \new_[26629]_  = ~A236 & A235;
  assign \new_[26632]_  = A267 & A266;
  assign \new_[26633]_  = \new_[26632]_  & \new_[26629]_ ;
  assign \new_[26634]_  = \new_[26633]_  & \new_[26626]_ ;
  assign \new_[26638]_  = ~A167 & A168;
  assign \new_[26639]_  = A170 & \new_[26638]_ ;
  assign \new_[26642]_  = ~A199 & A166;
  assign \new_[26645]_  = ~A201 & A200;
  assign \new_[26646]_  = \new_[26645]_  & \new_[26642]_ ;
  assign \new_[26647]_  = \new_[26646]_  & \new_[26639]_ ;
  assign \new_[26651]_  = A233 & ~A232;
  assign \new_[26652]_  = A202 & \new_[26651]_ ;
  assign \new_[26655]_  = A236 & ~A235;
  assign \new_[26658]_  = A300 & A299;
  assign \new_[26659]_  = \new_[26658]_  & \new_[26655]_ ;
  assign \new_[26660]_  = \new_[26659]_  & \new_[26652]_ ;
  assign \new_[26664]_  = ~A167 & A168;
  assign \new_[26665]_  = A170 & \new_[26664]_ ;
  assign \new_[26668]_  = ~A199 & A166;
  assign \new_[26671]_  = ~A201 & A200;
  assign \new_[26672]_  = \new_[26671]_  & \new_[26668]_ ;
  assign \new_[26673]_  = \new_[26672]_  & \new_[26665]_ ;
  assign \new_[26677]_  = A233 & ~A232;
  assign \new_[26678]_  = A202 & \new_[26677]_ ;
  assign \new_[26681]_  = A236 & ~A235;
  assign \new_[26684]_  = A300 & A298;
  assign \new_[26685]_  = \new_[26684]_  & \new_[26681]_ ;
  assign \new_[26686]_  = \new_[26685]_  & \new_[26678]_ ;
  assign \new_[26690]_  = ~A167 & A168;
  assign \new_[26691]_  = A170 & \new_[26690]_ ;
  assign \new_[26694]_  = ~A199 & A166;
  assign \new_[26697]_  = ~A201 & A200;
  assign \new_[26698]_  = \new_[26697]_  & \new_[26694]_ ;
  assign \new_[26699]_  = \new_[26698]_  & \new_[26691]_ ;
  assign \new_[26703]_  = A233 & ~A232;
  assign \new_[26704]_  = A202 & \new_[26703]_ ;
  assign \new_[26707]_  = A236 & ~A235;
  assign \new_[26710]_  = A267 & A265;
  assign \new_[26711]_  = \new_[26710]_  & \new_[26707]_ ;
  assign \new_[26712]_  = \new_[26711]_  & \new_[26704]_ ;
  assign \new_[26716]_  = ~A167 & A168;
  assign \new_[26717]_  = A170 & \new_[26716]_ ;
  assign \new_[26720]_  = ~A199 & A166;
  assign \new_[26723]_  = ~A201 & A200;
  assign \new_[26724]_  = \new_[26723]_  & \new_[26720]_ ;
  assign \new_[26725]_  = \new_[26724]_  & \new_[26717]_ ;
  assign \new_[26729]_  = A233 & ~A232;
  assign \new_[26730]_  = A202 & \new_[26729]_ ;
  assign \new_[26733]_  = A236 & ~A235;
  assign \new_[26736]_  = A267 & A266;
  assign \new_[26737]_  = \new_[26736]_  & \new_[26733]_ ;
  assign \new_[26738]_  = \new_[26737]_  & \new_[26730]_ ;
  assign \new_[26742]_  = ~A167 & A168;
  assign \new_[26743]_  = A170 & \new_[26742]_ ;
  assign \new_[26746]_  = ~A199 & A166;
  assign \new_[26749]_  = ~A201 & A200;
  assign \new_[26750]_  = \new_[26749]_  & \new_[26746]_ ;
  assign \new_[26751]_  = \new_[26750]_  & \new_[26743]_ ;
  assign \new_[26755]_  = ~A233 & A232;
  assign \new_[26756]_  = A202 & \new_[26755]_ ;
  assign \new_[26759]_  = A236 & ~A235;
  assign \new_[26762]_  = A300 & A299;
  assign \new_[26763]_  = \new_[26762]_  & \new_[26759]_ ;
  assign \new_[26764]_  = \new_[26763]_  & \new_[26756]_ ;
  assign \new_[26768]_  = ~A167 & A168;
  assign \new_[26769]_  = A170 & \new_[26768]_ ;
  assign \new_[26772]_  = ~A199 & A166;
  assign \new_[26775]_  = ~A201 & A200;
  assign \new_[26776]_  = \new_[26775]_  & \new_[26772]_ ;
  assign \new_[26777]_  = \new_[26776]_  & \new_[26769]_ ;
  assign \new_[26781]_  = ~A233 & A232;
  assign \new_[26782]_  = A202 & \new_[26781]_ ;
  assign \new_[26785]_  = A236 & ~A235;
  assign \new_[26788]_  = A300 & A298;
  assign \new_[26789]_  = \new_[26788]_  & \new_[26785]_ ;
  assign \new_[26790]_  = \new_[26789]_  & \new_[26782]_ ;
  assign \new_[26794]_  = ~A167 & A168;
  assign \new_[26795]_  = A170 & \new_[26794]_ ;
  assign \new_[26798]_  = ~A199 & A166;
  assign \new_[26801]_  = ~A201 & A200;
  assign \new_[26802]_  = \new_[26801]_  & \new_[26798]_ ;
  assign \new_[26803]_  = \new_[26802]_  & \new_[26795]_ ;
  assign \new_[26807]_  = ~A233 & A232;
  assign \new_[26808]_  = A202 & \new_[26807]_ ;
  assign \new_[26811]_  = A236 & ~A235;
  assign \new_[26814]_  = A267 & A265;
  assign \new_[26815]_  = \new_[26814]_  & \new_[26811]_ ;
  assign \new_[26816]_  = \new_[26815]_  & \new_[26808]_ ;
  assign \new_[26820]_  = ~A167 & A168;
  assign \new_[26821]_  = A170 & \new_[26820]_ ;
  assign \new_[26824]_  = ~A199 & A166;
  assign \new_[26827]_  = ~A201 & A200;
  assign \new_[26828]_  = \new_[26827]_  & \new_[26824]_ ;
  assign \new_[26829]_  = \new_[26828]_  & \new_[26821]_ ;
  assign \new_[26833]_  = ~A233 & A232;
  assign \new_[26834]_  = A202 & \new_[26833]_ ;
  assign \new_[26837]_  = A236 & ~A235;
  assign \new_[26840]_  = A267 & A266;
  assign \new_[26841]_  = \new_[26840]_  & \new_[26837]_ ;
  assign \new_[26842]_  = \new_[26841]_  & \new_[26834]_ ;
  assign \new_[26846]_  = ~A167 & A168;
  assign \new_[26847]_  = A170 & \new_[26846]_ ;
  assign \new_[26850]_  = ~A199 & A166;
  assign \new_[26853]_  = ~A201 & A200;
  assign \new_[26854]_  = \new_[26853]_  & \new_[26850]_ ;
  assign \new_[26855]_  = \new_[26854]_  & \new_[26847]_ ;
  assign \new_[26859]_  = ~A233 & ~A232;
  assign \new_[26860]_  = A202 & \new_[26859]_ ;
  assign \new_[26863]_  = ~A236 & A235;
  assign \new_[26866]_  = A300 & A299;
  assign \new_[26867]_  = \new_[26866]_  & \new_[26863]_ ;
  assign \new_[26868]_  = \new_[26867]_  & \new_[26860]_ ;
  assign \new_[26872]_  = ~A167 & A168;
  assign \new_[26873]_  = A170 & \new_[26872]_ ;
  assign \new_[26876]_  = ~A199 & A166;
  assign \new_[26879]_  = ~A201 & A200;
  assign \new_[26880]_  = \new_[26879]_  & \new_[26876]_ ;
  assign \new_[26881]_  = \new_[26880]_  & \new_[26873]_ ;
  assign \new_[26885]_  = ~A233 & ~A232;
  assign \new_[26886]_  = A202 & \new_[26885]_ ;
  assign \new_[26889]_  = ~A236 & A235;
  assign \new_[26892]_  = A300 & A298;
  assign \new_[26893]_  = \new_[26892]_  & \new_[26889]_ ;
  assign \new_[26894]_  = \new_[26893]_  & \new_[26886]_ ;
  assign \new_[26898]_  = ~A167 & A168;
  assign \new_[26899]_  = A170 & \new_[26898]_ ;
  assign \new_[26902]_  = ~A199 & A166;
  assign \new_[26905]_  = ~A201 & A200;
  assign \new_[26906]_  = \new_[26905]_  & \new_[26902]_ ;
  assign \new_[26907]_  = \new_[26906]_  & \new_[26899]_ ;
  assign \new_[26911]_  = ~A233 & ~A232;
  assign \new_[26912]_  = A202 & \new_[26911]_ ;
  assign \new_[26915]_  = ~A236 & A235;
  assign \new_[26918]_  = A267 & A265;
  assign \new_[26919]_  = \new_[26918]_  & \new_[26915]_ ;
  assign \new_[26920]_  = \new_[26919]_  & \new_[26912]_ ;
  assign \new_[26924]_  = ~A167 & A168;
  assign \new_[26925]_  = A170 & \new_[26924]_ ;
  assign \new_[26928]_  = ~A199 & A166;
  assign \new_[26931]_  = ~A201 & A200;
  assign \new_[26932]_  = \new_[26931]_  & \new_[26928]_ ;
  assign \new_[26933]_  = \new_[26932]_  & \new_[26925]_ ;
  assign \new_[26937]_  = ~A233 & ~A232;
  assign \new_[26938]_  = A202 & \new_[26937]_ ;
  assign \new_[26941]_  = ~A236 & A235;
  assign \new_[26944]_  = A267 & A266;
  assign \new_[26945]_  = \new_[26944]_  & \new_[26941]_ ;
  assign \new_[26946]_  = \new_[26945]_  & \new_[26938]_ ;
  assign \new_[26950]_  = ~A167 & A168;
  assign \new_[26951]_  = A170 & \new_[26950]_ ;
  assign \new_[26954]_  = ~A199 & A166;
  assign \new_[26957]_  = ~A201 & A200;
  assign \new_[26958]_  = \new_[26957]_  & \new_[26954]_ ;
  assign \new_[26959]_  = \new_[26958]_  & \new_[26951]_ ;
  assign \new_[26963]_  = A234 & A232;
  assign \new_[26964]_  = ~A203 & \new_[26963]_ ;
  assign \new_[26967]_  = A299 & A298;
  assign \new_[26970]_  = ~A302 & A301;
  assign \new_[26971]_  = \new_[26970]_  & \new_[26967]_ ;
  assign \new_[26972]_  = \new_[26971]_  & \new_[26964]_ ;
  assign \new_[26976]_  = ~A167 & A168;
  assign \new_[26977]_  = A170 & \new_[26976]_ ;
  assign \new_[26980]_  = ~A199 & A166;
  assign \new_[26983]_  = ~A201 & A200;
  assign \new_[26984]_  = \new_[26983]_  & \new_[26980]_ ;
  assign \new_[26985]_  = \new_[26984]_  & \new_[26977]_ ;
  assign \new_[26989]_  = A234 & A232;
  assign \new_[26990]_  = ~A203 & \new_[26989]_ ;
  assign \new_[26993]_  = ~A299 & A298;
  assign \new_[26996]_  = A302 & ~A301;
  assign \new_[26997]_  = \new_[26996]_  & \new_[26993]_ ;
  assign \new_[26998]_  = \new_[26997]_  & \new_[26990]_ ;
  assign \new_[27002]_  = ~A167 & A168;
  assign \new_[27003]_  = A170 & \new_[27002]_ ;
  assign \new_[27006]_  = ~A199 & A166;
  assign \new_[27009]_  = ~A201 & A200;
  assign \new_[27010]_  = \new_[27009]_  & \new_[27006]_ ;
  assign \new_[27011]_  = \new_[27010]_  & \new_[27003]_ ;
  assign \new_[27015]_  = A234 & A232;
  assign \new_[27016]_  = ~A203 & \new_[27015]_ ;
  assign \new_[27019]_  = A299 & ~A298;
  assign \new_[27022]_  = A302 & ~A301;
  assign \new_[27023]_  = \new_[27022]_  & \new_[27019]_ ;
  assign \new_[27024]_  = \new_[27023]_  & \new_[27016]_ ;
  assign \new_[27028]_  = ~A167 & A168;
  assign \new_[27029]_  = A170 & \new_[27028]_ ;
  assign \new_[27032]_  = ~A199 & A166;
  assign \new_[27035]_  = ~A201 & A200;
  assign \new_[27036]_  = \new_[27035]_  & \new_[27032]_ ;
  assign \new_[27037]_  = \new_[27036]_  & \new_[27029]_ ;
  assign \new_[27041]_  = A234 & A232;
  assign \new_[27042]_  = ~A203 & \new_[27041]_ ;
  assign \new_[27045]_  = ~A299 & ~A298;
  assign \new_[27048]_  = ~A302 & A301;
  assign \new_[27049]_  = \new_[27048]_  & \new_[27045]_ ;
  assign \new_[27050]_  = \new_[27049]_  & \new_[27042]_ ;
  assign \new_[27054]_  = ~A167 & A168;
  assign \new_[27055]_  = A170 & \new_[27054]_ ;
  assign \new_[27058]_  = ~A199 & A166;
  assign \new_[27061]_  = ~A201 & A200;
  assign \new_[27062]_  = \new_[27061]_  & \new_[27058]_ ;
  assign \new_[27063]_  = \new_[27062]_  & \new_[27055]_ ;
  assign \new_[27067]_  = A234 & A232;
  assign \new_[27068]_  = ~A203 & \new_[27067]_ ;
  assign \new_[27071]_  = A266 & A265;
  assign \new_[27074]_  = ~A269 & A268;
  assign \new_[27075]_  = \new_[27074]_  & \new_[27071]_ ;
  assign \new_[27076]_  = \new_[27075]_  & \new_[27068]_ ;
  assign \new_[27080]_  = ~A167 & A168;
  assign \new_[27081]_  = A170 & \new_[27080]_ ;
  assign \new_[27084]_  = ~A199 & A166;
  assign \new_[27087]_  = ~A201 & A200;
  assign \new_[27088]_  = \new_[27087]_  & \new_[27084]_ ;
  assign \new_[27089]_  = \new_[27088]_  & \new_[27081]_ ;
  assign \new_[27093]_  = A234 & A232;
  assign \new_[27094]_  = ~A203 & \new_[27093]_ ;
  assign \new_[27097]_  = A266 & ~A265;
  assign \new_[27100]_  = A269 & ~A268;
  assign \new_[27101]_  = \new_[27100]_  & \new_[27097]_ ;
  assign \new_[27102]_  = \new_[27101]_  & \new_[27094]_ ;
  assign \new_[27106]_  = ~A167 & A168;
  assign \new_[27107]_  = A170 & \new_[27106]_ ;
  assign \new_[27110]_  = ~A199 & A166;
  assign \new_[27113]_  = ~A201 & A200;
  assign \new_[27114]_  = \new_[27113]_  & \new_[27110]_ ;
  assign \new_[27115]_  = \new_[27114]_  & \new_[27107]_ ;
  assign \new_[27119]_  = A234 & A232;
  assign \new_[27120]_  = ~A203 & \new_[27119]_ ;
  assign \new_[27123]_  = ~A266 & A265;
  assign \new_[27126]_  = A269 & ~A268;
  assign \new_[27127]_  = \new_[27126]_  & \new_[27123]_ ;
  assign \new_[27128]_  = \new_[27127]_  & \new_[27120]_ ;
  assign \new_[27132]_  = ~A167 & A168;
  assign \new_[27133]_  = A170 & \new_[27132]_ ;
  assign \new_[27136]_  = ~A199 & A166;
  assign \new_[27139]_  = ~A201 & A200;
  assign \new_[27140]_  = \new_[27139]_  & \new_[27136]_ ;
  assign \new_[27141]_  = \new_[27140]_  & \new_[27133]_ ;
  assign \new_[27145]_  = A234 & A232;
  assign \new_[27146]_  = ~A203 & \new_[27145]_ ;
  assign \new_[27149]_  = ~A266 & ~A265;
  assign \new_[27152]_  = ~A269 & A268;
  assign \new_[27153]_  = \new_[27152]_  & \new_[27149]_ ;
  assign \new_[27154]_  = \new_[27153]_  & \new_[27146]_ ;
  assign \new_[27158]_  = ~A167 & A168;
  assign \new_[27159]_  = A170 & \new_[27158]_ ;
  assign \new_[27162]_  = ~A199 & A166;
  assign \new_[27165]_  = ~A201 & A200;
  assign \new_[27166]_  = \new_[27165]_  & \new_[27162]_ ;
  assign \new_[27167]_  = \new_[27166]_  & \new_[27159]_ ;
  assign \new_[27171]_  = A234 & A233;
  assign \new_[27172]_  = ~A203 & \new_[27171]_ ;
  assign \new_[27175]_  = A299 & A298;
  assign \new_[27178]_  = ~A302 & A301;
  assign \new_[27179]_  = \new_[27178]_  & \new_[27175]_ ;
  assign \new_[27180]_  = \new_[27179]_  & \new_[27172]_ ;
  assign \new_[27184]_  = ~A167 & A168;
  assign \new_[27185]_  = A170 & \new_[27184]_ ;
  assign \new_[27188]_  = ~A199 & A166;
  assign \new_[27191]_  = ~A201 & A200;
  assign \new_[27192]_  = \new_[27191]_  & \new_[27188]_ ;
  assign \new_[27193]_  = \new_[27192]_  & \new_[27185]_ ;
  assign \new_[27197]_  = A234 & A233;
  assign \new_[27198]_  = ~A203 & \new_[27197]_ ;
  assign \new_[27201]_  = ~A299 & A298;
  assign \new_[27204]_  = A302 & ~A301;
  assign \new_[27205]_  = \new_[27204]_  & \new_[27201]_ ;
  assign \new_[27206]_  = \new_[27205]_  & \new_[27198]_ ;
  assign \new_[27210]_  = ~A167 & A168;
  assign \new_[27211]_  = A170 & \new_[27210]_ ;
  assign \new_[27214]_  = ~A199 & A166;
  assign \new_[27217]_  = ~A201 & A200;
  assign \new_[27218]_  = \new_[27217]_  & \new_[27214]_ ;
  assign \new_[27219]_  = \new_[27218]_  & \new_[27211]_ ;
  assign \new_[27223]_  = A234 & A233;
  assign \new_[27224]_  = ~A203 & \new_[27223]_ ;
  assign \new_[27227]_  = A299 & ~A298;
  assign \new_[27230]_  = A302 & ~A301;
  assign \new_[27231]_  = \new_[27230]_  & \new_[27227]_ ;
  assign \new_[27232]_  = \new_[27231]_  & \new_[27224]_ ;
  assign \new_[27236]_  = ~A167 & A168;
  assign \new_[27237]_  = A170 & \new_[27236]_ ;
  assign \new_[27240]_  = ~A199 & A166;
  assign \new_[27243]_  = ~A201 & A200;
  assign \new_[27244]_  = \new_[27243]_  & \new_[27240]_ ;
  assign \new_[27245]_  = \new_[27244]_  & \new_[27237]_ ;
  assign \new_[27249]_  = A234 & A233;
  assign \new_[27250]_  = ~A203 & \new_[27249]_ ;
  assign \new_[27253]_  = ~A299 & ~A298;
  assign \new_[27256]_  = ~A302 & A301;
  assign \new_[27257]_  = \new_[27256]_  & \new_[27253]_ ;
  assign \new_[27258]_  = \new_[27257]_  & \new_[27250]_ ;
  assign \new_[27262]_  = ~A167 & A168;
  assign \new_[27263]_  = A170 & \new_[27262]_ ;
  assign \new_[27266]_  = ~A199 & A166;
  assign \new_[27269]_  = ~A201 & A200;
  assign \new_[27270]_  = \new_[27269]_  & \new_[27266]_ ;
  assign \new_[27271]_  = \new_[27270]_  & \new_[27263]_ ;
  assign \new_[27275]_  = A234 & A233;
  assign \new_[27276]_  = ~A203 & \new_[27275]_ ;
  assign \new_[27279]_  = A266 & A265;
  assign \new_[27282]_  = ~A269 & A268;
  assign \new_[27283]_  = \new_[27282]_  & \new_[27279]_ ;
  assign \new_[27284]_  = \new_[27283]_  & \new_[27276]_ ;
  assign \new_[27288]_  = ~A167 & A168;
  assign \new_[27289]_  = A170 & \new_[27288]_ ;
  assign \new_[27292]_  = ~A199 & A166;
  assign \new_[27295]_  = ~A201 & A200;
  assign \new_[27296]_  = \new_[27295]_  & \new_[27292]_ ;
  assign \new_[27297]_  = \new_[27296]_  & \new_[27289]_ ;
  assign \new_[27301]_  = A234 & A233;
  assign \new_[27302]_  = ~A203 & \new_[27301]_ ;
  assign \new_[27305]_  = A266 & ~A265;
  assign \new_[27308]_  = A269 & ~A268;
  assign \new_[27309]_  = \new_[27308]_  & \new_[27305]_ ;
  assign \new_[27310]_  = \new_[27309]_  & \new_[27302]_ ;
  assign \new_[27314]_  = ~A167 & A168;
  assign \new_[27315]_  = A170 & \new_[27314]_ ;
  assign \new_[27318]_  = ~A199 & A166;
  assign \new_[27321]_  = ~A201 & A200;
  assign \new_[27322]_  = \new_[27321]_  & \new_[27318]_ ;
  assign \new_[27323]_  = \new_[27322]_  & \new_[27315]_ ;
  assign \new_[27327]_  = A234 & A233;
  assign \new_[27328]_  = ~A203 & \new_[27327]_ ;
  assign \new_[27331]_  = ~A266 & A265;
  assign \new_[27334]_  = A269 & ~A268;
  assign \new_[27335]_  = \new_[27334]_  & \new_[27331]_ ;
  assign \new_[27336]_  = \new_[27335]_  & \new_[27328]_ ;
  assign \new_[27340]_  = ~A167 & A168;
  assign \new_[27341]_  = A170 & \new_[27340]_ ;
  assign \new_[27344]_  = ~A199 & A166;
  assign \new_[27347]_  = ~A201 & A200;
  assign \new_[27348]_  = \new_[27347]_  & \new_[27344]_ ;
  assign \new_[27349]_  = \new_[27348]_  & \new_[27341]_ ;
  assign \new_[27353]_  = A234 & A233;
  assign \new_[27354]_  = ~A203 & \new_[27353]_ ;
  assign \new_[27357]_  = ~A266 & ~A265;
  assign \new_[27360]_  = ~A269 & A268;
  assign \new_[27361]_  = \new_[27360]_  & \new_[27357]_ ;
  assign \new_[27362]_  = \new_[27361]_  & \new_[27354]_ ;
  assign \new_[27366]_  = ~A167 & A168;
  assign \new_[27367]_  = A170 & \new_[27366]_ ;
  assign \new_[27370]_  = ~A199 & A166;
  assign \new_[27373]_  = ~A201 & A200;
  assign \new_[27374]_  = \new_[27373]_  & \new_[27370]_ ;
  assign \new_[27375]_  = \new_[27374]_  & \new_[27367]_ ;
  assign \new_[27379]_  = A233 & A232;
  assign \new_[27380]_  = ~A203 & \new_[27379]_ ;
  assign \new_[27383]_  = ~A236 & A235;
  assign \new_[27386]_  = A300 & A299;
  assign \new_[27387]_  = \new_[27386]_  & \new_[27383]_ ;
  assign \new_[27388]_  = \new_[27387]_  & \new_[27380]_ ;
  assign \new_[27392]_  = ~A167 & A168;
  assign \new_[27393]_  = A170 & \new_[27392]_ ;
  assign \new_[27396]_  = ~A199 & A166;
  assign \new_[27399]_  = ~A201 & A200;
  assign \new_[27400]_  = \new_[27399]_  & \new_[27396]_ ;
  assign \new_[27401]_  = \new_[27400]_  & \new_[27393]_ ;
  assign \new_[27405]_  = A233 & A232;
  assign \new_[27406]_  = ~A203 & \new_[27405]_ ;
  assign \new_[27409]_  = ~A236 & A235;
  assign \new_[27412]_  = A300 & A298;
  assign \new_[27413]_  = \new_[27412]_  & \new_[27409]_ ;
  assign \new_[27414]_  = \new_[27413]_  & \new_[27406]_ ;
  assign \new_[27418]_  = ~A167 & A168;
  assign \new_[27419]_  = A170 & \new_[27418]_ ;
  assign \new_[27422]_  = ~A199 & A166;
  assign \new_[27425]_  = ~A201 & A200;
  assign \new_[27426]_  = \new_[27425]_  & \new_[27422]_ ;
  assign \new_[27427]_  = \new_[27426]_  & \new_[27419]_ ;
  assign \new_[27431]_  = A233 & A232;
  assign \new_[27432]_  = ~A203 & \new_[27431]_ ;
  assign \new_[27435]_  = ~A236 & A235;
  assign \new_[27438]_  = A267 & A265;
  assign \new_[27439]_  = \new_[27438]_  & \new_[27435]_ ;
  assign \new_[27440]_  = \new_[27439]_  & \new_[27432]_ ;
  assign \new_[27444]_  = ~A167 & A168;
  assign \new_[27445]_  = A170 & \new_[27444]_ ;
  assign \new_[27448]_  = ~A199 & A166;
  assign \new_[27451]_  = ~A201 & A200;
  assign \new_[27452]_  = \new_[27451]_  & \new_[27448]_ ;
  assign \new_[27453]_  = \new_[27452]_  & \new_[27445]_ ;
  assign \new_[27457]_  = A233 & A232;
  assign \new_[27458]_  = ~A203 & \new_[27457]_ ;
  assign \new_[27461]_  = ~A236 & A235;
  assign \new_[27464]_  = A267 & A266;
  assign \new_[27465]_  = \new_[27464]_  & \new_[27461]_ ;
  assign \new_[27466]_  = \new_[27465]_  & \new_[27458]_ ;
  assign \new_[27470]_  = ~A167 & A168;
  assign \new_[27471]_  = A170 & \new_[27470]_ ;
  assign \new_[27474]_  = ~A199 & A166;
  assign \new_[27477]_  = ~A201 & A200;
  assign \new_[27478]_  = \new_[27477]_  & \new_[27474]_ ;
  assign \new_[27479]_  = \new_[27478]_  & \new_[27471]_ ;
  assign \new_[27483]_  = A233 & ~A232;
  assign \new_[27484]_  = ~A203 & \new_[27483]_ ;
  assign \new_[27487]_  = A236 & ~A235;
  assign \new_[27490]_  = A300 & A299;
  assign \new_[27491]_  = \new_[27490]_  & \new_[27487]_ ;
  assign \new_[27492]_  = \new_[27491]_  & \new_[27484]_ ;
  assign \new_[27496]_  = ~A167 & A168;
  assign \new_[27497]_  = A170 & \new_[27496]_ ;
  assign \new_[27500]_  = ~A199 & A166;
  assign \new_[27503]_  = ~A201 & A200;
  assign \new_[27504]_  = \new_[27503]_  & \new_[27500]_ ;
  assign \new_[27505]_  = \new_[27504]_  & \new_[27497]_ ;
  assign \new_[27509]_  = A233 & ~A232;
  assign \new_[27510]_  = ~A203 & \new_[27509]_ ;
  assign \new_[27513]_  = A236 & ~A235;
  assign \new_[27516]_  = A300 & A298;
  assign \new_[27517]_  = \new_[27516]_  & \new_[27513]_ ;
  assign \new_[27518]_  = \new_[27517]_  & \new_[27510]_ ;
  assign \new_[27522]_  = ~A167 & A168;
  assign \new_[27523]_  = A170 & \new_[27522]_ ;
  assign \new_[27526]_  = ~A199 & A166;
  assign \new_[27529]_  = ~A201 & A200;
  assign \new_[27530]_  = \new_[27529]_  & \new_[27526]_ ;
  assign \new_[27531]_  = \new_[27530]_  & \new_[27523]_ ;
  assign \new_[27535]_  = A233 & ~A232;
  assign \new_[27536]_  = ~A203 & \new_[27535]_ ;
  assign \new_[27539]_  = A236 & ~A235;
  assign \new_[27542]_  = A267 & A265;
  assign \new_[27543]_  = \new_[27542]_  & \new_[27539]_ ;
  assign \new_[27544]_  = \new_[27543]_  & \new_[27536]_ ;
  assign \new_[27548]_  = ~A167 & A168;
  assign \new_[27549]_  = A170 & \new_[27548]_ ;
  assign \new_[27552]_  = ~A199 & A166;
  assign \new_[27555]_  = ~A201 & A200;
  assign \new_[27556]_  = \new_[27555]_  & \new_[27552]_ ;
  assign \new_[27557]_  = \new_[27556]_  & \new_[27549]_ ;
  assign \new_[27561]_  = A233 & ~A232;
  assign \new_[27562]_  = ~A203 & \new_[27561]_ ;
  assign \new_[27565]_  = A236 & ~A235;
  assign \new_[27568]_  = A267 & A266;
  assign \new_[27569]_  = \new_[27568]_  & \new_[27565]_ ;
  assign \new_[27570]_  = \new_[27569]_  & \new_[27562]_ ;
  assign \new_[27574]_  = ~A167 & A168;
  assign \new_[27575]_  = A170 & \new_[27574]_ ;
  assign \new_[27578]_  = ~A199 & A166;
  assign \new_[27581]_  = ~A201 & A200;
  assign \new_[27582]_  = \new_[27581]_  & \new_[27578]_ ;
  assign \new_[27583]_  = \new_[27582]_  & \new_[27575]_ ;
  assign \new_[27587]_  = ~A233 & A232;
  assign \new_[27588]_  = ~A203 & \new_[27587]_ ;
  assign \new_[27591]_  = A236 & ~A235;
  assign \new_[27594]_  = A300 & A299;
  assign \new_[27595]_  = \new_[27594]_  & \new_[27591]_ ;
  assign \new_[27596]_  = \new_[27595]_  & \new_[27588]_ ;
  assign \new_[27600]_  = ~A167 & A168;
  assign \new_[27601]_  = A170 & \new_[27600]_ ;
  assign \new_[27604]_  = ~A199 & A166;
  assign \new_[27607]_  = ~A201 & A200;
  assign \new_[27608]_  = \new_[27607]_  & \new_[27604]_ ;
  assign \new_[27609]_  = \new_[27608]_  & \new_[27601]_ ;
  assign \new_[27613]_  = ~A233 & A232;
  assign \new_[27614]_  = ~A203 & \new_[27613]_ ;
  assign \new_[27617]_  = A236 & ~A235;
  assign \new_[27620]_  = A300 & A298;
  assign \new_[27621]_  = \new_[27620]_  & \new_[27617]_ ;
  assign \new_[27622]_  = \new_[27621]_  & \new_[27614]_ ;
  assign \new_[27626]_  = ~A167 & A168;
  assign \new_[27627]_  = A170 & \new_[27626]_ ;
  assign \new_[27630]_  = ~A199 & A166;
  assign \new_[27633]_  = ~A201 & A200;
  assign \new_[27634]_  = \new_[27633]_  & \new_[27630]_ ;
  assign \new_[27635]_  = \new_[27634]_  & \new_[27627]_ ;
  assign \new_[27639]_  = ~A233 & A232;
  assign \new_[27640]_  = ~A203 & \new_[27639]_ ;
  assign \new_[27643]_  = A236 & ~A235;
  assign \new_[27646]_  = A267 & A265;
  assign \new_[27647]_  = \new_[27646]_  & \new_[27643]_ ;
  assign \new_[27648]_  = \new_[27647]_  & \new_[27640]_ ;
  assign \new_[27652]_  = ~A167 & A168;
  assign \new_[27653]_  = A170 & \new_[27652]_ ;
  assign \new_[27656]_  = ~A199 & A166;
  assign \new_[27659]_  = ~A201 & A200;
  assign \new_[27660]_  = \new_[27659]_  & \new_[27656]_ ;
  assign \new_[27661]_  = \new_[27660]_  & \new_[27653]_ ;
  assign \new_[27665]_  = ~A233 & A232;
  assign \new_[27666]_  = ~A203 & \new_[27665]_ ;
  assign \new_[27669]_  = A236 & ~A235;
  assign \new_[27672]_  = A267 & A266;
  assign \new_[27673]_  = \new_[27672]_  & \new_[27669]_ ;
  assign \new_[27674]_  = \new_[27673]_  & \new_[27666]_ ;
  assign \new_[27678]_  = ~A167 & A168;
  assign \new_[27679]_  = A170 & \new_[27678]_ ;
  assign \new_[27682]_  = ~A199 & A166;
  assign \new_[27685]_  = ~A201 & A200;
  assign \new_[27686]_  = \new_[27685]_  & \new_[27682]_ ;
  assign \new_[27687]_  = \new_[27686]_  & \new_[27679]_ ;
  assign \new_[27691]_  = ~A233 & ~A232;
  assign \new_[27692]_  = ~A203 & \new_[27691]_ ;
  assign \new_[27695]_  = ~A236 & A235;
  assign \new_[27698]_  = A300 & A299;
  assign \new_[27699]_  = \new_[27698]_  & \new_[27695]_ ;
  assign \new_[27700]_  = \new_[27699]_  & \new_[27692]_ ;
  assign \new_[27704]_  = ~A167 & A168;
  assign \new_[27705]_  = A170 & \new_[27704]_ ;
  assign \new_[27708]_  = ~A199 & A166;
  assign \new_[27711]_  = ~A201 & A200;
  assign \new_[27712]_  = \new_[27711]_  & \new_[27708]_ ;
  assign \new_[27713]_  = \new_[27712]_  & \new_[27705]_ ;
  assign \new_[27717]_  = ~A233 & ~A232;
  assign \new_[27718]_  = ~A203 & \new_[27717]_ ;
  assign \new_[27721]_  = ~A236 & A235;
  assign \new_[27724]_  = A300 & A298;
  assign \new_[27725]_  = \new_[27724]_  & \new_[27721]_ ;
  assign \new_[27726]_  = \new_[27725]_  & \new_[27718]_ ;
  assign \new_[27730]_  = ~A167 & A168;
  assign \new_[27731]_  = A170 & \new_[27730]_ ;
  assign \new_[27734]_  = ~A199 & A166;
  assign \new_[27737]_  = ~A201 & A200;
  assign \new_[27738]_  = \new_[27737]_  & \new_[27734]_ ;
  assign \new_[27739]_  = \new_[27738]_  & \new_[27731]_ ;
  assign \new_[27743]_  = ~A233 & ~A232;
  assign \new_[27744]_  = ~A203 & \new_[27743]_ ;
  assign \new_[27747]_  = ~A236 & A235;
  assign \new_[27750]_  = A267 & A265;
  assign \new_[27751]_  = \new_[27750]_  & \new_[27747]_ ;
  assign \new_[27752]_  = \new_[27751]_  & \new_[27744]_ ;
  assign \new_[27756]_  = ~A167 & A168;
  assign \new_[27757]_  = A170 & \new_[27756]_ ;
  assign \new_[27760]_  = ~A199 & A166;
  assign \new_[27763]_  = ~A201 & A200;
  assign \new_[27764]_  = \new_[27763]_  & \new_[27760]_ ;
  assign \new_[27765]_  = \new_[27764]_  & \new_[27757]_ ;
  assign \new_[27769]_  = ~A233 & ~A232;
  assign \new_[27770]_  = ~A203 & \new_[27769]_ ;
  assign \new_[27773]_  = ~A236 & A235;
  assign \new_[27776]_  = A267 & A266;
  assign \new_[27777]_  = \new_[27776]_  & \new_[27773]_ ;
  assign \new_[27778]_  = \new_[27777]_  & \new_[27770]_ ;
  assign \new_[27782]_  = ~A167 & A168;
  assign \new_[27783]_  = A170 & \new_[27782]_ ;
  assign \new_[27786]_  = A199 & A166;
  assign \new_[27789]_  = ~A201 & ~A200;
  assign \new_[27790]_  = \new_[27789]_  & \new_[27786]_ ;
  assign \new_[27791]_  = \new_[27790]_  & \new_[27783]_ ;
  assign \new_[27795]_  = A234 & A232;
  assign \new_[27796]_  = A202 & \new_[27795]_ ;
  assign \new_[27799]_  = A299 & A298;
  assign \new_[27802]_  = ~A302 & A301;
  assign \new_[27803]_  = \new_[27802]_  & \new_[27799]_ ;
  assign \new_[27804]_  = \new_[27803]_  & \new_[27796]_ ;
  assign \new_[27808]_  = ~A167 & A168;
  assign \new_[27809]_  = A170 & \new_[27808]_ ;
  assign \new_[27812]_  = A199 & A166;
  assign \new_[27815]_  = ~A201 & ~A200;
  assign \new_[27816]_  = \new_[27815]_  & \new_[27812]_ ;
  assign \new_[27817]_  = \new_[27816]_  & \new_[27809]_ ;
  assign \new_[27821]_  = A234 & A232;
  assign \new_[27822]_  = A202 & \new_[27821]_ ;
  assign \new_[27825]_  = ~A299 & A298;
  assign \new_[27828]_  = A302 & ~A301;
  assign \new_[27829]_  = \new_[27828]_  & \new_[27825]_ ;
  assign \new_[27830]_  = \new_[27829]_  & \new_[27822]_ ;
  assign \new_[27834]_  = ~A167 & A168;
  assign \new_[27835]_  = A170 & \new_[27834]_ ;
  assign \new_[27838]_  = A199 & A166;
  assign \new_[27841]_  = ~A201 & ~A200;
  assign \new_[27842]_  = \new_[27841]_  & \new_[27838]_ ;
  assign \new_[27843]_  = \new_[27842]_  & \new_[27835]_ ;
  assign \new_[27847]_  = A234 & A232;
  assign \new_[27848]_  = A202 & \new_[27847]_ ;
  assign \new_[27851]_  = A299 & ~A298;
  assign \new_[27854]_  = A302 & ~A301;
  assign \new_[27855]_  = \new_[27854]_  & \new_[27851]_ ;
  assign \new_[27856]_  = \new_[27855]_  & \new_[27848]_ ;
  assign \new_[27860]_  = ~A167 & A168;
  assign \new_[27861]_  = A170 & \new_[27860]_ ;
  assign \new_[27864]_  = A199 & A166;
  assign \new_[27867]_  = ~A201 & ~A200;
  assign \new_[27868]_  = \new_[27867]_  & \new_[27864]_ ;
  assign \new_[27869]_  = \new_[27868]_  & \new_[27861]_ ;
  assign \new_[27873]_  = A234 & A232;
  assign \new_[27874]_  = A202 & \new_[27873]_ ;
  assign \new_[27877]_  = ~A299 & ~A298;
  assign \new_[27880]_  = ~A302 & A301;
  assign \new_[27881]_  = \new_[27880]_  & \new_[27877]_ ;
  assign \new_[27882]_  = \new_[27881]_  & \new_[27874]_ ;
  assign \new_[27886]_  = ~A167 & A168;
  assign \new_[27887]_  = A170 & \new_[27886]_ ;
  assign \new_[27890]_  = A199 & A166;
  assign \new_[27893]_  = ~A201 & ~A200;
  assign \new_[27894]_  = \new_[27893]_  & \new_[27890]_ ;
  assign \new_[27895]_  = \new_[27894]_  & \new_[27887]_ ;
  assign \new_[27899]_  = A234 & A232;
  assign \new_[27900]_  = A202 & \new_[27899]_ ;
  assign \new_[27903]_  = A266 & A265;
  assign \new_[27906]_  = ~A269 & A268;
  assign \new_[27907]_  = \new_[27906]_  & \new_[27903]_ ;
  assign \new_[27908]_  = \new_[27907]_  & \new_[27900]_ ;
  assign \new_[27912]_  = ~A167 & A168;
  assign \new_[27913]_  = A170 & \new_[27912]_ ;
  assign \new_[27916]_  = A199 & A166;
  assign \new_[27919]_  = ~A201 & ~A200;
  assign \new_[27920]_  = \new_[27919]_  & \new_[27916]_ ;
  assign \new_[27921]_  = \new_[27920]_  & \new_[27913]_ ;
  assign \new_[27925]_  = A234 & A232;
  assign \new_[27926]_  = A202 & \new_[27925]_ ;
  assign \new_[27929]_  = A266 & ~A265;
  assign \new_[27932]_  = A269 & ~A268;
  assign \new_[27933]_  = \new_[27932]_  & \new_[27929]_ ;
  assign \new_[27934]_  = \new_[27933]_  & \new_[27926]_ ;
  assign \new_[27938]_  = ~A167 & A168;
  assign \new_[27939]_  = A170 & \new_[27938]_ ;
  assign \new_[27942]_  = A199 & A166;
  assign \new_[27945]_  = ~A201 & ~A200;
  assign \new_[27946]_  = \new_[27945]_  & \new_[27942]_ ;
  assign \new_[27947]_  = \new_[27946]_  & \new_[27939]_ ;
  assign \new_[27951]_  = A234 & A232;
  assign \new_[27952]_  = A202 & \new_[27951]_ ;
  assign \new_[27955]_  = ~A266 & A265;
  assign \new_[27958]_  = A269 & ~A268;
  assign \new_[27959]_  = \new_[27958]_  & \new_[27955]_ ;
  assign \new_[27960]_  = \new_[27959]_  & \new_[27952]_ ;
  assign \new_[27964]_  = ~A167 & A168;
  assign \new_[27965]_  = A170 & \new_[27964]_ ;
  assign \new_[27968]_  = A199 & A166;
  assign \new_[27971]_  = ~A201 & ~A200;
  assign \new_[27972]_  = \new_[27971]_  & \new_[27968]_ ;
  assign \new_[27973]_  = \new_[27972]_  & \new_[27965]_ ;
  assign \new_[27977]_  = A234 & A232;
  assign \new_[27978]_  = A202 & \new_[27977]_ ;
  assign \new_[27981]_  = ~A266 & ~A265;
  assign \new_[27984]_  = ~A269 & A268;
  assign \new_[27985]_  = \new_[27984]_  & \new_[27981]_ ;
  assign \new_[27986]_  = \new_[27985]_  & \new_[27978]_ ;
  assign \new_[27990]_  = ~A167 & A168;
  assign \new_[27991]_  = A170 & \new_[27990]_ ;
  assign \new_[27994]_  = A199 & A166;
  assign \new_[27997]_  = ~A201 & ~A200;
  assign \new_[27998]_  = \new_[27997]_  & \new_[27994]_ ;
  assign \new_[27999]_  = \new_[27998]_  & \new_[27991]_ ;
  assign \new_[28003]_  = A234 & A233;
  assign \new_[28004]_  = A202 & \new_[28003]_ ;
  assign \new_[28007]_  = A299 & A298;
  assign \new_[28010]_  = ~A302 & A301;
  assign \new_[28011]_  = \new_[28010]_  & \new_[28007]_ ;
  assign \new_[28012]_  = \new_[28011]_  & \new_[28004]_ ;
  assign \new_[28016]_  = ~A167 & A168;
  assign \new_[28017]_  = A170 & \new_[28016]_ ;
  assign \new_[28020]_  = A199 & A166;
  assign \new_[28023]_  = ~A201 & ~A200;
  assign \new_[28024]_  = \new_[28023]_  & \new_[28020]_ ;
  assign \new_[28025]_  = \new_[28024]_  & \new_[28017]_ ;
  assign \new_[28029]_  = A234 & A233;
  assign \new_[28030]_  = A202 & \new_[28029]_ ;
  assign \new_[28033]_  = ~A299 & A298;
  assign \new_[28036]_  = A302 & ~A301;
  assign \new_[28037]_  = \new_[28036]_  & \new_[28033]_ ;
  assign \new_[28038]_  = \new_[28037]_  & \new_[28030]_ ;
  assign \new_[28042]_  = ~A167 & A168;
  assign \new_[28043]_  = A170 & \new_[28042]_ ;
  assign \new_[28046]_  = A199 & A166;
  assign \new_[28049]_  = ~A201 & ~A200;
  assign \new_[28050]_  = \new_[28049]_  & \new_[28046]_ ;
  assign \new_[28051]_  = \new_[28050]_  & \new_[28043]_ ;
  assign \new_[28055]_  = A234 & A233;
  assign \new_[28056]_  = A202 & \new_[28055]_ ;
  assign \new_[28059]_  = A299 & ~A298;
  assign \new_[28062]_  = A302 & ~A301;
  assign \new_[28063]_  = \new_[28062]_  & \new_[28059]_ ;
  assign \new_[28064]_  = \new_[28063]_  & \new_[28056]_ ;
  assign \new_[28068]_  = ~A167 & A168;
  assign \new_[28069]_  = A170 & \new_[28068]_ ;
  assign \new_[28072]_  = A199 & A166;
  assign \new_[28075]_  = ~A201 & ~A200;
  assign \new_[28076]_  = \new_[28075]_  & \new_[28072]_ ;
  assign \new_[28077]_  = \new_[28076]_  & \new_[28069]_ ;
  assign \new_[28081]_  = A234 & A233;
  assign \new_[28082]_  = A202 & \new_[28081]_ ;
  assign \new_[28085]_  = ~A299 & ~A298;
  assign \new_[28088]_  = ~A302 & A301;
  assign \new_[28089]_  = \new_[28088]_  & \new_[28085]_ ;
  assign \new_[28090]_  = \new_[28089]_  & \new_[28082]_ ;
  assign \new_[28094]_  = ~A167 & A168;
  assign \new_[28095]_  = A170 & \new_[28094]_ ;
  assign \new_[28098]_  = A199 & A166;
  assign \new_[28101]_  = ~A201 & ~A200;
  assign \new_[28102]_  = \new_[28101]_  & \new_[28098]_ ;
  assign \new_[28103]_  = \new_[28102]_  & \new_[28095]_ ;
  assign \new_[28107]_  = A234 & A233;
  assign \new_[28108]_  = A202 & \new_[28107]_ ;
  assign \new_[28111]_  = A266 & A265;
  assign \new_[28114]_  = ~A269 & A268;
  assign \new_[28115]_  = \new_[28114]_  & \new_[28111]_ ;
  assign \new_[28116]_  = \new_[28115]_  & \new_[28108]_ ;
  assign \new_[28120]_  = ~A167 & A168;
  assign \new_[28121]_  = A170 & \new_[28120]_ ;
  assign \new_[28124]_  = A199 & A166;
  assign \new_[28127]_  = ~A201 & ~A200;
  assign \new_[28128]_  = \new_[28127]_  & \new_[28124]_ ;
  assign \new_[28129]_  = \new_[28128]_  & \new_[28121]_ ;
  assign \new_[28133]_  = A234 & A233;
  assign \new_[28134]_  = A202 & \new_[28133]_ ;
  assign \new_[28137]_  = A266 & ~A265;
  assign \new_[28140]_  = A269 & ~A268;
  assign \new_[28141]_  = \new_[28140]_  & \new_[28137]_ ;
  assign \new_[28142]_  = \new_[28141]_  & \new_[28134]_ ;
  assign \new_[28146]_  = ~A167 & A168;
  assign \new_[28147]_  = A170 & \new_[28146]_ ;
  assign \new_[28150]_  = A199 & A166;
  assign \new_[28153]_  = ~A201 & ~A200;
  assign \new_[28154]_  = \new_[28153]_  & \new_[28150]_ ;
  assign \new_[28155]_  = \new_[28154]_  & \new_[28147]_ ;
  assign \new_[28159]_  = A234 & A233;
  assign \new_[28160]_  = A202 & \new_[28159]_ ;
  assign \new_[28163]_  = ~A266 & A265;
  assign \new_[28166]_  = A269 & ~A268;
  assign \new_[28167]_  = \new_[28166]_  & \new_[28163]_ ;
  assign \new_[28168]_  = \new_[28167]_  & \new_[28160]_ ;
  assign \new_[28172]_  = ~A167 & A168;
  assign \new_[28173]_  = A170 & \new_[28172]_ ;
  assign \new_[28176]_  = A199 & A166;
  assign \new_[28179]_  = ~A201 & ~A200;
  assign \new_[28180]_  = \new_[28179]_  & \new_[28176]_ ;
  assign \new_[28181]_  = \new_[28180]_  & \new_[28173]_ ;
  assign \new_[28185]_  = A234 & A233;
  assign \new_[28186]_  = A202 & \new_[28185]_ ;
  assign \new_[28189]_  = ~A266 & ~A265;
  assign \new_[28192]_  = ~A269 & A268;
  assign \new_[28193]_  = \new_[28192]_  & \new_[28189]_ ;
  assign \new_[28194]_  = \new_[28193]_  & \new_[28186]_ ;
  assign \new_[28198]_  = ~A167 & A168;
  assign \new_[28199]_  = A170 & \new_[28198]_ ;
  assign \new_[28202]_  = A199 & A166;
  assign \new_[28205]_  = ~A201 & ~A200;
  assign \new_[28206]_  = \new_[28205]_  & \new_[28202]_ ;
  assign \new_[28207]_  = \new_[28206]_  & \new_[28199]_ ;
  assign \new_[28211]_  = A233 & A232;
  assign \new_[28212]_  = A202 & \new_[28211]_ ;
  assign \new_[28215]_  = ~A236 & A235;
  assign \new_[28218]_  = A300 & A299;
  assign \new_[28219]_  = \new_[28218]_  & \new_[28215]_ ;
  assign \new_[28220]_  = \new_[28219]_  & \new_[28212]_ ;
  assign \new_[28224]_  = ~A167 & A168;
  assign \new_[28225]_  = A170 & \new_[28224]_ ;
  assign \new_[28228]_  = A199 & A166;
  assign \new_[28231]_  = ~A201 & ~A200;
  assign \new_[28232]_  = \new_[28231]_  & \new_[28228]_ ;
  assign \new_[28233]_  = \new_[28232]_  & \new_[28225]_ ;
  assign \new_[28237]_  = A233 & A232;
  assign \new_[28238]_  = A202 & \new_[28237]_ ;
  assign \new_[28241]_  = ~A236 & A235;
  assign \new_[28244]_  = A300 & A298;
  assign \new_[28245]_  = \new_[28244]_  & \new_[28241]_ ;
  assign \new_[28246]_  = \new_[28245]_  & \new_[28238]_ ;
  assign \new_[28250]_  = ~A167 & A168;
  assign \new_[28251]_  = A170 & \new_[28250]_ ;
  assign \new_[28254]_  = A199 & A166;
  assign \new_[28257]_  = ~A201 & ~A200;
  assign \new_[28258]_  = \new_[28257]_  & \new_[28254]_ ;
  assign \new_[28259]_  = \new_[28258]_  & \new_[28251]_ ;
  assign \new_[28263]_  = A233 & A232;
  assign \new_[28264]_  = A202 & \new_[28263]_ ;
  assign \new_[28267]_  = ~A236 & A235;
  assign \new_[28270]_  = A267 & A265;
  assign \new_[28271]_  = \new_[28270]_  & \new_[28267]_ ;
  assign \new_[28272]_  = \new_[28271]_  & \new_[28264]_ ;
  assign \new_[28276]_  = ~A167 & A168;
  assign \new_[28277]_  = A170 & \new_[28276]_ ;
  assign \new_[28280]_  = A199 & A166;
  assign \new_[28283]_  = ~A201 & ~A200;
  assign \new_[28284]_  = \new_[28283]_  & \new_[28280]_ ;
  assign \new_[28285]_  = \new_[28284]_  & \new_[28277]_ ;
  assign \new_[28289]_  = A233 & A232;
  assign \new_[28290]_  = A202 & \new_[28289]_ ;
  assign \new_[28293]_  = ~A236 & A235;
  assign \new_[28296]_  = A267 & A266;
  assign \new_[28297]_  = \new_[28296]_  & \new_[28293]_ ;
  assign \new_[28298]_  = \new_[28297]_  & \new_[28290]_ ;
  assign \new_[28302]_  = ~A167 & A168;
  assign \new_[28303]_  = A170 & \new_[28302]_ ;
  assign \new_[28306]_  = A199 & A166;
  assign \new_[28309]_  = ~A201 & ~A200;
  assign \new_[28310]_  = \new_[28309]_  & \new_[28306]_ ;
  assign \new_[28311]_  = \new_[28310]_  & \new_[28303]_ ;
  assign \new_[28315]_  = A233 & ~A232;
  assign \new_[28316]_  = A202 & \new_[28315]_ ;
  assign \new_[28319]_  = A236 & ~A235;
  assign \new_[28322]_  = A300 & A299;
  assign \new_[28323]_  = \new_[28322]_  & \new_[28319]_ ;
  assign \new_[28324]_  = \new_[28323]_  & \new_[28316]_ ;
  assign \new_[28328]_  = ~A167 & A168;
  assign \new_[28329]_  = A170 & \new_[28328]_ ;
  assign \new_[28332]_  = A199 & A166;
  assign \new_[28335]_  = ~A201 & ~A200;
  assign \new_[28336]_  = \new_[28335]_  & \new_[28332]_ ;
  assign \new_[28337]_  = \new_[28336]_  & \new_[28329]_ ;
  assign \new_[28341]_  = A233 & ~A232;
  assign \new_[28342]_  = A202 & \new_[28341]_ ;
  assign \new_[28345]_  = A236 & ~A235;
  assign \new_[28348]_  = A300 & A298;
  assign \new_[28349]_  = \new_[28348]_  & \new_[28345]_ ;
  assign \new_[28350]_  = \new_[28349]_  & \new_[28342]_ ;
  assign \new_[28354]_  = ~A167 & A168;
  assign \new_[28355]_  = A170 & \new_[28354]_ ;
  assign \new_[28358]_  = A199 & A166;
  assign \new_[28361]_  = ~A201 & ~A200;
  assign \new_[28362]_  = \new_[28361]_  & \new_[28358]_ ;
  assign \new_[28363]_  = \new_[28362]_  & \new_[28355]_ ;
  assign \new_[28367]_  = A233 & ~A232;
  assign \new_[28368]_  = A202 & \new_[28367]_ ;
  assign \new_[28371]_  = A236 & ~A235;
  assign \new_[28374]_  = A267 & A265;
  assign \new_[28375]_  = \new_[28374]_  & \new_[28371]_ ;
  assign \new_[28376]_  = \new_[28375]_  & \new_[28368]_ ;
  assign \new_[28380]_  = ~A167 & A168;
  assign \new_[28381]_  = A170 & \new_[28380]_ ;
  assign \new_[28384]_  = A199 & A166;
  assign \new_[28387]_  = ~A201 & ~A200;
  assign \new_[28388]_  = \new_[28387]_  & \new_[28384]_ ;
  assign \new_[28389]_  = \new_[28388]_  & \new_[28381]_ ;
  assign \new_[28393]_  = A233 & ~A232;
  assign \new_[28394]_  = A202 & \new_[28393]_ ;
  assign \new_[28397]_  = A236 & ~A235;
  assign \new_[28400]_  = A267 & A266;
  assign \new_[28401]_  = \new_[28400]_  & \new_[28397]_ ;
  assign \new_[28402]_  = \new_[28401]_  & \new_[28394]_ ;
  assign \new_[28406]_  = ~A167 & A168;
  assign \new_[28407]_  = A170 & \new_[28406]_ ;
  assign \new_[28410]_  = A199 & A166;
  assign \new_[28413]_  = ~A201 & ~A200;
  assign \new_[28414]_  = \new_[28413]_  & \new_[28410]_ ;
  assign \new_[28415]_  = \new_[28414]_  & \new_[28407]_ ;
  assign \new_[28419]_  = ~A233 & A232;
  assign \new_[28420]_  = A202 & \new_[28419]_ ;
  assign \new_[28423]_  = A236 & ~A235;
  assign \new_[28426]_  = A300 & A299;
  assign \new_[28427]_  = \new_[28426]_  & \new_[28423]_ ;
  assign \new_[28428]_  = \new_[28427]_  & \new_[28420]_ ;
  assign \new_[28432]_  = ~A167 & A168;
  assign \new_[28433]_  = A170 & \new_[28432]_ ;
  assign \new_[28436]_  = A199 & A166;
  assign \new_[28439]_  = ~A201 & ~A200;
  assign \new_[28440]_  = \new_[28439]_  & \new_[28436]_ ;
  assign \new_[28441]_  = \new_[28440]_  & \new_[28433]_ ;
  assign \new_[28445]_  = ~A233 & A232;
  assign \new_[28446]_  = A202 & \new_[28445]_ ;
  assign \new_[28449]_  = A236 & ~A235;
  assign \new_[28452]_  = A300 & A298;
  assign \new_[28453]_  = \new_[28452]_  & \new_[28449]_ ;
  assign \new_[28454]_  = \new_[28453]_  & \new_[28446]_ ;
  assign \new_[28458]_  = ~A167 & A168;
  assign \new_[28459]_  = A170 & \new_[28458]_ ;
  assign \new_[28462]_  = A199 & A166;
  assign \new_[28465]_  = ~A201 & ~A200;
  assign \new_[28466]_  = \new_[28465]_  & \new_[28462]_ ;
  assign \new_[28467]_  = \new_[28466]_  & \new_[28459]_ ;
  assign \new_[28471]_  = ~A233 & A232;
  assign \new_[28472]_  = A202 & \new_[28471]_ ;
  assign \new_[28475]_  = A236 & ~A235;
  assign \new_[28478]_  = A267 & A265;
  assign \new_[28479]_  = \new_[28478]_  & \new_[28475]_ ;
  assign \new_[28480]_  = \new_[28479]_  & \new_[28472]_ ;
  assign \new_[28484]_  = ~A167 & A168;
  assign \new_[28485]_  = A170 & \new_[28484]_ ;
  assign \new_[28488]_  = A199 & A166;
  assign \new_[28491]_  = ~A201 & ~A200;
  assign \new_[28492]_  = \new_[28491]_  & \new_[28488]_ ;
  assign \new_[28493]_  = \new_[28492]_  & \new_[28485]_ ;
  assign \new_[28497]_  = ~A233 & A232;
  assign \new_[28498]_  = A202 & \new_[28497]_ ;
  assign \new_[28501]_  = A236 & ~A235;
  assign \new_[28504]_  = A267 & A266;
  assign \new_[28505]_  = \new_[28504]_  & \new_[28501]_ ;
  assign \new_[28506]_  = \new_[28505]_  & \new_[28498]_ ;
  assign \new_[28510]_  = ~A167 & A168;
  assign \new_[28511]_  = A170 & \new_[28510]_ ;
  assign \new_[28514]_  = A199 & A166;
  assign \new_[28517]_  = ~A201 & ~A200;
  assign \new_[28518]_  = \new_[28517]_  & \new_[28514]_ ;
  assign \new_[28519]_  = \new_[28518]_  & \new_[28511]_ ;
  assign \new_[28523]_  = ~A233 & ~A232;
  assign \new_[28524]_  = A202 & \new_[28523]_ ;
  assign \new_[28527]_  = ~A236 & A235;
  assign \new_[28530]_  = A300 & A299;
  assign \new_[28531]_  = \new_[28530]_  & \new_[28527]_ ;
  assign \new_[28532]_  = \new_[28531]_  & \new_[28524]_ ;
  assign \new_[28536]_  = ~A167 & A168;
  assign \new_[28537]_  = A170 & \new_[28536]_ ;
  assign \new_[28540]_  = A199 & A166;
  assign \new_[28543]_  = ~A201 & ~A200;
  assign \new_[28544]_  = \new_[28543]_  & \new_[28540]_ ;
  assign \new_[28545]_  = \new_[28544]_  & \new_[28537]_ ;
  assign \new_[28549]_  = ~A233 & ~A232;
  assign \new_[28550]_  = A202 & \new_[28549]_ ;
  assign \new_[28553]_  = ~A236 & A235;
  assign \new_[28556]_  = A300 & A298;
  assign \new_[28557]_  = \new_[28556]_  & \new_[28553]_ ;
  assign \new_[28558]_  = \new_[28557]_  & \new_[28550]_ ;
  assign \new_[28562]_  = ~A167 & A168;
  assign \new_[28563]_  = A170 & \new_[28562]_ ;
  assign \new_[28566]_  = A199 & A166;
  assign \new_[28569]_  = ~A201 & ~A200;
  assign \new_[28570]_  = \new_[28569]_  & \new_[28566]_ ;
  assign \new_[28571]_  = \new_[28570]_  & \new_[28563]_ ;
  assign \new_[28575]_  = ~A233 & ~A232;
  assign \new_[28576]_  = A202 & \new_[28575]_ ;
  assign \new_[28579]_  = ~A236 & A235;
  assign \new_[28582]_  = A267 & A265;
  assign \new_[28583]_  = \new_[28582]_  & \new_[28579]_ ;
  assign \new_[28584]_  = \new_[28583]_  & \new_[28576]_ ;
  assign \new_[28588]_  = ~A167 & A168;
  assign \new_[28589]_  = A170 & \new_[28588]_ ;
  assign \new_[28592]_  = A199 & A166;
  assign \new_[28595]_  = ~A201 & ~A200;
  assign \new_[28596]_  = \new_[28595]_  & \new_[28592]_ ;
  assign \new_[28597]_  = \new_[28596]_  & \new_[28589]_ ;
  assign \new_[28601]_  = ~A233 & ~A232;
  assign \new_[28602]_  = A202 & \new_[28601]_ ;
  assign \new_[28605]_  = ~A236 & A235;
  assign \new_[28608]_  = A267 & A266;
  assign \new_[28609]_  = \new_[28608]_  & \new_[28605]_ ;
  assign \new_[28610]_  = \new_[28609]_  & \new_[28602]_ ;
  assign \new_[28614]_  = ~A167 & A168;
  assign \new_[28615]_  = A170 & \new_[28614]_ ;
  assign \new_[28618]_  = A199 & A166;
  assign \new_[28621]_  = ~A201 & ~A200;
  assign \new_[28622]_  = \new_[28621]_  & \new_[28618]_ ;
  assign \new_[28623]_  = \new_[28622]_  & \new_[28615]_ ;
  assign \new_[28627]_  = A234 & A232;
  assign \new_[28628]_  = ~A203 & \new_[28627]_ ;
  assign \new_[28631]_  = A299 & A298;
  assign \new_[28634]_  = ~A302 & A301;
  assign \new_[28635]_  = \new_[28634]_  & \new_[28631]_ ;
  assign \new_[28636]_  = \new_[28635]_  & \new_[28628]_ ;
  assign \new_[28640]_  = ~A167 & A168;
  assign \new_[28641]_  = A170 & \new_[28640]_ ;
  assign \new_[28644]_  = A199 & A166;
  assign \new_[28647]_  = ~A201 & ~A200;
  assign \new_[28648]_  = \new_[28647]_  & \new_[28644]_ ;
  assign \new_[28649]_  = \new_[28648]_  & \new_[28641]_ ;
  assign \new_[28653]_  = A234 & A232;
  assign \new_[28654]_  = ~A203 & \new_[28653]_ ;
  assign \new_[28657]_  = ~A299 & A298;
  assign \new_[28660]_  = A302 & ~A301;
  assign \new_[28661]_  = \new_[28660]_  & \new_[28657]_ ;
  assign \new_[28662]_  = \new_[28661]_  & \new_[28654]_ ;
  assign \new_[28666]_  = ~A167 & A168;
  assign \new_[28667]_  = A170 & \new_[28666]_ ;
  assign \new_[28670]_  = A199 & A166;
  assign \new_[28673]_  = ~A201 & ~A200;
  assign \new_[28674]_  = \new_[28673]_  & \new_[28670]_ ;
  assign \new_[28675]_  = \new_[28674]_  & \new_[28667]_ ;
  assign \new_[28679]_  = A234 & A232;
  assign \new_[28680]_  = ~A203 & \new_[28679]_ ;
  assign \new_[28683]_  = A299 & ~A298;
  assign \new_[28686]_  = A302 & ~A301;
  assign \new_[28687]_  = \new_[28686]_  & \new_[28683]_ ;
  assign \new_[28688]_  = \new_[28687]_  & \new_[28680]_ ;
  assign \new_[28692]_  = ~A167 & A168;
  assign \new_[28693]_  = A170 & \new_[28692]_ ;
  assign \new_[28696]_  = A199 & A166;
  assign \new_[28699]_  = ~A201 & ~A200;
  assign \new_[28700]_  = \new_[28699]_  & \new_[28696]_ ;
  assign \new_[28701]_  = \new_[28700]_  & \new_[28693]_ ;
  assign \new_[28705]_  = A234 & A232;
  assign \new_[28706]_  = ~A203 & \new_[28705]_ ;
  assign \new_[28709]_  = ~A299 & ~A298;
  assign \new_[28712]_  = ~A302 & A301;
  assign \new_[28713]_  = \new_[28712]_  & \new_[28709]_ ;
  assign \new_[28714]_  = \new_[28713]_  & \new_[28706]_ ;
  assign \new_[28718]_  = ~A167 & A168;
  assign \new_[28719]_  = A170 & \new_[28718]_ ;
  assign \new_[28722]_  = A199 & A166;
  assign \new_[28725]_  = ~A201 & ~A200;
  assign \new_[28726]_  = \new_[28725]_  & \new_[28722]_ ;
  assign \new_[28727]_  = \new_[28726]_  & \new_[28719]_ ;
  assign \new_[28731]_  = A234 & A232;
  assign \new_[28732]_  = ~A203 & \new_[28731]_ ;
  assign \new_[28735]_  = A266 & A265;
  assign \new_[28738]_  = ~A269 & A268;
  assign \new_[28739]_  = \new_[28738]_  & \new_[28735]_ ;
  assign \new_[28740]_  = \new_[28739]_  & \new_[28732]_ ;
  assign \new_[28744]_  = ~A167 & A168;
  assign \new_[28745]_  = A170 & \new_[28744]_ ;
  assign \new_[28748]_  = A199 & A166;
  assign \new_[28751]_  = ~A201 & ~A200;
  assign \new_[28752]_  = \new_[28751]_  & \new_[28748]_ ;
  assign \new_[28753]_  = \new_[28752]_  & \new_[28745]_ ;
  assign \new_[28757]_  = A234 & A232;
  assign \new_[28758]_  = ~A203 & \new_[28757]_ ;
  assign \new_[28761]_  = A266 & ~A265;
  assign \new_[28764]_  = A269 & ~A268;
  assign \new_[28765]_  = \new_[28764]_  & \new_[28761]_ ;
  assign \new_[28766]_  = \new_[28765]_  & \new_[28758]_ ;
  assign \new_[28770]_  = ~A167 & A168;
  assign \new_[28771]_  = A170 & \new_[28770]_ ;
  assign \new_[28774]_  = A199 & A166;
  assign \new_[28777]_  = ~A201 & ~A200;
  assign \new_[28778]_  = \new_[28777]_  & \new_[28774]_ ;
  assign \new_[28779]_  = \new_[28778]_  & \new_[28771]_ ;
  assign \new_[28783]_  = A234 & A232;
  assign \new_[28784]_  = ~A203 & \new_[28783]_ ;
  assign \new_[28787]_  = ~A266 & A265;
  assign \new_[28790]_  = A269 & ~A268;
  assign \new_[28791]_  = \new_[28790]_  & \new_[28787]_ ;
  assign \new_[28792]_  = \new_[28791]_  & \new_[28784]_ ;
  assign \new_[28796]_  = ~A167 & A168;
  assign \new_[28797]_  = A170 & \new_[28796]_ ;
  assign \new_[28800]_  = A199 & A166;
  assign \new_[28803]_  = ~A201 & ~A200;
  assign \new_[28804]_  = \new_[28803]_  & \new_[28800]_ ;
  assign \new_[28805]_  = \new_[28804]_  & \new_[28797]_ ;
  assign \new_[28809]_  = A234 & A232;
  assign \new_[28810]_  = ~A203 & \new_[28809]_ ;
  assign \new_[28813]_  = ~A266 & ~A265;
  assign \new_[28816]_  = ~A269 & A268;
  assign \new_[28817]_  = \new_[28816]_  & \new_[28813]_ ;
  assign \new_[28818]_  = \new_[28817]_  & \new_[28810]_ ;
  assign \new_[28822]_  = ~A167 & A168;
  assign \new_[28823]_  = A170 & \new_[28822]_ ;
  assign \new_[28826]_  = A199 & A166;
  assign \new_[28829]_  = ~A201 & ~A200;
  assign \new_[28830]_  = \new_[28829]_  & \new_[28826]_ ;
  assign \new_[28831]_  = \new_[28830]_  & \new_[28823]_ ;
  assign \new_[28835]_  = A234 & A233;
  assign \new_[28836]_  = ~A203 & \new_[28835]_ ;
  assign \new_[28839]_  = A299 & A298;
  assign \new_[28842]_  = ~A302 & A301;
  assign \new_[28843]_  = \new_[28842]_  & \new_[28839]_ ;
  assign \new_[28844]_  = \new_[28843]_  & \new_[28836]_ ;
  assign \new_[28848]_  = ~A167 & A168;
  assign \new_[28849]_  = A170 & \new_[28848]_ ;
  assign \new_[28852]_  = A199 & A166;
  assign \new_[28855]_  = ~A201 & ~A200;
  assign \new_[28856]_  = \new_[28855]_  & \new_[28852]_ ;
  assign \new_[28857]_  = \new_[28856]_  & \new_[28849]_ ;
  assign \new_[28861]_  = A234 & A233;
  assign \new_[28862]_  = ~A203 & \new_[28861]_ ;
  assign \new_[28865]_  = ~A299 & A298;
  assign \new_[28868]_  = A302 & ~A301;
  assign \new_[28869]_  = \new_[28868]_  & \new_[28865]_ ;
  assign \new_[28870]_  = \new_[28869]_  & \new_[28862]_ ;
  assign \new_[28874]_  = ~A167 & A168;
  assign \new_[28875]_  = A170 & \new_[28874]_ ;
  assign \new_[28878]_  = A199 & A166;
  assign \new_[28881]_  = ~A201 & ~A200;
  assign \new_[28882]_  = \new_[28881]_  & \new_[28878]_ ;
  assign \new_[28883]_  = \new_[28882]_  & \new_[28875]_ ;
  assign \new_[28887]_  = A234 & A233;
  assign \new_[28888]_  = ~A203 & \new_[28887]_ ;
  assign \new_[28891]_  = A299 & ~A298;
  assign \new_[28894]_  = A302 & ~A301;
  assign \new_[28895]_  = \new_[28894]_  & \new_[28891]_ ;
  assign \new_[28896]_  = \new_[28895]_  & \new_[28888]_ ;
  assign \new_[28900]_  = ~A167 & A168;
  assign \new_[28901]_  = A170 & \new_[28900]_ ;
  assign \new_[28904]_  = A199 & A166;
  assign \new_[28907]_  = ~A201 & ~A200;
  assign \new_[28908]_  = \new_[28907]_  & \new_[28904]_ ;
  assign \new_[28909]_  = \new_[28908]_  & \new_[28901]_ ;
  assign \new_[28913]_  = A234 & A233;
  assign \new_[28914]_  = ~A203 & \new_[28913]_ ;
  assign \new_[28917]_  = ~A299 & ~A298;
  assign \new_[28920]_  = ~A302 & A301;
  assign \new_[28921]_  = \new_[28920]_  & \new_[28917]_ ;
  assign \new_[28922]_  = \new_[28921]_  & \new_[28914]_ ;
  assign \new_[28926]_  = ~A167 & A168;
  assign \new_[28927]_  = A170 & \new_[28926]_ ;
  assign \new_[28930]_  = A199 & A166;
  assign \new_[28933]_  = ~A201 & ~A200;
  assign \new_[28934]_  = \new_[28933]_  & \new_[28930]_ ;
  assign \new_[28935]_  = \new_[28934]_  & \new_[28927]_ ;
  assign \new_[28939]_  = A234 & A233;
  assign \new_[28940]_  = ~A203 & \new_[28939]_ ;
  assign \new_[28943]_  = A266 & A265;
  assign \new_[28946]_  = ~A269 & A268;
  assign \new_[28947]_  = \new_[28946]_  & \new_[28943]_ ;
  assign \new_[28948]_  = \new_[28947]_  & \new_[28940]_ ;
  assign \new_[28952]_  = ~A167 & A168;
  assign \new_[28953]_  = A170 & \new_[28952]_ ;
  assign \new_[28956]_  = A199 & A166;
  assign \new_[28959]_  = ~A201 & ~A200;
  assign \new_[28960]_  = \new_[28959]_  & \new_[28956]_ ;
  assign \new_[28961]_  = \new_[28960]_  & \new_[28953]_ ;
  assign \new_[28965]_  = A234 & A233;
  assign \new_[28966]_  = ~A203 & \new_[28965]_ ;
  assign \new_[28969]_  = A266 & ~A265;
  assign \new_[28972]_  = A269 & ~A268;
  assign \new_[28973]_  = \new_[28972]_  & \new_[28969]_ ;
  assign \new_[28974]_  = \new_[28973]_  & \new_[28966]_ ;
  assign \new_[28978]_  = ~A167 & A168;
  assign \new_[28979]_  = A170 & \new_[28978]_ ;
  assign \new_[28982]_  = A199 & A166;
  assign \new_[28985]_  = ~A201 & ~A200;
  assign \new_[28986]_  = \new_[28985]_  & \new_[28982]_ ;
  assign \new_[28987]_  = \new_[28986]_  & \new_[28979]_ ;
  assign \new_[28991]_  = A234 & A233;
  assign \new_[28992]_  = ~A203 & \new_[28991]_ ;
  assign \new_[28995]_  = ~A266 & A265;
  assign \new_[28998]_  = A269 & ~A268;
  assign \new_[28999]_  = \new_[28998]_  & \new_[28995]_ ;
  assign \new_[29000]_  = \new_[28999]_  & \new_[28992]_ ;
  assign \new_[29004]_  = ~A167 & A168;
  assign \new_[29005]_  = A170 & \new_[29004]_ ;
  assign \new_[29008]_  = A199 & A166;
  assign \new_[29011]_  = ~A201 & ~A200;
  assign \new_[29012]_  = \new_[29011]_  & \new_[29008]_ ;
  assign \new_[29013]_  = \new_[29012]_  & \new_[29005]_ ;
  assign \new_[29017]_  = A234 & A233;
  assign \new_[29018]_  = ~A203 & \new_[29017]_ ;
  assign \new_[29021]_  = ~A266 & ~A265;
  assign \new_[29024]_  = ~A269 & A268;
  assign \new_[29025]_  = \new_[29024]_  & \new_[29021]_ ;
  assign \new_[29026]_  = \new_[29025]_  & \new_[29018]_ ;
  assign \new_[29030]_  = ~A167 & A168;
  assign \new_[29031]_  = A170 & \new_[29030]_ ;
  assign \new_[29034]_  = A199 & A166;
  assign \new_[29037]_  = ~A201 & ~A200;
  assign \new_[29038]_  = \new_[29037]_  & \new_[29034]_ ;
  assign \new_[29039]_  = \new_[29038]_  & \new_[29031]_ ;
  assign \new_[29043]_  = A233 & A232;
  assign \new_[29044]_  = ~A203 & \new_[29043]_ ;
  assign \new_[29047]_  = ~A236 & A235;
  assign \new_[29050]_  = A300 & A299;
  assign \new_[29051]_  = \new_[29050]_  & \new_[29047]_ ;
  assign \new_[29052]_  = \new_[29051]_  & \new_[29044]_ ;
  assign \new_[29056]_  = ~A167 & A168;
  assign \new_[29057]_  = A170 & \new_[29056]_ ;
  assign \new_[29060]_  = A199 & A166;
  assign \new_[29063]_  = ~A201 & ~A200;
  assign \new_[29064]_  = \new_[29063]_  & \new_[29060]_ ;
  assign \new_[29065]_  = \new_[29064]_  & \new_[29057]_ ;
  assign \new_[29069]_  = A233 & A232;
  assign \new_[29070]_  = ~A203 & \new_[29069]_ ;
  assign \new_[29073]_  = ~A236 & A235;
  assign \new_[29076]_  = A300 & A298;
  assign \new_[29077]_  = \new_[29076]_  & \new_[29073]_ ;
  assign \new_[29078]_  = \new_[29077]_  & \new_[29070]_ ;
  assign \new_[29082]_  = ~A167 & A168;
  assign \new_[29083]_  = A170 & \new_[29082]_ ;
  assign \new_[29086]_  = A199 & A166;
  assign \new_[29089]_  = ~A201 & ~A200;
  assign \new_[29090]_  = \new_[29089]_  & \new_[29086]_ ;
  assign \new_[29091]_  = \new_[29090]_  & \new_[29083]_ ;
  assign \new_[29095]_  = A233 & A232;
  assign \new_[29096]_  = ~A203 & \new_[29095]_ ;
  assign \new_[29099]_  = ~A236 & A235;
  assign \new_[29102]_  = A267 & A265;
  assign \new_[29103]_  = \new_[29102]_  & \new_[29099]_ ;
  assign \new_[29104]_  = \new_[29103]_  & \new_[29096]_ ;
  assign \new_[29108]_  = ~A167 & A168;
  assign \new_[29109]_  = A170 & \new_[29108]_ ;
  assign \new_[29112]_  = A199 & A166;
  assign \new_[29115]_  = ~A201 & ~A200;
  assign \new_[29116]_  = \new_[29115]_  & \new_[29112]_ ;
  assign \new_[29117]_  = \new_[29116]_  & \new_[29109]_ ;
  assign \new_[29121]_  = A233 & A232;
  assign \new_[29122]_  = ~A203 & \new_[29121]_ ;
  assign \new_[29125]_  = ~A236 & A235;
  assign \new_[29128]_  = A267 & A266;
  assign \new_[29129]_  = \new_[29128]_  & \new_[29125]_ ;
  assign \new_[29130]_  = \new_[29129]_  & \new_[29122]_ ;
  assign \new_[29134]_  = ~A167 & A168;
  assign \new_[29135]_  = A170 & \new_[29134]_ ;
  assign \new_[29138]_  = A199 & A166;
  assign \new_[29141]_  = ~A201 & ~A200;
  assign \new_[29142]_  = \new_[29141]_  & \new_[29138]_ ;
  assign \new_[29143]_  = \new_[29142]_  & \new_[29135]_ ;
  assign \new_[29147]_  = A233 & ~A232;
  assign \new_[29148]_  = ~A203 & \new_[29147]_ ;
  assign \new_[29151]_  = A236 & ~A235;
  assign \new_[29154]_  = A300 & A299;
  assign \new_[29155]_  = \new_[29154]_  & \new_[29151]_ ;
  assign \new_[29156]_  = \new_[29155]_  & \new_[29148]_ ;
  assign \new_[29160]_  = ~A167 & A168;
  assign \new_[29161]_  = A170 & \new_[29160]_ ;
  assign \new_[29164]_  = A199 & A166;
  assign \new_[29167]_  = ~A201 & ~A200;
  assign \new_[29168]_  = \new_[29167]_  & \new_[29164]_ ;
  assign \new_[29169]_  = \new_[29168]_  & \new_[29161]_ ;
  assign \new_[29173]_  = A233 & ~A232;
  assign \new_[29174]_  = ~A203 & \new_[29173]_ ;
  assign \new_[29177]_  = A236 & ~A235;
  assign \new_[29180]_  = A300 & A298;
  assign \new_[29181]_  = \new_[29180]_  & \new_[29177]_ ;
  assign \new_[29182]_  = \new_[29181]_  & \new_[29174]_ ;
  assign \new_[29186]_  = ~A167 & A168;
  assign \new_[29187]_  = A170 & \new_[29186]_ ;
  assign \new_[29190]_  = A199 & A166;
  assign \new_[29193]_  = ~A201 & ~A200;
  assign \new_[29194]_  = \new_[29193]_  & \new_[29190]_ ;
  assign \new_[29195]_  = \new_[29194]_  & \new_[29187]_ ;
  assign \new_[29199]_  = A233 & ~A232;
  assign \new_[29200]_  = ~A203 & \new_[29199]_ ;
  assign \new_[29203]_  = A236 & ~A235;
  assign \new_[29206]_  = A267 & A265;
  assign \new_[29207]_  = \new_[29206]_  & \new_[29203]_ ;
  assign \new_[29208]_  = \new_[29207]_  & \new_[29200]_ ;
  assign \new_[29212]_  = ~A167 & A168;
  assign \new_[29213]_  = A170 & \new_[29212]_ ;
  assign \new_[29216]_  = A199 & A166;
  assign \new_[29219]_  = ~A201 & ~A200;
  assign \new_[29220]_  = \new_[29219]_  & \new_[29216]_ ;
  assign \new_[29221]_  = \new_[29220]_  & \new_[29213]_ ;
  assign \new_[29225]_  = A233 & ~A232;
  assign \new_[29226]_  = ~A203 & \new_[29225]_ ;
  assign \new_[29229]_  = A236 & ~A235;
  assign \new_[29232]_  = A267 & A266;
  assign \new_[29233]_  = \new_[29232]_  & \new_[29229]_ ;
  assign \new_[29234]_  = \new_[29233]_  & \new_[29226]_ ;
  assign \new_[29238]_  = ~A167 & A168;
  assign \new_[29239]_  = A170 & \new_[29238]_ ;
  assign \new_[29242]_  = A199 & A166;
  assign \new_[29245]_  = ~A201 & ~A200;
  assign \new_[29246]_  = \new_[29245]_  & \new_[29242]_ ;
  assign \new_[29247]_  = \new_[29246]_  & \new_[29239]_ ;
  assign \new_[29251]_  = ~A233 & A232;
  assign \new_[29252]_  = ~A203 & \new_[29251]_ ;
  assign \new_[29255]_  = A236 & ~A235;
  assign \new_[29258]_  = A300 & A299;
  assign \new_[29259]_  = \new_[29258]_  & \new_[29255]_ ;
  assign \new_[29260]_  = \new_[29259]_  & \new_[29252]_ ;
  assign \new_[29264]_  = ~A167 & A168;
  assign \new_[29265]_  = A170 & \new_[29264]_ ;
  assign \new_[29268]_  = A199 & A166;
  assign \new_[29271]_  = ~A201 & ~A200;
  assign \new_[29272]_  = \new_[29271]_  & \new_[29268]_ ;
  assign \new_[29273]_  = \new_[29272]_  & \new_[29265]_ ;
  assign \new_[29277]_  = ~A233 & A232;
  assign \new_[29278]_  = ~A203 & \new_[29277]_ ;
  assign \new_[29281]_  = A236 & ~A235;
  assign \new_[29284]_  = A300 & A298;
  assign \new_[29285]_  = \new_[29284]_  & \new_[29281]_ ;
  assign \new_[29286]_  = \new_[29285]_  & \new_[29278]_ ;
  assign \new_[29290]_  = ~A167 & A168;
  assign \new_[29291]_  = A170 & \new_[29290]_ ;
  assign \new_[29294]_  = A199 & A166;
  assign \new_[29297]_  = ~A201 & ~A200;
  assign \new_[29298]_  = \new_[29297]_  & \new_[29294]_ ;
  assign \new_[29299]_  = \new_[29298]_  & \new_[29291]_ ;
  assign \new_[29303]_  = ~A233 & A232;
  assign \new_[29304]_  = ~A203 & \new_[29303]_ ;
  assign \new_[29307]_  = A236 & ~A235;
  assign \new_[29310]_  = A267 & A265;
  assign \new_[29311]_  = \new_[29310]_  & \new_[29307]_ ;
  assign \new_[29312]_  = \new_[29311]_  & \new_[29304]_ ;
  assign \new_[29316]_  = ~A167 & A168;
  assign \new_[29317]_  = A170 & \new_[29316]_ ;
  assign \new_[29320]_  = A199 & A166;
  assign \new_[29323]_  = ~A201 & ~A200;
  assign \new_[29324]_  = \new_[29323]_  & \new_[29320]_ ;
  assign \new_[29325]_  = \new_[29324]_  & \new_[29317]_ ;
  assign \new_[29329]_  = ~A233 & A232;
  assign \new_[29330]_  = ~A203 & \new_[29329]_ ;
  assign \new_[29333]_  = A236 & ~A235;
  assign \new_[29336]_  = A267 & A266;
  assign \new_[29337]_  = \new_[29336]_  & \new_[29333]_ ;
  assign \new_[29338]_  = \new_[29337]_  & \new_[29330]_ ;
  assign \new_[29342]_  = ~A167 & A168;
  assign \new_[29343]_  = A170 & \new_[29342]_ ;
  assign \new_[29346]_  = A199 & A166;
  assign \new_[29349]_  = ~A201 & ~A200;
  assign \new_[29350]_  = \new_[29349]_  & \new_[29346]_ ;
  assign \new_[29351]_  = \new_[29350]_  & \new_[29343]_ ;
  assign \new_[29355]_  = ~A233 & ~A232;
  assign \new_[29356]_  = ~A203 & \new_[29355]_ ;
  assign \new_[29359]_  = ~A236 & A235;
  assign \new_[29362]_  = A300 & A299;
  assign \new_[29363]_  = \new_[29362]_  & \new_[29359]_ ;
  assign \new_[29364]_  = \new_[29363]_  & \new_[29356]_ ;
  assign \new_[29368]_  = ~A167 & A168;
  assign \new_[29369]_  = A170 & \new_[29368]_ ;
  assign \new_[29372]_  = A199 & A166;
  assign \new_[29375]_  = ~A201 & ~A200;
  assign \new_[29376]_  = \new_[29375]_  & \new_[29372]_ ;
  assign \new_[29377]_  = \new_[29376]_  & \new_[29369]_ ;
  assign \new_[29381]_  = ~A233 & ~A232;
  assign \new_[29382]_  = ~A203 & \new_[29381]_ ;
  assign \new_[29385]_  = ~A236 & A235;
  assign \new_[29388]_  = A300 & A298;
  assign \new_[29389]_  = \new_[29388]_  & \new_[29385]_ ;
  assign \new_[29390]_  = \new_[29389]_  & \new_[29382]_ ;
  assign \new_[29394]_  = ~A167 & A168;
  assign \new_[29395]_  = A170 & \new_[29394]_ ;
  assign \new_[29398]_  = A199 & A166;
  assign \new_[29401]_  = ~A201 & ~A200;
  assign \new_[29402]_  = \new_[29401]_  & \new_[29398]_ ;
  assign \new_[29403]_  = \new_[29402]_  & \new_[29395]_ ;
  assign \new_[29407]_  = ~A233 & ~A232;
  assign \new_[29408]_  = ~A203 & \new_[29407]_ ;
  assign \new_[29411]_  = ~A236 & A235;
  assign \new_[29414]_  = A267 & A265;
  assign \new_[29415]_  = \new_[29414]_  & \new_[29411]_ ;
  assign \new_[29416]_  = \new_[29415]_  & \new_[29408]_ ;
  assign \new_[29420]_  = ~A167 & A168;
  assign \new_[29421]_  = A170 & \new_[29420]_ ;
  assign \new_[29424]_  = A199 & A166;
  assign \new_[29427]_  = ~A201 & ~A200;
  assign \new_[29428]_  = \new_[29427]_  & \new_[29424]_ ;
  assign \new_[29429]_  = \new_[29428]_  & \new_[29421]_ ;
  assign \new_[29433]_  = ~A233 & ~A232;
  assign \new_[29434]_  = ~A203 & \new_[29433]_ ;
  assign \new_[29437]_  = ~A236 & A235;
  assign \new_[29440]_  = A267 & A266;
  assign \new_[29441]_  = \new_[29440]_  & \new_[29437]_ ;
  assign \new_[29442]_  = \new_[29441]_  & \new_[29434]_ ;
  assign \new_[29446]_  = ~A167 & A168;
  assign \new_[29447]_  = A169 & \new_[29446]_ ;
  assign \new_[29450]_  = A199 & A166;
  assign \new_[29453]_  = ~A201 & A200;
  assign \new_[29454]_  = \new_[29453]_  & \new_[29450]_ ;
  assign \new_[29455]_  = \new_[29454]_  & \new_[29447]_ ;
  assign \new_[29459]_  = A234 & A232;
  assign \new_[29460]_  = ~A202 & \new_[29459]_ ;
  assign \new_[29463]_  = A299 & A298;
  assign \new_[29466]_  = ~A302 & A301;
  assign \new_[29467]_  = \new_[29466]_  & \new_[29463]_ ;
  assign \new_[29468]_  = \new_[29467]_  & \new_[29460]_ ;
  assign \new_[29472]_  = ~A167 & A168;
  assign \new_[29473]_  = A169 & \new_[29472]_ ;
  assign \new_[29476]_  = A199 & A166;
  assign \new_[29479]_  = ~A201 & A200;
  assign \new_[29480]_  = \new_[29479]_  & \new_[29476]_ ;
  assign \new_[29481]_  = \new_[29480]_  & \new_[29473]_ ;
  assign \new_[29485]_  = A234 & A232;
  assign \new_[29486]_  = ~A202 & \new_[29485]_ ;
  assign \new_[29489]_  = ~A299 & A298;
  assign \new_[29492]_  = A302 & ~A301;
  assign \new_[29493]_  = \new_[29492]_  & \new_[29489]_ ;
  assign \new_[29494]_  = \new_[29493]_  & \new_[29486]_ ;
  assign \new_[29498]_  = ~A167 & A168;
  assign \new_[29499]_  = A169 & \new_[29498]_ ;
  assign \new_[29502]_  = A199 & A166;
  assign \new_[29505]_  = ~A201 & A200;
  assign \new_[29506]_  = \new_[29505]_  & \new_[29502]_ ;
  assign \new_[29507]_  = \new_[29506]_  & \new_[29499]_ ;
  assign \new_[29511]_  = A234 & A232;
  assign \new_[29512]_  = ~A202 & \new_[29511]_ ;
  assign \new_[29515]_  = A299 & ~A298;
  assign \new_[29518]_  = A302 & ~A301;
  assign \new_[29519]_  = \new_[29518]_  & \new_[29515]_ ;
  assign \new_[29520]_  = \new_[29519]_  & \new_[29512]_ ;
  assign \new_[29524]_  = ~A167 & A168;
  assign \new_[29525]_  = A169 & \new_[29524]_ ;
  assign \new_[29528]_  = A199 & A166;
  assign \new_[29531]_  = ~A201 & A200;
  assign \new_[29532]_  = \new_[29531]_  & \new_[29528]_ ;
  assign \new_[29533]_  = \new_[29532]_  & \new_[29525]_ ;
  assign \new_[29537]_  = A234 & A232;
  assign \new_[29538]_  = ~A202 & \new_[29537]_ ;
  assign \new_[29541]_  = ~A299 & ~A298;
  assign \new_[29544]_  = ~A302 & A301;
  assign \new_[29545]_  = \new_[29544]_  & \new_[29541]_ ;
  assign \new_[29546]_  = \new_[29545]_  & \new_[29538]_ ;
  assign \new_[29550]_  = ~A167 & A168;
  assign \new_[29551]_  = A169 & \new_[29550]_ ;
  assign \new_[29554]_  = A199 & A166;
  assign \new_[29557]_  = ~A201 & A200;
  assign \new_[29558]_  = \new_[29557]_  & \new_[29554]_ ;
  assign \new_[29559]_  = \new_[29558]_  & \new_[29551]_ ;
  assign \new_[29563]_  = A234 & A232;
  assign \new_[29564]_  = ~A202 & \new_[29563]_ ;
  assign \new_[29567]_  = A266 & A265;
  assign \new_[29570]_  = ~A269 & A268;
  assign \new_[29571]_  = \new_[29570]_  & \new_[29567]_ ;
  assign \new_[29572]_  = \new_[29571]_  & \new_[29564]_ ;
  assign \new_[29576]_  = ~A167 & A168;
  assign \new_[29577]_  = A169 & \new_[29576]_ ;
  assign \new_[29580]_  = A199 & A166;
  assign \new_[29583]_  = ~A201 & A200;
  assign \new_[29584]_  = \new_[29583]_  & \new_[29580]_ ;
  assign \new_[29585]_  = \new_[29584]_  & \new_[29577]_ ;
  assign \new_[29589]_  = A234 & A232;
  assign \new_[29590]_  = ~A202 & \new_[29589]_ ;
  assign \new_[29593]_  = A266 & ~A265;
  assign \new_[29596]_  = A269 & ~A268;
  assign \new_[29597]_  = \new_[29596]_  & \new_[29593]_ ;
  assign \new_[29598]_  = \new_[29597]_  & \new_[29590]_ ;
  assign \new_[29602]_  = ~A167 & A168;
  assign \new_[29603]_  = A169 & \new_[29602]_ ;
  assign \new_[29606]_  = A199 & A166;
  assign \new_[29609]_  = ~A201 & A200;
  assign \new_[29610]_  = \new_[29609]_  & \new_[29606]_ ;
  assign \new_[29611]_  = \new_[29610]_  & \new_[29603]_ ;
  assign \new_[29615]_  = A234 & A232;
  assign \new_[29616]_  = ~A202 & \new_[29615]_ ;
  assign \new_[29619]_  = ~A266 & A265;
  assign \new_[29622]_  = A269 & ~A268;
  assign \new_[29623]_  = \new_[29622]_  & \new_[29619]_ ;
  assign \new_[29624]_  = \new_[29623]_  & \new_[29616]_ ;
  assign \new_[29628]_  = ~A167 & A168;
  assign \new_[29629]_  = A169 & \new_[29628]_ ;
  assign \new_[29632]_  = A199 & A166;
  assign \new_[29635]_  = ~A201 & A200;
  assign \new_[29636]_  = \new_[29635]_  & \new_[29632]_ ;
  assign \new_[29637]_  = \new_[29636]_  & \new_[29629]_ ;
  assign \new_[29641]_  = A234 & A232;
  assign \new_[29642]_  = ~A202 & \new_[29641]_ ;
  assign \new_[29645]_  = ~A266 & ~A265;
  assign \new_[29648]_  = ~A269 & A268;
  assign \new_[29649]_  = \new_[29648]_  & \new_[29645]_ ;
  assign \new_[29650]_  = \new_[29649]_  & \new_[29642]_ ;
  assign \new_[29654]_  = ~A167 & A168;
  assign \new_[29655]_  = A169 & \new_[29654]_ ;
  assign \new_[29658]_  = A199 & A166;
  assign \new_[29661]_  = ~A201 & A200;
  assign \new_[29662]_  = \new_[29661]_  & \new_[29658]_ ;
  assign \new_[29663]_  = \new_[29662]_  & \new_[29655]_ ;
  assign \new_[29667]_  = A234 & A233;
  assign \new_[29668]_  = ~A202 & \new_[29667]_ ;
  assign \new_[29671]_  = A299 & A298;
  assign \new_[29674]_  = ~A302 & A301;
  assign \new_[29675]_  = \new_[29674]_  & \new_[29671]_ ;
  assign \new_[29676]_  = \new_[29675]_  & \new_[29668]_ ;
  assign \new_[29680]_  = ~A167 & A168;
  assign \new_[29681]_  = A169 & \new_[29680]_ ;
  assign \new_[29684]_  = A199 & A166;
  assign \new_[29687]_  = ~A201 & A200;
  assign \new_[29688]_  = \new_[29687]_  & \new_[29684]_ ;
  assign \new_[29689]_  = \new_[29688]_  & \new_[29681]_ ;
  assign \new_[29693]_  = A234 & A233;
  assign \new_[29694]_  = ~A202 & \new_[29693]_ ;
  assign \new_[29697]_  = ~A299 & A298;
  assign \new_[29700]_  = A302 & ~A301;
  assign \new_[29701]_  = \new_[29700]_  & \new_[29697]_ ;
  assign \new_[29702]_  = \new_[29701]_  & \new_[29694]_ ;
  assign \new_[29706]_  = ~A167 & A168;
  assign \new_[29707]_  = A169 & \new_[29706]_ ;
  assign \new_[29710]_  = A199 & A166;
  assign \new_[29713]_  = ~A201 & A200;
  assign \new_[29714]_  = \new_[29713]_  & \new_[29710]_ ;
  assign \new_[29715]_  = \new_[29714]_  & \new_[29707]_ ;
  assign \new_[29719]_  = A234 & A233;
  assign \new_[29720]_  = ~A202 & \new_[29719]_ ;
  assign \new_[29723]_  = A299 & ~A298;
  assign \new_[29726]_  = A302 & ~A301;
  assign \new_[29727]_  = \new_[29726]_  & \new_[29723]_ ;
  assign \new_[29728]_  = \new_[29727]_  & \new_[29720]_ ;
  assign \new_[29732]_  = ~A167 & A168;
  assign \new_[29733]_  = A169 & \new_[29732]_ ;
  assign \new_[29736]_  = A199 & A166;
  assign \new_[29739]_  = ~A201 & A200;
  assign \new_[29740]_  = \new_[29739]_  & \new_[29736]_ ;
  assign \new_[29741]_  = \new_[29740]_  & \new_[29733]_ ;
  assign \new_[29745]_  = A234 & A233;
  assign \new_[29746]_  = ~A202 & \new_[29745]_ ;
  assign \new_[29749]_  = ~A299 & ~A298;
  assign \new_[29752]_  = ~A302 & A301;
  assign \new_[29753]_  = \new_[29752]_  & \new_[29749]_ ;
  assign \new_[29754]_  = \new_[29753]_  & \new_[29746]_ ;
  assign \new_[29758]_  = ~A167 & A168;
  assign \new_[29759]_  = A169 & \new_[29758]_ ;
  assign \new_[29762]_  = A199 & A166;
  assign \new_[29765]_  = ~A201 & A200;
  assign \new_[29766]_  = \new_[29765]_  & \new_[29762]_ ;
  assign \new_[29767]_  = \new_[29766]_  & \new_[29759]_ ;
  assign \new_[29771]_  = A234 & A233;
  assign \new_[29772]_  = ~A202 & \new_[29771]_ ;
  assign \new_[29775]_  = A266 & A265;
  assign \new_[29778]_  = ~A269 & A268;
  assign \new_[29779]_  = \new_[29778]_  & \new_[29775]_ ;
  assign \new_[29780]_  = \new_[29779]_  & \new_[29772]_ ;
  assign \new_[29784]_  = ~A167 & A168;
  assign \new_[29785]_  = A169 & \new_[29784]_ ;
  assign \new_[29788]_  = A199 & A166;
  assign \new_[29791]_  = ~A201 & A200;
  assign \new_[29792]_  = \new_[29791]_  & \new_[29788]_ ;
  assign \new_[29793]_  = \new_[29792]_  & \new_[29785]_ ;
  assign \new_[29797]_  = A234 & A233;
  assign \new_[29798]_  = ~A202 & \new_[29797]_ ;
  assign \new_[29801]_  = A266 & ~A265;
  assign \new_[29804]_  = A269 & ~A268;
  assign \new_[29805]_  = \new_[29804]_  & \new_[29801]_ ;
  assign \new_[29806]_  = \new_[29805]_  & \new_[29798]_ ;
  assign \new_[29810]_  = ~A167 & A168;
  assign \new_[29811]_  = A169 & \new_[29810]_ ;
  assign \new_[29814]_  = A199 & A166;
  assign \new_[29817]_  = ~A201 & A200;
  assign \new_[29818]_  = \new_[29817]_  & \new_[29814]_ ;
  assign \new_[29819]_  = \new_[29818]_  & \new_[29811]_ ;
  assign \new_[29823]_  = A234 & A233;
  assign \new_[29824]_  = ~A202 & \new_[29823]_ ;
  assign \new_[29827]_  = ~A266 & A265;
  assign \new_[29830]_  = A269 & ~A268;
  assign \new_[29831]_  = \new_[29830]_  & \new_[29827]_ ;
  assign \new_[29832]_  = \new_[29831]_  & \new_[29824]_ ;
  assign \new_[29836]_  = ~A167 & A168;
  assign \new_[29837]_  = A169 & \new_[29836]_ ;
  assign \new_[29840]_  = A199 & A166;
  assign \new_[29843]_  = ~A201 & A200;
  assign \new_[29844]_  = \new_[29843]_  & \new_[29840]_ ;
  assign \new_[29845]_  = \new_[29844]_  & \new_[29837]_ ;
  assign \new_[29849]_  = A234 & A233;
  assign \new_[29850]_  = ~A202 & \new_[29849]_ ;
  assign \new_[29853]_  = ~A266 & ~A265;
  assign \new_[29856]_  = ~A269 & A268;
  assign \new_[29857]_  = \new_[29856]_  & \new_[29853]_ ;
  assign \new_[29858]_  = \new_[29857]_  & \new_[29850]_ ;
  assign \new_[29862]_  = ~A167 & A168;
  assign \new_[29863]_  = A169 & \new_[29862]_ ;
  assign \new_[29866]_  = A199 & A166;
  assign \new_[29869]_  = ~A201 & A200;
  assign \new_[29870]_  = \new_[29869]_  & \new_[29866]_ ;
  assign \new_[29871]_  = \new_[29870]_  & \new_[29863]_ ;
  assign \new_[29875]_  = A233 & A232;
  assign \new_[29876]_  = ~A202 & \new_[29875]_ ;
  assign \new_[29879]_  = ~A236 & A235;
  assign \new_[29882]_  = A300 & A299;
  assign \new_[29883]_  = \new_[29882]_  & \new_[29879]_ ;
  assign \new_[29884]_  = \new_[29883]_  & \new_[29876]_ ;
  assign \new_[29888]_  = ~A167 & A168;
  assign \new_[29889]_  = A169 & \new_[29888]_ ;
  assign \new_[29892]_  = A199 & A166;
  assign \new_[29895]_  = ~A201 & A200;
  assign \new_[29896]_  = \new_[29895]_  & \new_[29892]_ ;
  assign \new_[29897]_  = \new_[29896]_  & \new_[29889]_ ;
  assign \new_[29901]_  = A233 & A232;
  assign \new_[29902]_  = ~A202 & \new_[29901]_ ;
  assign \new_[29905]_  = ~A236 & A235;
  assign \new_[29908]_  = A300 & A298;
  assign \new_[29909]_  = \new_[29908]_  & \new_[29905]_ ;
  assign \new_[29910]_  = \new_[29909]_  & \new_[29902]_ ;
  assign \new_[29914]_  = ~A167 & A168;
  assign \new_[29915]_  = A169 & \new_[29914]_ ;
  assign \new_[29918]_  = A199 & A166;
  assign \new_[29921]_  = ~A201 & A200;
  assign \new_[29922]_  = \new_[29921]_  & \new_[29918]_ ;
  assign \new_[29923]_  = \new_[29922]_  & \new_[29915]_ ;
  assign \new_[29927]_  = A233 & A232;
  assign \new_[29928]_  = ~A202 & \new_[29927]_ ;
  assign \new_[29931]_  = ~A236 & A235;
  assign \new_[29934]_  = A267 & A265;
  assign \new_[29935]_  = \new_[29934]_  & \new_[29931]_ ;
  assign \new_[29936]_  = \new_[29935]_  & \new_[29928]_ ;
  assign \new_[29940]_  = ~A167 & A168;
  assign \new_[29941]_  = A169 & \new_[29940]_ ;
  assign \new_[29944]_  = A199 & A166;
  assign \new_[29947]_  = ~A201 & A200;
  assign \new_[29948]_  = \new_[29947]_  & \new_[29944]_ ;
  assign \new_[29949]_  = \new_[29948]_  & \new_[29941]_ ;
  assign \new_[29953]_  = A233 & A232;
  assign \new_[29954]_  = ~A202 & \new_[29953]_ ;
  assign \new_[29957]_  = ~A236 & A235;
  assign \new_[29960]_  = A267 & A266;
  assign \new_[29961]_  = \new_[29960]_  & \new_[29957]_ ;
  assign \new_[29962]_  = \new_[29961]_  & \new_[29954]_ ;
  assign \new_[29966]_  = ~A167 & A168;
  assign \new_[29967]_  = A169 & \new_[29966]_ ;
  assign \new_[29970]_  = A199 & A166;
  assign \new_[29973]_  = ~A201 & A200;
  assign \new_[29974]_  = \new_[29973]_  & \new_[29970]_ ;
  assign \new_[29975]_  = \new_[29974]_  & \new_[29967]_ ;
  assign \new_[29979]_  = A233 & ~A232;
  assign \new_[29980]_  = ~A202 & \new_[29979]_ ;
  assign \new_[29983]_  = A236 & ~A235;
  assign \new_[29986]_  = A300 & A299;
  assign \new_[29987]_  = \new_[29986]_  & \new_[29983]_ ;
  assign \new_[29988]_  = \new_[29987]_  & \new_[29980]_ ;
  assign \new_[29992]_  = ~A167 & A168;
  assign \new_[29993]_  = A169 & \new_[29992]_ ;
  assign \new_[29996]_  = A199 & A166;
  assign \new_[29999]_  = ~A201 & A200;
  assign \new_[30000]_  = \new_[29999]_  & \new_[29996]_ ;
  assign \new_[30001]_  = \new_[30000]_  & \new_[29993]_ ;
  assign \new_[30005]_  = A233 & ~A232;
  assign \new_[30006]_  = ~A202 & \new_[30005]_ ;
  assign \new_[30009]_  = A236 & ~A235;
  assign \new_[30012]_  = A300 & A298;
  assign \new_[30013]_  = \new_[30012]_  & \new_[30009]_ ;
  assign \new_[30014]_  = \new_[30013]_  & \new_[30006]_ ;
  assign \new_[30018]_  = ~A167 & A168;
  assign \new_[30019]_  = A169 & \new_[30018]_ ;
  assign \new_[30022]_  = A199 & A166;
  assign \new_[30025]_  = ~A201 & A200;
  assign \new_[30026]_  = \new_[30025]_  & \new_[30022]_ ;
  assign \new_[30027]_  = \new_[30026]_  & \new_[30019]_ ;
  assign \new_[30031]_  = A233 & ~A232;
  assign \new_[30032]_  = ~A202 & \new_[30031]_ ;
  assign \new_[30035]_  = A236 & ~A235;
  assign \new_[30038]_  = A267 & A265;
  assign \new_[30039]_  = \new_[30038]_  & \new_[30035]_ ;
  assign \new_[30040]_  = \new_[30039]_  & \new_[30032]_ ;
  assign \new_[30044]_  = ~A167 & A168;
  assign \new_[30045]_  = A169 & \new_[30044]_ ;
  assign \new_[30048]_  = A199 & A166;
  assign \new_[30051]_  = ~A201 & A200;
  assign \new_[30052]_  = \new_[30051]_  & \new_[30048]_ ;
  assign \new_[30053]_  = \new_[30052]_  & \new_[30045]_ ;
  assign \new_[30057]_  = A233 & ~A232;
  assign \new_[30058]_  = ~A202 & \new_[30057]_ ;
  assign \new_[30061]_  = A236 & ~A235;
  assign \new_[30064]_  = A267 & A266;
  assign \new_[30065]_  = \new_[30064]_  & \new_[30061]_ ;
  assign \new_[30066]_  = \new_[30065]_  & \new_[30058]_ ;
  assign \new_[30070]_  = ~A167 & A168;
  assign \new_[30071]_  = A169 & \new_[30070]_ ;
  assign \new_[30074]_  = A199 & A166;
  assign \new_[30077]_  = ~A201 & A200;
  assign \new_[30078]_  = \new_[30077]_  & \new_[30074]_ ;
  assign \new_[30079]_  = \new_[30078]_  & \new_[30071]_ ;
  assign \new_[30083]_  = ~A233 & A232;
  assign \new_[30084]_  = ~A202 & \new_[30083]_ ;
  assign \new_[30087]_  = A236 & ~A235;
  assign \new_[30090]_  = A300 & A299;
  assign \new_[30091]_  = \new_[30090]_  & \new_[30087]_ ;
  assign \new_[30092]_  = \new_[30091]_  & \new_[30084]_ ;
  assign \new_[30096]_  = ~A167 & A168;
  assign \new_[30097]_  = A169 & \new_[30096]_ ;
  assign \new_[30100]_  = A199 & A166;
  assign \new_[30103]_  = ~A201 & A200;
  assign \new_[30104]_  = \new_[30103]_  & \new_[30100]_ ;
  assign \new_[30105]_  = \new_[30104]_  & \new_[30097]_ ;
  assign \new_[30109]_  = ~A233 & A232;
  assign \new_[30110]_  = ~A202 & \new_[30109]_ ;
  assign \new_[30113]_  = A236 & ~A235;
  assign \new_[30116]_  = A300 & A298;
  assign \new_[30117]_  = \new_[30116]_  & \new_[30113]_ ;
  assign \new_[30118]_  = \new_[30117]_  & \new_[30110]_ ;
  assign \new_[30122]_  = ~A167 & A168;
  assign \new_[30123]_  = A169 & \new_[30122]_ ;
  assign \new_[30126]_  = A199 & A166;
  assign \new_[30129]_  = ~A201 & A200;
  assign \new_[30130]_  = \new_[30129]_  & \new_[30126]_ ;
  assign \new_[30131]_  = \new_[30130]_  & \new_[30123]_ ;
  assign \new_[30135]_  = ~A233 & A232;
  assign \new_[30136]_  = ~A202 & \new_[30135]_ ;
  assign \new_[30139]_  = A236 & ~A235;
  assign \new_[30142]_  = A267 & A265;
  assign \new_[30143]_  = \new_[30142]_  & \new_[30139]_ ;
  assign \new_[30144]_  = \new_[30143]_  & \new_[30136]_ ;
  assign \new_[30148]_  = ~A167 & A168;
  assign \new_[30149]_  = A169 & \new_[30148]_ ;
  assign \new_[30152]_  = A199 & A166;
  assign \new_[30155]_  = ~A201 & A200;
  assign \new_[30156]_  = \new_[30155]_  & \new_[30152]_ ;
  assign \new_[30157]_  = \new_[30156]_  & \new_[30149]_ ;
  assign \new_[30161]_  = ~A233 & A232;
  assign \new_[30162]_  = ~A202 & \new_[30161]_ ;
  assign \new_[30165]_  = A236 & ~A235;
  assign \new_[30168]_  = A267 & A266;
  assign \new_[30169]_  = \new_[30168]_  & \new_[30165]_ ;
  assign \new_[30170]_  = \new_[30169]_  & \new_[30162]_ ;
  assign \new_[30174]_  = ~A167 & A168;
  assign \new_[30175]_  = A169 & \new_[30174]_ ;
  assign \new_[30178]_  = A199 & A166;
  assign \new_[30181]_  = ~A201 & A200;
  assign \new_[30182]_  = \new_[30181]_  & \new_[30178]_ ;
  assign \new_[30183]_  = \new_[30182]_  & \new_[30175]_ ;
  assign \new_[30187]_  = ~A233 & ~A232;
  assign \new_[30188]_  = ~A202 & \new_[30187]_ ;
  assign \new_[30191]_  = ~A236 & A235;
  assign \new_[30194]_  = A300 & A299;
  assign \new_[30195]_  = \new_[30194]_  & \new_[30191]_ ;
  assign \new_[30196]_  = \new_[30195]_  & \new_[30188]_ ;
  assign \new_[30200]_  = ~A167 & A168;
  assign \new_[30201]_  = A169 & \new_[30200]_ ;
  assign \new_[30204]_  = A199 & A166;
  assign \new_[30207]_  = ~A201 & A200;
  assign \new_[30208]_  = \new_[30207]_  & \new_[30204]_ ;
  assign \new_[30209]_  = \new_[30208]_  & \new_[30201]_ ;
  assign \new_[30213]_  = ~A233 & ~A232;
  assign \new_[30214]_  = ~A202 & \new_[30213]_ ;
  assign \new_[30217]_  = ~A236 & A235;
  assign \new_[30220]_  = A300 & A298;
  assign \new_[30221]_  = \new_[30220]_  & \new_[30217]_ ;
  assign \new_[30222]_  = \new_[30221]_  & \new_[30214]_ ;
  assign \new_[30226]_  = ~A167 & A168;
  assign \new_[30227]_  = A169 & \new_[30226]_ ;
  assign \new_[30230]_  = A199 & A166;
  assign \new_[30233]_  = ~A201 & A200;
  assign \new_[30234]_  = \new_[30233]_  & \new_[30230]_ ;
  assign \new_[30235]_  = \new_[30234]_  & \new_[30227]_ ;
  assign \new_[30239]_  = ~A233 & ~A232;
  assign \new_[30240]_  = ~A202 & \new_[30239]_ ;
  assign \new_[30243]_  = ~A236 & A235;
  assign \new_[30246]_  = A267 & A265;
  assign \new_[30247]_  = \new_[30246]_  & \new_[30243]_ ;
  assign \new_[30248]_  = \new_[30247]_  & \new_[30240]_ ;
  assign \new_[30252]_  = ~A167 & A168;
  assign \new_[30253]_  = A169 & \new_[30252]_ ;
  assign \new_[30256]_  = A199 & A166;
  assign \new_[30259]_  = ~A201 & A200;
  assign \new_[30260]_  = \new_[30259]_  & \new_[30256]_ ;
  assign \new_[30261]_  = \new_[30260]_  & \new_[30253]_ ;
  assign \new_[30265]_  = ~A233 & ~A232;
  assign \new_[30266]_  = ~A202 & \new_[30265]_ ;
  assign \new_[30269]_  = ~A236 & A235;
  assign \new_[30272]_  = A267 & A266;
  assign \new_[30273]_  = \new_[30272]_  & \new_[30269]_ ;
  assign \new_[30274]_  = \new_[30273]_  & \new_[30266]_ ;
  assign \new_[30278]_  = ~A167 & A168;
  assign \new_[30279]_  = A169 & \new_[30278]_ ;
  assign \new_[30282]_  = A199 & A166;
  assign \new_[30285]_  = ~A201 & A200;
  assign \new_[30286]_  = \new_[30285]_  & \new_[30282]_ ;
  assign \new_[30287]_  = \new_[30286]_  & \new_[30279]_ ;
  assign \new_[30291]_  = A234 & A232;
  assign \new_[30292]_  = A203 & \new_[30291]_ ;
  assign \new_[30295]_  = A299 & A298;
  assign \new_[30298]_  = ~A302 & A301;
  assign \new_[30299]_  = \new_[30298]_  & \new_[30295]_ ;
  assign \new_[30300]_  = \new_[30299]_  & \new_[30292]_ ;
  assign \new_[30304]_  = ~A167 & A168;
  assign \new_[30305]_  = A169 & \new_[30304]_ ;
  assign \new_[30308]_  = A199 & A166;
  assign \new_[30311]_  = ~A201 & A200;
  assign \new_[30312]_  = \new_[30311]_  & \new_[30308]_ ;
  assign \new_[30313]_  = \new_[30312]_  & \new_[30305]_ ;
  assign \new_[30317]_  = A234 & A232;
  assign \new_[30318]_  = A203 & \new_[30317]_ ;
  assign \new_[30321]_  = ~A299 & A298;
  assign \new_[30324]_  = A302 & ~A301;
  assign \new_[30325]_  = \new_[30324]_  & \new_[30321]_ ;
  assign \new_[30326]_  = \new_[30325]_  & \new_[30318]_ ;
  assign \new_[30330]_  = ~A167 & A168;
  assign \new_[30331]_  = A169 & \new_[30330]_ ;
  assign \new_[30334]_  = A199 & A166;
  assign \new_[30337]_  = ~A201 & A200;
  assign \new_[30338]_  = \new_[30337]_  & \new_[30334]_ ;
  assign \new_[30339]_  = \new_[30338]_  & \new_[30331]_ ;
  assign \new_[30343]_  = A234 & A232;
  assign \new_[30344]_  = A203 & \new_[30343]_ ;
  assign \new_[30347]_  = A299 & ~A298;
  assign \new_[30350]_  = A302 & ~A301;
  assign \new_[30351]_  = \new_[30350]_  & \new_[30347]_ ;
  assign \new_[30352]_  = \new_[30351]_  & \new_[30344]_ ;
  assign \new_[30356]_  = ~A167 & A168;
  assign \new_[30357]_  = A169 & \new_[30356]_ ;
  assign \new_[30360]_  = A199 & A166;
  assign \new_[30363]_  = ~A201 & A200;
  assign \new_[30364]_  = \new_[30363]_  & \new_[30360]_ ;
  assign \new_[30365]_  = \new_[30364]_  & \new_[30357]_ ;
  assign \new_[30369]_  = A234 & A232;
  assign \new_[30370]_  = A203 & \new_[30369]_ ;
  assign \new_[30373]_  = ~A299 & ~A298;
  assign \new_[30376]_  = ~A302 & A301;
  assign \new_[30377]_  = \new_[30376]_  & \new_[30373]_ ;
  assign \new_[30378]_  = \new_[30377]_  & \new_[30370]_ ;
  assign \new_[30382]_  = ~A167 & A168;
  assign \new_[30383]_  = A169 & \new_[30382]_ ;
  assign \new_[30386]_  = A199 & A166;
  assign \new_[30389]_  = ~A201 & A200;
  assign \new_[30390]_  = \new_[30389]_  & \new_[30386]_ ;
  assign \new_[30391]_  = \new_[30390]_  & \new_[30383]_ ;
  assign \new_[30395]_  = A234 & A232;
  assign \new_[30396]_  = A203 & \new_[30395]_ ;
  assign \new_[30399]_  = A266 & A265;
  assign \new_[30402]_  = ~A269 & A268;
  assign \new_[30403]_  = \new_[30402]_  & \new_[30399]_ ;
  assign \new_[30404]_  = \new_[30403]_  & \new_[30396]_ ;
  assign \new_[30408]_  = ~A167 & A168;
  assign \new_[30409]_  = A169 & \new_[30408]_ ;
  assign \new_[30412]_  = A199 & A166;
  assign \new_[30415]_  = ~A201 & A200;
  assign \new_[30416]_  = \new_[30415]_  & \new_[30412]_ ;
  assign \new_[30417]_  = \new_[30416]_  & \new_[30409]_ ;
  assign \new_[30421]_  = A234 & A232;
  assign \new_[30422]_  = A203 & \new_[30421]_ ;
  assign \new_[30425]_  = A266 & ~A265;
  assign \new_[30428]_  = A269 & ~A268;
  assign \new_[30429]_  = \new_[30428]_  & \new_[30425]_ ;
  assign \new_[30430]_  = \new_[30429]_  & \new_[30422]_ ;
  assign \new_[30434]_  = ~A167 & A168;
  assign \new_[30435]_  = A169 & \new_[30434]_ ;
  assign \new_[30438]_  = A199 & A166;
  assign \new_[30441]_  = ~A201 & A200;
  assign \new_[30442]_  = \new_[30441]_  & \new_[30438]_ ;
  assign \new_[30443]_  = \new_[30442]_  & \new_[30435]_ ;
  assign \new_[30447]_  = A234 & A232;
  assign \new_[30448]_  = A203 & \new_[30447]_ ;
  assign \new_[30451]_  = ~A266 & A265;
  assign \new_[30454]_  = A269 & ~A268;
  assign \new_[30455]_  = \new_[30454]_  & \new_[30451]_ ;
  assign \new_[30456]_  = \new_[30455]_  & \new_[30448]_ ;
  assign \new_[30460]_  = ~A167 & A168;
  assign \new_[30461]_  = A169 & \new_[30460]_ ;
  assign \new_[30464]_  = A199 & A166;
  assign \new_[30467]_  = ~A201 & A200;
  assign \new_[30468]_  = \new_[30467]_  & \new_[30464]_ ;
  assign \new_[30469]_  = \new_[30468]_  & \new_[30461]_ ;
  assign \new_[30473]_  = A234 & A232;
  assign \new_[30474]_  = A203 & \new_[30473]_ ;
  assign \new_[30477]_  = ~A266 & ~A265;
  assign \new_[30480]_  = ~A269 & A268;
  assign \new_[30481]_  = \new_[30480]_  & \new_[30477]_ ;
  assign \new_[30482]_  = \new_[30481]_  & \new_[30474]_ ;
  assign \new_[30486]_  = ~A167 & A168;
  assign \new_[30487]_  = A169 & \new_[30486]_ ;
  assign \new_[30490]_  = A199 & A166;
  assign \new_[30493]_  = ~A201 & A200;
  assign \new_[30494]_  = \new_[30493]_  & \new_[30490]_ ;
  assign \new_[30495]_  = \new_[30494]_  & \new_[30487]_ ;
  assign \new_[30499]_  = A234 & A233;
  assign \new_[30500]_  = A203 & \new_[30499]_ ;
  assign \new_[30503]_  = A299 & A298;
  assign \new_[30506]_  = ~A302 & A301;
  assign \new_[30507]_  = \new_[30506]_  & \new_[30503]_ ;
  assign \new_[30508]_  = \new_[30507]_  & \new_[30500]_ ;
  assign \new_[30512]_  = ~A167 & A168;
  assign \new_[30513]_  = A169 & \new_[30512]_ ;
  assign \new_[30516]_  = A199 & A166;
  assign \new_[30519]_  = ~A201 & A200;
  assign \new_[30520]_  = \new_[30519]_  & \new_[30516]_ ;
  assign \new_[30521]_  = \new_[30520]_  & \new_[30513]_ ;
  assign \new_[30525]_  = A234 & A233;
  assign \new_[30526]_  = A203 & \new_[30525]_ ;
  assign \new_[30529]_  = ~A299 & A298;
  assign \new_[30532]_  = A302 & ~A301;
  assign \new_[30533]_  = \new_[30532]_  & \new_[30529]_ ;
  assign \new_[30534]_  = \new_[30533]_  & \new_[30526]_ ;
  assign \new_[30538]_  = ~A167 & A168;
  assign \new_[30539]_  = A169 & \new_[30538]_ ;
  assign \new_[30542]_  = A199 & A166;
  assign \new_[30545]_  = ~A201 & A200;
  assign \new_[30546]_  = \new_[30545]_  & \new_[30542]_ ;
  assign \new_[30547]_  = \new_[30546]_  & \new_[30539]_ ;
  assign \new_[30551]_  = A234 & A233;
  assign \new_[30552]_  = A203 & \new_[30551]_ ;
  assign \new_[30555]_  = A299 & ~A298;
  assign \new_[30558]_  = A302 & ~A301;
  assign \new_[30559]_  = \new_[30558]_  & \new_[30555]_ ;
  assign \new_[30560]_  = \new_[30559]_  & \new_[30552]_ ;
  assign \new_[30564]_  = ~A167 & A168;
  assign \new_[30565]_  = A169 & \new_[30564]_ ;
  assign \new_[30568]_  = A199 & A166;
  assign \new_[30571]_  = ~A201 & A200;
  assign \new_[30572]_  = \new_[30571]_  & \new_[30568]_ ;
  assign \new_[30573]_  = \new_[30572]_  & \new_[30565]_ ;
  assign \new_[30577]_  = A234 & A233;
  assign \new_[30578]_  = A203 & \new_[30577]_ ;
  assign \new_[30581]_  = ~A299 & ~A298;
  assign \new_[30584]_  = ~A302 & A301;
  assign \new_[30585]_  = \new_[30584]_  & \new_[30581]_ ;
  assign \new_[30586]_  = \new_[30585]_  & \new_[30578]_ ;
  assign \new_[30590]_  = ~A167 & A168;
  assign \new_[30591]_  = A169 & \new_[30590]_ ;
  assign \new_[30594]_  = A199 & A166;
  assign \new_[30597]_  = ~A201 & A200;
  assign \new_[30598]_  = \new_[30597]_  & \new_[30594]_ ;
  assign \new_[30599]_  = \new_[30598]_  & \new_[30591]_ ;
  assign \new_[30603]_  = A234 & A233;
  assign \new_[30604]_  = A203 & \new_[30603]_ ;
  assign \new_[30607]_  = A266 & A265;
  assign \new_[30610]_  = ~A269 & A268;
  assign \new_[30611]_  = \new_[30610]_  & \new_[30607]_ ;
  assign \new_[30612]_  = \new_[30611]_  & \new_[30604]_ ;
  assign \new_[30616]_  = ~A167 & A168;
  assign \new_[30617]_  = A169 & \new_[30616]_ ;
  assign \new_[30620]_  = A199 & A166;
  assign \new_[30623]_  = ~A201 & A200;
  assign \new_[30624]_  = \new_[30623]_  & \new_[30620]_ ;
  assign \new_[30625]_  = \new_[30624]_  & \new_[30617]_ ;
  assign \new_[30629]_  = A234 & A233;
  assign \new_[30630]_  = A203 & \new_[30629]_ ;
  assign \new_[30633]_  = A266 & ~A265;
  assign \new_[30636]_  = A269 & ~A268;
  assign \new_[30637]_  = \new_[30636]_  & \new_[30633]_ ;
  assign \new_[30638]_  = \new_[30637]_  & \new_[30630]_ ;
  assign \new_[30642]_  = ~A167 & A168;
  assign \new_[30643]_  = A169 & \new_[30642]_ ;
  assign \new_[30646]_  = A199 & A166;
  assign \new_[30649]_  = ~A201 & A200;
  assign \new_[30650]_  = \new_[30649]_  & \new_[30646]_ ;
  assign \new_[30651]_  = \new_[30650]_  & \new_[30643]_ ;
  assign \new_[30655]_  = A234 & A233;
  assign \new_[30656]_  = A203 & \new_[30655]_ ;
  assign \new_[30659]_  = ~A266 & A265;
  assign \new_[30662]_  = A269 & ~A268;
  assign \new_[30663]_  = \new_[30662]_  & \new_[30659]_ ;
  assign \new_[30664]_  = \new_[30663]_  & \new_[30656]_ ;
  assign \new_[30668]_  = ~A167 & A168;
  assign \new_[30669]_  = A169 & \new_[30668]_ ;
  assign \new_[30672]_  = A199 & A166;
  assign \new_[30675]_  = ~A201 & A200;
  assign \new_[30676]_  = \new_[30675]_  & \new_[30672]_ ;
  assign \new_[30677]_  = \new_[30676]_  & \new_[30669]_ ;
  assign \new_[30681]_  = A234 & A233;
  assign \new_[30682]_  = A203 & \new_[30681]_ ;
  assign \new_[30685]_  = ~A266 & ~A265;
  assign \new_[30688]_  = ~A269 & A268;
  assign \new_[30689]_  = \new_[30688]_  & \new_[30685]_ ;
  assign \new_[30690]_  = \new_[30689]_  & \new_[30682]_ ;
  assign \new_[30694]_  = ~A167 & A168;
  assign \new_[30695]_  = A169 & \new_[30694]_ ;
  assign \new_[30698]_  = A199 & A166;
  assign \new_[30701]_  = ~A201 & A200;
  assign \new_[30702]_  = \new_[30701]_  & \new_[30698]_ ;
  assign \new_[30703]_  = \new_[30702]_  & \new_[30695]_ ;
  assign \new_[30707]_  = A233 & A232;
  assign \new_[30708]_  = A203 & \new_[30707]_ ;
  assign \new_[30711]_  = ~A236 & A235;
  assign \new_[30714]_  = A300 & A299;
  assign \new_[30715]_  = \new_[30714]_  & \new_[30711]_ ;
  assign \new_[30716]_  = \new_[30715]_  & \new_[30708]_ ;
  assign \new_[30720]_  = ~A167 & A168;
  assign \new_[30721]_  = A169 & \new_[30720]_ ;
  assign \new_[30724]_  = A199 & A166;
  assign \new_[30727]_  = ~A201 & A200;
  assign \new_[30728]_  = \new_[30727]_  & \new_[30724]_ ;
  assign \new_[30729]_  = \new_[30728]_  & \new_[30721]_ ;
  assign \new_[30733]_  = A233 & A232;
  assign \new_[30734]_  = A203 & \new_[30733]_ ;
  assign \new_[30737]_  = ~A236 & A235;
  assign \new_[30740]_  = A300 & A298;
  assign \new_[30741]_  = \new_[30740]_  & \new_[30737]_ ;
  assign \new_[30742]_  = \new_[30741]_  & \new_[30734]_ ;
  assign \new_[30746]_  = ~A167 & A168;
  assign \new_[30747]_  = A169 & \new_[30746]_ ;
  assign \new_[30750]_  = A199 & A166;
  assign \new_[30753]_  = ~A201 & A200;
  assign \new_[30754]_  = \new_[30753]_  & \new_[30750]_ ;
  assign \new_[30755]_  = \new_[30754]_  & \new_[30747]_ ;
  assign \new_[30759]_  = A233 & A232;
  assign \new_[30760]_  = A203 & \new_[30759]_ ;
  assign \new_[30763]_  = ~A236 & A235;
  assign \new_[30766]_  = A267 & A265;
  assign \new_[30767]_  = \new_[30766]_  & \new_[30763]_ ;
  assign \new_[30768]_  = \new_[30767]_  & \new_[30760]_ ;
  assign \new_[30772]_  = ~A167 & A168;
  assign \new_[30773]_  = A169 & \new_[30772]_ ;
  assign \new_[30776]_  = A199 & A166;
  assign \new_[30779]_  = ~A201 & A200;
  assign \new_[30780]_  = \new_[30779]_  & \new_[30776]_ ;
  assign \new_[30781]_  = \new_[30780]_  & \new_[30773]_ ;
  assign \new_[30785]_  = A233 & A232;
  assign \new_[30786]_  = A203 & \new_[30785]_ ;
  assign \new_[30789]_  = ~A236 & A235;
  assign \new_[30792]_  = A267 & A266;
  assign \new_[30793]_  = \new_[30792]_  & \new_[30789]_ ;
  assign \new_[30794]_  = \new_[30793]_  & \new_[30786]_ ;
  assign \new_[30798]_  = ~A167 & A168;
  assign \new_[30799]_  = A169 & \new_[30798]_ ;
  assign \new_[30802]_  = A199 & A166;
  assign \new_[30805]_  = ~A201 & A200;
  assign \new_[30806]_  = \new_[30805]_  & \new_[30802]_ ;
  assign \new_[30807]_  = \new_[30806]_  & \new_[30799]_ ;
  assign \new_[30811]_  = A233 & ~A232;
  assign \new_[30812]_  = A203 & \new_[30811]_ ;
  assign \new_[30815]_  = A236 & ~A235;
  assign \new_[30818]_  = A300 & A299;
  assign \new_[30819]_  = \new_[30818]_  & \new_[30815]_ ;
  assign \new_[30820]_  = \new_[30819]_  & \new_[30812]_ ;
  assign \new_[30824]_  = ~A167 & A168;
  assign \new_[30825]_  = A169 & \new_[30824]_ ;
  assign \new_[30828]_  = A199 & A166;
  assign \new_[30831]_  = ~A201 & A200;
  assign \new_[30832]_  = \new_[30831]_  & \new_[30828]_ ;
  assign \new_[30833]_  = \new_[30832]_  & \new_[30825]_ ;
  assign \new_[30837]_  = A233 & ~A232;
  assign \new_[30838]_  = A203 & \new_[30837]_ ;
  assign \new_[30841]_  = A236 & ~A235;
  assign \new_[30844]_  = A300 & A298;
  assign \new_[30845]_  = \new_[30844]_  & \new_[30841]_ ;
  assign \new_[30846]_  = \new_[30845]_  & \new_[30838]_ ;
  assign \new_[30850]_  = ~A167 & A168;
  assign \new_[30851]_  = A169 & \new_[30850]_ ;
  assign \new_[30854]_  = A199 & A166;
  assign \new_[30857]_  = ~A201 & A200;
  assign \new_[30858]_  = \new_[30857]_  & \new_[30854]_ ;
  assign \new_[30859]_  = \new_[30858]_  & \new_[30851]_ ;
  assign \new_[30863]_  = A233 & ~A232;
  assign \new_[30864]_  = A203 & \new_[30863]_ ;
  assign \new_[30867]_  = A236 & ~A235;
  assign \new_[30870]_  = A267 & A265;
  assign \new_[30871]_  = \new_[30870]_  & \new_[30867]_ ;
  assign \new_[30872]_  = \new_[30871]_  & \new_[30864]_ ;
  assign \new_[30876]_  = ~A167 & A168;
  assign \new_[30877]_  = A169 & \new_[30876]_ ;
  assign \new_[30880]_  = A199 & A166;
  assign \new_[30883]_  = ~A201 & A200;
  assign \new_[30884]_  = \new_[30883]_  & \new_[30880]_ ;
  assign \new_[30885]_  = \new_[30884]_  & \new_[30877]_ ;
  assign \new_[30889]_  = A233 & ~A232;
  assign \new_[30890]_  = A203 & \new_[30889]_ ;
  assign \new_[30893]_  = A236 & ~A235;
  assign \new_[30896]_  = A267 & A266;
  assign \new_[30897]_  = \new_[30896]_  & \new_[30893]_ ;
  assign \new_[30898]_  = \new_[30897]_  & \new_[30890]_ ;
  assign \new_[30902]_  = ~A167 & A168;
  assign \new_[30903]_  = A169 & \new_[30902]_ ;
  assign \new_[30906]_  = A199 & A166;
  assign \new_[30909]_  = ~A201 & A200;
  assign \new_[30910]_  = \new_[30909]_  & \new_[30906]_ ;
  assign \new_[30911]_  = \new_[30910]_  & \new_[30903]_ ;
  assign \new_[30915]_  = ~A233 & A232;
  assign \new_[30916]_  = A203 & \new_[30915]_ ;
  assign \new_[30919]_  = A236 & ~A235;
  assign \new_[30922]_  = A300 & A299;
  assign \new_[30923]_  = \new_[30922]_  & \new_[30919]_ ;
  assign \new_[30924]_  = \new_[30923]_  & \new_[30916]_ ;
  assign \new_[30928]_  = ~A167 & A168;
  assign \new_[30929]_  = A169 & \new_[30928]_ ;
  assign \new_[30932]_  = A199 & A166;
  assign \new_[30935]_  = ~A201 & A200;
  assign \new_[30936]_  = \new_[30935]_  & \new_[30932]_ ;
  assign \new_[30937]_  = \new_[30936]_  & \new_[30929]_ ;
  assign \new_[30941]_  = ~A233 & A232;
  assign \new_[30942]_  = A203 & \new_[30941]_ ;
  assign \new_[30945]_  = A236 & ~A235;
  assign \new_[30948]_  = A300 & A298;
  assign \new_[30949]_  = \new_[30948]_  & \new_[30945]_ ;
  assign \new_[30950]_  = \new_[30949]_  & \new_[30942]_ ;
  assign \new_[30954]_  = ~A167 & A168;
  assign \new_[30955]_  = A169 & \new_[30954]_ ;
  assign \new_[30958]_  = A199 & A166;
  assign \new_[30961]_  = ~A201 & A200;
  assign \new_[30962]_  = \new_[30961]_  & \new_[30958]_ ;
  assign \new_[30963]_  = \new_[30962]_  & \new_[30955]_ ;
  assign \new_[30967]_  = ~A233 & A232;
  assign \new_[30968]_  = A203 & \new_[30967]_ ;
  assign \new_[30971]_  = A236 & ~A235;
  assign \new_[30974]_  = A267 & A265;
  assign \new_[30975]_  = \new_[30974]_  & \new_[30971]_ ;
  assign \new_[30976]_  = \new_[30975]_  & \new_[30968]_ ;
  assign \new_[30980]_  = ~A167 & A168;
  assign \new_[30981]_  = A169 & \new_[30980]_ ;
  assign \new_[30984]_  = A199 & A166;
  assign \new_[30987]_  = ~A201 & A200;
  assign \new_[30988]_  = \new_[30987]_  & \new_[30984]_ ;
  assign \new_[30989]_  = \new_[30988]_  & \new_[30981]_ ;
  assign \new_[30993]_  = ~A233 & A232;
  assign \new_[30994]_  = A203 & \new_[30993]_ ;
  assign \new_[30997]_  = A236 & ~A235;
  assign \new_[31000]_  = A267 & A266;
  assign \new_[31001]_  = \new_[31000]_  & \new_[30997]_ ;
  assign \new_[31002]_  = \new_[31001]_  & \new_[30994]_ ;
  assign \new_[31006]_  = ~A167 & A168;
  assign \new_[31007]_  = A169 & \new_[31006]_ ;
  assign \new_[31010]_  = A199 & A166;
  assign \new_[31013]_  = ~A201 & A200;
  assign \new_[31014]_  = \new_[31013]_  & \new_[31010]_ ;
  assign \new_[31015]_  = \new_[31014]_  & \new_[31007]_ ;
  assign \new_[31019]_  = ~A233 & ~A232;
  assign \new_[31020]_  = A203 & \new_[31019]_ ;
  assign \new_[31023]_  = ~A236 & A235;
  assign \new_[31026]_  = A300 & A299;
  assign \new_[31027]_  = \new_[31026]_  & \new_[31023]_ ;
  assign \new_[31028]_  = \new_[31027]_  & \new_[31020]_ ;
  assign \new_[31032]_  = ~A167 & A168;
  assign \new_[31033]_  = A169 & \new_[31032]_ ;
  assign \new_[31036]_  = A199 & A166;
  assign \new_[31039]_  = ~A201 & A200;
  assign \new_[31040]_  = \new_[31039]_  & \new_[31036]_ ;
  assign \new_[31041]_  = \new_[31040]_  & \new_[31033]_ ;
  assign \new_[31045]_  = ~A233 & ~A232;
  assign \new_[31046]_  = A203 & \new_[31045]_ ;
  assign \new_[31049]_  = ~A236 & A235;
  assign \new_[31052]_  = A300 & A298;
  assign \new_[31053]_  = \new_[31052]_  & \new_[31049]_ ;
  assign \new_[31054]_  = \new_[31053]_  & \new_[31046]_ ;
  assign \new_[31058]_  = ~A167 & A168;
  assign \new_[31059]_  = A169 & \new_[31058]_ ;
  assign \new_[31062]_  = A199 & A166;
  assign \new_[31065]_  = ~A201 & A200;
  assign \new_[31066]_  = \new_[31065]_  & \new_[31062]_ ;
  assign \new_[31067]_  = \new_[31066]_  & \new_[31059]_ ;
  assign \new_[31071]_  = ~A233 & ~A232;
  assign \new_[31072]_  = A203 & \new_[31071]_ ;
  assign \new_[31075]_  = ~A236 & A235;
  assign \new_[31078]_  = A267 & A265;
  assign \new_[31079]_  = \new_[31078]_  & \new_[31075]_ ;
  assign \new_[31080]_  = \new_[31079]_  & \new_[31072]_ ;
  assign \new_[31084]_  = ~A167 & A168;
  assign \new_[31085]_  = A169 & \new_[31084]_ ;
  assign \new_[31088]_  = A199 & A166;
  assign \new_[31091]_  = ~A201 & A200;
  assign \new_[31092]_  = \new_[31091]_  & \new_[31088]_ ;
  assign \new_[31093]_  = \new_[31092]_  & \new_[31085]_ ;
  assign \new_[31097]_  = ~A233 & ~A232;
  assign \new_[31098]_  = A203 & \new_[31097]_ ;
  assign \new_[31101]_  = ~A236 & A235;
  assign \new_[31104]_  = A267 & A266;
  assign \new_[31105]_  = \new_[31104]_  & \new_[31101]_ ;
  assign \new_[31106]_  = \new_[31105]_  & \new_[31098]_ ;
  assign \new_[31110]_  = ~A167 & A168;
  assign \new_[31111]_  = A169 & \new_[31110]_ ;
  assign \new_[31114]_  = ~A199 & A166;
  assign \new_[31117]_  = ~A201 & A200;
  assign \new_[31118]_  = \new_[31117]_  & \new_[31114]_ ;
  assign \new_[31119]_  = \new_[31118]_  & \new_[31111]_ ;
  assign \new_[31123]_  = A234 & A232;
  assign \new_[31124]_  = A202 & \new_[31123]_ ;
  assign \new_[31127]_  = A299 & A298;
  assign \new_[31130]_  = ~A302 & A301;
  assign \new_[31131]_  = \new_[31130]_  & \new_[31127]_ ;
  assign \new_[31132]_  = \new_[31131]_  & \new_[31124]_ ;
  assign \new_[31136]_  = ~A167 & A168;
  assign \new_[31137]_  = A169 & \new_[31136]_ ;
  assign \new_[31140]_  = ~A199 & A166;
  assign \new_[31143]_  = ~A201 & A200;
  assign \new_[31144]_  = \new_[31143]_  & \new_[31140]_ ;
  assign \new_[31145]_  = \new_[31144]_  & \new_[31137]_ ;
  assign \new_[31149]_  = A234 & A232;
  assign \new_[31150]_  = A202 & \new_[31149]_ ;
  assign \new_[31153]_  = ~A299 & A298;
  assign \new_[31156]_  = A302 & ~A301;
  assign \new_[31157]_  = \new_[31156]_  & \new_[31153]_ ;
  assign \new_[31158]_  = \new_[31157]_  & \new_[31150]_ ;
  assign \new_[31162]_  = ~A167 & A168;
  assign \new_[31163]_  = A169 & \new_[31162]_ ;
  assign \new_[31166]_  = ~A199 & A166;
  assign \new_[31169]_  = ~A201 & A200;
  assign \new_[31170]_  = \new_[31169]_  & \new_[31166]_ ;
  assign \new_[31171]_  = \new_[31170]_  & \new_[31163]_ ;
  assign \new_[31175]_  = A234 & A232;
  assign \new_[31176]_  = A202 & \new_[31175]_ ;
  assign \new_[31179]_  = A299 & ~A298;
  assign \new_[31182]_  = A302 & ~A301;
  assign \new_[31183]_  = \new_[31182]_  & \new_[31179]_ ;
  assign \new_[31184]_  = \new_[31183]_  & \new_[31176]_ ;
  assign \new_[31188]_  = ~A167 & A168;
  assign \new_[31189]_  = A169 & \new_[31188]_ ;
  assign \new_[31192]_  = ~A199 & A166;
  assign \new_[31195]_  = ~A201 & A200;
  assign \new_[31196]_  = \new_[31195]_  & \new_[31192]_ ;
  assign \new_[31197]_  = \new_[31196]_  & \new_[31189]_ ;
  assign \new_[31201]_  = A234 & A232;
  assign \new_[31202]_  = A202 & \new_[31201]_ ;
  assign \new_[31205]_  = ~A299 & ~A298;
  assign \new_[31208]_  = ~A302 & A301;
  assign \new_[31209]_  = \new_[31208]_  & \new_[31205]_ ;
  assign \new_[31210]_  = \new_[31209]_  & \new_[31202]_ ;
  assign \new_[31214]_  = ~A167 & A168;
  assign \new_[31215]_  = A169 & \new_[31214]_ ;
  assign \new_[31218]_  = ~A199 & A166;
  assign \new_[31221]_  = ~A201 & A200;
  assign \new_[31222]_  = \new_[31221]_  & \new_[31218]_ ;
  assign \new_[31223]_  = \new_[31222]_  & \new_[31215]_ ;
  assign \new_[31227]_  = A234 & A232;
  assign \new_[31228]_  = A202 & \new_[31227]_ ;
  assign \new_[31231]_  = A266 & A265;
  assign \new_[31234]_  = ~A269 & A268;
  assign \new_[31235]_  = \new_[31234]_  & \new_[31231]_ ;
  assign \new_[31236]_  = \new_[31235]_  & \new_[31228]_ ;
  assign \new_[31240]_  = ~A167 & A168;
  assign \new_[31241]_  = A169 & \new_[31240]_ ;
  assign \new_[31244]_  = ~A199 & A166;
  assign \new_[31247]_  = ~A201 & A200;
  assign \new_[31248]_  = \new_[31247]_  & \new_[31244]_ ;
  assign \new_[31249]_  = \new_[31248]_  & \new_[31241]_ ;
  assign \new_[31253]_  = A234 & A232;
  assign \new_[31254]_  = A202 & \new_[31253]_ ;
  assign \new_[31257]_  = A266 & ~A265;
  assign \new_[31260]_  = A269 & ~A268;
  assign \new_[31261]_  = \new_[31260]_  & \new_[31257]_ ;
  assign \new_[31262]_  = \new_[31261]_  & \new_[31254]_ ;
  assign \new_[31266]_  = ~A167 & A168;
  assign \new_[31267]_  = A169 & \new_[31266]_ ;
  assign \new_[31270]_  = ~A199 & A166;
  assign \new_[31273]_  = ~A201 & A200;
  assign \new_[31274]_  = \new_[31273]_  & \new_[31270]_ ;
  assign \new_[31275]_  = \new_[31274]_  & \new_[31267]_ ;
  assign \new_[31279]_  = A234 & A232;
  assign \new_[31280]_  = A202 & \new_[31279]_ ;
  assign \new_[31283]_  = ~A266 & A265;
  assign \new_[31286]_  = A269 & ~A268;
  assign \new_[31287]_  = \new_[31286]_  & \new_[31283]_ ;
  assign \new_[31288]_  = \new_[31287]_  & \new_[31280]_ ;
  assign \new_[31292]_  = ~A167 & A168;
  assign \new_[31293]_  = A169 & \new_[31292]_ ;
  assign \new_[31296]_  = ~A199 & A166;
  assign \new_[31299]_  = ~A201 & A200;
  assign \new_[31300]_  = \new_[31299]_  & \new_[31296]_ ;
  assign \new_[31301]_  = \new_[31300]_  & \new_[31293]_ ;
  assign \new_[31305]_  = A234 & A232;
  assign \new_[31306]_  = A202 & \new_[31305]_ ;
  assign \new_[31309]_  = ~A266 & ~A265;
  assign \new_[31312]_  = ~A269 & A268;
  assign \new_[31313]_  = \new_[31312]_  & \new_[31309]_ ;
  assign \new_[31314]_  = \new_[31313]_  & \new_[31306]_ ;
  assign \new_[31318]_  = ~A167 & A168;
  assign \new_[31319]_  = A169 & \new_[31318]_ ;
  assign \new_[31322]_  = ~A199 & A166;
  assign \new_[31325]_  = ~A201 & A200;
  assign \new_[31326]_  = \new_[31325]_  & \new_[31322]_ ;
  assign \new_[31327]_  = \new_[31326]_  & \new_[31319]_ ;
  assign \new_[31331]_  = A234 & A233;
  assign \new_[31332]_  = A202 & \new_[31331]_ ;
  assign \new_[31335]_  = A299 & A298;
  assign \new_[31338]_  = ~A302 & A301;
  assign \new_[31339]_  = \new_[31338]_  & \new_[31335]_ ;
  assign \new_[31340]_  = \new_[31339]_  & \new_[31332]_ ;
  assign \new_[31344]_  = ~A167 & A168;
  assign \new_[31345]_  = A169 & \new_[31344]_ ;
  assign \new_[31348]_  = ~A199 & A166;
  assign \new_[31351]_  = ~A201 & A200;
  assign \new_[31352]_  = \new_[31351]_  & \new_[31348]_ ;
  assign \new_[31353]_  = \new_[31352]_  & \new_[31345]_ ;
  assign \new_[31357]_  = A234 & A233;
  assign \new_[31358]_  = A202 & \new_[31357]_ ;
  assign \new_[31361]_  = ~A299 & A298;
  assign \new_[31364]_  = A302 & ~A301;
  assign \new_[31365]_  = \new_[31364]_  & \new_[31361]_ ;
  assign \new_[31366]_  = \new_[31365]_  & \new_[31358]_ ;
  assign \new_[31370]_  = ~A167 & A168;
  assign \new_[31371]_  = A169 & \new_[31370]_ ;
  assign \new_[31374]_  = ~A199 & A166;
  assign \new_[31377]_  = ~A201 & A200;
  assign \new_[31378]_  = \new_[31377]_  & \new_[31374]_ ;
  assign \new_[31379]_  = \new_[31378]_  & \new_[31371]_ ;
  assign \new_[31383]_  = A234 & A233;
  assign \new_[31384]_  = A202 & \new_[31383]_ ;
  assign \new_[31387]_  = A299 & ~A298;
  assign \new_[31390]_  = A302 & ~A301;
  assign \new_[31391]_  = \new_[31390]_  & \new_[31387]_ ;
  assign \new_[31392]_  = \new_[31391]_  & \new_[31384]_ ;
  assign \new_[31396]_  = ~A167 & A168;
  assign \new_[31397]_  = A169 & \new_[31396]_ ;
  assign \new_[31400]_  = ~A199 & A166;
  assign \new_[31403]_  = ~A201 & A200;
  assign \new_[31404]_  = \new_[31403]_  & \new_[31400]_ ;
  assign \new_[31405]_  = \new_[31404]_  & \new_[31397]_ ;
  assign \new_[31409]_  = A234 & A233;
  assign \new_[31410]_  = A202 & \new_[31409]_ ;
  assign \new_[31413]_  = ~A299 & ~A298;
  assign \new_[31416]_  = ~A302 & A301;
  assign \new_[31417]_  = \new_[31416]_  & \new_[31413]_ ;
  assign \new_[31418]_  = \new_[31417]_  & \new_[31410]_ ;
  assign \new_[31422]_  = ~A167 & A168;
  assign \new_[31423]_  = A169 & \new_[31422]_ ;
  assign \new_[31426]_  = ~A199 & A166;
  assign \new_[31429]_  = ~A201 & A200;
  assign \new_[31430]_  = \new_[31429]_  & \new_[31426]_ ;
  assign \new_[31431]_  = \new_[31430]_  & \new_[31423]_ ;
  assign \new_[31435]_  = A234 & A233;
  assign \new_[31436]_  = A202 & \new_[31435]_ ;
  assign \new_[31439]_  = A266 & A265;
  assign \new_[31442]_  = ~A269 & A268;
  assign \new_[31443]_  = \new_[31442]_  & \new_[31439]_ ;
  assign \new_[31444]_  = \new_[31443]_  & \new_[31436]_ ;
  assign \new_[31448]_  = ~A167 & A168;
  assign \new_[31449]_  = A169 & \new_[31448]_ ;
  assign \new_[31452]_  = ~A199 & A166;
  assign \new_[31455]_  = ~A201 & A200;
  assign \new_[31456]_  = \new_[31455]_  & \new_[31452]_ ;
  assign \new_[31457]_  = \new_[31456]_  & \new_[31449]_ ;
  assign \new_[31461]_  = A234 & A233;
  assign \new_[31462]_  = A202 & \new_[31461]_ ;
  assign \new_[31465]_  = A266 & ~A265;
  assign \new_[31468]_  = A269 & ~A268;
  assign \new_[31469]_  = \new_[31468]_  & \new_[31465]_ ;
  assign \new_[31470]_  = \new_[31469]_  & \new_[31462]_ ;
  assign \new_[31474]_  = ~A167 & A168;
  assign \new_[31475]_  = A169 & \new_[31474]_ ;
  assign \new_[31478]_  = ~A199 & A166;
  assign \new_[31481]_  = ~A201 & A200;
  assign \new_[31482]_  = \new_[31481]_  & \new_[31478]_ ;
  assign \new_[31483]_  = \new_[31482]_  & \new_[31475]_ ;
  assign \new_[31487]_  = A234 & A233;
  assign \new_[31488]_  = A202 & \new_[31487]_ ;
  assign \new_[31491]_  = ~A266 & A265;
  assign \new_[31494]_  = A269 & ~A268;
  assign \new_[31495]_  = \new_[31494]_  & \new_[31491]_ ;
  assign \new_[31496]_  = \new_[31495]_  & \new_[31488]_ ;
  assign \new_[31500]_  = ~A167 & A168;
  assign \new_[31501]_  = A169 & \new_[31500]_ ;
  assign \new_[31504]_  = ~A199 & A166;
  assign \new_[31507]_  = ~A201 & A200;
  assign \new_[31508]_  = \new_[31507]_  & \new_[31504]_ ;
  assign \new_[31509]_  = \new_[31508]_  & \new_[31501]_ ;
  assign \new_[31513]_  = A234 & A233;
  assign \new_[31514]_  = A202 & \new_[31513]_ ;
  assign \new_[31517]_  = ~A266 & ~A265;
  assign \new_[31520]_  = ~A269 & A268;
  assign \new_[31521]_  = \new_[31520]_  & \new_[31517]_ ;
  assign \new_[31522]_  = \new_[31521]_  & \new_[31514]_ ;
  assign \new_[31526]_  = ~A167 & A168;
  assign \new_[31527]_  = A169 & \new_[31526]_ ;
  assign \new_[31530]_  = ~A199 & A166;
  assign \new_[31533]_  = ~A201 & A200;
  assign \new_[31534]_  = \new_[31533]_  & \new_[31530]_ ;
  assign \new_[31535]_  = \new_[31534]_  & \new_[31527]_ ;
  assign \new_[31539]_  = A233 & A232;
  assign \new_[31540]_  = A202 & \new_[31539]_ ;
  assign \new_[31543]_  = ~A236 & A235;
  assign \new_[31546]_  = A300 & A299;
  assign \new_[31547]_  = \new_[31546]_  & \new_[31543]_ ;
  assign \new_[31548]_  = \new_[31547]_  & \new_[31540]_ ;
  assign \new_[31552]_  = ~A167 & A168;
  assign \new_[31553]_  = A169 & \new_[31552]_ ;
  assign \new_[31556]_  = ~A199 & A166;
  assign \new_[31559]_  = ~A201 & A200;
  assign \new_[31560]_  = \new_[31559]_  & \new_[31556]_ ;
  assign \new_[31561]_  = \new_[31560]_  & \new_[31553]_ ;
  assign \new_[31565]_  = A233 & A232;
  assign \new_[31566]_  = A202 & \new_[31565]_ ;
  assign \new_[31569]_  = ~A236 & A235;
  assign \new_[31572]_  = A300 & A298;
  assign \new_[31573]_  = \new_[31572]_  & \new_[31569]_ ;
  assign \new_[31574]_  = \new_[31573]_  & \new_[31566]_ ;
  assign \new_[31578]_  = ~A167 & A168;
  assign \new_[31579]_  = A169 & \new_[31578]_ ;
  assign \new_[31582]_  = ~A199 & A166;
  assign \new_[31585]_  = ~A201 & A200;
  assign \new_[31586]_  = \new_[31585]_  & \new_[31582]_ ;
  assign \new_[31587]_  = \new_[31586]_  & \new_[31579]_ ;
  assign \new_[31591]_  = A233 & A232;
  assign \new_[31592]_  = A202 & \new_[31591]_ ;
  assign \new_[31595]_  = ~A236 & A235;
  assign \new_[31598]_  = A267 & A265;
  assign \new_[31599]_  = \new_[31598]_  & \new_[31595]_ ;
  assign \new_[31600]_  = \new_[31599]_  & \new_[31592]_ ;
  assign \new_[31604]_  = ~A167 & A168;
  assign \new_[31605]_  = A169 & \new_[31604]_ ;
  assign \new_[31608]_  = ~A199 & A166;
  assign \new_[31611]_  = ~A201 & A200;
  assign \new_[31612]_  = \new_[31611]_  & \new_[31608]_ ;
  assign \new_[31613]_  = \new_[31612]_  & \new_[31605]_ ;
  assign \new_[31617]_  = A233 & A232;
  assign \new_[31618]_  = A202 & \new_[31617]_ ;
  assign \new_[31621]_  = ~A236 & A235;
  assign \new_[31624]_  = A267 & A266;
  assign \new_[31625]_  = \new_[31624]_  & \new_[31621]_ ;
  assign \new_[31626]_  = \new_[31625]_  & \new_[31618]_ ;
  assign \new_[31630]_  = ~A167 & A168;
  assign \new_[31631]_  = A169 & \new_[31630]_ ;
  assign \new_[31634]_  = ~A199 & A166;
  assign \new_[31637]_  = ~A201 & A200;
  assign \new_[31638]_  = \new_[31637]_  & \new_[31634]_ ;
  assign \new_[31639]_  = \new_[31638]_  & \new_[31631]_ ;
  assign \new_[31643]_  = A233 & ~A232;
  assign \new_[31644]_  = A202 & \new_[31643]_ ;
  assign \new_[31647]_  = A236 & ~A235;
  assign \new_[31650]_  = A300 & A299;
  assign \new_[31651]_  = \new_[31650]_  & \new_[31647]_ ;
  assign \new_[31652]_  = \new_[31651]_  & \new_[31644]_ ;
  assign \new_[31656]_  = ~A167 & A168;
  assign \new_[31657]_  = A169 & \new_[31656]_ ;
  assign \new_[31660]_  = ~A199 & A166;
  assign \new_[31663]_  = ~A201 & A200;
  assign \new_[31664]_  = \new_[31663]_  & \new_[31660]_ ;
  assign \new_[31665]_  = \new_[31664]_  & \new_[31657]_ ;
  assign \new_[31669]_  = A233 & ~A232;
  assign \new_[31670]_  = A202 & \new_[31669]_ ;
  assign \new_[31673]_  = A236 & ~A235;
  assign \new_[31676]_  = A300 & A298;
  assign \new_[31677]_  = \new_[31676]_  & \new_[31673]_ ;
  assign \new_[31678]_  = \new_[31677]_  & \new_[31670]_ ;
  assign \new_[31682]_  = ~A167 & A168;
  assign \new_[31683]_  = A169 & \new_[31682]_ ;
  assign \new_[31686]_  = ~A199 & A166;
  assign \new_[31689]_  = ~A201 & A200;
  assign \new_[31690]_  = \new_[31689]_  & \new_[31686]_ ;
  assign \new_[31691]_  = \new_[31690]_  & \new_[31683]_ ;
  assign \new_[31695]_  = A233 & ~A232;
  assign \new_[31696]_  = A202 & \new_[31695]_ ;
  assign \new_[31699]_  = A236 & ~A235;
  assign \new_[31702]_  = A267 & A265;
  assign \new_[31703]_  = \new_[31702]_  & \new_[31699]_ ;
  assign \new_[31704]_  = \new_[31703]_  & \new_[31696]_ ;
  assign \new_[31708]_  = ~A167 & A168;
  assign \new_[31709]_  = A169 & \new_[31708]_ ;
  assign \new_[31712]_  = ~A199 & A166;
  assign \new_[31715]_  = ~A201 & A200;
  assign \new_[31716]_  = \new_[31715]_  & \new_[31712]_ ;
  assign \new_[31717]_  = \new_[31716]_  & \new_[31709]_ ;
  assign \new_[31721]_  = A233 & ~A232;
  assign \new_[31722]_  = A202 & \new_[31721]_ ;
  assign \new_[31725]_  = A236 & ~A235;
  assign \new_[31728]_  = A267 & A266;
  assign \new_[31729]_  = \new_[31728]_  & \new_[31725]_ ;
  assign \new_[31730]_  = \new_[31729]_  & \new_[31722]_ ;
  assign \new_[31734]_  = ~A167 & A168;
  assign \new_[31735]_  = A169 & \new_[31734]_ ;
  assign \new_[31738]_  = ~A199 & A166;
  assign \new_[31741]_  = ~A201 & A200;
  assign \new_[31742]_  = \new_[31741]_  & \new_[31738]_ ;
  assign \new_[31743]_  = \new_[31742]_  & \new_[31735]_ ;
  assign \new_[31747]_  = ~A233 & A232;
  assign \new_[31748]_  = A202 & \new_[31747]_ ;
  assign \new_[31751]_  = A236 & ~A235;
  assign \new_[31754]_  = A300 & A299;
  assign \new_[31755]_  = \new_[31754]_  & \new_[31751]_ ;
  assign \new_[31756]_  = \new_[31755]_  & \new_[31748]_ ;
  assign \new_[31760]_  = ~A167 & A168;
  assign \new_[31761]_  = A169 & \new_[31760]_ ;
  assign \new_[31764]_  = ~A199 & A166;
  assign \new_[31767]_  = ~A201 & A200;
  assign \new_[31768]_  = \new_[31767]_  & \new_[31764]_ ;
  assign \new_[31769]_  = \new_[31768]_  & \new_[31761]_ ;
  assign \new_[31773]_  = ~A233 & A232;
  assign \new_[31774]_  = A202 & \new_[31773]_ ;
  assign \new_[31777]_  = A236 & ~A235;
  assign \new_[31780]_  = A300 & A298;
  assign \new_[31781]_  = \new_[31780]_  & \new_[31777]_ ;
  assign \new_[31782]_  = \new_[31781]_  & \new_[31774]_ ;
  assign \new_[31786]_  = ~A167 & A168;
  assign \new_[31787]_  = A169 & \new_[31786]_ ;
  assign \new_[31790]_  = ~A199 & A166;
  assign \new_[31793]_  = ~A201 & A200;
  assign \new_[31794]_  = \new_[31793]_  & \new_[31790]_ ;
  assign \new_[31795]_  = \new_[31794]_  & \new_[31787]_ ;
  assign \new_[31799]_  = ~A233 & A232;
  assign \new_[31800]_  = A202 & \new_[31799]_ ;
  assign \new_[31803]_  = A236 & ~A235;
  assign \new_[31806]_  = A267 & A265;
  assign \new_[31807]_  = \new_[31806]_  & \new_[31803]_ ;
  assign \new_[31808]_  = \new_[31807]_  & \new_[31800]_ ;
  assign \new_[31812]_  = ~A167 & A168;
  assign \new_[31813]_  = A169 & \new_[31812]_ ;
  assign \new_[31816]_  = ~A199 & A166;
  assign \new_[31819]_  = ~A201 & A200;
  assign \new_[31820]_  = \new_[31819]_  & \new_[31816]_ ;
  assign \new_[31821]_  = \new_[31820]_  & \new_[31813]_ ;
  assign \new_[31825]_  = ~A233 & A232;
  assign \new_[31826]_  = A202 & \new_[31825]_ ;
  assign \new_[31829]_  = A236 & ~A235;
  assign \new_[31832]_  = A267 & A266;
  assign \new_[31833]_  = \new_[31832]_  & \new_[31829]_ ;
  assign \new_[31834]_  = \new_[31833]_  & \new_[31826]_ ;
  assign \new_[31838]_  = ~A167 & A168;
  assign \new_[31839]_  = A169 & \new_[31838]_ ;
  assign \new_[31842]_  = ~A199 & A166;
  assign \new_[31845]_  = ~A201 & A200;
  assign \new_[31846]_  = \new_[31845]_  & \new_[31842]_ ;
  assign \new_[31847]_  = \new_[31846]_  & \new_[31839]_ ;
  assign \new_[31851]_  = ~A233 & ~A232;
  assign \new_[31852]_  = A202 & \new_[31851]_ ;
  assign \new_[31855]_  = ~A236 & A235;
  assign \new_[31858]_  = A300 & A299;
  assign \new_[31859]_  = \new_[31858]_  & \new_[31855]_ ;
  assign \new_[31860]_  = \new_[31859]_  & \new_[31852]_ ;
  assign \new_[31864]_  = ~A167 & A168;
  assign \new_[31865]_  = A169 & \new_[31864]_ ;
  assign \new_[31868]_  = ~A199 & A166;
  assign \new_[31871]_  = ~A201 & A200;
  assign \new_[31872]_  = \new_[31871]_  & \new_[31868]_ ;
  assign \new_[31873]_  = \new_[31872]_  & \new_[31865]_ ;
  assign \new_[31877]_  = ~A233 & ~A232;
  assign \new_[31878]_  = A202 & \new_[31877]_ ;
  assign \new_[31881]_  = ~A236 & A235;
  assign \new_[31884]_  = A300 & A298;
  assign \new_[31885]_  = \new_[31884]_  & \new_[31881]_ ;
  assign \new_[31886]_  = \new_[31885]_  & \new_[31878]_ ;
  assign \new_[31890]_  = ~A167 & A168;
  assign \new_[31891]_  = A169 & \new_[31890]_ ;
  assign \new_[31894]_  = ~A199 & A166;
  assign \new_[31897]_  = ~A201 & A200;
  assign \new_[31898]_  = \new_[31897]_  & \new_[31894]_ ;
  assign \new_[31899]_  = \new_[31898]_  & \new_[31891]_ ;
  assign \new_[31903]_  = ~A233 & ~A232;
  assign \new_[31904]_  = A202 & \new_[31903]_ ;
  assign \new_[31907]_  = ~A236 & A235;
  assign \new_[31910]_  = A267 & A265;
  assign \new_[31911]_  = \new_[31910]_  & \new_[31907]_ ;
  assign \new_[31912]_  = \new_[31911]_  & \new_[31904]_ ;
  assign \new_[31916]_  = ~A167 & A168;
  assign \new_[31917]_  = A169 & \new_[31916]_ ;
  assign \new_[31920]_  = ~A199 & A166;
  assign \new_[31923]_  = ~A201 & A200;
  assign \new_[31924]_  = \new_[31923]_  & \new_[31920]_ ;
  assign \new_[31925]_  = \new_[31924]_  & \new_[31917]_ ;
  assign \new_[31929]_  = ~A233 & ~A232;
  assign \new_[31930]_  = A202 & \new_[31929]_ ;
  assign \new_[31933]_  = ~A236 & A235;
  assign \new_[31936]_  = A267 & A266;
  assign \new_[31937]_  = \new_[31936]_  & \new_[31933]_ ;
  assign \new_[31938]_  = \new_[31937]_  & \new_[31930]_ ;
  assign \new_[31942]_  = ~A167 & A168;
  assign \new_[31943]_  = A169 & \new_[31942]_ ;
  assign \new_[31946]_  = ~A199 & A166;
  assign \new_[31949]_  = ~A201 & A200;
  assign \new_[31950]_  = \new_[31949]_  & \new_[31946]_ ;
  assign \new_[31951]_  = \new_[31950]_  & \new_[31943]_ ;
  assign \new_[31955]_  = A234 & A232;
  assign \new_[31956]_  = ~A203 & \new_[31955]_ ;
  assign \new_[31959]_  = A299 & A298;
  assign \new_[31962]_  = ~A302 & A301;
  assign \new_[31963]_  = \new_[31962]_  & \new_[31959]_ ;
  assign \new_[31964]_  = \new_[31963]_  & \new_[31956]_ ;
  assign \new_[31968]_  = ~A167 & A168;
  assign \new_[31969]_  = A169 & \new_[31968]_ ;
  assign \new_[31972]_  = ~A199 & A166;
  assign \new_[31975]_  = ~A201 & A200;
  assign \new_[31976]_  = \new_[31975]_  & \new_[31972]_ ;
  assign \new_[31977]_  = \new_[31976]_  & \new_[31969]_ ;
  assign \new_[31981]_  = A234 & A232;
  assign \new_[31982]_  = ~A203 & \new_[31981]_ ;
  assign \new_[31985]_  = ~A299 & A298;
  assign \new_[31988]_  = A302 & ~A301;
  assign \new_[31989]_  = \new_[31988]_  & \new_[31985]_ ;
  assign \new_[31990]_  = \new_[31989]_  & \new_[31982]_ ;
  assign \new_[31994]_  = ~A167 & A168;
  assign \new_[31995]_  = A169 & \new_[31994]_ ;
  assign \new_[31998]_  = ~A199 & A166;
  assign \new_[32001]_  = ~A201 & A200;
  assign \new_[32002]_  = \new_[32001]_  & \new_[31998]_ ;
  assign \new_[32003]_  = \new_[32002]_  & \new_[31995]_ ;
  assign \new_[32007]_  = A234 & A232;
  assign \new_[32008]_  = ~A203 & \new_[32007]_ ;
  assign \new_[32011]_  = A299 & ~A298;
  assign \new_[32014]_  = A302 & ~A301;
  assign \new_[32015]_  = \new_[32014]_  & \new_[32011]_ ;
  assign \new_[32016]_  = \new_[32015]_  & \new_[32008]_ ;
  assign \new_[32020]_  = ~A167 & A168;
  assign \new_[32021]_  = A169 & \new_[32020]_ ;
  assign \new_[32024]_  = ~A199 & A166;
  assign \new_[32027]_  = ~A201 & A200;
  assign \new_[32028]_  = \new_[32027]_  & \new_[32024]_ ;
  assign \new_[32029]_  = \new_[32028]_  & \new_[32021]_ ;
  assign \new_[32033]_  = A234 & A232;
  assign \new_[32034]_  = ~A203 & \new_[32033]_ ;
  assign \new_[32037]_  = ~A299 & ~A298;
  assign \new_[32040]_  = ~A302 & A301;
  assign \new_[32041]_  = \new_[32040]_  & \new_[32037]_ ;
  assign \new_[32042]_  = \new_[32041]_  & \new_[32034]_ ;
  assign \new_[32046]_  = ~A167 & A168;
  assign \new_[32047]_  = A169 & \new_[32046]_ ;
  assign \new_[32050]_  = ~A199 & A166;
  assign \new_[32053]_  = ~A201 & A200;
  assign \new_[32054]_  = \new_[32053]_  & \new_[32050]_ ;
  assign \new_[32055]_  = \new_[32054]_  & \new_[32047]_ ;
  assign \new_[32059]_  = A234 & A232;
  assign \new_[32060]_  = ~A203 & \new_[32059]_ ;
  assign \new_[32063]_  = A266 & A265;
  assign \new_[32066]_  = ~A269 & A268;
  assign \new_[32067]_  = \new_[32066]_  & \new_[32063]_ ;
  assign \new_[32068]_  = \new_[32067]_  & \new_[32060]_ ;
  assign \new_[32072]_  = ~A167 & A168;
  assign \new_[32073]_  = A169 & \new_[32072]_ ;
  assign \new_[32076]_  = ~A199 & A166;
  assign \new_[32079]_  = ~A201 & A200;
  assign \new_[32080]_  = \new_[32079]_  & \new_[32076]_ ;
  assign \new_[32081]_  = \new_[32080]_  & \new_[32073]_ ;
  assign \new_[32085]_  = A234 & A232;
  assign \new_[32086]_  = ~A203 & \new_[32085]_ ;
  assign \new_[32089]_  = A266 & ~A265;
  assign \new_[32092]_  = A269 & ~A268;
  assign \new_[32093]_  = \new_[32092]_  & \new_[32089]_ ;
  assign \new_[32094]_  = \new_[32093]_  & \new_[32086]_ ;
  assign \new_[32098]_  = ~A167 & A168;
  assign \new_[32099]_  = A169 & \new_[32098]_ ;
  assign \new_[32102]_  = ~A199 & A166;
  assign \new_[32105]_  = ~A201 & A200;
  assign \new_[32106]_  = \new_[32105]_  & \new_[32102]_ ;
  assign \new_[32107]_  = \new_[32106]_  & \new_[32099]_ ;
  assign \new_[32111]_  = A234 & A232;
  assign \new_[32112]_  = ~A203 & \new_[32111]_ ;
  assign \new_[32115]_  = ~A266 & A265;
  assign \new_[32118]_  = A269 & ~A268;
  assign \new_[32119]_  = \new_[32118]_  & \new_[32115]_ ;
  assign \new_[32120]_  = \new_[32119]_  & \new_[32112]_ ;
  assign \new_[32124]_  = ~A167 & A168;
  assign \new_[32125]_  = A169 & \new_[32124]_ ;
  assign \new_[32128]_  = ~A199 & A166;
  assign \new_[32131]_  = ~A201 & A200;
  assign \new_[32132]_  = \new_[32131]_  & \new_[32128]_ ;
  assign \new_[32133]_  = \new_[32132]_  & \new_[32125]_ ;
  assign \new_[32137]_  = A234 & A232;
  assign \new_[32138]_  = ~A203 & \new_[32137]_ ;
  assign \new_[32141]_  = ~A266 & ~A265;
  assign \new_[32144]_  = ~A269 & A268;
  assign \new_[32145]_  = \new_[32144]_  & \new_[32141]_ ;
  assign \new_[32146]_  = \new_[32145]_  & \new_[32138]_ ;
  assign \new_[32150]_  = ~A167 & A168;
  assign \new_[32151]_  = A169 & \new_[32150]_ ;
  assign \new_[32154]_  = ~A199 & A166;
  assign \new_[32157]_  = ~A201 & A200;
  assign \new_[32158]_  = \new_[32157]_  & \new_[32154]_ ;
  assign \new_[32159]_  = \new_[32158]_  & \new_[32151]_ ;
  assign \new_[32163]_  = A234 & A233;
  assign \new_[32164]_  = ~A203 & \new_[32163]_ ;
  assign \new_[32167]_  = A299 & A298;
  assign \new_[32170]_  = ~A302 & A301;
  assign \new_[32171]_  = \new_[32170]_  & \new_[32167]_ ;
  assign \new_[32172]_  = \new_[32171]_  & \new_[32164]_ ;
  assign \new_[32176]_  = ~A167 & A168;
  assign \new_[32177]_  = A169 & \new_[32176]_ ;
  assign \new_[32180]_  = ~A199 & A166;
  assign \new_[32183]_  = ~A201 & A200;
  assign \new_[32184]_  = \new_[32183]_  & \new_[32180]_ ;
  assign \new_[32185]_  = \new_[32184]_  & \new_[32177]_ ;
  assign \new_[32189]_  = A234 & A233;
  assign \new_[32190]_  = ~A203 & \new_[32189]_ ;
  assign \new_[32193]_  = ~A299 & A298;
  assign \new_[32196]_  = A302 & ~A301;
  assign \new_[32197]_  = \new_[32196]_  & \new_[32193]_ ;
  assign \new_[32198]_  = \new_[32197]_  & \new_[32190]_ ;
  assign \new_[32202]_  = ~A167 & A168;
  assign \new_[32203]_  = A169 & \new_[32202]_ ;
  assign \new_[32206]_  = ~A199 & A166;
  assign \new_[32209]_  = ~A201 & A200;
  assign \new_[32210]_  = \new_[32209]_  & \new_[32206]_ ;
  assign \new_[32211]_  = \new_[32210]_  & \new_[32203]_ ;
  assign \new_[32215]_  = A234 & A233;
  assign \new_[32216]_  = ~A203 & \new_[32215]_ ;
  assign \new_[32219]_  = A299 & ~A298;
  assign \new_[32222]_  = A302 & ~A301;
  assign \new_[32223]_  = \new_[32222]_  & \new_[32219]_ ;
  assign \new_[32224]_  = \new_[32223]_  & \new_[32216]_ ;
  assign \new_[32228]_  = ~A167 & A168;
  assign \new_[32229]_  = A169 & \new_[32228]_ ;
  assign \new_[32232]_  = ~A199 & A166;
  assign \new_[32235]_  = ~A201 & A200;
  assign \new_[32236]_  = \new_[32235]_  & \new_[32232]_ ;
  assign \new_[32237]_  = \new_[32236]_  & \new_[32229]_ ;
  assign \new_[32241]_  = A234 & A233;
  assign \new_[32242]_  = ~A203 & \new_[32241]_ ;
  assign \new_[32245]_  = ~A299 & ~A298;
  assign \new_[32248]_  = ~A302 & A301;
  assign \new_[32249]_  = \new_[32248]_  & \new_[32245]_ ;
  assign \new_[32250]_  = \new_[32249]_  & \new_[32242]_ ;
  assign \new_[32254]_  = ~A167 & A168;
  assign \new_[32255]_  = A169 & \new_[32254]_ ;
  assign \new_[32258]_  = ~A199 & A166;
  assign \new_[32261]_  = ~A201 & A200;
  assign \new_[32262]_  = \new_[32261]_  & \new_[32258]_ ;
  assign \new_[32263]_  = \new_[32262]_  & \new_[32255]_ ;
  assign \new_[32267]_  = A234 & A233;
  assign \new_[32268]_  = ~A203 & \new_[32267]_ ;
  assign \new_[32271]_  = A266 & A265;
  assign \new_[32274]_  = ~A269 & A268;
  assign \new_[32275]_  = \new_[32274]_  & \new_[32271]_ ;
  assign \new_[32276]_  = \new_[32275]_  & \new_[32268]_ ;
  assign \new_[32280]_  = ~A167 & A168;
  assign \new_[32281]_  = A169 & \new_[32280]_ ;
  assign \new_[32284]_  = ~A199 & A166;
  assign \new_[32287]_  = ~A201 & A200;
  assign \new_[32288]_  = \new_[32287]_  & \new_[32284]_ ;
  assign \new_[32289]_  = \new_[32288]_  & \new_[32281]_ ;
  assign \new_[32293]_  = A234 & A233;
  assign \new_[32294]_  = ~A203 & \new_[32293]_ ;
  assign \new_[32297]_  = A266 & ~A265;
  assign \new_[32300]_  = A269 & ~A268;
  assign \new_[32301]_  = \new_[32300]_  & \new_[32297]_ ;
  assign \new_[32302]_  = \new_[32301]_  & \new_[32294]_ ;
  assign \new_[32306]_  = ~A167 & A168;
  assign \new_[32307]_  = A169 & \new_[32306]_ ;
  assign \new_[32310]_  = ~A199 & A166;
  assign \new_[32313]_  = ~A201 & A200;
  assign \new_[32314]_  = \new_[32313]_  & \new_[32310]_ ;
  assign \new_[32315]_  = \new_[32314]_  & \new_[32307]_ ;
  assign \new_[32319]_  = A234 & A233;
  assign \new_[32320]_  = ~A203 & \new_[32319]_ ;
  assign \new_[32323]_  = ~A266 & A265;
  assign \new_[32326]_  = A269 & ~A268;
  assign \new_[32327]_  = \new_[32326]_  & \new_[32323]_ ;
  assign \new_[32328]_  = \new_[32327]_  & \new_[32320]_ ;
  assign \new_[32332]_  = ~A167 & A168;
  assign \new_[32333]_  = A169 & \new_[32332]_ ;
  assign \new_[32336]_  = ~A199 & A166;
  assign \new_[32339]_  = ~A201 & A200;
  assign \new_[32340]_  = \new_[32339]_  & \new_[32336]_ ;
  assign \new_[32341]_  = \new_[32340]_  & \new_[32333]_ ;
  assign \new_[32345]_  = A234 & A233;
  assign \new_[32346]_  = ~A203 & \new_[32345]_ ;
  assign \new_[32349]_  = ~A266 & ~A265;
  assign \new_[32352]_  = ~A269 & A268;
  assign \new_[32353]_  = \new_[32352]_  & \new_[32349]_ ;
  assign \new_[32354]_  = \new_[32353]_  & \new_[32346]_ ;
  assign \new_[32358]_  = ~A167 & A168;
  assign \new_[32359]_  = A169 & \new_[32358]_ ;
  assign \new_[32362]_  = ~A199 & A166;
  assign \new_[32365]_  = ~A201 & A200;
  assign \new_[32366]_  = \new_[32365]_  & \new_[32362]_ ;
  assign \new_[32367]_  = \new_[32366]_  & \new_[32359]_ ;
  assign \new_[32371]_  = A233 & A232;
  assign \new_[32372]_  = ~A203 & \new_[32371]_ ;
  assign \new_[32375]_  = ~A236 & A235;
  assign \new_[32378]_  = A300 & A299;
  assign \new_[32379]_  = \new_[32378]_  & \new_[32375]_ ;
  assign \new_[32380]_  = \new_[32379]_  & \new_[32372]_ ;
  assign \new_[32384]_  = ~A167 & A168;
  assign \new_[32385]_  = A169 & \new_[32384]_ ;
  assign \new_[32388]_  = ~A199 & A166;
  assign \new_[32391]_  = ~A201 & A200;
  assign \new_[32392]_  = \new_[32391]_  & \new_[32388]_ ;
  assign \new_[32393]_  = \new_[32392]_  & \new_[32385]_ ;
  assign \new_[32397]_  = A233 & A232;
  assign \new_[32398]_  = ~A203 & \new_[32397]_ ;
  assign \new_[32401]_  = ~A236 & A235;
  assign \new_[32404]_  = A300 & A298;
  assign \new_[32405]_  = \new_[32404]_  & \new_[32401]_ ;
  assign \new_[32406]_  = \new_[32405]_  & \new_[32398]_ ;
  assign \new_[32410]_  = ~A167 & A168;
  assign \new_[32411]_  = A169 & \new_[32410]_ ;
  assign \new_[32414]_  = ~A199 & A166;
  assign \new_[32417]_  = ~A201 & A200;
  assign \new_[32418]_  = \new_[32417]_  & \new_[32414]_ ;
  assign \new_[32419]_  = \new_[32418]_  & \new_[32411]_ ;
  assign \new_[32423]_  = A233 & A232;
  assign \new_[32424]_  = ~A203 & \new_[32423]_ ;
  assign \new_[32427]_  = ~A236 & A235;
  assign \new_[32430]_  = A267 & A265;
  assign \new_[32431]_  = \new_[32430]_  & \new_[32427]_ ;
  assign \new_[32432]_  = \new_[32431]_  & \new_[32424]_ ;
  assign \new_[32436]_  = ~A167 & A168;
  assign \new_[32437]_  = A169 & \new_[32436]_ ;
  assign \new_[32440]_  = ~A199 & A166;
  assign \new_[32443]_  = ~A201 & A200;
  assign \new_[32444]_  = \new_[32443]_  & \new_[32440]_ ;
  assign \new_[32445]_  = \new_[32444]_  & \new_[32437]_ ;
  assign \new_[32449]_  = A233 & A232;
  assign \new_[32450]_  = ~A203 & \new_[32449]_ ;
  assign \new_[32453]_  = ~A236 & A235;
  assign \new_[32456]_  = A267 & A266;
  assign \new_[32457]_  = \new_[32456]_  & \new_[32453]_ ;
  assign \new_[32458]_  = \new_[32457]_  & \new_[32450]_ ;
  assign \new_[32462]_  = ~A167 & A168;
  assign \new_[32463]_  = A169 & \new_[32462]_ ;
  assign \new_[32466]_  = ~A199 & A166;
  assign \new_[32469]_  = ~A201 & A200;
  assign \new_[32470]_  = \new_[32469]_  & \new_[32466]_ ;
  assign \new_[32471]_  = \new_[32470]_  & \new_[32463]_ ;
  assign \new_[32475]_  = A233 & ~A232;
  assign \new_[32476]_  = ~A203 & \new_[32475]_ ;
  assign \new_[32479]_  = A236 & ~A235;
  assign \new_[32482]_  = A300 & A299;
  assign \new_[32483]_  = \new_[32482]_  & \new_[32479]_ ;
  assign \new_[32484]_  = \new_[32483]_  & \new_[32476]_ ;
  assign \new_[32488]_  = ~A167 & A168;
  assign \new_[32489]_  = A169 & \new_[32488]_ ;
  assign \new_[32492]_  = ~A199 & A166;
  assign \new_[32495]_  = ~A201 & A200;
  assign \new_[32496]_  = \new_[32495]_  & \new_[32492]_ ;
  assign \new_[32497]_  = \new_[32496]_  & \new_[32489]_ ;
  assign \new_[32501]_  = A233 & ~A232;
  assign \new_[32502]_  = ~A203 & \new_[32501]_ ;
  assign \new_[32505]_  = A236 & ~A235;
  assign \new_[32508]_  = A300 & A298;
  assign \new_[32509]_  = \new_[32508]_  & \new_[32505]_ ;
  assign \new_[32510]_  = \new_[32509]_  & \new_[32502]_ ;
  assign \new_[32514]_  = ~A167 & A168;
  assign \new_[32515]_  = A169 & \new_[32514]_ ;
  assign \new_[32518]_  = ~A199 & A166;
  assign \new_[32521]_  = ~A201 & A200;
  assign \new_[32522]_  = \new_[32521]_  & \new_[32518]_ ;
  assign \new_[32523]_  = \new_[32522]_  & \new_[32515]_ ;
  assign \new_[32527]_  = A233 & ~A232;
  assign \new_[32528]_  = ~A203 & \new_[32527]_ ;
  assign \new_[32531]_  = A236 & ~A235;
  assign \new_[32534]_  = A267 & A265;
  assign \new_[32535]_  = \new_[32534]_  & \new_[32531]_ ;
  assign \new_[32536]_  = \new_[32535]_  & \new_[32528]_ ;
  assign \new_[32540]_  = ~A167 & A168;
  assign \new_[32541]_  = A169 & \new_[32540]_ ;
  assign \new_[32544]_  = ~A199 & A166;
  assign \new_[32547]_  = ~A201 & A200;
  assign \new_[32548]_  = \new_[32547]_  & \new_[32544]_ ;
  assign \new_[32549]_  = \new_[32548]_  & \new_[32541]_ ;
  assign \new_[32553]_  = A233 & ~A232;
  assign \new_[32554]_  = ~A203 & \new_[32553]_ ;
  assign \new_[32557]_  = A236 & ~A235;
  assign \new_[32560]_  = A267 & A266;
  assign \new_[32561]_  = \new_[32560]_  & \new_[32557]_ ;
  assign \new_[32562]_  = \new_[32561]_  & \new_[32554]_ ;
  assign \new_[32566]_  = ~A167 & A168;
  assign \new_[32567]_  = A169 & \new_[32566]_ ;
  assign \new_[32570]_  = ~A199 & A166;
  assign \new_[32573]_  = ~A201 & A200;
  assign \new_[32574]_  = \new_[32573]_  & \new_[32570]_ ;
  assign \new_[32575]_  = \new_[32574]_  & \new_[32567]_ ;
  assign \new_[32579]_  = ~A233 & A232;
  assign \new_[32580]_  = ~A203 & \new_[32579]_ ;
  assign \new_[32583]_  = A236 & ~A235;
  assign \new_[32586]_  = A300 & A299;
  assign \new_[32587]_  = \new_[32586]_  & \new_[32583]_ ;
  assign \new_[32588]_  = \new_[32587]_  & \new_[32580]_ ;
  assign \new_[32592]_  = ~A167 & A168;
  assign \new_[32593]_  = A169 & \new_[32592]_ ;
  assign \new_[32596]_  = ~A199 & A166;
  assign \new_[32599]_  = ~A201 & A200;
  assign \new_[32600]_  = \new_[32599]_  & \new_[32596]_ ;
  assign \new_[32601]_  = \new_[32600]_  & \new_[32593]_ ;
  assign \new_[32605]_  = ~A233 & A232;
  assign \new_[32606]_  = ~A203 & \new_[32605]_ ;
  assign \new_[32609]_  = A236 & ~A235;
  assign \new_[32612]_  = A300 & A298;
  assign \new_[32613]_  = \new_[32612]_  & \new_[32609]_ ;
  assign \new_[32614]_  = \new_[32613]_  & \new_[32606]_ ;
  assign \new_[32618]_  = ~A167 & A168;
  assign \new_[32619]_  = A169 & \new_[32618]_ ;
  assign \new_[32622]_  = ~A199 & A166;
  assign \new_[32625]_  = ~A201 & A200;
  assign \new_[32626]_  = \new_[32625]_  & \new_[32622]_ ;
  assign \new_[32627]_  = \new_[32626]_  & \new_[32619]_ ;
  assign \new_[32631]_  = ~A233 & A232;
  assign \new_[32632]_  = ~A203 & \new_[32631]_ ;
  assign \new_[32635]_  = A236 & ~A235;
  assign \new_[32638]_  = A267 & A265;
  assign \new_[32639]_  = \new_[32638]_  & \new_[32635]_ ;
  assign \new_[32640]_  = \new_[32639]_  & \new_[32632]_ ;
  assign \new_[32644]_  = ~A167 & A168;
  assign \new_[32645]_  = A169 & \new_[32644]_ ;
  assign \new_[32648]_  = ~A199 & A166;
  assign \new_[32651]_  = ~A201 & A200;
  assign \new_[32652]_  = \new_[32651]_  & \new_[32648]_ ;
  assign \new_[32653]_  = \new_[32652]_  & \new_[32645]_ ;
  assign \new_[32657]_  = ~A233 & A232;
  assign \new_[32658]_  = ~A203 & \new_[32657]_ ;
  assign \new_[32661]_  = A236 & ~A235;
  assign \new_[32664]_  = A267 & A266;
  assign \new_[32665]_  = \new_[32664]_  & \new_[32661]_ ;
  assign \new_[32666]_  = \new_[32665]_  & \new_[32658]_ ;
  assign \new_[32670]_  = ~A167 & A168;
  assign \new_[32671]_  = A169 & \new_[32670]_ ;
  assign \new_[32674]_  = ~A199 & A166;
  assign \new_[32677]_  = ~A201 & A200;
  assign \new_[32678]_  = \new_[32677]_  & \new_[32674]_ ;
  assign \new_[32679]_  = \new_[32678]_  & \new_[32671]_ ;
  assign \new_[32683]_  = ~A233 & ~A232;
  assign \new_[32684]_  = ~A203 & \new_[32683]_ ;
  assign \new_[32687]_  = ~A236 & A235;
  assign \new_[32690]_  = A300 & A299;
  assign \new_[32691]_  = \new_[32690]_  & \new_[32687]_ ;
  assign \new_[32692]_  = \new_[32691]_  & \new_[32684]_ ;
  assign \new_[32696]_  = ~A167 & A168;
  assign \new_[32697]_  = A169 & \new_[32696]_ ;
  assign \new_[32700]_  = ~A199 & A166;
  assign \new_[32703]_  = ~A201 & A200;
  assign \new_[32704]_  = \new_[32703]_  & \new_[32700]_ ;
  assign \new_[32705]_  = \new_[32704]_  & \new_[32697]_ ;
  assign \new_[32709]_  = ~A233 & ~A232;
  assign \new_[32710]_  = ~A203 & \new_[32709]_ ;
  assign \new_[32713]_  = ~A236 & A235;
  assign \new_[32716]_  = A300 & A298;
  assign \new_[32717]_  = \new_[32716]_  & \new_[32713]_ ;
  assign \new_[32718]_  = \new_[32717]_  & \new_[32710]_ ;
  assign \new_[32722]_  = ~A167 & A168;
  assign \new_[32723]_  = A169 & \new_[32722]_ ;
  assign \new_[32726]_  = ~A199 & A166;
  assign \new_[32729]_  = ~A201 & A200;
  assign \new_[32730]_  = \new_[32729]_  & \new_[32726]_ ;
  assign \new_[32731]_  = \new_[32730]_  & \new_[32723]_ ;
  assign \new_[32735]_  = ~A233 & ~A232;
  assign \new_[32736]_  = ~A203 & \new_[32735]_ ;
  assign \new_[32739]_  = ~A236 & A235;
  assign \new_[32742]_  = A267 & A265;
  assign \new_[32743]_  = \new_[32742]_  & \new_[32739]_ ;
  assign \new_[32744]_  = \new_[32743]_  & \new_[32736]_ ;
  assign \new_[32748]_  = ~A167 & A168;
  assign \new_[32749]_  = A169 & \new_[32748]_ ;
  assign \new_[32752]_  = ~A199 & A166;
  assign \new_[32755]_  = ~A201 & A200;
  assign \new_[32756]_  = \new_[32755]_  & \new_[32752]_ ;
  assign \new_[32757]_  = \new_[32756]_  & \new_[32749]_ ;
  assign \new_[32761]_  = ~A233 & ~A232;
  assign \new_[32762]_  = ~A203 & \new_[32761]_ ;
  assign \new_[32765]_  = ~A236 & A235;
  assign \new_[32768]_  = A267 & A266;
  assign \new_[32769]_  = \new_[32768]_  & \new_[32765]_ ;
  assign \new_[32770]_  = \new_[32769]_  & \new_[32762]_ ;
  assign \new_[32774]_  = ~A167 & A168;
  assign \new_[32775]_  = A169 & \new_[32774]_ ;
  assign \new_[32778]_  = A199 & A166;
  assign \new_[32781]_  = ~A201 & ~A200;
  assign \new_[32782]_  = \new_[32781]_  & \new_[32778]_ ;
  assign \new_[32783]_  = \new_[32782]_  & \new_[32775]_ ;
  assign \new_[32787]_  = A234 & A232;
  assign \new_[32788]_  = A202 & \new_[32787]_ ;
  assign \new_[32791]_  = A299 & A298;
  assign \new_[32794]_  = ~A302 & A301;
  assign \new_[32795]_  = \new_[32794]_  & \new_[32791]_ ;
  assign \new_[32796]_  = \new_[32795]_  & \new_[32788]_ ;
  assign \new_[32800]_  = ~A167 & A168;
  assign \new_[32801]_  = A169 & \new_[32800]_ ;
  assign \new_[32804]_  = A199 & A166;
  assign \new_[32807]_  = ~A201 & ~A200;
  assign \new_[32808]_  = \new_[32807]_  & \new_[32804]_ ;
  assign \new_[32809]_  = \new_[32808]_  & \new_[32801]_ ;
  assign \new_[32813]_  = A234 & A232;
  assign \new_[32814]_  = A202 & \new_[32813]_ ;
  assign \new_[32817]_  = ~A299 & A298;
  assign \new_[32820]_  = A302 & ~A301;
  assign \new_[32821]_  = \new_[32820]_  & \new_[32817]_ ;
  assign \new_[32822]_  = \new_[32821]_  & \new_[32814]_ ;
  assign \new_[32826]_  = ~A167 & A168;
  assign \new_[32827]_  = A169 & \new_[32826]_ ;
  assign \new_[32830]_  = A199 & A166;
  assign \new_[32833]_  = ~A201 & ~A200;
  assign \new_[32834]_  = \new_[32833]_  & \new_[32830]_ ;
  assign \new_[32835]_  = \new_[32834]_  & \new_[32827]_ ;
  assign \new_[32839]_  = A234 & A232;
  assign \new_[32840]_  = A202 & \new_[32839]_ ;
  assign \new_[32843]_  = A299 & ~A298;
  assign \new_[32846]_  = A302 & ~A301;
  assign \new_[32847]_  = \new_[32846]_  & \new_[32843]_ ;
  assign \new_[32848]_  = \new_[32847]_  & \new_[32840]_ ;
  assign \new_[32852]_  = ~A167 & A168;
  assign \new_[32853]_  = A169 & \new_[32852]_ ;
  assign \new_[32856]_  = A199 & A166;
  assign \new_[32859]_  = ~A201 & ~A200;
  assign \new_[32860]_  = \new_[32859]_  & \new_[32856]_ ;
  assign \new_[32861]_  = \new_[32860]_  & \new_[32853]_ ;
  assign \new_[32865]_  = A234 & A232;
  assign \new_[32866]_  = A202 & \new_[32865]_ ;
  assign \new_[32869]_  = ~A299 & ~A298;
  assign \new_[32872]_  = ~A302 & A301;
  assign \new_[32873]_  = \new_[32872]_  & \new_[32869]_ ;
  assign \new_[32874]_  = \new_[32873]_  & \new_[32866]_ ;
  assign \new_[32878]_  = ~A167 & A168;
  assign \new_[32879]_  = A169 & \new_[32878]_ ;
  assign \new_[32882]_  = A199 & A166;
  assign \new_[32885]_  = ~A201 & ~A200;
  assign \new_[32886]_  = \new_[32885]_  & \new_[32882]_ ;
  assign \new_[32887]_  = \new_[32886]_  & \new_[32879]_ ;
  assign \new_[32891]_  = A234 & A232;
  assign \new_[32892]_  = A202 & \new_[32891]_ ;
  assign \new_[32895]_  = A266 & A265;
  assign \new_[32898]_  = ~A269 & A268;
  assign \new_[32899]_  = \new_[32898]_  & \new_[32895]_ ;
  assign \new_[32900]_  = \new_[32899]_  & \new_[32892]_ ;
  assign \new_[32904]_  = ~A167 & A168;
  assign \new_[32905]_  = A169 & \new_[32904]_ ;
  assign \new_[32908]_  = A199 & A166;
  assign \new_[32911]_  = ~A201 & ~A200;
  assign \new_[32912]_  = \new_[32911]_  & \new_[32908]_ ;
  assign \new_[32913]_  = \new_[32912]_  & \new_[32905]_ ;
  assign \new_[32917]_  = A234 & A232;
  assign \new_[32918]_  = A202 & \new_[32917]_ ;
  assign \new_[32921]_  = A266 & ~A265;
  assign \new_[32924]_  = A269 & ~A268;
  assign \new_[32925]_  = \new_[32924]_  & \new_[32921]_ ;
  assign \new_[32926]_  = \new_[32925]_  & \new_[32918]_ ;
  assign \new_[32930]_  = ~A167 & A168;
  assign \new_[32931]_  = A169 & \new_[32930]_ ;
  assign \new_[32934]_  = A199 & A166;
  assign \new_[32937]_  = ~A201 & ~A200;
  assign \new_[32938]_  = \new_[32937]_  & \new_[32934]_ ;
  assign \new_[32939]_  = \new_[32938]_  & \new_[32931]_ ;
  assign \new_[32943]_  = A234 & A232;
  assign \new_[32944]_  = A202 & \new_[32943]_ ;
  assign \new_[32947]_  = ~A266 & A265;
  assign \new_[32950]_  = A269 & ~A268;
  assign \new_[32951]_  = \new_[32950]_  & \new_[32947]_ ;
  assign \new_[32952]_  = \new_[32951]_  & \new_[32944]_ ;
  assign \new_[32956]_  = ~A167 & A168;
  assign \new_[32957]_  = A169 & \new_[32956]_ ;
  assign \new_[32960]_  = A199 & A166;
  assign \new_[32963]_  = ~A201 & ~A200;
  assign \new_[32964]_  = \new_[32963]_  & \new_[32960]_ ;
  assign \new_[32965]_  = \new_[32964]_  & \new_[32957]_ ;
  assign \new_[32969]_  = A234 & A232;
  assign \new_[32970]_  = A202 & \new_[32969]_ ;
  assign \new_[32973]_  = ~A266 & ~A265;
  assign \new_[32976]_  = ~A269 & A268;
  assign \new_[32977]_  = \new_[32976]_  & \new_[32973]_ ;
  assign \new_[32978]_  = \new_[32977]_  & \new_[32970]_ ;
  assign \new_[32982]_  = ~A167 & A168;
  assign \new_[32983]_  = A169 & \new_[32982]_ ;
  assign \new_[32986]_  = A199 & A166;
  assign \new_[32989]_  = ~A201 & ~A200;
  assign \new_[32990]_  = \new_[32989]_  & \new_[32986]_ ;
  assign \new_[32991]_  = \new_[32990]_  & \new_[32983]_ ;
  assign \new_[32995]_  = A234 & A233;
  assign \new_[32996]_  = A202 & \new_[32995]_ ;
  assign \new_[32999]_  = A299 & A298;
  assign \new_[33002]_  = ~A302 & A301;
  assign \new_[33003]_  = \new_[33002]_  & \new_[32999]_ ;
  assign \new_[33004]_  = \new_[33003]_  & \new_[32996]_ ;
  assign \new_[33008]_  = ~A167 & A168;
  assign \new_[33009]_  = A169 & \new_[33008]_ ;
  assign \new_[33012]_  = A199 & A166;
  assign \new_[33015]_  = ~A201 & ~A200;
  assign \new_[33016]_  = \new_[33015]_  & \new_[33012]_ ;
  assign \new_[33017]_  = \new_[33016]_  & \new_[33009]_ ;
  assign \new_[33021]_  = A234 & A233;
  assign \new_[33022]_  = A202 & \new_[33021]_ ;
  assign \new_[33025]_  = ~A299 & A298;
  assign \new_[33028]_  = A302 & ~A301;
  assign \new_[33029]_  = \new_[33028]_  & \new_[33025]_ ;
  assign \new_[33030]_  = \new_[33029]_  & \new_[33022]_ ;
  assign \new_[33034]_  = ~A167 & A168;
  assign \new_[33035]_  = A169 & \new_[33034]_ ;
  assign \new_[33038]_  = A199 & A166;
  assign \new_[33041]_  = ~A201 & ~A200;
  assign \new_[33042]_  = \new_[33041]_  & \new_[33038]_ ;
  assign \new_[33043]_  = \new_[33042]_  & \new_[33035]_ ;
  assign \new_[33047]_  = A234 & A233;
  assign \new_[33048]_  = A202 & \new_[33047]_ ;
  assign \new_[33051]_  = A299 & ~A298;
  assign \new_[33054]_  = A302 & ~A301;
  assign \new_[33055]_  = \new_[33054]_  & \new_[33051]_ ;
  assign \new_[33056]_  = \new_[33055]_  & \new_[33048]_ ;
  assign \new_[33060]_  = ~A167 & A168;
  assign \new_[33061]_  = A169 & \new_[33060]_ ;
  assign \new_[33064]_  = A199 & A166;
  assign \new_[33067]_  = ~A201 & ~A200;
  assign \new_[33068]_  = \new_[33067]_  & \new_[33064]_ ;
  assign \new_[33069]_  = \new_[33068]_  & \new_[33061]_ ;
  assign \new_[33073]_  = A234 & A233;
  assign \new_[33074]_  = A202 & \new_[33073]_ ;
  assign \new_[33077]_  = ~A299 & ~A298;
  assign \new_[33080]_  = ~A302 & A301;
  assign \new_[33081]_  = \new_[33080]_  & \new_[33077]_ ;
  assign \new_[33082]_  = \new_[33081]_  & \new_[33074]_ ;
  assign \new_[33086]_  = ~A167 & A168;
  assign \new_[33087]_  = A169 & \new_[33086]_ ;
  assign \new_[33090]_  = A199 & A166;
  assign \new_[33093]_  = ~A201 & ~A200;
  assign \new_[33094]_  = \new_[33093]_  & \new_[33090]_ ;
  assign \new_[33095]_  = \new_[33094]_  & \new_[33087]_ ;
  assign \new_[33099]_  = A234 & A233;
  assign \new_[33100]_  = A202 & \new_[33099]_ ;
  assign \new_[33103]_  = A266 & A265;
  assign \new_[33106]_  = ~A269 & A268;
  assign \new_[33107]_  = \new_[33106]_  & \new_[33103]_ ;
  assign \new_[33108]_  = \new_[33107]_  & \new_[33100]_ ;
  assign \new_[33112]_  = ~A167 & A168;
  assign \new_[33113]_  = A169 & \new_[33112]_ ;
  assign \new_[33116]_  = A199 & A166;
  assign \new_[33119]_  = ~A201 & ~A200;
  assign \new_[33120]_  = \new_[33119]_  & \new_[33116]_ ;
  assign \new_[33121]_  = \new_[33120]_  & \new_[33113]_ ;
  assign \new_[33125]_  = A234 & A233;
  assign \new_[33126]_  = A202 & \new_[33125]_ ;
  assign \new_[33129]_  = A266 & ~A265;
  assign \new_[33132]_  = A269 & ~A268;
  assign \new_[33133]_  = \new_[33132]_  & \new_[33129]_ ;
  assign \new_[33134]_  = \new_[33133]_  & \new_[33126]_ ;
  assign \new_[33138]_  = ~A167 & A168;
  assign \new_[33139]_  = A169 & \new_[33138]_ ;
  assign \new_[33142]_  = A199 & A166;
  assign \new_[33145]_  = ~A201 & ~A200;
  assign \new_[33146]_  = \new_[33145]_  & \new_[33142]_ ;
  assign \new_[33147]_  = \new_[33146]_  & \new_[33139]_ ;
  assign \new_[33151]_  = A234 & A233;
  assign \new_[33152]_  = A202 & \new_[33151]_ ;
  assign \new_[33155]_  = ~A266 & A265;
  assign \new_[33158]_  = A269 & ~A268;
  assign \new_[33159]_  = \new_[33158]_  & \new_[33155]_ ;
  assign \new_[33160]_  = \new_[33159]_  & \new_[33152]_ ;
  assign \new_[33164]_  = ~A167 & A168;
  assign \new_[33165]_  = A169 & \new_[33164]_ ;
  assign \new_[33168]_  = A199 & A166;
  assign \new_[33171]_  = ~A201 & ~A200;
  assign \new_[33172]_  = \new_[33171]_  & \new_[33168]_ ;
  assign \new_[33173]_  = \new_[33172]_  & \new_[33165]_ ;
  assign \new_[33177]_  = A234 & A233;
  assign \new_[33178]_  = A202 & \new_[33177]_ ;
  assign \new_[33181]_  = ~A266 & ~A265;
  assign \new_[33184]_  = ~A269 & A268;
  assign \new_[33185]_  = \new_[33184]_  & \new_[33181]_ ;
  assign \new_[33186]_  = \new_[33185]_  & \new_[33178]_ ;
  assign \new_[33190]_  = ~A167 & A168;
  assign \new_[33191]_  = A169 & \new_[33190]_ ;
  assign \new_[33194]_  = A199 & A166;
  assign \new_[33197]_  = ~A201 & ~A200;
  assign \new_[33198]_  = \new_[33197]_  & \new_[33194]_ ;
  assign \new_[33199]_  = \new_[33198]_  & \new_[33191]_ ;
  assign \new_[33203]_  = A233 & A232;
  assign \new_[33204]_  = A202 & \new_[33203]_ ;
  assign \new_[33207]_  = ~A236 & A235;
  assign \new_[33210]_  = A300 & A299;
  assign \new_[33211]_  = \new_[33210]_  & \new_[33207]_ ;
  assign \new_[33212]_  = \new_[33211]_  & \new_[33204]_ ;
  assign \new_[33216]_  = ~A167 & A168;
  assign \new_[33217]_  = A169 & \new_[33216]_ ;
  assign \new_[33220]_  = A199 & A166;
  assign \new_[33223]_  = ~A201 & ~A200;
  assign \new_[33224]_  = \new_[33223]_  & \new_[33220]_ ;
  assign \new_[33225]_  = \new_[33224]_  & \new_[33217]_ ;
  assign \new_[33229]_  = A233 & A232;
  assign \new_[33230]_  = A202 & \new_[33229]_ ;
  assign \new_[33233]_  = ~A236 & A235;
  assign \new_[33236]_  = A300 & A298;
  assign \new_[33237]_  = \new_[33236]_  & \new_[33233]_ ;
  assign \new_[33238]_  = \new_[33237]_  & \new_[33230]_ ;
  assign \new_[33242]_  = ~A167 & A168;
  assign \new_[33243]_  = A169 & \new_[33242]_ ;
  assign \new_[33246]_  = A199 & A166;
  assign \new_[33249]_  = ~A201 & ~A200;
  assign \new_[33250]_  = \new_[33249]_  & \new_[33246]_ ;
  assign \new_[33251]_  = \new_[33250]_  & \new_[33243]_ ;
  assign \new_[33255]_  = A233 & A232;
  assign \new_[33256]_  = A202 & \new_[33255]_ ;
  assign \new_[33259]_  = ~A236 & A235;
  assign \new_[33262]_  = A267 & A265;
  assign \new_[33263]_  = \new_[33262]_  & \new_[33259]_ ;
  assign \new_[33264]_  = \new_[33263]_  & \new_[33256]_ ;
  assign \new_[33268]_  = ~A167 & A168;
  assign \new_[33269]_  = A169 & \new_[33268]_ ;
  assign \new_[33272]_  = A199 & A166;
  assign \new_[33275]_  = ~A201 & ~A200;
  assign \new_[33276]_  = \new_[33275]_  & \new_[33272]_ ;
  assign \new_[33277]_  = \new_[33276]_  & \new_[33269]_ ;
  assign \new_[33281]_  = A233 & A232;
  assign \new_[33282]_  = A202 & \new_[33281]_ ;
  assign \new_[33285]_  = ~A236 & A235;
  assign \new_[33288]_  = A267 & A266;
  assign \new_[33289]_  = \new_[33288]_  & \new_[33285]_ ;
  assign \new_[33290]_  = \new_[33289]_  & \new_[33282]_ ;
  assign \new_[33294]_  = ~A167 & A168;
  assign \new_[33295]_  = A169 & \new_[33294]_ ;
  assign \new_[33298]_  = A199 & A166;
  assign \new_[33301]_  = ~A201 & ~A200;
  assign \new_[33302]_  = \new_[33301]_  & \new_[33298]_ ;
  assign \new_[33303]_  = \new_[33302]_  & \new_[33295]_ ;
  assign \new_[33307]_  = A233 & ~A232;
  assign \new_[33308]_  = A202 & \new_[33307]_ ;
  assign \new_[33311]_  = A236 & ~A235;
  assign \new_[33314]_  = A300 & A299;
  assign \new_[33315]_  = \new_[33314]_  & \new_[33311]_ ;
  assign \new_[33316]_  = \new_[33315]_  & \new_[33308]_ ;
  assign \new_[33320]_  = ~A167 & A168;
  assign \new_[33321]_  = A169 & \new_[33320]_ ;
  assign \new_[33324]_  = A199 & A166;
  assign \new_[33327]_  = ~A201 & ~A200;
  assign \new_[33328]_  = \new_[33327]_  & \new_[33324]_ ;
  assign \new_[33329]_  = \new_[33328]_  & \new_[33321]_ ;
  assign \new_[33333]_  = A233 & ~A232;
  assign \new_[33334]_  = A202 & \new_[33333]_ ;
  assign \new_[33337]_  = A236 & ~A235;
  assign \new_[33340]_  = A300 & A298;
  assign \new_[33341]_  = \new_[33340]_  & \new_[33337]_ ;
  assign \new_[33342]_  = \new_[33341]_  & \new_[33334]_ ;
  assign \new_[33346]_  = ~A167 & A168;
  assign \new_[33347]_  = A169 & \new_[33346]_ ;
  assign \new_[33350]_  = A199 & A166;
  assign \new_[33353]_  = ~A201 & ~A200;
  assign \new_[33354]_  = \new_[33353]_  & \new_[33350]_ ;
  assign \new_[33355]_  = \new_[33354]_  & \new_[33347]_ ;
  assign \new_[33359]_  = A233 & ~A232;
  assign \new_[33360]_  = A202 & \new_[33359]_ ;
  assign \new_[33363]_  = A236 & ~A235;
  assign \new_[33366]_  = A267 & A265;
  assign \new_[33367]_  = \new_[33366]_  & \new_[33363]_ ;
  assign \new_[33368]_  = \new_[33367]_  & \new_[33360]_ ;
  assign \new_[33372]_  = ~A167 & A168;
  assign \new_[33373]_  = A169 & \new_[33372]_ ;
  assign \new_[33376]_  = A199 & A166;
  assign \new_[33379]_  = ~A201 & ~A200;
  assign \new_[33380]_  = \new_[33379]_  & \new_[33376]_ ;
  assign \new_[33381]_  = \new_[33380]_  & \new_[33373]_ ;
  assign \new_[33385]_  = A233 & ~A232;
  assign \new_[33386]_  = A202 & \new_[33385]_ ;
  assign \new_[33389]_  = A236 & ~A235;
  assign \new_[33392]_  = A267 & A266;
  assign \new_[33393]_  = \new_[33392]_  & \new_[33389]_ ;
  assign \new_[33394]_  = \new_[33393]_  & \new_[33386]_ ;
  assign \new_[33398]_  = ~A167 & A168;
  assign \new_[33399]_  = A169 & \new_[33398]_ ;
  assign \new_[33402]_  = A199 & A166;
  assign \new_[33405]_  = ~A201 & ~A200;
  assign \new_[33406]_  = \new_[33405]_  & \new_[33402]_ ;
  assign \new_[33407]_  = \new_[33406]_  & \new_[33399]_ ;
  assign \new_[33411]_  = ~A233 & A232;
  assign \new_[33412]_  = A202 & \new_[33411]_ ;
  assign \new_[33415]_  = A236 & ~A235;
  assign \new_[33418]_  = A300 & A299;
  assign \new_[33419]_  = \new_[33418]_  & \new_[33415]_ ;
  assign \new_[33420]_  = \new_[33419]_  & \new_[33412]_ ;
  assign \new_[33424]_  = ~A167 & A168;
  assign \new_[33425]_  = A169 & \new_[33424]_ ;
  assign \new_[33428]_  = A199 & A166;
  assign \new_[33431]_  = ~A201 & ~A200;
  assign \new_[33432]_  = \new_[33431]_  & \new_[33428]_ ;
  assign \new_[33433]_  = \new_[33432]_  & \new_[33425]_ ;
  assign \new_[33437]_  = ~A233 & A232;
  assign \new_[33438]_  = A202 & \new_[33437]_ ;
  assign \new_[33441]_  = A236 & ~A235;
  assign \new_[33444]_  = A300 & A298;
  assign \new_[33445]_  = \new_[33444]_  & \new_[33441]_ ;
  assign \new_[33446]_  = \new_[33445]_  & \new_[33438]_ ;
  assign \new_[33450]_  = ~A167 & A168;
  assign \new_[33451]_  = A169 & \new_[33450]_ ;
  assign \new_[33454]_  = A199 & A166;
  assign \new_[33457]_  = ~A201 & ~A200;
  assign \new_[33458]_  = \new_[33457]_  & \new_[33454]_ ;
  assign \new_[33459]_  = \new_[33458]_  & \new_[33451]_ ;
  assign \new_[33463]_  = ~A233 & A232;
  assign \new_[33464]_  = A202 & \new_[33463]_ ;
  assign \new_[33467]_  = A236 & ~A235;
  assign \new_[33470]_  = A267 & A265;
  assign \new_[33471]_  = \new_[33470]_  & \new_[33467]_ ;
  assign \new_[33472]_  = \new_[33471]_  & \new_[33464]_ ;
  assign \new_[33476]_  = ~A167 & A168;
  assign \new_[33477]_  = A169 & \new_[33476]_ ;
  assign \new_[33480]_  = A199 & A166;
  assign \new_[33483]_  = ~A201 & ~A200;
  assign \new_[33484]_  = \new_[33483]_  & \new_[33480]_ ;
  assign \new_[33485]_  = \new_[33484]_  & \new_[33477]_ ;
  assign \new_[33489]_  = ~A233 & A232;
  assign \new_[33490]_  = A202 & \new_[33489]_ ;
  assign \new_[33493]_  = A236 & ~A235;
  assign \new_[33496]_  = A267 & A266;
  assign \new_[33497]_  = \new_[33496]_  & \new_[33493]_ ;
  assign \new_[33498]_  = \new_[33497]_  & \new_[33490]_ ;
  assign \new_[33502]_  = ~A167 & A168;
  assign \new_[33503]_  = A169 & \new_[33502]_ ;
  assign \new_[33506]_  = A199 & A166;
  assign \new_[33509]_  = ~A201 & ~A200;
  assign \new_[33510]_  = \new_[33509]_  & \new_[33506]_ ;
  assign \new_[33511]_  = \new_[33510]_  & \new_[33503]_ ;
  assign \new_[33515]_  = ~A233 & ~A232;
  assign \new_[33516]_  = A202 & \new_[33515]_ ;
  assign \new_[33519]_  = ~A236 & A235;
  assign \new_[33522]_  = A300 & A299;
  assign \new_[33523]_  = \new_[33522]_  & \new_[33519]_ ;
  assign \new_[33524]_  = \new_[33523]_  & \new_[33516]_ ;
  assign \new_[33528]_  = ~A167 & A168;
  assign \new_[33529]_  = A169 & \new_[33528]_ ;
  assign \new_[33532]_  = A199 & A166;
  assign \new_[33535]_  = ~A201 & ~A200;
  assign \new_[33536]_  = \new_[33535]_  & \new_[33532]_ ;
  assign \new_[33537]_  = \new_[33536]_  & \new_[33529]_ ;
  assign \new_[33541]_  = ~A233 & ~A232;
  assign \new_[33542]_  = A202 & \new_[33541]_ ;
  assign \new_[33545]_  = ~A236 & A235;
  assign \new_[33548]_  = A300 & A298;
  assign \new_[33549]_  = \new_[33548]_  & \new_[33545]_ ;
  assign \new_[33550]_  = \new_[33549]_  & \new_[33542]_ ;
  assign \new_[33554]_  = ~A167 & A168;
  assign \new_[33555]_  = A169 & \new_[33554]_ ;
  assign \new_[33558]_  = A199 & A166;
  assign \new_[33561]_  = ~A201 & ~A200;
  assign \new_[33562]_  = \new_[33561]_  & \new_[33558]_ ;
  assign \new_[33563]_  = \new_[33562]_  & \new_[33555]_ ;
  assign \new_[33567]_  = ~A233 & ~A232;
  assign \new_[33568]_  = A202 & \new_[33567]_ ;
  assign \new_[33571]_  = ~A236 & A235;
  assign \new_[33574]_  = A267 & A265;
  assign \new_[33575]_  = \new_[33574]_  & \new_[33571]_ ;
  assign \new_[33576]_  = \new_[33575]_  & \new_[33568]_ ;
  assign \new_[33580]_  = ~A167 & A168;
  assign \new_[33581]_  = A169 & \new_[33580]_ ;
  assign \new_[33584]_  = A199 & A166;
  assign \new_[33587]_  = ~A201 & ~A200;
  assign \new_[33588]_  = \new_[33587]_  & \new_[33584]_ ;
  assign \new_[33589]_  = \new_[33588]_  & \new_[33581]_ ;
  assign \new_[33593]_  = ~A233 & ~A232;
  assign \new_[33594]_  = A202 & \new_[33593]_ ;
  assign \new_[33597]_  = ~A236 & A235;
  assign \new_[33600]_  = A267 & A266;
  assign \new_[33601]_  = \new_[33600]_  & \new_[33597]_ ;
  assign \new_[33602]_  = \new_[33601]_  & \new_[33594]_ ;
  assign \new_[33606]_  = ~A167 & A168;
  assign \new_[33607]_  = A169 & \new_[33606]_ ;
  assign \new_[33610]_  = A199 & A166;
  assign \new_[33613]_  = ~A201 & ~A200;
  assign \new_[33614]_  = \new_[33613]_  & \new_[33610]_ ;
  assign \new_[33615]_  = \new_[33614]_  & \new_[33607]_ ;
  assign \new_[33619]_  = A234 & A232;
  assign \new_[33620]_  = ~A203 & \new_[33619]_ ;
  assign \new_[33623]_  = A299 & A298;
  assign \new_[33626]_  = ~A302 & A301;
  assign \new_[33627]_  = \new_[33626]_  & \new_[33623]_ ;
  assign \new_[33628]_  = \new_[33627]_  & \new_[33620]_ ;
  assign \new_[33632]_  = ~A167 & A168;
  assign \new_[33633]_  = A169 & \new_[33632]_ ;
  assign \new_[33636]_  = A199 & A166;
  assign \new_[33639]_  = ~A201 & ~A200;
  assign \new_[33640]_  = \new_[33639]_  & \new_[33636]_ ;
  assign \new_[33641]_  = \new_[33640]_  & \new_[33633]_ ;
  assign \new_[33645]_  = A234 & A232;
  assign \new_[33646]_  = ~A203 & \new_[33645]_ ;
  assign \new_[33649]_  = ~A299 & A298;
  assign \new_[33652]_  = A302 & ~A301;
  assign \new_[33653]_  = \new_[33652]_  & \new_[33649]_ ;
  assign \new_[33654]_  = \new_[33653]_  & \new_[33646]_ ;
  assign \new_[33658]_  = ~A167 & A168;
  assign \new_[33659]_  = A169 & \new_[33658]_ ;
  assign \new_[33662]_  = A199 & A166;
  assign \new_[33665]_  = ~A201 & ~A200;
  assign \new_[33666]_  = \new_[33665]_  & \new_[33662]_ ;
  assign \new_[33667]_  = \new_[33666]_  & \new_[33659]_ ;
  assign \new_[33671]_  = A234 & A232;
  assign \new_[33672]_  = ~A203 & \new_[33671]_ ;
  assign \new_[33675]_  = A299 & ~A298;
  assign \new_[33678]_  = A302 & ~A301;
  assign \new_[33679]_  = \new_[33678]_  & \new_[33675]_ ;
  assign \new_[33680]_  = \new_[33679]_  & \new_[33672]_ ;
  assign \new_[33684]_  = ~A167 & A168;
  assign \new_[33685]_  = A169 & \new_[33684]_ ;
  assign \new_[33688]_  = A199 & A166;
  assign \new_[33691]_  = ~A201 & ~A200;
  assign \new_[33692]_  = \new_[33691]_  & \new_[33688]_ ;
  assign \new_[33693]_  = \new_[33692]_  & \new_[33685]_ ;
  assign \new_[33697]_  = A234 & A232;
  assign \new_[33698]_  = ~A203 & \new_[33697]_ ;
  assign \new_[33701]_  = ~A299 & ~A298;
  assign \new_[33704]_  = ~A302 & A301;
  assign \new_[33705]_  = \new_[33704]_  & \new_[33701]_ ;
  assign \new_[33706]_  = \new_[33705]_  & \new_[33698]_ ;
  assign \new_[33710]_  = ~A167 & A168;
  assign \new_[33711]_  = A169 & \new_[33710]_ ;
  assign \new_[33714]_  = A199 & A166;
  assign \new_[33717]_  = ~A201 & ~A200;
  assign \new_[33718]_  = \new_[33717]_  & \new_[33714]_ ;
  assign \new_[33719]_  = \new_[33718]_  & \new_[33711]_ ;
  assign \new_[33723]_  = A234 & A232;
  assign \new_[33724]_  = ~A203 & \new_[33723]_ ;
  assign \new_[33727]_  = A266 & A265;
  assign \new_[33730]_  = ~A269 & A268;
  assign \new_[33731]_  = \new_[33730]_  & \new_[33727]_ ;
  assign \new_[33732]_  = \new_[33731]_  & \new_[33724]_ ;
  assign \new_[33736]_  = ~A167 & A168;
  assign \new_[33737]_  = A169 & \new_[33736]_ ;
  assign \new_[33740]_  = A199 & A166;
  assign \new_[33743]_  = ~A201 & ~A200;
  assign \new_[33744]_  = \new_[33743]_  & \new_[33740]_ ;
  assign \new_[33745]_  = \new_[33744]_  & \new_[33737]_ ;
  assign \new_[33749]_  = A234 & A232;
  assign \new_[33750]_  = ~A203 & \new_[33749]_ ;
  assign \new_[33753]_  = A266 & ~A265;
  assign \new_[33756]_  = A269 & ~A268;
  assign \new_[33757]_  = \new_[33756]_  & \new_[33753]_ ;
  assign \new_[33758]_  = \new_[33757]_  & \new_[33750]_ ;
  assign \new_[33762]_  = ~A167 & A168;
  assign \new_[33763]_  = A169 & \new_[33762]_ ;
  assign \new_[33766]_  = A199 & A166;
  assign \new_[33769]_  = ~A201 & ~A200;
  assign \new_[33770]_  = \new_[33769]_  & \new_[33766]_ ;
  assign \new_[33771]_  = \new_[33770]_  & \new_[33763]_ ;
  assign \new_[33775]_  = A234 & A232;
  assign \new_[33776]_  = ~A203 & \new_[33775]_ ;
  assign \new_[33779]_  = ~A266 & A265;
  assign \new_[33782]_  = A269 & ~A268;
  assign \new_[33783]_  = \new_[33782]_  & \new_[33779]_ ;
  assign \new_[33784]_  = \new_[33783]_  & \new_[33776]_ ;
  assign \new_[33788]_  = ~A167 & A168;
  assign \new_[33789]_  = A169 & \new_[33788]_ ;
  assign \new_[33792]_  = A199 & A166;
  assign \new_[33795]_  = ~A201 & ~A200;
  assign \new_[33796]_  = \new_[33795]_  & \new_[33792]_ ;
  assign \new_[33797]_  = \new_[33796]_  & \new_[33789]_ ;
  assign \new_[33801]_  = A234 & A232;
  assign \new_[33802]_  = ~A203 & \new_[33801]_ ;
  assign \new_[33805]_  = ~A266 & ~A265;
  assign \new_[33808]_  = ~A269 & A268;
  assign \new_[33809]_  = \new_[33808]_  & \new_[33805]_ ;
  assign \new_[33810]_  = \new_[33809]_  & \new_[33802]_ ;
  assign \new_[33814]_  = ~A167 & A168;
  assign \new_[33815]_  = A169 & \new_[33814]_ ;
  assign \new_[33818]_  = A199 & A166;
  assign \new_[33821]_  = ~A201 & ~A200;
  assign \new_[33822]_  = \new_[33821]_  & \new_[33818]_ ;
  assign \new_[33823]_  = \new_[33822]_  & \new_[33815]_ ;
  assign \new_[33827]_  = A234 & A233;
  assign \new_[33828]_  = ~A203 & \new_[33827]_ ;
  assign \new_[33831]_  = A299 & A298;
  assign \new_[33834]_  = ~A302 & A301;
  assign \new_[33835]_  = \new_[33834]_  & \new_[33831]_ ;
  assign \new_[33836]_  = \new_[33835]_  & \new_[33828]_ ;
  assign \new_[33840]_  = ~A167 & A168;
  assign \new_[33841]_  = A169 & \new_[33840]_ ;
  assign \new_[33844]_  = A199 & A166;
  assign \new_[33847]_  = ~A201 & ~A200;
  assign \new_[33848]_  = \new_[33847]_  & \new_[33844]_ ;
  assign \new_[33849]_  = \new_[33848]_  & \new_[33841]_ ;
  assign \new_[33853]_  = A234 & A233;
  assign \new_[33854]_  = ~A203 & \new_[33853]_ ;
  assign \new_[33857]_  = ~A299 & A298;
  assign \new_[33860]_  = A302 & ~A301;
  assign \new_[33861]_  = \new_[33860]_  & \new_[33857]_ ;
  assign \new_[33862]_  = \new_[33861]_  & \new_[33854]_ ;
  assign \new_[33866]_  = ~A167 & A168;
  assign \new_[33867]_  = A169 & \new_[33866]_ ;
  assign \new_[33870]_  = A199 & A166;
  assign \new_[33873]_  = ~A201 & ~A200;
  assign \new_[33874]_  = \new_[33873]_  & \new_[33870]_ ;
  assign \new_[33875]_  = \new_[33874]_  & \new_[33867]_ ;
  assign \new_[33879]_  = A234 & A233;
  assign \new_[33880]_  = ~A203 & \new_[33879]_ ;
  assign \new_[33883]_  = A299 & ~A298;
  assign \new_[33886]_  = A302 & ~A301;
  assign \new_[33887]_  = \new_[33886]_  & \new_[33883]_ ;
  assign \new_[33888]_  = \new_[33887]_  & \new_[33880]_ ;
  assign \new_[33892]_  = ~A167 & A168;
  assign \new_[33893]_  = A169 & \new_[33892]_ ;
  assign \new_[33896]_  = A199 & A166;
  assign \new_[33899]_  = ~A201 & ~A200;
  assign \new_[33900]_  = \new_[33899]_  & \new_[33896]_ ;
  assign \new_[33901]_  = \new_[33900]_  & \new_[33893]_ ;
  assign \new_[33905]_  = A234 & A233;
  assign \new_[33906]_  = ~A203 & \new_[33905]_ ;
  assign \new_[33909]_  = ~A299 & ~A298;
  assign \new_[33912]_  = ~A302 & A301;
  assign \new_[33913]_  = \new_[33912]_  & \new_[33909]_ ;
  assign \new_[33914]_  = \new_[33913]_  & \new_[33906]_ ;
  assign \new_[33918]_  = ~A167 & A168;
  assign \new_[33919]_  = A169 & \new_[33918]_ ;
  assign \new_[33922]_  = A199 & A166;
  assign \new_[33925]_  = ~A201 & ~A200;
  assign \new_[33926]_  = \new_[33925]_  & \new_[33922]_ ;
  assign \new_[33927]_  = \new_[33926]_  & \new_[33919]_ ;
  assign \new_[33931]_  = A234 & A233;
  assign \new_[33932]_  = ~A203 & \new_[33931]_ ;
  assign \new_[33935]_  = A266 & A265;
  assign \new_[33938]_  = ~A269 & A268;
  assign \new_[33939]_  = \new_[33938]_  & \new_[33935]_ ;
  assign \new_[33940]_  = \new_[33939]_  & \new_[33932]_ ;
  assign \new_[33944]_  = ~A167 & A168;
  assign \new_[33945]_  = A169 & \new_[33944]_ ;
  assign \new_[33948]_  = A199 & A166;
  assign \new_[33951]_  = ~A201 & ~A200;
  assign \new_[33952]_  = \new_[33951]_  & \new_[33948]_ ;
  assign \new_[33953]_  = \new_[33952]_  & \new_[33945]_ ;
  assign \new_[33957]_  = A234 & A233;
  assign \new_[33958]_  = ~A203 & \new_[33957]_ ;
  assign \new_[33961]_  = A266 & ~A265;
  assign \new_[33964]_  = A269 & ~A268;
  assign \new_[33965]_  = \new_[33964]_  & \new_[33961]_ ;
  assign \new_[33966]_  = \new_[33965]_  & \new_[33958]_ ;
  assign \new_[33970]_  = ~A167 & A168;
  assign \new_[33971]_  = A169 & \new_[33970]_ ;
  assign \new_[33974]_  = A199 & A166;
  assign \new_[33977]_  = ~A201 & ~A200;
  assign \new_[33978]_  = \new_[33977]_  & \new_[33974]_ ;
  assign \new_[33979]_  = \new_[33978]_  & \new_[33971]_ ;
  assign \new_[33983]_  = A234 & A233;
  assign \new_[33984]_  = ~A203 & \new_[33983]_ ;
  assign \new_[33987]_  = ~A266 & A265;
  assign \new_[33990]_  = A269 & ~A268;
  assign \new_[33991]_  = \new_[33990]_  & \new_[33987]_ ;
  assign \new_[33992]_  = \new_[33991]_  & \new_[33984]_ ;
  assign \new_[33996]_  = ~A167 & A168;
  assign \new_[33997]_  = A169 & \new_[33996]_ ;
  assign \new_[34000]_  = A199 & A166;
  assign \new_[34003]_  = ~A201 & ~A200;
  assign \new_[34004]_  = \new_[34003]_  & \new_[34000]_ ;
  assign \new_[34005]_  = \new_[34004]_  & \new_[33997]_ ;
  assign \new_[34009]_  = A234 & A233;
  assign \new_[34010]_  = ~A203 & \new_[34009]_ ;
  assign \new_[34013]_  = ~A266 & ~A265;
  assign \new_[34016]_  = ~A269 & A268;
  assign \new_[34017]_  = \new_[34016]_  & \new_[34013]_ ;
  assign \new_[34018]_  = \new_[34017]_  & \new_[34010]_ ;
  assign \new_[34022]_  = ~A167 & A168;
  assign \new_[34023]_  = A169 & \new_[34022]_ ;
  assign \new_[34026]_  = A199 & A166;
  assign \new_[34029]_  = ~A201 & ~A200;
  assign \new_[34030]_  = \new_[34029]_  & \new_[34026]_ ;
  assign \new_[34031]_  = \new_[34030]_  & \new_[34023]_ ;
  assign \new_[34035]_  = A233 & A232;
  assign \new_[34036]_  = ~A203 & \new_[34035]_ ;
  assign \new_[34039]_  = ~A236 & A235;
  assign \new_[34042]_  = A300 & A299;
  assign \new_[34043]_  = \new_[34042]_  & \new_[34039]_ ;
  assign \new_[34044]_  = \new_[34043]_  & \new_[34036]_ ;
  assign \new_[34048]_  = ~A167 & A168;
  assign \new_[34049]_  = A169 & \new_[34048]_ ;
  assign \new_[34052]_  = A199 & A166;
  assign \new_[34055]_  = ~A201 & ~A200;
  assign \new_[34056]_  = \new_[34055]_  & \new_[34052]_ ;
  assign \new_[34057]_  = \new_[34056]_  & \new_[34049]_ ;
  assign \new_[34061]_  = A233 & A232;
  assign \new_[34062]_  = ~A203 & \new_[34061]_ ;
  assign \new_[34065]_  = ~A236 & A235;
  assign \new_[34068]_  = A300 & A298;
  assign \new_[34069]_  = \new_[34068]_  & \new_[34065]_ ;
  assign \new_[34070]_  = \new_[34069]_  & \new_[34062]_ ;
  assign \new_[34074]_  = ~A167 & A168;
  assign \new_[34075]_  = A169 & \new_[34074]_ ;
  assign \new_[34078]_  = A199 & A166;
  assign \new_[34081]_  = ~A201 & ~A200;
  assign \new_[34082]_  = \new_[34081]_  & \new_[34078]_ ;
  assign \new_[34083]_  = \new_[34082]_  & \new_[34075]_ ;
  assign \new_[34087]_  = A233 & A232;
  assign \new_[34088]_  = ~A203 & \new_[34087]_ ;
  assign \new_[34091]_  = ~A236 & A235;
  assign \new_[34094]_  = A267 & A265;
  assign \new_[34095]_  = \new_[34094]_  & \new_[34091]_ ;
  assign \new_[34096]_  = \new_[34095]_  & \new_[34088]_ ;
  assign \new_[34100]_  = ~A167 & A168;
  assign \new_[34101]_  = A169 & \new_[34100]_ ;
  assign \new_[34104]_  = A199 & A166;
  assign \new_[34107]_  = ~A201 & ~A200;
  assign \new_[34108]_  = \new_[34107]_  & \new_[34104]_ ;
  assign \new_[34109]_  = \new_[34108]_  & \new_[34101]_ ;
  assign \new_[34113]_  = A233 & A232;
  assign \new_[34114]_  = ~A203 & \new_[34113]_ ;
  assign \new_[34117]_  = ~A236 & A235;
  assign \new_[34120]_  = A267 & A266;
  assign \new_[34121]_  = \new_[34120]_  & \new_[34117]_ ;
  assign \new_[34122]_  = \new_[34121]_  & \new_[34114]_ ;
  assign \new_[34126]_  = ~A167 & A168;
  assign \new_[34127]_  = A169 & \new_[34126]_ ;
  assign \new_[34130]_  = A199 & A166;
  assign \new_[34133]_  = ~A201 & ~A200;
  assign \new_[34134]_  = \new_[34133]_  & \new_[34130]_ ;
  assign \new_[34135]_  = \new_[34134]_  & \new_[34127]_ ;
  assign \new_[34139]_  = A233 & ~A232;
  assign \new_[34140]_  = ~A203 & \new_[34139]_ ;
  assign \new_[34143]_  = A236 & ~A235;
  assign \new_[34146]_  = A300 & A299;
  assign \new_[34147]_  = \new_[34146]_  & \new_[34143]_ ;
  assign \new_[34148]_  = \new_[34147]_  & \new_[34140]_ ;
  assign \new_[34152]_  = ~A167 & A168;
  assign \new_[34153]_  = A169 & \new_[34152]_ ;
  assign \new_[34156]_  = A199 & A166;
  assign \new_[34159]_  = ~A201 & ~A200;
  assign \new_[34160]_  = \new_[34159]_  & \new_[34156]_ ;
  assign \new_[34161]_  = \new_[34160]_  & \new_[34153]_ ;
  assign \new_[34165]_  = A233 & ~A232;
  assign \new_[34166]_  = ~A203 & \new_[34165]_ ;
  assign \new_[34169]_  = A236 & ~A235;
  assign \new_[34172]_  = A300 & A298;
  assign \new_[34173]_  = \new_[34172]_  & \new_[34169]_ ;
  assign \new_[34174]_  = \new_[34173]_  & \new_[34166]_ ;
  assign \new_[34178]_  = ~A167 & A168;
  assign \new_[34179]_  = A169 & \new_[34178]_ ;
  assign \new_[34182]_  = A199 & A166;
  assign \new_[34185]_  = ~A201 & ~A200;
  assign \new_[34186]_  = \new_[34185]_  & \new_[34182]_ ;
  assign \new_[34187]_  = \new_[34186]_  & \new_[34179]_ ;
  assign \new_[34191]_  = A233 & ~A232;
  assign \new_[34192]_  = ~A203 & \new_[34191]_ ;
  assign \new_[34195]_  = A236 & ~A235;
  assign \new_[34198]_  = A267 & A265;
  assign \new_[34199]_  = \new_[34198]_  & \new_[34195]_ ;
  assign \new_[34200]_  = \new_[34199]_  & \new_[34192]_ ;
  assign \new_[34204]_  = ~A167 & A168;
  assign \new_[34205]_  = A169 & \new_[34204]_ ;
  assign \new_[34208]_  = A199 & A166;
  assign \new_[34211]_  = ~A201 & ~A200;
  assign \new_[34212]_  = \new_[34211]_  & \new_[34208]_ ;
  assign \new_[34213]_  = \new_[34212]_  & \new_[34205]_ ;
  assign \new_[34217]_  = A233 & ~A232;
  assign \new_[34218]_  = ~A203 & \new_[34217]_ ;
  assign \new_[34221]_  = A236 & ~A235;
  assign \new_[34224]_  = A267 & A266;
  assign \new_[34225]_  = \new_[34224]_  & \new_[34221]_ ;
  assign \new_[34226]_  = \new_[34225]_  & \new_[34218]_ ;
  assign \new_[34230]_  = ~A167 & A168;
  assign \new_[34231]_  = A169 & \new_[34230]_ ;
  assign \new_[34234]_  = A199 & A166;
  assign \new_[34237]_  = ~A201 & ~A200;
  assign \new_[34238]_  = \new_[34237]_  & \new_[34234]_ ;
  assign \new_[34239]_  = \new_[34238]_  & \new_[34231]_ ;
  assign \new_[34243]_  = ~A233 & A232;
  assign \new_[34244]_  = ~A203 & \new_[34243]_ ;
  assign \new_[34247]_  = A236 & ~A235;
  assign \new_[34250]_  = A300 & A299;
  assign \new_[34251]_  = \new_[34250]_  & \new_[34247]_ ;
  assign \new_[34252]_  = \new_[34251]_  & \new_[34244]_ ;
  assign \new_[34256]_  = ~A167 & A168;
  assign \new_[34257]_  = A169 & \new_[34256]_ ;
  assign \new_[34260]_  = A199 & A166;
  assign \new_[34263]_  = ~A201 & ~A200;
  assign \new_[34264]_  = \new_[34263]_  & \new_[34260]_ ;
  assign \new_[34265]_  = \new_[34264]_  & \new_[34257]_ ;
  assign \new_[34269]_  = ~A233 & A232;
  assign \new_[34270]_  = ~A203 & \new_[34269]_ ;
  assign \new_[34273]_  = A236 & ~A235;
  assign \new_[34276]_  = A300 & A298;
  assign \new_[34277]_  = \new_[34276]_  & \new_[34273]_ ;
  assign \new_[34278]_  = \new_[34277]_  & \new_[34270]_ ;
  assign \new_[34282]_  = ~A167 & A168;
  assign \new_[34283]_  = A169 & \new_[34282]_ ;
  assign \new_[34286]_  = A199 & A166;
  assign \new_[34289]_  = ~A201 & ~A200;
  assign \new_[34290]_  = \new_[34289]_  & \new_[34286]_ ;
  assign \new_[34291]_  = \new_[34290]_  & \new_[34283]_ ;
  assign \new_[34295]_  = ~A233 & A232;
  assign \new_[34296]_  = ~A203 & \new_[34295]_ ;
  assign \new_[34299]_  = A236 & ~A235;
  assign \new_[34302]_  = A267 & A265;
  assign \new_[34303]_  = \new_[34302]_  & \new_[34299]_ ;
  assign \new_[34304]_  = \new_[34303]_  & \new_[34296]_ ;
  assign \new_[34308]_  = ~A167 & A168;
  assign \new_[34309]_  = A169 & \new_[34308]_ ;
  assign \new_[34312]_  = A199 & A166;
  assign \new_[34315]_  = ~A201 & ~A200;
  assign \new_[34316]_  = \new_[34315]_  & \new_[34312]_ ;
  assign \new_[34317]_  = \new_[34316]_  & \new_[34309]_ ;
  assign \new_[34321]_  = ~A233 & A232;
  assign \new_[34322]_  = ~A203 & \new_[34321]_ ;
  assign \new_[34325]_  = A236 & ~A235;
  assign \new_[34328]_  = A267 & A266;
  assign \new_[34329]_  = \new_[34328]_  & \new_[34325]_ ;
  assign \new_[34330]_  = \new_[34329]_  & \new_[34322]_ ;
  assign \new_[34334]_  = ~A167 & A168;
  assign \new_[34335]_  = A169 & \new_[34334]_ ;
  assign \new_[34338]_  = A199 & A166;
  assign \new_[34341]_  = ~A201 & ~A200;
  assign \new_[34342]_  = \new_[34341]_  & \new_[34338]_ ;
  assign \new_[34343]_  = \new_[34342]_  & \new_[34335]_ ;
  assign \new_[34347]_  = ~A233 & ~A232;
  assign \new_[34348]_  = ~A203 & \new_[34347]_ ;
  assign \new_[34351]_  = ~A236 & A235;
  assign \new_[34354]_  = A300 & A299;
  assign \new_[34355]_  = \new_[34354]_  & \new_[34351]_ ;
  assign \new_[34356]_  = \new_[34355]_  & \new_[34348]_ ;
  assign \new_[34360]_  = ~A167 & A168;
  assign \new_[34361]_  = A169 & \new_[34360]_ ;
  assign \new_[34364]_  = A199 & A166;
  assign \new_[34367]_  = ~A201 & ~A200;
  assign \new_[34368]_  = \new_[34367]_  & \new_[34364]_ ;
  assign \new_[34369]_  = \new_[34368]_  & \new_[34361]_ ;
  assign \new_[34373]_  = ~A233 & ~A232;
  assign \new_[34374]_  = ~A203 & \new_[34373]_ ;
  assign \new_[34377]_  = ~A236 & A235;
  assign \new_[34380]_  = A300 & A298;
  assign \new_[34381]_  = \new_[34380]_  & \new_[34377]_ ;
  assign \new_[34382]_  = \new_[34381]_  & \new_[34374]_ ;
  assign \new_[34386]_  = ~A167 & A168;
  assign \new_[34387]_  = A169 & \new_[34386]_ ;
  assign \new_[34390]_  = A199 & A166;
  assign \new_[34393]_  = ~A201 & ~A200;
  assign \new_[34394]_  = \new_[34393]_  & \new_[34390]_ ;
  assign \new_[34395]_  = \new_[34394]_  & \new_[34387]_ ;
  assign \new_[34399]_  = ~A233 & ~A232;
  assign \new_[34400]_  = ~A203 & \new_[34399]_ ;
  assign \new_[34403]_  = ~A236 & A235;
  assign \new_[34406]_  = A267 & A265;
  assign \new_[34407]_  = \new_[34406]_  & \new_[34403]_ ;
  assign \new_[34408]_  = \new_[34407]_  & \new_[34400]_ ;
  assign \new_[34412]_  = ~A167 & A168;
  assign \new_[34413]_  = A169 & \new_[34412]_ ;
  assign \new_[34416]_  = A199 & A166;
  assign \new_[34419]_  = ~A201 & ~A200;
  assign \new_[34420]_  = \new_[34419]_  & \new_[34416]_ ;
  assign \new_[34421]_  = \new_[34420]_  & \new_[34413]_ ;
  assign \new_[34425]_  = ~A233 & ~A232;
  assign \new_[34426]_  = ~A203 & \new_[34425]_ ;
  assign \new_[34429]_  = ~A236 & A235;
  assign \new_[34432]_  = A267 & A266;
  assign \new_[34433]_  = \new_[34432]_  & \new_[34429]_ ;
  assign \new_[34434]_  = \new_[34433]_  & \new_[34426]_ ;
  assign \new_[34438]_  = ~A167 & A168;
  assign \new_[34439]_  = A170 & \new_[34438]_ ;
  assign \new_[34442]_  = ~A199 & A166;
  assign \new_[34445]_  = ~A202 & ~A200;
  assign \new_[34446]_  = \new_[34445]_  & \new_[34442]_ ;
  assign \new_[34447]_  = \new_[34446]_  & \new_[34439]_ ;
  assign \new_[34450]_  = A233 & A232;
  assign \new_[34453]_  = ~A236 & A235;
  assign \new_[34454]_  = \new_[34453]_  & \new_[34450]_ ;
  assign \new_[34457]_  = A299 & A298;
  assign \new_[34460]_  = ~A302 & A301;
  assign \new_[34461]_  = \new_[34460]_  & \new_[34457]_ ;
  assign \new_[34462]_  = \new_[34461]_  & \new_[34454]_ ;
  assign \new_[34466]_  = ~A167 & A168;
  assign \new_[34467]_  = A170 & \new_[34466]_ ;
  assign \new_[34470]_  = ~A199 & A166;
  assign \new_[34473]_  = ~A202 & ~A200;
  assign \new_[34474]_  = \new_[34473]_  & \new_[34470]_ ;
  assign \new_[34475]_  = \new_[34474]_  & \new_[34467]_ ;
  assign \new_[34478]_  = A233 & A232;
  assign \new_[34481]_  = ~A236 & A235;
  assign \new_[34482]_  = \new_[34481]_  & \new_[34478]_ ;
  assign \new_[34485]_  = ~A299 & A298;
  assign \new_[34488]_  = A302 & ~A301;
  assign \new_[34489]_  = \new_[34488]_  & \new_[34485]_ ;
  assign \new_[34490]_  = \new_[34489]_  & \new_[34482]_ ;
  assign \new_[34494]_  = ~A167 & A168;
  assign \new_[34495]_  = A170 & \new_[34494]_ ;
  assign \new_[34498]_  = ~A199 & A166;
  assign \new_[34501]_  = ~A202 & ~A200;
  assign \new_[34502]_  = \new_[34501]_  & \new_[34498]_ ;
  assign \new_[34503]_  = \new_[34502]_  & \new_[34495]_ ;
  assign \new_[34506]_  = A233 & A232;
  assign \new_[34509]_  = ~A236 & A235;
  assign \new_[34510]_  = \new_[34509]_  & \new_[34506]_ ;
  assign \new_[34513]_  = A299 & ~A298;
  assign \new_[34516]_  = A302 & ~A301;
  assign \new_[34517]_  = \new_[34516]_  & \new_[34513]_ ;
  assign \new_[34518]_  = \new_[34517]_  & \new_[34510]_ ;
  assign \new_[34522]_  = ~A167 & A168;
  assign \new_[34523]_  = A170 & \new_[34522]_ ;
  assign \new_[34526]_  = ~A199 & A166;
  assign \new_[34529]_  = ~A202 & ~A200;
  assign \new_[34530]_  = \new_[34529]_  & \new_[34526]_ ;
  assign \new_[34531]_  = \new_[34530]_  & \new_[34523]_ ;
  assign \new_[34534]_  = A233 & A232;
  assign \new_[34537]_  = ~A236 & A235;
  assign \new_[34538]_  = \new_[34537]_  & \new_[34534]_ ;
  assign \new_[34541]_  = ~A299 & ~A298;
  assign \new_[34544]_  = ~A302 & A301;
  assign \new_[34545]_  = \new_[34544]_  & \new_[34541]_ ;
  assign \new_[34546]_  = \new_[34545]_  & \new_[34538]_ ;
  assign \new_[34550]_  = ~A167 & A168;
  assign \new_[34551]_  = A170 & \new_[34550]_ ;
  assign \new_[34554]_  = ~A199 & A166;
  assign \new_[34557]_  = ~A202 & ~A200;
  assign \new_[34558]_  = \new_[34557]_  & \new_[34554]_ ;
  assign \new_[34559]_  = \new_[34558]_  & \new_[34551]_ ;
  assign \new_[34562]_  = A233 & A232;
  assign \new_[34565]_  = ~A236 & A235;
  assign \new_[34566]_  = \new_[34565]_  & \new_[34562]_ ;
  assign \new_[34569]_  = A266 & A265;
  assign \new_[34572]_  = ~A269 & A268;
  assign \new_[34573]_  = \new_[34572]_  & \new_[34569]_ ;
  assign \new_[34574]_  = \new_[34573]_  & \new_[34566]_ ;
  assign \new_[34578]_  = ~A167 & A168;
  assign \new_[34579]_  = A170 & \new_[34578]_ ;
  assign \new_[34582]_  = ~A199 & A166;
  assign \new_[34585]_  = ~A202 & ~A200;
  assign \new_[34586]_  = \new_[34585]_  & \new_[34582]_ ;
  assign \new_[34587]_  = \new_[34586]_  & \new_[34579]_ ;
  assign \new_[34590]_  = A233 & A232;
  assign \new_[34593]_  = ~A236 & A235;
  assign \new_[34594]_  = \new_[34593]_  & \new_[34590]_ ;
  assign \new_[34597]_  = A266 & ~A265;
  assign \new_[34600]_  = A269 & ~A268;
  assign \new_[34601]_  = \new_[34600]_  & \new_[34597]_ ;
  assign \new_[34602]_  = \new_[34601]_  & \new_[34594]_ ;
  assign \new_[34606]_  = ~A167 & A168;
  assign \new_[34607]_  = A170 & \new_[34606]_ ;
  assign \new_[34610]_  = ~A199 & A166;
  assign \new_[34613]_  = ~A202 & ~A200;
  assign \new_[34614]_  = \new_[34613]_  & \new_[34610]_ ;
  assign \new_[34615]_  = \new_[34614]_  & \new_[34607]_ ;
  assign \new_[34618]_  = A233 & A232;
  assign \new_[34621]_  = ~A236 & A235;
  assign \new_[34622]_  = \new_[34621]_  & \new_[34618]_ ;
  assign \new_[34625]_  = ~A266 & A265;
  assign \new_[34628]_  = A269 & ~A268;
  assign \new_[34629]_  = \new_[34628]_  & \new_[34625]_ ;
  assign \new_[34630]_  = \new_[34629]_  & \new_[34622]_ ;
  assign \new_[34634]_  = ~A167 & A168;
  assign \new_[34635]_  = A170 & \new_[34634]_ ;
  assign \new_[34638]_  = ~A199 & A166;
  assign \new_[34641]_  = ~A202 & ~A200;
  assign \new_[34642]_  = \new_[34641]_  & \new_[34638]_ ;
  assign \new_[34643]_  = \new_[34642]_  & \new_[34635]_ ;
  assign \new_[34646]_  = A233 & A232;
  assign \new_[34649]_  = ~A236 & A235;
  assign \new_[34650]_  = \new_[34649]_  & \new_[34646]_ ;
  assign \new_[34653]_  = ~A266 & ~A265;
  assign \new_[34656]_  = ~A269 & A268;
  assign \new_[34657]_  = \new_[34656]_  & \new_[34653]_ ;
  assign \new_[34658]_  = \new_[34657]_  & \new_[34650]_ ;
  assign \new_[34662]_  = ~A167 & A168;
  assign \new_[34663]_  = A170 & \new_[34662]_ ;
  assign \new_[34666]_  = ~A199 & A166;
  assign \new_[34669]_  = ~A202 & ~A200;
  assign \new_[34670]_  = \new_[34669]_  & \new_[34666]_ ;
  assign \new_[34671]_  = \new_[34670]_  & \new_[34663]_ ;
  assign \new_[34674]_  = A233 & ~A232;
  assign \new_[34677]_  = A236 & ~A235;
  assign \new_[34678]_  = \new_[34677]_  & \new_[34674]_ ;
  assign \new_[34681]_  = A299 & A298;
  assign \new_[34684]_  = ~A302 & A301;
  assign \new_[34685]_  = \new_[34684]_  & \new_[34681]_ ;
  assign \new_[34686]_  = \new_[34685]_  & \new_[34678]_ ;
  assign \new_[34690]_  = ~A167 & A168;
  assign \new_[34691]_  = A170 & \new_[34690]_ ;
  assign \new_[34694]_  = ~A199 & A166;
  assign \new_[34697]_  = ~A202 & ~A200;
  assign \new_[34698]_  = \new_[34697]_  & \new_[34694]_ ;
  assign \new_[34699]_  = \new_[34698]_  & \new_[34691]_ ;
  assign \new_[34702]_  = A233 & ~A232;
  assign \new_[34705]_  = A236 & ~A235;
  assign \new_[34706]_  = \new_[34705]_  & \new_[34702]_ ;
  assign \new_[34709]_  = ~A299 & A298;
  assign \new_[34712]_  = A302 & ~A301;
  assign \new_[34713]_  = \new_[34712]_  & \new_[34709]_ ;
  assign \new_[34714]_  = \new_[34713]_  & \new_[34706]_ ;
  assign \new_[34718]_  = ~A167 & A168;
  assign \new_[34719]_  = A170 & \new_[34718]_ ;
  assign \new_[34722]_  = ~A199 & A166;
  assign \new_[34725]_  = ~A202 & ~A200;
  assign \new_[34726]_  = \new_[34725]_  & \new_[34722]_ ;
  assign \new_[34727]_  = \new_[34726]_  & \new_[34719]_ ;
  assign \new_[34730]_  = A233 & ~A232;
  assign \new_[34733]_  = A236 & ~A235;
  assign \new_[34734]_  = \new_[34733]_  & \new_[34730]_ ;
  assign \new_[34737]_  = A299 & ~A298;
  assign \new_[34740]_  = A302 & ~A301;
  assign \new_[34741]_  = \new_[34740]_  & \new_[34737]_ ;
  assign \new_[34742]_  = \new_[34741]_  & \new_[34734]_ ;
  assign \new_[34746]_  = ~A167 & A168;
  assign \new_[34747]_  = A170 & \new_[34746]_ ;
  assign \new_[34750]_  = ~A199 & A166;
  assign \new_[34753]_  = ~A202 & ~A200;
  assign \new_[34754]_  = \new_[34753]_  & \new_[34750]_ ;
  assign \new_[34755]_  = \new_[34754]_  & \new_[34747]_ ;
  assign \new_[34758]_  = A233 & ~A232;
  assign \new_[34761]_  = A236 & ~A235;
  assign \new_[34762]_  = \new_[34761]_  & \new_[34758]_ ;
  assign \new_[34765]_  = ~A299 & ~A298;
  assign \new_[34768]_  = ~A302 & A301;
  assign \new_[34769]_  = \new_[34768]_  & \new_[34765]_ ;
  assign \new_[34770]_  = \new_[34769]_  & \new_[34762]_ ;
  assign \new_[34774]_  = ~A167 & A168;
  assign \new_[34775]_  = A170 & \new_[34774]_ ;
  assign \new_[34778]_  = ~A199 & A166;
  assign \new_[34781]_  = ~A202 & ~A200;
  assign \new_[34782]_  = \new_[34781]_  & \new_[34778]_ ;
  assign \new_[34783]_  = \new_[34782]_  & \new_[34775]_ ;
  assign \new_[34786]_  = A233 & ~A232;
  assign \new_[34789]_  = A236 & ~A235;
  assign \new_[34790]_  = \new_[34789]_  & \new_[34786]_ ;
  assign \new_[34793]_  = A266 & A265;
  assign \new_[34796]_  = ~A269 & A268;
  assign \new_[34797]_  = \new_[34796]_  & \new_[34793]_ ;
  assign \new_[34798]_  = \new_[34797]_  & \new_[34790]_ ;
  assign \new_[34802]_  = ~A167 & A168;
  assign \new_[34803]_  = A170 & \new_[34802]_ ;
  assign \new_[34806]_  = ~A199 & A166;
  assign \new_[34809]_  = ~A202 & ~A200;
  assign \new_[34810]_  = \new_[34809]_  & \new_[34806]_ ;
  assign \new_[34811]_  = \new_[34810]_  & \new_[34803]_ ;
  assign \new_[34814]_  = A233 & ~A232;
  assign \new_[34817]_  = A236 & ~A235;
  assign \new_[34818]_  = \new_[34817]_  & \new_[34814]_ ;
  assign \new_[34821]_  = A266 & ~A265;
  assign \new_[34824]_  = A269 & ~A268;
  assign \new_[34825]_  = \new_[34824]_  & \new_[34821]_ ;
  assign \new_[34826]_  = \new_[34825]_  & \new_[34818]_ ;
  assign \new_[34830]_  = ~A167 & A168;
  assign \new_[34831]_  = A170 & \new_[34830]_ ;
  assign \new_[34834]_  = ~A199 & A166;
  assign \new_[34837]_  = ~A202 & ~A200;
  assign \new_[34838]_  = \new_[34837]_  & \new_[34834]_ ;
  assign \new_[34839]_  = \new_[34838]_  & \new_[34831]_ ;
  assign \new_[34842]_  = A233 & ~A232;
  assign \new_[34845]_  = A236 & ~A235;
  assign \new_[34846]_  = \new_[34845]_  & \new_[34842]_ ;
  assign \new_[34849]_  = ~A266 & A265;
  assign \new_[34852]_  = A269 & ~A268;
  assign \new_[34853]_  = \new_[34852]_  & \new_[34849]_ ;
  assign \new_[34854]_  = \new_[34853]_  & \new_[34846]_ ;
  assign \new_[34858]_  = ~A167 & A168;
  assign \new_[34859]_  = A170 & \new_[34858]_ ;
  assign \new_[34862]_  = ~A199 & A166;
  assign \new_[34865]_  = ~A202 & ~A200;
  assign \new_[34866]_  = \new_[34865]_  & \new_[34862]_ ;
  assign \new_[34867]_  = \new_[34866]_  & \new_[34859]_ ;
  assign \new_[34870]_  = A233 & ~A232;
  assign \new_[34873]_  = A236 & ~A235;
  assign \new_[34874]_  = \new_[34873]_  & \new_[34870]_ ;
  assign \new_[34877]_  = ~A266 & ~A265;
  assign \new_[34880]_  = ~A269 & A268;
  assign \new_[34881]_  = \new_[34880]_  & \new_[34877]_ ;
  assign \new_[34882]_  = \new_[34881]_  & \new_[34874]_ ;
  assign \new_[34886]_  = ~A167 & A168;
  assign \new_[34887]_  = A170 & \new_[34886]_ ;
  assign \new_[34890]_  = ~A199 & A166;
  assign \new_[34893]_  = ~A202 & ~A200;
  assign \new_[34894]_  = \new_[34893]_  & \new_[34890]_ ;
  assign \new_[34895]_  = \new_[34894]_  & \new_[34887]_ ;
  assign \new_[34898]_  = ~A233 & A232;
  assign \new_[34901]_  = A236 & ~A235;
  assign \new_[34902]_  = \new_[34901]_  & \new_[34898]_ ;
  assign \new_[34905]_  = A299 & A298;
  assign \new_[34908]_  = ~A302 & A301;
  assign \new_[34909]_  = \new_[34908]_  & \new_[34905]_ ;
  assign \new_[34910]_  = \new_[34909]_  & \new_[34902]_ ;
  assign \new_[34914]_  = ~A167 & A168;
  assign \new_[34915]_  = A170 & \new_[34914]_ ;
  assign \new_[34918]_  = ~A199 & A166;
  assign \new_[34921]_  = ~A202 & ~A200;
  assign \new_[34922]_  = \new_[34921]_  & \new_[34918]_ ;
  assign \new_[34923]_  = \new_[34922]_  & \new_[34915]_ ;
  assign \new_[34926]_  = ~A233 & A232;
  assign \new_[34929]_  = A236 & ~A235;
  assign \new_[34930]_  = \new_[34929]_  & \new_[34926]_ ;
  assign \new_[34933]_  = ~A299 & A298;
  assign \new_[34936]_  = A302 & ~A301;
  assign \new_[34937]_  = \new_[34936]_  & \new_[34933]_ ;
  assign \new_[34938]_  = \new_[34937]_  & \new_[34930]_ ;
  assign \new_[34942]_  = ~A167 & A168;
  assign \new_[34943]_  = A170 & \new_[34942]_ ;
  assign \new_[34946]_  = ~A199 & A166;
  assign \new_[34949]_  = ~A202 & ~A200;
  assign \new_[34950]_  = \new_[34949]_  & \new_[34946]_ ;
  assign \new_[34951]_  = \new_[34950]_  & \new_[34943]_ ;
  assign \new_[34954]_  = ~A233 & A232;
  assign \new_[34957]_  = A236 & ~A235;
  assign \new_[34958]_  = \new_[34957]_  & \new_[34954]_ ;
  assign \new_[34961]_  = A299 & ~A298;
  assign \new_[34964]_  = A302 & ~A301;
  assign \new_[34965]_  = \new_[34964]_  & \new_[34961]_ ;
  assign \new_[34966]_  = \new_[34965]_  & \new_[34958]_ ;
  assign \new_[34970]_  = ~A167 & A168;
  assign \new_[34971]_  = A170 & \new_[34970]_ ;
  assign \new_[34974]_  = ~A199 & A166;
  assign \new_[34977]_  = ~A202 & ~A200;
  assign \new_[34978]_  = \new_[34977]_  & \new_[34974]_ ;
  assign \new_[34979]_  = \new_[34978]_  & \new_[34971]_ ;
  assign \new_[34982]_  = ~A233 & A232;
  assign \new_[34985]_  = A236 & ~A235;
  assign \new_[34986]_  = \new_[34985]_  & \new_[34982]_ ;
  assign \new_[34989]_  = ~A299 & ~A298;
  assign \new_[34992]_  = ~A302 & A301;
  assign \new_[34993]_  = \new_[34992]_  & \new_[34989]_ ;
  assign \new_[34994]_  = \new_[34993]_  & \new_[34986]_ ;
  assign \new_[34998]_  = ~A167 & A168;
  assign \new_[34999]_  = A170 & \new_[34998]_ ;
  assign \new_[35002]_  = ~A199 & A166;
  assign \new_[35005]_  = ~A202 & ~A200;
  assign \new_[35006]_  = \new_[35005]_  & \new_[35002]_ ;
  assign \new_[35007]_  = \new_[35006]_  & \new_[34999]_ ;
  assign \new_[35010]_  = ~A233 & A232;
  assign \new_[35013]_  = A236 & ~A235;
  assign \new_[35014]_  = \new_[35013]_  & \new_[35010]_ ;
  assign \new_[35017]_  = A266 & A265;
  assign \new_[35020]_  = ~A269 & A268;
  assign \new_[35021]_  = \new_[35020]_  & \new_[35017]_ ;
  assign \new_[35022]_  = \new_[35021]_  & \new_[35014]_ ;
  assign \new_[35026]_  = ~A167 & A168;
  assign \new_[35027]_  = A170 & \new_[35026]_ ;
  assign \new_[35030]_  = ~A199 & A166;
  assign \new_[35033]_  = ~A202 & ~A200;
  assign \new_[35034]_  = \new_[35033]_  & \new_[35030]_ ;
  assign \new_[35035]_  = \new_[35034]_  & \new_[35027]_ ;
  assign \new_[35038]_  = ~A233 & A232;
  assign \new_[35041]_  = A236 & ~A235;
  assign \new_[35042]_  = \new_[35041]_  & \new_[35038]_ ;
  assign \new_[35045]_  = A266 & ~A265;
  assign \new_[35048]_  = A269 & ~A268;
  assign \new_[35049]_  = \new_[35048]_  & \new_[35045]_ ;
  assign \new_[35050]_  = \new_[35049]_  & \new_[35042]_ ;
  assign \new_[35054]_  = ~A167 & A168;
  assign \new_[35055]_  = A170 & \new_[35054]_ ;
  assign \new_[35058]_  = ~A199 & A166;
  assign \new_[35061]_  = ~A202 & ~A200;
  assign \new_[35062]_  = \new_[35061]_  & \new_[35058]_ ;
  assign \new_[35063]_  = \new_[35062]_  & \new_[35055]_ ;
  assign \new_[35066]_  = ~A233 & A232;
  assign \new_[35069]_  = A236 & ~A235;
  assign \new_[35070]_  = \new_[35069]_  & \new_[35066]_ ;
  assign \new_[35073]_  = ~A266 & A265;
  assign \new_[35076]_  = A269 & ~A268;
  assign \new_[35077]_  = \new_[35076]_  & \new_[35073]_ ;
  assign \new_[35078]_  = \new_[35077]_  & \new_[35070]_ ;
  assign \new_[35082]_  = ~A167 & A168;
  assign \new_[35083]_  = A170 & \new_[35082]_ ;
  assign \new_[35086]_  = ~A199 & A166;
  assign \new_[35089]_  = ~A202 & ~A200;
  assign \new_[35090]_  = \new_[35089]_  & \new_[35086]_ ;
  assign \new_[35091]_  = \new_[35090]_  & \new_[35083]_ ;
  assign \new_[35094]_  = ~A233 & A232;
  assign \new_[35097]_  = A236 & ~A235;
  assign \new_[35098]_  = \new_[35097]_  & \new_[35094]_ ;
  assign \new_[35101]_  = ~A266 & ~A265;
  assign \new_[35104]_  = ~A269 & A268;
  assign \new_[35105]_  = \new_[35104]_  & \new_[35101]_ ;
  assign \new_[35106]_  = \new_[35105]_  & \new_[35098]_ ;
  assign \new_[35110]_  = ~A167 & A168;
  assign \new_[35111]_  = A170 & \new_[35110]_ ;
  assign \new_[35114]_  = ~A199 & A166;
  assign \new_[35117]_  = ~A202 & ~A200;
  assign \new_[35118]_  = \new_[35117]_  & \new_[35114]_ ;
  assign \new_[35119]_  = \new_[35118]_  & \new_[35111]_ ;
  assign \new_[35122]_  = ~A233 & ~A232;
  assign \new_[35125]_  = ~A236 & A235;
  assign \new_[35126]_  = \new_[35125]_  & \new_[35122]_ ;
  assign \new_[35129]_  = A299 & A298;
  assign \new_[35132]_  = ~A302 & A301;
  assign \new_[35133]_  = \new_[35132]_  & \new_[35129]_ ;
  assign \new_[35134]_  = \new_[35133]_  & \new_[35126]_ ;
  assign \new_[35138]_  = ~A167 & A168;
  assign \new_[35139]_  = A170 & \new_[35138]_ ;
  assign \new_[35142]_  = ~A199 & A166;
  assign \new_[35145]_  = ~A202 & ~A200;
  assign \new_[35146]_  = \new_[35145]_  & \new_[35142]_ ;
  assign \new_[35147]_  = \new_[35146]_  & \new_[35139]_ ;
  assign \new_[35150]_  = ~A233 & ~A232;
  assign \new_[35153]_  = ~A236 & A235;
  assign \new_[35154]_  = \new_[35153]_  & \new_[35150]_ ;
  assign \new_[35157]_  = ~A299 & A298;
  assign \new_[35160]_  = A302 & ~A301;
  assign \new_[35161]_  = \new_[35160]_  & \new_[35157]_ ;
  assign \new_[35162]_  = \new_[35161]_  & \new_[35154]_ ;
  assign \new_[35166]_  = ~A167 & A168;
  assign \new_[35167]_  = A170 & \new_[35166]_ ;
  assign \new_[35170]_  = ~A199 & A166;
  assign \new_[35173]_  = ~A202 & ~A200;
  assign \new_[35174]_  = \new_[35173]_  & \new_[35170]_ ;
  assign \new_[35175]_  = \new_[35174]_  & \new_[35167]_ ;
  assign \new_[35178]_  = ~A233 & ~A232;
  assign \new_[35181]_  = ~A236 & A235;
  assign \new_[35182]_  = \new_[35181]_  & \new_[35178]_ ;
  assign \new_[35185]_  = A299 & ~A298;
  assign \new_[35188]_  = A302 & ~A301;
  assign \new_[35189]_  = \new_[35188]_  & \new_[35185]_ ;
  assign \new_[35190]_  = \new_[35189]_  & \new_[35182]_ ;
  assign \new_[35194]_  = ~A167 & A168;
  assign \new_[35195]_  = A170 & \new_[35194]_ ;
  assign \new_[35198]_  = ~A199 & A166;
  assign \new_[35201]_  = ~A202 & ~A200;
  assign \new_[35202]_  = \new_[35201]_  & \new_[35198]_ ;
  assign \new_[35203]_  = \new_[35202]_  & \new_[35195]_ ;
  assign \new_[35206]_  = ~A233 & ~A232;
  assign \new_[35209]_  = ~A236 & A235;
  assign \new_[35210]_  = \new_[35209]_  & \new_[35206]_ ;
  assign \new_[35213]_  = ~A299 & ~A298;
  assign \new_[35216]_  = ~A302 & A301;
  assign \new_[35217]_  = \new_[35216]_  & \new_[35213]_ ;
  assign \new_[35218]_  = \new_[35217]_  & \new_[35210]_ ;
  assign \new_[35222]_  = ~A167 & A168;
  assign \new_[35223]_  = A170 & \new_[35222]_ ;
  assign \new_[35226]_  = ~A199 & A166;
  assign \new_[35229]_  = ~A202 & ~A200;
  assign \new_[35230]_  = \new_[35229]_  & \new_[35226]_ ;
  assign \new_[35231]_  = \new_[35230]_  & \new_[35223]_ ;
  assign \new_[35234]_  = ~A233 & ~A232;
  assign \new_[35237]_  = ~A236 & A235;
  assign \new_[35238]_  = \new_[35237]_  & \new_[35234]_ ;
  assign \new_[35241]_  = A266 & A265;
  assign \new_[35244]_  = ~A269 & A268;
  assign \new_[35245]_  = \new_[35244]_  & \new_[35241]_ ;
  assign \new_[35246]_  = \new_[35245]_  & \new_[35238]_ ;
  assign \new_[35250]_  = ~A167 & A168;
  assign \new_[35251]_  = A170 & \new_[35250]_ ;
  assign \new_[35254]_  = ~A199 & A166;
  assign \new_[35257]_  = ~A202 & ~A200;
  assign \new_[35258]_  = \new_[35257]_  & \new_[35254]_ ;
  assign \new_[35259]_  = \new_[35258]_  & \new_[35251]_ ;
  assign \new_[35262]_  = ~A233 & ~A232;
  assign \new_[35265]_  = ~A236 & A235;
  assign \new_[35266]_  = \new_[35265]_  & \new_[35262]_ ;
  assign \new_[35269]_  = A266 & ~A265;
  assign \new_[35272]_  = A269 & ~A268;
  assign \new_[35273]_  = \new_[35272]_  & \new_[35269]_ ;
  assign \new_[35274]_  = \new_[35273]_  & \new_[35266]_ ;
  assign \new_[35278]_  = ~A167 & A168;
  assign \new_[35279]_  = A170 & \new_[35278]_ ;
  assign \new_[35282]_  = ~A199 & A166;
  assign \new_[35285]_  = ~A202 & ~A200;
  assign \new_[35286]_  = \new_[35285]_  & \new_[35282]_ ;
  assign \new_[35287]_  = \new_[35286]_  & \new_[35279]_ ;
  assign \new_[35290]_  = ~A233 & ~A232;
  assign \new_[35293]_  = ~A236 & A235;
  assign \new_[35294]_  = \new_[35293]_  & \new_[35290]_ ;
  assign \new_[35297]_  = ~A266 & A265;
  assign \new_[35300]_  = A269 & ~A268;
  assign \new_[35301]_  = \new_[35300]_  & \new_[35297]_ ;
  assign \new_[35302]_  = \new_[35301]_  & \new_[35294]_ ;
  assign \new_[35306]_  = ~A167 & A168;
  assign \new_[35307]_  = A170 & \new_[35306]_ ;
  assign \new_[35310]_  = ~A199 & A166;
  assign \new_[35313]_  = ~A202 & ~A200;
  assign \new_[35314]_  = \new_[35313]_  & \new_[35310]_ ;
  assign \new_[35315]_  = \new_[35314]_  & \new_[35307]_ ;
  assign \new_[35318]_  = ~A233 & ~A232;
  assign \new_[35321]_  = ~A236 & A235;
  assign \new_[35322]_  = \new_[35321]_  & \new_[35318]_ ;
  assign \new_[35325]_  = ~A266 & ~A265;
  assign \new_[35328]_  = ~A269 & A268;
  assign \new_[35329]_  = \new_[35328]_  & \new_[35325]_ ;
  assign \new_[35330]_  = \new_[35329]_  & \new_[35322]_ ;
  assign \new_[35334]_  = ~A167 & A168;
  assign \new_[35335]_  = A170 & \new_[35334]_ ;
  assign \new_[35338]_  = ~A199 & A166;
  assign \new_[35341]_  = A203 & ~A200;
  assign \new_[35342]_  = \new_[35341]_  & \new_[35338]_ ;
  assign \new_[35343]_  = \new_[35342]_  & \new_[35335]_ ;
  assign \new_[35346]_  = A233 & A232;
  assign \new_[35349]_  = ~A236 & A235;
  assign \new_[35350]_  = \new_[35349]_  & \new_[35346]_ ;
  assign \new_[35353]_  = A299 & A298;
  assign \new_[35356]_  = ~A302 & A301;
  assign \new_[35357]_  = \new_[35356]_  & \new_[35353]_ ;
  assign \new_[35358]_  = \new_[35357]_  & \new_[35350]_ ;
  assign \new_[35362]_  = ~A167 & A168;
  assign \new_[35363]_  = A170 & \new_[35362]_ ;
  assign \new_[35366]_  = ~A199 & A166;
  assign \new_[35369]_  = A203 & ~A200;
  assign \new_[35370]_  = \new_[35369]_  & \new_[35366]_ ;
  assign \new_[35371]_  = \new_[35370]_  & \new_[35363]_ ;
  assign \new_[35374]_  = A233 & A232;
  assign \new_[35377]_  = ~A236 & A235;
  assign \new_[35378]_  = \new_[35377]_  & \new_[35374]_ ;
  assign \new_[35381]_  = ~A299 & A298;
  assign \new_[35384]_  = A302 & ~A301;
  assign \new_[35385]_  = \new_[35384]_  & \new_[35381]_ ;
  assign \new_[35386]_  = \new_[35385]_  & \new_[35378]_ ;
  assign \new_[35390]_  = ~A167 & A168;
  assign \new_[35391]_  = A170 & \new_[35390]_ ;
  assign \new_[35394]_  = ~A199 & A166;
  assign \new_[35397]_  = A203 & ~A200;
  assign \new_[35398]_  = \new_[35397]_  & \new_[35394]_ ;
  assign \new_[35399]_  = \new_[35398]_  & \new_[35391]_ ;
  assign \new_[35402]_  = A233 & A232;
  assign \new_[35405]_  = ~A236 & A235;
  assign \new_[35406]_  = \new_[35405]_  & \new_[35402]_ ;
  assign \new_[35409]_  = A299 & ~A298;
  assign \new_[35412]_  = A302 & ~A301;
  assign \new_[35413]_  = \new_[35412]_  & \new_[35409]_ ;
  assign \new_[35414]_  = \new_[35413]_  & \new_[35406]_ ;
  assign \new_[35418]_  = ~A167 & A168;
  assign \new_[35419]_  = A170 & \new_[35418]_ ;
  assign \new_[35422]_  = ~A199 & A166;
  assign \new_[35425]_  = A203 & ~A200;
  assign \new_[35426]_  = \new_[35425]_  & \new_[35422]_ ;
  assign \new_[35427]_  = \new_[35426]_  & \new_[35419]_ ;
  assign \new_[35430]_  = A233 & A232;
  assign \new_[35433]_  = ~A236 & A235;
  assign \new_[35434]_  = \new_[35433]_  & \new_[35430]_ ;
  assign \new_[35437]_  = ~A299 & ~A298;
  assign \new_[35440]_  = ~A302 & A301;
  assign \new_[35441]_  = \new_[35440]_  & \new_[35437]_ ;
  assign \new_[35442]_  = \new_[35441]_  & \new_[35434]_ ;
  assign \new_[35446]_  = ~A167 & A168;
  assign \new_[35447]_  = A170 & \new_[35446]_ ;
  assign \new_[35450]_  = ~A199 & A166;
  assign \new_[35453]_  = A203 & ~A200;
  assign \new_[35454]_  = \new_[35453]_  & \new_[35450]_ ;
  assign \new_[35455]_  = \new_[35454]_  & \new_[35447]_ ;
  assign \new_[35458]_  = A233 & A232;
  assign \new_[35461]_  = ~A236 & A235;
  assign \new_[35462]_  = \new_[35461]_  & \new_[35458]_ ;
  assign \new_[35465]_  = A266 & A265;
  assign \new_[35468]_  = ~A269 & A268;
  assign \new_[35469]_  = \new_[35468]_  & \new_[35465]_ ;
  assign \new_[35470]_  = \new_[35469]_  & \new_[35462]_ ;
  assign \new_[35474]_  = ~A167 & A168;
  assign \new_[35475]_  = A170 & \new_[35474]_ ;
  assign \new_[35478]_  = ~A199 & A166;
  assign \new_[35481]_  = A203 & ~A200;
  assign \new_[35482]_  = \new_[35481]_  & \new_[35478]_ ;
  assign \new_[35483]_  = \new_[35482]_  & \new_[35475]_ ;
  assign \new_[35486]_  = A233 & A232;
  assign \new_[35489]_  = ~A236 & A235;
  assign \new_[35490]_  = \new_[35489]_  & \new_[35486]_ ;
  assign \new_[35493]_  = A266 & ~A265;
  assign \new_[35496]_  = A269 & ~A268;
  assign \new_[35497]_  = \new_[35496]_  & \new_[35493]_ ;
  assign \new_[35498]_  = \new_[35497]_  & \new_[35490]_ ;
  assign \new_[35502]_  = ~A167 & A168;
  assign \new_[35503]_  = A170 & \new_[35502]_ ;
  assign \new_[35506]_  = ~A199 & A166;
  assign \new_[35509]_  = A203 & ~A200;
  assign \new_[35510]_  = \new_[35509]_  & \new_[35506]_ ;
  assign \new_[35511]_  = \new_[35510]_  & \new_[35503]_ ;
  assign \new_[35514]_  = A233 & A232;
  assign \new_[35517]_  = ~A236 & A235;
  assign \new_[35518]_  = \new_[35517]_  & \new_[35514]_ ;
  assign \new_[35521]_  = ~A266 & A265;
  assign \new_[35524]_  = A269 & ~A268;
  assign \new_[35525]_  = \new_[35524]_  & \new_[35521]_ ;
  assign \new_[35526]_  = \new_[35525]_  & \new_[35518]_ ;
  assign \new_[35530]_  = ~A167 & A168;
  assign \new_[35531]_  = A170 & \new_[35530]_ ;
  assign \new_[35534]_  = ~A199 & A166;
  assign \new_[35537]_  = A203 & ~A200;
  assign \new_[35538]_  = \new_[35537]_  & \new_[35534]_ ;
  assign \new_[35539]_  = \new_[35538]_  & \new_[35531]_ ;
  assign \new_[35542]_  = A233 & A232;
  assign \new_[35545]_  = ~A236 & A235;
  assign \new_[35546]_  = \new_[35545]_  & \new_[35542]_ ;
  assign \new_[35549]_  = ~A266 & ~A265;
  assign \new_[35552]_  = ~A269 & A268;
  assign \new_[35553]_  = \new_[35552]_  & \new_[35549]_ ;
  assign \new_[35554]_  = \new_[35553]_  & \new_[35546]_ ;
  assign \new_[35558]_  = ~A167 & A168;
  assign \new_[35559]_  = A170 & \new_[35558]_ ;
  assign \new_[35562]_  = ~A199 & A166;
  assign \new_[35565]_  = A203 & ~A200;
  assign \new_[35566]_  = \new_[35565]_  & \new_[35562]_ ;
  assign \new_[35567]_  = \new_[35566]_  & \new_[35559]_ ;
  assign \new_[35570]_  = A233 & ~A232;
  assign \new_[35573]_  = A236 & ~A235;
  assign \new_[35574]_  = \new_[35573]_  & \new_[35570]_ ;
  assign \new_[35577]_  = A299 & A298;
  assign \new_[35580]_  = ~A302 & A301;
  assign \new_[35581]_  = \new_[35580]_  & \new_[35577]_ ;
  assign \new_[35582]_  = \new_[35581]_  & \new_[35574]_ ;
  assign \new_[35586]_  = ~A167 & A168;
  assign \new_[35587]_  = A170 & \new_[35586]_ ;
  assign \new_[35590]_  = ~A199 & A166;
  assign \new_[35593]_  = A203 & ~A200;
  assign \new_[35594]_  = \new_[35593]_  & \new_[35590]_ ;
  assign \new_[35595]_  = \new_[35594]_  & \new_[35587]_ ;
  assign \new_[35598]_  = A233 & ~A232;
  assign \new_[35601]_  = A236 & ~A235;
  assign \new_[35602]_  = \new_[35601]_  & \new_[35598]_ ;
  assign \new_[35605]_  = ~A299 & A298;
  assign \new_[35608]_  = A302 & ~A301;
  assign \new_[35609]_  = \new_[35608]_  & \new_[35605]_ ;
  assign \new_[35610]_  = \new_[35609]_  & \new_[35602]_ ;
  assign \new_[35614]_  = ~A167 & A168;
  assign \new_[35615]_  = A170 & \new_[35614]_ ;
  assign \new_[35618]_  = ~A199 & A166;
  assign \new_[35621]_  = A203 & ~A200;
  assign \new_[35622]_  = \new_[35621]_  & \new_[35618]_ ;
  assign \new_[35623]_  = \new_[35622]_  & \new_[35615]_ ;
  assign \new_[35626]_  = A233 & ~A232;
  assign \new_[35629]_  = A236 & ~A235;
  assign \new_[35630]_  = \new_[35629]_  & \new_[35626]_ ;
  assign \new_[35633]_  = A299 & ~A298;
  assign \new_[35636]_  = A302 & ~A301;
  assign \new_[35637]_  = \new_[35636]_  & \new_[35633]_ ;
  assign \new_[35638]_  = \new_[35637]_  & \new_[35630]_ ;
  assign \new_[35642]_  = ~A167 & A168;
  assign \new_[35643]_  = A170 & \new_[35642]_ ;
  assign \new_[35646]_  = ~A199 & A166;
  assign \new_[35649]_  = A203 & ~A200;
  assign \new_[35650]_  = \new_[35649]_  & \new_[35646]_ ;
  assign \new_[35651]_  = \new_[35650]_  & \new_[35643]_ ;
  assign \new_[35654]_  = A233 & ~A232;
  assign \new_[35657]_  = A236 & ~A235;
  assign \new_[35658]_  = \new_[35657]_  & \new_[35654]_ ;
  assign \new_[35661]_  = ~A299 & ~A298;
  assign \new_[35664]_  = ~A302 & A301;
  assign \new_[35665]_  = \new_[35664]_  & \new_[35661]_ ;
  assign \new_[35666]_  = \new_[35665]_  & \new_[35658]_ ;
  assign \new_[35670]_  = ~A167 & A168;
  assign \new_[35671]_  = A170 & \new_[35670]_ ;
  assign \new_[35674]_  = ~A199 & A166;
  assign \new_[35677]_  = A203 & ~A200;
  assign \new_[35678]_  = \new_[35677]_  & \new_[35674]_ ;
  assign \new_[35679]_  = \new_[35678]_  & \new_[35671]_ ;
  assign \new_[35682]_  = A233 & ~A232;
  assign \new_[35685]_  = A236 & ~A235;
  assign \new_[35686]_  = \new_[35685]_  & \new_[35682]_ ;
  assign \new_[35689]_  = A266 & A265;
  assign \new_[35692]_  = ~A269 & A268;
  assign \new_[35693]_  = \new_[35692]_  & \new_[35689]_ ;
  assign \new_[35694]_  = \new_[35693]_  & \new_[35686]_ ;
  assign \new_[35698]_  = ~A167 & A168;
  assign \new_[35699]_  = A170 & \new_[35698]_ ;
  assign \new_[35702]_  = ~A199 & A166;
  assign \new_[35705]_  = A203 & ~A200;
  assign \new_[35706]_  = \new_[35705]_  & \new_[35702]_ ;
  assign \new_[35707]_  = \new_[35706]_  & \new_[35699]_ ;
  assign \new_[35710]_  = A233 & ~A232;
  assign \new_[35713]_  = A236 & ~A235;
  assign \new_[35714]_  = \new_[35713]_  & \new_[35710]_ ;
  assign \new_[35717]_  = A266 & ~A265;
  assign \new_[35720]_  = A269 & ~A268;
  assign \new_[35721]_  = \new_[35720]_  & \new_[35717]_ ;
  assign \new_[35722]_  = \new_[35721]_  & \new_[35714]_ ;
  assign \new_[35726]_  = ~A167 & A168;
  assign \new_[35727]_  = A170 & \new_[35726]_ ;
  assign \new_[35730]_  = ~A199 & A166;
  assign \new_[35733]_  = A203 & ~A200;
  assign \new_[35734]_  = \new_[35733]_  & \new_[35730]_ ;
  assign \new_[35735]_  = \new_[35734]_  & \new_[35727]_ ;
  assign \new_[35738]_  = A233 & ~A232;
  assign \new_[35741]_  = A236 & ~A235;
  assign \new_[35742]_  = \new_[35741]_  & \new_[35738]_ ;
  assign \new_[35745]_  = ~A266 & A265;
  assign \new_[35748]_  = A269 & ~A268;
  assign \new_[35749]_  = \new_[35748]_  & \new_[35745]_ ;
  assign \new_[35750]_  = \new_[35749]_  & \new_[35742]_ ;
  assign \new_[35754]_  = ~A167 & A168;
  assign \new_[35755]_  = A170 & \new_[35754]_ ;
  assign \new_[35758]_  = ~A199 & A166;
  assign \new_[35761]_  = A203 & ~A200;
  assign \new_[35762]_  = \new_[35761]_  & \new_[35758]_ ;
  assign \new_[35763]_  = \new_[35762]_  & \new_[35755]_ ;
  assign \new_[35766]_  = A233 & ~A232;
  assign \new_[35769]_  = A236 & ~A235;
  assign \new_[35770]_  = \new_[35769]_  & \new_[35766]_ ;
  assign \new_[35773]_  = ~A266 & ~A265;
  assign \new_[35776]_  = ~A269 & A268;
  assign \new_[35777]_  = \new_[35776]_  & \new_[35773]_ ;
  assign \new_[35778]_  = \new_[35777]_  & \new_[35770]_ ;
  assign \new_[35782]_  = ~A167 & A168;
  assign \new_[35783]_  = A170 & \new_[35782]_ ;
  assign \new_[35786]_  = ~A199 & A166;
  assign \new_[35789]_  = A203 & ~A200;
  assign \new_[35790]_  = \new_[35789]_  & \new_[35786]_ ;
  assign \new_[35791]_  = \new_[35790]_  & \new_[35783]_ ;
  assign \new_[35794]_  = ~A233 & A232;
  assign \new_[35797]_  = A236 & ~A235;
  assign \new_[35798]_  = \new_[35797]_  & \new_[35794]_ ;
  assign \new_[35801]_  = A299 & A298;
  assign \new_[35804]_  = ~A302 & A301;
  assign \new_[35805]_  = \new_[35804]_  & \new_[35801]_ ;
  assign \new_[35806]_  = \new_[35805]_  & \new_[35798]_ ;
  assign \new_[35810]_  = ~A167 & A168;
  assign \new_[35811]_  = A170 & \new_[35810]_ ;
  assign \new_[35814]_  = ~A199 & A166;
  assign \new_[35817]_  = A203 & ~A200;
  assign \new_[35818]_  = \new_[35817]_  & \new_[35814]_ ;
  assign \new_[35819]_  = \new_[35818]_  & \new_[35811]_ ;
  assign \new_[35822]_  = ~A233 & A232;
  assign \new_[35825]_  = A236 & ~A235;
  assign \new_[35826]_  = \new_[35825]_  & \new_[35822]_ ;
  assign \new_[35829]_  = ~A299 & A298;
  assign \new_[35832]_  = A302 & ~A301;
  assign \new_[35833]_  = \new_[35832]_  & \new_[35829]_ ;
  assign \new_[35834]_  = \new_[35833]_  & \new_[35826]_ ;
  assign \new_[35838]_  = ~A167 & A168;
  assign \new_[35839]_  = A170 & \new_[35838]_ ;
  assign \new_[35842]_  = ~A199 & A166;
  assign \new_[35845]_  = A203 & ~A200;
  assign \new_[35846]_  = \new_[35845]_  & \new_[35842]_ ;
  assign \new_[35847]_  = \new_[35846]_  & \new_[35839]_ ;
  assign \new_[35850]_  = ~A233 & A232;
  assign \new_[35853]_  = A236 & ~A235;
  assign \new_[35854]_  = \new_[35853]_  & \new_[35850]_ ;
  assign \new_[35857]_  = A299 & ~A298;
  assign \new_[35860]_  = A302 & ~A301;
  assign \new_[35861]_  = \new_[35860]_  & \new_[35857]_ ;
  assign \new_[35862]_  = \new_[35861]_  & \new_[35854]_ ;
  assign \new_[35866]_  = ~A167 & A168;
  assign \new_[35867]_  = A170 & \new_[35866]_ ;
  assign \new_[35870]_  = ~A199 & A166;
  assign \new_[35873]_  = A203 & ~A200;
  assign \new_[35874]_  = \new_[35873]_  & \new_[35870]_ ;
  assign \new_[35875]_  = \new_[35874]_  & \new_[35867]_ ;
  assign \new_[35878]_  = ~A233 & A232;
  assign \new_[35881]_  = A236 & ~A235;
  assign \new_[35882]_  = \new_[35881]_  & \new_[35878]_ ;
  assign \new_[35885]_  = ~A299 & ~A298;
  assign \new_[35888]_  = ~A302 & A301;
  assign \new_[35889]_  = \new_[35888]_  & \new_[35885]_ ;
  assign \new_[35890]_  = \new_[35889]_  & \new_[35882]_ ;
  assign \new_[35894]_  = ~A167 & A168;
  assign \new_[35895]_  = A170 & \new_[35894]_ ;
  assign \new_[35898]_  = ~A199 & A166;
  assign \new_[35901]_  = A203 & ~A200;
  assign \new_[35902]_  = \new_[35901]_  & \new_[35898]_ ;
  assign \new_[35903]_  = \new_[35902]_  & \new_[35895]_ ;
  assign \new_[35906]_  = ~A233 & A232;
  assign \new_[35909]_  = A236 & ~A235;
  assign \new_[35910]_  = \new_[35909]_  & \new_[35906]_ ;
  assign \new_[35913]_  = A266 & A265;
  assign \new_[35916]_  = ~A269 & A268;
  assign \new_[35917]_  = \new_[35916]_  & \new_[35913]_ ;
  assign \new_[35918]_  = \new_[35917]_  & \new_[35910]_ ;
  assign \new_[35922]_  = ~A167 & A168;
  assign \new_[35923]_  = A170 & \new_[35922]_ ;
  assign \new_[35926]_  = ~A199 & A166;
  assign \new_[35929]_  = A203 & ~A200;
  assign \new_[35930]_  = \new_[35929]_  & \new_[35926]_ ;
  assign \new_[35931]_  = \new_[35930]_  & \new_[35923]_ ;
  assign \new_[35934]_  = ~A233 & A232;
  assign \new_[35937]_  = A236 & ~A235;
  assign \new_[35938]_  = \new_[35937]_  & \new_[35934]_ ;
  assign \new_[35941]_  = A266 & ~A265;
  assign \new_[35944]_  = A269 & ~A268;
  assign \new_[35945]_  = \new_[35944]_  & \new_[35941]_ ;
  assign \new_[35946]_  = \new_[35945]_  & \new_[35938]_ ;
  assign \new_[35950]_  = ~A167 & A168;
  assign \new_[35951]_  = A170 & \new_[35950]_ ;
  assign \new_[35954]_  = ~A199 & A166;
  assign \new_[35957]_  = A203 & ~A200;
  assign \new_[35958]_  = \new_[35957]_  & \new_[35954]_ ;
  assign \new_[35959]_  = \new_[35958]_  & \new_[35951]_ ;
  assign \new_[35962]_  = ~A233 & A232;
  assign \new_[35965]_  = A236 & ~A235;
  assign \new_[35966]_  = \new_[35965]_  & \new_[35962]_ ;
  assign \new_[35969]_  = ~A266 & A265;
  assign \new_[35972]_  = A269 & ~A268;
  assign \new_[35973]_  = \new_[35972]_  & \new_[35969]_ ;
  assign \new_[35974]_  = \new_[35973]_  & \new_[35966]_ ;
  assign \new_[35978]_  = ~A167 & A168;
  assign \new_[35979]_  = A170 & \new_[35978]_ ;
  assign \new_[35982]_  = ~A199 & A166;
  assign \new_[35985]_  = A203 & ~A200;
  assign \new_[35986]_  = \new_[35985]_  & \new_[35982]_ ;
  assign \new_[35987]_  = \new_[35986]_  & \new_[35979]_ ;
  assign \new_[35990]_  = ~A233 & A232;
  assign \new_[35993]_  = A236 & ~A235;
  assign \new_[35994]_  = \new_[35993]_  & \new_[35990]_ ;
  assign \new_[35997]_  = ~A266 & ~A265;
  assign \new_[36000]_  = ~A269 & A268;
  assign \new_[36001]_  = \new_[36000]_  & \new_[35997]_ ;
  assign \new_[36002]_  = \new_[36001]_  & \new_[35994]_ ;
  assign \new_[36006]_  = ~A167 & A168;
  assign \new_[36007]_  = A170 & \new_[36006]_ ;
  assign \new_[36010]_  = ~A199 & A166;
  assign \new_[36013]_  = A203 & ~A200;
  assign \new_[36014]_  = \new_[36013]_  & \new_[36010]_ ;
  assign \new_[36015]_  = \new_[36014]_  & \new_[36007]_ ;
  assign \new_[36018]_  = ~A233 & ~A232;
  assign \new_[36021]_  = ~A236 & A235;
  assign \new_[36022]_  = \new_[36021]_  & \new_[36018]_ ;
  assign \new_[36025]_  = A299 & A298;
  assign \new_[36028]_  = ~A302 & A301;
  assign \new_[36029]_  = \new_[36028]_  & \new_[36025]_ ;
  assign \new_[36030]_  = \new_[36029]_  & \new_[36022]_ ;
  assign \new_[36034]_  = ~A167 & A168;
  assign \new_[36035]_  = A170 & \new_[36034]_ ;
  assign \new_[36038]_  = ~A199 & A166;
  assign \new_[36041]_  = A203 & ~A200;
  assign \new_[36042]_  = \new_[36041]_  & \new_[36038]_ ;
  assign \new_[36043]_  = \new_[36042]_  & \new_[36035]_ ;
  assign \new_[36046]_  = ~A233 & ~A232;
  assign \new_[36049]_  = ~A236 & A235;
  assign \new_[36050]_  = \new_[36049]_  & \new_[36046]_ ;
  assign \new_[36053]_  = ~A299 & A298;
  assign \new_[36056]_  = A302 & ~A301;
  assign \new_[36057]_  = \new_[36056]_  & \new_[36053]_ ;
  assign \new_[36058]_  = \new_[36057]_  & \new_[36050]_ ;
  assign \new_[36062]_  = ~A167 & A168;
  assign \new_[36063]_  = A170 & \new_[36062]_ ;
  assign \new_[36066]_  = ~A199 & A166;
  assign \new_[36069]_  = A203 & ~A200;
  assign \new_[36070]_  = \new_[36069]_  & \new_[36066]_ ;
  assign \new_[36071]_  = \new_[36070]_  & \new_[36063]_ ;
  assign \new_[36074]_  = ~A233 & ~A232;
  assign \new_[36077]_  = ~A236 & A235;
  assign \new_[36078]_  = \new_[36077]_  & \new_[36074]_ ;
  assign \new_[36081]_  = A299 & ~A298;
  assign \new_[36084]_  = A302 & ~A301;
  assign \new_[36085]_  = \new_[36084]_  & \new_[36081]_ ;
  assign \new_[36086]_  = \new_[36085]_  & \new_[36078]_ ;
  assign \new_[36090]_  = ~A167 & A168;
  assign \new_[36091]_  = A170 & \new_[36090]_ ;
  assign \new_[36094]_  = ~A199 & A166;
  assign \new_[36097]_  = A203 & ~A200;
  assign \new_[36098]_  = \new_[36097]_  & \new_[36094]_ ;
  assign \new_[36099]_  = \new_[36098]_  & \new_[36091]_ ;
  assign \new_[36102]_  = ~A233 & ~A232;
  assign \new_[36105]_  = ~A236 & A235;
  assign \new_[36106]_  = \new_[36105]_  & \new_[36102]_ ;
  assign \new_[36109]_  = ~A299 & ~A298;
  assign \new_[36112]_  = ~A302 & A301;
  assign \new_[36113]_  = \new_[36112]_  & \new_[36109]_ ;
  assign \new_[36114]_  = \new_[36113]_  & \new_[36106]_ ;
  assign \new_[36118]_  = ~A167 & A168;
  assign \new_[36119]_  = A170 & \new_[36118]_ ;
  assign \new_[36122]_  = ~A199 & A166;
  assign \new_[36125]_  = A203 & ~A200;
  assign \new_[36126]_  = \new_[36125]_  & \new_[36122]_ ;
  assign \new_[36127]_  = \new_[36126]_  & \new_[36119]_ ;
  assign \new_[36130]_  = ~A233 & ~A232;
  assign \new_[36133]_  = ~A236 & A235;
  assign \new_[36134]_  = \new_[36133]_  & \new_[36130]_ ;
  assign \new_[36137]_  = A266 & A265;
  assign \new_[36140]_  = ~A269 & A268;
  assign \new_[36141]_  = \new_[36140]_  & \new_[36137]_ ;
  assign \new_[36142]_  = \new_[36141]_  & \new_[36134]_ ;
  assign \new_[36146]_  = ~A167 & A168;
  assign \new_[36147]_  = A170 & \new_[36146]_ ;
  assign \new_[36150]_  = ~A199 & A166;
  assign \new_[36153]_  = A203 & ~A200;
  assign \new_[36154]_  = \new_[36153]_  & \new_[36150]_ ;
  assign \new_[36155]_  = \new_[36154]_  & \new_[36147]_ ;
  assign \new_[36158]_  = ~A233 & ~A232;
  assign \new_[36161]_  = ~A236 & A235;
  assign \new_[36162]_  = \new_[36161]_  & \new_[36158]_ ;
  assign \new_[36165]_  = A266 & ~A265;
  assign \new_[36168]_  = A269 & ~A268;
  assign \new_[36169]_  = \new_[36168]_  & \new_[36165]_ ;
  assign \new_[36170]_  = \new_[36169]_  & \new_[36162]_ ;
  assign \new_[36174]_  = ~A167 & A168;
  assign \new_[36175]_  = A170 & \new_[36174]_ ;
  assign \new_[36178]_  = ~A199 & A166;
  assign \new_[36181]_  = A203 & ~A200;
  assign \new_[36182]_  = \new_[36181]_  & \new_[36178]_ ;
  assign \new_[36183]_  = \new_[36182]_  & \new_[36175]_ ;
  assign \new_[36186]_  = ~A233 & ~A232;
  assign \new_[36189]_  = ~A236 & A235;
  assign \new_[36190]_  = \new_[36189]_  & \new_[36186]_ ;
  assign \new_[36193]_  = ~A266 & A265;
  assign \new_[36196]_  = A269 & ~A268;
  assign \new_[36197]_  = \new_[36196]_  & \new_[36193]_ ;
  assign \new_[36198]_  = \new_[36197]_  & \new_[36190]_ ;
  assign \new_[36202]_  = ~A167 & A168;
  assign \new_[36203]_  = A170 & \new_[36202]_ ;
  assign \new_[36206]_  = ~A199 & A166;
  assign \new_[36209]_  = A203 & ~A200;
  assign \new_[36210]_  = \new_[36209]_  & \new_[36206]_ ;
  assign \new_[36211]_  = \new_[36210]_  & \new_[36203]_ ;
  assign \new_[36214]_  = ~A233 & ~A232;
  assign \new_[36217]_  = ~A236 & A235;
  assign \new_[36218]_  = \new_[36217]_  & \new_[36214]_ ;
  assign \new_[36221]_  = ~A266 & ~A265;
  assign \new_[36224]_  = ~A269 & A268;
  assign \new_[36225]_  = \new_[36224]_  & \new_[36221]_ ;
  assign \new_[36226]_  = \new_[36225]_  & \new_[36218]_ ;
  assign \new_[36230]_  = ~A167 & A168;
  assign \new_[36231]_  = A169 & \new_[36230]_ ;
  assign \new_[36234]_  = ~A199 & A166;
  assign \new_[36237]_  = ~A202 & ~A200;
  assign \new_[36238]_  = \new_[36237]_  & \new_[36234]_ ;
  assign \new_[36239]_  = \new_[36238]_  & \new_[36231]_ ;
  assign \new_[36242]_  = A233 & A232;
  assign \new_[36245]_  = ~A236 & A235;
  assign \new_[36246]_  = \new_[36245]_  & \new_[36242]_ ;
  assign \new_[36249]_  = A299 & A298;
  assign \new_[36252]_  = ~A302 & A301;
  assign \new_[36253]_  = \new_[36252]_  & \new_[36249]_ ;
  assign \new_[36254]_  = \new_[36253]_  & \new_[36246]_ ;
  assign \new_[36258]_  = ~A167 & A168;
  assign \new_[36259]_  = A169 & \new_[36258]_ ;
  assign \new_[36262]_  = ~A199 & A166;
  assign \new_[36265]_  = ~A202 & ~A200;
  assign \new_[36266]_  = \new_[36265]_  & \new_[36262]_ ;
  assign \new_[36267]_  = \new_[36266]_  & \new_[36259]_ ;
  assign \new_[36270]_  = A233 & A232;
  assign \new_[36273]_  = ~A236 & A235;
  assign \new_[36274]_  = \new_[36273]_  & \new_[36270]_ ;
  assign \new_[36277]_  = ~A299 & A298;
  assign \new_[36280]_  = A302 & ~A301;
  assign \new_[36281]_  = \new_[36280]_  & \new_[36277]_ ;
  assign \new_[36282]_  = \new_[36281]_  & \new_[36274]_ ;
  assign \new_[36286]_  = ~A167 & A168;
  assign \new_[36287]_  = A169 & \new_[36286]_ ;
  assign \new_[36290]_  = ~A199 & A166;
  assign \new_[36293]_  = ~A202 & ~A200;
  assign \new_[36294]_  = \new_[36293]_  & \new_[36290]_ ;
  assign \new_[36295]_  = \new_[36294]_  & \new_[36287]_ ;
  assign \new_[36298]_  = A233 & A232;
  assign \new_[36301]_  = ~A236 & A235;
  assign \new_[36302]_  = \new_[36301]_  & \new_[36298]_ ;
  assign \new_[36305]_  = A299 & ~A298;
  assign \new_[36308]_  = A302 & ~A301;
  assign \new_[36309]_  = \new_[36308]_  & \new_[36305]_ ;
  assign \new_[36310]_  = \new_[36309]_  & \new_[36302]_ ;
  assign \new_[36314]_  = ~A167 & A168;
  assign \new_[36315]_  = A169 & \new_[36314]_ ;
  assign \new_[36318]_  = ~A199 & A166;
  assign \new_[36321]_  = ~A202 & ~A200;
  assign \new_[36322]_  = \new_[36321]_  & \new_[36318]_ ;
  assign \new_[36323]_  = \new_[36322]_  & \new_[36315]_ ;
  assign \new_[36326]_  = A233 & A232;
  assign \new_[36329]_  = ~A236 & A235;
  assign \new_[36330]_  = \new_[36329]_  & \new_[36326]_ ;
  assign \new_[36333]_  = ~A299 & ~A298;
  assign \new_[36336]_  = ~A302 & A301;
  assign \new_[36337]_  = \new_[36336]_  & \new_[36333]_ ;
  assign \new_[36338]_  = \new_[36337]_  & \new_[36330]_ ;
  assign \new_[36342]_  = ~A167 & A168;
  assign \new_[36343]_  = A169 & \new_[36342]_ ;
  assign \new_[36346]_  = ~A199 & A166;
  assign \new_[36349]_  = ~A202 & ~A200;
  assign \new_[36350]_  = \new_[36349]_  & \new_[36346]_ ;
  assign \new_[36351]_  = \new_[36350]_  & \new_[36343]_ ;
  assign \new_[36354]_  = A233 & A232;
  assign \new_[36357]_  = ~A236 & A235;
  assign \new_[36358]_  = \new_[36357]_  & \new_[36354]_ ;
  assign \new_[36361]_  = A266 & A265;
  assign \new_[36364]_  = ~A269 & A268;
  assign \new_[36365]_  = \new_[36364]_  & \new_[36361]_ ;
  assign \new_[36366]_  = \new_[36365]_  & \new_[36358]_ ;
  assign \new_[36370]_  = ~A167 & A168;
  assign \new_[36371]_  = A169 & \new_[36370]_ ;
  assign \new_[36374]_  = ~A199 & A166;
  assign \new_[36377]_  = ~A202 & ~A200;
  assign \new_[36378]_  = \new_[36377]_  & \new_[36374]_ ;
  assign \new_[36379]_  = \new_[36378]_  & \new_[36371]_ ;
  assign \new_[36382]_  = A233 & A232;
  assign \new_[36385]_  = ~A236 & A235;
  assign \new_[36386]_  = \new_[36385]_  & \new_[36382]_ ;
  assign \new_[36389]_  = A266 & ~A265;
  assign \new_[36392]_  = A269 & ~A268;
  assign \new_[36393]_  = \new_[36392]_  & \new_[36389]_ ;
  assign \new_[36394]_  = \new_[36393]_  & \new_[36386]_ ;
  assign \new_[36398]_  = ~A167 & A168;
  assign \new_[36399]_  = A169 & \new_[36398]_ ;
  assign \new_[36402]_  = ~A199 & A166;
  assign \new_[36405]_  = ~A202 & ~A200;
  assign \new_[36406]_  = \new_[36405]_  & \new_[36402]_ ;
  assign \new_[36407]_  = \new_[36406]_  & \new_[36399]_ ;
  assign \new_[36410]_  = A233 & A232;
  assign \new_[36413]_  = ~A236 & A235;
  assign \new_[36414]_  = \new_[36413]_  & \new_[36410]_ ;
  assign \new_[36417]_  = ~A266 & A265;
  assign \new_[36420]_  = A269 & ~A268;
  assign \new_[36421]_  = \new_[36420]_  & \new_[36417]_ ;
  assign \new_[36422]_  = \new_[36421]_  & \new_[36414]_ ;
  assign \new_[36426]_  = ~A167 & A168;
  assign \new_[36427]_  = A169 & \new_[36426]_ ;
  assign \new_[36430]_  = ~A199 & A166;
  assign \new_[36433]_  = ~A202 & ~A200;
  assign \new_[36434]_  = \new_[36433]_  & \new_[36430]_ ;
  assign \new_[36435]_  = \new_[36434]_  & \new_[36427]_ ;
  assign \new_[36438]_  = A233 & A232;
  assign \new_[36441]_  = ~A236 & A235;
  assign \new_[36442]_  = \new_[36441]_  & \new_[36438]_ ;
  assign \new_[36445]_  = ~A266 & ~A265;
  assign \new_[36448]_  = ~A269 & A268;
  assign \new_[36449]_  = \new_[36448]_  & \new_[36445]_ ;
  assign \new_[36450]_  = \new_[36449]_  & \new_[36442]_ ;
  assign \new_[36454]_  = ~A167 & A168;
  assign \new_[36455]_  = A169 & \new_[36454]_ ;
  assign \new_[36458]_  = ~A199 & A166;
  assign \new_[36461]_  = ~A202 & ~A200;
  assign \new_[36462]_  = \new_[36461]_  & \new_[36458]_ ;
  assign \new_[36463]_  = \new_[36462]_  & \new_[36455]_ ;
  assign \new_[36466]_  = A233 & ~A232;
  assign \new_[36469]_  = A236 & ~A235;
  assign \new_[36470]_  = \new_[36469]_  & \new_[36466]_ ;
  assign \new_[36473]_  = A299 & A298;
  assign \new_[36476]_  = ~A302 & A301;
  assign \new_[36477]_  = \new_[36476]_  & \new_[36473]_ ;
  assign \new_[36478]_  = \new_[36477]_  & \new_[36470]_ ;
  assign \new_[36482]_  = ~A167 & A168;
  assign \new_[36483]_  = A169 & \new_[36482]_ ;
  assign \new_[36486]_  = ~A199 & A166;
  assign \new_[36489]_  = ~A202 & ~A200;
  assign \new_[36490]_  = \new_[36489]_  & \new_[36486]_ ;
  assign \new_[36491]_  = \new_[36490]_  & \new_[36483]_ ;
  assign \new_[36494]_  = A233 & ~A232;
  assign \new_[36497]_  = A236 & ~A235;
  assign \new_[36498]_  = \new_[36497]_  & \new_[36494]_ ;
  assign \new_[36501]_  = ~A299 & A298;
  assign \new_[36504]_  = A302 & ~A301;
  assign \new_[36505]_  = \new_[36504]_  & \new_[36501]_ ;
  assign \new_[36506]_  = \new_[36505]_  & \new_[36498]_ ;
  assign \new_[36510]_  = ~A167 & A168;
  assign \new_[36511]_  = A169 & \new_[36510]_ ;
  assign \new_[36514]_  = ~A199 & A166;
  assign \new_[36517]_  = ~A202 & ~A200;
  assign \new_[36518]_  = \new_[36517]_  & \new_[36514]_ ;
  assign \new_[36519]_  = \new_[36518]_  & \new_[36511]_ ;
  assign \new_[36522]_  = A233 & ~A232;
  assign \new_[36525]_  = A236 & ~A235;
  assign \new_[36526]_  = \new_[36525]_  & \new_[36522]_ ;
  assign \new_[36529]_  = A299 & ~A298;
  assign \new_[36532]_  = A302 & ~A301;
  assign \new_[36533]_  = \new_[36532]_  & \new_[36529]_ ;
  assign \new_[36534]_  = \new_[36533]_  & \new_[36526]_ ;
  assign \new_[36538]_  = ~A167 & A168;
  assign \new_[36539]_  = A169 & \new_[36538]_ ;
  assign \new_[36542]_  = ~A199 & A166;
  assign \new_[36545]_  = ~A202 & ~A200;
  assign \new_[36546]_  = \new_[36545]_  & \new_[36542]_ ;
  assign \new_[36547]_  = \new_[36546]_  & \new_[36539]_ ;
  assign \new_[36550]_  = A233 & ~A232;
  assign \new_[36553]_  = A236 & ~A235;
  assign \new_[36554]_  = \new_[36553]_  & \new_[36550]_ ;
  assign \new_[36557]_  = ~A299 & ~A298;
  assign \new_[36560]_  = ~A302 & A301;
  assign \new_[36561]_  = \new_[36560]_  & \new_[36557]_ ;
  assign \new_[36562]_  = \new_[36561]_  & \new_[36554]_ ;
  assign \new_[36566]_  = ~A167 & A168;
  assign \new_[36567]_  = A169 & \new_[36566]_ ;
  assign \new_[36570]_  = ~A199 & A166;
  assign \new_[36573]_  = ~A202 & ~A200;
  assign \new_[36574]_  = \new_[36573]_  & \new_[36570]_ ;
  assign \new_[36575]_  = \new_[36574]_  & \new_[36567]_ ;
  assign \new_[36578]_  = A233 & ~A232;
  assign \new_[36581]_  = A236 & ~A235;
  assign \new_[36582]_  = \new_[36581]_  & \new_[36578]_ ;
  assign \new_[36585]_  = A266 & A265;
  assign \new_[36588]_  = ~A269 & A268;
  assign \new_[36589]_  = \new_[36588]_  & \new_[36585]_ ;
  assign \new_[36590]_  = \new_[36589]_  & \new_[36582]_ ;
  assign \new_[36594]_  = ~A167 & A168;
  assign \new_[36595]_  = A169 & \new_[36594]_ ;
  assign \new_[36598]_  = ~A199 & A166;
  assign \new_[36601]_  = ~A202 & ~A200;
  assign \new_[36602]_  = \new_[36601]_  & \new_[36598]_ ;
  assign \new_[36603]_  = \new_[36602]_  & \new_[36595]_ ;
  assign \new_[36606]_  = A233 & ~A232;
  assign \new_[36609]_  = A236 & ~A235;
  assign \new_[36610]_  = \new_[36609]_  & \new_[36606]_ ;
  assign \new_[36613]_  = A266 & ~A265;
  assign \new_[36616]_  = A269 & ~A268;
  assign \new_[36617]_  = \new_[36616]_  & \new_[36613]_ ;
  assign \new_[36618]_  = \new_[36617]_  & \new_[36610]_ ;
  assign \new_[36622]_  = ~A167 & A168;
  assign \new_[36623]_  = A169 & \new_[36622]_ ;
  assign \new_[36626]_  = ~A199 & A166;
  assign \new_[36629]_  = ~A202 & ~A200;
  assign \new_[36630]_  = \new_[36629]_  & \new_[36626]_ ;
  assign \new_[36631]_  = \new_[36630]_  & \new_[36623]_ ;
  assign \new_[36634]_  = A233 & ~A232;
  assign \new_[36637]_  = A236 & ~A235;
  assign \new_[36638]_  = \new_[36637]_  & \new_[36634]_ ;
  assign \new_[36641]_  = ~A266 & A265;
  assign \new_[36644]_  = A269 & ~A268;
  assign \new_[36645]_  = \new_[36644]_  & \new_[36641]_ ;
  assign \new_[36646]_  = \new_[36645]_  & \new_[36638]_ ;
  assign \new_[36650]_  = ~A167 & A168;
  assign \new_[36651]_  = A169 & \new_[36650]_ ;
  assign \new_[36654]_  = ~A199 & A166;
  assign \new_[36657]_  = ~A202 & ~A200;
  assign \new_[36658]_  = \new_[36657]_  & \new_[36654]_ ;
  assign \new_[36659]_  = \new_[36658]_  & \new_[36651]_ ;
  assign \new_[36662]_  = A233 & ~A232;
  assign \new_[36665]_  = A236 & ~A235;
  assign \new_[36666]_  = \new_[36665]_  & \new_[36662]_ ;
  assign \new_[36669]_  = ~A266 & ~A265;
  assign \new_[36672]_  = ~A269 & A268;
  assign \new_[36673]_  = \new_[36672]_  & \new_[36669]_ ;
  assign \new_[36674]_  = \new_[36673]_  & \new_[36666]_ ;
  assign \new_[36678]_  = ~A167 & A168;
  assign \new_[36679]_  = A169 & \new_[36678]_ ;
  assign \new_[36682]_  = ~A199 & A166;
  assign \new_[36685]_  = ~A202 & ~A200;
  assign \new_[36686]_  = \new_[36685]_  & \new_[36682]_ ;
  assign \new_[36687]_  = \new_[36686]_  & \new_[36679]_ ;
  assign \new_[36690]_  = ~A233 & A232;
  assign \new_[36693]_  = A236 & ~A235;
  assign \new_[36694]_  = \new_[36693]_  & \new_[36690]_ ;
  assign \new_[36697]_  = A299 & A298;
  assign \new_[36700]_  = ~A302 & A301;
  assign \new_[36701]_  = \new_[36700]_  & \new_[36697]_ ;
  assign \new_[36702]_  = \new_[36701]_  & \new_[36694]_ ;
  assign \new_[36706]_  = ~A167 & A168;
  assign \new_[36707]_  = A169 & \new_[36706]_ ;
  assign \new_[36710]_  = ~A199 & A166;
  assign \new_[36713]_  = ~A202 & ~A200;
  assign \new_[36714]_  = \new_[36713]_  & \new_[36710]_ ;
  assign \new_[36715]_  = \new_[36714]_  & \new_[36707]_ ;
  assign \new_[36718]_  = ~A233 & A232;
  assign \new_[36721]_  = A236 & ~A235;
  assign \new_[36722]_  = \new_[36721]_  & \new_[36718]_ ;
  assign \new_[36725]_  = ~A299 & A298;
  assign \new_[36728]_  = A302 & ~A301;
  assign \new_[36729]_  = \new_[36728]_  & \new_[36725]_ ;
  assign \new_[36730]_  = \new_[36729]_  & \new_[36722]_ ;
  assign \new_[36734]_  = ~A167 & A168;
  assign \new_[36735]_  = A169 & \new_[36734]_ ;
  assign \new_[36738]_  = ~A199 & A166;
  assign \new_[36741]_  = ~A202 & ~A200;
  assign \new_[36742]_  = \new_[36741]_  & \new_[36738]_ ;
  assign \new_[36743]_  = \new_[36742]_  & \new_[36735]_ ;
  assign \new_[36746]_  = ~A233 & A232;
  assign \new_[36749]_  = A236 & ~A235;
  assign \new_[36750]_  = \new_[36749]_  & \new_[36746]_ ;
  assign \new_[36753]_  = A299 & ~A298;
  assign \new_[36756]_  = A302 & ~A301;
  assign \new_[36757]_  = \new_[36756]_  & \new_[36753]_ ;
  assign \new_[36758]_  = \new_[36757]_  & \new_[36750]_ ;
  assign \new_[36762]_  = ~A167 & A168;
  assign \new_[36763]_  = A169 & \new_[36762]_ ;
  assign \new_[36766]_  = ~A199 & A166;
  assign \new_[36769]_  = ~A202 & ~A200;
  assign \new_[36770]_  = \new_[36769]_  & \new_[36766]_ ;
  assign \new_[36771]_  = \new_[36770]_  & \new_[36763]_ ;
  assign \new_[36774]_  = ~A233 & A232;
  assign \new_[36777]_  = A236 & ~A235;
  assign \new_[36778]_  = \new_[36777]_  & \new_[36774]_ ;
  assign \new_[36781]_  = ~A299 & ~A298;
  assign \new_[36784]_  = ~A302 & A301;
  assign \new_[36785]_  = \new_[36784]_  & \new_[36781]_ ;
  assign \new_[36786]_  = \new_[36785]_  & \new_[36778]_ ;
  assign \new_[36790]_  = ~A167 & A168;
  assign \new_[36791]_  = A169 & \new_[36790]_ ;
  assign \new_[36794]_  = ~A199 & A166;
  assign \new_[36797]_  = ~A202 & ~A200;
  assign \new_[36798]_  = \new_[36797]_  & \new_[36794]_ ;
  assign \new_[36799]_  = \new_[36798]_  & \new_[36791]_ ;
  assign \new_[36802]_  = ~A233 & A232;
  assign \new_[36805]_  = A236 & ~A235;
  assign \new_[36806]_  = \new_[36805]_  & \new_[36802]_ ;
  assign \new_[36809]_  = A266 & A265;
  assign \new_[36812]_  = ~A269 & A268;
  assign \new_[36813]_  = \new_[36812]_  & \new_[36809]_ ;
  assign \new_[36814]_  = \new_[36813]_  & \new_[36806]_ ;
  assign \new_[36818]_  = ~A167 & A168;
  assign \new_[36819]_  = A169 & \new_[36818]_ ;
  assign \new_[36822]_  = ~A199 & A166;
  assign \new_[36825]_  = ~A202 & ~A200;
  assign \new_[36826]_  = \new_[36825]_  & \new_[36822]_ ;
  assign \new_[36827]_  = \new_[36826]_  & \new_[36819]_ ;
  assign \new_[36830]_  = ~A233 & A232;
  assign \new_[36833]_  = A236 & ~A235;
  assign \new_[36834]_  = \new_[36833]_  & \new_[36830]_ ;
  assign \new_[36837]_  = A266 & ~A265;
  assign \new_[36840]_  = A269 & ~A268;
  assign \new_[36841]_  = \new_[36840]_  & \new_[36837]_ ;
  assign \new_[36842]_  = \new_[36841]_  & \new_[36834]_ ;
  assign \new_[36846]_  = ~A167 & A168;
  assign \new_[36847]_  = A169 & \new_[36846]_ ;
  assign \new_[36850]_  = ~A199 & A166;
  assign \new_[36853]_  = ~A202 & ~A200;
  assign \new_[36854]_  = \new_[36853]_  & \new_[36850]_ ;
  assign \new_[36855]_  = \new_[36854]_  & \new_[36847]_ ;
  assign \new_[36858]_  = ~A233 & A232;
  assign \new_[36861]_  = A236 & ~A235;
  assign \new_[36862]_  = \new_[36861]_  & \new_[36858]_ ;
  assign \new_[36865]_  = ~A266 & A265;
  assign \new_[36868]_  = A269 & ~A268;
  assign \new_[36869]_  = \new_[36868]_  & \new_[36865]_ ;
  assign \new_[36870]_  = \new_[36869]_  & \new_[36862]_ ;
  assign \new_[36874]_  = ~A167 & A168;
  assign \new_[36875]_  = A169 & \new_[36874]_ ;
  assign \new_[36878]_  = ~A199 & A166;
  assign \new_[36881]_  = ~A202 & ~A200;
  assign \new_[36882]_  = \new_[36881]_  & \new_[36878]_ ;
  assign \new_[36883]_  = \new_[36882]_  & \new_[36875]_ ;
  assign \new_[36886]_  = ~A233 & A232;
  assign \new_[36889]_  = A236 & ~A235;
  assign \new_[36890]_  = \new_[36889]_  & \new_[36886]_ ;
  assign \new_[36893]_  = ~A266 & ~A265;
  assign \new_[36896]_  = ~A269 & A268;
  assign \new_[36897]_  = \new_[36896]_  & \new_[36893]_ ;
  assign \new_[36898]_  = \new_[36897]_  & \new_[36890]_ ;
  assign \new_[36902]_  = ~A167 & A168;
  assign \new_[36903]_  = A169 & \new_[36902]_ ;
  assign \new_[36906]_  = ~A199 & A166;
  assign \new_[36909]_  = ~A202 & ~A200;
  assign \new_[36910]_  = \new_[36909]_  & \new_[36906]_ ;
  assign \new_[36911]_  = \new_[36910]_  & \new_[36903]_ ;
  assign \new_[36914]_  = ~A233 & ~A232;
  assign \new_[36917]_  = ~A236 & A235;
  assign \new_[36918]_  = \new_[36917]_  & \new_[36914]_ ;
  assign \new_[36921]_  = A299 & A298;
  assign \new_[36924]_  = ~A302 & A301;
  assign \new_[36925]_  = \new_[36924]_  & \new_[36921]_ ;
  assign \new_[36926]_  = \new_[36925]_  & \new_[36918]_ ;
  assign \new_[36930]_  = ~A167 & A168;
  assign \new_[36931]_  = A169 & \new_[36930]_ ;
  assign \new_[36934]_  = ~A199 & A166;
  assign \new_[36937]_  = ~A202 & ~A200;
  assign \new_[36938]_  = \new_[36937]_  & \new_[36934]_ ;
  assign \new_[36939]_  = \new_[36938]_  & \new_[36931]_ ;
  assign \new_[36942]_  = ~A233 & ~A232;
  assign \new_[36945]_  = ~A236 & A235;
  assign \new_[36946]_  = \new_[36945]_  & \new_[36942]_ ;
  assign \new_[36949]_  = ~A299 & A298;
  assign \new_[36952]_  = A302 & ~A301;
  assign \new_[36953]_  = \new_[36952]_  & \new_[36949]_ ;
  assign \new_[36954]_  = \new_[36953]_  & \new_[36946]_ ;
  assign \new_[36958]_  = ~A167 & A168;
  assign \new_[36959]_  = A169 & \new_[36958]_ ;
  assign \new_[36962]_  = ~A199 & A166;
  assign \new_[36965]_  = ~A202 & ~A200;
  assign \new_[36966]_  = \new_[36965]_  & \new_[36962]_ ;
  assign \new_[36967]_  = \new_[36966]_  & \new_[36959]_ ;
  assign \new_[36970]_  = ~A233 & ~A232;
  assign \new_[36973]_  = ~A236 & A235;
  assign \new_[36974]_  = \new_[36973]_  & \new_[36970]_ ;
  assign \new_[36977]_  = A299 & ~A298;
  assign \new_[36980]_  = A302 & ~A301;
  assign \new_[36981]_  = \new_[36980]_  & \new_[36977]_ ;
  assign \new_[36982]_  = \new_[36981]_  & \new_[36974]_ ;
  assign \new_[36986]_  = ~A167 & A168;
  assign \new_[36987]_  = A169 & \new_[36986]_ ;
  assign \new_[36990]_  = ~A199 & A166;
  assign \new_[36993]_  = ~A202 & ~A200;
  assign \new_[36994]_  = \new_[36993]_  & \new_[36990]_ ;
  assign \new_[36995]_  = \new_[36994]_  & \new_[36987]_ ;
  assign \new_[36998]_  = ~A233 & ~A232;
  assign \new_[37001]_  = ~A236 & A235;
  assign \new_[37002]_  = \new_[37001]_  & \new_[36998]_ ;
  assign \new_[37005]_  = ~A299 & ~A298;
  assign \new_[37008]_  = ~A302 & A301;
  assign \new_[37009]_  = \new_[37008]_  & \new_[37005]_ ;
  assign \new_[37010]_  = \new_[37009]_  & \new_[37002]_ ;
  assign \new_[37014]_  = ~A167 & A168;
  assign \new_[37015]_  = A169 & \new_[37014]_ ;
  assign \new_[37018]_  = ~A199 & A166;
  assign \new_[37021]_  = ~A202 & ~A200;
  assign \new_[37022]_  = \new_[37021]_  & \new_[37018]_ ;
  assign \new_[37023]_  = \new_[37022]_  & \new_[37015]_ ;
  assign \new_[37026]_  = ~A233 & ~A232;
  assign \new_[37029]_  = ~A236 & A235;
  assign \new_[37030]_  = \new_[37029]_  & \new_[37026]_ ;
  assign \new_[37033]_  = A266 & A265;
  assign \new_[37036]_  = ~A269 & A268;
  assign \new_[37037]_  = \new_[37036]_  & \new_[37033]_ ;
  assign \new_[37038]_  = \new_[37037]_  & \new_[37030]_ ;
  assign \new_[37042]_  = ~A167 & A168;
  assign \new_[37043]_  = A169 & \new_[37042]_ ;
  assign \new_[37046]_  = ~A199 & A166;
  assign \new_[37049]_  = ~A202 & ~A200;
  assign \new_[37050]_  = \new_[37049]_  & \new_[37046]_ ;
  assign \new_[37051]_  = \new_[37050]_  & \new_[37043]_ ;
  assign \new_[37054]_  = ~A233 & ~A232;
  assign \new_[37057]_  = ~A236 & A235;
  assign \new_[37058]_  = \new_[37057]_  & \new_[37054]_ ;
  assign \new_[37061]_  = A266 & ~A265;
  assign \new_[37064]_  = A269 & ~A268;
  assign \new_[37065]_  = \new_[37064]_  & \new_[37061]_ ;
  assign \new_[37066]_  = \new_[37065]_  & \new_[37058]_ ;
  assign \new_[37070]_  = ~A167 & A168;
  assign \new_[37071]_  = A169 & \new_[37070]_ ;
  assign \new_[37074]_  = ~A199 & A166;
  assign \new_[37077]_  = ~A202 & ~A200;
  assign \new_[37078]_  = \new_[37077]_  & \new_[37074]_ ;
  assign \new_[37079]_  = \new_[37078]_  & \new_[37071]_ ;
  assign \new_[37082]_  = ~A233 & ~A232;
  assign \new_[37085]_  = ~A236 & A235;
  assign \new_[37086]_  = \new_[37085]_  & \new_[37082]_ ;
  assign \new_[37089]_  = ~A266 & A265;
  assign \new_[37092]_  = A269 & ~A268;
  assign \new_[37093]_  = \new_[37092]_  & \new_[37089]_ ;
  assign \new_[37094]_  = \new_[37093]_  & \new_[37086]_ ;
  assign \new_[37098]_  = ~A167 & A168;
  assign \new_[37099]_  = A169 & \new_[37098]_ ;
  assign \new_[37102]_  = ~A199 & A166;
  assign \new_[37105]_  = ~A202 & ~A200;
  assign \new_[37106]_  = \new_[37105]_  & \new_[37102]_ ;
  assign \new_[37107]_  = \new_[37106]_  & \new_[37099]_ ;
  assign \new_[37110]_  = ~A233 & ~A232;
  assign \new_[37113]_  = ~A236 & A235;
  assign \new_[37114]_  = \new_[37113]_  & \new_[37110]_ ;
  assign \new_[37117]_  = ~A266 & ~A265;
  assign \new_[37120]_  = ~A269 & A268;
  assign \new_[37121]_  = \new_[37120]_  & \new_[37117]_ ;
  assign \new_[37122]_  = \new_[37121]_  & \new_[37114]_ ;
  assign \new_[37126]_  = ~A167 & A168;
  assign \new_[37127]_  = A169 & \new_[37126]_ ;
  assign \new_[37130]_  = ~A199 & A166;
  assign \new_[37133]_  = A203 & ~A200;
  assign \new_[37134]_  = \new_[37133]_  & \new_[37130]_ ;
  assign \new_[37135]_  = \new_[37134]_  & \new_[37127]_ ;
  assign \new_[37138]_  = A233 & A232;
  assign \new_[37141]_  = ~A236 & A235;
  assign \new_[37142]_  = \new_[37141]_  & \new_[37138]_ ;
  assign \new_[37145]_  = A299 & A298;
  assign \new_[37148]_  = ~A302 & A301;
  assign \new_[37149]_  = \new_[37148]_  & \new_[37145]_ ;
  assign \new_[37150]_  = \new_[37149]_  & \new_[37142]_ ;
  assign \new_[37154]_  = ~A167 & A168;
  assign \new_[37155]_  = A169 & \new_[37154]_ ;
  assign \new_[37158]_  = ~A199 & A166;
  assign \new_[37161]_  = A203 & ~A200;
  assign \new_[37162]_  = \new_[37161]_  & \new_[37158]_ ;
  assign \new_[37163]_  = \new_[37162]_  & \new_[37155]_ ;
  assign \new_[37166]_  = A233 & A232;
  assign \new_[37169]_  = ~A236 & A235;
  assign \new_[37170]_  = \new_[37169]_  & \new_[37166]_ ;
  assign \new_[37173]_  = ~A299 & A298;
  assign \new_[37176]_  = A302 & ~A301;
  assign \new_[37177]_  = \new_[37176]_  & \new_[37173]_ ;
  assign \new_[37178]_  = \new_[37177]_  & \new_[37170]_ ;
  assign \new_[37182]_  = ~A167 & A168;
  assign \new_[37183]_  = A169 & \new_[37182]_ ;
  assign \new_[37186]_  = ~A199 & A166;
  assign \new_[37189]_  = A203 & ~A200;
  assign \new_[37190]_  = \new_[37189]_  & \new_[37186]_ ;
  assign \new_[37191]_  = \new_[37190]_  & \new_[37183]_ ;
  assign \new_[37194]_  = A233 & A232;
  assign \new_[37197]_  = ~A236 & A235;
  assign \new_[37198]_  = \new_[37197]_  & \new_[37194]_ ;
  assign \new_[37201]_  = A299 & ~A298;
  assign \new_[37204]_  = A302 & ~A301;
  assign \new_[37205]_  = \new_[37204]_  & \new_[37201]_ ;
  assign \new_[37206]_  = \new_[37205]_  & \new_[37198]_ ;
  assign \new_[37210]_  = ~A167 & A168;
  assign \new_[37211]_  = A169 & \new_[37210]_ ;
  assign \new_[37214]_  = ~A199 & A166;
  assign \new_[37217]_  = A203 & ~A200;
  assign \new_[37218]_  = \new_[37217]_  & \new_[37214]_ ;
  assign \new_[37219]_  = \new_[37218]_  & \new_[37211]_ ;
  assign \new_[37222]_  = A233 & A232;
  assign \new_[37225]_  = ~A236 & A235;
  assign \new_[37226]_  = \new_[37225]_  & \new_[37222]_ ;
  assign \new_[37229]_  = ~A299 & ~A298;
  assign \new_[37232]_  = ~A302 & A301;
  assign \new_[37233]_  = \new_[37232]_  & \new_[37229]_ ;
  assign \new_[37234]_  = \new_[37233]_  & \new_[37226]_ ;
  assign \new_[37238]_  = ~A167 & A168;
  assign \new_[37239]_  = A169 & \new_[37238]_ ;
  assign \new_[37242]_  = ~A199 & A166;
  assign \new_[37245]_  = A203 & ~A200;
  assign \new_[37246]_  = \new_[37245]_  & \new_[37242]_ ;
  assign \new_[37247]_  = \new_[37246]_  & \new_[37239]_ ;
  assign \new_[37250]_  = A233 & A232;
  assign \new_[37253]_  = ~A236 & A235;
  assign \new_[37254]_  = \new_[37253]_  & \new_[37250]_ ;
  assign \new_[37257]_  = A266 & A265;
  assign \new_[37260]_  = ~A269 & A268;
  assign \new_[37261]_  = \new_[37260]_  & \new_[37257]_ ;
  assign \new_[37262]_  = \new_[37261]_  & \new_[37254]_ ;
  assign \new_[37266]_  = ~A167 & A168;
  assign \new_[37267]_  = A169 & \new_[37266]_ ;
  assign \new_[37270]_  = ~A199 & A166;
  assign \new_[37273]_  = A203 & ~A200;
  assign \new_[37274]_  = \new_[37273]_  & \new_[37270]_ ;
  assign \new_[37275]_  = \new_[37274]_  & \new_[37267]_ ;
  assign \new_[37278]_  = A233 & A232;
  assign \new_[37281]_  = ~A236 & A235;
  assign \new_[37282]_  = \new_[37281]_  & \new_[37278]_ ;
  assign \new_[37285]_  = A266 & ~A265;
  assign \new_[37288]_  = A269 & ~A268;
  assign \new_[37289]_  = \new_[37288]_  & \new_[37285]_ ;
  assign \new_[37290]_  = \new_[37289]_  & \new_[37282]_ ;
  assign \new_[37294]_  = ~A167 & A168;
  assign \new_[37295]_  = A169 & \new_[37294]_ ;
  assign \new_[37298]_  = ~A199 & A166;
  assign \new_[37301]_  = A203 & ~A200;
  assign \new_[37302]_  = \new_[37301]_  & \new_[37298]_ ;
  assign \new_[37303]_  = \new_[37302]_  & \new_[37295]_ ;
  assign \new_[37306]_  = A233 & A232;
  assign \new_[37309]_  = ~A236 & A235;
  assign \new_[37310]_  = \new_[37309]_  & \new_[37306]_ ;
  assign \new_[37313]_  = ~A266 & A265;
  assign \new_[37316]_  = A269 & ~A268;
  assign \new_[37317]_  = \new_[37316]_  & \new_[37313]_ ;
  assign \new_[37318]_  = \new_[37317]_  & \new_[37310]_ ;
  assign \new_[37322]_  = ~A167 & A168;
  assign \new_[37323]_  = A169 & \new_[37322]_ ;
  assign \new_[37326]_  = ~A199 & A166;
  assign \new_[37329]_  = A203 & ~A200;
  assign \new_[37330]_  = \new_[37329]_  & \new_[37326]_ ;
  assign \new_[37331]_  = \new_[37330]_  & \new_[37323]_ ;
  assign \new_[37334]_  = A233 & A232;
  assign \new_[37337]_  = ~A236 & A235;
  assign \new_[37338]_  = \new_[37337]_  & \new_[37334]_ ;
  assign \new_[37341]_  = ~A266 & ~A265;
  assign \new_[37344]_  = ~A269 & A268;
  assign \new_[37345]_  = \new_[37344]_  & \new_[37341]_ ;
  assign \new_[37346]_  = \new_[37345]_  & \new_[37338]_ ;
  assign \new_[37350]_  = ~A167 & A168;
  assign \new_[37351]_  = A169 & \new_[37350]_ ;
  assign \new_[37354]_  = ~A199 & A166;
  assign \new_[37357]_  = A203 & ~A200;
  assign \new_[37358]_  = \new_[37357]_  & \new_[37354]_ ;
  assign \new_[37359]_  = \new_[37358]_  & \new_[37351]_ ;
  assign \new_[37362]_  = A233 & ~A232;
  assign \new_[37365]_  = A236 & ~A235;
  assign \new_[37366]_  = \new_[37365]_  & \new_[37362]_ ;
  assign \new_[37369]_  = A299 & A298;
  assign \new_[37372]_  = ~A302 & A301;
  assign \new_[37373]_  = \new_[37372]_  & \new_[37369]_ ;
  assign \new_[37374]_  = \new_[37373]_  & \new_[37366]_ ;
  assign \new_[37378]_  = ~A167 & A168;
  assign \new_[37379]_  = A169 & \new_[37378]_ ;
  assign \new_[37382]_  = ~A199 & A166;
  assign \new_[37385]_  = A203 & ~A200;
  assign \new_[37386]_  = \new_[37385]_  & \new_[37382]_ ;
  assign \new_[37387]_  = \new_[37386]_  & \new_[37379]_ ;
  assign \new_[37390]_  = A233 & ~A232;
  assign \new_[37393]_  = A236 & ~A235;
  assign \new_[37394]_  = \new_[37393]_  & \new_[37390]_ ;
  assign \new_[37397]_  = ~A299 & A298;
  assign \new_[37400]_  = A302 & ~A301;
  assign \new_[37401]_  = \new_[37400]_  & \new_[37397]_ ;
  assign \new_[37402]_  = \new_[37401]_  & \new_[37394]_ ;
  assign \new_[37406]_  = ~A167 & A168;
  assign \new_[37407]_  = A169 & \new_[37406]_ ;
  assign \new_[37410]_  = ~A199 & A166;
  assign \new_[37413]_  = A203 & ~A200;
  assign \new_[37414]_  = \new_[37413]_  & \new_[37410]_ ;
  assign \new_[37415]_  = \new_[37414]_  & \new_[37407]_ ;
  assign \new_[37418]_  = A233 & ~A232;
  assign \new_[37421]_  = A236 & ~A235;
  assign \new_[37422]_  = \new_[37421]_  & \new_[37418]_ ;
  assign \new_[37425]_  = A299 & ~A298;
  assign \new_[37428]_  = A302 & ~A301;
  assign \new_[37429]_  = \new_[37428]_  & \new_[37425]_ ;
  assign \new_[37430]_  = \new_[37429]_  & \new_[37422]_ ;
  assign \new_[37434]_  = ~A167 & A168;
  assign \new_[37435]_  = A169 & \new_[37434]_ ;
  assign \new_[37438]_  = ~A199 & A166;
  assign \new_[37441]_  = A203 & ~A200;
  assign \new_[37442]_  = \new_[37441]_  & \new_[37438]_ ;
  assign \new_[37443]_  = \new_[37442]_  & \new_[37435]_ ;
  assign \new_[37446]_  = A233 & ~A232;
  assign \new_[37449]_  = A236 & ~A235;
  assign \new_[37450]_  = \new_[37449]_  & \new_[37446]_ ;
  assign \new_[37453]_  = ~A299 & ~A298;
  assign \new_[37456]_  = ~A302 & A301;
  assign \new_[37457]_  = \new_[37456]_  & \new_[37453]_ ;
  assign \new_[37458]_  = \new_[37457]_  & \new_[37450]_ ;
  assign \new_[37462]_  = ~A167 & A168;
  assign \new_[37463]_  = A169 & \new_[37462]_ ;
  assign \new_[37466]_  = ~A199 & A166;
  assign \new_[37469]_  = A203 & ~A200;
  assign \new_[37470]_  = \new_[37469]_  & \new_[37466]_ ;
  assign \new_[37471]_  = \new_[37470]_  & \new_[37463]_ ;
  assign \new_[37474]_  = A233 & ~A232;
  assign \new_[37477]_  = A236 & ~A235;
  assign \new_[37478]_  = \new_[37477]_  & \new_[37474]_ ;
  assign \new_[37481]_  = A266 & A265;
  assign \new_[37484]_  = ~A269 & A268;
  assign \new_[37485]_  = \new_[37484]_  & \new_[37481]_ ;
  assign \new_[37486]_  = \new_[37485]_  & \new_[37478]_ ;
  assign \new_[37490]_  = ~A167 & A168;
  assign \new_[37491]_  = A169 & \new_[37490]_ ;
  assign \new_[37494]_  = ~A199 & A166;
  assign \new_[37497]_  = A203 & ~A200;
  assign \new_[37498]_  = \new_[37497]_  & \new_[37494]_ ;
  assign \new_[37499]_  = \new_[37498]_  & \new_[37491]_ ;
  assign \new_[37502]_  = A233 & ~A232;
  assign \new_[37505]_  = A236 & ~A235;
  assign \new_[37506]_  = \new_[37505]_  & \new_[37502]_ ;
  assign \new_[37509]_  = A266 & ~A265;
  assign \new_[37512]_  = A269 & ~A268;
  assign \new_[37513]_  = \new_[37512]_  & \new_[37509]_ ;
  assign \new_[37514]_  = \new_[37513]_  & \new_[37506]_ ;
  assign \new_[37518]_  = ~A167 & A168;
  assign \new_[37519]_  = A169 & \new_[37518]_ ;
  assign \new_[37522]_  = ~A199 & A166;
  assign \new_[37525]_  = A203 & ~A200;
  assign \new_[37526]_  = \new_[37525]_  & \new_[37522]_ ;
  assign \new_[37527]_  = \new_[37526]_  & \new_[37519]_ ;
  assign \new_[37530]_  = A233 & ~A232;
  assign \new_[37533]_  = A236 & ~A235;
  assign \new_[37534]_  = \new_[37533]_  & \new_[37530]_ ;
  assign \new_[37537]_  = ~A266 & A265;
  assign \new_[37540]_  = A269 & ~A268;
  assign \new_[37541]_  = \new_[37540]_  & \new_[37537]_ ;
  assign \new_[37542]_  = \new_[37541]_  & \new_[37534]_ ;
  assign \new_[37546]_  = ~A167 & A168;
  assign \new_[37547]_  = A169 & \new_[37546]_ ;
  assign \new_[37550]_  = ~A199 & A166;
  assign \new_[37553]_  = A203 & ~A200;
  assign \new_[37554]_  = \new_[37553]_  & \new_[37550]_ ;
  assign \new_[37555]_  = \new_[37554]_  & \new_[37547]_ ;
  assign \new_[37558]_  = A233 & ~A232;
  assign \new_[37561]_  = A236 & ~A235;
  assign \new_[37562]_  = \new_[37561]_  & \new_[37558]_ ;
  assign \new_[37565]_  = ~A266 & ~A265;
  assign \new_[37568]_  = ~A269 & A268;
  assign \new_[37569]_  = \new_[37568]_  & \new_[37565]_ ;
  assign \new_[37570]_  = \new_[37569]_  & \new_[37562]_ ;
  assign \new_[37574]_  = ~A167 & A168;
  assign \new_[37575]_  = A169 & \new_[37574]_ ;
  assign \new_[37578]_  = ~A199 & A166;
  assign \new_[37581]_  = A203 & ~A200;
  assign \new_[37582]_  = \new_[37581]_  & \new_[37578]_ ;
  assign \new_[37583]_  = \new_[37582]_  & \new_[37575]_ ;
  assign \new_[37586]_  = ~A233 & A232;
  assign \new_[37589]_  = A236 & ~A235;
  assign \new_[37590]_  = \new_[37589]_  & \new_[37586]_ ;
  assign \new_[37593]_  = A299 & A298;
  assign \new_[37596]_  = ~A302 & A301;
  assign \new_[37597]_  = \new_[37596]_  & \new_[37593]_ ;
  assign \new_[37598]_  = \new_[37597]_  & \new_[37590]_ ;
  assign \new_[37602]_  = ~A167 & A168;
  assign \new_[37603]_  = A169 & \new_[37602]_ ;
  assign \new_[37606]_  = ~A199 & A166;
  assign \new_[37609]_  = A203 & ~A200;
  assign \new_[37610]_  = \new_[37609]_  & \new_[37606]_ ;
  assign \new_[37611]_  = \new_[37610]_  & \new_[37603]_ ;
  assign \new_[37614]_  = ~A233 & A232;
  assign \new_[37617]_  = A236 & ~A235;
  assign \new_[37618]_  = \new_[37617]_  & \new_[37614]_ ;
  assign \new_[37621]_  = ~A299 & A298;
  assign \new_[37624]_  = A302 & ~A301;
  assign \new_[37625]_  = \new_[37624]_  & \new_[37621]_ ;
  assign \new_[37626]_  = \new_[37625]_  & \new_[37618]_ ;
  assign \new_[37630]_  = ~A167 & A168;
  assign \new_[37631]_  = A169 & \new_[37630]_ ;
  assign \new_[37634]_  = ~A199 & A166;
  assign \new_[37637]_  = A203 & ~A200;
  assign \new_[37638]_  = \new_[37637]_  & \new_[37634]_ ;
  assign \new_[37639]_  = \new_[37638]_  & \new_[37631]_ ;
  assign \new_[37642]_  = ~A233 & A232;
  assign \new_[37645]_  = A236 & ~A235;
  assign \new_[37646]_  = \new_[37645]_  & \new_[37642]_ ;
  assign \new_[37649]_  = A299 & ~A298;
  assign \new_[37652]_  = A302 & ~A301;
  assign \new_[37653]_  = \new_[37652]_  & \new_[37649]_ ;
  assign \new_[37654]_  = \new_[37653]_  & \new_[37646]_ ;
  assign \new_[37658]_  = ~A167 & A168;
  assign \new_[37659]_  = A169 & \new_[37658]_ ;
  assign \new_[37662]_  = ~A199 & A166;
  assign \new_[37665]_  = A203 & ~A200;
  assign \new_[37666]_  = \new_[37665]_  & \new_[37662]_ ;
  assign \new_[37667]_  = \new_[37666]_  & \new_[37659]_ ;
  assign \new_[37670]_  = ~A233 & A232;
  assign \new_[37673]_  = A236 & ~A235;
  assign \new_[37674]_  = \new_[37673]_  & \new_[37670]_ ;
  assign \new_[37677]_  = ~A299 & ~A298;
  assign \new_[37680]_  = ~A302 & A301;
  assign \new_[37681]_  = \new_[37680]_  & \new_[37677]_ ;
  assign \new_[37682]_  = \new_[37681]_  & \new_[37674]_ ;
  assign \new_[37686]_  = ~A167 & A168;
  assign \new_[37687]_  = A169 & \new_[37686]_ ;
  assign \new_[37690]_  = ~A199 & A166;
  assign \new_[37693]_  = A203 & ~A200;
  assign \new_[37694]_  = \new_[37693]_  & \new_[37690]_ ;
  assign \new_[37695]_  = \new_[37694]_  & \new_[37687]_ ;
  assign \new_[37698]_  = ~A233 & A232;
  assign \new_[37701]_  = A236 & ~A235;
  assign \new_[37702]_  = \new_[37701]_  & \new_[37698]_ ;
  assign \new_[37705]_  = A266 & A265;
  assign \new_[37708]_  = ~A269 & A268;
  assign \new_[37709]_  = \new_[37708]_  & \new_[37705]_ ;
  assign \new_[37710]_  = \new_[37709]_  & \new_[37702]_ ;
  assign \new_[37714]_  = ~A167 & A168;
  assign \new_[37715]_  = A169 & \new_[37714]_ ;
  assign \new_[37718]_  = ~A199 & A166;
  assign \new_[37721]_  = A203 & ~A200;
  assign \new_[37722]_  = \new_[37721]_  & \new_[37718]_ ;
  assign \new_[37723]_  = \new_[37722]_  & \new_[37715]_ ;
  assign \new_[37726]_  = ~A233 & A232;
  assign \new_[37729]_  = A236 & ~A235;
  assign \new_[37730]_  = \new_[37729]_  & \new_[37726]_ ;
  assign \new_[37733]_  = A266 & ~A265;
  assign \new_[37736]_  = A269 & ~A268;
  assign \new_[37737]_  = \new_[37736]_  & \new_[37733]_ ;
  assign \new_[37738]_  = \new_[37737]_  & \new_[37730]_ ;
  assign \new_[37742]_  = ~A167 & A168;
  assign \new_[37743]_  = A169 & \new_[37742]_ ;
  assign \new_[37746]_  = ~A199 & A166;
  assign \new_[37749]_  = A203 & ~A200;
  assign \new_[37750]_  = \new_[37749]_  & \new_[37746]_ ;
  assign \new_[37751]_  = \new_[37750]_  & \new_[37743]_ ;
  assign \new_[37754]_  = ~A233 & A232;
  assign \new_[37757]_  = A236 & ~A235;
  assign \new_[37758]_  = \new_[37757]_  & \new_[37754]_ ;
  assign \new_[37761]_  = ~A266 & A265;
  assign \new_[37764]_  = A269 & ~A268;
  assign \new_[37765]_  = \new_[37764]_  & \new_[37761]_ ;
  assign \new_[37766]_  = \new_[37765]_  & \new_[37758]_ ;
  assign \new_[37770]_  = ~A167 & A168;
  assign \new_[37771]_  = A169 & \new_[37770]_ ;
  assign \new_[37774]_  = ~A199 & A166;
  assign \new_[37777]_  = A203 & ~A200;
  assign \new_[37778]_  = \new_[37777]_  & \new_[37774]_ ;
  assign \new_[37779]_  = \new_[37778]_  & \new_[37771]_ ;
  assign \new_[37782]_  = ~A233 & A232;
  assign \new_[37785]_  = A236 & ~A235;
  assign \new_[37786]_  = \new_[37785]_  & \new_[37782]_ ;
  assign \new_[37789]_  = ~A266 & ~A265;
  assign \new_[37792]_  = ~A269 & A268;
  assign \new_[37793]_  = \new_[37792]_  & \new_[37789]_ ;
  assign \new_[37794]_  = \new_[37793]_  & \new_[37786]_ ;
  assign \new_[37798]_  = ~A167 & A168;
  assign \new_[37799]_  = A169 & \new_[37798]_ ;
  assign \new_[37802]_  = ~A199 & A166;
  assign \new_[37805]_  = A203 & ~A200;
  assign \new_[37806]_  = \new_[37805]_  & \new_[37802]_ ;
  assign \new_[37807]_  = \new_[37806]_  & \new_[37799]_ ;
  assign \new_[37810]_  = ~A233 & ~A232;
  assign \new_[37813]_  = ~A236 & A235;
  assign \new_[37814]_  = \new_[37813]_  & \new_[37810]_ ;
  assign \new_[37817]_  = A299 & A298;
  assign \new_[37820]_  = ~A302 & A301;
  assign \new_[37821]_  = \new_[37820]_  & \new_[37817]_ ;
  assign \new_[37822]_  = \new_[37821]_  & \new_[37814]_ ;
  assign \new_[37826]_  = ~A167 & A168;
  assign \new_[37827]_  = A169 & \new_[37826]_ ;
  assign \new_[37830]_  = ~A199 & A166;
  assign \new_[37833]_  = A203 & ~A200;
  assign \new_[37834]_  = \new_[37833]_  & \new_[37830]_ ;
  assign \new_[37835]_  = \new_[37834]_  & \new_[37827]_ ;
  assign \new_[37838]_  = ~A233 & ~A232;
  assign \new_[37841]_  = ~A236 & A235;
  assign \new_[37842]_  = \new_[37841]_  & \new_[37838]_ ;
  assign \new_[37845]_  = ~A299 & A298;
  assign \new_[37848]_  = A302 & ~A301;
  assign \new_[37849]_  = \new_[37848]_  & \new_[37845]_ ;
  assign \new_[37850]_  = \new_[37849]_  & \new_[37842]_ ;
  assign \new_[37854]_  = ~A167 & A168;
  assign \new_[37855]_  = A169 & \new_[37854]_ ;
  assign \new_[37858]_  = ~A199 & A166;
  assign \new_[37861]_  = A203 & ~A200;
  assign \new_[37862]_  = \new_[37861]_  & \new_[37858]_ ;
  assign \new_[37863]_  = \new_[37862]_  & \new_[37855]_ ;
  assign \new_[37866]_  = ~A233 & ~A232;
  assign \new_[37869]_  = ~A236 & A235;
  assign \new_[37870]_  = \new_[37869]_  & \new_[37866]_ ;
  assign \new_[37873]_  = A299 & ~A298;
  assign \new_[37876]_  = A302 & ~A301;
  assign \new_[37877]_  = \new_[37876]_  & \new_[37873]_ ;
  assign \new_[37878]_  = \new_[37877]_  & \new_[37870]_ ;
  assign \new_[37882]_  = ~A167 & A168;
  assign \new_[37883]_  = A169 & \new_[37882]_ ;
  assign \new_[37886]_  = ~A199 & A166;
  assign \new_[37889]_  = A203 & ~A200;
  assign \new_[37890]_  = \new_[37889]_  & \new_[37886]_ ;
  assign \new_[37891]_  = \new_[37890]_  & \new_[37883]_ ;
  assign \new_[37894]_  = ~A233 & ~A232;
  assign \new_[37897]_  = ~A236 & A235;
  assign \new_[37898]_  = \new_[37897]_  & \new_[37894]_ ;
  assign \new_[37901]_  = ~A299 & ~A298;
  assign \new_[37904]_  = ~A302 & A301;
  assign \new_[37905]_  = \new_[37904]_  & \new_[37901]_ ;
  assign \new_[37906]_  = \new_[37905]_  & \new_[37898]_ ;
  assign \new_[37910]_  = ~A167 & A168;
  assign \new_[37911]_  = A169 & \new_[37910]_ ;
  assign \new_[37914]_  = ~A199 & A166;
  assign \new_[37917]_  = A203 & ~A200;
  assign \new_[37918]_  = \new_[37917]_  & \new_[37914]_ ;
  assign \new_[37919]_  = \new_[37918]_  & \new_[37911]_ ;
  assign \new_[37922]_  = ~A233 & ~A232;
  assign \new_[37925]_  = ~A236 & A235;
  assign \new_[37926]_  = \new_[37925]_  & \new_[37922]_ ;
  assign \new_[37929]_  = A266 & A265;
  assign \new_[37932]_  = ~A269 & A268;
  assign \new_[37933]_  = \new_[37932]_  & \new_[37929]_ ;
  assign \new_[37934]_  = \new_[37933]_  & \new_[37926]_ ;
  assign \new_[37938]_  = ~A167 & A168;
  assign \new_[37939]_  = A169 & \new_[37938]_ ;
  assign \new_[37942]_  = ~A199 & A166;
  assign \new_[37945]_  = A203 & ~A200;
  assign \new_[37946]_  = \new_[37945]_  & \new_[37942]_ ;
  assign \new_[37947]_  = \new_[37946]_  & \new_[37939]_ ;
  assign \new_[37950]_  = ~A233 & ~A232;
  assign \new_[37953]_  = ~A236 & A235;
  assign \new_[37954]_  = \new_[37953]_  & \new_[37950]_ ;
  assign \new_[37957]_  = A266 & ~A265;
  assign \new_[37960]_  = A269 & ~A268;
  assign \new_[37961]_  = \new_[37960]_  & \new_[37957]_ ;
  assign \new_[37962]_  = \new_[37961]_  & \new_[37954]_ ;
  assign \new_[37966]_  = ~A167 & A168;
  assign \new_[37967]_  = A169 & \new_[37966]_ ;
  assign \new_[37970]_  = ~A199 & A166;
  assign \new_[37973]_  = A203 & ~A200;
  assign \new_[37974]_  = \new_[37973]_  & \new_[37970]_ ;
  assign \new_[37975]_  = \new_[37974]_  & \new_[37967]_ ;
  assign \new_[37978]_  = ~A233 & ~A232;
  assign \new_[37981]_  = ~A236 & A235;
  assign \new_[37982]_  = \new_[37981]_  & \new_[37978]_ ;
  assign \new_[37985]_  = ~A266 & A265;
  assign \new_[37988]_  = A269 & ~A268;
  assign \new_[37989]_  = \new_[37988]_  & \new_[37985]_ ;
  assign \new_[37990]_  = \new_[37989]_  & \new_[37982]_ ;
  assign \new_[37994]_  = ~A167 & A168;
  assign \new_[37995]_  = A169 & \new_[37994]_ ;
  assign \new_[37998]_  = ~A199 & A166;
  assign \new_[38001]_  = A203 & ~A200;
  assign \new_[38002]_  = \new_[38001]_  & \new_[37998]_ ;
  assign \new_[38003]_  = \new_[38002]_  & \new_[37995]_ ;
  assign \new_[38006]_  = ~A233 & ~A232;
  assign \new_[38009]_  = ~A236 & A235;
  assign \new_[38010]_  = \new_[38009]_  & \new_[38006]_ ;
  assign \new_[38013]_  = ~A266 & ~A265;
  assign \new_[38016]_  = ~A269 & A268;
  assign \new_[38017]_  = \new_[38016]_  & \new_[38013]_ ;
  assign \new_[38018]_  = \new_[38017]_  & \new_[38010]_ ;
  assign \new_[38021]_  = A168 & A170;
  assign \new_[38024]_  = A166 & ~A167;
  assign \new_[38025]_  = \new_[38024]_  & \new_[38021]_ ;
  assign \new_[38028]_  = A200 & A199;
  assign \new_[38031]_  = ~A202 & ~A201;
  assign \new_[38032]_  = \new_[38031]_  & \new_[38028]_ ;
  assign \new_[38033]_  = \new_[38032]_  & \new_[38025]_ ;
  assign \new_[38036]_  = A233 & A232;
  assign \new_[38039]_  = ~A236 & A235;
  assign \new_[38040]_  = \new_[38039]_  & \new_[38036]_ ;
  assign \new_[38043]_  = A299 & A298;
  assign \new_[38046]_  = ~A302 & A301;
  assign \new_[38047]_  = \new_[38046]_  & \new_[38043]_ ;
  assign \new_[38048]_  = \new_[38047]_  & \new_[38040]_ ;
  assign \new_[38051]_  = A168 & A170;
  assign \new_[38054]_  = A166 & ~A167;
  assign \new_[38055]_  = \new_[38054]_  & \new_[38051]_ ;
  assign \new_[38058]_  = A200 & A199;
  assign \new_[38061]_  = ~A202 & ~A201;
  assign \new_[38062]_  = \new_[38061]_  & \new_[38058]_ ;
  assign \new_[38063]_  = \new_[38062]_  & \new_[38055]_ ;
  assign \new_[38066]_  = A233 & A232;
  assign \new_[38069]_  = ~A236 & A235;
  assign \new_[38070]_  = \new_[38069]_  & \new_[38066]_ ;
  assign \new_[38073]_  = ~A299 & A298;
  assign \new_[38076]_  = A302 & ~A301;
  assign \new_[38077]_  = \new_[38076]_  & \new_[38073]_ ;
  assign \new_[38078]_  = \new_[38077]_  & \new_[38070]_ ;
  assign \new_[38081]_  = A168 & A170;
  assign \new_[38084]_  = A166 & ~A167;
  assign \new_[38085]_  = \new_[38084]_  & \new_[38081]_ ;
  assign \new_[38088]_  = A200 & A199;
  assign \new_[38091]_  = ~A202 & ~A201;
  assign \new_[38092]_  = \new_[38091]_  & \new_[38088]_ ;
  assign \new_[38093]_  = \new_[38092]_  & \new_[38085]_ ;
  assign \new_[38096]_  = A233 & A232;
  assign \new_[38099]_  = ~A236 & A235;
  assign \new_[38100]_  = \new_[38099]_  & \new_[38096]_ ;
  assign \new_[38103]_  = A299 & ~A298;
  assign \new_[38106]_  = A302 & ~A301;
  assign \new_[38107]_  = \new_[38106]_  & \new_[38103]_ ;
  assign \new_[38108]_  = \new_[38107]_  & \new_[38100]_ ;
  assign \new_[38111]_  = A168 & A170;
  assign \new_[38114]_  = A166 & ~A167;
  assign \new_[38115]_  = \new_[38114]_  & \new_[38111]_ ;
  assign \new_[38118]_  = A200 & A199;
  assign \new_[38121]_  = ~A202 & ~A201;
  assign \new_[38122]_  = \new_[38121]_  & \new_[38118]_ ;
  assign \new_[38123]_  = \new_[38122]_  & \new_[38115]_ ;
  assign \new_[38126]_  = A233 & A232;
  assign \new_[38129]_  = ~A236 & A235;
  assign \new_[38130]_  = \new_[38129]_  & \new_[38126]_ ;
  assign \new_[38133]_  = ~A299 & ~A298;
  assign \new_[38136]_  = ~A302 & A301;
  assign \new_[38137]_  = \new_[38136]_  & \new_[38133]_ ;
  assign \new_[38138]_  = \new_[38137]_  & \new_[38130]_ ;
  assign \new_[38141]_  = A168 & A170;
  assign \new_[38144]_  = A166 & ~A167;
  assign \new_[38145]_  = \new_[38144]_  & \new_[38141]_ ;
  assign \new_[38148]_  = A200 & A199;
  assign \new_[38151]_  = ~A202 & ~A201;
  assign \new_[38152]_  = \new_[38151]_  & \new_[38148]_ ;
  assign \new_[38153]_  = \new_[38152]_  & \new_[38145]_ ;
  assign \new_[38156]_  = A233 & A232;
  assign \new_[38159]_  = ~A236 & A235;
  assign \new_[38160]_  = \new_[38159]_  & \new_[38156]_ ;
  assign \new_[38163]_  = A266 & A265;
  assign \new_[38166]_  = ~A269 & A268;
  assign \new_[38167]_  = \new_[38166]_  & \new_[38163]_ ;
  assign \new_[38168]_  = \new_[38167]_  & \new_[38160]_ ;
  assign \new_[38171]_  = A168 & A170;
  assign \new_[38174]_  = A166 & ~A167;
  assign \new_[38175]_  = \new_[38174]_  & \new_[38171]_ ;
  assign \new_[38178]_  = A200 & A199;
  assign \new_[38181]_  = ~A202 & ~A201;
  assign \new_[38182]_  = \new_[38181]_  & \new_[38178]_ ;
  assign \new_[38183]_  = \new_[38182]_  & \new_[38175]_ ;
  assign \new_[38186]_  = A233 & A232;
  assign \new_[38189]_  = ~A236 & A235;
  assign \new_[38190]_  = \new_[38189]_  & \new_[38186]_ ;
  assign \new_[38193]_  = A266 & ~A265;
  assign \new_[38196]_  = A269 & ~A268;
  assign \new_[38197]_  = \new_[38196]_  & \new_[38193]_ ;
  assign \new_[38198]_  = \new_[38197]_  & \new_[38190]_ ;
  assign \new_[38201]_  = A168 & A170;
  assign \new_[38204]_  = A166 & ~A167;
  assign \new_[38205]_  = \new_[38204]_  & \new_[38201]_ ;
  assign \new_[38208]_  = A200 & A199;
  assign \new_[38211]_  = ~A202 & ~A201;
  assign \new_[38212]_  = \new_[38211]_  & \new_[38208]_ ;
  assign \new_[38213]_  = \new_[38212]_  & \new_[38205]_ ;
  assign \new_[38216]_  = A233 & A232;
  assign \new_[38219]_  = ~A236 & A235;
  assign \new_[38220]_  = \new_[38219]_  & \new_[38216]_ ;
  assign \new_[38223]_  = ~A266 & A265;
  assign \new_[38226]_  = A269 & ~A268;
  assign \new_[38227]_  = \new_[38226]_  & \new_[38223]_ ;
  assign \new_[38228]_  = \new_[38227]_  & \new_[38220]_ ;
  assign \new_[38231]_  = A168 & A170;
  assign \new_[38234]_  = A166 & ~A167;
  assign \new_[38235]_  = \new_[38234]_  & \new_[38231]_ ;
  assign \new_[38238]_  = A200 & A199;
  assign \new_[38241]_  = ~A202 & ~A201;
  assign \new_[38242]_  = \new_[38241]_  & \new_[38238]_ ;
  assign \new_[38243]_  = \new_[38242]_  & \new_[38235]_ ;
  assign \new_[38246]_  = A233 & A232;
  assign \new_[38249]_  = ~A236 & A235;
  assign \new_[38250]_  = \new_[38249]_  & \new_[38246]_ ;
  assign \new_[38253]_  = ~A266 & ~A265;
  assign \new_[38256]_  = ~A269 & A268;
  assign \new_[38257]_  = \new_[38256]_  & \new_[38253]_ ;
  assign \new_[38258]_  = \new_[38257]_  & \new_[38250]_ ;
  assign \new_[38261]_  = A168 & A170;
  assign \new_[38264]_  = A166 & ~A167;
  assign \new_[38265]_  = \new_[38264]_  & \new_[38261]_ ;
  assign \new_[38268]_  = A200 & A199;
  assign \new_[38271]_  = ~A202 & ~A201;
  assign \new_[38272]_  = \new_[38271]_  & \new_[38268]_ ;
  assign \new_[38273]_  = \new_[38272]_  & \new_[38265]_ ;
  assign \new_[38276]_  = A233 & ~A232;
  assign \new_[38279]_  = A236 & ~A235;
  assign \new_[38280]_  = \new_[38279]_  & \new_[38276]_ ;
  assign \new_[38283]_  = A299 & A298;
  assign \new_[38286]_  = ~A302 & A301;
  assign \new_[38287]_  = \new_[38286]_  & \new_[38283]_ ;
  assign \new_[38288]_  = \new_[38287]_  & \new_[38280]_ ;
  assign \new_[38291]_  = A168 & A170;
  assign \new_[38294]_  = A166 & ~A167;
  assign \new_[38295]_  = \new_[38294]_  & \new_[38291]_ ;
  assign \new_[38298]_  = A200 & A199;
  assign \new_[38301]_  = ~A202 & ~A201;
  assign \new_[38302]_  = \new_[38301]_  & \new_[38298]_ ;
  assign \new_[38303]_  = \new_[38302]_  & \new_[38295]_ ;
  assign \new_[38306]_  = A233 & ~A232;
  assign \new_[38309]_  = A236 & ~A235;
  assign \new_[38310]_  = \new_[38309]_  & \new_[38306]_ ;
  assign \new_[38313]_  = ~A299 & A298;
  assign \new_[38316]_  = A302 & ~A301;
  assign \new_[38317]_  = \new_[38316]_  & \new_[38313]_ ;
  assign \new_[38318]_  = \new_[38317]_  & \new_[38310]_ ;
  assign \new_[38321]_  = A168 & A170;
  assign \new_[38324]_  = A166 & ~A167;
  assign \new_[38325]_  = \new_[38324]_  & \new_[38321]_ ;
  assign \new_[38328]_  = A200 & A199;
  assign \new_[38331]_  = ~A202 & ~A201;
  assign \new_[38332]_  = \new_[38331]_  & \new_[38328]_ ;
  assign \new_[38333]_  = \new_[38332]_  & \new_[38325]_ ;
  assign \new_[38336]_  = A233 & ~A232;
  assign \new_[38339]_  = A236 & ~A235;
  assign \new_[38340]_  = \new_[38339]_  & \new_[38336]_ ;
  assign \new_[38343]_  = A299 & ~A298;
  assign \new_[38346]_  = A302 & ~A301;
  assign \new_[38347]_  = \new_[38346]_  & \new_[38343]_ ;
  assign \new_[38348]_  = \new_[38347]_  & \new_[38340]_ ;
  assign \new_[38351]_  = A168 & A170;
  assign \new_[38354]_  = A166 & ~A167;
  assign \new_[38355]_  = \new_[38354]_  & \new_[38351]_ ;
  assign \new_[38358]_  = A200 & A199;
  assign \new_[38361]_  = ~A202 & ~A201;
  assign \new_[38362]_  = \new_[38361]_  & \new_[38358]_ ;
  assign \new_[38363]_  = \new_[38362]_  & \new_[38355]_ ;
  assign \new_[38366]_  = A233 & ~A232;
  assign \new_[38369]_  = A236 & ~A235;
  assign \new_[38370]_  = \new_[38369]_  & \new_[38366]_ ;
  assign \new_[38373]_  = ~A299 & ~A298;
  assign \new_[38376]_  = ~A302 & A301;
  assign \new_[38377]_  = \new_[38376]_  & \new_[38373]_ ;
  assign \new_[38378]_  = \new_[38377]_  & \new_[38370]_ ;
  assign \new_[38381]_  = A168 & A170;
  assign \new_[38384]_  = A166 & ~A167;
  assign \new_[38385]_  = \new_[38384]_  & \new_[38381]_ ;
  assign \new_[38388]_  = A200 & A199;
  assign \new_[38391]_  = ~A202 & ~A201;
  assign \new_[38392]_  = \new_[38391]_  & \new_[38388]_ ;
  assign \new_[38393]_  = \new_[38392]_  & \new_[38385]_ ;
  assign \new_[38396]_  = A233 & ~A232;
  assign \new_[38399]_  = A236 & ~A235;
  assign \new_[38400]_  = \new_[38399]_  & \new_[38396]_ ;
  assign \new_[38403]_  = A266 & A265;
  assign \new_[38406]_  = ~A269 & A268;
  assign \new_[38407]_  = \new_[38406]_  & \new_[38403]_ ;
  assign \new_[38408]_  = \new_[38407]_  & \new_[38400]_ ;
  assign \new_[38411]_  = A168 & A170;
  assign \new_[38414]_  = A166 & ~A167;
  assign \new_[38415]_  = \new_[38414]_  & \new_[38411]_ ;
  assign \new_[38418]_  = A200 & A199;
  assign \new_[38421]_  = ~A202 & ~A201;
  assign \new_[38422]_  = \new_[38421]_  & \new_[38418]_ ;
  assign \new_[38423]_  = \new_[38422]_  & \new_[38415]_ ;
  assign \new_[38426]_  = A233 & ~A232;
  assign \new_[38429]_  = A236 & ~A235;
  assign \new_[38430]_  = \new_[38429]_  & \new_[38426]_ ;
  assign \new_[38433]_  = A266 & ~A265;
  assign \new_[38436]_  = A269 & ~A268;
  assign \new_[38437]_  = \new_[38436]_  & \new_[38433]_ ;
  assign \new_[38438]_  = \new_[38437]_  & \new_[38430]_ ;
  assign \new_[38441]_  = A168 & A170;
  assign \new_[38444]_  = A166 & ~A167;
  assign \new_[38445]_  = \new_[38444]_  & \new_[38441]_ ;
  assign \new_[38448]_  = A200 & A199;
  assign \new_[38451]_  = ~A202 & ~A201;
  assign \new_[38452]_  = \new_[38451]_  & \new_[38448]_ ;
  assign \new_[38453]_  = \new_[38452]_  & \new_[38445]_ ;
  assign \new_[38456]_  = A233 & ~A232;
  assign \new_[38459]_  = A236 & ~A235;
  assign \new_[38460]_  = \new_[38459]_  & \new_[38456]_ ;
  assign \new_[38463]_  = ~A266 & A265;
  assign \new_[38466]_  = A269 & ~A268;
  assign \new_[38467]_  = \new_[38466]_  & \new_[38463]_ ;
  assign \new_[38468]_  = \new_[38467]_  & \new_[38460]_ ;
  assign \new_[38471]_  = A168 & A170;
  assign \new_[38474]_  = A166 & ~A167;
  assign \new_[38475]_  = \new_[38474]_  & \new_[38471]_ ;
  assign \new_[38478]_  = A200 & A199;
  assign \new_[38481]_  = ~A202 & ~A201;
  assign \new_[38482]_  = \new_[38481]_  & \new_[38478]_ ;
  assign \new_[38483]_  = \new_[38482]_  & \new_[38475]_ ;
  assign \new_[38486]_  = A233 & ~A232;
  assign \new_[38489]_  = A236 & ~A235;
  assign \new_[38490]_  = \new_[38489]_  & \new_[38486]_ ;
  assign \new_[38493]_  = ~A266 & ~A265;
  assign \new_[38496]_  = ~A269 & A268;
  assign \new_[38497]_  = \new_[38496]_  & \new_[38493]_ ;
  assign \new_[38498]_  = \new_[38497]_  & \new_[38490]_ ;
  assign \new_[38501]_  = A168 & A170;
  assign \new_[38504]_  = A166 & ~A167;
  assign \new_[38505]_  = \new_[38504]_  & \new_[38501]_ ;
  assign \new_[38508]_  = A200 & A199;
  assign \new_[38511]_  = ~A202 & ~A201;
  assign \new_[38512]_  = \new_[38511]_  & \new_[38508]_ ;
  assign \new_[38513]_  = \new_[38512]_  & \new_[38505]_ ;
  assign \new_[38516]_  = ~A233 & A232;
  assign \new_[38519]_  = A236 & ~A235;
  assign \new_[38520]_  = \new_[38519]_  & \new_[38516]_ ;
  assign \new_[38523]_  = A299 & A298;
  assign \new_[38526]_  = ~A302 & A301;
  assign \new_[38527]_  = \new_[38526]_  & \new_[38523]_ ;
  assign \new_[38528]_  = \new_[38527]_  & \new_[38520]_ ;
  assign \new_[38531]_  = A168 & A170;
  assign \new_[38534]_  = A166 & ~A167;
  assign \new_[38535]_  = \new_[38534]_  & \new_[38531]_ ;
  assign \new_[38538]_  = A200 & A199;
  assign \new_[38541]_  = ~A202 & ~A201;
  assign \new_[38542]_  = \new_[38541]_  & \new_[38538]_ ;
  assign \new_[38543]_  = \new_[38542]_  & \new_[38535]_ ;
  assign \new_[38546]_  = ~A233 & A232;
  assign \new_[38549]_  = A236 & ~A235;
  assign \new_[38550]_  = \new_[38549]_  & \new_[38546]_ ;
  assign \new_[38553]_  = ~A299 & A298;
  assign \new_[38556]_  = A302 & ~A301;
  assign \new_[38557]_  = \new_[38556]_  & \new_[38553]_ ;
  assign \new_[38558]_  = \new_[38557]_  & \new_[38550]_ ;
  assign \new_[38561]_  = A168 & A170;
  assign \new_[38564]_  = A166 & ~A167;
  assign \new_[38565]_  = \new_[38564]_  & \new_[38561]_ ;
  assign \new_[38568]_  = A200 & A199;
  assign \new_[38571]_  = ~A202 & ~A201;
  assign \new_[38572]_  = \new_[38571]_  & \new_[38568]_ ;
  assign \new_[38573]_  = \new_[38572]_  & \new_[38565]_ ;
  assign \new_[38576]_  = ~A233 & A232;
  assign \new_[38579]_  = A236 & ~A235;
  assign \new_[38580]_  = \new_[38579]_  & \new_[38576]_ ;
  assign \new_[38583]_  = A299 & ~A298;
  assign \new_[38586]_  = A302 & ~A301;
  assign \new_[38587]_  = \new_[38586]_  & \new_[38583]_ ;
  assign \new_[38588]_  = \new_[38587]_  & \new_[38580]_ ;
  assign \new_[38591]_  = A168 & A170;
  assign \new_[38594]_  = A166 & ~A167;
  assign \new_[38595]_  = \new_[38594]_  & \new_[38591]_ ;
  assign \new_[38598]_  = A200 & A199;
  assign \new_[38601]_  = ~A202 & ~A201;
  assign \new_[38602]_  = \new_[38601]_  & \new_[38598]_ ;
  assign \new_[38603]_  = \new_[38602]_  & \new_[38595]_ ;
  assign \new_[38606]_  = ~A233 & A232;
  assign \new_[38609]_  = A236 & ~A235;
  assign \new_[38610]_  = \new_[38609]_  & \new_[38606]_ ;
  assign \new_[38613]_  = ~A299 & ~A298;
  assign \new_[38616]_  = ~A302 & A301;
  assign \new_[38617]_  = \new_[38616]_  & \new_[38613]_ ;
  assign \new_[38618]_  = \new_[38617]_  & \new_[38610]_ ;
  assign \new_[38621]_  = A168 & A170;
  assign \new_[38624]_  = A166 & ~A167;
  assign \new_[38625]_  = \new_[38624]_  & \new_[38621]_ ;
  assign \new_[38628]_  = A200 & A199;
  assign \new_[38631]_  = ~A202 & ~A201;
  assign \new_[38632]_  = \new_[38631]_  & \new_[38628]_ ;
  assign \new_[38633]_  = \new_[38632]_  & \new_[38625]_ ;
  assign \new_[38636]_  = ~A233 & A232;
  assign \new_[38639]_  = A236 & ~A235;
  assign \new_[38640]_  = \new_[38639]_  & \new_[38636]_ ;
  assign \new_[38643]_  = A266 & A265;
  assign \new_[38646]_  = ~A269 & A268;
  assign \new_[38647]_  = \new_[38646]_  & \new_[38643]_ ;
  assign \new_[38648]_  = \new_[38647]_  & \new_[38640]_ ;
  assign \new_[38651]_  = A168 & A170;
  assign \new_[38654]_  = A166 & ~A167;
  assign \new_[38655]_  = \new_[38654]_  & \new_[38651]_ ;
  assign \new_[38658]_  = A200 & A199;
  assign \new_[38661]_  = ~A202 & ~A201;
  assign \new_[38662]_  = \new_[38661]_  & \new_[38658]_ ;
  assign \new_[38663]_  = \new_[38662]_  & \new_[38655]_ ;
  assign \new_[38666]_  = ~A233 & A232;
  assign \new_[38669]_  = A236 & ~A235;
  assign \new_[38670]_  = \new_[38669]_  & \new_[38666]_ ;
  assign \new_[38673]_  = A266 & ~A265;
  assign \new_[38676]_  = A269 & ~A268;
  assign \new_[38677]_  = \new_[38676]_  & \new_[38673]_ ;
  assign \new_[38678]_  = \new_[38677]_  & \new_[38670]_ ;
  assign \new_[38681]_  = A168 & A170;
  assign \new_[38684]_  = A166 & ~A167;
  assign \new_[38685]_  = \new_[38684]_  & \new_[38681]_ ;
  assign \new_[38688]_  = A200 & A199;
  assign \new_[38691]_  = ~A202 & ~A201;
  assign \new_[38692]_  = \new_[38691]_  & \new_[38688]_ ;
  assign \new_[38693]_  = \new_[38692]_  & \new_[38685]_ ;
  assign \new_[38696]_  = ~A233 & A232;
  assign \new_[38699]_  = A236 & ~A235;
  assign \new_[38700]_  = \new_[38699]_  & \new_[38696]_ ;
  assign \new_[38703]_  = ~A266 & A265;
  assign \new_[38706]_  = A269 & ~A268;
  assign \new_[38707]_  = \new_[38706]_  & \new_[38703]_ ;
  assign \new_[38708]_  = \new_[38707]_  & \new_[38700]_ ;
  assign \new_[38711]_  = A168 & A170;
  assign \new_[38714]_  = A166 & ~A167;
  assign \new_[38715]_  = \new_[38714]_  & \new_[38711]_ ;
  assign \new_[38718]_  = A200 & A199;
  assign \new_[38721]_  = ~A202 & ~A201;
  assign \new_[38722]_  = \new_[38721]_  & \new_[38718]_ ;
  assign \new_[38723]_  = \new_[38722]_  & \new_[38715]_ ;
  assign \new_[38726]_  = ~A233 & A232;
  assign \new_[38729]_  = A236 & ~A235;
  assign \new_[38730]_  = \new_[38729]_  & \new_[38726]_ ;
  assign \new_[38733]_  = ~A266 & ~A265;
  assign \new_[38736]_  = ~A269 & A268;
  assign \new_[38737]_  = \new_[38736]_  & \new_[38733]_ ;
  assign \new_[38738]_  = \new_[38737]_  & \new_[38730]_ ;
  assign \new_[38741]_  = A168 & A170;
  assign \new_[38744]_  = A166 & ~A167;
  assign \new_[38745]_  = \new_[38744]_  & \new_[38741]_ ;
  assign \new_[38748]_  = A200 & A199;
  assign \new_[38751]_  = ~A202 & ~A201;
  assign \new_[38752]_  = \new_[38751]_  & \new_[38748]_ ;
  assign \new_[38753]_  = \new_[38752]_  & \new_[38745]_ ;
  assign \new_[38756]_  = ~A233 & ~A232;
  assign \new_[38759]_  = ~A236 & A235;
  assign \new_[38760]_  = \new_[38759]_  & \new_[38756]_ ;
  assign \new_[38763]_  = A299 & A298;
  assign \new_[38766]_  = ~A302 & A301;
  assign \new_[38767]_  = \new_[38766]_  & \new_[38763]_ ;
  assign \new_[38768]_  = \new_[38767]_  & \new_[38760]_ ;
  assign \new_[38771]_  = A168 & A170;
  assign \new_[38774]_  = A166 & ~A167;
  assign \new_[38775]_  = \new_[38774]_  & \new_[38771]_ ;
  assign \new_[38778]_  = A200 & A199;
  assign \new_[38781]_  = ~A202 & ~A201;
  assign \new_[38782]_  = \new_[38781]_  & \new_[38778]_ ;
  assign \new_[38783]_  = \new_[38782]_  & \new_[38775]_ ;
  assign \new_[38786]_  = ~A233 & ~A232;
  assign \new_[38789]_  = ~A236 & A235;
  assign \new_[38790]_  = \new_[38789]_  & \new_[38786]_ ;
  assign \new_[38793]_  = ~A299 & A298;
  assign \new_[38796]_  = A302 & ~A301;
  assign \new_[38797]_  = \new_[38796]_  & \new_[38793]_ ;
  assign \new_[38798]_  = \new_[38797]_  & \new_[38790]_ ;
  assign \new_[38801]_  = A168 & A170;
  assign \new_[38804]_  = A166 & ~A167;
  assign \new_[38805]_  = \new_[38804]_  & \new_[38801]_ ;
  assign \new_[38808]_  = A200 & A199;
  assign \new_[38811]_  = ~A202 & ~A201;
  assign \new_[38812]_  = \new_[38811]_  & \new_[38808]_ ;
  assign \new_[38813]_  = \new_[38812]_  & \new_[38805]_ ;
  assign \new_[38816]_  = ~A233 & ~A232;
  assign \new_[38819]_  = ~A236 & A235;
  assign \new_[38820]_  = \new_[38819]_  & \new_[38816]_ ;
  assign \new_[38823]_  = A299 & ~A298;
  assign \new_[38826]_  = A302 & ~A301;
  assign \new_[38827]_  = \new_[38826]_  & \new_[38823]_ ;
  assign \new_[38828]_  = \new_[38827]_  & \new_[38820]_ ;
  assign \new_[38831]_  = A168 & A170;
  assign \new_[38834]_  = A166 & ~A167;
  assign \new_[38835]_  = \new_[38834]_  & \new_[38831]_ ;
  assign \new_[38838]_  = A200 & A199;
  assign \new_[38841]_  = ~A202 & ~A201;
  assign \new_[38842]_  = \new_[38841]_  & \new_[38838]_ ;
  assign \new_[38843]_  = \new_[38842]_  & \new_[38835]_ ;
  assign \new_[38846]_  = ~A233 & ~A232;
  assign \new_[38849]_  = ~A236 & A235;
  assign \new_[38850]_  = \new_[38849]_  & \new_[38846]_ ;
  assign \new_[38853]_  = ~A299 & ~A298;
  assign \new_[38856]_  = ~A302 & A301;
  assign \new_[38857]_  = \new_[38856]_  & \new_[38853]_ ;
  assign \new_[38858]_  = \new_[38857]_  & \new_[38850]_ ;
  assign \new_[38861]_  = A168 & A170;
  assign \new_[38864]_  = A166 & ~A167;
  assign \new_[38865]_  = \new_[38864]_  & \new_[38861]_ ;
  assign \new_[38868]_  = A200 & A199;
  assign \new_[38871]_  = ~A202 & ~A201;
  assign \new_[38872]_  = \new_[38871]_  & \new_[38868]_ ;
  assign \new_[38873]_  = \new_[38872]_  & \new_[38865]_ ;
  assign \new_[38876]_  = ~A233 & ~A232;
  assign \new_[38879]_  = ~A236 & A235;
  assign \new_[38880]_  = \new_[38879]_  & \new_[38876]_ ;
  assign \new_[38883]_  = A266 & A265;
  assign \new_[38886]_  = ~A269 & A268;
  assign \new_[38887]_  = \new_[38886]_  & \new_[38883]_ ;
  assign \new_[38888]_  = \new_[38887]_  & \new_[38880]_ ;
  assign \new_[38891]_  = A168 & A170;
  assign \new_[38894]_  = A166 & ~A167;
  assign \new_[38895]_  = \new_[38894]_  & \new_[38891]_ ;
  assign \new_[38898]_  = A200 & A199;
  assign \new_[38901]_  = ~A202 & ~A201;
  assign \new_[38902]_  = \new_[38901]_  & \new_[38898]_ ;
  assign \new_[38903]_  = \new_[38902]_  & \new_[38895]_ ;
  assign \new_[38906]_  = ~A233 & ~A232;
  assign \new_[38909]_  = ~A236 & A235;
  assign \new_[38910]_  = \new_[38909]_  & \new_[38906]_ ;
  assign \new_[38913]_  = A266 & ~A265;
  assign \new_[38916]_  = A269 & ~A268;
  assign \new_[38917]_  = \new_[38916]_  & \new_[38913]_ ;
  assign \new_[38918]_  = \new_[38917]_  & \new_[38910]_ ;
  assign \new_[38921]_  = A168 & A170;
  assign \new_[38924]_  = A166 & ~A167;
  assign \new_[38925]_  = \new_[38924]_  & \new_[38921]_ ;
  assign \new_[38928]_  = A200 & A199;
  assign \new_[38931]_  = ~A202 & ~A201;
  assign \new_[38932]_  = \new_[38931]_  & \new_[38928]_ ;
  assign \new_[38933]_  = \new_[38932]_  & \new_[38925]_ ;
  assign \new_[38936]_  = ~A233 & ~A232;
  assign \new_[38939]_  = ~A236 & A235;
  assign \new_[38940]_  = \new_[38939]_  & \new_[38936]_ ;
  assign \new_[38943]_  = ~A266 & A265;
  assign \new_[38946]_  = A269 & ~A268;
  assign \new_[38947]_  = \new_[38946]_  & \new_[38943]_ ;
  assign \new_[38948]_  = \new_[38947]_  & \new_[38940]_ ;
  assign \new_[38951]_  = A168 & A170;
  assign \new_[38954]_  = A166 & ~A167;
  assign \new_[38955]_  = \new_[38954]_  & \new_[38951]_ ;
  assign \new_[38958]_  = A200 & A199;
  assign \new_[38961]_  = ~A202 & ~A201;
  assign \new_[38962]_  = \new_[38961]_  & \new_[38958]_ ;
  assign \new_[38963]_  = \new_[38962]_  & \new_[38955]_ ;
  assign \new_[38966]_  = ~A233 & ~A232;
  assign \new_[38969]_  = ~A236 & A235;
  assign \new_[38970]_  = \new_[38969]_  & \new_[38966]_ ;
  assign \new_[38973]_  = ~A266 & ~A265;
  assign \new_[38976]_  = ~A269 & A268;
  assign \new_[38977]_  = \new_[38976]_  & \new_[38973]_ ;
  assign \new_[38978]_  = \new_[38977]_  & \new_[38970]_ ;
  assign \new_[38981]_  = A168 & A170;
  assign \new_[38984]_  = A166 & ~A167;
  assign \new_[38985]_  = \new_[38984]_  & \new_[38981]_ ;
  assign \new_[38988]_  = A200 & A199;
  assign \new_[38991]_  = A203 & ~A201;
  assign \new_[38992]_  = \new_[38991]_  & \new_[38988]_ ;
  assign \new_[38993]_  = \new_[38992]_  & \new_[38985]_ ;
  assign \new_[38996]_  = A233 & A232;
  assign \new_[38999]_  = ~A236 & A235;
  assign \new_[39000]_  = \new_[38999]_  & \new_[38996]_ ;
  assign \new_[39003]_  = A299 & A298;
  assign \new_[39006]_  = ~A302 & A301;
  assign \new_[39007]_  = \new_[39006]_  & \new_[39003]_ ;
  assign \new_[39008]_  = \new_[39007]_  & \new_[39000]_ ;
  assign \new_[39011]_  = A168 & A170;
  assign \new_[39014]_  = A166 & ~A167;
  assign \new_[39015]_  = \new_[39014]_  & \new_[39011]_ ;
  assign \new_[39018]_  = A200 & A199;
  assign \new_[39021]_  = A203 & ~A201;
  assign \new_[39022]_  = \new_[39021]_  & \new_[39018]_ ;
  assign \new_[39023]_  = \new_[39022]_  & \new_[39015]_ ;
  assign \new_[39026]_  = A233 & A232;
  assign \new_[39029]_  = ~A236 & A235;
  assign \new_[39030]_  = \new_[39029]_  & \new_[39026]_ ;
  assign \new_[39033]_  = ~A299 & A298;
  assign \new_[39036]_  = A302 & ~A301;
  assign \new_[39037]_  = \new_[39036]_  & \new_[39033]_ ;
  assign \new_[39038]_  = \new_[39037]_  & \new_[39030]_ ;
  assign \new_[39041]_  = A168 & A170;
  assign \new_[39044]_  = A166 & ~A167;
  assign \new_[39045]_  = \new_[39044]_  & \new_[39041]_ ;
  assign \new_[39048]_  = A200 & A199;
  assign \new_[39051]_  = A203 & ~A201;
  assign \new_[39052]_  = \new_[39051]_  & \new_[39048]_ ;
  assign \new_[39053]_  = \new_[39052]_  & \new_[39045]_ ;
  assign \new_[39056]_  = A233 & A232;
  assign \new_[39059]_  = ~A236 & A235;
  assign \new_[39060]_  = \new_[39059]_  & \new_[39056]_ ;
  assign \new_[39063]_  = A299 & ~A298;
  assign \new_[39066]_  = A302 & ~A301;
  assign \new_[39067]_  = \new_[39066]_  & \new_[39063]_ ;
  assign \new_[39068]_  = \new_[39067]_  & \new_[39060]_ ;
  assign \new_[39071]_  = A168 & A170;
  assign \new_[39074]_  = A166 & ~A167;
  assign \new_[39075]_  = \new_[39074]_  & \new_[39071]_ ;
  assign \new_[39078]_  = A200 & A199;
  assign \new_[39081]_  = A203 & ~A201;
  assign \new_[39082]_  = \new_[39081]_  & \new_[39078]_ ;
  assign \new_[39083]_  = \new_[39082]_  & \new_[39075]_ ;
  assign \new_[39086]_  = A233 & A232;
  assign \new_[39089]_  = ~A236 & A235;
  assign \new_[39090]_  = \new_[39089]_  & \new_[39086]_ ;
  assign \new_[39093]_  = ~A299 & ~A298;
  assign \new_[39096]_  = ~A302 & A301;
  assign \new_[39097]_  = \new_[39096]_  & \new_[39093]_ ;
  assign \new_[39098]_  = \new_[39097]_  & \new_[39090]_ ;
  assign \new_[39101]_  = A168 & A170;
  assign \new_[39104]_  = A166 & ~A167;
  assign \new_[39105]_  = \new_[39104]_  & \new_[39101]_ ;
  assign \new_[39108]_  = A200 & A199;
  assign \new_[39111]_  = A203 & ~A201;
  assign \new_[39112]_  = \new_[39111]_  & \new_[39108]_ ;
  assign \new_[39113]_  = \new_[39112]_  & \new_[39105]_ ;
  assign \new_[39116]_  = A233 & A232;
  assign \new_[39119]_  = ~A236 & A235;
  assign \new_[39120]_  = \new_[39119]_  & \new_[39116]_ ;
  assign \new_[39123]_  = A266 & A265;
  assign \new_[39126]_  = ~A269 & A268;
  assign \new_[39127]_  = \new_[39126]_  & \new_[39123]_ ;
  assign \new_[39128]_  = \new_[39127]_  & \new_[39120]_ ;
  assign \new_[39131]_  = A168 & A170;
  assign \new_[39134]_  = A166 & ~A167;
  assign \new_[39135]_  = \new_[39134]_  & \new_[39131]_ ;
  assign \new_[39138]_  = A200 & A199;
  assign \new_[39141]_  = A203 & ~A201;
  assign \new_[39142]_  = \new_[39141]_  & \new_[39138]_ ;
  assign \new_[39143]_  = \new_[39142]_  & \new_[39135]_ ;
  assign \new_[39146]_  = A233 & A232;
  assign \new_[39149]_  = ~A236 & A235;
  assign \new_[39150]_  = \new_[39149]_  & \new_[39146]_ ;
  assign \new_[39153]_  = A266 & ~A265;
  assign \new_[39156]_  = A269 & ~A268;
  assign \new_[39157]_  = \new_[39156]_  & \new_[39153]_ ;
  assign \new_[39158]_  = \new_[39157]_  & \new_[39150]_ ;
  assign \new_[39161]_  = A168 & A170;
  assign \new_[39164]_  = A166 & ~A167;
  assign \new_[39165]_  = \new_[39164]_  & \new_[39161]_ ;
  assign \new_[39168]_  = A200 & A199;
  assign \new_[39171]_  = A203 & ~A201;
  assign \new_[39172]_  = \new_[39171]_  & \new_[39168]_ ;
  assign \new_[39173]_  = \new_[39172]_  & \new_[39165]_ ;
  assign \new_[39176]_  = A233 & A232;
  assign \new_[39179]_  = ~A236 & A235;
  assign \new_[39180]_  = \new_[39179]_  & \new_[39176]_ ;
  assign \new_[39183]_  = ~A266 & A265;
  assign \new_[39186]_  = A269 & ~A268;
  assign \new_[39187]_  = \new_[39186]_  & \new_[39183]_ ;
  assign \new_[39188]_  = \new_[39187]_  & \new_[39180]_ ;
  assign \new_[39191]_  = A168 & A170;
  assign \new_[39194]_  = A166 & ~A167;
  assign \new_[39195]_  = \new_[39194]_  & \new_[39191]_ ;
  assign \new_[39198]_  = A200 & A199;
  assign \new_[39201]_  = A203 & ~A201;
  assign \new_[39202]_  = \new_[39201]_  & \new_[39198]_ ;
  assign \new_[39203]_  = \new_[39202]_  & \new_[39195]_ ;
  assign \new_[39206]_  = A233 & A232;
  assign \new_[39209]_  = ~A236 & A235;
  assign \new_[39210]_  = \new_[39209]_  & \new_[39206]_ ;
  assign \new_[39213]_  = ~A266 & ~A265;
  assign \new_[39216]_  = ~A269 & A268;
  assign \new_[39217]_  = \new_[39216]_  & \new_[39213]_ ;
  assign \new_[39218]_  = \new_[39217]_  & \new_[39210]_ ;
  assign \new_[39221]_  = A168 & A170;
  assign \new_[39224]_  = A166 & ~A167;
  assign \new_[39225]_  = \new_[39224]_  & \new_[39221]_ ;
  assign \new_[39228]_  = A200 & A199;
  assign \new_[39231]_  = A203 & ~A201;
  assign \new_[39232]_  = \new_[39231]_  & \new_[39228]_ ;
  assign \new_[39233]_  = \new_[39232]_  & \new_[39225]_ ;
  assign \new_[39236]_  = A233 & ~A232;
  assign \new_[39239]_  = A236 & ~A235;
  assign \new_[39240]_  = \new_[39239]_  & \new_[39236]_ ;
  assign \new_[39243]_  = A299 & A298;
  assign \new_[39246]_  = ~A302 & A301;
  assign \new_[39247]_  = \new_[39246]_  & \new_[39243]_ ;
  assign \new_[39248]_  = \new_[39247]_  & \new_[39240]_ ;
  assign \new_[39251]_  = A168 & A170;
  assign \new_[39254]_  = A166 & ~A167;
  assign \new_[39255]_  = \new_[39254]_  & \new_[39251]_ ;
  assign \new_[39258]_  = A200 & A199;
  assign \new_[39261]_  = A203 & ~A201;
  assign \new_[39262]_  = \new_[39261]_  & \new_[39258]_ ;
  assign \new_[39263]_  = \new_[39262]_  & \new_[39255]_ ;
  assign \new_[39266]_  = A233 & ~A232;
  assign \new_[39269]_  = A236 & ~A235;
  assign \new_[39270]_  = \new_[39269]_  & \new_[39266]_ ;
  assign \new_[39273]_  = ~A299 & A298;
  assign \new_[39276]_  = A302 & ~A301;
  assign \new_[39277]_  = \new_[39276]_  & \new_[39273]_ ;
  assign \new_[39278]_  = \new_[39277]_  & \new_[39270]_ ;
  assign \new_[39281]_  = A168 & A170;
  assign \new_[39284]_  = A166 & ~A167;
  assign \new_[39285]_  = \new_[39284]_  & \new_[39281]_ ;
  assign \new_[39288]_  = A200 & A199;
  assign \new_[39291]_  = A203 & ~A201;
  assign \new_[39292]_  = \new_[39291]_  & \new_[39288]_ ;
  assign \new_[39293]_  = \new_[39292]_  & \new_[39285]_ ;
  assign \new_[39296]_  = A233 & ~A232;
  assign \new_[39299]_  = A236 & ~A235;
  assign \new_[39300]_  = \new_[39299]_  & \new_[39296]_ ;
  assign \new_[39303]_  = A299 & ~A298;
  assign \new_[39306]_  = A302 & ~A301;
  assign \new_[39307]_  = \new_[39306]_  & \new_[39303]_ ;
  assign \new_[39308]_  = \new_[39307]_  & \new_[39300]_ ;
  assign \new_[39311]_  = A168 & A170;
  assign \new_[39314]_  = A166 & ~A167;
  assign \new_[39315]_  = \new_[39314]_  & \new_[39311]_ ;
  assign \new_[39318]_  = A200 & A199;
  assign \new_[39321]_  = A203 & ~A201;
  assign \new_[39322]_  = \new_[39321]_  & \new_[39318]_ ;
  assign \new_[39323]_  = \new_[39322]_  & \new_[39315]_ ;
  assign \new_[39326]_  = A233 & ~A232;
  assign \new_[39329]_  = A236 & ~A235;
  assign \new_[39330]_  = \new_[39329]_  & \new_[39326]_ ;
  assign \new_[39333]_  = ~A299 & ~A298;
  assign \new_[39336]_  = ~A302 & A301;
  assign \new_[39337]_  = \new_[39336]_  & \new_[39333]_ ;
  assign \new_[39338]_  = \new_[39337]_  & \new_[39330]_ ;
  assign \new_[39341]_  = A168 & A170;
  assign \new_[39344]_  = A166 & ~A167;
  assign \new_[39345]_  = \new_[39344]_  & \new_[39341]_ ;
  assign \new_[39348]_  = A200 & A199;
  assign \new_[39351]_  = A203 & ~A201;
  assign \new_[39352]_  = \new_[39351]_  & \new_[39348]_ ;
  assign \new_[39353]_  = \new_[39352]_  & \new_[39345]_ ;
  assign \new_[39356]_  = A233 & ~A232;
  assign \new_[39359]_  = A236 & ~A235;
  assign \new_[39360]_  = \new_[39359]_  & \new_[39356]_ ;
  assign \new_[39363]_  = A266 & A265;
  assign \new_[39366]_  = ~A269 & A268;
  assign \new_[39367]_  = \new_[39366]_  & \new_[39363]_ ;
  assign \new_[39368]_  = \new_[39367]_  & \new_[39360]_ ;
  assign \new_[39371]_  = A168 & A170;
  assign \new_[39374]_  = A166 & ~A167;
  assign \new_[39375]_  = \new_[39374]_  & \new_[39371]_ ;
  assign \new_[39378]_  = A200 & A199;
  assign \new_[39381]_  = A203 & ~A201;
  assign \new_[39382]_  = \new_[39381]_  & \new_[39378]_ ;
  assign \new_[39383]_  = \new_[39382]_  & \new_[39375]_ ;
  assign \new_[39386]_  = A233 & ~A232;
  assign \new_[39389]_  = A236 & ~A235;
  assign \new_[39390]_  = \new_[39389]_  & \new_[39386]_ ;
  assign \new_[39393]_  = A266 & ~A265;
  assign \new_[39396]_  = A269 & ~A268;
  assign \new_[39397]_  = \new_[39396]_  & \new_[39393]_ ;
  assign \new_[39398]_  = \new_[39397]_  & \new_[39390]_ ;
  assign \new_[39401]_  = A168 & A170;
  assign \new_[39404]_  = A166 & ~A167;
  assign \new_[39405]_  = \new_[39404]_  & \new_[39401]_ ;
  assign \new_[39408]_  = A200 & A199;
  assign \new_[39411]_  = A203 & ~A201;
  assign \new_[39412]_  = \new_[39411]_  & \new_[39408]_ ;
  assign \new_[39413]_  = \new_[39412]_  & \new_[39405]_ ;
  assign \new_[39416]_  = A233 & ~A232;
  assign \new_[39419]_  = A236 & ~A235;
  assign \new_[39420]_  = \new_[39419]_  & \new_[39416]_ ;
  assign \new_[39423]_  = ~A266 & A265;
  assign \new_[39426]_  = A269 & ~A268;
  assign \new_[39427]_  = \new_[39426]_  & \new_[39423]_ ;
  assign \new_[39428]_  = \new_[39427]_  & \new_[39420]_ ;
  assign \new_[39431]_  = A168 & A170;
  assign \new_[39434]_  = A166 & ~A167;
  assign \new_[39435]_  = \new_[39434]_  & \new_[39431]_ ;
  assign \new_[39438]_  = A200 & A199;
  assign \new_[39441]_  = A203 & ~A201;
  assign \new_[39442]_  = \new_[39441]_  & \new_[39438]_ ;
  assign \new_[39443]_  = \new_[39442]_  & \new_[39435]_ ;
  assign \new_[39446]_  = A233 & ~A232;
  assign \new_[39449]_  = A236 & ~A235;
  assign \new_[39450]_  = \new_[39449]_  & \new_[39446]_ ;
  assign \new_[39453]_  = ~A266 & ~A265;
  assign \new_[39456]_  = ~A269 & A268;
  assign \new_[39457]_  = \new_[39456]_  & \new_[39453]_ ;
  assign \new_[39458]_  = \new_[39457]_  & \new_[39450]_ ;
  assign \new_[39461]_  = A168 & A170;
  assign \new_[39464]_  = A166 & ~A167;
  assign \new_[39465]_  = \new_[39464]_  & \new_[39461]_ ;
  assign \new_[39468]_  = A200 & A199;
  assign \new_[39471]_  = A203 & ~A201;
  assign \new_[39472]_  = \new_[39471]_  & \new_[39468]_ ;
  assign \new_[39473]_  = \new_[39472]_  & \new_[39465]_ ;
  assign \new_[39476]_  = ~A233 & A232;
  assign \new_[39479]_  = A236 & ~A235;
  assign \new_[39480]_  = \new_[39479]_  & \new_[39476]_ ;
  assign \new_[39483]_  = A299 & A298;
  assign \new_[39486]_  = ~A302 & A301;
  assign \new_[39487]_  = \new_[39486]_  & \new_[39483]_ ;
  assign \new_[39488]_  = \new_[39487]_  & \new_[39480]_ ;
  assign \new_[39491]_  = A168 & A170;
  assign \new_[39494]_  = A166 & ~A167;
  assign \new_[39495]_  = \new_[39494]_  & \new_[39491]_ ;
  assign \new_[39498]_  = A200 & A199;
  assign \new_[39501]_  = A203 & ~A201;
  assign \new_[39502]_  = \new_[39501]_  & \new_[39498]_ ;
  assign \new_[39503]_  = \new_[39502]_  & \new_[39495]_ ;
  assign \new_[39506]_  = ~A233 & A232;
  assign \new_[39509]_  = A236 & ~A235;
  assign \new_[39510]_  = \new_[39509]_  & \new_[39506]_ ;
  assign \new_[39513]_  = ~A299 & A298;
  assign \new_[39516]_  = A302 & ~A301;
  assign \new_[39517]_  = \new_[39516]_  & \new_[39513]_ ;
  assign \new_[39518]_  = \new_[39517]_  & \new_[39510]_ ;
  assign \new_[39521]_  = A168 & A170;
  assign \new_[39524]_  = A166 & ~A167;
  assign \new_[39525]_  = \new_[39524]_  & \new_[39521]_ ;
  assign \new_[39528]_  = A200 & A199;
  assign \new_[39531]_  = A203 & ~A201;
  assign \new_[39532]_  = \new_[39531]_  & \new_[39528]_ ;
  assign \new_[39533]_  = \new_[39532]_  & \new_[39525]_ ;
  assign \new_[39536]_  = ~A233 & A232;
  assign \new_[39539]_  = A236 & ~A235;
  assign \new_[39540]_  = \new_[39539]_  & \new_[39536]_ ;
  assign \new_[39543]_  = A299 & ~A298;
  assign \new_[39546]_  = A302 & ~A301;
  assign \new_[39547]_  = \new_[39546]_  & \new_[39543]_ ;
  assign \new_[39548]_  = \new_[39547]_  & \new_[39540]_ ;
  assign \new_[39551]_  = A168 & A170;
  assign \new_[39554]_  = A166 & ~A167;
  assign \new_[39555]_  = \new_[39554]_  & \new_[39551]_ ;
  assign \new_[39558]_  = A200 & A199;
  assign \new_[39561]_  = A203 & ~A201;
  assign \new_[39562]_  = \new_[39561]_  & \new_[39558]_ ;
  assign \new_[39563]_  = \new_[39562]_  & \new_[39555]_ ;
  assign \new_[39566]_  = ~A233 & A232;
  assign \new_[39569]_  = A236 & ~A235;
  assign \new_[39570]_  = \new_[39569]_  & \new_[39566]_ ;
  assign \new_[39573]_  = ~A299 & ~A298;
  assign \new_[39576]_  = ~A302 & A301;
  assign \new_[39577]_  = \new_[39576]_  & \new_[39573]_ ;
  assign \new_[39578]_  = \new_[39577]_  & \new_[39570]_ ;
  assign \new_[39581]_  = A168 & A170;
  assign \new_[39584]_  = A166 & ~A167;
  assign \new_[39585]_  = \new_[39584]_  & \new_[39581]_ ;
  assign \new_[39588]_  = A200 & A199;
  assign \new_[39591]_  = A203 & ~A201;
  assign \new_[39592]_  = \new_[39591]_  & \new_[39588]_ ;
  assign \new_[39593]_  = \new_[39592]_  & \new_[39585]_ ;
  assign \new_[39596]_  = ~A233 & A232;
  assign \new_[39599]_  = A236 & ~A235;
  assign \new_[39600]_  = \new_[39599]_  & \new_[39596]_ ;
  assign \new_[39603]_  = A266 & A265;
  assign \new_[39606]_  = ~A269 & A268;
  assign \new_[39607]_  = \new_[39606]_  & \new_[39603]_ ;
  assign \new_[39608]_  = \new_[39607]_  & \new_[39600]_ ;
  assign \new_[39611]_  = A168 & A170;
  assign \new_[39614]_  = A166 & ~A167;
  assign \new_[39615]_  = \new_[39614]_  & \new_[39611]_ ;
  assign \new_[39618]_  = A200 & A199;
  assign \new_[39621]_  = A203 & ~A201;
  assign \new_[39622]_  = \new_[39621]_  & \new_[39618]_ ;
  assign \new_[39623]_  = \new_[39622]_  & \new_[39615]_ ;
  assign \new_[39626]_  = ~A233 & A232;
  assign \new_[39629]_  = A236 & ~A235;
  assign \new_[39630]_  = \new_[39629]_  & \new_[39626]_ ;
  assign \new_[39633]_  = A266 & ~A265;
  assign \new_[39636]_  = A269 & ~A268;
  assign \new_[39637]_  = \new_[39636]_  & \new_[39633]_ ;
  assign \new_[39638]_  = \new_[39637]_  & \new_[39630]_ ;
  assign \new_[39641]_  = A168 & A170;
  assign \new_[39644]_  = A166 & ~A167;
  assign \new_[39645]_  = \new_[39644]_  & \new_[39641]_ ;
  assign \new_[39648]_  = A200 & A199;
  assign \new_[39651]_  = A203 & ~A201;
  assign \new_[39652]_  = \new_[39651]_  & \new_[39648]_ ;
  assign \new_[39653]_  = \new_[39652]_  & \new_[39645]_ ;
  assign \new_[39656]_  = ~A233 & A232;
  assign \new_[39659]_  = A236 & ~A235;
  assign \new_[39660]_  = \new_[39659]_  & \new_[39656]_ ;
  assign \new_[39663]_  = ~A266 & A265;
  assign \new_[39666]_  = A269 & ~A268;
  assign \new_[39667]_  = \new_[39666]_  & \new_[39663]_ ;
  assign \new_[39668]_  = \new_[39667]_  & \new_[39660]_ ;
  assign \new_[39671]_  = A168 & A170;
  assign \new_[39674]_  = A166 & ~A167;
  assign \new_[39675]_  = \new_[39674]_  & \new_[39671]_ ;
  assign \new_[39678]_  = A200 & A199;
  assign \new_[39681]_  = A203 & ~A201;
  assign \new_[39682]_  = \new_[39681]_  & \new_[39678]_ ;
  assign \new_[39683]_  = \new_[39682]_  & \new_[39675]_ ;
  assign \new_[39686]_  = ~A233 & A232;
  assign \new_[39689]_  = A236 & ~A235;
  assign \new_[39690]_  = \new_[39689]_  & \new_[39686]_ ;
  assign \new_[39693]_  = ~A266 & ~A265;
  assign \new_[39696]_  = ~A269 & A268;
  assign \new_[39697]_  = \new_[39696]_  & \new_[39693]_ ;
  assign \new_[39698]_  = \new_[39697]_  & \new_[39690]_ ;
  assign \new_[39701]_  = A168 & A170;
  assign \new_[39704]_  = A166 & ~A167;
  assign \new_[39705]_  = \new_[39704]_  & \new_[39701]_ ;
  assign \new_[39708]_  = A200 & A199;
  assign \new_[39711]_  = A203 & ~A201;
  assign \new_[39712]_  = \new_[39711]_  & \new_[39708]_ ;
  assign \new_[39713]_  = \new_[39712]_  & \new_[39705]_ ;
  assign \new_[39716]_  = ~A233 & ~A232;
  assign \new_[39719]_  = ~A236 & A235;
  assign \new_[39720]_  = \new_[39719]_  & \new_[39716]_ ;
  assign \new_[39723]_  = A299 & A298;
  assign \new_[39726]_  = ~A302 & A301;
  assign \new_[39727]_  = \new_[39726]_  & \new_[39723]_ ;
  assign \new_[39728]_  = \new_[39727]_  & \new_[39720]_ ;
  assign \new_[39731]_  = A168 & A170;
  assign \new_[39734]_  = A166 & ~A167;
  assign \new_[39735]_  = \new_[39734]_  & \new_[39731]_ ;
  assign \new_[39738]_  = A200 & A199;
  assign \new_[39741]_  = A203 & ~A201;
  assign \new_[39742]_  = \new_[39741]_  & \new_[39738]_ ;
  assign \new_[39743]_  = \new_[39742]_  & \new_[39735]_ ;
  assign \new_[39746]_  = ~A233 & ~A232;
  assign \new_[39749]_  = ~A236 & A235;
  assign \new_[39750]_  = \new_[39749]_  & \new_[39746]_ ;
  assign \new_[39753]_  = ~A299 & A298;
  assign \new_[39756]_  = A302 & ~A301;
  assign \new_[39757]_  = \new_[39756]_  & \new_[39753]_ ;
  assign \new_[39758]_  = \new_[39757]_  & \new_[39750]_ ;
  assign \new_[39761]_  = A168 & A170;
  assign \new_[39764]_  = A166 & ~A167;
  assign \new_[39765]_  = \new_[39764]_  & \new_[39761]_ ;
  assign \new_[39768]_  = A200 & A199;
  assign \new_[39771]_  = A203 & ~A201;
  assign \new_[39772]_  = \new_[39771]_  & \new_[39768]_ ;
  assign \new_[39773]_  = \new_[39772]_  & \new_[39765]_ ;
  assign \new_[39776]_  = ~A233 & ~A232;
  assign \new_[39779]_  = ~A236 & A235;
  assign \new_[39780]_  = \new_[39779]_  & \new_[39776]_ ;
  assign \new_[39783]_  = A299 & ~A298;
  assign \new_[39786]_  = A302 & ~A301;
  assign \new_[39787]_  = \new_[39786]_  & \new_[39783]_ ;
  assign \new_[39788]_  = \new_[39787]_  & \new_[39780]_ ;
  assign \new_[39791]_  = A168 & A170;
  assign \new_[39794]_  = A166 & ~A167;
  assign \new_[39795]_  = \new_[39794]_  & \new_[39791]_ ;
  assign \new_[39798]_  = A200 & A199;
  assign \new_[39801]_  = A203 & ~A201;
  assign \new_[39802]_  = \new_[39801]_  & \new_[39798]_ ;
  assign \new_[39803]_  = \new_[39802]_  & \new_[39795]_ ;
  assign \new_[39806]_  = ~A233 & ~A232;
  assign \new_[39809]_  = ~A236 & A235;
  assign \new_[39810]_  = \new_[39809]_  & \new_[39806]_ ;
  assign \new_[39813]_  = ~A299 & ~A298;
  assign \new_[39816]_  = ~A302 & A301;
  assign \new_[39817]_  = \new_[39816]_  & \new_[39813]_ ;
  assign \new_[39818]_  = \new_[39817]_  & \new_[39810]_ ;
  assign \new_[39821]_  = A168 & A170;
  assign \new_[39824]_  = A166 & ~A167;
  assign \new_[39825]_  = \new_[39824]_  & \new_[39821]_ ;
  assign \new_[39828]_  = A200 & A199;
  assign \new_[39831]_  = A203 & ~A201;
  assign \new_[39832]_  = \new_[39831]_  & \new_[39828]_ ;
  assign \new_[39833]_  = \new_[39832]_  & \new_[39825]_ ;
  assign \new_[39836]_  = ~A233 & ~A232;
  assign \new_[39839]_  = ~A236 & A235;
  assign \new_[39840]_  = \new_[39839]_  & \new_[39836]_ ;
  assign \new_[39843]_  = A266 & A265;
  assign \new_[39846]_  = ~A269 & A268;
  assign \new_[39847]_  = \new_[39846]_  & \new_[39843]_ ;
  assign \new_[39848]_  = \new_[39847]_  & \new_[39840]_ ;
  assign \new_[39851]_  = A168 & A170;
  assign \new_[39854]_  = A166 & ~A167;
  assign \new_[39855]_  = \new_[39854]_  & \new_[39851]_ ;
  assign \new_[39858]_  = A200 & A199;
  assign \new_[39861]_  = A203 & ~A201;
  assign \new_[39862]_  = \new_[39861]_  & \new_[39858]_ ;
  assign \new_[39863]_  = \new_[39862]_  & \new_[39855]_ ;
  assign \new_[39866]_  = ~A233 & ~A232;
  assign \new_[39869]_  = ~A236 & A235;
  assign \new_[39870]_  = \new_[39869]_  & \new_[39866]_ ;
  assign \new_[39873]_  = A266 & ~A265;
  assign \new_[39876]_  = A269 & ~A268;
  assign \new_[39877]_  = \new_[39876]_  & \new_[39873]_ ;
  assign \new_[39878]_  = \new_[39877]_  & \new_[39870]_ ;
  assign \new_[39881]_  = A168 & A170;
  assign \new_[39884]_  = A166 & ~A167;
  assign \new_[39885]_  = \new_[39884]_  & \new_[39881]_ ;
  assign \new_[39888]_  = A200 & A199;
  assign \new_[39891]_  = A203 & ~A201;
  assign \new_[39892]_  = \new_[39891]_  & \new_[39888]_ ;
  assign \new_[39893]_  = \new_[39892]_  & \new_[39885]_ ;
  assign \new_[39896]_  = ~A233 & ~A232;
  assign \new_[39899]_  = ~A236 & A235;
  assign \new_[39900]_  = \new_[39899]_  & \new_[39896]_ ;
  assign \new_[39903]_  = ~A266 & A265;
  assign \new_[39906]_  = A269 & ~A268;
  assign \new_[39907]_  = \new_[39906]_  & \new_[39903]_ ;
  assign \new_[39908]_  = \new_[39907]_  & \new_[39900]_ ;
  assign \new_[39911]_  = A168 & A170;
  assign \new_[39914]_  = A166 & ~A167;
  assign \new_[39915]_  = \new_[39914]_  & \new_[39911]_ ;
  assign \new_[39918]_  = A200 & A199;
  assign \new_[39921]_  = A203 & ~A201;
  assign \new_[39922]_  = \new_[39921]_  & \new_[39918]_ ;
  assign \new_[39923]_  = \new_[39922]_  & \new_[39915]_ ;
  assign \new_[39926]_  = ~A233 & ~A232;
  assign \new_[39929]_  = ~A236 & A235;
  assign \new_[39930]_  = \new_[39929]_  & \new_[39926]_ ;
  assign \new_[39933]_  = ~A266 & ~A265;
  assign \new_[39936]_  = ~A269 & A268;
  assign \new_[39937]_  = \new_[39936]_  & \new_[39933]_ ;
  assign \new_[39938]_  = \new_[39937]_  & \new_[39930]_ ;
  assign \new_[39941]_  = A168 & A170;
  assign \new_[39944]_  = A166 & ~A167;
  assign \new_[39945]_  = \new_[39944]_  & \new_[39941]_ ;
  assign \new_[39948]_  = A200 & ~A199;
  assign \new_[39951]_  = A202 & ~A201;
  assign \new_[39952]_  = \new_[39951]_  & \new_[39948]_ ;
  assign \new_[39953]_  = \new_[39952]_  & \new_[39945]_ ;
  assign \new_[39956]_  = A233 & A232;
  assign \new_[39959]_  = ~A236 & A235;
  assign \new_[39960]_  = \new_[39959]_  & \new_[39956]_ ;
  assign \new_[39963]_  = A299 & A298;
  assign \new_[39966]_  = ~A302 & A301;
  assign \new_[39967]_  = \new_[39966]_  & \new_[39963]_ ;
  assign \new_[39968]_  = \new_[39967]_  & \new_[39960]_ ;
  assign \new_[39971]_  = A168 & A170;
  assign \new_[39974]_  = A166 & ~A167;
  assign \new_[39975]_  = \new_[39974]_  & \new_[39971]_ ;
  assign \new_[39978]_  = A200 & ~A199;
  assign \new_[39981]_  = A202 & ~A201;
  assign \new_[39982]_  = \new_[39981]_  & \new_[39978]_ ;
  assign \new_[39983]_  = \new_[39982]_  & \new_[39975]_ ;
  assign \new_[39986]_  = A233 & A232;
  assign \new_[39989]_  = ~A236 & A235;
  assign \new_[39990]_  = \new_[39989]_  & \new_[39986]_ ;
  assign \new_[39993]_  = ~A299 & A298;
  assign \new_[39996]_  = A302 & ~A301;
  assign \new_[39997]_  = \new_[39996]_  & \new_[39993]_ ;
  assign \new_[39998]_  = \new_[39997]_  & \new_[39990]_ ;
  assign \new_[40001]_  = A168 & A170;
  assign \new_[40004]_  = A166 & ~A167;
  assign \new_[40005]_  = \new_[40004]_  & \new_[40001]_ ;
  assign \new_[40008]_  = A200 & ~A199;
  assign \new_[40011]_  = A202 & ~A201;
  assign \new_[40012]_  = \new_[40011]_  & \new_[40008]_ ;
  assign \new_[40013]_  = \new_[40012]_  & \new_[40005]_ ;
  assign \new_[40016]_  = A233 & A232;
  assign \new_[40019]_  = ~A236 & A235;
  assign \new_[40020]_  = \new_[40019]_  & \new_[40016]_ ;
  assign \new_[40023]_  = A299 & ~A298;
  assign \new_[40026]_  = A302 & ~A301;
  assign \new_[40027]_  = \new_[40026]_  & \new_[40023]_ ;
  assign \new_[40028]_  = \new_[40027]_  & \new_[40020]_ ;
  assign \new_[40031]_  = A168 & A170;
  assign \new_[40034]_  = A166 & ~A167;
  assign \new_[40035]_  = \new_[40034]_  & \new_[40031]_ ;
  assign \new_[40038]_  = A200 & ~A199;
  assign \new_[40041]_  = A202 & ~A201;
  assign \new_[40042]_  = \new_[40041]_  & \new_[40038]_ ;
  assign \new_[40043]_  = \new_[40042]_  & \new_[40035]_ ;
  assign \new_[40046]_  = A233 & A232;
  assign \new_[40049]_  = ~A236 & A235;
  assign \new_[40050]_  = \new_[40049]_  & \new_[40046]_ ;
  assign \new_[40053]_  = ~A299 & ~A298;
  assign \new_[40056]_  = ~A302 & A301;
  assign \new_[40057]_  = \new_[40056]_  & \new_[40053]_ ;
  assign \new_[40058]_  = \new_[40057]_  & \new_[40050]_ ;
  assign \new_[40061]_  = A168 & A170;
  assign \new_[40064]_  = A166 & ~A167;
  assign \new_[40065]_  = \new_[40064]_  & \new_[40061]_ ;
  assign \new_[40068]_  = A200 & ~A199;
  assign \new_[40071]_  = A202 & ~A201;
  assign \new_[40072]_  = \new_[40071]_  & \new_[40068]_ ;
  assign \new_[40073]_  = \new_[40072]_  & \new_[40065]_ ;
  assign \new_[40076]_  = A233 & A232;
  assign \new_[40079]_  = ~A236 & A235;
  assign \new_[40080]_  = \new_[40079]_  & \new_[40076]_ ;
  assign \new_[40083]_  = A266 & A265;
  assign \new_[40086]_  = ~A269 & A268;
  assign \new_[40087]_  = \new_[40086]_  & \new_[40083]_ ;
  assign \new_[40088]_  = \new_[40087]_  & \new_[40080]_ ;
  assign \new_[40091]_  = A168 & A170;
  assign \new_[40094]_  = A166 & ~A167;
  assign \new_[40095]_  = \new_[40094]_  & \new_[40091]_ ;
  assign \new_[40098]_  = A200 & ~A199;
  assign \new_[40101]_  = A202 & ~A201;
  assign \new_[40102]_  = \new_[40101]_  & \new_[40098]_ ;
  assign \new_[40103]_  = \new_[40102]_  & \new_[40095]_ ;
  assign \new_[40106]_  = A233 & A232;
  assign \new_[40109]_  = ~A236 & A235;
  assign \new_[40110]_  = \new_[40109]_  & \new_[40106]_ ;
  assign \new_[40113]_  = A266 & ~A265;
  assign \new_[40116]_  = A269 & ~A268;
  assign \new_[40117]_  = \new_[40116]_  & \new_[40113]_ ;
  assign \new_[40118]_  = \new_[40117]_  & \new_[40110]_ ;
  assign \new_[40121]_  = A168 & A170;
  assign \new_[40124]_  = A166 & ~A167;
  assign \new_[40125]_  = \new_[40124]_  & \new_[40121]_ ;
  assign \new_[40128]_  = A200 & ~A199;
  assign \new_[40131]_  = A202 & ~A201;
  assign \new_[40132]_  = \new_[40131]_  & \new_[40128]_ ;
  assign \new_[40133]_  = \new_[40132]_  & \new_[40125]_ ;
  assign \new_[40136]_  = A233 & A232;
  assign \new_[40139]_  = ~A236 & A235;
  assign \new_[40140]_  = \new_[40139]_  & \new_[40136]_ ;
  assign \new_[40143]_  = ~A266 & A265;
  assign \new_[40146]_  = A269 & ~A268;
  assign \new_[40147]_  = \new_[40146]_  & \new_[40143]_ ;
  assign \new_[40148]_  = \new_[40147]_  & \new_[40140]_ ;
  assign \new_[40151]_  = A168 & A170;
  assign \new_[40154]_  = A166 & ~A167;
  assign \new_[40155]_  = \new_[40154]_  & \new_[40151]_ ;
  assign \new_[40158]_  = A200 & ~A199;
  assign \new_[40161]_  = A202 & ~A201;
  assign \new_[40162]_  = \new_[40161]_  & \new_[40158]_ ;
  assign \new_[40163]_  = \new_[40162]_  & \new_[40155]_ ;
  assign \new_[40166]_  = A233 & A232;
  assign \new_[40169]_  = ~A236 & A235;
  assign \new_[40170]_  = \new_[40169]_  & \new_[40166]_ ;
  assign \new_[40173]_  = ~A266 & ~A265;
  assign \new_[40176]_  = ~A269 & A268;
  assign \new_[40177]_  = \new_[40176]_  & \new_[40173]_ ;
  assign \new_[40178]_  = \new_[40177]_  & \new_[40170]_ ;
  assign \new_[40181]_  = A168 & A170;
  assign \new_[40184]_  = A166 & ~A167;
  assign \new_[40185]_  = \new_[40184]_  & \new_[40181]_ ;
  assign \new_[40188]_  = A200 & ~A199;
  assign \new_[40191]_  = A202 & ~A201;
  assign \new_[40192]_  = \new_[40191]_  & \new_[40188]_ ;
  assign \new_[40193]_  = \new_[40192]_  & \new_[40185]_ ;
  assign \new_[40196]_  = A233 & ~A232;
  assign \new_[40199]_  = A236 & ~A235;
  assign \new_[40200]_  = \new_[40199]_  & \new_[40196]_ ;
  assign \new_[40203]_  = A299 & A298;
  assign \new_[40206]_  = ~A302 & A301;
  assign \new_[40207]_  = \new_[40206]_  & \new_[40203]_ ;
  assign \new_[40208]_  = \new_[40207]_  & \new_[40200]_ ;
  assign \new_[40211]_  = A168 & A170;
  assign \new_[40214]_  = A166 & ~A167;
  assign \new_[40215]_  = \new_[40214]_  & \new_[40211]_ ;
  assign \new_[40218]_  = A200 & ~A199;
  assign \new_[40221]_  = A202 & ~A201;
  assign \new_[40222]_  = \new_[40221]_  & \new_[40218]_ ;
  assign \new_[40223]_  = \new_[40222]_  & \new_[40215]_ ;
  assign \new_[40226]_  = A233 & ~A232;
  assign \new_[40229]_  = A236 & ~A235;
  assign \new_[40230]_  = \new_[40229]_  & \new_[40226]_ ;
  assign \new_[40233]_  = ~A299 & A298;
  assign \new_[40236]_  = A302 & ~A301;
  assign \new_[40237]_  = \new_[40236]_  & \new_[40233]_ ;
  assign \new_[40238]_  = \new_[40237]_  & \new_[40230]_ ;
  assign \new_[40241]_  = A168 & A170;
  assign \new_[40244]_  = A166 & ~A167;
  assign \new_[40245]_  = \new_[40244]_  & \new_[40241]_ ;
  assign \new_[40248]_  = A200 & ~A199;
  assign \new_[40251]_  = A202 & ~A201;
  assign \new_[40252]_  = \new_[40251]_  & \new_[40248]_ ;
  assign \new_[40253]_  = \new_[40252]_  & \new_[40245]_ ;
  assign \new_[40256]_  = A233 & ~A232;
  assign \new_[40259]_  = A236 & ~A235;
  assign \new_[40260]_  = \new_[40259]_  & \new_[40256]_ ;
  assign \new_[40263]_  = A299 & ~A298;
  assign \new_[40266]_  = A302 & ~A301;
  assign \new_[40267]_  = \new_[40266]_  & \new_[40263]_ ;
  assign \new_[40268]_  = \new_[40267]_  & \new_[40260]_ ;
  assign \new_[40271]_  = A168 & A170;
  assign \new_[40274]_  = A166 & ~A167;
  assign \new_[40275]_  = \new_[40274]_  & \new_[40271]_ ;
  assign \new_[40278]_  = A200 & ~A199;
  assign \new_[40281]_  = A202 & ~A201;
  assign \new_[40282]_  = \new_[40281]_  & \new_[40278]_ ;
  assign \new_[40283]_  = \new_[40282]_  & \new_[40275]_ ;
  assign \new_[40286]_  = A233 & ~A232;
  assign \new_[40289]_  = A236 & ~A235;
  assign \new_[40290]_  = \new_[40289]_  & \new_[40286]_ ;
  assign \new_[40293]_  = ~A299 & ~A298;
  assign \new_[40296]_  = ~A302 & A301;
  assign \new_[40297]_  = \new_[40296]_  & \new_[40293]_ ;
  assign \new_[40298]_  = \new_[40297]_  & \new_[40290]_ ;
  assign \new_[40301]_  = A168 & A170;
  assign \new_[40304]_  = A166 & ~A167;
  assign \new_[40305]_  = \new_[40304]_  & \new_[40301]_ ;
  assign \new_[40308]_  = A200 & ~A199;
  assign \new_[40311]_  = A202 & ~A201;
  assign \new_[40312]_  = \new_[40311]_  & \new_[40308]_ ;
  assign \new_[40313]_  = \new_[40312]_  & \new_[40305]_ ;
  assign \new_[40316]_  = A233 & ~A232;
  assign \new_[40319]_  = A236 & ~A235;
  assign \new_[40320]_  = \new_[40319]_  & \new_[40316]_ ;
  assign \new_[40323]_  = A266 & A265;
  assign \new_[40326]_  = ~A269 & A268;
  assign \new_[40327]_  = \new_[40326]_  & \new_[40323]_ ;
  assign \new_[40328]_  = \new_[40327]_  & \new_[40320]_ ;
  assign \new_[40331]_  = A168 & A170;
  assign \new_[40334]_  = A166 & ~A167;
  assign \new_[40335]_  = \new_[40334]_  & \new_[40331]_ ;
  assign \new_[40338]_  = A200 & ~A199;
  assign \new_[40341]_  = A202 & ~A201;
  assign \new_[40342]_  = \new_[40341]_  & \new_[40338]_ ;
  assign \new_[40343]_  = \new_[40342]_  & \new_[40335]_ ;
  assign \new_[40346]_  = A233 & ~A232;
  assign \new_[40349]_  = A236 & ~A235;
  assign \new_[40350]_  = \new_[40349]_  & \new_[40346]_ ;
  assign \new_[40353]_  = A266 & ~A265;
  assign \new_[40356]_  = A269 & ~A268;
  assign \new_[40357]_  = \new_[40356]_  & \new_[40353]_ ;
  assign \new_[40358]_  = \new_[40357]_  & \new_[40350]_ ;
  assign \new_[40361]_  = A168 & A170;
  assign \new_[40364]_  = A166 & ~A167;
  assign \new_[40365]_  = \new_[40364]_  & \new_[40361]_ ;
  assign \new_[40368]_  = A200 & ~A199;
  assign \new_[40371]_  = A202 & ~A201;
  assign \new_[40372]_  = \new_[40371]_  & \new_[40368]_ ;
  assign \new_[40373]_  = \new_[40372]_  & \new_[40365]_ ;
  assign \new_[40376]_  = A233 & ~A232;
  assign \new_[40379]_  = A236 & ~A235;
  assign \new_[40380]_  = \new_[40379]_  & \new_[40376]_ ;
  assign \new_[40383]_  = ~A266 & A265;
  assign \new_[40386]_  = A269 & ~A268;
  assign \new_[40387]_  = \new_[40386]_  & \new_[40383]_ ;
  assign \new_[40388]_  = \new_[40387]_  & \new_[40380]_ ;
  assign \new_[40391]_  = A168 & A170;
  assign \new_[40394]_  = A166 & ~A167;
  assign \new_[40395]_  = \new_[40394]_  & \new_[40391]_ ;
  assign \new_[40398]_  = A200 & ~A199;
  assign \new_[40401]_  = A202 & ~A201;
  assign \new_[40402]_  = \new_[40401]_  & \new_[40398]_ ;
  assign \new_[40403]_  = \new_[40402]_  & \new_[40395]_ ;
  assign \new_[40406]_  = A233 & ~A232;
  assign \new_[40409]_  = A236 & ~A235;
  assign \new_[40410]_  = \new_[40409]_  & \new_[40406]_ ;
  assign \new_[40413]_  = ~A266 & ~A265;
  assign \new_[40416]_  = ~A269 & A268;
  assign \new_[40417]_  = \new_[40416]_  & \new_[40413]_ ;
  assign \new_[40418]_  = \new_[40417]_  & \new_[40410]_ ;
  assign \new_[40421]_  = A168 & A170;
  assign \new_[40424]_  = A166 & ~A167;
  assign \new_[40425]_  = \new_[40424]_  & \new_[40421]_ ;
  assign \new_[40428]_  = A200 & ~A199;
  assign \new_[40431]_  = A202 & ~A201;
  assign \new_[40432]_  = \new_[40431]_  & \new_[40428]_ ;
  assign \new_[40433]_  = \new_[40432]_  & \new_[40425]_ ;
  assign \new_[40436]_  = ~A233 & A232;
  assign \new_[40439]_  = A236 & ~A235;
  assign \new_[40440]_  = \new_[40439]_  & \new_[40436]_ ;
  assign \new_[40443]_  = A299 & A298;
  assign \new_[40446]_  = ~A302 & A301;
  assign \new_[40447]_  = \new_[40446]_  & \new_[40443]_ ;
  assign \new_[40448]_  = \new_[40447]_  & \new_[40440]_ ;
  assign \new_[40451]_  = A168 & A170;
  assign \new_[40454]_  = A166 & ~A167;
  assign \new_[40455]_  = \new_[40454]_  & \new_[40451]_ ;
  assign \new_[40458]_  = A200 & ~A199;
  assign \new_[40461]_  = A202 & ~A201;
  assign \new_[40462]_  = \new_[40461]_  & \new_[40458]_ ;
  assign \new_[40463]_  = \new_[40462]_  & \new_[40455]_ ;
  assign \new_[40466]_  = ~A233 & A232;
  assign \new_[40469]_  = A236 & ~A235;
  assign \new_[40470]_  = \new_[40469]_  & \new_[40466]_ ;
  assign \new_[40473]_  = ~A299 & A298;
  assign \new_[40476]_  = A302 & ~A301;
  assign \new_[40477]_  = \new_[40476]_  & \new_[40473]_ ;
  assign \new_[40478]_  = \new_[40477]_  & \new_[40470]_ ;
  assign \new_[40481]_  = A168 & A170;
  assign \new_[40484]_  = A166 & ~A167;
  assign \new_[40485]_  = \new_[40484]_  & \new_[40481]_ ;
  assign \new_[40488]_  = A200 & ~A199;
  assign \new_[40491]_  = A202 & ~A201;
  assign \new_[40492]_  = \new_[40491]_  & \new_[40488]_ ;
  assign \new_[40493]_  = \new_[40492]_  & \new_[40485]_ ;
  assign \new_[40496]_  = ~A233 & A232;
  assign \new_[40499]_  = A236 & ~A235;
  assign \new_[40500]_  = \new_[40499]_  & \new_[40496]_ ;
  assign \new_[40503]_  = A299 & ~A298;
  assign \new_[40506]_  = A302 & ~A301;
  assign \new_[40507]_  = \new_[40506]_  & \new_[40503]_ ;
  assign \new_[40508]_  = \new_[40507]_  & \new_[40500]_ ;
  assign \new_[40511]_  = A168 & A170;
  assign \new_[40514]_  = A166 & ~A167;
  assign \new_[40515]_  = \new_[40514]_  & \new_[40511]_ ;
  assign \new_[40518]_  = A200 & ~A199;
  assign \new_[40521]_  = A202 & ~A201;
  assign \new_[40522]_  = \new_[40521]_  & \new_[40518]_ ;
  assign \new_[40523]_  = \new_[40522]_  & \new_[40515]_ ;
  assign \new_[40526]_  = ~A233 & A232;
  assign \new_[40529]_  = A236 & ~A235;
  assign \new_[40530]_  = \new_[40529]_  & \new_[40526]_ ;
  assign \new_[40533]_  = ~A299 & ~A298;
  assign \new_[40536]_  = ~A302 & A301;
  assign \new_[40537]_  = \new_[40536]_  & \new_[40533]_ ;
  assign \new_[40538]_  = \new_[40537]_  & \new_[40530]_ ;
  assign \new_[40541]_  = A168 & A170;
  assign \new_[40544]_  = A166 & ~A167;
  assign \new_[40545]_  = \new_[40544]_  & \new_[40541]_ ;
  assign \new_[40548]_  = A200 & ~A199;
  assign \new_[40551]_  = A202 & ~A201;
  assign \new_[40552]_  = \new_[40551]_  & \new_[40548]_ ;
  assign \new_[40553]_  = \new_[40552]_  & \new_[40545]_ ;
  assign \new_[40556]_  = ~A233 & A232;
  assign \new_[40559]_  = A236 & ~A235;
  assign \new_[40560]_  = \new_[40559]_  & \new_[40556]_ ;
  assign \new_[40563]_  = A266 & A265;
  assign \new_[40566]_  = ~A269 & A268;
  assign \new_[40567]_  = \new_[40566]_  & \new_[40563]_ ;
  assign \new_[40568]_  = \new_[40567]_  & \new_[40560]_ ;
  assign \new_[40571]_  = A168 & A170;
  assign \new_[40574]_  = A166 & ~A167;
  assign \new_[40575]_  = \new_[40574]_  & \new_[40571]_ ;
  assign \new_[40578]_  = A200 & ~A199;
  assign \new_[40581]_  = A202 & ~A201;
  assign \new_[40582]_  = \new_[40581]_  & \new_[40578]_ ;
  assign \new_[40583]_  = \new_[40582]_  & \new_[40575]_ ;
  assign \new_[40586]_  = ~A233 & A232;
  assign \new_[40589]_  = A236 & ~A235;
  assign \new_[40590]_  = \new_[40589]_  & \new_[40586]_ ;
  assign \new_[40593]_  = A266 & ~A265;
  assign \new_[40596]_  = A269 & ~A268;
  assign \new_[40597]_  = \new_[40596]_  & \new_[40593]_ ;
  assign \new_[40598]_  = \new_[40597]_  & \new_[40590]_ ;
  assign \new_[40601]_  = A168 & A170;
  assign \new_[40604]_  = A166 & ~A167;
  assign \new_[40605]_  = \new_[40604]_  & \new_[40601]_ ;
  assign \new_[40608]_  = A200 & ~A199;
  assign \new_[40611]_  = A202 & ~A201;
  assign \new_[40612]_  = \new_[40611]_  & \new_[40608]_ ;
  assign \new_[40613]_  = \new_[40612]_  & \new_[40605]_ ;
  assign \new_[40616]_  = ~A233 & A232;
  assign \new_[40619]_  = A236 & ~A235;
  assign \new_[40620]_  = \new_[40619]_  & \new_[40616]_ ;
  assign \new_[40623]_  = ~A266 & A265;
  assign \new_[40626]_  = A269 & ~A268;
  assign \new_[40627]_  = \new_[40626]_  & \new_[40623]_ ;
  assign \new_[40628]_  = \new_[40627]_  & \new_[40620]_ ;
  assign \new_[40631]_  = A168 & A170;
  assign \new_[40634]_  = A166 & ~A167;
  assign \new_[40635]_  = \new_[40634]_  & \new_[40631]_ ;
  assign \new_[40638]_  = A200 & ~A199;
  assign \new_[40641]_  = A202 & ~A201;
  assign \new_[40642]_  = \new_[40641]_  & \new_[40638]_ ;
  assign \new_[40643]_  = \new_[40642]_  & \new_[40635]_ ;
  assign \new_[40646]_  = ~A233 & A232;
  assign \new_[40649]_  = A236 & ~A235;
  assign \new_[40650]_  = \new_[40649]_  & \new_[40646]_ ;
  assign \new_[40653]_  = ~A266 & ~A265;
  assign \new_[40656]_  = ~A269 & A268;
  assign \new_[40657]_  = \new_[40656]_  & \new_[40653]_ ;
  assign \new_[40658]_  = \new_[40657]_  & \new_[40650]_ ;
  assign \new_[40661]_  = A168 & A170;
  assign \new_[40664]_  = A166 & ~A167;
  assign \new_[40665]_  = \new_[40664]_  & \new_[40661]_ ;
  assign \new_[40668]_  = A200 & ~A199;
  assign \new_[40671]_  = A202 & ~A201;
  assign \new_[40672]_  = \new_[40671]_  & \new_[40668]_ ;
  assign \new_[40673]_  = \new_[40672]_  & \new_[40665]_ ;
  assign \new_[40676]_  = ~A233 & ~A232;
  assign \new_[40679]_  = ~A236 & A235;
  assign \new_[40680]_  = \new_[40679]_  & \new_[40676]_ ;
  assign \new_[40683]_  = A299 & A298;
  assign \new_[40686]_  = ~A302 & A301;
  assign \new_[40687]_  = \new_[40686]_  & \new_[40683]_ ;
  assign \new_[40688]_  = \new_[40687]_  & \new_[40680]_ ;
  assign \new_[40691]_  = A168 & A170;
  assign \new_[40694]_  = A166 & ~A167;
  assign \new_[40695]_  = \new_[40694]_  & \new_[40691]_ ;
  assign \new_[40698]_  = A200 & ~A199;
  assign \new_[40701]_  = A202 & ~A201;
  assign \new_[40702]_  = \new_[40701]_  & \new_[40698]_ ;
  assign \new_[40703]_  = \new_[40702]_  & \new_[40695]_ ;
  assign \new_[40706]_  = ~A233 & ~A232;
  assign \new_[40709]_  = ~A236 & A235;
  assign \new_[40710]_  = \new_[40709]_  & \new_[40706]_ ;
  assign \new_[40713]_  = ~A299 & A298;
  assign \new_[40716]_  = A302 & ~A301;
  assign \new_[40717]_  = \new_[40716]_  & \new_[40713]_ ;
  assign \new_[40718]_  = \new_[40717]_  & \new_[40710]_ ;
  assign \new_[40721]_  = A168 & A170;
  assign \new_[40724]_  = A166 & ~A167;
  assign \new_[40725]_  = \new_[40724]_  & \new_[40721]_ ;
  assign \new_[40728]_  = A200 & ~A199;
  assign \new_[40731]_  = A202 & ~A201;
  assign \new_[40732]_  = \new_[40731]_  & \new_[40728]_ ;
  assign \new_[40733]_  = \new_[40732]_  & \new_[40725]_ ;
  assign \new_[40736]_  = ~A233 & ~A232;
  assign \new_[40739]_  = ~A236 & A235;
  assign \new_[40740]_  = \new_[40739]_  & \new_[40736]_ ;
  assign \new_[40743]_  = A299 & ~A298;
  assign \new_[40746]_  = A302 & ~A301;
  assign \new_[40747]_  = \new_[40746]_  & \new_[40743]_ ;
  assign \new_[40748]_  = \new_[40747]_  & \new_[40740]_ ;
  assign \new_[40751]_  = A168 & A170;
  assign \new_[40754]_  = A166 & ~A167;
  assign \new_[40755]_  = \new_[40754]_  & \new_[40751]_ ;
  assign \new_[40758]_  = A200 & ~A199;
  assign \new_[40761]_  = A202 & ~A201;
  assign \new_[40762]_  = \new_[40761]_  & \new_[40758]_ ;
  assign \new_[40763]_  = \new_[40762]_  & \new_[40755]_ ;
  assign \new_[40766]_  = ~A233 & ~A232;
  assign \new_[40769]_  = ~A236 & A235;
  assign \new_[40770]_  = \new_[40769]_  & \new_[40766]_ ;
  assign \new_[40773]_  = ~A299 & ~A298;
  assign \new_[40776]_  = ~A302 & A301;
  assign \new_[40777]_  = \new_[40776]_  & \new_[40773]_ ;
  assign \new_[40778]_  = \new_[40777]_  & \new_[40770]_ ;
  assign \new_[40781]_  = A168 & A170;
  assign \new_[40784]_  = A166 & ~A167;
  assign \new_[40785]_  = \new_[40784]_  & \new_[40781]_ ;
  assign \new_[40788]_  = A200 & ~A199;
  assign \new_[40791]_  = A202 & ~A201;
  assign \new_[40792]_  = \new_[40791]_  & \new_[40788]_ ;
  assign \new_[40793]_  = \new_[40792]_  & \new_[40785]_ ;
  assign \new_[40796]_  = ~A233 & ~A232;
  assign \new_[40799]_  = ~A236 & A235;
  assign \new_[40800]_  = \new_[40799]_  & \new_[40796]_ ;
  assign \new_[40803]_  = A266 & A265;
  assign \new_[40806]_  = ~A269 & A268;
  assign \new_[40807]_  = \new_[40806]_  & \new_[40803]_ ;
  assign \new_[40808]_  = \new_[40807]_  & \new_[40800]_ ;
  assign \new_[40811]_  = A168 & A170;
  assign \new_[40814]_  = A166 & ~A167;
  assign \new_[40815]_  = \new_[40814]_  & \new_[40811]_ ;
  assign \new_[40818]_  = A200 & ~A199;
  assign \new_[40821]_  = A202 & ~A201;
  assign \new_[40822]_  = \new_[40821]_  & \new_[40818]_ ;
  assign \new_[40823]_  = \new_[40822]_  & \new_[40815]_ ;
  assign \new_[40826]_  = ~A233 & ~A232;
  assign \new_[40829]_  = ~A236 & A235;
  assign \new_[40830]_  = \new_[40829]_  & \new_[40826]_ ;
  assign \new_[40833]_  = A266 & ~A265;
  assign \new_[40836]_  = A269 & ~A268;
  assign \new_[40837]_  = \new_[40836]_  & \new_[40833]_ ;
  assign \new_[40838]_  = \new_[40837]_  & \new_[40830]_ ;
  assign \new_[40841]_  = A168 & A170;
  assign \new_[40844]_  = A166 & ~A167;
  assign \new_[40845]_  = \new_[40844]_  & \new_[40841]_ ;
  assign \new_[40848]_  = A200 & ~A199;
  assign \new_[40851]_  = A202 & ~A201;
  assign \new_[40852]_  = \new_[40851]_  & \new_[40848]_ ;
  assign \new_[40853]_  = \new_[40852]_  & \new_[40845]_ ;
  assign \new_[40856]_  = ~A233 & ~A232;
  assign \new_[40859]_  = ~A236 & A235;
  assign \new_[40860]_  = \new_[40859]_  & \new_[40856]_ ;
  assign \new_[40863]_  = ~A266 & A265;
  assign \new_[40866]_  = A269 & ~A268;
  assign \new_[40867]_  = \new_[40866]_  & \new_[40863]_ ;
  assign \new_[40868]_  = \new_[40867]_  & \new_[40860]_ ;
  assign \new_[40871]_  = A168 & A170;
  assign \new_[40874]_  = A166 & ~A167;
  assign \new_[40875]_  = \new_[40874]_  & \new_[40871]_ ;
  assign \new_[40878]_  = A200 & ~A199;
  assign \new_[40881]_  = A202 & ~A201;
  assign \new_[40882]_  = \new_[40881]_  & \new_[40878]_ ;
  assign \new_[40883]_  = \new_[40882]_  & \new_[40875]_ ;
  assign \new_[40886]_  = ~A233 & ~A232;
  assign \new_[40889]_  = ~A236 & A235;
  assign \new_[40890]_  = \new_[40889]_  & \new_[40886]_ ;
  assign \new_[40893]_  = ~A266 & ~A265;
  assign \new_[40896]_  = ~A269 & A268;
  assign \new_[40897]_  = \new_[40896]_  & \new_[40893]_ ;
  assign \new_[40898]_  = \new_[40897]_  & \new_[40890]_ ;
  assign \new_[40901]_  = A168 & A170;
  assign \new_[40904]_  = A166 & ~A167;
  assign \new_[40905]_  = \new_[40904]_  & \new_[40901]_ ;
  assign \new_[40908]_  = A200 & ~A199;
  assign \new_[40911]_  = ~A203 & ~A201;
  assign \new_[40912]_  = \new_[40911]_  & \new_[40908]_ ;
  assign \new_[40913]_  = \new_[40912]_  & \new_[40905]_ ;
  assign \new_[40916]_  = A233 & A232;
  assign \new_[40919]_  = ~A236 & A235;
  assign \new_[40920]_  = \new_[40919]_  & \new_[40916]_ ;
  assign \new_[40923]_  = A299 & A298;
  assign \new_[40926]_  = ~A302 & A301;
  assign \new_[40927]_  = \new_[40926]_  & \new_[40923]_ ;
  assign \new_[40928]_  = \new_[40927]_  & \new_[40920]_ ;
  assign \new_[40931]_  = A168 & A170;
  assign \new_[40934]_  = A166 & ~A167;
  assign \new_[40935]_  = \new_[40934]_  & \new_[40931]_ ;
  assign \new_[40938]_  = A200 & ~A199;
  assign \new_[40941]_  = ~A203 & ~A201;
  assign \new_[40942]_  = \new_[40941]_  & \new_[40938]_ ;
  assign \new_[40943]_  = \new_[40942]_  & \new_[40935]_ ;
  assign \new_[40946]_  = A233 & A232;
  assign \new_[40949]_  = ~A236 & A235;
  assign \new_[40950]_  = \new_[40949]_  & \new_[40946]_ ;
  assign \new_[40953]_  = ~A299 & A298;
  assign \new_[40956]_  = A302 & ~A301;
  assign \new_[40957]_  = \new_[40956]_  & \new_[40953]_ ;
  assign \new_[40958]_  = \new_[40957]_  & \new_[40950]_ ;
  assign \new_[40961]_  = A168 & A170;
  assign \new_[40964]_  = A166 & ~A167;
  assign \new_[40965]_  = \new_[40964]_  & \new_[40961]_ ;
  assign \new_[40968]_  = A200 & ~A199;
  assign \new_[40971]_  = ~A203 & ~A201;
  assign \new_[40972]_  = \new_[40971]_  & \new_[40968]_ ;
  assign \new_[40973]_  = \new_[40972]_  & \new_[40965]_ ;
  assign \new_[40976]_  = A233 & A232;
  assign \new_[40979]_  = ~A236 & A235;
  assign \new_[40980]_  = \new_[40979]_  & \new_[40976]_ ;
  assign \new_[40983]_  = A299 & ~A298;
  assign \new_[40986]_  = A302 & ~A301;
  assign \new_[40987]_  = \new_[40986]_  & \new_[40983]_ ;
  assign \new_[40988]_  = \new_[40987]_  & \new_[40980]_ ;
  assign \new_[40991]_  = A168 & A170;
  assign \new_[40994]_  = A166 & ~A167;
  assign \new_[40995]_  = \new_[40994]_  & \new_[40991]_ ;
  assign \new_[40998]_  = A200 & ~A199;
  assign \new_[41001]_  = ~A203 & ~A201;
  assign \new_[41002]_  = \new_[41001]_  & \new_[40998]_ ;
  assign \new_[41003]_  = \new_[41002]_  & \new_[40995]_ ;
  assign \new_[41006]_  = A233 & A232;
  assign \new_[41009]_  = ~A236 & A235;
  assign \new_[41010]_  = \new_[41009]_  & \new_[41006]_ ;
  assign \new_[41013]_  = ~A299 & ~A298;
  assign \new_[41016]_  = ~A302 & A301;
  assign \new_[41017]_  = \new_[41016]_  & \new_[41013]_ ;
  assign \new_[41018]_  = \new_[41017]_  & \new_[41010]_ ;
  assign \new_[41021]_  = A168 & A170;
  assign \new_[41024]_  = A166 & ~A167;
  assign \new_[41025]_  = \new_[41024]_  & \new_[41021]_ ;
  assign \new_[41028]_  = A200 & ~A199;
  assign \new_[41031]_  = ~A203 & ~A201;
  assign \new_[41032]_  = \new_[41031]_  & \new_[41028]_ ;
  assign \new_[41033]_  = \new_[41032]_  & \new_[41025]_ ;
  assign \new_[41036]_  = A233 & A232;
  assign \new_[41039]_  = ~A236 & A235;
  assign \new_[41040]_  = \new_[41039]_  & \new_[41036]_ ;
  assign \new_[41043]_  = A266 & A265;
  assign \new_[41046]_  = ~A269 & A268;
  assign \new_[41047]_  = \new_[41046]_  & \new_[41043]_ ;
  assign \new_[41048]_  = \new_[41047]_  & \new_[41040]_ ;
  assign \new_[41051]_  = A168 & A170;
  assign \new_[41054]_  = A166 & ~A167;
  assign \new_[41055]_  = \new_[41054]_  & \new_[41051]_ ;
  assign \new_[41058]_  = A200 & ~A199;
  assign \new_[41061]_  = ~A203 & ~A201;
  assign \new_[41062]_  = \new_[41061]_  & \new_[41058]_ ;
  assign \new_[41063]_  = \new_[41062]_  & \new_[41055]_ ;
  assign \new_[41066]_  = A233 & A232;
  assign \new_[41069]_  = ~A236 & A235;
  assign \new_[41070]_  = \new_[41069]_  & \new_[41066]_ ;
  assign \new_[41073]_  = A266 & ~A265;
  assign \new_[41076]_  = A269 & ~A268;
  assign \new_[41077]_  = \new_[41076]_  & \new_[41073]_ ;
  assign \new_[41078]_  = \new_[41077]_  & \new_[41070]_ ;
  assign \new_[41081]_  = A168 & A170;
  assign \new_[41084]_  = A166 & ~A167;
  assign \new_[41085]_  = \new_[41084]_  & \new_[41081]_ ;
  assign \new_[41088]_  = A200 & ~A199;
  assign \new_[41091]_  = ~A203 & ~A201;
  assign \new_[41092]_  = \new_[41091]_  & \new_[41088]_ ;
  assign \new_[41093]_  = \new_[41092]_  & \new_[41085]_ ;
  assign \new_[41096]_  = A233 & A232;
  assign \new_[41099]_  = ~A236 & A235;
  assign \new_[41100]_  = \new_[41099]_  & \new_[41096]_ ;
  assign \new_[41103]_  = ~A266 & A265;
  assign \new_[41106]_  = A269 & ~A268;
  assign \new_[41107]_  = \new_[41106]_  & \new_[41103]_ ;
  assign \new_[41108]_  = \new_[41107]_  & \new_[41100]_ ;
  assign \new_[41111]_  = A168 & A170;
  assign \new_[41114]_  = A166 & ~A167;
  assign \new_[41115]_  = \new_[41114]_  & \new_[41111]_ ;
  assign \new_[41118]_  = A200 & ~A199;
  assign \new_[41121]_  = ~A203 & ~A201;
  assign \new_[41122]_  = \new_[41121]_  & \new_[41118]_ ;
  assign \new_[41123]_  = \new_[41122]_  & \new_[41115]_ ;
  assign \new_[41126]_  = A233 & A232;
  assign \new_[41129]_  = ~A236 & A235;
  assign \new_[41130]_  = \new_[41129]_  & \new_[41126]_ ;
  assign \new_[41133]_  = ~A266 & ~A265;
  assign \new_[41136]_  = ~A269 & A268;
  assign \new_[41137]_  = \new_[41136]_  & \new_[41133]_ ;
  assign \new_[41138]_  = \new_[41137]_  & \new_[41130]_ ;
  assign \new_[41141]_  = A168 & A170;
  assign \new_[41144]_  = A166 & ~A167;
  assign \new_[41145]_  = \new_[41144]_  & \new_[41141]_ ;
  assign \new_[41148]_  = A200 & ~A199;
  assign \new_[41151]_  = ~A203 & ~A201;
  assign \new_[41152]_  = \new_[41151]_  & \new_[41148]_ ;
  assign \new_[41153]_  = \new_[41152]_  & \new_[41145]_ ;
  assign \new_[41156]_  = A233 & ~A232;
  assign \new_[41159]_  = A236 & ~A235;
  assign \new_[41160]_  = \new_[41159]_  & \new_[41156]_ ;
  assign \new_[41163]_  = A299 & A298;
  assign \new_[41166]_  = ~A302 & A301;
  assign \new_[41167]_  = \new_[41166]_  & \new_[41163]_ ;
  assign \new_[41168]_  = \new_[41167]_  & \new_[41160]_ ;
  assign \new_[41171]_  = A168 & A170;
  assign \new_[41174]_  = A166 & ~A167;
  assign \new_[41175]_  = \new_[41174]_  & \new_[41171]_ ;
  assign \new_[41178]_  = A200 & ~A199;
  assign \new_[41181]_  = ~A203 & ~A201;
  assign \new_[41182]_  = \new_[41181]_  & \new_[41178]_ ;
  assign \new_[41183]_  = \new_[41182]_  & \new_[41175]_ ;
  assign \new_[41186]_  = A233 & ~A232;
  assign \new_[41189]_  = A236 & ~A235;
  assign \new_[41190]_  = \new_[41189]_  & \new_[41186]_ ;
  assign \new_[41193]_  = ~A299 & A298;
  assign \new_[41196]_  = A302 & ~A301;
  assign \new_[41197]_  = \new_[41196]_  & \new_[41193]_ ;
  assign \new_[41198]_  = \new_[41197]_  & \new_[41190]_ ;
  assign \new_[41201]_  = A168 & A170;
  assign \new_[41204]_  = A166 & ~A167;
  assign \new_[41205]_  = \new_[41204]_  & \new_[41201]_ ;
  assign \new_[41208]_  = A200 & ~A199;
  assign \new_[41211]_  = ~A203 & ~A201;
  assign \new_[41212]_  = \new_[41211]_  & \new_[41208]_ ;
  assign \new_[41213]_  = \new_[41212]_  & \new_[41205]_ ;
  assign \new_[41216]_  = A233 & ~A232;
  assign \new_[41219]_  = A236 & ~A235;
  assign \new_[41220]_  = \new_[41219]_  & \new_[41216]_ ;
  assign \new_[41223]_  = A299 & ~A298;
  assign \new_[41226]_  = A302 & ~A301;
  assign \new_[41227]_  = \new_[41226]_  & \new_[41223]_ ;
  assign \new_[41228]_  = \new_[41227]_  & \new_[41220]_ ;
  assign \new_[41231]_  = A168 & A170;
  assign \new_[41234]_  = A166 & ~A167;
  assign \new_[41235]_  = \new_[41234]_  & \new_[41231]_ ;
  assign \new_[41238]_  = A200 & ~A199;
  assign \new_[41241]_  = ~A203 & ~A201;
  assign \new_[41242]_  = \new_[41241]_  & \new_[41238]_ ;
  assign \new_[41243]_  = \new_[41242]_  & \new_[41235]_ ;
  assign \new_[41246]_  = A233 & ~A232;
  assign \new_[41249]_  = A236 & ~A235;
  assign \new_[41250]_  = \new_[41249]_  & \new_[41246]_ ;
  assign \new_[41253]_  = ~A299 & ~A298;
  assign \new_[41256]_  = ~A302 & A301;
  assign \new_[41257]_  = \new_[41256]_  & \new_[41253]_ ;
  assign \new_[41258]_  = \new_[41257]_  & \new_[41250]_ ;
  assign \new_[41261]_  = A168 & A170;
  assign \new_[41264]_  = A166 & ~A167;
  assign \new_[41265]_  = \new_[41264]_  & \new_[41261]_ ;
  assign \new_[41268]_  = A200 & ~A199;
  assign \new_[41271]_  = ~A203 & ~A201;
  assign \new_[41272]_  = \new_[41271]_  & \new_[41268]_ ;
  assign \new_[41273]_  = \new_[41272]_  & \new_[41265]_ ;
  assign \new_[41276]_  = A233 & ~A232;
  assign \new_[41279]_  = A236 & ~A235;
  assign \new_[41280]_  = \new_[41279]_  & \new_[41276]_ ;
  assign \new_[41283]_  = A266 & A265;
  assign \new_[41286]_  = ~A269 & A268;
  assign \new_[41287]_  = \new_[41286]_  & \new_[41283]_ ;
  assign \new_[41288]_  = \new_[41287]_  & \new_[41280]_ ;
  assign \new_[41291]_  = A168 & A170;
  assign \new_[41294]_  = A166 & ~A167;
  assign \new_[41295]_  = \new_[41294]_  & \new_[41291]_ ;
  assign \new_[41298]_  = A200 & ~A199;
  assign \new_[41301]_  = ~A203 & ~A201;
  assign \new_[41302]_  = \new_[41301]_  & \new_[41298]_ ;
  assign \new_[41303]_  = \new_[41302]_  & \new_[41295]_ ;
  assign \new_[41306]_  = A233 & ~A232;
  assign \new_[41309]_  = A236 & ~A235;
  assign \new_[41310]_  = \new_[41309]_  & \new_[41306]_ ;
  assign \new_[41313]_  = A266 & ~A265;
  assign \new_[41316]_  = A269 & ~A268;
  assign \new_[41317]_  = \new_[41316]_  & \new_[41313]_ ;
  assign \new_[41318]_  = \new_[41317]_  & \new_[41310]_ ;
  assign \new_[41321]_  = A168 & A170;
  assign \new_[41324]_  = A166 & ~A167;
  assign \new_[41325]_  = \new_[41324]_  & \new_[41321]_ ;
  assign \new_[41328]_  = A200 & ~A199;
  assign \new_[41331]_  = ~A203 & ~A201;
  assign \new_[41332]_  = \new_[41331]_  & \new_[41328]_ ;
  assign \new_[41333]_  = \new_[41332]_  & \new_[41325]_ ;
  assign \new_[41336]_  = A233 & ~A232;
  assign \new_[41339]_  = A236 & ~A235;
  assign \new_[41340]_  = \new_[41339]_  & \new_[41336]_ ;
  assign \new_[41343]_  = ~A266 & A265;
  assign \new_[41346]_  = A269 & ~A268;
  assign \new_[41347]_  = \new_[41346]_  & \new_[41343]_ ;
  assign \new_[41348]_  = \new_[41347]_  & \new_[41340]_ ;
  assign \new_[41351]_  = A168 & A170;
  assign \new_[41354]_  = A166 & ~A167;
  assign \new_[41355]_  = \new_[41354]_  & \new_[41351]_ ;
  assign \new_[41358]_  = A200 & ~A199;
  assign \new_[41361]_  = ~A203 & ~A201;
  assign \new_[41362]_  = \new_[41361]_  & \new_[41358]_ ;
  assign \new_[41363]_  = \new_[41362]_  & \new_[41355]_ ;
  assign \new_[41366]_  = A233 & ~A232;
  assign \new_[41369]_  = A236 & ~A235;
  assign \new_[41370]_  = \new_[41369]_  & \new_[41366]_ ;
  assign \new_[41373]_  = ~A266 & ~A265;
  assign \new_[41376]_  = ~A269 & A268;
  assign \new_[41377]_  = \new_[41376]_  & \new_[41373]_ ;
  assign \new_[41378]_  = \new_[41377]_  & \new_[41370]_ ;
  assign \new_[41381]_  = A168 & A170;
  assign \new_[41384]_  = A166 & ~A167;
  assign \new_[41385]_  = \new_[41384]_  & \new_[41381]_ ;
  assign \new_[41388]_  = A200 & ~A199;
  assign \new_[41391]_  = ~A203 & ~A201;
  assign \new_[41392]_  = \new_[41391]_  & \new_[41388]_ ;
  assign \new_[41393]_  = \new_[41392]_  & \new_[41385]_ ;
  assign \new_[41396]_  = ~A233 & A232;
  assign \new_[41399]_  = A236 & ~A235;
  assign \new_[41400]_  = \new_[41399]_  & \new_[41396]_ ;
  assign \new_[41403]_  = A299 & A298;
  assign \new_[41406]_  = ~A302 & A301;
  assign \new_[41407]_  = \new_[41406]_  & \new_[41403]_ ;
  assign \new_[41408]_  = \new_[41407]_  & \new_[41400]_ ;
  assign \new_[41411]_  = A168 & A170;
  assign \new_[41414]_  = A166 & ~A167;
  assign \new_[41415]_  = \new_[41414]_  & \new_[41411]_ ;
  assign \new_[41418]_  = A200 & ~A199;
  assign \new_[41421]_  = ~A203 & ~A201;
  assign \new_[41422]_  = \new_[41421]_  & \new_[41418]_ ;
  assign \new_[41423]_  = \new_[41422]_  & \new_[41415]_ ;
  assign \new_[41426]_  = ~A233 & A232;
  assign \new_[41429]_  = A236 & ~A235;
  assign \new_[41430]_  = \new_[41429]_  & \new_[41426]_ ;
  assign \new_[41433]_  = ~A299 & A298;
  assign \new_[41436]_  = A302 & ~A301;
  assign \new_[41437]_  = \new_[41436]_  & \new_[41433]_ ;
  assign \new_[41438]_  = \new_[41437]_  & \new_[41430]_ ;
  assign \new_[41441]_  = A168 & A170;
  assign \new_[41444]_  = A166 & ~A167;
  assign \new_[41445]_  = \new_[41444]_  & \new_[41441]_ ;
  assign \new_[41448]_  = A200 & ~A199;
  assign \new_[41451]_  = ~A203 & ~A201;
  assign \new_[41452]_  = \new_[41451]_  & \new_[41448]_ ;
  assign \new_[41453]_  = \new_[41452]_  & \new_[41445]_ ;
  assign \new_[41456]_  = ~A233 & A232;
  assign \new_[41459]_  = A236 & ~A235;
  assign \new_[41460]_  = \new_[41459]_  & \new_[41456]_ ;
  assign \new_[41463]_  = A299 & ~A298;
  assign \new_[41466]_  = A302 & ~A301;
  assign \new_[41467]_  = \new_[41466]_  & \new_[41463]_ ;
  assign \new_[41468]_  = \new_[41467]_  & \new_[41460]_ ;
  assign \new_[41471]_  = A168 & A170;
  assign \new_[41474]_  = A166 & ~A167;
  assign \new_[41475]_  = \new_[41474]_  & \new_[41471]_ ;
  assign \new_[41478]_  = A200 & ~A199;
  assign \new_[41481]_  = ~A203 & ~A201;
  assign \new_[41482]_  = \new_[41481]_  & \new_[41478]_ ;
  assign \new_[41483]_  = \new_[41482]_  & \new_[41475]_ ;
  assign \new_[41486]_  = ~A233 & A232;
  assign \new_[41489]_  = A236 & ~A235;
  assign \new_[41490]_  = \new_[41489]_  & \new_[41486]_ ;
  assign \new_[41493]_  = ~A299 & ~A298;
  assign \new_[41496]_  = ~A302 & A301;
  assign \new_[41497]_  = \new_[41496]_  & \new_[41493]_ ;
  assign \new_[41498]_  = \new_[41497]_  & \new_[41490]_ ;
  assign \new_[41501]_  = A168 & A170;
  assign \new_[41504]_  = A166 & ~A167;
  assign \new_[41505]_  = \new_[41504]_  & \new_[41501]_ ;
  assign \new_[41508]_  = A200 & ~A199;
  assign \new_[41511]_  = ~A203 & ~A201;
  assign \new_[41512]_  = \new_[41511]_  & \new_[41508]_ ;
  assign \new_[41513]_  = \new_[41512]_  & \new_[41505]_ ;
  assign \new_[41516]_  = ~A233 & A232;
  assign \new_[41519]_  = A236 & ~A235;
  assign \new_[41520]_  = \new_[41519]_  & \new_[41516]_ ;
  assign \new_[41523]_  = A266 & A265;
  assign \new_[41526]_  = ~A269 & A268;
  assign \new_[41527]_  = \new_[41526]_  & \new_[41523]_ ;
  assign \new_[41528]_  = \new_[41527]_  & \new_[41520]_ ;
  assign \new_[41531]_  = A168 & A170;
  assign \new_[41534]_  = A166 & ~A167;
  assign \new_[41535]_  = \new_[41534]_  & \new_[41531]_ ;
  assign \new_[41538]_  = A200 & ~A199;
  assign \new_[41541]_  = ~A203 & ~A201;
  assign \new_[41542]_  = \new_[41541]_  & \new_[41538]_ ;
  assign \new_[41543]_  = \new_[41542]_  & \new_[41535]_ ;
  assign \new_[41546]_  = ~A233 & A232;
  assign \new_[41549]_  = A236 & ~A235;
  assign \new_[41550]_  = \new_[41549]_  & \new_[41546]_ ;
  assign \new_[41553]_  = A266 & ~A265;
  assign \new_[41556]_  = A269 & ~A268;
  assign \new_[41557]_  = \new_[41556]_  & \new_[41553]_ ;
  assign \new_[41558]_  = \new_[41557]_  & \new_[41550]_ ;
  assign \new_[41561]_  = A168 & A170;
  assign \new_[41564]_  = A166 & ~A167;
  assign \new_[41565]_  = \new_[41564]_  & \new_[41561]_ ;
  assign \new_[41568]_  = A200 & ~A199;
  assign \new_[41571]_  = ~A203 & ~A201;
  assign \new_[41572]_  = \new_[41571]_  & \new_[41568]_ ;
  assign \new_[41573]_  = \new_[41572]_  & \new_[41565]_ ;
  assign \new_[41576]_  = ~A233 & A232;
  assign \new_[41579]_  = A236 & ~A235;
  assign \new_[41580]_  = \new_[41579]_  & \new_[41576]_ ;
  assign \new_[41583]_  = ~A266 & A265;
  assign \new_[41586]_  = A269 & ~A268;
  assign \new_[41587]_  = \new_[41586]_  & \new_[41583]_ ;
  assign \new_[41588]_  = \new_[41587]_  & \new_[41580]_ ;
  assign \new_[41591]_  = A168 & A170;
  assign \new_[41594]_  = A166 & ~A167;
  assign \new_[41595]_  = \new_[41594]_  & \new_[41591]_ ;
  assign \new_[41598]_  = A200 & ~A199;
  assign \new_[41601]_  = ~A203 & ~A201;
  assign \new_[41602]_  = \new_[41601]_  & \new_[41598]_ ;
  assign \new_[41603]_  = \new_[41602]_  & \new_[41595]_ ;
  assign \new_[41606]_  = ~A233 & A232;
  assign \new_[41609]_  = A236 & ~A235;
  assign \new_[41610]_  = \new_[41609]_  & \new_[41606]_ ;
  assign \new_[41613]_  = ~A266 & ~A265;
  assign \new_[41616]_  = ~A269 & A268;
  assign \new_[41617]_  = \new_[41616]_  & \new_[41613]_ ;
  assign \new_[41618]_  = \new_[41617]_  & \new_[41610]_ ;
  assign \new_[41621]_  = A168 & A170;
  assign \new_[41624]_  = A166 & ~A167;
  assign \new_[41625]_  = \new_[41624]_  & \new_[41621]_ ;
  assign \new_[41628]_  = A200 & ~A199;
  assign \new_[41631]_  = ~A203 & ~A201;
  assign \new_[41632]_  = \new_[41631]_  & \new_[41628]_ ;
  assign \new_[41633]_  = \new_[41632]_  & \new_[41625]_ ;
  assign \new_[41636]_  = ~A233 & ~A232;
  assign \new_[41639]_  = ~A236 & A235;
  assign \new_[41640]_  = \new_[41639]_  & \new_[41636]_ ;
  assign \new_[41643]_  = A299 & A298;
  assign \new_[41646]_  = ~A302 & A301;
  assign \new_[41647]_  = \new_[41646]_  & \new_[41643]_ ;
  assign \new_[41648]_  = \new_[41647]_  & \new_[41640]_ ;
  assign \new_[41651]_  = A168 & A170;
  assign \new_[41654]_  = A166 & ~A167;
  assign \new_[41655]_  = \new_[41654]_  & \new_[41651]_ ;
  assign \new_[41658]_  = A200 & ~A199;
  assign \new_[41661]_  = ~A203 & ~A201;
  assign \new_[41662]_  = \new_[41661]_  & \new_[41658]_ ;
  assign \new_[41663]_  = \new_[41662]_  & \new_[41655]_ ;
  assign \new_[41666]_  = ~A233 & ~A232;
  assign \new_[41669]_  = ~A236 & A235;
  assign \new_[41670]_  = \new_[41669]_  & \new_[41666]_ ;
  assign \new_[41673]_  = ~A299 & A298;
  assign \new_[41676]_  = A302 & ~A301;
  assign \new_[41677]_  = \new_[41676]_  & \new_[41673]_ ;
  assign \new_[41678]_  = \new_[41677]_  & \new_[41670]_ ;
  assign \new_[41681]_  = A168 & A170;
  assign \new_[41684]_  = A166 & ~A167;
  assign \new_[41685]_  = \new_[41684]_  & \new_[41681]_ ;
  assign \new_[41688]_  = A200 & ~A199;
  assign \new_[41691]_  = ~A203 & ~A201;
  assign \new_[41692]_  = \new_[41691]_  & \new_[41688]_ ;
  assign \new_[41693]_  = \new_[41692]_  & \new_[41685]_ ;
  assign \new_[41696]_  = ~A233 & ~A232;
  assign \new_[41699]_  = ~A236 & A235;
  assign \new_[41700]_  = \new_[41699]_  & \new_[41696]_ ;
  assign \new_[41703]_  = A299 & ~A298;
  assign \new_[41706]_  = A302 & ~A301;
  assign \new_[41707]_  = \new_[41706]_  & \new_[41703]_ ;
  assign \new_[41708]_  = \new_[41707]_  & \new_[41700]_ ;
  assign \new_[41711]_  = A168 & A170;
  assign \new_[41714]_  = A166 & ~A167;
  assign \new_[41715]_  = \new_[41714]_  & \new_[41711]_ ;
  assign \new_[41718]_  = A200 & ~A199;
  assign \new_[41721]_  = ~A203 & ~A201;
  assign \new_[41722]_  = \new_[41721]_  & \new_[41718]_ ;
  assign \new_[41723]_  = \new_[41722]_  & \new_[41715]_ ;
  assign \new_[41726]_  = ~A233 & ~A232;
  assign \new_[41729]_  = ~A236 & A235;
  assign \new_[41730]_  = \new_[41729]_  & \new_[41726]_ ;
  assign \new_[41733]_  = ~A299 & ~A298;
  assign \new_[41736]_  = ~A302 & A301;
  assign \new_[41737]_  = \new_[41736]_  & \new_[41733]_ ;
  assign \new_[41738]_  = \new_[41737]_  & \new_[41730]_ ;
  assign \new_[41741]_  = A168 & A170;
  assign \new_[41744]_  = A166 & ~A167;
  assign \new_[41745]_  = \new_[41744]_  & \new_[41741]_ ;
  assign \new_[41748]_  = A200 & ~A199;
  assign \new_[41751]_  = ~A203 & ~A201;
  assign \new_[41752]_  = \new_[41751]_  & \new_[41748]_ ;
  assign \new_[41753]_  = \new_[41752]_  & \new_[41745]_ ;
  assign \new_[41756]_  = ~A233 & ~A232;
  assign \new_[41759]_  = ~A236 & A235;
  assign \new_[41760]_  = \new_[41759]_  & \new_[41756]_ ;
  assign \new_[41763]_  = A266 & A265;
  assign \new_[41766]_  = ~A269 & A268;
  assign \new_[41767]_  = \new_[41766]_  & \new_[41763]_ ;
  assign \new_[41768]_  = \new_[41767]_  & \new_[41760]_ ;
  assign \new_[41771]_  = A168 & A170;
  assign \new_[41774]_  = A166 & ~A167;
  assign \new_[41775]_  = \new_[41774]_  & \new_[41771]_ ;
  assign \new_[41778]_  = A200 & ~A199;
  assign \new_[41781]_  = ~A203 & ~A201;
  assign \new_[41782]_  = \new_[41781]_  & \new_[41778]_ ;
  assign \new_[41783]_  = \new_[41782]_  & \new_[41775]_ ;
  assign \new_[41786]_  = ~A233 & ~A232;
  assign \new_[41789]_  = ~A236 & A235;
  assign \new_[41790]_  = \new_[41789]_  & \new_[41786]_ ;
  assign \new_[41793]_  = A266 & ~A265;
  assign \new_[41796]_  = A269 & ~A268;
  assign \new_[41797]_  = \new_[41796]_  & \new_[41793]_ ;
  assign \new_[41798]_  = \new_[41797]_  & \new_[41790]_ ;
  assign \new_[41801]_  = A168 & A170;
  assign \new_[41804]_  = A166 & ~A167;
  assign \new_[41805]_  = \new_[41804]_  & \new_[41801]_ ;
  assign \new_[41808]_  = A200 & ~A199;
  assign \new_[41811]_  = ~A203 & ~A201;
  assign \new_[41812]_  = \new_[41811]_  & \new_[41808]_ ;
  assign \new_[41813]_  = \new_[41812]_  & \new_[41805]_ ;
  assign \new_[41816]_  = ~A233 & ~A232;
  assign \new_[41819]_  = ~A236 & A235;
  assign \new_[41820]_  = \new_[41819]_  & \new_[41816]_ ;
  assign \new_[41823]_  = ~A266 & A265;
  assign \new_[41826]_  = A269 & ~A268;
  assign \new_[41827]_  = \new_[41826]_  & \new_[41823]_ ;
  assign \new_[41828]_  = \new_[41827]_  & \new_[41820]_ ;
  assign \new_[41831]_  = A168 & A170;
  assign \new_[41834]_  = A166 & ~A167;
  assign \new_[41835]_  = \new_[41834]_  & \new_[41831]_ ;
  assign \new_[41838]_  = A200 & ~A199;
  assign \new_[41841]_  = ~A203 & ~A201;
  assign \new_[41842]_  = \new_[41841]_  & \new_[41838]_ ;
  assign \new_[41843]_  = \new_[41842]_  & \new_[41835]_ ;
  assign \new_[41846]_  = ~A233 & ~A232;
  assign \new_[41849]_  = ~A236 & A235;
  assign \new_[41850]_  = \new_[41849]_  & \new_[41846]_ ;
  assign \new_[41853]_  = ~A266 & ~A265;
  assign \new_[41856]_  = ~A269 & A268;
  assign \new_[41857]_  = \new_[41856]_  & \new_[41853]_ ;
  assign \new_[41858]_  = \new_[41857]_  & \new_[41850]_ ;
  assign \new_[41861]_  = A168 & A170;
  assign \new_[41864]_  = A166 & ~A167;
  assign \new_[41865]_  = \new_[41864]_  & \new_[41861]_ ;
  assign \new_[41868]_  = ~A200 & A199;
  assign \new_[41871]_  = A202 & ~A201;
  assign \new_[41872]_  = \new_[41871]_  & \new_[41868]_ ;
  assign \new_[41873]_  = \new_[41872]_  & \new_[41865]_ ;
  assign \new_[41876]_  = A233 & A232;
  assign \new_[41879]_  = ~A236 & A235;
  assign \new_[41880]_  = \new_[41879]_  & \new_[41876]_ ;
  assign \new_[41883]_  = A299 & A298;
  assign \new_[41886]_  = ~A302 & A301;
  assign \new_[41887]_  = \new_[41886]_  & \new_[41883]_ ;
  assign \new_[41888]_  = \new_[41887]_  & \new_[41880]_ ;
  assign \new_[41891]_  = A168 & A170;
  assign \new_[41894]_  = A166 & ~A167;
  assign \new_[41895]_  = \new_[41894]_  & \new_[41891]_ ;
  assign \new_[41898]_  = ~A200 & A199;
  assign \new_[41901]_  = A202 & ~A201;
  assign \new_[41902]_  = \new_[41901]_  & \new_[41898]_ ;
  assign \new_[41903]_  = \new_[41902]_  & \new_[41895]_ ;
  assign \new_[41906]_  = A233 & A232;
  assign \new_[41909]_  = ~A236 & A235;
  assign \new_[41910]_  = \new_[41909]_  & \new_[41906]_ ;
  assign \new_[41913]_  = ~A299 & A298;
  assign \new_[41916]_  = A302 & ~A301;
  assign \new_[41917]_  = \new_[41916]_  & \new_[41913]_ ;
  assign \new_[41918]_  = \new_[41917]_  & \new_[41910]_ ;
  assign \new_[41921]_  = A168 & A170;
  assign \new_[41924]_  = A166 & ~A167;
  assign \new_[41925]_  = \new_[41924]_  & \new_[41921]_ ;
  assign \new_[41928]_  = ~A200 & A199;
  assign \new_[41931]_  = A202 & ~A201;
  assign \new_[41932]_  = \new_[41931]_  & \new_[41928]_ ;
  assign \new_[41933]_  = \new_[41932]_  & \new_[41925]_ ;
  assign \new_[41936]_  = A233 & A232;
  assign \new_[41939]_  = ~A236 & A235;
  assign \new_[41940]_  = \new_[41939]_  & \new_[41936]_ ;
  assign \new_[41943]_  = A299 & ~A298;
  assign \new_[41946]_  = A302 & ~A301;
  assign \new_[41947]_  = \new_[41946]_  & \new_[41943]_ ;
  assign \new_[41948]_  = \new_[41947]_  & \new_[41940]_ ;
  assign \new_[41951]_  = A168 & A170;
  assign \new_[41954]_  = A166 & ~A167;
  assign \new_[41955]_  = \new_[41954]_  & \new_[41951]_ ;
  assign \new_[41958]_  = ~A200 & A199;
  assign \new_[41961]_  = A202 & ~A201;
  assign \new_[41962]_  = \new_[41961]_  & \new_[41958]_ ;
  assign \new_[41963]_  = \new_[41962]_  & \new_[41955]_ ;
  assign \new_[41966]_  = A233 & A232;
  assign \new_[41969]_  = ~A236 & A235;
  assign \new_[41970]_  = \new_[41969]_  & \new_[41966]_ ;
  assign \new_[41973]_  = ~A299 & ~A298;
  assign \new_[41976]_  = ~A302 & A301;
  assign \new_[41977]_  = \new_[41976]_  & \new_[41973]_ ;
  assign \new_[41978]_  = \new_[41977]_  & \new_[41970]_ ;
  assign \new_[41981]_  = A168 & A170;
  assign \new_[41984]_  = A166 & ~A167;
  assign \new_[41985]_  = \new_[41984]_  & \new_[41981]_ ;
  assign \new_[41988]_  = ~A200 & A199;
  assign \new_[41991]_  = A202 & ~A201;
  assign \new_[41992]_  = \new_[41991]_  & \new_[41988]_ ;
  assign \new_[41993]_  = \new_[41992]_  & \new_[41985]_ ;
  assign \new_[41996]_  = A233 & A232;
  assign \new_[41999]_  = ~A236 & A235;
  assign \new_[42000]_  = \new_[41999]_  & \new_[41996]_ ;
  assign \new_[42003]_  = A266 & A265;
  assign \new_[42006]_  = ~A269 & A268;
  assign \new_[42007]_  = \new_[42006]_  & \new_[42003]_ ;
  assign \new_[42008]_  = \new_[42007]_  & \new_[42000]_ ;
  assign \new_[42011]_  = A168 & A170;
  assign \new_[42014]_  = A166 & ~A167;
  assign \new_[42015]_  = \new_[42014]_  & \new_[42011]_ ;
  assign \new_[42018]_  = ~A200 & A199;
  assign \new_[42021]_  = A202 & ~A201;
  assign \new_[42022]_  = \new_[42021]_  & \new_[42018]_ ;
  assign \new_[42023]_  = \new_[42022]_  & \new_[42015]_ ;
  assign \new_[42026]_  = A233 & A232;
  assign \new_[42029]_  = ~A236 & A235;
  assign \new_[42030]_  = \new_[42029]_  & \new_[42026]_ ;
  assign \new_[42033]_  = A266 & ~A265;
  assign \new_[42036]_  = A269 & ~A268;
  assign \new_[42037]_  = \new_[42036]_  & \new_[42033]_ ;
  assign \new_[42038]_  = \new_[42037]_  & \new_[42030]_ ;
  assign \new_[42041]_  = A168 & A170;
  assign \new_[42044]_  = A166 & ~A167;
  assign \new_[42045]_  = \new_[42044]_  & \new_[42041]_ ;
  assign \new_[42048]_  = ~A200 & A199;
  assign \new_[42051]_  = A202 & ~A201;
  assign \new_[42052]_  = \new_[42051]_  & \new_[42048]_ ;
  assign \new_[42053]_  = \new_[42052]_  & \new_[42045]_ ;
  assign \new_[42056]_  = A233 & A232;
  assign \new_[42059]_  = ~A236 & A235;
  assign \new_[42060]_  = \new_[42059]_  & \new_[42056]_ ;
  assign \new_[42063]_  = ~A266 & A265;
  assign \new_[42066]_  = A269 & ~A268;
  assign \new_[42067]_  = \new_[42066]_  & \new_[42063]_ ;
  assign \new_[42068]_  = \new_[42067]_  & \new_[42060]_ ;
  assign \new_[42071]_  = A168 & A170;
  assign \new_[42074]_  = A166 & ~A167;
  assign \new_[42075]_  = \new_[42074]_  & \new_[42071]_ ;
  assign \new_[42078]_  = ~A200 & A199;
  assign \new_[42081]_  = A202 & ~A201;
  assign \new_[42082]_  = \new_[42081]_  & \new_[42078]_ ;
  assign \new_[42083]_  = \new_[42082]_  & \new_[42075]_ ;
  assign \new_[42086]_  = A233 & A232;
  assign \new_[42089]_  = ~A236 & A235;
  assign \new_[42090]_  = \new_[42089]_  & \new_[42086]_ ;
  assign \new_[42093]_  = ~A266 & ~A265;
  assign \new_[42096]_  = ~A269 & A268;
  assign \new_[42097]_  = \new_[42096]_  & \new_[42093]_ ;
  assign \new_[42098]_  = \new_[42097]_  & \new_[42090]_ ;
  assign \new_[42101]_  = A168 & A170;
  assign \new_[42104]_  = A166 & ~A167;
  assign \new_[42105]_  = \new_[42104]_  & \new_[42101]_ ;
  assign \new_[42108]_  = ~A200 & A199;
  assign \new_[42111]_  = A202 & ~A201;
  assign \new_[42112]_  = \new_[42111]_  & \new_[42108]_ ;
  assign \new_[42113]_  = \new_[42112]_  & \new_[42105]_ ;
  assign \new_[42116]_  = A233 & ~A232;
  assign \new_[42119]_  = A236 & ~A235;
  assign \new_[42120]_  = \new_[42119]_  & \new_[42116]_ ;
  assign \new_[42123]_  = A299 & A298;
  assign \new_[42126]_  = ~A302 & A301;
  assign \new_[42127]_  = \new_[42126]_  & \new_[42123]_ ;
  assign \new_[42128]_  = \new_[42127]_  & \new_[42120]_ ;
  assign \new_[42131]_  = A168 & A170;
  assign \new_[42134]_  = A166 & ~A167;
  assign \new_[42135]_  = \new_[42134]_  & \new_[42131]_ ;
  assign \new_[42138]_  = ~A200 & A199;
  assign \new_[42141]_  = A202 & ~A201;
  assign \new_[42142]_  = \new_[42141]_  & \new_[42138]_ ;
  assign \new_[42143]_  = \new_[42142]_  & \new_[42135]_ ;
  assign \new_[42146]_  = A233 & ~A232;
  assign \new_[42149]_  = A236 & ~A235;
  assign \new_[42150]_  = \new_[42149]_  & \new_[42146]_ ;
  assign \new_[42153]_  = ~A299 & A298;
  assign \new_[42156]_  = A302 & ~A301;
  assign \new_[42157]_  = \new_[42156]_  & \new_[42153]_ ;
  assign \new_[42158]_  = \new_[42157]_  & \new_[42150]_ ;
  assign \new_[42161]_  = A168 & A170;
  assign \new_[42164]_  = A166 & ~A167;
  assign \new_[42165]_  = \new_[42164]_  & \new_[42161]_ ;
  assign \new_[42168]_  = ~A200 & A199;
  assign \new_[42171]_  = A202 & ~A201;
  assign \new_[42172]_  = \new_[42171]_  & \new_[42168]_ ;
  assign \new_[42173]_  = \new_[42172]_  & \new_[42165]_ ;
  assign \new_[42176]_  = A233 & ~A232;
  assign \new_[42179]_  = A236 & ~A235;
  assign \new_[42180]_  = \new_[42179]_  & \new_[42176]_ ;
  assign \new_[42183]_  = A299 & ~A298;
  assign \new_[42186]_  = A302 & ~A301;
  assign \new_[42187]_  = \new_[42186]_  & \new_[42183]_ ;
  assign \new_[42188]_  = \new_[42187]_  & \new_[42180]_ ;
  assign \new_[42191]_  = A168 & A170;
  assign \new_[42194]_  = A166 & ~A167;
  assign \new_[42195]_  = \new_[42194]_  & \new_[42191]_ ;
  assign \new_[42198]_  = ~A200 & A199;
  assign \new_[42201]_  = A202 & ~A201;
  assign \new_[42202]_  = \new_[42201]_  & \new_[42198]_ ;
  assign \new_[42203]_  = \new_[42202]_  & \new_[42195]_ ;
  assign \new_[42206]_  = A233 & ~A232;
  assign \new_[42209]_  = A236 & ~A235;
  assign \new_[42210]_  = \new_[42209]_  & \new_[42206]_ ;
  assign \new_[42213]_  = ~A299 & ~A298;
  assign \new_[42216]_  = ~A302 & A301;
  assign \new_[42217]_  = \new_[42216]_  & \new_[42213]_ ;
  assign \new_[42218]_  = \new_[42217]_  & \new_[42210]_ ;
  assign \new_[42221]_  = A168 & A170;
  assign \new_[42224]_  = A166 & ~A167;
  assign \new_[42225]_  = \new_[42224]_  & \new_[42221]_ ;
  assign \new_[42228]_  = ~A200 & A199;
  assign \new_[42231]_  = A202 & ~A201;
  assign \new_[42232]_  = \new_[42231]_  & \new_[42228]_ ;
  assign \new_[42233]_  = \new_[42232]_  & \new_[42225]_ ;
  assign \new_[42236]_  = A233 & ~A232;
  assign \new_[42239]_  = A236 & ~A235;
  assign \new_[42240]_  = \new_[42239]_  & \new_[42236]_ ;
  assign \new_[42243]_  = A266 & A265;
  assign \new_[42246]_  = ~A269 & A268;
  assign \new_[42247]_  = \new_[42246]_  & \new_[42243]_ ;
  assign \new_[42248]_  = \new_[42247]_  & \new_[42240]_ ;
  assign \new_[42251]_  = A168 & A170;
  assign \new_[42254]_  = A166 & ~A167;
  assign \new_[42255]_  = \new_[42254]_  & \new_[42251]_ ;
  assign \new_[42258]_  = ~A200 & A199;
  assign \new_[42261]_  = A202 & ~A201;
  assign \new_[42262]_  = \new_[42261]_  & \new_[42258]_ ;
  assign \new_[42263]_  = \new_[42262]_  & \new_[42255]_ ;
  assign \new_[42266]_  = A233 & ~A232;
  assign \new_[42269]_  = A236 & ~A235;
  assign \new_[42270]_  = \new_[42269]_  & \new_[42266]_ ;
  assign \new_[42273]_  = A266 & ~A265;
  assign \new_[42276]_  = A269 & ~A268;
  assign \new_[42277]_  = \new_[42276]_  & \new_[42273]_ ;
  assign \new_[42278]_  = \new_[42277]_  & \new_[42270]_ ;
  assign \new_[42281]_  = A168 & A170;
  assign \new_[42284]_  = A166 & ~A167;
  assign \new_[42285]_  = \new_[42284]_  & \new_[42281]_ ;
  assign \new_[42288]_  = ~A200 & A199;
  assign \new_[42291]_  = A202 & ~A201;
  assign \new_[42292]_  = \new_[42291]_  & \new_[42288]_ ;
  assign \new_[42293]_  = \new_[42292]_  & \new_[42285]_ ;
  assign \new_[42296]_  = A233 & ~A232;
  assign \new_[42299]_  = A236 & ~A235;
  assign \new_[42300]_  = \new_[42299]_  & \new_[42296]_ ;
  assign \new_[42303]_  = ~A266 & A265;
  assign \new_[42306]_  = A269 & ~A268;
  assign \new_[42307]_  = \new_[42306]_  & \new_[42303]_ ;
  assign \new_[42308]_  = \new_[42307]_  & \new_[42300]_ ;
  assign \new_[42311]_  = A168 & A170;
  assign \new_[42314]_  = A166 & ~A167;
  assign \new_[42315]_  = \new_[42314]_  & \new_[42311]_ ;
  assign \new_[42318]_  = ~A200 & A199;
  assign \new_[42321]_  = A202 & ~A201;
  assign \new_[42322]_  = \new_[42321]_  & \new_[42318]_ ;
  assign \new_[42323]_  = \new_[42322]_  & \new_[42315]_ ;
  assign \new_[42326]_  = A233 & ~A232;
  assign \new_[42329]_  = A236 & ~A235;
  assign \new_[42330]_  = \new_[42329]_  & \new_[42326]_ ;
  assign \new_[42333]_  = ~A266 & ~A265;
  assign \new_[42336]_  = ~A269 & A268;
  assign \new_[42337]_  = \new_[42336]_  & \new_[42333]_ ;
  assign \new_[42338]_  = \new_[42337]_  & \new_[42330]_ ;
  assign \new_[42341]_  = A168 & A170;
  assign \new_[42344]_  = A166 & ~A167;
  assign \new_[42345]_  = \new_[42344]_  & \new_[42341]_ ;
  assign \new_[42348]_  = ~A200 & A199;
  assign \new_[42351]_  = A202 & ~A201;
  assign \new_[42352]_  = \new_[42351]_  & \new_[42348]_ ;
  assign \new_[42353]_  = \new_[42352]_  & \new_[42345]_ ;
  assign \new_[42356]_  = ~A233 & A232;
  assign \new_[42359]_  = A236 & ~A235;
  assign \new_[42360]_  = \new_[42359]_  & \new_[42356]_ ;
  assign \new_[42363]_  = A299 & A298;
  assign \new_[42366]_  = ~A302 & A301;
  assign \new_[42367]_  = \new_[42366]_  & \new_[42363]_ ;
  assign \new_[42368]_  = \new_[42367]_  & \new_[42360]_ ;
  assign \new_[42371]_  = A168 & A170;
  assign \new_[42374]_  = A166 & ~A167;
  assign \new_[42375]_  = \new_[42374]_  & \new_[42371]_ ;
  assign \new_[42378]_  = ~A200 & A199;
  assign \new_[42381]_  = A202 & ~A201;
  assign \new_[42382]_  = \new_[42381]_  & \new_[42378]_ ;
  assign \new_[42383]_  = \new_[42382]_  & \new_[42375]_ ;
  assign \new_[42386]_  = ~A233 & A232;
  assign \new_[42389]_  = A236 & ~A235;
  assign \new_[42390]_  = \new_[42389]_  & \new_[42386]_ ;
  assign \new_[42393]_  = ~A299 & A298;
  assign \new_[42396]_  = A302 & ~A301;
  assign \new_[42397]_  = \new_[42396]_  & \new_[42393]_ ;
  assign \new_[42398]_  = \new_[42397]_  & \new_[42390]_ ;
  assign \new_[42401]_  = A168 & A170;
  assign \new_[42404]_  = A166 & ~A167;
  assign \new_[42405]_  = \new_[42404]_  & \new_[42401]_ ;
  assign \new_[42408]_  = ~A200 & A199;
  assign \new_[42411]_  = A202 & ~A201;
  assign \new_[42412]_  = \new_[42411]_  & \new_[42408]_ ;
  assign \new_[42413]_  = \new_[42412]_  & \new_[42405]_ ;
  assign \new_[42416]_  = ~A233 & A232;
  assign \new_[42419]_  = A236 & ~A235;
  assign \new_[42420]_  = \new_[42419]_  & \new_[42416]_ ;
  assign \new_[42423]_  = A299 & ~A298;
  assign \new_[42426]_  = A302 & ~A301;
  assign \new_[42427]_  = \new_[42426]_  & \new_[42423]_ ;
  assign \new_[42428]_  = \new_[42427]_  & \new_[42420]_ ;
  assign \new_[42431]_  = A168 & A170;
  assign \new_[42434]_  = A166 & ~A167;
  assign \new_[42435]_  = \new_[42434]_  & \new_[42431]_ ;
  assign \new_[42438]_  = ~A200 & A199;
  assign \new_[42441]_  = A202 & ~A201;
  assign \new_[42442]_  = \new_[42441]_  & \new_[42438]_ ;
  assign \new_[42443]_  = \new_[42442]_  & \new_[42435]_ ;
  assign \new_[42446]_  = ~A233 & A232;
  assign \new_[42449]_  = A236 & ~A235;
  assign \new_[42450]_  = \new_[42449]_  & \new_[42446]_ ;
  assign \new_[42453]_  = ~A299 & ~A298;
  assign \new_[42456]_  = ~A302 & A301;
  assign \new_[42457]_  = \new_[42456]_  & \new_[42453]_ ;
  assign \new_[42458]_  = \new_[42457]_  & \new_[42450]_ ;
  assign \new_[42461]_  = A168 & A170;
  assign \new_[42464]_  = A166 & ~A167;
  assign \new_[42465]_  = \new_[42464]_  & \new_[42461]_ ;
  assign \new_[42468]_  = ~A200 & A199;
  assign \new_[42471]_  = A202 & ~A201;
  assign \new_[42472]_  = \new_[42471]_  & \new_[42468]_ ;
  assign \new_[42473]_  = \new_[42472]_  & \new_[42465]_ ;
  assign \new_[42476]_  = ~A233 & A232;
  assign \new_[42479]_  = A236 & ~A235;
  assign \new_[42480]_  = \new_[42479]_  & \new_[42476]_ ;
  assign \new_[42483]_  = A266 & A265;
  assign \new_[42486]_  = ~A269 & A268;
  assign \new_[42487]_  = \new_[42486]_  & \new_[42483]_ ;
  assign \new_[42488]_  = \new_[42487]_  & \new_[42480]_ ;
  assign \new_[42491]_  = A168 & A170;
  assign \new_[42494]_  = A166 & ~A167;
  assign \new_[42495]_  = \new_[42494]_  & \new_[42491]_ ;
  assign \new_[42498]_  = ~A200 & A199;
  assign \new_[42501]_  = A202 & ~A201;
  assign \new_[42502]_  = \new_[42501]_  & \new_[42498]_ ;
  assign \new_[42503]_  = \new_[42502]_  & \new_[42495]_ ;
  assign \new_[42506]_  = ~A233 & A232;
  assign \new_[42509]_  = A236 & ~A235;
  assign \new_[42510]_  = \new_[42509]_  & \new_[42506]_ ;
  assign \new_[42513]_  = A266 & ~A265;
  assign \new_[42516]_  = A269 & ~A268;
  assign \new_[42517]_  = \new_[42516]_  & \new_[42513]_ ;
  assign \new_[42518]_  = \new_[42517]_  & \new_[42510]_ ;
  assign \new_[42521]_  = A168 & A170;
  assign \new_[42524]_  = A166 & ~A167;
  assign \new_[42525]_  = \new_[42524]_  & \new_[42521]_ ;
  assign \new_[42528]_  = ~A200 & A199;
  assign \new_[42531]_  = A202 & ~A201;
  assign \new_[42532]_  = \new_[42531]_  & \new_[42528]_ ;
  assign \new_[42533]_  = \new_[42532]_  & \new_[42525]_ ;
  assign \new_[42536]_  = ~A233 & A232;
  assign \new_[42539]_  = A236 & ~A235;
  assign \new_[42540]_  = \new_[42539]_  & \new_[42536]_ ;
  assign \new_[42543]_  = ~A266 & A265;
  assign \new_[42546]_  = A269 & ~A268;
  assign \new_[42547]_  = \new_[42546]_  & \new_[42543]_ ;
  assign \new_[42548]_  = \new_[42547]_  & \new_[42540]_ ;
  assign \new_[42551]_  = A168 & A170;
  assign \new_[42554]_  = A166 & ~A167;
  assign \new_[42555]_  = \new_[42554]_  & \new_[42551]_ ;
  assign \new_[42558]_  = ~A200 & A199;
  assign \new_[42561]_  = A202 & ~A201;
  assign \new_[42562]_  = \new_[42561]_  & \new_[42558]_ ;
  assign \new_[42563]_  = \new_[42562]_  & \new_[42555]_ ;
  assign \new_[42566]_  = ~A233 & A232;
  assign \new_[42569]_  = A236 & ~A235;
  assign \new_[42570]_  = \new_[42569]_  & \new_[42566]_ ;
  assign \new_[42573]_  = ~A266 & ~A265;
  assign \new_[42576]_  = ~A269 & A268;
  assign \new_[42577]_  = \new_[42576]_  & \new_[42573]_ ;
  assign \new_[42578]_  = \new_[42577]_  & \new_[42570]_ ;
  assign \new_[42581]_  = A168 & A170;
  assign \new_[42584]_  = A166 & ~A167;
  assign \new_[42585]_  = \new_[42584]_  & \new_[42581]_ ;
  assign \new_[42588]_  = ~A200 & A199;
  assign \new_[42591]_  = A202 & ~A201;
  assign \new_[42592]_  = \new_[42591]_  & \new_[42588]_ ;
  assign \new_[42593]_  = \new_[42592]_  & \new_[42585]_ ;
  assign \new_[42596]_  = ~A233 & ~A232;
  assign \new_[42599]_  = ~A236 & A235;
  assign \new_[42600]_  = \new_[42599]_  & \new_[42596]_ ;
  assign \new_[42603]_  = A299 & A298;
  assign \new_[42606]_  = ~A302 & A301;
  assign \new_[42607]_  = \new_[42606]_  & \new_[42603]_ ;
  assign \new_[42608]_  = \new_[42607]_  & \new_[42600]_ ;
  assign \new_[42611]_  = A168 & A170;
  assign \new_[42614]_  = A166 & ~A167;
  assign \new_[42615]_  = \new_[42614]_  & \new_[42611]_ ;
  assign \new_[42618]_  = ~A200 & A199;
  assign \new_[42621]_  = A202 & ~A201;
  assign \new_[42622]_  = \new_[42621]_  & \new_[42618]_ ;
  assign \new_[42623]_  = \new_[42622]_  & \new_[42615]_ ;
  assign \new_[42626]_  = ~A233 & ~A232;
  assign \new_[42629]_  = ~A236 & A235;
  assign \new_[42630]_  = \new_[42629]_  & \new_[42626]_ ;
  assign \new_[42633]_  = ~A299 & A298;
  assign \new_[42636]_  = A302 & ~A301;
  assign \new_[42637]_  = \new_[42636]_  & \new_[42633]_ ;
  assign \new_[42638]_  = \new_[42637]_  & \new_[42630]_ ;
  assign \new_[42641]_  = A168 & A170;
  assign \new_[42644]_  = A166 & ~A167;
  assign \new_[42645]_  = \new_[42644]_  & \new_[42641]_ ;
  assign \new_[42648]_  = ~A200 & A199;
  assign \new_[42651]_  = A202 & ~A201;
  assign \new_[42652]_  = \new_[42651]_  & \new_[42648]_ ;
  assign \new_[42653]_  = \new_[42652]_  & \new_[42645]_ ;
  assign \new_[42656]_  = ~A233 & ~A232;
  assign \new_[42659]_  = ~A236 & A235;
  assign \new_[42660]_  = \new_[42659]_  & \new_[42656]_ ;
  assign \new_[42663]_  = A299 & ~A298;
  assign \new_[42666]_  = A302 & ~A301;
  assign \new_[42667]_  = \new_[42666]_  & \new_[42663]_ ;
  assign \new_[42668]_  = \new_[42667]_  & \new_[42660]_ ;
  assign \new_[42671]_  = A168 & A170;
  assign \new_[42674]_  = A166 & ~A167;
  assign \new_[42675]_  = \new_[42674]_  & \new_[42671]_ ;
  assign \new_[42678]_  = ~A200 & A199;
  assign \new_[42681]_  = A202 & ~A201;
  assign \new_[42682]_  = \new_[42681]_  & \new_[42678]_ ;
  assign \new_[42683]_  = \new_[42682]_  & \new_[42675]_ ;
  assign \new_[42686]_  = ~A233 & ~A232;
  assign \new_[42689]_  = ~A236 & A235;
  assign \new_[42690]_  = \new_[42689]_  & \new_[42686]_ ;
  assign \new_[42693]_  = ~A299 & ~A298;
  assign \new_[42696]_  = ~A302 & A301;
  assign \new_[42697]_  = \new_[42696]_  & \new_[42693]_ ;
  assign \new_[42698]_  = \new_[42697]_  & \new_[42690]_ ;
  assign \new_[42701]_  = A168 & A170;
  assign \new_[42704]_  = A166 & ~A167;
  assign \new_[42705]_  = \new_[42704]_  & \new_[42701]_ ;
  assign \new_[42708]_  = ~A200 & A199;
  assign \new_[42711]_  = A202 & ~A201;
  assign \new_[42712]_  = \new_[42711]_  & \new_[42708]_ ;
  assign \new_[42713]_  = \new_[42712]_  & \new_[42705]_ ;
  assign \new_[42716]_  = ~A233 & ~A232;
  assign \new_[42719]_  = ~A236 & A235;
  assign \new_[42720]_  = \new_[42719]_  & \new_[42716]_ ;
  assign \new_[42723]_  = A266 & A265;
  assign \new_[42726]_  = ~A269 & A268;
  assign \new_[42727]_  = \new_[42726]_  & \new_[42723]_ ;
  assign \new_[42728]_  = \new_[42727]_  & \new_[42720]_ ;
  assign \new_[42731]_  = A168 & A170;
  assign \new_[42734]_  = A166 & ~A167;
  assign \new_[42735]_  = \new_[42734]_  & \new_[42731]_ ;
  assign \new_[42738]_  = ~A200 & A199;
  assign \new_[42741]_  = A202 & ~A201;
  assign \new_[42742]_  = \new_[42741]_  & \new_[42738]_ ;
  assign \new_[42743]_  = \new_[42742]_  & \new_[42735]_ ;
  assign \new_[42746]_  = ~A233 & ~A232;
  assign \new_[42749]_  = ~A236 & A235;
  assign \new_[42750]_  = \new_[42749]_  & \new_[42746]_ ;
  assign \new_[42753]_  = A266 & ~A265;
  assign \new_[42756]_  = A269 & ~A268;
  assign \new_[42757]_  = \new_[42756]_  & \new_[42753]_ ;
  assign \new_[42758]_  = \new_[42757]_  & \new_[42750]_ ;
  assign \new_[42761]_  = A168 & A170;
  assign \new_[42764]_  = A166 & ~A167;
  assign \new_[42765]_  = \new_[42764]_  & \new_[42761]_ ;
  assign \new_[42768]_  = ~A200 & A199;
  assign \new_[42771]_  = A202 & ~A201;
  assign \new_[42772]_  = \new_[42771]_  & \new_[42768]_ ;
  assign \new_[42773]_  = \new_[42772]_  & \new_[42765]_ ;
  assign \new_[42776]_  = ~A233 & ~A232;
  assign \new_[42779]_  = ~A236 & A235;
  assign \new_[42780]_  = \new_[42779]_  & \new_[42776]_ ;
  assign \new_[42783]_  = ~A266 & A265;
  assign \new_[42786]_  = A269 & ~A268;
  assign \new_[42787]_  = \new_[42786]_  & \new_[42783]_ ;
  assign \new_[42788]_  = \new_[42787]_  & \new_[42780]_ ;
  assign \new_[42791]_  = A168 & A170;
  assign \new_[42794]_  = A166 & ~A167;
  assign \new_[42795]_  = \new_[42794]_  & \new_[42791]_ ;
  assign \new_[42798]_  = ~A200 & A199;
  assign \new_[42801]_  = A202 & ~A201;
  assign \new_[42802]_  = \new_[42801]_  & \new_[42798]_ ;
  assign \new_[42803]_  = \new_[42802]_  & \new_[42795]_ ;
  assign \new_[42806]_  = ~A233 & ~A232;
  assign \new_[42809]_  = ~A236 & A235;
  assign \new_[42810]_  = \new_[42809]_  & \new_[42806]_ ;
  assign \new_[42813]_  = ~A266 & ~A265;
  assign \new_[42816]_  = ~A269 & A268;
  assign \new_[42817]_  = \new_[42816]_  & \new_[42813]_ ;
  assign \new_[42818]_  = \new_[42817]_  & \new_[42810]_ ;
  assign \new_[42821]_  = A168 & A170;
  assign \new_[42824]_  = A166 & ~A167;
  assign \new_[42825]_  = \new_[42824]_  & \new_[42821]_ ;
  assign \new_[42828]_  = ~A200 & A199;
  assign \new_[42831]_  = ~A203 & ~A201;
  assign \new_[42832]_  = \new_[42831]_  & \new_[42828]_ ;
  assign \new_[42833]_  = \new_[42832]_  & \new_[42825]_ ;
  assign \new_[42836]_  = A233 & A232;
  assign \new_[42839]_  = ~A236 & A235;
  assign \new_[42840]_  = \new_[42839]_  & \new_[42836]_ ;
  assign \new_[42843]_  = A299 & A298;
  assign \new_[42846]_  = ~A302 & A301;
  assign \new_[42847]_  = \new_[42846]_  & \new_[42843]_ ;
  assign \new_[42848]_  = \new_[42847]_  & \new_[42840]_ ;
  assign \new_[42851]_  = A168 & A170;
  assign \new_[42854]_  = A166 & ~A167;
  assign \new_[42855]_  = \new_[42854]_  & \new_[42851]_ ;
  assign \new_[42858]_  = ~A200 & A199;
  assign \new_[42861]_  = ~A203 & ~A201;
  assign \new_[42862]_  = \new_[42861]_  & \new_[42858]_ ;
  assign \new_[42863]_  = \new_[42862]_  & \new_[42855]_ ;
  assign \new_[42866]_  = A233 & A232;
  assign \new_[42869]_  = ~A236 & A235;
  assign \new_[42870]_  = \new_[42869]_  & \new_[42866]_ ;
  assign \new_[42873]_  = ~A299 & A298;
  assign \new_[42876]_  = A302 & ~A301;
  assign \new_[42877]_  = \new_[42876]_  & \new_[42873]_ ;
  assign \new_[42878]_  = \new_[42877]_  & \new_[42870]_ ;
  assign \new_[42881]_  = A168 & A170;
  assign \new_[42884]_  = A166 & ~A167;
  assign \new_[42885]_  = \new_[42884]_  & \new_[42881]_ ;
  assign \new_[42888]_  = ~A200 & A199;
  assign \new_[42891]_  = ~A203 & ~A201;
  assign \new_[42892]_  = \new_[42891]_  & \new_[42888]_ ;
  assign \new_[42893]_  = \new_[42892]_  & \new_[42885]_ ;
  assign \new_[42896]_  = A233 & A232;
  assign \new_[42899]_  = ~A236 & A235;
  assign \new_[42900]_  = \new_[42899]_  & \new_[42896]_ ;
  assign \new_[42903]_  = A299 & ~A298;
  assign \new_[42906]_  = A302 & ~A301;
  assign \new_[42907]_  = \new_[42906]_  & \new_[42903]_ ;
  assign \new_[42908]_  = \new_[42907]_  & \new_[42900]_ ;
  assign \new_[42911]_  = A168 & A170;
  assign \new_[42914]_  = A166 & ~A167;
  assign \new_[42915]_  = \new_[42914]_  & \new_[42911]_ ;
  assign \new_[42918]_  = ~A200 & A199;
  assign \new_[42921]_  = ~A203 & ~A201;
  assign \new_[42922]_  = \new_[42921]_  & \new_[42918]_ ;
  assign \new_[42923]_  = \new_[42922]_  & \new_[42915]_ ;
  assign \new_[42926]_  = A233 & A232;
  assign \new_[42929]_  = ~A236 & A235;
  assign \new_[42930]_  = \new_[42929]_  & \new_[42926]_ ;
  assign \new_[42933]_  = ~A299 & ~A298;
  assign \new_[42936]_  = ~A302 & A301;
  assign \new_[42937]_  = \new_[42936]_  & \new_[42933]_ ;
  assign \new_[42938]_  = \new_[42937]_  & \new_[42930]_ ;
  assign \new_[42941]_  = A168 & A170;
  assign \new_[42944]_  = A166 & ~A167;
  assign \new_[42945]_  = \new_[42944]_  & \new_[42941]_ ;
  assign \new_[42948]_  = ~A200 & A199;
  assign \new_[42951]_  = ~A203 & ~A201;
  assign \new_[42952]_  = \new_[42951]_  & \new_[42948]_ ;
  assign \new_[42953]_  = \new_[42952]_  & \new_[42945]_ ;
  assign \new_[42956]_  = A233 & A232;
  assign \new_[42959]_  = ~A236 & A235;
  assign \new_[42960]_  = \new_[42959]_  & \new_[42956]_ ;
  assign \new_[42963]_  = A266 & A265;
  assign \new_[42966]_  = ~A269 & A268;
  assign \new_[42967]_  = \new_[42966]_  & \new_[42963]_ ;
  assign \new_[42968]_  = \new_[42967]_  & \new_[42960]_ ;
  assign \new_[42971]_  = A168 & A170;
  assign \new_[42974]_  = A166 & ~A167;
  assign \new_[42975]_  = \new_[42974]_  & \new_[42971]_ ;
  assign \new_[42978]_  = ~A200 & A199;
  assign \new_[42981]_  = ~A203 & ~A201;
  assign \new_[42982]_  = \new_[42981]_  & \new_[42978]_ ;
  assign \new_[42983]_  = \new_[42982]_  & \new_[42975]_ ;
  assign \new_[42986]_  = A233 & A232;
  assign \new_[42989]_  = ~A236 & A235;
  assign \new_[42990]_  = \new_[42989]_  & \new_[42986]_ ;
  assign \new_[42993]_  = A266 & ~A265;
  assign \new_[42996]_  = A269 & ~A268;
  assign \new_[42997]_  = \new_[42996]_  & \new_[42993]_ ;
  assign \new_[42998]_  = \new_[42997]_  & \new_[42990]_ ;
  assign \new_[43001]_  = A168 & A170;
  assign \new_[43004]_  = A166 & ~A167;
  assign \new_[43005]_  = \new_[43004]_  & \new_[43001]_ ;
  assign \new_[43008]_  = ~A200 & A199;
  assign \new_[43011]_  = ~A203 & ~A201;
  assign \new_[43012]_  = \new_[43011]_  & \new_[43008]_ ;
  assign \new_[43013]_  = \new_[43012]_  & \new_[43005]_ ;
  assign \new_[43016]_  = A233 & A232;
  assign \new_[43019]_  = ~A236 & A235;
  assign \new_[43020]_  = \new_[43019]_  & \new_[43016]_ ;
  assign \new_[43023]_  = ~A266 & A265;
  assign \new_[43026]_  = A269 & ~A268;
  assign \new_[43027]_  = \new_[43026]_  & \new_[43023]_ ;
  assign \new_[43028]_  = \new_[43027]_  & \new_[43020]_ ;
  assign \new_[43031]_  = A168 & A170;
  assign \new_[43034]_  = A166 & ~A167;
  assign \new_[43035]_  = \new_[43034]_  & \new_[43031]_ ;
  assign \new_[43038]_  = ~A200 & A199;
  assign \new_[43041]_  = ~A203 & ~A201;
  assign \new_[43042]_  = \new_[43041]_  & \new_[43038]_ ;
  assign \new_[43043]_  = \new_[43042]_  & \new_[43035]_ ;
  assign \new_[43046]_  = A233 & A232;
  assign \new_[43049]_  = ~A236 & A235;
  assign \new_[43050]_  = \new_[43049]_  & \new_[43046]_ ;
  assign \new_[43053]_  = ~A266 & ~A265;
  assign \new_[43056]_  = ~A269 & A268;
  assign \new_[43057]_  = \new_[43056]_  & \new_[43053]_ ;
  assign \new_[43058]_  = \new_[43057]_  & \new_[43050]_ ;
  assign \new_[43061]_  = A168 & A170;
  assign \new_[43064]_  = A166 & ~A167;
  assign \new_[43065]_  = \new_[43064]_  & \new_[43061]_ ;
  assign \new_[43068]_  = ~A200 & A199;
  assign \new_[43071]_  = ~A203 & ~A201;
  assign \new_[43072]_  = \new_[43071]_  & \new_[43068]_ ;
  assign \new_[43073]_  = \new_[43072]_  & \new_[43065]_ ;
  assign \new_[43076]_  = A233 & ~A232;
  assign \new_[43079]_  = A236 & ~A235;
  assign \new_[43080]_  = \new_[43079]_  & \new_[43076]_ ;
  assign \new_[43083]_  = A299 & A298;
  assign \new_[43086]_  = ~A302 & A301;
  assign \new_[43087]_  = \new_[43086]_  & \new_[43083]_ ;
  assign \new_[43088]_  = \new_[43087]_  & \new_[43080]_ ;
  assign \new_[43091]_  = A168 & A170;
  assign \new_[43094]_  = A166 & ~A167;
  assign \new_[43095]_  = \new_[43094]_  & \new_[43091]_ ;
  assign \new_[43098]_  = ~A200 & A199;
  assign \new_[43101]_  = ~A203 & ~A201;
  assign \new_[43102]_  = \new_[43101]_  & \new_[43098]_ ;
  assign \new_[43103]_  = \new_[43102]_  & \new_[43095]_ ;
  assign \new_[43106]_  = A233 & ~A232;
  assign \new_[43109]_  = A236 & ~A235;
  assign \new_[43110]_  = \new_[43109]_  & \new_[43106]_ ;
  assign \new_[43113]_  = ~A299 & A298;
  assign \new_[43116]_  = A302 & ~A301;
  assign \new_[43117]_  = \new_[43116]_  & \new_[43113]_ ;
  assign \new_[43118]_  = \new_[43117]_  & \new_[43110]_ ;
  assign \new_[43121]_  = A168 & A170;
  assign \new_[43124]_  = A166 & ~A167;
  assign \new_[43125]_  = \new_[43124]_  & \new_[43121]_ ;
  assign \new_[43128]_  = ~A200 & A199;
  assign \new_[43131]_  = ~A203 & ~A201;
  assign \new_[43132]_  = \new_[43131]_  & \new_[43128]_ ;
  assign \new_[43133]_  = \new_[43132]_  & \new_[43125]_ ;
  assign \new_[43136]_  = A233 & ~A232;
  assign \new_[43139]_  = A236 & ~A235;
  assign \new_[43140]_  = \new_[43139]_  & \new_[43136]_ ;
  assign \new_[43143]_  = A299 & ~A298;
  assign \new_[43146]_  = A302 & ~A301;
  assign \new_[43147]_  = \new_[43146]_  & \new_[43143]_ ;
  assign \new_[43148]_  = \new_[43147]_  & \new_[43140]_ ;
  assign \new_[43151]_  = A168 & A170;
  assign \new_[43154]_  = A166 & ~A167;
  assign \new_[43155]_  = \new_[43154]_  & \new_[43151]_ ;
  assign \new_[43158]_  = ~A200 & A199;
  assign \new_[43161]_  = ~A203 & ~A201;
  assign \new_[43162]_  = \new_[43161]_  & \new_[43158]_ ;
  assign \new_[43163]_  = \new_[43162]_  & \new_[43155]_ ;
  assign \new_[43166]_  = A233 & ~A232;
  assign \new_[43169]_  = A236 & ~A235;
  assign \new_[43170]_  = \new_[43169]_  & \new_[43166]_ ;
  assign \new_[43173]_  = ~A299 & ~A298;
  assign \new_[43176]_  = ~A302 & A301;
  assign \new_[43177]_  = \new_[43176]_  & \new_[43173]_ ;
  assign \new_[43178]_  = \new_[43177]_  & \new_[43170]_ ;
  assign \new_[43181]_  = A168 & A170;
  assign \new_[43184]_  = A166 & ~A167;
  assign \new_[43185]_  = \new_[43184]_  & \new_[43181]_ ;
  assign \new_[43188]_  = ~A200 & A199;
  assign \new_[43191]_  = ~A203 & ~A201;
  assign \new_[43192]_  = \new_[43191]_  & \new_[43188]_ ;
  assign \new_[43193]_  = \new_[43192]_  & \new_[43185]_ ;
  assign \new_[43196]_  = A233 & ~A232;
  assign \new_[43199]_  = A236 & ~A235;
  assign \new_[43200]_  = \new_[43199]_  & \new_[43196]_ ;
  assign \new_[43203]_  = A266 & A265;
  assign \new_[43206]_  = ~A269 & A268;
  assign \new_[43207]_  = \new_[43206]_  & \new_[43203]_ ;
  assign \new_[43208]_  = \new_[43207]_  & \new_[43200]_ ;
  assign \new_[43211]_  = A168 & A170;
  assign \new_[43214]_  = A166 & ~A167;
  assign \new_[43215]_  = \new_[43214]_  & \new_[43211]_ ;
  assign \new_[43218]_  = ~A200 & A199;
  assign \new_[43221]_  = ~A203 & ~A201;
  assign \new_[43222]_  = \new_[43221]_  & \new_[43218]_ ;
  assign \new_[43223]_  = \new_[43222]_  & \new_[43215]_ ;
  assign \new_[43226]_  = A233 & ~A232;
  assign \new_[43229]_  = A236 & ~A235;
  assign \new_[43230]_  = \new_[43229]_  & \new_[43226]_ ;
  assign \new_[43233]_  = A266 & ~A265;
  assign \new_[43236]_  = A269 & ~A268;
  assign \new_[43237]_  = \new_[43236]_  & \new_[43233]_ ;
  assign \new_[43238]_  = \new_[43237]_  & \new_[43230]_ ;
  assign \new_[43241]_  = A168 & A170;
  assign \new_[43244]_  = A166 & ~A167;
  assign \new_[43245]_  = \new_[43244]_  & \new_[43241]_ ;
  assign \new_[43248]_  = ~A200 & A199;
  assign \new_[43251]_  = ~A203 & ~A201;
  assign \new_[43252]_  = \new_[43251]_  & \new_[43248]_ ;
  assign \new_[43253]_  = \new_[43252]_  & \new_[43245]_ ;
  assign \new_[43256]_  = A233 & ~A232;
  assign \new_[43259]_  = A236 & ~A235;
  assign \new_[43260]_  = \new_[43259]_  & \new_[43256]_ ;
  assign \new_[43263]_  = ~A266 & A265;
  assign \new_[43266]_  = A269 & ~A268;
  assign \new_[43267]_  = \new_[43266]_  & \new_[43263]_ ;
  assign \new_[43268]_  = \new_[43267]_  & \new_[43260]_ ;
  assign \new_[43271]_  = A168 & A170;
  assign \new_[43274]_  = A166 & ~A167;
  assign \new_[43275]_  = \new_[43274]_  & \new_[43271]_ ;
  assign \new_[43278]_  = ~A200 & A199;
  assign \new_[43281]_  = ~A203 & ~A201;
  assign \new_[43282]_  = \new_[43281]_  & \new_[43278]_ ;
  assign \new_[43283]_  = \new_[43282]_  & \new_[43275]_ ;
  assign \new_[43286]_  = A233 & ~A232;
  assign \new_[43289]_  = A236 & ~A235;
  assign \new_[43290]_  = \new_[43289]_  & \new_[43286]_ ;
  assign \new_[43293]_  = ~A266 & ~A265;
  assign \new_[43296]_  = ~A269 & A268;
  assign \new_[43297]_  = \new_[43296]_  & \new_[43293]_ ;
  assign \new_[43298]_  = \new_[43297]_  & \new_[43290]_ ;
  assign \new_[43301]_  = A168 & A170;
  assign \new_[43304]_  = A166 & ~A167;
  assign \new_[43305]_  = \new_[43304]_  & \new_[43301]_ ;
  assign \new_[43308]_  = ~A200 & A199;
  assign \new_[43311]_  = ~A203 & ~A201;
  assign \new_[43312]_  = \new_[43311]_  & \new_[43308]_ ;
  assign \new_[43313]_  = \new_[43312]_  & \new_[43305]_ ;
  assign \new_[43316]_  = ~A233 & A232;
  assign \new_[43319]_  = A236 & ~A235;
  assign \new_[43320]_  = \new_[43319]_  & \new_[43316]_ ;
  assign \new_[43323]_  = A299 & A298;
  assign \new_[43326]_  = ~A302 & A301;
  assign \new_[43327]_  = \new_[43326]_  & \new_[43323]_ ;
  assign \new_[43328]_  = \new_[43327]_  & \new_[43320]_ ;
  assign \new_[43331]_  = A168 & A170;
  assign \new_[43334]_  = A166 & ~A167;
  assign \new_[43335]_  = \new_[43334]_  & \new_[43331]_ ;
  assign \new_[43338]_  = ~A200 & A199;
  assign \new_[43341]_  = ~A203 & ~A201;
  assign \new_[43342]_  = \new_[43341]_  & \new_[43338]_ ;
  assign \new_[43343]_  = \new_[43342]_  & \new_[43335]_ ;
  assign \new_[43346]_  = ~A233 & A232;
  assign \new_[43349]_  = A236 & ~A235;
  assign \new_[43350]_  = \new_[43349]_  & \new_[43346]_ ;
  assign \new_[43353]_  = ~A299 & A298;
  assign \new_[43356]_  = A302 & ~A301;
  assign \new_[43357]_  = \new_[43356]_  & \new_[43353]_ ;
  assign \new_[43358]_  = \new_[43357]_  & \new_[43350]_ ;
  assign \new_[43361]_  = A168 & A170;
  assign \new_[43364]_  = A166 & ~A167;
  assign \new_[43365]_  = \new_[43364]_  & \new_[43361]_ ;
  assign \new_[43368]_  = ~A200 & A199;
  assign \new_[43371]_  = ~A203 & ~A201;
  assign \new_[43372]_  = \new_[43371]_  & \new_[43368]_ ;
  assign \new_[43373]_  = \new_[43372]_  & \new_[43365]_ ;
  assign \new_[43376]_  = ~A233 & A232;
  assign \new_[43379]_  = A236 & ~A235;
  assign \new_[43380]_  = \new_[43379]_  & \new_[43376]_ ;
  assign \new_[43383]_  = A299 & ~A298;
  assign \new_[43386]_  = A302 & ~A301;
  assign \new_[43387]_  = \new_[43386]_  & \new_[43383]_ ;
  assign \new_[43388]_  = \new_[43387]_  & \new_[43380]_ ;
  assign \new_[43391]_  = A168 & A170;
  assign \new_[43394]_  = A166 & ~A167;
  assign \new_[43395]_  = \new_[43394]_  & \new_[43391]_ ;
  assign \new_[43398]_  = ~A200 & A199;
  assign \new_[43401]_  = ~A203 & ~A201;
  assign \new_[43402]_  = \new_[43401]_  & \new_[43398]_ ;
  assign \new_[43403]_  = \new_[43402]_  & \new_[43395]_ ;
  assign \new_[43406]_  = ~A233 & A232;
  assign \new_[43409]_  = A236 & ~A235;
  assign \new_[43410]_  = \new_[43409]_  & \new_[43406]_ ;
  assign \new_[43413]_  = ~A299 & ~A298;
  assign \new_[43416]_  = ~A302 & A301;
  assign \new_[43417]_  = \new_[43416]_  & \new_[43413]_ ;
  assign \new_[43418]_  = \new_[43417]_  & \new_[43410]_ ;
  assign \new_[43421]_  = A168 & A170;
  assign \new_[43424]_  = A166 & ~A167;
  assign \new_[43425]_  = \new_[43424]_  & \new_[43421]_ ;
  assign \new_[43428]_  = ~A200 & A199;
  assign \new_[43431]_  = ~A203 & ~A201;
  assign \new_[43432]_  = \new_[43431]_  & \new_[43428]_ ;
  assign \new_[43433]_  = \new_[43432]_  & \new_[43425]_ ;
  assign \new_[43436]_  = ~A233 & A232;
  assign \new_[43439]_  = A236 & ~A235;
  assign \new_[43440]_  = \new_[43439]_  & \new_[43436]_ ;
  assign \new_[43443]_  = A266 & A265;
  assign \new_[43446]_  = ~A269 & A268;
  assign \new_[43447]_  = \new_[43446]_  & \new_[43443]_ ;
  assign \new_[43448]_  = \new_[43447]_  & \new_[43440]_ ;
  assign \new_[43451]_  = A168 & A170;
  assign \new_[43454]_  = A166 & ~A167;
  assign \new_[43455]_  = \new_[43454]_  & \new_[43451]_ ;
  assign \new_[43458]_  = ~A200 & A199;
  assign \new_[43461]_  = ~A203 & ~A201;
  assign \new_[43462]_  = \new_[43461]_  & \new_[43458]_ ;
  assign \new_[43463]_  = \new_[43462]_  & \new_[43455]_ ;
  assign \new_[43466]_  = ~A233 & A232;
  assign \new_[43469]_  = A236 & ~A235;
  assign \new_[43470]_  = \new_[43469]_  & \new_[43466]_ ;
  assign \new_[43473]_  = A266 & ~A265;
  assign \new_[43476]_  = A269 & ~A268;
  assign \new_[43477]_  = \new_[43476]_  & \new_[43473]_ ;
  assign \new_[43478]_  = \new_[43477]_  & \new_[43470]_ ;
  assign \new_[43481]_  = A168 & A170;
  assign \new_[43484]_  = A166 & ~A167;
  assign \new_[43485]_  = \new_[43484]_  & \new_[43481]_ ;
  assign \new_[43488]_  = ~A200 & A199;
  assign \new_[43491]_  = ~A203 & ~A201;
  assign \new_[43492]_  = \new_[43491]_  & \new_[43488]_ ;
  assign \new_[43493]_  = \new_[43492]_  & \new_[43485]_ ;
  assign \new_[43496]_  = ~A233 & A232;
  assign \new_[43499]_  = A236 & ~A235;
  assign \new_[43500]_  = \new_[43499]_  & \new_[43496]_ ;
  assign \new_[43503]_  = ~A266 & A265;
  assign \new_[43506]_  = A269 & ~A268;
  assign \new_[43507]_  = \new_[43506]_  & \new_[43503]_ ;
  assign \new_[43508]_  = \new_[43507]_  & \new_[43500]_ ;
  assign \new_[43511]_  = A168 & A170;
  assign \new_[43514]_  = A166 & ~A167;
  assign \new_[43515]_  = \new_[43514]_  & \new_[43511]_ ;
  assign \new_[43518]_  = ~A200 & A199;
  assign \new_[43521]_  = ~A203 & ~A201;
  assign \new_[43522]_  = \new_[43521]_  & \new_[43518]_ ;
  assign \new_[43523]_  = \new_[43522]_  & \new_[43515]_ ;
  assign \new_[43526]_  = ~A233 & A232;
  assign \new_[43529]_  = A236 & ~A235;
  assign \new_[43530]_  = \new_[43529]_  & \new_[43526]_ ;
  assign \new_[43533]_  = ~A266 & ~A265;
  assign \new_[43536]_  = ~A269 & A268;
  assign \new_[43537]_  = \new_[43536]_  & \new_[43533]_ ;
  assign \new_[43538]_  = \new_[43537]_  & \new_[43530]_ ;
  assign \new_[43541]_  = A168 & A170;
  assign \new_[43544]_  = A166 & ~A167;
  assign \new_[43545]_  = \new_[43544]_  & \new_[43541]_ ;
  assign \new_[43548]_  = ~A200 & A199;
  assign \new_[43551]_  = ~A203 & ~A201;
  assign \new_[43552]_  = \new_[43551]_  & \new_[43548]_ ;
  assign \new_[43553]_  = \new_[43552]_  & \new_[43545]_ ;
  assign \new_[43556]_  = ~A233 & ~A232;
  assign \new_[43559]_  = ~A236 & A235;
  assign \new_[43560]_  = \new_[43559]_  & \new_[43556]_ ;
  assign \new_[43563]_  = A299 & A298;
  assign \new_[43566]_  = ~A302 & A301;
  assign \new_[43567]_  = \new_[43566]_  & \new_[43563]_ ;
  assign \new_[43568]_  = \new_[43567]_  & \new_[43560]_ ;
  assign \new_[43571]_  = A168 & A170;
  assign \new_[43574]_  = A166 & ~A167;
  assign \new_[43575]_  = \new_[43574]_  & \new_[43571]_ ;
  assign \new_[43578]_  = ~A200 & A199;
  assign \new_[43581]_  = ~A203 & ~A201;
  assign \new_[43582]_  = \new_[43581]_  & \new_[43578]_ ;
  assign \new_[43583]_  = \new_[43582]_  & \new_[43575]_ ;
  assign \new_[43586]_  = ~A233 & ~A232;
  assign \new_[43589]_  = ~A236 & A235;
  assign \new_[43590]_  = \new_[43589]_  & \new_[43586]_ ;
  assign \new_[43593]_  = ~A299 & A298;
  assign \new_[43596]_  = A302 & ~A301;
  assign \new_[43597]_  = \new_[43596]_  & \new_[43593]_ ;
  assign \new_[43598]_  = \new_[43597]_  & \new_[43590]_ ;
  assign \new_[43601]_  = A168 & A170;
  assign \new_[43604]_  = A166 & ~A167;
  assign \new_[43605]_  = \new_[43604]_  & \new_[43601]_ ;
  assign \new_[43608]_  = ~A200 & A199;
  assign \new_[43611]_  = ~A203 & ~A201;
  assign \new_[43612]_  = \new_[43611]_  & \new_[43608]_ ;
  assign \new_[43613]_  = \new_[43612]_  & \new_[43605]_ ;
  assign \new_[43616]_  = ~A233 & ~A232;
  assign \new_[43619]_  = ~A236 & A235;
  assign \new_[43620]_  = \new_[43619]_  & \new_[43616]_ ;
  assign \new_[43623]_  = A299 & ~A298;
  assign \new_[43626]_  = A302 & ~A301;
  assign \new_[43627]_  = \new_[43626]_  & \new_[43623]_ ;
  assign \new_[43628]_  = \new_[43627]_  & \new_[43620]_ ;
  assign \new_[43631]_  = A168 & A170;
  assign \new_[43634]_  = A166 & ~A167;
  assign \new_[43635]_  = \new_[43634]_  & \new_[43631]_ ;
  assign \new_[43638]_  = ~A200 & A199;
  assign \new_[43641]_  = ~A203 & ~A201;
  assign \new_[43642]_  = \new_[43641]_  & \new_[43638]_ ;
  assign \new_[43643]_  = \new_[43642]_  & \new_[43635]_ ;
  assign \new_[43646]_  = ~A233 & ~A232;
  assign \new_[43649]_  = ~A236 & A235;
  assign \new_[43650]_  = \new_[43649]_  & \new_[43646]_ ;
  assign \new_[43653]_  = ~A299 & ~A298;
  assign \new_[43656]_  = ~A302 & A301;
  assign \new_[43657]_  = \new_[43656]_  & \new_[43653]_ ;
  assign \new_[43658]_  = \new_[43657]_  & \new_[43650]_ ;
  assign \new_[43661]_  = A168 & A170;
  assign \new_[43664]_  = A166 & ~A167;
  assign \new_[43665]_  = \new_[43664]_  & \new_[43661]_ ;
  assign \new_[43668]_  = ~A200 & A199;
  assign \new_[43671]_  = ~A203 & ~A201;
  assign \new_[43672]_  = \new_[43671]_  & \new_[43668]_ ;
  assign \new_[43673]_  = \new_[43672]_  & \new_[43665]_ ;
  assign \new_[43676]_  = ~A233 & ~A232;
  assign \new_[43679]_  = ~A236 & A235;
  assign \new_[43680]_  = \new_[43679]_  & \new_[43676]_ ;
  assign \new_[43683]_  = A266 & A265;
  assign \new_[43686]_  = ~A269 & A268;
  assign \new_[43687]_  = \new_[43686]_  & \new_[43683]_ ;
  assign \new_[43688]_  = \new_[43687]_  & \new_[43680]_ ;
  assign \new_[43691]_  = A168 & A170;
  assign \new_[43694]_  = A166 & ~A167;
  assign \new_[43695]_  = \new_[43694]_  & \new_[43691]_ ;
  assign \new_[43698]_  = ~A200 & A199;
  assign \new_[43701]_  = ~A203 & ~A201;
  assign \new_[43702]_  = \new_[43701]_  & \new_[43698]_ ;
  assign \new_[43703]_  = \new_[43702]_  & \new_[43695]_ ;
  assign \new_[43706]_  = ~A233 & ~A232;
  assign \new_[43709]_  = ~A236 & A235;
  assign \new_[43710]_  = \new_[43709]_  & \new_[43706]_ ;
  assign \new_[43713]_  = A266 & ~A265;
  assign \new_[43716]_  = A269 & ~A268;
  assign \new_[43717]_  = \new_[43716]_  & \new_[43713]_ ;
  assign \new_[43718]_  = \new_[43717]_  & \new_[43710]_ ;
  assign \new_[43721]_  = A168 & A170;
  assign \new_[43724]_  = A166 & ~A167;
  assign \new_[43725]_  = \new_[43724]_  & \new_[43721]_ ;
  assign \new_[43728]_  = ~A200 & A199;
  assign \new_[43731]_  = ~A203 & ~A201;
  assign \new_[43732]_  = \new_[43731]_  & \new_[43728]_ ;
  assign \new_[43733]_  = \new_[43732]_  & \new_[43725]_ ;
  assign \new_[43736]_  = ~A233 & ~A232;
  assign \new_[43739]_  = ~A236 & A235;
  assign \new_[43740]_  = \new_[43739]_  & \new_[43736]_ ;
  assign \new_[43743]_  = ~A266 & A265;
  assign \new_[43746]_  = A269 & ~A268;
  assign \new_[43747]_  = \new_[43746]_  & \new_[43743]_ ;
  assign \new_[43748]_  = \new_[43747]_  & \new_[43740]_ ;
  assign \new_[43751]_  = A168 & A170;
  assign \new_[43754]_  = A166 & ~A167;
  assign \new_[43755]_  = \new_[43754]_  & \new_[43751]_ ;
  assign \new_[43758]_  = ~A200 & A199;
  assign \new_[43761]_  = ~A203 & ~A201;
  assign \new_[43762]_  = \new_[43761]_  & \new_[43758]_ ;
  assign \new_[43763]_  = \new_[43762]_  & \new_[43755]_ ;
  assign \new_[43766]_  = ~A233 & ~A232;
  assign \new_[43769]_  = ~A236 & A235;
  assign \new_[43770]_  = \new_[43769]_  & \new_[43766]_ ;
  assign \new_[43773]_  = ~A266 & ~A265;
  assign \new_[43776]_  = ~A269 & A268;
  assign \new_[43777]_  = \new_[43776]_  & \new_[43773]_ ;
  assign \new_[43778]_  = \new_[43777]_  & \new_[43770]_ ;
  assign \new_[43781]_  = A168 & A169;
  assign \new_[43784]_  = A166 & ~A167;
  assign \new_[43785]_  = \new_[43784]_  & \new_[43781]_ ;
  assign \new_[43788]_  = A200 & A199;
  assign \new_[43791]_  = ~A202 & ~A201;
  assign \new_[43792]_  = \new_[43791]_  & \new_[43788]_ ;
  assign \new_[43793]_  = \new_[43792]_  & \new_[43785]_ ;
  assign \new_[43796]_  = A233 & A232;
  assign \new_[43799]_  = ~A236 & A235;
  assign \new_[43800]_  = \new_[43799]_  & \new_[43796]_ ;
  assign \new_[43803]_  = A299 & A298;
  assign \new_[43806]_  = ~A302 & A301;
  assign \new_[43807]_  = \new_[43806]_  & \new_[43803]_ ;
  assign \new_[43808]_  = \new_[43807]_  & \new_[43800]_ ;
  assign \new_[43811]_  = A168 & A169;
  assign \new_[43814]_  = A166 & ~A167;
  assign \new_[43815]_  = \new_[43814]_  & \new_[43811]_ ;
  assign \new_[43818]_  = A200 & A199;
  assign \new_[43821]_  = ~A202 & ~A201;
  assign \new_[43822]_  = \new_[43821]_  & \new_[43818]_ ;
  assign \new_[43823]_  = \new_[43822]_  & \new_[43815]_ ;
  assign \new_[43826]_  = A233 & A232;
  assign \new_[43829]_  = ~A236 & A235;
  assign \new_[43830]_  = \new_[43829]_  & \new_[43826]_ ;
  assign \new_[43833]_  = ~A299 & A298;
  assign \new_[43836]_  = A302 & ~A301;
  assign \new_[43837]_  = \new_[43836]_  & \new_[43833]_ ;
  assign \new_[43838]_  = \new_[43837]_  & \new_[43830]_ ;
  assign \new_[43841]_  = A168 & A169;
  assign \new_[43844]_  = A166 & ~A167;
  assign \new_[43845]_  = \new_[43844]_  & \new_[43841]_ ;
  assign \new_[43848]_  = A200 & A199;
  assign \new_[43851]_  = ~A202 & ~A201;
  assign \new_[43852]_  = \new_[43851]_  & \new_[43848]_ ;
  assign \new_[43853]_  = \new_[43852]_  & \new_[43845]_ ;
  assign \new_[43856]_  = A233 & A232;
  assign \new_[43859]_  = ~A236 & A235;
  assign \new_[43860]_  = \new_[43859]_  & \new_[43856]_ ;
  assign \new_[43863]_  = A299 & ~A298;
  assign \new_[43866]_  = A302 & ~A301;
  assign \new_[43867]_  = \new_[43866]_  & \new_[43863]_ ;
  assign \new_[43868]_  = \new_[43867]_  & \new_[43860]_ ;
  assign \new_[43871]_  = A168 & A169;
  assign \new_[43874]_  = A166 & ~A167;
  assign \new_[43875]_  = \new_[43874]_  & \new_[43871]_ ;
  assign \new_[43878]_  = A200 & A199;
  assign \new_[43881]_  = ~A202 & ~A201;
  assign \new_[43882]_  = \new_[43881]_  & \new_[43878]_ ;
  assign \new_[43883]_  = \new_[43882]_  & \new_[43875]_ ;
  assign \new_[43886]_  = A233 & A232;
  assign \new_[43889]_  = ~A236 & A235;
  assign \new_[43890]_  = \new_[43889]_  & \new_[43886]_ ;
  assign \new_[43893]_  = ~A299 & ~A298;
  assign \new_[43896]_  = ~A302 & A301;
  assign \new_[43897]_  = \new_[43896]_  & \new_[43893]_ ;
  assign \new_[43898]_  = \new_[43897]_  & \new_[43890]_ ;
  assign \new_[43901]_  = A168 & A169;
  assign \new_[43904]_  = A166 & ~A167;
  assign \new_[43905]_  = \new_[43904]_  & \new_[43901]_ ;
  assign \new_[43908]_  = A200 & A199;
  assign \new_[43911]_  = ~A202 & ~A201;
  assign \new_[43912]_  = \new_[43911]_  & \new_[43908]_ ;
  assign \new_[43913]_  = \new_[43912]_  & \new_[43905]_ ;
  assign \new_[43916]_  = A233 & A232;
  assign \new_[43919]_  = ~A236 & A235;
  assign \new_[43920]_  = \new_[43919]_  & \new_[43916]_ ;
  assign \new_[43923]_  = A266 & A265;
  assign \new_[43926]_  = ~A269 & A268;
  assign \new_[43927]_  = \new_[43926]_  & \new_[43923]_ ;
  assign \new_[43928]_  = \new_[43927]_  & \new_[43920]_ ;
  assign \new_[43931]_  = A168 & A169;
  assign \new_[43934]_  = A166 & ~A167;
  assign \new_[43935]_  = \new_[43934]_  & \new_[43931]_ ;
  assign \new_[43938]_  = A200 & A199;
  assign \new_[43941]_  = ~A202 & ~A201;
  assign \new_[43942]_  = \new_[43941]_  & \new_[43938]_ ;
  assign \new_[43943]_  = \new_[43942]_  & \new_[43935]_ ;
  assign \new_[43946]_  = A233 & A232;
  assign \new_[43949]_  = ~A236 & A235;
  assign \new_[43950]_  = \new_[43949]_  & \new_[43946]_ ;
  assign \new_[43953]_  = A266 & ~A265;
  assign \new_[43956]_  = A269 & ~A268;
  assign \new_[43957]_  = \new_[43956]_  & \new_[43953]_ ;
  assign \new_[43958]_  = \new_[43957]_  & \new_[43950]_ ;
  assign \new_[43961]_  = A168 & A169;
  assign \new_[43964]_  = A166 & ~A167;
  assign \new_[43965]_  = \new_[43964]_  & \new_[43961]_ ;
  assign \new_[43968]_  = A200 & A199;
  assign \new_[43971]_  = ~A202 & ~A201;
  assign \new_[43972]_  = \new_[43971]_  & \new_[43968]_ ;
  assign \new_[43973]_  = \new_[43972]_  & \new_[43965]_ ;
  assign \new_[43976]_  = A233 & A232;
  assign \new_[43979]_  = ~A236 & A235;
  assign \new_[43980]_  = \new_[43979]_  & \new_[43976]_ ;
  assign \new_[43983]_  = ~A266 & A265;
  assign \new_[43986]_  = A269 & ~A268;
  assign \new_[43987]_  = \new_[43986]_  & \new_[43983]_ ;
  assign \new_[43988]_  = \new_[43987]_  & \new_[43980]_ ;
  assign \new_[43991]_  = A168 & A169;
  assign \new_[43994]_  = A166 & ~A167;
  assign \new_[43995]_  = \new_[43994]_  & \new_[43991]_ ;
  assign \new_[43998]_  = A200 & A199;
  assign \new_[44001]_  = ~A202 & ~A201;
  assign \new_[44002]_  = \new_[44001]_  & \new_[43998]_ ;
  assign \new_[44003]_  = \new_[44002]_  & \new_[43995]_ ;
  assign \new_[44006]_  = A233 & A232;
  assign \new_[44009]_  = ~A236 & A235;
  assign \new_[44010]_  = \new_[44009]_  & \new_[44006]_ ;
  assign \new_[44013]_  = ~A266 & ~A265;
  assign \new_[44016]_  = ~A269 & A268;
  assign \new_[44017]_  = \new_[44016]_  & \new_[44013]_ ;
  assign \new_[44018]_  = \new_[44017]_  & \new_[44010]_ ;
  assign \new_[44021]_  = A168 & A169;
  assign \new_[44024]_  = A166 & ~A167;
  assign \new_[44025]_  = \new_[44024]_  & \new_[44021]_ ;
  assign \new_[44028]_  = A200 & A199;
  assign \new_[44031]_  = ~A202 & ~A201;
  assign \new_[44032]_  = \new_[44031]_  & \new_[44028]_ ;
  assign \new_[44033]_  = \new_[44032]_  & \new_[44025]_ ;
  assign \new_[44036]_  = A233 & ~A232;
  assign \new_[44039]_  = A236 & ~A235;
  assign \new_[44040]_  = \new_[44039]_  & \new_[44036]_ ;
  assign \new_[44043]_  = A299 & A298;
  assign \new_[44046]_  = ~A302 & A301;
  assign \new_[44047]_  = \new_[44046]_  & \new_[44043]_ ;
  assign \new_[44048]_  = \new_[44047]_  & \new_[44040]_ ;
  assign \new_[44051]_  = A168 & A169;
  assign \new_[44054]_  = A166 & ~A167;
  assign \new_[44055]_  = \new_[44054]_  & \new_[44051]_ ;
  assign \new_[44058]_  = A200 & A199;
  assign \new_[44061]_  = ~A202 & ~A201;
  assign \new_[44062]_  = \new_[44061]_  & \new_[44058]_ ;
  assign \new_[44063]_  = \new_[44062]_  & \new_[44055]_ ;
  assign \new_[44066]_  = A233 & ~A232;
  assign \new_[44069]_  = A236 & ~A235;
  assign \new_[44070]_  = \new_[44069]_  & \new_[44066]_ ;
  assign \new_[44073]_  = ~A299 & A298;
  assign \new_[44076]_  = A302 & ~A301;
  assign \new_[44077]_  = \new_[44076]_  & \new_[44073]_ ;
  assign \new_[44078]_  = \new_[44077]_  & \new_[44070]_ ;
  assign \new_[44081]_  = A168 & A169;
  assign \new_[44084]_  = A166 & ~A167;
  assign \new_[44085]_  = \new_[44084]_  & \new_[44081]_ ;
  assign \new_[44088]_  = A200 & A199;
  assign \new_[44091]_  = ~A202 & ~A201;
  assign \new_[44092]_  = \new_[44091]_  & \new_[44088]_ ;
  assign \new_[44093]_  = \new_[44092]_  & \new_[44085]_ ;
  assign \new_[44096]_  = A233 & ~A232;
  assign \new_[44099]_  = A236 & ~A235;
  assign \new_[44100]_  = \new_[44099]_  & \new_[44096]_ ;
  assign \new_[44103]_  = A299 & ~A298;
  assign \new_[44106]_  = A302 & ~A301;
  assign \new_[44107]_  = \new_[44106]_  & \new_[44103]_ ;
  assign \new_[44108]_  = \new_[44107]_  & \new_[44100]_ ;
  assign \new_[44111]_  = A168 & A169;
  assign \new_[44114]_  = A166 & ~A167;
  assign \new_[44115]_  = \new_[44114]_  & \new_[44111]_ ;
  assign \new_[44118]_  = A200 & A199;
  assign \new_[44121]_  = ~A202 & ~A201;
  assign \new_[44122]_  = \new_[44121]_  & \new_[44118]_ ;
  assign \new_[44123]_  = \new_[44122]_  & \new_[44115]_ ;
  assign \new_[44126]_  = A233 & ~A232;
  assign \new_[44129]_  = A236 & ~A235;
  assign \new_[44130]_  = \new_[44129]_  & \new_[44126]_ ;
  assign \new_[44133]_  = ~A299 & ~A298;
  assign \new_[44136]_  = ~A302 & A301;
  assign \new_[44137]_  = \new_[44136]_  & \new_[44133]_ ;
  assign \new_[44138]_  = \new_[44137]_  & \new_[44130]_ ;
  assign \new_[44141]_  = A168 & A169;
  assign \new_[44144]_  = A166 & ~A167;
  assign \new_[44145]_  = \new_[44144]_  & \new_[44141]_ ;
  assign \new_[44148]_  = A200 & A199;
  assign \new_[44151]_  = ~A202 & ~A201;
  assign \new_[44152]_  = \new_[44151]_  & \new_[44148]_ ;
  assign \new_[44153]_  = \new_[44152]_  & \new_[44145]_ ;
  assign \new_[44156]_  = A233 & ~A232;
  assign \new_[44159]_  = A236 & ~A235;
  assign \new_[44160]_  = \new_[44159]_  & \new_[44156]_ ;
  assign \new_[44163]_  = A266 & A265;
  assign \new_[44166]_  = ~A269 & A268;
  assign \new_[44167]_  = \new_[44166]_  & \new_[44163]_ ;
  assign \new_[44168]_  = \new_[44167]_  & \new_[44160]_ ;
  assign \new_[44171]_  = A168 & A169;
  assign \new_[44174]_  = A166 & ~A167;
  assign \new_[44175]_  = \new_[44174]_  & \new_[44171]_ ;
  assign \new_[44178]_  = A200 & A199;
  assign \new_[44181]_  = ~A202 & ~A201;
  assign \new_[44182]_  = \new_[44181]_  & \new_[44178]_ ;
  assign \new_[44183]_  = \new_[44182]_  & \new_[44175]_ ;
  assign \new_[44186]_  = A233 & ~A232;
  assign \new_[44189]_  = A236 & ~A235;
  assign \new_[44190]_  = \new_[44189]_  & \new_[44186]_ ;
  assign \new_[44193]_  = A266 & ~A265;
  assign \new_[44196]_  = A269 & ~A268;
  assign \new_[44197]_  = \new_[44196]_  & \new_[44193]_ ;
  assign \new_[44198]_  = \new_[44197]_  & \new_[44190]_ ;
  assign \new_[44201]_  = A168 & A169;
  assign \new_[44204]_  = A166 & ~A167;
  assign \new_[44205]_  = \new_[44204]_  & \new_[44201]_ ;
  assign \new_[44208]_  = A200 & A199;
  assign \new_[44211]_  = ~A202 & ~A201;
  assign \new_[44212]_  = \new_[44211]_  & \new_[44208]_ ;
  assign \new_[44213]_  = \new_[44212]_  & \new_[44205]_ ;
  assign \new_[44216]_  = A233 & ~A232;
  assign \new_[44219]_  = A236 & ~A235;
  assign \new_[44220]_  = \new_[44219]_  & \new_[44216]_ ;
  assign \new_[44223]_  = ~A266 & A265;
  assign \new_[44226]_  = A269 & ~A268;
  assign \new_[44227]_  = \new_[44226]_  & \new_[44223]_ ;
  assign \new_[44228]_  = \new_[44227]_  & \new_[44220]_ ;
  assign \new_[44231]_  = A168 & A169;
  assign \new_[44234]_  = A166 & ~A167;
  assign \new_[44235]_  = \new_[44234]_  & \new_[44231]_ ;
  assign \new_[44238]_  = A200 & A199;
  assign \new_[44241]_  = ~A202 & ~A201;
  assign \new_[44242]_  = \new_[44241]_  & \new_[44238]_ ;
  assign \new_[44243]_  = \new_[44242]_  & \new_[44235]_ ;
  assign \new_[44246]_  = A233 & ~A232;
  assign \new_[44249]_  = A236 & ~A235;
  assign \new_[44250]_  = \new_[44249]_  & \new_[44246]_ ;
  assign \new_[44253]_  = ~A266 & ~A265;
  assign \new_[44256]_  = ~A269 & A268;
  assign \new_[44257]_  = \new_[44256]_  & \new_[44253]_ ;
  assign \new_[44258]_  = \new_[44257]_  & \new_[44250]_ ;
  assign \new_[44261]_  = A168 & A169;
  assign \new_[44264]_  = A166 & ~A167;
  assign \new_[44265]_  = \new_[44264]_  & \new_[44261]_ ;
  assign \new_[44268]_  = A200 & A199;
  assign \new_[44271]_  = ~A202 & ~A201;
  assign \new_[44272]_  = \new_[44271]_  & \new_[44268]_ ;
  assign \new_[44273]_  = \new_[44272]_  & \new_[44265]_ ;
  assign \new_[44276]_  = ~A233 & A232;
  assign \new_[44279]_  = A236 & ~A235;
  assign \new_[44280]_  = \new_[44279]_  & \new_[44276]_ ;
  assign \new_[44283]_  = A299 & A298;
  assign \new_[44286]_  = ~A302 & A301;
  assign \new_[44287]_  = \new_[44286]_  & \new_[44283]_ ;
  assign \new_[44288]_  = \new_[44287]_  & \new_[44280]_ ;
  assign \new_[44291]_  = A168 & A169;
  assign \new_[44294]_  = A166 & ~A167;
  assign \new_[44295]_  = \new_[44294]_  & \new_[44291]_ ;
  assign \new_[44298]_  = A200 & A199;
  assign \new_[44301]_  = ~A202 & ~A201;
  assign \new_[44302]_  = \new_[44301]_  & \new_[44298]_ ;
  assign \new_[44303]_  = \new_[44302]_  & \new_[44295]_ ;
  assign \new_[44306]_  = ~A233 & A232;
  assign \new_[44309]_  = A236 & ~A235;
  assign \new_[44310]_  = \new_[44309]_  & \new_[44306]_ ;
  assign \new_[44313]_  = ~A299 & A298;
  assign \new_[44316]_  = A302 & ~A301;
  assign \new_[44317]_  = \new_[44316]_  & \new_[44313]_ ;
  assign \new_[44318]_  = \new_[44317]_  & \new_[44310]_ ;
  assign \new_[44321]_  = A168 & A169;
  assign \new_[44324]_  = A166 & ~A167;
  assign \new_[44325]_  = \new_[44324]_  & \new_[44321]_ ;
  assign \new_[44328]_  = A200 & A199;
  assign \new_[44331]_  = ~A202 & ~A201;
  assign \new_[44332]_  = \new_[44331]_  & \new_[44328]_ ;
  assign \new_[44333]_  = \new_[44332]_  & \new_[44325]_ ;
  assign \new_[44336]_  = ~A233 & A232;
  assign \new_[44339]_  = A236 & ~A235;
  assign \new_[44340]_  = \new_[44339]_  & \new_[44336]_ ;
  assign \new_[44343]_  = A299 & ~A298;
  assign \new_[44346]_  = A302 & ~A301;
  assign \new_[44347]_  = \new_[44346]_  & \new_[44343]_ ;
  assign \new_[44348]_  = \new_[44347]_  & \new_[44340]_ ;
  assign \new_[44351]_  = A168 & A169;
  assign \new_[44354]_  = A166 & ~A167;
  assign \new_[44355]_  = \new_[44354]_  & \new_[44351]_ ;
  assign \new_[44358]_  = A200 & A199;
  assign \new_[44361]_  = ~A202 & ~A201;
  assign \new_[44362]_  = \new_[44361]_  & \new_[44358]_ ;
  assign \new_[44363]_  = \new_[44362]_  & \new_[44355]_ ;
  assign \new_[44366]_  = ~A233 & A232;
  assign \new_[44369]_  = A236 & ~A235;
  assign \new_[44370]_  = \new_[44369]_  & \new_[44366]_ ;
  assign \new_[44373]_  = ~A299 & ~A298;
  assign \new_[44376]_  = ~A302 & A301;
  assign \new_[44377]_  = \new_[44376]_  & \new_[44373]_ ;
  assign \new_[44378]_  = \new_[44377]_  & \new_[44370]_ ;
  assign \new_[44381]_  = A168 & A169;
  assign \new_[44384]_  = A166 & ~A167;
  assign \new_[44385]_  = \new_[44384]_  & \new_[44381]_ ;
  assign \new_[44388]_  = A200 & A199;
  assign \new_[44391]_  = ~A202 & ~A201;
  assign \new_[44392]_  = \new_[44391]_  & \new_[44388]_ ;
  assign \new_[44393]_  = \new_[44392]_  & \new_[44385]_ ;
  assign \new_[44396]_  = ~A233 & A232;
  assign \new_[44399]_  = A236 & ~A235;
  assign \new_[44400]_  = \new_[44399]_  & \new_[44396]_ ;
  assign \new_[44403]_  = A266 & A265;
  assign \new_[44406]_  = ~A269 & A268;
  assign \new_[44407]_  = \new_[44406]_  & \new_[44403]_ ;
  assign \new_[44408]_  = \new_[44407]_  & \new_[44400]_ ;
  assign \new_[44411]_  = A168 & A169;
  assign \new_[44414]_  = A166 & ~A167;
  assign \new_[44415]_  = \new_[44414]_  & \new_[44411]_ ;
  assign \new_[44418]_  = A200 & A199;
  assign \new_[44421]_  = ~A202 & ~A201;
  assign \new_[44422]_  = \new_[44421]_  & \new_[44418]_ ;
  assign \new_[44423]_  = \new_[44422]_  & \new_[44415]_ ;
  assign \new_[44426]_  = ~A233 & A232;
  assign \new_[44429]_  = A236 & ~A235;
  assign \new_[44430]_  = \new_[44429]_  & \new_[44426]_ ;
  assign \new_[44433]_  = A266 & ~A265;
  assign \new_[44436]_  = A269 & ~A268;
  assign \new_[44437]_  = \new_[44436]_  & \new_[44433]_ ;
  assign \new_[44438]_  = \new_[44437]_  & \new_[44430]_ ;
  assign \new_[44441]_  = A168 & A169;
  assign \new_[44444]_  = A166 & ~A167;
  assign \new_[44445]_  = \new_[44444]_  & \new_[44441]_ ;
  assign \new_[44448]_  = A200 & A199;
  assign \new_[44451]_  = ~A202 & ~A201;
  assign \new_[44452]_  = \new_[44451]_  & \new_[44448]_ ;
  assign \new_[44453]_  = \new_[44452]_  & \new_[44445]_ ;
  assign \new_[44456]_  = ~A233 & A232;
  assign \new_[44459]_  = A236 & ~A235;
  assign \new_[44460]_  = \new_[44459]_  & \new_[44456]_ ;
  assign \new_[44463]_  = ~A266 & A265;
  assign \new_[44466]_  = A269 & ~A268;
  assign \new_[44467]_  = \new_[44466]_  & \new_[44463]_ ;
  assign \new_[44468]_  = \new_[44467]_  & \new_[44460]_ ;
  assign \new_[44471]_  = A168 & A169;
  assign \new_[44474]_  = A166 & ~A167;
  assign \new_[44475]_  = \new_[44474]_  & \new_[44471]_ ;
  assign \new_[44478]_  = A200 & A199;
  assign \new_[44481]_  = ~A202 & ~A201;
  assign \new_[44482]_  = \new_[44481]_  & \new_[44478]_ ;
  assign \new_[44483]_  = \new_[44482]_  & \new_[44475]_ ;
  assign \new_[44486]_  = ~A233 & A232;
  assign \new_[44489]_  = A236 & ~A235;
  assign \new_[44490]_  = \new_[44489]_  & \new_[44486]_ ;
  assign \new_[44493]_  = ~A266 & ~A265;
  assign \new_[44496]_  = ~A269 & A268;
  assign \new_[44497]_  = \new_[44496]_  & \new_[44493]_ ;
  assign \new_[44498]_  = \new_[44497]_  & \new_[44490]_ ;
  assign \new_[44501]_  = A168 & A169;
  assign \new_[44504]_  = A166 & ~A167;
  assign \new_[44505]_  = \new_[44504]_  & \new_[44501]_ ;
  assign \new_[44508]_  = A200 & A199;
  assign \new_[44511]_  = ~A202 & ~A201;
  assign \new_[44512]_  = \new_[44511]_  & \new_[44508]_ ;
  assign \new_[44513]_  = \new_[44512]_  & \new_[44505]_ ;
  assign \new_[44516]_  = ~A233 & ~A232;
  assign \new_[44519]_  = ~A236 & A235;
  assign \new_[44520]_  = \new_[44519]_  & \new_[44516]_ ;
  assign \new_[44523]_  = A299 & A298;
  assign \new_[44526]_  = ~A302 & A301;
  assign \new_[44527]_  = \new_[44526]_  & \new_[44523]_ ;
  assign \new_[44528]_  = \new_[44527]_  & \new_[44520]_ ;
  assign \new_[44531]_  = A168 & A169;
  assign \new_[44534]_  = A166 & ~A167;
  assign \new_[44535]_  = \new_[44534]_  & \new_[44531]_ ;
  assign \new_[44538]_  = A200 & A199;
  assign \new_[44541]_  = ~A202 & ~A201;
  assign \new_[44542]_  = \new_[44541]_  & \new_[44538]_ ;
  assign \new_[44543]_  = \new_[44542]_  & \new_[44535]_ ;
  assign \new_[44546]_  = ~A233 & ~A232;
  assign \new_[44549]_  = ~A236 & A235;
  assign \new_[44550]_  = \new_[44549]_  & \new_[44546]_ ;
  assign \new_[44553]_  = ~A299 & A298;
  assign \new_[44556]_  = A302 & ~A301;
  assign \new_[44557]_  = \new_[44556]_  & \new_[44553]_ ;
  assign \new_[44558]_  = \new_[44557]_  & \new_[44550]_ ;
  assign \new_[44561]_  = A168 & A169;
  assign \new_[44564]_  = A166 & ~A167;
  assign \new_[44565]_  = \new_[44564]_  & \new_[44561]_ ;
  assign \new_[44568]_  = A200 & A199;
  assign \new_[44571]_  = ~A202 & ~A201;
  assign \new_[44572]_  = \new_[44571]_  & \new_[44568]_ ;
  assign \new_[44573]_  = \new_[44572]_  & \new_[44565]_ ;
  assign \new_[44576]_  = ~A233 & ~A232;
  assign \new_[44579]_  = ~A236 & A235;
  assign \new_[44580]_  = \new_[44579]_  & \new_[44576]_ ;
  assign \new_[44583]_  = A299 & ~A298;
  assign \new_[44586]_  = A302 & ~A301;
  assign \new_[44587]_  = \new_[44586]_  & \new_[44583]_ ;
  assign \new_[44588]_  = \new_[44587]_  & \new_[44580]_ ;
  assign \new_[44591]_  = A168 & A169;
  assign \new_[44594]_  = A166 & ~A167;
  assign \new_[44595]_  = \new_[44594]_  & \new_[44591]_ ;
  assign \new_[44598]_  = A200 & A199;
  assign \new_[44601]_  = ~A202 & ~A201;
  assign \new_[44602]_  = \new_[44601]_  & \new_[44598]_ ;
  assign \new_[44603]_  = \new_[44602]_  & \new_[44595]_ ;
  assign \new_[44606]_  = ~A233 & ~A232;
  assign \new_[44609]_  = ~A236 & A235;
  assign \new_[44610]_  = \new_[44609]_  & \new_[44606]_ ;
  assign \new_[44613]_  = ~A299 & ~A298;
  assign \new_[44616]_  = ~A302 & A301;
  assign \new_[44617]_  = \new_[44616]_  & \new_[44613]_ ;
  assign \new_[44618]_  = \new_[44617]_  & \new_[44610]_ ;
  assign \new_[44621]_  = A168 & A169;
  assign \new_[44624]_  = A166 & ~A167;
  assign \new_[44625]_  = \new_[44624]_  & \new_[44621]_ ;
  assign \new_[44628]_  = A200 & A199;
  assign \new_[44631]_  = ~A202 & ~A201;
  assign \new_[44632]_  = \new_[44631]_  & \new_[44628]_ ;
  assign \new_[44633]_  = \new_[44632]_  & \new_[44625]_ ;
  assign \new_[44636]_  = ~A233 & ~A232;
  assign \new_[44639]_  = ~A236 & A235;
  assign \new_[44640]_  = \new_[44639]_  & \new_[44636]_ ;
  assign \new_[44643]_  = A266 & A265;
  assign \new_[44646]_  = ~A269 & A268;
  assign \new_[44647]_  = \new_[44646]_  & \new_[44643]_ ;
  assign \new_[44648]_  = \new_[44647]_  & \new_[44640]_ ;
  assign \new_[44651]_  = A168 & A169;
  assign \new_[44654]_  = A166 & ~A167;
  assign \new_[44655]_  = \new_[44654]_  & \new_[44651]_ ;
  assign \new_[44658]_  = A200 & A199;
  assign \new_[44661]_  = ~A202 & ~A201;
  assign \new_[44662]_  = \new_[44661]_  & \new_[44658]_ ;
  assign \new_[44663]_  = \new_[44662]_  & \new_[44655]_ ;
  assign \new_[44666]_  = ~A233 & ~A232;
  assign \new_[44669]_  = ~A236 & A235;
  assign \new_[44670]_  = \new_[44669]_  & \new_[44666]_ ;
  assign \new_[44673]_  = A266 & ~A265;
  assign \new_[44676]_  = A269 & ~A268;
  assign \new_[44677]_  = \new_[44676]_  & \new_[44673]_ ;
  assign \new_[44678]_  = \new_[44677]_  & \new_[44670]_ ;
  assign \new_[44681]_  = A168 & A169;
  assign \new_[44684]_  = A166 & ~A167;
  assign \new_[44685]_  = \new_[44684]_  & \new_[44681]_ ;
  assign \new_[44688]_  = A200 & A199;
  assign \new_[44691]_  = ~A202 & ~A201;
  assign \new_[44692]_  = \new_[44691]_  & \new_[44688]_ ;
  assign \new_[44693]_  = \new_[44692]_  & \new_[44685]_ ;
  assign \new_[44696]_  = ~A233 & ~A232;
  assign \new_[44699]_  = ~A236 & A235;
  assign \new_[44700]_  = \new_[44699]_  & \new_[44696]_ ;
  assign \new_[44703]_  = ~A266 & A265;
  assign \new_[44706]_  = A269 & ~A268;
  assign \new_[44707]_  = \new_[44706]_  & \new_[44703]_ ;
  assign \new_[44708]_  = \new_[44707]_  & \new_[44700]_ ;
  assign \new_[44711]_  = A168 & A169;
  assign \new_[44714]_  = A166 & ~A167;
  assign \new_[44715]_  = \new_[44714]_  & \new_[44711]_ ;
  assign \new_[44718]_  = A200 & A199;
  assign \new_[44721]_  = ~A202 & ~A201;
  assign \new_[44722]_  = \new_[44721]_  & \new_[44718]_ ;
  assign \new_[44723]_  = \new_[44722]_  & \new_[44715]_ ;
  assign \new_[44726]_  = ~A233 & ~A232;
  assign \new_[44729]_  = ~A236 & A235;
  assign \new_[44730]_  = \new_[44729]_  & \new_[44726]_ ;
  assign \new_[44733]_  = ~A266 & ~A265;
  assign \new_[44736]_  = ~A269 & A268;
  assign \new_[44737]_  = \new_[44736]_  & \new_[44733]_ ;
  assign \new_[44738]_  = \new_[44737]_  & \new_[44730]_ ;
  assign \new_[44741]_  = A168 & A169;
  assign \new_[44744]_  = A166 & ~A167;
  assign \new_[44745]_  = \new_[44744]_  & \new_[44741]_ ;
  assign \new_[44748]_  = A200 & A199;
  assign \new_[44751]_  = A203 & ~A201;
  assign \new_[44752]_  = \new_[44751]_  & \new_[44748]_ ;
  assign \new_[44753]_  = \new_[44752]_  & \new_[44745]_ ;
  assign \new_[44756]_  = A233 & A232;
  assign \new_[44759]_  = ~A236 & A235;
  assign \new_[44760]_  = \new_[44759]_  & \new_[44756]_ ;
  assign \new_[44763]_  = A299 & A298;
  assign \new_[44766]_  = ~A302 & A301;
  assign \new_[44767]_  = \new_[44766]_  & \new_[44763]_ ;
  assign \new_[44768]_  = \new_[44767]_  & \new_[44760]_ ;
  assign \new_[44771]_  = A168 & A169;
  assign \new_[44774]_  = A166 & ~A167;
  assign \new_[44775]_  = \new_[44774]_  & \new_[44771]_ ;
  assign \new_[44778]_  = A200 & A199;
  assign \new_[44781]_  = A203 & ~A201;
  assign \new_[44782]_  = \new_[44781]_  & \new_[44778]_ ;
  assign \new_[44783]_  = \new_[44782]_  & \new_[44775]_ ;
  assign \new_[44786]_  = A233 & A232;
  assign \new_[44789]_  = ~A236 & A235;
  assign \new_[44790]_  = \new_[44789]_  & \new_[44786]_ ;
  assign \new_[44793]_  = ~A299 & A298;
  assign \new_[44796]_  = A302 & ~A301;
  assign \new_[44797]_  = \new_[44796]_  & \new_[44793]_ ;
  assign \new_[44798]_  = \new_[44797]_  & \new_[44790]_ ;
  assign \new_[44801]_  = A168 & A169;
  assign \new_[44804]_  = A166 & ~A167;
  assign \new_[44805]_  = \new_[44804]_  & \new_[44801]_ ;
  assign \new_[44808]_  = A200 & A199;
  assign \new_[44811]_  = A203 & ~A201;
  assign \new_[44812]_  = \new_[44811]_  & \new_[44808]_ ;
  assign \new_[44813]_  = \new_[44812]_  & \new_[44805]_ ;
  assign \new_[44816]_  = A233 & A232;
  assign \new_[44819]_  = ~A236 & A235;
  assign \new_[44820]_  = \new_[44819]_  & \new_[44816]_ ;
  assign \new_[44823]_  = A299 & ~A298;
  assign \new_[44826]_  = A302 & ~A301;
  assign \new_[44827]_  = \new_[44826]_  & \new_[44823]_ ;
  assign \new_[44828]_  = \new_[44827]_  & \new_[44820]_ ;
  assign \new_[44831]_  = A168 & A169;
  assign \new_[44834]_  = A166 & ~A167;
  assign \new_[44835]_  = \new_[44834]_  & \new_[44831]_ ;
  assign \new_[44838]_  = A200 & A199;
  assign \new_[44841]_  = A203 & ~A201;
  assign \new_[44842]_  = \new_[44841]_  & \new_[44838]_ ;
  assign \new_[44843]_  = \new_[44842]_  & \new_[44835]_ ;
  assign \new_[44846]_  = A233 & A232;
  assign \new_[44849]_  = ~A236 & A235;
  assign \new_[44850]_  = \new_[44849]_  & \new_[44846]_ ;
  assign \new_[44853]_  = ~A299 & ~A298;
  assign \new_[44856]_  = ~A302 & A301;
  assign \new_[44857]_  = \new_[44856]_  & \new_[44853]_ ;
  assign \new_[44858]_  = \new_[44857]_  & \new_[44850]_ ;
  assign \new_[44861]_  = A168 & A169;
  assign \new_[44864]_  = A166 & ~A167;
  assign \new_[44865]_  = \new_[44864]_  & \new_[44861]_ ;
  assign \new_[44868]_  = A200 & A199;
  assign \new_[44871]_  = A203 & ~A201;
  assign \new_[44872]_  = \new_[44871]_  & \new_[44868]_ ;
  assign \new_[44873]_  = \new_[44872]_  & \new_[44865]_ ;
  assign \new_[44876]_  = A233 & A232;
  assign \new_[44879]_  = ~A236 & A235;
  assign \new_[44880]_  = \new_[44879]_  & \new_[44876]_ ;
  assign \new_[44883]_  = A266 & A265;
  assign \new_[44886]_  = ~A269 & A268;
  assign \new_[44887]_  = \new_[44886]_  & \new_[44883]_ ;
  assign \new_[44888]_  = \new_[44887]_  & \new_[44880]_ ;
  assign \new_[44891]_  = A168 & A169;
  assign \new_[44894]_  = A166 & ~A167;
  assign \new_[44895]_  = \new_[44894]_  & \new_[44891]_ ;
  assign \new_[44898]_  = A200 & A199;
  assign \new_[44901]_  = A203 & ~A201;
  assign \new_[44902]_  = \new_[44901]_  & \new_[44898]_ ;
  assign \new_[44903]_  = \new_[44902]_  & \new_[44895]_ ;
  assign \new_[44906]_  = A233 & A232;
  assign \new_[44909]_  = ~A236 & A235;
  assign \new_[44910]_  = \new_[44909]_  & \new_[44906]_ ;
  assign \new_[44913]_  = A266 & ~A265;
  assign \new_[44916]_  = A269 & ~A268;
  assign \new_[44917]_  = \new_[44916]_  & \new_[44913]_ ;
  assign \new_[44918]_  = \new_[44917]_  & \new_[44910]_ ;
  assign \new_[44921]_  = A168 & A169;
  assign \new_[44924]_  = A166 & ~A167;
  assign \new_[44925]_  = \new_[44924]_  & \new_[44921]_ ;
  assign \new_[44928]_  = A200 & A199;
  assign \new_[44931]_  = A203 & ~A201;
  assign \new_[44932]_  = \new_[44931]_  & \new_[44928]_ ;
  assign \new_[44933]_  = \new_[44932]_  & \new_[44925]_ ;
  assign \new_[44936]_  = A233 & A232;
  assign \new_[44939]_  = ~A236 & A235;
  assign \new_[44940]_  = \new_[44939]_  & \new_[44936]_ ;
  assign \new_[44943]_  = ~A266 & A265;
  assign \new_[44946]_  = A269 & ~A268;
  assign \new_[44947]_  = \new_[44946]_  & \new_[44943]_ ;
  assign \new_[44948]_  = \new_[44947]_  & \new_[44940]_ ;
  assign \new_[44951]_  = A168 & A169;
  assign \new_[44954]_  = A166 & ~A167;
  assign \new_[44955]_  = \new_[44954]_  & \new_[44951]_ ;
  assign \new_[44958]_  = A200 & A199;
  assign \new_[44961]_  = A203 & ~A201;
  assign \new_[44962]_  = \new_[44961]_  & \new_[44958]_ ;
  assign \new_[44963]_  = \new_[44962]_  & \new_[44955]_ ;
  assign \new_[44966]_  = A233 & A232;
  assign \new_[44969]_  = ~A236 & A235;
  assign \new_[44970]_  = \new_[44969]_  & \new_[44966]_ ;
  assign \new_[44973]_  = ~A266 & ~A265;
  assign \new_[44976]_  = ~A269 & A268;
  assign \new_[44977]_  = \new_[44976]_  & \new_[44973]_ ;
  assign \new_[44978]_  = \new_[44977]_  & \new_[44970]_ ;
  assign \new_[44981]_  = A168 & A169;
  assign \new_[44984]_  = A166 & ~A167;
  assign \new_[44985]_  = \new_[44984]_  & \new_[44981]_ ;
  assign \new_[44988]_  = A200 & A199;
  assign \new_[44991]_  = A203 & ~A201;
  assign \new_[44992]_  = \new_[44991]_  & \new_[44988]_ ;
  assign \new_[44993]_  = \new_[44992]_  & \new_[44985]_ ;
  assign \new_[44996]_  = A233 & ~A232;
  assign \new_[44999]_  = A236 & ~A235;
  assign \new_[45000]_  = \new_[44999]_  & \new_[44996]_ ;
  assign \new_[45003]_  = A299 & A298;
  assign \new_[45006]_  = ~A302 & A301;
  assign \new_[45007]_  = \new_[45006]_  & \new_[45003]_ ;
  assign \new_[45008]_  = \new_[45007]_  & \new_[45000]_ ;
  assign \new_[45011]_  = A168 & A169;
  assign \new_[45014]_  = A166 & ~A167;
  assign \new_[45015]_  = \new_[45014]_  & \new_[45011]_ ;
  assign \new_[45018]_  = A200 & A199;
  assign \new_[45021]_  = A203 & ~A201;
  assign \new_[45022]_  = \new_[45021]_  & \new_[45018]_ ;
  assign \new_[45023]_  = \new_[45022]_  & \new_[45015]_ ;
  assign \new_[45026]_  = A233 & ~A232;
  assign \new_[45029]_  = A236 & ~A235;
  assign \new_[45030]_  = \new_[45029]_  & \new_[45026]_ ;
  assign \new_[45033]_  = ~A299 & A298;
  assign \new_[45036]_  = A302 & ~A301;
  assign \new_[45037]_  = \new_[45036]_  & \new_[45033]_ ;
  assign \new_[45038]_  = \new_[45037]_  & \new_[45030]_ ;
  assign \new_[45041]_  = A168 & A169;
  assign \new_[45044]_  = A166 & ~A167;
  assign \new_[45045]_  = \new_[45044]_  & \new_[45041]_ ;
  assign \new_[45048]_  = A200 & A199;
  assign \new_[45051]_  = A203 & ~A201;
  assign \new_[45052]_  = \new_[45051]_  & \new_[45048]_ ;
  assign \new_[45053]_  = \new_[45052]_  & \new_[45045]_ ;
  assign \new_[45056]_  = A233 & ~A232;
  assign \new_[45059]_  = A236 & ~A235;
  assign \new_[45060]_  = \new_[45059]_  & \new_[45056]_ ;
  assign \new_[45063]_  = A299 & ~A298;
  assign \new_[45066]_  = A302 & ~A301;
  assign \new_[45067]_  = \new_[45066]_  & \new_[45063]_ ;
  assign \new_[45068]_  = \new_[45067]_  & \new_[45060]_ ;
  assign \new_[45071]_  = A168 & A169;
  assign \new_[45074]_  = A166 & ~A167;
  assign \new_[45075]_  = \new_[45074]_  & \new_[45071]_ ;
  assign \new_[45078]_  = A200 & A199;
  assign \new_[45081]_  = A203 & ~A201;
  assign \new_[45082]_  = \new_[45081]_  & \new_[45078]_ ;
  assign \new_[45083]_  = \new_[45082]_  & \new_[45075]_ ;
  assign \new_[45086]_  = A233 & ~A232;
  assign \new_[45089]_  = A236 & ~A235;
  assign \new_[45090]_  = \new_[45089]_  & \new_[45086]_ ;
  assign \new_[45093]_  = ~A299 & ~A298;
  assign \new_[45096]_  = ~A302 & A301;
  assign \new_[45097]_  = \new_[45096]_  & \new_[45093]_ ;
  assign \new_[45098]_  = \new_[45097]_  & \new_[45090]_ ;
  assign \new_[45101]_  = A168 & A169;
  assign \new_[45104]_  = A166 & ~A167;
  assign \new_[45105]_  = \new_[45104]_  & \new_[45101]_ ;
  assign \new_[45108]_  = A200 & A199;
  assign \new_[45111]_  = A203 & ~A201;
  assign \new_[45112]_  = \new_[45111]_  & \new_[45108]_ ;
  assign \new_[45113]_  = \new_[45112]_  & \new_[45105]_ ;
  assign \new_[45116]_  = A233 & ~A232;
  assign \new_[45119]_  = A236 & ~A235;
  assign \new_[45120]_  = \new_[45119]_  & \new_[45116]_ ;
  assign \new_[45123]_  = A266 & A265;
  assign \new_[45126]_  = ~A269 & A268;
  assign \new_[45127]_  = \new_[45126]_  & \new_[45123]_ ;
  assign \new_[45128]_  = \new_[45127]_  & \new_[45120]_ ;
  assign \new_[45131]_  = A168 & A169;
  assign \new_[45134]_  = A166 & ~A167;
  assign \new_[45135]_  = \new_[45134]_  & \new_[45131]_ ;
  assign \new_[45138]_  = A200 & A199;
  assign \new_[45141]_  = A203 & ~A201;
  assign \new_[45142]_  = \new_[45141]_  & \new_[45138]_ ;
  assign \new_[45143]_  = \new_[45142]_  & \new_[45135]_ ;
  assign \new_[45146]_  = A233 & ~A232;
  assign \new_[45149]_  = A236 & ~A235;
  assign \new_[45150]_  = \new_[45149]_  & \new_[45146]_ ;
  assign \new_[45153]_  = A266 & ~A265;
  assign \new_[45156]_  = A269 & ~A268;
  assign \new_[45157]_  = \new_[45156]_  & \new_[45153]_ ;
  assign \new_[45158]_  = \new_[45157]_  & \new_[45150]_ ;
  assign \new_[45161]_  = A168 & A169;
  assign \new_[45164]_  = A166 & ~A167;
  assign \new_[45165]_  = \new_[45164]_  & \new_[45161]_ ;
  assign \new_[45168]_  = A200 & A199;
  assign \new_[45171]_  = A203 & ~A201;
  assign \new_[45172]_  = \new_[45171]_  & \new_[45168]_ ;
  assign \new_[45173]_  = \new_[45172]_  & \new_[45165]_ ;
  assign \new_[45176]_  = A233 & ~A232;
  assign \new_[45179]_  = A236 & ~A235;
  assign \new_[45180]_  = \new_[45179]_  & \new_[45176]_ ;
  assign \new_[45183]_  = ~A266 & A265;
  assign \new_[45186]_  = A269 & ~A268;
  assign \new_[45187]_  = \new_[45186]_  & \new_[45183]_ ;
  assign \new_[45188]_  = \new_[45187]_  & \new_[45180]_ ;
  assign \new_[45191]_  = A168 & A169;
  assign \new_[45194]_  = A166 & ~A167;
  assign \new_[45195]_  = \new_[45194]_  & \new_[45191]_ ;
  assign \new_[45198]_  = A200 & A199;
  assign \new_[45201]_  = A203 & ~A201;
  assign \new_[45202]_  = \new_[45201]_  & \new_[45198]_ ;
  assign \new_[45203]_  = \new_[45202]_  & \new_[45195]_ ;
  assign \new_[45206]_  = A233 & ~A232;
  assign \new_[45209]_  = A236 & ~A235;
  assign \new_[45210]_  = \new_[45209]_  & \new_[45206]_ ;
  assign \new_[45213]_  = ~A266 & ~A265;
  assign \new_[45216]_  = ~A269 & A268;
  assign \new_[45217]_  = \new_[45216]_  & \new_[45213]_ ;
  assign \new_[45218]_  = \new_[45217]_  & \new_[45210]_ ;
  assign \new_[45221]_  = A168 & A169;
  assign \new_[45224]_  = A166 & ~A167;
  assign \new_[45225]_  = \new_[45224]_  & \new_[45221]_ ;
  assign \new_[45228]_  = A200 & A199;
  assign \new_[45231]_  = A203 & ~A201;
  assign \new_[45232]_  = \new_[45231]_  & \new_[45228]_ ;
  assign \new_[45233]_  = \new_[45232]_  & \new_[45225]_ ;
  assign \new_[45236]_  = ~A233 & A232;
  assign \new_[45239]_  = A236 & ~A235;
  assign \new_[45240]_  = \new_[45239]_  & \new_[45236]_ ;
  assign \new_[45243]_  = A299 & A298;
  assign \new_[45246]_  = ~A302 & A301;
  assign \new_[45247]_  = \new_[45246]_  & \new_[45243]_ ;
  assign \new_[45248]_  = \new_[45247]_  & \new_[45240]_ ;
  assign \new_[45251]_  = A168 & A169;
  assign \new_[45254]_  = A166 & ~A167;
  assign \new_[45255]_  = \new_[45254]_  & \new_[45251]_ ;
  assign \new_[45258]_  = A200 & A199;
  assign \new_[45261]_  = A203 & ~A201;
  assign \new_[45262]_  = \new_[45261]_  & \new_[45258]_ ;
  assign \new_[45263]_  = \new_[45262]_  & \new_[45255]_ ;
  assign \new_[45266]_  = ~A233 & A232;
  assign \new_[45269]_  = A236 & ~A235;
  assign \new_[45270]_  = \new_[45269]_  & \new_[45266]_ ;
  assign \new_[45273]_  = ~A299 & A298;
  assign \new_[45276]_  = A302 & ~A301;
  assign \new_[45277]_  = \new_[45276]_  & \new_[45273]_ ;
  assign \new_[45278]_  = \new_[45277]_  & \new_[45270]_ ;
  assign \new_[45281]_  = A168 & A169;
  assign \new_[45284]_  = A166 & ~A167;
  assign \new_[45285]_  = \new_[45284]_  & \new_[45281]_ ;
  assign \new_[45288]_  = A200 & A199;
  assign \new_[45291]_  = A203 & ~A201;
  assign \new_[45292]_  = \new_[45291]_  & \new_[45288]_ ;
  assign \new_[45293]_  = \new_[45292]_  & \new_[45285]_ ;
  assign \new_[45296]_  = ~A233 & A232;
  assign \new_[45299]_  = A236 & ~A235;
  assign \new_[45300]_  = \new_[45299]_  & \new_[45296]_ ;
  assign \new_[45303]_  = A299 & ~A298;
  assign \new_[45306]_  = A302 & ~A301;
  assign \new_[45307]_  = \new_[45306]_  & \new_[45303]_ ;
  assign \new_[45308]_  = \new_[45307]_  & \new_[45300]_ ;
  assign \new_[45311]_  = A168 & A169;
  assign \new_[45314]_  = A166 & ~A167;
  assign \new_[45315]_  = \new_[45314]_  & \new_[45311]_ ;
  assign \new_[45318]_  = A200 & A199;
  assign \new_[45321]_  = A203 & ~A201;
  assign \new_[45322]_  = \new_[45321]_  & \new_[45318]_ ;
  assign \new_[45323]_  = \new_[45322]_  & \new_[45315]_ ;
  assign \new_[45326]_  = ~A233 & A232;
  assign \new_[45329]_  = A236 & ~A235;
  assign \new_[45330]_  = \new_[45329]_  & \new_[45326]_ ;
  assign \new_[45333]_  = ~A299 & ~A298;
  assign \new_[45336]_  = ~A302 & A301;
  assign \new_[45337]_  = \new_[45336]_  & \new_[45333]_ ;
  assign \new_[45338]_  = \new_[45337]_  & \new_[45330]_ ;
  assign \new_[45341]_  = A168 & A169;
  assign \new_[45344]_  = A166 & ~A167;
  assign \new_[45345]_  = \new_[45344]_  & \new_[45341]_ ;
  assign \new_[45348]_  = A200 & A199;
  assign \new_[45351]_  = A203 & ~A201;
  assign \new_[45352]_  = \new_[45351]_  & \new_[45348]_ ;
  assign \new_[45353]_  = \new_[45352]_  & \new_[45345]_ ;
  assign \new_[45356]_  = ~A233 & A232;
  assign \new_[45359]_  = A236 & ~A235;
  assign \new_[45360]_  = \new_[45359]_  & \new_[45356]_ ;
  assign \new_[45363]_  = A266 & A265;
  assign \new_[45366]_  = ~A269 & A268;
  assign \new_[45367]_  = \new_[45366]_  & \new_[45363]_ ;
  assign \new_[45368]_  = \new_[45367]_  & \new_[45360]_ ;
  assign \new_[45371]_  = A168 & A169;
  assign \new_[45374]_  = A166 & ~A167;
  assign \new_[45375]_  = \new_[45374]_  & \new_[45371]_ ;
  assign \new_[45378]_  = A200 & A199;
  assign \new_[45381]_  = A203 & ~A201;
  assign \new_[45382]_  = \new_[45381]_  & \new_[45378]_ ;
  assign \new_[45383]_  = \new_[45382]_  & \new_[45375]_ ;
  assign \new_[45386]_  = ~A233 & A232;
  assign \new_[45389]_  = A236 & ~A235;
  assign \new_[45390]_  = \new_[45389]_  & \new_[45386]_ ;
  assign \new_[45393]_  = A266 & ~A265;
  assign \new_[45396]_  = A269 & ~A268;
  assign \new_[45397]_  = \new_[45396]_  & \new_[45393]_ ;
  assign \new_[45398]_  = \new_[45397]_  & \new_[45390]_ ;
  assign \new_[45401]_  = A168 & A169;
  assign \new_[45404]_  = A166 & ~A167;
  assign \new_[45405]_  = \new_[45404]_  & \new_[45401]_ ;
  assign \new_[45408]_  = A200 & A199;
  assign \new_[45411]_  = A203 & ~A201;
  assign \new_[45412]_  = \new_[45411]_  & \new_[45408]_ ;
  assign \new_[45413]_  = \new_[45412]_  & \new_[45405]_ ;
  assign \new_[45416]_  = ~A233 & A232;
  assign \new_[45419]_  = A236 & ~A235;
  assign \new_[45420]_  = \new_[45419]_  & \new_[45416]_ ;
  assign \new_[45423]_  = ~A266 & A265;
  assign \new_[45426]_  = A269 & ~A268;
  assign \new_[45427]_  = \new_[45426]_  & \new_[45423]_ ;
  assign \new_[45428]_  = \new_[45427]_  & \new_[45420]_ ;
  assign \new_[45431]_  = A168 & A169;
  assign \new_[45434]_  = A166 & ~A167;
  assign \new_[45435]_  = \new_[45434]_  & \new_[45431]_ ;
  assign \new_[45438]_  = A200 & A199;
  assign \new_[45441]_  = A203 & ~A201;
  assign \new_[45442]_  = \new_[45441]_  & \new_[45438]_ ;
  assign \new_[45443]_  = \new_[45442]_  & \new_[45435]_ ;
  assign \new_[45446]_  = ~A233 & A232;
  assign \new_[45449]_  = A236 & ~A235;
  assign \new_[45450]_  = \new_[45449]_  & \new_[45446]_ ;
  assign \new_[45453]_  = ~A266 & ~A265;
  assign \new_[45456]_  = ~A269 & A268;
  assign \new_[45457]_  = \new_[45456]_  & \new_[45453]_ ;
  assign \new_[45458]_  = \new_[45457]_  & \new_[45450]_ ;
  assign \new_[45461]_  = A168 & A169;
  assign \new_[45464]_  = A166 & ~A167;
  assign \new_[45465]_  = \new_[45464]_  & \new_[45461]_ ;
  assign \new_[45468]_  = A200 & A199;
  assign \new_[45471]_  = A203 & ~A201;
  assign \new_[45472]_  = \new_[45471]_  & \new_[45468]_ ;
  assign \new_[45473]_  = \new_[45472]_  & \new_[45465]_ ;
  assign \new_[45476]_  = ~A233 & ~A232;
  assign \new_[45479]_  = ~A236 & A235;
  assign \new_[45480]_  = \new_[45479]_  & \new_[45476]_ ;
  assign \new_[45483]_  = A299 & A298;
  assign \new_[45486]_  = ~A302 & A301;
  assign \new_[45487]_  = \new_[45486]_  & \new_[45483]_ ;
  assign \new_[45488]_  = \new_[45487]_  & \new_[45480]_ ;
  assign \new_[45491]_  = A168 & A169;
  assign \new_[45494]_  = A166 & ~A167;
  assign \new_[45495]_  = \new_[45494]_  & \new_[45491]_ ;
  assign \new_[45498]_  = A200 & A199;
  assign \new_[45501]_  = A203 & ~A201;
  assign \new_[45502]_  = \new_[45501]_  & \new_[45498]_ ;
  assign \new_[45503]_  = \new_[45502]_  & \new_[45495]_ ;
  assign \new_[45506]_  = ~A233 & ~A232;
  assign \new_[45509]_  = ~A236 & A235;
  assign \new_[45510]_  = \new_[45509]_  & \new_[45506]_ ;
  assign \new_[45513]_  = ~A299 & A298;
  assign \new_[45516]_  = A302 & ~A301;
  assign \new_[45517]_  = \new_[45516]_  & \new_[45513]_ ;
  assign \new_[45518]_  = \new_[45517]_  & \new_[45510]_ ;
  assign \new_[45521]_  = A168 & A169;
  assign \new_[45524]_  = A166 & ~A167;
  assign \new_[45525]_  = \new_[45524]_  & \new_[45521]_ ;
  assign \new_[45528]_  = A200 & A199;
  assign \new_[45531]_  = A203 & ~A201;
  assign \new_[45532]_  = \new_[45531]_  & \new_[45528]_ ;
  assign \new_[45533]_  = \new_[45532]_  & \new_[45525]_ ;
  assign \new_[45536]_  = ~A233 & ~A232;
  assign \new_[45539]_  = ~A236 & A235;
  assign \new_[45540]_  = \new_[45539]_  & \new_[45536]_ ;
  assign \new_[45543]_  = A299 & ~A298;
  assign \new_[45546]_  = A302 & ~A301;
  assign \new_[45547]_  = \new_[45546]_  & \new_[45543]_ ;
  assign \new_[45548]_  = \new_[45547]_  & \new_[45540]_ ;
  assign \new_[45551]_  = A168 & A169;
  assign \new_[45554]_  = A166 & ~A167;
  assign \new_[45555]_  = \new_[45554]_  & \new_[45551]_ ;
  assign \new_[45558]_  = A200 & A199;
  assign \new_[45561]_  = A203 & ~A201;
  assign \new_[45562]_  = \new_[45561]_  & \new_[45558]_ ;
  assign \new_[45563]_  = \new_[45562]_  & \new_[45555]_ ;
  assign \new_[45566]_  = ~A233 & ~A232;
  assign \new_[45569]_  = ~A236 & A235;
  assign \new_[45570]_  = \new_[45569]_  & \new_[45566]_ ;
  assign \new_[45573]_  = ~A299 & ~A298;
  assign \new_[45576]_  = ~A302 & A301;
  assign \new_[45577]_  = \new_[45576]_  & \new_[45573]_ ;
  assign \new_[45578]_  = \new_[45577]_  & \new_[45570]_ ;
  assign \new_[45581]_  = A168 & A169;
  assign \new_[45584]_  = A166 & ~A167;
  assign \new_[45585]_  = \new_[45584]_  & \new_[45581]_ ;
  assign \new_[45588]_  = A200 & A199;
  assign \new_[45591]_  = A203 & ~A201;
  assign \new_[45592]_  = \new_[45591]_  & \new_[45588]_ ;
  assign \new_[45593]_  = \new_[45592]_  & \new_[45585]_ ;
  assign \new_[45596]_  = ~A233 & ~A232;
  assign \new_[45599]_  = ~A236 & A235;
  assign \new_[45600]_  = \new_[45599]_  & \new_[45596]_ ;
  assign \new_[45603]_  = A266 & A265;
  assign \new_[45606]_  = ~A269 & A268;
  assign \new_[45607]_  = \new_[45606]_  & \new_[45603]_ ;
  assign \new_[45608]_  = \new_[45607]_  & \new_[45600]_ ;
  assign \new_[45611]_  = A168 & A169;
  assign \new_[45614]_  = A166 & ~A167;
  assign \new_[45615]_  = \new_[45614]_  & \new_[45611]_ ;
  assign \new_[45618]_  = A200 & A199;
  assign \new_[45621]_  = A203 & ~A201;
  assign \new_[45622]_  = \new_[45621]_  & \new_[45618]_ ;
  assign \new_[45623]_  = \new_[45622]_  & \new_[45615]_ ;
  assign \new_[45626]_  = ~A233 & ~A232;
  assign \new_[45629]_  = ~A236 & A235;
  assign \new_[45630]_  = \new_[45629]_  & \new_[45626]_ ;
  assign \new_[45633]_  = A266 & ~A265;
  assign \new_[45636]_  = A269 & ~A268;
  assign \new_[45637]_  = \new_[45636]_  & \new_[45633]_ ;
  assign \new_[45638]_  = \new_[45637]_  & \new_[45630]_ ;
  assign \new_[45641]_  = A168 & A169;
  assign \new_[45644]_  = A166 & ~A167;
  assign \new_[45645]_  = \new_[45644]_  & \new_[45641]_ ;
  assign \new_[45648]_  = A200 & A199;
  assign \new_[45651]_  = A203 & ~A201;
  assign \new_[45652]_  = \new_[45651]_  & \new_[45648]_ ;
  assign \new_[45653]_  = \new_[45652]_  & \new_[45645]_ ;
  assign \new_[45656]_  = ~A233 & ~A232;
  assign \new_[45659]_  = ~A236 & A235;
  assign \new_[45660]_  = \new_[45659]_  & \new_[45656]_ ;
  assign \new_[45663]_  = ~A266 & A265;
  assign \new_[45666]_  = A269 & ~A268;
  assign \new_[45667]_  = \new_[45666]_  & \new_[45663]_ ;
  assign \new_[45668]_  = \new_[45667]_  & \new_[45660]_ ;
  assign \new_[45671]_  = A168 & A169;
  assign \new_[45674]_  = A166 & ~A167;
  assign \new_[45675]_  = \new_[45674]_  & \new_[45671]_ ;
  assign \new_[45678]_  = A200 & A199;
  assign \new_[45681]_  = A203 & ~A201;
  assign \new_[45682]_  = \new_[45681]_  & \new_[45678]_ ;
  assign \new_[45683]_  = \new_[45682]_  & \new_[45675]_ ;
  assign \new_[45686]_  = ~A233 & ~A232;
  assign \new_[45689]_  = ~A236 & A235;
  assign \new_[45690]_  = \new_[45689]_  & \new_[45686]_ ;
  assign \new_[45693]_  = ~A266 & ~A265;
  assign \new_[45696]_  = ~A269 & A268;
  assign \new_[45697]_  = \new_[45696]_  & \new_[45693]_ ;
  assign \new_[45698]_  = \new_[45697]_  & \new_[45690]_ ;
  assign \new_[45701]_  = A168 & A169;
  assign \new_[45704]_  = A166 & ~A167;
  assign \new_[45705]_  = \new_[45704]_  & \new_[45701]_ ;
  assign \new_[45708]_  = A200 & ~A199;
  assign \new_[45711]_  = A202 & ~A201;
  assign \new_[45712]_  = \new_[45711]_  & \new_[45708]_ ;
  assign \new_[45713]_  = \new_[45712]_  & \new_[45705]_ ;
  assign \new_[45716]_  = A233 & A232;
  assign \new_[45719]_  = ~A236 & A235;
  assign \new_[45720]_  = \new_[45719]_  & \new_[45716]_ ;
  assign \new_[45723]_  = A299 & A298;
  assign \new_[45726]_  = ~A302 & A301;
  assign \new_[45727]_  = \new_[45726]_  & \new_[45723]_ ;
  assign \new_[45728]_  = \new_[45727]_  & \new_[45720]_ ;
  assign \new_[45731]_  = A168 & A169;
  assign \new_[45734]_  = A166 & ~A167;
  assign \new_[45735]_  = \new_[45734]_  & \new_[45731]_ ;
  assign \new_[45738]_  = A200 & ~A199;
  assign \new_[45741]_  = A202 & ~A201;
  assign \new_[45742]_  = \new_[45741]_  & \new_[45738]_ ;
  assign \new_[45743]_  = \new_[45742]_  & \new_[45735]_ ;
  assign \new_[45746]_  = A233 & A232;
  assign \new_[45749]_  = ~A236 & A235;
  assign \new_[45750]_  = \new_[45749]_  & \new_[45746]_ ;
  assign \new_[45753]_  = ~A299 & A298;
  assign \new_[45756]_  = A302 & ~A301;
  assign \new_[45757]_  = \new_[45756]_  & \new_[45753]_ ;
  assign \new_[45758]_  = \new_[45757]_  & \new_[45750]_ ;
  assign \new_[45761]_  = A168 & A169;
  assign \new_[45764]_  = A166 & ~A167;
  assign \new_[45765]_  = \new_[45764]_  & \new_[45761]_ ;
  assign \new_[45768]_  = A200 & ~A199;
  assign \new_[45771]_  = A202 & ~A201;
  assign \new_[45772]_  = \new_[45771]_  & \new_[45768]_ ;
  assign \new_[45773]_  = \new_[45772]_  & \new_[45765]_ ;
  assign \new_[45776]_  = A233 & A232;
  assign \new_[45779]_  = ~A236 & A235;
  assign \new_[45780]_  = \new_[45779]_  & \new_[45776]_ ;
  assign \new_[45783]_  = A299 & ~A298;
  assign \new_[45786]_  = A302 & ~A301;
  assign \new_[45787]_  = \new_[45786]_  & \new_[45783]_ ;
  assign \new_[45788]_  = \new_[45787]_  & \new_[45780]_ ;
  assign \new_[45791]_  = A168 & A169;
  assign \new_[45794]_  = A166 & ~A167;
  assign \new_[45795]_  = \new_[45794]_  & \new_[45791]_ ;
  assign \new_[45798]_  = A200 & ~A199;
  assign \new_[45801]_  = A202 & ~A201;
  assign \new_[45802]_  = \new_[45801]_  & \new_[45798]_ ;
  assign \new_[45803]_  = \new_[45802]_  & \new_[45795]_ ;
  assign \new_[45806]_  = A233 & A232;
  assign \new_[45809]_  = ~A236 & A235;
  assign \new_[45810]_  = \new_[45809]_  & \new_[45806]_ ;
  assign \new_[45813]_  = ~A299 & ~A298;
  assign \new_[45816]_  = ~A302 & A301;
  assign \new_[45817]_  = \new_[45816]_  & \new_[45813]_ ;
  assign \new_[45818]_  = \new_[45817]_  & \new_[45810]_ ;
  assign \new_[45821]_  = A168 & A169;
  assign \new_[45824]_  = A166 & ~A167;
  assign \new_[45825]_  = \new_[45824]_  & \new_[45821]_ ;
  assign \new_[45828]_  = A200 & ~A199;
  assign \new_[45831]_  = A202 & ~A201;
  assign \new_[45832]_  = \new_[45831]_  & \new_[45828]_ ;
  assign \new_[45833]_  = \new_[45832]_  & \new_[45825]_ ;
  assign \new_[45836]_  = A233 & A232;
  assign \new_[45839]_  = ~A236 & A235;
  assign \new_[45840]_  = \new_[45839]_  & \new_[45836]_ ;
  assign \new_[45843]_  = A266 & A265;
  assign \new_[45846]_  = ~A269 & A268;
  assign \new_[45847]_  = \new_[45846]_  & \new_[45843]_ ;
  assign \new_[45848]_  = \new_[45847]_  & \new_[45840]_ ;
  assign \new_[45851]_  = A168 & A169;
  assign \new_[45854]_  = A166 & ~A167;
  assign \new_[45855]_  = \new_[45854]_  & \new_[45851]_ ;
  assign \new_[45858]_  = A200 & ~A199;
  assign \new_[45861]_  = A202 & ~A201;
  assign \new_[45862]_  = \new_[45861]_  & \new_[45858]_ ;
  assign \new_[45863]_  = \new_[45862]_  & \new_[45855]_ ;
  assign \new_[45866]_  = A233 & A232;
  assign \new_[45869]_  = ~A236 & A235;
  assign \new_[45870]_  = \new_[45869]_  & \new_[45866]_ ;
  assign \new_[45873]_  = A266 & ~A265;
  assign \new_[45876]_  = A269 & ~A268;
  assign \new_[45877]_  = \new_[45876]_  & \new_[45873]_ ;
  assign \new_[45878]_  = \new_[45877]_  & \new_[45870]_ ;
  assign \new_[45881]_  = A168 & A169;
  assign \new_[45884]_  = A166 & ~A167;
  assign \new_[45885]_  = \new_[45884]_  & \new_[45881]_ ;
  assign \new_[45888]_  = A200 & ~A199;
  assign \new_[45891]_  = A202 & ~A201;
  assign \new_[45892]_  = \new_[45891]_  & \new_[45888]_ ;
  assign \new_[45893]_  = \new_[45892]_  & \new_[45885]_ ;
  assign \new_[45896]_  = A233 & A232;
  assign \new_[45899]_  = ~A236 & A235;
  assign \new_[45900]_  = \new_[45899]_  & \new_[45896]_ ;
  assign \new_[45903]_  = ~A266 & A265;
  assign \new_[45906]_  = A269 & ~A268;
  assign \new_[45907]_  = \new_[45906]_  & \new_[45903]_ ;
  assign \new_[45908]_  = \new_[45907]_  & \new_[45900]_ ;
  assign \new_[45911]_  = A168 & A169;
  assign \new_[45914]_  = A166 & ~A167;
  assign \new_[45915]_  = \new_[45914]_  & \new_[45911]_ ;
  assign \new_[45918]_  = A200 & ~A199;
  assign \new_[45921]_  = A202 & ~A201;
  assign \new_[45922]_  = \new_[45921]_  & \new_[45918]_ ;
  assign \new_[45923]_  = \new_[45922]_  & \new_[45915]_ ;
  assign \new_[45926]_  = A233 & A232;
  assign \new_[45929]_  = ~A236 & A235;
  assign \new_[45930]_  = \new_[45929]_  & \new_[45926]_ ;
  assign \new_[45933]_  = ~A266 & ~A265;
  assign \new_[45936]_  = ~A269 & A268;
  assign \new_[45937]_  = \new_[45936]_  & \new_[45933]_ ;
  assign \new_[45938]_  = \new_[45937]_  & \new_[45930]_ ;
  assign \new_[45941]_  = A168 & A169;
  assign \new_[45944]_  = A166 & ~A167;
  assign \new_[45945]_  = \new_[45944]_  & \new_[45941]_ ;
  assign \new_[45948]_  = A200 & ~A199;
  assign \new_[45951]_  = A202 & ~A201;
  assign \new_[45952]_  = \new_[45951]_  & \new_[45948]_ ;
  assign \new_[45953]_  = \new_[45952]_  & \new_[45945]_ ;
  assign \new_[45956]_  = A233 & ~A232;
  assign \new_[45959]_  = A236 & ~A235;
  assign \new_[45960]_  = \new_[45959]_  & \new_[45956]_ ;
  assign \new_[45963]_  = A299 & A298;
  assign \new_[45966]_  = ~A302 & A301;
  assign \new_[45967]_  = \new_[45966]_  & \new_[45963]_ ;
  assign \new_[45968]_  = \new_[45967]_  & \new_[45960]_ ;
  assign \new_[45971]_  = A168 & A169;
  assign \new_[45974]_  = A166 & ~A167;
  assign \new_[45975]_  = \new_[45974]_  & \new_[45971]_ ;
  assign \new_[45978]_  = A200 & ~A199;
  assign \new_[45981]_  = A202 & ~A201;
  assign \new_[45982]_  = \new_[45981]_  & \new_[45978]_ ;
  assign \new_[45983]_  = \new_[45982]_  & \new_[45975]_ ;
  assign \new_[45986]_  = A233 & ~A232;
  assign \new_[45989]_  = A236 & ~A235;
  assign \new_[45990]_  = \new_[45989]_  & \new_[45986]_ ;
  assign \new_[45993]_  = ~A299 & A298;
  assign \new_[45996]_  = A302 & ~A301;
  assign \new_[45997]_  = \new_[45996]_  & \new_[45993]_ ;
  assign \new_[45998]_  = \new_[45997]_  & \new_[45990]_ ;
  assign \new_[46001]_  = A168 & A169;
  assign \new_[46004]_  = A166 & ~A167;
  assign \new_[46005]_  = \new_[46004]_  & \new_[46001]_ ;
  assign \new_[46008]_  = A200 & ~A199;
  assign \new_[46011]_  = A202 & ~A201;
  assign \new_[46012]_  = \new_[46011]_  & \new_[46008]_ ;
  assign \new_[46013]_  = \new_[46012]_  & \new_[46005]_ ;
  assign \new_[46016]_  = A233 & ~A232;
  assign \new_[46019]_  = A236 & ~A235;
  assign \new_[46020]_  = \new_[46019]_  & \new_[46016]_ ;
  assign \new_[46023]_  = A299 & ~A298;
  assign \new_[46026]_  = A302 & ~A301;
  assign \new_[46027]_  = \new_[46026]_  & \new_[46023]_ ;
  assign \new_[46028]_  = \new_[46027]_  & \new_[46020]_ ;
  assign \new_[46031]_  = A168 & A169;
  assign \new_[46034]_  = A166 & ~A167;
  assign \new_[46035]_  = \new_[46034]_  & \new_[46031]_ ;
  assign \new_[46038]_  = A200 & ~A199;
  assign \new_[46041]_  = A202 & ~A201;
  assign \new_[46042]_  = \new_[46041]_  & \new_[46038]_ ;
  assign \new_[46043]_  = \new_[46042]_  & \new_[46035]_ ;
  assign \new_[46046]_  = A233 & ~A232;
  assign \new_[46049]_  = A236 & ~A235;
  assign \new_[46050]_  = \new_[46049]_  & \new_[46046]_ ;
  assign \new_[46053]_  = ~A299 & ~A298;
  assign \new_[46056]_  = ~A302 & A301;
  assign \new_[46057]_  = \new_[46056]_  & \new_[46053]_ ;
  assign \new_[46058]_  = \new_[46057]_  & \new_[46050]_ ;
  assign \new_[46061]_  = A168 & A169;
  assign \new_[46064]_  = A166 & ~A167;
  assign \new_[46065]_  = \new_[46064]_  & \new_[46061]_ ;
  assign \new_[46068]_  = A200 & ~A199;
  assign \new_[46071]_  = A202 & ~A201;
  assign \new_[46072]_  = \new_[46071]_  & \new_[46068]_ ;
  assign \new_[46073]_  = \new_[46072]_  & \new_[46065]_ ;
  assign \new_[46076]_  = A233 & ~A232;
  assign \new_[46079]_  = A236 & ~A235;
  assign \new_[46080]_  = \new_[46079]_  & \new_[46076]_ ;
  assign \new_[46083]_  = A266 & A265;
  assign \new_[46086]_  = ~A269 & A268;
  assign \new_[46087]_  = \new_[46086]_  & \new_[46083]_ ;
  assign \new_[46088]_  = \new_[46087]_  & \new_[46080]_ ;
  assign \new_[46091]_  = A168 & A169;
  assign \new_[46094]_  = A166 & ~A167;
  assign \new_[46095]_  = \new_[46094]_  & \new_[46091]_ ;
  assign \new_[46098]_  = A200 & ~A199;
  assign \new_[46101]_  = A202 & ~A201;
  assign \new_[46102]_  = \new_[46101]_  & \new_[46098]_ ;
  assign \new_[46103]_  = \new_[46102]_  & \new_[46095]_ ;
  assign \new_[46106]_  = A233 & ~A232;
  assign \new_[46109]_  = A236 & ~A235;
  assign \new_[46110]_  = \new_[46109]_  & \new_[46106]_ ;
  assign \new_[46113]_  = A266 & ~A265;
  assign \new_[46116]_  = A269 & ~A268;
  assign \new_[46117]_  = \new_[46116]_  & \new_[46113]_ ;
  assign \new_[46118]_  = \new_[46117]_  & \new_[46110]_ ;
  assign \new_[46121]_  = A168 & A169;
  assign \new_[46124]_  = A166 & ~A167;
  assign \new_[46125]_  = \new_[46124]_  & \new_[46121]_ ;
  assign \new_[46128]_  = A200 & ~A199;
  assign \new_[46131]_  = A202 & ~A201;
  assign \new_[46132]_  = \new_[46131]_  & \new_[46128]_ ;
  assign \new_[46133]_  = \new_[46132]_  & \new_[46125]_ ;
  assign \new_[46136]_  = A233 & ~A232;
  assign \new_[46139]_  = A236 & ~A235;
  assign \new_[46140]_  = \new_[46139]_  & \new_[46136]_ ;
  assign \new_[46143]_  = ~A266 & A265;
  assign \new_[46146]_  = A269 & ~A268;
  assign \new_[46147]_  = \new_[46146]_  & \new_[46143]_ ;
  assign \new_[46148]_  = \new_[46147]_  & \new_[46140]_ ;
  assign \new_[46151]_  = A168 & A169;
  assign \new_[46154]_  = A166 & ~A167;
  assign \new_[46155]_  = \new_[46154]_  & \new_[46151]_ ;
  assign \new_[46158]_  = A200 & ~A199;
  assign \new_[46161]_  = A202 & ~A201;
  assign \new_[46162]_  = \new_[46161]_  & \new_[46158]_ ;
  assign \new_[46163]_  = \new_[46162]_  & \new_[46155]_ ;
  assign \new_[46166]_  = A233 & ~A232;
  assign \new_[46169]_  = A236 & ~A235;
  assign \new_[46170]_  = \new_[46169]_  & \new_[46166]_ ;
  assign \new_[46173]_  = ~A266 & ~A265;
  assign \new_[46176]_  = ~A269 & A268;
  assign \new_[46177]_  = \new_[46176]_  & \new_[46173]_ ;
  assign \new_[46178]_  = \new_[46177]_  & \new_[46170]_ ;
  assign \new_[46181]_  = A168 & A169;
  assign \new_[46184]_  = A166 & ~A167;
  assign \new_[46185]_  = \new_[46184]_  & \new_[46181]_ ;
  assign \new_[46188]_  = A200 & ~A199;
  assign \new_[46191]_  = A202 & ~A201;
  assign \new_[46192]_  = \new_[46191]_  & \new_[46188]_ ;
  assign \new_[46193]_  = \new_[46192]_  & \new_[46185]_ ;
  assign \new_[46196]_  = ~A233 & A232;
  assign \new_[46199]_  = A236 & ~A235;
  assign \new_[46200]_  = \new_[46199]_  & \new_[46196]_ ;
  assign \new_[46203]_  = A299 & A298;
  assign \new_[46206]_  = ~A302 & A301;
  assign \new_[46207]_  = \new_[46206]_  & \new_[46203]_ ;
  assign \new_[46208]_  = \new_[46207]_  & \new_[46200]_ ;
  assign \new_[46211]_  = A168 & A169;
  assign \new_[46214]_  = A166 & ~A167;
  assign \new_[46215]_  = \new_[46214]_  & \new_[46211]_ ;
  assign \new_[46218]_  = A200 & ~A199;
  assign \new_[46221]_  = A202 & ~A201;
  assign \new_[46222]_  = \new_[46221]_  & \new_[46218]_ ;
  assign \new_[46223]_  = \new_[46222]_  & \new_[46215]_ ;
  assign \new_[46226]_  = ~A233 & A232;
  assign \new_[46229]_  = A236 & ~A235;
  assign \new_[46230]_  = \new_[46229]_  & \new_[46226]_ ;
  assign \new_[46233]_  = ~A299 & A298;
  assign \new_[46236]_  = A302 & ~A301;
  assign \new_[46237]_  = \new_[46236]_  & \new_[46233]_ ;
  assign \new_[46238]_  = \new_[46237]_  & \new_[46230]_ ;
  assign \new_[46241]_  = A168 & A169;
  assign \new_[46244]_  = A166 & ~A167;
  assign \new_[46245]_  = \new_[46244]_  & \new_[46241]_ ;
  assign \new_[46248]_  = A200 & ~A199;
  assign \new_[46251]_  = A202 & ~A201;
  assign \new_[46252]_  = \new_[46251]_  & \new_[46248]_ ;
  assign \new_[46253]_  = \new_[46252]_  & \new_[46245]_ ;
  assign \new_[46256]_  = ~A233 & A232;
  assign \new_[46259]_  = A236 & ~A235;
  assign \new_[46260]_  = \new_[46259]_  & \new_[46256]_ ;
  assign \new_[46263]_  = A299 & ~A298;
  assign \new_[46266]_  = A302 & ~A301;
  assign \new_[46267]_  = \new_[46266]_  & \new_[46263]_ ;
  assign \new_[46268]_  = \new_[46267]_  & \new_[46260]_ ;
  assign \new_[46271]_  = A168 & A169;
  assign \new_[46274]_  = A166 & ~A167;
  assign \new_[46275]_  = \new_[46274]_  & \new_[46271]_ ;
  assign \new_[46278]_  = A200 & ~A199;
  assign \new_[46281]_  = A202 & ~A201;
  assign \new_[46282]_  = \new_[46281]_  & \new_[46278]_ ;
  assign \new_[46283]_  = \new_[46282]_  & \new_[46275]_ ;
  assign \new_[46286]_  = ~A233 & A232;
  assign \new_[46289]_  = A236 & ~A235;
  assign \new_[46290]_  = \new_[46289]_  & \new_[46286]_ ;
  assign \new_[46293]_  = ~A299 & ~A298;
  assign \new_[46296]_  = ~A302 & A301;
  assign \new_[46297]_  = \new_[46296]_  & \new_[46293]_ ;
  assign \new_[46298]_  = \new_[46297]_  & \new_[46290]_ ;
  assign \new_[46301]_  = A168 & A169;
  assign \new_[46304]_  = A166 & ~A167;
  assign \new_[46305]_  = \new_[46304]_  & \new_[46301]_ ;
  assign \new_[46308]_  = A200 & ~A199;
  assign \new_[46311]_  = A202 & ~A201;
  assign \new_[46312]_  = \new_[46311]_  & \new_[46308]_ ;
  assign \new_[46313]_  = \new_[46312]_  & \new_[46305]_ ;
  assign \new_[46316]_  = ~A233 & A232;
  assign \new_[46319]_  = A236 & ~A235;
  assign \new_[46320]_  = \new_[46319]_  & \new_[46316]_ ;
  assign \new_[46323]_  = A266 & A265;
  assign \new_[46326]_  = ~A269 & A268;
  assign \new_[46327]_  = \new_[46326]_  & \new_[46323]_ ;
  assign \new_[46328]_  = \new_[46327]_  & \new_[46320]_ ;
  assign \new_[46331]_  = A168 & A169;
  assign \new_[46334]_  = A166 & ~A167;
  assign \new_[46335]_  = \new_[46334]_  & \new_[46331]_ ;
  assign \new_[46338]_  = A200 & ~A199;
  assign \new_[46341]_  = A202 & ~A201;
  assign \new_[46342]_  = \new_[46341]_  & \new_[46338]_ ;
  assign \new_[46343]_  = \new_[46342]_  & \new_[46335]_ ;
  assign \new_[46346]_  = ~A233 & A232;
  assign \new_[46349]_  = A236 & ~A235;
  assign \new_[46350]_  = \new_[46349]_  & \new_[46346]_ ;
  assign \new_[46353]_  = A266 & ~A265;
  assign \new_[46356]_  = A269 & ~A268;
  assign \new_[46357]_  = \new_[46356]_  & \new_[46353]_ ;
  assign \new_[46358]_  = \new_[46357]_  & \new_[46350]_ ;
  assign \new_[46361]_  = A168 & A169;
  assign \new_[46364]_  = A166 & ~A167;
  assign \new_[46365]_  = \new_[46364]_  & \new_[46361]_ ;
  assign \new_[46368]_  = A200 & ~A199;
  assign \new_[46371]_  = A202 & ~A201;
  assign \new_[46372]_  = \new_[46371]_  & \new_[46368]_ ;
  assign \new_[46373]_  = \new_[46372]_  & \new_[46365]_ ;
  assign \new_[46376]_  = ~A233 & A232;
  assign \new_[46379]_  = A236 & ~A235;
  assign \new_[46380]_  = \new_[46379]_  & \new_[46376]_ ;
  assign \new_[46383]_  = ~A266 & A265;
  assign \new_[46386]_  = A269 & ~A268;
  assign \new_[46387]_  = \new_[46386]_  & \new_[46383]_ ;
  assign \new_[46388]_  = \new_[46387]_  & \new_[46380]_ ;
  assign \new_[46391]_  = A168 & A169;
  assign \new_[46394]_  = A166 & ~A167;
  assign \new_[46395]_  = \new_[46394]_  & \new_[46391]_ ;
  assign \new_[46398]_  = A200 & ~A199;
  assign \new_[46401]_  = A202 & ~A201;
  assign \new_[46402]_  = \new_[46401]_  & \new_[46398]_ ;
  assign \new_[46403]_  = \new_[46402]_  & \new_[46395]_ ;
  assign \new_[46406]_  = ~A233 & A232;
  assign \new_[46409]_  = A236 & ~A235;
  assign \new_[46410]_  = \new_[46409]_  & \new_[46406]_ ;
  assign \new_[46413]_  = ~A266 & ~A265;
  assign \new_[46416]_  = ~A269 & A268;
  assign \new_[46417]_  = \new_[46416]_  & \new_[46413]_ ;
  assign \new_[46418]_  = \new_[46417]_  & \new_[46410]_ ;
  assign \new_[46421]_  = A168 & A169;
  assign \new_[46424]_  = A166 & ~A167;
  assign \new_[46425]_  = \new_[46424]_  & \new_[46421]_ ;
  assign \new_[46428]_  = A200 & ~A199;
  assign \new_[46431]_  = A202 & ~A201;
  assign \new_[46432]_  = \new_[46431]_  & \new_[46428]_ ;
  assign \new_[46433]_  = \new_[46432]_  & \new_[46425]_ ;
  assign \new_[46436]_  = ~A233 & ~A232;
  assign \new_[46439]_  = ~A236 & A235;
  assign \new_[46440]_  = \new_[46439]_  & \new_[46436]_ ;
  assign \new_[46443]_  = A299 & A298;
  assign \new_[46446]_  = ~A302 & A301;
  assign \new_[46447]_  = \new_[46446]_  & \new_[46443]_ ;
  assign \new_[46448]_  = \new_[46447]_  & \new_[46440]_ ;
  assign \new_[46451]_  = A168 & A169;
  assign \new_[46454]_  = A166 & ~A167;
  assign \new_[46455]_  = \new_[46454]_  & \new_[46451]_ ;
  assign \new_[46458]_  = A200 & ~A199;
  assign \new_[46461]_  = A202 & ~A201;
  assign \new_[46462]_  = \new_[46461]_  & \new_[46458]_ ;
  assign \new_[46463]_  = \new_[46462]_  & \new_[46455]_ ;
  assign \new_[46466]_  = ~A233 & ~A232;
  assign \new_[46469]_  = ~A236 & A235;
  assign \new_[46470]_  = \new_[46469]_  & \new_[46466]_ ;
  assign \new_[46473]_  = ~A299 & A298;
  assign \new_[46476]_  = A302 & ~A301;
  assign \new_[46477]_  = \new_[46476]_  & \new_[46473]_ ;
  assign \new_[46478]_  = \new_[46477]_  & \new_[46470]_ ;
  assign \new_[46481]_  = A168 & A169;
  assign \new_[46484]_  = A166 & ~A167;
  assign \new_[46485]_  = \new_[46484]_  & \new_[46481]_ ;
  assign \new_[46488]_  = A200 & ~A199;
  assign \new_[46491]_  = A202 & ~A201;
  assign \new_[46492]_  = \new_[46491]_  & \new_[46488]_ ;
  assign \new_[46493]_  = \new_[46492]_  & \new_[46485]_ ;
  assign \new_[46496]_  = ~A233 & ~A232;
  assign \new_[46499]_  = ~A236 & A235;
  assign \new_[46500]_  = \new_[46499]_  & \new_[46496]_ ;
  assign \new_[46503]_  = A299 & ~A298;
  assign \new_[46506]_  = A302 & ~A301;
  assign \new_[46507]_  = \new_[46506]_  & \new_[46503]_ ;
  assign \new_[46508]_  = \new_[46507]_  & \new_[46500]_ ;
  assign \new_[46511]_  = A168 & A169;
  assign \new_[46514]_  = A166 & ~A167;
  assign \new_[46515]_  = \new_[46514]_  & \new_[46511]_ ;
  assign \new_[46518]_  = A200 & ~A199;
  assign \new_[46521]_  = A202 & ~A201;
  assign \new_[46522]_  = \new_[46521]_  & \new_[46518]_ ;
  assign \new_[46523]_  = \new_[46522]_  & \new_[46515]_ ;
  assign \new_[46526]_  = ~A233 & ~A232;
  assign \new_[46529]_  = ~A236 & A235;
  assign \new_[46530]_  = \new_[46529]_  & \new_[46526]_ ;
  assign \new_[46533]_  = ~A299 & ~A298;
  assign \new_[46536]_  = ~A302 & A301;
  assign \new_[46537]_  = \new_[46536]_  & \new_[46533]_ ;
  assign \new_[46538]_  = \new_[46537]_  & \new_[46530]_ ;
  assign \new_[46541]_  = A168 & A169;
  assign \new_[46544]_  = A166 & ~A167;
  assign \new_[46545]_  = \new_[46544]_  & \new_[46541]_ ;
  assign \new_[46548]_  = A200 & ~A199;
  assign \new_[46551]_  = A202 & ~A201;
  assign \new_[46552]_  = \new_[46551]_  & \new_[46548]_ ;
  assign \new_[46553]_  = \new_[46552]_  & \new_[46545]_ ;
  assign \new_[46556]_  = ~A233 & ~A232;
  assign \new_[46559]_  = ~A236 & A235;
  assign \new_[46560]_  = \new_[46559]_  & \new_[46556]_ ;
  assign \new_[46563]_  = A266 & A265;
  assign \new_[46566]_  = ~A269 & A268;
  assign \new_[46567]_  = \new_[46566]_  & \new_[46563]_ ;
  assign \new_[46568]_  = \new_[46567]_  & \new_[46560]_ ;
  assign \new_[46571]_  = A168 & A169;
  assign \new_[46574]_  = A166 & ~A167;
  assign \new_[46575]_  = \new_[46574]_  & \new_[46571]_ ;
  assign \new_[46578]_  = A200 & ~A199;
  assign \new_[46581]_  = A202 & ~A201;
  assign \new_[46582]_  = \new_[46581]_  & \new_[46578]_ ;
  assign \new_[46583]_  = \new_[46582]_  & \new_[46575]_ ;
  assign \new_[46586]_  = ~A233 & ~A232;
  assign \new_[46589]_  = ~A236 & A235;
  assign \new_[46590]_  = \new_[46589]_  & \new_[46586]_ ;
  assign \new_[46593]_  = A266 & ~A265;
  assign \new_[46596]_  = A269 & ~A268;
  assign \new_[46597]_  = \new_[46596]_  & \new_[46593]_ ;
  assign \new_[46598]_  = \new_[46597]_  & \new_[46590]_ ;
  assign \new_[46601]_  = A168 & A169;
  assign \new_[46604]_  = A166 & ~A167;
  assign \new_[46605]_  = \new_[46604]_  & \new_[46601]_ ;
  assign \new_[46608]_  = A200 & ~A199;
  assign \new_[46611]_  = A202 & ~A201;
  assign \new_[46612]_  = \new_[46611]_  & \new_[46608]_ ;
  assign \new_[46613]_  = \new_[46612]_  & \new_[46605]_ ;
  assign \new_[46616]_  = ~A233 & ~A232;
  assign \new_[46619]_  = ~A236 & A235;
  assign \new_[46620]_  = \new_[46619]_  & \new_[46616]_ ;
  assign \new_[46623]_  = ~A266 & A265;
  assign \new_[46626]_  = A269 & ~A268;
  assign \new_[46627]_  = \new_[46626]_  & \new_[46623]_ ;
  assign \new_[46628]_  = \new_[46627]_  & \new_[46620]_ ;
  assign \new_[46631]_  = A168 & A169;
  assign \new_[46634]_  = A166 & ~A167;
  assign \new_[46635]_  = \new_[46634]_  & \new_[46631]_ ;
  assign \new_[46638]_  = A200 & ~A199;
  assign \new_[46641]_  = A202 & ~A201;
  assign \new_[46642]_  = \new_[46641]_  & \new_[46638]_ ;
  assign \new_[46643]_  = \new_[46642]_  & \new_[46635]_ ;
  assign \new_[46646]_  = ~A233 & ~A232;
  assign \new_[46649]_  = ~A236 & A235;
  assign \new_[46650]_  = \new_[46649]_  & \new_[46646]_ ;
  assign \new_[46653]_  = ~A266 & ~A265;
  assign \new_[46656]_  = ~A269 & A268;
  assign \new_[46657]_  = \new_[46656]_  & \new_[46653]_ ;
  assign \new_[46658]_  = \new_[46657]_  & \new_[46650]_ ;
  assign \new_[46661]_  = A168 & A169;
  assign \new_[46664]_  = A166 & ~A167;
  assign \new_[46665]_  = \new_[46664]_  & \new_[46661]_ ;
  assign \new_[46668]_  = A200 & ~A199;
  assign \new_[46671]_  = ~A203 & ~A201;
  assign \new_[46672]_  = \new_[46671]_  & \new_[46668]_ ;
  assign \new_[46673]_  = \new_[46672]_  & \new_[46665]_ ;
  assign \new_[46676]_  = A233 & A232;
  assign \new_[46679]_  = ~A236 & A235;
  assign \new_[46680]_  = \new_[46679]_  & \new_[46676]_ ;
  assign \new_[46683]_  = A299 & A298;
  assign \new_[46686]_  = ~A302 & A301;
  assign \new_[46687]_  = \new_[46686]_  & \new_[46683]_ ;
  assign \new_[46688]_  = \new_[46687]_  & \new_[46680]_ ;
  assign \new_[46691]_  = A168 & A169;
  assign \new_[46694]_  = A166 & ~A167;
  assign \new_[46695]_  = \new_[46694]_  & \new_[46691]_ ;
  assign \new_[46698]_  = A200 & ~A199;
  assign \new_[46701]_  = ~A203 & ~A201;
  assign \new_[46702]_  = \new_[46701]_  & \new_[46698]_ ;
  assign \new_[46703]_  = \new_[46702]_  & \new_[46695]_ ;
  assign \new_[46706]_  = A233 & A232;
  assign \new_[46709]_  = ~A236 & A235;
  assign \new_[46710]_  = \new_[46709]_  & \new_[46706]_ ;
  assign \new_[46713]_  = ~A299 & A298;
  assign \new_[46716]_  = A302 & ~A301;
  assign \new_[46717]_  = \new_[46716]_  & \new_[46713]_ ;
  assign \new_[46718]_  = \new_[46717]_  & \new_[46710]_ ;
  assign \new_[46721]_  = A168 & A169;
  assign \new_[46724]_  = A166 & ~A167;
  assign \new_[46725]_  = \new_[46724]_  & \new_[46721]_ ;
  assign \new_[46728]_  = A200 & ~A199;
  assign \new_[46731]_  = ~A203 & ~A201;
  assign \new_[46732]_  = \new_[46731]_  & \new_[46728]_ ;
  assign \new_[46733]_  = \new_[46732]_  & \new_[46725]_ ;
  assign \new_[46736]_  = A233 & A232;
  assign \new_[46739]_  = ~A236 & A235;
  assign \new_[46740]_  = \new_[46739]_  & \new_[46736]_ ;
  assign \new_[46743]_  = A299 & ~A298;
  assign \new_[46746]_  = A302 & ~A301;
  assign \new_[46747]_  = \new_[46746]_  & \new_[46743]_ ;
  assign \new_[46748]_  = \new_[46747]_  & \new_[46740]_ ;
  assign \new_[46751]_  = A168 & A169;
  assign \new_[46754]_  = A166 & ~A167;
  assign \new_[46755]_  = \new_[46754]_  & \new_[46751]_ ;
  assign \new_[46758]_  = A200 & ~A199;
  assign \new_[46761]_  = ~A203 & ~A201;
  assign \new_[46762]_  = \new_[46761]_  & \new_[46758]_ ;
  assign \new_[46763]_  = \new_[46762]_  & \new_[46755]_ ;
  assign \new_[46766]_  = A233 & A232;
  assign \new_[46769]_  = ~A236 & A235;
  assign \new_[46770]_  = \new_[46769]_  & \new_[46766]_ ;
  assign \new_[46773]_  = ~A299 & ~A298;
  assign \new_[46776]_  = ~A302 & A301;
  assign \new_[46777]_  = \new_[46776]_  & \new_[46773]_ ;
  assign \new_[46778]_  = \new_[46777]_  & \new_[46770]_ ;
  assign \new_[46781]_  = A168 & A169;
  assign \new_[46784]_  = A166 & ~A167;
  assign \new_[46785]_  = \new_[46784]_  & \new_[46781]_ ;
  assign \new_[46788]_  = A200 & ~A199;
  assign \new_[46791]_  = ~A203 & ~A201;
  assign \new_[46792]_  = \new_[46791]_  & \new_[46788]_ ;
  assign \new_[46793]_  = \new_[46792]_  & \new_[46785]_ ;
  assign \new_[46796]_  = A233 & A232;
  assign \new_[46799]_  = ~A236 & A235;
  assign \new_[46800]_  = \new_[46799]_  & \new_[46796]_ ;
  assign \new_[46803]_  = A266 & A265;
  assign \new_[46806]_  = ~A269 & A268;
  assign \new_[46807]_  = \new_[46806]_  & \new_[46803]_ ;
  assign \new_[46808]_  = \new_[46807]_  & \new_[46800]_ ;
  assign \new_[46811]_  = A168 & A169;
  assign \new_[46814]_  = A166 & ~A167;
  assign \new_[46815]_  = \new_[46814]_  & \new_[46811]_ ;
  assign \new_[46818]_  = A200 & ~A199;
  assign \new_[46821]_  = ~A203 & ~A201;
  assign \new_[46822]_  = \new_[46821]_  & \new_[46818]_ ;
  assign \new_[46823]_  = \new_[46822]_  & \new_[46815]_ ;
  assign \new_[46826]_  = A233 & A232;
  assign \new_[46829]_  = ~A236 & A235;
  assign \new_[46830]_  = \new_[46829]_  & \new_[46826]_ ;
  assign \new_[46833]_  = A266 & ~A265;
  assign \new_[46836]_  = A269 & ~A268;
  assign \new_[46837]_  = \new_[46836]_  & \new_[46833]_ ;
  assign \new_[46838]_  = \new_[46837]_  & \new_[46830]_ ;
  assign \new_[46841]_  = A168 & A169;
  assign \new_[46844]_  = A166 & ~A167;
  assign \new_[46845]_  = \new_[46844]_  & \new_[46841]_ ;
  assign \new_[46848]_  = A200 & ~A199;
  assign \new_[46851]_  = ~A203 & ~A201;
  assign \new_[46852]_  = \new_[46851]_  & \new_[46848]_ ;
  assign \new_[46853]_  = \new_[46852]_  & \new_[46845]_ ;
  assign \new_[46856]_  = A233 & A232;
  assign \new_[46859]_  = ~A236 & A235;
  assign \new_[46860]_  = \new_[46859]_  & \new_[46856]_ ;
  assign \new_[46863]_  = ~A266 & A265;
  assign \new_[46866]_  = A269 & ~A268;
  assign \new_[46867]_  = \new_[46866]_  & \new_[46863]_ ;
  assign \new_[46868]_  = \new_[46867]_  & \new_[46860]_ ;
  assign \new_[46871]_  = A168 & A169;
  assign \new_[46874]_  = A166 & ~A167;
  assign \new_[46875]_  = \new_[46874]_  & \new_[46871]_ ;
  assign \new_[46878]_  = A200 & ~A199;
  assign \new_[46881]_  = ~A203 & ~A201;
  assign \new_[46882]_  = \new_[46881]_  & \new_[46878]_ ;
  assign \new_[46883]_  = \new_[46882]_  & \new_[46875]_ ;
  assign \new_[46886]_  = A233 & A232;
  assign \new_[46889]_  = ~A236 & A235;
  assign \new_[46890]_  = \new_[46889]_  & \new_[46886]_ ;
  assign \new_[46893]_  = ~A266 & ~A265;
  assign \new_[46896]_  = ~A269 & A268;
  assign \new_[46897]_  = \new_[46896]_  & \new_[46893]_ ;
  assign \new_[46898]_  = \new_[46897]_  & \new_[46890]_ ;
  assign \new_[46901]_  = A168 & A169;
  assign \new_[46904]_  = A166 & ~A167;
  assign \new_[46905]_  = \new_[46904]_  & \new_[46901]_ ;
  assign \new_[46908]_  = A200 & ~A199;
  assign \new_[46911]_  = ~A203 & ~A201;
  assign \new_[46912]_  = \new_[46911]_  & \new_[46908]_ ;
  assign \new_[46913]_  = \new_[46912]_  & \new_[46905]_ ;
  assign \new_[46916]_  = A233 & ~A232;
  assign \new_[46919]_  = A236 & ~A235;
  assign \new_[46920]_  = \new_[46919]_  & \new_[46916]_ ;
  assign \new_[46923]_  = A299 & A298;
  assign \new_[46926]_  = ~A302 & A301;
  assign \new_[46927]_  = \new_[46926]_  & \new_[46923]_ ;
  assign \new_[46928]_  = \new_[46927]_  & \new_[46920]_ ;
  assign \new_[46931]_  = A168 & A169;
  assign \new_[46934]_  = A166 & ~A167;
  assign \new_[46935]_  = \new_[46934]_  & \new_[46931]_ ;
  assign \new_[46938]_  = A200 & ~A199;
  assign \new_[46941]_  = ~A203 & ~A201;
  assign \new_[46942]_  = \new_[46941]_  & \new_[46938]_ ;
  assign \new_[46943]_  = \new_[46942]_  & \new_[46935]_ ;
  assign \new_[46946]_  = A233 & ~A232;
  assign \new_[46949]_  = A236 & ~A235;
  assign \new_[46950]_  = \new_[46949]_  & \new_[46946]_ ;
  assign \new_[46953]_  = ~A299 & A298;
  assign \new_[46956]_  = A302 & ~A301;
  assign \new_[46957]_  = \new_[46956]_  & \new_[46953]_ ;
  assign \new_[46958]_  = \new_[46957]_  & \new_[46950]_ ;
  assign \new_[46961]_  = A168 & A169;
  assign \new_[46964]_  = A166 & ~A167;
  assign \new_[46965]_  = \new_[46964]_  & \new_[46961]_ ;
  assign \new_[46968]_  = A200 & ~A199;
  assign \new_[46971]_  = ~A203 & ~A201;
  assign \new_[46972]_  = \new_[46971]_  & \new_[46968]_ ;
  assign \new_[46973]_  = \new_[46972]_  & \new_[46965]_ ;
  assign \new_[46976]_  = A233 & ~A232;
  assign \new_[46979]_  = A236 & ~A235;
  assign \new_[46980]_  = \new_[46979]_  & \new_[46976]_ ;
  assign \new_[46983]_  = A299 & ~A298;
  assign \new_[46986]_  = A302 & ~A301;
  assign \new_[46987]_  = \new_[46986]_  & \new_[46983]_ ;
  assign \new_[46988]_  = \new_[46987]_  & \new_[46980]_ ;
  assign \new_[46991]_  = A168 & A169;
  assign \new_[46994]_  = A166 & ~A167;
  assign \new_[46995]_  = \new_[46994]_  & \new_[46991]_ ;
  assign \new_[46998]_  = A200 & ~A199;
  assign \new_[47001]_  = ~A203 & ~A201;
  assign \new_[47002]_  = \new_[47001]_  & \new_[46998]_ ;
  assign \new_[47003]_  = \new_[47002]_  & \new_[46995]_ ;
  assign \new_[47006]_  = A233 & ~A232;
  assign \new_[47009]_  = A236 & ~A235;
  assign \new_[47010]_  = \new_[47009]_  & \new_[47006]_ ;
  assign \new_[47013]_  = ~A299 & ~A298;
  assign \new_[47016]_  = ~A302 & A301;
  assign \new_[47017]_  = \new_[47016]_  & \new_[47013]_ ;
  assign \new_[47018]_  = \new_[47017]_  & \new_[47010]_ ;
  assign \new_[47021]_  = A168 & A169;
  assign \new_[47024]_  = A166 & ~A167;
  assign \new_[47025]_  = \new_[47024]_  & \new_[47021]_ ;
  assign \new_[47028]_  = A200 & ~A199;
  assign \new_[47031]_  = ~A203 & ~A201;
  assign \new_[47032]_  = \new_[47031]_  & \new_[47028]_ ;
  assign \new_[47033]_  = \new_[47032]_  & \new_[47025]_ ;
  assign \new_[47036]_  = A233 & ~A232;
  assign \new_[47039]_  = A236 & ~A235;
  assign \new_[47040]_  = \new_[47039]_  & \new_[47036]_ ;
  assign \new_[47043]_  = A266 & A265;
  assign \new_[47046]_  = ~A269 & A268;
  assign \new_[47047]_  = \new_[47046]_  & \new_[47043]_ ;
  assign \new_[47048]_  = \new_[47047]_  & \new_[47040]_ ;
  assign \new_[47051]_  = A168 & A169;
  assign \new_[47054]_  = A166 & ~A167;
  assign \new_[47055]_  = \new_[47054]_  & \new_[47051]_ ;
  assign \new_[47058]_  = A200 & ~A199;
  assign \new_[47061]_  = ~A203 & ~A201;
  assign \new_[47062]_  = \new_[47061]_  & \new_[47058]_ ;
  assign \new_[47063]_  = \new_[47062]_  & \new_[47055]_ ;
  assign \new_[47066]_  = A233 & ~A232;
  assign \new_[47069]_  = A236 & ~A235;
  assign \new_[47070]_  = \new_[47069]_  & \new_[47066]_ ;
  assign \new_[47073]_  = A266 & ~A265;
  assign \new_[47076]_  = A269 & ~A268;
  assign \new_[47077]_  = \new_[47076]_  & \new_[47073]_ ;
  assign \new_[47078]_  = \new_[47077]_  & \new_[47070]_ ;
  assign \new_[47081]_  = A168 & A169;
  assign \new_[47084]_  = A166 & ~A167;
  assign \new_[47085]_  = \new_[47084]_  & \new_[47081]_ ;
  assign \new_[47088]_  = A200 & ~A199;
  assign \new_[47091]_  = ~A203 & ~A201;
  assign \new_[47092]_  = \new_[47091]_  & \new_[47088]_ ;
  assign \new_[47093]_  = \new_[47092]_  & \new_[47085]_ ;
  assign \new_[47096]_  = A233 & ~A232;
  assign \new_[47099]_  = A236 & ~A235;
  assign \new_[47100]_  = \new_[47099]_  & \new_[47096]_ ;
  assign \new_[47103]_  = ~A266 & A265;
  assign \new_[47106]_  = A269 & ~A268;
  assign \new_[47107]_  = \new_[47106]_  & \new_[47103]_ ;
  assign \new_[47108]_  = \new_[47107]_  & \new_[47100]_ ;
  assign \new_[47111]_  = A168 & A169;
  assign \new_[47114]_  = A166 & ~A167;
  assign \new_[47115]_  = \new_[47114]_  & \new_[47111]_ ;
  assign \new_[47118]_  = A200 & ~A199;
  assign \new_[47121]_  = ~A203 & ~A201;
  assign \new_[47122]_  = \new_[47121]_  & \new_[47118]_ ;
  assign \new_[47123]_  = \new_[47122]_  & \new_[47115]_ ;
  assign \new_[47126]_  = A233 & ~A232;
  assign \new_[47129]_  = A236 & ~A235;
  assign \new_[47130]_  = \new_[47129]_  & \new_[47126]_ ;
  assign \new_[47133]_  = ~A266 & ~A265;
  assign \new_[47136]_  = ~A269 & A268;
  assign \new_[47137]_  = \new_[47136]_  & \new_[47133]_ ;
  assign \new_[47138]_  = \new_[47137]_  & \new_[47130]_ ;
  assign \new_[47141]_  = A168 & A169;
  assign \new_[47144]_  = A166 & ~A167;
  assign \new_[47145]_  = \new_[47144]_  & \new_[47141]_ ;
  assign \new_[47148]_  = A200 & ~A199;
  assign \new_[47151]_  = ~A203 & ~A201;
  assign \new_[47152]_  = \new_[47151]_  & \new_[47148]_ ;
  assign \new_[47153]_  = \new_[47152]_  & \new_[47145]_ ;
  assign \new_[47156]_  = ~A233 & A232;
  assign \new_[47159]_  = A236 & ~A235;
  assign \new_[47160]_  = \new_[47159]_  & \new_[47156]_ ;
  assign \new_[47163]_  = A299 & A298;
  assign \new_[47166]_  = ~A302 & A301;
  assign \new_[47167]_  = \new_[47166]_  & \new_[47163]_ ;
  assign \new_[47168]_  = \new_[47167]_  & \new_[47160]_ ;
  assign \new_[47171]_  = A168 & A169;
  assign \new_[47174]_  = A166 & ~A167;
  assign \new_[47175]_  = \new_[47174]_  & \new_[47171]_ ;
  assign \new_[47178]_  = A200 & ~A199;
  assign \new_[47181]_  = ~A203 & ~A201;
  assign \new_[47182]_  = \new_[47181]_  & \new_[47178]_ ;
  assign \new_[47183]_  = \new_[47182]_  & \new_[47175]_ ;
  assign \new_[47186]_  = ~A233 & A232;
  assign \new_[47189]_  = A236 & ~A235;
  assign \new_[47190]_  = \new_[47189]_  & \new_[47186]_ ;
  assign \new_[47193]_  = ~A299 & A298;
  assign \new_[47196]_  = A302 & ~A301;
  assign \new_[47197]_  = \new_[47196]_  & \new_[47193]_ ;
  assign \new_[47198]_  = \new_[47197]_  & \new_[47190]_ ;
  assign \new_[47201]_  = A168 & A169;
  assign \new_[47204]_  = A166 & ~A167;
  assign \new_[47205]_  = \new_[47204]_  & \new_[47201]_ ;
  assign \new_[47208]_  = A200 & ~A199;
  assign \new_[47211]_  = ~A203 & ~A201;
  assign \new_[47212]_  = \new_[47211]_  & \new_[47208]_ ;
  assign \new_[47213]_  = \new_[47212]_  & \new_[47205]_ ;
  assign \new_[47216]_  = ~A233 & A232;
  assign \new_[47219]_  = A236 & ~A235;
  assign \new_[47220]_  = \new_[47219]_  & \new_[47216]_ ;
  assign \new_[47223]_  = A299 & ~A298;
  assign \new_[47226]_  = A302 & ~A301;
  assign \new_[47227]_  = \new_[47226]_  & \new_[47223]_ ;
  assign \new_[47228]_  = \new_[47227]_  & \new_[47220]_ ;
  assign \new_[47231]_  = A168 & A169;
  assign \new_[47234]_  = A166 & ~A167;
  assign \new_[47235]_  = \new_[47234]_  & \new_[47231]_ ;
  assign \new_[47238]_  = A200 & ~A199;
  assign \new_[47241]_  = ~A203 & ~A201;
  assign \new_[47242]_  = \new_[47241]_  & \new_[47238]_ ;
  assign \new_[47243]_  = \new_[47242]_  & \new_[47235]_ ;
  assign \new_[47246]_  = ~A233 & A232;
  assign \new_[47249]_  = A236 & ~A235;
  assign \new_[47250]_  = \new_[47249]_  & \new_[47246]_ ;
  assign \new_[47253]_  = ~A299 & ~A298;
  assign \new_[47256]_  = ~A302 & A301;
  assign \new_[47257]_  = \new_[47256]_  & \new_[47253]_ ;
  assign \new_[47258]_  = \new_[47257]_  & \new_[47250]_ ;
  assign \new_[47261]_  = A168 & A169;
  assign \new_[47264]_  = A166 & ~A167;
  assign \new_[47265]_  = \new_[47264]_  & \new_[47261]_ ;
  assign \new_[47268]_  = A200 & ~A199;
  assign \new_[47271]_  = ~A203 & ~A201;
  assign \new_[47272]_  = \new_[47271]_  & \new_[47268]_ ;
  assign \new_[47273]_  = \new_[47272]_  & \new_[47265]_ ;
  assign \new_[47276]_  = ~A233 & A232;
  assign \new_[47279]_  = A236 & ~A235;
  assign \new_[47280]_  = \new_[47279]_  & \new_[47276]_ ;
  assign \new_[47283]_  = A266 & A265;
  assign \new_[47286]_  = ~A269 & A268;
  assign \new_[47287]_  = \new_[47286]_  & \new_[47283]_ ;
  assign \new_[47288]_  = \new_[47287]_  & \new_[47280]_ ;
  assign \new_[47291]_  = A168 & A169;
  assign \new_[47294]_  = A166 & ~A167;
  assign \new_[47295]_  = \new_[47294]_  & \new_[47291]_ ;
  assign \new_[47298]_  = A200 & ~A199;
  assign \new_[47301]_  = ~A203 & ~A201;
  assign \new_[47302]_  = \new_[47301]_  & \new_[47298]_ ;
  assign \new_[47303]_  = \new_[47302]_  & \new_[47295]_ ;
  assign \new_[47306]_  = ~A233 & A232;
  assign \new_[47309]_  = A236 & ~A235;
  assign \new_[47310]_  = \new_[47309]_  & \new_[47306]_ ;
  assign \new_[47313]_  = A266 & ~A265;
  assign \new_[47316]_  = A269 & ~A268;
  assign \new_[47317]_  = \new_[47316]_  & \new_[47313]_ ;
  assign \new_[47318]_  = \new_[47317]_  & \new_[47310]_ ;
  assign \new_[47321]_  = A168 & A169;
  assign \new_[47324]_  = A166 & ~A167;
  assign \new_[47325]_  = \new_[47324]_  & \new_[47321]_ ;
  assign \new_[47328]_  = A200 & ~A199;
  assign \new_[47331]_  = ~A203 & ~A201;
  assign \new_[47332]_  = \new_[47331]_  & \new_[47328]_ ;
  assign \new_[47333]_  = \new_[47332]_  & \new_[47325]_ ;
  assign \new_[47336]_  = ~A233 & A232;
  assign \new_[47339]_  = A236 & ~A235;
  assign \new_[47340]_  = \new_[47339]_  & \new_[47336]_ ;
  assign \new_[47343]_  = ~A266 & A265;
  assign \new_[47346]_  = A269 & ~A268;
  assign \new_[47347]_  = \new_[47346]_  & \new_[47343]_ ;
  assign \new_[47348]_  = \new_[47347]_  & \new_[47340]_ ;
  assign \new_[47351]_  = A168 & A169;
  assign \new_[47354]_  = A166 & ~A167;
  assign \new_[47355]_  = \new_[47354]_  & \new_[47351]_ ;
  assign \new_[47358]_  = A200 & ~A199;
  assign \new_[47361]_  = ~A203 & ~A201;
  assign \new_[47362]_  = \new_[47361]_  & \new_[47358]_ ;
  assign \new_[47363]_  = \new_[47362]_  & \new_[47355]_ ;
  assign \new_[47366]_  = ~A233 & A232;
  assign \new_[47369]_  = A236 & ~A235;
  assign \new_[47370]_  = \new_[47369]_  & \new_[47366]_ ;
  assign \new_[47373]_  = ~A266 & ~A265;
  assign \new_[47376]_  = ~A269 & A268;
  assign \new_[47377]_  = \new_[47376]_  & \new_[47373]_ ;
  assign \new_[47378]_  = \new_[47377]_  & \new_[47370]_ ;
  assign \new_[47381]_  = A168 & A169;
  assign \new_[47384]_  = A166 & ~A167;
  assign \new_[47385]_  = \new_[47384]_  & \new_[47381]_ ;
  assign \new_[47388]_  = A200 & ~A199;
  assign \new_[47391]_  = ~A203 & ~A201;
  assign \new_[47392]_  = \new_[47391]_  & \new_[47388]_ ;
  assign \new_[47393]_  = \new_[47392]_  & \new_[47385]_ ;
  assign \new_[47396]_  = ~A233 & ~A232;
  assign \new_[47399]_  = ~A236 & A235;
  assign \new_[47400]_  = \new_[47399]_  & \new_[47396]_ ;
  assign \new_[47403]_  = A299 & A298;
  assign \new_[47406]_  = ~A302 & A301;
  assign \new_[47407]_  = \new_[47406]_  & \new_[47403]_ ;
  assign \new_[47408]_  = \new_[47407]_  & \new_[47400]_ ;
  assign \new_[47411]_  = A168 & A169;
  assign \new_[47414]_  = A166 & ~A167;
  assign \new_[47415]_  = \new_[47414]_  & \new_[47411]_ ;
  assign \new_[47418]_  = A200 & ~A199;
  assign \new_[47421]_  = ~A203 & ~A201;
  assign \new_[47422]_  = \new_[47421]_  & \new_[47418]_ ;
  assign \new_[47423]_  = \new_[47422]_  & \new_[47415]_ ;
  assign \new_[47426]_  = ~A233 & ~A232;
  assign \new_[47429]_  = ~A236 & A235;
  assign \new_[47430]_  = \new_[47429]_  & \new_[47426]_ ;
  assign \new_[47433]_  = ~A299 & A298;
  assign \new_[47436]_  = A302 & ~A301;
  assign \new_[47437]_  = \new_[47436]_  & \new_[47433]_ ;
  assign \new_[47438]_  = \new_[47437]_  & \new_[47430]_ ;
  assign \new_[47441]_  = A168 & A169;
  assign \new_[47444]_  = A166 & ~A167;
  assign \new_[47445]_  = \new_[47444]_  & \new_[47441]_ ;
  assign \new_[47448]_  = A200 & ~A199;
  assign \new_[47451]_  = ~A203 & ~A201;
  assign \new_[47452]_  = \new_[47451]_  & \new_[47448]_ ;
  assign \new_[47453]_  = \new_[47452]_  & \new_[47445]_ ;
  assign \new_[47456]_  = ~A233 & ~A232;
  assign \new_[47459]_  = ~A236 & A235;
  assign \new_[47460]_  = \new_[47459]_  & \new_[47456]_ ;
  assign \new_[47463]_  = A299 & ~A298;
  assign \new_[47466]_  = A302 & ~A301;
  assign \new_[47467]_  = \new_[47466]_  & \new_[47463]_ ;
  assign \new_[47468]_  = \new_[47467]_  & \new_[47460]_ ;
  assign \new_[47471]_  = A168 & A169;
  assign \new_[47474]_  = A166 & ~A167;
  assign \new_[47475]_  = \new_[47474]_  & \new_[47471]_ ;
  assign \new_[47478]_  = A200 & ~A199;
  assign \new_[47481]_  = ~A203 & ~A201;
  assign \new_[47482]_  = \new_[47481]_  & \new_[47478]_ ;
  assign \new_[47483]_  = \new_[47482]_  & \new_[47475]_ ;
  assign \new_[47486]_  = ~A233 & ~A232;
  assign \new_[47489]_  = ~A236 & A235;
  assign \new_[47490]_  = \new_[47489]_  & \new_[47486]_ ;
  assign \new_[47493]_  = ~A299 & ~A298;
  assign \new_[47496]_  = ~A302 & A301;
  assign \new_[47497]_  = \new_[47496]_  & \new_[47493]_ ;
  assign \new_[47498]_  = \new_[47497]_  & \new_[47490]_ ;
  assign \new_[47501]_  = A168 & A169;
  assign \new_[47504]_  = A166 & ~A167;
  assign \new_[47505]_  = \new_[47504]_  & \new_[47501]_ ;
  assign \new_[47508]_  = A200 & ~A199;
  assign \new_[47511]_  = ~A203 & ~A201;
  assign \new_[47512]_  = \new_[47511]_  & \new_[47508]_ ;
  assign \new_[47513]_  = \new_[47512]_  & \new_[47505]_ ;
  assign \new_[47516]_  = ~A233 & ~A232;
  assign \new_[47519]_  = ~A236 & A235;
  assign \new_[47520]_  = \new_[47519]_  & \new_[47516]_ ;
  assign \new_[47523]_  = A266 & A265;
  assign \new_[47526]_  = ~A269 & A268;
  assign \new_[47527]_  = \new_[47526]_  & \new_[47523]_ ;
  assign \new_[47528]_  = \new_[47527]_  & \new_[47520]_ ;
  assign \new_[47531]_  = A168 & A169;
  assign \new_[47534]_  = A166 & ~A167;
  assign \new_[47535]_  = \new_[47534]_  & \new_[47531]_ ;
  assign \new_[47538]_  = A200 & ~A199;
  assign \new_[47541]_  = ~A203 & ~A201;
  assign \new_[47542]_  = \new_[47541]_  & \new_[47538]_ ;
  assign \new_[47543]_  = \new_[47542]_  & \new_[47535]_ ;
  assign \new_[47546]_  = ~A233 & ~A232;
  assign \new_[47549]_  = ~A236 & A235;
  assign \new_[47550]_  = \new_[47549]_  & \new_[47546]_ ;
  assign \new_[47553]_  = A266 & ~A265;
  assign \new_[47556]_  = A269 & ~A268;
  assign \new_[47557]_  = \new_[47556]_  & \new_[47553]_ ;
  assign \new_[47558]_  = \new_[47557]_  & \new_[47550]_ ;
  assign \new_[47561]_  = A168 & A169;
  assign \new_[47564]_  = A166 & ~A167;
  assign \new_[47565]_  = \new_[47564]_  & \new_[47561]_ ;
  assign \new_[47568]_  = A200 & ~A199;
  assign \new_[47571]_  = ~A203 & ~A201;
  assign \new_[47572]_  = \new_[47571]_  & \new_[47568]_ ;
  assign \new_[47573]_  = \new_[47572]_  & \new_[47565]_ ;
  assign \new_[47576]_  = ~A233 & ~A232;
  assign \new_[47579]_  = ~A236 & A235;
  assign \new_[47580]_  = \new_[47579]_  & \new_[47576]_ ;
  assign \new_[47583]_  = ~A266 & A265;
  assign \new_[47586]_  = A269 & ~A268;
  assign \new_[47587]_  = \new_[47586]_  & \new_[47583]_ ;
  assign \new_[47588]_  = \new_[47587]_  & \new_[47580]_ ;
  assign \new_[47591]_  = A168 & A169;
  assign \new_[47594]_  = A166 & ~A167;
  assign \new_[47595]_  = \new_[47594]_  & \new_[47591]_ ;
  assign \new_[47598]_  = A200 & ~A199;
  assign \new_[47601]_  = ~A203 & ~A201;
  assign \new_[47602]_  = \new_[47601]_  & \new_[47598]_ ;
  assign \new_[47603]_  = \new_[47602]_  & \new_[47595]_ ;
  assign \new_[47606]_  = ~A233 & ~A232;
  assign \new_[47609]_  = ~A236 & A235;
  assign \new_[47610]_  = \new_[47609]_  & \new_[47606]_ ;
  assign \new_[47613]_  = ~A266 & ~A265;
  assign \new_[47616]_  = ~A269 & A268;
  assign \new_[47617]_  = \new_[47616]_  & \new_[47613]_ ;
  assign \new_[47618]_  = \new_[47617]_  & \new_[47610]_ ;
  assign \new_[47621]_  = A168 & A169;
  assign \new_[47624]_  = A166 & ~A167;
  assign \new_[47625]_  = \new_[47624]_  & \new_[47621]_ ;
  assign \new_[47628]_  = ~A200 & A199;
  assign \new_[47631]_  = A202 & ~A201;
  assign \new_[47632]_  = \new_[47631]_  & \new_[47628]_ ;
  assign \new_[47633]_  = \new_[47632]_  & \new_[47625]_ ;
  assign \new_[47636]_  = A233 & A232;
  assign \new_[47639]_  = ~A236 & A235;
  assign \new_[47640]_  = \new_[47639]_  & \new_[47636]_ ;
  assign \new_[47643]_  = A299 & A298;
  assign \new_[47646]_  = ~A302 & A301;
  assign \new_[47647]_  = \new_[47646]_  & \new_[47643]_ ;
  assign \new_[47648]_  = \new_[47647]_  & \new_[47640]_ ;
  assign \new_[47651]_  = A168 & A169;
  assign \new_[47654]_  = A166 & ~A167;
  assign \new_[47655]_  = \new_[47654]_  & \new_[47651]_ ;
  assign \new_[47658]_  = ~A200 & A199;
  assign \new_[47661]_  = A202 & ~A201;
  assign \new_[47662]_  = \new_[47661]_  & \new_[47658]_ ;
  assign \new_[47663]_  = \new_[47662]_  & \new_[47655]_ ;
  assign \new_[47666]_  = A233 & A232;
  assign \new_[47669]_  = ~A236 & A235;
  assign \new_[47670]_  = \new_[47669]_  & \new_[47666]_ ;
  assign \new_[47673]_  = ~A299 & A298;
  assign \new_[47676]_  = A302 & ~A301;
  assign \new_[47677]_  = \new_[47676]_  & \new_[47673]_ ;
  assign \new_[47678]_  = \new_[47677]_  & \new_[47670]_ ;
  assign \new_[47681]_  = A168 & A169;
  assign \new_[47684]_  = A166 & ~A167;
  assign \new_[47685]_  = \new_[47684]_  & \new_[47681]_ ;
  assign \new_[47688]_  = ~A200 & A199;
  assign \new_[47691]_  = A202 & ~A201;
  assign \new_[47692]_  = \new_[47691]_  & \new_[47688]_ ;
  assign \new_[47693]_  = \new_[47692]_  & \new_[47685]_ ;
  assign \new_[47696]_  = A233 & A232;
  assign \new_[47699]_  = ~A236 & A235;
  assign \new_[47700]_  = \new_[47699]_  & \new_[47696]_ ;
  assign \new_[47703]_  = A299 & ~A298;
  assign \new_[47706]_  = A302 & ~A301;
  assign \new_[47707]_  = \new_[47706]_  & \new_[47703]_ ;
  assign \new_[47708]_  = \new_[47707]_  & \new_[47700]_ ;
  assign \new_[47711]_  = A168 & A169;
  assign \new_[47714]_  = A166 & ~A167;
  assign \new_[47715]_  = \new_[47714]_  & \new_[47711]_ ;
  assign \new_[47718]_  = ~A200 & A199;
  assign \new_[47721]_  = A202 & ~A201;
  assign \new_[47722]_  = \new_[47721]_  & \new_[47718]_ ;
  assign \new_[47723]_  = \new_[47722]_  & \new_[47715]_ ;
  assign \new_[47726]_  = A233 & A232;
  assign \new_[47729]_  = ~A236 & A235;
  assign \new_[47730]_  = \new_[47729]_  & \new_[47726]_ ;
  assign \new_[47733]_  = ~A299 & ~A298;
  assign \new_[47736]_  = ~A302 & A301;
  assign \new_[47737]_  = \new_[47736]_  & \new_[47733]_ ;
  assign \new_[47738]_  = \new_[47737]_  & \new_[47730]_ ;
  assign \new_[47741]_  = A168 & A169;
  assign \new_[47744]_  = A166 & ~A167;
  assign \new_[47745]_  = \new_[47744]_  & \new_[47741]_ ;
  assign \new_[47748]_  = ~A200 & A199;
  assign \new_[47751]_  = A202 & ~A201;
  assign \new_[47752]_  = \new_[47751]_  & \new_[47748]_ ;
  assign \new_[47753]_  = \new_[47752]_  & \new_[47745]_ ;
  assign \new_[47756]_  = A233 & A232;
  assign \new_[47759]_  = ~A236 & A235;
  assign \new_[47760]_  = \new_[47759]_  & \new_[47756]_ ;
  assign \new_[47763]_  = A266 & A265;
  assign \new_[47766]_  = ~A269 & A268;
  assign \new_[47767]_  = \new_[47766]_  & \new_[47763]_ ;
  assign \new_[47768]_  = \new_[47767]_  & \new_[47760]_ ;
  assign \new_[47771]_  = A168 & A169;
  assign \new_[47774]_  = A166 & ~A167;
  assign \new_[47775]_  = \new_[47774]_  & \new_[47771]_ ;
  assign \new_[47778]_  = ~A200 & A199;
  assign \new_[47781]_  = A202 & ~A201;
  assign \new_[47782]_  = \new_[47781]_  & \new_[47778]_ ;
  assign \new_[47783]_  = \new_[47782]_  & \new_[47775]_ ;
  assign \new_[47786]_  = A233 & A232;
  assign \new_[47789]_  = ~A236 & A235;
  assign \new_[47790]_  = \new_[47789]_  & \new_[47786]_ ;
  assign \new_[47793]_  = A266 & ~A265;
  assign \new_[47796]_  = A269 & ~A268;
  assign \new_[47797]_  = \new_[47796]_  & \new_[47793]_ ;
  assign \new_[47798]_  = \new_[47797]_  & \new_[47790]_ ;
  assign \new_[47801]_  = A168 & A169;
  assign \new_[47804]_  = A166 & ~A167;
  assign \new_[47805]_  = \new_[47804]_  & \new_[47801]_ ;
  assign \new_[47808]_  = ~A200 & A199;
  assign \new_[47811]_  = A202 & ~A201;
  assign \new_[47812]_  = \new_[47811]_  & \new_[47808]_ ;
  assign \new_[47813]_  = \new_[47812]_  & \new_[47805]_ ;
  assign \new_[47816]_  = A233 & A232;
  assign \new_[47819]_  = ~A236 & A235;
  assign \new_[47820]_  = \new_[47819]_  & \new_[47816]_ ;
  assign \new_[47823]_  = ~A266 & A265;
  assign \new_[47826]_  = A269 & ~A268;
  assign \new_[47827]_  = \new_[47826]_  & \new_[47823]_ ;
  assign \new_[47828]_  = \new_[47827]_  & \new_[47820]_ ;
  assign \new_[47831]_  = A168 & A169;
  assign \new_[47834]_  = A166 & ~A167;
  assign \new_[47835]_  = \new_[47834]_  & \new_[47831]_ ;
  assign \new_[47838]_  = ~A200 & A199;
  assign \new_[47841]_  = A202 & ~A201;
  assign \new_[47842]_  = \new_[47841]_  & \new_[47838]_ ;
  assign \new_[47843]_  = \new_[47842]_  & \new_[47835]_ ;
  assign \new_[47846]_  = A233 & A232;
  assign \new_[47849]_  = ~A236 & A235;
  assign \new_[47850]_  = \new_[47849]_  & \new_[47846]_ ;
  assign \new_[47853]_  = ~A266 & ~A265;
  assign \new_[47856]_  = ~A269 & A268;
  assign \new_[47857]_  = \new_[47856]_  & \new_[47853]_ ;
  assign \new_[47858]_  = \new_[47857]_  & \new_[47850]_ ;
  assign \new_[47861]_  = A168 & A169;
  assign \new_[47864]_  = A166 & ~A167;
  assign \new_[47865]_  = \new_[47864]_  & \new_[47861]_ ;
  assign \new_[47868]_  = ~A200 & A199;
  assign \new_[47871]_  = A202 & ~A201;
  assign \new_[47872]_  = \new_[47871]_  & \new_[47868]_ ;
  assign \new_[47873]_  = \new_[47872]_  & \new_[47865]_ ;
  assign \new_[47876]_  = A233 & ~A232;
  assign \new_[47879]_  = A236 & ~A235;
  assign \new_[47880]_  = \new_[47879]_  & \new_[47876]_ ;
  assign \new_[47883]_  = A299 & A298;
  assign \new_[47886]_  = ~A302 & A301;
  assign \new_[47887]_  = \new_[47886]_  & \new_[47883]_ ;
  assign \new_[47888]_  = \new_[47887]_  & \new_[47880]_ ;
  assign \new_[47891]_  = A168 & A169;
  assign \new_[47894]_  = A166 & ~A167;
  assign \new_[47895]_  = \new_[47894]_  & \new_[47891]_ ;
  assign \new_[47898]_  = ~A200 & A199;
  assign \new_[47901]_  = A202 & ~A201;
  assign \new_[47902]_  = \new_[47901]_  & \new_[47898]_ ;
  assign \new_[47903]_  = \new_[47902]_  & \new_[47895]_ ;
  assign \new_[47906]_  = A233 & ~A232;
  assign \new_[47909]_  = A236 & ~A235;
  assign \new_[47910]_  = \new_[47909]_  & \new_[47906]_ ;
  assign \new_[47913]_  = ~A299 & A298;
  assign \new_[47916]_  = A302 & ~A301;
  assign \new_[47917]_  = \new_[47916]_  & \new_[47913]_ ;
  assign \new_[47918]_  = \new_[47917]_  & \new_[47910]_ ;
  assign \new_[47921]_  = A168 & A169;
  assign \new_[47924]_  = A166 & ~A167;
  assign \new_[47925]_  = \new_[47924]_  & \new_[47921]_ ;
  assign \new_[47928]_  = ~A200 & A199;
  assign \new_[47931]_  = A202 & ~A201;
  assign \new_[47932]_  = \new_[47931]_  & \new_[47928]_ ;
  assign \new_[47933]_  = \new_[47932]_  & \new_[47925]_ ;
  assign \new_[47936]_  = A233 & ~A232;
  assign \new_[47939]_  = A236 & ~A235;
  assign \new_[47940]_  = \new_[47939]_  & \new_[47936]_ ;
  assign \new_[47943]_  = A299 & ~A298;
  assign \new_[47946]_  = A302 & ~A301;
  assign \new_[47947]_  = \new_[47946]_  & \new_[47943]_ ;
  assign \new_[47948]_  = \new_[47947]_  & \new_[47940]_ ;
  assign \new_[47951]_  = A168 & A169;
  assign \new_[47954]_  = A166 & ~A167;
  assign \new_[47955]_  = \new_[47954]_  & \new_[47951]_ ;
  assign \new_[47958]_  = ~A200 & A199;
  assign \new_[47961]_  = A202 & ~A201;
  assign \new_[47962]_  = \new_[47961]_  & \new_[47958]_ ;
  assign \new_[47963]_  = \new_[47962]_  & \new_[47955]_ ;
  assign \new_[47966]_  = A233 & ~A232;
  assign \new_[47969]_  = A236 & ~A235;
  assign \new_[47970]_  = \new_[47969]_  & \new_[47966]_ ;
  assign \new_[47973]_  = ~A299 & ~A298;
  assign \new_[47976]_  = ~A302 & A301;
  assign \new_[47977]_  = \new_[47976]_  & \new_[47973]_ ;
  assign \new_[47978]_  = \new_[47977]_  & \new_[47970]_ ;
  assign \new_[47981]_  = A168 & A169;
  assign \new_[47984]_  = A166 & ~A167;
  assign \new_[47985]_  = \new_[47984]_  & \new_[47981]_ ;
  assign \new_[47988]_  = ~A200 & A199;
  assign \new_[47991]_  = A202 & ~A201;
  assign \new_[47992]_  = \new_[47991]_  & \new_[47988]_ ;
  assign \new_[47993]_  = \new_[47992]_  & \new_[47985]_ ;
  assign \new_[47996]_  = A233 & ~A232;
  assign \new_[47999]_  = A236 & ~A235;
  assign \new_[48000]_  = \new_[47999]_  & \new_[47996]_ ;
  assign \new_[48003]_  = A266 & A265;
  assign \new_[48006]_  = ~A269 & A268;
  assign \new_[48007]_  = \new_[48006]_  & \new_[48003]_ ;
  assign \new_[48008]_  = \new_[48007]_  & \new_[48000]_ ;
  assign \new_[48011]_  = A168 & A169;
  assign \new_[48014]_  = A166 & ~A167;
  assign \new_[48015]_  = \new_[48014]_  & \new_[48011]_ ;
  assign \new_[48018]_  = ~A200 & A199;
  assign \new_[48021]_  = A202 & ~A201;
  assign \new_[48022]_  = \new_[48021]_  & \new_[48018]_ ;
  assign \new_[48023]_  = \new_[48022]_  & \new_[48015]_ ;
  assign \new_[48026]_  = A233 & ~A232;
  assign \new_[48029]_  = A236 & ~A235;
  assign \new_[48030]_  = \new_[48029]_  & \new_[48026]_ ;
  assign \new_[48033]_  = A266 & ~A265;
  assign \new_[48036]_  = A269 & ~A268;
  assign \new_[48037]_  = \new_[48036]_  & \new_[48033]_ ;
  assign \new_[48038]_  = \new_[48037]_  & \new_[48030]_ ;
  assign \new_[48041]_  = A168 & A169;
  assign \new_[48044]_  = A166 & ~A167;
  assign \new_[48045]_  = \new_[48044]_  & \new_[48041]_ ;
  assign \new_[48048]_  = ~A200 & A199;
  assign \new_[48051]_  = A202 & ~A201;
  assign \new_[48052]_  = \new_[48051]_  & \new_[48048]_ ;
  assign \new_[48053]_  = \new_[48052]_  & \new_[48045]_ ;
  assign \new_[48056]_  = A233 & ~A232;
  assign \new_[48059]_  = A236 & ~A235;
  assign \new_[48060]_  = \new_[48059]_  & \new_[48056]_ ;
  assign \new_[48063]_  = ~A266 & A265;
  assign \new_[48066]_  = A269 & ~A268;
  assign \new_[48067]_  = \new_[48066]_  & \new_[48063]_ ;
  assign \new_[48068]_  = \new_[48067]_  & \new_[48060]_ ;
  assign \new_[48071]_  = A168 & A169;
  assign \new_[48074]_  = A166 & ~A167;
  assign \new_[48075]_  = \new_[48074]_  & \new_[48071]_ ;
  assign \new_[48078]_  = ~A200 & A199;
  assign \new_[48081]_  = A202 & ~A201;
  assign \new_[48082]_  = \new_[48081]_  & \new_[48078]_ ;
  assign \new_[48083]_  = \new_[48082]_  & \new_[48075]_ ;
  assign \new_[48086]_  = A233 & ~A232;
  assign \new_[48089]_  = A236 & ~A235;
  assign \new_[48090]_  = \new_[48089]_  & \new_[48086]_ ;
  assign \new_[48093]_  = ~A266 & ~A265;
  assign \new_[48096]_  = ~A269 & A268;
  assign \new_[48097]_  = \new_[48096]_  & \new_[48093]_ ;
  assign \new_[48098]_  = \new_[48097]_  & \new_[48090]_ ;
  assign \new_[48101]_  = A168 & A169;
  assign \new_[48104]_  = A166 & ~A167;
  assign \new_[48105]_  = \new_[48104]_  & \new_[48101]_ ;
  assign \new_[48108]_  = ~A200 & A199;
  assign \new_[48111]_  = A202 & ~A201;
  assign \new_[48112]_  = \new_[48111]_  & \new_[48108]_ ;
  assign \new_[48113]_  = \new_[48112]_  & \new_[48105]_ ;
  assign \new_[48116]_  = ~A233 & A232;
  assign \new_[48119]_  = A236 & ~A235;
  assign \new_[48120]_  = \new_[48119]_  & \new_[48116]_ ;
  assign \new_[48123]_  = A299 & A298;
  assign \new_[48126]_  = ~A302 & A301;
  assign \new_[48127]_  = \new_[48126]_  & \new_[48123]_ ;
  assign \new_[48128]_  = \new_[48127]_  & \new_[48120]_ ;
  assign \new_[48131]_  = A168 & A169;
  assign \new_[48134]_  = A166 & ~A167;
  assign \new_[48135]_  = \new_[48134]_  & \new_[48131]_ ;
  assign \new_[48138]_  = ~A200 & A199;
  assign \new_[48141]_  = A202 & ~A201;
  assign \new_[48142]_  = \new_[48141]_  & \new_[48138]_ ;
  assign \new_[48143]_  = \new_[48142]_  & \new_[48135]_ ;
  assign \new_[48146]_  = ~A233 & A232;
  assign \new_[48149]_  = A236 & ~A235;
  assign \new_[48150]_  = \new_[48149]_  & \new_[48146]_ ;
  assign \new_[48153]_  = ~A299 & A298;
  assign \new_[48156]_  = A302 & ~A301;
  assign \new_[48157]_  = \new_[48156]_  & \new_[48153]_ ;
  assign \new_[48158]_  = \new_[48157]_  & \new_[48150]_ ;
  assign \new_[48161]_  = A168 & A169;
  assign \new_[48164]_  = A166 & ~A167;
  assign \new_[48165]_  = \new_[48164]_  & \new_[48161]_ ;
  assign \new_[48168]_  = ~A200 & A199;
  assign \new_[48171]_  = A202 & ~A201;
  assign \new_[48172]_  = \new_[48171]_  & \new_[48168]_ ;
  assign \new_[48173]_  = \new_[48172]_  & \new_[48165]_ ;
  assign \new_[48176]_  = ~A233 & A232;
  assign \new_[48179]_  = A236 & ~A235;
  assign \new_[48180]_  = \new_[48179]_  & \new_[48176]_ ;
  assign \new_[48183]_  = A299 & ~A298;
  assign \new_[48186]_  = A302 & ~A301;
  assign \new_[48187]_  = \new_[48186]_  & \new_[48183]_ ;
  assign \new_[48188]_  = \new_[48187]_  & \new_[48180]_ ;
  assign \new_[48191]_  = A168 & A169;
  assign \new_[48194]_  = A166 & ~A167;
  assign \new_[48195]_  = \new_[48194]_  & \new_[48191]_ ;
  assign \new_[48198]_  = ~A200 & A199;
  assign \new_[48201]_  = A202 & ~A201;
  assign \new_[48202]_  = \new_[48201]_  & \new_[48198]_ ;
  assign \new_[48203]_  = \new_[48202]_  & \new_[48195]_ ;
  assign \new_[48206]_  = ~A233 & A232;
  assign \new_[48209]_  = A236 & ~A235;
  assign \new_[48210]_  = \new_[48209]_  & \new_[48206]_ ;
  assign \new_[48213]_  = ~A299 & ~A298;
  assign \new_[48216]_  = ~A302 & A301;
  assign \new_[48217]_  = \new_[48216]_  & \new_[48213]_ ;
  assign \new_[48218]_  = \new_[48217]_  & \new_[48210]_ ;
  assign \new_[48221]_  = A168 & A169;
  assign \new_[48224]_  = A166 & ~A167;
  assign \new_[48225]_  = \new_[48224]_  & \new_[48221]_ ;
  assign \new_[48228]_  = ~A200 & A199;
  assign \new_[48231]_  = A202 & ~A201;
  assign \new_[48232]_  = \new_[48231]_  & \new_[48228]_ ;
  assign \new_[48233]_  = \new_[48232]_  & \new_[48225]_ ;
  assign \new_[48236]_  = ~A233 & A232;
  assign \new_[48239]_  = A236 & ~A235;
  assign \new_[48240]_  = \new_[48239]_  & \new_[48236]_ ;
  assign \new_[48243]_  = A266 & A265;
  assign \new_[48246]_  = ~A269 & A268;
  assign \new_[48247]_  = \new_[48246]_  & \new_[48243]_ ;
  assign \new_[48248]_  = \new_[48247]_  & \new_[48240]_ ;
  assign \new_[48251]_  = A168 & A169;
  assign \new_[48254]_  = A166 & ~A167;
  assign \new_[48255]_  = \new_[48254]_  & \new_[48251]_ ;
  assign \new_[48258]_  = ~A200 & A199;
  assign \new_[48261]_  = A202 & ~A201;
  assign \new_[48262]_  = \new_[48261]_  & \new_[48258]_ ;
  assign \new_[48263]_  = \new_[48262]_  & \new_[48255]_ ;
  assign \new_[48266]_  = ~A233 & A232;
  assign \new_[48269]_  = A236 & ~A235;
  assign \new_[48270]_  = \new_[48269]_  & \new_[48266]_ ;
  assign \new_[48273]_  = A266 & ~A265;
  assign \new_[48276]_  = A269 & ~A268;
  assign \new_[48277]_  = \new_[48276]_  & \new_[48273]_ ;
  assign \new_[48278]_  = \new_[48277]_  & \new_[48270]_ ;
  assign \new_[48281]_  = A168 & A169;
  assign \new_[48284]_  = A166 & ~A167;
  assign \new_[48285]_  = \new_[48284]_  & \new_[48281]_ ;
  assign \new_[48288]_  = ~A200 & A199;
  assign \new_[48291]_  = A202 & ~A201;
  assign \new_[48292]_  = \new_[48291]_  & \new_[48288]_ ;
  assign \new_[48293]_  = \new_[48292]_  & \new_[48285]_ ;
  assign \new_[48296]_  = ~A233 & A232;
  assign \new_[48299]_  = A236 & ~A235;
  assign \new_[48300]_  = \new_[48299]_  & \new_[48296]_ ;
  assign \new_[48303]_  = ~A266 & A265;
  assign \new_[48306]_  = A269 & ~A268;
  assign \new_[48307]_  = \new_[48306]_  & \new_[48303]_ ;
  assign \new_[48308]_  = \new_[48307]_  & \new_[48300]_ ;
  assign \new_[48311]_  = A168 & A169;
  assign \new_[48314]_  = A166 & ~A167;
  assign \new_[48315]_  = \new_[48314]_  & \new_[48311]_ ;
  assign \new_[48318]_  = ~A200 & A199;
  assign \new_[48321]_  = A202 & ~A201;
  assign \new_[48322]_  = \new_[48321]_  & \new_[48318]_ ;
  assign \new_[48323]_  = \new_[48322]_  & \new_[48315]_ ;
  assign \new_[48326]_  = ~A233 & A232;
  assign \new_[48329]_  = A236 & ~A235;
  assign \new_[48330]_  = \new_[48329]_  & \new_[48326]_ ;
  assign \new_[48333]_  = ~A266 & ~A265;
  assign \new_[48336]_  = ~A269 & A268;
  assign \new_[48337]_  = \new_[48336]_  & \new_[48333]_ ;
  assign \new_[48338]_  = \new_[48337]_  & \new_[48330]_ ;
  assign \new_[48341]_  = A168 & A169;
  assign \new_[48344]_  = A166 & ~A167;
  assign \new_[48345]_  = \new_[48344]_  & \new_[48341]_ ;
  assign \new_[48348]_  = ~A200 & A199;
  assign \new_[48351]_  = A202 & ~A201;
  assign \new_[48352]_  = \new_[48351]_  & \new_[48348]_ ;
  assign \new_[48353]_  = \new_[48352]_  & \new_[48345]_ ;
  assign \new_[48356]_  = ~A233 & ~A232;
  assign \new_[48359]_  = ~A236 & A235;
  assign \new_[48360]_  = \new_[48359]_  & \new_[48356]_ ;
  assign \new_[48363]_  = A299 & A298;
  assign \new_[48366]_  = ~A302 & A301;
  assign \new_[48367]_  = \new_[48366]_  & \new_[48363]_ ;
  assign \new_[48368]_  = \new_[48367]_  & \new_[48360]_ ;
  assign \new_[48371]_  = A168 & A169;
  assign \new_[48374]_  = A166 & ~A167;
  assign \new_[48375]_  = \new_[48374]_  & \new_[48371]_ ;
  assign \new_[48378]_  = ~A200 & A199;
  assign \new_[48381]_  = A202 & ~A201;
  assign \new_[48382]_  = \new_[48381]_  & \new_[48378]_ ;
  assign \new_[48383]_  = \new_[48382]_  & \new_[48375]_ ;
  assign \new_[48386]_  = ~A233 & ~A232;
  assign \new_[48389]_  = ~A236 & A235;
  assign \new_[48390]_  = \new_[48389]_  & \new_[48386]_ ;
  assign \new_[48393]_  = ~A299 & A298;
  assign \new_[48396]_  = A302 & ~A301;
  assign \new_[48397]_  = \new_[48396]_  & \new_[48393]_ ;
  assign \new_[48398]_  = \new_[48397]_  & \new_[48390]_ ;
  assign \new_[48401]_  = A168 & A169;
  assign \new_[48404]_  = A166 & ~A167;
  assign \new_[48405]_  = \new_[48404]_  & \new_[48401]_ ;
  assign \new_[48408]_  = ~A200 & A199;
  assign \new_[48411]_  = A202 & ~A201;
  assign \new_[48412]_  = \new_[48411]_  & \new_[48408]_ ;
  assign \new_[48413]_  = \new_[48412]_  & \new_[48405]_ ;
  assign \new_[48416]_  = ~A233 & ~A232;
  assign \new_[48419]_  = ~A236 & A235;
  assign \new_[48420]_  = \new_[48419]_  & \new_[48416]_ ;
  assign \new_[48423]_  = A299 & ~A298;
  assign \new_[48426]_  = A302 & ~A301;
  assign \new_[48427]_  = \new_[48426]_  & \new_[48423]_ ;
  assign \new_[48428]_  = \new_[48427]_  & \new_[48420]_ ;
  assign \new_[48431]_  = A168 & A169;
  assign \new_[48434]_  = A166 & ~A167;
  assign \new_[48435]_  = \new_[48434]_  & \new_[48431]_ ;
  assign \new_[48438]_  = ~A200 & A199;
  assign \new_[48441]_  = A202 & ~A201;
  assign \new_[48442]_  = \new_[48441]_  & \new_[48438]_ ;
  assign \new_[48443]_  = \new_[48442]_  & \new_[48435]_ ;
  assign \new_[48446]_  = ~A233 & ~A232;
  assign \new_[48449]_  = ~A236 & A235;
  assign \new_[48450]_  = \new_[48449]_  & \new_[48446]_ ;
  assign \new_[48453]_  = ~A299 & ~A298;
  assign \new_[48456]_  = ~A302 & A301;
  assign \new_[48457]_  = \new_[48456]_  & \new_[48453]_ ;
  assign \new_[48458]_  = \new_[48457]_  & \new_[48450]_ ;
  assign \new_[48461]_  = A168 & A169;
  assign \new_[48464]_  = A166 & ~A167;
  assign \new_[48465]_  = \new_[48464]_  & \new_[48461]_ ;
  assign \new_[48468]_  = ~A200 & A199;
  assign \new_[48471]_  = A202 & ~A201;
  assign \new_[48472]_  = \new_[48471]_  & \new_[48468]_ ;
  assign \new_[48473]_  = \new_[48472]_  & \new_[48465]_ ;
  assign \new_[48476]_  = ~A233 & ~A232;
  assign \new_[48479]_  = ~A236 & A235;
  assign \new_[48480]_  = \new_[48479]_  & \new_[48476]_ ;
  assign \new_[48483]_  = A266 & A265;
  assign \new_[48486]_  = ~A269 & A268;
  assign \new_[48487]_  = \new_[48486]_  & \new_[48483]_ ;
  assign \new_[48488]_  = \new_[48487]_  & \new_[48480]_ ;
  assign \new_[48491]_  = A168 & A169;
  assign \new_[48494]_  = A166 & ~A167;
  assign \new_[48495]_  = \new_[48494]_  & \new_[48491]_ ;
  assign \new_[48498]_  = ~A200 & A199;
  assign \new_[48501]_  = A202 & ~A201;
  assign \new_[48502]_  = \new_[48501]_  & \new_[48498]_ ;
  assign \new_[48503]_  = \new_[48502]_  & \new_[48495]_ ;
  assign \new_[48506]_  = ~A233 & ~A232;
  assign \new_[48509]_  = ~A236 & A235;
  assign \new_[48510]_  = \new_[48509]_  & \new_[48506]_ ;
  assign \new_[48513]_  = A266 & ~A265;
  assign \new_[48516]_  = A269 & ~A268;
  assign \new_[48517]_  = \new_[48516]_  & \new_[48513]_ ;
  assign \new_[48518]_  = \new_[48517]_  & \new_[48510]_ ;
  assign \new_[48521]_  = A168 & A169;
  assign \new_[48524]_  = A166 & ~A167;
  assign \new_[48525]_  = \new_[48524]_  & \new_[48521]_ ;
  assign \new_[48528]_  = ~A200 & A199;
  assign \new_[48531]_  = A202 & ~A201;
  assign \new_[48532]_  = \new_[48531]_  & \new_[48528]_ ;
  assign \new_[48533]_  = \new_[48532]_  & \new_[48525]_ ;
  assign \new_[48536]_  = ~A233 & ~A232;
  assign \new_[48539]_  = ~A236 & A235;
  assign \new_[48540]_  = \new_[48539]_  & \new_[48536]_ ;
  assign \new_[48543]_  = ~A266 & A265;
  assign \new_[48546]_  = A269 & ~A268;
  assign \new_[48547]_  = \new_[48546]_  & \new_[48543]_ ;
  assign \new_[48548]_  = \new_[48547]_  & \new_[48540]_ ;
  assign \new_[48551]_  = A168 & A169;
  assign \new_[48554]_  = A166 & ~A167;
  assign \new_[48555]_  = \new_[48554]_  & \new_[48551]_ ;
  assign \new_[48558]_  = ~A200 & A199;
  assign \new_[48561]_  = A202 & ~A201;
  assign \new_[48562]_  = \new_[48561]_  & \new_[48558]_ ;
  assign \new_[48563]_  = \new_[48562]_  & \new_[48555]_ ;
  assign \new_[48566]_  = ~A233 & ~A232;
  assign \new_[48569]_  = ~A236 & A235;
  assign \new_[48570]_  = \new_[48569]_  & \new_[48566]_ ;
  assign \new_[48573]_  = ~A266 & ~A265;
  assign \new_[48576]_  = ~A269 & A268;
  assign \new_[48577]_  = \new_[48576]_  & \new_[48573]_ ;
  assign \new_[48578]_  = \new_[48577]_  & \new_[48570]_ ;
  assign \new_[48581]_  = A168 & A169;
  assign \new_[48584]_  = A166 & ~A167;
  assign \new_[48585]_  = \new_[48584]_  & \new_[48581]_ ;
  assign \new_[48588]_  = ~A200 & A199;
  assign \new_[48591]_  = ~A203 & ~A201;
  assign \new_[48592]_  = \new_[48591]_  & \new_[48588]_ ;
  assign \new_[48593]_  = \new_[48592]_  & \new_[48585]_ ;
  assign \new_[48596]_  = A233 & A232;
  assign \new_[48599]_  = ~A236 & A235;
  assign \new_[48600]_  = \new_[48599]_  & \new_[48596]_ ;
  assign \new_[48603]_  = A299 & A298;
  assign \new_[48606]_  = ~A302 & A301;
  assign \new_[48607]_  = \new_[48606]_  & \new_[48603]_ ;
  assign \new_[48608]_  = \new_[48607]_  & \new_[48600]_ ;
  assign \new_[48611]_  = A168 & A169;
  assign \new_[48614]_  = A166 & ~A167;
  assign \new_[48615]_  = \new_[48614]_  & \new_[48611]_ ;
  assign \new_[48618]_  = ~A200 & A199;
  assign \new_[48621]_  = ~A203 & ~A201;
  assign \new_[48622]_  = \new_[48621]_  & \new_[48618]_ ;
  assign \new_[48623]_  = \new_[48622]_  & \new_[48615]_ ;
  assign \new_[48626]_  = A233 & A232;
  assign \new_[48629]_  = ~A236 & A235;
  assign \new_[48630]_  = \new_[48629]_  & \new_[48626]_ ;
  assign \new_[48633]_  = ~A299 & A298;
  assign \new_[48636]_  = A302 & ~A301;
  assign \new_[48637]_  = \new_[48636]_  & \new_[48633]_ ;
  assign \new_[48638]_  = \new_[48637]_  & \new_[48630]_ ;
  assign \new_[48641]_  = A168 & A169;
  assign \new_[48644]_  = A166 & ~A167;
  assign \new_[48645]_  = \new_[48644]_  & \new_[48641]_ ;
  assign \new_[48648]_  = ~A200 & A199;
  assign \new_[48651]_  = ~A203 & ~A201;
  assign \new_[48652]_  = \new_[48651]_  & \new_[48648]_ ;
  assign \new_[48653]_  = \new_[48652]_  & \new_[48645]_ ;
  assign \new_[48656]_  = A233 & A232;
  assign \new_[48659]_  = ~A236 & A235;
  assign \new_[48660]_  = \new_[48659]_  & \new_[48656]_ ;
  assign \new_[48663]_  = A299 & ~A298;
  assign \new_[48666]_  = A302 & ~A301;
  assign \new_[48667]_  = \new_[48666]_  & \new_[48663]_ ;
  assign \new_[48668]_  = \new_[48667]_  & \new_[48660]_ ;
  assign \new_[48671]_  = A168 & A169;
  assign \new_[48674]_  = A166 & ~A167;
  assign \new_[48675]_  = \new_[48674]_  & \new_[48671]_ ;
  assign \new_[48678]_  = ~A200 & A199;
  assign \new_[48681]_  = ~A203 & ~A201;
  assign \new_[48682]_  = \new_[48681]_  & \new_[48678]_ ;
  assign \new_[48683]_  = \new_[48682]_  & \new_[48675]_ ;
  assign \new_[48686]_  = A233 & A232;
  assign \new_[48689]_  = ~A236 & A235;
  assign \new_[48690]_  = \new_[48689]_  & \new_[48686]_ ;
  assign \new_[48693]_  = ~A299 & ~A298;
  assign \new_[48696]_  = ~A302 & A301;
  assign \new_[48697]_  = \new_[48696]_  & \new_[48693]_ ;
  assign \new_[48698]_  = \new_[48697]_  & \new_[48690]_ ;
  assign \new_[48701]_  = A168 & A169;
  assign \new_[48704]_  = A166 & ~A167;
  assign \new_[48705]_  = \new_[48704]_  & \new_[48701]_ ;
  assign \new_[48708]_  = ~A200 & A199;
  assign \new_[48711]_  = ~A203 & ~A201;
  assign \new_[48712]_  = \new_[48711]_  & \new_[48708]_ ;
  assign \new_[48713]_  = \new_[48712]_  & \new_[48705]_ ;
  assign \new_[48716]_  = A233 & A232;
  assign \new_[48719]_  = ~A236 & A235;
  assign \new_[48720]_  = \new_[48719]_  & \new_[48716]_ ;
  assign \new_[48723]_  = A266 & A265;
  assign \new_[48726]_  = ~A269 & A268;
  assign \new_[48727]_  = \new_[48726]_  & \new_[48723]_ ;
  assign \new_[48728]_  = \new_[48727]_  & \new_[48720]_ ;
  assign \new_[48731]_  = A168 & A169;
  assign \new_[48734]_  = A166 & ~A167;
  assign \new_[48735]_  = \new_[48734]_  & \new_[48731]_ ;
  assign \new_[48738]_  = ~A200 & A199;
  assign \new_[48741]_  = ~A203 & ~A201;
  assign \new_[48742]_  = \new_[48741]_  & \new_[48738]_ ;
  assign \new_[48743]_  = \new_[48742]_  & \new_[48735]_ ;
  assign \new_[48746]_  = A233 & A232;
  assign \new_[48749]_  = ~A236 & A235;
  assign \new_[48750]_  = \new_[48749]_  & \new_[48746]_ ;
  assign \new_[48753]_  = A266 & ~A265;
  assign \new_[48756]_  = A269 & ~A268;
  assign \new_[48757]_  = \new_[48756]_  & \new_[48753]_ ;
  assign \new_[48758]_  = \new_[48757]_  & \new_[48750]_ ;
  assign \new_[48761]_  = A168 & A169;
  assign \new_[48764]_  = A166 & ~A167;
  assign \new_[48765]_  = \new_[48764]_  & \new_[48761]_ ;
  assign \new_[48768]_  = ~A200 & A199;
  assign \new_[48771]_  = ~A203 & ~A201;
  assign \new_[48772]_  = \new_[48771]_  & \new_[48768]_ ;
  assign \new_[48773]_  = \new_[48772]_  & \new_[48765]_ ;
  assign \new_[48776]_  = A233 & A232;
  assign \new_[48779]_  = ~A236 & A235;
  assign \new_[48780]_  = \new_[48779]_  & \new_[48776]_ ;
  assign \new_[48783]_  = ~A266 & A265;
  assign \new_[48786]_  = A269 & ~A268;
  assign \new_[48787]_  = \new_[48786]_  & \new_[48783]_ ;
  assign \new_[48788]_  = \new_[48787]_  & \new_[48780]_ ;
  assign \new_[48791]_  = A168 & A169;
  assign \new_[48794]_  = A166 & ~A167;
  assign \new_[48795]_  = \new_[48794]_  & \new_[48791]_ ;
  assign \new_[48798]_  = ~A200 & A199;
  assign \new_[48801]_  = ~A203 & ~A201;
  assign \new_[48802]_  = \new_[48801]_  & \new_[48798]_ ;
  assign \new_[48803]_  = \new_[48802]_  & \new_[48795]_ ;
  assign \new_[48806]_  = A233 & A232;
  assign \new_[48809]_  = ~A236 & A235;
  assign \new_[48810]_  = \new_[48809]_  & \new_[48806]_ ;
  assign \new_[48813]_  = ~A266 & ~A265;
  assign \new_[48816]_  = ~A269 & A268;
  assign \new_[48817]_  = \new_[48816]_  & \new_[48813]_ ;
  assign \new_[48818]_  = \new_[48817]_  & \new_[48810]_ ;
  assign \new_[48821]_  = A168 & A169;
  assign \new_[48824]_  = A166 & ~A167;
  assign \new_[48825]_  = \new_[48824]_  & \new_[48821]_ ;
  assign \new_[48828]_  = ~A200 & A199;
  assign \new_[48831]_  = ~A203 & ~A201;
  assign \new_[48832]_  = \new_[48831]_  & \new_[48828]_ ;
  assign \new_[48833]_  = \new_[48832]_  & \new_[48825]_ ;
  assign \new_[48836]_  = A233 & ~A232;
  assign \new_[48839]_  = A236 & ~A235;
  assign \new_[48840]_  = \new_[48839]_  & \new_[48836]_ ;
  assign \new_[48843]_  = A299 & A298;
  assign \new_[48846]_  = ~A302 & A301;
  assign \new_[48847]_  = \new_[48846]_  & \new_[48843]_ ;
  assign \new_[48848]_  = \new_[48847]_  & \new_[48840]_ ;
  assign \new_[48851]_  = A168 & A169;
  assign \new_[48854]_  = A166 & ~A167;
  assign \new_[48855]_  = \new_[48854]_  & \new_[48851]_ ;
  assign \new_[48858]_  = ~A200 & A199;
  assign \new_[48861]_  = ~A203 & ~A201;
  assign \new_[48862]_  = \new_[48861]_  & \new_[48858]_ ;
  assign \new_[48863]_  = \new_[48862]_  & \new_[48855]_ ;
  assign \new_[48866]_  = A233 & ~A232;
  assign \new_[48869]_  = A236 & ~A235;
  assign \new_[48870]_  = \new_[48869]_  & \new_[48866]_ ;
  assign \new_[48873]_  = ~A299 & A298;
  assign \new_[48876]_  = A302 & ~A301;
  assign \new_[48877]_  = \new_[48876]_  & \new_[48873]_ ;
  assign \new_[48878]_  = \new_[48877]_  & \new_[48870]_ ;
  assign \new_[48881]_  = A168 & A169;
  assign \new_[48884]_  = A166 & ~A167;
  assign \new_[48885]_  = \new_[48884]_  & \new_[48881]_ ;
  assign \new_[48888]_  = ~A200 & A199;
  assign \new_[48891]_  = ~A203 & ~A201;
  assign \new_[48892]_  = \new_[48891]_  & \new_[48888]_ ;
  assign \new_[48893]_  = \new_[48892]_  & \new_[48885]_ ;
  assign \new_[48896]_  = A233 & ~A232;
  assign \new_[48899]_  = A236 & ~A235;
  assign \new_[48900]_  = \new_[48899]_  & \new_[48896]_ ;
  assign \new_[48903]_  = A299 & ~A298;
  assign \new_[48906]_  = A302 & ~A301;
  assign \new_[48907]_  = \new_[48906]_  & \new_[48903]_ ;
  assign \new_[48908]_  = \new_[48907]_  & \new_[48900]_ ;
  assign \new_[48911]_  = A168 & A169;
  assign \new_[48914]_  = A166 & ~A167;
  assign \new_[48915]_  = \new_[48914]_  & \new_[48911]_ ;
  assign \new_[48918]_  = ~A200 & A199;
  assign \new_[48921]_  = ~A203 & ~A201;
  assign \new_[48922]_  = \new_[48921]_  & \new_[48918]_ ;
  assign \new_[48923]_  = \new_[48922]_  & \new_[48915]_ ;
  assign \new_[48926]_  = A233 & ~A232;
  assign \new_[48929]_  = A236 & ~A235;
  assign \new_[48930]_  = \new_[48929]_  & \new_[48926]_ ;
  assign \new_[48933]_  = ~A299 & ~A298;
  assign \new_[48936]_  = ~A302 & A301;
  assign \new_[48937]_  = \new_[48936]_  & \new_[48933]_ ;
  assign \new_[48938]_  = \new_[48937]_  & \new_[48930]_ ;
  assign \new_[48941]_  = A168 & A169;
  assign \new_[48944]_  = A166 & ~A167;
  assign \new_[48945]_  = \new_[48944]_  & \new_[48941]_ ;
  assign \new_[48948]_  = ~A200 & A199;
  assign \new_[48951]_  = ~A203 & ~A201;
  assign \new_[48952]_  = \new_[48951]_  & \new_[48948]_ ;
  assign \new_[48953]_  = \new_[48952]_  & \new_[48945]_ ;
  assign \new_[48956]_  = A233 & ~A232;
  assign \new_[48959]_  = A236 & ~A235;
  assign \new_[48960]_  = \new_[48959]_  & \new_[48956]_ ;
  assign \new_[48963]_  = A266 & A265;
  assign \new_[48966]_  = ~A269 & A268;
  assign \new_[48967]_  = \new_[48966]_  & \new_[48963]_ ;
  assign \new_[48968]_  = \new_[48967]_  & \new_[48960]_ ;
  assign \new_[48971]_  = A168 & A169;
  assign \new_[48974]_  = A166 & ~A167;
  assign \new_[48975]_  = \new_[48974]_  & \new_[48971]_ ;
  assign \new_[48978]_  = ~A200 & A199;
  assign \new_[48981]_  = ~A203 & ~A201;
  assign \new_[48982]_  = \new_[48981]_  & \new_[48978]_ ;
  assign \new_[48983]_  = \new_[48982]_  & \new_[48975]_ ;
  assign \new_[48986]_  = A233 & ~A232;
  assign \new_[48989]_  = A236 & ~A235;
  assign \new_[48990]_  = \new_[48989]_  & \new_[48986]_ ;
  assign \new_[48993]_  = A266 & ~A265;
  assign \new_[48996]_  = A269 & ~A268;
  assign \new_[48997]_  = \new_[48996]_  & \new_[48993]_ ;
  assign \new_[48998]_  = \new_[48997]_  & \new_[48990]_ ;
  assign \new_[49001]_  = A168 & A169;
  assign \new_[49004]_  = A166 & ~A167;
  assign \new_[49005]_  = \new_[49004]_  & \new_[49001]_ ;
  assign \new_[49008]_  = ~A200 & A199;
  assign \new_[49011]_  = ~A203 & ~A201;
  assign \new_[49012]_  = \new_[49011]_  & \new_[49008]_ ;
  assign \new_[49013]_  = \new_[49012]_  & \new_[49005]_ ;
  assign \new_[49016]_  = A233 & ~A232;
  assign \new_[49019]_  = A236 & ~A235;
  assign \new_[49020]_  = \new_[49019]_  & \new_[49016]_ ;
  assign \new_[49023]_  = ~A266 & A265;
  assign \new_[49026]_  = A269 & ~A268;
  assign \new_[49027]_  = \new_[49026]_  & \new_[49023]_ ;
  assign \new_[49028]_  = \new_[49027]_  & \new_[49020]_ ;
  assign \new_[49031]_  = A168 & A169;
  assign \new_[49034]_  = A166 & ~A167;
  assign \new_[49035]_  = \new_[49034]_  & \new_[49031]_ ;
  assign \new_[49038]_  = ~A200 & A199;
  assign \new_[49041]_  = ~A203 & ~A201;
  assign \new_[49042]_  = \new_[49041]_  & \new_[49038]_ ;
  assign \new_[49043]_  = \new_[49042]_  & \new_[49035]_ ;
  assign \new_[49046]_  = A233 & ~A232;
  assign \new_[49049]_  = A236 & ~A235;
  assign \new_[49050]_  = \new_[49049]_  & \new_[49046]_ ;
  assign \new_[49053]_  = ~A266 & ~A265;
  assign \new_[49056]_  = ~A269 & A268;
  assign \new_[49057]_  = \new_[49056]_  & \new_[49053]_ ;
  assign \new_[49058]_  = \new_[49057]_  & \new_[49050]_ ;
  assign \new_[49061]_  = A168 & A169;
  assign \new_[49064]_  = A166 & ~A167;
  assign \new_[49065]_  = \new_[49064]_  & \new_[49061]_ ;
  assign \new_[49068]_  = ~A200 & A199;
  assign \new_[49071]_  = ~A203 & ~A201;
  assign \new_[49072]_  = \new_[49071]_  & \new_[49068]_ ;
  assign \new_[49073]_  = \new_[49072]_  & \new_[49065]_ ;
  assign \new_[49076]_  = ~A233 & A232;
  assign \new_[49079]_  = A236 & ~A235;
  assign \new_[49080]_  = \new_[49079]_  & \new_[49076]_ ;
  assign \new_[49083]_  = A299 & A298;
  assign \new_[49086]_  = ~A302 & A301;
  assign \new_[49087]_  = \new_[49086]_  & \new_[49083]_ ;
  assign \new_[49088]_  = \new_[49087]_  & \new_[49080]_ ;
  assign \new_[49091]_  = A168 & A169;
  assign \new_[49094]_  = A166 & ~A167;
  assign \new_[49095]_  = \new_[49094]_  & \new_[49091]_ ;
  assign \new_[49098]_  = ~A200 & A199;
  assign \new_[49101]_  = ~A203 & ~A201;
  assign \new_[49102]_  = \new_[49101]_  & \new_[49098]_ ;
  assign \new_[49103]_  = \new_[49102]_  & \new_[49095]_ ;
  assign \new_[49106]_  = ~A233 & A232;
  assign \new_[49109]_  = A236 & ~A235;
  assign \new_[49110]_  = \new_[49109]_  & \new_[49106]_ ;
  assign \new_[49113]_  = ~A299 & A298;
  assign \new_[49116]_  = A302 & ~A301;
  assign \new_[49117]_  = \new_[49116]_  & \new_[49113]_ ;
  assign \new_[49118]_  = \new_[49117]_  & \new_[49110]_ ;
  assign \new_[49121]_  = A168 & A169;
  assign \new_[49124]_  = A166 & ~A167;
  assign \new_[49125]_  = \new_[49124]_  & \new_[49121]_ ;
  assign \new_[49128]_  = ~A200 & A199;
  assign \new_[49131]_  = ~A203 & ~A201;
  assign \new_[49132]_  = \new_[49131]_  & \new_[49128]_ ;
  assign \new_[49133]_  = \new_[49132]_  & \new_[49125]_ ;
  assign \new_[49136]_  = ~A233 & A232;
  assign \new_[49139]_  = A236 & ~A235;
  assign \new_[49140]_  = \new_[49139]_  & \new_[49136]_ ;
  assign \new_[49143]_  = A299 & ~A298;
  assign \new_[49146]_  = A302 & ~A301;
  assign \new_[49147]_  = \new_[49146]_  & \new_[49143]_ ;
  assign \new_[49148]_  = \new_[49147]_  & \new_[49140]_ ;
  assign \new_[49151]_  = A168 & A169;
  assign \new_[49154]_  = A166 & ~A167;
  assign \new_[49155]_  = \new_[49154]_  & \new_[49151]_ ;
  assign \new_[49158]_  = ~A200 & A199;
  assign \new_[49161]_  = ~A203 & ~A201;
  assign \new_[49162]_  = \new_[49161]_  & \new_[49158]_ ;
  assign \new_[49163]_  = \new_[49162]_  & \new_[49155]_ ;
  assign \new_[49166]_  = ~A233 & A232;
  assign \new_[49169]_  = A236 & ~A235;
  assign \new_[49170]_  = \new_[49169]_  & \new_[49166]_ ;
  assign \new_[49173]_  = ~A299 & ~A298;
  assign \new_[49176]_  = ~A302 & A301;
  assign \new_[49177]_  = \new_[49176]_  & \new_[49173]_ ;
  assign \new_[49178]_  = \new_[49177]_  & \new_[49170]_ ;
  assign \new_[49181]_  = A168 & A169;
  assign \new_[49184]_  = A166 & ~A167;
  assign \new_[49185]_  = \new_[49184]_  & \new_[49181]_ ;
  assign \new_[49188]_  = ~A200 & A199;
  assign \new_[49191]_  = ~A203 & ~A201;
  assign \new_[49192]_  = \new_[49191]_  & \new_[49188]_ ;
  assign \new_[49193]_  = \new_[49192]_  & \new_[49185]_ ;
  assign \new_[49196]_  = ~A233 & A232;
  assign \new_[49199]_  = A236 & ~A235;
  assign \new_[49200]_  = \new_[49199]_  & \new_[49196]_ ;
  assign \new_[49203]_  = A266 & A265;
  assign \new_[49206]_  = ~A269 & A268;
  assign \new_[49207]_  = \new_[49206]_  & \new_[49203]_ ;
  assign \new_[49208]_  = \new_[49207]_  & \new_[49200]_ ;
  assign \new_[49211]_  = A168 & A169;
  assign \new_[49214]_  = A166 & ~A167;
  assign \new_[49215]_  = \new_[49214]_  & \new_[49211]_ ;
  assign \new_[49218]_  = ~A200 & A199;
  assign \new_[49221]_  = ~A203 & ~A201;
  assign \new_[49222]_  = \new_[49221]_  & \new_[49218]_ ;
  assign \new_[49223]_  = \new_[49222]_  & \new_[49215]_ ;
  assign \new_[49226]_  = ~A233 & A232;
  assign \new_[49229]_  = A236 & ~A235;
  assign \new_[49230]_  = \new_[49229]_  & \new_[49226]_ ;
  assign \new_[49233]_  = A266 & ~A265;
  assign \new_[49236]_  = A269 & ~A268;
  assign \new_[49237]_  = \new_[49236]_  & \new_[49233]_ ;
  assign \new_[49238]_  = \new_[49237]_  & \new_[49230]_ ;
  assign \new_[49241]_  = A168 & A169;
  assign \new_[49244]_  = A166 & ~A167;
  assign \new_[49245]_  = \new_[49244]_  & \new_[49241]_ ;
  assign \new_[49248]_  = ~A200 & A199;
  assign \new_[49251]_  = ~A203 & ~A201;
  assign \new_[49252]_  = \new_[49251]_  & \new_[49248]_ ;
  assign \new_[49253]_  = \new_[49252]_  & \new_[49245]_ ;
  assign \new_[49256]_  = ~A233 & A232;
  assign \new_[49259]_  = A236 & ~A235;
  assign \new_[49260]_  = \new_[49259]_  & \new_[49256]_ ;
  assign \new_[49263]_  = ~A266 & A265;
  assign \new_[49266]_  = A269 & ~A268;
  assign \new_[49267]_  = \new_[49266]_  & \new_[49263]_ ;
  assign \new_[49268]_  = \new_[49267]_  & \new_[49260]_ ;
  assign \new_[49271]_  = A168 & A169;
  assign \new_[49274]_  = A166 & ~A167;
  assign \new_[49275]_  = \new_[49274]_  & \new_[49271]_ ;
  assign \new_[49278]_  = ~A200 & A199;
  assign \new_[49281]_  = ~A203 & ~A201;
  assign \new_[49282]_  = \new_[49281]_  & \new_[49278]_ ;
  assign \new_[49283]_  = \new_[49282]_  & \new_[49275]_ ;
  assign \new_[49286]_  = ~A233 & A232;
  assign \new_[49289]_  = A236 & ~A235;
  assign \new_[49290]_  = \new_[49289]_  & \new_[49286]_ ;
  assign \new_[49293]_  = ~A266 & ~A265;
  assign \new_[49296]_  = ~A269 & A268;
  assign \new_[49297]_  = \new_[49296]_  & \new_[49293]_ ;
  assign \new_[49298]_  = \new_[49297]_  & \new_[49290]_ ;
  assign \new_[49301]_  = A168 & A169;
  assign \new_[49304]_  = A166 & ~A167;
  assign \new_[49305]_  = \new_[49304]_  & \new_[49301]_ ;
  assign \new_[49308]_  = ~A200 & A199;
  assign \new_[49311]_  = ~A203 & ~A201;
  assign \new_[49312]_  = \new_[49311]_  & \new_[49308]_ ;
  assign \new_[49313]_  = \new_[49312]_  & \new_[49305]_ ;
  assign \new_[49316]_  = ~A233 & ~A232;
  assign \new_[49319]_  = ~A236 & A235;
  assign \new_[49320]_  = \new_[49319]_  & \new_[49316]_ ;
  assign \new_[49323]_  = A299 & A298;
  assign \new_[49326]_  = ~A302 & A301;
  assign \new_[49327]_  = \new_[49326]_  & \new_[49323]_ ;
  assign \new_[49328]_  = \new_[49327]_  & \new_[49320]_ ;
  assign \new_[49331]_  = A168 & A169;
  assign \new_[49334]_  = A166 & ~A167;
  assign \new_[49335]_  = \new_[49334]_  & \new_[49331]_ ;
  assign \new_[49338]_  = ~A200 & A199;
  assign \new_[49341]_  = ~A203 & ~A201;
  assign \new_[49342]_  = \new_[49341]_  & \new_[49338]_ ;
  assign \new_[49343]_  = \new_[49342]_  & \new_[49335]_ ;
  assign \new_[49346]_  = ~A233 & ~A232;
  assign \new_[49349]_  = ~A236 & A235;
  assign \new_[49350]_  = \new_[49349]_  & \new_[49346]_ ;
  assign \new_[49353]_  = ~A299 & A298;
  assign \new_[49356]_  = A302 & ~A301;
  assign \new_[49357]_  = \new_[49356]_  & \new_[49353]_ ;
  assign \new_[49358]_  = \new_[49357]_  & \new_[49350]_ ;
  assign \new_[49361]_  = A168 & A169;
  assign \new_[49364]_  = A166 & ~A167;
  assign \new_[49365]_  = \new_[49364]_  & \new_[49361]_ ;
  assign \new_[49368]_  = ~A200 & A199;
  assign \new_[49371]_  = ~A203 & ~A201;
  assign \new_[49372]_  = \new_[49371]_  & \new_[49368]_ ;
  assign \new_[49373]_  = \new_[49372]_  & \new_[49365]_ ;
  assign \new_[49376]_  = ~A233 & ~A232;
  assign \new_[49379]_  = ~A236 & A235;
  assign \new_[49380]_  = \new_[49379]_  & \new_[49376]_ ;
  assign \new_[49383]_  = A299 & ~A298;
  assign \new_[49386]_  = A302 & ~A301;
  assign \new_[49387]_  = \new_[49386]_  & \new_[49383]_ ;
  assign \new_[49388]_  = \new_[49387]_  & \new_[49380]_ ;
  assign \new_[49391]_  = A168 & A169;
  assign \new_[49394]_  = A166 & ~A167;
  assign \new_[49395]_  = \new_[49394]_  & \new_[49391]_ ;
  assign \new_[49398]_  = ~A200 & A199;
  assign \new_[49401]_  = ~A203 & ~A201;
  assign \new_[49402]_  = \new_[49401]_  & \new_[49398]_ ;
  assign \new_[49403]_  = \new_[49402]_  & \new_[49395]_ ;
  assign \new_[49406]_  = ~A233 & ~A232;
  assign \new_[49409]_  = ~A236 & A235;
  assign \new_[49410]_  = \new_[49409]_  & \new_[49406]_ ;
  assign \new_[49413]_  = ~A299 & ~A298;
  assign \new_[49416]_  = ~A302 & A301;
  assign \new_[49417]_  = \new_[49416]_  & \new_[49413]_ ;
  assign \new_[49418]_  = \new_[49417]_  & \new_[49410]_ ;
  assign \new_[49421]_  = A168 & A169;
  assign \new_[49424]_  = A166 & ~A167;
  assign \new_[49425]_  = \new_[49424]_  & \new_[49421]_ ;
  assign \new_[49428]_  = ~A200 & A199;
  assign \new_[49431]_  = ~A203 & ~A201;
  assign \new_[49432]_  = \new_[49431]_  & \new_[49428]_ ;
  assign \new_[49433]_  = \new_[49432]_  & \new_[49425]_ ;
  assign \new_[49436]_  = ~A233 & ~A232;
  assign \new_[49439]_  = ~A236 & A235;
  assign \new_[49440]_  = \new_[49439]_  & \new_[49436]_ ;
  assign \new_[49443]_  = A266 & A265;
  assign \new_[49446]_  = ~A269 & A268;
  assign \new_[49447]_  = \new_[49446]_  & \new_[49443]_ ;
  assign \new_[49448]_  = \new_[49447]_  & \new_[49440]_ ;
  assign \new_[49451]_  = A168 & A169;
  assign \new_[49454]_  = A166 & ~A167;
  assign \new_[49455]_  = \new_[49454]_  & \new_[49451]_ ;
  assign \new_[49458]_  = ~A200 & A199;
  assign \new_[49461]_  = ~A203 & ~A201;
  assign \new_[49462]_  = \new_[49461]_  & \new_[49458]_ ;
  assign \new_[49463]_  = \new_[49462]_  & \new_[49455]_ ;
  assign \new_[49466]_  = ~A233 & ~A232;
  assign \new_[49469]_  = ~A236 & A235;
  assign \new_[49470]_  = \new_[49469]_  & \new_[49466]_ ;
  assign \new_[49473]_  = A266 & ~A265;
  assign \new_[49476]_  = A269 & ~A268;
  assign \new_[49477]_  = \new_[49476]_  & \new_[49473]_ ;
  assign \new_[49478]_  = \new_[49477]_  & \new_[49470]_ ;
  assign \new_[49481]_  = A168 & A169;
  assign \new_[49484]_  = A166 & ~A167;
  assign \new_[49485]_  = \new_[49484]_  & \new_[49481]_ ;
  assign \new_[49488]_  = ~A200 & A199;
  assign \new_[49491]_  = ~A203 & ~A201;
  assign \new_[49492]_  = \new_[49491]_  & \new_[49488]_ ;
  assign \new_[49493]_  = \new_[49492]_  & \new_[49485]_ ;
  assign \new_[49496]_  = ~A233 & ~A232;
  assign \new_[49499]_  = ~A236 & A235;
  assign \new_[49500]_  = \new_[49499]_  & \new_[49496]_ ;
  assign \new_[49503]_  = ~A266 & A265;
  assign \new_[49506]_  = A269 & ~A268;
  assign \new_[49507]_  = \new_[49506]_  & \new_[49503]_ ;
  assign \new_[49508]_  = \new_[49507]_  & \new_[49500]_ ;
  assign \new_[49511]_  = A168 & A169;
  assign \new_[49514]_  = A166 & ~A167;
  assign \new_[49515]_  = \new_[49514]_  & \new_[49511]_ ;
  assign \new_[49518]_  = ~A200 & A199;
  assign \new_[49521]_  = ~A203 & ~A201;
  assign \new_[49522]_  = \new_[49521]_  & \new_[49518]_ ;
  assign \new_[49523]_  = \new_[49522]_  & \new_[49515]_ ;
  assign \new_[49526]_  = ~A233 & ~A232;
  assign \new_[49529]_  = ~A236 & A235;
  assign \new_[49530]_  = \new_[49529]_  & \new_[49526]_ ;
  assign \new_[49533]_  = ~A266 & ~A265;
  assign \new_[49536]_  = ~A269 & A268;
  assign \new_[49537]_  = \new_[49536]_  & \new_[49533]_ ;
  assign \new_[49538]_  = \new_[49537]_  & \new_[49530]_ ;
endmodule


