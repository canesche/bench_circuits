module bigkey ( clock, 
    \key<255> , \key<254> , \key<253> , \key<252> , \key<251> , \key<250> ,
    \key<249> , \key<248> , \key<247> , \key<246> , \key<245> , \key<244> ,
    \key<243> , \key<242> , \key<241> , \key<240> , \key<239> , \key<238> ,
    \key<237> , \key<236> , \key<235> , \key<234> , \key<233> , \key<232> ,
    \key<231> , \key<230> , \key<229> , \key<228> , \key<227> , \key<226> ,
    \key<225> , \key<224> , \key<223> , \key<222> , \key<221> , \key<220> ,
    \key<219> , \key<218> , \key<217> , \key<216> , \key<215> , \key<214> ,
    \key<213> , \key<212> , \key<211> , \key<210> , \key<209> , \key<208> ,
    \key<207> , \key<206> , \key<205> , \key<204> , \key<203> , \key<202> ,
    \key<201> , \key<200> , \key<199> , \key<198> , \key<197> , \key<196> ,
    \key<195> , \key<194> , \key<193> , \key<192> , \key<191> , \key<190> ,
    \key<189> , \key<188> , \key<187> , \key<186> , \key<185> , \key<184> ,
    \key<183> , \key<182> , \key<181> , \key<180> , \key<179> , \key<178> ,
    \key<177> , \key<176> , \key<175> , \key<174> , \key<173> , \key<172> ,
    \key<171> , \key<170> , \key<169> , \key<168> , \key<167> , \key<166> ,
    \key<165> , \key<164> , \key<163> , \key<162> , \key<161> , \key<160> ,
    \key<159> , \key<158> , \key<157> , \key<156> , \key<155> , \key<154> ,
    \key<153> , \key<152> , \key<151> , \key<150> , \key<149> , \key<148> ,
    \key<147> , \key<146> , \key<145> , \key<144> , \key<143> , \key<142> ,
    \key<141> , \key<140> , \key<139> , \key<138> , \key<137> , \key<136> ,
    \key<135> , \key<134> , \key<133> , \key<132> , \key<131> , \key<130> ,
    \key<129> , \key<128> , \key<127> , \key<126> , \key<125> , \key<124> ,
    \key<123> , \key<122> , \key<121> , \key<120> , \key<119> , \key<118> ,
    \key<117> , \key<116> , \key<115> , \key<114> , \key<113> , \key<112> ,
    \key<111> , \key<110> , \key<109> , \key<108> , \key<107> , \key<106> ,
    \key<105> , \key<104> , \key<103> , \key<102> , \key<101> , \key<100> ,
    \key<99> , \key<98> , \key<97> , \key<96> , \key<95> , \key<94> ,
    \key<93> , \key<92> , \key<91> , \key<90> , \key<89> , \key<88> ,
    \key<87> , \key<86> , \key<85> , \key<84> , \key<83> , \key<82> ,
    \key<81> , \key<80> , \key<79> , \key<78> , \key<77> , \key<76> ,
    \key<75> , \key<74> , \key<73> , \key<72> , \key<71> , \key<70> ,
    \key<69> , \key<68> , \key<67> , \key<66> , \key<65> , \key<64> ,
    \key<63> , \key<62> , \key<61> , \key<60> , \key<59> , \key<58> ,
    \key<57> , \key<56> , \key<55> , \key<54> , \key<53> , \key<52> ,
    \key<51> , \key<50> , \key<49> , \key<48> , \key<47> , \key<46> ,
    \key<45> , \key<44> , \key<43> , \key<42> , \key<41> , \key<40> ,
    \key<39> , \key<38> , \key<37> , \key<36> , \key<35> , \key<34> ,
    \key<33> , \key<32> , \key<31> , \key<30> , \key<29> , \key<28> ,
    \key<27> , \key<26> , \key<25> , \key<24> , \key<23> , \key<22> ,
    \key<21> , \key<20> , \key<19> , \key<18> , \key<17> , \key<16> ,
    \key<15> , \key<14> , \key<13> , \key<12> , \key<11> , \key<10> ,
    \key<9> , \key<8> , \key<7> , \key<6> , \key<5> , \key<4> , \key<3> ,
    \key<2> , \key<1> , \key<0> , \encrypt<0> , \start<0> , \count<3> ,
    \count<2> , \count<1> , \count<0> ,
    \new_count<3> , \new_count<2> , \new_count<1> , \new_count<0> ,
    \data_ready<0> , \KSi<191> , \KSi<190> , \KSi<189> , \KSi<188> ,
    \KSi<187> , \KSi<186> , \KSi<185> , \KSi<184> , \KSi<183> , \KSi<182> ,
    \KSi<181> , \KSi<180> , \KSi<179> , \KSi<178> , \KSi<177> , \KSi<176> ,
    \KSi<175> , \KSi<174> , \KSi<173> , \KSi<172> , \KSi<171> , \KSi<170> ,
    \KSi<169> , \KSi<168> , \KSi<167> , \KSi<166> , \KSi<165> , \KSi<164> ,
    \KSi<163> , \KSi<162> , \KSi<161> , \KSi<160> , \KSi<159> , \KSi<158> ,
    \KSi<157> , \KSi<156> , \KSi<155> , \KSi<154> , \KSi<153> , \KSi<152> ,
    \KSi<151> , \KSi<150> , \KSi<149> , \KSi<148> , \KSi<147> , \KSi<146> ,
    \KSi<145> , \KSi<144> , \KSi<143> , \KSi<142> , \KSi<141> , \KSi<140> ,
    \KSi<139> , \KSi<138> , \KSi<137> , \KSi<136> , \KSi<135> , \KSi<134> ,
    \KSi<133> , \KSi<132> , \KSi<131> , \KSi<130> , \KSi<129> , \KSi<128> ,
    \KSi<127> , \KSi<126> , \KSi<125> , \KSi<124> , \KSi<123> , \KSi<122> ,
    \KSi<121> , \KSi<120> , \KSi<119> , \KSi<118> , \KSi<117> , \KSi<116> ,
    \KSi<115> , \KSi<114> , \KSi<113> , \KSi<112> , \KSi<111> , \KSi<110> ,
    \KSi<109> , \KSi<108> , \KSi<107> , \KSi<106> , \KSi<105> , \KSi<104> ,
    \KSi<103> , \KSi<102> , \KSi<101> , \KSi<100> , \KSi<99> , \KSi<98> ,
    \KSi<97> , \KSi<96> , \KSi<95> , \KSi<94> , \KSi<93> , \KSi<92> ,
    \KSi<91> , \KSi<90> , \KSi<89> , \KSi<88> , \KSi<87> , \KSi<86> ,
    \KSi<85> , \KSi<84> , \KSi<83> , \KSi<82> , \KSi<81> , \KSi<80> ,
    \KSi<79> , \KSi<78> , \KSi<77> , \KSi<76> , \KSi<75> , \KSi<74> ,
    \KSi<73> , \KSi<72> , \KSi<71> , \KSi<70> , \KSi<69> , \KSi<68> ,
    \KSi<67> , \KSi<66> , \KSi<65> , \KSi<64> , \KSi<63> , \KSi<62> ,
    \KSi<61> , \KSi<60> , \KSi<59> , \KSi<58> , \KSi<57> , \KSi<56> ,
    \KSi<55> , \KSi<54> , \KSi<53> , \KSi<52> , \KSi<51> , \KSi<50> ,
    \KSi<49> , \KSi<48> , \KSi<47> , \KSi<46> , \KSi<45> , \KSi<44> ,
    \KSi<43> , \KSi<42> , \KSi<41> , \KSi<40> , \KSi<39> , \KSi<38> ,
    \KSi<37> , \KSi<36> , \KSi<35> , \KSi<34> , \KSi<33> , \KSi<32> ,
    \KSi<31> , \KSi<30> , \KSi<29> , \KSi<28> , \KSi<27> , \KSi<26> ,
    \KSi<25> , \KSi<24> , \KSi<23> , \KSi<22> , \KSi<21> , \KSi<20> ,
    \KSi<19> , \KSi<18> , \KSi<17> , \KSi<16> , \KSi<15> , \KSi<14> ,
    \KSi<13> , \KSi<12> , \KSi<11> , \KSi<10> , \KSi<9> , \KSi<8> ,
    \KSi<7> , \KSi<6> , \KSi<5> , \KSi<4> , \KSi<3> , \KSi<2> , \KSi<1> ,
    \KSi<0>   );
  input  clock;
  input  \key<255> , \key<254> , \key<253> , \key<252> , \key<251> ,
    \key<250> , \key<249> , \key<248> , \key<247> , \key<246> , \key<245> ,
    \key<244> , \key<243> , \key<242> , \key<241> , \key<240> , \key<239> ,
    \key<238> , \key<237> , \key<236> , \key<235> , \key<234> , \key<233> ,
    \key<232> , \key<231> , \key<230> , \key<229> , \key<228> , \key<227> ,
    \key<226> , \key<225> , \key<224> , \key<223> , \key<222> , \key<221> ,
    \key<220> , \key<219> , \key<218> , \key<217> , \key<216> , \key<215> ,
    \key<214> , \key<213> , \key<212> , \key<211> , \key<210> , \key<209> ,
    \key<208> , \key<207> , \key<206> , \key<205> , \key<204> , \key<203> ,
    \key<202> , \key<201> , \key<200> , \key<199> , \key<198> , \key<197> ,
    \key<196> , \key<195> , \key<194> , \key<193> , \key<192> , \key<191> ,
    \key<190> , \key<189> , \key<188> , \key<187> , \key<186> , \key<185> ,
    \key<184> , \key<183> , \key<182> , \key<181> , \key<180> , \key<179> ,
    \key<178> , \key<177> , \key<176> , \key<175> , \key<174> , \key<173> ,
    \key<172> , \key<171> , \key<170> , \key<169> , \key<168> , \key<167> ,
    \key<166> , \key<165> , \key<164> , \key<163> , \key<162> , \key<161> ,
    \key<160> , \key<159> , \key<158> , \key<157> , \key<156> , \key<155> ,
    \key<154> , \key<153> , \key<152> , \key<151> , \key<150> , \key<149> ,
    \key<148> , \key<147> , \key<146> , \key<145> , \key<144> , \key<143> ,
    \key<142> , \key<141> , \key<140> , \key<139> , \key<138> , \key<137> ,
    \key<136> , \key<135> , \key<134> , \key<133> , \key<132> , \key<131> ,
    \key<130> , \key<129> , \key<128> , \key<127> , \key<126> , \key<125> ,
    \key<124> , \key<123> , \key<122> , \key<121> , \key<120> , \key<119> ,
    \key<118> , \key<117> , \key<116> , \key<115> , \key<114> , \key<113> ,
    \key<112> , \key<111> , \key<110> , \key<109> , \key<108> , \key<107> ,
    \key<106> , \key<105> , \key<104> , \key<103> , \key<102> , \key<101> ,
    \key<100> , \key<99> , \key<98> , \key<97> , \key<96> , \key<95> ,
    \key<94> , \key<93> , \key<92> , \key<91> , \key<90> , \key<89> ,
    \key<88> , \key<87> , \key<86> , \key<85> , \key<84> , \key<83> ,
    \key<82> , \key<81> , \key<80> , \key<79> , \key<78> , \key<77> ,
    \key<76> , \key<75> , \key<74> , \key<73> , \key<72> , \key<71> ,
    \key<70> , \key<69> , \key<68> , \key<67> , \key<66> , \key<65> ,
    \key<64> , \key<63> , \key<62> , \key<61> , \key<60> , \key<59> ,
    \key<58> , \key<57> , \key<56> , \key<55> , \key<54> , \key<53> ,
    \key<52> , \key<51> , \key<50> , \key<49> , \key<48> , \key<47> ,
    \key<46> , \key<45> , \key<44> , \key<43> , \key<42> , \key<41> ,
    \key<40> , \key<39> , \key<38> , \key<37> , \key<36> , \key<35> ,
    \key<34> , \key<33> , \key<32> , \key<31> , \key<30> , \key<29> ,
    \key<28> , \key<27> , \key<26> , \key<25> , \key<24> , \key<23> ,
    \key<22> , \key<21> , \key<20> , \key<19> , \key<18> , \key<17> ,
    \key<16> , \key<15> , \key<14> , \key<13> , \key<12> , \key<11> ,
    \key<10> , \key<9> , \key<8> , \key<7> , \key<6> , \key<5> , \key<4> ,
    \key<3> , \key<2> , \key<1> , \key<0> , \encrypt<0> , \start<0> ,
    \count<3> , \count<2> , \count<1> , \count<0> ;
  output \new_count<3> , \new_count<2> , \new_count<1> , \new_count<0> ,
    \data_ready<0> , \KSi<191> , \KSi<190> , \KSi<189> , \KSi<188> ,
    \KSi<187> , \KSi<186> , \KSi<185> , \KSi<184> , \KSi<183> , \KSi<182> ,
    \KSi<181> , \KSi<180> , \KSi<179> , \KSi<178> , \KSi<177> , \KSi<176> ,
    \KSi<175> , \KSi<174> , \KSi<173> , \KSi<172> , \KSi<171> , \KSi<170> ,
    \KSi<169> , \KSi<168> , \KSi<167> , \KSi<166> , \KSi<165> , \KSi<164> ,
    \KSi<163> , \KSi<162> , \KSi<161> , \KSi<160> , \KSi<159> , \KSi<158> ,
    \KSi<157> , \KSi<156> , \KSi<155> , \KSi<154> , \KSi<153> , \KSi<152> ,
    \KSi<151> , \KSi<150> , \KSi<149> , \KSi<148> , \KSi<147> , \KSi<146> ,
    \KSi<145> , \KSi<144> , \KSi<143> , \KSi<142> , \KSi<141> , \KSi<140> ,
    \KSi<139> , \KSi<138> , \KSi<137> , \KSi<136> , \KSi<135> , \KSi<134> ,
    \KSi<133> , \KSi<132> , \KSi<131> , \KSi<130> , \KSi<129> , \KSi<128> ,
    \KSi<127> , \KSi<126> , \KSi<125> , \KSi<124> , \KSi<123> , \KSi<122> ,
    \KSi<121> , \KSi<120> , \KSi<119> , \KSi<118> , \KSi<117> , \KSi<116> ,
    \KSi<115> , \KSi<114> , \KSi<113> , \KSi<112> , \KSi<111> , \KSi<110> ,
    \KSi<109> , \KSi<108> , \KSi<107> , \KSi<106> , \KSi<105> , \KSi<104> ,
    \KSi<103> , \KSi<102> , \KSi<101> , \KSi<100> , \KSi<99> , \KSi<98> ,
    \KSi<97> , \KSi<96> , \KSi<95> , \KSi<94> , \KSi<93> , \KSi<92> ,
    \KSi<91> , \KSi<90> , \KSi<89> , \KSi<88> , \KSi<87> , \KSi<86> ,
    \KSi<85> , \KSi<84> , \KSi<83> , \KSi<82> , \KSi<81> , \KSi<80> ,
    \KSi<79> , \KSi<78> , \KSi<77> , \KSi<76> , \KSi<75> , \KSi<74> ,
    \KSi<73> , \KSi<72> , \KSi<71> , \KSi<70> , \KSi<69> , \KSi<68> ,
    \KSi<67> , \KSi<66> , \KSi<65> , \KSi<64> , \KSi<63> , \KSi<62> ,
    \KSi<61> , \KSi<60> , \KSi<59> , \KSi<58> , \KSi<57> , \KSi<56> ,
    \KSi<55> , \KSi<54> , \KSi<53> , \KSi<52> , \KSi<51> , \KSi<50> ,
    \KSi<49> , \KSi<48> , \KSi<47> , \KSi<46> , \KSi<45> , \KSi<44> ,
    \KSi<43> , \KSi<42> , \KSi<41> , \KSi<40> , \KSi<39> , \KSi<38> ,
    \KSi<37> , \KSi<36> , \KSi<35> , \KSi<34> , \KSi<33> , \KSi<32> ,
    \KSi<31> , \KSi<30> , \KSi<29> , \KSi<28> , \KSi<27> , \KSi<26> ,
    \KSi<25> , \KSi<24> , \KSi<23> , \KSi<22> , \KSi<21> , \KSi<20> ,
    \KSi<19> , \KSi<18> , \KSi<17> , \KSi<16> , \KSi<15> , \KSi<14> ,
    \KSi<13> , \KSi<12> , \KSi<11> , \KSi<10> , \KSi<9> , \KSi<8> ,
    \KSi<7> , \KSi<6> , \KSi<5> , \KSi<4> , \KSi<3> , \KSi<2> , \KSi<1> ,
    \KSi<0> ;
  reg \C<111> , \C<110> , \C<109> , \C<108> , \C<107> , \C<106> , \C<105> ,
    \C<104> , \C<103> , \C<102> , \C<101> , \C<100> , \C<99> , \C<98> ,
    \C<97> , \C<96> , \C<95> , \C<94> , \C<93> , \C<92> , \C<91> , \C<90> ,
    \C<89> , \C<88> , \C<87> , \C<86> , \C<85> , \C<84> , \C<83> , \C<82> ,
    \C<81> , \C<80> , \C<79> , \C<78> , \C<77> , \C<76> , \C<75> , \C<74> ,
    \C<73> , \C<72> , \C<71> , \C<70> , \C<69> , \C<68> , \C<67> , \C<66> ,
    \C<65> , \C<64> , \C<63> , \C<62> , \C<61> , \C<60> , \C<59> , \C<58> ,
    \C<57> , \C<56> , \C<55> , \C<54> , \C<53> , \C<52> , \C<51> , \C<50> ,
    \C<49> , \C<48> , \C<47> , \C<46> , \C<45> , \C<44> , \C<43> , \C<42> ,
    \C<41> , \C<40> , \C<39> , \C<38> , \C<37> , \C<36> , \C<35> , \C<34> ,
    \C<33> , \C<32> , \C<31> , \C<30> , \C<29> , \C<28> , \C<27> , \C<26> ,
    \C<25> , \C<24> , \C<23> , \C<22> , \C<21> , \C<20> , \C<19> , \C<18> ,
    \C<17> , \C<16> , \C<15> , \C<14> , \C<13> , \C<12> , \C<11> , \C<10> ,
    \C<9> , \C<8> , \C<7> , \C<6> , \C<5> , \C<4> , \C<3> , \C<2> , \C<1> ,
    \C<0> , \D<111> , \D<110> , \D<109> , \D<108> , \D<107> , \D<106> ,
    \D<105> , \D<104> , \D<103> , \D<102> , \D<101> , \D<100> , \D<99> ,
    \D<98> , \D<97> , \D<96> , \D<95> , \D<94> , \D<93> , \D<92> , \D<91> ,
    \D<90> , \D<89> , \D<88> , \D<87> , \D<86> , \D<85> , \D<84> , \D<83> ,
    \D<82> , \D<81> , \D<80> , \D<79> , \D<78> , \D<77> , \D<76> , \D<75> ,
    \D<74> , \D<73> , \D<72> , \D<71> , \D<70> , \D<69> , \D<68> , \D<67> ,
    \D<66> , \D<65> , \D<64> , \D<63> , \D<62> , \D<61> , \D<60> , \D<59> ,
    \D<58> , \D<57> , \D<56> , \D<55> , \D<54> , \D<53> , \D<52> , \D<51> ,
    \D<50> , \D<49> , \D<48> , \D<47> , \D<46> , \D<45> , \D<44> , \D<43> ,
    \D<42> , \D<41> , \D<40> , \D<39> , \D<38> , \D<37> , \D<36> , \D<35> ,
    \D<34> , \D<33> , \D<32> , \D<31> , \D<30> , \D<29> , \D<28> , \D<27> ,
    \D<26> , \D<25> , \D<24> , \D<23> , \D<22> , \D<21> , \D<20> , \D<19> ,
    \D<18> , \D<17> , \D<16> , \D<15> , \D<14> , \D<13> , \D<12> , \D<11> ,
    \D<10> , \D<9> , \D<8> , \D<7> , \D<6> , \D<5> , \D<4> , \D<3> ,
    \D<2> , \D<1> , \D<0> ;
  wire new_n1132_, new_n1133_, new_n1134_, new_n1135_1_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_1_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_1_, new_n1146_,
    new_n1148_, new_n1149_, new_n1150_1_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_1_, new_n1156_, new_n1158_,
    new_n1159_, new_n1160_1_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_1_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_1_, new_n1172_, new_n1173_, new_n1174_, new_n1175_1_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_1_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_1_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_1_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_1_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_1_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1210_1_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_1_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_1_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_1_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_1_, new_n1231_, new_n1232_, new_n1234_,
    new_n1235_1_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_1_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_1_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1250_1_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_1_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_1_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_1_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_1_,
    new_n1276_, new_n1278_, new_n1279_, new_n1280_1_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_1_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_1_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_1_, new_n1296_,
    new_n1297_, new_n1298_, new_n1300_1_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_1_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_1_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_1_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_1_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_1_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_1_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_1_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_1_, new_n1341_, new_n1342_, new_n1344_,
    new_n1345_1_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_1_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_1_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_1_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_1_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_1_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_1_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_1_,
    new_n1386_, new_n1388_, new_n1389_, new_n1390_1_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_1_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_1_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_1_, new_n1406_,
    new_n1407_, new_n1408_, new_n1410_1_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_1_, new_n1416_, new_n1417_,
    new_n1418_, new_n1419_, new_n1420_1_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_1_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_1_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_1_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_1_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_1_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_1_, new_n1451_, new_n1452_, new_n1454_,
    new_n1455_1_, new_n1456_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_1_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_1_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_1_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_1_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_1_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_1_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_1_,
    new_n1496_, new_n1498_, new_n1499_, new_n1500_1_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_1_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_1_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_1_, new_n1516_,
    new_n1517_, new_n1518_, new_n1520_1_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_1_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_1_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_1_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_1_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_1_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_1_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_1_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_1_, new_n1561_, new_n1562_, new_n1564_,
    new_n1565_1_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_1_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_1_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_1_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_1_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_1_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_1_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_1_,
    new_n1606_, new_n1608_, new_n1609_, new_n1610_1_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_1_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_1_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_1_, new_n1626_,
    new_n1627_, new_n1628_, new_n1630_1_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_1_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_1_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_1_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_1_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_1_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_1_, new_n1661_, new_n1662_, new_n1663_,
    new_n1664_, new_n1665_1_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_1_, new_n1671_, new_n1672_, new_n1674_,
    new_n1675_1_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_1_, new_n1681_, new_n1682_, new_n1683_, new_n1684_,
    new_n1685_1_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_1_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_1_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_1_,
    new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_1_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_1_,
    new_n1716_, new_n1718_, new_n1719_, new_n1720_1_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_1_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_1_, new_n1731_,
    new_n1732_, new_n1733_, new_n1734_, new_n1735_1_, new_n1736_,
    new_n1737_, new_n1738_, new_n1740_1_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_1_, new_n1746_, new_n1747_,
    new_n1748_, new_n1749_, new_n1750_1_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_1_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_1_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_1_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_1_, new_n1771_, new_n1772_, new_n1773_,
    new_n1774_, new_n1775_1_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_1_, new_n1781_, new_n1782_, new_n1784_,
    new_n1785_1_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1790_1_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_1_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_1_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_1_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_1_,
    new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_1_,
    new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_1_,
    new_n1826_, new_n1828_, new_n1829_, new_n1830_1_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_1_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_1_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_1_, new_n1846_,
    new_n1847_, new_n1848_, new_n1850_1_, new_n1851_, new_n1852_,
    new_n1853_, new_n1854_, new_n1855_1_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_1_, new_n1861_, new_n1862_,
    new_n1863_, new_n1864_, new_n1865_1_, new_n1866_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_1_, new_n1872_, new_n1873_,
    new_n1874_, new_n1875_1_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_1_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_1_, new_n1886_, new_n1887_, new_n1888_,
    new_n1889_, new_n1890_1_, new_n1891_, new_n1892_, new_n1894_,
    new_n1895_1_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_1_, new_n1901_, new_n1902_, new_n1903_, new_n1904_,
    new_n1905_1_, new_n1906_, new_n1907_, new_n1908_, new_n1909_,
    new_n1910_1_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_1_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_1_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_1_,
    new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_1_,
    new_n1936_, new_n1938_, new_n1939_, new_n1940_1_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_1_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_1_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_1_, new_n1956_,
    new_n1957_, new_n1958_, new_n1960_1_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_1_, new_n1966_, new_n1967_,
    new_n1968_, new_n1969_, new_n1970_1_, new_n1971_, new_n1972_,
    new_n1973_, new_n1974_, new_n1975_1_, new_n1976_, new_n1977_,
    new_n1978_, new_n1979_, new_n1980_1_, new_n1982_, new_n1983_,
    new_n1984_, new_n1985_1_, new_n1986_, new_n1987_, new_n1988_,
    new_n1989_, new_n1990_1_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_1_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_1_, new_n2001_, new_n2002_, new_n2004_,
    new_n2005_1_, new_n2006_, new_n2007_, new_n2008_, new_n2009_,
    new_n2010_1_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_1_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_1_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_1_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_1_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2070_, new_n2071_, new_n2072_, new_n2073_,
    new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_,
    new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_,
    new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2114_, new_n2115_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_,
    new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_,
    new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_,
    new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2180_,
    new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_,
    new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_,
    new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_,
    new_n2199_, new_n2200_, new_n2202_, new_n2203_, new_n2204_, new_n2205_,
    new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_,
    new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_,
    new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2224_,
    new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_,
    new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_,
    new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_,
    new_n2243_, new_n2244_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2290_, new_n2291_, new_n2292_, new_n2293_,
    new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_,
    new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_,
    new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2334_, new_n2335_, new_n2336_, new_n2337_,
    new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_,
    new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_,
    new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2356_,
    new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_,
    new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_,
    new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_,
    new_n2375_, new_n2376_, new_n2378_, new_n2379_, new_n2380_, new_n2381_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2422_, new_n2423_, new_n2424_, new_n2425_,
    new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_,
    new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_,
    new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2444_,
    new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_,
    new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_,
    new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_,
    new_n2463_, new_n2464_, new_n2466_, new_n2467_, new_n2468_, new_n2469_,
    new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_,
    new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_,
    new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2554_, new_n2555_, new_n2556_, new_n2557_,
    new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_,
    new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_,
    new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2576_,
    new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_,
    new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_,
    new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_,
    new_n2595_, new_n2596_, new_n2598_, new_n2599_, new_n2600_, new_n2601_,
    new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_,
    new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_,
    new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2686_, new_n2687_, new_n2688_, new_n2689_,
    new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_,
    new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_,
    new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2708_,
    new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_,
    new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_,
    new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_,
    new_n2727_, new_n2728_, new_n2730_, new_n2731_, new_n2732_, new_n2733_,
    new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_,
    new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_,
    new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2752_,
    new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_,
    new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_,
    new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_,
    new_n2771_, new_n2772_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2796_,
    new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_,
    new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2818_, new_n2819_, new_n2820_, new_n2821_,
    new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_,
    new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_,
    new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2840_,
    new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_,
    new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_,
    new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_,
    new_n2859_, new_n2860_, new_n2862_, new_n2863_, new_n2864_, new_n2865_,
    new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_,
    new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_,
    new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2884_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_,
    new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_,
    new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2904_, new_n2906_, new_n2907_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2928_,
    new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_,
    new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2950_, new_n2951_, new_n2952_, new_n2953_,
    new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_,
    new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_,
    new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2994_, new_n2995_, new_n2996_, new_n2997_,
    new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_,
    new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_,
    new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3016_,
    new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_,
    new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_,
    new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_,
    new_n3035_, new_n3036_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3060_,
    new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_,
    new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_,
    new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_,
    new_n3079_, new_n3080_, new_n3082_, new_n3083_, new_n3084_, new_n3085_,
    new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_,
    new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_,
    new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3104_,
    new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_,
    new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_,
    new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_,
    new_n3123_, new_n3124_, new_n3126_, new_n3127_, new_n3128_, new_n3129_,
    new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_,
    new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_,
    new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3148_,
    new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_,
    new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_,
    new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_,
    new_n3167_, new_n3168_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3192_,
    new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_,
    new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_,
    new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_,
    new_n3211_, new_n3212_, new_n3214_, new_n3215_, new_n3216_, new_n3217_,
    new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_,
    new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_,
    new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3236_,
    new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_,
    new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_,
    new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_,
    new_n3255_, new_n3256_, new_n3258_, new_n3259_, new_n3260_, new_n3261_,
    new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_,
    new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3280_,
    new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_,
    new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_,
    new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_,
    new_n3299_, new_n3300_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3324_,
    new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3346_, new_n3347_, new_n3348_, new_n3349_,
    new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_,
    new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_,
    new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3368_,
    new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_,
    new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_,
    new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_,
    new_n3387_, new_n3388_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3412_,
    new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_,
    new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_,
    new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_,
    new_n3431_, new_n3432_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3456_,
    new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_,
    new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_,
    new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_,
    new_n3475_, new_n3476_, new_n3478_, new_n3479_, new_n3480_, new_n3481_,
    new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_,
    new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_,
    new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3500_,
    new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_,
    new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_,
    new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_,
    new_n3519_, new_n3520_, new_n3522_, new_n3523_, new_n3524_, new_n3525_,
    new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_,
    new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_,
    new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3544_,
    new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_,
    new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_,
    new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_,
    new_n3563_, new_n3564_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3588_,
    new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_,
    new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_,
    new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_,
    new_n3607_, new_n3608_, new_n3610_, new_n3611_, new_n3612_, new_n3613_,
    new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_,
    new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_,
    new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3632_,
    new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_,
    new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_,
    new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_,
    new_n3651_, new_n3652_, new_n3654_, new_n3655_, new_n3656_, new_n3657_,
    new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_,
    new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_,
    new_n3670_, new_n3671_, new_n3673_, new_n3674_, new_n3675_, new_n3676_,
    new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_,
    new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_,
    new_n3689_, new_n3690_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3711_, new_n3712_, new_n3713_, new_n3714_,
    new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_,
    new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_,
    new_n3727_, new_n3728_, new_n3730_, new_n3731_, new_n3732_, new_n3733_,
    new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_,
    new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_,
    new_n3746_, new_n3747_, new_n3749_, new_n3750_, new_n3751_, new_n3752_,
    new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_,
    new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_,
    new_n3765_, new_n3766_, new_n3768_, new_n3769_, new_n3770_, new_n3771_,
    new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_,
    new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_,
    new_n3784_, new_n3785_, new_n3787_, new_n3788_, new_n3789_, new_n3790_,
    new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_,
    new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_,
    new_n3803_, new_n3804_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3825_, new_n3826_, new_n3827_, new_n3828_,
    new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_,
    new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_,
    new_n3841_, new_n3842_, new_n3844_, new_n3845_, new_n3846_, new_n3847_,
    new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_,
    new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_,
    new_n3860_, new_n3861_, new_n3863_, new_n3864_, new_n3865_, new_n3866_,
    new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_,
    new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_,
    new_n3879_, new_n3880_, new_n3882_, new_n3883_, new_n3884_, new_n3885_,
    new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3901_, new_n3902_, new_n3903_, new_n3904_,
    new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_,
    new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_,
    new_n3917_, new_n3918_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3939_, new_n3940_, new_n3941_, new_n3942_,
    new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_,
    new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_,
    new_n3955_, new_n3956_, new_n3958_, new_n3959_, new_n3960_, new_n3961_,
    new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_,
    new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_,
    new_n3974_, new_n3975_, new_n3977_, new_n3978_, new_n3979_, new_n3980_,
    new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_,
    new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_,
    new_n3993_, new_n3994_, new_n3996_, new_n3997_, new_n3998_, new_n3999_,
    new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_,
    new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_,
    new_n4012_, new_n4013_, new_n4015_, new_n4016_, new_n4017_, new_n4018_,
    new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_,
    new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_,
    new_n4031_, new_n4032_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4053_, new_n4054_, new_n4055_, new_n4056_,
    new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_,
    new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_,
    new_n4069_, new_n4070_, new_n4072_, new_n4073_, new_n4074_, new_n4075_,
    new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_,
    new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_,
    new_n4088_, new_n4089_, new_n4091_, new_n4092_, new_n4093_, new_n4094_,
    new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_,
    new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_,
    new_n4107_, new_n4108_, new_n4110_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4129_, new_n4130_, new_n4131_, new_n4132_,
    new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_,
    new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_,
    new_n4145_, new_n4146_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_,
    new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_,
    new_n4164_, new_n4165_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4186_, new_n4187_, new_n4188_, new_n4189_,
    new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_, new_n4195_,
    new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_, new_n4201_,
    new_n4202_, new_n4203_, new_n4205_, new_n4206_, new_n4207_, new_n4208_,
    new_n4209_, new_n4210_, new_n4211_, new_n4212_, new_n4213_, new_n4214_,
    new_n4215_, new_n4216_, new_n4217_, new_n4218_, new_n4219_, new_n4220_,
    new_n4221_, new_n4222_, new_n4224_, new_n4225_, new_n4226_, new_n4227_,
    new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_,
    new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_,
    new_n4240_, new_n4241_, new_n4243_, new_n4244_, new_n4245_, new_n4246_,
    new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_,
    new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_,
    new_n4259_, new_n4260_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4281_, new_n4282_, new_n4283_, new_n4284_,
    new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_,
    new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_,
    new_n4297_, new_n4298_, new_n4300_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4319_, new_n4320_, new_n4321_, new_n4322_,
    new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_, new_n4328_,
    new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_, new_n4334_,
    new_n4335_, new_n4336_, new_n4338_, new_n4339_, new_n4340_, new_n4341_,
    new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_,
    new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_,
    new_n4354_, new_n4355_, new_n4357_, new_n4358_, new_n4359_, new_n4360_,
    new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_,
    new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_,
    new_n4373_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_,
    new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_,
    new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_, new_n4436_,
    new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_, new_n4442_,
    new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_, new_n4448_,
    new_n4450_, new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_,
    new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_,
    new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_,
    new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_,
    new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_,
    new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_,
    new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_,
    new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_,
    new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_,
    new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_,
    new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_,
    new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_,
    new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_,
    new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_, new_n4575_,
    new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_,
    new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_,
    new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_,
    new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_,
    new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_,
    new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_,
    new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_,
    new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_,
    new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_,
    new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_,
    new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_,
    new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_,
    new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_,
    new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_,
    new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_,
    new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_,
    new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_,
    new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_,
    new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_,
    new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_,
    new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_,
    new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_,
    new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_,
    new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_,
    new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_,
    new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_,
    new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_,
    new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_,
    new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_,
    new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_,
    new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_,
    new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_,
    new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_,
    new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_,
    new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_,
    new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_,
    new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_,
    new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_,
    new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_,
    new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_,
    new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_,
    new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_,
    new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_,
    new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_,
    new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_,
    new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_,
    new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_,
    new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_,
    new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_,
    new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_,
    new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_,
    new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_,
    new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_,
    new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_,
    new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_,
    new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_,
    new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_,
    new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_,
    new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_,
    new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_,
    new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_,
    new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_,
    new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_,
    new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_,
    new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_,
    new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_,
    new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_,
    new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_,
    new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_,
    new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_,
    new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_,
    new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_,
    new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_,
    new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_,
    new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_,
    new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_,
    new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_,
    new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_,
    new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_,
    new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_,
    new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_,
    new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_,
    new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_,
    new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_,
    new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_,
    new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_,
    new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_,
    new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_,
    new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_,
    new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_,
    new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_,
    new_n5260_, new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_,
    new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_,
    new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_,
    new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_,
    new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_,
    new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_, new_n5348_,
    new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_, new_n5354_,
    new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_,
    new_n5362_, new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_,
    new_n5368_, new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_,
    new_n5374_, new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_,
    new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_,
    new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_,
    new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_,
    new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_,
    new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_,
    new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_,
    new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_,
    new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_,
    new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5437_,
    new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_,
    new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_,
    new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5455_, new_n5456_,
    new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_,
    new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_,
    new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5474_, new_n5475_,
    new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_,
    new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_,
    new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5493_, new_n5494_,
    new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_,
    new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_,
    new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5512_, new_n5513_,
    new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_,
    new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_,
    new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5531_, new_n5532_,
    new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_,
    new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_,
    new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5550_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5569_, new_n5570_,
    new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_,
    new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_,
    new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5588_, new_n5589_,
    new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_,
    new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_,
    new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5607_, new_n5608_,
    new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_,
    new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_,
    new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5626_, new_n5627_,
    new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5645_, new_n5646_,
    new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_,
    new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_,
    new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5664_, new_n5665_,
    new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_,
    new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_,
    new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5683_, new_n5684_,
    new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_,
    new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_,
    new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5702_, new_n5703_,
    new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_,
    new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_, new_n5715_,
    new_n5716_, new_n5717_, new_n5718_, new_n5719_, new_n5721_, new_n5722_,
    new_n5723_, new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_,
    new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_,
    new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5740_, new_n5741_,
    new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_,
    new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_,
    new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5759_, new_n5760_,
    new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_,
    new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_,
    new_n5773_, new_n5774_, new_n5775_, new_n5776_, n920, n925, n930, n935,
    n940, n945, n950, n955, n960, n965, n970, n975, n980, n985, n990, n995,
    n1000, n1005, n1010, n1015, n1020, n1025, n1030, n1035, n1040, n1045,
    n1050, n1055, n1060, n1065, n1070, n1075, n1080, n1085, n1090, n1095,
    n1100, n1105, n1110, n1115, n1120, n1125, n1130, n1135, n1140, n1145,
    n1150, n1155, n1160, n1165, n1170, n1175, n1180, n1185, n1190, n1195,
    n1200, n1205, n1210, n1215, n1220, n1225, n1230, n1235, n1240, n1245,
    n1250, n1255, n1260, n1265, n1270, n1275, n1280, n1285, n1290, n1295,
    n1300, n1305, n1310, n1315, n1320, n1325, n1330, n1335, n1340, n1345,
    n1350, n1355, n1360, n1365, n1370, n1375, n1380, n1385, n1390, n1395,
    n1400, n1405, n1410, n1415, n1420, n1425, n1430, n1435, n1440, n1445,
    n1450, n1455, n1460, n1465, n1470, n1475, n1480, n1485, n1490, n1495,
    n1500, n1505, n1510, n1515, n1520, n1525, n1530, n1535, n1540, n1545,
    n1550, n1555, n1560, n1565, n1570, n1575, n1580, n1585, n1590, n1595,
    n1600, n1605, n1610, n1615, n1620, n1625, n1630, n1635, n1640, n1645,
    n1650, n1655, n1660, n1665, n1670, n1675, n1680, n1685, n1690, n1695,
    n1700, n1705, n1710, n1715, n1720, n1725, n1730, n1735, n1740, n1745,
    n1750, n1755, n1760, n1765, n1770, n1775, n1780, n1785, n1790, n1795,
    n1800, n1805, n1810, n1815, n1820, n1825, n1830, n1835, n1840, n1845,
    n1850, n1855, n1860, n1865, n1870, n1875, n1880, n1885, n1890, n1895,
    n1900, n1905, n1910, n1915, n1920, n1925, n1930, n1935, n1940, n1945,
    n1950, n1955, n1960, n1965, n1970, n1975, n1980, n1985, n1990, n1995,
    n2000, n2005, n2010, n2015, n2020, n2025, n2030, n2035;
  assign new_n1132_ = ~\count<1>  & ~\count<0> ;
  assign new_n1133_ = ~\count<2>  & new_n1132_;
  assign new_n1134_ = \count<3>  & ~new_n1133_;
  assign new_n1135_1_ = ~\count<3>  & new_n1133_;
  assign new_n1136_ = ~new_n1134_ & ~new_n1135_1_;
  assign new_n1137_ = \count<1>  & \count<0> ;
  assign new_n1138_ = \count<2>  & new_n1137_;
  assign new_n1139_ = ~\count<3>  & new_n1138_;
  assign new_n1140_1_ = \count<3>  & ~new_n1138_;
  assign new_n1141_ = ~new_n1139_ & ~new_n1140_1_;
  assign new_n1142_ = ~\encrypt<0>  & \start<0> ;
  assign new_n1143_ = ~\encrypt<0>  & ~new_n1136_;
  assign new_n1144_ = \encrypt<0>  & ~new_n1141_;
  assign new_n1145_1_ = ~new_n1143_ & ~new_n1144_;
  assign new_n1146_ = ~\start<0>  & ~new_n1145_1_;
  assign \new_count<3>  = new_n1142_ | new_n1146_;
  assign new_n1148_ = \count<2>  & ~new_n1132_;
  assign new_n1149_ = ~new_n1133_ & ~new_n1148_;
  assign new_n1150_1_ = ~\count<2>  & new_n1137_;
  assign new_n1151_ = \count<2>  & ~new_n1137_;
  assign new_n1152_ = ~new_n1150_1_ & ~new_n1151_;
  assign new_n1153_ = ~\encrypt<0>  & ~new_n1149_;
  assign new_n1154_ = \encrypt<0>  & ~new_n1152_;
  assign new_n1155_1_ = ~new_n1153_ & ~new_n1154_;
  assign new_n1156_ = ~\start<0>  & ~new_n1155_1_;
  assign \new_count<2>  = new_n1142_ | new_n1156_;
  assign new_n1158_ = ~new_n1132_ & ~new_n1137_;
  assign new_n1159_ = ~\count<1>  & \count<0> ;
  assign new_n1160_1_ = \count<1>  & ~\count<0> ;
  assign new_n1161_ = ~new_n1159_ & ~new_n1160_1_;
  assign new_n1162_ = ~\encrypt<0>  & ~new_n1158_;
  assign new_n1163_ = \encrypt<0>  & ~new_n1161_;
  assign new_n1164_ = ~new_n1162_ & ~new_n1163_;
  assign new_n1165_1_ = ~\start<0>  & ~new_n1164_;
  assign \new_count<1>  = new_n1142_ | new_n1165_1_;
  assign new_n1167_ = ~\encrypt<0>  & ~\count<0> ;
  assign new_n1168_ = \encrypt<0>  & ~\count<0> ;
  assign new_n1169_ = ~new_n1167_ & ~new_n1168_;
  assign new_n1170_1_ = ~\start<0>  & ~new_n1169_;
  assign \new_count<0>  = new_n1142_ | new_n1170_1_;
  assign new_n1172_ = \encrypt<0>  & \count<0> ;
  assign new_n1173_ = \count<3>  & \count<2> ;
  assign new_n1174_ = \count<1>  & new_n1173_;
  assign new_n1175_1_ = new_n1172_ & new_n1174_;
  assign new_n1176_ = ~\count<3>  & ~\count<2> ;
  assign new_n1177_ = ~\count<1>  & new_n1176_;
  assign new_n1178_ = new_n1167_ & new_n1177_;
  assign new_n1179_ = ~new_n1175_1_ & ~new_n1178_;
  assign \data_ready<0>  = ~\start<0>  & ~new_n1179_;
  assign new_n1181_ = ~new_n1174_ & ~new_n1177_;
  assign new_n1182_ = \count<0>  & ~new_n1181_;
  assign new_n1183_ = ~\count<2>  & ~\count<1> ;
  assign new_n1184_ = ~\count<0>  & new_n1183_;
  assign new_n1185_1_ = ~new_n1182_ & ~new_n1184_;
  assign new_n1186_ = ~\count<0>  & ~new_n1181_;
  assign new_n1187_ = ~\count<3>  & \count<2> ;
  assign new_n1188_ = new_n1137_ & new_n1187_;
  assign new_n1189_ = ~new_n1186_ & ~new_n1188_;
  assign new_n1190_1_ = \key<227>  & ~\encrypt<0> ;
  assign new_n1191_ = \key<56>  & \encrypt<0> ;
  assign new_n1192_ = ~new_n1190_1_ & ~new_n1191_;
  assign new_n1193_ = \start<0>  & ~new_n1192_;
  assign new_n1194_ = ~\C<111>  & ~\D<111> ;
  assign new_n1195_1_ = \C<111>  & \D<111> ;
  assign new_n1196_ = ~new_n1194_ & ~new_n1195_1_;
  assign new_n1197_ = ~new_n1185_1_ & ~new_n1196_;
  assign new_n1198_ = new_n1185_1_ & ~new_n1194_;
  assign new_n1199_ = ~new_n1197_ & ~new_n1198_;
  assign new_n1200_1_ = ~\encrypt<0>  & ~new_n1199_;
  assign new_n1201_ = \D<111>  & ~new_n1189_;
  assign new_n1202_ = ~\D<111>  & new_n1189_;
  assign new_n1203_ = ~new_n1201_ & ~new_n1202_;
  assign new_n1204_ = \C<111>  & ~new_n1203_;
  assign new_n1205_1_ = \D<111>  & new_n1189_;
  assign new_n1206_ = ~\C<111>  & new_n1205_1_;
  assign new_n1207_ = ~new_n1204_ & ~new_n1206_;
  assign new_n1208_ = \encrypt<0>  & ~new_n1207_;
  assign new_n1209_ = ~new_n1200_1_ & ~new_n1208_;
  assign new_n1210_1_ = ~\start<0>  & ~new_n1209_;
  assign n920 = new_n1193_ | new_n1210_1_;
  assign new_n1212_ = \key<235>  & ~\encrypt<0> ;
  assign new_n1213_ = \key<227>  & \encrypt<0> ;
  assign new_n1214_ = ~new_n1212_ & ~new_n1213_;
  assign new_n1215_1_ = \start<0>  & ~new_n1214_;
  assign new_n1216_ = ~\C<110>  & ~\D<110> ;
  assign new_n1217_ = \C<110>  & \D<110> ;
  assign new_n1218_ = ~new_n1216_ & ~new_n1217_;
  assign new_n1219_ = ~new_n1185_1_ & ~new_n1218_;
  assign new_n1220_1_ = new_n1185_1_ & ~new_n1216_;
  assign new_n1221_ = ~new_n1219_ & ~new_n1220_1_;
  assign new_n1222_ = ~\encrypt<0>  & ~new_n1221_;
  assign new_n1223_ = \D<110>  & ~new_n1189_;
  assign new_n1224_ = ~\D<110>  & new_n1189_;
  assign new_n1225_1_ = ~new_n1223_ & ~new_n1224_;
  assign new_n1226_ = \C<110>  & ~new_n1225_1_;
  assign new_n1227_ = \D<110>  & new_n1189_;
  assign new_n1228_ = ~\C<110>  & new_n1227_;
  assign new_n1229_ = ~new_n1226_ & ~new_n1228_;
  assign new_n1230_1_ = \encrypt<0>  & ~new_n1229_;
  assign new_n1231_ = ~new_n1222_ & ~new_n1230_1_;
  assign new_n1232_ = ~\start<0>  & ~new_n1231_;
  assign n925 = new_n1215_1_ | new_n1232_;
  assign new_n1234_ = \key<243>  & ~\encrypt<0> ;
  assign new_n1235_1_ = \key<235>  & \encrypt<0> ;
  assign new_n1236_ = ~new_n1234_ & ~new_n1235_1_;
  assign new_n1237_ = \start<0>  & ~new_n1236_;
  assign new_n1238_ = ~\C<109>  & ~\D<109> ;
  assign new_n1239_ = \C<109>  & \D<109> ;
  assign new_n1240_1_ = ~new_n1238_ & ~new_n1239_;
  assign new_n1241_ = ~new_n1185_1_ & ~new_n1240_1_;
  assign new_n1242_ = new_n1185_1_ & ~new_n1238_;
  assign new_n1243_ = ~new_n1241_ & ~new_n1242_;
  assign new_n1244_ = ~\encrypt<0>  & ~new_n1243_;
  assign new_n1245_1_ = \D<109>  & ~new_n1189_;
  assign new_n1246_ = ~\D<109>  & new_n1189_;
  assign new_n1247_ = ~new_n1245_1_ & ~new_n1246_;
  assign new_n1248_ = \C<109>  & ~new_n1247_;
  assign new_n1249_ = \D<109>  & new_n1189_;
  assign new_n1250_1_ = ~\C<109>  & new_n1249_;
  assign new_n1251_ = ~new_n1248_ & ~new_n1250_1_;
  assign new_n1252_ = \encrypt<0>  & ~new_n1251_;
  assign new_n1253_ = ~new_n1244_ & ~new_n1252_;
  assign new_n1254_ = ~\start<0>  & ~new_n1253_;
  assign n930 = new_n1237_ | new_n1254_;
  assign new_n1256_ = \key<251>  & ~\encrypt<0> ;
  assign new_n1257_ = \key<243>  & \encrypt<0> ;
  assign new_n1258_ = ~new_n1256_ & ~new_n1257_;
  assign new_n1259_ = \start<0>  & ~new_n1258_;
  assign new_n1260_1_ = ~\C<108>  & ~\D<108> ;
  assign new_n1261_ = \C<108>  & \D<108> ;
  assign new_n1262_ = ~new_n1260_1_ & ~new_n1261_;
  assign new_n1263_ = ~new_n1185_1_ & ~new_n1262_;
  assign new_n1264_ = new_n1185_1_ & ~new_n1260_1_;
  assign new_n1265_1_ = ~new_n1263_ & ~new_n1264_;
  assign new_n1266_ = ~\encrypt<0>  & ~new_n1265_1_;
  assign new_n1267_ = \D<108>  & ~new_n1189_;
  assign new_n1268_ = ~\D<108>  & new_n1189_;
  assign new_n1269_ = ~new_n1267_ & ~new_n1268_;
  assign new_n1270_1_ = \C<108>  & ~new_n1269_;
  assign new_n1271_ = \D<108>  & new_n1189_;
  assign new_n1272_ = ~\C<108>  & new_n1271_;
  assign new_n1273_ = ~new_n1270_1_ & ~new_n1272_;
  assign new_n1274_ = \encrypt<0>  & ~new_n1273_;
  assign new_n1275_1_ = ~new_n1266_ & ~new_n1274_;
  assign new_n1276_ = ~\start<0>  & ~new_n1275_1_;
  assign n935 = new_n1259_ | new_n1276_;
  assign new_n1278_ = \key<194>  & ~\encrypt<0> ;
  assign new_n1279_ = \key<251>  & \encrypt<0> ;
  assign new_n1280_1_ = ~new_n1278_ & ~new_n1279_;
  assign new_n1281_ = \start<0>  & ~new_n1280_1_;
  assign new_n1282_ = ~\C<107>  & ~\D<107> ;
  assign new_n1283_ = \C<107>  & \D<107> ;
  assign new_n1284_ = ~new_n1282_ & ~new_n1283_;
  assign new_n1285_1_ = ~new_n1185_1_ & ~new_n1284_;
  assign new_n1286_ = new_n1185_1_ & ~new_n1282_;
  assign new_n1287_ = ~new_n1285_1_ & ~new_n1286_;
  assign new_n1288_ = ~\encrypt<0>  & ~new_n1287_;
  assign new_n1289_ = \D<107>  & ~new_n1189_;
  assign new_n1290_1_ = ~\D<107>  & new_n1189_;
  assign new_n1291_ = ~new_n1289_ & ~new_n1290_1_;
  assign new_n1292_ = \C<107>  & ~new_n1291_;
  assign new_n1293_ = \D<107>  & new_n1189_;
  assign new_n1294_ = ~\C<107>  & new_n1293_;
  assign new_n1295_1_ = ~new_n1292_ & ~new_n1294_;
  assign new_n1296_ = \encrypt<0>  & ~new_n1295_1_;
  assign new_n1297_ = ~new_n1288_ & ~new_n1296_;
  assign new_n1298_ = ~\start<0>  & ~new_n1297_;
  assign n940 = new_n1281_ | new_n1298_;
  assign new_n1300_1_ = \key<202>  & ~\encrypt<0> ;
  assign new_n1301_ = \key<194>  & \encrypt<0> ;
  assign new_n1302_ = ~new_n1300_1_ & ~new_n1301_;
  assign new_n1303_ = \start<0>  & ~new_n1302_;
  assign new_n1304_ = ~\C<106>  & ~\D<106> ;
  assign new_n1305_1_ = \C<106>  & \D<106> ;
  assign new_n1306_ = ~new_n1304_ & ~new_n1305_1_;
  assign new_n1307_ = ~new_n1185_1_ & ~new_n1306_;
  assign new_n1308_ = new_n1185_1_ & ~new_n1304_;
  assign new_n1309_ = ~new_n1307_ & ~new_n1308_;
  assign new_n1310_1_ = ~\encrypt<0>  & ~new_n1309_;
  assign new_n1311_ = \D<106>  & ~new_n1189_;
  assign new_n1312_ = ~\D<106>  & new_n1189_;
  assign new_n1313_ = ~new_n1311_ & ~new_n1312_;
  assign new_n1314_ = \C<106>  & ~new_n1313_;
  assign new_n1315_1_ = \D<106>  & new_n1189_;
  assign new_n1316_ = ~\C<106>  & new_n1315_1_;
  assign new_n1317_ = ~new_n1314_ & ~new_n1316_;
  assign new_n1318_ = \encrypt<0>  & ~new_n1317_;
  assign new_n1319_ = ~new_n1310_1_ & ~new_n1318_;
  assign new_n1320_1_ = ~\start<0>  & ~new_n1319_;
  assign n945 = new_n1303_ | new_n1320_1_;
  assign new_n1322_ = \key<210>  & ~\encrypt<0> ;
  assign new_n1323_ = \key<202>  & \encrypt<0> ;
  assign new_n1324_ = ~new_n1322_ & ~new_n1323_;
  assign new_n1325_1_ = \start<0>  & ~new_n1324_;
  assign new_n1326_ = ~\C<105>  & ~\D<105> ;
  assign new_n1327_ = \C<105>  & \D<105> ;
  assign new_n1328_ = ~new_n1326_ & ~new_n1327_;
  assign new_n1329_ = ~new_n1185_1_ & ~new_n1328_;
  assign new_n1330_1_ = new_n1185_1_ & ~new_n1326_;
  assign new_n1331_ = ~new_n1329_ & ~new_n1330_1_;
  assign new_n1332_ = ~\encrypt<0>  & ~new_n1331_;
  assign new_n1333_ = \D<105>  & ~new_n1189_;
  assign new_n1334_ = ~\D<105>  & new_n1189_;
  assign new_n1335_1_ = ~new_n1333_ & ~new_n1334_;
  assign new_n1336_ = \C<105>  & ~new_n1335_1_;
  assign new_n1337_ = \D<105>  & new_n1189_;
  assign new_n1338_ = ~\C<105>  & new_n1337_;
  assign new_n1339_ = ~new_n1336_ & ~new_n1338_;
  assign new_n1340_1_ = \encrypt<0>  & ~new_n1339_;
  assign new_n1341_ = ~new_n1332_ & ~new_n1340_1_;
  assign new_n1342_ = ~\start<0>  & ~new_n1341_;
  assign n950 = new_n1325_1_ | new_n1342_;
  assign new_n1344_ = \key<218>  & ~\encrypt<0> ;
  assign new_n1345_1_ = \key<210>  & \encrypt<0> ;
  assign new_n1346_ = ~new_n1344_ & ~new_n1345_1_;
  assign new_n1347_ = \start<0>  & ~new_n1346_;
  assign new_n1348_ = ~\C<104>  & ~\D<104> ;
  assign new_n1349_ = \C<104>  & \D<104> ;
  assign new_n1350_1_ = ~new_n1348_ & ~new_n1349_;
  assign new_n1351_ = ~new_n1185_1_ & ~new_n1350_1_;
  assign new_n1352_ = new_n1185_1_ & ~new_n1348_;
  assign new_n1353_ = ~new_n1351_ & ~new_n1352_;
  assign new_n1354_ = ~\encrypt<0>  & ~new_n1353_;
  assign new_n1355_1_ = \D<104>  & ~new_n1189_;
  assign new_n1356_ = ~\D<104>  & new_n1189_;
  assign new_n1357_ = ~new_n1355_1_ & ~new_n1356_;
  assign new_n1358_ = \C<104>  & ~new_n1357_;
  assign new_n1359_ = \D<104>  & new_n1189_;
  assign new_n1360_1_ = ~\C<104>  & new_n1359_;
  assign new_n1361_ = ~new_n1358_ & ~new_n1360_1_;
  assign new_n1362_ = \encrypt<0>  & ~new_n1361_;
  assign new_n1363_ = ~new_n1354_ & ~new_n1362_;
  assign new_n1364_ = ~\start<0>  & ~new_n1363_;
  assign n955 = new_n1347_ | new_n1364_;
  assign new_n1366_ = \key<226>  & ~\encrypt<0> ;
  assign new_n1367_ = \key<218>  & \encrypt<0> ;
  assign new_n1368_ = ~new_n1366_ & ~new_n1367_;
  assign new_n1369_ = \start<0>  & ~new_n1368_;
  assign new_n1370_1_ = ~\C<103>  & ~\D<103> ;
  assign new_n1371_ = \C<103>  & \D<103> ;
  assign new_n1372_ = ~new_n1370_1_ & ~new_n1371_;
  assign new_n1373_ = ~new_n1185_1_ & ~new_n1372_;
  assign new_n1374_ = new_n1185_1_ & ~new_n1370_1_;
  assign new_n1375_1_ = ~new_n1373_ & ~new_n1374_;
  assign new_n1376_ = ~\encrypt<0>  & ~new_n1375_1_;
  assign new_n1377_ = \D<103>  & ~new_n1189_;
  assign new_n1378_ = ~\D<103>  & new_n1189_;
  assign new_n1379_ = ~new_n1377_ & ~new_n1378_;
  assign new_n1380_1_ = \C<103>  & ~new_n1379_;
  assign new_n1381_ = \D<103>  & new_n1189_;
  assign new_n1382_ = ~\C<103>  & new_n1381_;
  assign new_n1383_ = ~new_n1380_1_ & ~new_n1382_;
  assign new_n1384_ = \encrypt<0>  & ~new_n1383_;
  assign new_n1385_1_ = ~new_n1376_ & ~new_n1384_;
  assign new_n1386_ = ~\start<0>  & ~new_n1385_1_;
  assign n960 = new_n1369_ | new_n1386_;
  assign new_n1388_ = \key<234>  & ~\encrypt<0> ;
  assign new_n1389_ = \key<226>  & \encrypt<0> ;
  assign new_n1390_1_ = ~new_n1388_ & ~new_n1389_;
  assign new_n1391_ = \start<0>  & ~new_n1390_1_;
  assign new_n1392_ = ~\C<102>  & ~\D<102> ;
  assign new_n1393_ = \C<102>  & \D<102> ;
  assign new_n1394_ = ~new_n1392_ & ~new_n1393_;
  assign new_n1395_1_ = ~new_n1185_1_ & ~new_n1394_;
  assign new_n1396_ = new_n1185_1_ & ~new_n1392_;
  assign new_n1397_ = ~new_n1395_1_ & ~new_n1396_;
  assign new_n1398_ = ~\encrypt<0>  & ~new_n1397_;
  assign new_n1399_ = \D<102>  & ~new_n1189_;
  assign new_n1400_1_ = ~\D<102>  & new_n1189_;
  assign new_n1401_ = ~new_n1399_ & ~new_n1400_1_;
  assign new_n1402_ = \C<102>  & ~new_n1401_;
  assign new_n1403_ = \D<102>  & new_n1189_;
  assign new_n1404_ = ~\C<102>  & new_n1403_;
  assign new_n1405_1_ = ~new_n1402_ & ~new_n1404_;
  assign new_n1406_ = \encrypt<0>  & ~new_n1405_1_;
  assign new_n1407_ = ~new_n1398_ & ~new_n1406_;
  assign new_n1408_ = ~\start<0>  & ~new_n1407_;
  assign n965 = new_n1391_ | new_n1408_;
  assign new_n1410_1_ = \key<242>  & ~\encrypt<0> ;
  assign new_n1411_ = \key<234>  & \encrypt<0> ;
  assign new_n1412_ = ~new_n1410_1_ & ~new_n1411_;
  assign new_n1413_ = \start<0>  & ~new_n1412_;
  assign new_n1414_ = ~\C<101>  & ~\D<101> ;
  assign new_n1415_1_ = \C<101>  & \D<101> ;
  assign new_n1416_ = ~new_n1414_ & ~new_n1415_1_;
  assign new_n1417_ = ~new_n1185_1_ & ~new_n1416_;
  assign new_n1418_ = new_n1185_1_ & ~new_n1414_;
  assign new_n1419_ = ~new_n1417_ & ~new_n1418_;
  assign new_n1420_1_ = ~\encrypt<0>  & ~new_n1419_;
  assign new_n1421_ = \D<101>  & ~new_n1189_;
  assign new_n1422_ = ~\D<101>  & new_n1189_;
  assign new_n1423_ = ~new_n1421_ & ~new_n1422_;
  assign new_n1424_ = \C<101>  & ~new_n1423_;
  assign new_n1425_1_ = \D<101>  & new_n1189_;
  assign new_n1426_ = ~\C<101>  & new_n1425_1_;
  assign new_n1427_ = ~new_n1424_ & ~new_n1426_;
  assign new_n1428_ = \encrypt<0>  & ~new_n1427_;
  assign new_n1429_ = ~new_n1420_1_ & ~new_n1428_;
  assign new_n1430_1_ = ~\start<0>  & ~new_n1429_;
  assign n970 = new_n1413_ | new_n1430_1_;
  assign new_n1432_ = \key<250>  & ~\encrypt<0> ;
  assign new_n1433_ = \key<242>  & \encrypt<0> ;
  assign new_n1434_ = ~new_n1432_ & ~new_n1433_;
  assign new_n1435_1_ = \start<0>  & ~new_n1434_;
  assign new_n1436_ = ~\C<100>  & ~\D<100> ;
  assign new_n1437_ = \C<100>  & \D<100> ;
  assign new_n1438_ = ~new_n1436_ & ~new_n1437_;
  assign new_n1439_ = ~new_n1185_1_ & ~new_n1438_;
  assign new_n1440_1_ = new_n1185_1_ & ~new_n1436_;
  assign new_n1441_ = ~new_n1439_ & ~new_n1440_1_;
  assign new_n1442_ = ~\encrypt<0>  & ~new_n1441_;
  assign new_n1443_ = \D<100>  & ~new_n1189_;
  assign new_n1444_ = ~\D<100>  & new_n1189_;
  assign new_n1445_1_ = ~new_n1443_ & ~new_n1444_;
  assign new_n1446_ = \C<100>  & ~new_n1445_1_;
  assign new_n1447_ = \D<100>  & new_n1189_;
  assign new_n1448_ = ~\C<100>  & new_n1447_;
  assign new_n1449_ = ~new_n1446_ & ~new_n1448_;
  assign new_n1450_1_ = \encrypt<0>  & ~new_n1449_;
  assign new_n1451_ = ~new_n1442_ & ~new_n1450_1_;
  assign new_n1452_ = ~\start<0>  & ~new_n1451_;
  assign n975 = new_n1435_1_ | new_n1452_;
  assign new_n1454_ = \key<193>  & ~\encrypt<0> ;
  assign new_n1455_1_ = \key<250>  & \encrypt<0> ;
  assign new_n1456_ = ~new_n1454_ & ~new_n1455_1_;
  assign new_n1457_ = \start<0>  & ~new_n1456_;
  assign new_n1458_ = ~\C<99>  & ~\D<99> ;
  assign new_n1459_ = \C<99>  & \D<99> ;
  assign new_n1460_1_ = ~new_n1458_ & ~new_n1459_;
  assign new_n1461_ = ~new_n1185_1_ & ~new_n1460_1_;
  assign new_n1462_ = new_n1185_1_ & ~new_n1458_;
  assign new_n1463_ = ~new_n1461_ & ~new_n1462_;
  assign new_n1464_ = ~\encrypt<0>  & ~new_n1463_;
  assign new_n1465_1_ = \D<99>  & ~new_n1189_;
  assign new_n1466_ = ~\D<99>  & new_n1189_;
  assign new_n1467_ = ~new_n1465_1_ & ~new_n1466_;
  assign new_n1468_ = \C<99>  & ~new_n1467_;
  assign new_n1469_ = \D<99>  & new_n1189_;
  assign new_n1470_1_ = ~\C<99>  & new_n1469_;
  assign new_n1471_ = ~new_n1468_ & ~new_n1470_1_;
  assign new_n1472_ = \encrypt<0>  & ~new_n1471_;
  assign new_n1473_ = ~new_n1464_ & ~new_n1472_;
  assign new_n1474_ = ~\start<0>  & ~new_n1473_;
  assign n980 = new_n1457_ | new_n1474_;
  assign new_n1476_ = \key<201>  & ~\encrypt<0> ;
  assign new_n1477_ = \key<193>  & \encrypt<0> ;
  assign new_n1478_ = ~new_n1476_ & ~new_n1477_;
  assign new_n1479_ = \start<0>  & ~new_n1478_;
  assign new_n1480_1_ = ~\C<98>  & ~\D<98> ;
  assign new_n1481_ = \C<98>  & \D<98> ;
  assign new_n1482_ = ~new_n1480_1_ & ~new_n1481_;
  assign new_n1483_ = ~new_n1185_1_ & ~new_n1482_;
  assign new_n1484_ = new_n1185_1_ & ~new_n1480_1_;
  assign new_n1485_1_ = ~new_n1483_ & ~new_n1484_;
  assign new_n1486_ = ~\encrypt<0>  & ~new_n1485_1_;
  assign new_n1487_ = \D<98>  & ~new_n1189_;
  assign new_n1488_ = ~\D<98>  & new_n1189_;
  assign new_n1489_ = ~new_n1487_ & ~new_n1488_;
  assign new_n1490_1_ = \C<98>  & ~new_n1489_;
  assign new_n1491_ = \D<98>  & new_n1189_;
  assign new_n1492_ = ~\C<98>  & new_n1491_;
  assign new_n1493_ = ~new_n1490_1_ & ~new_n1492_;
  assign new_n1494_ = \encrypt<0>  & ~new_n1493_;
  assign new_n1495_1_ = ~new_n1486_ & ~new_n1494_;
  assign new_n1496_ = ~\start<0>  & ~new_n1495_1_;
  assign n985 = new_n1479_ | new_n1496_;
  assign new_n1498_ = \key<209>  & ~\encrypt<0> ;
  assign new_n1499_ = \key<201>  & \encrypt<0> ;
  assign new_n1500_1_ = ~new_n1498_ & ~new_n1499_;
  assign new_n1501_ = \start<0>  & ~new_n1500_1_;
  assign new_n1502_ = ~\C<97>  & ~\D<97> ;
  assign new_n1503_ = \C<97>  & \D<97> ;
  assign new_n1504_ = ~new_n1502_ & ~new_n1503_;
  assign new_n1505_1_ = ~new_n1185_1_ & ~new_n1504_;
  assign new_n1506_ = new_n1185_1_ & ~new_n1502_;
  assign new_n1507_ = ~new_n1505_1_ & ~new_n1506_;
  assign new_n1508_ = ~\encrypt<0>  & ~new_n1507_;
  assign new_n1509_ = \D<97>  & ~new_n1189_;
  assign new_n1510_1_ = ~\D<97>  & new_n1189_;
  assign new_n1511_ = ~new_n1509_ & ~new_n1510_1_;
  assign new_n1512_ = \C<97>  & ~new_n1511_;
  assign new_n1513_ = \D<97>  & new_n1189_;
  assign new_n1514_ = ~\C<97>  & new_n1513_;
  assign new_n1515_1_ = ~new_n1512_ & ~new_n1514_;
  assign new_n1516_ = \encrypt<0>  & ~new_n1515_1_;
  assign new_n1517_ = ~new_n1508_ & ~new_n1516_;
  assign new_n1518_ = ~\start<0>  & ~new_n1517_;
  assign n990 = new_n1501_ | new_n1518_;
  assign new_n1520_1_ = \key<217>  & ~\encrypt<0> ;
  assign new_n1521_ = \key<209>  & \encrypt<0> ;
  assign new_n1522_ = ~new_n1520_1_ & ~new_n1521_;
  assign new_n1523_ = \start<0>  & ~new_n1522_;
  assign new_n1524_ = ~\C<96>  & ~\D<96> ;
  assign new_n1525_1_ = \C<96>  & \D<96> ;
  assign new_n1526_ = ~new_n1524_ & ~new_n1525_1_;
  assign new_n1527_ = ~new_n1185_1_ & ~new_n1526_;
  assign new_n1528_ = new_n1185_1_ & ~new_n1524_;
  assign new_n1529_ = ~new_n1527_ & ~new_n1528_;
  assign new_n1530_1_ = ~\encrypt<0>  & ~new_n1529_;
  assign new_n1531_ = \D<96>  & ~new_n1189_;
  assign new_n1532_ = ~\D<96>  & new_n1189_;
  assign new_n1533_ = ~new_n1531_ & ~new_n1532_;
  assign new_n1534_ = \C<96>  & ~new_n1533_;
  assign new_n1535_1_ = \D<96>  & new_n1189_;
  assign new_n1536_ = ~\C<96>  & new_n1535_1_;
  assign new_n1537_ = ~new_n1534_ & ~new_n1536_;
  assign new_n1538_ = \encrypt<0>  & ~new_n1537_;
  assign new_n1539_ = ~new_n1530_1_ & ~new_n1538_;
  assign new_n1540_1_ = ~\start<0>  & ~new_n1539_;
  assign n995 = new_n1523_ | new_n1540_1_;
  assign new_n1542_ = \key<225>  & ~\encrypt<0> ;
  assign new_n1543_ = \key<217>  & \encrypt<0> ;
  assign new_n1544_ = ~new_n1542_ & ~new_n1543_;
  assign new_n1545_1_ = \start<0>  & ~new_n1544_;
  assign new_n1546_ = ~\C<95>  & ~\D<95> ;
  assign new_n1547_ = \C<95>  & \D<95> ;
  assign new_n1548_ = ~new_n1546_ & ~new_n1547_;
  assign new_n1549_ = ~new_n1185_1_ & ~new_n1548_;
  assign new_n1550_1_ = new_n1185_1_ & ~new_n1546_;
  assign new_n1551_ = ~new_n1549_ & ~new_n1550_1_;
  assign new_n1552_ = ~\encrypt<0>  & ~new_n1551_;
  assign new_n1553_ = \D<95>  & ~new_n1189_;
  assign new_n1554_ = ~\D<95>  & new_n1189_;
  assign new_n1555_1_ = ~new_n1553_ & ~new_n1554_;
  assign new_n1556_ = \C<95>  & ~new_n1555_1_;
  assign new_n1557_ = \D<95>  & new_n1189_;
  assign new_n1558_ = ~\C<95>  & new_n1557_;
  assign new_n1559_ = ~new_n1556_ & ~new_n1558_;
  assign new_n1560_1_ = \encrypt<0>  & ~new_n1559_;
  assign new_n1561_ = ~new_n1552_ & ~new_n1560_1_;
  assign new_n1562_ = ~\start<0>  & ~new_n1561_;
  assign n1000 = new_n1545_1_ | new_n1562_;
  assign new_n1564_ = \key<233>  & ~\encrypt<0> ;
  assign new_n1565_1_ = \key<225>  & \encrypt<0> ;
  assign new_n1566_ = ~new_n1564_ & ~new_n1565_1_;
  assign new_n1567_ = \start<0>  & ~new_n1566_;
  assign new_n1568_ = ~\C<94>  & ~\D<94> ;
  assign new_n1569_ = \C<94>  & \D<94> ;
  assign new_n1570_1_ = ~new_n1568_ & ~new_n1569_;
  assign new_n1571_ = ~new_n1185_1_ & ~new_n1570_1_;
  assign new_n1572_ = new_n1185_1_ & ~new_n1568_;
  assign new_n1573_ = ~new_n1571_ & ~new_n1572_;
  assign new_n1574_ = ~\encrypt<0>  & ~new_n1573_;
  assign new_n1575_1_ = \D<94>  & ~new_n1189_;
  assign new_n1576_ = ~\D<94>  & new_n1189_;
  assign new_n1577_ = ~new_n1575_1_ & ~new_n1576_;
  assign new_n1578_ = \C<94>  & ~new_n1577_;
  assign new_n1579_ = \D<94>  & new_n1189_;
  assign new_n1580_1_ = ~\C<94>  & new_n1579_;
  assign new_n1581_ = ~new_n1578_ & ~new_n1580_1_;
  assign new_n1582_ = \encrypt<0>  & ~new_n1581_;
  assign new_n1583_ = ~new_n1574_ & ~new_n1582_;
  assign new_n1584_ = ~\start<0>  & ~new_n1583_;
  assign n1005 = new_n1567_ | new_n1584_;
  assign new_n1586_ = \key<241>  & ~\encrypt<0> ;
  assign new_n1587_ = \key<233>  & \encrypt<0> ;
  assign new_n1588_ = ~new_n1586_ & ~new_n1587_;
  assign new_n1589_ = \start<0>  & ~new_n1588_;
  assign new_n1590_1_ = ~\C<93>  & ~\D<93> ;
  assign new_n1591_ = \C<93>  & \D<93> ;
  assign new_n1592_ = ~new_n1590_1_ & ~new_n1591_;
  assign new_n1593_ = ~new_n1185_1_ & ~new_n1592_;
  assign new_n1594_ = new_n1185_1_ & ~new_n1590_1_;
  assign new_n1595_1_ = ~new_n1593_ & ~new_n1594_;
  assign new_n1596_ = ~\encrypt<0>  & ~new_n1595_1_;
  assign new_n1597_ = \D<93>  & ~new_n1189_;
  assign new_n1598_ = ~\D<93>  & new_n1189_;
  assign new_n1599_ = ~new_n1597_ & ~new_n1598_;
  assign new_n1600_1_ = \C<93>  & ~new_n1599_;
  assign new_n1601_ = \D<93>  & new_n1189_;
  assign new_n1602_ = ~\C<93>  & new_n1601_;
  assign new_n1603_ = ~new_n1600_1_ & ~new_n1602_;
  assign new_n1604_ = \encrypt<0>  & ~new_n1603_;
  assign new_n1605_1_ = ~new_n1596_ & ~new_n1604_;
  assign new_n1606_ = ~\start<0>  & ~new_n1605_1_;
  assign n1010 = new_n1589_ | new_n1606_;
  assign new_n1608_ = \key<249>  & ~\encrypt<0> ;
  assign new_n1609_ = \key<241>  & \encrypt<0> ;
  assign new_n1610_1_ = ~new_n1608_ & ~new_n1609_;
  assign new_n1611_ = \start<0>  & ~new_n1610_1_;
  assign new_n1612_ = ~\C<92>  & ~\D<92> ;
  assign new_n1613_ = \C<92>  & \D<92> ;
  assign new_n1614_ = ~new_n1612_ & ~new_n1613_;
  assign new_n1615_1_ = ~new_n1185_1_ & ~new_n1614_;
  assign new_n1616_ = new_n1185_1_ & ~new_n1612_;
  assign new_n1617_ = ~new_n1615_1_ & ~new_n1616_;
  assign new_n1618_ = ~\encrypt<0>  & ~new_n1617_;
  assign new_n1619_ = \D<92>  & ~new_n1189_;
  assign new_n1620_1_ = ~\D<92>  & new_n1189_;
  assign new_n1621_ = ~new_n1619_ & ~new_n1620_1_;
  assign new_n1622_ = \C<92>  & ~new_n1621_;
  assign new_n1623_ = \D<92>  & new_n1189_;
  assign new_n1624_ = ~\C<92>  & new_n1623_;
  assign new_n1625_1_ = ~new_n1622_ & ~new_n1624_;
  assign new_n1626_ = \encrypt<0>  & ~new_n1625_1_;
  assign new_n1627_ = ~new_n1618_ & ~new_n1626_;
  assign new_n1628_ = ~\start<0>  & ~new_n1627_;
  assign n1015 = new_n1611_ | new_n1628_;
  assign new_n1630_1_ = \key<192>  & ~\encrypt<0> ;
  assign new_n1631_ = \key<249>  & \encrypt<0> ;
  assign new_n1632_ = ~new_n1630_1_ & ~new_n1631_;
  assign new_n1633_ = \start<0>  & ~new_n1632_;
  assign new_n1634_ = ~\C<91>  & ~\D<91> ;
  assign new_n1635_1_ = \C<91>  & \D<91> ;
  assign new_n1636_ = ~new_n1634_ & ~new_n1635_1_;
  assign new_n1637_ = ~new_n1185_1_ & ~new_n1636_;
  assign new_n1638_ = new_n1185_1_ & ~new_n1634_;
  assign new_n1639_ = ~new_n1637_ & ~new_n1638_;
  assign new_n1640_1_ = ~\encrypt<0>  & ~new_n1639_;
  assign new_n1641_ = \D<91>  & ~new_n1189_;
  assign new_n1642_ = ~\D<91>  & new_n1189_;
  assign new_n1643_ = ~new_n1641_ & ~new_n1642_;
  assign new_n1644_ = \C<91>  & ~new_n1643_;
  assign new_n1645_1_ = \D<91>  & new_n1189_;
  assign new_n1646_ = ~\C<91>  & new_n1645_1_;
  assign new_n1647_ = ~new_n1644_ & ~new_n1646_;
  assign new_n1648_ = \encrypt<0>  & ~new_n1647_;
  assign new_n1649_ = ~new_n1640_1_ & ~new_n1648_;
  assign new_n1650_1_ = ~\start<0>  & ~new_n1649_;
  assign n1020 = new_n1633_ | new_n1650_1_;
  assign new_n1652_ = \key<200>  & ~\encrypt<0> ;
  assign new_n1653_ = \key<192>  & \encrypt<0> ;
  assign new_n1654_ = ~new_n1652_ & ~new_n1653_;
  assign new_n1655_1_ = \start<0>  & ~new_n1654_;
  assign new_n1656_ = ~\C<90>  & ~\D<90> ;
  assign new_n1657_ = \C<90>  & \D<90> ;
  assign new_n1658_ = ~new_n1656_ & ~new_n1657_;
  assign new_n1659_ = ~new_n1185_1_ & ~new_n1658_;
  assign new_n1660_1_ = new_n1185_1_ & ~new_n1656_;
  assign new_n1661_ = ~new_n1659_ & ~new_n1660_1_;
  assign new_n1662_ = ~\encrypt<0>  & ~new_n1661_;
  assign new_n1663_ = \D<90>  & ~new_n1189_;
  assign new_n1664_ = ~\D<90>  & new_n1189_;
  assign new_n1665_1_ = ~new_n1663_ & ~new_n1664_;
  assign new_n1666_ = \C<90>  & ~new_n1665_1_;
  assign new_n1667_ = \D<90>  & new_n1189_;
  assign new_n1668_ = ~\C<90>  & new_n1667_;
  assign new_n1669_ = ~new_n1666_ & ~new_n1668_;
  assign new_n1670_1_ = \encrypt<0>  & ~new_n1669_;
  assign new_n1671_ = ~new_n1662_ & ~new_n1670_1_;
  assign new_n1672_ = ~\start<0>  & ~new_n1671_;
  assign n1025 = new_n1655_1_ | new_n1672_;
  assign new_n1674_ = \key<208>  & ~\encrypt<0> ;
  assign new_n1675_1_ = \key<200>  & \encrypt<0> ;
  assign new_n1676_ = ~new_n1674_ & ~new_n1675_1_;
  assign new_n1677_ = \start<0>  & ~new_n1676_;
  assign new_n1678_ = ~\C<89>  & ~\D<89> ;
  assign new_n1679_ = \C<89>  & \D<89> ;
  assign new_n1680_1_ = ~new_n1678_ & ~new_n1679_;
  assign new_n1681_ = ~new_n1185_1_ & ~new_n1680_1_;
  assign new_n1682_ = new_n1185_1_ & ~new_n1678_;
  assign new_n1683_ = ~new_n1681_ & ~new_n1682_;
  assign new_n1684_ = ~\encrypt<0>  & ~new_n1683_;
  assign new_n1685_1_ = \D<89>  & ~new_n1189_;
  assign new_n1686_ = ~\D<89>  & new_n1189_;
  assign new_n1687_ = ~new_n1685_1_ & ~new_n1686_;
  assign new_n1688_ = \C<89>  & ~new_n1687_;
  assign new_n1689_ = \D<89>  & new_n1189_;
  assign new_n1690_1_ = ~\C<89>  & new_n1689_;
  assign new_n1691_ = ~new_n1688_ & ~new_n1690_1_;
  assign new_n1692_ = \encrypt<0>  & ~new_n1691_;
  assign new_n1693_ = ~new_n1684_ & ~new_n1692_;
  assign new_n1694_ = ~\start<0>  & ~new_n1693_;
  assign n1030 = new_n1677_ | new_n1694_;
  assign new_n1696_ = \key<216>  & ~\encrypt<0> ;
  assign new_n1697_ = \key<208>  & \encrypt<0> ;
  assign new_n1698_ = ~new_n1696_ & ~new_n1697_;
  assign new_n1699_ = \start<0>  & ~new_n1698_;
  assign new_n1700_1_ = ~\C<88>  & ~\D<88> ;
  assign new_n1701_ = \C<88>  & \D<88> ;
  assign new_n1702_ = ~new_n1700_1_ & ~new_n1701_;
  assign new_n1703_ = ~new_n1185_1_ & ~new_n1702_;
  assign new_n1704_ = new_n1185_1_ & ~new_n1700_1_;
  assign new_n1705_1_ = ~new_n1703_ & ~new_n1704_;
  assign new_n1706_ = ~\encrypt<0>  & ~new_n1705_1_;
  assign new_n1707_ = \D<88>  & ~new_n1189_;
  assign new_n1708_ = ~\D<88>  & new_n1189_;
  assign new_n1709_ = ~new_n1707_ & ~new_n1708_;
  assign new_n1710_1_ = \C<88>  & ~new_n1709_;
  assign new_n1711_ = \D<88>  & new_n1189_;
  assign new_n1712_ = ~\C<88>  & new_n1711_;
  assign new_n1713_ = ~new_n1710_1_ & ~new_n1712_;
  assign new_n1714_ = \encrypt<0>  & ~new_n1713_;
  assign new_n1715_1_ = ~new_n1706_ & ~new_n1714_;
  assign new_n1716_ = ~\start<0>  & ~new_n1715_1_;
  assign n1035 = new_n1699_ | new_n1716_;
  assign new_n1718_ = \key<224>  & ~\encrypt<0> ;
  assign new_n1719_ = \key<216>  & \encrypt<0> ;
  assign new_n1720_1_ = ~new_n1718_ & ~new_n1719_;
  assign new_n1721_ = \start<0>  & ~new_n1720_1_;
  assign new_n1722_ = ~\C<87>  & ~\D<87> ;
  assign new_n1723_ = \C<87>  & \D<87> ;
  assign new_n1724_ = ~new_n1722_ & ~new_n1723_;
  assign new_n1725_1_ = ~new_n1185_1_ & ~new_n1724_;
  assign new_n1726_ = new_n1185_1_ & ~new_n1722_;
  assign new_n1727_ = ~new_n1725_1_ & ~new_n1726_;
  assign new_n1728_ = ~\encrypt<0>  & ~new_n1727_;
  assign new_n1729_ = \D<87>  & ~new_n1189_;
  assign new_n1730_1_ = ~\D<87>  & new_n1189_;
  assign new_n1731_ = ~new_n1729_ & ~new_n1730_1_;
  assign new_n1732_ = \C<87>  & ~new_n1731_;
  assign new_n1733_ = \D<87>  & new_n1189_;
  assign new_n1734_ = ~\C<87>  & new_n1733_;
  assign new_n1735_1_ = ~new_n1732_ & ~new_n1734_;
  assign new_n1736_ = \encrypt<0>  & ~new_n1735_1_;
  assign new_n1737_ = ~new_n1728_ & ~new_n1736_;
  assign new_n1738_ = ~\start<0>  & ~new_n1737_;
  assign n1040 = new_n1721_ | new_n1738_;
  assign new_n1740_1_ = \key<232>  & ~\encrypt<0> ;
  assign new_n1741_ = \key<224>  & \encrypt<0> ;
  assign new_n1742_ = ~new_n1740_1_ & ~new_n1741_;
  assign new_n1743_ = \start<0>  & ~new_n1742_;
  assign new_n1744_ = ~\C<86>  & ~\D<86> ;
  assign new_n1745_1_ = \C<86>  & \D<86> ;
  assign new_n1746_ = ~new_n1744_ & ~new_n1745_1_;
  assign new_n1747_ = ~new_n1185_1_ & ~new_n1746_;
  assign new_n1748_ = new_n1185_1_ & ~new_n1744_;
  assign new_n1749_ = ~new_n1747_ & ~new_n1748_;
  assign new_n1750_1_ = ~\encrypt<0>  & ~new_n1749_;
  assign new_n1751_ = \D<86>  & ~new_n1189_;
  assign new_n1752_ = ~\D<86>  & new_n1189_;
  assign new_n1753_ = ~new_n1751_ & ~new_n1752_;
  assign new_n1754_ = \C<86>  & ~new_n1753_;
  assign new_n1755_1_ = \D<86>  & new_n1189_;
  assign new_n1756_ = ~\C<86>  & new_n1755_1_;
  assign new_n1757_ = ~new_n1754_ & ~new_n1756_;
  assign new_n1758_ = \encrypt<0>  & ~new_n1757_;
  assign new_n1759_ = ~new_n1750_1_ & ~new_n1758_;
  assign new_n1760_1_ = ~\start<0>  & ~new_n1759_;
  assign n1045 = new_n1743_ | new_n1760_1_;
  assign new_n1762_ = \key<240>  & ~\encrypt<0> ;
  assign new_n1763_ = \key<232>  & \encrypt<0> ;
  assign new_n1764_ = ~new_n1762_ & ~new_n1763_;
  assign new_n1765_1_ = \start<0>  & ~new_n1764_;
  assign new_n1766_ = ~\C<85>  & ~\D<85> ;
  assign new_n1767_ = \C<85>  & \D<85> ;
  assign new_n1768_ = ~new_n1766_ & ~new_n1767_;
  assign new_n1769_ = ~new_n1185_1_ & ~new_n1768_;
  assign new_n1770_1_ = new_n1185_1_ & ~new_n1766_;
  assign new_n1771_ = ~new_n1769_ & ~new_n1770_1_;
  assign new_n1772_ = ~\encrypt<0>  & ~new_n1771_;
  assign new_n1773_ = \D<85>  & ~new_n1189_;
  assign new_n1774_ = ~\D<85>  & new_n1189_;
  assign new_n1775_1_ = ~new_n1773_ & ~new_n1774_;
  assign new_n1776_ = \C<85>  & ~new_n1775_1_;
  assign new_n1777_ = \D<85>  & new_n1189_;
  assign new_n1778_ = ~\C<85>  & new_n1777_;
  assign new_n1779_ = ~new_n1776_ & ~new_n1778_;
  assign new_n1780_1_ = \encrypt<0>  & ~new_n1779_;
  assign new_n1781_ = ~new_n1772_ & ~new_n1780_1_;
  assign new_n1782_ = ~\start<0>  & ~new_n1781_;
  assign n1050 = new_n1765_1_ | new_n1782_;
  assign new_n1784_ = \key<248>  & ~\encrypt<0> ;
  assign new_n1785_1_ = \key<240>  & \encrypt<0> ;
  assign new_n1786_ = ~new_n1784_ & ~new_n1785_1_;
  assign new_n1787_ = \start<0>  & ~new_n1786_;
  assign new_n1788_ = ~\C<84>  & ~\D<84> ;
  assign new_n1789_ = \C<84>  & \D<84> ;
  assign new_n1790_1_ = ~new_n1788_ & ~new_n1789_;
  assign new_n1791_ = ~new_n1185_1_ & ~new_n1790_1_;
  assign new_n1792_ = new_n1185_1_ & ~new_n1788_;
  assign new_n1793_ = ~new_n1791_ & ~new_n1792_;
  assign new_n1794_ = ~\encrypt<0>  & ~new_n1793_;
  assign new_n1795_1_ = \D<84>  & ~new_n1189_;
  assign new_n1796_ = ~\D<84>  & new_n1189_;
  assign new_n1797_ = ~new_n1795_1_ & ~new_n1796_;
  assign new_n1798_ = \C<84>  & ~new_n1797_;
  assign new_n1799_ = \D<84>  & new_n1189_;
  assign new_n1800_1_ = ~\C<84>  & new_n1799_;
  assign new_n1801_ = ~new_n1798_ & ~new_n1800_1_;
  assign new_n1802_ = \encrypt<0>  & ~new_n1801_;
  assign new_n1803_ = ~new_n1794_ & ~new_n1802_;
  assign new_n1804_ = ~\start<0>  & ~new_n1803_;
  assign n1055 = new_n1787_ | new_n1804_;
  assign new_n1806_ = \key<163>  & ~\encrypt<0> ;
  assign new_n1807_ = \key<248>  & \encrypt<0> ;
  assign new_n1808_ = ~new_n1806_ & ~new_n1807_;
  assign new_n1809_ = \start<0>  & ~new_n1808_;
  assign new_n1810_1_ = ~\C<83>  & ~\D<83> ;
  assign new_n1811_ = \C<83>  & \D<83> ;
  assign new_n1812_ = ~new_n1810_1_ & ~new_n1811_;
  assign new_n1813_ = ~new_n1185_1_ & ~new_n1812_;
  assign new_n1814_ = new_n1185_1_ & ~new_n1810_1_;
  assign new_n1815_1_ = ~new_n1813_ & ~new_n1814_;
  assign new_n1816_ = ~\encrypt<0>  & ~new_n1815_1_;
  assign new_n1817_ = \D<83>  & ~new_n1189_;
  assign new_n1818_ = ~\D<83>  & new_n1189_;
  assign new_n1819_ = ~new_n1817_ & ~new_n1818_;
  assign new_n1820_1_ = \C<83>  & ~new_n1819_;
  assign new_n1821_ = \D<83>  & new_n1189_;
  assign new_n1822_ = ~\C<83>  & new_n1821_;
  assign new_n1823_ = ~new_n1820_1_ & ~new_n1822_;
  assign new_n1824_ = \encrypt<0>  & ~new_n1823_;
  assign new_n1825_1_ = ~new_n1816_ & ~new_n1824_;
  assign new_n1826_ = ~\start<0>  & ~new_n1825_1_;
  assign n1060 = new_n1809_ | new_n1826_;
  assign new_n1828_ = \key<171>  & ~\encrypt<0> ;
  assign new_n1829_ = \key<163>  & \encrypt<0> ;
  assign new_n1830_1_ = ~new_n1828_ & ~new_n1829_;
  assign new_n1831_ = \start<0>  & ~new_n1830_1_;
  assign new_n1832_ = ~\C<82>  & ~\D<82> ;
  assign new_n1833_ = \C<82>  & \D<82> ;
  assign new_n1834_ = ~new_n1832_ & ~new_n1833_;
  assign new_n1835_1_ = ~new_n1185_1_ & ~new_n1834_;
  assign new_n1836_ = new_n1185_1_ & ~new_n1832_;
  assign new_n1837_ = ~new_n1835_1_ & ~new_n1836_;
  assign new_n1838_ = ~\encrypt<0>  & ~new_n1837_;
  assign new_n1839_ = \D<82>  & ~new_n1189_;
  assign new_n1840_1_ = ~\D<82>  & new_n1189_;
  assign new_n1841_ = ~new_n1839_ & ~new_n1840_1_;
  assign new_n1842_ = \C<82>  & ~new_n1841_;
  assign new_n1843_ = \D<82>  & new_n1189_;
  assign new_n1844_ = ~\C<82>  & new_n1843_;
  assign new_n1845_1_ = ~new_n1842_ & ~new_n1844_;
  assign new_n1846_ = \encrypt<0>  & ~new_n1845_1_;
  assign new_n1847_ = ~new_n1838_ & ~new_n1846_;
  assign new_n1848_ = ~\start<0>  & ~new_n1847_;
  assign n1065 = new_n1831_ | new_n1848_;
  assign new_n1850_1_ = \key<179>  & ~\encrypt<0> ;
  assign new_n1851_ = \key<171>  & \encrypt<0> ;
  assign new_n1852_ = ~new_n1850_1_ & ~new_n1851_;
  assign new_n1853_ = \start<0>  & ~new_n1852_;
  assign new_n1854_ = ~\C<81>  & ~\D<81> ;
  assign new_n1855_1_ = \C<81>  & \D<81> ;
  assign new_n1856_ = ~new_n1854_ & ~new_n1855_1_;
  assign new_n1857_ = ~new_n1185_1_ & ~new_n1856_;
  assign new_n1858_ = new_n1185_1_ & ~new_n1854_;
  assign new_n1859_ = ~new_n1857_ & ~new_n1858_;
  assign new_n1860_1_ = ~\encrypt<0>  & ~new_n1859_;
  assign new_n1861_ = \D<81>  & ~new_n1189_;
  assign new_n1862_ = ~\D<81>  & new_n1189_;
  assign new_n1863_ = ~new_n1861_ & ~new_n1862_;
  assign new_n1864_ = \C<81>  & ~new_n1863_;
  assign new_n1865_1_ = \D<81>  & new_n1189_;
  assign new_n1866_ = ~\C<81>  & new_n1865_1_;
  assign new_n1867_ = ~new_n1864_ & ~new_n1866_;
  assign new_n1868_ = \encrypt<0>  & ~new_n1867_;
  assign new_n1869_ = ~new_n1860_1_ & ~new_n1868_;
  assign new_n1870_1_ = ~\start<0>  & ~new_n1869_;
  assign n1070 = new_n1853_ | new_n1870_1_;
  assign new_n1872_ = \key<187>  & ~\encrypt<0> ;
  assign new_n1873_ = \key<179>  & \encrypt<0> ;
  assign new_n1874_ = ~new_n1872_ & ~new_n1873_;
  assign new_n1875_1_ = \start<0>  & ~new_n1874_;
  assign new_n1876_ = ~\C<80>  & ~\D<80> ;
  assign new_n1877_ = \C<80>  & \D<80> ;
  assign new_n1878_ = ~new_n1876_ & ~new_n1877_;
  assign new_n1879_ = ~new_n1185_1_ & ~new_n1878_;
  assign new_n1880_1_ = new_n1185_1_ & ~new_n1876_;
  assign new_n1881_ = ~new_n1879_ & ~new_n1880_1_;
  assign new_n1882_ = ~\encrypt<0>  & ~new_n1881_;
  assign new_n1883_ = \D<80>  & ~new_n1189_;
  assign new_n1884_ = ~\D<80>  & new_n1189_;
  assign new_n1885_1_ = ~new_n1883_ & ~new_n1884_;
  assign new_n1886_ = \C<80>  & ~new_n1885_1_;
  assign new_n1887_ = \D<80>  & new_n1189_;
  assign new_n1888_ = ~\C<80>  & new_n1887_;
  assign new_n1889_ = ~new_n1886_ & ~new_n1888_;
  assign new_n1890_1_ = \encrypt<0>  & ~new_n1889_;
  assign new_n1891_ = ~new_n1882_ & ~new_n1890_1_;
  assign new_n1892_ = ~\start<0>  & ~new_n1891_;
  assign n1075 = new_n1875_1_ | new_n1892_;
  assign new_n1894_ = \key<130>  & ~\encrypt<0> ;
  assign new_n1895_1_ = \key<187>  & \encrypt<0> ;
  assign new_n1896_ = ~new_n1894_ & ~new_n1895_1_;
  assign new_n1897_ = \start<0>  & ~new_n1896_;
  assign new_n1898_ = ~\C<79>  & ~\D<79> ;
  assign new_n1899_ = \C<79>  & \D<79> ;
  assign new_n1900_1_ = ~new_n1898_ & ~new_n1899_;
  assign new_n1901_ = ~new_n1185_1_ & ~new_n1900_1_;
  assign new_n1902_ = new_n1185_1_ & ~new_n1898_;
  assign new_n1903_ = ~new_n1901_ & ~new_n1902_;
  assign new_n1904_ = ~\encrypt<0>  & ~new_n1903_;
  assign new_n1905_1_ = \D<79>  & ~new_n1189_;
  assign new_n1906_ = ~\D<79>  & new_n1189_;
  assign new_n1907_ = ~new_n1905_1_ & ~new_n1906_;
  assign new_n1908_ = \C<79>  & ~new_n1907_;
  assign new_n1909_ = \D<79>  & new_n1189_;
  assign new_n1910_1_ = ~\C<79>  & new_n1909_;
  assign new_n1911_ = ~new_n1908_ & ~new_n1910_1_;
  assign new_n1912_ = \encrypt<0>  & ~new_n1911_;
  assign new_n1913_ = ~new_n1904_ & ~new_n1912_;
  assign new_n1914_ = ~\start<0>  & ~new_n1913_;
  assign n1080 = new_n1897_ | new_n1914_;
  assign new_n1916_ = \key<138>  & ~\encrypt<0> ;
  assign new_n1917_ = \key<130>  & \encrypt<0> ;
  assign new_n1918_ = ~new_n1916_ & ~new_n1917_;
  assign new_n1919_ = \start<0>  & ~new_n1918_;
  assign new_n1920_1_ = ~\C<78>  & ~\D<78> ;
  assign new_n1921_ = \C<78>  & \D<78> ;
  assign new_n1922_ = ~new_n1920_1_ & ~new_n1921_;
  assign new_n1923_ = ~new_n1185_1_ & ~new_n1922_;
  assign new_n1924_ = new_n1185_1_ & ~new_n1920_1_;
  assign new_n1925_1_ = ~new_n1923_ & ~new_n1924_;
  assign new_n1926_ = ~\encrypt<0>  & ~new_n1925_1_;
  assign new_n1927_ = \D<78>  & ~new_n1189_;
  assign new_n1928_ = ~\D<78>  & new_n1189_;
  assign new_n1929_ = ~new_n1927_ & ~new_n1928_;
  assign new_n1930_1_ = \C<78>  & ~new_n1929_;
  assign new_n1931_ = \D<78>  & new_n1189_;
  assign new_n1932_ = ~\C<78>  & new_n1931_;
  assign new_n1933_ = ~new_n1930_1_ & ~new_n1932_;
  assign new_n1934_ = \encrypt<0>  & ~new_n1933_;
  assign new_n1935_1_ = ~new_n1926_ & ~new_n1934_;
  assign new_n1936_ = ~\start<0>  & ~new_n1935_1_;
  assign n1085 = new_n1919_ | new_n1936_;
  assign new_n1938_ = \key<146>  & ~\encrypt<0> ;
  assign new_n1939_ = \key<138>  & \encrypt<0> ;
  assign new_n1940_1_ = ~new_n1938_ & ~new_n1939_;
  assign new_n1941_ = \start<0>  & ~new_n1940_1_;
  assign new_n1942_ = ~\C<77>  & ~\D<77> ;
  assign new_n1943_ = \C<77>  & \D<77> ;
  assign new_n1944_ = ~new_n1942_ & ~new_n1943_;
  assign new_n1945_1_ = ~new_n1185_1_ & ~new_n1944_;
  assign new_n1946_ = new_n1185_1_ & ~new_n1942_;
  assign new_n1947_ = ~new_n1945_1_ & ~new_n1946_;
  assign new_n1948_ = ~\encrypt<0>  & ~new_n1947_;
  assign new_n1949_ = \D<77>  & ~new_n1189_;
  assign new_n1950_1_ = ~\D<77>  & new_n1189_;
  assign new_n1951_ = ~new_n1949_ & ~new_n1950_1_;
  assign new_n1952_ = \C<77>  & ~new_n1951_;
  assign new_n1953_ = \D<77>  & new_n1189_;
  assign new_n1954_ = ~\C<77>  & new_n1953_;
  assign new_n1955_1_ = ~new_n1952_ & ~new_n1954_;
  assign new_n1956_ = \encrypt<0>  & ~new_n1955_1_;
  assign new_n1957_ = ~new_n1948_ & ~new_n1956_;
  assign new_n1958_ = ~\start<0>  & ~new_n1957_;
  assign n1090 = new_n1941_ | new_n1958_;
  assign new_n1960_1_ = \key<154>  & ~\encrypt<0> ;
  assign new_n1961_ = \key<146>  & \encrypt<0> ;
  assign new_n1962_ = ~new_n1960_1_ & ~new_n1961_;
  assign new_n1963_ = \start<0>  & ~new_n1962_;
  assign new_n1964_ = ~\C<76>  & ~\D<76> ;
  assign new_n1965_1_ = \C<76>  & \D<76> ;
  assign new_n1966_ = ~new_n1964_ & ~new_n1965_1_;
  assign new_n1967_ = ~new_n1185_1_ & ~new_n1966_;
  assign new_n1968_ = new_n1185_1_ & ~new_n1964_;
  assign new_n1969_ = ~new_n1967_ & ~new_n1968_;
  assign new_n1970_1_ = ~\encrypt<0>  & ~new_n1969_;
  assign new_n1971_ = \D<76>  & ~new_n1189_;
  assign new_n1972_ = ~\D<76>  & new_n1189_;
  assign new_n1973_ = ~new_n1971_ & ~new_n1972_;
  assign new_n1974_ = \C<76>  & ~new_n1973_;
  assign new_n1975_1_ = \D<76>  & new_n1189_;
  assign new_n1976_ = ~\C<76>  & new_n1975_1_;
  assign new_n1977_ = ~new_n1974_ & ~new_n1976_;
  assign new_n1978_ = \encrypt<0>  & ~new_n1977_;
  assign new_n1979_ = ~new_n1970_1_ & ~new_n1978_;
  assign new_n1980_1_ = ~\start<0>  & ~new_n1979_;
  assign n1095 = new_n1963_ | new_n1980_1_;
  assign new_n1982_ = \key<162>  & ~\encrypt<0> ;
  assign new_n1983_ = \key<154>  & \encrypt<0> ;
  assign new_n1984_ = ~new_n1982_ & ~new_n1983_;
  assign new_n1985_1_ = \start<0>  & ~new_n1984_;
  assign new_n1986_ = ~\C<75>  & ~\D<75> ;
  assign new_n1987_ = \C<75>  & \D<75> ;
  assign new_n1988_ = ~new_n1986_ & ~new_n1987_;
  assign new_n1989_ = ~new_n1185_1_ & ~new_n1988_;
  assign new_n1990_1_ = new_n1185_1_ & ~new_n1986_;
  assign new_n1991_ = ~new_n1989_ & ~new_n1990_1_;
  assign new_n1992_ = ~\encrypt<0>  & ~new_n1991_;
  assign new_n1993_ = \D<75>  & ~new_n1189_;
  assign new_n1994_ = ~\D<75>  & new_n1189_;
  assign new_n1995_1_ = ~new_n1993_ & ~new_n1994_;
  assign new_n1996_ = \C<75>  & ~new_n1995_1_;
  assign new_n1997_ = \D<75>  & new_n1189_;
  assign new_n1998_ = ~\C<75>  & new_n1997_;
  assign new_n1999_ = ~new_n1996_ & ~new_n1998_;
  assign new_n2000_1_ = \encrypt<0>  & ~new_n1999_;
  assign new_n2001_ = ~new_n1992_ & ~new_n2000_1_;
  assign new_n2002_ = ~\start<0>  & ~new_n2001_;
  assign n1100 = new_n1985_1_ | new_n2002_;
  assign new_n2004_ = \key<170>  & ~\encrypt<0> ;
  assign new_n2005_1_ = \key<162>  & \encrypt<0> ;
  assign new_n2006_ = ~new_n2004_ & ~new_n2005_1_;
  assign new_n2007_ = \start<0>  & ~new_n2006_;
  assign new_n2008_ = ~\C<74>  & ~\D<74> ;
  assign new_n2009_ = \C<74>  & \D<74> ;
  assign new_n2010_1_ = ~new_n2008_ & ~new_n2009_;
  assign new_n2011_ = ~new_n1185_1_ & ~new_n2010_1_;
  assign new_n2012_ = new_n1185_1_ & ~new_n2008_;
  assign new_n2013_ = ~new_n2011_ & ~new_n2012_;
  assign new_n2014_ = ~\encrypt<0>  & ~new_n2013_;
  assign new_n2015_1_ = \D<74>  & ~new_n1189_;
  assign new_n2016_ = ~\D<74>  & new_n1189_;
  assign new_n2017_ = ~new_n2015_1_ & ~new_n2016_;
  assign new_n2018_ = \C<74>  & ~new_n2017_;
  assign new_n2019_ = \D<74>  & new_n1189_;
  assign new_n2020_1_ = ~\C<74>  & new_n2019_;
  assign new_n2021_ = ~new_n2018_ & ~new_n2020_1_;
  assign new_n2022_ = \encrypt<0>  & ~new_n2021_;
  assign new_n2023_ = ~new_n2014_ & ~new_n2022_;
  assign new_n2024_ = ~\start<0>  & ~new_n2023_;
  assign n1105 = new_n2007_ | new_n2024_;
  assign new_n2026_ = \key<178>  & ~\encrypt<0> ;
  assign new_n2027_ = \key<170>  & \encrypt<0> ;
  assign new_n2028_ = ~new_n2026_ & ~new_n2027_;
  assign new_n2029_ = \start<0>  & ~new_n2028_;
  assign new_n2030_1_ = ~\C<73>  & ~\D<73> ;
  assign new_n2031_ = \C<73>  & \D<73> ;
  assign new_n2032_ = ~new_n2030_1_ & ~new_n2031_;
  assign new_n2033_ = ~new_n1185_1_ & ~new_n2032_;
  assign new_n2034_ = new_n1185_1_ & ~new_n2030_1_;
  assign new_n2035_1_ = ~new_n2033_ & ~new_n2034_;
  assign new_n2036_ = ~\encrypt<0>  & ~new_n2035_1_;
  assign new_n2037_ = \D<73>  & ~new_n1189_;
  assign new_n2038_ = ~\D<73>  & new_n1189_;
  assign new_n2039_ = ~new_n2037_ & ~new_n2038_;
  assign new_n2040_ = \C<73>  & ~new_n2039_;
  assign new_n2041_ = \D<73>  & new_n1189_;
  assign new_n2042_ = ~\C<73>  & new_n2041_;
  assign new_n2043_ = ~new_n2040_ & ~new_n2042_;
  assign new_n2044_ = \encrypt<0>  & ~new_n2043_;
  assign new_n2045_ = ~new_n2036_ & ~new_n2044_;
  assign new_n2046_ = ~\start<0>  & ~new_n2045_;
  assign n1110 = new_n2029_ | new_n2046_;
  assign new_n2048_ = \key<186>  & ~\encrypt<0> ;
  assign new_n2049_ = \key<178>  & \encrypt<0> ;
  assign new_n2050_ = ~new_n2048_ & ~new_n2049_;
  assign new_n2051_ = \start<0>  & ~new_n2050_;
  assign new_n2052_ = ~\C<72>  & ~\D<72> ;
  assign new_n2053_ = \C<72>  & \D<72> ;
  assign new_n2054_ = ~new_n2052_ & ~new_n2053_;
  assign new_n2055_ = ~new_n1185_1_ & ~new_n2054_;
  assign new_n2056_ = new_n1185_1_ & ~new_n2052_;
  assign new_n2057_ = ~new_n2055_ & ~new_n2056_;
  assign new_n2058_ = ~\encrypt<0>  & ~new_n2057_;
  assign new_n2059_ = \D<72>  & ~new_n1189_;
  assign new_n2060_ = ~\D<72>  & new_n1189_;
  assign new_n2061_ = ~new_n2059_ & ~new_n2060_;
  assign new_n2062_ = \C<72>  & ~new_n2061_;
  assign new_n2063_ = \D<72>  & new_n1189_;
  assign new_n2064_ = ~\C<72>  & new_n2063_;
  assign new_n2065_ = ~new_n2062_ & ~new_n2064_;
  assign new_n2066_ = \encrypt<0>  & ~new_n2065_;
  assign new_n2067_ = ~new_n2058_ & ~new_n2066_;
  assign new_n2068_ = ~\start<0>  & ~new_n2067_;
  assign n1115 = new_n2051_ | new_n2068_;
  assign new_n2070_ = \key<129>  & ~\encrypt<0> ;
  assign new_n2071_ = \key<186>  & \encrypt<0> ;
  assign new_n2072_ = ~new_n2070_ & ~new_n2071_;
  assign new_n2073_ = \start<0>  & ~new_n2072_;
  assign new_n2074_ = ~\C<71>  & ~\D<71> ;
  assign new_n2075_ = \C<71>  & \D<71> ;
  assign new_n2076_ = ~new_n2074_ & ~new_n2075_;
  assign new_n2077_ = ~new_n1185_1_ & ~new_n2076_;
  assign new_n2078_ = new_n1185_1_ & ~new_n2074_;
  assign new_n2079_ = ~new_n2077_ & ~new_n2078_;
  assign new_n2080_ = ~\encrypt<0>  & ~new_n2079_;
  assign new_n2081_ = \D<71>  & ~new_n1189_;
  assign new_n2082_ = ~\D<71>  & new_n1189_;
  assign new_n2083_ = ~new_n2081_ & ~new_n2082_;
  assign new_n2084_ = \C<71>  & ~new_n2083_;
  assign new_n2085_ = \D<71>  & new_n1189_;
  assign new_n2086_ = ~\C<71>  & new_n2085_;
  assign new_n2087_ = ~new_n2084_ & ~new_n2086_;
  assign new_n2088_ = \encrypt<0>  & ~new_n2087_;
  assign new_n2089_ = ~new_n2080_ & ~new_n2088_;
  assign new_n2090_ = ~\start<0>  & ~new_n2089_;
  assign n1120 = new_n2073_ | new_n2090_;
  assign new_n2092_ = \key<137>  & ~\encrypt<0> ;
  assign new_n2093_ = \key<129>  & \encrypt<0> ;
  assign new_n2094_ = ~new_n2092_ & ~new_n2093_;
  assign new_n2095_ = \start<0>  & ~new_n2094_;
  assign new_n2096_ = ~\C<70>  & ~\D<70> ;
  assign new_n2097_ = \C<70>  & \D<70> ;
  assign new_n2098_ = ~new_n2096_ & ~new_n2097_;
  assign new_n2099_ = ~new_n1185_1_ & ~new_n2098_;
  assign new_n2100_ = new_n1185_1_ & ~new_n2096_;
  assign new_n2101_ = ~new_n2099_ & ~new_n2100_;
  assign new_n2102_ = ~\encrypt<0>  & ~new_n2101_;
  assign new_n2103_ = \D<70>  & ~new_n1189_;
  assign new_n2104_ = ~\D<70>  & new_n1189_;
  assign new_n2105_ = ~new_n2103_ & ~new_n2104_;
  assign new_n2106_ = \C<70>  & ~new_n2105_;
  assign new_n2107_ = \D<70>  & new_n1189_;
  assign new_n2108_ = ~\C<70>  & new_n2107_;
  assign new_n2109_ = ~new_n2106_ & ~new_n2108_;
  assign new_n2110_ = \encrypt<0>  & ~new_n2109_;
  assign new_n2111_ = ~new_n2102_ & ~new_n2110_;
  assign new_n2112_ = ~\start<0>  & ~new_n2111_;
  assign n1125 = new_n2095_ | new_n2112_;
  assign new_n2114_ = \key<145>  & ~\encrypt<0> ;
  assign new_n2115_ = \key<137>  & \encrypt<0> ;
  assign new_n2116_ = ~new_n2114_ & ~new_n2115_;
  assign new_n2117_ = \start<0>  & ~new_n2116_;
  assign new_n2118_ = ~\C<69>  & ~\D<69> ;
  assign new_n2119_ = \C<69>  & \D<69> ;
  assign new_n2120_ = ~new_n2118_ & ~new_n2119_;
  assign new_n2121_ = ~new_n1185_1_ & ~new_n2120_;
  assign new_n2122_ = new_n1185_1_ & ~new_n2118_;
  assign new_n2123_ = ~new_n2121_ & ~new_n2122_;
  assign new_n2124_ = ~\encrypt<0>  & ~new_n2123_;
  assign new_n2125_ = \D<69>  & ~new_n1189_;
  assign new_n2126_ = ~\D<69>  & new_n1189_;
  assign new_n2127_ = ~new_n2125_ & ~new_n2126_;
  assign new_n2128_ = \C<69>  & ~new_n2127_;
  assign new_n2129_ = \D<69>  & new_n1189_;
  assign new_n2130_ = ~\C<69>  & new_n2129_;
  assign new_n2131_ = ~new_n2128_ & ~new_n2130_;
  assign new_n2132_ = \encrypt<0>  & ~new_n2131_;
  assign new_n2133_ = ~new_n2124_ & ~new_n2132_;
  assign new_n2134_ = ~\start<0>  & ~new_n2133_;
  assign n1130 = new_n2117_ | new_n2134_;
  assign new_n2136_ = \key<153>  & ~\encrypt<0> ;
  assign new_n2137_ = \key<145>  & \encrypt<0> ;
  assign new_n2138_ = ~new_n2136_ & ~new_n2137_;
  assign new_n2139_ = \start<0>  & ~new_n2138_;
  assign new_n2140_ = ~\C<68>  & ~\D<68> ;
  assign new_n2141_ = \C<68>  & \D<68> ;
  assign new_n2142_ = ~new_n2140_ & ~new_n2141_;
  assign new_n2143_ = ~new_n1185_1_ & ~new_n2142_;
  assign new_n2144_ = new_n1185_1_ & ~new_n2140_;
  assign new_n2145_ = ~new_n2143_ & ~new_n2144_;
  assign new_n2146_ = ~\encrypt<0>  & ~new_n2145_;
  assign new_n2147_ = \D<68>  & ~new_n1189_;
  assign new_n2148_ = ~\D<68>  & new_n1189_;
  assign new_n2149_ = ~new_n2147_ & ~new_n2148_;
  assign new_n2150_ = \C<68>  & ~new_n2149_;
  assign new_n2151_ = \D<68>  & new_n1189_;
  assign new_n2152_ = ~\C<68>  & new_n2151_;
  assign new_n2153_ = ~new_n2150_ & ~new_n2152_;
  assign new_n2154_ = \encrypt<0>  & ~new_n2153_;
  assign new_n2155_ = ~new_n2146_ & ~new_n2154_;
  assign new_n2156_ = ~\start<0>  & ~new_n2155_;
  assign n1135 = new_n2139_ | new_n2156_;
  assign new_n2158_ = \key<161>  & ~\encrypt<0> ;
  assign new_n2159_ = \key<153>  & \encrypt<0> ;
  assign new_n2160_ = ~new_n2158_ & ~new_n2159_;
  assign new_n2161_ = \start<0>  & ~new_n2160_;
  assign new_n2162_ = ~\C<67>  & ~\D<67> ;
  assign new_n2163_ = \C<67>  & \D<67> ;
  assign new_n2164_ = ~new_n2162_ & ~new_n2163_;
  assign new_n2165_ = ~new_n1185_1_ & ~new_n2164_;
  assign new_n2166_ = new_n1185_1_ & ~new_n2162_;
  assign new_n2167_ = ~new_n2165_ & ~new_n2166_;
  assign new_n2168_ = ~\encrypt<0>  & ~new_n2167_;
  assign new_n2169_ = \D<67>  & ~new_n1189_;
  assign new_n2170_ = ~\D<67>  & new_n1189_;
  assign new_n2171_ = ~new_n2169_ & ~new_n2170_;
  assign new_n2172_ = \C<67>  & ~new_n2171_;
  assign new_n2173_ = \D<67>  & new_n1189_;
  assign new_n2174_ = ~\C<67>  & new_n2173_;
  assign new_n2175_ = ~new_n2172_ & ~new_n2174_;
  assign new_n2176_ = \encrypt<0>  & ~new_n2175_;
  assign new_n2177_ = ~new_n2168_ & ~new_n2176_;
  assign new_n2178_ = ~\start<0>  & ~new_n2177_;
  assign n1140 = new_n2161_ | new_n2178_;
  assign new_n2180_ = \key<169>  & ~\encrypt<0> ;
  assign new_n2181_ = \key<161>  & \encrypt<0> ;
  assign new_n2182_ = ~new_n2180_ & ~new_n2181_;
  assign new_n2183_ = \start<0>  & ~new_n2182_;
  assign new_n2184_ = ~\C<66>  & ~\D<66> ;
  assign new_n2185_ = \C<66>  & \D<66> ;
  assign new_n2186_ = ~new_n2184_ & ~new_n2185_;
  assign new_n2187_ = ~new_n1185_1_ & ~new_n2186_;
  assign new_n2188_ = new_n1185_1_ & ~new_n2184_;
  assign new_n2189_ = ~new_n2187_ & ~new_n2188_;
  assign new_n2190_ = ~\encrypt<0>  & ~new_n2189_;
  assign new_n2191_ = \D<66>  & ~new_n1189_;
  assign new_n2192_ = ~\D<66>  & new_n1189_;
  assign new_n2193_ = ~new_n2191_ & ~new_n2192_;
  assign new_n2194_ = \C<66>  & ~new_n2193_;
  assign new_n2195_ = \D<66>  & new_n1189_;
  assign new_n2196_ = ~\C<66>  & new_n2195_;
  assign new_n2197_ = ~new_n2194_ & ~new_n2196_;
  assign new_n2198_ = \encrypt<0>  & ~new_n2197_;
  assign new_n2199_ = ~new_n2190_ & ~new_n2198_;
  assign new_n2200_ = ~\start<0>  & ~new_n2199_;
  assign n1145 = new_n2183_ | new_n2200_;
  assign new_n2202_ = \key<177>  & ~\encrypt<0> ;
  assign new_n2203_ = \key<169>  & \encrypt<0> ;
  assign new_n2204_ = ~new_n2202_ & ~new_n2203_;
  assign new_n2205_ = \start<0>  & ~new_n2204_;
  assign new_n2206_ = ~\C<65>  & ~\D<65> ;
  assign new_n2207_ = \C<65>  & \D<65> ;
  assign new_n2208_ = ~new_n2206_ & ~new_n2207_;
  assign new_n2209_ = ~new_n1185_1_ & ~new_n2208_;
  assign new_n2210_ = new_n1185_1_ & ~new_n2206_;
  assign new_n2211_ = ~new_n2209_ & ~new_n2210_;
  assign new_n2212_ = ~\encrypt<0>  & ~new_n2211_;
  assign new_n2213_ = \D<65>  & ~new_n1189_;
  assign new_n2214_ = ~\D<65>  & new_n1189_;
  assign new_n2215_ = ~new_n2213_ & ~new_n2214_;
  assign new_n2216_ = \C<65>  & ~new_n2215_;
  assign new_n2217_ = \D<65>  & new_n1189_;
  assign new_n2218_ = ~\C<65>  & new_n2217_;
  assign new_n2219_ = ~new_n2216_ & ~new_n2218_;
  assign new_n2220_ = \encrypt<0>  & ~new_n2219_;
  assign new_n2221_ = ~new_n2212_ & ~new_n2220_;
  assign new_n2222_ = ~\start<0>  & ~new_n2221_;
  assign n1150 = new_n2205_ | new_n2222_;
  assign new_n2224_ = \key<185>  & ~\encrypt<0> ;
  assign new_n2225_ = \key<177>  & \encrypt<0> ;
  assign new_n2226_ = ~new_n2224_ & ~new_n2225_;
  assign new_n2227_ = \start<0>  & ~new_n2226_;
  assign new_n2228_ = ~\C<64>  & ~\D<64> ;
  assign new_n2229_ = \C<64>  & \D<64> ;
  assign new_n2230_ = ~new_n2228_ & ~new_n2229_;
  assign new_n2231_ = ~new_n1185_1_ & ~new_n2230_;
  assign new_n2232_ = new_n1185_1_ & ~new_n2228_;
  assign new_n2233_ = ~new_n2231_ & ~new_n2232_;
  assign new_n2234_ = ~\encrypt<0>  & ~new_n2233_;
  assign new_n2235_ = \D<64>  & ~new_n1189_;
  assign new_n2236_ = ~\D<64>  & new_n1189_;
  assign new_n2237_ = ~new_n2235_ & ~new_n2236_;
  assign new_n2238_ = \C<64>  & ~new_n2237_;
  assign new_n2239_ = \D<64>  & new_n1189_;
  assign new_n2240_ = ~\C<64>  & new_n2239_;
  assign new_n2241_ = ~new_n2238_ & ~new_n2240_;
  assign new_n2242_ = \encrypt<0>  & ~new_n2241_;
  assign new_n2243_ = ~new_n2234_ & ~new_n2242_;
  assign new_n2244_ = ~\start<0>  & ~new_n2243_;
  assign n1155 = new_n2227_ | new_n2244_;
  assign new_n2246_ = \key<128>  & ~\encrypt<0> ;
  assign new_n2247_ = \key<185>  & \encrypt<0> ;
  assign new_n2248_ = ~new_n2246_ & ~new_n2247_;
  assign new_n2249_ = \start<0>  & ~new_n2248_;
  assign new_n2250_ = ~\C<63>  & ~\D<63> ;
  assign new_n2251_ = \C<63>  & \D<63> ;
  assign new_n2252_ = ~new_n2250_ & ~new_n2251_;
  assign new_n2253_ = ~new_n1185_1_ & ~new_n2252_;
  assign new_n2254_ = new_n1185_1_ & ~new_n2250_;
  assign new_n2255_ = ~new_n2253_ & ~new_n2254_;
  assign new_n2256_ = ~\encrypt<0>  & ~new_n2255_;
  assign new_n2257_ = \D<63>  & ~new_n1189_;
  assign new_n2258_ = ~\D<63>  & new_n1189_;
  assign new_n2259_ = ~new_n2257_ & ~new_n2258_;
  assign new_n2260_ = \C<63>  & ~new_n2259_;
  assign new_n2261_ = \D<63>  & new_n1189_;
  assign new_n2262_ = ~\C<63>  & new_n2261_;
  assign new_n2263_ = ~new_n2260_ & ~new_n2262_;
  assign new_n2264_ = \encrypt<0>  & ~new_n2263_;
  assign new_n2265_ = ~new_n2256_ & ~new_n2264_;
  assign new_n2266_ = ~\start<0>  & ~new_n2265_;
  assign n1160 = new_n2249_ | new_n2266_;
  assign new_n2268_ = \key<136>  & ~\encrypt<0> ;
  assign new_n2269_ = \key<128>  & \encrypt<0> ;
  assign new_n2270_ = ~new_n2268_ & ~new_n2269_;
  assign new_n2271_ = \start<0>  & ~new_n2270_;
  assign new_n2272_ = ~\C<62>  & ~\D<62> ;
  assign new_n2273_ = \C<62>  & \D<62> ;
  assign new_n2274_ = ~new_n2272_ & ~new_n2273_;
  assign new_n2275_ = ~new_n1185_1_ & ~new_n2274_;
  assign new_n2276_ = new_n1185_1_ & ~new_n2272_;
  assign new_n2277_ = ~new_n2275_ & ~new_n2276_;
  assign new_n2278_ = ~\encrypt<0>  & ~new_n2277_;
  assign new_n2279_ = \D<62>  & ~new_n1189_;
  assign new_n2280_ = ~\D<62>  & new_n1189_;
  assign new_n2281_ = ~new_n2279_ & ~new_n2280_;
  assign new_n2282_ = \C<62>  & ~new_n2281_;
  assign new_n2283_ = \D<62>  & new_n1189_;
  assign new_n2284_ = ~\C<62>  & new_n2283_;
  assign new_n2285_ = ~new_n2282_ & ~new_n2284_;
  assign new_n2286_ = \encrypt<0>  & ~new_n2285_;
  assign new_n2287_ = ~new_n2278_ & ~new_n2286_;
  assign new_n2288_ = ~\start<0>  & ~new_n2287_;
  assign n1165 = new_n2271_ | new_n2288_;
  assign new_n2290_ = \key<144>  & ~\encrypt<0> ;
  assign new_n2291_ = \key<136>  & \encrypt<0> ;
  assign new_n2292_ = ~new_n2290_ & ~new_n2291_;
  assign new_n2293_ = \start<0>  & ~new_n2292_;
  assign new_n2294_ = ~\C<61>  & ~\D<61> ;
  assign new_n2295_ = \C<61>  & \D<61> ;
  assign new_n2296_ = ~new_n2294_ & ~new_n2295_;
  assign new_n2297_ = ~new_n1185_1_ & ~new_n2296_;
  assign new_n2298_ = new_n1185_1_ & ~new_n2294_;
  assign new_n2299_ = ~new_n2297_ & ~new_n2298_;
  assign new_n2300_ = ~\encrypt<0>  & ~new_n2299_;
  assign new_n2301_ = \D<61>  & ~new_n1189_;
  assign new_n2302_ = ~\D<61>  & new_n1189_;
  assign new_n2303_ = ~new_n2301_ & ~new_n2302_;
  assign new_n2304_ = \C<61>  & ~new_n2303_;
  assign new_n2305_ = \D<61>  & new_n1189_;
  assign new_n2306_ = ~\C<61>  & new_n2305_;
  assign new_n2307_ = ~new_n2304_ & ~new_n2306_;
  assign new_n2308_ = \encrypt<0>  & ~new_n2307_;
  assign new_n2309_ = ~new_n2300_ & ~new_n2308_;
  assign new_n2310_ = ~\start<0>  & ~new_n2309_;
  assign n1170 = new_n2293_ | new_n2310_;
  assign new_n2312_ = \key<152>  & ~\encrypt<0> ;
  assign new_n2313_ = \key<144>  & \encrypt<0> ;
  assign new_n2314_ = ~new_n2312_ & ~new_n2313_;
  assign new_n2315_ = \start<0>  & ~new_n2314_;
  assign new_n2316_ = ~\C<60>  & ~\D<60> ;
  assign new_n2317_ = \C<60>  & \D<60> ;
  assign new_n2318_ = ~new_n2316_ & ~new_n2317_;
  assign new_n2319_ = ~new_n1185_1_ & ~new_n2318_;
  assign new_n2320_ = new_n1185_1_ & ~new_n2316_;
  assign new_n2321_ = ~new_n2319_ & ~new_n2320_;
  assign new_n2322_ = ~\encrypt<0>  & ~new_n2321_;
  assign new_n2323_ = \D<60>  & ~new_n1189_;
  assign new_n2324_ = ~\D<60>  & new_n1189_;
  assign new_n2325_ = ~new_n2323_ & ~new_n2324_;
  assign new_n2326_ = \C<60>  & ~new_n2325_;
  assign new_n2327_ = \D<60>  & new_n1189_;
  assign new_n2328_ = ~\C<60>  & new_n2327_;
  assign new_n2329_ = ~new_n2326_ & ~new_n2328_;
  assign new_n2330_ = \encrypt<0>  & ~new_n2329_;
  assign new_n2331_ = ~new_n2322_ & ~new_n2330_;
  assign new_n2332_ = ~\start<0>  & ~new_n2331_;
  assign n1175 = new_n2315_ | new_n2332_;
  assign new_n2334_ = \key<160>  & ~\encrypt<0> ;
  assign new_n2335_ = \key<152>  & \encrypt<0> ;
  assign new_n2336_ = ~new_n2334_ & ~new_n2335_;
  assign new_n2337_ = \start<0>  & ~new_n2336_;
  assign new_n2338_ = ~\C<59>  & ~\D<59> ;
  assign new_n2339_ = \C<59>  & \D<59> ;
  assign new_n2340_ = ~new_n2338_ & ~new_n2339_;
  assign new_n2341_ = ~new_n1185_1_ & ~new_n2340_;
  assign new_n2342_ = new_n1185_1_ & ~new_n2338_;
  assign new_n2343_ = ~new_n2341_ & ~new_n2342_;
  assign new_n2344_ = ~\encrypt<0>  & ~new_n2343_;
  assign new_n2345_ = \D<59>  & ~new_n1189_;
  assign new_n2346_ = ~\D<59>  & new_n1189_;
  assign new_n2347_ = ~new_n2345_ & ~new_n2346_;
  assign new_n2348_ = \C<59>  & ~new_n2347_;
  assign new_n2349_ = \D<59>  & new_n1189_;
  assign new_n2350_ = ~\C<59>  & new_n2349_;
  assign new_n2351_ = ~new_n2348_ & ~new_n2350_;
  assign new_n2352_ = \encrypt<0>  & ~new_n2351_;
  assign new_n2353_ = ~new_n2344_ & ~new_n2352_;
  assign new_n2354_ = ~\start<0>  & ~new_n2353_;
  assign n1180 = new_n2337_ | new_n2354_;
  assign new_n2356_ = \key<168>  & ~\encrypt<0> ;
  assign new_n2357_ = \key<160>  & \encrypt<0> ;
  assign new_n2358_ = ~new_n2356_ & ~new_n2357_;
  assign new_n2359_ = \start<0>  & ~new_n2358_;
  assign new_n2360_ = ~\C<58>  & ~\D<58> ;
  assign new_n2361_ = \C<58>  & \D<58> ;
  assign new_n2362_ = ~new_n2360_ & ~new_n2361_;
  assign new_n2363_ = ~new_n1185_1_ & ~new_n2362_;
  assign new_n2364_ = new_n1185_1_ & ~new_n2360_;
  assign new_n2365_ = ~new_n2363_ & ~new_n2364_;
  assign new_n2366_ = ~\encrypt<0>  & ~new_n2365_;
  assign new_n2367_ = \D<58>  & ~new_n1189_;
  assign new_n2368_ = ~\D<58>  & new_n1189_;
  assign new_n2369_ = ~new_n2367_ & ~new_n2368_;
  assign new_n2370_ = \C<58>  & ~new_n2369_;
  assign new_n2371_ = \D<58>  & new_n1189_;
  assign new_n2372_ = ~\C<58>  & new_n2371_;
  assign new_n2373_ = ~new_n2370_ & ~new_n2372_;
  assign new_n2374_ = \encrypt<0>  & ~new_n2373_;
  assign new_n2375_ = ~new_n2366_ & ~new_n2374_;
  assign new_n2376_ = ~\start<0>  & ~new_n2375_;
  assign n1185 = new_n2359_ | new_n2376_;
  assign new_n2378_ = \key<176>  & ~\encrypt<0> ;
  assign new_n2379_ = \key<168>  & \encrypt<0> ;
  assign new_n2380_ = ~new_n2378_ & ~new_n2379_;
  assign new_n2381_ = \start<0>  & ~new_n2380_;
  assign new_n2382_ = ~\C<57>  & ~\D<57> ;
  assign new_n2383_ = \C<57>  & \D<57> ;
  assign new_n2384_ = ~new_n2382_ & ~new_n2383_;
  assign new_n2385_ = ~new_n1185_1_ & ~new_n2384_;
  assign new_n2386_ = new_n1185_1_ & ~new_n2382_;
  assign new_n2387_ = ~new_n2385_ & ~new_n2386_;
  assign new_n2388_ = ~\encrypt<0>  & ~new_n2387_;
  assign new_n2389_ = \D<57>  & ~new_n1189_;
  assign new_n2390_ = ~\D<57>  & new_n1189_;
  assign new_n2391_ = ~new_n2389_ & ~new_n2390_;
  assign new_n2392_ = \C<57>  & ~new_n2391_;
  assign new_n2393_ = \D<57>  & new_n1189_;
  assign new_n2394_ = ~\C<57>  & new_n2393_;
  assign new_n2395_ = ~new_n2392_ & ~new_n2394_;
  assign new_n2396_ = \encrypt<0>  & ~new_n2395_;
  assign new_n2397_ = ~new_n2388_ & ~new_n2396_;
  assign new_n2398_ = ~\start<0>  & ~new_n2397_;
  assign n1190 = new_n2381_ | new_n2398_;
  assign new_n2400_ = \key<184>  & ~\encrypt<0> ;
  assign new_n2401_ = \key<176>  & \encrypt<0> ;
  assign new_n2402_ = ~new_n2400_ & ~new_n2401_;
  assign new_n2403_ = \start<0>  & ~new_n2402_;
  assign new_n2404_ = ~\C<56>  & ~\D<56> ;
  assign new_n2405_ = \C<56>  & \D<56> ;
  assign new_n2406_ = ~new_n2404_ & ~new_n2405_;
  assign new_n2407_ = ~new_n1185_1_ & ~new_n2406_;
  assign new_n2408_ = new_n1185_1_ & ~new_n2404_;
  assign new_n2409_ = ~new_n2407_ & ~new_n2408_;
  assign new_n2410_ = ~\encrypt<0>  & ~new_n2409_;
  assign new_n2411_ = \D<56>  & ~new_n1189_;
  assign new_n2412_ = ~\D<56>  & new_n1189_;
  assign new_n2413_ = ~new_n2411_ & ~new_n2412_;
  assign new_n2414_ = \C<56>  & ~new_n2413_;
  assign new_n2415_ = \D<56>  & new_n1189_;
  assign new_n2416_ = ~\C<56>  & new_n2415_;
  assign new_n2417_ = ~new_n2414_ & ~new_n2416_;
  assign new_n2418_ = \encrypt<0>  & ~new_n2417_;
  assign new_n2419_ = ~new_n2410_ & ~new_n2418_;
  assign new_n2420_ = ~\start<0>  & ~new_n2419_;
  assign n1195 = new_n2403_ | new_n2420_;
  assign new_n2422_ = \key<99>  & ~\encrypt<0> ;
  assign new_n2423_ = \key<184>  & \encrypt<0> ;
  assign new_n2424_ = ~new_n2422_ & ~new_n2423_;
  assign new_n2425_ = \start<0>  & ~new_n2424_;
  assign new_n2426_ = ~\C<55>  & ~\D<55> ;
  assign new_n2427_ = \C<55>  & \D<55> ;
  assign new_n2428_ = ~new_n2426_ & ~new_n2427_;
  assign new_n2429_ = ~new_n1185_1_ & ~new_n2428_;
  assign new_n2430_ = new_n1185_1_ & ~new_n2426_;
  assign new_n2431_ = ~new_n2429_ & ~new_n2430_;
  assign new_n2432_ = ~\encrypt<0>  & ~new_n2431_;
  assign new_n2433_ = \D<55>  & ~new_n1189_;
  assign new_n2434_ = ~\D<55>  & new_n1189_;
  assign new_n2435_ = ~new_n2433_ & ~new_n2434_;
  assign new_n2436_ = \C<55>  & ~new_n2435_;
  assign new_n2437_ = \D<55>  & new_n1189_;
  assign new_n2438_ = ~\C<55>  & new_n2437_;
  assign new_n2439_ = ~new_n2436_ & ~new_n2438_;
  assign new_n2440_ = \encrypt<0>  & ~new_n2439_;
  assign new_n2441_ = ~new_n2432_ & ~new_n2440_;
  assign new_n2442_ = ~\start<0>  & ~new_n2441_;
  assign n1200 = new_n2425_ | new_n2442_;
  assign new_n2444_ = \key<107>  & ~\encrypt<0> ;
  assign new_n2445_ = \key<99>  & \encrypt<0> ;
  assign new_n2446_ = ~new_n2444_ & ~new_n2445_;
  assign new_n2447_ = \start<0>  & ~new_n2446_;
  assign new_n2448_ = ~\C<54>  & ~\D<54> ;
  assign new_n2449_ = \C<54>  & \D<54> ;
  assign new_n2450_ = ~new_n2448_ & ~new_n2449_;
  assign new_n2451_ = ~new_n1185_1_ & ~new_n2450_;
  assign new_n2452_ = new_n1185_1_ & ~new_n2448_;
  assign new_n2453_ = ~new_n2451_ & ~new_n2452_;
  assign new_n2454_ = ~\encrypt<0>  & ~new_n2453_;
  assign new_n2455_ = \D<54>  & ~new_n1189_;
  assign new_n2456_ = ~\D<54>  & new_n1189_;
  assign new_n2457_ = ~new_n2455_ & ~new_n2456_;
  assign new_n2458_ = \C<54>  & ~new_n2457_;
  assign new_n2459_ = \D<54>  & new_n1189_;
  assign new_n2460_ = ~\C<54>  & new_n2459_;
  assign new_n2461_ = ~new_n2458_ & ~new_n2460_;
  assign new_n2462_ = \encrypt<0>  & ~new_n2461_;
  assign new_n2463_ = ~new_n2454_ & ~new_n2462_;
  assign new_n2464_ = ~\start<0>  & ~new_n2463_;
  assign n1205 = new_n2447_ | new_n2464_;
  assign new_n2466_ = \key<115>  & ~\encrypt<0> ;
  assign new_n2467_ = \key<107>  & \encrypt<0> ;
  assign new_n2468_ = ~new_n2466_ & ~new_n2467_;
  assign new_n2469_ = \start<0>  & ~new_n2468_;
  assign new_n2470_ = ~\C<53>  & ~\D<53> ;
  assign new_n2471_ = \C<53>  & \D<53> ;
  assign new_n2472_ = ~new_n2470_ & ~new_n2471_;
  assign new_n2473_ = ~new_n1185_1_ & ~new_n2472_;
  assign new_n2474_ = new_n1185_1_ & ~new_n2470_;
  assign new_n2475_ = ~new_n2473_ & ~new_n2474_;
  assign new_n2476_ = ~\encrypt<0>  & ~new_n2475_;
  assign new_n2477_ = \D<53>  & ~new_n1189_;
  assign new_n2478_ = ~\D<53>  & new_n1189_;
  assign new_n2479_ = ~new_n2477_ & ~new_n2478_;
  assign new_n2480_ = \C<53>  & ~new_n2479_;
  assign new_n2481_ = \D<53>  & new_n1189_;
  assign new_n2482_ = ~\C<53>  & new_n2481_;
  assign new_n2483_ = ~new_n2480_ & ~new_n2482_;
  assign new_n2484_ = \encrypt<0>  & ~new_n2483_;
  assign new_n2485_ = ~new_n2476_ & ~new_n2484_;
  assign new_n2486_ = ~\start<0>  & ~new_n2485_;
  assign n1210 = new_n2469_ | new_n2486_;
  assign new_n2488_ = \key<123>  & ~\encrypt<0> ;
  assign new_n2489_ = \key<115>  & \encrypt<0> ;
  assign new_n2490_ = ~new_n2488_ & ~new_n2489_;
  assign new_n2491_ = \start<0>  & ~new_n2490_;
  assign new_n2492_ = ~\C<52>  & ~\D<52> ;
  assign new_n2493_ = \C<52>  & \D<52> ;
  assign new_n2494_ = ~new_n2492_ & ~new_n2493_;
  assign new_n2495_ = ~new_n1185_1_ & ~new_n2494_;
  assign new_n2496_ = new_n1185_1_ & ~new_n2492_;
  assign new_n2497_ = ~new_n2495_ & ~new_n2496_;
  assign new_n2498_ = ~\encrypt<0>  & ~new_n2497_;
  assign new_n2499_ = \D<52>  & ~new_n1189_;
  assign new_n2500_ = ~\D<52>  & new_n1189_;
  assign new_n2501_ = ~new_n2499_ & ~new_n2500_;
  assign new_n2502_ = \C<52>  & ~new_n2501_;
  assign new_n2503_ = \D<52>  & new_n1189_;
  assign new_n2504_ = ~\C<52>  & new_n2503_;
  assign new_n2505_ = ~new_n2502_ & ~new_n2504_;
  assign new_n2506_ = \encrypt<0>  & ~new_n2505_;
  assign new_n2507_ = ~new_n2498_ & ~new_n2506_;
  assign new_n2508_ = ~\start<0>  & ~new_n2507_;
  assign n1215 = new_n2491_ | new_n2508_;
  assign new_n2510_ = \key<66>  & ~\encrypt<0> ;
  assign new_n2511_ = \key<123>  & \encrypt<0> ;
  assign new_n2512_ = ~new_n2510_ & ~new_n2511_;
  assign new_n2513_ = \start<0>  & ~new_n2512_;
  assign new_n2514_ = ~\C<51>  & ~\D<51> ;
  assign new_n2515_ = \C<51>  & \D<51> ;
  assign new_n2516_ = ~new_n2514_ & ~new_n2515_;
  assign new_n2517_ = ~new_n1185_1_ & ~new_n2516_;
  assign new_n2518_ = new_n1185_1_ & ~new_n2514_;
  assign new_n2519_ = ~new_n2517_ & ~new_n2518_;
  assign new_n2520_ = ~\encrypt<0>  & ~new_n2519_;
  assign new_n2521_ = \D<51>  & ~new_n1189_;
  assign new_n2522_ = ~\D<51>  & new_n1189_;
  assign new_n2523_ = ~new_n2521_ & ~new_n2522_;
  assign new_n2524_ = \C<51>  & ~new_n2523_;
  assign new_n2525_ = \D<51>  & new_n1189_;
  assign new_n2526_ = ~\C<51>  & new_n2525_;
  assign new_n2527_ = ~new_n2524_ & ~new_n2526_;
  assign new_n2528_ = \encrypt<0>  & ~new_n2527_;
  assign new_n2529_ = ~new_n2520_ & ~new_n2528_;
  assign new_n2530_ = ~\start<0>  & ~new_n2529_;
  assign n1220 = new_n2513_ | new_n2530_;
  assign new_n2532_ = \key<74>  & ~\encrypt<0> ;
  assign new_n2533_ = \key<66>  & \encrypt<0> ;
  assign new_n2534_ = ~new_n2532_ & ~new_n2533_;
  assign new_n2535_ = \start<0>  & ~new_n2534_;
  assign new_n2536_ = ~\C<50>  & ~\D<50> ;
  assign new_n2537_ = \C<50>  & \D<50> ;
  assign new_n2538_ = ~new_n2536_ & ~new_n2537_;
  assign new_n2539_ = ~new_n1185_1_ & ~new_n2538_;
  assign new_n2540_ = new_n1185_1_ & ~new_n2536_;
  assign new_n2541_ = ~new_n2539_ & ~new_n2540_;
  assign new_n2542_ = ~\encrypt<0>  & ~new_n2541_;
  assign new_n2543_ = \D<50>  & ~new_n1189_;
  assign new_n2544_ = ~\D<50>  & new_n1189_;
  assign new_n2545_ = ~new_n2543_ & ~new_n2544_;
  assign new_n2546_ = \C<50>  & ~new_n2545_;
  assign new_n2547_ = \D<50>  & new_n1189_;
  assign new_n2548_ = ~\C<50>  & new_n2547_;
  assign new_n2549_ = ~new_n2546_ & ~new_n2548_;
  assign new_n2550_ = \encrypt<0>  & ~new_n2549_;
  assign new_n2551_ = ~new_n2542_ & ~new_n2550_;
  assign new_n2552_ = ~\start<0>  & ~new_n2551_;
  assign n1225 = new_n2535_ | new_n2552_;
  assign new_n2554_ = \key<82>  & ~\encrypt<0> ;
  assign new_n2555_ = \key<74>  & \encrypt<0> ;
  assign new_n2556_ = ~new_n2554_ & ~new_n2555_;
  assign new_n2557_ = \start<0>  & ~new_n2556_;
  assign new_n2558_ = ~\C<49>  & ~\D<49> ;
  assign new_n2559_ = \C<49>  & \D<49> ;
  assign new_n2560_ = ~new_n2558_ & ~new_n2559_;
  assign new_n2561_ = ~new_n1185_1_ & ~new_n2560_;
  assign new_n2562_ = new_n1185_1_ & ~new_n2558_;
  assign new_n2563_ = ~new_n2561_ & ~new_n2562_;
  assign new_n2564_ = ~\encrypt<0>  & ~new_n2563_;
  assign new_n2565_ = \D<49>  & ~new_n1189_;
  assign new_n2566_ = ~\D<49>  & new_n1189_;
  assign new_n2567_ = ~new_n2565_ & ~new_n2566_;
  assign new_n2568_ = \C<49>  & ~new_n2567_;
  assign new_n2569_ = \D<49>  & new_n1189_;
  assign new_n2570_ = ~\C<49>  & new_n2569_;
  assign new_n2571_ = ~new_n2568_ & ~new_n2570_;
  assign new_n2572_ = \encrypt<0>  & ~new_n2571_;
  assign new_n2573_ = ~new_n2564_ & ~new_n2572_;
  assign new_n2574_ = ~\start<0>  & ~new_n2573_;
  assign n1230 = new_n2557_ | new_n2574_;
  assign new_n2576_ = \key<90>  & ~\encrypt<0> ;
  assign new_n2577_ = \key<82>  & \encrypt<0> ;
  assign new_n2578_ = ~new_n2576_ & ~new_n2577_;
  assign new_n2579_ = \start<0>  & ~new_n2578_;
  assign new_n2580_ = ~\C<48>  & ~\D<48> ;
  assign new_n2581_ = \C<48>  & \D<48> ;
  assign new_n2582_ = ~new_n2580_ & ~new_n2581_;
  assign new_n2583_ = ~new_n1185_1_ & ~new_n2582_;
  assign new_n2584_ = new_n1185_1_ & ~new_n2580_;
  assign new_n2585_ = ~new_n2583_ & ~new_n2584_;
  assign new_n2586_ = ~\encrypt<0>  & ~new_n2585_;
  assign new_n2587_ = \D<48>  & ~new_n1189_;
  assign new_n2588_ = ~\D<48>  & new_n1189_;
  assign new_n2589_ = ~new_n2587_ & ~new_n2588_;
  assign new_n2590_ = \C<48>  & ~new_n2589_;
  assign new_n2591_ = \D<48>  & new_n1189_;
  assign new_n2592_ = ~\C<48>  & new_n2591_;
  assign new_n2593_ = ~new_n2590_ & ~new_n2592_;
  assign new_n2594_ = \encrypt<0>  & ~new_n2593_;
  assign new_n2595_ = ~new_n2586_ & ~new_n2594_;
  assign new_n2596_ = ~\start<0>  & ~new_n2595_;
  assign n1235 = new_n2579_ | new_n2596_;
  assign new_n2598_ = \key<98>  & ~\encrypt<0> ;
  assign new_n2599_ = \key<90>  & \encrypt<0> ;
  assign new_n2600_ = ~new_n2598_ & ~new_n2599_;
  assign new_n2601_ = \start<0>  & ~new_n2600_;
  assign new_n2602_ = ~\C<47>  & ~\D<47> ;
  assign new_n2603_ = \C<47>  & \D<47> ;
  assign new_n2604_ = ~new_n2602_ & ~new_n2603_;
  assign new_n2605_ = ~new_n1185_1_ & ~new_n2604_;
  assign new_n2606_ = new_n1185_1_ & ~new_n2602_;
  assign new_n2607_ = ~new_n2605_ & ~new_n2606_;
  assign new_n2608_ = ~\encrypt<0>  & ~new_n2607_;
  assign new_n2609_ = \D<47>  & ~new_n1189_;
  assign new_n2610_ = ~\D<47>  & new_n1189_;
  assign new_n2611_ = ~new_n2609_ & ~new_n2610_;
  assign new_n2612_ = \C<47>  & ~new_n2611_;
  assign new_n2613_ = \D<47>  & new_n1189_;
  assign new_n2614_ = ~\C<47>  & new_n2613_;
  assign new_n2615_ = ~new_n2612_ & ~new_n2614_;
  assign new_n2616_ = \encrypt<0>  & ~new_n2615_;
  assign new_n2617_ = ~new_n2608_ & ~new_n2616_;
  assign new_n2618_ = ~\start<0>  & ~new_n2617_;
  assign n1240 = new_n2601_ | new_n2618_;
  assign new_n2620_ = \key<106>  & ~\encrypt<0> ;
  assign new_n2621_ = \key<98>  & \encrypt<0> ;
  assign new_n2622_ = ~new_n2620_ & ~new_n2621_;
  assign new_n2623_ = \start<0>  & ~new_n2622_;
  assign new_n2624_ = ~\C<46>  & ~\D<46> ;
  assign new_n2625_ = \C<46>  & \D<46> ;
  assign new_n2626_ = ~new_n2624_ & ~new_n2625_;
  assign new_n2627_ = ~new_n1185_1_ & ~new_n2626_;
  assign new_n2628_ = new_n1185_1_ & ~new_n2624_;
  assign new_n2629_ = ~new_n2627_ & ~new_n2628_;
  assign new_n2630_ = ~\encrypt<0>  & ~new_n2629_;
  assign new_n2631_ = \D<46>  & ~new_n1189_;
  assign new_n2632_ = ~\D<46>  & new_n1189_;
  assign new_n2633_ = ~new_n2631_ & ~new_n2632_;
  assign new_n2634_ = \C<46>  & ~new_n2633_;
  assign new_n2635_ = \D<46>  & new_n1189_;
  assign new_n2636_ = ~\C<46>  & new_n2635_;
  assign new_n2637_ = ~new_n2634_ & ~new_n2636_;
  assign new_n2638_ = \encrypt<0>  & ~new_n2637_;
  assign new_n2639_ = ~new_n2630_ & ~new_n2638_;
  assign new_n2640_ = ~\start<0>  & ~new_n2639_;
  assign n1245 = new_n2623_ | new_n2640_;
  assign new_n2642_ = \key<114>  & ~\encrypt<0> ;
  assign new_n2643_ = \key<106>  & \encrypt<0> ;
  assign new_n2644_ = ~new_n2642_ & ~new_n2643_;
  assign new_n2645_ = \start<0>  & ~new_n2644_;
  assign new_n2646_ = ~\C<45>  & ~\D<45> ;
  assign new_n2647_ = \C<45>  & \D<45> ;
  assign new_n2648_ = ~new_n2646_ & ~new_n2647_;
  assign new_n2649_ = ~new_n1185_1_ & ~new_n2648_;
  assign new_n2650_ = new_n1185_1_ & ~new_n2646_;
  assign new_n2651_ = ~new_n2649_ & ~new_n2650_;
  assign new_n2652_ = ~\encrypt<0>  & ~new_n2651_;
  assign new_n2653_ = \D<45>  & ~new_n1189_;
  assign new_n2654_ = ~\D<45>  & new_n1189_;
  assign new_n2655_ = ~new_n2653_ & ~new_n2654_;
  assign new_n2656_ = \C<45>  & ~new_n2655_;
  assign new_n2657_ = \D<45>  & new_n1189_;
  assign new_n2658_ = ~\C<45>  & new_n2657_;
  assign new_n2659_ = ~new_n2656_ & ~new_n2658_;
  assign new_n2660_ = \encrypt<0>  & ~new_n2659_;
  assign new_n2661_ = ~new_n2652_ & ~new_n2660_;
  assign new_n2662_ = ~\start<0>  & ~new_n2661_;
  assign n1250 = new_n2645_ | new_n2662_;
  assign new_n2664_ = \key<122>  & ~\encrypt<0> ;
  assign new_n2665_ = \key<114>  & \encrypt<0> ;
  assign new_n2666_ = ~new_n2664_ & ~new_n2665_;
  assign new_n2667_ = \start<0>  & ~new_n2666_;
  assign new_n2668_ = ~\C<44>  & ~\D<44> ;
  assign new_n2669_ = \C<44>  & \D<44> ;
  assign new_n2670_ = ~new_n2668_ & ~new_n2669_;
  assign new_n2671_ = ~new_n1185_1_ & ~new_n2670_;
  assign new_n2672_ = new_n1185_1_ & ~new_n2668_;
  assign new_n2673_ = ~new_n2671_ & ~new_n2672_;
  assign new_n2674_ = ~\encrypt<0>  & ~new_n2673_;
  assign new_n2675_ = \D<44>  & ~new_n1189_;
  assign new_n2676_ = ~\D<44>  & new_n1189_;
  assign new_n2677_ = ~new_n2675_ & ~new_n2676_;
  assign new_n2678_ = \C<44>  & ~new_n2677_;
  assign new_n2679_ = \D<44>  & new_n1189_;
  assign new_n2680_ = ~\C<44>  & new_n2679_;
  assign new_n2681_ = ~new_n2678_ & ~new_n2680_;
  assign new_n2682_ = \encrypt<0>  & ~new_n2681_;
  assign new_n2683_ = ~new_n2674_ & ~new_n2682_;
  assign new_n2684_ = ~\start<0>  & ~new_n2683_;
  assign n1255 = new_n2667_ | new_n2684_;
  assign new_n2686_ = \key<65>  & ~\encrypt<0> ;
  assign new_n2687_ = \key<122>  & \encrypt<0> ;
  assign new_n2688_ = ~new_n2686_ & ~new_n2687_;
  assign new_n2689_ = \start<0>  & ~new_n2688_;
  assign new_n2690_ = ~\C<43>  & ~\D<43> ;
  assign new_n2691_ = \C<43>  & \D<43> ;
  assign new_n2692_ = ~new_n2690_ & ~new_n2691_;
  assign new_n2693_ = ~new_n1185_1_ & ~new_n2692_;
  assign new_n2694_ = new_n1185_1_ & ~new_n2690_;
  assign new_n2695_ = ~new_n2693_ & ~new_n2694_;
  assign new_n2696_ = ~\encrypt<0>  & ~new_n2695_;
  assign new_n2697_ = \D<43>  & ~new_n1189_;
  assign new_n2698_ = ~\D<43>  & new_n1189_;
  assign new_n2699_ = ~new_n2697_ & ~new_n2698_;
  assign new_n2700_ = \C<43>  & ~new_n2699_;
  assign new_n2701_ = \D<43>  & new_n1189_;
  assign new_n2702_ = ~\C<43>  & new_n2701_;
  assign new_n2703_ = ~new_n2700_ & ~new_n2702_;
  assign new_n2704_ = \encrypt<0>  & ~new_n2703_;
  assign new_n2705_ = ~new_n2696_ & ~new_n2704_;
  assign new_n2706_ = ~\start<0>  & ~new_n2705_;
  assign n1260 = new_n2689_ | new_n2706_;
  assign new_n2708_ = \key<73>  & ~\encrypt<0> ;
  assign new_n2709_ = \key<65>  & \encrypt<0> ;
  assign new_n2710_ = ~new_n2708_ & ~new_n2709_;
  assign new_n2711_ = \start<0>  & ~new_n2710_;
  assign new_n2712_ = ~\C<42>  & ~\D<42> ;
  assign new_n2713_ = \C<42>  & \D<42> ;
  assign new_n2714_ = ~new_n2712_ & ~new_n2713_;
  assign new_n2715_ = ~new_n1185_1_ & ~new_n2714_;
  assign new_n2716_ = new_n1185_1_ & ~new_n2712_;
  assign new_n2717_ = ~new_n2715_ & ~new_n2716_;
  assign new_n2718_ = ~\encrypt<0>  & ~new_n2717_;
  assign new_n2719_ = \D<42>  & ~new_n1189_;
  assign new_n2720_ = ~\D<42>  & new_n1189_;
  assign new_n2721_ = ~new_n2719_ & ~new_n2720_;
  assign new_n2722_ = \C<42>  & ~new_n2721_;
  assign new_n2723_ = \D<42>  & new_n1189_;
  assign new_n2724_ = ~\C<42>  & new_n2723_;
  assign new_n2725_ = ~new_n2722_ & ~new_n2724_;
  assign new_n2726_ = \encrypt<0>  & ~new_n2725_;
  assign new_n2727_ = ~new_n2718_ & ~new_n2726_;
  assign new_n2728_ = ~\start<0>  & ~new_n2727_;
  assign n1265 = new_n2711_ | new_n2728_;
  assign new_n2730_ = \key<81>  & ~\encrypt<0> ;
  assign new_n2731_ = \key<73>  & \encrypt<0> ;
  assign new_n2732_ = ~new_n2730_ & ~new_n2731_;
  assign new_n2733_ = \start<0>  & ~new_n2732_;
  assign new_n2734_ = ~\C<41>  & ~\D<41> ;
  assign new_n2735_ = \C<41>  & \D<41> ;
  assign new_n2736_ = ~new_n2734_ & ~new_n2735_;
  assign new_n2737_ = ~new_n1185_1_ & ~new_n2736_;
  assign new_n2738_ = new_n1185_1_ & ~new_n2734_;
  assign new_n2739_ = ~new_n2737_ & ~new_n2738_;
  assign new_n2740_ = ~\encrypt<0>  & ~new_n2739_;
  assign new_n2741_ = \D<41>  & ~new_n1189_;
  assign new_n2742_ = ~\D<41>  & new_n1189_;
  assign new_n2743_ = ~new_n2741_ & ~new_n2742_;
  assign new_n2744_ = \C<41>  & ~new_n2743_;
  assign new_n2745_ = \D<41>  & new_n1189_;
  assign new_n2746_ = ~\C<41>  & new_n2745_;
  assign new_n2747_ = ~new_n2744_ & ~new_n2746_;
  assign new_n2748_ = \encrypt<0>  & ~new_n2747_;
  assign new_n2749_ = ~new_n2740_ & ~new_n2748_;
  assign new_n2750_ = ~\start<0>  & ~new_n2749_;
  assign n1270 = new_n2733_ | new_n2750_;
  assign new_n2752_ = \key<89>  & ~\encrypt<0> ;
  assign new_n2753_ = \key<81>  & \encrypt<0> ;
  assign new_n2754_ = ~new_n2752_ & ~new_n2753_;
  assign new_n2755_ = \start<0>  & ~new_n2754_;
  assign new_n2756_ = ~\C<40>  & ~\D<40> ;
  assign new_n2757_ = \C<40>  & \D<40> ;
  assign new_n2758_ = ~new_n2756_ & ~new_n2757_;
  assign new_n2759_ = ~new_n1185_1_ & ~new_n2758_;
  assign new_n2760_ = new_n1185_1_ & ~new_n2756_;
  assign new_n2761_ = ~new_n2759_ & ~new_n2760_;
  assign new_n2762_ = ~\encrypt<0>  & ~new_n2761_;
  assign new_n2763_ = \D<40>  & ~new_n1189_;
  assign new_n2764_ = ~\D<40>  & new_n1189_;
  assign new_n2765_ = ~new_n2763_ & ~new_n2764_;
  assign new_n2766_ = \C<40>  & ~new_n2765_;
  assign new_n2767_ = \D<40>  & new_n1189_;
  assign new_n2768_ = ~\C<40>  & new_n2767_;
  assign new_n2769_ = ~new_n2766_ & ~new_n2768_;
  assign new_n2770_ = \encrypt<0>  & ~new_n2769_;
  assign new_n2771_ = ~new_n2762_ & ~new_n2770_;
  assign new_n2772_ = ~\start<0>  & ~new_n2771_;
  assign n1275 = new_n2755_ | new_n2772_;
  assign new_n2774_ = \key<97>  & ~\encrypt<0> ;
  assign new_n2775_ = \key<89>  & \encrypt<0> ;
  assign new_n2776_ = ~new_n2774_ & ~new_n2775_;
  assign new_n2777_ = \start<0>  & ~new_n2776_;
  assign new_n2778_ = ~\C<39>  & ~\D<39> ;
  assign new_n2779_ = \C<39>  & \D<39> ;
  assign new_n2780_ = ~new_n2778_ & ~new_n2779_;
  assign new_n2781_ = ~new_n1185_1_ & ~new_n2780_;
  assign new_n2782_ = new_n1185_1_ & ~new_n2778_;
  assign new_n2783_ = ~new_n2781_ & ~new_n2782_;
  assign new_n2784_ = ~\encrypt<0>  & ~new_n2783_;
  assign new_n2785_ = \D<39>  & ~new_n1189_;
  assign new_n2786_ = ~\D<39>  & new_n1189_;
  assign new_n2787_ = ~new_n2785_ & ~new_n2786_;
  assign new_n2788_ = \C<39>  & ~new_n2787_;
  assign new_n2789_ = \D<39>  & new_n1189_;
  assign new_n2790_ = ~\C<39>  & new_n2789_;
  assign new_n2791_ = ~new_n2788_ & ~new_n2790_;
  assign new_n2792_ = \encrypt<0>  & ~new_n2791_;
  assign new_n2793_ = ~new_n2784_ & ~new_n2792_;
  assign new_n2794_ = ~\start<0>  & ~new_n2793_;
  assign n1280 = new_n2777_ | new_n2794_;
  assign new_n2796_ = \key<105>  & ~\encrypt<0> ;
  assign new_n2797_ = \key<97>  & \encrypt<0> ;
  assign new_n2798_ = ~new_n2796_ & ~new_n2797_;
  assign new_n2799_ = \start<0>  & ~new_n2798_;
  assign new_n2800_ = ~\C<38>  & ~\D<38> ;
  assign new_n2801_ = \C<38>  & \D<38> ;
  assign new_n2802_ = ~new_n2800_ & ~new_n2801_;
  assign new_n2803_ = ~new_n1185_1_ & ~new_n2802_;
  assign new_n2804_ = new_n1185_1_ & ~new_n2800_;
  assign new_n2805_ = ~new_n2803_ & ~new_n2804_;
  assign new_n2806_ = ~\encrypt<0>  & ~new_n2805_;
  assign new_n2807_ = \D<38>  & ~new_n1189_;
  assign new_n2808_ = ~\D<38>  & new_n1189_;
  assign new_n2809_ = ~new_n2807_ & ~new_n2808_;
  assign new_n2810_ = \C<38>  & ~new_n2809_;
  assign new_n2811_ = \D<38>  & new_n1189_;
  assign new_n2812_ = ~\C<38>  & new_n2811_;
  assign new_n2813_ = ~new_n2810_ & ~new_n2812_;
  assign new_n2814_ = \encrypt<0>  & ~new_n2813_;
  assign new_n2815_ = ~new_n2806_ & ~new_n2814_;
  assign new_n2816_ = ~\start<0>  & ~new_n2815_;
  assign n1285 = new_n2799_ | new_n2816_;
  assign new_n2818_ = \key<113>  & ~\encrypt<0> ;
  assign new_n2819_ = \key<105>  & \encrypt<0> ;
  assign new_n2820_ = ~new_n2818_ & ~new_n2819_;
  assign new_n2821_ = \start<0>  & ~new_n2820_;
  assign new_n2822_ = ~\C<37>  & ~\D<37> ;
  assign new_n2823_ = \C<37>  & \D<37> ;
  assign new_n2824_ = ~new_n2822_ & ~new_n2823_;
  assign new_n2825_ = ~new_n1185_1_ & ~new_n2824_;
  assign new_n2826_ = new_n1185_1_ & ~new_n2822_;
  assign new_n2827_ = ~new_n2825_ & ~new_n2826_;
  assign new_n2828_ = ~\encrypt<0>  & ~new_n2827_;
  assign new_n2829_ = \D<37>  & ~new_n1189_;
  assign new_n2830_ = ~\D<37>  & new_n1189_;
  assign new_n2831_ = ~new_n2829_ & ~new_n2830_;
  assign new_n2832_ = \C<37>  & ~new_n2831_;
  assign new_n2833_ = \D<37>  & new_n1189_;
  assign new_n2834_ = ~\C<37>  & new_n2833_;
  assign new_n2835_ = ~new_n2832_ & ~new_n2834_;
  assign new_n2836_ = \encrypt<0>  & ~new_n2835_;
  assign new_n2837_ = ~new_n2828_ & ~new_n2836_;
  assign new_n2838_ = ~\start<0>  & ~new_n2837_;
  assign n1290 = new_n2821_ | new_n2838_;
  assign new_n2840_ = \key<121>  & ~\encrypt<0> ;
  assign new_n2841_ = \key<113>  & \encrypt<0> ;
  assign new_n2842_ = ~new_n2840_ & ~new_n2841_;
  assign new_n2843_ = \start<0>  & ~new_n2842_;
  assign new_n2844_ = ~\C<36>  & ~\D<36> ;
  assign new_n2845_ = \C<36>  & \D<36> ;
  assign new_n2846_ = ~new_n2844_ & ~new_n2845_;
  assign new_n2847_ = ~new_n1185_1_ & ~new_n2846_;
  assign new_n2848_ = new_n1185_1_ & ~new_n2844_;
  assign new_n2849_ = ~new_n2847_ & ~new_n2848_;
  assign new_n2850_ = ~\encrypt<0>  & ~new_n2849_;
  assign new_n2851_ = \D<36>  & ~new_n1189_;
  assign new_n2852_ = ~\D<36>  & new_n1189_;
  assign new_n2853_ = ~new_n2851_ & ~new_n2852_;
  assign new_n2854_ = \C<36>  & ~new_n2853_;
  assign new_n2855_ = \D<36>  & new_n1189_;
  assign new_n2856_ = ~\C<36>  & new_n2855_;
  assign new_n2857_ = ~new_n2854_ & ~new_n2856_;
  assign new_n2858_ = \encrypt<0>  & ~new_n2857_;
  assign new_n2859_ = ~new_n2850_ & ~new_n2858_;
  assign new_n2860_ = ~\start<0>  & ~new_n2859_;
  assign n1295 = new_n2843_ | new_n2860_;
  assign new_n2862_ = \key<64>  & ~\encrypt<0> ;
  assign new_n2863_ = \key<121>  & \encrypt<0> ;
  assign new_n2864_ = ~new_n2862_ & ~new_n2863_;
  assign new_n2865_ = \start<0>  & ~new_n2864_;
  assign new_n2866_ = ~\C<35>  & ~\D<35> ;
  assign new_n2867_ = \C<35>  & \D<35> ;
  assign new_n2868_ = ~new_n2866_ & ~new_n2867_;
  assign new_n2869_ = ~new_n1185_1_ & ~new_n2868_;
  assign new_n2870_ = new_n1185_1_ & ~new_n2866_;
  assign new_n2871_ = ~new_n2869_ & ~new_n2870_;
  assign new_n2872_ = ~\encrypt<0>  & ~new_n2871_;
  assign new_n2873_ = \D<35>  & ~new_n1189_;
  assign new_n2874_ = ~\D<35>  & new_n1189_;
  assign new_n2875_ = ~new_n2873_ & ~new_n2874_;
  assign new_n2876_ = \C<35>  & ~new_n2875_;
  assign new_n2877_ = \D<35>  & new_n1189_;
  assign new_n2878_ = ~\C<35>  & new_n2877_;
  assign new_n2879_ = ~new_n2876_ & ~new_n2878_;
  assign new_n2880_ = \encrypt<0>  & ~new_n2879_;
  assign new_n2881_ = ~new_n2872_ & ~new_n2880_;
  assign new_n2882_ = ~\start<0>  & ~new_n2881_;
  assign n1300 = new_n2865_ | new_n2882_;
  assign new_n2884_ = \key<72>  & ~\encrypt<0> ;
  assign new_n2885_ = \key<64>  & \encrypt<0> ;
  assign new_n2886_ = ~new_n2884_ & ~new_n2885_;
  assign new_n2887_ = \start<0>  & ~new_n2886_;
  assign new_n2888_ = ~\C<34>  & ~\D<34> ;
  assign new_n2889_ = \C<34>  & \D<34> ;
  assign new_n2890_ = ~new_n2888_ & ~new_n2889_;
  assign new_n2891_ = ~new_n1185_1_ & ~new_n2890_;
  assign new_n2892_ = new_n1185_1_ & ~new_n2888_;
  assign new_n2893_ = ~new_n2891_ & ~new_n2892_;
  assign new_n2894_ = ~\encrypt<0>  & ~new_n2893_;
  assign new_n2895_ = \D<34>  & ~new_n1189_;
  assign new_n2896_ = ~\D<34>  & new_n1189_;
  assign new_n2897_ = ~new_n2895_ & ~new_n2896_;
  assign new_n2898_ = \C<34>  & ~new_n2897_;
  assign new_n2899_ = \D<34>  & new_n1189_;
  assign new_n2900_ = ~\C<34>  & new_n2899_;
  assign new_n2901_ = ~new_n2898_ & ~new_n2900_;
  assign new_n2902_ = \encrypt<0>  & ~new_n2901_;
  assign new_n2903_ = ~new_n2894_ & ~new_n2902_;
  assign new_n2904_ = ~\start<0>  & ~new_n2903_;
  assign n1305 = new_n2887_ | new_n2904_;
  assign new_n2906_ = \key<80>  & ~\encrypt<0> ;
  assign new_n2907_ = \key<72>  & \encrypt<0> ;
  assign new_n2908_ = ~new_n2906_ & ~new_n2907_;
  assign new_n2909_ = \start<0>  & ~new_n2908_;
  assign new_n2910_ = ~\C<33>  & ~\D<33> ;
  assign new_n2911_ = \C<33>  & \D<33> ;
  assign new_n2912_ = ~new_n2910_ & ~new_n2911_;
  assign new_n2913_ = ~new_n1185_1_ & ~new_n2912_;
  assign new_n2914_ = new_n1185_1_ & ~new_n2910_;
  assign new_n2915_ = ~new_n2913_ & ~new_n2914_;
  assign new_n2916_ = ~\encrypt<0>  & ~new_n2915_;
  assign new_n2917_ = \D<33>  & ~new_n1189_;
  assign new_n2918_ = ~\D<33>  & new_n1189_;
  assign new_n2919_ = ~new_n2917_ & ~new_n2918_;
  assign new_n2920_ = \C<33>  & ~new_n2919_;
  assign new_n2921_ = \D<33>  & new_n1189_;
  assign new_n2922_ = ~\C<33>  & new_n2921_;
  assign new_n2923_ = ~new_n2920_ & ~new_n2922_;
  assign new_n2924_ = \encrypt<0>  & ~new_n2923_;
  assign new_n2925_ = ~new_n2916_ & ~new_n2924_;
  assign new_n2926_ = ~\start<0>  & ~new_n2925_;
  assign n1310 = new_n2909_ | new_n2926_;
  assign new_n2928_ = \key<88>  & ~\encrypt<0> ;
  assign new_n2929_ = \key<80>  & \encrypt<0> ;
  assign new_n2930_ = ~new_n2928_ & ~new_n2929_;
  assign new_n2931_ = \start<0>  & ~new_n2930_;
  assign new_n2932_ = ~\C<32>  & ~\D<32> ;
  assign new_n2933_ = \C<32>  & \D<32> ;
  assign new_n2934_ = ~new_n2932_ & ~new_n2933_;
  assign new_n2935_ = ~new_n1185_1_ & ~new_n2934_;
  assign new_n2936_ = new_n1185_1_ & ~new_n2932_;
  assign new_n2937_ = ~new_n2935_ & ~new_n2936_;
  assign new_n2938_ = ~\encrypt<0>  & ~new_n2937_;
  assign new_n2939_ = \D<32>  & ~new_n1189_;
  assign new_n2940_ = ~\D<32>  & new_n1189_;
  assign new_n2941_ = ~new_n2939_ & ~new_n2940_;
  assign new_n2942_ = \C<32>  & ~new_n2941_;
  assign new_n2943_ = \D<32>  & new_n1189_;
  assign new_n2944_ = ~\C<32>  & new_n2943_;
  assign new_n2945_ = ~new_n2942_ & ~new_n2944_;
  assign new_n2946_ = \encrypt<0>  & ~new_n2945_;
  assign new_n2947_ = ~new_n2938_ & ~new_n2946_;
  assign new_n2948_ = ~\start<0>  & ~new_n2947_;
  assign n1315 = new_n2931_ | new_n2948_;
  assign new_n2950_ = \key<96>  & ~\encrypt<0> ;
  assign new_n2951_ = \key<88>  & \encrypt<0> ;
  assign new_n2952_ = ~new_n2950_ & ~new_n2951_;
  assign new_n2953_ = \start<0>  & ~new_n2952_;
  assign new_n2954_ = ~\C<31>  & ~\D<31> ;
  assign new_n2955_ = \C<31>  & \D<31> ;
  assign new_n2956_ = ~new_n2954_ & ~new_n2955_;
  assign new_n2957_ = ~new_n1185_1_ & ~new_n2956_;
  assign new_n2958_ = new_n1185_1_ & ~new_n2954_;
  assign new_n2959_ = ~new_n2957_ & ~new_n2958_;
  assign new_n2960_ = ~\encrypt<0>  & ~new_n2959_;
  assign new_n2961_ = \D<31>  & ~new_n1189_;
  assign new_n2962_ = ~\D<31>  & new_n1189_;
  assign new_n2963_ = ~new_n2961_ & ~new_n2962_;
  assign new_n2964_ = \C<31>  & ~new_n2963_;
  assign new_n2965_ = \D<31>  & new_n1189_;
  assign new_n2966_ = ~\C<31>  & new_n2965_;
  assign new_n2967_ = ~new_n2964_ & ~new_n2966_;
  assign new_n2968_ = \encrypt<0>  & ~new_n2967_;
  assign new_n2969_ = ~new_n2960_ & ~new_n2968_;
  assign new_n2970_ = ~\start<0>  & ~new_n2969_;
  assign n1320 = new_n2953_ | new_n2970_;
  assign new_n2972_ = \key<104>  & ~\encrypt<0> ;
  assign new_n2973_ = \key<96>  & \encrypt<0> ;
  assign new_n2974_ = ~new_n2972_ & ~new_n2973_;
  assign new_n2975_ = \start<0>  & ~new_n2974_;
  assign new_n2976_ = ~\C<30>  & ~\D<30> ;
  assign new_n2977_ = \C<30>  & \D<30> ;
  assign new_n2978_ = ~new_n2976_ & ~new_n2977_;
  assign new_n2979_ = ~new_n1185_1_ & ~new_n2978_;
  assign new_n2980_ = new_n1185_1_ & ~new_n2976_;
  assign new_n2981_ = ~new_n2979_ & ~new_n2980_;
  assign new_n2982_ = ~\encrypt<0>  & ~new_n2981_;
  assign new_n2983_ = \D<30>  & ~new_n1189_;
  assign new_n2984_ = ~\D<30>  & new_n1189_;
  assign new_n2985_ = ~new_n2983_ & ~new_n2984_;
  assign new_n2986_ = \C<30>  & ~new_n2985_;
  assign new_n2987_ = \D<30>  & new_n1189_;
  assign new_n2988_ = ~\C<30>  & new_n2987_;
  assign new_n2989_ = ~new_n2986_ & ~new_n2988_;
  assign new_n2990_ = \encrypt<0>  & ~new_n2989_;
  assign new_n2991_ = ~new_n2982_ & ~new_n2990_;
  assign new_n2992_ = ~\start<0>  & ~new_n2991_;
  assign n1325 = new_n2975_ | new_n2992_;
  assign new_n2994_ = \key<112>  & ~\encrypt<0> ;
  assign new_n2995_ = \key<104>  & \encrypt<0> ;
  assign new_n2996_ = ~new_n2994_ & ~new_n2995_;
  assign new_n2997_ = \start<0>  & ~new_n2996_;
  assign new_n2998_ = ~\C<29>  & ~\D<29> ;
  assign new_n2999_ = \C<29>  & \D<29> ;
  assign new_n3000_ = ~new_n2998_ & ~new_n2999_;
  assign new_n3001_ = ~new_n1185_1_ & ~new_n3000_;
  assign new_n3002_ = new_n1185_1_ & ~new_n2998_;
  assign new_n3003_ = ~new_n3001_ & ~new_n3002_;
  assign new_n3004_ = ~\encrypt<0>  & ~new_n3003_;
  assign new_n3005_ = \D<29>  & ~new_n1189_;
  assign new_n3006_ = ~\D<29>  & new_n1189_;
  assign new_n3007_ = ~new_n3005_ & ~new_n3006_;
  assign new_n3008_ = \C<29>  & ~new_n3007_;
  assign new_n3009_ = \D<29>  & new_n1189_;
  assign new_n3010_ = ~\C<29>  & new_n3009_;
  assign new_n3011_ = ~new_n3008_ & ~new_n3010_;
  assign new_n3012_ = \encrypt<0>  & ~new_n3011_;
  assign new_n3013_ = ~new_n3004_ & ~new_n3012_;
  assign new_n3014_ = ~\start<0>  & ~new_n3013_;
  assign n1330 = new_n2997_ | new_n3014_;
  assign new_n3016_ = \key<120>  & ~\encrypt<0> ;
  assign new_n3017_ = \key<112>  & \encrypt<0> ;
  assign new_n3018_ = ~new_n3016_ & ~new_n3017_;
  assign new_n3019_ = \start<0>  & ~new_n3018_;
  assign new_n3020_ = ~\C<28>  & ~\D<28> ;
  assign new_n3021_ = \C<28>  & \D<28> ;
  assign new_n3022_ = ~new_n3020_ & ~new_n3021_;
  assign new_n3023_ = ~new_n1185_1_ & ~new_n3022_;
  assign new_n3024_ = new_n1185_1_ & ~new_n3020_;
  assign new_n3025_ = ~new_n3023_ & ~new_n3024_;
  assign new_n3026_ = ~\encrypt<0>  & ~new_n3025_;
  assign new_n3027_ = \D<28>  & ~new_n1189_;
  assign new_n3028_ = ~\D<28>  & new_n1189_;
  assign new_n3029_ = ~new_n3027_ & ~new_n3028_;
  assign new_n3030_ = \C<28>  & ~new_n3029_;
  assign new_n3031_ = \D<28>  & new_n1189_;
  assign new_n3032_ = ~\C<28>  & new_n3031_;
  assign new_n3033_ = ~new_n3030_ & ~new_n3032_;
  assign new_n3034_ = \encrypt<0>  & ~new_n3033_;
  assign new_n3035_ = ~new_n3026_ & ~new_n3034_;
  assign new_n3036_ = ~\start<0>  & ~new_n3035_;
  assign n1335 = new_n3019_ | new_n3036_;
  assign new_n3038_ = \key<35>  & ~\encrypt<0> ;
  assign new_n3039_ = \key<120>  & \encrypt<0> ;
  assign new_n3040_ = ~new_n3038_ & ~new_n3039_;
  assign new_n3041_ = \start<0>  & ~new_n3040_;
  assign new_n3042_ = ~\C<27>  & ~\D<27> ;
  assign new_n3043_ = \C<27>  & \D<27> ;
  assign new_n3044_ = ~new_n3042_ & ~new_n3043_;
  assign new_n3045_ = ~new_n1185_1_ & ~new_n3044_;
  assign new_n3046_ = new_n1185_1_ & ~new_n3042_;
  assign new_n3047_ = ~new_n3045_ & ~new_n3046_;
  assign new_n3048_ = ~\encrypt<0>  & ~new_n3047_;
  assign new_n3049_ = \D<27>  & ~new_n1189_;
  assign new_n3050_ = ~\D<27>  & new_n1189_;
  assign new_n3051_ = ~new_n3049_ & ~new_n3050_;
  assign new_n3052_ = \C<27>  & ~new_n3051_;
  assign new_n3053_ = \D<27>  & new_n1189_;
  assign new_n3054_ = ~\C<27>  & new_n3053_;
  assign new_n3055_ = ~new_n3052_ & ~new_n3054_;
  assign new_n3056_ = \encrypt<0>  & ~new_n3055_;
  assign new_n3057_ = ~new_n3048_ & ~new_n3056_;
  assign new_n3058_ = ~\start<0>  & ~new_n3057_;
  assign n1340 = new_n3041_ | new_n3058_;
  assign new_n3060_ = \key<43>  & ~\encrypt<0> ;
  assign new_n3061_ = \key<35>  & \encrypt<0> ;
  assign new_n3062_ = ~new_n3060_ & ~new_n3061_;
  assign new_n3063_ = \start<0>  & ~new_n3062_;
  assign new_n3064_ = ~\C<26>  & ~\D<26> ;
  assign new_n3065_ = \C<26>  & \D<26> ;
  assign new_n3066_ = ~new_n3064_ & ~new_n3065_;
  assign new_n3067_ = ~new_n1185_1_ & ~new_n3066_;
  assign new_n3068_ = new_n1185_1_ & ~new_n3064_;
  assign new_n3069_ = ~new_n3067_ & ~new_n3068_;
  assign new_n3070_ = ~\encrypt<0>  & ~new_n3069_;
  assign new_n3071_ = \D<26>  & ~new_n1189_;
  assign new_n3072_ = ~\D<26>  & new_n1189_;
  assign new_n3073_ = ~new_n3071_ & ~new_n3072_;
  assign new_n3074_ = \C<26>  & ~new_n3073_;
  assign new_n3075_ = \D<26>  & new_n1189_;
  assign new_n3076_ = ~\C<26>  & new_n3075_;
  assign new_n3077_ = ~new_n3074_ & ~new_n3076_;
  assign new_n3078_ = \encrypt<0>  & ~new_n3077_;
  assign new_n3079_ = ~new_n3070_ & ~new_n3078_;
  assign new_n3080_ = ~\start<0>  & ~new_n3079_;
  assign n1345 = new_n3063_ | new_n3080_;
  assign new_n3082_ = \key<51>  & ~\encrypt<0> ;
  assign new_n3083_ = \key<43>  & \encrypt<0> ;
  assign new_n3084_ = ~new_n3082_ & ~new_n3083_;
  assign new_n3085_ = \start<0>  & ~new_n3084_;
  assign new_n3086_ = ~\C<25>  & ~\D<25> ;
  assign new_n3087_ = \C<25>  & \D<25> ;
  assign new_n3088_ = ~new_n3086_ & ~new_n3087_;
  assign new_n3089_ = ~new_n1185_1_ & ~new_n3088_;
  assign new_n3090_ = new_n1185_1_ & ~new_n3086_;
  assign new_n3091_ = ~new_n3089_ & ~new_n3090_;
  assign new_n3092_ = ~\encrypt<0>  & ~new_n3091_;
  assign new_n3093_ = \D<25>  & ~new_n1189_;
  assign new_n3094_ = ~\D<25>  & new_n1189_;
  assign new_n3095_ = ~new_n3093_ & ~new_n3094_;
  assign new_n3096_ = \C<25>  & ~new_n3095_;
  assign new_n3097_ = \D<25>  & new_n1189_;
  assign new_n3098_ = ~\C<25>  & new_n3097_;
  assign new_n3099_ = ~new_n3096_ & ~new_n3098_;
  assign new_n3100_ = \encrypt<0>  & ~new_n3099_;
  assign new_n3101_ = ~new_n3092_ & ~new_n3100_;
  assign new_n3102_ = ~\start<0>  & ~new_n3101_;
  assign n1350 = new_n3085_ | new_n3102_;
  assign new_n3104_ = \key<59>  & ~\encrypt<0> ;
  assign new_n3105_ = \key<51>  & \encrypt<0> ;
  assign new_n3106_ = ~new_n3104_ & ~new_n3105_;
  assign new_n3107_ = \start<0>  & ~new_n3106_;
  assign new_n3108_ = ~\C<24>  & ~\D<24> ;
  assign new_n3109_ = \C<24>  & \D<24> ;
  assign new_n3110_ = ~new_n3108_ & ~new_n3109_;
  assign new_n3111_ = ~new_n1185_1_ & ~new_n3110_;
  assign new_n3112_ = new_n1185_1_ & ~new_n3108_;
  assign new_n3113_ = ~new_n3111_ & ~new_n3112_;
  assign new_n3114_ = ~\encrypt<0>  & ~new_n3113_;
  assign new_n3115_ = \D<24>  & ~new_n1189_;
  assign new_n3116_ = ~\D<24>  & new_n1189_;
  assign new_n3117_ = ~new_n3115_ & ~new_n3116_;
  assign new_n3118_ = \C<24>  & ~new_n3117_;
  assign new_n3119_ = \D<24>  & new_n1189_;
  assign new_n3120_ = ~\C<24>  & new_n3119_;
  assign new_n3121_ = ~new_n3118_ & ~new_n3120_;
  assign new_n3122_ = \encrypt<0>  & ~new_n3121_;
  assign new_n3123_ = ~new_n3114_ & ~new_n3122_;
  assign new_n3124_ = ~\start<0>  & ~new_n3123_;
  assign n1355 = new_n3107_ | new_n3124_;
  assign new_n3126_ = \key<2>  & ~\encrypt<0> ;
  assign new_n3127_ = \key<59>  & \encrypt<0> ;
  assign new_n3128_ = ~new_n3126_ & ~new_n3127_;
  assign new_n3129_ = \start<0>  & ~new_n3128_;
  assign new_n3130_ = ~\C<23>  & ~\D<23> ;
  assign new_n3131_ = \C<23>  & \D<23> ;
  assign new_n3132_ = ~new_n3130_ & ~new_n3131_;
  assign new_n3133_ = ~new_n1185_1_ & ~new_n3132_;
  assign new_n3134_ = new_n1185_1_ & ~new_n3130_;
  assign new_n3135_ = ~new_n3133_ & ~new_n3134_;
  assign new_n3136_ = ~\encrypt<0>  & ~new_n3135_;
  assign new_n3137_ = \D<23>  & ~new_n1189_;
  assign new_n3138_ = ~\D<23>  & new_n1189_;
  assign new_n3139_ = ~new_n3137_ & ~new_n3138_;
  assign new_n3140_ = \C<23>  & ~new_n3139_;
  assign new_n3141_ = \D<23>  & new_n1189_;
  assign new_n3142_ = ~\C<23>  & new_n3141_;
  assign new_n3143_ = ~new_n3140_ & ~new_n3142_;
  assign new_n3144_ = \encrypt<0>  & ~new_n3143_;
  assign new_n3145_ = ~new_n3136_ & ~new_n3144_;
  assign new_n3146_ = ~\start<0>  & ~new_n3145_;
  assign n1360 = new_n3129_ | new_n3146_;
  assign new_n3148_ = \key<10>  & ~\encrypt<0> ;
  assign new_n3149_ = \key<2>  & \encrypt<0> ;
  assign new_n3150_ = ~new_n3148_ & ~new_n3149_;
  assign new_n3151_ = \start<0>  & ~new_n3150_;
  assign new_n3152_ = ~\C<22>  & ~\D<22> ;
  assign new_n3153_ = \C<22>  & \D<22> ;
  assign new_n3154_ = ~new_n3152_ & ~new_n3153_;
  assign new_n3155_ = ~new_n1185_1_ & ~new_n3154_;
  assign new_n3156_ = new_n1185_1_ & ~new_n3152_;
  assign new_n3157_ = ~new_n3155_ & ~new_n3156_;
  assign new_n3158_ = ~\encrypt<0>  & ~new_n3157_;
  assign new_n3159_ = \D<22>  & ~new_n1189_;
  assign new_n3160_ = ~\D<22>  & new_n1189_;
  assign new_n3161_ = ~new_n3159_ & ~new_n3160_;
  assign new_n3162_ = \C<22>  & ~new_n3161_;
  assign new_n3163_ = \D<22>  & new_n1189_;
  assign new_n3164_ = ~\C<22>  & new_n3163_;
  assign new_n3165_ = ~new_n3162_ & ~new_n3164_;
  assign new_n3166_ = \encrypt<0>  & ~new_n3165_;
  assign new_n3167_ = ~new_n3158_ & ~new_n3166_;
  assign new_n3168_ = ~\start<0>  & ~new_n3167_;
  assign n1365 = new_n3151_ | new_n3168_;
  assign new_n3170_ = \key<18>  & ~\encrypt<0> ;
  assign new_n3171_ = \key<10>  & \encrypt<0> ;
  assign new_n3172_ = ~new_n3170_ & ~new_n3171_;
  assign new_n3173_ = \start<0>  & ~new_n3172_;
  assign new_n3174_ = ~\C<21>  & ~\D<21> ;
  assign new_n3175_ = \C<21>  & \D<21> ;
  assign new_n3176_ = ~new_n3174_ & ~new_n3175_;
  assign new_n3177_ = ~new_n1185_1_ & ~new_n3176_;
  assign new_n3178_ = new_n1185_1_ & ~new_n3174_;
  assign new_n3179_ = ~new_n3177_ & ~new_n3178_;
  assign new_n3180_ = ~\encrypt<0>  & ~new_n3179_;
  assign new_n3181_ = \D<21>  & ~new_n1189_;
  assign new_n3182_ = ~\D<21>  & new_n1189_;
  assign new_n3183_ = ~new_n3181_ & ~new_n3182_;
  assign new_n3184_ = \C<21>  & ~new_n3183_;
  assign new_n3185_ = \D<21>  & new_n1189_;
  assign new_n3186_ = ~\C<21>  & new_n3185_;
  assign new_n3187_ = ~new_n3184_ & ~new_n3186_;
  assign new_n3188_ = \encrypt<0>  & ~new_n3187_;
  assign new_n3189_ = ~new_n3180_ & ~new_n3188_;
  assign new_n3190_ = ~\start<0>  & ~new_n3189_;
  assign n1370 = new_n3173_ | new_n3190_;
  assign new_n3192_ = \key<26>  & ~\encrypt<0> ;
  assign new_n3193_ = \key<18>  & \encrypt<0> ;
  assign new_n3194_ = ~new_n3192_ & ~new_n3193_;
  assign new_n3195_ = \start<0>  & ~new_n3194_;
  assign new_n3196_ = ~\C<20>  & ~\D<20> ;
  assign new_n3197_ = \C<20>  & \D<20> ;
  assign new_n3198_ = ~new_n3196_ & ~new_n3197_;
  assign new_n3199_ = ~new_n1185_1_ & ~new_n3198_;
  assign new_n3200_ = new_n1185_1_ & ~new_n3196_;
  assign new_n3201_ = ~new_n3199_ & ~new_n3200_;
  assign new_n3202_ = ~\encrypt<0>  & ~new_n3201_;
  assign new_n3203_ = \D<20>  & ~new_n1189_;
  assign new_n3204_ = ~\D<20>  & new_n1189_;
  assign new_n3205_ = ~new_n3203_ & ~new_n3204_;
  assign new_n3206_ = \C<20>  & ~new_n3205_;
  assign new_n3207_ = \D<20>  & new_n1189_;
  assign new_n3208_ = ~\C<20>  & new_n3207_;
  assign new_n3209_ = ~new_n3206_ & ~new_n3208_;
  assign new_n3210_ = \encrypt<0>  & ~new_n3209_;
  assign new_n3211_ = ~new_n3202_ & ~new_n3210_;
  assign new_n3212_ = ~\start<0>  & ~new_n3211_;
  assign n1375 = new_n3195_ | new_n3212_;
  assign new_n3214_ = \key<34>  & ~\encrypt<0> ;
  assign new_n3215_ = \key<26>  & \encrypt<0> ;
  assign new_n3216_ = ~new_n3214_ & ~new_n3215_;
  assign new_n3217_ = \start<0>  & ~new_n3216_;
  assign new_n3218_ = ~\C<19>  & ~\D<19> ;
  assign new_n3219_ = \C<19>  & \D<19> ;
  assign new_n3220_ = ~new_n3218_ & ~new_n3219_;
  assign new_n3221_ = ~new_n1185_1_ & ~new_n3220_;
  assign new_n3222_ = new_n1185_1_ & ~new_n3218_;
  assign new_n3223_ = ~new_n3221_ & ~new_n3222_;
  assign new_n3224_ = ~\encrypt<0>  & ~new_n3223_;
  assign new_n3225_ = \D<19>  & ~new_n1189_;
  assign new_n3226_ = ~\D<19>  & new_n1189_;
  assign new_n3227_ = ~new_n3225_ & ~new_n3226_;
  assign new_n3228_ = \C<19>  & ~new_n3227_;
  assign new_n3229_ = \D<19>  & new_n1189_;
  assign new_n3230_ = ~\C<19>  & new_n3229_;
  assign new_n3231_ = ~new_n3228_ & ~new_n3230_;
  assign new_n3232_ = \encrypt<0>  & ~new_n3231_;
  assign new_n3233_ = ~new_n3224_ & ~new_n3232_;
  assign new_n3234_ = ~\start<0>  & ~new_n3233_;
  assign n1380 = new_n3217_ | new_n3234_;
  assign new_n3236_ = \key<42>  & ~\encrypt<0> ;
  assign new_n3237_ = \key<34>  & \encrypt<0> ;
  assign new_n3238_ = ~new_n3236_ & ~new_n3237_;
  assign new_n3239_ = \start<0>  & ~new_n3238_;
  assign new_n3240_ = ~\C<18>  & ~\D<18> ;
  assign new_n3241_ = \C<18>  & \D<18> ;
  assign new_n3242_ = ~new_n3240_ & ~new_n3241_;
  assign new_n3243_ = ~new_n1185_1_ & ~new_n3242_;
  assign new_n3244_ = new_n1185_1_ & ~new_n3240_;
  assign new_n3245_ = ~new_n3243_ & ~new_n3244_;
  assign new_n3246_ = ~\encrypt<0>  & ~new_n3245_;
  assign new_n3247_ = \D<18>  & ~new_n1189_;
  assign new_n3248_ = ~\D<18>  & new_n1189_;
  assign new_n3249_ = ~new_n3247_ & ~new_n3248_;
  assign new_n3250_ = \C<18>  & ~new_n3249_;
  assign new_n3251_ = \D<18>  & new_n1189_;
  assign new_n3252_ = ~\C<18>  & new_n3251_;
  assign new_n3253_ = ~new_n3250_ & ~new_n3252_;
  assign new_n3254_ = \encrypt<0>  & ~new_n3253_;
  assign new_n3255_ = ~new_n3246_ & ~new_n3254_;
  assign new_n3256_ = ~\start<0>  & ~new_n3255_;
  assign n1385 = new_n3239_ | new_n3256_;
  assign new_n3258_ = \key<50>  & ~\encrypt<0> ;
  assign new_n3259_ = \key<42>  & \encrypt<0> ;
  assign new_n3260_ = ~new_n3258_ & ~new_n3259_;
  assign new_n3261_ = \start<0>  & ~new_n3260_;
  assign new_n3262_ = ~\C<17>  & ~\D<17> ;
  assign new_n3263_ = \C<17>  & \D<17> ;
  assign new_n3264_ = ~new_n3262_ & ~new_n3263_;
  assign new_n3265_ = ~new_n1185_1_ & ~new_n3264_;
  assign new_n3266_ = new_n1185_1_ & ~new_n3262_;
  assign new_n3267_ = ~new_n3265_ & ~new_n3266_;
  assign new_n3268_ = ~\encrypt<0>  & ~new_n3267_;
  assign new_n3269_ = \D<17>  & ~new_n1189_;
  assign new_n3270_ = ~\D<17>  & new_n1189_;
  assign new_n3271_ = ~new_n3269_ & ~new_n3270_;
  assign new_n3272_ = \C<17>  & ~new_n3271_;
  assign new_n3273_ = \D<17>  & new_n1189_;
  assign new_n3274_ = ~\C<17>  & new_n3273_;
  assign new_n3275_ = ~new_n3272_ & ~new_n3274_;
  assign new_n3276_ = \encrypt<0>  & ~new_n3275_;
  assign new_n3277_ = ~new_n3268_ & ~new_n3276_;
  assign new_n3278_ = ~\start<0>  & ~new_n3277_;
  assign n1390 = new_n3261_ | new_n3278_;
  assign new_n3280_ = \key<58>  & ~\encrypt<0> ;
  assign new_n3281_ = \key<50>  & \encrypt<0> ;
  assign new_n3282_ = ~new_n3280_ & ~new_n3281_;
  assign new_n3283_ = \start<0>  & ~new_n3282_;
  assign new_n3284_ = ~\C<16>  & ~\D<16> ;
  assign new_n3285_ = \C<16>  & \D<16> ;
  assign new_n3286_ = ~new_n3284_ & ~new_n3285_;
  assign new_n3287_ = ~new_n1185_1_ & ~new_n3286_;
  assign new_n3288_ = new_n1185_1_ & ~new_n3284_;
  assign new_n3289_ = ~new_n3287_ & ~new_n3288_;
  assign new_n3290_ = ~\encrypt<0>  & ~new_n3289_;
  assign new_n3291_ = \D<16>  & ~new_n1189_;
  assign new_n3292_ = ~\D<16>  & new_n1189_;
  assign new_n3293_ = ~new_n3291_ & ~new_n3292_;
  assign new_n3294_ = \C<16>  & ~new_n3293_;
  assign new_n3295_ = \D<16>  & new_n1189_;
  assign new_n3296_ = ~\C<16>  & new_n3295_;
  assign new_n3297_ = ~new_n3294_ & ~new_n3296_;
  assign new_n3298_ = \encrypt<0>  & ~new_n3297_;
  assign new_n3299_ = ~new_n3290_ & ~new_n3298_;
  assign new_n3300_ = ~\start<0>  & ~new_n3299_;
  assign n1395 = new_n3283_ | new_n3300_;
  assign new_n3302_ = \key<1>  & ~\encrypt<0> ;
  assign new_n3303_ = \key<58>  & \encrypt<0> ;
  assign new_n3304_ = ~new_n3302_ & ~new_n3303_;
  assign new_n3305_ = \start<0>  & ~new_n3304_;
  assign new_n3306_ = ~\C<15>  & ~\D<15> ;
  assign new_n3307_ = \C<15>  & \D<15> ;
  assign new_n3308_ = ~new_n3306_ & ~new_n3307_;
  assign new_n3309_ = ~new_n1185_1_ & ~new_n3308_;
  assign new_n3310_ = new_n1185_1_ & ~new_n3306_;
  assign new_n3311_ = ~new_n3309_ & ~new_n3310_;
  assign new_n3312_ = ~\encrypt<0>  & ~new_n3311_;
  assign new_n3313_ = \D<15>  & ~new_n1189_;
  assign new_n3314_ = ~\D<15>  & new_n1189_;
  assign new_n3315_ = ~new_n3313_ & ~new_n3314_;
  assign new_n3316_ = \C<15>  & ~new_n3315_;
  assign new_n3317_ = \D<15>  & new_n1189_;
  assign new_n3318_ = ~\C<15>  & new_n3317_;
  assign new_n3319_ = ~new_n3316_ & ~new_n3318_;
  assign new_n3320_ = \encrypt<0>  & ~new_n3319_;
  assign new_n3321_ = ~new_n3312_ & ~new_n3320_;
  assign new_n3322_ = ~\start<0>  & ~new_n3321_;
  assign n1400 = new_n3305_ | new_n3322_;
  assign new_n3324_ = \key<9>  & ~\encrypt<0> ;
  assign new_n3325_ = \key<1>  & \encrypt<0> ;
  assign new_n3326_ = ~new_n3324_ & ~new_n3325_;
  assign new_n3327_ = \start<0>  & ~new_n3326_;
  assign new_n3328_ = ~\C<14>  & ~\D<14> ;
  assign new_n3329_ = \C<14>  & \D<14> ;
  assign new_n3330_ = ~new_n3328_ & ~new_n3329_;
  assign new_n3331_ = ~new_n1185_1_ & ~new_n3330_;
  assign new_n3332_ = new_n1185_1_ & ~new_n3328_;
  assign new_n3333_ = ~new_n3331_ & ~new_n3332_;
  assign new_n3334_ = ~\encrypt<0>  & ~new_n3333_;
  assign new_n3335_ = \D<14>  & ~new_n1189_;
  assign new_n3336_ = ~\D<14>  & new_n1189_;
  assign new_n3337_ = ~new_n3335_ & ~new_n3336_;
  assign new_n3338_ = \C<14>  & ~new_n3337_;
  assign new_n3339_ = \D<14>  & new_n1189_;
  assign new_n3340_ = ~\C<14>  & new_n3339_;
  assign new_n3341_ = ~new_n3338_ & ~new_n3340_;
  assign new_n3342_ = \encrypt<0>  & ~new_n3341_;
  assign new_n3343_ = ~new_n3334_ & ~new_n3342_;
  assign new_n3344_ = ~\start<0>  & ~new_n3343_;
  assign n1405 = new_n3327_ | new_n3344_;
  assign new_n3346_ = \key<17>  & ~\encrypt<0> ;
  assign new_n3347_ = \key<9>  & \encrypt<0> ;
  assign new_n3348_ = ~new_n3346_ & ~new_n3347_;
  assign new_n3349_ = \start<0>  & ~new_n3348_;
  assign new_n3350_ = ~\C<13>  & ~\D<13> ;
  assign new_n3351_ = \C<13>  & \D<13> ;
  assign new_n3352_ = ~new_n3350_ & ~new_n3351_;
  assign new_n3353_ = ~new_n1185_1_ & ~new_n3352_;
  assign new_n3354_ = new_n1185_1_ & ~new_n3350_;
  assign new_n3355_ = ~new_n3353_ & ~new_n3354_;
  assign new_n3356_ = ~\encrypt<0>  & ~new_n3355_;
  assign new_n3357_ = \D<13>  & ~new_n1189_;
  assign new_n3358_ = ~\D<13>  & new_n1189_;
  assign new_n3359_ = ~new_n3357_ & ~new_n3358_;
  assign new_n3360_ = \C<13>  & ~new_n3359_;
  assign new_n3361_ = \D<13>  & new_n1189_;
  assign new_n3362_ = ~\C<13>  & new_n3361_;
  assign new_n3363_ = ~new_n3360_ & ~new_n3362_;
  assign new_n3364_ = \encrypt<0>  & ~new_n3363_;
  assign new_n3365_ = ~new_n3356_ & ~new_n3364_;
  assign new_n3366_ = ~\start<0>  & ~new_n3365_;
  assign n1410 = new_n3349_ | new_n3366_;
  assign new_n3368_ = \key<25>  & ~\encrypt<0> ;
  assign new_n3369_ = \key<17>  & \encrypt<0> ;
  assign new_n3370_ = ~new_n3368_ & ~new_n3369_;
  assign new_n3371_ = \start<0>  & ~new_n3370_;
  assign new_n3372_ = ~\C<12>  & ~\D<12> ;
  assign new_n3373_ = \C<12>  & \D<12> ;
  assign new_n3374_ = ~new_n3372_ & ~new_n3373_;
  assign new_n3375_ = ~new_n1185_1_ & ~new_n3374_;
  assign new_n3376_ = new_n1185_1_ & ~new_n3372_;
  assign new_n3377_ = ~new_n3375_ & ~new_n3376_;
  assign new_n3378_ = ~\encrypt<0>  & ~new_n3377_;
  assign new_n3379_ = \D<12>  & ~new_n1189_;
  assign new_n3380_ = ~\D<12>  & new_n1189_;
  assign new_n3381_ = ~new_n3379_ & ~new_n3380_;
  assign new_n3382_ = \C<12>  & ~new_n3381_;
  assign new_n3383_ = \D<12>  & new_n1189_;
  assign new_n3384_ = ~\C<12>  & new_n3383_;
  assign new_n3385_ = ~new_n3382_ & ~new_n3384_;
  assign new_n3386_ = \encrypt<0>  & ~new_n3385_;
  assign new_n3387_ = ~new_n3378_ & ~new_n3386_;
  assign new_n3388_ = ~\start<0>  & ~new_n3387_;
  assign n1415 = new_n3371_ | new_n3388_;
  assign new_n3390_ = \key<33>  & ~\encrypt<0> ;
  assign new_n3391_ = \key<25>  & \encrypt<0> ;
  assign new_n3392_ = ~new_n3390_ & ~new_n3391_;
  assign new_n3393_ = \start<0>  & ~new_n3392_;
  assign new_n3394_ = ~\C<11>  & ~\D<11> ;
  assign new_n3395_ = \C<11>  & \D<11> ;
  assign new_n3396_ = ~new_n3394_ & ~new_n3395_;
  assign new_n3397_ = ~new_n1185_1_ & ~new_n3396_;
  assign new_n3398_ = new_n1185_1_ & ~new_n3394_;
  assign new_n3399_ = ~new_n3397_ & ~new_n3398_;
  assign new_n3400_ = ~\encrypt<0>  & ~new_n3399_;
  assign new_n3401_ = \D<11>  & ~new_n1189_;
  assign new_n3402_ = ~\D<11>  & new_n1189_;
  assign new_n3403_ = ~new_n3401_ & ~new_n3402_;
  assign new_n3404_ = \C<11>  & ~new_n3403_;
  assign new_n3405_ = \D<11>  & new_n1189_;
  assign new_n3406_ = ~\C<11>  & new_n3405_;
  assign new_n3407_ = ~new_n3404_ & ~new_n3406_;
  assign new_n3408_ = \encrypt<0>  & ~new_n3407_;
  assign new_n3409_ = ~new_n3400_ & ~new_n3408_;
  assign new_n3410_ = ~\start<0>  & ~new_n3409_;
  assign n1420 = new_n3393_ | new_n3410_;
  assign new_n3412_ = \key<41>  & ~\encrypt<0> ;
  assign new_n3413_ = \key<33>  & \encrypt<0> ;
  assign new_n3414_ = ~new_n3412_ & ~new_n3413_;
  assign new_n3415_ = \start<0>  & ~new_n3414_;
  assign new_n3416_ = ~\C<10>  & ~\D<10> ;
  assign new_n3417_ = \C<10>  & \D<10> ;
  assign new_n3418_ = ~new_n3416_ & ~new_n3417_;
  assign new_n3419_ = ~new_n1185_1_ & ~new_n3418_;
  assign new_n3420_ = new_n1185_1_ & ~new_n3416_;
  assign new_n3421_ = ~new_n3419_ & ~new_n3420_;
  assign new_n3422_ = ~\encrypt<0>  & ~new_n3421_;
  assign new_n3423_ = \D<10>  & ~new_n1189_;
  assign new_n3424_ = ~\D<10>  & new_n1189_;
  assign new_n3425_ = ~new_n3423_ & ~new_n3424_;
  assign new_n3426_ = \C<10>  & ~new_n3425_;
  assign new_n3427_ = \D<10>  & new_n1189_;
  assign new_n3428_ = ~\C<10>  & new_n3427_;
  assign new_n3429_ = ~new_n3426_ & ~new_n3428_;
  assign new_n3430_ = \encrypt<0>  & ~new_n3429_;
  assign new_n3431_ = ~new_n3422_ & ~new_n3430_;
  assign new_n3432_ = ~\start<0>  & ~new_n3431_;
  assign n1425 = new_n3415_ | new_n3432_;
  assign new_n3434_ = \key<49>  & ~\encrypt<0> ;
  assign new_n3435_ = \key<41>  & \encrypt<0> ;
  assign new_n3436_ = ~new_n3434_ & ~new_n3435_;
  assign new_n3437_ = \start<0>  & ~new_n3436_;
  assign new_n3438_ = ~\C<9>  & ~\D<9> ;
  assign new_n3439_ = \C<9>  & \D<9> ;
  assign new_n3440_ = ~new_n3438_ & ~new_n3439_;
  assign new_n3441_ = ~new_n1185_1_ & ~new_n3440_;
  assign new_n3442_ = new_n1185_1_ & ~new_n3438_;
  assign new_n3443_ = ~new_n3441_ & ~new_n3442_;
  assign new_n3444_ = ~\encrypt<0>  & ~new_n3443_;
  assign new_n3445_ = \D<9>  & ~new_n1189_;
  assign new_n3446_ = ~\D<9>  & new_n1189_;
  assign new_n3447_ = ~new_n3445_ & ~new_n3446_;
  assign new_n3448_ = \C<9>  & ~new_n3447_;
  assign new_n3449_ = \D<9>  & new_n1189_;
  assign new_n3450_ = ~\C<9>  & new_n3449_;
  assign new_n3451_ = ~new_n3448_ & ~new_n3450_;
  assign new_n3452_ = \encrypt<0>  & ~new_n3451_;
  assign new_n3453_ = ~new_n3444_ & ~new_n3452_;
  assign new_n3454_ = ~\start<0>  & ~new_n3453_;
  assign n1430 = new_n3437_ | new_n3454_;
  assign new_n3456_ = \key<57>  & ~\encrypt<0> ;
  assign new_n3457_ = \key<49>  & \encrypt<0> ;
  assign new_n3458_ = ~new_n3456_ & ~new_n3457_;
  assign new_n3459_ = \start<0>  & ~new_n3458_;
  assign new_n3460_ = ~\C<8>  & ~\D<8> ;
  assign new_n3461_ = \C<8>  & \D<8> ;
  assign new_n3462_ = ~new_n3460_ & ~new_n3461_;
  assign new_n3463_ = ~new_n1185_1_ & ~new_n3462_;
  assign new_n3464_ = new_n1185_1_ & ~new_n3460_;
  assign new_n3465_ = ~new_n3463_ & ~new_n3464_;
  assign new_n3466_ = ~\encrypt<0>  & ~new_n3465_;
  assign new_n3467_ = \D<8>  & ~new_n1189_;
  assign new_n3468_ = ~\D<8>  & new_n1189_;
  assign new_n3469_ = ~new_n3467_ & ~new_n3468_;
  assign new_n3470_ = \C<8>  & ~new_n3469_;
  assign new_n3471_ = \D<8>  & new_n1189_;
  assign new_n3472_ = ~\C<8>  & new_n3471_;
  assign new_n3473_ = ~new_n3470_ & ~new_n3472_;
  assign new_n3474_ = \encrypt<0>  & ~new_n3473_;
  assign new_n3475_ = ~new_n3466_ & ~new_n3474_;
  assign new_n3476_ = ~\start<0>  & ~new_n3475_;
  assign n1435 = new_n3459_ | new_n3476_;
  assign new_n3478_ = \key<0>  & ~\encrypt<0> ;
  assign new_n3479_ = \key<57>  & \encrypt<0> ;
  assign new_n3480_ = ~new_n3478_ & ~new_n3479_;
  assign new_n3481_ = \start<0>  & ~new_n3480_;
  assign new_n3482_ = ~\C<7>  & ~\D<7> ;
  assign new_n3483_ = \C<7>  & \D<7> ;
  assign new_n3484_ = ~new_n3482_ & ~new_n3483_;
  assign new_n3485_ = ~new_n1185_1_ & ~new_n3484_;
  assign new_n3486_ = new_n1185_1_ & ~new_n3482_;
  assign new_n3487_ = ~new_n3485_ & ~new_n3486_;
  assign new_n3488_ = ~\encrypt<0>  & ~new_n3487_;
  assign new_n3489_ = \D<7>  & ~new_n1189_;
  assign new_n3490_ = ~\D<7>  & new_n1189_;
  assign new_n3491_ = ~new_n3489_ & ~new_n3490_;
  assign new_n3492_ = \C<7>  & ~new_n3491_;
  assign new_n3493_ = \D<7>  & new_n1189_;
  assign new_n3494_ = ~\C<7>  & new_n3493_;
  assign new_n3495_ = ~new_n3492_ & ~new_n3494_;
  assign new_n3496_ = \encrypt<0>  & ~new_n3495_;
  assign new_n3497_ = ~new_n3488_ & ~new_n3496_;
  assign new_n3498_ = ~\start<0>  & ~new_n3497_;
  assign n1440 = new_n3481_ | new_n3498_;
  assign new_n3500_ = \key<8>  & ~\encrypt<0> ;
  assign new_n3501_ = \key<0>  & \encrypt<0> ;
  assign new_n3502_ = ~new_n3500_ & ~new_n3501_;
  assign new_n3503_ = \start<0>  & ~new_n3502_;
  assign new_n3504_ = ~\C<6>  & ~\D<6> ;
  assign new_n3505_ = \C<6>  & \D<6> ;
  assign new_n3506_ = ~new_n3504_ & ~new_n3505_;
  assign new_n3507_ = ~new_n1185_1_ & ~new_n3506_;
  assign new_n3508_ = new_n1185_1_ & ~new_n3504_;
  assign new_n3509_ = ~new_n3507_ & ~new_n3508_;
  assign new_n3510_ = ~\encrypt<0>  & ~new_n3509_;
  assign new_n3511_ = \D<6>  & ~new_n1189_;
  assign new_n3512_ = ~\D<6>  & new_n1189_;
  assign new_n3513_ = ~new_n3511_ & ~new_n3512_;
  assign new_n3514_ = \C<6>  & ~new_n3513_;
  assign new_n3515_ = \D<6>  & new_n1189_;
  assign new_n3516_ = ~\C<6>  & new_n3515_;
  assign new_n3517_ = ~new_n3514_ & ~new_n3516_;
  assign new_n3518_ = \encrypt<0>  & ~new_n3517_;
  assign new_n3519_ = ~new_n3510_ & ~new_n3518_;
  assign new_n3520_ = ~\start<0>  & ~new_n3519_;
  assign n1445 = new_n3503_ | new_n3520_;
  assign new_n3522_ = \key<16>  & ~\encrypt<0> ;
  assign new_n3523_ = \key<8>  & \encrypt<0> ;
  assign new_n3524_ = ~new_n3522_ & ~new_n3523_;
  assign new_n3525_ = \start<0>  & ~new_n3524_;
  assign new_n3526_ = ~\C<5>  & ~\D<5> ;
  assign new_n3527_ = \C<5>  & \D<5> ;
  assign new_n3528_ = ~new_n3526_ & ~new_n3527_;
  assign new_n3529_ = ~new_n1185_1_ & ~new_n3528_;
  assign new_n3530_ = new_n1185_1_ & ~new_n3526_;
  assign new_n3531_ = ~new_n3529_ & ~new_n3530_;
  assign new_n3532_ = ~\encrypt<0>  & ~new_n3531_;
  assign new_n3533_ = \D<5>  & ~new_n1189_;
  assign new_n3534_ = ~\D<5>  & new_n1189_;
  assign new_n3535_ = ~new_n3533_ & ~new_n3534_;
  assign new_n3536_ = \C<5>  & ~new_n3535_;
  assign new_n3537_ = \D<5>  & new_n1189_;
  assign new_n3538_ = ~\C<5>  & new_n3537_;
  assign new_n3539_ = ~new_n3536_ & ~new_n3538_;
  assign new_n3540_ = \encrypt<0>  & ~new_n3539_;
  assign new_n3541_ = ~new_n3532_ & ~new_n3540_;
  assign new_n3542_ = ~\start<0>  & ~new_n3541_;
  assign n1450 = new_n3525_ | new_n3542_;
  assign new_n3544_ = \key<24>  & ~\encrypt<0> ;
  assign new_n3545_ = \key<16>  & \encrypt<0> ;
  assign new_n3546_ = ~new_n3544_ & ~new_n3545_;
  assign new_n3547_ = \start<0>  & ~new_n3546_;
  assign new_n3548_ = ~\C<4>  & ~\D<4> ;
  assign new_n3549_ = \C<4>  & \D<4> ;
  assign new_n3550_ = ~new_n3548_ & ~new_n3549_;
  assign new_n3551_ = ~new_n1185_1_ & ~new_n3550_;
  assign new_n3552_ = new_n1185_1_ & ~new_n3548_;
  assign new_n3553_ = ~new_n3551_ & ~new_n3552_;
  assign new_n3554_ = ~\encrypt<0>  & ~new_n3553_;
  assign new_n3555_ = \D<4>  & ~new_n1189_;
  assign new_n3556_ = ~\D<4>  & new_n1189_;
  assign new_n3557_ = ~new_n3555_ & ~new_n3556_;
  assign new_n3558_ = \C<4>  & ~new_n3557_;
  assign new_n3559_ = \D<4>  & new_n1189_;
  assign new_n3560_ = ~\C<4>  & new_n3559_;
  assign new_n3561_ = ~new_n3558_ & ~new_n3560_;
  assign new_n3562_ = \encrypt<0>  & ~new_n3561_;
  assign new_n3563_ = ~new_n3554_ & ~new_n3562_;
  assign new_n3564_ = ~\start<0>  & ~new_n3563_;
  assign n1455 = new_n3547_ | new_n3564_;
  assign new_n3566_ = \key<32>  & ~\encrypt<0> ;
  assign new_n3567_ = \key<24>  & \encrypt<0> ;
  assign new_n3568_ = ~new_n3566_ & ~new_n3567_;
  assign new_n3569_ = \start<0>  & ~new_n3568_;
  assign new_n3570_ = ~\C<3>  & ~\D<3> ;
  assign new_n3571_ = \C<3>  & \D<3> ;
  assign new_n3572_ = ~new_n3570_ & ~new_n3571_;
  assign new_n3573_ = ~new_n1185_1_ & ~new_n3572_;
  assign new_n3574_ = new_n1185_1_ & ~new_n3570_;
  assign new_n3575_ = ~new_n3573_ & ~new_n3574_;
  assign new_n3576_ = ~\encrypt<0>  & ~new_n3575_;
  assign new_n3577_ = \D<3>  & ~new_n1189_;
  assign new_n3578_ = ~\D<3>  & new_n1189_;
  assign new_n3579_ = ~new_n3577_ & ~new_n3578_;
  assign new_n3580_ = \C<3>  & ~new_n3579_;
  assign new_n3581_ = \D<3>  & new_n1189_;
  assign new_n3582_ = ~\C<3>  & new_n3581_;
  assign new_n3583_ = ~new_n3580_ & ~new_n3582_;
  assign new_n3584_ = \encrypt<0>  & ~new_n3583_;
  assign new_n3585_ = ~new_n3576_ & ~new_n3584_;
  assign new_n3586_ = ~\start<0>  & ~new_n3585_;
  assign n1460 = new_n3569_ | new_n3586_;
  assign new_n3588_ = \key<40>  & ~\encrypt<0> ;
  assign new_n3589_ = \key<32>  & \encrypt<0> ;
  assign new_n3590_ = ~new_n3588_ & ~new_n3589_;
  assign new_n3591_ = \start<0>  & ~new_n3590_;
  assign new_n3592_ = ~\C<2>  & ~\D<2> ;
  assign new_n3593_ = \C<2>  & \D<2> ;
  assign new_n3594_ = ~new_n3592_ & ~new_n3593_;
  assign new_n3595_ = ~new_n1185_1_ & ~new_n3594_;
  assign new_n3596_ = new_n1185_1_ & ~new_n3592_;
  assign new_n3597_ = ~new_n3595_ & ~new_n3596_;
  assign new_n3598_ = ~\encrypt<0>  & ~new_n3597_;
  assign new_n3599_ = \D<2>  & ~new_n1189_;
  assign new_n3600_ = ~\D<2>  & new_n1189_;
  assign new_n3601_ = ~new_n3599_ & ~new_n3600_;
  assign new_n3602_ = \C<2>  & ~new_n3601_;
  assign new_n3603_ = \D<2>  & new_n1189_;
  assign new_n3604_ = ~\C<2>  & new_n3603_;
  assign new_n3605_ = ~new_n3602_ & ~new_n3604_;
  assign new_n3606_ = \encrypt<0>  & ~new_n3605_;
  assign new_n3607_ = ~new_n3598_ & ~new_n3606_;
  assign new_n3608_ = ~\start<0>  & ~new_n3607_;
  assign n1465 = new_n3591_ | new_n3608_;
  assign new_n3610_ = \key<48>  & ~\encrypt<0> ;
  assign new_n3611_ = \key<40>  & \encrypt<0> ;
  assign new_n3612_ = ~new_n3610_ & ~new_n3611_;
  assign new_n3613_ = \start<0>  & ~new_n3612_;
  assign new_n3614_ = ~\C<1>  & ~\D<1> ;
  assign new_n3615_ = \C<1>  & \D<1> ;
  assign new_n3616_ = ~new_n3614_ & ~new_n3615_;
  assign new_n3617_ = ~new_n1185_1_ & ~new_n3616_;
  assign new_n3618_ = new_n1185_1_ & ~new_n3614_;
  assign new_n3619_ = ~new_n3617_ & ~new_n3618_;
  assign new_n3620_ = ~\encrypt<0>  & ~new_n3619_;
  assign new_n3621_ = \D<1>  & ~new_n1189_;
  assign new_n3622_ = ~\D<1>  & new_n1189_;
  assign new_n3623_ = ~new_n3621_ & ~new_n3622_;
  assign new_n3624_ = \C<1>  & ~new_n3623_;
  assign new_n3625_ = \D<1>  & new_n1189_;
  assign new_n3626_ = ~\C<1>  & new_n3625_;
  assign new_n3627_ = ~new_n3624_ & ~new_n3626_;
  assign new_n3628_ = \encrypt<0>  & ~new_n3627_;
  assign new_n3629_ = ~new_n3620_ & ~new_n3628_;
  assign new_n3630_ = ~\start<0>  & ~new_n3629_;
  assign n1470 = new_n3613_ | new_n3630_;
  assign new_n3632_ = \key<56>  & ~\encrypt<0> ;
  assign new_n3633_ = \key<48>  & \encrypt<0> ;
  assign new_n3634_ = ~new_n3632_ & ~new_n3633_;
  assign new_n3635_ = \start<0>  & ~new_n3634_;
  assign new_n3636_ = ~\C<0>  & ~\D<0> ;
  assign new_n3637_ = \C<0>  & \D<0> ;
  assign new_n3638_ = ~new_n3636_ & ~new_n3637_;
  assign new_n3639_ = ~new_n1185_1_ & ~new_n3638_;
  assign new_n3640_ = new_n1185_1_ & ~new_n3636_;
  assign new_n3641_ = ~new_n3639_ & ~new_n3640_;
  assign new_n3642_ = ~\encrypt<0>  & ~new_n3641_;
  assign new_n3643_ = \D<0>  & ~new_n1189_;
  assign new_n3644_ = ~\D<0>  & new_n1189_;
  assign new_n3645_ = ~new_n3643_ & ~new_n3644_;
  assign new_n3646_ = \C<0>  & ~new_n3645_;
  assign new_n3647_ = \D<0>  & new_n1189_;
  assign new_n3648_ = ~\C<0>  & new_n3647_;
  assign new_n3649_ = ~new_n3646_ & ~new_n3648_;
  assign new_n3650_ = \encrypt<0>  & ~new_n3649_;
  assign new_n3651_ = ~new_n3642_ & ~new_n3650_;
  assign new_n3652_ = ~\start<0>  & ~new_n3651_;
  assign n1475 = new_n3635_ | new_n3652_;
  assign new_n3654_ = \key<195>  & ~\encrypt<0> ;
  assign new_n3655_ = \key<62>  & \encrypt<0> ;
  assign new_n3656_ = ~new_n3654_ & ~new_n3655_;
  assign new_n3657_ = \start<0>  & ~new_n3656_;
  assign new_n3658_ = ~new_n1185_1_ & ~new_n1194_;
  assign new_n3659_ = new_n1185_1_ & ~new_n1196_;
  assign new_n3660_ = ~new_n3658_ & ~new_n3659_;
  assign new_n3661_ = ~\encrypt<0>  & ~new_n3660_;
  assign new_n3662_ = ~\C<111>  & ~new_n1189_;
  assign new_n3663_ = \C<111>  & new_n1189_;
  assign new_n3664_ = ~new_n3662_ & ~new_n3663_;
  assign new_n3665_ = \D<111>  & ~new_n3664_;
  assign new_n3666_ = \C<111>  & ~new_n1189_;
  assign new_n3667_ = ~\D<111>  & new_n3666_;
  assign new_n3668_ = ~new_n3665_ & ~new_n3667_;
  assign new_n3669_ = \encrypt<0>  & ~new_n3668_;
  assign new_n3670_ = ~new_n3661_ & ~new_n3669_;
  assign new_n3671_ = ~\start<0>  & ~new_n3670_;
  assign n1480 = new_n3657_ | new_n3671_;
  assign new_n3673_ = \key<203>  & ~\encrypt<0> ;
  assign new_n3674_ = \key<195>  & \encrypt<0> ;
  assign new_n3675_ = ~new_n3673_ & ~new_n3674_;
  assign new_n3676_ = \start<0>  & ~new_n3675_;
  assign new_n3677_ = ~new_n1185_1_ & ~new_n1216_;
  assign new_n3678_ = new_n1185_1_ & ~new_n1218_;
  assign new_n3679_ = ~new_n3677_ & ~new_n3678_;
  assign new_n3680_ = ~\encrypt<0>  & ~new_n3679_;
  assign new_n3681_ = ~\C<110>  & ~new_n1189_;
  assign new_n3682_ = \C<110>  & new_n1189_;
  assign new_n3683_ = ~new_n3681_ & ~new_n3682_;
  assign new_n3684_ = \D<110>  & ~new_n3683_;
  assign new_n3685_ = \C<110>  & ~new_n1189_;
  assign new_n3686_ = ~\D<110>  & new_n3685_;
  assign new_n3687_ = ~new_n3684_ & ~new_n3686_;
  assign new_n3688_ = \encrypt<0>  & ~new_n3687_;
  assign new_n3689_ = ~new_n3680_ & ~new_n3688_;
  assign new_n3690_ = ~\start<0>  & ~new_n3689_;
  assign n1485 = new_n3676_ | new_n3690_;
  assign new_n3692_ = \key<211>  & ~\encrypt<0> ;
  assign new_n3693_ = \key<203>  & \encrypt<0> ;
  assign new_n3694_ = ~new_n3692_ & ~new_n3693_;
  assign new_n3695_ = \start<0>  & ~new_n3694_;
  assign new_n3696_ = ~new_n1185_1_ & ~new_n1238_;
  assign new_n3697_ = new_n1185_1_ & ~new_n1240_1_;
  assign new_n3698_ = ~new_n3696_ & ~new_n3697_;
  assign new_n3699_ = ~\encrypt<0>  & ~new_n3698_;
  assign new_n3700_ = ~\C<109>  & ~new_n1189_;
  assign new_n3701_ = \C<109>  & new_n1189_;
  assign new_n3702_ = ~new_n3700_ & ~new_n3701_;
  assign new_n3703_ = \D<109>  & ~new_n3702_;
  assign new_n3704_ = \C<109>  & ~new_n1189_;
  assign new_n3705_ = ~\D<109>  & new_n3704_;
  assign new_n3706_ = ~new_n3703_ & ~new_n3705_;
  assign new_n3707_ = \encrypt<0>  & ~new_n3706_;
  assign new_n3708_ = ~new_n3699_ & ~new_n3707_;
  assign new_n3709_ = ~\start<0>  & ~new_n3708_;
  assign n1490 = new_n3695_ | new_n3709_;
  assign new_n3711_ = \key<219>  & ~\encrypt<0> ;
  assign new_n3712_ = \key<211>  & \encrypt<0> ;
  assign new_n3713_ = ~new_n3711_ & ~new_n3712_;
  assign new_n3714_ = \start<0>  & ~new_n3713_;
  assign new_n3715_ = ~new_n1185_1_ & ~new_n1260_1_;
  assign new_n3716_ = new_n1185_1_ & ~new_n1262_;
  assign new_n3717_ = ~new_n3715_ & ~new_n3716_;
  assign new_n3718_ = ~\encrypt<0>  & ~new_n3717_;
  assign new_n3719_ = ~\C<108>  & ~new_n1189_;
  assign new_n3720_ = \C<108>  & new_n1189_;
  assign new_n3721_ = ~new_n3719_ & ~new_n3720_;
  assign new_n3722_ = \D<108>  & ~new_n3721_;
  assign new_n3723_ = \C<108>  & ~new_n1189_;
  assign new_n3724_ = ~\D<108>  & new_n3723_;
  assign new_n3725_ = ~new_n3722_ & ~new_n3724_;
  assign new_n3726_ = \encrypt<0>  & ~new_n3725_;
  assign new_n3727_ = ~new_n3718_ & ~new_n3726_;
  assign new_n3728_ = ~\start<0>  & ~new_n3727_;
  assign n1495 = new_n3714_ | new_n3728_;
  assign new_n3730_ = \key<196>  & ~\encrypt<0> ;
  assign new_n3731_ = \key<219>  & \encrypt<0> ;
  assign new_n3732_ = ~new_n3730_ & ~new_n3731_;
  assign new_n3733_ = \start<0>  & ~new_n3732_;
  assign new_n3734_ = ~new_n1185_1_ & ~new_n1282_;
  assign new_n3735_ = new_n1185_1_ & ~new_n1284_;
  assign new_n3736_ = ~new_n3734_ & ~new_n3735_;
  assign new_n3737_ = ~\encrypt<0>  & ~new_n3736_;
  assign new_n3738_ = ~\C<107>  & ~new_n1189_;
  assign new_n3739_ = \C<107>  & new_n1189_;
  assign new_n3740_ = ~new_n3738_ & ~new_n3739_;
  assign new_n3741_ = \D<107>  & ~new_n3740_;
  assign new_n3742_ = \C<107>  & ~new_n1189_;
  assign new_n3743_ = ~\D<107>  & new_n3742_;
  assign new_n3744_ = ~new_n3741_ & ~new_n3743_;
  assign new_n3745_ = \encrypt<0>  & ~new_n3744_;
  assign new_n3746_ = ~new_n3737_ & ~new_n3745_;
  assign new_n3747_ = ~\start<0>  & ~new_n3746_;
  assign n1500 = new_n3733_ | new_n3747_;
  assign new_n3749_ = \key<204>  & ~\encrypt<0> ;
  assign new_n3750_ = \key<196>  & \encrypt<0> ;
  assign new_n3751_ = ~new_n3749_ & ~new_n3750_;
  assign new_n3752_ = \start<0>  & ~new_n3751_;
  assign new_n3753_ = ~new_n1185_1_ & ~new_n1304_;
  assign new_n3754_ = new_n1185_1_ & ~new_n1306_;
  assign new_n3755_ = ~new_n3753_ & ~new_n3754_;
  assign new_n3756_ = ~\encrypt<0>  & ~new_n3755_;
  assign new_n3757_ = ~\C<106>  & ~new_n1189_;
  assign new_n3758_ = \C<106>  & new_n1189_;
  assign new_n3759_ = ~new_n3757_ & ~new_n3758_;
  assign new_n3760_ = \D<106>  & ~new_n3759_;
  assign new_n3761_ = \C<106>  & ~new_n1189_;
  assign new_n3762_ = ~\D<106>  & new_n3761_;
  assign new_n3763_ = ~new_n3760_ & ~new_n3762_;
  assign new_n3764_ = \encrypt<0>  & ~new_n3763_;
  assign new_n3765_ = ~new_n3756_ & ~new_n3764_;
  assign new_n3766_ = ~\start<0>  & ~new_n3765_;
  assign n1505 = new_n3752_ | new_n3766_;
  assign new_n3768_ = \key<212>  & ~\encrypt<0> ;
  assign new_n3769_ = \key<204>  & \encrypt<0> ;
  assign new_n3770_ = ~new_n3768_ & ~new_n3769_;
  assign new_n3771_ = \start<0>  & ~new_n3770_;
  assign new_n3772_ = ~new_n1185_1_ & ~new_n1326_;
  assign new_n3773_ = new_n1185_1_ & ~new_n1328_;
  assign new_n3774_ = ~new_n3772_ & ~new_n3773_;
  assign new_n3775_ = ~\encrypt<0>  & ~new_n3774_;
  assign new_n3776_ = ~\C<105>  & ~new_n1189_;
  assign new_n3777_ = \C<105>  & new_n1189_;
  assign new_n3778_ = ~new_n3776_ & ~new_n3777_;
  assign new_n3779_ = \D<105>  & ~new_n3778_;
  assign new_n3780_ = \C<105>  & ~new_n1189_;
  assign new_n3781_ = ~\D<105>  & new_n3780_;
  assign new_n3782_ = ~new_n3779_ & ~new_n3781_;
  assign new_n3783_ = \encrypt<0>  & ~new_n3782_;
  assign new_n3784_ = ~new_n3775_ & ~new_n3783_;
  assign new_n3785_ = ~\start<0>  & ~new_n3784_;
  assign n1510 = new_n3771_ | new_n3785_;
  assign new_n3787_ = \key<220>  & ~\encrypt<0> ;
  assign new_n3788_ = \key<212>  & \encrypt<0> ;
  assign new_n3789_ = ~new_n3787_ & ~new_n3788_;
  assign new_n3790_ = \start<0>  & ~new_n3789_;
  assign new_n3791_ = ~new_n1185_1_ & ~new_n1348_;
  assign new_n3792_ = new_n1185_1_ & ~new_n1350_1_;
  assign new_n3793_ = ~new_n3791_ & ~new_n3792_;
  assign new_n3794_ = ~\encrypt<0>  & ~new_n3793_;
  assign new_n3795_ = ~\C<104>  & ~new_n1189_;
  assign new_n3796_ = \C<104>  & new_n1189_;
  assign new_n3797_ = ~new_n3795_ & ~new_n3796_;
  assign new_n3798_ = \D<104>  & ~new_n3797_;
  assign new_n3799_ = \C<104>  & ~new_n1189_;
  assign new_n3800_ = ~\D<104>  & new_n3799_;
  assign new_n3801_ = ~new_n3798_ & ~new_n3800_;
  assign new_n3802_ = \encrypt<0>  & ~new_n3801_;
  assign new_n3803_ = ~new_n3794_ & ~new_n3802_;
  assign new_n3804_ = ~\start<0>  & ~new_n3803_;
  assign n1515 = new_n3790_ | new_n3804_;
  assign new_n3806_ = \key<228>  & ~\encrypt<0> ;
  assign new_n3807_ = \key<220>  & \encrypt<0> ;
  assign new_n3808_ = ~new_n3806_ & ~new_n3807_;
  assign new_n3809_ = \start<0>  & ~new_n3808_;
  assign new_n3810_ = ~new_n1185_1_ & ~new_n1370_1_;
  assign new_n3811_ = new_n1185_1_ & ~new_n1372_;
  assign new_n3812_ = ~new_n3810_ & ~new_n3811_;
  assign new_n3813_ = ~\encrypt<0>  & ~new_n3812_;
  assign new_n3814_ = ~\C<103>  & ~new_n1189_;
  assign new_n3815_ = \C<103>  & new_n1189_;
  assign new_n3816_ = ~new_n3814_ & ~new_n3815_;
  assign new_n3817_ = \D<103>  & ~new_n3816_;
  assign new_n3818_ = \C<103>  & ~new_n1189_;
  assign new_n3819_ = ~\D<103>  & new_n3818_;
  assign new_n3820_ = ~new_n3817_ & ~new_n3819_;
  assign new_n3821_ = \encrypt<0>  & ~new_n3820_;
  assign new_n3822_ = ~new_n3813_ & ~new_n3821_;
  assign new_n3823_ = ~\start<0>  & ~new_n3822_;
  assign n1520 = new_n3809_ | new_n3823_;
  assign new_n3825_ = \key<172>  & ~\encrypt<0> ;
  assign new_n3826_ = \key<228>  & \encrypt<0> ;
  assign new_n3827_ = ~new_n3825_ & ~new_n3826_;
  assign new_n3828_ = \start<0>  & ~new_n3827_;
  assign new_n3829_ = ~new_n1185_1_ & ~new_n1392_;
  assign new_n3830_ = new_n1185_1_ & ~new_n1394_;
  assign new_n3831_ = ~new_n3829_ & ~new_n3830_;
  assign new_n3832_ = ~\encrypt<0>  & ~new_n3831_;
  assign new_n3833_ = ~\C<102>  & ~new_n1189_;
  assign new_n3834_ = \C<102>  & new_n1189_;
  assign new_n3835_ = ~new_n3833_ & ~new_n3834_;
  assign new_n3836_ = \D<102>  & ~new_n3835_;
  assign new_n3837_ = \C<102>  & ~new_n1189_;
  assign new_n3838_ = ~\D<102>  & new_n3837_;
  assign new_n3839_ = ~new_n3836_ & ~new_n3838_;
  assign new_n3840_ = \encrypt<0>  & ~new_n3839_;
  assign new_n3841_ = ~new_n3832_ & ~new_n3840_;
  assign new_n3842_ = ~\start<0>  & ~new_n3841_;
  assign n1525 = new_n3828_ | new_n3842_;
  assign new_n3844_ = \key<244>  & ~\encrypt<0> ;
  assign new_n3845_ = \key<172>  & \encrypt<0> ;
  assign new_n3846_ = ~new_n3844_ & ~new_n3845_;
  assign new_n3847_ = \start<0>  & ~new_n3846_;
  assign new_n3848_ = ~new_n1185_1_ & ~new_n1414_;
  assign new_n3849_ = new_n1185_1_ & ~new_n1416_;
  assign new_n3850_ = ~new_n3848_ & ~new_n3849_;
  assign new_n3851_ = ~\encrypt<0>  & ~new_n3850_;
  assign new_n3852_ = ~\C<101>  & ~new_n1189_;
  assign new_n3853_ = \C<101>  & new_n1189_;
  assign new_n3854_ = ~new_n3852_ & ~new_n3853_;
  assign new_n3855_ = \D<101>  & ~new_n3854_;
  assign new_n3856_ = \C<101>  & ~new_n1189_;
  assign new_n3857_ = ~\D<101>  & new_n3856_;
  assign new_n3858_ = ~new_n3855_ & ~new_n3857_;
  assign new_n3859_ = \encrypt<0>  & ~new_n3858_;
  assign new_n3860_ = ~new_n3851_ & ~new_n3859_;
  assign new_n3861_ = ~\start<0>  & ~new_n3860_;
  assign n1530 = new_n3847_ | new_n3861_;
  assign new_n3863_ = \key<252>  & ~\encrypt<0> ;
  assign new_n3864_ = \key<244>  & \encrypt<0> ;
  assign new_n3865_ = ~new_n3863_ & ~new_n3864_;
  assign new_n3866_ = \start<0>  & ~new_n3865_;
  assign new_n3867_ = ~new_n1185_1_ & ~new_n1436_;
  assign new_n3868_ = new_n1185_1_ & ~new_n1438_;
  assign new_n3869_ = ~new_n3867_ & ~new_n3868_;
  assign new_n3870_ = ~\encrypt<0>  & ~new_n3869_;
  assign new_n3871_ = ~\C<100>  & ~new_n1189_;
  assign new_n3872_ = \C<100>  & new_n1189_;
  assign new_n3873_ = ~new_n3871_ & ~new_n3872_;
  assign new_n3874_ = \D<100>  & ~new_n3873_;
  assign new_n3875_ = \C<100>  & ~new_n1189_;
  assign new_n3876_ = ~\D<100>  & new_n3875_;
  assign new_n3877_ = ~new_n3874_ & ~new_n3876_;
  assign new_n3878_ = \encrypt<0>  & ~new_n3877_;
  assign new_n3879_ = ~new_n3870_ & ~new_n3878_;
  assign new_n3880_ = ~\start<0>  & ~new_n3879_;
  assign n1535 = new_n3866_ | new_n3880_;
  assign new_n3882_ = \key<197>  & ~\encrypt<0> ;
  assign new_n3883_ = \key<252>  & \encrypt<0> ;
  assign new_n3884_ = ~new_n3882_ & ~new_n3883_;
  assign new_n3885_ = \start<0>  & ~new_n3884_;
  assign new_n3886_ = ~new_n1185_1_ & ~new_n1458_;
  assign new_n3887_ = new_n1185_1_ & ~new_n1460_1_;
  assign new_n3888_ = ~new_n3886_ & ~new_n3887_;
  assign new_n3889_ = ~\encrypt<0>  & ~new_n3888_;
  assign new_n3890_ = ~\C<99>  & ~new_n1189_;
  assign new_n3891_ = \C<99>  & new_n1189_;
  assign new_n3892_ = ~new_n3890_ & ~new_n3891_;
  assign new_n3893_ = \D<99>  & ~new_n3892_;
  assign new_n3894_ = \C<99>  & ~new_n1189_;
  assign new_n3895_ = ~\D<99>  & new_n3894_;
  assign new_n3896_ = ~new_n3893_ & ~new_n3895_;
  assign new_n3897_ = \encrypt<0>  & ~new_n3896_;
  assign new_n3898_ = ~new_n3889_ & ~new_n3897_;
  assign new_n3899_ = ~\start<0>  & ~new_n3898_;
  assign n1540 = new_n3885_ | new_n3899_;
  assign new_n3901_ = \key<205>  & ~\encrypt<0> ;
  assign new_n3902_ = \key<197>  & \encrypt<0> ;
  assign new_n3903_ = ~new_n3901_ & ~new_n3902_;
  assign new_n3904_ = \start<0>  & ~new_n3903_;
  assign new_n3905_ = ~new_n1185_1_ & ~new_n1480_1_;
  assign new_n3906_ = new_n1185_1_ & ~new_n1482_;
  assign new_n3907_ = ~new_n3905_ & ~new_n3906_;
  assign new_n3908_ = ~\encrypt<0>  & ~new_n3907_;
  assign new_n3909_ = ~\C<98>  & ~new_n1189_;
  assign new_n3910_ = \C<98>  & new_n1189_;
  assign new_n3911_ = ~new_n3909_ & ~new_n3910_;
  assign new_n3912_ = \D<98>  & ~new_n3911_;
  assign new_n3913_ = \C<98>  & ~new_n1189_;
  assign new_n3914_ = ~\D<98>  & new_n3913_;
  assign new_n3915_ = ~new_n3912_ & ~new_n3914_;
  assign new_n3916_ = \encrypt<0>  & ~new_n3915_;
  assign new_n3917_ = ~new_n3908_ & ~new_n3916_;
  assign new_n3918_ = ~\start<0>  & ~new_n3917_;
  assign n1545 = new_n3904_ | new_n3918_;
  assign new_n3920_ = \key<213>  & ~\encrypt<0> ;
  assign new_n3921_ = \key<205>  & \encrypt<0> ;
  assign new_n3922_ = ~new_n3920_ & ~new_n3921_;
  assign new_n3923_ = \start<0>  & ~new_n3922_;
  assign new_n3924_ = ~new_n1185_1_ & ~new_n1502_;
  assign new_n3925_ = new_n1185_1_ & ~new_n1504_;
  assign new_n3926_ = ~new_n3924_ & ~new_n3925_;
  assign new_n3927_ = ~\encrypt<0>  & ~new_n3926_;
  assign new_n3928_ = ~\C<97>  & ~new_n1189_;
  assign new_n3929_ = \C<97>  & new_n1189_;
  assign new_n3930_ = ~new_n3928_ & ~new_n3929_;
  assign new_n3931_ = \D<97>  & ~new_n3930_;
  assign new_n3932_ = \C<97>  & ~new_n1189_;
  assign new_n3933_ = ~\D<97>  & new_n3932_;
  assign new_n3934_ = ~new_n3931_ & ~new_n3933_;
  assign new_n3935_ = \encrypt<0>  & ~new_n3934_;
  assign new_n3936_ = ~new_n3927_ & ~new_n3935_;
  assign new_n3937_ = ~\start<0>  & ~new_n3936_;
  assign n1550 = new_n3923_ | new_n3937_;
  assign new_n3939_ = \key<221>  & ~\encrypt<0> ;
  assign new_n3940_ = \key<213>  & \encrypt<0> ;
  assign new_n3941_ = ~new_n3939_ & ~new_n3940_;
  assign new_n3942_ = \start<0>  & ~new_n3941_;
  assign new_n3943_ = ~new_n1185_1_ & ~new_n1524_;
  assign new_n3944_ = new_n1185_1_ & ~new_n1526_;
  assign new_n3945_ = ~new_n3943_ & ~new_n3944_;
  assign new_n3946_ = ~\encrypt<0>  & ~new_n3945_;
  assign new_n3947_ = ~\C<96>  & ~new_n1189_;
  assign new_n3948_ = \C<96>  & new_n1189_;
  assign new_n3949_ = ~new_n3947_ & ~new_n3948_;
  assign new_n3950_ = \D<96>  & ~new_n3949_;
  assign new_n3951_ = \C<96>  & ~new_n1189_;
  assign new_n3952_ = ~\D<96>  & new_n3951_;
  assign new_n3953_ = ~new_n3950_ & ~new_n3952_;
  assign new_n3954_ = \encrypt<0>  & ~new_n3953_;
  assign new_n3955_ = ~new_n3946_ & ~new_n3954_;
  assign new_n3956_ = ~\start<0>  & ~new_n3955_;
  assign n1555 = new_n3942_ | new_n3956_;
  assign new_n3958_ = \key<229>  & ~\encrypt<0> ;
  assign new_n3959_ = \key<221>  & \encrypt<0> ;
  assign new_n3960_ = ~new_n3958_ & ~new_n3959_;
  assign new_n3961_ = \start<0>  & ~new_n3960_;
  assign new_n3962_ = ~new_n1185_1_ & ~new_n1546_;
  assign new_n3963_ = new_n1185_1_ & ~new_n1548_;
  assign new_n3964_ = ~new_n3962_ & ~new_n3963_;
  assign new_n3965_ = ~\encrypt<0>  & ~new_n3964_;
  assign new_n3966_ = ~\C<95>  & ~new_n1189_;
  assign new_n3967_ = \C<95>  & new_n1189_;
  assign new_n3968_ = ~new_n3966_ & ~new_n3967_;
  assign new_n3969_ = \D<95>  & ~new_n3968_;
  assign new_n3970_ = \C<95>  & ~new_n1189_;
  assign new_n3971_ = ~\D<95>  & new_n3970_;
  assign new_n3972_ = ~new_n3969_ & ~new_n3971_;
  assign new_n3973_ = \encrypt<0>  & ~new_n3972_;
  assign new_n3974_ = ~new_n3965_ & ~new_n3973_;
  assign new_n3975_ = ~\start<0>  & ~new_n3974_;
  assign n1560 = new_n3961_ | new_n3975_;
  assign new_n3977_ = \key<237>  & ~\encrypt<0> ;
  assign new_n3978_ = \key<229>  & \encrypt<0> ;
  assign new_n3979_ = ~new_n3977_ & ~new_n3978_;
  assign new_n3980_ = \start<0>  & ~new_n3979_;
  assign new_n3981_ = ~new_n1185_1_ & ~new_n1568_;
  assign new_n3982_ = new_n1185_1_ & ~new_n1570_1_;
  assign new_n3983_ = ~new_n3981_ & ~new_n3982_;
  assign new_n3984_ = ~\encrypt<0>  & ~new_n3983_;
  assign new_n3985_ = ~\C<94>  & ~new_n1189_;
  assign new_n3986_ = \C<94>  & new_n1189_;
  assign new_n3987_ = ~new_n3985_ & ~new_n3986_;
  assign new_n3988_ = \D<94>  & ~new_n3987_;
  assign new_n3989_ = \C<94>  & ~new_n1189_;
  assign new_n3990_ = ~\D<94>  & new_n3989_;
  assign new_n3991_ = ~new_n3988_ & ~new_n3990_;
  assign new_n3992_ = \encrypt<0>  & ~new_n3991_;
  assign new_n3993_ = ~new_n3984_ & ~new_n3992_;
  assign new_n3994_ = ~\start<0>  & ~new_n3993_;
  assign n1565 = new_n3980_ | new_n3994_;
  assign new_n3996_ = \key<245>  & ~\encrypt<0> ;
  assign new_n3997_ = \key<237>  & \encrypt<0> ;
  assign new_n3998_ = ~new_n3996_ & ~new_n3997_;
  assign new_n3999_ = \start<0>  & ~new_n3998_;
  assign new_n4000_ = ~new_n1185_1_ & ~new_n1590_1_;
  assign new_n4001_ = new_n1185_1_ & ~new_n1592_;
  assign new_n4002_ = ~new_n4000_ & ~new_n4001_;
  assign new_n4003_ = ~\encrypt<0>  & ~new_n4002_;
  assign new_n4004_ = ~\C<93>  & ~new_n1189_;
  assign new_n4005_ = \C<93>  & new_n1189_;
  assign new_n4006_ = ~new_n4004_ & ~new_n4005_;
  assign new_n4007_ = \D<93>  & ~new_n4006_;
  assign new_n4008_ = \C<93>  & ~new_n1189_;
  assign new_n4009_ = ~\D<93>  & new_n4008_;
  assign new_n4010_ = ~new_n4007_ & ~new_n4009_;
  assign new_n4011_ = \encrypt<0>  & ~new_n4010_;
  assign new_n4012_ = ~new_n4003_ & ~new_n4011_;
  assign new_n4013_ = ~\start<0>  & ~new_n4012_;
  assign n1570 = new_n3999_ | new_n4013_;
  assign new_n4015_ = \key<253>  & ~\encrypt<0> ;
  assign new_n4016_ = \key<245>  & \encrypt<0> ;
  assign new_n4017_ = ~new_n4015_ & ~new_n4016_;
  assign new_n4018_ = \start<0>  & ~new_n4017_;
  assign new_n4019_ = ~new_n1185_1_ & ~new_n1612_;
  assign new_n4020_ = new_n1185_1_ & ~new_n1614_;
  assign new_n4021_ = ~new_n4019_ & ~new_n4020_;
  assign new_n4022_ = ~\encrypt<0>  & ~new_n4021_;
  assign new_n4023_ = ~\C<92>  & ~new_n1189_;
  assign new_n4024_ = \C<92>  & new_n1189_;
  assign new_n4025_ = ~new_n4023_ & ~new_n4024_;
  assign new_n4026_ = \D<92>  & ~new_n4025_;
  assign new_n4027_ = \C<92>  & ~new_n1189_;
  assign new_n4028_ = ~\D<92>  & new_n4027_;
  assign new_n4029_ = ~new_n4026_ & ~new_n4028_;
  assign new_n4030_ = \encrypt<0>  & ~new_n4029_;
  assign new_n4031_ = ~new_n4022_ & ~new_n4030_;
  assign new_n4032_ = ~\start<0>  & ~new_n4031_;
  assign n1575 = new_n4018_ | new_n4032_;
  assign new_n4034_ = \key<198>  & ~\encrypt<0> ;
  assign new_n4035_ = \key<253>  & \encrypt<0> ;
  assign new_n4036_ = ~new_n4034_ & ~new_n4035_;
  assign new_n4037_ = \start<0>  & ~new_n4036_;
  assign new_n4038_ = ~new_n1185_1_ & ~new_n1634_;
  assign new_n4039_ = new_n1185_1_ & ~new_n1636_;
  assign new_n4040_ = ~new_n4038_ & ~new_n4039_;
  assign new_n4041_ = ~\encrypt<0>  & ~new_n4040_;
  assign new_n4042_ = ~\C<91>  & ~new_n1189_;
  assign new_n4043_ = \C<91>  & new_n1189_;
  assign new_n4044_ = ~new_n4042_ & ~new_n4043_;
  assign new_n4045_ = \D<91>  & ~new_n4044_;
  assign new_n4046_ = \C<91>  & ~new_n1189_;
  assign new_n4047_ = ~\D<91>  & new_n4046_;
  assign new_n4048_ = ~new_n4045_ & ~new_n4047_;
  assign new_n4049_ = \encrypt<0>  & ~new_n4048_;
  assign new_n4050_ = ~new_n4041_ & ~new_n4049_;
  assign new_n4051_ = ~\start<0>  & ~new_n4050_;
  assign n1580 = new_n4037_ | new_n4051_;
  assign new_n4053_ = \key<206>  & ~\encrypt<0> ;
  assign new_n4054_ = \key<198>  & \encrypt<0> ;
  assign new_n4055_ = ~new_n4053_ & ~new_n4054_;
  assign new_n4056_ = \start<0>  & ~new_n4055_;
  assign new_n4057_ = ~new_n1185_1_ & ~new_n1656_;
  assign new_n4058_ = new_n1185_1_ & ~new_n1658_;
  assign new_n4059_ = ~new_n4057_ & ~new_n4058_;
  assign new_n4060_ = ~\encrypt<0>  & ~new_n4059_;
  assign new_n4061_ = ~\C<90>  & ~new_n1189_;
  assign new_n4062_ = \C<90>  & new_n1189_;
  assign new_n4063_ = ~new_n4061_ & ~new_n4062_;
  assign new_n4064_ = \D<90>  & ~new_n4063_;
  assign new_n4065_ = \C<90>  & ~new_n1189_;
  assign new_n4066_ = ~\D<90>  & new_n4065_;
  assign new_n4067_ = ~new_n4064_ & ~new_n4066_;
  assign new_n4068_ = \encrypt<0>  & ~new_n4067_;
  assign new_n4069_ = ~new_n4060_ & ~new_n4068_;
  assign new_n4070_ = ~\start<0>  & ~new_n4069_;
  assign n1585 = new_n4056_ | new_n4070_;
  assign new_n4072_ = \key<214>  & ~\encrypt<0> ;
  assign new_n4073_ = \key<206>  & \encrypt<0> ;
  assign new_n4074_ = ~new_n4072_ & ~new_n4073_;
  assign new_n4075_ = \start<0>  & ~new_n4074_;
  assign new_n4076_ = ~new_n1185_1_ & ~new_n1678_;
  assign new_n4077_ = new_n1185_1_ & ~new_n1680_1_;
  assign new_n4078_ = ~new_n4076_ & ~new_n4077_;
  assign new_n4079_ = ~\encrypt<0>  & ~new_n4078_;
  assign new_n4080_ = ~\C<89>  & ~new_n1189_;
  assign new_n4081_ = \C<89>  & new_n1189_;
  assign new_n4082_ = ~new_n4080_ & ~new_n4081_;
  assign new_n4083_ = \D<89>  & ~new_n4082_;
  assign new_n4084_ = \C<89>  & ~new_n1189_;
  assign new_n4085_ = ~\D<89>  & new_n4084_;
  assign new_n4086_ = ~new_n4083_ & ~new_n4085_;
  assign new_n4087_ = \encrypt<0>  & ~new_n4086_;
  assign new_n4088_ = ~new_n4079_ & ~new_n4087_;
  assign new_n4089_ = ~\start<0>  & ~new_n4088_;
  assign n1590 = new_n4075_ | new_n4089_;
  assign new_n4091_ = \key<222>  & ~\encrypt<0> ;
  assign new_n4092_ = \key<214>  & \encrypt<0> ;
  assign new_n4093_ = ~new_n4091_ & ~new_n4092_;
  assign new_n4094_ = \start<0>  & ~new_n4093_;
  assign new_n4095_ = ~new_n1185_1_ & ~new_n1700_1_;
  assign new_n4096_ = new_n1185_1_ & ~new_n1702_;
  assign new_n4097_ = ~new_n4095_ & ~new_n4096_;
  assign new_n4098_ = ~\encrypt<0>  & ~new_n4097_;
  assign new_n4099_ = ~\C<88>  & ~new_n1189_;
  assign new_n4100_ = \C<88>  & new_n1189_;
  assign new_n4101_ = ~new_n4099_ & ~new_n4100_;
  assign new_n4102_ = \D<88>  & ~new_n4101_;
  assign new_n4103_ = \C<88>  & ~new_n1189_;
  assign new_n4104_ = ~\D<88>  & new_n4103_;
  assign new_n4105_ = ~new_n4102_ & ~new_n4104_;
  assign new_n4106_ = \encrypt<0>  & ~new_n4105_;
  assign new_n4107_ = ~new_n4098_ & ~new_n4106_;
  assign new_n4108_ = ~\start<0>  & ~new_n4107_;
  assign n1595 = new_n4094_ | new_n4108_;
  assign new_n4110_ = \key<230>  & ~\encrypt<0> ;
  assign new_n4111_ = \key<222>  & \encrypt<0> ;
  assign new_n4112_ = ~new_n4110_ & ~new_n4111_;
  assign new_n4113_ = \start<0>  & ~new_n4112_;
  assign new_n4114_ = ~new_n1185_1_ & ~new_n1722_;
  assign new_n4115_ = new_n1185_1_ & ~new_n1724_;
  assign new_n4116_ = ~new_n4114_ & ~new_n4115_;
  assign new_n4117_ = ~\encrypt<0>  & ~new_n4116_;
  assign new_n4118_ = ~\C<87>  & ~new_n1189_;
  assign new_n4119_ = \C<87>  & new_n1189_;
  assign new_n4120_ = ~new_n4118_ & ~new_n4119_;
  assign new_n4121_ = \D<87>  & ~new_n4120_;
  assign new_n4122_ = \C<87>  & ~new_n1189_;
  assign new_n4123_ = ~\D<87>  & new_n4122_;
  assign new_n4124_ = ~new_n4121_ & ~new_n4123_;
  assign new_n4125_ = \encrypt<0>  & ~new_n4124_;
  assign new_n4126_ = ~new_n4117_ & ~new_n4125_;
  assign new_n4127_ = ~\start<0>  & ~new_n4126_;
  assign n1600 = new_n4113_ | new_n4127_;
  assign new_n4129_ = \key<238>  & ~\encrypt<0> ;
  assign new_n4130_ = \key<230>  & \encrypt<0> ;
  assign new_n4131_ = ~new_n4129_ & ~new_n4130_;
  assign new_n4132_ = \start<0>  & ~new_n4131_;
  assign new_n4133_ = ~new_n1185_1_ & ~new_n1744_;
  assign new_n4134_ = new_n1185_1_ & ~new_n1746_;
  assign new_n4135_ = ~new_n4133_ & ~new_n4134_;
  assign new_n4136_ = ~\encrypt<0>  & ~new_n4135_;
  assign new_n4137_ = ~\C<86>  & ~new_n1189_;
  assign new_n4138_ = \C<86>  & new_n1189_;
  assign new_n4139_ = ~new_n4137_ & ~new_n4138_;
  assign new_n4140_ = \D<86>  & ~new_n4139_;
  assign new_n4141_ = \C<86>  & ~new_n1189_;
  assign new_n4142_ = ~\D<86>  & new_n4141_;
  assign new_n4143_ = ~new_n4140_ & ~new_n4142_;
  assign new_n4144_ = \encrypt<0>  & ~new_n4143_;
  assign new_n4145_ = ~new_n4136_ & ~new_n4144_;
  assign new_n4146_ = ~\start<0>  & ~new_n4145_;
  assign n1605 = new_n4132_ | new_n4146_;
  assign new_n4148_ = \key<246>  & ~\encrypt<0> ;
  assign new_n4149_ = \key<238>  & \encrypt<0> ;
  assign new_n4150_ = ~new_n4148_ & ~new_n4149_;
  assign new_n4151_ = \start<0>  & ~new_n4150_;
  assign new_n4152_ = ~new_n1185_1_ & ~new_n1766_;
  assign new_n4153_ = new_n1185_1_ & ~new_n1768_;
  assign new_n4154_ = ~new_n4152_ & ~new_n4153_;
  assign new_n4155_ = ~\encrypt<0>  & ~new_n4154_;
  assign new_n4156_ = ~\C<85>  & ~new_n1189_;
  assign new_n4157_ = \C<85>  & new_n1189_;
  assign new_n4158_ = ~new_n4156_ & ~new_n4157_;
  assign new_n4159_ = \D<85>  & ~new_n4158_;
  assign new_n4160_ = \C<85>  & ~new_n1189_;
  assign new_n4161_ = ~\D<85>  & new_n4160_;
  assign new_n4162_ = ~new_n4159_ & ~new_n4161_;
  assign new_n4163_ = \encrypt<0>  & ~new_n4162_;
  assign new_n4164_ = ~new_n4155_ & ~new_n4163_;
  assign new_n4165_ = ~\start<0>  & ~new_n4164_;
  assign n1610 = new_n4151_ | new_n4165_;
  assign new_n4167_ = \key<254>  & ~\encrypt<0> ;
  assign new_n4168_ = \key<246>  & \encrypt<0> ;
  assign new_n4169_ = ~new_n4167_ & ~new_n4168_;
  assign new_n4170_ = \start<0>  & ~new_n4169_;
  assign new_n4171_ = ~new_n1185_1_ & ~new_n1788_;
  assign new_n4172_ = new_n1185_1_ & ~new_n1790_1_;
  assign new_n4173_ = ~new_n4171_ & ~new_n4172_;
  assign new_n4174_ = ~\encrypt<0>  & ~new_n4173_;
  assign new_n4175_ = ~\C<84>  & ~new_n1189_;
  assign new_n4176_ = \C<84>  & new_n1189_;
  assign new_n4177_ = ~new_n4175_ & ~new_n4176_;
  assign new_n4178_ = \D<84>  & ~new_n4177_;
  assign new_n4179_ = \C<84>  & ~new_n1189_;
  assign new_n4180_ = ~\D<84>  & new_n4179_;
  assign new_n4181_ = ~new_n4178_ & ~new_n4180_;
  assign new_n4182_ = \encrypt<0>  & ~new_n4181_;
  assign new_n4183_ = ~new_n4174_ & ~new_n4182_;
  assign new_n4184_ = ~\start<0>  & ~new_n4183_;
  assign n1615 = new_n4170_ | new_n4184_;
  assign new_n4186_ = \key<131>  & ~\encrypt<0> ;
  assign new_n4187_ = \key<254>  & \encrypt<0> ;
  assign new_n4188_ = ~new_n4186_ & ~new_n4187_;
  assign new_n4189_ = \start<0>  & ~new_n4188_;
  assign new_n4190_ = ~new_n1185_1_ & ~new_n1810_1_;
  assign new_n4191_ = new_n1185_1_ & ~new_n1812_;
  assign new_n4192_ = ~new_n4190_ & ~new_n4191_;
  assign new_n4193_ = ~\encrypt<0>  & ~new_n4192_;
  assign new_n4194_ = ~\C<83>  & ~new_n1189_;
  assign new_n4195_ = \C<83>  & new_n1189_;
  assign new_n4196_ = ~new_n4194_ & ~new_n4195_;
  assign new_n4197_ = \D<83>  & ~new_n4196_;
  assign new_n4198_ = \C<83>  & ~new_n1189_;
  assign new_n4199_ = ~\D<83>  & new_n4198_;
  assign new_n4200_ = ~new_n4197_ & ~new_n4199_;
  assign new_n4201_ = \encrypt<0>  & ~new_n4200_;
  assign new_n4202_ = ~new_n4193_ & ~new_n4201_;
  assign new_n4203_ = ~\start<0>  & ~new_n4202_;
  assign n1620 = new_n4189_ | new_n4203_;
  assign new_n4205_ = \key<139>  & ~\encrypt<0> ;
  assign new_n4206_ = \key<131>  & \encrypt<0> ;
  assign new_n4207_ = ~new_n4205_ & ~new_n4206_;
  assign new_n4208_ = \start<0>  & ~new_n4207_;
  assign new_n4209_ = ~new_n1185_1_ & ~new_n1832_;
  assign new_n4210_ = new_n1185_1_ & ~new_n1834_;
  assign new_n4211_ = ~new_n4209_ & ~new_n4210_;
  assign new_n4212_ = ~\encrypt<0>  & ~new_n4211_;
  assign new_n4213_ = ~\C<82>  & ~new_n1189_;
  assign new_n4214_ = \C<82>  & new_n1189_;
  assign new_n4215_ = ~new_n4213_ & ~new_n4214_;
  assign new_n4216_ = \D<82>  & ~new_n4215_;
  assign new_n4217_ = \C<82>  & ~new_n1189_;
  assign new_n4218_ = ~\D<82>  & new_n4217_;
  assign new_n4219_ = ~new_n4216_ & ~new_n4218_;
  assign new_n4220_ = \encrypt<0>  & ~new_n4219_;
  assign new_n4221_ = ~new_n4212_ & ~new_n4220_;
  assign new_n4222_ = ~\start<0>  & ~new_n4221_;
  assign n1625 = new_n4208_ | new_n4222_;
  assign new_n4224_ = \key<147>  & ~\encrypt<0> ;
  assign new_n4225_ = \key<139>  & \encrypt<0> ;
  assign new_n4226_ = ~new_n4224_ & ~new_n4225_;
  assign new_n4227_ = \start<0>  & ~new_n4226_;
  assign new_n4228_ = ~new_n1185_1_ & ~new_n1854_;
  assign new_n4229_ = new_n1185_1_ & ~new_n1856_;
  assign new_n4230_ = ~new_n4228_ & ~new_n4229_;
  assign new_n4231_ = ~\encrypt<0>  & ~new_n4230_;
  assign new_n4232_ = ~\C<81>  & ~new_n1189_;
  assign new_n4233_ = \C<81>  & new_n1189_;
  assign new_n4234_ = ~new_n4232_ & ~new_n4233_;
  assign new_n4235_ = \D<81>  & ~new_n4234_;
  assign new_n4236_ = \C<81>  & ~new_n1189_;
  assign new_n4237_ = ~\D<81>  & new_n4236_;
  assign new_n4238_ = ~new_n4235_ & ~new_n4237_;
  assign new_n4239_ = \encrypt<0>  & ~new_n4238_;
  assign new_n4240_ = ~new_n4231_ & ~new_n4239_;
  assign new_n4241_ = ~\start<0>  & ~new_n4240_;
  assign n1630 = new_n4227_ | new_n4241_;
  assign new_n4243_ = \key<155>  & ~\encrypt<0> ;
  assign new_n4244_ = \key<147>  & \encrypt<0> ;
  assign new_n4245_ = ~new_n4243_ & ~new_n4244_;
  assign new_n4246_ = \start<0>  & ~new_n4245_;
  assign new_n4247_ = ~new_n1185_1_ & ~new_n1876_;
  assign new_n4248_ = new_n1185_1_ & ~new_n1878_;
  assign new_n4249_ = ~new_n4247_ & ~new_n4248_;
  assign new_n4250_ = ~\encrypt<0>  & ~new_n4249_;
  assign new_n4251_ = ~\C<80>  & ~new_n1189_;
  assign new_n4252_ = \C<80>  & new_n1189_;
  assign new_n4253_ = ~new_n4251_ & ~new_n4252_;
  assign new_n4254_ = \D<80>  & ~new_n4253_;
  assign new_n4255_ = \C<80>  & ~new_n1189_;
  assign new_n4256_ = ~\D<80>  & new_n4255_;
  assign new_n4257_ = ~new_n4254_ & ~new_n4256_;
  assign new_n4258_ = \encrypt<0>  & ~new_n4257_;
  assign new_n4259_ = ~new_n4250_ & ~new_n4258_;
  assign new_n4260_ = ~\start<0>  & ~new_n4259_;
  assign n1635 = new_n4246_ | new_n4260_;
  assign new_n4262_ = \key<132>  & ~\encrypt<0> ;
  assign new_n4263_ = \key<155>  & \encrypt<0> ;
  assign new_n4264_ = ~new_n4262_ & ~new_n4263_;
  assign new_n4265_ = \start<0>  & ~new_n4264_;
  assign new_n4266_ = ~new_n1185_1_ & ~new_n1898_;
  assign new_n4267_ = new_n1185_1_ & ~new_n1900_1_;
  assign new_n4268_ = ~new_n4266_ & ~new_n4267_;
  assign new_n4269_ = ~\encrypt<0>  & ~new_n4268_;
  assign new_n4270_ = ~\C<79>  & ~new_n1189_;
  assign new_n4271_ = \C<79>  & new_n1189_;
  assign new_n4272_ = ~new_n4270_ & ~new_n4271_;
  assign new_n4273_ = \D<79>  & ~new_n4272_;
  assign new_n4274_ = \C<79>  & ~new_n1189_;
  assign new_n4275_ = ~\D<79>  & new_n4274_;
  assign new_n4276_ = ~new_n4273_ & ~new_n4275_;
  assign new_n4277_ = \encrypt<0>  & ~new_n4276_;
  assign new_n4278_ = ~new_n4269_ & ~new_n4277_;
  assign new_n4279_ = ~\start<0>  & ~new_n4278_;
  assign n1640 = new_n4265_ | new_n4279_;
  assign new_n4281_ = \key<140>  & ~\encrypt<0> ;
  assign new_n4282_ = \key<132>  & \encrypt<0> ;
  assign new_n4283_ = ~new_n4281_ & ~new_n4282_;
  assign new_n4284_ = \start<0>  & ~new_n4283_;
  assign new_n4285_ = ~new_n1185_1_ & ~new_n1920_1_;
  assign new_n4286_ = new_n1185_1_ & ~new_n1922_;
  assign new_n4287_ = ~new_n4285_ & ~new_n4286_;
  assign new_n4288_ = ~\encrypt<0>  & ~new_n4287_;
  assign new_n4289_ = ~\C<78>  & ~new_n1189_;
  assign new_n4290_ = \C<78>  & new_n1189_;
  assign new_n4291_ = ~new_n4289_ & ~new_n4290_;
  assign new_n4292_ = \D<78>  & ~new_n4291_;
  assign new_n4293_ = \C<78>  & ~new_n1189_;
  assign new_n4294_ = ~\D<78>  & new_n4293_;
  assign new_n4295_ = ~new_n4292_ & ~new_n4294_;
  assign new_n4296_ = \encrypt<0>  & ~new_n4295_;
  assign new_n4297_ = ~new_n4288_ & ~new_n4296_;
  assign new_n4298_ = ~\start<0>  & ~new_n4297_;
  assign n1645 = new_n4284_ | new_n4298_;
  assign new_n4300_ = \key<148>  & ~\encrypt<0> ;
  assign new_n4301_ = \key<140>  & \encrypt<0> ;
  assign new_n4302_ = ~new_n4300_ & ~new_n4301_;
  assign new_n4303_ = \start<0>  & ~new_n4302_;
  assign new_n4304_ = ~new_n1185_1_ & ~new_n1942_;
  assign new_n4305_ = new_n1185_1_ & ~new_n1944_;
  assign new_n4306_ = ~new_n4304_ & ~new_n4305_;
  assign new_n4307_ = ~\encrypt<0>  & ~new_n4306_;
  assign new_n4308_ = ~\C<77>  & ~new_n1189_;
  assign new_n4309_ = \C<77>  & new_n1189_;
  assign new_n4310_ = ~new_n4308_ & ~new_n4309_;
  assign new_n4311_ = \D<77>  & ~new_n4310_;
  assign new_n4312_ = \C<77>  & ~new_n1189_;
  assign new_n4313_ = ~\D<77>  & new_n4312_;
  assign new_n4314_ = ~new_n4311_ & ~new_n4313_;
  assign new_n4315_ = \encrypt<0>  & ~new_n4314_;
  assign new_n4316_ = ~new_n4307_ & ~new_n4315_;
  assign new_n4317_ = ~\start<0>  & ~new_n4316_;
  assign n1650 = new_n4303_ | new_n4317_;
  assign new_n4319_ = \key<156>  & ~\encrypt<0> ;
  assign new_n4320_ = \key<148>  & \encrypt<0> ;
  assign new_n4321_ = ~new_n4319_ & ~new_n4320_;
  assign new_n4322_ = \start<0>  & ~new_n4321_;
  assign new_n4323_ = ~new_n1185_1_ & ~new_n1964_;
  assign new_n4324_ = new_n1185_1_ & ~new_n1966_;
  assign new_n4325_ = ~new_n4323_ & ~new_n4324_;
  assign new_n4326_ = ~\encrypt<0>  & ~new_n4325_;
  assign new_n4327_ = ~\C<76>  & ~new_n1189_;
  assign new_n4328_ = \C<76>  & new_n1189_;
  assign new_n4329_ = ~new_n4327_ & ~new_n4328_;
  assign new_n4330_ = \D<76>  & ~new_n4329_;
  assign new_n4331_ = \C<76>  & ~new_n1189_;
  assign new_n4332_ = ~\D<76>  & new_n4331_;
  assign new_n4333_ = ~new_n4330_ & ~new_n4332_;
  assign new_n4334_ = \encrypt<0>  & ~new_n4333_;
  assign new_n4335_ = ~new_n4326_ & ~new_n4334_;
  assign new_n4336_ = ~\start<0>  & ~new_n4335_;
  assign n1655 = new_n4322_ | new_n4336_;
  assign new_n4338_ = \key<164>  & ~\encrypt<0> ;
  assign new_n4339_ = \key<156>  & \encrypt<0> ;
  assign new_n4340_ = ~new_n4338_ & ~new_n4339_;
  assign new_n4341_ = \start<0>  & ~new_n4340_;
  assign new_n4342_ = ~new_n1185_1_ & ~new_n1986_;
  assign new_n4343_ = new_n1185_1_ & ~new_n1988_;
  assign new_n4344_ = ~new_n4342_ & ~new_n4343_;
  assign new_n4345_ = ~\encrypt<0>  & ~new_n4344_;
  assign new_n4346_ = ~\C<75>  & ~new_n1189_;
  assign new_n4347_ = \C<75>  & new_n1189_;
  assign new_n4348_ = ~new_n4346_ & ~new_n4347_;
  assign new_n4349_ = \D<75>  & ~new_n4348_;
  assign new_n4350_ = \C<75>  & ~new_n1189_;
  assign new_n4351_ = ~\D<75>  & new_n4350_;
  assign new_n4352_ = ~new_n4349_ & ~new_n4351_;
  assign new_n4353_ = \encrypt<0>  & ~new_n4352_;
  assign new_n4354_ = ~new_n4345_ & ~new_n4353_;
  assign new_n4355_ = ~\start<0>  & ~new_n4354_;
  assign n1660 = new_n4341_ | new_n4355_;
  assign new_n4357_ = \key<164>  & \encrypt<0> ;
  assign new_n4358_ = ~new_n3825_ & ~new_n4357_;
  assign new_n4359_ = \start<0>  & ~new_n4358_;
  assign new_n4360_ = ~new_n1185_1_ & ~new_n2008_;
  assign new_n4361_ = new_n1185_1_ & ~new_n2010_1_;
  assign new_n4362_ = ~new_n4360_ & ~new_n4361_;
  assign new_n4363_ = ~\encrypt<0>  & ~new_n4362_;
  assign new_n4364_ = ~\C<74>  & ~new_n1189_;
  assign new_n4365_ = \C<74>  & new_n1189_;
  assign new_n4366_ = ~new_n4364_ & ~new_n4365_;
  assign new_n4367_ = \D<74>  & ~new_n4366_;
  assign new_n4368_ = \C<74>  & ~new_n1189_;
  assign new_n4369_ = ~\D<74>  & new_n4368_;
  assign new_n4370_ = ~new_n4367_ & ~new_n4369_;
  assign new_n4371_ = \encrypt<0>  & ~new_n4370_;
  assign new_n4372_ = ~new_n4363_ & ~new_n4371_;
  assign new_n4373_ = ~\start<0>  & ~new_n4372_;
  assign n1665 = new_n4359_ | new_n4373_;
  assign new_n4375_ = \key<180>  & ~\encrypt<0> ;
  assign new_n4376_ = ~new_n3845_ & ~new_n4375_;
  assign new_n4377_ = \start<0>  & ~new_n4376_;
  assign new_n4378_ = ~new_n1185_1_ & ~new_n2030_1_;
  assign new_n4379_ = new_n1185_1_ & ~new_n2032_;
  assign new_n4380_ = ~new_n4378_ & ~new_n4379_;
  assign new_n4381_ = ~\encrypt<0>  & ~new_n4380_;
  assign new_n4382_ = ~\C<73>  & ~new_n1189_;
  assign new_n4383_ = \C<73>  & new_n1189_;
  assign new_n4384_ = ~new_n4382_ & ~new_n4383_;
  assign new_n4385_ = \D<73>  & ~new_n4384_;
  assign new_n4386_ = \C<73>  & ~new_n1189_;
  assign new_n4387_ = ~\D<73>  & new_n4386_;
  assign new_n4388_ = ~new_n4385_ & ~new_n4387_;
  assign new_n4389_ = \encrypt<0>  & ~new_n4388_;
  assign new_n4390_ = ~new_n4381_ & ~new_n4389_;
  assign new_n4391_ = ~\start<0>  & ~new_n4390_;
  assign n1670 = new_n4377_ | new_n4391_;
  assign new_n4393_ = \key<188>  & ~\encrypt<0> ;
  assign new_n4394_ = \key<180>  & \encrypt<0> ;
  assign new_n4395_ = ~new_n4393_ & ~new_n4394_;
  assign new_n4396_ = \start<0>  & ~new_n4395_;
  assign new_n4397_ = ~new_n1185_1_ & ~new_n2052_;
  assign new_n4398_ = new_n1185_1_ & ~new_n2054_;
  assign new_n4399_ = ~new_n4397_ & ~new_n4398_;
  assign new_n4400_ = ~\encrypt<0>  & ~new_n4399_;
  assign new_n4401_ = ~\C<72>  & ~new_n1189_;
  assign new_n4402_ = \C<72>  & new_n1189_;
  assign new_n4403_ = ~new_n4401_ & ~new_n4402_;
  assign new_n4404_ = \D<72>  & ~new_n4403_;
  assign new_n4405_ = \C<72>  & ~new_n1189_;
  assign new_n4406_ = ~\D<72>  & new_n4405_;
  assign new_n4407_ = ~new_n4404_ & ~new_n4406_;
  assign new_n4408_ = \encrypt<0>  & ~new_n4407_;
  assign new_n4409_ = ~new_n4400_ & ~new_n4408_;
  assign new_n4410_ = ~\start<0>  & ~new_n4409_;
  assign n1675 = new_n4396_ | new_n4410_;
  assign new_n4412_ = \key<133>  & ~\encrypt<0> ;
  assign new_n4413_ = \key<188>  & \encrypt<0> ;
  assign new_n4414_ = ~new_n4412_ & ~new_n4413_;
  assign new_n4415_ = \start<0>  & ~new_n4414_;
  assign new_n4416_ = ~new_n1185_1_ & ~new_n2074_;
  assign new_n4417_ = new_n1185_1_ & ~new_n2076_;
  assign new_n4418_ = ~new_n4416_ & ~new_n4417_;
  assign new_n4419_ = ~\encrypt<0>  & ~new_n4418_;
  assign new_n4420_ = ~\C<71>  & ~new_n1189_;
  assign new_n4421_ = \C<71>  & new_n1189_;
  assign new_n4422_ = ~new_n4420_ & ~new_n4421_;
  assign new_n4423_ = \D<71>  & ~new_n4422_;
  assign new_n4424_ = \C<71>  & ~new_n1189_;
  assign new_n4425_ = ~\D<71>  & new_n4424_;
  assign new_n4426_ = ~new_n4423_ & ~new_n4425_;
  assign new_n4427_ = \encrypt<0>  & ~new_n4426_;
  assign new_n4428_ = ~new_n4419_ & ~new_n4427_;
  assign new_n4429_ = ~\start<0>  & ~new_n4428_;
  assign n1680 = new_n4415_ | new_n4429_;
  assign new_n4431_ = \key<141>  & ~\encrypt<0> ;
  assign new_n4432_ = \key<133>  & \encrypt<0> ;
  assign new_n4433_ = ~new_n4431_ & ~new_n4432_;
  assign new_n4434_ = \start<0>  & ~new_n4433_;
  assign new_n4435_ = ~new_n1185_1_ & ~new_n2096_;
  assign new_n4436_ = new_n1185_1_ & ~new_n2098_;
  assign new_n4437_ = ~new_n4435_ & ~new_n4436_;
  assign new_n4438_ = ~\encrypt<0>  & ~new_n4437_;
  assign new_n4439_ = ~\C<70>  & ~new_n1189_;
  assign new_n4440_ = \C<70>  & new_n1189_;
  assign new_n4441_ = ~new_n4439_ & ~new_n4440_;
  assign new_n4442_ = \D<70>  & ~new_n4441_;
  assign new_n4443_ = \C<70>  & ~new_n1189_;
  assign new_n4444_ = ~\D<70>  & new_n4443_;
  assign new_n4445_ = ~new_n4442_ & ~new_n4444_;
  assign new_n4446_ = \encrypt<0>  & ~new_n4445_;
  assign new_n4447_ = ~new_n4438_ & ~new_n4446_;
  assign new_n4448_ = ~\start<0>  & ~new_n4447_;
  assign n1685 = new_n4434_ | new_n4448_;
  assign new_n4450_ = \key<149>  & ~\encrypt<0> ;
  assign new_n4451_ = \key<141>  & \encrypt<0> ;
  assign new_n4452_ = ~new_n4450_ & ~new_n4451_;
  assign new_n4453_ = \start<0>  & ~new_n4452_;
  assign new_n4454_ = ~new_n1185_1_ & ~new_n2118_;
  assign new_n4455_ = new_n1185_1_ & ~new_n2120_;
  assign new_n4456_ = ~new_n4454_ & ~new_n4455_;
  assign new_n4457_ = ~\encrypt<0>  & ~new_n4456_;
  assign new_n4458_ = ~\C<69>  & ~new_n1189_;
  assign new_n4459_ = \C<69>  & new_n1189_;
  assign new_n4460_ = ~new_n4458_ & ~new_n4459_;
  assign new_n4461_ = \D<69>  & ~new_n4460_;
  assign new_n4462_ = \C<69>  & ~new_n1189_;
  assign new_n4463_ = ~\D<69>  & new_n4462_;
  assign new_n4464_ = ~new_n4461_ & ~new_n4463_;
  assign new_n4465_ = \encrypt<0>  & ~new_n4464_;
  assign new_n4466_ = ~new_n4457_ & ~new_n4465_;
  assign new_n4467_ = ~\start<0>  & ~new_n4466_;
  assign n1690 = new_n4453_ | new_n4467_;
  assign new_n4469_ = \key<157>  & ~\encrypt<0> ;
  assign new_n4470_ = \key<149>  & \encrypt<0> ;
  assign new_n4471_ = ~new_n4469_ & ~new_n4470_;
  assign new_n4472_ = \start<0>  & ~new_n4471_;
  assign new_n4473_ = ~new_n1185_1_ & ~new_n2140_;
  assign new_n4474_ = new_n1185_1_ & ~new_n2142_;
  assign new_n4475_ = ~new_n4473_ & ~new_n4474_;
  assign new_n4476_ = ~\encrypt<0>  & ~new_n4475_;
  assign new_n4477_ = ~\C<68>  & ~new_n1189_;
  assign new_n4478_ = \C<68>  & new_n1189_;
  assign new_n4479_ = ~new_n4477_ & ~new_n4478_;
  assign new_n4480_ = \D<68>  & ~new_n4479_;
  assign new_n4481_ = \C<68>  & ~new_n1189_;
  assign new_n4482_ = ~\D<68>  & new_n4481_;
  assign new_n4483_ = ~new_n4480_ & ~new_n4482_;
  assign new_n4484_ = \encrypt<0>  & ~new_n4483_;
  assign new_n4485_ = ~new_n4476_ & ~new_n4484_;
  assign new_n4486_ = ~\start<0>  & ~new_n4485_;
  assign n1695 = new_n4472_ | new_n4486_;
  assign new_n4488_ = \key<165>  & ~\encrypt<0> ;
  assign new_n4489_ = \key<157>  & \encrypt<0> ;
  assign new_n4490_ = ~new_n4488_ & ~new_n4489_;
  assign new_n4491_ = \start<0>  & ~new_n4490_;
  assign new_n4492_ = ~new_n1185_1_ & ~new_n2162_;
  assign new_n4493_ = new_n1185_1_ & ~new_n2164_;
  assign new_n4494_ = ~new_n4492_ & ~new_n4493_;
  assign new_n4495_ = ~\encrypt<0>  & ~new_n4494_;
  assign new_n4496_ = ~\C<67>  & ~new_n1189_;
  assign new_n4497_ = \C<67>  & new_n1189_;
  assign new_n4498_ = ~new_n4496_ & ~new_n4497_;
  assign new_n4499_ = \D<67>  & ~new_n4498_;
  assign new_n4500_ = \C<67>  & ~new_n1189_;
  assign new_n4501_ = ~\D<67>  & new_n4500_;
  assign new_n4502_ = ~new_n4499_ & ~new_n4501_;
  assign new_n4503_ = \encrypt<0>  & ~new_n4502_;
  assign new_n4504_ = ~new_n4495_ & ~new_n4503_;
  assign new_n4505_ = ~\start<0>  & ~new_n4504_;
  assign n1700 = new_n4491_ | new_n4505_;
  assign new_n4507_ = \key<173>  & ~\encrypt<0> ;
  assign new_n4508_ = \key<165>  & \encrypt<0> ;
  assign new_n4509_ = ~new_n4507_ & ~new_n4508_;
  assign new_n4510_ = \start<0>  & ~new_n4509_;
  assign new_n4511_ = ~new_n1185_1_ & ~new_n2184_;
  assign new_n4512_ = new_n1185_1_ & ~new_n2186_;
  assign new_n4513_ = ~new_n4511_ & ~new_n4512_;
  assign new_n4514_ = ~\encrypt<0>  & ~new_n4513_;
  assign new_n4515_ = ~\C<66>  & ~new_n1189_;
  assign new_n4516_ = \C<66>  & new_n1189_;
  assign new_n4517_ = ~new_n4515_ & ~new_n4516_;
  assign new_n4518_ = \D<66>  & ~new_n4517_;
  assign new_n4519_ = \C<66>  & ~new_n1189_;
  assign new_n4520_ = ~\D<66>  & new_n4519_;
  assign new_n4521_ = ~new_n4518_ & ~new_n4520_;
  assign new_n4522_ = \encrypt<0>  & ~new_n4521_;
  assign new_n4523_ = ~new_n4514_ & ~new_n4522_;
  assign new_n4524_ = ~\start<0>  & ~new_n4523_;
  assign n1705 = new_n4510_ | new_n4524_;
  assign new_n4526_ = \key<181>  & ~\encrypt<0> ;
  assign new_n4527_ = \key<173>  & \encrypt<0> ;
  assign new_n4528_ = ~new_n4526_ & ~new_n4527_;
  assign new_n4529_ = \start<0>  & ~new_n4528_;
  assign new_n4530_ = ~new_n1185_1_ & ~new_n2206_;
  assign new_n4531_ = new_n1185_1_ & ~new_n2208_;
  assign new_n4532_ = ~new_n4530_ & ~new_n4531_;
  assign new_n4533_ = ~\encrypt<0>  & ~new_n4532_;
  assign new_n4534_ = ~\C<65>  & ~new_n1189_;
  assign new_n4535_ = \C<65>  & new_n1189_;
  assign new_n4536_ = ~new_n4534_ & ~new_n4535_;
  assign new_n4537_ = \D<65>  & ~new_n4536_;
  assign new_n4538_ = \C<65>  & ~new_n1189_;
  assign new_n4539_ = ~\D<65>  & new_n4538_;
  assign new_n4540_ = ~new_n4537_ & ~new_n4539_;
  assign new_n4541_ = \encrypt<0>  & ~new_n4540_;
  assign new_n4542_ = ~new_n4533_ & ~new_n4541_;
  assign new_n4543_ = ~\start<0>  & ~new_n4542_;
  assign n1710 = new_n4529_ | new_n4543_;
  assign new_n4545_ = \key<189>  & ~\encrypt<0> ;
  assign new_n4546_ = \key<181>  & \encrypt<0> ;
  assign new_n4547_ = ~new_n4545_ & ~new_n4546_;
  assign new_n4548_ = \start<0>  & ~new_n4547_;
  assign new_n4549_ = ~new_n1185_1_ & ~new_n2228_;
  assign new_n4550_ = new_n1185_1_ & ~new_n2230_;
  assign new_n4551_ = ~new_n4549_ & ~new_n4550_;
  assign new_n4552_ = ~\encrypt<0>  & ~new_n4551_;
  assign new_n4553_ = ~\C<64>  & ~new_n1189_;
  assign new_n4554_ = \C<64>  & new_n1189_;
  assign new_n4555_ = ~new_n4553_ & ~new_n4554_;
  assign new_n4556_ = \D<64>  & ~new_n4555_;
  assign new_n4557_ = \C<64>  & ~new_n1189_;
  assign new_n4558_ = ~\D<64>  & new_n4557_;
  assign new_n4559_ = ~new_n4556_ & ~new_n4558_;
  assign new_n4560_ = \encrypt<0>  & ~new_n4559_;
  assign new_n4561_ = ~new_n4552_ & ~new_n4560_;
  assign new_n4562_ = ~\start<0>  & ~new_n4561_;
  assign n1715 = new_n4548_ | new_n4562_;
  assign new_n4564_ = \key<134>  & ~\encrypt<0> ;
  assign new_n4565_ = \key<189>  & \encrypt<0> ;
  assign new_n4566_ = ~new_n4564_ & ~new_n4565_;
  assign new_n4567_ = \start<0>  & ~new_n4566_;
  assign new_n4568_ = ~new_n1185_1_ & ~new_n2250_;
  assign new_n4569_ = new_n1185_1_ & ~new_n2252_;
  assign new_n4570_ = ~new_n4568_ & ~new_n4569_;
  assign new_n4571_ = ~\encrypt<0>  & ~new_n4570_;
  assign new_n4572_ = ~\C<63>  & ~new_n1189_;
  assign new_n4573_ = \C<63>  & new_n1189_;
  assign new_n4574_ = ~new_n4572_ & ~new_n4573_;
  assign new_n4575_ = \D<63>  & ~new_n4574_;
  assign new_n4576_ = \C<63>  & ~new_n1189_;
  assign new_n4577_ = ~\D<63>  & new_n4576_;
  assign new_n4578_ = ~new_n4575_ & ~new_n4577_;
  assign new_n4579_ = \encrypt<0>  & ~new_n4578_;
  assign new_n4580_ = ~new_n4571_ & ~new_n4579_;
  assign new_n4581_ = ~\start<0>  & ~new_n4580_;
  assign n1720 = new_n4567_ | new_n4581_;
  assign new_n4583_ = \key<142>  & ~\encrypt<0> ;
  assign new_n4584_ = \key<134>  & \encrypt<0> ;
  assign new_n4585_ = ~new_n4583_ & ~new_n4584_;
  assign new_n4586_ = \start<0>  & ~new_n4585_;
  assign new_n4587_ = ~new_n1185_1_ & ~new_n2272_;
  assign new_n4588_ = new_n1185_1_ & ~new_n2274_;
  assign new_n4589_ = ~new_n4587_ & ~new_n4588_;
  assign new_n4590_ = ~\encrypt<0>  & ~new_n4589_;
  assign new_n4591_ = ~\C<62>  & ~new_n1189_;
  assign new_n4592_ = \C<62>  & new_n1189_;
  assign new_n4593_ = ~new_n4591_ & ~new_n4592_;
  assign new_n4594_ = \D<62>  & ~new_n4593_;
  assign new_n4595_ = \C<62>  & ~new_n1189_;
  assign new_n4596_ = ~\D<62>  & new_n4595_;
  assign new_n4597_ = ~new_n4594_ & ~new_n4596_;
  assign new_n4598_ = \encrypt<0>  & ~new_n4597_;
  assign new_n4599_ = ~new_n4590_ & ~new_n4598_;
  assign new_n4600_ = ~\start<0>  & ~new_n4599_;
  assign n1725 = new_n4586_ | new_n4600_;
  assign new_n4602_ = \key<150>  & ~\encrypt<0> ;
  assign new_n4603_ = \key<142>  & \encrypt<0> ;
  assign new_n4604_ = ~new_n4602_ & ~new_n4603_;
  assign new_n4605_ = \start<0>  & ~new_n4604_;
  assign new_n4606_ = ~new_n1185_1_ & ~new_n2294_;
  assign new_n4607_ = new_n1185_1_ & ~new_n2296_;
  assign new_n4608_ = ~new_n4606_ & ~new_n4607_;
  assign new_n4609_ = ~\encrypt<0>  & ~new_n4608_;
  assign new_n4610_ = ~\C<61>  & ~new_n1189_;
  assign new_n4611_ = \C<61>  & new_n1189_;
  assign new_n4612_ = ~new_n4610_ & ~new_n4611_;
  assign new_n4613_ = \D<61>  & ~new_n4612_;
  assign new_n4614_ = \C<61>  & ~new_n1189_;
  assign new_n4615_ = ~\D<61>  & new_n4614_;
  assign new_n4616_ = ~new_n4613_ & ~new_n4615_;
  assign new_n4617_ = \encrypt<0>  & ~new_n4616_;
  assign new_n4618_ = ~new_n4609_ & ~new_n4617_;
  assign new_n4619_ = ~\start<0>  & ~new_n4618_;
  assign n1730 = new_n4605_ | new_n4619_;
  assign new_n4621_ = \key<158>  & ~\encrypt<0> ;
  assign new_n4622_ = \key<150>  & \encrypt<0> ;
  assign new_n4623_ = ~new_n4621_ & ~new_n4622_;
  assign new_n4624_ = \start<0>  & ~new_n4623_;
  assign new_n4625_ = ~new_n1185_1_ & ~new_n2316_;
  assign new_n4626_ = new_n1185_1_ & ~new_n2318_;
  assign new_n4627_ = ~new_n4625_ & ~new_n4626_;
  assign new_n4628_ = ~\encrypt<0>  & ~new_n4627_;
  assign new_n4629_ = ~\C<60>  & ~new_n1189_;
  assign new_n4630_ = \C<60>  & new_n1189_;
  assign new_n4631_ = ~new_n4629_ & ~new_n4630_;
  assign new_n4632_ = \D<60>  & ~new_n4631_;
  assign new_n4633_ = \C<60>  & ~new_n1189_;
  assign new_n4634_ = ~\D<60>  & new_n4633_;
  assign new_n4635_ = ~new_n4632_ & ~new_n4634_;
  assign new_n4636_ = \encrypt<0>  & ~new_n4635_;
  assign new_n4637_ = ~new_n4628_ & ~new_n4636_;
  assign new_n4638_ = ~\start<0>  & ~new_n4637_;
  assign n1735 = new_n4624_ | new_n4638_;
  assign new_n4640_ = \key<166>  & ~\encrypt<0> ;
  assign new_n4641_ = \key<158>  & \encrypt<0> ;
  assign new_n4642_ = ~new_n4640_ & ~new_n4641_;
  assign new_n4643_ = \start<0>  & ~new_n4642_;
  assign new_n4644_ = ~new_n1185_1_ & ~new_n2338_;
  assign new_n4645_ = new_n1185_1_ & ~new_n2340_;
  assign new_n4646_ = ~new_n4644_ & ~new_n4645_;
  assign new_n4647_ = ~\encrypt<0>  & ~new_n4646_;
  assign new_n4648_ = ~\C<59>  & ~new_n1189_;
  assign new_n4649_ = \C<59>  & new_n1189_;
  assign new_n4650_ = ~new_n4648_ & ~new_n4649_;
  assign new_n4651_ = \D<59>  & ~new_n4650_;
  assign new_n4652_ = \C<59>  & ~new_n1189_;
  assign new_n4653_ = ~\D<59>  & new_n4652_;
  assign new_n4654_ = ~new_n4651_ & ~new_n4653_;
  assign new_n4655_ = \encrypt<0>  & ~new_n4654_;
  assign new_n4656_ = ~new_n4647_ & ~new_n4655_;
  assign new_n4657_ = ~\start<0>  & ~new_n4656_;
  assign n1740 = new_n4643_ | new_n4657_;
  assign new_n4659_ = \key<174>  & ~\encrypt<0> ;
  assign new_n4660_ = \key<166>  & \encrypt<0> ;
  assign new_n4661_ = ~new_n4659_ & ~new_n4660_;
  assign new_n4662_ = \start<0>  & ~new_n4661_;
  assign new_n4663_ = ~new_n1185_1_ & ~new_n2360_;
  assign new_n4664_ = new_n1185_1_ & ~new_n2362_;
  assign new_n4665_ = ~new_n4663_ & ~new_n4664_;
  assign new_n4666_ = ~\encrypt<0>  & ~new_n4665_;
  assign new_n4667_ = ~\C<58>  & ~new_n1189_;
  assign new_n4668_ = \C<58>  & new_n1189_;
  assign new_n4669_ = ~new_n4667_ & ~new_n4668_;
  assign new_n4670_ = \D<58>  & ~new_n4669_;
  assign new_n4671_ = \C<58>  & ~new_n1189_;
  assign new_n4672_ = ~\D<58>  & new_n4671_;
  assign new_n4673_ = ~new_n4670_ & ~new_n4672_;
  assign new_n4674_ = \encrypt<0>  & ~new_n4673_;
  assign new_n4675_ = ~new_n4666_ & ~new_n4674_;
  assign new_n4676_ = ~\start<0>  & ~new_n4675_;
  assign n1745 = new_n4662_ | new_n4676_;
  assign new_n4678_ = \key<182>  & ~\encrypt<0> ;
  assign new_n4679_ = \key<174>  & \encrypt<0> ;
  assign new_n4680_ = ~new_n4678_ & ~new_n4679_;
  assign new_n4681_ = \start<0>  & ~new_n4680_;
  assign new_n4682_ = ~new_n1185_1_ & ~new_n2382_;
  assign new_n4683_ = new_n1185_1_ & ~new_n2384_;
  assign new_n4684_ = ~new_n4682_ & ~new_n4683_;
  assign new_n4685_ = ~\encrypt<0>  & ~new_n4684_;
  assign new_n4686_ = ~\C<57>  & ~new_n1189_;
  assign new_n4687_ = \C<57>  & new_n1189_;
  assign new_n4688_ = ~new_n4686_ & ~new_n4687_;
  assign new_n4689_ = \D<57>  & ~new_n4688_;
  assign new_n4690_ = \C<57>  & ~new_n1189_;
  assign new_n4691_ = ~\D<57>  & new_n4690_;
  assign new_n4692_ = ~new_n4689_ & ~new_n4691_;
  assign new_n4693_ = \encrypt<0>  & ~new_n4692_;
  assign new_n4694_ = ~new_n4685_ & ~new_n4693_;
  assign new_n4695_ = ~\start<0>  & ~new_n4694_;
  assign n1750 = new_n4681_ | new_n4695_;
  assign new_n4697_ = \key<190>  & ~\encrypt<0> ;
  assign new_n4698_ = \key<182>  & \encrypt<0> ;
  assign new_n4699_ = ~new_n4697_ & ~new_n4698_;
  assign new_n4700_ = \start<0>  & ~new_n4699_;
  assign new_n4701_ = ~new_n1185_1_ & ~new_n2404_;
  assign new_n4702_ = new_n1185_1_ & ~new_n2406_;
  assign new_n4703_ = ~new_n4701_ & ~new_n4702_;
  assign new_n4704_ = ~\encrypt<0>  & ~new_n4703_;
  assign new_n4705_ = ~\C<56>  & ~new_n1189_;
  assign new_n4706_ = \C<56>  & new_n1189_;
  assign new_n4707_ = ~new_n4705_ & ~new_n4706_;
  assign new_n4708_ = \D<56>  & ~new_n4707_;
  assign new_n4709_ = \C<56>  & ~new_n1189_;
  assign new_n4710_ = ~\D<56>  & new_n4709_;
  assign new_n4711_ = ~new_n4708_ & ~new_n4710_;
  assign new_n4712_ = \encrypt<0>  & ~new_n4711_;
  assign new_n4713_ = ~new_n4704_ & ~new_n4712_;
  assign new_n4714_ = ~\start<0>  & ~new_n4713_;
  assign n1755 = new_n4700_ | new_n4714_;
  assign new_n4716_ = \key<67>  & ~\encrypt<0> ;
  assign new_n4717_ = \key<190>  & \encrypt<0> ;
  assign new_n4718_ = ~new_n4716_ & ~new_n4717_;
  assign new_n4719_ = \start<0>  & ~new_n4718_;
  assign new_n4720_ = ~new_n1185_1_ & ~new_n2426_;
  assign new_n4721_ = new_n1185_1_ & ~new_n2428_;
  assign new_n4722_ = ~new_n4720_ & ~new_n4721_;
  assign new_n4723_ = ~\encrypt<0>  & ~new_n4722_;
  assign new_n4724_ = ~\C<55>  & ~new_n1189_;
  assign new_n4725_ = \C<55>  & new_n1189_;
  assign new_n4726_ = ~new_n4724_ & ~new_n4725_;
  assign new_n4727_ = \D<55>  & ~new_n4726_;
  assign new_n4728_ = \C<55>  & ~new_n1189_;
  assign new_n4729_ = ~\D<55>  & new_n4728_;
  assign new_n4730_ = ~new_n4727_ & ~new_n4729_;
  assign new_n4731_ = \encrypt<0>  & ~new_n4730_;
  assign new_n4732_ = ~new_n4723_ & ~new_n4731_;
  assign new_n4733_ = ~\start<0>  & ~new_n4732_;
  assign n1760 = new_n4719_ | new_n4733_;
  assign new_n4735_ = \key<75>  & ~\encrypt<0> ;
  assign new_n4736_ = \key<67>  & \encrypt<0> ;
  assign new_n4737_ = ~new_n4735_ & ~new_n4736_;
  assign new_n4738_ = \start<0>  & ~new_n4737_;
  assign new_n4739_ = ~new_n1185_1_ & ~new_n2448_;
  assign new_n4740_ = new_n1185_1_ & ~new_n2450_;
  assign new_n4741_ = ~new_n4739_ & ~new_n4740_;
  assign new_n4742_ = ~\encrypt<0>  & ~new_n4741_;
  assign new_n4743_ = ~\C<54>  & ~new_n1189_;
  assign new_n4744_ = \C<54>  & new_n1189_;
  assign new_n4745_ = ~new_n4743_ & ~new_n4744_;
  assign new_n4746_ = \D<54>  & ~new_n4745_;
  assign new_n4747_ = \C<54>  & ~new_n1189_;
  assign new_n4748_ = ~\D<54>  & new_n4747_;
  assign new_n4749_ = ~new_n4746_ & ~new_n4748_;
  assign new_n4750_ = \encrypt<0>  & ~new_n4749_;
  assign new_n4751_ = ~new_n4742_ & ~new_n4750_;
  assign new_n4752_ = ~\start<0>  & ~new_n4751_;
  assign n1765 = new_n4738_ | new_n4752_;
  assign new_n4754_ = \key<83>  & ~\encrypt<0> ;
  assign new_n4755_ = \key<75>  & \encrypt<0> ;
  assign new_n4756_ = ~new_n4754_ & ~new_n4755_;
  assign new_n4757_ = \start<0>  & ~new_n4756_;
  assign new_n4758_ = ~new_n1185_1_ & ~new_n2470_;
  assign new_n4759_ = new_n1185_1_ & ~new_n2472_;
  assign new_n4760_ = ~new_n4758_ & ~new_n4759_;
  assign new_n4761_ = ~\encrypt<0>  & ~new_n4760_;
  assign new_n4762_ = ~\C<53>  & ~new_n1189_;
  assign new_n4763_ = \C<53>  & new_n1189_;
  assign new_n4764_ = ~new_n4762_ & ~new_n4763_;
  assign new_n4765_ = \D<53>  & ~new_n4764_;
  assign new_n4766_ = \C<53>  & ~new_n1189_;
  assign new_n4767_ = ~\D<53>  & new_n4766_;
  assign new_n4768_ = ~new_n4765_ & ~new_n4767_;
  assign new_n4769_ = \encrypt<0>  & ~new_n4768_;
  assign new_n4770_ = ~new_n4761_ & ~new_n4769_;
  assign new_n4771_ = ~\start<0>  & ~new_n4770_;
  assign n1770 = new_n4757_ | new_n4771_;
  assign new_n4773_ = \key<91>  & ~\encrypt<0> ;
  assign new_n4774_ = \key<83>  & \encrypt<0> ;
  assign new_n4775_ = ~new_n4773_ & ~new_n4774_;
  assign new_n4776_ = \start<0>  & ~new_n4775_;
  assign new_n4777_ = ~new_n1185_1_ & ~new_n2492_;
  assign new_n4778_ = new_n1185_1_ & ~new_n2494_;
  assign new_n4779_ = ~new_n4777_ & ~new_n4778_;
  assign new_n4780_ = ~\encrypt<0>  & ~new_n4779_;
  assign new_n4781_ = ~\C<52>  & ~new_n1189_;
  assign new_n4782_ = \C<52>  & new_n1189_;
  assign new_n4783_ = ~new_n4781_ & ~new_n4782_;
  assign new_n4784_ = \D<52>  & ~new_n4783_;
  assign new_n4785_ = \C<52>  & ~new_n1189_;
  assign new_n4786_ = ~\D<52>  & new_n4785_;
  assign new_n4787_ = ~new_n4784_ & ~new_n4786_;
  assign new_n4788_ = \encrypt<0>  & ~new_n4787_;
  assign new_n4789_ = ~new_n4780_ & ~new_n4788_;
  assign new_n4790_ = ~\start<0>  & ~new_n4789_;
  assign n1775 = new_n4776_ | new_n4790_;
  assign new_n4792_ = \key<68>  & ~\encrypt<0> ;
  assign new_n4793_ = \key<91>  & \encrypt<0> ;
  assign new_n4794_ = ~new_n4792_ & ~new_n4793_;
  assign new_n4795_ = \start<0>  & ~new_n4794_;
  assign new_n4796_ = ~new_n1185_1_ & ~new_n2514_;
  assign new_n4797_ = new_n1185_1_ & ~new_n2516_;
  assign new_n4798_ = ~new_n4796_ & ~new_n4797_;
  assign new_n4799_ = ~\encrypt<0>  & ~new_n4798_;
  assign new_n4800_ = ~\C<51>  & ~new_n1189_;
  assign new_n4801_ = \C<51>  & new_n1189_;
  assign new_n4802_ = ~new_n4800_ & ~new_n4801_;
  assign new_n4803_ = \D<51>  & ~new_n4802_;
  assign new_n4804_ = \C<51>  & ~new_n1189_;
  assign new_n4805_ = ~\D<51>  & new_n4804_;
  assign new_n4806_ = ~new_n4803_ & ~new_n4805_;
  assign new_n4807_ = \encrypt<0>  & ~new_n4806_;
  assign new_n4808_ = ~new_n4799_ & ~new_n4807_;
  assign new_n4809_ = ~\start<0>  & ~new_n4808_;
  assign n1780 = new_n4795_ | new_n4809_;
  assign new_n4811_ = \key<76>  & ~\encrypt<0> ;
  assign new_n4812_ = \key<68>  & \encrypt<0> ;
  assign new_n4813_ = ~new_n4811_ & ~new_n4812_;
  assign new_n4814_ = \start<0>  & ~new_n4813_;
  assign new_n4815_ = ~new_n1185_1_ & ~new_n2536_;
  assign new_n4816_ = new_n1185_1_ & ~new_n2538_;
  assign new_n4817_ = ~new_n4815_ & ~new_n4816_;
  assign new_n4818_ = ~\encrypt<0>  & ~new_n4817_;
  assign new_n4819_ = ~\C<50>  & ~new_n1189_;
  assign new_n4820_ = \C<50>  & new_n1189_;
  assign new_n4821_ = ~new_n4819_ & ~new_n4820_;
  assign new_n4822_ = \D<50>  & ~new_n4821_;
  assign new_n4823_ = \C<50>  & ~new_n1189_;
  assign new_n4824_ = ~\D<50>  & new_n4823_;
  assign new_n4825_ = ~new_n4822_ & ~new_n4824_;
  assign new_n4826_ = \encrypt<0>  & ~new_n4825_;
  assign new_n4827_ = ~new_n4818_ & ~new_n4826_;
  assign new_n4828_ = ~\start<0>  & ~new_n4827_;
  assign n1785 = new_n4814_ | new_n4828_;
  assign new_n4830_ = \key<84>  & ~\encrypt<0> ;
  assign new_n4831_ = \key<76>  & \encrypt<0> ;
  assign new_n4832_ = ~new_n4830_ & ~new_n4831_;
  assign new_n4833_ = \start<0>  & ~new_n4832_;
  assign new_n4834_ = ~new_n1185_1_ & ~new_n2558_;
  assign new_n4835_ = new_n1185_1_ & ~new_n2560_;
  assign new_n4836_ = ~new_n4834_ & ~new_n4835_;
  assign new_n4837_ = ~\encrypt<0>  & ~new_n4836_;
  assign new_n4838_ = ~\C<49>  & ~new_n1189_;
  assign new_n4839_ = \C<49>  & new_n1189_;
  assign new_n4840_ = ~new_n4838_ & ~new_n4839_;
  assign new_n4841_ = \D<49>  & ~new_n4840_;
  assign new_n4842_ = \C<49>  & ~new_n1189_;
  assign new_n4843_ = ~\D<49>  & new_n4842_;
  assign new_n4844_ = ~new_n4841_ & ~new_n4843_;
  assign new_n4845_ = \encrypt<0>  & ~new_n4844_;
  assign new_n4846_ = ~new_n4837_ & ~new_n4845_;
  assign new_n4847_ = ~\start<0>  & ~new_n4846_;
  assign n1790 = new_n4833_ | new_n4847_;
  assign new_n4849_ = \key<92>  & ~\encrypt<0> ;
  assign new_n4850_ = \key<84>  & \encrypt<0> ;
  assign new_n4851_ = ~new_n4849_ & ~new_n4850_;
  assign new_n4852_ = \start<0>  & ~new_n4851_;
  assign new_n4853_ = ~new_n1185_1_ & ~new_n2580_;
  assign new_n4854_ = new_n1185_1_ & ~new_n2582_;
  assign new_n4855_ = ~new_n4853_ & ~new_n4854_;
  assign new_n4856_ = ~\encrypt<0>  & ~new_n4855_;
  assign new_n4857_ = ~\C<48>  & ~new_n1189_;
  assign new_n4858_ = \C<48>  & new_n1189_;
  assign new_n4859_ = ~new_n4857_ & ~new_n4858_;
  assign new_n4860_ = \D<48>  & ~new_n4859_;
  assign new_n4861_ = \C<48>  & ~new_n1189_;
  assign new_n4862_ = ~\D<48>  & new_n4861_;
  assign new_n4863_ = ~new_n4860_ & ~new_n4862_;
  assign new_n4864_ = \encrypt<0>  & ~new_n4863_;
  assign new_n4865_ = ~new_n4856_ & ~new_n4864_;
  assign new_n4866_ = ~\start<0>  & ~new_n4865_;
  assign n1795 = new_n4852_ | new_n4866_;
  assign new_n4868_ = \key<100>  & ~\encrypt<0> ;
  assign new_n4869_ = \key<92>  & \encrypt<0> ;
  assign new_n4870_ = ~new_n4868_ & ~new_n4869_;
  assign new_n4871_ = \start<0>  & ~new_n4870_;
  assign new_n4872_ = ~new_n1185_1_ & ~new_n2602_;
  assign new_n4873_ = new_n1185_1_ & ~new_n2604_;
  assign new_n4874_ = ~new_n4872_ & ~new_n4873_;
  assign new_n4875_ = ~\encrypt<0>  & ~new_n4874_;
  assign new_n4876_ = ~\C<47>  & ~new_n1189_;
  assign new_n4877_ = \C<47>  & new_n1189_;
  assign new_n4878_ = ~new_n4876_ & ~new_n4877_;
  assign new_n4879_ = \D<47>  & ~new_n4878_;
  assign new_n4880_ = \C<47>  & ~new_n1189_;
  assign new_n4881_ = ~\D<47>  & new_n4880_;
  assign new_n4882_ = ~new_n4879_ & ~new_n4881_;
  assign new_n4883_ = \encrypt<0>  & ~new_n4882_;
  assign new_n4884_ = ~new_n4875_ & ~new_n4883_;
  assign new_n4885_ = ~\start<0>  & ~new_n4884_;
  assign n1800 = new_n4871_ | new_n4885_;
  assign new_n4887_ = \key<44>  & ~\encrypt<0> ;
  assign new_n4888_ = \key<100>  & \encrypt<0> ;
  assign new_n4889_ = ~new_n4887_ & ~new_n4888_;
  assign new_n4890_ = \start<0>  & ~new_n4889_;
  assign new_n4891_ = ~new_n1185_1_ & ~new_n2624_;
  assign new_n4892_ = new_n1185_1_ & ~new_n2626_;
  assign new_n4893_ = ~new_n4891_ & ~new_n4892_;
  assign new_n4894_ = ~\encrypt<0>  & ~new_n4893_;
  assign new_n4895_ = ~\C<46>  & ~new_n1189_;
  assign new_n4896_ = \C<46>  & new_n1189_;
  assign new_n4897_ = ~new_n4895_ & ~new_n4896_;
  assign new_n4898_ = \D<46>  & ~new_n4897_;
  assign new_n4899_ = \C<46>  & ~new_n1189_;
  assign new_n4900_ = ~\D<46>  & new_n4899_;
  assign new_n4901_ = ~new_n4898_ & ~new_n4900_;
  assign new_n4902_ = \encrypt<0>  & ~new_n4901_;
  assign new_n4903_ = ~new_n4894_ & ~new_n4902_;
  assign new_n4904_ = ~\start<0>  & ~new_n4903_;
  assign n1805 = new_n4890_ | new_n4904_;
  assign new_n4906_ = \key<116>  & ~\encrypt<0> ;
  assign new_n4907_ = \key<44>  & \encrypt<0> ;
  assign new_n4908_ = ~new_n4906_ & ~new_n4907_;
  assign new_n4909_ = \start<0>  & ~new_n4908_;
  assign new_n4910_ = ~new_n1185_1_ & ~new_n2646_;
  assign new_n4911_ = new_n1185_1_ & ~new_n2648_;
  assign new_n4912_ = ~new_n4910_ & ~new_n4911_;
  assign new_n4913_ = ~\encrypt<0>  & ~new_n4912_;
  assign new_n4914_ = ~\C<45>  & ~new_n1189_;
  assign new_n4915_ = \C<45>  & new_n1189_;
  assign new_n4916_ = ~new_n4914_ & ~new_n4915_;
  assign new_n4917_ = \D<45>  & ~new_n4916_;
  assign new_n4918_ = \C<45>  & ~new_n1189_;
  assign new_n4919_ = ~\D<45>  & new_n4918_;
  assign new_n4920_ = ~new_n4917_ & ~new_n4919_;
  assign new_n4921_ = \encrypt<0>  & ~new_n4920_;
  assign new_n4922_ = ~new_n4913_ & ~new_n4921_;
  assign new_n4923_ = ~\start<0>  & ~new_n4922_;
  assign n1810 = new_n4909_ | new_n4923_;
  assign new_n4925_ = \key<124>  & ~\encrypt<0> ;
  assign new_n4926_ = \key<116>  & \encrypt<0> ;
  assign new_n4927_ = ~new_n4925_ & ~new_n4926_;
  assign new_n4928_ = \start<0>  & ~new_n4927_;
  assign new_n4929_ = ~new_n1185_1_ & ~new_n2668_;
  assign new_n4930_ = new_n1185_1_ & ~new_n2670_;
  assign new_n4931_ = ~new_n4929_ & ~new_n4930_;
  assign new_n4932_ = ~\encrypt<0>  & ~new_n4931_;
  assign new_n4933_ = ~\C<44>  & ~new_n1189_;
  assign new_n4934_ = \C<44>  & new_n1189_;
  assign new_n4935_ = ~new_n4933_ & ~new_n4934_;
  assign new_n4936_ = \D<44>  & ~new_n4935_;
  assign new_n4937_ = \C<44>  & ~new_n1189_;
  assign new_n4938_ = ~\D<44>  & new_n4937_;
  assign new_n4939_ = ~new_n4936_ & ~new_n4938_;
  assign new_n4940_ = \encrypt<0>  & ~new_n4939_;
  assign new_n4941_ = ~new_n4932_ & ~new_n4940_;
  assign new_n4942_ = ~\start<0>  & ~new_n4941_;
  assign n1815 = new_n4928_ | new_n4942_;
  assign new_n4944_ = \key<69>  & ~\encrypt<0> ;
  assign new_n4945_ = \key<124>  & \encrypt<0> ;
  assign new_n4946_ = ~new_n4944_ & ~new_n4945_;
  assign new_n4947_ = \start<0>  & ~new_n4946_;
  assign new_n4948_ = ~new_n1185_1_ & ~new_n2690_;
  assign new_n4949_ = new_n1185_1_ & ~new_n2692_;
  assign new_n4950_ = ~new_n4948_ & ~new_n4949_;
  assign new_n4951_ = ~\encrypt<0>  & ~new_n4950_;
  assign new_n4952_ = ~\C<43>  & ~new_n1189_;
  assign new_n4953_ = \C<43>  & new_n1189_;
  assign new_n4954_ = ~new_n4952_ & ~new_n4953_;
  assign new_n4955_ = \D<43>  & ~new_n4954_;
  assign new_n4956_ = \C<43>  & ~new_n1189_;
  assign new_n4957_ = ~\D<43>  & new_n4956_;
  assign new_n4958_ = ~new_n4955_ & ~new_n4957_;
  assign new_n4959_ = \encrypt<0>  & ~new_n4958_;
  assign new_n4960_ = ~new_n4951_ & ~new_n4959_;
  assign new_n4961_ = ~\start<0>  & ~new_n4960_;
  assign n1820 = new_n4947_ | new_n4961_;
  assign new_n4963_ = \key<77>  & ~\encrypt<0> ;
  assign new_n4964_ = \key<69>  & \encrypt<0> ;
  assign new_n4965_ = ~new_n4963_ & ~new_n4964_;
  assign new_n4966_ = \start<0>  & ~new_n4965_;
  assign new_n4967_ = ~new_n1185_1_ & ~new_n2712_;
  assign new_n4968_ = new_n1185_1_ & ~new_n2714_;
  assign new_n4969_ = ~new_n4967_ & ~new_n4968_;
  assign new_n4970_ = ~\encrypt<0>  & ~new_n4969_;
  assign new_n4971_ = ~\C<42>  & ~new_n1189_;
  assign new_n4972_ = \C<42>  & new_n1189_;
  assign new_n4973_ = ~new_n4971_ & ~new_n4972_;
  assign new_n4974_ = \D<42>  & ~new_n4973_;
  assign new_n4975_ = \C<42>  & ~new_n1189_;
  assign new_n4976_ = ~\D<42>  & new_n4975_;
  assign new_n4977_ = ~new_n4974_ & ~new_n4976_;
  assign new_n4978_ = \encrypt<0>  & ~new_n4977_;
  assign new_n4979_ = ~new_n4970_ & ~new_n4978_;
  assign new_n4980_ = ~\start<0>  & ~new_n4979_;
  assign n1825 = new_n4966_ | new_n4980_;
  assign new_n4982_ = \key<85>  & ~\encrypt<0> ;
  assign new_n4983_ = \key<77>  & \encrypt<0> ;
  assign new_n4984_ = ~new_n4982_ & ~new_n4983_;
  assign new_n4985_ = \start<0>  & ~new_n4984_;
  assign new_n4986_ = ~new_n1185_1_ & ~new_n2734_;
  assign new_n4987_ = new_n1185_1_ & ~new_n2736_;
  assign new_n4988_ = ~new_n4986_ & ~new_n4987_;
  assign new_n4989_ = ~\encrypt<0>  & ~new_n4988_;
  assign new_n4990_ = ~\C<41>  & ~new_n1189_;
  assign new_n4991_ = \C<41>  & new_n1189_;
  assign new_n4992_ = ~new_n4990_ & ~new_n4991_;
  assign new_n4993_ = \D<41>  & ~new_n4992_;
  assign new_n4994_ = \C<41>  & ~new_n1189_;
  assign new_n4995_ = ~\D<41>  & new_n4994_;
  assign new_n4996_ = ~new_n4993_ & ~new_n4995_;
  assign new_n4997_ = \encrypt<0>  & ~new_n4996_;
  assign new_n4998_ = ~new_n4989_ & ~new_n4997_;
  assign new_n4999_ = ~\start<0>  & ~new_n4998_;
  assign n1830 = new_n4985_ | new_n4999_;
  assign new_n5001_ = \key<93>  & ~\encrypt<0> ;
  assign new_n5002_ = \key<85>  & \encrypt<0> ;
  assign new_n5003_ = ~new_n5001_ & ~new_n5002_;
  assign new_n5004_ = \start<0>  & ~new_n5003_;
  assign new_n5005_ = ~new_n1185_1_ & ~new_n2756_;
  assign new_n5006_ = new_n1185_1_ & ~new_n2758_;
  assign new_n5007_ = ~new_n5005_ & ~new_n5006_;
  assign new_n5008_ = ~\encrypt<0>  & ~new_n5007_;
  assign new_n5009_ = ~\C<40>  & ~new_n1189_;
  assign new_n5010_ = \C<40>  & new_n1189_;
  assign new_n5011_ = ~new_n5009_ & ~new_n5010_;
  assign new_n5012_ = \D<40>  & ~new_n5011_;
  assign new_n5013_ = \C<40>  & ~new_n1189_;
  assign new_n5014_ = ~\D<40>  & new_n5013_;
  assign new_n5015_ = ~new_n5012_ & ~new_n5014_;
  assign new_n5016_ = \encrypt<0>  & ~new_n5015_;
  assign new_n5017_ = ~new_n5008_ & ~new_n5016_;
  assign new_n5018_ = ~\start<0>  & ~new_n5017_;
  assign n1835 = new_n5004_ | new_n5018_;
  assign new_n5020_ = \key<101>  & ~\encrypt<0> ;
  assign new_n5021_ = \key<93>  & \encrypt<0> ;
  assign new_n5022_ = ~new_n5020_ & ~new_n5021_;
  assign new_n5023_ = \start<0>  & ~new_n5022_;
  assign new_n5024_ = ~new_n1185_1_ & ~new_n2778_;
  assign new_n5025_ = new_n1185_1_ & ~new_n2780_;
  assign new_n5026_ = ~new_n5024_ & ~new_n5025_;
  assign new_n5027_ = ~\encrypt<0>  & ~new_n5026_;
  assign new_n5028_ = ~\C<39>  & ~new_n1189_;
  assign new_n5029_ = \C<39>  & new_n1189_;
  assign new_n5030_ = ~new_n5028_ & ~new_n5029_;
  assign new_n5031_ = \D<39>  & ~new_n5030_;
  assign new_n5032_ = \C<39>  & ~new_n1189_;
  assign new_n5033_ = ~\D<39>  & new_n5032_;
  assign new_n5034_ = ~new_n5031_ & ~new_n5033_;
  assign new_n5035_ = \encrypt<0>  & ~new_n5034_;
  assign new_n5036_ = ~new_n5027_ & ~new_n5035_;
  assign new_n5037_ = ~\start<0>  & ~new_n5036_;
  assign n1840 = new_n5023_ | new_n5037_;
  assign new_n5039_ = \key<109>  & ~\encrypt<0> ;
  assign new_n5040_ = \key<101>  & \encrypt<0> ;
  assign new_n5041_ = ~new_n5039_ & ~new_n5040_;
  assign new_n5042_ = \start<0>  & ~new_n5041_;
  assign new_n5043_ = ~new_n1185_1_ & ~new_n2800_;
  assign new_n5044_ = new_n1185_1_ & ~new_n2802_;
  assign new_n5045_ = ~new_n5043_ & ~new_n5044_;
  assign new_n5046_ = ~\encrypt<0>  & ~new_n5045_;
  assign new_n5047_ = ~\C<38>  & ~new_n1189_;
  assign new_n5048_ = \C<38>  & new_n1189_;
  assign new_n5049_ = ~new_n5047_ & ~new_n5048_;
  assign new_n5050_ = \D<38>  & ~new_n5049_;
  assign new_n5051_ = \C<38>  & ~new_n1189_;
  assign new_n5052_ = ~\D<38>  & new_n5051_;
  assign new_n5053_ = ~new_n5050_ & ~new_n5052_;
  assign new_n5054_ = \encrypt<0>  & ~new_n5053_;
  assign new_n5055_ = ~new_n5046_ & ~new_n5054_;
  assign new_n5056_ = ~\start<0>  & ~new_n5055_;
  assign n1845 = new_n5042_ | new_n5056_;
  assign new_n5058_ = \key<117>  & ~\encrypt<0> ;
  assign new_n5059_ = \key<109>  & \encrypt<0> ;
  assign new_n5060_ = ~new_n5058_ & ~new_n5059_;
  assign new_n5061_ = \start<0>  & ~new_n5060_;
  assign new_n5062_ = ~new_n1185_1_ & ~new_n2822_;
  assign new_n5063_ = new_n1185_1_ & ~new_n2824_;
  assign new_n5064_ = ~new_n5062_ & ~new_n5063_;
  assign new_n5065_ = ~\encrypt<0>  & ~new_n5064_;
  assign new_n5066_ = ~\C<37>  & ~new_n1189_;
  assign new_n5067_ = \C<37>  & new_n1189_;
  assign new_n5068_ = ~new_n5066_ & ~new_n5067_;
  assign new_n5069_ = \D<37>  & ~new_n5068_;
  assign new_n5070_ = \C<37>  & ~new_n1189_;
  assign new_n5071_ = ~\D<37>  & new_n5070_;
  assign new_n5072_ = ~new_n5069_ & ~new_n5071_;
  assign new_n5073_ = \encrypt<0>  & ~new_n5072_;
  assign new_n5074_ = ~new_n5065_ & ~new_n5073_;
  assign new_n5075_ = ~\start<0>  & ~new_n5074_;
  assign n1850 = new_n5061_ | new_n5075_;
  assign new_n5077_ = \key<125>  & ~\encrypt<0> ;
  assign new_n5078_ = \key<117>  & \encrypt<0> ;
  assign new_n5079_ = ~new_n5077_ & ~new_n5078_;
  assign new_n5080_ = \start<0>  & ~new_n5079_;
  assign new_n5081_ = ~new_n1185_1_ & ~new_n2844_;
  assign new_n5082_ = new_n1185_1_ & ~new_n2846_;
  assign new_n5083_ = ~new_n5081_ & ~new_n5082_;
  assign new_n5084_ = ~\encrypt<0>  & ~new_n5083_;
  assign new_n5085_ = ~\C<36>  & ~new_n1189_;
  assign new_n5086_ = \C<36>  & new_n1189_;
  assign new_n5087_ = ~new_n5085_ & ~new_n5086_;
  assign new_n5088_ = \D<36>  & ~new_n5087_;
  assign new_n5089_ = \C<36>  & ~new_n1189_;
  assign new_n5090_ = ~\D<36>  & new_n5089_;
  assign new_n5091_ = ~new_n5088_ & ~new_n5090_;
  assign new_n5092_ = \encrypt<0>  & ~new_n5091_;
  assign new_n5093_ = ~new_n5084_ & ~new_n5092_;
  assign new_n5094_ = ~\start<0>  & ~new_n5093_;
  assign n1855 = new_n5080_ | new_n5094_;
  assign new_n5096_ = \key<70>  & ~\encrypt<0> ;
  assign new_n5097_ = \key<125>  & \encrypt<0> ;
  assign new_n5098_ = ~new_n5096_ & ~new_n5097_;
  assign new_n5099_ = \start<0>  & ~new_n5098_;
  assign new_n5100_ = ~new_n1185_1_ & ~new_n2866_;
  assign new_n5101_ = new_n1185_1_ & ~new_n2868_;
  assign new_n5102_ = ~new_n5100_ & ~new_n5101_;
  assign new_n5103_ = ~\encrypt<0>  & ~new_n5102_;
  assign new_n5104_ = ~\C<35>  & ~new_n1189_;
  assign new_n5105_ = \C<35>  & new_n1189_;
  assign new_n5106_ = ~new_n5104_ & ~new_n5105_;
  assign new_n5107_ = \D<35>  & ~new_n5106_;
  assign new_n5108_ = \C<35>  & ~new_n1189_;
  assign new_n5109_ = ~\D<35>  & new_n5108_;
  assign new_n5110_ = ~new_n5107_ & ~new_n5109_;
  assign new_n5111_ = \encrypt<0>  & ~new_n5110_;
  assign new_n5112_ = ~new_n5103_ & ~new_n5111_;
  assign new_n5113_ = ~\start<0>  & ~new_n5112_;
  assign n1860 = new_n5099_ | new_n5113_;
  assign new_n5115_ = \key<78>  & ~\encrypt<0> ;
  assign new_n5116_ = \key<70>  & \encrypt<0> ;
  assign new_n5117_ = ~new_n5115_ & ~new_n5116_;
  assign new_n5118_ = \start<0>  & ~new_n5117_;
  assign new_n5119_ = ~new_n1185_1_ & ~new_n2888_;
  assign new_n5120_ = new_n1185_1_ & ~new_n2890_;
  assign new_n5121_ = ~new_n5119_ & ~new_n5120_;
  assign new_n5122_ = ~\encrypt<0>  & ~new_n5121_;
  assign new_n5123_ = ~\C<34>  & ~new_n1189_;
  assign new_n5124_ = \C<34>  & new_n1189_;
  assign new_n5125_ = ~new_n5123_ & ~new_n5124_;
  assign new_n5126_ = \D<34>  & ~new_n5125_;
  assign new_n5127_ = \C<34>  & ~new_n1189_;
  assign new_n5128_ = ~\D<34>  & new_n5127_;
  assign new_n5129_ = ~new_n5126_ & ~new_n5128_;
  assign new_n5130_ = \encrypt<0>  & ~new_n5129_;
  assign new_n5131_ = ~new_n5122_ & ~new_n5130_;
  assign new_n5132_ = ~\start<0>  & ~new_n5131_;
  assign n1865 = new_n5118_ | new_n5132_;
  assign new_n5134_ = \key<86>  & ~\encrypt<0> ;
  assign new_n5135_ = \key<78>  & \encrypt<0> ;
  assign new_n5136_ = ~new_n5134_ & ~new_n5135_;
  assign new_n5137_ = \start<0>  & ~new_n5136_;
  assign new_n5138_ = ~new_n1185_1_ & ~new_n2910_;
  assign new_n5139_ = new_n1185_1_ & ~new_n2912_;
  assign new_n5140_ = ~new_n5138_ & ~new_n5139_;
  assign new_n5141_ = ~\encrypt<0>  & ~new_n5140_;
  assign new_n5142_ = ~\C<33>  & ~new_n1189_;
  assign new_n5143_ = \C<33>  & new_n1189_;
  assign new_n5144_ = ~new_n5142_ & ~new_n5143_;
  assign new_n5145_ = \D<33>  & ~new_n5144_;
  assign new_n5146_ = \C<33>  & ~new_n1189_;
  assign new_n5147_ = ~\D<33>  & new_n5146_;
  assign new_n5148_ = ~new_n5145_ & ~new_n5147_;
  assign new_n5149_ = \encrypt<0>  & ~new_n5148_;
  assign new_n5150_ = ~new_n5141_ & ~new_n5149_;
  assign new_n5151_ = ~\start<0>  & ~new_n5150_;
  assign n1870 = new_n5137_ | new_n5151_;
  assign new_n5153_ = \key<94>  & ~\encrypt<0> ;
  assign new_n5154_ = \key<86>  & \encrypt<0> ;
  assign new_n5155_ = ~new_n5153_ & ~new_n5154_;
  assign new_n5156_ = \start<0>  & ~new_n5155_;
  assign new_n5157_ = ~new_n1185_1_ & ~new_n2932_;
  assign new_n5158_ = new_n1185_1_ & ~new_n2934_;
  assign new_n5159_ = ~new_n5157_ & ~new_n5158_;
  assign new_n5160_ = ~\encrypt<0>  & ~new_n5159_;
  assign new_n5161_ = ~\C<32>  & ~new_n1189_;
  assign new_n5162_ = \C<32>  & new_n1189_;
  assign new_n5163_ = ~new_n5161_ & ~new_n5162_;
  assign new_n5164_ = \D<32>  & ~new_n5163_;
  assign new_n5165_ = \C<32>  & ~new_n1189_;
  assign new_n5166_ = ~\D<32>  & new_n5165_;
  assign new_n5167_ = ~new_n5164_ & ~new_n5166_;
  assign new_n5168_ = \encrypt<0>  & ~new_n5167_;
  assign new_n5169_ = ~new_n5160_ & ~new_n5168_;
  assign new_n5170_ = ~\start<0>  & ~new_n5169_;
  assign n1875 = new_n5156_ | new_n5170_;
  assign new_n5172_ = \key<102>  & ~\encrypt<0> ;
  assign new_n5173_ = \key<94>  & \encrypt<0> ;
  assign new_n5174_ = ~new_n5172_ & ~new_n5173_;
  assign new_n5175_ = \start<0>  & ~new_n5174_;
  assign new_n5176_ = ~new_n1185_1_ & ~new_n2954_;
  assign new_n5177_ = new_n1185_1_ & ~new_n2956_;
  assign new_n5178_ = ~new_n5176_ & ~new_n5177_;
  assign new_n5179_ = ~\encrypt<0>  & ~new_n5178_;
  assign new_n5180_ = ~\C<31>  & ~new_n1189_;
  assign new_n5181_ = \C<31>  & new_n1189_;
  assign new_n5182_ = ~new_n5180_ & ~new_n5181_;
  assign new_n5183_ = \D<31>  & ~new_n5182_;
  assign new_n5184_ = \C<31>  & ~new_n1189_;
  assign new_n5185_ = ~\D<31>  & new_n5184_;
  assign new_n5186_ = ~new_n5183_ & ~new_n5185_;
  assign new_n5187_ = \encrypt<0>  & ~new_n5186_;
  assign new_n5188_ = ~new_n5179_ & ~new_n5187_;
  assign new_n5189_ = ~\start<0>  & ~new_n5188_;
  assign n1880 = new_n5175_ | new_n5189_;
  assign new_n5191_ = \key<110>  & ~\encrypt<0> ;
  assign new_n5192_ = \key<102>  & \encrypt<0> ;
  assign new_n5193_ = ~new_n5191_ & ~new_n5192_;
  assign new_n5194_ = \start<0>  & ~new_n5193_;
  assign new_n5195_ = ~new_n1185_1_ & ~new_n2976_;
  assign new_n5196_ = new_n1185_1_ & ~new_n2978_;
  assign new_n5197_ = ~new_n5195_ & ~new_n5196_;
  assign new_n5198_ = ~\encrypt<0>  & ~new_n5197_;
  assign new_n5199_ = ~\C<30>  & ~new_n1189_;
  assign new_n5200_ = \C<30>  & new_n1189_;
  assign new_n5201_ = ~new_n5199_ & ~new_n5200_;
  assign new_n5202_ = \D<30>  & ~new_n5201_;
  assign new_n5203_ = \C<30>  & ~new_n1189_;
  assign new_n5204_ = ~\D<30>  & new_n5203_;
  assign new_n5205_ = ~new_n5202_ & ~new_n5204_;
  assign new_n5206_ = \encrypt<0>  & ~new_n5205_;
  assign new_n5207_ = ~new_n5198_ & ~new_n5206_;
  assign new_n5208_ = ~\start<0>  & ~new_n5207_;
  assign n1885 = new_n5194_ | new_n5208_;
  assign new_n5210_ = \key<118>  & ~\encrypt<0> ;
  assign new_n5211_ = \key<110>  & \encrypt<0> ;
  assign new_n5212_ = ~new_n5210_ & ~new_n5211_;
  assign new_n5213_ = \start<0>  & ~new_n5212_;
  assign new_n5214_ = ~new_n1185_1_ & ~new_n2998_;
  assign new_n5215_ = new_n1185_1_ & ~new_n3000_;
  assign new_n5216_ = ~new_n5214_ & ~new_n5215_;
  assign new_n5217_ = ~\encrypt<0>  & ~new_n5216_;
  assign new_n5218_ = ~\C<29>  & ~new_n1189_;
  assign new_n5219_ = \C<29>  & new_n1189_;
  assign new_n5220_ = ~new_n5218_ & ~new_n5219_;
  assign new_n5221_ = \D<29>  & ~new_n5220_;
  assign new_n5222_ = \C<29>  & ~new_n1189_;
  assign new_n5223_ = ~\D<29>  & new_n5222_;
  assign new_n5224_ = ~new_n5221_ & ~new_n5223_;
  assign new_n5225_ = \encrypt<0>  & ~new_n5224_;
  assign new_n5226_ = ~new_n5217_ & ~new_n5225_;
  assign new_n5227_ = ~\start<0>  & ~new_n5226_;
  assign n1890 = new_n5213_ | new_n5227_;
  assign new_n5229_ = \key<126>  & ~\encrypt<0> ;
  assign new_n5230_ = \key<118>  & \encrypt<0> ;
  assign new_n5231_ = ~new_n5229_ & ~new_n5230_;
  assign new_n5232_ = \start<0>  & ~new_n5231_;
  assign new_n5233_ = ~new_n1185_1_ & ~new_n3020_;
  assign new_n5234_ = new_n1185_1_ & ~new_n3022_;
  assign new_n5235_ = ~new_n5233_ & ~new_n5234_;
  assign new_n5236_ = ~\encrypt<0>  & ~new_n5235_;
  assign new_n5237_ = ~\C<28>  & ~new_n1189_;
  assign new_n5238_ = \C<28>  & new_n1189_;
  assign new_n5239_ = ~new_n5237_ & ~new_n5238_;
  assign new_n5240_ = \D<28>  & ~new_n5239_;
  assign new_n5241_ = \C<28>  & ~new_n1189_;
  assign new_n5242_ = ~\D<28>  & new_n5241_;
  assign new_n5243_ = ~new_n5240_ & ~new_n5242_;
  assign new_n5244_ = \encrypt<0>  & ~new_n5243_;
  assign new_n5245_ = ~new_n5236_ & ~new_n5244_;
  assign new_n5246_ = ~\start<0>  & ~new_n5245_;
  assign n1895 = new_n5232_ | new_n5246_;
  assign new_n5248_ = \key<3>  & ~\encrypt<0> ;
  assign new_n5249_ = \key<126>  & \encrypt<0> ;
  assign new_n5250_ = ~new_n5248_ & ~new_n5249_;
  assign new_n5251_ = \start<0>  & ~new_n5250_;
  assign new_n5252_ = ~new_n1185_1_ & ~new_n3042_;
  assign new_n5253_ = new_n1185_1_ & ~new_n3044_;
  assign new_n5254_ = ~new_n5252_ & ~new_n5253_;
  assign new_n5255_ = ~\encrypt<0>  & ~new_n5254_;
  assign new_n5256_ = ~\C<27>  & ~new_n1189_;
  assign new_n5257_ = \C<27>  & new_n1189_;
  assign new_n5258_ = ~new_n5256_ & ~new_n5257_;
  assign new_n5259_ = \D<27>  & ~new_n5258_;
  assign new_n5260_ = \C<27>  & ~new_n1189_;
  assign new_n5261_ = ~\D<27>  & new_n5260_;
  assign new_n5262_ = ~new_n5259_ & ~new_n5261_;
  assign new_n5263_ = \encrypt<0>  & ~new_n5262_;
  assign new_n5264_ = ~new_n5255_ & ~new_n5263_;
  assign new_n5265_ = ~\start<0>  & ~new_n5264_;
  assign n1900 = new_n5251_ | new_n5265_;
  assign new_n5267_ = \key<11>  & ~\encrypt<0> ;
  assign new_n5268_ = \key<3>  & \encrypt<0> ;
  assign new_n5269_ = ~new_n5267_ & ~new_n5268_;
  assign new_n5270_ = \start<0>  & ~new_n5269_;
  assign new_n5271_ = ~new_n1185_1_ & ~new_n3064_;
  assign new_n5272_ = new_n1185_1_ & ~new_n3066_;
  assign new_n5273_ = ~new_n5271_ & ~new_n5272_;
  assign new_n5274_ = ~\encrypt<0>  & ~new_n5273_;
  assign new_n5275_ = ~\C<26>  & ~new_n1189_;
  assign new_n5276_ = \C<26>  & new_n1189_;
  assign new_n5277_ = ~new_n5275_ & ~new_n5276_;
  assign new_n5278_ = \D<26>  & ~new_n5277_;
  assign new_n5279_ = \C<26>  & ~new_n1189_;
  assign new_n5280_ = ~\D<26>  & new_n5279_;
  assign new_n5281_ = ~new_n5278_ & ~new_n5280_;
  assign new_n5282_ = \encrypt<0>  & ~new_n5281_;
  assign new_n5283_ = ~new_n5274_ & ~new_n5282_;
  assign new_n5284_ = ~\start<0>  & ~new_n5283_;
  assign n1905 = new_n5270_ | new_n5284_;
  assign new_n5286_ = \key<19>  & ~\encrypt<0> ;
  assign new_n5287_ = \key<11>  & \encrypt<0> ;
  assign new_n5288_ = ~new_n5286_ & ~new_n5287_;
  assign new_n5289_ = \start<0>  & ~new_n5288_;
  assign new_n5290_ = ~new_n1185_1_ & ~new_n3086_;
  assign new_n5291_ = new_n1185_1_ & ~new_n3088_;
  assign new_n5292_ = ~new_n5290_ & ~new_n5291_;
  assign new_n5293_ = ~\encrypt<0>  & ~new_n5292_;
  assign new_n5294_ = ~\C<25>  & ~new_n1189_;
  assign new_n5295_ = \C<25>  & new_n1189_;
  assign new_n5296_ = ~new_n5294_ & ~new_n5295_;
  assign new_n5297_ = \D<25>  & ~new_n5296_;
  assign new_n5298_ = \C<25>  & ~new_n1189_;
  assign new_n5299_ = ~\D<25>  & new_n5298_;
  assign new_n5300_ = ~new_n5297_ & ~new_n5299_;
  assign new_n5301_ = \encrypt<0>  & ~new_n5300_;
  assign new_n5302_ = ~new_n5293_ & ~new_n5301_;
  assign new_n5303_ = ~\start<0>  & ~new_n5302_;
  assign n1910 = new_n5289_ | new_n5303_;
  assign new_n5305_ = \key<27>  & ~\encrypt<0> ;
  assign new_n5306_ = \key<19>  & \encrypt<0> ;
  assign new_n5307_ = ~new_n5305_ & ~new_n5306_;
  assign new_n5308_ = \start<0>  & ~new_n5307_;
  assign new_n5309_ = ~new_n1185_1_ & ~new_n3108_;
  assign new_n5310_ = new_n1185_1_ & ~new_n3110_;
  assign new_n5311_ = ~new_n5309_ & ~new_n5310_;
  assign new_n5312_ = ~\encrypt<0>  & ~new_n5311_;
  assign new_n5313_ = ~\C<24>  & ~new_n1189_;
  assign new_n5314_ = \C<24>  & new_n1189_;
  assign new_n5315_ = ~new_n5313_ & ~new_n5314_;
  assign new_n5316_ = \D<24>  & ~new_n5315_;
  assign new_n5317_ = \C<24>  & ~new_n1189_;
  assign new_n5318_ = ~\D<24>  & new_n5317_;
  assign new_n5319_ = ~new_n5316_ & ~new_n5318_;
  assign new_n5320_ = \encrypt<0>  & ~new_n5319_;
  assign new_n5321_ = ~new_n5312_ & ~new_n5320_;
  assign new_n5322_ = ~\start<0>  & ~new_n5321_;
  assign n1915 = new_n5308_ | new_n5322_;
  assign new_n5324_ = \key<4>  & ~\encrypt<0> ;
  assign new_n5325_ = \key<27>  & \encrypt<0> ;
  assign new_n5326_ = ~new_n5324_ & ~new_n5325_;
  assign new_n5327_ = \start<0>  & ~new_n5326_;
  assign new_n5328_ = ~new_n1185_1_ & ~new_n3130_;
  assign new_n5329_ = new_n1185_1_ & ~new_n3132_;
  assign new_n5330_ = ~new_n5328_ & ~new_n5329_;
  assign new_n5331_ = ~\encrypt<0>  & ~new_n5330_;
  assign new_n5332_ = ~\C<23>  & ~new_n1189_;
  assign new_n5333_ = \C<23>  & new_n1189_;
  assign new_n5334_ = ~new_n5332_ & ~new_n5333_;
  assign new_n5335_ = \D<23>  & ~new_n5334_;
  assign new_n5336_ = \C<23>  & ~new_n1189_;
  assign new_n5337_ = ~\D<23>  & new_n5336_;
  assign new_n5338_ = ~new_n5335_ & ~new_n5337_;
  assign new_n5339_ = \encrypt<0>  & ~new_n5338_;
  assign new_n5340_ = ~new_n5331_ & ~new_n5339_;
  assign new_n5341_ = ~\start<0>  & ~new_n5340_;
  assign n1920 = new_n5327_ | new_n5341_;
  assign new_n5343_ = \key<12>  & ~\encrypt<0> ;
  assign new_n5344_ = \key<4>  & \encrypt<0> ;
  assign new_n5345_ = ~new_n5343_ & ~new_n5344_;
  assign new_n5346_ = \start<0>  & ~new_n5345_;
  assign new_n5347_ = ~new_n1185_1_ & ~new_n3152_;
  assign new_n5348_ = new_n1185_1_ & ~new_n3154_;
  assign new_n5349_ = ~new_n5347_ & ~new_n5348_;
  assign new_n5350_ = ~\encrypt<0>  & ~new_n5349_;
  assign new_n5351_ = ~\C<22>  & ~new_n1189_;
  assign new_n5352_ = \C<22>  & new_n1189_;
  assign new_n5353_ = ~new_n5351_ & ~new_n5352_;
  assign new_n5354_ = \D<22>  & ~new_n5353_;
  assign new_n5355_ = \C<22>  & ~new_n1189_;
  assign new_n5356_ = ~\D<22>  & new_n5355_;
  assign new_n5357_ = ~new_n5354_ & ~new_n5356_;
  assign new_n5358_ = \encrypt<0>  & ~new_n5357_;
  assign new_n5359_ = ~new_n5350_ & ~new_n5358_;
  assign new_n5360_ = ~\start<0>  & ~new_n5359_;
  assign n1925 = new_n5346_ | new_n5360_;
  assign new_n5362_ = \key<20>  & ~\encrypt<0> ;
  assign new_n5363_ = \key<12>  & \encrypt<0> ;
  assign new_n5364_ = ~new_n5362_ & ~new_n5363_;
  assign new_n5365_ = \start<0>  & ~new_n5364_;
  assign new_n5366_ = ~new_n1185_1_ & ~new_n3174_;
  assign new_n5367_ = new_n1185_1_ & ~new_n3176_;
  assign new_n5368_ = ~new_n5366_ & ~new_n5367_;
  assign new_n5369_ = ~\encrypt<0>  & ~new_n5368_;
  assign new_n5370_ = ~\C<21>  & ~new_n1189_;
  assign new_n5371_ = \C<21>  & new_n1189_;
  assign new_n5372_ = ~new_n5370_ & ~new_n5371_;
  assign new_n5373_ = \D<21>  & ~new_n5372_;
  assign new_n5374_ = \C<21>  & ~new_n1189_;
  assign new_n5375_ = ~\D<21>  & new_n5374_;
  assign new_n5376_ = ~new_n5373_ & ~new_n5375_;
  assign new_n5377_ = \encrypt<0>  & ~new_n5376_;
  assign new_n5378_ = ~new_n5369_ & ~new_n5377_;
  assign new_n5379_ = ~\start<0>  & ~new_n5378_;
  assign n1930 = new_n5365_ | new_n5379_;
  assign new_n5381_ = \key<28>  & ~\encrypt<0> ;
  assign new_n5382_ = \key<20>  & \encrypt<0> ;
  assign new_n5383_ = ~new_n5381_ & ~new_n5382_;
  assign new_n5384_ = \start<0>  & ~new_n5383_;
  assign new_n5385_ = ~new_n1185_1_ & ~new_n3196_;
  assign new_n5386_ = new_n1185_1_ & ~new_n3198_;
  assign new_n5387_ = ~new_n5385_ & ~new_n5386_;
  assign new_n5388_ = ~\encrypt<0>  & ~new_n5387_;
  assign new_n5389_ = ~\C<20>  & ~new_n1189_;
  assign new_n5390_ = \C<20>  & new_n1189_;
  assign new_n5391_ = ~new_n5389_ & ~new_n5390_;
  assign new_n5392_ = \D<20>  & ~new_n5391_;
  assign new_n5393_ = \C<20>  & ~new_n1189_;
  assign new_n5394_ = ~\D<20>  & new_n5393_;
  assign new_n5395_ = ~new_n5392_ & ~new_n5394_;
  assign new_n5396_ = \encrypt<0>  & ~new_n5395_;
  assign new_n5397_ = ~new_n5388_ & ~new_n5396_;
  assign new_n5398_ = ~\start<0>  & ~new_n5397_;
  assign n1935 = new_n5384_ | new_n5398_;
  assign new_n5400_ = \key<36>  & ~\encrypt<0> ;
  assign new_n5401_ = \key<28>  & \encrypt<0> ;
  assign new_n5402_ = ~new_n5400_ & ~new_n5401_;
  assign new_n5403_ = \start<0>  & ~new_n5402_;
  assign new_n5404_ = ~new_n1185_1_ & ~new_n3218_;
  assign new_n5405_ = new_n1185_1_ & ~new_n3220_;
  assign new_n5406_ = ~new_n5404_ & ~new_n5405_;
  assign new_n5407_ = ~\encrypt<0>  & ~new_n5406_;
  assign new_n5408_ = ~\C<19>  & ~new_n1189_;
  assign new_n5409_ = \C<19>  & new_n1189_;
  assign new_n5410_ = ~new_n5408_ & ~new_n5409_;
  assign new_n5411_ = \D<19>  & ~new_n5410_;
  assign new_n5412_ = \C<19>  & ~new_n1189_;
  assign new_n5413_ = ~\D<19>  & new_n5412_;
  assign new_n5414_ = ~new_n5411_ & ~new_n5413_;
  assign new_n5415_ = \encrypt<0>  & ~new_n5414_;
  assign new_n5416_ = ~new_n5407_ & ~new_n5415_;
  assign new_n5417_ = ~\start<0>  & ~new_n5416_;
  assign n1940 = new_n5403_ | new_n5417_;
  assign new_n5419_ = \key<36>  & \encrypt<0> ;
  assign new_n5420_ = ~new_n4887_ & ~new_n5419_;
  assign new_n5421_ = \start<0>  & ~new_n5420_;
  assign new_n5422_ = ~new_n1185_1_ & ~new_n3240_;
  assign new_n5423_ = new_n1185_1_ & ~new_n3242_;
  assign new_n5424_ = ~new_n5422_ & ~new_n5423_;
  assign new_n5425_ = ~\encrypt<0>  & ~new_n5424_;
  assign new_n5426_ = ~\C<18>  & ~new_n1189_;
  assign new_n5427_ = \C<18>  & new_n1189_;
  assign new_n5428_ = ~new_n5426_ & ~new_n5427_;
  assign new_n5429_ = \D<18>  & ~new_n5428_;
  assign new_n5430_ = \C<18>  & ~new_n1189_;
  assign new_n5431_ = ~\D<18>  & new_n5430_;
  assign new_n5432_ = ~new_n5429_ & ~new_n5431_;
  assign new_n5433_ = \encrypt<0>  & ~new_n5432_;
  assign new_n5434_ = ~new_n5425_ & ~new_n5433_;
  assign new_n5435_ = ~\start<0>  & ~new_n5434_;
  assign n1945 = new_n5421_ | new_n5435_;
  assign new_n5437_ = \key<52>  & ~\encrypt<0> ;
  assign new_n5438_ = ~new_n4907_ & ~new_n5437_;
  assign new_n5439_ = \start<0>  & ~new_n5438_;
  assign new_n5440_ = ~new_n1185_1_ & ~new_n3262_;
  assign new_n5441_ = new_n1185_1_ & ~new_n3264_;
  assign new_n5442_ = ~new_n5440_ & ~new_n5441_;
  assign new_n5443_ = ~\encrypt<0>  & ~new_n5442_;
  assign new_n5444_ = ~\C<17>  & ~new_n1189_;
  assign new_n5445_ = \C<17>  & new_n1189_;
  assign new_n5446_ = ~new_n5444_ & ~new_n5445_;
  assign new_n5447_ = \D<17>  & ~new_n5446_;
  assign new_n5448_ = \C<17>  & ~new_n1189_;
  assign new_n5449_ = ~\D<17>  & new_n5448_;
  assign new_n5450_ = ~new_n5447_ & ~new_n5449_;
  assign new_n5451_ = \encrypt<0>  & ~new_n5450_;
  assign new_n5452_ = ~new_n5443_ & ~new_n5451_;
  assign new_n5453_ = ~\start<0>  & ~new_n5452_;
  assign n1950 = new_n5439_ | new_n5453_;
  assign new_n5455_ = \key<60>  & ~\encrypt<0> ;
  assign new_n5456_ = \key<52>  & \encrypt<0> ;
  assign new_n5457_ = ~new_n5455_ & ~new_n5456_;
  assign new_n5458_ = \start<0>  & ~new_n5457_;
  assign new_n5459_ = ~new_n1185_1_ & ~new_n3284_;
  assign new_n5460_ = new_n1185_1_ & ~new_n3286_;
  assign new_n5461_ = ~new_n5459_ & ~new_n5460_;
  assign new_n5462_ = ~\encrypt<0>  & ~new_n5461_;
  assign new_n5463_ = ~\C<16>  & ~new_n1189_;
  assign new_n5464_ = \C<16>  & new_n1189_;
  assign new_n5465_ = ~new_n5463_ & ~new_n5464_;
  assign new_n5466_ = \D<16>  & ~new_n5465_;
  assign new_n5467_ = \C<16>  & ~new_n1189_;
  assign new_n5468_ = ~\D<16>  & new_n5467_;
  assign new_n5469_ = ~new_n5466_ & ~new_n5468_;
  assign new_n5470_ = \encrypt<0>  & ~new_n5469_;
  assign new_n5471_ = ~new_n5462_ & ~new_n5470_;
  assign new_n5472_ = ~\start<0>  & ~new_n5471_;
  assign n1955 = new_n5458_ | new_n5472_;
  assign new_n5474_ = \key<5>  & ~\encrypt<0> ;
  assign new_n5475_ = \key<60>  & \encrypt<0> ;
  assign new_n5476_ = ~new_n5474_ & ~new_n5475_;
  assign new_n5477_ = \start<0>  & ~new_n5476_;
  assign new_n5478_ = ~new_n1185_1_ & ~new_n3306_;
  assign new_n5479_ = new_n1185_1_ & ~new_n3308_;
  assign new_n5480_ = ~new_n5478_ & ~new_n5479_;
  assign new_n5481_ = ~\encrypt<0>  & ~new_n5480_;
  assign new_n5482_ = ~\C<15>  & ~new_n1189_;
  assign new_n5483_ = \C<15>  & new_n1189_;
  assign new_n5484_ = ~new_n5482_ & ~new_n5483_;
  assign new_n5485_ = \D<15>  & ~new_n5484_;
  assign new_n5486_ = \C<15>  & ~new_n1189_;
  assign new_n5487_ = ~\D<15>  & new_n5486_;
  assign new_n5488_ = ~new_n5485_ & ~new_n5487_;
  assign new_n5489_ = \encrypt<0>  & ~new_n5488_;
  assign new_n5490_ = ~new_n5481_ & ~new_n5489_;
  assign new_n5491_ = ~\start<0>  & ~new_n5490_;
  assign n1960 = new_n5477_ | new_n5491_;
  assign new_n5493_ = \key<13>  & ~\encrypt<0> ;
  assign new_n5494_ = \key<5>  & \encrypt<0> ;
  assign new_n5495_ = ~new_n5493_ & ~new_n5494_;
  assign new_n5496_ = \start<0>  & ~new_n5495_;
  assign new_n5497_ = ~new_n1185_1_ & ~new_n3328_;
  assign new_n5498_ = new_n1185_1_ & ~new_n3330_;
  assign new_n5499_ = ~new_n5497_ & ~new_n5498_;
  assign new_n5500_ = ~\encrypt<0>  & ~new_n5499_;
  assign new_n5501_ = ~\C<14>  & ~new_n1189_;
  assign new_n5502_ = \C<14>  & new_n1189_;
  assign new_n5503_ = ~new_n5501_ & ~new_n5502_;
  assign new_n5504_ = \D<14>  & ~new_n5503_;
  assign new_n5505_ = \C<14>  & ~new_n1189_;
  assign new_n5506_ = ~\D<14>  & new_n5505_;
  assign new_n5507_ = ~new_n5504_ & ~new_n5506_;
  assign new_n5508_ = \encrypt<0>  & ~new_n5507_;
  assign new_n5509_ = ~new_n5500_ & ~new_n5508_;
  assign new_n5510_ = ~\start<0>  & ~new_n5509_;
  assign n1965 = new_n5496_ | new_n5510_;
  assign new_n5512_ = \key<21>  & ~\encrypt<0> ;
  assign new_n5513_ = \key<13>  & \encrypt<0> ;
  assign new_n5514_ = ~new_n5512_ & ~new_n5513_;
  assign new_n5515_ = \start<0>  & ~new_n5514_;
  assign new_n5516_ = ~new_n1185_1_ & ~new_n3350_;
  assign new_n5517_ = new_n1185_1_ & ~new_n3352_;
  assign new_n5518_ = ~new_n5516_ & ~new_n5517_;
  assign new_n5519_ = ~\encrypt<0>  & ~new_n5518_;
  assign new_n5520_ = ~\C<13>  & ~new_n1189_;
  assign new_n5521_ = \C<13>  & new_n1189_;
  assign new_n5522_ = ~new_n5520_ & ~new_n5521_;
  assign new_n5523_ = \D<13>  & ~new_n5522_;
  assign new_n5524_ = \C<13>  & ~new_n1189_;
  assign new_n5525_ = ~\D<13>  & new_n5524_;
  assign new_n5526_ = ~new_n5523_ & ~new_n5525_;
  assign new_n5527_ = \encrypt<0>  & ~new_n5526_;
  assign new_n5528_ = ~new_n5519_ & ~new_n5527_;
  assign new_n5529_ = ~\start<0>  & ~new_n5528_;
  assign n1970 = new_n5515_ | new_n5529_;
  assign new_n5531_ = \key<29>  & ~\encrypt<0> ;
  assign new_n5532_ = \key<21>  & \encrypt<0> ;
  assign new_n5533_ = ~new_n5531_ & ~new_n5532_;
  assign new_n5534_ = \start<0>  & ~new_n5533_;
  assign new_n5535_ = ~new_n1185_1_ & ~new_n3372_;
  assign new_n5536_ = new_n1185_1_ & ~new_n3374_;
  assign new_n5537_ = ~new_n5535_ & ~new_n5536_;
  assign new_n5538_ = ~\encrypt<0>  & ~new_n5537_;
  assign new_n5539_ = ~\C<12>  & ~new_n1189_;
  assign new_n5540_ = \C<12>  & new_n1189_;
  assign new_n5541_ = ~new_n5539_ & ~new_n5540_;
  assign new_n5542_ = \D<12>  & ~new_n5541_;
  assign new_n5543_ = \C<12>  & ~new_n1189_;
  assign new_n5544_ = ~\D<12>  & new_n5543_;
  assign new_n5545_ = ~new_n5542_ & ~new_n5544_;
  assign new_n5546_ = \encrypt<0>  & ~new_n5545_;
  assign new_n5547_ = ~new_n5538_ & ~new_n5546_;
  assign new_n5548_ = ~\start<0>  & ~new_n5547_;
  assign n1975 = new_n5534_ | new_n5548_;
  assign new_n5550_ = \key<37>  & ~\encrypt<0> ;
  assign new_n5551_ = \key<29>  & \encrypt<0> ;
  assign new_n5552_ = ~new_n5550_ & ~new_n5551_;
  assign new_n5553_ = \start<0>  & ~new_n5552_;
  assign new_n5554_ = ~new_n1185_1_ & ~new_n3394_;
  assign new_n5555_ = new_n1185_1_ & ~new_n3396_;
  assign new_n5556_ = ~new_n5554_ & ~new_n5555_;
  assign new_n5557_ = ~\encrypt<0>  & ~new_n5556_;
  assign new_n5558_ = ~\C<11>  & ~new_n1189_;
  assign new_n5559_ = \C<11>  & new_n1189_;
  assign new_n5560_ = ~new_n5558_ & ~new_n5559_;
  assign new_n5561_ = \D<11>  & ~new_n5560_;
  assign new_n5562_ = \C<11>  & ~new_n1189_;
  assign new_n5563_ = ~\D<11>  & new_n5562_;
  assign new_n5564_ = ~new_n5561_ & ~new_n5563_;
  assign new_n5565_ = \encrypt<0>  & ~new_n5564_;
  assign new_n5566_ = ~new_n5557_ & ~new_n5565_;
  assign new_n5567_ = ~\start<0>  & ~new_n5566_;
  assign n1980 = new_n5553_ | new_n5567_;
  assign new_n5569_ = \key<45>  & ~\encrypt<0> ;
  assign new_n5570_ = \key<37>  & \encrypt<0> ;
  assign new_n5571_ = ~new_n5569_ & ~new_n5570_;
  assign new_n5572_ = \start<0>  & ~new_n5571_;
  assign new_n5573_ = ~new_n1185_1_ & ~new_n3416_;
  assign new_n5574_ = new_n1185_1_ & ~new_n3418_;
  assign new_n5575_ = ~new_n5573_ & ~new_n5574_;
  assign new_n5576_ = ~\encrypt<0>  & ~new_n5575_;
  assign new_n5577_ = ~\C<10>  & ~new_n1189_;
  assign new_n5578_ = \C<10>  & new_n1189_;
  assign new_n5579_ = ~new_n5577_ & ~new_n5578_;
  assign new_n5580_ = \D<10>  & ~new_n5579_;
  assign new_n5581_ = \C<10>  & ~new_n1189_;
  assign new_n5582_ = ~\D<10>  & new_n5581_;
  assign new_n5583_ = ~new_n5580_ & ~new_n5582_;
  assign new_n5584_ = \encrypt<0>  & ~new_n5583_;
  assign new_n5585_ = ~new_n5576_ & ~new_n5584_;
  assign new_n5586_ = ~\start<0>  & ~new_n5585_;
  assign n1985 = new_n5572_ | new_n5586_;
  assign new_n5588_ = \key<53>  & ~\encrypt<0> ;
  assign new_n5589_ = \key<45>  & \encrypt<0> ;
  assign new_n5590_ = ~new_n5588_ & ~new_n5589_;
  assign new_n5591_ = \start<0>  & ~new_n5590_;
  assign new_n5592_ = ~new_n1185_1_ & ~new_n3438_;
  assign new_n5593_ = new_n1185_1_ & ~new_n3440_;
  assign new_n5594_ = ~new_n5592_ & ~new_n5593_;
  assign new_n5595_ = ~\encrypt<0>  & ~new_n5594_;
  assign new_n5596_ = ~\C<9>  & ~new_n1189_;
  assign new_n5597_ = \C<9>  & new_n1189_;
  assign new_n5598_ = ~new_n5596_ & ~new_n5597_;
  assign new_n5599_ = \D<9>  & ~new_n5598_;
  assign new_n5600_ = \C<9>  & ~new_n1189_;
  assign new_n5601_ = ~\D<9>  & new_n5600_;
  assign new_n5602_ = ~new_n5599_ & ~new_n5601_;
  assign new_n5603_ = \encrypt<0>  & ~new_n5602_;
  assign new_n5604_ = ~new_n5595_ & ~new_n5603_;
  assign new_n5605_ = ~\start<0>  & ~new_n5604_;
  assign n1990 = new_n5591_ | new_n5605_;
  assign new_n5607_ = \key<61>  & ~\encrypt<0> ;
  assign new_n5608_ = \key<53>  & \encrypt<0> ;
  assign new_n5609_ = ~new_n5607_ & ~new_n5608_;
  assign new_n5610_ = \start<0>  & ~new_n5609_;
  assign new_n5611_ = ~new_n1185_1_ & ~new_n3460_;
  assign new_n5612_ = new_n1185_1_ & ~new_n3462_;
  assign new_n5613_ = ~new_n5611_ & ~new_n5612_;
  assign new_n5614_ = ~\encrypt<0>  & ~new_n5613_;
  assign new_n5615_ = ~\C<8>  & ~new_n1189_;
  assign new_n5616_ = \C<8>  & new_n1189_;
  assign new_n5617_ = ~new_n5615_ & ~new_n5616_;
  assign new_n5618_ = \D<8>  & ~new_n5617_;
  assign new_n5619_ = \C<8>  & ~new_n1189_;
  assign new_n5620_ = ~\D<8>  & new_n5619_;
  assign new_n5621_ = ~new_n5618_ & ~new_n5620_;
  assign new_n5622_ = \encrypt<0>  & ~new_n5621_;
  assign new_n5623_ = ~new_n5614_ & ~new_n5622_;
  assign new_n5624_ = ~\start<0>  & ~new_n5623_;
  assign n1995 = new_n5610_ | new_n5624_;
  assign new_n5626_ = \key<6>  & ~\encrypt<0> ;
  assign new_n5627_ = \key<61>  & \encrypt<0> ;
  assign new_n5628_ = ~new_n5626_ & ~new_n5627_;
  assign new_n5629_ = \start<0>  & ~new_n5628_;
  assign new_n5630_ = ~new_n1185_1_ & ~new_n3482_;
  assign new_n5631_ = new_n1185_1_ & ~new_n3484_;
  assign new_n5632_ = ~new_n5630_ & ~new_n5631_;
  assign new_n5633_ = ~\encrypt<0>  & ~new_n5632_;
  assign new_n5634_ = ~\C<7>  & ~new_n1189_;
  assign new_n5635_ = \C<7>  & new_n1189_;
  assign new_n5636_ = ~new_n5634_ & ~new_n5635_;
  assign new_n5637_ = \D<7>  & ~new_n5636_;
  assign new_n5638_ = \C<7>  & ~new_n1189_;
  assign new_n5639_ = ~\D<7>  & new_n5638_;
  assign new_n5640_ = ~new_n5637_ & ~new_n5639_;
  assign new_n5641_ = \encrypt<0>  & ~new_n5640_;
  assign new_n5642_ = ~new_n5633_ & ~new_n5641_;
  assign new_n5643_ = ~\start<0>  & ~new_n5642_;
  assign n2000 = new_n5629_ | new_n5643_;
  assign new_n5645_ = \key<14>  & ~\encrypt<0> ;
  assign new_n5646_ = \key<6>  & \encrypt<0> ;
  assign new_n5647_ = ~new_n5645_ & ~new_n5646_;
  assign new_n5648_ = \start<0>  & ~new_n5647_;
  assign new_n5649_ = ~new_n1185_1_ & ~new_n3504_;
  assign new_n5650_ = new_n1185_1_ & ~new_n3506_;
  assign new_n5651_ = ~new_n5649_ & ~new_n5650_;
  assign new_n5652_ = ~\encrypt<0>  & ~new_n5651_;
  assign new_n5653_ = ~\C<6>  & ~new_n1189_;
  assign new_n5654_ = \C<6>  & new_n1189_;
  assign new_n5655_ = ~new_n5653_ & ~new_n5654_;
  assign new_n5656_ = \D<6>  & ~new_n5655_;
  assign new_n5657_ = \C<6>  & ~new_n1189_;
  assign new_n5658_ = ~\D<6>  & new_n5657_;
  assign new_n5659_ = ~new_n5656_ & ~new_n5658_;
  assign new_n5660_ = \encrypt<0>  & ~new_n5659_;
  assign new_n5661_ = ~new_n5652_ & ~new_n5660_;
  assign new_n5662_ = ~\start<0>  & ~new_n5661_;
  assign n2005 = new_n5648_ | new_n5662_;
  assign new_n5664_ = \key<22>  & ~\encrypt<0> ;
  assign new_n5665_ = \key<14>  & \encrypt<0> ;
  assign new_n5666_ = ~new_n5664_ & ~new_n5665_;
  assign new_n5667_ = \start<0>  & ~new_n5666_;
  assign new_n5668_ = ~new_n1185_1_ & ~new_n3526_;
  assign new_n5669_ = new_n1185_1_ & ~new_n3528_;
  assign new_n5670_ = ~new_n5668_ & ~new_n5669_;
  assign new_n5671_ = ~\encrypt<0>  & ~new_n5670_;
  assign new_n5672_ = ~\C<5>  & ~new_n1189_;
  assign new_n5673_ = \C<5>  & new_n1189_;
  assign new_n5674_ = ~new_n5672_ & ~new_n5673_;
  assign new_n5675_ = \D<5>  & ~new_n5674_;
  assign new_n5676_ = \C<5>  & ~new_n1189_;
  assign new_n5677_ = ~\D<5>  & new_n5676_;
  assign new_n5678_ = ~new_n5675_ & ~new_n5677_;
  assign new_n5679_ = \encrypt<0>  & ~new_n5678_;
  assign new_n5680_ = ~new_n5671_ & ~new_n5679_;
  assign new_n5681_ = ~\start<0>  & ~new_n5680_;
  assign n2010 = new_n5667_ | new_n5681_;
  assign new_n5683_ = \key<30>  & ~\encrypt<0> ;
  assign new_n5684_ = \key<22>  & \encrypt<0> ;
  assign new_n5685_ = ~new_n5683_ & ~new_n5684_;
  assign new_n5686_ = \start<0>  & ~new_n5685_;
  assign new_n5687_ = ~new_n1185_1_ & ~new_n3548_;
  assign new_n5688_ = new_n1185_1_ & ~new_n3550_;
  assign new_n5689_ = ~new_n5687_ & ~new_n5688_;
  assign new_n5690_ = ~\encrypt<0>  & ~new_n5689_;
  assign new_n5691_ = ~\C<4>  & ~new_n1189_;
  assign new_n5692_ = \C<4>  & new_n1189_;
  assign new_n5693_ = ~new_n5691_ & ~new_n5692_;
  assign new_n5694_ = \D<4>  & ~new_n5693_;
  assign new_n5695_ = \C<4>  & ~new_n1189_;
  assign new_n5696_ = ~\D<4>  & new_n5695_;
  assign new_n5697_ = ~new_n5694_ & ~new_n5696_;
  assign new_n5698_ = \encrypt<0>  & ~new_n5697_;
  assign new_n5699_ = ~new_n5690_ & ~new_n5698_;
  assign new_n5700_ = ~\start<0>  & ~new_n5699_;
  assign n2015 = new_n5686_ | new_n5700_;
  assign new_n5702_ = \key<38>  & ~\encrypt<0> ;
  assign new_n5703_ = \key<30>  & \encrypt<0> ;
  assign new_n5704_ = ~new_n5702_ & ~new_n5703_;
  assign new_n5705_ = \start<0>  & ~new_n5704_;
  assign new_n5706_ = ~new_n1185_1_ & ~new_n3570_;
  assign new_n5707_ = new_n1185_1_ & ~new_n3572_;
  assign new_n5708_ = ~new_n5706_ & ~new_n5707_;
  assign new_n5709_ = ~\encrypt<0>  & ~new_n5708_;
  assign new_n5710_ = ~\C<3>  & ~new_n1189_;
  assign new_n5711_ = \C<3>  & new_n1189_;
  assign new_n5712_ = ~new_n5710_ & ~new_n5711_;
  assign new_n5713_ = \D<3>  & ~new_n5712_;
  assign new_n5714_ = \C<3>  & ~new_n1189_;
  assign new_n5715_ = ~\D<3>  & new_n5714_;
  assign new_n5716_ = ~new_n5713_ & ~new_n5715_;
  assign new_n5717_ = \encrypt<0>  & ~new_n5716_;
  assign new_n5718_ = ~new_n5709_ & ~new_n5717_;
  assign new_n5719_ = ~\start<0>  & ~new_n5718_;
  assign n2020 = new_n5705_ | new_n5719_;
  assign new_n5721_ = \key<46>  & ~\encrypt<0> ;
  assign new_n5722_ = \key<38>  & \encrypt<0> ;
  assign new_n5723_ = ~new_n5721_ & ~new_n5722_;
  assign new_n5724_ = \start<0>  & ~new_n5723_;
  assign new_n5725_ = ~new_n1185_1_ & ~new_n3592_;
  assign new_n5726_ = new_n1185_1_ & ~new_n3594_;
  assign new_n5727_ = ~new_n5725_ & ~new_n5726_;
  assign new_n5728_ = ~\encrypt<0>  & ~new_n5727_;
  assign new_n5729_ = ~\C<2>  & ~new_n1189_;
  assign new_n5730_ = \C<2>  & new_n1189_;
  assign new_n5731_ = ~new_n5729_ & ~new_n5730_;
  assign new_n5732_ = \D<2>  & ~new_n5731_;
  assign new_n5733_ = \C<2>  & ~new_n1189_;
  assign new_n5734_ = ~\D<2>  & new_n5733_;
  assign new_n5735_ = ~new_n5732_ & ~new_n5734_;
  assign new_n5736_ = \encrypt<0>  & ~new_n5735_;
  assign new_n5737_ = ~new_n5728_ & ~new_n5736_;
  assign new_n5738_ = ~\start<0>  & ~new_n5737_;
  assign n2025 = new_n5724_ | new_n5738_;
  assign new_n5740_ = \key<54>  & ~\encrypt<0> ;
  assign new_n5741_ = \key<46>  & \encrypt<0> ;
  assign new_n5742_ = ~new_n5740_ & ~new_n5741_;
  assign new_n5743_ = \start<0>  & ~new_n5742_;
  assign new_n5744_ = ~new_n1185_1_ & ~new_n3614_;
  assign new_n5745_ = new_n1185_1_ & ~new_n3616_;
  assign new_n5746_ = ~new_n5744_ & ~new_n5745_;
  assign new_n5747_ = ~\encrypt<0>  & ~new_n5746_;
  assign new_n5748_ = ~\C<1>  & ~new_n1189_;
  assign new_n5749_ = \C<1>  & new_n1189_;
  assign new_n5750_ = ~new_n5748_ & ~new_n5749_;
  assign new_n5751_ = \D<1>  & ~new_n5750_;
  assign new_n5752_ = \C<1>  & ~new_n1189_;
  assign new_n5753_ = ~\D<1>  & new_n5752_;
  assign new_n5754_ = ~new_n5751_ & ~new_n5753_;
  assign new_n5755_ = \encrypt<0>  & ~new_n5754_;
  assign new_n5756_ = ~new_n5747_ & ~new_n5755_;
  assign new_n5757_ = ~\start<0>  & ~new_n5756_;
  assign n2030 = new_n5743_ | new_n5757_;
  assign new_n5759_ = \key<62>  & ~\encrypt<0> ;
  assign new_n5760_ = \key<54>  & \encrypt<0> ;
  assign new_n5761_ = ~new_n5759_ & ~new_n5760_;
  assign new_n5762_ = \start<0>  & ~new_n5761_;
  assign new_n5763_ = ~new_n1185_1_ & ~new_n3636_;
  assign new_n5764_ = new_n1185_1_ & ~new_n3638_;
  assign new_n5765_ = ~new_n5763_ & ~new_n5764_;
  assign new_n5766_ = ~\encrypt<0>  & ~new_n5765_;
  assign new_n5767_ = ~\C<0>  & ~new_n1189_;
  assign new_n5768_ = \C<0>  & new_n1189_;
  assign new_n5769_ = ~new_n5767_ & ~new_n5768_;
  assign new_n5770_ = \D<0>  & ~new_n5769_;
  assign new_n5771_ = \C<0>  & ~new_n1189_;
  assign new_n5772_ = ~\D<0>  & new_n5771_;
  assign new_n5773_ = ~new_n5770_ & ~new_n5772_;
  assign new_n5774_ = \encrypt<0>  & ~new_n5773_;
  assign new_n5775_ = ~new_n5766_ & ~new_n5774_;
  assign new_n5776_ = ~\start<0>  & ~new_n5775_;
  assign n2035 = new_n5762_ | new_n5776_;
  assign \KSi<191>  = \D<87> ;
  assign \KSi<190>  = \D<84> ;
  assign \KSi<189>  = \D<91> ;
  assign \KSi<188>  = \D<105> ;
  assign \KSi<187>  = \D<87> ;
  assign \KSi<186>  = \D<101> ;
  assign \KSi<185>  = \D<108> ;
  assign \KSi<184>  = \D<89> ;
  assign \KSi<183>  = \D<111> ;
  assign \KSi<182>  = \D<94> ;
  assign \KSi<181>  = \D<104> ;
  assign \KSi<180>  = \D<99> ;
  assign \KSi<179>  = \D<103> ;
  assign \KSi<178>  = \D<88> ;
  assign \KSi<177>  = \D<100> ;
  assign \KSi<176>  = \D<106> ;
  assign \KSi<175>  = \D<95> ;
  assign \KSi<174>  = \D<85> ;
  assign \KSi<173>  = \D<110> ;
  assign \KSi<172>  = \D<102> ;
  assign \KSi<171>  = \D<92> ;
  assign \KSi<170>  = \D<86> ;
  assign \KSi<169>  = \D<107> ;
  assign \KSi<168>  = \D<104> ;
  assign \KSi<167>  = \D<59> ;
  assign \KSi<166>  = \D<56> ;
  assign \KSi<165>  = \D<63> ;
  assign \KSi<164>  = \D<77> ;
  assign \KSi<163>  = \D<69> ;
  assign \KSi<162>  = \D<73> ;
  assign \KSi<161>  = \D<80> ;
  assign \KSi<160>  = \D<61> ;
  assign \KSi<159>  = \D<83> ;
  assign \KSi<158>  = \D<66> ;
  assign \KSi<157>  = \D<76> ;
  assign \KSi<156>  = \D<71> ;
  assign \KSi<155>  = \D<75> ;
  assign \KSi<154>  = \D<60> ;
  assign \KSi<153>  = \D<70> ;
  assign \KSi<152>  = \D<78> ;
  assign \KSi<151>  = \D<67> ;
  assign \KSi<150>  = \D<57> ;
  assign \KSi<149>  = \D<82> ;
  assign \KSi<148>  = \D<74> ;
  assign \KSi<147>  = \D<64> ;
  assign \KSi<146>  = \D<58> ;
  assign \KSi<145>  = \D<79> ;
  assign \KSi<144>  = \D<68> ;
  assign \KSi<143>  = \D<31> ;
  assign \KSi<142>  = \D<28> ;
  assign \KSi<141>  = \D<35> ;
  assign \KSi<140>  = \D<49> ;
  assign \KSi<139>  = \D<31> ;
  assign \KSi<138>  = \D<45> ;
  assign \KSi<137>  = \D<52> ;
  assign \KSi<136>  = \D<33> ;
  assign \KSi<135>  = \D<55> ;
  assign \KSi<134>  = \D<38> ;
  assign \KSi<133>  = \D<48> ;
  assign \KSi<132>  = \D<43> ;
  assign \KSi<131>  = \D<47> ;
  assign \KSi<130>  = \D<32> ;
  assign \KSi<129>  = \D<44> ;
  assign \KSi<128>  = \D<50> ;
  assign \KSi<127>  = \D<39> ;
  assign \KSi<126>  = \D<29> ;
  assign \KSi<125>  = \D<54> ;
  assign \KSi<124>  = \D<46> ;
  assign \KSi<123>  = \D<36> ;
  assign \KSi<122>  = \D<30> ;
  assign \KSi<121>  = \D<51> ;
  assign \KSi<120>  = \D<40> ;
  assign \KSi<119>  = \D<3> ;
  assign \KSi<118>  = \D<0> ;
  assign \KSi<117>  = \D<7> ;
  assign \KSi<116>  = \D<21> ;
  assign \KSi<115>  = \D<13> ;
  assign \KSi<114>  = \D<17> ;
  assign \KSi<113>  = \D<24> ;
  assign \KSi<112>  = \D<5> ;
  assign \KSi<111>  = \D<27> ;
  assign \KSi<110>  = \D<10> ;
  assign \KSi<109>  = \D<20> ;
  assign \KSi<108>  = \D<15> ;
  assign \KSi<107>  = \D<19> ;
  assign \KSi<106>  = \D<4> ;
  assign \KSi<105>  = \D<16> ;
  assign \KSi<104>  = \D<22> ;
  assign \KSi<103>  = \D<11> ;
  assign \KSi<102>  = \D<1> ;
  assign \KSi<101>  = \D<26> ;
  assign \KSi<100>  = \D<18> ;
  assign \KSi<99>  = \D<8> ;
  assign \KSi<98>  = \D<2> ;
  assign \KSi<97>  = \D<23> ;
  assign \KSi<96>  = \D<12> ;
  assign \KSi<95>  = \C<85> ;
  assign \KSi<94>  = \C<96> ;
  assign \KSi<93>  = \C<103> ;
  assign \KSi<92>  = \C<110> ;
  assign \KSi<91>  = \C<90> ;
  assign \KSi<90>  = \C<109> ;
  assign \KSi<89>  = \C<91> ;
  assign \KSi<88>  = \C<109> ;
  assign \KSi<87>  = \C<87> ;
  assign \KSi<86>  = \C<95> ;
  assign \KSi<85>  = \C<102> ;
  assign \KSi<84>  = \C<106> ;
  assign \KSi<83>  = \C<93> ;
  assign \KSi<82>  = \C<104> ;
  assign \KSi<81>  = \C<89> ;
  assign \KSi<80>  = \C<98> ;
  assign \KSi<79>  = \C<111> ;
  assign \KSi<78>  = \C<86> ;
  assign \KSi<77>  = \C<88> ;
  assign \KSi<76>  = \C<84> ;
  assign \KSi<75>  = \C<107> ;
  assign \KSi<74>  = \C<94> ;
  assign \KSi<73>  = \C<100> ;
  assign \KSi<72>  = \C<97> ;
  assign \KSi<71>  = \C<57> ;
  assign \KSi<70>  = \C<68> ;
  assign \KSi<69>  = \C<75> ;
  assign \KSi<68>  = \C<82> ;
  assign \KSi<67>  = \C<62> ;
  assign \KSi<66>  = \C<71> ;
  assign \KSi<65>  = \C<63> ;
  assign \KSi<64>  = \C<81> ;
  assign \KSi<63>  = \C<59> ;
  assign \KSi<62>  = \C<67> ;
  assign \KSi<61>  = \C<74> ;
  assign \KSi<60>  = \C<78> ;
  assign \KSi<59>  = \C<65> ;
  assign \KSi<58>  = \C<76> ;
  assign \KSi<57>  = \C<61> ;
  assign \KSi<56>  = \C<70> ;
  assign \KSi<55>  = \C<83> ;
  assign \KSi<54>  = \C<58> ;
  assign \KSi<53>  = \C<60> ;
  assign \KSi<52>  = \C<56> ;
  assign \KSi<51>  = \C<79> ;
  assign \KSi<50>  = \C<66> ;
  assign \KSi<49>  = \C<72> ;
  assign \KSi<48>  = \C<69> ;
  assign \KSi<47>  = \C<29> ;
  assign \KSi<46>  = \C<40> ;
  assign \KSi<45>  = \C<47> ;
  assign \KSi<44>  = \C<54> ;
  assign \KSi<43>  = \C<34> ;
  assign \KSi<42>  = \C<43> ;
  assign \KSi<41>  = \C<35> ;
  assign \KSi<40>  = \C<53> ;
  assign \KSi<39>  = \C<31> ;
  assign \KSi<38>  = \C<39> ;
  assign \KSi<37>  = \C<46> ;
  assign \KSi<36>  = \C<50> ;
  assign \KSi<35>  = \C<37> ;
  assign \KSi<34>  = \C<48> ;
  assign \KSi<33>  = \C<33> ;
  assign \KSi<32>  = \C<42> ;
  assign \KSi<31>  = \C<55> ;
  assign \KSi<30>  = \C<30> ;
  assign \KSi<29>  = \C<32> ;
  assign \KSi<28>  = \C<28> ;
  assign \KSi<27>  = \C<51> ;
  assign \KSi<26>  = \C<38> ;
  assign \KSi<25>  = \C<44> ;
  assign \KSi<24>  = \C<41> ;
  assign \KSi<23>  = \C<1> ;
  assign \KSi<22>  = \C<12> ;
  assign \KSi<21>  = \C<19> ;
  assign \KSi<20>  = \C<26> ;
  assign \KSi<19>  = \C<6> ;
  assign \KSi<18>  = \C<15> ;
  assign \KSi<17>  = \C<7> ;
  assign \KSi<16>  = \C<25> ;
  assign \KSi<15>  = \C<3> ;
  assign \KSi<14>  = \C<11> ;
  assign \KSi<13>  = \C<18> ;
  assign \KSi<12>  = \C<22> ;
  assign \KSi<11>  = \C<9> ;
  assign \KSi<10>  = \C<20> ;
  assign \KSi<9>  = \C<5> ;
  assign \KSi<8>  = \C<14> ;
  assign \KSi<7>  = \C<27> ;
  assign \KSi<6>  = \C<2> ;
  assign \KSi<5>  = \C<4> ;
  assign \KSi<4>  = \C<0> ;
  assign \KSi<3>  = \C<23> ;
  assign \KSi<2>  = \C<10> ;
  assign \KSi<1>  = \C<16> ;
  assign \KSi<0>  = \C<13> ;
  always @ (posedge clock) begin
    \C<111>  <= n920;
    \C<110>  <= n925;
    \C<109>  <= n930;
    \C<108>  <= n935;
    \C<107>  <= n940;
    \C<106>  <= n945;
    \C<105>  <= n950;
    \C<104>  <= n955;
    \C<103>  <= n960;
    \C<102>  <= n965;
    \C<101>  <= n970;
    \C<100>  <= n975;
    \C<99>  <= n980;
    \C<98>  <= n985;
    \C<97>  <= n990;
    \C<96>  <= n995;
    \C<95>  <= n1000;
    \C<94>  <= n1005;
    \C<93>  <= n1010;
    \C<92>  <= n1015;
    \C<91>  <= n1020;
    \C<90>  <= n1025;
    \C<89>  <= n1030;
    \C<88>  <= n1035;
    \C<87>  <= n1040;
    \C<86>  <= n1045;
    \C<85>  <= n1050;
    \C<84>  <= n1055;
    \C<83>  <= n1060;
    \C<82>  <= n1065;
    \C<81>  <= n1070;
    \C<80>  <= n1075;
    \C<79>  <= n1080;
    \C<78>  <= n1085;
    \C<77>  <= n1090;
    \C<76>  <= n1095;
    \C<75>  <= n1100;
    \C<74>  <= n1105;
    \C<73>  <= n1110;
    \C<72>  <= n1115;
    \C<71>  <= n1120;
    \C<70>  <= n1125;
    \C<69>  <= n1130;
    \C<68>  <= n1135;
    \C<67>  <= n1140;
    \C<66>  <= n1145;
    \C<65>  <= n1150;
    \C<64>  <= n1155;
    \C<63>  <= n1160;
    \C<62>  <= n1165;
    \C<61>  <= n1170;
    \C<60>  <= n1175;
    \C<59>  <= n1180;
    \C<58>  <= n1185;
    \C<57>  <= n1190;
    \C<56>  <= n1195;
    \C<55>  <= n1200;
    \C<54>  <= n1205;
    \C<53>  <= n1210;
    \C<52>  <= n1215;
    \C<51>  <= n1220;
    \C<50>  <= n1225;
    \C<49>  <= n1230;
    \C<48>  <= n1235;
    \C<47>  <= n1240;
    \C<46>  <= n1245;
    \C<45>  <= n1250;
    \C<44>  <= n1255;
    \C<43>  <= n1260;
    \C<42>  <= n1265;
    \C<41>  <= n1270;
    \C<40>  <= n1275;
    \C<39>  <= n1280;
    \C<38>  <= n1285;
    \C<37>  <= n1290;
    \C<36>  <= n1295;
    \C<35>  <= n1300;
    \C<34>  <= n1305;
    \C<33>  <= n1310;
    \C<32>  <= n1315;
    \C<31>  <= n1320;
    \C<30>  <= n1325;
    \C<29>  <= n1330;
    \C<28>  <= n1335;
    \C<27>  <= n1340;
    \C<26>  <= n1345;
    \C<25>  <= n1350;
    \C<24>  <= n1355;
    \C<23>  <= n1360;
    \C<22>  <= n1365;
    \C<21>  <= n1370;
    \C<20>  <= n1375;
    \C<19>  <= n1380;
    \C<18>  <= n1385;
    \C<17>  <= n1390;
    \C<16>  <= n1395;
    \C<15>  <= n1400;
    \C<14>  <= n1405;
    \C<13>  <= n1410;
    \C<12>  <= n1415;
    \C<11>  <= n1420;
    \C<10>  <= n1425;
    \C<9>  <= n1430;
    \C<8>  <= n1435;
    \C<7>  <= n1440;
    \C<6>  <= n1445;
    \C<5>  <= n1450;
    \C<4>  <= n1455;
    \C<3>  <= n1460;
    \C<2>  <= n1465;
    \C<1>  <= n1470;
    \C<0>  <= n1475;
    \D<111>  <= n1480;
    \D<110>  <= n1485;
    \D<109>  <= n1490;
    \D<108>  <= n1495;
    \D<107>  <= n1500;
    \D<106>  <= n1505;
    \D<105>  <= n1510;
    \D<104>  <= n1515;
    \D<103>  <= n1520;
    \D<102>  <= n1525;
    \D<101>  <= n1530;
    \D<100>  <= n1535;
    \D<99>  <= n1540;
    \D<98>  <= n1545;
    \D<97>  <= n1550;
    \D<96>  <= n1555;
    \D<95>  <= n1560;
    \D<94>  <= n1565;
    \D<93>  <= n1570;
    \D<92>  <= n1575;
    \D<91>  <= n1580;
    \D<90>  <= n1585;
    \D<89>  <= n1590;
    \D<88>  <= n1595;
    \D<87>  <= n1600;
    \D<86>  <= n1605;
    \D<85>  <= n1610;
    \D<84>  <= n1615;
    \D<83>  <= n1620;
    \D<82>  <= n1625;
    \D<81>  <= n1630;
    \D<80>  <= n1635;
    \D<79>  <= n1640;
    \D<78>  <= n1645;
    \D<77>  <= n1650;
    \D<76>  <= n1655;
    \D<75>  <= n1660;
    \D<74>  <= n1665;
    \D<73>  <= n1670;
    \D<72>  <= n1675;
    \D<71>  <= n1680;
    \D<70>  <= n1685;
    \D<69>  <= n1690;
    \D<68>  <= n1695;
    \D<67>  <= n1700;
    \D<66>  <= n1705;
    \D<65>  <= n1710;
    \D<64>  <= n1715;
    \D<63>  <= n1720;
    \D<62>  <= n1725;
    \D<61>  <= n1730;
    \D<60>  <= n1735;
    \D<59>  <= n1740;
    \D<58>  <= n1745;
    \D<57>  <= n1750;
    \D<56>  <= n1755;
    \D<55>  <= n1760;
    \D<54>  <= n1765;
    \D<53>  <= n1770;
    \D<52>  <= n1775;
    \D<51>  <= n1780;
    \D<50>  <= n1785;
    \D<49>  <= n1790;
    \D<48>  <= n1795;
    \D<47>  <= n1800;
    \D<46>  <= n1805;
    \D<45>  <= n1810;
    \D<44>  <= n1815;
    \D<43>  <= n1820;
    \D<42>  <= n1825;
    \D<41>  <= n1830;
    \D<40>  <= n1835;
    \D<39>  <= n1840;
    \D<38>  <= n1845;
    \D<37>  <= n1850;
    \D<36>  <= n1855;
    \D<35>  <= n1860;
    \D<34>  <= n1865;
    \D<33>  <= n1870;
    \D<32>  <= n1875;
    \D<31>  <= n1880;
    \D<30>  <= n1885;
    \D<29>  <= n1890;
    \D<28>  <= n1895;
    \D<27>  <= n1900;
    \D<26>  <= n1905;
    \D<25>  <= n1910;
    \D<24>  <= n1915;
    \D<23>  <= n1920;
    \D<22>  <= n1925;
    \D<21>  <= n1930;
    \D<20>  <= n1935;
    \D<19>  <= n1940;
    \D<18>  <= n1945;
    \D<17>  <= n1950;
    \D<16>  <= n1955;
    \D<15>  <= n1960;
    \D<14>  <= n1965;
    \D<13>  <= n1970;
    \D<12>  <= n1975;
    \D<11>  <= n1980;
    \D<10>  <= n1985;
    \D<9>  <= n1990;
    \D<8>  <= n1995;
    \D<7>  <= n2000;
    \D<6>  <= n2005;
    \D<5>  <= n2010;
    \D<4>  <= n2015;
    \D<3>  <= n2020;
    \D<2>  <= n2025;
    \D<1>  <= n2030;
    \D<0>  <= n2035;
  end
  initial begin
    \C<111>  <= 1'b0;
    \C<110>  <= 1'b0;
    \C<109>  <= 1'b0;
    \C<108>  <= 1'b0;
    \C<107>  <= 1'b0;
    \C<106>  <= 1'b0;
    \C<105>  <= 1'b0;
    \C<104>  <= 1'b0;
    \C<103>  <= 1'b0;
    \C<102>  <= 1'b0;
    \C<101>  <= 1'b0;
    \C<100>  <= 1'b0;
    \C<99>  <= 1'b0;
    \C<98>  <= 1'b0;
    \C<97>  <= 1'b0;
    \C<96>  <= 1'b0;
    \C<95>  <= 1'b0;
    \C<94>  <= 1'b0;
    \C<93>  <= 1'b0;
    \C<92>  <= 1'b0;
    \C<91>  <= 1'b0;
    \C<90>  <= 1'b0;
    \C<89>  <= 1'b0;
    \C<88>  <= 1'b0;
    \C<87>  <= 1'b0;
    \C<86>  <= 1'b0;
    \C<85>  <= 1'b0;
    \C<84>  <= 1'b0;
    \C<83>  <= 1'b0;
    \C<82>  <= 1'b0;
    \C<81>  <= 1'b0;
    \C<80>  <= 1'b0;
    \C<79>  <= 1'b0;
    \C<78>  <= 1'b0;
    \C<77>  <= 1'b0;
    \C<76>  <= 1'b0;
    \C<75>  <= 1'b0;
    \C<74>  <= 1'b0;
    \C<73>  <= 1'b0;
    \C<72>  <= 1'b0;
    \C<71>  <= 1'b0;
    \C<70>  <= 1'b0;
    \C<69>  <= 1'b0;
    \C<68>  <= 1'b0;
    \C<67>  <= 1'b0;
    \C<66>  <= 1'b0;
    \C<65>  <= 1'b0;
    \C<64>  <= 1'b0;
    \C<63>  <= 1'b0;
    \C<62>  <= 1'b0;
    \C<61>  <= 1'b0;
    \C<60>  <= 1'b0;
    \C<59>  <= 1'b0;
    \C<58>  <= 1'b0;
    \C<57>  <= 1'b0;
    \C<56>  <= 1'b0;
    \C<55>  <= 1'b0;
    \C<54>  <= 1'b0;
    \C<53>  <= 1'b0;
    \C<52>  <= 1'b0;
    \C<51>  <= 1'b0;
    \C<50>  <= 1'b0;
    \C<49>  <= 1'b0;
    \C<48>  <= 1'b0;
    \C<47>  <= 1'b0;
    \C<46>  <= 1'b0;
    \C<45>  <= 1'b0;
    \C<44>  <= 1'b0;
    \C<43>  <= 1'b0;
    \C<42>  <= 1'b0;
    \C<41>  <= 1'b0;
    \C<40>  <= 1'b0;
    \C<39>  <= 1'b0;
    \C<38>  <= 1'b0;
    \C<37>  <= 1'b0;
    \C<36>  <= 1'b0;
    \C<35>  <= 1'b0;
    \C<34>  <= 1'b0;
    \C<33>  <= 1'b0;
    \C<32>  <= 1'b0;
    \C<31>  <= 1'b0;
    \C<30>  <= 1'b0;
    \C<29>  <= 1'b0;
    \C<28>  <= 1'b0;
    \C<27>  <= 1'b0;
    \C<26>  <= 1'b0;
    \C<25>  <= 1'b0;
    \C<24>  <= 1'b0;
    \C<23>  <= 1'b0;
    \C<22>  <= 1'b0;
    \C<21>  <= 1'b0;
    \C<20>  <= 1'b0;
    \C<19>  <= 1'b0;
    \C<18>  <= 1'b0;
    \C<17>  <= 1'b0;
    \C<16>  <= 1'b0;
    \C<15>  <= 1'b0;
    \C<14>  <= 1'b0;
    \C<13>  <= 1'b0;
    \C<12>  <= 1'b0;
    \C<11>  <= 1'b0;
    \C<10>  <= 1'b0;
    \C<9>  <= 1'b0;
    \C<8>  <= 1'b0;
    \C<7>  <= 1'b0;
    \C<6>  <= 1'b0;
    \C<5>  <= 1'b0;
    \C<4>  <= 1'b0;
    \C<3>  <= 1'b0;
    \C<2>  <= 1'b0;
    \C<1>  <= 1'b0;
    \C<0>  <= 1'b0;
    \D<111>  <= 1'b0;
    \D<110>  <= 1'b0;
    \D<109>  <= 1'b0;
    \D<108>  <= 1'b0;
    \D<107>  <= 1'b0;
    \D<106>  <= 1'b0;
    \D<105>  <= 1'b0;
    \D<104>  <= 1'b0;
    \D<103>  <= 1'b0;
    \D<102>  <= 1'b0;
    \D<101>  <= 1'b0;
    \D<100>  <= 1'b0;
    \D<99>  <= 1'b0;
    \D<98>  <= 1'b0;
    \D<97>  <= 1'b0;
    \D<96>  <= 1'b0;
    \D<95>  <= 1'b0;
    \D<94>  <= 1'b0;
    \D<93>  <= 1'b0;
    \D<92>  <= 1'b0;
    \D<91>  <= 1'b0;
    \D<90>  <= 1'b0;
    \D<89>  <= 1'b0;
    \D<88>  <= 1'b0;
    \D<87>  <= 1'b0;
    \D<86>  <= 1'b0;
    \D<85>  <= 1'b0;
    \D<84>  <= 1'b0;
    \D<83>  <= 1'b0;
    \D<82>  <= 1'b0;
    \D<81>  <= 1'b0;
    \D<80>  <= 1'b0;
    \D<79>  <= 1'b0;
    \D<78>  <= 1'b0;
    \D<77>  <= 1'b0;
    \D<76>  <= 1'b0;
    \D<75>  <= 1'b0;
    \D<74>  <= 1'b0;
    \D<73>  <= 1'b0;
    \D<72>  <= 1'b0;
    \D<71>  <= 1'b0;
    \D<70>  <= 1'b0;
    \D<69>  <= 1'b0;
    \D<68>  <= 1'b0;
    \D<67>  <= 1'b0;
    \D<66>  <= 1'b0;
    \D<65>  <= 1'b0;
    \D<64>  <= 1'b0;
    \D<63>  <= 1'b0;
    \D<62>  <= 1'b0;
    \D<61>  <= 1'b0;
    \D<60>  <= 1'b0;
    \D<59>  <= 1'b0;
    \D<58>  <= 1'b0;
    \D<57>  <= 1'b0;
    \D<56>  <= 1'b0;
    \D<55>  <= 1'b0;
    \D<54>  <= 1'b0;
    \D<53>  <= 1'b0;
    \D<52>  <= 1'b0;
    \D<51>  <= 1'b0;
    \D<50>  <= 1'b0;
    \D<49>  <= 1'b0;
    \D<48>  <= 1'b0;
    \D<47>  <= 1'b0;
    \D<46>  <= 1'b0;
    \D<45>  <= 1'b0;
    \D<44>  <= 1'b0;
    \D<43>  <= 1'b0;
    \D<42>  <= 1'b0;
    \D<41>  <= 1'b0;
    \D<40>  <= 1'b0;
    \D<39>  <= 1'b0;
    \D<38>  <= 1'b0;
    \D<37>  <= 1'b0;
    \D<36>  <= 1'b0;
    \D<35>  <= 1'b0;
    \D<34>  <= 1'b0;
    \D<33>  <= 1'b0;
    \D<32>  <= 1'b0;
    \D<31>  <= 1'b0;
    \D<30>  <= 1'b0;
    \D<29>  <= 1'b0;
    \D<28>  <= 1'b0;
    \D<27>  <= 1'b0;
    \D<26>  <= 1'b0;
    \D<25>  <= 1'b0;
    \D<24>  <= 1'b0;
    \D<23>  <= 1'b0;
    \D<22>  <= 1'b0;
    \D<21>  <= 1'b0;
    \D<20>  <= 1'b0;
    \D<19>  <= 1'b0;
    \D<18>  <= 1'b0;
    \D<17>  <= 1'b0;
    \D<16>  <= 1'b0;
    \D<15>  <= 1'b0;
    \D<14>  <= 1'b0;
    \D<13>  <= 1'b0;
    \D<12>  <= 1'b0;
    \D<11>  <= 1'b0;
    \D<10>  <= 1'b0;
    \D<9>  <= 1'b0;
    \D<8>  <= 1'b0;
    \D<7>  <= 1'b0;
    \D<6>  <= 1'b0;
    \D<5>  <= 1'b0;
    \D<4>  <= 1'b0;
    \D<3>  <= 1'b0;
    \D<2>  <= 1'b0;
    \D<1>  <= 1'b0;
    \D<0>  <= 1'b0;
  end
endmodule

