module cht ( 
    a, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y,
    z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0,
    r0, s0, t0, u0, v0,
    w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1,
    o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2  );
  input  a, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v,
    w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0,
    p0, q0, r0, s0, t0, u0, v0;
  output w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1,
    n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2,
    f2;
  wire new_n84_, new_n85_, new_n86_, new_n87_, new_n89_, new_n90_, new_n91_,
    new_n92_, new_n94_, new_n95_, new_n96_, new_n97_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n114_, new_n115_,
    new_n116_, new_n117_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n124_, new_n125_, new_n126_, new_n127_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n154_, new_n155_, new_n156_, new_n157_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n244_, new_n245_, new_n246_, new_n247_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n259_, new_n260_, new_n261_, new_n262_, new_n264_,
    new_n265_, new_n266_, new_n267_;
  assign new_n84_ = ~f & i;
  assign new_n85_ = m & ~new_n84_;
  assign new_n86_ = f & i;
  assign new_n87_ = ~new_n85_ & ~new_n86_;
  assign w0 = ~l & ~new_n87_;
  assign new_n89_ = ~g & i;
  assign new_n90_ = n & ~new_n89_;
  assign new_n91_ = g & i;
  assign new_n92_ = ~new_n90_ & ~new_n91_;
  assign x0 = ~l & ~new_n92_;
  assign new_n94_ = ~h & i;
  assign new_n95_ = o & ~new_n94_;
  assign new_n96_ = h & i;
  assign new_n97_ = ~new_n95_ & ~new_n96_;
  assign y0 = ~l & ~new_n97_;
  assign new_n99_ = ~c & i;
  assign new_n100_ = p & ~new_n99_;
  assign new_n101_ = c & i;
  assign new_n102_ = ~new_n100_ & ~new_n101_;
  assign z0 = ~l & ~new_n102_;
  assign new_n104_ = ~d & i;
  assign new_n105_ = q & ~new_n104_;
  assign new_n106_ = d & i;
  assign new_n107_ = ~new_n105_ & ~new_n106_;
  assign a1 = ~l & ~new_n107_;
  assign new_n109_ = ~e & i;
  assign new_n110_ = r & ~new_n109_;
  assign new_n111_ = e & i;
  assign new_n112_ = ~new_n110_ & ~new_n111_;
  assign b1 = ~l & ~new_n112_;
  assign new_n114_ = ~j & ~s;
  assign new_n115_ = t & ~new_n114_;
  assign new_n116_ = ~j & s;
  assign new_n117_ = ~new_n115_ & ~new_n116_;
  assign c1 = ~l & ~new_n117_;
  assign new_n119_ = ~j & ~t;
  assign new_n120_ = u & ~new_n119_;
  assign new_n121_ = ~j & t;
  assign new_n122_ = ~new_n120_ & ~new_n121_;
  assign d1 = ~l & ~new_n122_;
  assign new_n124_ = ~j & ~u;
  assign new_n125_ = v & ~new_n124_;
  assign new_n126_ = ~j & u;
  assign new_n127_ = ~new_n125_ & ~new_n126_;
  assign e1 = ~l & ~new_n127_;
  assign new_n129_ = ~j & ~v;
  assign new_n130_ = w & ~new_n129_;
  assign new_n131_ = ~j & v;
  assign new_n132_ = ~new_n130_ & ~new_n131_;
  assign f1 = ~l & ~new_n132_;
  assign new_n134_ = ~j & ~w;
  assign new_n135_ = x & ~new_n134_;
  assign new_n136_ = ~j & w;
  assign new_n137_ = ~new_n135_ & ~new_n136_;
  assign g1 = ~l & ~new_n137_;
  assign new_n139_ = ~j & ~x;
  assign new_n140_ = y & ~new_n139_;
  assign new_n141_ = ~j & x;
  assign new_n142_ = ~new_n140_ & ~new_n141_;
  assign h1 = ~l & ~new_n142_;
  assign new_n144_ = ~j & ~y;
  assign new_n145_ = z & ~new_n144_;
  assign new_n146_ = ~j & y;
  assign new_n147_ = ~new_n145_ & ~new_n146_;
  assign i1 = ~l & ~new_n147_;
  assign new_n149_ = ~j & ~z;
  assign new_n150_ = a0 & ~new_n149_;
  assign new_n151_ = ~j & z;
  assign new_n152_ = ~new_n150_ & ~new_n151_;
  assign j1 = ~l & ~new_n152_;
  assign new_n154_ = ~j & ~a0;
  assign new_n155_ = b0 & ~new_n154_;
  assign new_n156_ = ~j & a0;
  assign new_n157_ = ~new_n155_ & ~new_n156_;
  assign k1 = ~l & ~new_n157_;
  assign new_n159_ = ~j & ~b0;
  assign new_n160_ = c0 & ~new_n159_;
  assign new_n161_ = ~j & b0;
  assign new_n162_ = ~new_n160_ & ~new_n161_;
  assign l1 = ~l & ~new_n162_;
  assign new_n164_ = ~j & ~c0;
  assign new_n165_ = d0 & ~new_n164_;
  assign new_n166_ = ~j & c0;
  assign new_n167_ = ~new_n165_ & ~new_n166_;
  assign m1 = ~l & ~new_n167_;
  assign new_n169_ = ~j & ~d0;
  assign new_n170_ = e0 & ~new_n169_;
  assign new_n171_ = ~j & d0;
  assign new_n172_ = ~new_n170_ & ~new_n171_;
  assign n1 = ~l & ~new_n172_;
  assign new_n174_ = ~j & ~e0;
  assign new_n175_ = f0 & ~new_n174_;
  assign new_n176_ = ~j & e0;
  assign new_n177_ = ~new_n175_ & ~new_n176_;
  assign o1 = ~l & ~new_n177_;
  assign new_n179_ = ~a & j;
  assign new_n180_ = f0 & ~new_n179_;
  assign new_n181_ = a & j;
  assign new_n182_ = ~new_n180_ & ~new_n181_;
  assign p1 = ~l & ~new_n182_;
  assign new_n184_ = ~k & ~g0;
  assign new_n185_ = h0 & ~new_n184_;
  assign new_n186_ = ~k & g0;
  assign new_n187_ = ~new_n185_ & ~new_n186_;
  assign q1 = ~l & ~new_n187_;
  assign new_n189_ = ~k & ~h0;
  assign new_n190_ = i0 & ~new_n189_;
  assign new_n191_ = ~k & h0;
  assign new_n192_ = ~new_n190_ & ~new_n191_;
  assign r1 = ~l & ~new_n192_;
  assign new_n194_ = ~k & ~i0;
  assign new_n195_ = j0 & ~new_n194_;
  assign new_n196_ = ~k & i0;
  assign new_n197_ = ~new_n195_ & ~new_n196_;
  assign s1 = ~l & ~new_n197_;
  assign new_n199_ = ~k & ~j0;
  assign new_n200_ = k0 & ~new_n199_;
  assign new_n201_ = ~k & j0;
  assign new_n202_ = ~new_n200_ & ~new_n201_;
  assign t1 = ~l & ~new_n202_;
  assign new_n204_ = ~k & ~k0;
  assign new_n205_ = l0 & ~new_n204_;
  assign new_n206_ = ~k & k0;
  assign new_n207_ = ~new_n205_ & ~new_n206_;
  assign u1 = ~l & ~new_n207_;
  assign new_n209_ = ~k & ~l0;
  assign new_n210_ = m0 & ~new_n209_;
  assign new_n211_ = ~k & l0;
  assign new_n212_ = ~new_n210_ & ~new_n211_;
  assign v1 = ~l & ~new_n212_;
  assign new_n214_ = ~k & ~m0;
  assign new_n215_ = n0 & ~new_n214_;
  assign new_n216_ = ~k & m0;
  assign new_n217_ = ~new_n215_ & ~new_n216_;
  assign w1 = ~l & ~new_n217_;
  assign new_n219_ = ~k & ~n0;
  assign new_n220_ = ~p & ~o0;
  assign new_n221_ = a & ~new_n220_;
  assign new_n222_ = ~p & o0;
  assign new_n223_ = ~new_n221_ & ~new_n222_;
  assign new_n224_ = ~new_n219_ & ~new_n223_;
  assign new_n225_ = ~k & n0;
  assign new_n226_ = ~new_n224_ & ~new_n225_;
  assign x1 = ~l & ~new_n226_;
  assign new_n228_ = k & ~p;
  assign new_n229_ = ~o0 & ~new_n228_;
  assign new_n230_ = p0 & ~new_n229_;
  assign new_n231_ = o0 & ~new_n228_;
  assign new_n232_ = ~new_n230_ & ~new_n231_;
  assign y1 = ~l & ~new_n232_;
  assign new_n234_ = ~p0 & ~new_n228_;
  assign new_n235_ = q0 & ~new_n234_;
  assign new_n236_ = p0 & ~new_n228_;
  assign new_n237_ = ~new_n235_ & ~new_n236_;
  assign z1 = ~l & ~new_n237_;
  assign new_n239_ = ~q0 & ~new_n228_;
  assign new_n240_ = r0 & ~new_n239_;
  assign new_n241_ = q0 & ~new_n228_;
  assign new_n242_ = ~new_n240_ & ~new_n241_;
  assign a2 = ~l & ~new_n242_;
  assign new_n244_ = ~r0 & ~new_n228_;
  assign new_n245_ = s0 & ~new_n244_;
  assign new_n246_ = r0 & ~new_n228_;
  assign new_n247_ = ~new_n245_ & ~new_n246_;
  assign b2 = ~l & ~new_n247_;
  assign new_n249_ = ~s0 & ~new_n228_;
  assign new_n250_ = t0 & ~new_n249_;
  assign new_n251_ = s0 & ~new_n228_;
  assign new_n252_ = ~new_n250_ & ~new_n251_;
  assign c2 = ~l & ~new_n252_;
  assign new_n254_ = ~t0 & ~new_n228_;
  assign new_n255_ = u0 & ~new_n254_;
  assign new_n256_ = t0 & ~new_n228_;
  assign new_n257_ = ~new_n255_ & ~new_n256_;
  assign d2 = ~l & ~new_n257_;
  assign new_n259_ = ~u0 & ~new_n228_;
  assign new_n260_ = v0 & ~new_n259_;
  assign new_n261_ = u0 & ~new_n228_;
  assign new_n262_ = ~new_n260_ & ~new_n261_;
  assign e2 = ~l & ~new_n262_;
  assign new_n264_ = ~v0 & ~new_n228_;
  assign new_n265_ = a & ~new_n264_;
  assign new_n266_ = v0 & ~new_n228_;
  assign new_n267_ = ~new_n265_ & ~new_n266_;
  assign f2 = ~l & ~new_n267_;
endmodule

