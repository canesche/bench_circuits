module top ( clock, 
    pg6, pg19, pg5, pg29, pg4, pg3, pg2, pg1, pg9, pg8, pclk, pg30, pg20,
    pg10, pg12, pg23, pg34, pg11, pg24, pg33, pg14, pg21, pg32, pg13, pg22,
    pg31, pg16, pg27, pg15, pg28, pg18, pg25, pg36, pg17, pg26, pg35,
    pg100bf, pg106bf, pg107, pg92, pg91, pg103bf, pg83, pg94, pg104bf,
    pg84, pg85, pg105bf, pg98bf, pg86bf, pg97bf, pg99bf, pg101bf, pg89bf,
    pg87bf, pg90, pg96bf, pg88bf, pg95bf  );
  input  clock;
  input  pg6, pg19, pg5, pg29, pg4, pg3, pg2, pg1, pg9, pg8, pclk, pg30,
    pg20, pg10, pg12, pg23, pg34, pg11, pg24, pg33, pg14, pg21, pg32, pg13,
    pg22, pg31, pg16, pg27, pg15, pg28, pg18, pg25, pg36, pg17, pg26, pg35;
  output pg100bf, pg106bf, pg107, pg92, pg91, pg103bf, pg83, pg94, pg104bf,
    pg84, pg85, pg105bf, pg98bf, pg86bf, pg97bf, pg99bf, pg101bf, pg89bf,
    pg87bf, pg90, pg96bf, pg88bf, pg95bf;
  reg ng73, ng69, ng70, ng71, ng72, ng65, ng66, ng67, ng68, ng64, ng74,
    ng75, ng76, ng77, ng78, ng79, ng80, ng81, ng82;
  wire new_n117_, new_n119_, new_n120_1_, new_n121_, new_n122_, new_n123_,
    new_n124_, new_n126_, new_n127_, new_n129_, new_n131_, new_n132_,
    new_n134_, new_n135_1_, new_n136_, new_n137_, new_n138_, new_n139_,
    new_n140_1_, new_n142_, new_n143_, new_n144_, new_n145_1_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_1_, new_n151_, new_n153_,
    new_n155_1_, new_n156_, new_n157_, new_n158_, new_n160_1_, new_n163_,
    new_n166_, new_n168_, new_n171_, new_n173_, new_n175_1_, new_n177_,
    new_n179_, new_n180_1_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_1_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_1_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_1_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_1_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_1_, new_n206_, new_n207_, new_n211_,
    new_n212_, new_n213_, new_n215_, new_n216_, new_n217_, new_n219_,
    new_n220_, new_n222_, new_n223_, new_n224_, new_n226_, new_n227_,
    new_n229_, new_n230_, new_n233_, new_n235_, new_n236_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n271_, new_n272_,
    new_n273_, new_n275_, n120, n125, n130, n135, n140, n145, n150, n155,
    n160, n165, n170, n175, n180, n185, n190, n195, n200, n205, n210;
  assign new_n117_ = ~pg4 & ng69;
  assign pg100bf = ~pg35 | ~new_n117_;
  assign new_n119_ = pg9 & ~pg13;
  assign new_n120_1_ = pg10 & new_n119_;
  assign new_n121_ = ~pg3 & new_n120_1_;
  assign new_n122_ = ~pg3 & ~pg11;
  assign new_n123_ = ~ng67 & ~new_n121_;
  assign new_n124_ = ~new_n122_ & new_n123_;
  assign pg89bf = ~pg25 | ~new_n124_;
  assign new_n126_ = ~pg3 & pg89bf;
  assign new_n127_ = ng78 & ~new_n126_;
  assign pg106bf = ~pg17 | ~new_n127_;
  assign new_n129_ = ~pg4 & ng79;
  assign pg107 = pg18 & new_n129_;
  assign new_n131_ = pg12 & pg13;
  assign new_n132_ = pg11 & new_n131_;
  assign pg92 = pg28 & new_n132_;
  assign new_n134_ = ~pg9 & ~pg13;
  assign new_n135_1_ = ~pg10 & new_n134_;
  assign new_n136_ = ~pg3 & new_n135_1_;
  assign new_n137_ = pg10 & new_n134_;
  assign new_n138_ = ~pg3 & new_n137_;
  assign new_n139_ = ~ng65 & ~new_n138_;
  assign new_n140_1_ = ~new_n122_ & new_n139_;
  assign pg87bf = ~pg23 | ~new_n140_1_;
  assign new_n142_ = ~pg3 & pg87bf;
  assign new_n143_ = ng76 & ~new_n142_;
  assign new_n144_ = ng64 & ~new_n143_;
  assign new_n145_1_ = ~pg2 & new_n144_;
  assign new_n146_ = ng66 & ~new_n127_;
  assign new_n147_ = ~pg2 & new_n146_;
  assign new_n148_ = ~pg10 & new_n119_;
  assign new_n149_ = ~pg3 & new_n148_;
  assign new_n150_1_ = ~new_n147_ & ~new_n149_;
  assign new_n151_ = ~new_n122_ & new_n150_1_;
  assign pg88bf = ~pg24 | ~new_n151_;
  assign new_n153_ = ~pg3 & pg88bf;
  assign n150 = ng77 & ~new_n153_;
  assign new_n155_1_ = ~new_n127_ & new_n145_1_;
  assign new_n156_ = ~n150 & new_n155_1_;
  assign new_n157_ = ~new_n136_ & ~new_n156_;
  assign new_n158_ = ~new_n122_ & new_n157_;
  assign pg86bf = ~pg22 | ~new_n158_;
  assign new_n160_1_ = ~pg3 & pg86bf;
  assign n165 = ng75 & ~new_n160_1_;
  assign pg103bf = ~pg14 | ~n165;
  assign new_n163_ = ~pg4 & ng80;
  assign pg83 = pg19 & new_n163_;
  assign pg104bf = ~pg15 | ~new_n143_;
  assign new_n166_ = ~pg4 & ng81;
  assign pg84 = pg20 & new_n166_;
  assign new_n168_ = ~pg4 & ng82;
  assign pg85 = pg21 & new_n168_;
  assign pg105bf = ~pg16 | ~n150;
  assign new_n171_ = ~pg4 & ng71;
  assign pg98bf = ~pg33 | ~new_n171_;
  assign new_n173_ = ng72 & ~pg87bf;
  assign pg97bf = ~pg32 | ~new_n173_;
  assign new_n175_1_ = ng70 & ~pg88bf;
  assign pg99bf = ~pg34 | ~new_n175_1_;
  assign new_n177_ = ng68 & ~pg89bf;
  assign pg101bf = ~pg36 | ~new_n177_;
  assign new_n179_ = ng74 & ~pg86bf;
  assign new_n180_1_ = ~pg10 & new_n179_;
  assign new_n181_ = ~pg9 & new_n180_1_;
  assign new_n182_ = ~pg4 & ng73;
  assign new_n183_ = ~pg13 & new_n181_;
  assign new_n184_ = new_n182_ & new_n183_;
  assign new_n185_1_ = ~pg10 & new_n175_1_;
  assign new_n186_ = pg9 & new_n185_1_;
  assign new_n187_ = ~pg13 & new_n186_;
  assign new_n188_ = new_n117_ & new_n187_;
  assign new_n189_ = ~new_n184_ & ~new_n188_;
  assign new_n190_1_ = pg12 & new_n189_;
  assign new_n191_ = pg10 & ~pg13;
  assign new_n192_ = new_n177_ & new_n191_;
  assign new_n193_ = pg9 & new_n192_;
  assign new_n194_ = ~pg11 & new_n117_;
  assign new_n195_1_ = new_n177_ & new_n194_;
  assign new_n196_ = new_n175_1_ & new_n195_1_;
  assign new_n197_ = new_n171_ & new_n182_;
  assign new_n198_ = new_n173_ & new_n197_;
  assign new_n199_ = new_n179_ & new_n198_;
  assign new_n200_1_ = new_n196_ & new_n199_;
  assign new_n201_ = pg10 & new_n173_;
  assign new_n202_ = ~pg9 & new_n201_;
  assign new_n203_ = ~pg13 & new_n202_;
  assign new_n204_ = new_n171_ & new_n203_;
  assign new_n205_1_ = new_n190_1_ & ~new_n193_;
  assign new_n206_ = ~new_n200_1_ & ~new_n204_;
  assign new_n207_ = new_n205_1_ & new_n206_;
  assign pg90 = pg26 & new_n207_;
  assign pg96bf = ~pg31 | ~new_n182_;
  assign pg95bf = ~pg30 | ~new_n179_;
  assign new_n211_ = ~new_n179_ & new_n182_;
  assign new_n212_ = ~pg86bf & new_n211_;
  assign new_n213_ = ~new_n179_ & ~new_n182_;
  assign n120 = ~new_n212_ & ~new_n213_;
  assign new_n215_ = new_n117_ & ~new_n175_1_;
  assign new_n216_ = ~pg88bf & new_n215_;
  assign new_n217_ = ~new_n117_ & ~new_n175_1_;
  assign n125 = ~new_n216_ & ~new_n217_;
  assign new_n219_ = new_n117_ & new_n175_1_;
  assign new_n220_ = pg88bf & new_n219_;
  assign n130 = ~new_n215_ & ~new_n220_;
  assign new_n222_ = new_n171_ & ~new_n173_;
  assign new_n223_ = ~pg87bf & new_n222_;
  assign new_n224_ = ~new_n171_ & ~new_n173_;
  assign n135 = ~new_n223_ & ~new_n224_;
  assign new_n226_ = new_n171_ & new_n173_;
  assign new_n227_ = pg87bf & new_n226_;
  assign n140 = ~new_n222_ & ~new_n227_;
  assign new_n229_ = ~new_n127_ & new_n143_;
  assign new_n230_ = ~n150 & new_n229_;
  assign n145 = ~pg2 & new_n230_;
  assign n155 = ~pg2 & new_n127_;
  assign new_n233_ = pg89bf & new_n177_;
  assign n160 = new_n177_ & ~new_n233_;
  assign new_n235_ = new_n179_ & new_n182_;
  assign new_n236_ = pg86bf & new_n235_;
  assign n170 = ~new_n211_ & ~new_n236_;
  assign new_n238_ = pg8 & n165;
  assign new_n239_ = ~new_n127_ & ~n150;
  assign new_n240_ = ~new_n143_ & new_n239_;
  assign new_n241_ = new_n179_ & new_n240_;
  assign new_n242_ = new_n182_ & new_n241_;
  assign new_n243_ = pg8 & new_n242_;
  assign new_n244_ = ~pg2 & n165;
  assign new_n245_ = ~new_n238_ & ~new_n243_;
  assign n175 = new_n244_ | ~new_n245_;
  assign new_n247_ = pg5 & new_n143_;
  assign new_n248_ = ~n165 & new_n239_;
  assign new_n249_ = new_n173_ & new_n248_;
  assign new_n250_ = new_n171_ & new_n249_;
  assign new_n251_ = pg5 & new_n250_;
  assign new_n252_ = ~pg2 & new_n143_;
  assign new_n253_ = ~new_n247_ & ~new_n251_;
  assign n180 = new_n252_ | ~new_n253_;
  assign new_n255_ = pg6 & n150;
  assign new_n256_ = ~new_n127_ & ~new_n143_;
  assign new_n257_ = ~n165 & new_n256_;
  assign new_n258_ = new_n175_1_ & new_n257_;
  assign new_n259_ = new_n117_ & new_n258_;
  assign new_n260_ = pg6 & new_n259_;
  assign new_n261_ = ~pg2 & n150;
  assign new_n262_ = ~new_n255_ & ~new_n260_;
  assign n185 = new_n261_ | ~new_n262_;
  assign new_n264_ = pg1 & new_n127_;
  assign new_n265_ = ~new_n143_ & ~n165;
  assign new_n266_ = pg1 & new_n265_;
  assign new_n267_ = new_n177_ & new_n266_;
  assign new_n268_ = ~n150 & new_n267_;
  assign new_n269_ = ~new_n264_ & ~new_n268_;
  assign n190 = n155 | ~new_n269_;
  assign new_n271_ = ~new_n143_ & n165;
  assign new_n272_ = ~pg2 & new_n271_;
  assign new_n273_ = ~new_n127_ & new_n272_;
  assign n195 = ~n150 & new_n273_;
  assign new_n275_ = ~new_n127_ & n150;
  assign n205 = ~pg2 & new_n275_;
  assign pg91 = pg27;
  assign pg94 = pg29;
  assign n200 = n145;
  assign n210 = n155;
  always @ (posedge clock) begin
    ng73 <= n120;
    ng69 <= n125;
    ng70 <= n130;
    ng71 <= n135;
    ng72 <= n140;
    ng65 <= n145;
    ng66 <= n150;
    ng67 <= n155;
    ng68 <= n160;
    ng64 <= n165;
    ng74 <= n170;
    ng75 <= n175;
    ng76 <= n180;
    ng77 <= n185;
    ng78 <= n190;
    ng79 <= n195;
    ng80 <= n200;
    ng81 <= n205;
    ng82 <= n210;
  end
endmodule

