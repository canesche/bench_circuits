module x1 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, y,
    z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0,
    r0, s0, t0, u0, v0, w0, x0, y0, z0,
    a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1,
    s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0,
    p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0;
  output a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1,
    r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2;
  wire new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n118_, new_n119_, new_n121_,
    new_n122_, new_n123_, new_n124_, new_n125_, new_n126_, new_n127_,
    new_n128_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n144_, new_n145_, new_n146_, new_n147_,
    new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n324_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n337_, new_n338_,
    new_n340_, new_n341_, new_n342_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_;
  assign a2 = f0 | r0;
  assign new_n88_ = ~a0 & ~a2;
  assign new_n89_ = ~b & ~new_n88_;
  assign new_n90_ = ~r & ~v;
  assign new_n91_ = ~j & new_n90_;
  assign new_n92_ = ~n & ~new_n91_;
  assign new_n93_ = l & ~m;
  assign new_n94_ = new_n92_ & new_n93_;
  assign new_n95_ = a0 & ~new_n94_;
  assign a1 = new_n89_ | new_n95_;
  assign new_n97_ = b & ~m;
  assign new_n98_ = ~a & new_n97_;
  assign new_n99_ = ~k & ~n;
  assign new_n100_ = l & a0;
  assign new_n101_ = new_n99_ & new_n100_;
  assign new_n102_ = new_n98_ & new_n101_;
  assign new_n103_ = ~w & g0;
  assign new_n104_ = c & new_n103_;
  assign new_n105_ = ~new_n102_ & ~new_n104_;
  assign new_n106_ = j & ~new_n105_;
  assign new_n107_ = ~k & new_n100_;
  assign new_n108_ = ~k0 & ~new_n107_;
  assign new_n109_ = v & ~new_n108_;
  assign new_n110_ = ~n & new_n109_;
  assign new_n111_ = ~m & new_n110_;
  assign new_n112_ = ~j & new_n111_;
  assign new_n113_ = b & new_n112_;
  assign new_n114_ = ~a & new_n113_;
  assign new_n115_ = o0 & t0;
  assign new_n116_ = ~new_n114_ & ~new_n115_;
  assign b1 = new_n106_ | ~new_n116_;
  assign new_n118_ = ~m & ~v;
  assign new_n119_ = ~v & ~new_n118_;
  assign c1 = b0 & ~new_n119_;
  assign new_n121_ = c0 & ~new_n119_;
  assign new_n122_ = o & p;
  assign new_n123_ = d0 & ~new_n122_;
  assign new_n124_ = ~h & new_n123_;
  assign new_n125_ = ~d & new_n124_;
  assign new_n126_ = ~a & new_n125_;
  assign new_n127_ = ~m & new_n126_;
  assign new_n128_ = ~v & new_n127_;
  assign d1 = new_n121_ | new_n128_;
  assign new_n130_ = ~e & ~u;
  assign new_n131_ = g & ~new_n130_;
  assign new_n132_ = ~e & ~w;
  assign new_n133_ = ~u & new_n132_;
  assign new_n134_ = ~new_n131_ & ~new_n133_;
  assign new_n135_ = d0 & ~new_n134_;
  assign new_n136_ = d & new_n135_;
  assign new_n137_ = ~h & e0;
  assign new_n138_ = ~a & new_n137_;
  assign new_n139_ = ~new_n136_ & ~new_n138_;
  assign new_n140_ = ~o & ~new_n139_;
  assign new_n141_ = ~m & new_n140_;
  assign new_n142_ = o0 & u0;
  assign e1 = new_n141_ | new_n142_;
  assign new_n144_ = o & q;
  assign new_n145_ = g & i;
  assign new_n146_ = ~new_n144_ & ~new_n145_;
  assign new_n147_ = q0 & new_n146_;
  assign new_n148_ = ~a & ~h;
  assign new_n149_ = o & new_n148_;
  assign new_n150_ = p & e0;
  assign new_n151_ = ~m & new_n150_;
  assign new_n152_ = new_n149_ & new_n151_;
  assign f1 = new_n147_ | new_n152_;
  assign new_n154_ = ~new_n130_ & ~new_n131_;
  assign new_n155_ = d0 & ~new_n154_;
  assign new_n156_ = p & new_n155_;
  assign new_n157_ = o & new_n156_;
  assign new_n158_ = r & s;
  assign new_n159_ = c & d;
  assign new_n160_ = p & q;
  assign new_n161_ = o & new_n160_;
  assign new_n162_ = ~new_n159_ & ~new_n161_;
  assign new_n163_ = ~new_n158_ & new_n162_;
  assign new_n164_ = p0 & new_n163_;
  assign new_n165_ = ~h & new_n164_;
  assign new_n166_ = ~g & new_n165_;
  assign new_n167_ = ~a & new_n166_;
  assign new_n168_ = ~new_n157_ & ~new_n167_;
  assign new_n169_ = ~v & ~new_n168_;
  assign new_n170_ = ~m & new_n169_;
  assign new_n171_ = ~g & ~v;
  assign new_n172_ = ~new_n161_ & ~new_n171_;
  assign new_n173_ = ~new_n158_ & new_n172_;
  assign new_n174_ = ~i & new_n173_;
  assign new_n175_ = p0 & new_n174_;
  assign new_n176_ = ~h & new_n175_;
  assign new_n177_ = ~a & new_n176_;
  assign new_n178_ = v & d0;
  assign new_n179_ = o0 & v0;
  assign new_n180_ = ~new_n178_ & ~new_n179_;
  assign new_n181_ = ~new_n177_ & new_n180_;
  assign g1 = new_n170_ | ~new_n181_;
  assign new_n183_ = ~d & d0;
  assign new_n184_ = ~s0 & ~new_n183_;
  assign new_n185_ = ~o & e0;
  assign new_n186_ = ~p0 & ~new_n185_;
  assign new_n187_ = new_n184_ & new_n186_;
  assign new_n188_ = ~w & ~new_n187_;
  assign new_n189_ = ~u & new_n188_;
  assign new_n190_ = h & new_n189_;
  assign new_n191_ = ~e & new_n190_;
  assign h1 = ~a & new_n191_;
  assign new_n193_ = ~a & ~m;
  assign new_n194_ = ~e0 & ~h0;
  assign new_n195_ = ~q0 & ~s0;
  assign new_n196_ = ~k0 & new_n195_;
  assign new_n197_ = new_n194_ & new_n196_;
  assign new_n198_ = ~new_n193_ & ~new_n197_;
  assign new_n199_ = a & ~j;
  assign new_n200_ = ~m & ~new_n199_;
  assign new_n201_ = g0 & ~new_n200_;
  assign new_n202_ = ~l0 & ~p0;
  assign new_n203_ = s & ~new_n202_;
  assign new_n204_ = r & new_n203_;
  assign new_n205_ = m & ~v;
  assign new_n206_ = ~a & ~new_n205_;
  assign new_n207_ = ~d0 & ~p0;
  assign new_n208_ = ~new_n206_ & ~new_n207_;
  assign new_n209_ = ~b0 & ~c0;
  assign new_n210_ = m & ~new_n209_;
  assign new_n211_ = w & d0;
  assign new_n212_ = d & new_n211_;
  assign new_n213_ = ~new_n210_ & ~new_n212_;
  assign new_n214_ = ~v & ~new_n213_;
  assign new_n215_ = b & r0;
  assign new_n216_ = t & i0;
  assign new_n217_ = ~j0 & ~new_n216_;
  assign new_n218_ = ~a0 & new_n217_;
  assign new_n219_ = a & ~new_n218_;
  assign new_n220_ = ~new_n215_ & ~new_n219_;
  assign new_n221_ = ~new_n214_ & new_n220_;
  assign new_n222_ = ~new_n208_ & new_n221_;
  assign new_n223_ = ~new_n204_ & new_n222_;
  assign new_n224_ = ~new_n201_ & new_n223_;
  assign k1 = new_n198_ | ~new_n224_;
  assign new_n226_ = ~d0 & ~e0;
  assign new_n227_ = h & ~new_n226_;
  assign new_n228_ = o & ~p;
  assign new_n229_ = g & ~new_n228_;
  assign new_n230_ = d & d0;
  assign new_n231_ = ~e0 & ~new_n230_;
  assign new_n232_ = ~new_n229_ & ~new_n231_;
  assign new_n233_ = ~g & new_n122_;
  assign new_n234_ = new_n183_ & new_n233_;
  assign new_n235_ = ~new_n232_ & ~new_n234_;
  assign new_n236_ = ~v & ~new_n235_;
  assign new_n237_ = ~a & new_n236_;
  assign new_n238_ = ~h & new_n237_;
  assign new_n239_ = ~h0 & ~new_n238_;
  assign new_n240_ = ~new_n227_ & new_n239_;
  assign new_n241_ = ~new_n130_ & ~new_n240_;
  assign new_n242_ = ~p0 & ~q0;
  assign new_n243_ = q & ~new_n242_;
  assign new_n244_ = p & new_n243_;
  assign new_n245_ = o & new_n244_;
  assign new_n246_ = k & a0;
  assign new_n247_ = ~f0 & ~new_n246_;
  assign new_n248_ = b & ~new_n247_;
  assign new_n249_ = w & h0;
  assign new_n250_ = ~new_n248_ & ~new_n249_;
  assign new_n251_ = ~new_n245_ & new_n250_;
  assign l1 = new_n241_ | ~new_n251_;
  assign new_n253_ = j & h0;
  assign new_n254_ = ~a & d;
  assign new_n255_ = ~m & o;
  assign new_n256_ = ~e & new_n255_;
  assign new_n257_ = new_n254_ & new_n256_;
  assign new_n258_ = ~p & ~u;
  assign new_n259_ = ~w & d0;
  assign new_n260_ = ~v & new_n259_;
  assign new_n261_ = new_n258_ & new_n260_;
  assign new_n262_ = new_n257_ & new_n261_;
  assign m1 = new_n253_ | new_n262_;
  assign new_n264_ = v & g0;
  assign new_n265_ = f & new_n264_;
  assign new_n266_ = ~e & ~m;
  assign new_n267_ = ~w & h0;
  assign new_n268_ = ~u & new_n267_;
  assign new_n269_ = new_n266_ & new_n268_;
  assign new_n270_ = ~new_n265_ & ~new_n269_;
  assign new_n271_ = ~j & ~new_n270_;
  assign new_n272_ = ~c & g0;
  assign new_n273_ = j & new_n272_;
  assign new_n274_ = ~w & s0;
  assign new_n275_ = new_n130_ & new_n274_;
  assign new_n276_ = ~new_n273_ & ~new_n275_;
  assign new_n277_ = ~h & ~new_n276_;
  assign new_n278_ = ~p & e0;
  assign new_n279_ = ~g & p;
  assign new_n280_ = ~q & q0;
  assign new_n281_ = new_n279_ & new_n280_;
  assign new_n282_ = ~new_n278_ & ~new_n281_;
  assign new_n283_ = o & ~new_n282_;
  assign new_n284_ = o0 & w0;
  assign new_n285_ = c & ~v;
  assign new_n286_ = d & p0;
  assign new_n287_ = ~g & new_n286_;
  assign new_n288_ = new_n285_ & new_n287_;
  assign new_n289_ = ~new_n284_ & ~new_n288_;
  assign new_n290_ = ~new_n283_ & new_n289_;
  assign new_n291_ = ~w & ~new_n290_;
  assign new_n292_ = ~u & new_n291_;
  assign new_n293_ = ~e & new_n292_;
  assign new_n294_ = ~new_n277_ & ~new_n293_;
  assign new_n295_ = ~m & ~new_n294_;
  assign new_n296_ = ~new_n271_ & ~new_n295_;
  assign n1 = ~a & ~new_n296_;
  assign new_n298_ = q & new_n122_;
  assign new_n299_ = ~new_n242_ & ~new_n298_;
  assign new_n300_ = g & new_n299_;
  assign new_n301_ = ~v & new_n300_;
  assign new_n302_ = ~h & i0;
  assign new_n303_ = v & p0;
  assign new_n304_ = ~new_n302_ & ~new_n303_;
  assign new_n305_ = ~new_n301_ & new_n304_;
  assign new_n306_ = i & ~new_n305_;
  assign o1 = ~a & new_n306_;
  assign new_n308_ = ~v & ~new_n108_;
  assign new_n309_ = ~s & new_n308_;
  assign new_n310_ = r & new_n309_;
  assign new_n311_ = ~m & new_n310_;
  assign new_n312_ = ~j & new_n311_;
  assign new_n313_ = b & new_n312_;
  assign new_n314_ = ~i & i0;
  assign new_n315_ = ~h & new_n314_;
  assign new_n316_ = ~j0 & ~new_n315_;
  assign new_n317_ = ~new_n313_ & new_n316_;
  assign new_n318_ = ~a & ~new_n317_;
  assign new_n319_ = a & ~h;
  assign new_n320_ = ~t & i0;
  assign new_n321_ = ~i & new_n320_;
  assign new_n322_ = new_n319_ & new_n321_;
  assign r1 = new_n318_ | new_n322_;
  assign new_n324_ = h & t;
  assign s1 = i0 & new_n324_;
  assign new_n326_ = ~f & g0;
  assign new_n327_ = n & k0;
  assign new_n328_ = ~new_n326_ & ~new_n327_;
  assign new_n329_ = v & ~new_n328_;
  assign new_n330_ = ~r & k0;
  assign new_n331_ = ~g0 & ~new_n330_;
  assign new_n332_ = ~v & ~new_n331_;
  assign new_n333_ = ~new_n329_ & ~new_n332_;
  assign new_n334_ = ~m & ~new_n333_;
  assign new_n335_ = ~j & new_n334_;
  assign v1 = ~a & new_n335_;
  assign new_n337_ = ~a0 & ~k0;
  assign new_n338_ = s & ~new_n337_;
  assign w1 = r & new_n338_;
  assign new_n340_ = ~g0 & ~a2;
  assign new_n341_ = ~j & ~new_n340_;
  assign new_n342_ = ~z & ~h0;
  assign x1 = new_n341_ | ~new_n342_;
  assign new_n344_ = ~g0 & ~r0;
  assign new_n345_ = ~f0 & new_n344_;
  assign new_n346_ = ~j & ~new_n345_;
  assign new_n347_ = ~h0 & ~new_n346_;
  assign y1 = ~z & new_n347_;
  assign z1 = c0 | d0;
  assign new_n350_ = ~e0 & ~p0;
  assign new_n351_ = p & ~new_n279_;
  assign new_n352_ = ~new_n350_ & ~new_n351_;
  assign new_n353_ = ~w & new_n352_;
  assign new_n354_ = ~v & new_n353_;
  assign new_n355_ = ~u & new_n354_;
  assign new_n356_ = o & new_n355_;
  assign new_n357_ = ~m & new_n356_;
  assign new_n358_ = ~e & new_n357_;
  assign b2 = ~a & new_n358_;
  assign new_n360_ = ~v & q0;
  assign new_n361_ = ~p0 & ~new_n360_;
  assign new_n362_ = ~new_n298_ & ~new_n361_;
  assign new_n363_ = g & new_n362_;
  assign new_n364_ = ~new_n303_ & ~new_n363_;
  assign new_n365_ = i & ~new_n364_;
  assign new_n366_ = ~a & new_n365_;
  assign new_n367_ = ~y & ~z;
  assign new_n368_ = ~h0 & ~i0;
  assign new_n369_ = new_n367_ & new_n368_;
  assign d2 = new_n366_ | ~new_n369_;
  assign new_n371_ = g & ~new_n161_;
  assign new_n372_ = ~new_n303_ & ~new_n371_;
  assign new_n373_ = ~a & i;
  assign new_n374_ = ~new_n361_ & new_n373_;
  assign new_n375_ = ~new_n372_ & new_n374_;
  assign new_n376_ = ~i0 & ~new_n375_;
  assign new_n377_ = ~h0 & new_n376_;
  assign new_n378_ = ~z & new_n377_;
  assign e2 = ~y & new_n378_;
  assign new_n380_ = ~m & r;
  assign new_n381_ = ~j & new_n380_;
  assign new_n382_ = ~z0 & ~new_n381_;
  assign new_n383_ = l & ~new_n382_;
  assign new_n384_ = b & new_n383_;
  assign new_n385_ = a0 & ~new_n384_;
  assign new_n386_ = ~new_n183_ & ~new_n185_;
  assign new_n387_ = ~new_n216_ & new_n386_;
  assign new_n388_ = ~s0 & new_n387_;
  assign new_n389_ = ~p0 & new_n388_;
  assign new_n390_ = h & ~new_n389_;
  assign new_n391_ = ~new_n385_ & ~new_n390_;
  assign new_n392_ = ~x0 & new_n391_;
  assign new_n393_ = ~r0 & new_n392_;
  assign new_n394_ = ~m0 & new_n393_;
  assign f2 = ~f0 & new_n394_;
  assign new_n396_ = ~j & ~m;
  assign new_n397_ = r & new_n396_;
  assign new_n398_ = ~z0 & ~new_n397_;
  assign new_n399_ = l & ~new_n398_;
  assign new_n400_ = b & ~new_n399_;
  assign new_n401_ = b & ~new_n400_;
  assign new_n402_ = a0 & ~new_n401_;
  assign new_n403_ = ~m0 & ~x0;
  assign new_n404_ = ~a2 & new_n403_;
  assign new_n405_ = ~new_n185_ & ~new_n216_;
  assign new_n406_ = ~p0 & new_n184_;
  assign new_n407_ = new_n405_ & new_n406_;
  assign new_n408_ = h & ~new_n407_;
  assign new_n409_ = new_n404_ & ~new_n408_;
  assign g2 = new_n402_ | ~new_n409_;
  assign new_n411_ = c & g0;
  assign new_n412_ = i & i0;
  assign new_n413_ = ~d & h;
  assign new_n414_ = d0 & ~new_n413_;
  assign new_n415_ = v & k0;
  assign new_n416_ = ~j & new_n415_;
  assign new_n417_ = ~a0 & ~new_n416_;
  assign new_n418_ = b & l;
  assign new_n419_ = ~m & ~n;
  assign new_n420_ = ~a & new_n419_;
  assign new_n421_ = new_n418_ & new_n420_;
  assign new_n422_ = ~new_n417_ & new_n421_;
  assign new_n423_ = ~new_n414_ & ~new_n422_;
  assign new_n424_ = ~new_n412_ & new_n423_;
  assign new_n425_ = ~new_n411_ & new_n424_;
  assign new_n426_ = b & v;
  assign new_n427_ = l & new_n426_;
  assign new_n428_ = ~n & ~new_n337_;
  assign new_n429_ = new_n193_ & new_n428_;
  assign new_n430_ = new_n427_ & new_n429_;
  assign new_n431_ = ~new_n414_ & ~new_n430_;
  assign new_n432_ = ~new_n412_ & new_n431_;
  assign new_n433_ = ~j & new_n432_;
  assign new_n434_ = ~new_n425_ & ~new_n433_;
  assign new_n435_ = ~h0 & ~new_n434_;
  assign new_n436_ = ~c0 & new_n435_;
  assign new_n437_ = ~b0 & new_n436_;
  assign new_n438_ = ~z & new_n437_;
  assign h2 = ~y & new_n438_;
  assign new_n440_ = ~a & new_n418_;
  assign new_n441_ = new_n415_ & new_n419_;
  assign new_n442_ = new_n440_ & new_n441_;
  assign new_n443_ = ~j & ~new_n442_;
  assign new_n444_ = g0 & ~new_n443_;
  assign new_n445_ = c & new_n444_;
  assign new_n446_ = ~j & k0;
  assign new_n447_ = ~a0 & ~new_n446_;
  assign new_n448_ = v & ~new_n447_;
  assign new_n449_ = j & a0;
  assign new_n450_ = ~new_n448_ & ~new_n449_;
  assign new_n451_ = ~n & ~new_n450_;
  assign new_n452_ = ~m & new_n451_;
  assign new_n453_ = l & new_n452_;
  assign new_n454_ = b & new_n453_;
  assign new_n455_ = ~a & new_n454_;
  assign new_n456_ = ~c0 & ~h0;
  assign new_n457_ = ~z & new_n456_;
  assign new_n458_ = ~y & ~new_n412_;
  assign new_n459_ = ~b0 & new_n458_;
  assign new_n460_ = new_n457_ & new_n459_;
  assign new_n461_ = ~new_n414_ & new_n460_;
  assign new_n462_ = ~new_n455_ & new_n461_;
  assign i2 = new_n445_ | ~new_n462_;
  assign i1 = m0;
  assign j1 = n0;
  assign p1 = y;
  assign q1 = z;
  assign t1 = x0;
  assign u1 = y0;
  assign c2 = h0;
endmodule

