module top ( 
    pv108_3_, pv109_0_, pv118_4_, pv149_4_, pv257_2_, pv268_0_, pv288_2_,
    pv108_4_, pv118_3_, pv149_5_, pv216_0_, pv257_1_, pv268_1_, pv278_0_,
    pv288_3_, pv289_0_, pv2_0_, pv108_5_, pv118_6_, pv149_6_, pv248_0_,
    pv257_4_, pv288_4_, pv118_5_, pv149_7_, pv207_0_, pv257_3_, pv258_0_,
    pv288_5_, pv60_0_, pv78_1_, pv88_2_, pv118_0_, pv172_0_, pv189_4_,
    pv215_0_, pv257_6_, pv259_0_, pv268_4_, pv78_0_, pv88_3_, pv108_0_,
    pv189_5_, pv199_4_, pv205_0_, pv213_5_, pv234_4_, pv249_0_, pv257_5_,
    pv268_5_, pv302_0_, pv108_1_, pv118_2_, pv223_5_, pv234_3_, pv268_2_,
    pv279_0_, pv288_0_, pv1_0_, pv108_2_, pv118_1_, pv171_0_, pv234_2_,
    pv257_7_, pv268_3_, pv269_0_, pv288_1_, pv4_0_, pv32_7_, pv39_0_,
    pv100_3_, pv101_0_, pv132_0_, pv189_0_, pv199_1_, pv229_1_, pv239_2_,
    pv32_6_, pv38_0_, pv65_0_, pv100_4_, pv189_1_, pv199_0_, pv229_2_,
    pv239_1_, pv245_0_, pv32_5_, pv37_0_, pv62_0_, pv100_5_, pv189_2_,
    pv199_3_, pv239_0_, pv275_0_, pv5_0_, pv32_4_, pv63_0_, pv102_0_,
    pv189_3_, pv199_2_, pv229_0_, pv32_3_, pv35_0_, pv68_0_, pv71_0_,
    pv110_0_, pv149_0_, pv246_0_, pv277_0_, pv295_0_, pv3_0_, pv32_2_,
    pv34_0_, pv69_0_, pv70_0_, pv100_0_, pv118_7_, pv149_1_, pv32_1_,
    pv33_0_, pv66_0_, pv100_1_, pv149_2_, pv169_0_, pv257_0_, pv32_0_,
    pv67_0_, pv100_2_, pv149_3_, pv169_1_, pv247_0_, pv32_10_, pv53_0_,
    pv124_1_, pv165_2_, pv242_0_, pv7_0_, pv32_11_, pv52_0_, pv124_2_,
    pv132_7_, pv134_1_, pv165_3_, pv11_0_, pv55_0_, pv132_6_, pv134_0_,
    pv165_0_, pv262_0_, pv10_0_, pv124_0_, pv132_5_, pv165_1_, pv175_0_,
    pv243_0_, pv272_0_, pv294_0_, pv57_0_, pv132_4_, pv165_6_, pv194_4_,
    pv229_5_, pv56_0_, pv91_1_, pv132_3_, pv165_7_, pv177_0_, pv194_3_,
    pv274_0_, pv292_0_, pv6_0_, pv32_9_, pv40_0_, pv59_0_, pv94_1_,
    pv132_2_, pv165_4_, pv229_3_, pv239_4_, pv244_0_, pv293_0_, pv32_8_,
    pv41_0_, pv94_0_, pv132_1_, pv165_5_, pv229_4_, pv239_3_, pv42_0_,
    pv78_5_, pv84_2_, pv183_2_, pv194_0_, pv213_2_, pv223_3_, pv234_1_,
    pv260_0_, pv291_0_, pv16_0_, pv43_0_, pv78_4_, pv84_3_, pv183_3_,
    pv213_1_, pv223_4_, pv234_0_, pv270_0_, pv44_0_, pv78_3_, pv84_4_,
    pv88_0_, pv91_0_, pv183_4_, pv194_2_, pv204_0_, pv213_4_, pv223_1_,
    pv240_0_, pv301_0_, pv45_0_, pv78_2_, pv84_5_, pv88_1_, pv183_5_,
    pv194_1_, pv213_3_, pv214_0_, pv223_2_, pv8_0_, pv13_0_, pv46_0_,
    pv124_5_, pv202_0_, pv288_6_, pv12_0_, pv223_0_, pv241_0_, pv288_7_,
    pv15_0_, pv48_0_, pv51_0_, pv84_0_, pv124_3_, pv174_0_, pv183_0_,
    pv213_0_, pv271_0_, pv280_0_, pv9_0_, pv14_0_, pv50_0_, pv84_1_,
    pv124_4_, pv183_1_, pv203_0_, pv261_0_, pv290_0_,
    pv778, pv789, pv1213_5_, pv1243_0_, pv1261, pv1371, pv1382, pv1470,
    pv1512_3_, pv1613_1_, pv1757_0_, pv1781_1_, pv1829_2_, pv1953_2_,
    pv375_0_, pv410_0_, pv508_0_, pv539, pv1213_6_, pv1260, pv1372,
    pv1440_0_, pv1758_0_, pv1781_0_, pv1829_1_, pv1953_3_, pv657, pv787,
    pv1213_7_, pv1263, pv1380, pv1759_0_, pv1829_4_, pv1953_4_, pv656,
    pv779, pv1213_8_, pv1262, pv1370, pv1829_3_, pv1953_5_, pv763,
    pv1213_9_, pv1243_4_, pv1265, pv1375, pv1386, pv1481_0_, pv1717_0_,
    pv1829_6_, pv634_0_, pv1243_3_, pv1264, pv1480_0_, pv1741_0_,
    pv1829_5_, pv321_2_, pv512, pv783, pv1243_2_, pv1256, pv1267,
    pv1281_0_, pv1373, pv1384, pv1829_8_, pv1953_0_, pv775, pv784,
    pv1243_1_, pv1257, pv1266, pv1365, pv1374, pv1459_0_, pv1829_7_,
    pv1953_1_, pv543, pv587, pv651, pv781, pv1297_1_, pv1423, pv1771_0_,
    pv1900_0_, pv1921_1_, pv393_0_, pv500_0_, pv544, pv650, pv782,
    pv1213_11_, pv1297_2_, pv1771_1_, pv1921_0_, pv1992_0_, pv541, pv620,
    pv707, pv802_0_, pv1213_10_, pv1274_0_, pv1297_3_, pv1432, pv1726_0_,
    pv1921_3_, pv1968_0_, pv1992_1_, pv357, pv423_0_, pv542, pv621, pv630,
    pv780, pv1297_4_, pv1671_0_, pv1921_2_, pv547, pv655, pv1467_0_,
    pv1629_0_, pv1863_0_, pv1896_0_, pv1921_5_, pv1953_6_, pv377, pv548,
    pv654, pv821_0_, pv1431, pv1897_0_, pv1921_4_, pv1953_7_, pv1960_1_,
    pv527, pv538, pv545, pv653, pv1829_0_, pv1898_0_, pv537, pv546,
    pv597_0_, pv652, pv801, pv1864_0_, pv1899_0_, pv572_8_, pv585_0_,
    pv1709_1_, pv1760_0_, pv373, pv572_7_, pv1439_0_, pv1709_0_, pv572_6_,
    pv1539, pv1719, pv1960_0_, pv572_5_, pv1392_0_, pv1536_0_, pv1679_0_,
    pv1833_0_, pv356, pv435_0_, pv1492_0_, pv1537, pv511_0_, pv540,
    pv609_0_, pv1426, pv1620_0_, pv1736, pv1429, pv1832, pv432, pv572_9_,
    pv1297_0_, pv1428, pv1495_0_, pv1693_0_, pv1901_0_, pv572_0_,
    pv1243_8_, pv1258, pv1243_7_, pv1259, pv1552_0_, pv1745_0_, pv1829_9_,
    pv798_0_, pv1243_6_, pv1552_1_, pv1645_0_, pv1652_0_, pv603_0_,
    pv1213_0_, pv1243_5_, pv1378, pv1387, pv572_4_, pv826_0_, pv1213_1_,
    pv1669, pv572_3_, pv591_0_, pv966, pv1213_2_, pv1709_4_, pv398_0_,
    pv572_2_, pv640_0_, pv1213_3_, pv1512_1_, pv1709_3_, pv572_1_, pv986,
    pv1213_4_, pv1243_9_, pv1451_0_, pv1512_2_, pv1613_0_, pv1709_2_  );
  input  pv108_3_, pv109_0_, pv118_4_, pv149_4_, pv257_2_, pv268_0_,
    pv288_2_, pv108_4_, pv118_3_, pv149_5_, pv216_0_, pv257_1_, pv268_1_,
    pv278_0_, pv288_3_, pv289_0_, pv2_0_, pv108_5_, pv118_6_, pv149_6_,
    pv248_0_, pv257_4_, pv288_4_, pv118_5_, pv149_7_, pv207_0_, pv257_3_,
    pv258_0_, pv288_5_, pv60_0_, pv78_1_, pv88_2_, pv118_0_, pv172_0_,
    pv189_4_, pv215_0_, pv257_6_, pv259_0_, pv268_4_, pv78_0_, pv88_3_,
    pv108_0_, pv189_5_, pv199_4_, pv205_0_, pv213_5_, pv234_4_, pv249_0_,
    pv257_5_, pv268_5_, pv302_0_, pv108_1_, pv118_2_, pv223_5_, pv234_3_,
    pv268_2_, pv279_0_, pv288_0_, pv1_0_, pv108_2_, pv118_1_, pv171_0_,
    pv234_2_, pv257_7_, pv268_3_, pv269_0_, pv288_1_, pv4_0_, pv32_7_,
    pv39_0_, pv100_3_, pv101_0_, pv132_0_, pv189_0_, pv199_1_, pv229_1_,
    pv239_2_, pv32_6_, pv38_0_, pv65_0_, pv100_4_, pv189_1_, pv199_0_,
    pv229_2_, pv239_1_, pv245_0_, pv32_5_, pv37_0_, pv62_0_, pv100_5_,
    pv189_2_, pv199_3_, pv239_0_, pv275_0_, pv5_0_, pv32_4_, pv63_0_,
    pv102_0_, pv189_3_, pv199_2_, pv229_0_, pv32_3_, pv35_0_, pv68_0_,
    pv71_0_, pv110_0_, pv149_0_, pv246_0_, pv277_0_, pv295_0_, pv3_0_,
    pv32_2_, pv34_0_, pv69_0_, pv70_0_, pv100_0_, pv118_7_, pv149_1_,
    pv32_1_, pv33_0_, pv66_0_, pv100_1_, pv149_2_, pv169_0_, pv257_0_,
    pv32_0_, pv67_0_, pv100_2_, pv149_3_, pv169_1_, pv247_0_, pv32_10_,
    pv53_0_, pv124_1_, pv165_2_, pv242_0_, pv7_0_, pv32_11_, pv52_0_,
    pv124_2_, pv132_7_, pv134_1_, pv165_3_, pv11_0_, pv55_0_, pv132_6_,
    pv134_0_, pv165_0_, pv262_0_, pv10_0_, pv124_0_, pv132_5_, pv165_1_,
    pv175_0_, pv243_0_, pv272_0_, pv294_0_, pv57_0_, pv132_4_, pv165_6_,
    pv194_4_, pv229_5_, pv56_0_, pv91_1_, pv132_3_, pv165_7_, pv177_0_,
    pv194_3_, pv274_0_, pv292_0_, pv6_0_, pv32_9_, pv40_0_, pv59_0_,
    pv94_1_, pv132_2_, pv165_4_, pv229_3_, pv239_4_, pv244_0_, pv293_0_,
    pv32_8_, pv41_0_, pv94_0_, pv132_1_, pv165_5_, pv229_4_, pv239_3_,
    pv42_0_, pv78_5_, pv84_2_, pv183_2_, pv194_0_, pv213_2_, pv223_3_,
    pv234_1_, pv260_0_, pv291_0_, pv16_0_, pv43_0_, pv78_4_, pv84_3_,
    pv183_3_, pv213_1_, pv223_4_, pv234_0_, pv270_0_, pv44_0_, pv78_3_,
    pv84_4_, pv88_0_, pv91_0_, pv183_4_, pv194_2_, pv204_0_, pv213_4_,
    pv223_1_, pv240_0_, pv301_0_, pv45_0_, pv78_2_, pv84_5_, pv88_1_,
    pv183_5_, pv194_1_, pv213_3_, pv214_0_, pv223_2_, pv8_0_, pv13_0_,
    pv46_0_, pv124_5_, pv202_0_, pv288_6_, pv12_0_, pv223_0_, pv241_0_,
    pv288_7_, pv15_0_, pv48_0_, pv51_0_, pv84_0_, pv124_3_, pv174_0_,
    pv183_0_, pv213_0_, pv271_0_, pv280_0_, pv9_0_, pv14_0_, pv50_0_,
    pv84_1_, pv124_4_, pv183_1_, pv203_0_, pv261_0_, pv290_0_;
  output pv778, pv789, pv1213_5_, pv1243_0_, pv1261, pv1371, pv1382, pv1470,
    pv1512_3_, pv1613_1_, pv1757_0_, pv1781_1_, pv1829_2_, pv1953_2_,
    pv375_0_, pv410_0_, pv508_0_, pv539, pv1213_6_, pv1260, pv1372,
    pv1440_0_, pv1758_0_, pv1781_0_, pv1829_1_, pv1953_3_, pv657, pv787,
    pv1213_7_, pv1263, pv1380, pv1759_0_, pv1829_4_, pv1953_4_, pv656,
    pv779, pv1213_8_, pv1262, pv1370, pv1829_3_, pv1953_5_, pv763,
    pv1213_9_, pv1243_4_, pv1265, pv1375, pv1386, pv1481_0_, pv1717_0_,
    pv1829_6_, pv634_0_, pv1243_3_, pv1264, pv1480_0_, pv1741_0_,
    pv1829_5_, pv321_2_, pv512, pv783, pv1243_2_, pv1256, pv1267,
    pv1281_0_, pv1373, pv1384, pv1829_8_, pv1953_0_, pv775, pv784,
    pv1243_1_, pv1257, pv1266, pv1365, pv1374, pv1459_0_, pv1829_7_,
    pv1953_1_, pv543, pv587, pv651, pv781, pv1297_1_, pv1423, pv1771_0_,
    pv1900_0_, pv1921_1_, pv393_0_, pv500_0_, pv544, pv650, pv782,
    pv1213_11_, pv1297_2_, pv1771_1_, pv1921_0_, pv1992_0_, pv541, pv620,
    pv707, pv802_0_, pv1213_10_, pv1274_0_, pv1297_3_, pv1432, pv1726_0_,
    pv1921_3_, pv1968_0_, pv1992_1_, pv357, pv423_0_, pv542, pv621, pv630,
    pv780, pv1297_4_, pv1671_0_, pv1921_2_, pv547, pv655, pv1467_0_,
    pv1629_0_, pv1863_0_, pv1896_0_, pv1921_5_, pv1953_6_, pv377, pv548,
    pv654, pv821_0_, pv1431, pv1897_0_, pv1921_4_, pv1953_7_, pv1960_1_,
    pv527, pv538, pv545, pv653, pv1829_0_, pv1898_0_, pv537, pv546,
    pv597_0_, pv652, pv801, pv1864_0_, pv1899_0_, pv572_8_, pv585_0_,
    pv1709_1_, pv1760_0_, pv373, pv572_7_, pv1439_0_, pv1709_0_, pv572_6_,
    pv1539, pv1719, pv1960_0_, pv572_5_, pv1392_0_, pv1536_0_, pv1679_0_,
    pv1833_0_, pv356, pv435_0_, pv1492_0_, pv1537, pv511_0_, pv540,
    pv609_0_, pv1426, pv1620_0_, pv1736, pv1429, pv1832, pv432, pv572_9_,
    pv1297_0_, pv1428, pv1495_0_, pv1693_0_, pv1901_0_, pv572_0_,
    pv1243_8_, pv1258, pv1243_7_, pv1259, pv1552_0_, pv1745_0_, pv1829_9_,
    pv798_0_, pv1243_6_, pv1552_1_, pv1645_0_, pv1652_0_, pv603_0_,
    pv1213_0_, pv1243_5_, pv1378, pv1387, pv572_4_, pv826_0_, pv1213_1_,
    pv1669, pv572_3_, pv591_0_, pv966, pv1213_2_, pv1709_4_, pv398_0_,
    pv572_2_, pv640_0_, pv1213_3_, pv1512_1_, pv1709_3_, pv572_1_, pv986,
    pv1213_4_, pv1243_9_, pv1451_0_, pv1512_2_, pv1613_0_, pv1709_2_;
  wire new_n483_, new_n484_, new_n485_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_,
    new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1104_, new_n1105_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1113_, new_n1114_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1125_, new_n1126_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1140_, new_n1141_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1152_, new_n1153_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1170_, new_n1171_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1189_, new_n1190_, new_n1192_,
    new_n1193_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1303_, new_n1304_, new_n1305_, new_n1308_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1325_, new_n1326_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1355_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1425_, new_n1426_, new_n1428_,
    new_n1429_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1470_,
    new_n1471_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1489_, new_n1490_, new_n1491_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1521_, new_n1522_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1559_, new_n1560_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1598_, new_n1599_, new_n1600_, new_n1602_, new_n1603_,
    new_n1604_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1620_, new_n1621_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1628_, new_n1629_, new_n1630_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1656_, new_n1658_, new_n1659_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1684_, new_n1685_, new_n1689_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1704_, new_n1705_,
    new_n1706_, new_n1707_, new_n1709_, new_n1710_, new_n1712_, new_n1713_,
    new_n1714_, new_n1715_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2046_, new_n2047_, new_n2048_, new_n2050_, new_n2051_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2104_, new_n2105_, new_n2106_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2114_, new_n2115_,
    new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2121_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2131_, new_n2132_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2165_, new_n2166_, new_n2167_, new_n2169_, new_n2170_,
    new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2182_, new_n2183_,
    new_n2184_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2194_, new_n2195_, new_n2196_, new_n2198_, new_n2199_,
    new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2206_,
    new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_,
    new_n2214_, new_n2215_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2222_, new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2230_,
    new_n2231_, new_n2232_, new_n2234_, new_n2235_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2260_,
    new_n2261_, new_n2262_, new_n2263_, new_n2265_, new_n2266_, new_n2268_,
    new_n2269_, new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2278_,
    new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2286_,
    new_n2287_, new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_,
    new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_,
    new_n2300_, new_n2301_, new_n2302_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2314_,
    new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2321_,
    new_n2322_, new_n2323_, new_n2325_, new_n2326_, new_n2327_, new_n2329_,
    new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_,
    new_n2337_, new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_,
    new_n2344_, new_n2345_, new_n2347_, new_n2348_, new_n2349_, new_n2350_,
    new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_,
    new_n2357_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2374_, new_n2375_, new_n2376_, new_n2377_,
    new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_,
    new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_,
    new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_,
    new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_,
    new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_,
    new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_,
    new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_,
    new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_,
    new_n2426_, new_n2427_, new_n2428_, new_n2431_, new_n2432_, new_n2433_,
    new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2440_, new_n2443_,
    new_n2444_, new_n2445_, new_n2446_, new_n2449_, new_n2450_, new_n2451_,
    new_n2452_, new_n2453_, new_n2455_, new_n2456_, new_n2457_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2465_, new_n2466_, new_n2468_,
    new_n2469_, new_n2470_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2480_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2503_, new_n2504_,
    new_n2506_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2559_, new_n2560_, new_n2562_,
    new_n2563_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_,
    new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2576_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_,
    new_n2585_, new_n2586_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2617_,
    new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_,
    new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2630_,
    new_n2631_, new_n2632_, new_n2634_, new_n2635_, new_n2636_, new_n2637_,
    new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2644_,
    new_n2645_, new_n2646_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_,
    new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2684_, new_n2685_,
    new_n2686_, new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_,
    new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_,
    new_n2699_, new_n2700_, new_n2701_, new_n2703_, new_n2704_, new_n2705_,
    new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2730_, new_n2731_, new_n2732_,
    new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_,
    new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_,
    new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2751_,
    new_n2752_, new_n2753_;
  assign pv778 = pv5_0_ & pv9_0_;
  assign new_n483_ = pv71_0_ & pv202_0_;
  assign new_n484_ = ~pv13_0_ & new_n483_;
  assign new_n485_ = pv4_0_ & ~new_n484_;
  assign pv789 = pv9_0_ & new_n485_;
  assign new_n487_ = pv149_2_ & ~pv149_3_;
  assign new_n488_ = ~pv149_0_ & new_n487_;
  assign new_n489_ = pv149_1_ & new_n488_;
  assign new_n490_ = pv149_4_ & new_n489_;
  assign new_n491_ = ~pv174_0_ & new_n490_;
  assign new_n492_ = ~pv149_0_ & pv149_2_;
  assign new_n493_ = ~pv149_1_ & new_n492_;
  assign new_n494_ = pv149_3_ & new_n493_;
  assign new_n495_ = ~new_n491_ & ~new_n494_;
  assign new_n496_ = pv60_0_ & ~new_n495_;
  assign new_n497_ = ~pv149_4_ & ~pv149_3_;
  assign new_n498_ = new_n493_ & new_n497_;
  assign new_n499_ = ~pv149_5_ & new_n498_;
  assign new_n500_ = pv149_4_ & ~pv149_3_;
  assign new_n501_ = new_n493_ & new_n500_;
  assign new_n502_ = ~pv149_5_ & new_n501_;
  assign new_n503_ = pv149_5_ & new_n498_;
  assign new_n504_ = ~new_n499_ & ~new_n502_;
  assign new_n505_ = ~new_n503_ & new_n504_;
  assign new_n506_ = pv277_0_ & new_n491_;
  assign new_n507_ = pv278_0_ & ~new_n506_;
  assign new_n508_ = new_n491_ & ~new_n507_;
  assign new_n509_ = ~pv149_0_ & ~pv149_1_;
  assign new_n510_ = ~pv149_2_ & new_n509_;
  assign new_n511_ = ~pv174_0_ & new_n510_;
  assign pv707 = ~pv149_3_ & new_n511_;
  assign new_n513_ = pv149_4_ & pv707;
  assign new_n514_ = ~pv149_5_ & new_n513_;
  assign new_n515_ = pv149_5_ & new_n513_;
  assign new_n516_ = pv88_2_ & pv88_3_;
  assign new_n517_ = ~pv149_4_ & new_n516_;
  assign new_n518_ = pv707 & new_n517_;
  assign new_n519_ = ~pv149_5_ & new_n518_;
  assign new_n520_ = ~pv88_2_ & pv88_3_;
  assign new_n521_ = ~pv149_4_ & new_n520_;
  assign new_n522_ = pv707 & new_n521_;
  assign new_n523_ = ~pv149_5_ & new_n522_;
  assign new_n524_ = pv149_5_ & ~pv88_2_;
  assign new_n525_ = ~pv149_3_ & new_n524_;
  assign new_n526_ = new_n511_ & new_n525_;
  assign new_n527_ = ~pv149_4_ & new_n526_;
  assign new_n528_ = pv88_3_ & new_n527_;
  assign new_n529_ = pv149_5_ & pv88_2_;
  assign new_n530_ = ~pv149_3_ & new_n529_;
  assign new_n531_ = new_n511_ & new_n530_;
  assign new_n532_ = ~pv149_4_ & new_n531_;
  assign new_n533_ = ~pv88_3_ & new_n532_;
  assign new_n534_ = pv88_2_ & ~pv88_3_;
  assign new_n535_ = ~pv149_4_ & new_n534_;
  assign new_n536_ = pv707 & new_n535_;
  assign new_n537_ = ~pv149_5_ & new_n536_;
  assign new_n538_ = ~pv88_3_ & new_n527_;
  assign new_n539_ = ~new_n514_ & ~new_n515_;
  assign new_n540_ = ~new_n519_ & ~new_n523_;
  assign new_n541_ = new_n539_ & new_n540_;
  assign new_n542_ = ~new_n528_ & ~new_n533_;
  assign new_n543_ = ~new_n537_ & ~new_n538_;
  assign new_n544_ = new_n542_ & new_n543_;
  assign new_n545_ = new_n541_ & new_n544_;
  assign new_n546_ = pv149_3_ & new_n511_;
  assign new_n547_ = new_n505_ & ~new_n508_;
  assign new_n548_ = new_n545_ & new_n547_;
  assign new_n549_ = ~new_n494_ & ~new_n546_;
  assign new_n550_ = new_n548_ & new_n549_;
  assign new_n551_ = ~pv53_0_ & ~pv56_0_;
  assign new_n552_ = ~pv57_0_ & new_n551_;
  assign new_n553_ = ~new_n493_ & ~new_n510_;
  assign new_n554_ = pv169_1_ & ~new_n553_;
  assign new_n555_ = ~new_n545_ & new_n554_;
  assign new_n556_ = pv60_0_ & new_n555_;
  assign new_n557_ = new_n546_ & new_n554_;
  assign new_n558_ = pv56_0_ & new_n557_;
  assign new_n559_ = pv60_0_ & new_n557_;
  assign new_n560_ = pv56_0_ & new_n555_;
  assign new_n561_ = ~new_n556_ & ~new_n558_;
  assign new_n562_ = ~new_n559_ & ~new_n560_;
  assign new_n563_ = new_n561_ & new_n562_;
  assign new_n564_ = ~new_n550_ & ~new_n552_;
  assign new_n565_ = new_n563_ & new_n564_;
  assign new_n566_ = ~pv149_0_ & pv149_1_;
  assign new_n567_ = ~pv149_2_ & new_n566_;
  assign new_n568_ = pv149_4_ & new_n567_;
  assign new_n569_ = ~pv149_5_ & new_n568_;
  assign new_n570_ = ~pv149_3_ & new_n569_;
  assign new_n571_ = pv149_7_ & new_n570_;
  assign new_n572_ = pv149_6_ & new_n571_;
  assign new_n573_ = ~pv149_4_ & new_n489_;
  assign new_n574_ = pv149_1_ & new_n492_;
  assign new_n575_ = pv149_3_ & new_n574_;
  assign new_n576_ = ~pv165_6_ & ~pv165_4_;
  assign new_n577_ = ~pv165_5_ & new_n576_;
  assign new_n578_ = pv165_3_ & new_n577_;
  assign new_n579_ = pv70_0_ & new_n578_;
  assign new_n580_ = pv149_5_ & new_n568_;
  assign new_n581_ = ~pv149_3_ & new_n580_;
  assign new_n582_ = pv149_7_ & new_n581_;
  assign new_n583_ = pv149_6_ & new_n582_;
  assign new_n584_ = ~pv149_7_ & new_n581_;
  assign new_n585_ = pv149_6_ & new_n584_;
  assign new_n586_ = ~new_n583_ & ~new_n585_;
  assign pv802_0_ = pv52_0_ | pv51_0_;
  assign new_n588_ = ~new_n586_ & ~pv802_0_;
  assign new_n589_ = ~pv55_0_ & new_n588_;
  assign new_n590_ = ~new_n490_ & ~new_n510_;
  assign new_n591_ = ~new_n589_ & new_n590_;
  assign new_n592_ = ~pv292_0_ & ~new_n579_;
  assign new_n593_ = ~new_n591_ & new_n592_;
  assign new_n594_ = ~pv291_0_ & new_n593_;
  assign pv763 = pv169_0_ & new_n594_;
  assign new_n596_ = pv165_3_ & pv165_5_;
  assign new_n597_ = pv165_7_ & new_n596_;
  assign new_n598_ = pv261_0_ & new_n597_;
  assign new_n599_ = pv70_0_ & new_n598_;
  assign new_n600_ = pv763 & new_n599_;
  assign new_n601_ = pv165_2_ & new_n600_;
  assign new_n602_ = pv165_0_ & new_n601_;
  assign new_n603_ = pv165_1_ & new_n602_;
  assign new_n604_ = pv165_4_ & new_n603_;
  assign new_n605_ = pv165_6_ & new_n604_;
  assign new_n606_ = pv165_3_ & pv165_4_;
  assign new_n607_ = pv165_6_ & new_n606_;
  assign new_n608_ = pv165_5_ & new_n607_;
  assign new_n609_ = pv165_7_ & new_n608_;
  assign new_n610_ = pv165_2_ & new_n609_;
  assign new_n611_ = pv165_0_ & new_n610_;
  assign new_n612_ = pv165_1_ & new_n611_;
  assign new_n613_ = pv261_0_ & new_n612_;
  assign new_n614_ = ~pv204_0_ & new_n613_;
  assign new_n615_ = ~new_n605_ & ~new_n614_;
  assign new_n616_ = ~pv262_0_ & new_n615_;
  assign new_n617_ = pv53_0_ & ~pv56_0_;
  assign new_n618_ = ~new_n573_ & new_n617_;
  assign new_n619_ = ~new_n575_ & new_n618_;
  assign new_n620_ = new_n616_ & new_n619_;
  assign new_n621_ = ~new_n565_ & ~new_n572_;
  assign new_n622_ = ~new_n620_ & new_n621_;
  assign new_n623_ = ~new_n496_ & ~new_n622_;
  assign new_n624_ = pv763 & new_n616_;
  assign new_n625_ = new_n507_ & new_n575_;
  assign new_n626_ = ~new_n491_ & new_n553_;
  assign new_n627_ = ~new_n573_ & new_n626_;
  assign new_n628_ = ~pv174_0_ & ~new_n627_;
  assign new_n629_ = ~pv60_0_ & ~pv59_0_;
  assign new_n630_ = ~new_n507_ & ~new_n629_;
  assign new_n631_ = new_n575_ & new_n630_;
  assign new_n632_ = ~new_n625_ & ~new_n628_;
  assign new_n633_ = ~new_n631_ & new_n632_;
  assign new_n634_ = ~new_n507_ & new_n575_;
  assign new_n635_ = ~pv59_0_ & new_n634_;
  assign new_n636_ = ~new_n616_ & new_n633_;
  assign new_n637_ = ~new_n635_ & new_n636_;
  assign new_n638_ = pv257_0_ & new_n637_;
  assign new_n639_ = ~new_n491_ & ~new_n575_;
  assign new_n640_ = ~new_n573_ & new_n639_;
  assign new_n641_ = ~new_n553_ & new_n640_;
  assign new_n642_ = pv223_5_ & new_n641_;
  assign new_n643_ = new_n553_ & ~new_n640_;
  assign new_n644_ = pv183_5_ & new_n643_;
  assign new_n645_ = ~new_n642_ & ~new_n644_;
  assign new_n646_ = new_n616_ & ~new_n633_;
  assign new_n647_ = ~new_n635_ & new_n646_;
  assign new_n648_ = ~new_n645_ & new_n647_;
  assign new_n649_ = ~new_n638_ & ~new_n648_;
  assign new_n650_ = ~new_n624_ & ~new_n649_;
  assign new_n651_ = ~pv56_0_ & ~pv59_0_;
  assign new_n652_ = ~pv60_0_ & new_n651_;
  assign new_n653_ = pv763 & ~new_n652_;
  assign new_n654_ = new_n624_ & ~new_n653_;
  assign new_n655_ = new_n624_ & new_n654_;
  assign new_n656_ = ~new_n653_ & new_n655_;
  assign new_n657_ = ~new_n650_ & ~new_n656_;
  assign new_n658_ = new_n622_ & ~new_n623_;
  assign new_n659_ = ~new_n657_ & new_n658_;
  assign new_n660_ = ~new_n622_ & new_n623_;
  assign new_n661_ = pv32_5_ & new_n660_;
  assign pv1213_5_ = new_n659_ | new_n661_;
  assign new_n663_ = new_n575_ & new_n616_;
  assign new_n664_ = ~pv59_0_ & new_n663_;
  assign new_n665_ = ~new_n507_ & new_n664_;
  assign new_n666_ = pv149_4_ & new_n665_;
  assign new_n667_ = new_n633_ & new_n666_;
  assign new_n668_ = pv257_7_ & new_n637_;
  assign new_n669_ = pv234_0_ & new_n641_;
  assign new_n670_ = pv194_0_ & new_n643_;
  assign new_n671_ = ~new_n669_ & ~new_n670_;
  assign new_n672_ = new_n647_ & ~new_n671_;
  assign new_n673_ = ~new_n667_ & ~new_n668_;
  assign new_n674_ = ~new_n672_ & new_n673_;
  assign new_n675_ = ~new_n624_ & ~new_n674_;
  assign new_n676_ = pv32_2_ & new_n653_;
  assign new_n677_ = pv32_5_ & ~new_n653_;
  assign new_n678_ = ~new_n676_ & ~new_n677_;
  assign new_n679_ = new_n624_ & ~new_n678_;
  assign new_n680_ = ~new_n675_ & ~new_n679_;
  assign new_n681_ = new_n658_ & ~new_n680_;
  assign new_n682_ = pv78_4_ & new_n660_;
  assign pv321_2_ = ~new_n681_ & ~new_n682_;
  assign pv1260 = pv3_0_ & pv11_0_;
  assign pv1261 = ~pv62_0_ & pv1260;
  assign new_n686_ = pv268_4_ & pv268_3_;
  assign new_n687_ = pv268_2_ & new_n686_;
  assign new_n688_ = pv268_5_ & new_n687_;
  assign new_n689_ = pv268_1_ & ~new_n688_;
  assign new_n690_ = ~pv268_1_ & new_n688_;
  assign pv1371 = new_n689_ | new_n690_;
  assign new_n692_ = pv10_0_ & ~pv13_0_;
  assign new_n693_ = ~new_n493_ & ~new_n511_;
  assign new_n694_ = pv802_0_ & ~new_n693_;
  assign new_n695_ = ~new_n494_ & ~new_n694_;
  assign pv782 = pv7_0_ & new_n692_;
  assign pv1382 = ~new_n695_ & pv782;
  assign new_n698_ = pv165_0_ & pv165_1_;
  assign new_n699_ = ~pv165_2_ & new_n698_;
  assign new_n700_ = pv165_7_ & new_n699_;
  assign new_n701_ = ~pv290_0_ & new_n700_;
  assign new_n702_ = ~pv165_7_ & new_n699_;
  assign new_n703_ = pv172_0_ & pv56_0_;
  assign new_n704_ = pv207_0_ & ~new_n703_;
  assign new_n705_ = pv59_0_ & new_n554_;
  assign new_n706_ = new_n704_ & new_n705_;
  assign new_n707_ = ~new_n493_ & new_n706_;
  assign new_n708_ = ~pv149_4_ & new_n567_;
  assign new_n709_ = pv149_5_ & new_n708_;
  assign new_n710_ = ~pv149_3_ & new_n709_;
  assign new_n711_ = ~pv149_7_ & new_n710_;
  assign new_n712_ = ~pv149_6_ & new_n711_;
  assign new_n713_ = ~pv174_0_ & new_n583_;
  assign new_n714_ = ~new_n554_ & ~new_n712_;
  assign new_n715_ = new_n704_ & new_n714_;
  assign new_n716_ = ~new_n713_ & new_n715_;
  assign new_n717_ = ~new_n493_ & new_n716_;
  assign new_n718_ = pv172_0_ & pv215_0_;
  assign new_n719_ = pv67_0_ & new_n718_;
  assign new_n720_ = pv59_0_ & new_n713_;
  assign new_n721_ = new_n704_ & new_n720_;
  assign new_n722_ = ~new_n493_ & new_n721_;
  assign new_n723_ = pv62_0_ & new_n712_;
  assign new_n724_ = new_n704_ & new_n723_;
  assign new_n725_ = ~new_n493_ & new_n724_;
  assign new_n726_ = ~pv214_0_ & ~new_n707_;
  assign new_n727_ = ~new_n717_ & new_n726_;
  assign new_n728_ = ~new_n719_ & ~new_n722_;
  assign new_n729_ = ~new_n725_ & new_n728_;
  assign new_n730_ = new_n727_ & new_n729_;
  assign new_n731_ = pv241_0_ & ~new_n639_;
  assign new_n732_ = ~new_n573_ & ~new_n731_;
  assign new_n733_ = ~pv275_0_ & pv272_0_;
  assign new_n734_ = ~new_n732_ & new_n733_;
  assign new_n735_ = ~pv802_0_ & new_n734_;
  assign new_n736_ = pv261_0_ & new_n735_;
  assign new_n737_ = new_n507_ & new_n736_;
  assign new_n738_ = pv261_0_ & ~pv802_0_;
  assign new_n739_ = ~new_n732_ & new_n738_;
  assign new_n740_ = ~new_n507_ & new_n739_;
  assign new_n741_ = pv56_0_ & ~new_n639_;
  assign new_n742_ = ~pv802_0_ & ~new_n640_;
  assign new_n743_ = ~new_n507_ & new_n742_;
  assign new_n744_ = pv242_0_ & new_n743_;
  assign new_n745_ = ~new_n741_ & new_n744_;
  assign new_n746_ = pv272_0_ & ~pv802_0_;
  assign new_n747_ = pv134_0_ & new_n746_;
  assign new_n748_ = pv242_0_ & new_n747_;
  assign new_n749_ = pv134_1_ & new_n748_;
  assign new_n750_ = ~pv275_0_ & new_n749_;
  assign new_n751_ = new_n507_ & new_n750_;
  assign new_n752_ = new_n730_ & ~new_n737_;
  assign new_n753_ = ~new_n740_ & new_n752_;
  assign new_n754_ = ~new_n745_ & ~new_n751_;
  assign new_n755_ = new_n753_ & new_n754_;
  assign new_n756_ = ~new_n701_ & ~new_n702_;
  assign new_n757_ = ~pv302_0_ & new_n755_;
  assign new_n758_ = new_n756_ & new_n757_;
  assign new_n759_ = ~pv149_5_ & new_n708_;
  assign new_n760_ = ~pv149_3_ & new_n759_;
  assign new_n761_ = pv149_7_ & new_n760_;
  assign new_n762_ = pv149_6_ & new_n761_;
  assign new_n763_ = pv67_0_ & pv14_0_;
  assign new_n764_ = new_n758_ & new_n763_;
  assign pv1470 = ~new_n762_ & new_n764_;
  assign new_n766_ = pv149_5_ & new_n501_;
  assign new_n767_ = pv88_3_ & new_n532_;
  assign new_n768_ = ~pv88_2_ & ~pv88_3_;
  assign new_n769_ = ~pv149_4_ & new_n768_;
  assign new_n770_ = pv707 & new_n769_;
  assign new_n771_ = ~pv149_5_ & new_n770_;
  assign new_n772_ = ~new_n767_ & ~new_n771_;
  assign new_n773_ = ~new_n554_ & ~new_n772_;
  assign new_n774_ = ~new_n766_ & ~new_n773_;
  assign new_n775_ = pv56_0_ & ~new_n774_;
  assign new_n776_ = ~pv172_0_ & new_n775_;
  assign new_n777_ = pv278_0_ & ~new_n640_;
  assign new_n778_ = pv171_0_ & ~new_n553_;
  assign new_n779_ = pv56_0_ & new_n778_;
  assign new_n780_ = ~pv248_0_ & ~new_n703_;
  assign new_n781_ = ~new_n777_ & new_n780_;
  assign new_n782_ = pv177_0_ & new_n781_;
  assign new_n783_ = ~new_n779_ & new_n782_;
  assign new_n784_ = ~pv274_0_ & ~pv271_0_;
  assign new_n785_ = new_n554_ & ~new_n772_;
  assign new_n786_ = pv59_0_ & new_n785_;
  assign new_n787_ = ~new_n776_ & ~new_n783_;
  assign new_n788_ = ~new_n784_ & new_n787_;
  assign new_n789_ = ~new_n786_ & new_n788_;
  assign new_n790_ = new_n493_ & new_n704_;
  assign new_n791_ = pv149_7_ & new_n493_;
  assign new_n792_ = pv56_0_ & new_n791_;
  assign new_n793_ = ~new_n790_ & ~new_n792_;
  assign new_n794_ = ~new_n789_ & new_n793_;
  assign pv1536_0_ = ~new_n755_ | ~new_n794_;
  assign new_n796_ = new_n755_ & pv1536_0_;
  assign new_n797_ = pv223_2_ & new_n641_;
  assign new_n798_ = pv183_2_ & new_n643_;
  assign new_n799_ = ~new_n797_ & ~new_n798_;
  assign new_n800_ = new_n616_ & ~new_n635_;
  assign new_n801_ = ~new_n633_ & new_n800_;
  assign new_n802_ = ~new_n799_ & new_n801_;
  assign new_n803_ = ~new_n624_ & new_n802_;
  assign new_n804_ = new_n622_ & new_n803_;
  assign new_n805_ = ~new_n624_ & new_n804_;
  assign new_n806_ = ~new_n623_ & new_n805_;
  assign new_n807_ = pv32_2_ & new_n660_;
  assign pv1213_2_ = new_n806_ | new_n807_;
  assign new_n809_ = pv223_3_ & new_n641_;
  assign new_n810_ = pv183_3_ & new_n643_;
  assign new_n811_ = ~new_n809_ & ~new_n810_;
  assign new_n812_ = new_n801_ & ~new_n811_;
  assign new_n813_ = ~new_n624_ & new_n812_;
  assign new_n814_ = new_n622_ & new_n813_;
  assign new_n815_ = ~new_n624_ & new_n814_;
  assign new_n816_ = ~new_n623_ & new_n815_;
  assign new_n817_ = pv32_3_ & new_n660_;
  assign pv1213_3_ = new_n816_ | new_n817_;
  assign new_n819_ = pv223_1_ & new_n641_;
  assign new_n820_ = pv183_1_ & new_n643_;
  assign new_n821_ = ~new_n819_ & ~new_n820_;
  assign new_n822_ = new_n801_ & ~new_n821_;
  assign new_n823_ = ~new_n624_ & new_n822_;
  assign new_n824_ = new_n622_ & new_n823_;
  assign new_n825_ = ~new_n624_ & new_n824_;
  assign new_n826_ = ~new_n623_ & new_n825_;
  assign new_n827_ = pv32_1_ & new_n660_;
  assign pv1213_1_ = new_n826_ | new_n827_;
  assign new_n829_ = pv223_0_ & new_n641_;
  assign new_n830_ = pv183_0_ & new_n643_;
  assign new_n831_ = ~new_n829_ & ~new_n830_;
  assign new_n832_ = new_n801_ & ~new_n831_;
  assign new_n833_ = ~new_n624_ & new_n832_;
  assign new_n834_ = new_n622_ & new_n833_;
  assign new_n835_ = ~new_n624_ & new_n834_;
  assign new_n836_ = ~new_n623_ & new_n835_;
  assign new_n837_ = pv32_0_ & new_n660_;
  assign pv1213_0_ = new_n836_ | new_n837_;
  assign new_n839_ = pv149_3_ & new_n759_;
  assign new_n840_ = ~pv149_7_ & new_n839_;
  assign new_n841_ = ~pv149_6_ & new_n840_;
  assign new_n842_ = ~pv802_0_ & new_n841_;
  assign new_n843_ = pv1213_2_ & pv1213_3_;
  assign new_n844_ = ~pv1213_1_ & new_n843_;
  assign new_n845_ = ~pv1213_0_ & new_n844_;
  assign new_n846_ = ~new_n842_ & new_n845_;
  assign new_n847_ = pv288_6_ & new_n846_;
  assign new_n848_ = pv288_7_ & new_n847_;
  assign new_n849_ = ~pv1213_3_ & ~pv1213_0_;
  assign new_n850_ = pv1213_2_ & new_n849_;
  assign new_n851_ = ~pv1213_1_ & new_n850_;
  assign new_n852_ = ~new_n842_ & new_n851_;
  assign new_n853_ = pv288_6_ & new_n852_;
  assign new_n854_ = pv288_7_ & new_n853_;
  assign new_n855_ = ~pv288_6_ & pv288_7_;
  assign new_n856_ = ~pv288_4_ & pv288_5_;
  assign new_n857_ = new_n855_ & new_n856_;
  assign new_n858_ = ~new_n855_ & ~new_n856_;
  assign new_n859_ = ~new_n857_ & ~new_n858_;
  assign new_n860_ = ~pv288_2_ & pv288_3_;
  assign new_n861_ = ~new_n859_ & new_n860_;
  assign new_n862_ = pv288_2_ & ~pv288_3_;
  assign new_n863_ = new_n861_ & new_n862_;
  assign new_n864_ = ~new_n855_ & new_n856_;
  assign new_n865_ = pv288_6_ & ~pv288_7_;
  assign new_n866_ = ~new_n855_ & ~new_n865_;
  assign new_n867_ = pv288_4_ & ~pv288_5_;
  assign new_n868_ = ~new_n866_ & new_n867_;
  assign new_n869_ = new_n866_ & ~new_n867_;
  assign new_n870_ = ~new_n868_ & ~new_n869_;
  assign new_n871_ = ~new_n864_ & ~new_n870_;
  assign new_n872_ = new_n864_ & new_n870_;
  assign new_n873_ = ~new_n871_ & ~new_n872_;
  assign new_n874_ = new_n862_ & ~new_n873_;
  assign new_n875_ = new_n861_ & ~new_n873_;
  assign new_n876_ = ~new_n863_ & ~new_n874_;
  assign new_n877_ = ~new_n875_ & new_n876_;
  assign new_n878_ = pv288_2_ & pv288_3_;
  assign new_n879_ = ~new_n877_ & new_n878_;
  assign new_n880_ = ~pv288_6_ & ~pv288_7_;
  assign new_n881_ = pv288_4_ & pv288_5_;
  assign new_n882_ = ~new_n880_ & new_n881_;
  assign new_n883_ = new_n880_ & ~new_n881_;
  assign new_n884_ = ~new_n882_ & ~new_n883_;
  assign new_n885_ = new_n864_ & new_n867_;
  assign new_n886_ = new_n866_ & new_n867_;
  assign new_n887_ = new_n864_ & new_n866_;
  assign new_n888_ = ~new_n885_ & ~new_n886_;
  assign new_n889_ = ~new_n887_ & new_n888_;
  assign new_n890_ = new_n884_ & ~new_n889_;
  assign new_n891_ = ~new_n884_ & new_n889_;
  assign new_n892_ = ~new_n890_ & ~new_n891_;
  assign new_n893_ = new_n878_ & ~new_n892_;
  assign new_n894_ = ~new_n877_ & ~new_n892_;
  assign new_n895_ = ~new_n879_ & ~new_n893_;
  assign new_n896_ = ~new_n894_ & new_n895_;
  assign new_n897_ = new_n881_ & ~new_n889_;
  assign new_n898_ = new_n880_ & new_n881_;
  assign new_n899_ = new_n880_ & ~new_n889_;
  assign new_n900_ = ~new_n897_ & ~new_n898_;
  assign new_n901_ = ~new_n899_ & new_n900_;
  assign new_n902_ = new_n880_ & new_n901_;
  assign new_n903_ = ~new_n880_ & ~new_n901_;
  assign new_n904_ = ~new_n902_ & ~new_n903_;
  assign new_n905_ = new_n896_ & ~new_n904_;
  assign new_n906_ = ~new_n896_ & new_n904_;
  assign new_n907_ = ~new_n905_ & ~new_n906_;
  assign new_n908_ = ~pv1213_0_ & ~new_n907_;
  assign new_n909_ = pv1213_0_ & new_n907_;
  assign new_n910_ = ~new_n908_ & ~new_n909_;
  assign new_n911_ = new_n862_ & new_n873_;
  assign new_n912_ = ~new_n862_ & ~new_n873_;
  assign new_n913_ = ~new_n911_ & ~new_n912_;
  assign new_n914_ = ~new_n861_ & ~new_n913_;
  assign new_n915_ = new_n861_ & new_n913_;
  assign new_n916_ = ~new_n914_ & ~new_n915_;
  assign new_n917_ = ~pv1213_2_ & ~new_n916_;
  assign new_n918_ = pv1213_2_ & new_n916_;
  assign new_n919_ = ~new_n917_ & ~new_n918_;
  assign new_n920_ = new_n859_ & new_n860_;
  assign new_n921_ = ~new_n859_ & ~new_n860_;
  assign new_n922_ = ~new_n920_ & ~new_n921_;
  assign new_n923_ = ~pv1213_3_ & ~new_n922_;
  assign new_n924_ = pv1213_3_ & new_n922_;
  assign new_n925_ = ~new_n923_ & ~new_n924_;
  assign new_n926_ = new_n878_ & new_n892_;
  assign new_n927_ = ~new_n878_ & ~new_n892_;
  assign new_n928_ = ~new_n926_ & ~new_n927_;
  assign new_n929_ = ~new_n877_ & new_n928_;
  assign new_n930_ = new_n877_ & ~new_n928_;
  assign new_n931_ = ~new_n929_ & ~new_n930_;
  assign new_n932_ = ~pv1213_1_ & ~new_n931_;
  assign new_n933_ = pv1213_1_ & new_n931_;
  assign new_n934_ = ~new_n932_ & ~new_n933_;
  assign new_n935_ = new_n910_ & new_n919_;
  assign new_n936_ = new_n925_ & new_n935_;
  assign new_n937_ = new_n934_ & new_n936_;
  assign new_n938_ = ~new_n842_ & new_n937_;
  assign new_n939_ = new_n878_ & new_n938_;
  assign new_n940_ = ~pv1213_0_ & ~new_n904_;
  assign new_n941_ = pv1213_0_ & new_n904_;
  assign new_n942_ = ~new_n940_ & ~new_n941_;
  assign new_n943_ = ~pv1213_2_ & ~new_n873_;
  assign new_n944_ = pv1213_2_ & new_n873_;
  assign new_n945_ = ~new_n943_ & ~new_n944_;
  assign new_n946_ = ~pv1213_3_ & ~new_n859_;
  assign new_n947_ = pv1213_3_ & new_n859_;
  assign new_n948_ = ~new_n946_ & ~new_n947_;
  assign new_n949_ = ~pv1213_1_ & ~new_n892_;
  assign new_n950_ = pv1213_1_ & new_n892_;
  assign new_n951_ = ~new_n949_ & ~new_n950_;
  assign new_n952_ = new_n942_ & new_n945_;
  assign new_n953_ = new_n948_ & new_n952_;
  assign new_n954_ = new_n951_ & new_n953_;
  assign new_n955_ = ~new_n842_ & new_n954_;
  assign new_n956_ = new_n881_ & new_n955_;
  assign new_n957_ = ~pv288_0_ & pv288_1_;
  assign new_n958_ = ~new_n922_ & new_n957_;
  assign new_n959_ = pv288_0_ & ~pv288_1_;
  assign new_n960_ = new_n958_ & new_n959_;
  assign new_n961_ = ~new_n916_ & new_n959_;
  assign new_n962_ = ~new_n916_ & new_n958_;
  assign new_n963_ = ~new_n960_ & ~new_n961_;
  assign new_n964_ = ~new_n962_ & new_n963_;
  assign new_n965_ = pv288_0_ & pv288_1_;
  assign new_n966_ = ~new_n964_ & new_n965_;
  assign new_n967_ = ~new_n931_ & new_n965_;
  assign new_n968_ = ~new_n931_ & ~new_n964_;
  assign new_n969_ = ~new_n966_ & ~new_n967_;
  assign new_n970_ = ~new_n968_ & new_n969_;
  assign new_n971_ = ~new_n907_ & new_n970_;
  assign new_n972_ = new_n907_ & ~new_n970_;
  assign new_n973_ = ~new_n971_ & ~new_n972_;
  assign new_n974_ = ~pv1213_0_ & ~new_n973_;
  assign new_n975_ = pv1213_0_ & new_n973_;
  assign new_n976_ = ~new_n974_ & ~new_n975_;
  assign new_n977_ = new_n916_ & new_n959_;
  assign new_n978_ = ~new_n916_ & ~new_n959_;
  assign new_n979_ = ~new_n977_ & ~new_n978_;
  assign new_n980_ = ~new_n958_ & ~new_n979_;
  assign new_n981_ = new_n958_ & new_n979_;
  assign new_n982_ = ~new_n980_ & ~new_n981_;
  assign new_n983_ = ~pv1213_2_ & ~new_n982_;
  assign new_n984_ = pv1213_2_ & new_n982_;
  assign new_n985_ = ~new_n983_ & ~new_n984_;
  assign new_n986_ = new_n922_ & new_n957_;
  assign new_n987_ = ~new_n922_ & ~new_n957_;
  assign new_n988_ = ~new_n986_ & ~new_n987_;
  assign new_n989_ = ~pv1213_3_ & ~new_n988_;
  assign new_n990_ = pv1213_3_ & new_n988_;
  assign new_n991_ = ~new_n989_ & ~new_n990_;
  assign new_n992_ = new_n931_ & new_n965_;
  assign new_n993_ = ~new_n931_ & ~new_n965_;
  assign new_n994_ = ~new_n992_ & ~new_n993_;
  assign new_n995_ = ~new_n964_ & new_n994_;
  assign new_n996_ = new_n964_ & ~new_n994_;
  assign new_n997_ = ~new_n995_ & ~new_n996_;
  assign new_n998_ = ~pv1213_1_ & ~new_n997_;
  assign new_n999_ = pv1213_1_ & new_n997_;
  assign new_n1000_ = ~new_n998_ & ~new_n999_;
  assign new_n1001_ = new_n976_ & new_n985_;
  assign new_n1002_ = new_n991_ & new_n1001_;
  assign new_n1003_ = new_n1000_ & new_n1002_;
  assign new_n1004_ = ~new_n842_ & new_n1003_;
  assign new_n1005_ = new_n965_ & new_n1004_;
  assign new_n1006_ = new_n982_ & new_n988_;
  assign new_n1007_ = new_n997_ & new_n1006_;
  assign new_n1008_ = ~new_n973_ & ~new_n1007_;
  assign new_n1009_ = new_n973_ & new_n1007_;
  assign new_n1010_ = ~new_n1008_ & ~new_n1009_;
  assign new_n1011_ = ~pv1213_0_ & ~new_n1010_;
  assign new_n1012_ = pv1213_0_ & new_n1010_;
  assign new_n1013_ = ~new_n1011_ & ~new_n1012_;
  assign new_n1014_ = ~new_n982_ & ~new_n988_;
  assign new_n1015_ = ~new_n1006_ & ~new_n1014_;
  assign new_n1016_ = ~pv1213_2_ & ~new_n1015_;
  assign new_n1017_ = pv1213_2_ & new_n1015_;
  assign new_n1018_ = ~new_n1016_ & ~new_n1017_;
  assign new_n1019_ = ~pv1213_3_ & new_n988_;
  assign new_n1020_ = pv1213_3_ & ~new_n988_;
  assign new_n1021_ = ~new_n1019_ & ~new_n1020_;
  assign new_n1022_ = ~new_n997_ & ~new_n1006_;
  assign new_n1023_ = ~new_n1007_ & ~new_n1022_;
  assign new_n1024_ = ~pv1213_1_ & ~new_n1023_;
  assign new_n1025_ = pv1213_1_ & new_n1023_;
  assign new_n1026_ = ~new_n1024_ & ~new_n1025_;
  assign new_n1027_ = new_n1013_ & new_n1018_;
  assign new_n1028_ = new_n1021_ & new_n1027_;
  assign new_n1029_ = new_n1026_ & new_n1028_;
  assign new_n1030_ = ~new_n842_ & new_n1029_;
  assign new_n1031_ = new_n965_ & new_n1030_;
  assign new_n1032_ = new_n859_ & new_n873_;
  assign new_n1033_ = new_n892_ & new_n1032_;
  assign new_n1034_ = ~new_n904_ & ~new_n1033_;
  assign new_n1035_ = new_n904_ & new_n1033_;
  assign new_n1036_ = ~new_n1034_ & ~new_n1035_;
  assign new_n1037_ = ~pv1213_0_ & ~new_n1036_;
  assign new_n1038_ = pv1213_0_ & new_n1036_;
  assign new_n1039_ = ~new_n1037_ & ~new_n1038_;
  assign new_n1040_ = ~new_n859_ & ~new_n873_;
  assign new_n1041_ = ~new_n1032_ & ~new_n1040_;
  assign new_n1042_ = ~pv1213_2_ & ~new_n1041_;
  assign new_n1043_ = pv1213_2_ & new_n1041_;
  assign new_n1044_ = ~new_n1042_ & ~new_n1043_;
  assign new_n1045_ = ~pv1213_3_ & new_n859_;
  assign new_n1046_ = pv1213_3_ & ~new_n859_;
  assign new_n1047_ = ~new_n1045_ & ~new_n1046_;
  assign new_n1048_ = ~new_n892_ & ~new_n1032_;
  assign new_n1049_ = ~new_n1033_ & ~new_n1048_;
  assign new_n1050_ = ~pv1213_1_ & ~new_n1049_;
  assign new_n1051_ = pv1213_1_ & new_n1049_;
  assign new_n1052_ = ~new_n1050_ & ~new_n1051_;
  assign new_n1053_ = new_n1039_ & new_n1044_;
  assign new_n1054_ = new_n1047_ & new_n1053_;
  assign new_n1055_ = new_n1052_ & new_n1054_;
  assign new_n1056_ = ~new_n842_ & new_n1055_;
  assign new_n1057_ = new_n881_ & new_n1056_;
  assign new_n1058_ = new_n916_ & new_n922_;
  assign new_n1059_ = new_n931_ & new_n1058_;
  assign new_n1060_ = ~new_n907_ & ~new_n1059_;
  assign new_n1061_ = new_n907_ & new_n1059_;
  assign new_n1062_ = ~new_n1060_ & ~new_n1061_;
  assign new_n1063_ = ~pv1213_0_ & ~new_n1062_;
  assign new_n1064_ = pv1213_0_ & new_n1062_;
  assign new_n1065_ = ~new_n1063_ & ~new_n1064_;
  assign new_n1066_ = ~new_n916_ & ~new_n922_;
  assign new_n1067_ = ~new_n1058_ & ~new_n1066_;
  assign new_n1068_ = ~pv1213_2_ & ~new_n1067_;
  assign new_n1069_ = pv1213_2_ & new_n1067_;
  assign new_n1070_ = ~new_n1068_ & ~new_n1069_;
  assign new_n1071_ = ~pv1213_3_ & new_n922_;
  assign new_n1072_ = pv1213_3_ & ~new_n922_;
  assign new_n1073_ = ~new_n1071_ & ~new_n1072_;
  assign new_n1074_ = ~new_n931_ & ~new_n1058_;
  assign new_n1075_ = ~new_n1059_ & ~new_n1074_;
  assign new_n1076_ = ~pv1213_1_ & ~new_n1075_;
  assign new_n1077_ = pv1213_1_ & new_n1075_;
  assign new_n1078_ = ~new_n1076_ & ~new_n1077_;
  assign new_n1079_ = new_n1065_ & new_n1070_;
  assign new_n1080_ = new_n1073_ & new_n1079_;
  assign new_n1081_ = new_n1078_ & new_n1080_;
  assign new_n1082_ = ~new_n842_ & new_n1081_;
  assign new_n1083_ = new_n878_ & new_n1082_;
  assign new_n1084_ = ~new_n848_ & ~new_n854_;
  assign new_n1085_ = ~new_n939_ & new_n1084_;
  assign new_n1086_ = ~new_n956_ & new_n1085_;
  assign new_n1087_ = ~new_n1005_ & new_n1086_;
  assign new_n1088_ = ~new_n1031_ & new_n1087_;
  assign new_n1089_ = ~new_n1057_ & new_n1088_;
  assign new_n1090_ = ~new_n1083_ & new_n1089_;
  assign new_n1091_ = ~pv1536_0_ & ~new_n1090_;
  assign pv1512_3_ = new_n796_ | new_n1091_;
  assign new_n1093_ = pv149_6_ & new_n840_;
  assign new_n1094_ = ~pv149_7_ & new_n570_;
  assign new_n1095_ = ~pv149_6_ & new_n1094_;
  assign new_n1096_ = ~pv149_6_ & new_n571_;
  assign new_n1097_ = ~new_n1093_ & new_n1095_;
  assign new_n1098_ = ~new_n1096_ & new_n1097_;
  assign new_n1099_ = pv132_2_ & new_n1098_;
  assign new_n1100_ = ~new_n1093_ & ~new_n1095_;
  assign new_n1101_ = new_n1096_ & new_n1100_;
  assign new_n1102_ = pv118_0_ & new_n1101_;
  assign pv1953_2_ = new_n1099_ | new_n1102_;
  assign new_n1104_ = pv132_3_ & new_n1098_;
  assign new_n1105_ = pv118_1_ & new_n1101_;
  assign pv1953_3_ = new_n1104_ | new_n1105_;
  assign new_n1107_ = ~pv1953_2_ & pv1953_3_;
  assign new_n1108_ = pv1953_2_ & ~pv1953_3_;
  assign new_n1109_ = ~new_n1107_ & ~new_n1108_;
  assign new_n1110_ = pv132_4_ & new_n1098_;
  assign new_n1111_ = pv118_2_ & new_n1101_;
  assign pv1953_4_ = new_n1110_ | new_n1111_;
  assign new_n1113_ = pv132_5_ & new_n1098_;
  assign new_n1114_ = pv118_3_ & new_n1101_;
  assign pv1953_5_ = new_n1113_ | new_n1114_;
  assign new_n1116_ = ~pv1953_4_ & pv1953_5_;
  assign new_n1117_ = pv1953_4_ & ~pv1953_5_;
  assign new_n1118_ = ~new_n1116_ & ~new_n1117_;
  assign new_n1119_ = new_n1109_ & ~new_n1118_;
  assign new_n1120_ = ~new_n1109_ & new_n1118_;
  assign new_n1121_ = ~new_n1119_ & ~new_n1120_;
  assign new_n1122_ = pv132_6_ & new_n1098_;
  assign new_n1123_ = pv118_4_ & new_n1101_;
  assign pv1953_6_ = new_n1122_ | new_n1123_;
  assign new_n1125_ = pv132_7_ & new_n1098_;
  assign new_n1126_ = pv118_5_ & new_n1101_;
  assign pv1953_7_ = new_n1125_ | new_n1126_;
  assign new_n1128_ = ~pv1953_6_ & pv1953_7_;
  assign new_n1129_ = pv1953_6_ & ~pv1953_7_;
  assign new_n1130_ = ~new_n1128_ & ~new_n1129_;
  assign new_n1131_ = pv149_7_ & new_n710_;
  assign new_n1132_ = pv149_6_ & new_n1131_;
  assign new_n1133_ = pv149_6_ & new_n711_;
  assign new_n1134_ = ~new_n1132_ & ~new_n1133_;
  assign new_n1135_ = new_n1096_ & new_n1134_;
  assign new_n1136_ = pv118_6_ & new_n1135_;
  assign new_n1137_ = ~new_n1096_ & ~new_n1134_;
  assign new_n1138_ = pv48_0_ & new_n1137_;
  assign pv1960_0_ = new_n1136_ | new_n1138_;
  assign new_n1140_ = pv118_7_ & new_n1135_;
  assign new_n1141_ = pv46_0_ & new_n1137_;
  assign pv1960_1_ = new_n1140_ | new_n1141_;
  assign new_n1143_ = ~pv1960_0_ & pv1960_1_;
  assign new_n1144_ = pv1960_0_ & ~pv1960_1_;
  assign new_n1145_ = ~new_n1143_ & ~new_n1144_;
  assign new_n1146_ = new_n1130_ & ~new_n1145_;
  assign new_n1147_ = ~new_n1130_ & new_n1145_;
  assign new_n1148_ = ~new_n1146_ & ~new_n1147_;
  assign new_n1149_ = new_n1121_ & ~new_n1148_;
  assign new_n1150_ = ~new_n1121_ & new_n1148_;
  assign pv1613_1_ = ~new_n1149_ & ~new_n1150_;
  assign new_n1152_ = ~pv16_0_ & pv15_0_;
  assign new_n1153_ = pv16_0_ & pv15_0_;
  assign pv1757_0_ = new_n1152_ | new_n1153_;
  assign new_n1155_ = pv257_6_ & new_n637_;
  assign new_n1156_ = pv229_5_ & new_n641_;
  assign new_n1157_ = pv189_5_ & new_n643_;
  assign new_n1158_ = ~new_n1156_ & ~new_n1157_;
  assign new_n1159_ = new_n647_ & ~new_n1158_;
  assign new_n1160_ = ~new_n1155_ & ~new_n1159_;
  assign new_n1161_ = ~new_n624_ & ~new_n1160_;
  assign new_n1162_ = pv32_1_ & new_n653_;
  assign new_n1163_ = pv32_4_ & ~new_n653_;
  assign new_n1164_ = ~new_n1162_ & ~new_n1163_;
  assign new_n1165_ = new_n624_ & ~new_n1164_;
  assign new_n1166_ = ~new_n1161_ & ~new_n1165_;
  assign new_n1167_ = new_n658_ & ~new_n1166_;
  assign new_n1168_ = pv32_11_ & new_n660_;
  assign pv1213_11_ = new_n1167_ | new_n1168_;
  assign new_n1170_ = ~new_n572_ & ~pv1213_11_;
  assign new_n1171_ = ~pv78_3_ & new_n572_;
  assign pv1781_1_ = new_n1170_ | new_n1171_;
  assign new_n1173_ = pv234_2_ & new_n641_;
  assign new_n1174_ = pv194_2_ & new_n643_;
  assign new_n1175_ = ~new_n1173_ & ~new_n1174_;
  assign new_n1176_ = new_n647_ & ~new_n1175_;
  assign new_n1177_ = pv149_6_ & new_n665_;
  assign new_n1178_ = new_n633_ & new_n1177_;
  assign new_n1179_ = ~new_n1176_ & ~new_n1178_;
  assign new_n1180_ = ~new_n624_ & ~new_n1179_;
  assign new_n1181_ = pv32_4_ & new_n653_;
  assign new_n1182_ = pv32_7_ & ~new_n653_;
  assign new_n1183_ = ~new_n1181_ & ~new_n1182_;
  assign new_n1184_ = new_n624_ & ~new_n1183_;
  assign new_n1185_ = ~new_n1180_ & ~new_n1184_;
  assign new_n1186_ = new_n658_ & ~new_n1185_;
  assign new_n1187_ = pv84_0_ & new_n660_;
  assign pv1243_2_ = new_n1186_ | new_n1187_;
  assign new_n1189_ = pv37_0_ & ~pv1243_2_;
  assign new_n1190_ = ~pv37_0_ & ~pv1213_5_;
  assign pv1829_2_ = new_n1189_ | new_n1190_;
  assign new_n1192_ = pv109_0_ & ~pv13_0_;
  assign new_n1193_ = pv1_0_ & ~new_n1192_;
  assign pv1431 = pv9_0_ & new_n1193_;
  assign pv787 = pv7_0_ & pv9_0_;
  assign pv1423 = pv1_0_ & pv9_0_;
  assign pv1258 = pv2_0_ & pv9_0_;
  assign pv1263 = pv4_0_ & pv9_0_;
  assign pv1387 = pv8_0_ & pv9_0_;
  assign pv1259 = pv3_0_ & pv9_0_;
  assign pv780 = pv6_0_ & pv9_0_;
  assign new_n1202_ = ~pv1431 & ~pv787;
  assign new_n1203_ = ~pv1423 & new_n1202_;
  assign new_n1204_ = ~pv1423 & ~pv1258;
  assign new_n1205_ = ~pv789 & new_n1204_;
  assign new_n1206_ = new_n1203_ & new_n1205_;
  assign new_n1207_ = ~pv778 & ~pv780;
  assign new_n1208_ = ~pv1263 & ~pv1387;
  assign new_n1209_ = ~pv1259 & new_n1208_;
  assign new_n1210_ = new_n1207_ & new_n1209_;
  assign pv375_0_ = ~new_n1206_ | ~new_n1210_;
  assign new_n1212_ = pv62_0_ & new_n555_;
  assign new_n1213_ = ~new_n545_ & ~new_n554_;
  assign new_n1214_ = new_n505_ & ~new_n785_;
  assign new_n1215_ = ~new_n1213_ & new_n1214_;
  assign new_n1216_ = pv59_0_ & ~new_n1215_;
  assign new_n1217_ = ~new_n775_ & ~new_n1212_;
  assign new_n1218_ = ~new_n1216_ & new_n1217_;
  assign new_n1219_ = ~new_n699_ & ~pv1757_0_;
  assign pv410_0_ = new_n1218_ | ~new_n1219_;
  assign new_n1221_ = pv59_0_ & new_n557_;
  assign new_n1222_ = pv62_0_ & new_n1132_;
  assign new_n1223_ = ~pv149_6_ & new_n1131_;
  assign new_n1224_ = pv149_6_ & new_n1094_;
  assign new_n1225_ = ~new_n572_ & ~new_n1223_;
  assign new_n1226_ = ~new_n1224_ & new_n1225_;
  assign new_n1227_ = pv56_0_ & ~new_n1226_;
  assign new_n1228_ = ~new_n491_ & new_n693_;
  assign new_n1229_ = pv802_0_ & ~new_n1228_;
  assign new_n1230_ = ~new_n1227_ & ~new_n1229_;
  assign new_n1231_ = ~pv84_2_ & pv84_3_;
  assign new_n1232_ = pv84_2_ & ~pv84_3_;
  assign new_n1233_ = ~new_n1231_ & ~new_n1232_;
  assign new_n1234_ = ~pv84_4_ & pv84_5_;
  assign new_n1235_ = pv84_4_ & ~pv84_5_;
  assign new_n1236_ = ~new_n1234_ & ~new_n1235_;
  assign new_n1237_ = new_n1233_ & ~new_n1236_;
  assign new_n1238_ = ~new_n1233_ & new_n1236_;
  assign new_n1239_ = ~new_n1237_ & ~new_n1238_;
  assign new_n1240_ = ~pv88_0_ & pv88_1_;
  assign new_n1241_ = pv88_0_ & ~pv88_1_;
  assign new_n1242_ = ~new_n1240_ & ~new_n1241_;
  assign new_n1243_ = ~new_n520_ & ~new_n534_;
  assign new_n1244_ = new_n1242_ & ~new_n1243_;
  assign new_n1245_ = ~new_n1242_ & new_n1243_;
  assign new_n1246_ = ~new_n1244_ & ~new_n1245_;
  assign new_n1247_ = new_n1239_ & ~new_n1246_;
  assign new_n1248_ = ~new_n1239_ & new_n1246_;
  assign new_n1249_ = ~new_n1247_ & ~new_n1248_;
  assign new_n1250_ = pv94_1_ & new_n1249_;
  assign new_n1251_ = ~pv94_1_ & ~new_n1249_;
  assign new_n1252_ = ~new_n1250_ & ~new_n1251_;
  assign new_n1253_ = pv78_1_ & ~pv78_0_;
  assign new_n1254_ = ~pv78_1_ & pv78_0_;
  assign new_n1255_ = ~new_n1253_ & ~new_n1254_;
  assign new_n1256_ = pv78_3_ & ~pv78_2_;
  assign new_n1257_ = ~pv78_3_ & pv78_2_;
  assign new_n1258_ = ~new_n1256_ & ~new_n1257_;
  assign new_n1259_ = new_n1255_ & ~new_n1258_;
  assign new_n1260_ = ~new_n1255_ & new_n1258_;
  assign new_n1261_ = ~new_n1259_ & ~new_n1260_;
  assign new_n1262_ = pv78_5_ & ~pv78_4_;
  assign new_n1263_ = ~pv78_5_ & pv78_4_;
  assign new_n1264_ = ~new_n1262_ & ~new_n1263_;
  assign new_n1265_ = ~pv84_0_ & pv84_1_;
  assign new_n1266_ = pv84_0_ & ~pv84_1_;
  assign new_n1267_ = ~new_n1265_ & ~new_n1266_;
  assign new_n1268_ = new_n1264_ & ~new_n1267_;
  assign new_n1269_ = ~new_n1264_ & new_n1267_;
  assign new_n1270_ = ~new_n1268_ & ~new_n1269_;
  assign new_n1271_ = new_n1261_ & ~new_n1270_;
  assign new_n1272_ = ~new_n1261_ & new_n1270_;
  assign new_n1273_ = ~new_n1271_ & ~new_n1272_;
  assign new_n1274_ = pv94_0_ & new_n1273_;
  assign new_n1275_ = ~pv94_0_ & ~new_n1273_;
  assign new_n1276_ = ~new_n1274_ & ~new_n1275_;
  assign new_n1277_ = ~new_n1252_ & ~new_n1276_;
  assign new_n1278_ = ~new_n1230_ & ~new_n1277_;
  assign new_n1279_ = new_n1223_ & ~new_n1278_;
  assign new_n1280_ = new_n546_ & ~new_n554_;
  assign new_n1281_ = ~new_n491_ & ~new_n1279_;
  assign new_n1282_ = ~new_n494_ & new_n1281_;
  assign new_n1283_ = ~new_n575_ & ~new_n1280_;
  assign new_n1284_ = new_n1282_ & new_n1283_;
  assign new_n1285_ = pv56_0_ & ~new_n1284_;
  assign new_n1286_ = pv56_0_ & ~new_n1134_;
  assign new_n1287_ = ~new_n1221_ & ~new_n1222_;
  assign new_n1288_ = ~new_n1285_ & ~new_n1286_;
  assign pv508_0_ = ~new_n1287_ | ~new_n1288_;
  assign pv539 = new_n491_ & pv1213_2_;
  assign new_n1291_ = pv257_1_ & new_n637_;
  assign new_n1292_ = pv229_0_ & new_n641_;
  assign new_n1293_ = pv189_0_ & new_n643_;
  assign new_n1294_ = ~new_n1292_ & ~new_n1293_;
  assign new_n1295_ = new_n647_ & ~new_n1294_;
  assign new_n1296_ = ~new_n1291_ & ~new_n1295_;
  assign new_n1297_ = ~new_n624_ & ~new_n1296_;
  assign new_n1298_ = new_n624_ & new_n653_;
  assign new_n1299_ = ~new_n1297_ & ~new_n1298_;
  assign new_n1300_ = new_n658_ & ~new_n1299_;
  assign new_n1301_ = pv32_6_ & new_n660_;
  assign pv1213_6_ = new_n1300_ | new_n1301_;
  assign new_n1303_ = pv268_5_ & new_n686_;
  assign new_n1304_ = pv268_2_ & ~new_n1303_;
  assign new_n1305_ = ~pv268_2_ & new_n1303_;
  assign pv1372 = new_n1304_ | new_n1305_;
  assign pv1440_0_ = ~pv14_0_ | new_n507_;
  assign new_n1308_ = pv16_0_ & ~pv15_0_;
  assign pv1758_0_ = new_n1152_ | new_n1308_;
  assign new_n1310_ = pv257_5_ & new_n637_;
  assign new_n1311_ = pv229_4_ & new_n641_;
  assign new_n1312_ = pv189_4_ & new_n643_;
  assign new_n1313_ = ~new_n1311_ & ~new_n1312_;
  assign new_n1314_ = new_n647_ & ~new_n1313_;
  assign new_n1315_ = ~new_n1310_ & ~new_n1314_;
  assign new_n1316_ = ~new_n624_ & ~new_n1315_;
  assign new_n1317_ = pv32_0_ & new_n653_;
  assign new_n1318_ = pv32_3_ & ~new_n653_;
  assign new_n1319_ = ~new_n1317_ & ~new_n1318_;
  assign new_n1320_ = new_n624_ & ~new_n1319_;
  assign new_n1321_ = ~new_n1316_ & ~new_n1320_;
  assign new_n1322_ = new_n658_ & ~new_n1321_;
  assign new_n1323_ = pv32_10_ & new_n660_;
  assign pv1213_10_ = new_n1322_ | new_n1323_;
  assign new_n1325_ = ~new_n572_ & ~pv1213_10_;
  assign new_n1326_ = ~pv78_2_ & new_n572_;
  assign pv1781_0_ = new_n1325_ | new_n1326_;
  assign new_n1328_ = pv234_1_ & new_n641_;
  assign new_n1329_ = pv194_1_ & new_n643_;
  assign new_n1330_ = ~new_n1328_ & ~new_n1329_;
  assign new_n1331_ = new_n647_ & ~new_n1330_;
  assign new_n1332_ = pv149_5_ & new_n665_;
  assign new_n1333_ = new_n633_ & new_n1332_;
  assign new_n1334_ = ~new_n1331_ & ~new_n1333_;
  assign new_n1335_ = ~new_n624_ & ~new_n1334_;
  assign new_n1336_ = pv32_3_ & new_n653_;
  assign new_n1337_ = pv32_6_ & ~new_n653_;
  assign new_n1338_ = ~new_n1336_ & ~new_n1337_;
  assign new_n1339_ = new_n624_ & ~new_n1338_;
  assign new_n1340_ = ~new_n1335_ & ~new_n1339_;
  assign new_n1341_ = new_n658_ & ~new_n1340_;
  assign new_n1342_ = pv78_5_ & new_n660_;
  assign pv1243_1_ = new_n1341_ | new_n1342_;
  assign new_n1344_ = pv37_0_ & ~pv1243_1_;
  assign new_n1345_ = pv223_4_ & new_n641_;
  assign new_n1346_ = pv183_4_ & new_n643_;
  assign new_n1347_ = ~new_n1345_ & ~new_n1346_;
  assign new_n1348_ = new_n647_ & ~new_n1347_;
  assign new_n1349_ = ~new_n1155_ & ~new_n1348_;
  assign new_n1350_ = new_n658_ & ~new_n1349_;
  assign new_n1351_ = ~new_n624_ & new_n1350_;
  assign new_n1352_ = ~new_n624_ & new_n1351_;
  assign new_n1353_ = pv32_4_ & new_n660_;
  assign pv1213_4_ = new_n1352_ | new_n1353_;
  assign new_n1355_ = ~pv37_0_ & ~pv1213_4_;
  assign pv1829_1_ = new_n1344_ | new_n1355_;
  assign new_n1357_ = pv257_2_ & new_n637_;
  assign new_n1358_ = pv229_1_ & new_n641_;
  assign new_n1359_ = pv189_1_ & new_n643_;
  assign new_n1360_ = ~new_n1358_ & ~new_n1359_;
  assign new_n1361_ = new_n647_ & ~new_n1360_;
  assign new_n1362_ = ~new_n1357_ & ~new_n1361_;
  assign new_n1363_ = ~new_n624_ & ~new_n1362_;
  assign new_n1364_ = pv32_0_ & ~new_n653_;
  assign new_n1365_ = ~new_n653_ & ~new_n1364_;
  assign new_n1366_ = new_n624_ & ~new_n1365_;
  assign new_n1367_ = ~new_n1363_ & ~new_n1366_;
  assign new_n1368_ = new_n658_ & ~new_n1367_;
  assign new_n1369_ = pv32_7_ & new_n660_;
  assign pv1213_7_ = new_n1368_ | new_n1369_;
  assign new_n1371_ = new_n507_ & ~pv802_0_;
  assign new_n1372_ = pv248_0_ & ~pv802_0_;
  assign new_n1373_ = pv194_3_ & pv194_1_;
  assign new_n1374_ = pv199_2_ & new_n1373_;
  assign new_n1375_ = pv199_0_ & new_n1374_;
  assign new_n1376_ = pv199_4_ & new_n1375_;
  assign new_n1377_ = pv199_1_ & new_n1376_;
  assign new_n1378_ = pv199_3_ & new_n1377_;
  assign new_n1379_ = pv194_2_ & new_n1378_;
  assign new_n1380_ = pv194_4_ & new_n1379_;
  assign new_n1381_ = pv194_0_ & new_n1380_;
  assign new_n1382_ = ~pv802_0_ & new_n1381_;
  assign new_n1383_ = ~new_n1371_ & ~new_n1372_;
  assign new_n1384_ = ~new_n1382_ & new_n1383_;
  assign new_n1385_ = ~new_n639_ & new_n1384_;
  assign new_n1386_ = ~new_n740_ & new_n1385_;
  assign new_n1387_ = ~pv274_0_ & pv271_0_;
  assign new_n1388_ = ~new_n572_ & new_n1387_;
  assign new_n1389_ = pv134_1_ & pv134_0_;
  assign new_n1390_ = new_n1388_ & new_n1389_;
  assign new_n1391_ = new_n507_ & new_n1390_;
  assign new_n1392_ = ~new_n1381_ & new_n1391_;
  assign new_n1393_ = new_n573_ & ~pv802_0_;
  assign new_n1394_ = ~new_n1372_ & new_n1393_;
  assign new_n1395_ = ~new_n507_ & new_n1394_;
  assign new_n1396_ = ~new_n740_ & new_n1395_;
  assign new_n1397_ = ~new_n1381_ & new_n1396_;
  assign new_n1398_ = ~new_n1386_ & ~new_n1392_;
  assign new_n1399_ = ~new_n1397_ & new_n1398_;
  assign new_n1400_ = pv7_0_ & ~new_n1399_;
  assign pv1380 = new_n692_ & new_n1400_;
  assign new_n1402_ = new_n510_ & new_n1308_;
  assign new_n1403_ = new_n490_ & new_n1308_;
  assign new_n1404_ = pv56_0_ & new_n1093_;
  assign new_n1405_ = pv14_0_ & ~new_n1404_;
  assign new_n1406_ = pv101_0_ & new_n1405_;
  assign new_n1407_ = ~new_n1402_ & ~new_n1403_;
  assign pv1759_0_ = new_n1406_ | ~new_n1407_;
  assign new_n1409_ = pv234_4_ & new_n641_;
  assign new_n1410_ = pv194_4_ & new_n643_;
  assign new_n1411_ = ~new_n1409_ & ~new_n1410_;
  assign new_n1412_ = ~new_n624_ & ~new_n635_;
  assign new_n1413_ = ~new_n1411_ & new_n1412_;
  assign new_n1414_ = new_n616_ & new_n1413_;
  assign new_n1415_ = ~new_n633_ & new_n1414_;
  assign new_n1416_ = ~new_n624_ & new_n1415_;
  assign new_n1417_ = pv32_6_ & new_n653_;
  assign new_n1418_ = pv32_9_ & ~new_n653_;
  assign new_n1419_ = ~new_n1417_ & ~new_n1418_;
  assign new_n1420_ = new_n624_ & ~new_n1419_;
  assign new_n1421_ = ~new_n1416_ & ~new_n1420_;
  assign new_n1422_ = new_n658_ & ~new_n1421_;
  assign new_n1423_ = pv84_2_ & new_n660_;
  assign pv1243_4_ = new_n1422_ | new_n1423_;
  assign new_n1425_ = pv37_0_ & ~pv1243_4_;
  assign new_n1426_ = ~pv37_0_ & ~pv1213_7_;
  assign pv1829_4_ = new_n1425_ | new_n1426_;
  assign new_n1428_ = pv257_6_ & ~pv257_7_;
  assign new_n1429_ = ~pv257_6_ & pv257_7_;
  assign pv656 = new_n1428_ | new_n1429_;
  assign pv779 = pv6_0_ & new_n692_;
  assign new_n1432_ = pv257_3_ & new_n637_;
  assign new_n1433_ = pv229_2_ & new_n641_;
  assign new_n1434_ = pv189_2_ & new_n643_;
  assign new_n1435_ = ~new_n1433_ & ~new_n1434_;
  assign new_n1436_ = new_n647_ & ~new_n1435_;
  assign new_n1437_ = ~new_n1432_ & ~new_n1436_;
  assign new_n1438_ = ~new_n624_ & ~new_n1437_;
  assign new_n1439_ = pv32_1_ & ~new_n653_;
  assign new_n1440_ = ~new_n653_ & ~new_n1439_;
  assign new_n1441_ = new_n624_ & ~new_n1440_;
  assign new_n1442_ = ~new_n1438_ & ~new_n1441_;
  assign new_n1443_ = new_n658_ & ~new_n1442_;
  assign new_n1444_ = pv32_8_ & new_n660_;
  assign pv1213_8_ = new_n1443_ | new_n1444_;
  assign pv1262 = pv4_0_ & new_n692_;
  assign new_n1447_ = pv268_4_ & pv268_2_;
  assign new_n1448_ = pv268_3_ & new_n1447_;
  assign new_n1449_ = pv268_1_ & new_n1448_;
  assign new_n1450_ = pv268_5_ & new_n1449_;
  assign new_n1451_ = pv268_0_ & ~new_n1450_;
  assign new_n1452_ = ~pv268_0_ & new_n1450_;
  assign pv1370 = new_n1451_ | new_n1452_;
  assign new_n1454_ = pv234_3_ & new_n641_;
  assign new_n1455_ = pv194_3_ & new_n643_;
  assign new_n1456_ = ~new_n1454_ & ~new_n1455_;
  assign new_n1457_ = new_n647_ & ~new_n1456_;
  assign new_n1458_ = pv149_7_ & new_n665_;
  assign new_n1459_ = new_n633_ & new_n1458_;
  assign new_n1460_ = ~new_n1457_ & ~new_n1459_;
  assign new_n1461_ = ~new_n624_ & ~new_n1460_;
  assign new_n1462_ = pv32_5_ & new_n653_;
  assign new_n1463_ = pv32_8_ & ~new_n653_;
  assign new_n1464_ = ~new_n1462_ & ~new_n1463_;
  assign new_n1465_ = new_n624_ & ~new_n1464_;
  assign new_n1466_ = ~new_n1461_ & ~new_n1465_;
  assign new_n1467_ = new_n658_ & ~new_n1466_;
  assign new_n1468_ = pv84_1_ & new_n660_;
  assign pv1243_3_ = new_n1467_ | new_n1468_;
  assign new_n1470_ = pv37_0_ & ~pv1243_3_;
  assign new_n1471_ = ~pv37_0_ & ~pv1213_6_;
  assign pv1829_3_ = new_n1470_ | new_n1471_;
  assign new_n1473_ = pv257_4_ & new_n637_;
  assign new_n1474_ = pv229_3_ & new_n641_;
  assign new_n1475_ = pv189_3_ & new_n643_;
  assign new_n1476_ = ~new_n1474_ & ~new_n1475_;
  assign new_n1477_ = new_n647_ & ~new_n1476_;
  assign new_n1478_ = ~new_n1473_ & ~new_n1477_;
  assign new_n1479_ = ~new_n624_ & ~new_n1478_;
  assign new_n1480_ = pv32_2_ & ~new_n653_;
  assign new_n1481_ = ~new_n653_ & ~new_n1480_;
  assign new_n1482_ = new_n624_ & ~new_n1481_;
  assign new_n1483_ = ~new_n1479_ & ~new_n1482_;
  assign new_n1484_ = new_n658_ & ~new_n1483_;
  assign new_n1485_ = pv32_9_ & new_n660_;
  assign pv1213_9_ = new_n1484_ | new_n1485_;
  assign pv1264 = pv4_0_ & pv12_0_;
  assign pv1265 = pv52_0_ & pv1264;
  assign new_n1489_ = ~pv56_0_ & ~pv50_0_;
  assign new_n1490_ = ~pv62_0_ & new_n1489_;
  assign new_n1491_ = ~new_n616_ & ~new_n1490_;
  assign pv1386 = pv782 & new_n1491_;
  assign new_n1493_ = ~pv280_0_ & new_n494_;
  assign new_n1494_ = pv165_2_ & pv165_1_;
  assign new_n1495_ = ~pv165_0_ & new_n1494_;
  assign new_n1496_ = pv203_0_ & new_n1495_;
  assign new_n1497_ = pv240_0_ & ~new_n1493_;
  assign new_n1498_ = ~new_n1496_ & new_n1497_;
  assign new_n1499_ = new_n758_ & new_n1498_;
  assign new_n1500_ = ~new_n699_ & new_n1499_;
  assign new_n1501_ = ~pv172_0_ & new_n1500_;
  assign new_n1502_ = ~new_n507_ & ~new_n640_;
  assign new_n1503_ = ~new_n494_ & ~new_n1502_;
  assign new_n1504_ = pv802_0_ & ~new_n1503_;
  assign pv1717_0_ = new_n1501_ | new_n1504_;
  assign new_n1506_ = pv239_1_ & new_n641_;
  assign new_n1507_ = pv199_1_ & new_n643_;
  assign new_n1508_ = ~new_n1506_ & ~new_n1507_;
  assign new_n1509_ = new_n1412_ & ~new_n1508_;
  assign new_n1510_ = new_n616_ & new_n1509_;
  assign new_n1511_ = ~new_n633_ & new_n1510_;
  assign new_n1512_ = ~new_n624_ & new_n1511_;
  assign new_n1513_ = pv32_8_ & new_n653_;
  assign new_n1514_ = pv32_11_ & ~new_n653_;
  assign new_n1515_ = ~new_n1513_ & ~new_n1514_;
  assign new_n1516_ = new_n624_ & ~new_n1515_;
  assign new_n1517_ = ~new_n1512_ & ~new_n1516_;
  assign new_n1518_ = new_n658_ & ~new_n1517_;
  assign new_n1519_ = pv84_4_ & new_n660_;
  assign pv1243_6_ = new_n1518_ | new_n1519_;
  assign new_n1521_ = pv37_0_ & ~pv1243_6_;
  assign new_n1522_ = ~pv37_0_ & ~pv1213_9_;
  assign pv1829_6_ = new_n1521_ | new_n1522_;
  assign new_n1524_ = ~pv202_0_ & ~pv271_0_;
  assign new_n1525_ = pv274_0_ & new_n1524_;
  assign new_n1526_ = pv274_0_ & ~new_n1525_;
  assign new_n1527_ = ~pv271_0_ & new_n1526_;
  assign new_n1528_ = pv269_0_ & ~new_n1525_;
  assign new_n1529_ = pv271_0_ & new_n1528_;
  assign pv634_0_ = ~new_n1527_ & ~new_n1529_;
  assign new_n1531_ = new_n493_ & pv1757_0_;
  assign new_n1532_ = pv802_0_ & new_n1531_;
  assign new_n1533_ = ~new_n493_ & pv1757_0_;
  assign new_n1534_ = ~new_n1278_ & ~new_n1532_;
  assign pv1480_0_ = new_n1533_ | ~new_n1534_;
  assign new_n1536_ = ~new_n699_ & new_n707_;
  assign new_n1537_ = ~new_n699_ & new_n717_;
  assign new_n1538_ = pv290_0_ & new_n699_;
  assign new_n1539_ = ~new_n699_ & new_n722_;
  assign new_n1540_ = ~new_n725_ & ~new_n1536_;
  assign new_n1541_ = ~new_n1537_ & new_n1540_;
  assign new_n1542_ = ~new_n1538_ & ~new_n1539_;
  assign pv1741_0_ = ~new_n1541_ | ~new_n1542_;
  assign new_n1544_ = pv239_0_ & new_n641_;
  assign new_n1545_ = pv199_0_ & new_n643_;
  assign new_n1546_ = ~new_n1544_ & ~new_n1545_;
  assign new_n1547_ = new_n1412_ & ~new_n1546_;
  assign new_n1548_ = new_n616_ & new_n1547_;
  assign new_n1549_ = ~new_n633_ & new_n1548_;
  assign new_n1550_ = ~new_n624_ & new_n1549_;
  assign new_n1551_ = pv32_7_ & new_n653_;
  assign new_n1552_ = pv32_10_ & ~new_n653_;
  assign new_n1553_ = ~new_n1551_ & ~new_n1552_;
  assign new_n1554_ = new_n624_ & ~new_n1553_;
  assign new_n1555_ = ~new_n1550_ & ~new_n1554_;
  assign new_n1556_ = new_n658_ & ~new_n1555_;
  assign new_n1557_ = pv84_3_ & new_n660_;
  assign pv1243_5_ = new_n1556_ | new_n1557_;
  assign new_n1559_ = pv37_0_ & ~pv1243_5_;
  assign new_n1560_ = ~pv37_0_ & ~pv1213_8_;
  assign pv1829_5_ = new_n1559_ | new_n1560_;
  assign new_n1562_ = pv39_0_ & ~pv38_0_;
  assign new_n1563_ = ~pv39_0_ & pv38_0_;
  assign new_n1564_ = ~new_n1562_ & ~new_n1563_;
  assign new_n1565_ = pv42_0_ & ~pv44_0_;
  assign new_n1566_ = ~pv42_0_ & pv44_0_;
  assign new_n1567_ = ~new_n1565_ & ~new_n1566_;
  assign pv512 = new_n1564_ & new_n1567_;
  assign pv783 = pv5_0_ & pv11_0_;
  assign pv1256 = pv2_0_ & new_n692_;
  assign pv1267 = pv2_0_ & pv11_0_;
  assign new_n1572_ = ~pv302_0_ & new_n493_;
  assign new_n1573_ = new_n511_ & new_n554_;
  assign new_n1574_ = ~new_n1572_ & ~new_n1573_;
  assign new_n1575_ = ~new_n712_ & ~new_n713_;
  assign new_n1576_ = new_n1574_ & new_n1575_;
  assign new_n1577_ = ~new_n699_ & new_n704_;
  assign new_n1578_ = ~pv289_0_ & new_n1577_;
  assign new_n1579_ = ~new_n1576_ & new_n1578_;
  assign new_n1580_ = pv14_0_ & new_n1579_;
  assign new_n1581_ = ~new_n585_ & ~new_n1580_;
  assign new_n1582_ = ~new_n699_ & new_n1581_;
  assign new_n1583_ = new_n704_ & new_n1582_;
  assign new_n1584_ = new_n490_ & new_n1583_;
  assign new_n1585_ = pv290_0_ & new_n490_;
  assign new_n1586_ = new_n699_ & new_n1585_;
  assign new_n1587_ = ~new_n1584_ & ~new_n1586_;
  assign new_n1588_ = ~pv149_6_ & new_n761_;
  assign new_n1589_ = pv56_0_ & new_n1588_;
  assign new_n1590_ = pv14_0_ & new_n1587_;
  assign new_n1591_ = pv213_0_ & new_n1590_;
  assign new_n1592_ = ~new_n1589_ & new_n1591_;
  assign new_n1593_ = ~pv165_3_ & new_n577_;
  assign new_n1594_ = ~pv165_7_ & new_n1593_;
  assign new_n1595_ = ~new_n704_ & ~new_n1594_;
  assign new_n1596_ = ~new_n1587_ & ~new_n1595_;
  assign pv1281_0_ = new_n1592_ | new_n1596_;
  assign new_n1598_ = pv268_4_ & pv268_5_;
  assign new_n1599_ = pv268_3_ & ~new_n1598_;
  assign new_n1600_ = ~pv268_3_ & new_n1598_;
  assign pv1373 = new_n1599_ | new_n1600_;
  assign new_n1602_ = pv56_0_ & ~new_n1278_;
  assign new_n1603_ = new_n1224_ & new_n1602_;
  assign new_n1604_ = ~new_n699_ & new_n1603_;
  assign pv1384 = pv782 & new_n1604_;
  assign new_n1606_ = pv239_3_ & new_n641_;
  assign new_n1607_ = pv199_3_ & new_n643_;
  assign new_n1608_ = ~new_n1606_ & ~new_n1607_;
  assign new_n1609_ = new_n1412_ & ~new_n1608_;
  assign new_n1610_ = new_n616_ & new_n1609_;
  assign new_n1611_ = ~new_n633_ & new_n1610_;
  assign new_n1612_ = ~new_n624_ & new_n1611_;
  assign new_n1613_ = pv32_10_ & new_n624_;
  assign new_n1614_ = new_n624_ & new_n1613_;
  assign new_n1615_ = new_n653_ & new_n1614_;
  assign new_n1616_ = ~new_n1612_ & ~new_n1615_;
  assign new_n1617_ = new_n658_ & ~new_n1616_;
  assign new_n1618_ = pv88_0_ & new_n660_;
  assign pv1243_8_ = new_n1617_ | new_n1618_;
  assign new_n1620_ = pv37_0_ & ~pv1243_8_;
  assign new_n1621_ = ~pv37_0_ & ~pv1213_11_;
  assign pv1829_8_ = new_n1620_ | new_n1621_;
  assign new_n1623_ = pv132_0_ & new_n1098_;
  assign new_n1624_ = new_n1093_ & ~new_n1095_;
  assign new_n1625_ = ~new_n1096_ & new_n1624_;
  assign new_n1626_ = pv108_5_ & new_n1625_;
  assign pv1953_0_ = new_n1623_ | new_n1626_;
  assign new_n1628_ = pv14_0_ & new_n758_;
  assign new_n1629_ = ~new_n615_ & new_n1628_;
  assign new_n1630_ = pv763 & new_n1629_;
  assign pv775 = pv70_0_ & new_n1630_;
  assign pv784 = pv7_0_ & pv11_0_;
  assign new_n1633_ = ~pv57_0_ & new_n1223_;
  assign new_n1634_ = ~new_n494_ & new_n545_;
  assign new_n1635_ = new_n505_ & new_n1634_;
  assign new_n1636_ = ~new_n491_ & ~new_n546_;
  assign new_n1637_ = new_n772_ & new_n1636_;
  assign new_n1638_ = new_n1635_ & new_n1637_;
  assign new_n1639_ = pv57_0_ & ~new_n1638_;
  assign new_n1640_ = ~pv60_0_ & ~pv63_0_;
  assign new_n1641_ = new_n572_ & ~new_n1640_;
  assign new_n1642_ = ~new_n1633_ & ~new_n1639_;
  assign new_n1643_ = pv12_0_ & new_n1642_;
  assign new_n1644_ = ~pv174_0_ & new_n1643_;
  assign new_n1645_ = pv2_0_ & new_n1644_;
  assign new_n1646_ = ~new_n1641_ & new_n1645_;
  assign pv1257 = ~pv35_0_ & new_n1646_;
  assign pv1266 = pv4_0_ & pv11_0_;
  assign new_n1649_ = ~new_n712_ & ~new_n785_;
  assign new_n1650_ = new_n758_ & new_n1649_;
  assign new_n1651_ = ~new_n1223_ & new_n1650_;
  assign new_n1652_ = pv14_0_ & new_n1651_;
  assign new_n1653_ = pv62_0_ & new_n1652_;
  assign new_n1654_ = new_n505_ & new_n1653_;
  assign new_n1655_ = ~new_n1133_ & new_n1654_;
  assign new_n1656_ = new_n616_ & new_n1655_;
  assign pv1365 = ~new_n1213_ & new_n1656_;
  assign new_n1658_ = pv268_4_ & ~pv268_5_;
  assign new_n1659_ = ~pv268_4_ & pv268_5_;
  assign pv1374 = new_n1658_ | new_n1659_;
  assign new_n1661_ = ~pv258_0_ & new_n1491_;
  assign new_n1662_ = pv268_0_ & new_n1450_;
  assign new_n1663_ = pv258_0_ & new_n1662_;
  assign new_n1664_ = ~new_n1661_ & ~new_n1663_;
  assign new_n1665_ = pv14_0_ & new_n1664_;
  assign new_n1666_ = pv259_0_ & new_n1665_;
  assign new_n1667_ = pv14_0_ & ~new_n1664_;
  assign new_n1668_ = ~pv259_0_ & new_n1667_;
  assign pv1459_0_ = new_n1666_ | new_n1668_;
  assign new_n1670_ = pv239_2_ & new_n641_;
  assign new_n1671_ = pv199_2_ & new_n643_;
  assign new_n1672_ = ~new_n1670_ & ~new_n1671_;
  assign new_n1673_ = new_n1412_ & ~new_n1672_;
  assign new_n1674_ = new_n616_ & new_n1673_;
  assign new_n1675_ = ~new_n633_ & new_n1674_;
  assign new_n1676_ = ~new_n624_ & new_n1675_;
  assign new_n1677_ = pv32_9_ & new_n624_;
  assign new_n1678_ = new_n624_ & new_n1677_;
  assign new_n1679_ = new_n653_ & new_n1678_;
  assign new_n1680_ = ~new_n1676_ & ~new_n1679_;
  assign new_n1681_ = new_n658_ & ~new_n1680_;
  assign new_n1682_ = pv84_5_ & new_n660_;
  assign pv1243_7_ = new_n1681_ | new_n1682_;
  assign new_n1684_ = pv37_0_ & ~pv1243_7_;
  assign new_n1685_ = ~pv37_0_ & ~pv1213_10_;
  assign pv1829_7_ = new_n1684_ | new_n1685_;
  assign pv1953_1_ = pv132_1_ & new_n1098_;
  assign pv543 = new_n491_ & pv1213_6_;
  assign new_n1689_ = pv802_0_ & ~new_n640_;
  assign pv587 = ~pv243_0_ & ~new_n1689_;
  assign new_n1691_ = pv257_2_ & pv257_4_;
  assign new_n1692_ = pv257_5_ & new_n1691_;
  assign new_n1693_ = pv257_3_ & new_n1692_;
  assign new_n1694_ = pv257_7_ & new_n1693_;
  assign new_n1695_ = pv257_6_ & new_n1694_;
  assign new_n1696_ = pv257_1_ & ~new_n1695_;
  assign new_n1697_ = ~pv257_1_ & new_n1695_;
  assign pv651 = new_n1696_ | new_n1697_;
  assign new_n1699_ = pv56_0_ & ~new_n586_;
  assign new_n1700_ = ~pv174_0_ & new_n1699_;
  assign new_n1701_ = ~pv52_0_ & ~new_n1700_;
  assign new_n1702_ = pv6_0_ & pv12_0_;
  assign pv781 = ~new_n1701_ & new_n1702_;
  assign new_n1704_ = pv14_0_ & ~new_n1586_;
  assign new_n1705_ = pv213_2_ & new_n1704_;
  assign new_n1706_ = ~new_n1589_ & new_n1705_;
  assign new_n1707_ = pv165_4_ & new_n1586_;
  assign pv1297_1_ = new_n1706_ | new_n1707_;
  assign new_n1709_ = ~pv88_2_ & new_n572_;
  assign new_n1710_ = ~pv134_0_ & ~new_n572_;
  assign pv1771_0_ = new_n1709_ | new_n1710_;
  assign new_n1712_ = pv149_7_ & new_n839_;
  assign new_n1713_ = ~pv149_6_ & new_n1712_;
  assign new_n1714_ = pv56_0_ & new_n1713_;
  assign new_n1715_ = pv108_4_ & ~new_n1714_;
  assign pv1900_0_ = new_n1152_ | new_n1715_;
  assign new_n1717_ = ~pv149_7_ & new_n760_;
  assign new_n1718_ = pv149_6_ & new_n1717_;
  assign new_n1719_ = ~new_n1095_ & ~new_n1713_;
  assign new_n1720_ = new_n1718_ & new_n1719_;
  assign new_n1721_ = ~new_n1588_ & new_n1720_;
  assign new_n1722_ = pv100_1_ & new_n1721_;
  assign new_n1723_ = new_n1095_ & ~new_n1713_;
  assign new_n1724_ = ~new_n1718_ & new_n1723_;
  assign new_n1725_ = ~new_n1588_ & new_n1724_;
  assign new_n1726_ = pv124_1_ & new_n1725_;
  assign new_n1727_ = ~new_n1718_ & new_n1719_;
  assign new_n1728_ = new_n1588_ & new_n1727_;
  assign new_n1729_ = pv213_1_ & new_n1728_;
  assign new_n1730_ = ~new_n1095_ & new_n1713_;
  assign new_n1731_ = ~new_n1718_ & new_n1730_;
  assign new_n1732_ = ~new_n1588_ & new_n1731_;
  assign new_n1733_ = pv108_1_ & new_n1732_;
  assign new_n1734_ = ~new_n1722_ & ~new_n1726_;
  assign new_n1735_ = ~new_n1729_ & ~new_n1733_;
  assign pv1921_1_ = ~new_n1734_ | ~new_n1735_;
  assign new_n1737_ = pv239_4_ & new_n641_;
  assign new_n1738_ = pv199_4_ & new_n643_;
  assign new_n1739_ = ~new_n1737_ & ~new_n1738_;
  assign new_n1740_ = new_n1412_ & ~new_n1739_;
  assign new_n1741_ = new_n616_ & new_n1740_;
  assign new_n1742_ = ~new_n633_ & new_n1741_;
  assign new_n1743_ = ~new_n624_ & new_n1742_;
  assign new_n1744_ = pv32_11_ & new_n624_;
  assign new_n1745_ = new_n624_ & new_n1744_;
  assign new_n1746_ = new_n653_ & new_n1745_;
  assign new_n1747_ = ~new_n1743_ & ~new_n1746_;
  assign new_n1748_ = new_n658_ & ~new_n1747_;
  assign new_n1749_ = pv88_1_ & new_n660_;
  assign pv1243_9_ = new_n1748_ | new_n1749_;
  assign new_n1751_ = ~pv1213_2_ & ~pv1213_0_;
  assign new_n1752_ = ~pv1213_3_ & new_n1751_;
  assign new_n1753_ = ~pv1213_1_ & new_n1752_;
  assign new_n1754_ = ~new_n842_ & new_n1753_;
  assign new_n1755_ = ~new_n880_ & new_n1754_;
  assign new_n1756_ = pv1213_3_ & new_n1751_;
  assign new_n1757_ = ~pv1213_1_ & new_n1756_;
  assign new_n1758_ = ~new_n842_ & new_n1757_;
  assign new_n1759_ = pv288_6_ & new_n1758_;
  assign new_n1760_ = ~new_n1755_ & ~new_n1759_;
  assign new_n1761_ = new_n616_ & new_n1760_;
  assign new_n1762_ = new_n616_ & new_n1084_;
  assign new_n1763_ = new_n1761_ & new_n1762_;
  assign new_n1764_ = pv288_6_ & pv288_7_;
  assign new_n1765_ = ~new_n1763_ & new_n1764_;
  assign new_n1766_ = new_n957_ & ~new_n973_;
  assign new_n1767_ = new_n959_ & ~new_n988_;
  assign new_n1768_ = ~new_n959_ & ~new_n988_;
  assign new_n1769_ = ~new_n1767_ & ~new_n1768_;
  assign new_n1770_ = new_n959_ & ~new_n982_;
  assign new_n1771_ = new_n988_ & ~new_n1015_;
  assign new_n1772_ = ~new_n988_ & new_n1015_;
  assign new_n1773_ = ~new_n1771_ & ~new_n1772_;
  assign new_n1774_ = ~new_n959_ & ~new_n1773_;
  assign new_n1775_ = ~new_n1770_ & ~new_n1774_;
  assign new_n1776_ = new_n1769_ & new_n1775_;
  assign new_n1777_ = new_n959_ & ~new_n997_;
  assign new_n1778_ = ~new_n1023_ & ~new_n1772_;
  assign new_n1779_ = new_n1023_ & new_n1772_;
  assign new_n1780_ = ~new_n1778_ & ~new_n1779_;
  assign new_n1781_ = ~new_n959_ & ~new_n1780_;
  assign new_n1782_ = ~new_n1777_ & ~new_n1781_;
  assign new_n1783_ = new_n1776_ & new_n1782_;
  assign new_n1784_ = new_n959_ & ~new_n973_;
  assign new_n1785_ = ~new_n1010_ & ~new_n1779_;
  assign new_n1786_ = new_n1010_ & new_n1779_;
  assign new_n1787_ = ~new_n1785_ & ~new_n1786_;
  assign new_n1788_ = ~new_n959_ & ~new_n1787_;
  assign new_n1789_ = ~new_n1784_ & ~new_n1788_;
  assign new_n1790_ = ~new_n1783_ & ~new_n1789_;
  assign new_n1791_ = new_n1783_ & new_n1789_;
  assign new_n1792_ = ~new_n1790_ & ~new_n1791_;
  assign new_n1793_ = ~new_n957_ & ~new_n1792_;
  assign new_n1794_ = ~new_n1766_ & ~new_n1793_;
  assign new_n1795_ = ~pv1213_0_ & ~new_n1794_;
  assign new_n1796_ = pv1213_0_ & new_n1794_;
  assign new_n1797_ = ~new_n1795_ & ~new_n1796_;
  assign new_n1798_ = new_n957_ & ~new_n982_;
  assign new_n1799_ = ~new_n1769_ & ~new_n1775_;
  assign new_n1800_ = ~new_n1776_ & ~new_n1799_;
  assign new_n1801_ = ~new_n957_ & ~new_n1800_;
  assign new_n1802_ = ~new_n1798_ & ~new_n1801_;
  assign new_n1803_ = ~pv1213_2_ & ~new_n1802_;
  assign new_n1804_ = pv1213_2_ & new_n1802_;
  assign new_n1805_ = ~new_n1803_ & ~new_n1804_;
  assign new_n1806_ = new_n957_ & ~new_n988_;
  assign new_n1807_ = ~new_n957_ & new_n1769_;
  assign new_n1808_ = ~new_n1806_ & ~new_n1807_;
  assign new_n1809_ = ~pv1213_3_ & ~new_n1808_;
  assign new_n1810_ = pv1213_3_ & new_n1808_;
  assign new_n1811_ = ~new_n1809_ & ~new_n1810_;
  assign new_n1812_ = new_n957_ & ~new_n997_;
  assign new_n1813_ = ~new_n1776_ & ~new_n1782_;
  assign new_n1814_ = ~new_n1783_ & ~new_n1813_;
  assign new_n1815_ = ~new_n957_ & ~new_n1814_;
  assign new_n1816_ = ~new_n1812_ & ~new_n1815_;
  assign new_n1817_ = ~pv1213_1_ & ~new_n1816_;
  assign new_n1818_ = pv1213_1_ & new_n1816_;
  assign new_n1819_ = ~new_n1817_ & ~new_n1818_;
  assign new_n1820_ = ~pv288_0_ & ~pv288_1_;
  assign new_n1821_ = new_n1797_ & new_n1805_;
  assign new_n1822_ = new_n1811_ & new_n1821_;
  assign new_n1823_ = new_n1819_ & new_n1822_;
  assign new_n1824_ = ~new_n842_ & new_n1823_;
  assign new_n1825_ = ~new_n1820_ & new_n1824_;
  assign new_n1826_ = ~pv1213_0_ & ~new_n1789_;
  assign new_n1827_ = pv1213_0_ & new_n1789_;
  assign new_n1828_ = ~new_n1826_ & ~new_n1827_;
  assign new_n1829_ = ~pv1213_2_ & ~new_n1775_;
  assign new_n1830_ = pv1213_2_ & new_n1775_;
  assign new_n1831_ = ~new_n1829_ & ~new_n1830_;
  assign new_n1832_ = ~pv1213_3_ & ~new_n1769_;
  assign new_n1833_ = pv1213_3_ & new_n1769_;
  assign new_n1834_ = ~new_n1832_ & ~new_n1833_;
  assign new_n1835_ = ~pv1213_1_ & ~new_n1782_;
  assign new_n1836_ = pv1213_1_ & new_n1782_;
  assign new_n1837_ = ~new_n1835_ & ~new_n1836_;
  assign new_n1838_ = new_n1828_ & new_n1831_;
  assign new_n1839_ = new_n1834_ & new_n1838_;
  assign new_n1840_ = new_n1837_ & new_n1839_;
  assign new_n1841_ = ~new_n842_ & new_n1840_;
  assign new_n1842_ = pv288_0_ & new_n1841_;
  assign new_n1843_ = ~new_n1825_ & ~new_n1842_;
  assign new_n1844_ = new_n616_ & new_n1843_;
  assign new_n1845_ = ~new_n1005_ & ~new_n1031_;
  assign new_n1846_ = new_n616_ & new_n1845_;
  assign new_n1847_ = new_n1844_ & new_n1846_;
  assign new_n1848_ = new_n965_ & ~new_n1847_;
  assign new_n1849_ = new_n860_ & ~new_n907_;
  assign new_n1850_ = new_n862_ & ~new_n922_;
  assign new_n1851_ = ~new_n862_ & ~new_n922_;
  assign new_n1852_ = ~new_n1850_ & ~new_n1851_;
  assign new_n1853_ = new_n862_ & ~new_n916_;
  assign new_n1854_ = new_n922_ & ~new_n1067_;
  assign new_n1855_ = ~new_n922_ & new_n1067_;
  assign new_n1856_ = ~new_n1854_ & ~new_n1855_;
  assign new_n1857_ = ~new_n862_ & ~new_n1856_;
  assign new_n1858_ = ~new_n1853_ & ~new_n1857_;
  assign new_n1859_ = new_n1852_ & new_n1858_;
  assign new_n1860_ = new_n862_ & ~new_n931_;
  assign new_n1861_ = ~new_n1075_ & ~new_n1855_;
  assign new_n1862_ = new_n1075_ & new_n1855_;
  assign new_n1863_ = ~new_n1861_ & ~new_n1862_;
  assign new_n1864_ = ~new_n862_ & ~new_n1863_;
  assign new_n1865_ = ~new_n1860_ & ~new_n1864_;
  assign new_n1866_ = new_n1859_ & new_n1865_;
  assign new_n1867_ = new_n862_ & ~new_n907_;
  assign new_n1868_ = ~new_n1062_ & ~new_n1862_;
  assign new_n1869_ = new_n1062_ & new_n1862_;
  assign new_n1870_ = ~new_n1868_ & ~new_n1869_;
  assign new_n1871_ = ~new_n862_ & ~new_n1870_;
  assign new_n1872_ = ~new_n1867_ & ~new_n1871_;
  assign new_n1873_ = ~new_n1866_ & ~new_n1872_;
  assign new_n1874_ = new_n1866_ & new_n1872_;
  assign new_n1875_ = ~new_n1873_ & ~new_n1874_;
  assign new_n1876_ = ~new_n860_ & ~new_n1875_;
  assign new_n1877_ = ~new_n1849_ & ~new_n1876_;
  assign new_n1878_ = ~pv1213_0_ & ~new_n1877_;
  assign new_n1879_ = pv1213_0_ & new_n1877_;
  assign new_n1880_ = ~new_n1878_ & ~new_n1879_;
  assign new_n1881_ = new_n860_ & ~new_n916_;
  assign new_n1882_ = ~new_n1852_ & ~new_n1858_;
  assign new_n1883_ = ~new_n1859_ & ~new_n1882_;
  assign new_n1884_ = ~new_n860_ & ~new_n1883_;
  assign new_n1885_ = ~new_n1881_ & ~new_n1884_;
  assign new_n1886_ = ~pv1213_2_ & ~new_n1885_;
  assign new_n1887_ = pv1213_2_ & new_n1885_;
  assign new_n1888_ = ~new_n1886_ & ~new_n1887_;
  assign new_n1889_ = new_n860_ & ~new_n922_;
  assign new_n1890_ = ~new_n860_ & new_n1852_;
  assign new_n1891_ = ~new_n1889_ & ~new_n1890_;
  assign new_n1892_ = ~pv1213_3_ & ~new_n1891_;
  assign new_n1893_ = pv1213_3_ & new_n1891_;
  assign new_n1894_ = ~new_n1892_ & ~new_n1893_;
  assign new_n1895_ = new_n860_ & ~new_n931_;
  assign new_n1896_ = ~new_n1859_ & ~new_n1865_;
  assign new_n1897_ = ~new_n1866_ & ~new_n1896_;
  assign new_n1898_ = ~new_n860_ & ~new_n1897_;
  assign new_n1899_ = ~new_n1895_ & ~new_n1898_;
  assign new_n1900_ = ~pv1213_1_ & ~new_n1899_;
  assign new_n1901_ = pv1213_1_ & new_n1899_;
  assign new_n1902_ = ~new_n1900_ & ~new_n1901_;
  assign new_n1903_ = ~pv288_2_ & ~pv288_3_;
  assign new_n1904_ = new_n1880_ & new_n1888_;
  assign new_n1905_ = new_n1894_ & new_n1904_;
  assign new_n1906_ = new_n1902_ & new_n1905_;
  assign new_n1907_ = ~new_n842_ & new_n1906_;
  assign new_n1908_ = ~new_n1903_ & new_n1907_;
  assign new_n1909_ = ~pv1213_0_ & ~new_n1872_;
  assign new_n1910_ = pv1213_0_ & new_n1872_;
  assign new_n1911_ = ~new_n1909_ & ~new_n1910_;
  assign new_n1912_ = ~pv1213_2_ & ~new_n1858_;
  assign new_n1913_ = pv1213_2_ & new_n1858_;
  assign new_n1914_ = ~new_n1912_ & ~new_n1913_;
  assign new_n1915_ = ~pv1213_3_ & ~new_n1852_;
  assign new_n1916_ = pv1213_3_ & new_n1852_;
  assign new_n1917_ = ~new_n1915_ & ~new_n1916_;
  assign new_n1918_ = ~pv1213_1_ & ~new_n1865_;
  assign new_n1919_ = pv1213_1_ & new_n1865_;
  assign new_n1920_ = ~new_n1918_ & ~new_n1919_;
  assign new_n1921_ = new_n1911_ & new_n1914_;
  assign new_n1922_ = new_n1917_ & new_n1921_;
  assign new_n1923_ = new_n1920_ & new_n1922_;
  assign new_n1924_ = ~new_n842_ & new_n1923_;
  assign new_n1925_ = pv288_2_ & new_n1924_;
  assign new_n1926_ = ~new_n1908_ & ~new_n1925_;
  assign new_n1927_ = new_n616_ & new_n1926_;
  assign new_n1928_ = ~new_n939_ & ~new_n1083_;
  assign new_n1929_ = new_n616_ & new_n1928_;
  assign new_n1930_ = new_n1927_ & new_n1929_;
  assign new_n1931_ = new_n878_ & ~new_n1930_;
  assign new_n1932_ = new_n856_ & ~new_n904_;
  assign new_n1933_ = ~new_n859_ & new_n867_;
  assign new_n1934_ = ~new_n859_ & ~new_n867_;
  assign new_n1935_ = ~new_n1933_ & ~new_n1934_;
  assign new_n1936_ = new_n867_ & ~new_n873_;
  assign new_n1937_ = new_n859_ & ~new_n1041_;
  assign new_n1938_ = ~new_n859_ & new_n1041_;
  assign new_n1939_ = ~new_n1937_ & ~new_n1938_;
  assign new_n1940_ = ~new_n867_ & ~new_n1939_;
  assign new_n1941_ = ~new_n1936_ & ~new_n1940_;
  assign new_n1942_ = new_n1935_ & new_n1941_;
  assign new_n1943_ = new_n867_ & ~new_n892_;
  assign new_n1944_ = ~new_n1049_ & ~new_n1938_;
  assign new_n1945_ = new_n1049_ & new_n1938_;
  assign new_n1946_ = ~new_n1944_ & ~new_n1945_;
  assign new_n1947_ = ~new_n867_ & ~new_n1946_;
  assign new_n1948_ = ~new_n1943_ & ~new_n1947_;
  assign new_n1949_ = new_n1942_ & new_n1948_;
  assign new_n1950_ = new_n867_ & ~new_n904_;
  assign new_n1951_ = ~new_n1036_ & ~new_n1945_;
  assign new_n1952_ = new_n1036_ & new_n1945_;
  assign new_n1953_ = ~new_n1951_ & ~new_n1952_;
  assign new_n1954_ = ~new_n867_ & ~new_n1953_;
  assign new_n1955_ = ~new_n1950_ & ~new_n1954_;
  assign new_n1956_ = ~new_n1949_ & ~new_n1955_;
  assign new_n1957_ = new_n1949_ & new_n1955_;
  assign new_n1958_ = ~new_n1956_ & ~new_n1957_;
  assign new_n1959_ = ~new_n856_ & ~new_n1958_;
  assign new_n1960_ = ~new_n1932_ & ~new_n1959_;
  assign new_n1961_ = ~pv1213_0_ & ~new_n1960_;
  assign new_n1962_ = pv1213_0_ & new_n1960_;
  assign new_n1963_ = ~new_n1961_ & ~new_n1962_;
  assign new_n1964_ = new_n856_ & ~new_n873_;
  assign new_n1965_ = ~new_n1935_ & ~new_n1941_;
  assign new_n1966_ = ~new_n1942_ & ~new_n1965_;
  assign new_n1967_ = ~new_n856_ & ~new_n1966_;
  assign new_n1968_ = ~new_n1964_ & ~new_n1967_;
  assign new_n1969_ = ~pv1213_2_ & ~new_n1968_;
  assign new_n1970_ = pv1213_2_ & new_n1968_;
  assign new_n1971_ = ~new_n1969_ & ~new_n1970_;
  assign new_n1972_ = new_n856_ & ~new_n859_;
  assign new_n1973_ = ~new_n856_ & new_n1935_;
  assign new_n1974_ = ~new_n1972_ & ~new_n1973_;
  assign new_n1975_ = ~pv1213_3_ & ~new_n1974_;
  assign new_n1976_ = pv1213_3_ & new_n1974_;
  assign new_n1977_ = ~new_n1975_ & ~new_n1976_;
  assign new_n1978_ = new_n856_ & ~new_n892_;
  assign new_n1979_ = ~new_n1942_ & ~new_n1948_;
  assign new_n1980_ = ~new_n1949_ & ~new_n1979_;
  assign new_n1981_ = ~new_n856_ & ~new_n1980_;
  assign new_n1982_ = ~new_n1978_ & ~new_n1981_;
  assign new_n1983_ = ~pv1213_1_ & ~new_n1982_;
  assign new_n1984_ = pv1213_1_ & new_n1982_;
  assign new_n1985_ = ~new_n1983_ & ~new_n1984_;
  assign new_n1986_ = ~pv288_4_ & ~pv288_5_;
  assign new_n1987_ = new_n1963_ & new_n1971_;
  assign new_n1988_ = new_n1977_ & new_n1987_;
  assign new_n1989_ = new_n1985_ & new_n1988_;
  assign new_n1990_ = ~new_n842_ & new_n1989_;
  assign new_n1991_ = ~new_n1986_ & new_n1990_;
  assign new_n1992_ = ~pv1213_0_ & ~new_n1955_;
  assign new_n1993_ = pv1213_0_ & new_n1955_;
  assign new_n1994_ = ~new_n1992_ & ~new_n1993_;
  assign new_n1995_ = ~pv1213_2_ & ~new_n1941_;
  assign new_n1996_ = pv1213_2_ & new_n1941_;
  assign new_n1997_ = ~new_n1995_ & ~new_n1996_;
  assign new_n1998_ = ~pv1213_3_ & ~new_n1935_;
  assign new_n1999_ = pv1213_3_ & new_n1935_;
  assign new_n2000_ = ~new_n1998_ & ~new_n1999_;
  assign new_n2001_ = ~pv1213_1_ & ~new_n1948_;
  assign new_n2002_ = pv1213_1_ & new_n1948_;
  assign new_n2003_ = ~new_n2001_ & ~new_n2002_;
  assign new_n2004_ = new_n1994_ & new_n1997_;
  assign new_n2005_ = new_n2000_ & new_n2004_;
  assign new_n2006_ = new_n2003_ & new_n2005_;
  assign new_n2007_ = ~new_n842_ & new_n2006_;
  assign new_n2008_ = pv288_4_ & new_n2007_;
  assign new_n2009_ = ~new_n1991_ & ~new_n2008_;
  assign new_n2010_ = new_n616_ & new_n2009_;
  assign new_n2011_ = ~new_n956_ & ~new_n1057_;
  assign new_n2012_ = new_n616_ & new_n2011_;
  assign new_n2013_ = new_n2010_ & new_n2012_;
  assign new_n2014_ = new_n881_ & ~new_n2013_;
  assign new_n2015_ = ~new_n1765_ & ~new_n1848_;
  assign new_n2016_ = ~new_n1931_ & ~new_n2014_;
  assign new_n2017_ = new_n2015_ & new_n2016_;
  assign new_n2018_ = ~pv172_0_ & pv240_0_;
  assign pv1719 = ~new_n699_ & new_n2018_;
  assign new_n2020_ = pv1243_7_ & pv1243_9_;
  assign new_n2021_ = ~new_n2017_ & new_n2020_;
  assign new_n2022_ = pv1243_8_ & new_n2021_;
  assign new_n2023_ = ~pv248_0_ & new_n2022_;
  assign new_n2024_ = pv1719 & new_n2023_;
  assign new_n2025_ = pv243_0_ & pv244_0_;
  assign new_n2026_ = pv245_0_ & new_n2025_;
  assign new_n2027_ = pv246_0_ & new_n2026_;
  assign new_n2028_ = pv247_0_ & new_n2027_;
  assign new_n2029_ = pv1719 & new_n2028_;
  assign new_n2030_ = ~pv248_0_ & new_n2029_;
  assign new_n2031_ = new_n1380_ & pv1719;
  assign new_n2032_ = ~pv248_0_ & new_n2031_;
  assign new_n2033_ = ~new_n2024_ & ~new_n2030_;
  assign pv393_0_ = new_n2032_ | ~new_n2033_;
  assign pv500_0_ = pv271_0_ | ~pv14_0_;
  assign pv544 = new_n491_ & pv1213_7_;
  assign new_n2037_ = pv257_2_ & pv257_1_;
  assign new_n2038_ = pv257_5_ & new_n2037_;
  assign new_n2039_ = pv257_3_ & new_n2038_;
  assign new_n2040_ = pv257_7_ & new_n2039_;
  assign new_n2041_ = pv257_4_ & new_n2040_;
  assign new_n2042_ = pv257_6_ & new_n2041_;
  assign new_n2043_ = pv257_0_ & ~new_n2042_;
  assign new_n2044_ = ~pv257_0_ & new_n2042_;
  assign pv650 = new_n2043_ | new_n2044_;
  assign new_n2046_ = pv213_3_ & new_n1704_;
  assign new_n2047_ = ~new_n1589_ & new_n2046_;
  assign new_n2048_ = pv165_5_ & new_n1586_;
  assign pv1297_2_ = new_n2047_ | new_n2048_;
  assign new_n2050_ = ~pv88_3_ & new_n572_;
  assign new_n2051_ = ~pv134_1_ & ~new_n572_;
  assign pv1771_1_ = new_n2050_ | new_n2051_;
  assign new_n2053_ = pv100_0_ & new_n1721_;
  assign new_n2054_ = pv124_0_ & new_n1725_;
  assign new_n2055_ = pv213_0_ & new_n1728_;
  assign new_n2056_ = pv108_0_ & new_n1732_;
  assign new_n2057_ = ~new_n2053_ & ~new_n2054_;
  assign new_n2058_ = ~new_n2055_ & ~new_n2056_;
  assign pv1921_0_ = ~new_n2057_ | ~new_n2058_;
  assign new_n2060_ = pv802_0_ & ~new_n639_;
  assign new_n2061_ = ~new_n1388_ & ~new_n2060_;
  assign new_n2062_ = pv134_1_ & ~pv134_0_;
  assign new_n2063_ = ~pv134_1_ & pv134_0_;
  assign new_n2064_ = ~new_n2062_ & ~new_n2063_;
  assign new_n2065_ = ~new_n2060_ & ~new_n2061_;
  assign new_n2066_ = new_n1388_ & new_n2065_;
  assign new_n2067_ = ~new_n2064_ & new_n2066_;
  assign new_n2068_ = new_n1388_ & ~new_n2060_;
  assign new_n2069_ = ~new_n1388_ & ~new_n2068_;
  assign new_n2070_ = ~new_n2060_ & new_n2069_;
  assign new_n2071_ = pv134_0_ & new_n2070_;
  assign pv1992_0_ = new_n2067_ | new_n2071_;
  assign pv541 = new_n491_ & pv1213_4_;
  assign new_n2074_ = ~pv214_0_ & ~new_n699_;
  assign new_n2075_ = new_n1285_ & new_n2074_;
  assign new_n2076_ = ~new_n704_ & new_n2075_;
  assign new_n2077_ = ~new_n557_ & ~new_n1279_;
  assign new_n2078_ = pv59_0_ & ~new_n699_;
  assign new_n2079_ = ~new_n2077_ & new_n2078_;
  assign new_n2080_ = ~pv214_0_ & new_n2079_;
  assign new_n2081_ = pv62_0_ & ~new_n699_;
  assign new_n2082_ = new_n1132_ & new_n2081_;
  assign new_n2083_ = ~pv214_0_ & new_n2082_;
  assign new_n2084_ = ~new_n2076_ & ~new_n2080_;
  assign pv620 = ~new_n2083_ & new_n2084_;
  assign new_n2086_ = pv62_0_ & new_n758_;
  assign new_n2087_ = new_n557_ & new_n2086_;
  assign new_n2088_ = pv14_0_ & new_n2087_;
  assign new_n2089_ = ~new_n491_ & ~new_n1280_;
  assign new_n2090_ = ~new_n573_ & ~new_n773_;
  assign new_n2091_ = new_n2089_ & new_n2090_;
  assign new_n2092_ = ~new_n494_ & ~new_n575_;
  assign new_n2093_ = ~new_n766_ & new_n2092_;
  assign new_n2094_ = new_n2091_ & new_n2093_;
  assign new_n2095_ = ~pv174_0_ & new_n585_;
  assign new_n2096_ = new_n2094_ & ~new_n2095_;
  assign new_n2097_ = pv59_0_ & new_n2096_;
  assign new_n2098_ = ~new_n713_ & new_n2097_;
  assign new_n2099_ = ~pv1719 & new_n2098_;
  assign new_n2100_ = pv14_0_ & new_n2099_;
  assign new_n2101_ = ~new_n841_ & new_n2100_;
  assign new_n2102_ = new_n758_ & new_n2101_;
  assign pv1274_0_ = new_n2088_ | new_n2102_;
  assign new_n2104_ = pv213_4_ & new_n1704_;
  assign new_n2105_ = ~new_n1589_ & new_n2104_;
  assign new_n2106_ = pv165_6_ & new_n1586_;
  assign pv1297_3_ = new_n2105_ | new_n2106_;
  assign pv1432 = pv66_0_ & new_n1628_;
  assign new_n2109_ = pv242_0_ & new_n639_;
  assign new_n2110_ = pv14_0_ & new_n2109_;
  assign new_n2111_ = ~pv1536_0_ & new_n1381_;
  assign new_n2112_ = ~new_n640_ & new_n2111_;
  assign pv1726_0_ = new_n2110_ | new_n2112_;
  assign new_n2114_ = pv100_3_ & new_n1721_;
  assign new_n2115_ = pv124_3_ & new_n1725_;
  assign new_n2116_ = pv213_3_ & new_n1728_;
  assign new_n2117_ = pv108_3_ & new_n1732_;
  assign new_n2118_ = ~new_n2114_ & ~new_n2115_;
  assign new_n2119_ = ~new_n2116_ & ~new_n2117_;
  assign pv1921_3_ = ~new_n2118_ | ~new_n2119_;
  assign new_n2121_ = pv101_0_ & new_n1152_;
  assign new_n2122_ = ~pv108_4_ & new_n2121_;
  assign new_n2123_ = pv56_0_ & new_n1096_;
  assign new_n2124_ = pv14_0_ & ~new_n2122_;
  assign new_n2125_ = ~new_n2123_ & new_n2124_;
  assign new_n2126_ = pv110_0_ & new_n2125_;
  assign new_n2127_ = ~pv102_0_ & ~pv1758_0_;
  assign new_n2128_ = new_n510_ & ~new_n2127_;
  assign new_n2129_ = ~pv110_0_ & new_n2128_;
  assign pv1968_0_ = new_n2126_ | new_n2129_;
  assign new_n2131_ = ~pv134_1_ & new_n2066_;
  assign new_n2132_ = pv134_1_ & new_n2070_;
  assign pv1992_1_ = new_n2131_ | new_n2132_;
  assign new_n2134_ = ~new_n1759_ & ~new_n2008_;
  assign new_n2135_ = ~new_n1842_ & new_n2134_;
  assign new_n2136_ = ~new_n1925_ & new_n2135_;
  assign new_n2137_ = new_n616_ & new_n2136_;
  assign new_n2138_ = ~new_n939_ & new_n2137_;
  assign new_n2139_ = ~new_n1005_ & new_n2138_;
  assign new_n2140_ = ~new_n848_ & new_n2139_;
  assign pv357 = ~new_n956_ & new_n2140_;
  assign new_n2142_ = new_n505_ & new_n616_;
  assign new_n2143_ = new_n545_ & new_n2142_;
  assign new_n2144_ = new_n549_ & new_n2143_;
  assign new_n2145_ = pv802_0_ & ~new_n2144_;
  assign new_n2146_ = ~new_n557_ & new_n774_;
  assign new_n2147_ = ~pv174_0_ & ~new_n555_;
  assign new_n2148_ = new_n2146_ & new_n2147_;
  assign new_n2149_ = pv56_0_ & ~new_n2148_;
  assign new_n2150_ = new_n616_ & new_n1215_;
  assign new_n2151_ = pv59_0_ & ~new_n2150_;
  assign new_n2152_ = pv70_0_ & ~new_n616_;
  assign new_n2153_ = pv802_0_ & new_n1502_;
  assign new_n2154_ = ~pv215_0_ & pv66_0_;
  assign new_n2155_ = pv763 & new_n2154_;
  assign new_n2156_ = ~new_n699_ & new_n2155_;
  assign new_n2157_ = ~new_n2145_ & ~new_n2149_;
  assign new_n2158_ = ~new_n1212_ & ~new_n2151_;
  assign new_n2159_ = new_n2157_ & new_n2158_;
  assign new_n2160_ = ~new_n2152_ & ~new_n2153_;
  assign new_n2161_ = ~pv1719 & ~new_n2156_;
  assign new_n2162_ = new_n2160_ & new_n2161_;
  assign pv423_0_ = ~new_n2159_ | ~new_n2162_;
  assign pv542 = new_n491_ & pv1213_5_;
  assign new_n2165_ = pv41_0_ & ~pv45_0_;
  assign new_n2166_ = ~pv41_0_ & pv45_0_;
  assign new_n2167_ = ~new_n2165_ & ~new_n2166_;
  assign pv621 = pv293_0_ & new_n2167_;
  assign new_n2169_ = pv62_0_ & new_n572_;
  assign new_n2170_ = pv56_0_ & new_n572_;
  assign new_n2171_ = ~new_n491_ & ~new_n573_;
  assign new_n2172_ = ~new_n575_ & new_n2171_;
  assign new_n2173_ = pv802_0_ & ~new_n2172_;
  assign new_n2174_ = new_n507_ & new_n2173_;
  assign new_n2175_ = new_n507_ & ~new_n732_;
  assign new_n2176_ = pv59_0_ & new_n2175_;
  assign new_n2177_ = ~new_n2170_ & ~new_n2174_;
  assign new_n2178_ = ~pv270_0_ & ~new_n2176_;
  assign new_n2179_ = new_n2177_ & new_n2178_;
  assign new_n2180_ = ~pv302_0_ & ~new_n2169_;
  assign pv630 = ~new_n2179_ & new_n2180_;
  assign new_n2182_ = pv213_5_ & new_n1704_;
  assign new_n2183_ = ~new_n1589_ & new_n2182_;
  assign new_n2184_ = pv165_7_ & new_n1586_;
  assign pv1297_4_ = new_n2183_ | new_n2184_;
  assign new_n2186_ = pv100_2_ & new_n1721_;
  assign new_n2187_ = pv124_2_ & new_n1725_;
  assign new_n2188_ = pv213_2_ & new_n1728_;
  assign new_n2189_ = pv108_2_ & new_n1732_;
  assign new_n2190_ = ~new_n2186_ & ~new_n2187_;
  assign new_n2191_ = ~new_n2188_ & ~new_n2189_;
  assign pv1921_2_ = ~new_n2190_ | ~new_n2191_;
  assign pv547 = new_n491_ & pv1213_10_;
  assign new_n2194_ = pv257_6_ & pv257_7_;
  assign new_n2195_ = pv257_5_ & ~new_n2194_;
  assign new_n2196_ = ~pv257_5_ & new_n2194_;
  assign pv655 = new_n2195_ | new_n2196_;
  assign new_n2198_ = ~pv259_0_ & new_n1661_;
  assign new_n2199_ = pv259_0_ & new_n1663_;
  assign new_n2200_ = ~new_n2198_ & ~new_n2199_;
  assign new_n2201_ = pv14_0_ & new_n2200_;
  assign new_n2202_ = pv260_0_ & new_n2201_;
  assign new_n2203_ = pv14_0_ & ~new_n2200_;
  assign new_n2204_ = ~pv260_0_ & new_n2203_;
  assign pv1467_0_ = new_n2202_ | new_n2204_;
  assign new_n2206_ = pv62_0_ & pv91_1_;
  assign new_n2207_ = pv59_0_ & pv91_0_;
  assign new_n2208_ = ~new_n2206_ & ~new_n2207_;
  assign new_n2209_ = new_n1223_ & ~new_n2208_;
  assign new_n2210_ = ~pv294_0_ & ~new_n1279_;
  assign new_n2211_ = ~new_n1132_ & new_n2210_;
  assign new_n2212_ = new_n2167_ & ~new_n2209_;
  assign pv1629_0_ = new_n2211_ | ~new_n2212_;
  assign new_n2214_ = pv108_0_ & ~new_n1714_;
  assign new_n2215_ = ~new_n1278_ & ~new_n2214_;
  assign pv1896_0_ = new_n1153_ | ~new_n2215_;
  assign new_n2217_ = pv213_5_ & new_n1728_;
  assign new_n2218_ = pv100_5_ & new_n1721_;
  assign new_n2219_ = pv124_5_ & new_n1725_;
  assign new_n2220_ = ~new_n2217_ & ~new_n2218_;
  assign pv1921_5_ = new_n2219_ | ~new_n2220_;
  assign new_n2222_ = ~pv35_0_ & ~new_n1496_;
  assign pv377 = pv203_0_ & ~new_n2222_;
  assign pv548 = new_n491_ & pv1213_11_;
  assign new_n2225_ = pv257_6_ & pv257_5_;
  assign new_n2226_ = pv257_7_ & new_n2225_;
  assign new_n2227_ = pv257_4_ & ~new_n2226_;
  assign new_n2228_ = ~pv257_4_ & new_n2226_;
  assign pv654 = new_n2227_ | new_n2228_;
  assign new_n2230_ = new_n494_ & pv802_0_;
  assign new_n2231_ = ~pv279_0_ & ~new_n2230_;
  assign new_n2232_ = pv149_5_ & new_n2230_;
  assign pv821_0_ = new_n2231_ | new_n2232_;
  assign new_n2234_ = new_n491_ & new_n1278_;
  assign new_n2235_ = pv108_1_ & ~new_n1714_;
  assign pv1897_0_ = new_n2234_ | new_n2235_;
  assign new_n2237_ = pv100_4_ & new_n1721_;
  assign new_n2238_ = pv124_4_ & new_n1725_;
  assign new_n2239_ = pv213_4_ & new_n1728_;
  assign new_n2240_ = pv108_4_ & new_n1732_;
  assign new_n2241_ = ~new_n2237_ & ~new_n2238_;
  assign new_n2242_ = ~new_n2239_ & ~new_n2240_;
  assign pv1921_4_ = ~new_n2241_ | ~new_n2242_;
  assign new_n2244_ = pv56_0_ & new_n773_;
  assign new_n2245_ = pv59_0_ & ~new_n545_;
  assign new_n2246_ = ~new_n554_ & new_n2245_;
  assign new_n2247_ = pv56_0_ & new_n766_;
  assign new_n2248_ = pv59_0_ & ~new_n505_;
  assign new_n2249_ = ~new_n786_ & ~new_n2244_;
  assign new_n2250_ = ~new_n2246_ & new_n2249_;
  assign new_n2251_ = ~new_n2247_ & new_n2250_;
  assign new_n2252_ = ~new_n1212_ & new_n2251_;
  assign new_n2253_ = ~new_n2248_ & new_n2252_;
  assign new_n2254_ = ~pv43_0_ & ~new_n699_;
  assign new_n2255_ = ~pv214_0_ & new_n2254_;
  assign new_n2256_ = ~new_n2253_ & new_n2255_;
  assign pv527 = ~new_n704_ & new_n2256_;
  assign pv538 = new_n491_ & pv1213_1_;
  assign pv545 = new_n491_ & pv1213_8_;
  assign new_n2260_ = pv257_4_ & new_n2225_;
  assign new_n2261_ = pv257_7_ & new_n2260_;
  assign new_n2262_ = pv257_3_ & ~new_n2261_;
  assign new_n2263_ = ~pv257_3_ & new_n2261_;
  assign pv653 = new_n2262_ | new_n2263_;
  assign new_n2265_ = pv37_0_ & ~pv1213_2_;
  assign new_n2266_ = ~pv37_0_ & pv321_2_;
  assign pv1829_0_ = new_n2265_ | new_n2266_;
  assign new_n2268_ = new_n490_ & new_n719_;
  assign new_n2269_ = pv108_2_ & ~new_n1714_;
  assign pv1898_0_ = new_n2268_ | new_n2269_;
  assign pv537 = new_n491_ & pv1213_0_;
  assign pv546 = new_n491_ & pv1213_9_;
  assign new_n2273_ = ~new_n1689_ & ~new_n2025_;
  assign new_n2274_ = pv245_0_ & new_n2273_;
  assign new_n2275_ = ~new_n1689_ & new_n2025_;
  assign new_n2276_ = ~pv245_0_ & new_n2275_;
  assign pv597_0_ = new_n2274_ | new_n2276_;
  assign new_n2278_ = pv257_4_ & pv257_6_;
  assign new_n2279_ = pv257_5_ & new_n2278_;
  assign new_n2280_ = pv257_3_ & new_n2279_;
  assign new_n2281_ = pv257_7_ & new_n2280_;
  assign new_n2282_ = pv257_2_ & ~new_n2281_;
  assign new_n2283_ = ~pv257_2_ & new_n2281_;
  assign pv652 = new_n2282_ | new_n2283_;
  assign pv801 = new_n579_ & new_n586_;
  assign new_n2286_ = new_n510_ & new_n719_;
  assign new_n2287_ = pv108_3_ & ~new_n1714_;
  assign pv1899_0_ = new_n2286_ | new_n2287_;
  assign new_n2289_ = ~pv802_0_ & new_n1502_;
  assign new_n2290_ = ~new_n1392_ & ~new_n2289_;
  assign new_n2291_ = new_n575_ & pv802_0_;
  assign new_n2292_ = new_n2290_ & ~new_n2291_;
  assign new_n2293_ = pv802_0_ & new_n2292_;
  assign new_n2294_ = new_n491_ & new_n2293_;
  assign new_n2295_ = pv1243_8_ & new_n2294_;
  assign new_n2296_ = new_n491_ & pv802_0_;
  assign new_n2297_ = ~pv199_4_ & pv199_3_;
  assign new_n2298_ = pv199_4_ & ~pv199_3_;
  assign new_n2299_ = ~new_n2297_ & ~new_n2298_;
  assign new_n2300_ = ~new_n2291_ & ~new_n2296_;
  assign new_n2301_ = ~new_n2290_ & new_n2300_;
  assign new_n2302_ = ~new_n2299_ & new_n2301_;
  assign pv572_8_ = new_n2295_ | new_n2302_;
  assign new_n2304_ = ~new_n510_ & ~new_n567_;
  assign new_n2305_ = pv290_0_ & ~new_n2304_;
  assign new_n2306_ = new_n699_ & new_n2305_;
  assign new_n2307_ = pv56_0_ & new_n1718_;
  assign new_n2308_ = pv14_0_ & ~new_n2306_;
  assign new_n2309_ = pv100_2_ & new_n2308_;
  assign new_n2310_ = ~new_n2307_ & new_n2309_;
  assign new_n2311_ = pv165_4_ & new_n2306_;
  assign pv1709_1_ = new_n2310_ | new_n2311_;
  assign pv373 = pv10_0_ & pv13_0_;
  assign new_n2314_ = pv1243_7_ & new_n2294_;
  assign new_n2315_ = pv199_4_ & pv199_3_;
  assign new_n2316_ = pv199_2_ & ~new_n2315_;
  assign new_n2317_ = ~pv199_2_ & new_n2315_;
  assign new_n2318_ = ~new_n2316_ & ~new_n2317_;
  assign new_n2319_ = new_n2301_ & ~new_n2318_;
  assign pv572_7_ = new_n2314_ | new_n2319_;
  assign new_n2321_ = ~pv149_6_ & new_n582_;
  assign new_n2322_ = pv14_0_ & ~new_n491_;
  assign new_n2323_ = pv277_0_ & new_n2322_;
  assign pv1439_0_ = new_n2321_ | new_n2323_;
  assign new_n2325_ = pv100_1_ & new_n2308_;
  assign new_n2326_ = ~new_n2307_ & new_n2325_;
  assign new_n2327_ = pv165_3_ & new_n2306_;
  assign pv1709_0_ = new_n2326_ | new_n2327_;
  assign new_n2329_ = pv1243_6_ & new_n2294_;
  assign new_n2330_ = pv199_3_ & pv199_2_;
  assign new_n2331_ = pv199_4_ & new_n2330_;
  assign new_n2332_ = pv199_1_ & ~new_n2331_;
  assign new_n2333_ = ~pv199_1_ & new_n2331_;
  assign new_n2334_ = ~new_n2332_ & ~new_n2333_;
  assign new_n2335_ = new_n2301_ & ~new_n2334_;
  assign pv572_6_ = new_n2329_ | new_n2335_;
  assign new_n2337_ = ~pv69_0_ & ~pv50_0_;
  assign pv1539 = new_n1628_ & ~new_n2337_;
  assign new_n2339_ = pv1243_5_ & new_n2294_;
  assign new_n2340_ = pv199_1_ & new_n2330_;
  assign new_n2341_ = pv199_4_ & new_n2340_;
  assign new_n2342_ = pv199_0_ & ~new_n2341_;
  assign new_n2343_ = ~pv199_0_ & new_n2341_;
  assign new_n2344_ = ~new_n2342_ & ~new_n2343_;
  assign new_n2345_ = new_n2301_ & ~new_n2344_;
  assign pv572_5_ = new_n2339_ | new_n2345_;
  assign new_n2347_ = pv165_3_ & ~pv165_5_;
  assign new_n2348_ = new_n758_ & new_n2347_;
  assign new_n2349_ = pv763 & new_n2348_;
  assign new_n2350_ = pv14_0_ & new_n2349_;
  assign new_n2351_ = pv70_0_ & new_n2350_;
  assign new_n2352_ = ~pv165_4_ & new_n2351_;
  assign new_n2353_ = pv165_6_ & new_n2352_;
  assign new_n2354_ = pv65_0_ & ~new_n555_;
  assign new_n2355_ = new_n758_ & new_n2354_;
  assign new_n2356_ = ~new_n1132_ & new_n2355_;
  assign new_n2357_ = pv14_0_ & new_n2356_;
  assign pv1392_0_ = new_n2353_ | new_n2357_;
  assign new_n2359_ = pv258_0_ & ~pv259_0_;
  assign new_n2360_ = ~pv260_0_ & new_n2359_;
  assign new_n2361_ = ~pv59_0_ & new_n2360_;
  assign new_n2362_ = pv262_0_ & ~new_n2361_;
  assign new_n2363_ = pv14_0_ & new_n2362_;
  assign pv1679_0_ = ~new_n615_ | new_n2363_;
  assign new_n2365_ = new_n616_ & ~new_n842_;
  assign new_n2366_ = ~new_n1755_ & ~new_n1991_;
  assign new_n2367_ = ~new_n1825_ & new_n2366_;
  assign new_n2368_ = ~new_n1908_ & new_n2367_;
  assign new_n2369_ = new_n2365_ & new_n2368_;
  assign new_n2370_ = ~new_n1083_ & new_n2369_;
  assign new_n2371_ = ~new_n1031_ & new_n2370_;
  assign new_n2372_ = ~new_n854_ & new_n2371_;
  assign pv356 = ~new_n1057_ & new_n2372_;
  assign new_n2374_ = pv215_0_ & pv66_0_;
  assign new_n2375_ = pv66_0_ & new_n762_;
  assign new_n2376_ = pv66_0_ & pv763;
  assign new_n2377_ = new_n493_ & pv802_0_;
  assign new_n2378_ = ~new_n491_ & ~new_n511_;
  assign new_n2379_ = ~pv763 & ~new_n2378_;
  assign new_n2380_ = pv802_0_ & new_n2379_;
  assign new_n2381_ = ~new_n713_ & ~new_n1132_;
  assign new_n2382_ = ~new_n1133_ & ~new_n1223_;
  assign new_n2383_ = new_n2381_ & new_n2382_;
  assign new_n2384_ = pv56_0_ & ~new_n2383_;
  assign new_n2385_ = ~new_n2375_ & ~new_n2376_;
  assign new_n2386_ = ~new_n2377_ & new_n2385_;
  assign new_n2387_ = ~new_n2380_ & ~new_n2384_;
  assign new_n2388_ = new_n2386_ & new_n2387_;
  assign new_n2389_ = ~pv32_1_ & ~new_n997_;
  assign new_n2390_ = pv32_1_ & new_n997_;
  assign new_n2391_ = ~new_n2389_ & ~new_n2390_;
  assign new_n2392_ = ~pv32_0_ & ~new_n973_;
  assign new_n2393_ = pv32_0_ & new_n973_;
  assign new_n2394_ = ~new_n2392_ & ~new_n2393_;
  assign new_n2395_ = ~pv32_2_ & ~new_n982_;
  assign new_n2396_ = pv32_2_ & new_n982_;
  assign new_n2397_ = ~new_n2395_ & ~new_n2396_;
  assign new_n2398_ = new_n988_ & new_n2391_;
  assign new_n2399_ = new_n2394_ & new_n2398_;
  assign new_n2400_ = pv32_3_ & new_n2399_;
  assign new_n2401_ = new_n2397_ & new_n2400_;
  assign new_n2402_ = new_n2390_ & new_n2394_;
  assign new_n2403_ = new_n982_ & new_n2394_;
  assign new_n2404_ = pv32_2_ & new_n2403_;
  assign new_n2405_ = new_n2391_ & new_n2404_;
  assign new_n2406_ = ~new_n2393_ & ~new_n2401_;
  assign new_n2407_ = ~new_n2402_ & ~new_n2405_;
  assign new_n2408_ = new_n2406_ & new_n2407_;
  assign new_n2409_ = ~new_n2388_ & ~new_n2408_;
  assign new_n2410_ = new_n1496_ & pv1719;
  assign new_n2411_ = new_n702_ & pv1719;
  assign new_n2412_ = pv302_0_ & pv1719;
  assign new_n2413_ = ~new_n554_ & ~pv763;
  assign new_n2414_ = pv802_0_ & ~new_n2413_;
  assign new_n2415_ = ~new_n2374_ & ~new_n2409_;
  assign new_n2416_ = ~pv43_0_ & new_n2415_;
  assign new_n2417_ = new_n616_ & new_n2416_;
  assign new_n2418_ = ~pv214_0_ & new_n2417_;
  assign new_n2419_ = ~new_n2032_ & new_n2418_;
  assign new_n2420_ = ~new_n2024_ & new_n2419_;
  assign new_n2421_ = ~new_n2410_ & new_n2420_;
  assign new_n2422_ = ~new_n2030_ & new_n2421_;
  assign new_n2423_ = ~new_n2411_ & new_n2422_;
  assign new_n2424_ = ~new_n2412_ & new_n2423_;
  assign new_n2425_ = pv423_0_ & new_n2424_;
  assign new_n2426_ = ~new_n1278_ & new_n2425_;
  assign new_n2427_ = ~new_n704_ & new_n2426_;
  assign new_n2428_ = ~pv1757_0_ & new_n2427_;
  assign pv432 = ~new_n2414_ & new_n2428_;
  assign pv435_0_ = pv630 | pv432;
  assign new_n2431_ = pv216_0_ & ~pv214_0_;
  assign new_n2432_ = ~pv68_0_ & ~pv69_0_;
  assign new_n2433_ = ~pv66_0_ & new_n2432_;
  assign new_n2434_ = ~pv70_0_ & new_n2433_;
  assign new_n2435_ = pv14_0_ & new_n730_;
  assign new_n2436_ = ~new_n2434_ & new_n2435_;
  assign new_n2437_ = pv215_0_ & new_n2436_;
  assign pv1492_0_ = new_n2431_ | new_n2437_;
  assign pv1537 = pv68_0_ & new_n1628_;
  assign new_n2440_ = ~pv43_0_ & pv45_0_;
  assign pv511_0_ = pv40_0_ | new_n2440_;
  assign pv540 = new_n491_ & pv1213_3_;
  assign new_n2443_ = ~new_n1689_ & ~new_n2027_;
  assign new_n2444_ = pv247_0_ & new_n2443_;
  assign new_n2445_ = ~new_n1689_ & new_n2027_;
  assign new_n2446_ = ~pv247_0_ & new_n2445_;
  assign pv609_0_ = new_n2444_ | new_n2446_;
  assign pv1426 = pv1_0_ & new_n692_;
  assign new_n2449_ = ~pv302_0_ & pv292_0_;
  assign new_n2450_ = pv174_0_ & new_n699_;
  assign new_n2451_ = pv174_0_ & ~new_n755_;
  assign new_n2452_ = ~new_n579_ & ~new_n2449_;
  assign new_n2453_ = ~new_n2450_ & ~new_n2451_;
  assign pv1620_0_ = ~new_n2452_ | ~new_n2453_;
  assign new_n2455_ = ~pv290_0_ & ~pv802_0_;
  assign new_n2456_ = new_n702_ & new_n2455_;
  assign new_n2457_ = new_n732_ & new_n2456_;
  assign pv1736 = ~pv289_0_ & new_n2457_;
  assign pv1429 = pv1_0_ & pv12_0_;
  assign new_n2460_ = ~new_n1490_ & ~new_n2363_;
  assign new_n2461_ = pv262_0_ & new_n2460_;
  assign new_n2462_ = pv261_0_ & ~new_n2461_;
  assign new_n2463_ = ~new_n1662_ & ~new_n2462_;
  assign pv1832 = pv14_0_ & ~new_n2463_;
  assign new_n2465_ = pv1243_9_ & new_n2294_;
  assign new_n2466_ = ~pv199_4_ & new_n2301_;
  assign pv572_9_ = new_n2465_ | new_n2466_;
  assign new_n2468_ = pv213_1_ & new_n1704_;
  assign new_n2469_ = ~new_n1589_ & new_n2468_;
  assign new_n2470_ = pv165_3_ & new_n1586_;
  assign pv1297_0_ = new_n2469_ | new_n2470_;
  assign pv1428 = pv1_0_ & pv11_0_;
  assign new_n2473_ = new_n1583_ & ~new_n2304_;
  assign new_n2474_ = ~new_n2306_ & ~new_n2473_;
  assign new_n2475_ = pv14_0_ & new_n2474_;
  assign new_n2476_ = pv100_0_ & new_n2475_;
  assign new_n2477_ = ~new_n2307_ & new_n2476_;
  assign new_n2478_ = ~new_n1595_ & ~new_n2474_;
  assign pv1693_0_ = new_n2477_ | new_n2478_;
  assign new_n2480_ = pv108_5_ & ~new_n1404_;
  assign pv1901_0_ = new_n1308_ | new_n2480_;
  assign new_n2482_ = pv194_0_ & ~new_n1380_;
  assign new_n2483_ = ~pv194_0_ & new_n1380_;
  assign new_n2484_ = ~new_n2482_ & ~new_n2483_;
  assign new_n2485_ = new_n2301_ & ~new_n2484_;
  assign new_n2486_ = new_n2290_ & ~new_n2296_;
  assign new_n2487_ = pv802_0_ & new_n2486_;
  assign new_n2488_ = new_n575_ & new_n2487_;
  assign new_n2489_ = pv149_4_ & new_n2488_;
  assign new_n2490_ = ~pv321_2_ & new_n2294_;
  assign new_n2491_ = ~new_n2485_ & ~new_n2489_;
  assign pv572_0_ = new_n2490_ | ~new_n2491_;
  assign new_n2493_ = pv239_4_ & ~pv239_3_;
  assign new_n2494_ = ~pv239_4_ & pv239_3_;
  assign new_n2495_ = ~new_n2493_ & ~new_n2494_;
  assign new_n2496_ = ~pv802_0_ & ~new_n694_;
  assign new_n2497_ = new_n494_ & new_n2496_;
  assign new_n2498_ = ~new_n2495_ & new_n2497_;
  assign new_n2499_ = new_n494_ & ~pv802_0_;
  assign new_n2500_ = new_n694_ & ~new_n2499_;
  assign new_n2501_ = pv1243_8_ & new_n2500_;
  assign pv1552_0_ = new_n2498_ | new_n2501_;
  assign new_n2503_ = pv33_0_ & ~new_n490_;
  assign new_n2504_ = pv289_0_ & new_n2503_;
  assign pv1745_0_ = new_n585_ | ~new_n2504_;
  assign new_n2506_ = pv37_0_ & ~pv1243_9_;
  assign pv1829_9_ = new_n2266_ | new_n2506_;
  assign new_n2508_ = pv149_3_ & ~new_n1093_;
  assign new_n2509_ = ~new_n1713_ & new_n2508_;
  assign new_n2510_ = new_n567_ & new_n2509_;
  assign new_n2511_ = ~new_n841_ & new_n2510_;
  assign new_n2512_ = pv149_5_ & new_n567_;
  assign new_n2513_ = ~pv149_3_ & new_n2512_;
  assign new_n2514_ = pv149_4_ & new_n2513_;
  assign new_n2515_ = ~pv149_7_ & new_n2514_;
  assign new_n2516_ = ~pv149_6_ & new_n2515_;
  assign new_n2517_ = ~pv149_6_ & new_n1717_;
  assign new_n2518_ = ~new_n2511_ & ~new_n2516_;
  assign new_n2519_ = ~new_n2517_ & new_n2518_;
  assign new_n2520_ = ~pv302_0_ & ~new_n2519_;
  assign new_n2521_ = pv149_0_ & pv149_1_;
  assign new_n2522_ = ~pv149_2_ & new_n2521_;
  assign new_n2523_ = pv149_0_ & pv149_2_;
  assign new_n2524_ = ~pv149_1_ & new_n2523_;
  assign new_n2525_ = pv149_2_ & new_n2521_;
  assign new_n2526_ = ~new_n2522_ & ~new_n2524_;
  assign new_n2527_ = new_n2519_ & new_n2526_;
  assign new_n2528_ = ~new_n2525_ & new_n2527_;
  assign new_n2529_ = ~new_n2520_ & ~new_n2528_;
  assign new_n2530_ = new_n616_ & new_n2529_;
  assign new_n2531_ = pv65_0_ & new_n1132_;
  assign new_n2532_ = pv258_0_ & ~pv260_0_;
  assign new_n2533_ = ~new_n616_ & new_n2532_;
  assign new_n2534_ = ~pv259_0_ & new_n2533_;
  assign new_n2535_ = ~pv59_0_ & new_n2534_;
  assign new_n2536_ = ~new_n1718_ & ~new_n2535_;
  assign new_n2537_ = ~new_n1224_ & new_n2536_;
  assign new_n2538_ = ~new_n1095_ & new_n2537_;
  assign new_n2539_ = ~new_n2321_ & new_n2538_;
  assign new_n2540_ = ~new_n1096_ & new_n2539_;
  assign new_n2541_ = ~new_n1588_ & new_n2540_;
  assign new_n2542_ = pv56_0_ & ~new_n2541_;
  assign new_n2543_ = pv62_0_ & ~new_n2382_;
  assign new_n2544_ = ~new_n2531_ & ~new_n2542_;
  assign new_n2545_ = ~new_n2543_ & new_n2544_;
  assign new_n2546_ = ~pv1741_0_ & ~new_n2545_;
  assign new_n2547_ = ~new_n702_ & new_n2546_;
  assign new_n2548_ = new_n758_ & ~new_n1496_;
  assign new_n2549_ = ~new_n732_ & ~new_n2548_;
  assign new_n2550_ = pv290_0_ & ~new_n699_;
  assign new_n2551_ = ~pv289_0_ & ~new_n2547_;
  assign new_n2552_ = ~pv214_0_ & ~new_n2549_;
  assign new_n2553_ = new_n2551_ & new_n2552_;
  assign new_n2554_ = ~pv302_0_ & ~new_n701_;
  assign new_n2555_ = ~new_n2550_ & new_n2554_;
  assign new_n2556_ = new_n2553_ & new_n2555_;
  assign new_n2557_ = ~new_n2530_ & new_n2556_;
  assign pv798_0_ = ~pv14_0_ | ~new_n2557_;
  assign new_n2559_ = ~pv239_4_ & new_n2497_;
  assign new_n2560_ = pv1243_9_ & new_n2500_;
  assign pv1552_1_ = new_n2559_ | new_n2560_;
  assign new_n2562_ = pv802_0_ & new_n791_;
  assign new_n2563_ = ~new_n1580_ & ~new_n2562_;
  assign pv1645_0_ = new_n2409_ | ~new_n2563_;
  assign new_n2565_ = new_n507_ & ~new_n2172_;
  assign new_n2566_ = pv295_0_ & ~new_n2565_;
  assign new_n2567_ = new_n616_ & new_n2566_;
  assign new_n2568_ = ~pv249_0_ & new_n2567_;
  assign new_n2569_ = ~pv289_0_ & new_n2568_;
  assign pv1652_0_ = pv290_0_ | ~new_n2569_;
  assign new_n2571_ = ~new_n1689_ & ~new_n2026_;
  assign new_n2572_ = pv246_0_ & new_n2571_;
  assign new_n2573_ = ~new_n1689_ & new_n2026_;
  assign new_n2574_ = ~pv246_0_ & new_n2573_;
  assign pv603_0_ = new_n2572_ | new_n2574_;
  assign new_n2576_ = pv7_0_ & new_n2060_;
  assign pv1378 = new_n692_ & new_n2576_;
  assign new_n2578_ = pv1243_4_ & new_n2294_;
  assign new_n2579_ = pv199_1_ & pv199_3_;
  assign new_n2580_ = pv199_2_ & new_n2579_;
  assign new_n2581_ = pv199_0_ & new_n2580_;
  assign new_n2582_ = pv199_4_ & new_n2581_;
  assign new_n2583_ = pv194_4_ & ~new_n2582_;
  assign new_n2584_ = ~pv194_4_ & new_n2582_;
  assign new_n2585_ = ~new_n2583_ & ~new_n2584_;
  assign new_n2586_ = new_n2301_ & ~new_n2585_;
  assign pv572_4_ = new_n2578_ | new_n2586_;
  assign new_n2588_ = pv149_4_ & new_n2230_;
  assign new_n2589_ = pv279_0_ & ~new_n2230_;
  assign new_n2590_ = pv280_0_ & new_n2589_;
  assign new_n2591_ = ~pv280_0_ & new_n2231_;
  assign new_n2592_ = ~new_n2588_ & ~new_n2590_;
  assign pv826_0_ = new_n2591_ | ~new_n2592_;
  assign new_n2594_ = ~pv802_0_ & new_n702_;
  assign new_n2595_ = ~pv289_0_ & new_n2594_;
  assign new_n2596_ = pv262_0_ & new_n2363_;
  assign new_n2597_ = new_n615_ & ~new_n2596_;
  assign new_n2598_ = ~new_n1095_ & ~new_n1588_;
  assign new_n2599_ = ~new_n1096_ & ~new_n1718_;
  assign new_n2600_ = new_n2598_ & new_n2599_;
  assign new_n2601_ = ~new_n1224_ & ~new_n2321_;
  assign new_n2602_ = new_n2597_ & new_n2601_;
  assign new_n2603_ = new_n2600_ & new_n2602_;
  assign new_n2604_ = pv1741_0_ & new_n2603_;
  assign new_n2605_ = ~pv289_0_ & new_n2604_;
  assign new_n2606_ = ~new_n1132_ & new_n2597_;
  assign new_n2607_ = ~new_n1133_ & new_n2606_;
  assign new_n2608_ = new_n2603_ & new_n2607_;
  assign new_n2609_ = ~new_n1223_ & new_n2608_;
  assign new_n2610_ = ~new_n701_ & ~new_n2609_;
  assign new_n2611_ = new_n2545_ & new_n2610_;
  assign new_n2612_ = new_n755_ & new_n2611_;
  assign new_n2613_ = ~pv289_0_ & new_n2612_;
  assign new_n2614_ = ~new_n2595_ & ~new_n2605_;
  assign new_n2615_ = ~new_n2613_ & new_n2614_;
  assign pv1669 = ~new_n2375_ & new_n2615_;
  assign new_n2617_ = pv199_1_ & pv194_4_;
  assign new_n2618_ = pv199_2_ & new_n2617_;
  assign new_n2619_ = pv199_0_ & new_n2618_;
  assign new_n2620_ = pv199_4_ & new_n2619_;
  assign new_n2621_ = pv199_3_ & new_n2620_;
  assign new_n2622_ = pv194_3_ & ~new_n2621_;
  assign new_n2623_ = ~pv194_3_ & new_n2621_;
  assign new_n2624_ = ~new_n2622_ & ~new_n2623_;
  assign new_n2625_ = new_n2301_ & ~new_n2624_;
  assign new_n2626_ = pv149_7_ & new_n2488_;
  assign new_n2627_ = pv1243_3_ & new_n2294_;
  assign new_n2628_ = ~new_n2625_ & ~new_n2626_;
  assign pv572_3_ = new_n2627_ | ~new_n2628_;
  assign new_n2630_ = pv244_0_ & pv587;
  assign new_n2631_ = pv243_0_ & ~new_n1689_;
  assign new_n2632_ = ~pv244_0_ & new_n2631_;
  assign pv591_0_ = new_n2630_ | new_n2632_;
  assign new_n2634_ = new_n579_ & ~new_n586_;
  assign new_n2635_ = pv802_0_ & ~new_n2530_;
  assign new_n2636_ = pv763 & ~new_n1701_;
  assign new_n2637_ = ~new_n586_ & new_n2636_;
  assign new_n2638_ = pv56_0_ & new_n2637_;
  assign new_n2639_ = pv56_0_ & ~new_n2519_;
  assign new_n2640_ = ~new_n2634_ & ~new_n2635_;
  assign new_n2641_ = ~new_n2638_ & ~new_n2639_;
  assign new_n2642_ = new_n2640_ & new_n2641_;
  assign pv966 = new_n1628_ & ~new_n2642_;
  assign new_n2644_ = pv100_5_ & new_n2308_;
  assign new_n2645_ = ~new_n2307_ & new_n2644_;
  assign new_n2646_ = pv165_7_ & new_n2306_;
  assign pv1709_4_ = new_n2645_ | new_n2646_;
  assign new_n2648_ = pv248_0_ & pv1719;
  assign new_n2649_ = ~pv423_0_ & ~new_n2648_;
  assign new_n2650_ = ~pv43_0_ & ~new_n2411_;
  assign new_n2651_ = ~new_n2414_ & new_n2650_;
  assign new_n2652_ = ~new_n2649_ & new_n2651_;
  assign new_n2653_ = ~pv214_0_ & new_n2652_;
  assign new_n2654_ = ~new_n2030_ & new_n2653_;
  assign new_n2655_ = ~new_n2024_ & new_n2654_;
  assign new_n2656_ = ~new_n2410_ & new_n2655_;
  assign new_n2657_ = ~new_n2412_ & new_n2656_;
  assign pv398_0_ = new_n2032_ | ~new_n2657_;
  assign new_n2659_ = pv194_4_ & pv194_3_;
  assign new_n2660_ = pv199_2_ & new_n2659_;
  assign new_n2661_ = pv199_0_ & new_n2660_;
  assign new_n2662_ = pv199_4_ & new_n2661_;
  assign new_n2663_ = pv199_1_ & new_n2662_;
  assign new_n2664_ = pv199_3_ & new_n2663_;
  assign new_n2665_ = pv194_2_ & ~new_n2664_;
  assign new_n2666_ = ~pv194_2_ & new_n2664_;
  assign new_n2667_ = ~new_n2665_ & ~new_n2666_;
  assign new_n2668_ = new_n2301_ & ~new_n2667_;
  assign new_n2669_ = pv149_6_ & new_n2488_;
  assign new_n2670_ = pv1243_2_ & new_n2294_;
  assign new_n2671_ = ~new_n2668_ & ~new_n2669_;
  assign pv572_2_ = new_n2670_ | ~new_n2671_;
  assign pv640_0_ = pv271_0_ | new_n1525_;
  assign new_n2674_ = new_n755_ & new_n1699_;
  assign new_n2675_ = pv1536_0_ & ~new_n2674_;
  assign new_n2676_ = ~new_n1842_ & new_n1926_;
  assign new_n2677_ = ~new_n939_ & new_n2676_;
  assign new_n2678_ = ~new_n1005_ & new_n2677_;
  assign new_n2679_ = ~new_n1031_ & new_n2678_;
  assign new_n2680_ = ~new_n1083_ & new_n2679_;
  assign new_n2681_ = ~new_n1825_ & new_n2680_;
  assign new_n2682_ = ~pv1536_0_ & ~new_n2681_;
  assign pv1512_1_ = new_n2675_ | new_n2682_;
  assign new_n2684_ = pv100_4_ & new_n2308_;
  assign new_n2685_ = ~new_n2307_ & new_n2684_;
  assign new_n2686_ = pv165_6_ & new_n2306_;
  assign pv1709_3_ = new_n2685_ | new_n2686_;
  assign new_n2688_ = pv194_3_ & pv194_2_;
  assign new_n2689_ = pv199_2_ & new_n2688_;
  assign new_n2690_ = pv199_0_ & new_n2689_;
  assign new_n2691_ = pv199_4_ & new_n2690_;
  assign new_n2692_ = pv199_3_ & new_n2691_;
  assign new_n2693_ = pv194_4_ & new_n2692_;
  assign new_n2694_ = pv199_1_ & new_n2693_;
  assign new_n2695_ = pv194_1_ & ~new_n2694_;
  assign new_n2696_ = ~pv194_1_ & new_n2694_;
  assign new_n2697_ = ~new_n2695_ & ~new_n2696_;
  assign new_n2698_ = new_n2301_ & ~new_n2697_;
  assign new_n2699_ = pv149_5_ & new_n2488_;
  assign new_n2700_ = pv1243_1_ & new_n2294_;
  assign new_n2701_ = ~new_n2698_ & ~new_n2699_;
  assign pv572_1_ = new_n2700_ | ~new_n2701_;
  assign new_n2703_ = new_n2519_ & ~new_n2638_;
  assign new_n2704_ = new_n2541_ & new_n2703_;
  assign new_n2705_ = pv56_0_ & new_n2704_;
  assign new_n2706_ = pv62_0_ & ~new_n616_;
  assign new_n2707_ = ~new_n494_ & new_n640_;
  assign new_n2708_ = ~new_n1280_ & new_n2707_;
  assign new_n2709_ = pv59_0_ & ~new_n2708_;
  assign new_n2710_ = ~new_n2705_ & ~new_n2706_;
  assign new_n2711_ = ~new_n2709_ & new_n2710_;
  assign pv986 = new_n1628_ & ~new_n2711_;
  assign new_n2713_ = ~new_n1491_ & ~new_n1662_;
  assign new_n2714_ = pv258_0_ & pv14_0_;
  assign new_n2715_ = new_n2713_ & new_n2714_;
  assign new_n2716_ = ~pv258_0_ & pv14_0_;
  assign new_n2717_ = ~new_n2713_ & new_n2716_;
  assign pv1451_0_ = new_n2715_ | new_n2717_;
  assign new_n2719_ = new_n755_ & ~new_n793_;
  assign new_n2720_ = ~new_n1699_ & new_n2719_;
  assign new_n2721_ = pv1536_0_ & ~new_n2720_;
  assign new_n2722_ = ~new_n1842_ & new_n2009_;
  assign new_n2723_ = ~new_n956_ & new_n2722_;
  assign new_n2724_ = ~new_n1005_ & new_n2723_;
  assign new_n2725_ = ~new_n1031_ & new_n2724_;
  assign new_n2726_ = ~new_n1057_ & new_n2725_;
  assign new_n2727_ = ~new_n1825_ & new_n2726_;
  assign new_n2728_ = ~pv1536_0_ & ~new_n2727_;
  assign pv1512_2_ = new_n2721_ | new_n2728_;
  assign new_n2730_ = pv1921_1_ & ~pv1921_0_;
  assign new_n2731_ = ~pv1921_1_ & pv1921_0_;
  assign new_n2732_ = ~new_n2730_ & ~new_n2731_;
  assign new_n2733_ = pv1921_3_ & ~pv1921_2_;
  assign new_n2734_ = ~pv1921_3_ & pv1921_2_;
  assign new_n2735_ = ~new_n2733_ & ~new_n2734_;
  assign new_n2736_ = new_n2732_ & ~new_n2735_;
  assign new_n2737_ = ~new_n2732_ & new_n2735_;
  assign new_n2738_ = ~new_n2736_ & ~new_n2737_;
  assign new_n2739_ = pv1921_5_ & ~pv1921_4_;
  assign new_n2740_ = ~pv1921_5_ & pv1921_4_;
  assign new_n2741_ = ~new_n2739_ & ~new_n2740_;
  assign new_n2742_ = ~pv1953_0_ & pv1953_1_;
  assign new_n2743_ = pv1953_0_ & ~pv1953_1_;
  assign new_n2744_ = ~new_n2742_ & ~new_n2743_;
  assign new_n2745_ = new_n2741_ & ~new_n2744_;
  assign new_n2746_ = ~new_n2741_ & new_n2744_;
  assign new_n2747_ = ~new_n2745_ & ~new_n2746_;
  assign new_n2748_ = new_n2738_ & ~new_n2747_;
  assign new_n2749_ = ~new_n2738_ & new_n2747_;
  assign pv1613_0_ = ~new_n2748_ & ~new_n2749_;
  assign new_n2751_ = pv100_3_ & new_n2308_;
  assign new_n2752_ = ~new_n2307_ & new_n2751_;
  assign new_n2753_ = pv165_5_ & new_n2306_;
  assign pv1709_2_ = new_n2752_ | new_n2753_;
  assign pv1243_0_ = ~pv321_2_;
  assign pv657 = ~pv257_7_;
  assign pv1375 = ~pv268_5_;
  assign pv1481_0_ = ~pv214_0_;
  assign pv1671_0_ = ~pv205_0_;
  assign pv1863_0_ = ~pv301_0_;
  assign pv1864_0_ = ~pv302_0_;
  assign pv585_0_ = ~pv34_0_;
  assign pv1760_0_ = ~pv101_0_;
  assign pv1833_0_ = ~pv261_0_;
  assign pv1495_0_ = ~pv175_0_;
endmodule

