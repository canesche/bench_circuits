module i7 ( 
    \V199(1) , \V32(27) , \V199(0) , \V32(26) , \V32(25) , \V32(24) ,
    \V32(23) , \V32(22) , \V32(21) , \V32(20) , \V32(19) , \V32(18) ,
    \V32(17) , \V32(16) , \V32(15) , \V32(14) , \V32(13) , \V32(12) ,
    \V32(11) , \V32(10) , \V32(9) , \V32(8) , \V32(7) , \V32(6) , \V32(5) ,
    \V32(4) , \V32(3) , \V32(2) , \V32(1) , \V32(0) , \V96(27) , \V96(26) ,
    \V96(25) , \V96(24) , \V96(23) , \V96(22) , \V96(21) , \V96(20) ,
    \V96(19) , \V96(18) , \V96(17) , \V96(16) , \V96(15) , \V96(14) ,
    \V96(13) , \V96(12) , \V96(11) , \V96(10) , \V96(9) , \V96(8) ,
    \V96(7) , \V96(6) , \V96(5) , \V96(4) , \V96(3) , \V96(2) , \V96(1) ,
    \V96(0) , \V64(27) , \V64(26) , \V64(25) , \V64(24) , \V64(23) ,
    \V64(22) , \V64(21) , \V64(20) , \V64(19) , \V64(18) , \V64(17) ,
    \V64(16) , \V64(15) , \V64(14) , \V64(13) , \V64(12) , \V64(11) ,
    \V64(10) , \V64(9) , \V64(8) , \V64(7) , \V64(6) , \V64(5) , \V64(4) ,
    \V64(3) , \V64(2) , \V64(1) , \V64(0) , \V128(27) , \V199(4) ,
    \V128(26) , \V128(25) , \V128(24) , \V128(23) , \V128(22) , \V128(21) ,
    \V128(20) , \V128(19) , \V128(18) , \V128(17) , \V128(16) , \V128(15) ,
    \V128(14) , \V128(13) , \V128(12) , \V128(11) , \V128(10) , \V128(9) ,
    \V128(8) , \V128(7) , \V128(6) , \V128(5) , \V128(4) , \V128(3) ,
    \V128(2) , \V128(1) , \V128(0) , \V32(31) , \V32(30) , \V32(29) ,
    \V32(28) , \V192(27) , \V192(26) , \V192(25) , \V192(24) , \V192(23) ,
    \V192(22) , \V192(21) , \V192(20) , \V192(19) , \V192(18) , \V192(17) ,
    \V192(16) , \V192(15) , \V192(14) , \V192(13) , \V192(12) , \V192(11) ,
    \V192(10) , \V192(9) , \V192(8) , \V192(7) , \V192(6) , \V192(5) ,
    \V192(4) , \V192(3) , \V192(2) , \V192(1) , \V192(0) , \V96(31) ,
    \V96(30) , \V96(29) , \V96(28) , \V160(27) , \V160(26) , \V160(25) ,
    \V160(24) , \V160(23) , \V160(22) , \V160(21) , \V160(20) , \V160(19) ,
    \V160(18) , \V160(17) , \V160(16) , \V160(15) , \V160(14) , \V160(13) ,
    \V160(12) , \V160(11) , \V160(10) , \V160(9) , \V160(8) , \V160(7) ,
    \V160(6) , \V160(5) , \V160(4) , \V160(3) , \V160(2) , \V160(1) ,
    \V160(0) , \V64(31) , \V64(30) , \V64(29) , \V64(28) , \V128(31) ,
    \V199(3) , \V128(30) , \V128(29) , \V128(28) , \V195(0) , \V194(1) ,
    \V194(0) , \V192(31) , \V192(30) , \V192(29) , \V192(28) , \V160(31) ,
    \V160(30) , \V160(29) , \V160(28) ,
    \V227(27) , \V227(26) , \V227(25) , \V227(24) , \V227(23) , \V227(22) ,
    \V227(21) , \V227(20) , \V227(19) , \V227(18) , \V227(17) , \V227(16) ,
    \V227(15) , \V227(14) , \V227(13) , \V227(12) , \V227(11) , \V227(10) ,
    \V227(9) , \V227(8) , \V227(7) , \V227(6) , \V227(5) , \V227(4) ,
    \V227(3) , \V227(2) , \V227(1) , \V227(0) , \V259(31) , \V259(30) ,
    \V259(29) , \V259(28) , \V259(27) , \V259(26) , \V259(25) , \V259(24) ,
    \V259(23) , \V259(22) , \V259(21) , \V259(20) , \V259(19) , \V259(18) ,
    \V259(17) , \V259(16) , \V259(15) , \V259(14) , \V259(13) , \V259(12) ,
    \V259(11) , \V259(10) , \V259(9) , \V259(8) , \V259(7) , \V259(6) ,
    \V259(5) , \V259(4) , \V259(3) , \V259(2) , \V259(1) , \V259(0) ,
    \V266(6) , \V266(5) , \V266(4) , \V266(3) , \V266(2) , \V266(1) ,
    \V266(0)   );
  input  \V199(1) , \V32(27) , \V199(0) , \V32(26) , \V32(25) ,
    \V32(24) , \V32(23) , \V32(22) , \V32(21) , \V32(20) , \V32(19) ,
    \V32(18) , \V32(17) , \V32(16) , \V32(15) , \V32(14) , \V32(13) ,
    \V32(12) , \V32(11) , \V32(10) , \V32(9) , \V32(8) , \V32(7) ,
    \V32(6) , \V32(5) , \V32(4) , \V32(3) , \V32(2) , \V32(1) , \V32(0) ,
    \V96(27) , \V96(26) , \V96(25) , \V96(24) , \V96(23) , \V96(22) ,
    \V96(21) , \V96(20) , \V96(19) , \V96(18) , \V96(17) , \V96(16) ,
    \V96(15) , \V96(14) , \V96(13) , \V96(12) , \V96(11) , \V96(10) ,
    \V96(9) , \V96(8) , \V96(7) , \V96(6) , \V96(5) , \V96(4) , \V96(3) ,
    \V96(2) , \V96(1) , \V96(0) , \V64(27) , \V64(26) , \V64(25) ,
    \V64(24) , \V64(23) , \V64(22) , \V64(21) , \V64(20) , \V64(19) ,
    \V64(18) , \V64(17) , \V64(16) , \V64(15) , \V64(14) , \V64(13) ,
    \V64(12) , \V64(11) , \V64(10) , \V64(9) , \V64(8) , \V64(7) ,
    \V64(6) , \V64(5) , \V64(4) , \V64(3) , \V64(2) , \V64(1) , \V64(0) ,
    \V128(27) , \V199(4) , \V128(26) , \V128(25) , \V128(24) , \V128(23) ,
    \V128(22) , \V128(21) , \V128(20) , \V128(19) , \V128(18) , \V128(17) ,
    \V128(16) , \V128(15) , \V128(14) , \V128(13) , \V128(12) , \V128(11) ,
    \V128(10) , \V128(9) , \V128(8) , \V128(7) , \V128(6) , \V128(5) ,
    \V128(4) , \V128(3) , \V128(2) , \V128(1) , \V128(0) , \V32(31) ,
    \V32(30) , \V32(29) , \V32(28) , \V192(27) , \V192(26) , \V192(25) ,
    \V192(24) , \V192(23) , \V192(22) , \V192(21) , \V192(20) , \V192(19) ,
    \V192(18) , \V192(17) , \V192(16) , \V192(15) , \V192(14) , \V192(13) ,
    \V192(12) , \V192(11) , \V192(10) , \V192(9) , \V192(8) , \V192(7) ,
    \V192(6) , \V192(5) , \V192(4) , \V192(3) , \V192(2) , \V192(1) ,
    \V192(0) , \V96(31) , \V96(30) , \V96(29) , \V96(28) , \V160(27) ,
    \V160(26) , \V160(25) , \V160(24) , \V160(23) , \V160(22) , \V160(21) ,
    \V160(20) , \V160(19) , \V160(18) , \V160(17) , \V160(16) , \V160(15) ,
    \V160(14) , \V160(13) , \V160(12) , \V160(11) , \V160(10) , \V160(9) ,
    \V160(8) , \V160(7) , \V160(6) , \V160(5) , \V160(4) , \V160(3) ,
    \V160(2) , \V160(1) , \V160(0) , \V64(31) , \V64(30) , \V64(29) ,
    \V64(28) , \V128(31) , \V199(3) , \V128(30) , \V128(29) , \V128(28) ,
    \V195(0) , \V194(1) , \V194(0) , \V192(31) , \V192(30) , \V192(29) ,
    \V192(28) , \V160(31) , \V160(30) , \V160(29) , \V160(28) ;
  output \V227(27) , \V227(26) , \V227(25) , \V227(24) , \V227(23) ,
    \V227(22) , \V227(21) , \V227(20) , \V227(19) , \V227(18) , \V227(17) ,
    \V227(16) , \V227(15) , \V227(14) , \V227(13) , \V227(12) , \V227(11) ,
    \V227(10) , \V227(9) , \V227(8) , \V227(7) , \V227(6) , \V227(5) ,
    \V227(4) , \V227(3) , \V227(2) , \V227(1) , \V227(0) , \V259(31) ,
    \V259(30) , \V259(29) , \V259(28) , \V259(27) , \V259(26) , \V259(25) ,
    \V259(24) , \V259(23) , \V259(22) , \V259(21) , \V259(20) , \V259(19) ,
    \V259(18) , \V259(17) , \V259(16) , \V259(15) , \V259(14) , \V259(13) ,
    \V259(12) , \V259(11) , \V259(10) , \V259(9) , \V259(8) , \V259(7) ,
    \V259(6) , \V259(5) , \V259(4) , \V259(3) , \V259(2) , \V259(1) ,
    \V259(0) , \V266(6) , \V266(5) , \V266(4) , \V266(3) , \V266(2) ,
    \V266(1) , \V266(0) ;
  wire new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_;
  assign new_n267_ = ~\V199(1)  & \V32(27) ;
  assign new_n268_ = \V199(0)  & new_n267_;
  assign new_n269_ = ~\V199(1)  & \V96(27) ;
  assign new_n270_ = ~\V199(0)  & new_n269_;
  assign new_n271_ = \V199(1)  & \V64(27) ;
  assign new_n272_ = \V199(0)  & new_n271_;
  assign new_n273_ = \V199(1)  & ~\V96(27) ;
  assign new_n274_ = ~\V199(0)  & new_n273_;
  assign new_n275_ = ~new_n272_ & ~new_n274_;
  assign new_n276_ = ~new_n268_ & ~new_n270_;
  assign \V227(27)  = ~new_n275_ | ~new_n276_;
  assign new_n278_ = ~\V199(1)  & \V32(26) ;
  assign new_n279_ = \V199(0)  & new_n278_;
  assign new_n280_ = ~\V199(1)  & \V96(26) ;
  assign new_n281_ = ~\V199(0)  & new_n280_;
  assign new_n282_ = \V199(1)  & \V64(26) ;
  assign new_n283_ = \V199(0)  & new_n282_;
  assign new_n284_ = \V199(1)  & ~\V96(26) ;
  assign new_n285_ = ~\V199(0)  & new_n284_;
  assign new_n286_ = ~new_n283_ & ~new_n285_;
  assign new_n287_ = ~new_n279_ & ~new_n281_;
  assign \V227(26)  = ~new_n286_ | ~new_n287_;
  assign new_n289_ = ~\V199(1)  & \V32(25) ;
  assign new_n290_ = \V199(0)  & new_n289_;
  assign new_n291_ = ~\V199(1)  & \V96(25) ;
  assign new_n292_ = ~\V199(0)  & new_n291_;
  assign new_n293_ = \V199(1)  & \V64(25) ;
  assign new_n294_ = \V199(0)  & new_n293_;
  assign new_n295_ = \V199(1)  & ~\V96(25) ;
  assign new_n296_ = ~\V199(0)  & new_n295_;
  assign new_n297_ = ~new_n294_ & ~new_n296_;
  assign new_n298_ = ~new_n290_ & ~new_n292_;
  assign \V227(25)  = ~new_n297_ | ~new_n298_;
  assign new_n300_ = ~\V199(1)  & \V32(24) ;
  assign new_n301_ = \V199(0)  & new_n300_;
  assign new_n302_ = ~\V199(1)  & \V96(24) ;
  assign new_n303_ = ~\V199(0)  & new_n302_;
  assign new_n304_ = \V199(1)  & \V64(24) ;
  assign new_n305_ = \V199(0)  & new_n304_;
  assign new_n306_ = \V199(1)  & ~\V96(24) ;
  assign new_n307_ = ~\V199(0)  & new_n306_;
  assign new_n308_ = ~new_n305_ & ~new_n307_;
  assign new_n309_ = ~new_n301_ & ~new_n303_;
  assign \V227(24)  = ~new_n308_ | ~new_n309_;
  assign new_n311_ = ~\V199(1)  & \V32(23) ;
  assign new_n312_ = \V199(0)  & new_n311_;
  assign new_n313_ = ~\V199(1)  & \V96(23) ;
  assign new_n314_ = ~\V199(0)  & new_n313_;
  assign new_n315_ = \V199(1)  & \V64(23) ;
  assign new_n316_ = \V199(0)  & new_n315_;
  assign new_n317_ = \V199(1)  & ~\V96(23) ;
  assign new_n318_ = ~\V199(0)  & new_n317_;
  assign new_n319_ = ~new_n316_ & ~new_n318_;
  assign new_n320_ = ~new_n312_ & ~new_n314_;
  assign \V227(23)  = ~new_n319_ | ~new_n320_;
  assign new_n322_ = ~\V199(1)  & \V32(22) ;
  assign new_n323_ = \V199(0)  & new_n322_;
  assign new_n324_ = ~\V199(1)  & \V96(22) ;
  assign new_n325_ = ~\V199(0)  & new_n324_;
  assign new_n326_ = \V199(1)  & \V64(22) ;
  assign new_n327_ = \V199(0)  & new_n326_;
  assign new_n328_ = \V199(1)  & ~\V96(22) ;
  assign new_n329_ = ~\V199(0)  & new_n328_;
  assign new_n330_ = ~new_n327_ & ~new_n329_;
  assign new_n331_ = ~new_n323_ & ~new_n325_;
  assign \V227(22)  = ~new_n330_ | ~new_n331_;
  assign new_n333_ = ~\V199(1)  & \V32(21) ;
  assign new_n334_ = \V199(0)  & new_n333_;
  assign new_n335_ = ~\V199(1)  & \V96(21) ;
  assign new_n336_ = ~\V199(0)  & new_n335_;
  assign new_n337_ = \V199(1)  & \V64(21) ;
  assign new_n338_ = \V199(0)  & new_n337_;
  assign new_n339_ = \V199(1)  & ~\V96(21) ;
  assign new_n340_ = ~\V199(0)  & new_n339_;
  assign new_n341_ = ~new_n338_ & ~new_n340_;
  assign new_n342_ = ~new_n334_ & ~new_n336_;
  assign \V227(21)  = ~new_n341_ | ~new_n342_;
  assign new_n344_ = ~\V199(1)  & \V32(20) ;
  assign new_n345_ = \V199(0)  & new_n344_;
  assign new_n346_ = ~\V199(1)  & \V96(20) ;
  assign new_n347_ = ~\V199(0)  & new_n346_;
  assign new_n348_ = \V199(1)  & \V64(20) ;
  assign new_n349_ = \V199(0)  & new_n348_;
  assign new_n350_ = \V199(1)  & ~\V96(20) ;
  assign new_n351_ = ~\V199(0)  & new_n350_;
  assign new_n352_ = ~new_n349_ & ~new_n351_;
  assign new_n353_ = ~new_n345_ & ~new_n347_;
  assign \V227(20)  = ~new_n352_ | ~new_n353_;
  assign new_n355_ = ~\V199(1)  & \V32(19) ;
  assign new_n356_ = \V199(0)  & new_n355_;
  assign new_n357_ = ~\V199(1)  & \V96(19) ;
  assign new_n358_ = ~\V199(0)  & new_n357_;
  assign new_n359_ = \V199(1)  & \V64(19) ;
  assign new_n360_ = \V199(0)  & new_n359_;
  assign new_n361_ = \V199(1)  & ~\V96(19) ;
  assign new_n362_ = ~\V199(0)  & new_n361_;
  assign new_n363_ = ~new_n360_ & ~new_n362_;
  assign new_n364_ = ~new_n356_ & ~new_n358_;
  assign \V227(19)  = ~new_n363_ | ~new_n364_;
  assign new_n366_ = ~\V199(1)  & \V32(18) ;
  assign new_n367_ = \V199(0)  & new_n366_;
  assign new_n368_ = ~\V199(1)  & \V96(18) ;
  assign new_n369_ = ~\V199(0)  & new_n368_;
  assign new_n370_ = \V199(1)  & \V64(18) ;
  assign new_n371_ = \V199(0)  & new_n370_;
  assign new_n372_ = \V199(1)  & ~\V96(18) ;
  assign new_n373_ = ~\V199(0)  & new_n372_;
  assign new_n374_ = ~new_n371_ & ~new_n373_;
  assign new_n375_ = ~new_n367_ & ~new_n369_;
  assign \V227(18)  = ~new_n374_ | ~new_n375_;
  assign new_n377_ = ~\V199(1)  & \V32(17) ;
  assign new_n378_ = \V199(0)  & new_n377_;
  assign new_n379_ = ~\V199(1)  & \V96(17) ;
  assign new_n380_ = ~\V199(0)  & new_n379_;
  assign new_n381_ = \V199(1)  & \V64(17) ;
  assign new_n382_ = \V199(0)  & new_n381_;
  assign new_n383_ = \V199(1)  & ~\V96(17) ;
  assign new_n384_ = ~\V199(0)  & new_n383_;
  assign new_n385_ = ~new_n382_ & ~new_n384_;
  assign new_n386_ = ~new_n378_ & ~new_n380_;
  assign \V227(17)  = ~new_n385_ | ~new_n386_;
  assign new_n388_ = ~\V199(1)  & \V32(16) ;
  assign new_n389_ = \V199(0)  & new_n388_;
  assign new_n390_ = ~\V199(1)  & \V96(16) ;
  assign new_n391_ = ~\V199(0)  & new_n390_;
  assign new_n392_ = \V199(1)  & \V64(16) ;
  assign new_n393_ = \V199(0)  & new_n392_;
  assign new_n394_ = \V199(1)  & ~\V96(16) ;
  assign new_n395_ = ~\V199(0)  & new_n394_;
  assign new_n396_ = ~new_n393_ & ~new_n395_;
  assign new_n397_ = ~new_n389_ & ~new_n391_;
  assign \V227(16)  = ~new_n396_ | ~new_n397_;
  assign new_n399_ = ~\V199(1)  & \V32(15) ;
  assign new_n400_ = \V199(0)  & new_n399_;
  assign new_n401_ = ~\V199(1)  & \V96(15) ;
  assign new_n402_ = ~\V199(0)  & new_n401_;
  assign new_n403_ = \V199(1)  & \V64(15) ;
  assign new_n404_ = \V199(0)  & new_n403_;
  assign new_n405_ = \V199(1)  & ~\V96(15) ;
  assign new_n406_ = ~\V199(0)  & new_n405_;
  assign new_n407_ = ~new_n404_ & ~new_n406_;
  assign new_n408_ = ~new_n400_ & ~new_n402_;
  assign \V227(15)  = ~new_n407_ | ~new_n408_;
  assign new_n410_ = ~\V199(1)  & \V32(14) ;
  assign new_n411_ = \V199(0)  & new_n410_;
  assign new_n412_ = ~\V199(1)  & \V96(14) ;
  assign new_n413_ = ~\V199(0)  & new_n412_;
  assign new_n414_ = \V199(1)  & \V64(14) ;
  assign new_n415_ = \V199(0)  & new_n414_;
  assign new_n416_ = \V199(1)  & ~\V96(14) ;
  assign new_n417_ = ~\V199(0)  & new_n416_;
  assign new_n418_ = ~new_n415_ & ~new_n417_;
  assign new_n419_ = ~new_n411_ & ~new_n413_;
  assign \V227(14)  = ~new_n418_ | ~new_n419_;
  assign new_n421_ = ~\V199(1)  & \V32(13) ;
  assign new_n422_ = \V199(0)  & new_n421_;
  assign new_n423_ = ~\V199(1)  & \V96(13) ;
  assign new_n424_ = ~\V199(0)  & new_n423_;
  assign new_n425_ = \V199(1)  & \V64(13) ;
  assign new_n426_ = \V199(0)  & new_n425_;
  assign new_n427_ = \V199(1)  & ~\V96(13) ;
  assign new_n428_ = ~\V199(0)  & new_n427_;
  assign new_n429_ = ~new_n426_ & ~new_n428_;
  assign new_n430_ = ~new_n422_ & ~new_n424_;
  assign \V227(13)  = ~new_n429_ | ~new_n430_;
  assign new_n432_ = ~\V199(1)  & \V32(12) ;
  assign new_n433_ = \V199(0)  & new_n432_;
  assign new_n434_ = ~\V199(1)  & \V96(12) ;
  assign new_n435_ = ~\V199(0)  & new_n434_;
  assign new_n436_ = \V199(1)  & \V64(12) ;
  assign new_n437_ = \V199(0)  & new_n436_;
  assign new_n438_ = \V199(1)  & ~\V96(12) ;
  assign new_n439_ = ~\V199(0)  & new_n438_;
  assign new_n440_ = ~new_n437_ & ~new_n439_;
  assign new_n441_ = ~new_n433_ & ~new_n435_;
  assign \V227(12)  = ~new_n440_ | ~new_n441_;
  assign new_n443_ = ~\V199(1)  & \V32(11) ;
  assign new_n444_ = \V199(0)  & new_n443_;
  assign new_n445_ = ~\V199(1)  & \V96(11) ;
  assign new_n446_ = ~\V199(0)  & new_n445_;
  assign new_n447_ = \V199(1)  & \V64(11) ;
  assign new_n448_ = \V199(0)  & new_n447_;
  assign new_n449_ = \V199(1)  & ~\V96(11) ;
  assign new_n450_ = ~\V199(0)  & new_n449_;
  assign new_n451_ = ~new_n448_ & ~new_n450_;
  assign new_n452_ = ~new_n444_ & ~new_n446_;
  assign \V227(11)  = ~new_n451_ | ~new_n452_;
  assign new_n454_ = ~\V199(1)  & \V32(10) ;
  assign new_n455_ = \V199(0)  & new_n454_;
  assign new_n456_ = ~\V199(1)  & \V96(10) ;
  assign new_n457_ = ~\V199(0)  & new_n456_;
  assign new_n458_ = \V199(1)  & \V64(10) ;
  assign new_n459_ = \V199(0)  & new_n458_;
  assign new_n460_ = \V199(1)  & ~\V96(10) ;
  assign new_n461_ = ~\V199(0)  & new_n460_;
  assign new_n462_ = ~new_n459_ & ~new_n461_;
  assign new_n463_ = ~new_n455_ & ~new_n457_;
  assign \V227(10)  = ~new_n462_ | ~new_n463_;
  assign new_n465_ = ~\V199(1)  & \V32(9) ;
  assign new_n466_ = \V199(0)  & new_n465_;
  assign new_n467_ = ~\V199(1)  & \V96(9) ;
  assign new_n468_ = ~\V199(0)  & new_n467_;
  assign new_n469_ = \V199(1)  & \V64(9) ;
  assign new_n470_ = \V199(0)  & new_n469_;
  assign new_n471_ = \V199(1)  & ~\V96(9) ;
  assign new_n472_ = ~\V199(0)  & new_n471_;
  assign new_n473_ = ~new_n470_ & ~new_n472_;
  assign new_n474_ = ~new_n466_ & ~new_n468_;
  assign \V227(9)  = ~new_n473_ | ~new_n474_;
  assign new_n476_ = ~\V199(1)  & \V32(8) ;
  assign new_n477_ = \V199(0)  & new_n476_;
  assign new_n478_ = ~\V199(1)  & \V96(8) ;
  assign new_n479_ = ~\V199(0)  & new_n478_;
  assign new_n480_ = \V199(1)  & \V64(8) ;
  assign new_n481_ = \V199(0)  & new_n480_;
  assign new_n482_ = \V199(1)  & ~\V96(8) ;
  assign new_n483_ = ~\V199(0)  & new_n482_;
  assign new_n484_ = ~new_n481_ & ~new_n483_;
  assign new_n485_ = ~new_n477_ & ~new_n479_;
  assign \V227(8)  = ~new_n484_ | ~new_n485_;
  assign new_n487_ = ~\V199(1)  & \V32(7) ;
  assign new_n488_ = \V199(0)  & new_n487_;
  assign new_n489_ = ~\V199(1)  & \V96(7) ;
  assign new_n490_ = ~\V199(0)  & new_n489_;
  assign new_n491_ = \V199(1)  & \V64(7) ;
  assign new_n492_ = \V199(0)  & new_n491_;
  assign new_n493_ = \V199(1)  & ~\V96(7) ;
  assign new_n494_ = ~\V199(0)  & new_n493_;
  assign new_n495_ = ~new_n492_ & ~new_n494_;
  assign new_n496_ = ~new_n488_ & ~new_n490_;
  assign \V227(7)  = ~new_n495_ | ~new_n496_;
  assign new_n498_ = ~\V199(1)  & \V32(6) ;
  assign new_n499_ = \V199(0)  & new_n498_;
  assign new_n500_ = ~\V199(1)  & \V96(6) ;
  assign new_n501_ = ~\V199(0)  & new_n500_;
  assign new_n502_ = \V199(1)  & \V64(6) ;
  assign new_n503_ = \V199(0)  & new_n502_;
  assign new_n504_ = \V199(1)  & ~\V96(6) ;
  assign new_n505_ = ~\V199(0)  & new_n504_;
  assign new_n506_ = ~new_n503_ & ~new_n505_;
  assign new_n507_ = ~new_n499_ & ~new_n501_;
  assign \V227(6)  = ~new_n506_ | ~new_n507_;
  assign new_n509_ = ~\V199(1)  & \V32(5) ;
  assign new_n510_ = \V199(0)  & new_n509_;
  assign new_n511_ = ~\V199(1)  & \V96(5) ;
  assign new_n512_ = ~\V199(0)  & new_n511_;
  assign new_n513_ = \V199(1)  & \V64(5) ;
  assign new_n514_ = \V199(0)  & new_n513_;
  assign new_n515_ = \V199(1)  & ~\V96(5) ;
  assign new_n516_ = ~\V199(0)  & new_n515_;
  assign new_n517_ = ~new_n514_ & ~new_n516_;
  assign new_n518_ = ~new_n510_ & ~new_n512_;
  assign \V227(5)  = ~new_n517_ | ~new_n518_;
  assign new_n520_ = ~\V199(1)  & \V32(4) ;
  assign new_n521_ = \V199(0)  & new_n520_;
  assign new_n522_ = ~\V199(1)  & \V96(4) ;
  assign new_n523_ = ~\V199(0)  & new_n522_;
  assign new_n524_ = \V199(1)  & \V64(4) ;
  assign new_n525_ = \V199(0)  & new_n524_;
  assign new_n526_ = \V199(1)  & ~\V96(4) ;
  assign new_n527_ = ~\V199(0)  & new_n526_;
  assign new_n528_ = ~new_n525_ & ~new_n527_;
  assign new_n529_ = ~new_n521_ & ~new_n523_;
  assign \V227(4)  = ~new_n528_ | ~new_n529_;
  assign new_n531_ = ~\V199(1)  & \V32(3) ;
  assign new_n532_ = \V199(0)  & new_n531_;
  assign new_n533_ = ~\V199(1)  & \V96(3) ;
  assign new_n534_ = ~\V199(0)  & new_n533_;
  assign new_n535_ = \V199(1)  & \V64(3) ;
  assign new_n536_ = \V199(0)  & new_n535_;
  assign new_n537_ = \V199(1)  & ~\V96(3) ;
  assign new_n538_ = ~\V199(0)  & new_n537_;
  assign new_n539_ = ~new_n536_ & ~new_n538_;
  assign new_n540_ = ~new_n532_ & ~new_n534_;
  assign \V227(3)  = ~new_n539_ | ~new_n540_;
  assign new_n542_ = ~\V199(1)  & \V32(2) ;
  assign new_n543_ = \V199(0)  & new_n542_;
  assign new_n544_ = ~\V199(1)  & \V96(2) ;
  assign new_n545_ = ~\V199(0)  & new_n544_;
  assign new_n546_ = \V199(1)  & \V64(2) ;
  assign new_n547_ = \V199(0)  & new_n546_;
  assign new_n548_ = \V199(1)  & ~\V96(2) ;
  assign new_n549_ = ~\V199(0)  & new_n548_;
  assign new_n550_ = ~new_n547_ & ~new_n549_;
  assign new_n551_ = ~new_n543_ & ~new_n545_;
  assign \V227(2)  = ~new_n550_ | ~new_n551_;
  assign new_n553_ = ~\V199(1)  & \V32(1) ;
  assign new_n554_ = \V199(0)  & new_n553_;
  assign new_n555_ = ~\V199(1)  & \V96(1) ;
  assign new_n556_ = ~\V199(0)  & new_n555_;
  assign new_n557_ = \V199(1)  & \V64(1) ;
  assign new_n558_ = \V199(0)  & new_n557_;
  assign new_n559_ = \V199(1)  & ~\V96(1) ;
  assign new_n560_ = ~\V199(0)  & new_n559_;
  assign new_n561_ = ~new_n558_ & ~new_n560_;
  assign new_n562_ = ~new_n554_ & ~new_n556_;
  assign \V227(1)  = ~new_n561_ | ~new_n562_;
  assign new_n564_ = ~\V199(1)  & \V32(0) ;
  assign new_n565_ = \V199(0)  & new_n564_;
  assign new_n566_ = ~\V199(1)  & \V96(0) ;
  assign new_n567_ = ~\V199(0)  & new_n566_;
  assign new_n568_ = \V199(1)  & \V64(0) ;
  assign new_n569_ = \V199(0)  & new_n568_;
  assign new_n570_ = \V199(1)  & ~\V96(0) ;
  assign new_n571_ = ~\V199(0)  & new_n570_;
  assign new_n572_ = ~new_n569_ & ~new_n571_;
  assign new_n573_ = ~new_n565_ & ~new_n567_;
  assign \V227(0)  = ~new_n572_ | ~new_n573_;
  assign new_n575_ = \V199(0)  & \V128(27) ;
  assign new_n576_ = ~\V199(1)  & new_n575_;
  assign new_n577_ = \V199(4)  & new_n576_;
  assign new_n578_ = ~\V199(0)  & \V192(27) ;
  assign new_n579_ = ~\V199(1)  & new_n578_;
  assign new_n580_ = \V199(4)  & new_n579_;
  assign new_n581_ = \V199(0)  & \V160(27) ;
  assign new_n582_ = \V199(1)  & new_n581_;
  assign new_n583_ = \V199(4)  & new_n582_;
  assign new_n584_ = ~\V199(0)  & ~\V192(27) ;
  assign new_n585_ = \V199(1)  & new_n584_;
  assign new_n586_ = \V199(4)  & new_n585_;
  assign new_n587_ = \V199(1)  & ~\V199(4) ;
  assign new_n588_ = ~new_n586_ & ~new_n587_;
  assign new_n589_ = ~new_n577_ & ~new_n580_;
  assign new_n590_ = ~new_n583_ & new_n589_;
  assign \V259(31)  = ~new_n588_ | ~new_n590_;
  assign new_n592_ = \V199(0)  & \V128(26) ;
  assign new_n593_ = ~\V199(1)  & new_n592_;
  assign new_n594_ = \V199(4)  & new_n593_;
  assign new_n595_ = ~\V199(0)  & \V192(26) ;
  assign new_n596_ = ~\V199(1)  & new_n595_;
  assign new_n597_ = \V199(4)  & new_n596_;
  assign new_n598_ = \V199(0)  & \V160(26) ;
  assign new_n599_ = \V199(1)  & new_n598_;
  assign new_n600_ = \V199(4)  & new_n599_;
  assign new_n601_ = ~\V199(0)  & ~\V192(26) ;
  assign new_n602_ = \V199(1)  & new_n601_;
  assign new_n603_ = \V199(4)  & new_n602_;
  assign new_n604_ = ~new_n587_ & ~new_n603_;
  assign new_n605_ = ~new_n594_ & ~new_n597_;
  assign new_n606_ = ~new_n600_ & new_n605_;
  assign \V259(30)  = ~new_n604_ | ~new_n606_;
  assign new_n608_ = \V199(0)  & \V128(25) ;
  assign new_n609_ = ~\V199(1)  & new_n608_;
  assign new_n610_ = \V199(4)  & new_n609_;
  assign new_n611_ = ~\V199(0)  & \V192(25) ;
  assign new_n612_ = ~\V199(1)  & new_n611_;
  assign new_n613_ = \V199(4)  & new_n612_;
  assign new_n614_ = \V199(0)  & \V160(25) ;
  assign new_n615_ = \V199(1)  & new_n614_;
  assign new_n616_ = \V199(4)  & new_n615_;
  assign new_n617_ = ~\V199(0)  & ~\V192(25) ;
  assign new_n618_ = \V199(1)  & new_n617_;
  assign new_n619_ = \V199(4)  & new_n618_;
  assign new_n620_ = ~new_n587_ & ~new_n619_;
  assign new_n621_ = ~new_n610_ & ~new_n613_;
  assign new_n622_ = ~new_n616_ & new_n621_;
  assign \V259(29)  = ~new_n620_ | ~new_n622_;
  assign new_n624_ = \V199(0)  & \V128(24) ;
  assign new_n625_ = ~\V199(1)  & new_n624_;
  assign new_n626_ = \V199(4)  & new_n625_;
  assign new_n627_ = ~\V199(0)  & \V192(24) ;
  assign new_n628_ = ~\V199(1)  & new_n627_;
  assign new_n629_ = \V199(4)  & new_n628_;
  assign new_n630_ = \V199(0)  & \V160(24) ;
  assign new_n631_ = \V199(1)  & new_n630_;
  assign new_n632_ = \V199(4)  & new_n631_;
  assign new_n633_ = ~\V199(0)  & ~\V192(24) ;
  assign new_n634_ = \V199(1)  & new_n633_;
  assign new_n635_ = \V199(4)  & new_n634_;
  assign new_n636_ = ~new_n587_ & ~new_n635_;
  assign new_n637_ = ~new_n626_ & ~new_n629_;
  assign new_n638_ = ~new_n632_ & new_n637_;
  assign \V259(28)  = ~new_n636_ | ~new_n638_;
  assign new_n640_ = \V199(0)  & \V128(23) ;
  assign new_n641_ = ~\V199(1)  & new_n640_;
  assign new_n642_ = \V199(4)  & new_n641_;
  assign new_n643_ = ~\V199(0)  & \V192(23) ;
  assign new_n644_ = ~\V199(1)  & new_n643_;
  assign new_n645_ = \V199(4)  & new_n644_;
  assign new_n646_ = \V199(0)  & \V160(23) ;
  assign new_n647_ = \V199(1)  & new_n646_;
  assign new_n648_ = \V199(4)  & new_n647_;
  assign new_n649_ = ~\V199(0)  & ~\V192(23) ;
  assign new_n650_ = \V199(1)  & new_n649_;
  assign new_n651_ = \V199(4)  & new_n650_;
  assign new_n652_ = ~new_n587_ & ~new_n651_;
  assign new_n653_ = ~new_n642_ & ~new_n645_;
  assign new_n654_ = ~new_n648_ & new_n653_;
  assign \V259(27)  = ~new_n652_ | ~new_n654_;
  assign new_n656_ = \V199(0)  & \V128(22) ;
  assign new_n657_ = ~\V199(1)  & new_n656_;
  assign new_n658_ = \V199(4)  & new_n657_;
  assign new_n659_ = ~\V199(0)  & \V192(22) ;
  assign new_n660_ = ~\V199(1)  & new_n659_;
  assign new_n661_ = \V199(4)  & new_n660_;
  assign new_n662_ = \V199(0)  & \V160(22) ;
  assign new_n663_ = \V199(1)  & new_n662_;
  assign new_n664_ = \V199(4)  & new_n663_;
  assign new_n665_ = ~\V199(0)  & ~\V192(22) ;
  assign new_n666_ = \V199(1)  & new_n665_;
  assign new_n667_ = \V199(4)  & new_n666_;
  assign new_n668_ = ~new_n587_ & ~new_n667_;
  assign new_n669_ = ~new_n658_ & ~new_n661_;
  assign new_n670_ = ~new_n664_ & new_n669_;
  assign \V259(26)  = ~new_n668_ | ~new_n670_;
  assign new_n672_ = \V199(0)  & \V128(21) ;
  assign new_n673_ = ~\V199(1)  & new_n672_;
  assign new_n674_ = \V199(4)  & new_n673_;
  assign new_n675_ = ~\V199(0)  & \V192(21) ;
  assign new_n676_ = ~\V199(1)  & new_n675_;
  assign new_n677_ = \V199(4)  & new_n676_;
  assign new_n678_ = \V199(0)  & \V160(21) ;
  assign new_n679_ = \V199(1)  & new_n678_;
  assign new_n680_ = \V199(4)  & new_n679_;
  assign new_n681_ = ~\V199(0)  & ~\V192(21) ;
  assign new_n682_ = \V199(1)  & new_n681_;
  assign new_n683_ = \V199(4)  & new_n682_;
  assign new_n684_ = ~new_n587_ & ~new_n683_;
  assign new_n685_ = ~new_n674_ & ~new_n677_;
  assign new_n686_ = ~new_n680_ & new_n685_;
  assign \V259(25)  = ~new_n684_ | ~new_n686_;
  assign new_n688_ = \V199(0)  & \V128(20) ;
  assign new_n689_ = ~\V199(1)  & new_n688_;
  assign new_n690_ = \V199(4)  & new_n689_;
  assign new_n691_ = ~\V199(0)  & \V192(20) ;
  assign new_n692_ = ~\V199(1)  & new_n691_;
  assign new_n693_ = \V199(4)  & new_n692_;
  assign new_n694_ = \V199(0)  & \V160(20) ;
  assign new_n695_ = \V199(1)  & new_n694_;
  assign new_n696_ = \V199(4)  & new_n695_;
  assign new_n697_ = ~\V199(0)  & ~\V192(20) ;
  assign new_n698_ = \V199(1)  & new_n697_;
  assign new_n699_ = \V199(4)  & new_n698_;
  assign new_n700_ = ~new_n587_ & ~new_n699_;
  assign new_n701_ = ~new_n690_ & ~new_n693_;
  assign new_n702_ = ~new_n696_ & new_n701_;
  assign \V259(24)  = ~new_n700_ | ~new_n702_;
  assign new_n704_ = \V199(0)  & \V128(19) ;
  assign new_n705_ = ~\V199(1)  & new_n704_;
  assign new_n706_ = \V199(4)  & new_n705_;
  assign new_n707_ = ~\V199(0)  & \V192(19) ;
  assign new_n708_ = ~\V199(1)  & new_n707_;
  assign new_n709_ = \V199(4)  & new_n708_;
  assign new_n710_ = \V199(0)  & \V160(19) ;
  assign new_n711_ = \V199(1)  & new_n710_;
  assign new_n712_ = \V199(4)  & new_n711_;
  assign new_n713_ = ~\V199(0)  & ~\V192(19) ;
  assign new_n714_ = \V199(1)  & new_n713_;
  assign new_n715_ = \V199(4)  & new_n714_;
  assign new_n716_ = ~new_n587_ & ~new_n715_;
  assign new_n717_ = ~new_n706_ & ~new_n709_;
  assign new_n718_ = ~new_n712_ & new_n717_;
  assign \V259(23)  = ~new_n716_ | ~new_n718_;
  assign new_n720_ = \V199(0)  & \V128(18) ;
  assign new_n721_ = ~\V199(1)  & new_n720_;
  assign new_n722_ = \V199(4)  & new_n721_;
  assign new_n723_ = ~\V199(0)  & \V192(18) ;
  assign new_n724_ = ~\V199(1)  & new_n723_;
  assign new_n725_ = \V199(4)  & new_n724_;
  assign new_n726_ = \V199(0)  & \V160(18) ;
  assign new_n727_ = \V199(1)  & new_n726_;
  assign new_n728_ = \V199(4)  & new_n727_;
  assign new_n729_ = ~\V199(0)  & ~\V192(18) ;
  assign new_n730_ = \V199(1)  & new_n729_;
  assign new_n731_ = \V199(4)  & new_n730_;
  assign new_n732_ = ~new_n587_ & ~new_n731_;
  assign new_n733_ = ~new_n722_ & ~new_n725_;
  assign new_n734_ = ~new_n728_ & new_n733_;
  assign \V259(22)  = ~new_n732_ | ~new_n734_;
  assign new_n736_ = \V199(0)  & \V128(17) ;
  assign new_n737_ = ~\V199(1)  & new_n736_;
  assign new_n738_ = \V199(4)  & new_n737_;
  assign new_n739_ = ~\V199(0)  & \V192(17) ;
  assign new_n740_ = ~\V199(1)  & new_n739_;
  assign new_n741_ = \V199(4)  & new_n740_;
  assign new_n742_ = \V199(0)  & \V160(17) ;
  assign new_n743_ = \V199(1)  & new_n742_;
  assign new_n744_ = \V199(4)  & new_n743_;
  assign new_n745_ = ~\V199(0)  & ~\V192(17) ;
  assign new_n746_ = \V199(1)  & new_n745_;
  assign new_n747_ = \V199(4)  & new_n746_;
  assign new_n748_ = ~new_n587_ & ~new_n747_;
  assign new_n749_ = ~new_n738_ & ~new_n741_;
  assign new_n750_ = ~new_n744_ & new_n749_;
  assign \V259(21)  = ~new_n748_ | ~new_n750_;
  assign new_n752_ = \V199(0)  & \V128(16) ;
  assign new_n753_ = ~\V199(1)  & new_n752_;
  assign new_n754_ = \V199(4)  & new_n753_;
  assign new_n755_ = ~\V199(0)  & \V192(16) ;
  assign new_n756_ = ~\V199(1)  & new_n755_;
  assign new_n757_ = \V199(4)  & new_n756_;
  assign new_n758_ = \V199(0)  & \V160(16) ;
  assign new_n759_ = \V199(1)  & new_n758_;
  assign new_n760_ = \V199(4)  & new_n759_;
  assign new_n761_ = ~\V199(0)  & ~\V192(16) ;
  assign new_n762_ = \V199(1)  & new_n761_;
  assign new_n763_ = \V199(4)  & new_n762_;
  assign new_n764_ = ~new_n587_ & ~new_n763_;
  assign new_n765_ = ~new_n754_ & ~new_n757_;
  assign new_n766_ = ~new_n760_ & new_n765_;
  assign \V259(20)  = ~new_n764_ | ~new_n766_;
  assign new_n768_ = \V199(0)  & \V128(15) ;
  assign new_n769_ = ~\V199(1)  & new_n768_;
  assign new_n770_ = \V199(4)  & new_n769_;
  assign new_n771_ = ~\V199(0)  & \V192(15) ;
  assign new_n772_ = ~\V199(1)  & new_n771_;
  assign new_n773_ = \V199(4)  & new_n772_;
  assign new_n774_ = \V199(0)  & \V160(15) ;
  assign new_n775_ = \V199(1)  & new_n774_;
  assign new_n776_ = \V199(4)  & new_n775_;
  assign new_n777_ = ~\V199(0)  & ~\V192(15) ;
  assign new_n778_ = \V199(1)  & new_n777_;
  assign new_n779_ = \V199(4)  & new_n778_;
  assign new_n780_ = ~new_n587_ & ~new_n779_;
  assign new_n781_ = ~new_n770_ & ~new_n773_;
  assign new_n782_ = ~new_n776_ & new_n781_;
  assign \V259(19)  = ~new_n780_ | ~new_n782_;
  assign new_n784_ = \V199(0)  & \V128(14) ;
  assign new_n785_ = ~\V199(1)  & new_n784_;
  assign new_n786_ = \V199(4)  & new_n785_;
  assign new_n787_ = ~\V199(0)  & \V192(14) ;
  assign new_n788_ = ~\V199(1)  & new_n787_;
  assign new_n789_ = \V199(4)  & new_n788_;
  assign new_n790_ = \V199(0)  & \V160(14) ;
  assign new_n791_ = \V199(1)  & new_n790_;
  assign new_n792_ = \V199(4)  & new_n791_;
  assign new_n793_ = ~\V199(0)  & ~\V192(14) ;
  assign new_n794_ = \V199(1)  & new_n793_;
  assign new_n795_ = \V199(4)  & new_n794_;
  assign new_n796_ = ~new_n587_ & ~new_n795_;
  assign new_n797_ = ~new_n786_ & ~new_n789_;
  assign new_n798_ = ~new_n792_ & new_n797_;
  assign \V259(18)  = ~new_n796_ | ~new_n798_;
  assign new_n800_ = \V199(0)  & \V128(13) ;
  assign new_n801_ = ~\V199(1)  & new_n800_;
  assign new_n802_ = \V199(4)  & new_n801_;
  assign new_n803_ = ~\V199(0)  & \V192(13) ;
  assign new_n804_ = ~\V199(1)  & new_n803_;
  assign new_n805_ = \V199(4)  & new_n804_;
  assign new_n806_ = \V199(0)  & \V160(13) ;
  assign new_n807_ = \V199(1)  & new_n806_;
  assign new_n808_ = \V199(4)  & new_n807_;
  assign new_n809_ = ~\V199(0)  & ~\V192(13) ;
  assign new_n810_ = \V199(1)  & new_n809_;
  assign new_n811_ = \V199(4)  & new_n810_;
  assign new_n812_ = ~new_n587_ & ~new_n811_;
  assign new_n813_ = ~new_n802_ & ~new_n805_;
  assign new_n814_ = ~new_n808_ & new_n813_;
  assign \V259(17)  = ~new_n812_ | ~new_n814_;
  assign new_n816_ = \V199(0)  & \V128(12) ;
  assign new_n817_ = ~\V199(1)  & new_n816_;
  assign new_n818_ = \V199(4)  & new_n817_;
  assign new_n819_ = ~\V199(0)  & \V192(12) ;
  assign new_n820_ = ~\V199(1)  & new_n819_;
  assign new_n821_ = \V199(4)  & new_n820_;
  assign new_n822_ = \V199(0)  & \V160(12) ;
  assign new_n823_ = \V199(1)  & new_n822_;
  assign new_n824_ = \V199(4)  & new_n823_;
  assign new_n825_ = ~\V199(0)  & ~\V192(12) ;
  assign new_n826_ = \V199(1)  & new_n825_;
  assign new_n827_ = \V199(4)  & new_n826_;
  assign new_n828_ = ~new_n587_ & ~new_n827_;
  assign new_n829_ = ~new_n818_ & ~new_n821_;
  assign new_n830_ = ~new_n824_ & new_n829_;
  assign \V259(16)  = ~new_n828_ | ~new_n830_;
  assign new_n832_ = \V199(0)  & \V128(11) ;
  assign new_n833_ = ~\V199(1)  & new_n832_;
  assign new_n834_ = \V199(4)  & new_n833_;
  assign new_n835_ = ~\V199(0)  & \V192(11) ;
  assign new_n836_ = ~\V199(1)  & new_n835_;
  assign new_n837_ = \V199(4)  & new_n836_;
  assign new_n838_ = \V199(0)  & \V160(11) ;
  assign new_n839_ = \V199(1)  & new_n838_;
  assign new_n840_ = \V199(4)  & new_n839_;
  assign new_n841_ = ~\V199(0)  & ~\V192(11) ;
  assign new_n842_ = \V199(1)  & new_n841_;
  assign new_n843_ = \V199(4)  & new_n842_;
  assign new_n844_ = ~new_n587_ & ~new_n843_;
  assign new_n845_ = ~new_n834_ & ~new_n837_;
  assign new_n846_ = ~new_n840_ & new_n845_;
  assign \V259(15)  = ~new_n844_ | ~new_n846_;
  assign new_n848_ = \V199(0)  & \V128(10) ;
  assign new_n849_ = ~\V199(1)  & new_n848_;
  assign new_n850_ = \V199(4)  & new_n849_;
  assign new_n851_ = ~\V199(0)  & \V192(10) ;
  assign new_n852_ = ~\V199(1)  & new_n851_;
  assign new_n853_ = \V199(4)  & new_n852_;
  assign new_n854_ = \V199(0)  & \V160(10) ;
  assign new_n855_ = \V199(1)  & new_n854_;
  assign new_n856_ = \V199(4)  & new_n855_;
  assign new_n857_ = ~\V199(0)  & ~\V192(10) ;
  assign new_n858_ = \V199(1)  & new_n857_;
  assign new_n859_ = \V199(4)  & new_n858_;
  assign new_n860_ = ~new_n587_ & ~new_n859_;
  assign new_n861_ = ~new_n850_ & ~new_n853_;
  assign new_n862_ = ~new_n856_ & new_n861_;
  assign \V259(14)  = ~new_n860_ | ~new_n862_;
  assign new_n864_ = \V199(0)  & \V128(9) ;
  assign new_n865_ = ~\V199(1)  & new_n864_;
  assign new_n866_ = \V199(4)  & new_n865_;
  assign new_n867_ = ~\V199(0)  & \V192(9) ;
  assign new_n868_ = ~\V199(1)  & new_n867_;
  assign new_n869_ = \V199(4)  & new_n868_;
  assign new_n870_ = \V199(0)  & \V160(9) ;
  assign new_n871_ = \V199(1)  & new_n870_;
  assign new_n872_ = \V199(4)  & new_n871_;
  assign new_n873_ = ~\V199(0)  & ~\V192(9) ;
  assign new_n874_ = \V199(1)  & new_n873_;
  assign new_n875_ = \V199(4)  & new_n874_;
  assign new_n876_ = ~new_n587_ & ~new_n875_;
  assign new_n877_ = ~new_n866_ & ~new_n869_;
  assign new_n878_ = ~new_n872_ & new_n877_;
  assign \V259(13)  = ~new_n876_ | ~new_n878_;
  assign new_n880_ = \V199(0)  & \V128(8) ;
  assign new_n881_ = ~\V199(1)  & new_n880_;
  assign new_n882_ = \V199(4)  & new_n881_;
  assign new_n883_ = ~\V199(0)  & \V192(8) ;
  assign new_n884_ = ~\V199(1)  & new_n883_;
  assign new_n885_ = \V199(4)  & new_n884_;
  assign new_n886_ = \V199(0)  & \V160(8) ;
  assign new_n887_ = \V199(1)  & new_n886_;
  assign new_n888_ = \V199(4)  & new_n887_;
  assign new_n889_ = ~\V199(0)  & ~\V192(8) ;
  assign new_n890_ = \V199(1)  & new_n889_;
  assign new_n891_ = \V199(4)  & new_n890_;
  assign new_n892_ = ~new_n587_ & ~new_n891_;
  assign new_n893_ = ~new_n882_ & ~new_n885_;
  assign new_n894_ = ~new_n888_ & new_n893_;
  assign \V259(12)  = ~new_n892_ | ~new_n894_;
  assign new_n896_ = \V199(0)  & \V128(7) ;
  assign new_n897_ = ~\V199(1)  & new_n896_;
  assign new_n898_ = \V199(4)  & new_n897_;
  assign new_n899_ = ~\V199(0)  & \V192(7) ;
  assign new_n900_ = ~\V199(1)  & new_n899_;
  assign new_n901_ = \V199(4)  & new_n900_;
  assign new_n902_ = \V199(0)  & \V160(7) ;
  assign new_n903_ = \V199(1)  & new_n902_;
  assign new_n904_ = \V199(4)  & new_n903_;
  assign new_n905_ = ~\V199(0)  & ~\V192(7) ;
  assign new_n906_ = \V199(1)  & new_n905_;
  assign new_n907_ = \V199(4)  & new_n906_;
  assign new_n908_ = ~new_n587_ & ~new_n907_;
  assign new_n909_ = ~new_n898_ & ~new_n901_;
  assign new_n910_ = ~new_n904_ & new_n909_;
  assign \V259(11)  = ~new_n908_ | ~new_n910_;
  assign new_n912_ = \V199(0)  & \V128(6) ;
  assign new_n913_ = ~\V199(1)  & new_n912_;
  assign new_n914_ = \V199(4)  & new_n913_;
  assign new_n915_ = ~\V199(0)  & \V192(6) ;
  assign new_n916_ = ~\V199(1)  & new_n915_;
  assign new_n917_ = \V199(4)  & new_n916_;
  assign new_n918_ = \V199(0)  & \V160(6) ;
  assign new_n919_ = \V199(1)  & new_n918_;
  assign new_n920_ = \V199(4)  & new_n919_;
  assign new_n921_ = ~\V199(0)  & ~\V192(6) ;
  assign new_n922_ = \V199(1)  & new_n921_;
  assign new_n923_ = \V199(4)  & new_n922_;
  assign new_n924_ = ~new_n587_ & ~new_n923_;
  assign new_n925_ = ~new_n914_ & ~new_n917_;
  assign new_n926_ = ~new_n920_ & new_n925_;
  assign \V259(10)  = ~new_n924_ | ~new_n926_;
  assign new_n928_ = \V199(0)  & \V128(5) ;
  assign new_n929_ = ~\V199(1)  & new_n928_;
  assign new_n930_ = \V199(4)  & new_n929_;
  assign new_n931_ = ~\V199(0)  & \V192(5) ;
  assign new_n932_ = ~\V199(1)  & new_n931_;
  assign new_n933_ = \V199(4)  & new_n932_;
  assign new_n934_ = \V199(0)  & \V160(5) ;
  assign new_n935_ = \V199(1)  & new_n934_;
  assign new_n936_ = \V199(4)  & new_n935_;
  assign new_n937_ = ~\V199(0)  & ~\V192(5) ;
  assign new_n938_ = \V199(1)  & new_n937_;
  assign new_n939_ = \V199(4)  & new_n938_;
  assign new_n940_ = ~new_n587_ & ~new_n939_;
  assign new_n941_ = ~new_n930_ & ~new_n933_;
  assign new_n942_ = ~new_n936_ & new_n941_;
  assign \V259(9)  = ~new_n940_ | ~new_n942_;
  assign new_n944_ = \V199(0)  & \V128(4) ;
  assign new_n945_ = ~\V199(1)  & new_n944_;
  assign new_n946_ = \V199(4)  & new_n945_;
  assign new_n947_ = ~\V199(0)  & \V192(4) ;
  assign new_n948_ = ~\V199(1)  & new_n947_;
  assign new_n949_ = \V199(4)  & new_n948_;
  assign new_n950_ = \V199(0)  & \V160(4) ;
  assign new_n951_ = \V199(1)  & new_n950_;
  assign new_n952_ = \V199(4)  & new_n951_;
  assign new_n953_ = ~\V199(0)  & ~\V192(4) ;
  assign new_n954_ = \V199(1)  & new_n953_;
  assign new_n955_ = \V199(4)  & new_n954_;
  assign new_n956_ = ~new_n587_ & ~new_n955_;
  assign new_n957_ = ~new_n946_ & ~new_n949_;
  assign new_n958_ = ~new_n952_ & new_n957_;
  assign \V259(8)  = ~new_n956_ | ~new_n958_;
  assign new_n960_ = \V199(0)  & \V128(3) ;
  assign new_n961_ = ~\V199(1)  & new_n960_;
  assign new_n962_ = \V199(4)  & new_n961_;
  assign new_n963_ = ~\V199(0)  & \V192(3) ;
  assign new_n964_ = ~\V199(1)  & new_n963_;
  assign new_n965_ = \V199(4)  & new_n964_;
  assign new_n966_ = \V199(0)  & \V160(3) ;
  assign new_n967_ = \V199(1)  & new_n966_;
  assign new_n968_ = \V199(4)  & new_n967_;
  assign new_n969_ = ~\V199(0)  & ~\V192(3) ;
  assign new_n970_ = \V199(1)  & new_n969_;
  assign new_n971_ = \V199(4)  & new_n970_;
  assign new_n972_ = ~new_n587_ & ~new_n971_;
  assign new_n973_ = ~new_n962_ & ~new_n965_;
  assign new_n974_ = ~new_n968_ & new_n973_;
  assign \V259(7)  = ~new_n972_ | ~new_n974_;
  assign new_n976_ = \V199(0)  & \V128(2) ;
  assign new_n977_ = ~\V199(1)  & new_n976_;
  assign new_n978_ = \V199(4)  & new_n977_;
  assign new_n979_ = ~\V199(0)  & \V192(2) ;
  assign new_n980_ = ~\V199(1)  & new_n979_;
  assign new_n981_ = \V199(4)  & new_n980_;
  assign new_n982_ = \V199(0)  & \V160(2) ;
  assign new_n983_ = \V199(1)  & new_n982_;
  assign new_n984_ = \V199(4)  & new_n983_;
  assign new_n985_ = ~\V199(0)  & ~\V192(2) ;
  assign new_n986_ = \V199(1)  & new_n985_;
  assign new_n987_ = \V199(4)  & new_n986_;
  assign new_n988_ = ~new_n587_ & ~new_n987_;
  assign new_n989_ = ~new_n978_ & ~new_n981_;
  assign new_n990_ = ~new_n984_ & new_n989_;
  assign \V259(6)  = ~new_n988_ | ~new_n990_;
  assign new_n992_ = \V199(0)  & \V128(1) ;
  assign new_n993_ = ~\V199(1)  & new_n992_;
  assign new_n994_ = \V199(4)  & new_n993_;
  assign new_n995_ = ~\V199(0)  & \V192(1) ;
  assign new_n996_ = ~\V199(1)  & new_n995_;
  assign new_n997_ = \V199(4)  & new_n996_;
  assign new_n998_ = \V199(0)  & \V160(1) ;
  assign new_n999_ = \V199(1)  & new_n998_;
  assign new_n1000_ = \V199(4)  & new_n999_;
  assign new_n1001_ = ~\V199(0)  & ~\V192(1) ;
  assign new_n1002_ = \V199(1)  & new_n1001_;
  assign new_n1003_ = \V199(4)  & new_n1002_;
  assign new_n1004_ = ~new_n587_ & ~new_n1003_;
  assign new_n1005_ = ~new_n994_ & ~new_n997_;
  assign new_n1006_ = ~new_n1000_ & new_n1005_;
  assign \V259(5)  = ~new_n1004_ | ~new_n1006_;
  assign new_n1008_ = \V199(0)  & \V128(0) ;
  assign new_n1009_ = ~\V199(1)  & new_n1008_;
  assign new_n1010_ = \V199(4)  & new_n1009_;
  assign new_n1011_ = ~\V199(0)  & \V192(0) ;
  assign new_n1012_ = ~\V199(1)  & new_n1011_;
  assign new_n1013_ = \V199(4)  & new_n1012_;
  assign new_n1014_ = \V199(0)  & \V160(0) ;
  assign new_n1015_ = \V199(1)  & new_n1014_;
  assign new_n1016_ = \V199(4)  & new_n1015_;
  assign new_n1017_ = ~\V199(0)  & ~\V192(0) ;
  assign new_n1018_ = \V199(1)  & new_n1017_;
  assign new_n1019_ = \V199(4)  & new_n1018_;
  assign new_n1020_ = ~new_n587_ & ~new_n1019_;
  assign new_n1021_ = ~new_n1010_ & ~new_n1013_;
  assign new_n1022_ = ~new_n1016_ & new_n1021_;
  assign \V259(4)  = ~new_n1020_ | ~new_n1022_;
  assign new_n1024_ = \V199(0)  & \V32(31) ;
  assign new_n1025_ = ~\V199(1)  & new_n1024_;
  assign new_n1026_ = \V199(4)  & new_n1025_;
  assign new_n1027_ = ~\V199(0)  & \V96(31) ;
  assign new_n1028_ = ~\V199(1)  & new_n1027_;
  assign new_n1029_ = \V199(4)  & new_n1028_;
  assign new_n1030_ = \V199(0)  & \V64(31) ;
  assign new_n1031_ = \V199(1)  & new_n1030_;
  assign new_n1032_ = \V199(4)  & new_n1031_;
  assign new_n1033_ = ~\V199(0)  & ~\V96(31) ;
  assign new_n1034_ = \V199(1)  & new_n1033_;
  assign new_n1035_ = \V199(4)  & new_n1034_;
  assign new_n1036_ = ~new_n587_ & ~new_n1035_;
  assign new_n1037_ = ~new_n1026_ & ~new_n1029_;
  assign new_n1038_ = ~new_n1032_ & new_n1037_;
  assign \V259(3)  = ~new_n1036_ | ~new_n1038_;
  assign new_n1040_ = \V199(0)  & \V32(30) ;
  assign new_n1041_ = ~\V199(1)  & new_n1040_;
  assign new_n1042_ = \V199(4)  & new_n1041_;
  assign new_n1043_ = ~\V199(0)  & \V96(30) ;
  assign new_n1044_ = ~\V199(1)  & new_n1043_;
  assign new_n1045_ = \V199(4)  & new_n1044_;
  assign new_n1046_ = \V199(0)  & \V64(30) ;
  assign new_n1047_ = \V199(1)  & new_n1046_;
  assign new_n1048_ = \V199(4)  & new_n1047_;
  assign new_n1049_ = ~\V199(0)  & ~\V96(30) ;
  assign new_n1050_ = \V199(1)  & new_n1049_;
  assign new_n1051_ = \V199(4)  & new_n1050_;
  assign new_n1052_ = ~new_n587_ & ~new_n1051_;
  assign new_n1053_ = ~new_n1042_ & ~new_n1045_;
  assign new_n1054_ = ~new_n1048_ & new_n1053_;
  assign \V259(2)  = ~new_n1052_ | ~new_n1054_;
  assign new_n1056_ = \V199(0)  & \V32(29) ;
  assign new_n1057_ = ~\V199(1)  & new_n1056_;
  assign new_n1058_ = \V199(4)  & new_n1057_;
  assign new_n1059_ = ~\V199(0)  & \V96(29) ;
  assign new_n1060_ = ~\V199(1)  & new_n1059_;
  assign new_n1061_ = \V199(4)  & new_n1060_;
  assign new_n1062_ = \V199(0)  & \V64(29) ;
  assign new_n1063_ = \V199(1)  & new_n1062_;
  assign new_n1064_ = \V199(4)  & new_n1063_;
  assign new_n1065_ = ~\V199(0)  & ~\V96(29) ;
  assign new_n1066_ = \V199(1)  & new_n1065_;
  assign new_n1067_ = \V199(4)  & new_n1066_;
  assign new_n1068_ = ~new_n587_ & ~new_n1067_;
  assign new_n1069_ = ~new_n1058_ & ~new_n1061_;
  assign new_n1070_ = ~new_n1064_ & new_n1069_;
  assign \V259(1)  = ~new_n1068_ | ~new_n1070_;
  assign new_n1072_ = \V199(0)  & \V32(28) ;
  assign new_n1073_ = ~\V199(1)  & new_n1072_;
  assign new_n1074_ = \V199(4)  & new_n1073_;
  assign new_n1075_ = ~\V199(0)  & \V96(28) ;
  assign new_n1076_ = ~\V199(1)  & new_n1075_;
  assign new_n1077_ = \V199(4)  & new_n1076_;
  assign new_n1078_ = \V199(0)  & \V64(28) ;
  assign new_n1079_ = \V199(1)  & new_n1078_;
  assign new_n1080_ = \V199(4)  & new_n1079_;
  assign new_n1081_ = ~\V199(0)  & ~\V96(28) ;
  assign new_n1082_ = \V199(1)  & new_n1081_;
  assign new_n1083_ = \V199(4)  & new_n1082_;
  assign new_n1084_ = ~new_n587_ & ~new_n1083_;
  assign new_n1085_ = ~new_n1074_ & ~new_n1077_;
  assign new_n1086_ = ~new_n1080_ & new_n1085_;
  assign \V259(0)  = ~new_n1084_ | ~new_n1086_;
  assign new_n1088_ = ~\V199(0)  & \V195(0) ;
  assign new_n1089_ = \V199(1)  & new_n1088_;
  assign new_n1090_ = \V199(3)  & new_n1089_;
  assign new_n1091_ = ~\V199(1)  & new_n1088_;
  assign new_n1092_ = \V199(3)  & new_n1091_;
  assign \V266(6)  = new_n1090_ | new_n1092_;
  assign new_n1094_ = \V199(1)  & ~\V199(3) ;
  assign new_n1095_ = ~\V199(0)  & \V194(1) ;
  assign new_n1096_ = ~\V199(1)  & new_n1095_;
  assign new_n1097_ = \V199(3)  & new_n1096_;
  assign new_n1098_ = \V199(1)  & \V199(3) ;
  assign new_n1099_ = \V199(0)  & new_n1098_;
  assign new_n1100_ = ~\V199(0)  & ~\V194(1) ;
  assign new_n1101_ = \V199(1)  & new_n1100_;
  assign new_n1102_ = \V199(3)  & new_n1101_;
  assign new_n1103_ = ~new_n1099_ & ~new_n1102_;
  assign new_n1104_ = ~new_n1094_ & ~new_n1097_;
  assign \V266(5)  = ~new_n1103_ | ~new_n1104_;
  assign new_n1106_ = ~\V199(0)  & \V194(0) ;
  assign new_n1107_ = ~\V199(1)  & new_n1106_;
  assign new_n1108_ = \V199(3)  & new_n1107_;
  assign new_n1109_ = ~\V199(0)  & ~\V194(0) ;
  assign new_n1110_ = \V199(1)  & new_n1109_;
  assign new_n1111_ = \V199(3)  & new_n1110_;
  assign new_n1112_ = ~new_n1099_ & ~new_n1111_;
  assign new_n1113_ = ~new_n1094_ & ~new_n1108_;
  assign \V266(4)  = ~new_n1112_ | ~new_n1113_;
  assign new_n1115_ = \V199(0)  & \V128(31) ;
  assign new_n1116_ = ~\V199(1)  & new_n1115_;
  assign new_n1117_ = \V199(3)  & new_n1116_;
  assign new_n1118_ = ~\V199(0)  & \V192(31) ;
  assign new_n1119_ = ~\V199(1)  & new_n1118_;
  assign new_n1120_ = \V199(3)  & new_n1119_;
  assign new_n1121_ = \V160(31)  & new_n1099_;
  assign new_n1122_ = ~\V199(0)  & ~\V192(31) ;
  assign new_n1123_ = \V199(1)  & new_n1122_;
  assign new_n1124_ = \V199(3)  & new_n1123_;
  assign new_n1125_ = ~new_n1094_ & ~new_n1124_;
  assign new_n1126_ = ~new_n1117_ & ~new_n1120_;
  assign new_n1127_ = ~new_n1121_ & new_n1126_;
  assign \V266(3)  = ~new_n1125_ | ~new_n1127_;
  assign new_n1129_ = \V199(0)  & \V128(30) ;
  assign new_n1130_ = ~\V199(1)  & new_n1129_;
  assign new_n1131_ = \V199(3)  & new_n1130_;
  assign new_n1132_ = ~\V199(0)  & \V192(30) ;
  assign new_n1133_ = ~\V199(1)  & new_n1132_;
  assign new_n1134_ = \V199(3)  & new_n1133_;
  assign new_n1135_ = \V160(30)  & new_n1099_;
  assign new_n1136_ = ~\V199(0)  & ~\V192(30) ;
  assign new_n1137_ = \V199(1)  & new_n1136_;
  assign new_n1138_ = \V199(3)  & new_n1137_;
  assign new_n1139_ = ~new_n1094_ & ~new_n1138_;
  assign new_n1140_ = ~new_n1131_ & ~new_n1134_;
  assign new_n1141_ = ~new_n1135_ & new_n1140_;
  assign \V266(2)  = ~new_n1139_ | ~new_n1141_;
  assign new_n1143_ = \V199(0)  & \V128(29) ;
  assign new_n1144_ = ~\V199(1)  & new_n1143_;
  assign new_n1145_ = \V199(3)  & new_n1144_;
  assign new_n1146_ = ~\V199(0)  & \V192(29) ;
  assign new_n1147_ = ~\V199(1)  & new_n1146_;
  assign new_n1148_ = \V199(3)  & new_n1147_;
  assign new_n1149_ = \V160(29)  & new_n1099_;
  assign new_n1150_ = ~\V199(0)  & ~\V192(29) ;
  assign new_n1151_ = \V199(1)  & new_n1150_;
  assign new_n1152_ = \V199(3)  & new_n1151_;
  assign new_n1153_ = ~new_n1094_ & ~new_n1152_;
  assign new_n1154_ = ~new_n1145_ & ~new_n1148_;
  assign new_n1155_ = ~new_n1149_ & new_n1154_;
  assign \V266(1)  = ~new_n1153_ | ~new_n1155_;
  assign new_n1157_ = \V199(0)  & \V128(28) ;
  assign new_n1158_ = ~\V199(1)  & new_n1157_;
  assign new_n1159_ = \V199(3)  & new_n1158_;
  assign new_n1160_ = ~\V199(0)  & \V192(28) ;
  assign new_n1161_ = ~\V199(1)  & new_n1160_;
  assign new_n1162_ = \V199(3)  & new_n1161_;
  assign new_n1163_ = \V160(28)  & new_n1099_;
  assign new_n1164_ = ~\V199(0)  & ~\V192(28) ;
  assign new_n1165_ = \V199(1)  & new_n1164_;
  assign new_n1166_ = \V199(3)  & new_n1165_;
  assign new_n1167_ = ~new_n1094_ & ~new_n1166_;
  assign new_n1168_ = ~new_n1159_ & ~new_n1162_;
  assign new_n1169_ = ~new_n1163_ & new_n1168_;
  assign \V266(0)  = ~new_n1167_ | ~new_n1169_;
endmodule

